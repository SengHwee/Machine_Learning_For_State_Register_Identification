
module sha1_core(clk, reset_n, init, next, \block[0] , \block[1] , \block[2] , \block[3] , \block[4] , \block[5] , \block[6] , \block[7] , \block[8] , \block[9] , \block[10] , \block[11] , \block[12] , \block[13] , \block[14] , \block[15] , \block[16] , \block[17] , \block[18] , \block[19] , \block[20] , \block[21] , \block[22] , \block[23] , \block[24] , \block[25] , \block[26] , \block[27] , \block[28] , \block[29] , \block[30] , \block[31] , \block[32] , \block[33] , \block[34] , \block[35] , \block[36] , \block[37] , \block[38] , \block[39] , \block[40] , \block[41] , \block[42] , \block[43] , \block[44] , \block[45] , \block[46] , \block[47] , \block[48] , \block[49] , \block[50] , \block[51] , \block[52] , \block[53] , \block[54] , \block[55] , \block[56] , \block[57] , \block[58] , \block[59] , \block[60] , \block[61] , \block[62] , \block[63] , \block[64] , \block[65] , \block[66] , \block[67] , \block[68] , \block[69] , \block[70] , \block[71] , \block[72] , \block[73] , \block[74] , \block[75] , \block[76] , \block[77] , \block[78] , \block[79] , \block[80] , \block[81] , \block[82] , \block[83] , \block[84] , \block[85] , \block[86] , \block[87] , \block[88] , \block[89] , \block[90] , \block[91] , \block[92] , \block[93] , \block[94] , \block[95] , \block[96] , \block[97] , \block[98] , \block[99] , \block[100] , \block[101] , \block[102] , \block[103] , \block[104] , \block[105] , \block[106] , \block[107] , \block[108] , \block[109] , \block[110] , \block[111] , \block[112] , \block[113] , \block[114] , \block[115] , \block[116] , \block[117] , \block[118] , \block[119] , \block[120] , \block[121] , \block[122] , \block[123] , \block[124] , \block[125] , \block[126] , \block[127] , \block[128] , \block[129] , \block[130] , \block[131] , \block[132] , \block[133] , \block[134] , \block[135] , \block[136] , \block[137] , \block[138] , \block[139] , \block[140] , \block[141] , \block[142] , \block[143] , \block[144] , \block[145] , \block[146] , \block[147] , \block[148] , \block[149] , \block[150] , \block[151] , \block[152] , \block[153] , \block[154] , \block[155] , \block[156] , \block[157] , \block[158] , \block[159] , \block[160] , \block[161] , \block[162] , \block[163] , \block[164] , \block[165] , \block[166] , \block[167] , \block[168] , \block[169] , \block[170] , \block[171] , \block[172] , \block[173] , \block[174] , \block[175] , \block[176] , \block[177] , \block[178] , \block[179] , \block[180] , \block[181] , \block[182] , \block[183] , \block[184] , \block[185] , \block[186] , \block[187] , \block[188] , \block[189] , \block[190] , \block[191] , \block[192] , \block[193] , \block[194] , \block[195] , \block[196] , \block[197] , \block[198] , \block[199] , \block[200] , \block[201] , \block[202] , \block[203] , \block[204] , \block[205] , \block[206] , \block[207] , \block[208] , \block[209] , \block[210] , \block[211] , \block[212] , \block[213] , \block[214] , \block[215] , \block[216] , \block[217] , \block[218] , \block[219] , \block[220] , \block[221] , \block[222] , \block[223] , \block[224] , \block[225] , \block[226] , \block[227] , \block[228] , \block[229] , \block[230] , \block[231] , \block[232] , \block[233] , \block[234] , \block[235] , \block[236] , \block[237] , \block[238] , \block[239] , \block[240] , \block[241] , \block[242] , \block[243] , \block[244] , \block[245] , \block[246] , \block[247] , \block[248] , \block[249] , \block[250] , \block[251] , \block[252] , \block[253] , \block[254] , \block[255] , \block[256] , \block[257] , \block[258] , \block[259] , \block[260] , \block[261] , \block[262] , \block[263] , \block[264] , \block[265] , \block[266] , \block[267] , \block[268] , \block[269] , \block[270] , \block[271] , \block[272] , \block[273] , \block[274] , \block[275] , \block[276] , \block[277] , \block[278] , \block[279] , \block[280] , \block[281] , \block[282] , \block[283] , \block[284] , \block[285] , \block[286] , \block[287] , \block[288] , \block[289] , \block[290] , \block[291] , \block[292] , \block[293] , \block[294] , \block[295] , \block[296] , \block[297] , \block[298] , \block[299] , \block[300] , \block[301] , \block[302] , \block[303] , \block[304] , \block[305] , \block[306] , \block[307] , \block[308] , \block[309] , \block[310] , \block[311] , \block[312] , \block[313] , \block[314] , \block[315] , \block[316] , \block[317] , \block[318] , \block[319] , \block[320] , \block[321] , \block[322] , \block[323] , \block[324] , \block[325] , \block[326] , \block[327] , \block[328] , \block[329] , \block[330] , \block[331] , \block[332] , \block[333] , \block[334] , \block[335] , \block[336] , \block[337] , \block[338] , \block[339] , \block[340] , \block[341] , \block[342] , \block[343] , \block[344] , \block[345] , \block[346] , \block[347] , \block[348] , \block[349] , \block[350] , \block[351] , \block[352] , \block[353] , \block[354] , \block[355] , \block[356] , \block[357] , \block[358] , \block[359] , \block[360] , \block[361] , \block[362] , \block[363] , \block[364] , \block[365] , \block[366] , \block[367] , \block[368] , \block[369] , \block[370] , \block[371] , \block[372] , \block[373] , \block[374] , \block[375] , \block[376] , \block[377] , \block[378] , \block[379] , \block[380] , \block[381] , \block[382] , \block[383] , \block[384] , \block[385] , \block[386] , \block[387] , \block[388] , \block[389] , \block[390] , \block[391] , \block[392] , \block[393] , \block[394] , \block[395] , \block[396] , \block[397] , \block[398] , \block[399] , \block[400] , \block[401] , \block[402] , \block[403] , \block[404] , \block[405] , \block[406] , \block[407] , \block[408] , \block[409] , \block[410] , \block[411] , \block[412] , \block[413] , \block[414] , \block[415] , \block[416] , \block[417] , \block[418] , \block[419] , \block[420] , \block[421] , \block[422] , \block[423] , \block[424] , \block[425] , \block[426] , \block[427] , \block[428] , \block[429] , \block[430] , \block[431] , \block[432] , \block[433] , \block[434] , \block[435] , \block[436] , \block[437] , \block[438] , \block[439] , \block[440] , \block[441] , \block[442] , \block[443] , \block[444] , \block[445] , \block[446] , \block[447] , \block[448] , \block[449] , \block[450] , \block[451] , \block[452] , \block[453] , \block[454] , \block[455] , \block[456] , \block[457] , \block[458] , \block[459] , \block[460] , \block[461] , \block[462] , \block[463] , \block[464] , \block[465] , \block[466] , \block[467] , \block[468] , \block[469] , \block[470] , \block[471] , \block[472] , \block[473] , \block[474] , \block[475] , \block[476] , \block[477] , \block[478] , \block[479] , \block[480] , \block[481] , \block[482] , \block[483] , \block[484] , \block[485] , \block[486] , \block[487] , \block[488] , \block[489] , \block[490] , \block[491] , \block[492] , \block[493] , \block[494] , \block[495] , \block[496] , \block[497] , \block[498] , \block[499] , \block[500] , \block[501] , \block[502] , \block[503] , \block[504] , \block[505] , \block[506] , \block[507] , \block[508] , \block[509] , \block[510] , \block[511] , ready, \digest[0] , \digest[1] , \digest[2] , \digest[3] , \digest[4] , \digest[5] , \digest[6] , \digest[7] , \digest[8] , \digest[9] , \digest[10] , \digest[11] , \digest[12] , \digest[13] , \digest[14] , \digest[15] , \digest[16] , \digest[17] , \digest[18] , \digest[19] , \digest[20] , \digest[21] , \digest[22] , \digest[23] , \digest[24] , \digest[25] , \digest[26] , \digest[27] , \digest[28] , \digest[29] , \digest[30] , \digest[31] , \digest[32] , \digest[33] , \digest[34] , \digest[35] , \digest[36] , \digest[37] , \digest[38] , \digest[39] , \digest[40] , \digest[41] , \digest[42] , \digest[43] , \digest[44] , \digest[45] , \digest[46] , \digest[47] , \digest[48] , \digest[49] , \digest[50] , \digest[51] , \digest[52] , \digest[53] , \digest[54] , \digest[55] , \digest[56] , \digest[57] , \digest[58] , \digest[59] , \digest[60] , \digest[61] , \digest[62] , \digest[63] , \digest[64] , \digest[65] , \digest[66] , \digest[67] , \digest[68] , \digest[69] , \digest[70] , \digest[71] , \digest[72] , \digest[73] , \digest[74] , \digest[75] , \digest[76] , \digest[77] , \digest[78] , \digest[79] , \digest[80] , \digest[81] , \digest[82] , \digest[83] , \digest[84] , \digest[85] , \digest[86] , \digest[87] , \digest[88] , \digest[89] , \digest[90] , \digest[91] , \digest[92] , \digest[93] , \digest[94] , \digest[95] , \digest[96] , \digest[97] , \digest[98] , \digest[99] , \digest[100] , \digest[101] , \digest[102] , \digest[103] , \digest[104] , \digest[105] , \digest[106] , \digest[107] , \digest[108] , \digest[109] , \digest[110] , \digest[111] , \digest[112] , \digest[113] , \digest[114] , \digest[115] , \digest[116] , \digest[117] , \digest[118] , \digest[119] , \digest[120] , \digest[121] , \digest[122] , \digest[123] , \digest[124] , \digest[125] , \digest[126] , \digest[127] , \digest[128] , \digest[129] , \digest[130] , \digest[131] , \digest[132] , \digest[133] , \digest[134] , \digest[135] , \digest[136] , \digest[137] , \digest[138] , \digest[139] , \digest[140] , \digest[141] , \digest[142] , \digest[143] , \digest[144] , \digest[145] , \digest[146] , \digest[147] , \digest[148] , \digest[149] , \digest[150] , \digest[151] , \digest[152] , \digest[153] , \digest[154] , \digest[155] , \digest[156] , \digest[157] , \digest[158] , \digest[159] , digest_valid);
  wire H0_reg_0__FF_INPUT;
  wire H0_reg_10__FF_INPUT;
  wire H0_reg_11__FF_INPUT;
  wire H0_reg_12__FF_INPUT;
  wire H0_reg_13__FF_INPUT;
  wire H0_reg_14__FF_INPUT;
  wire H0_reg_15__FF_INPUT;
  wire H0_reg_16__FF_INPUT;
  wire H0_reg_17__FF_INPUT;
  wire H0_reg_18__FF_INPUT;
  wire H0_reg_19__FF_INPUT;
  wire H0_reg_1__FF_INPUT;
  wire H0_reg_20__FF_INPUT;
  wire H0_reg_21__FF_INPUT;
  wire H0_reg_22__FF_INPUT;
  wire H0_reg_23__FF_INPUT;
  wire H0_reg_24__FF_INPUT;
  wire H0_reg_25__FF_INPUT;
  wire H0_reg_26__FF_INPUT;
  wire H0_reg_27__FF_INPUT;
  wire H0_reg_28__FF_INPUT;
  wire H0_reg_29__FF_INPUT;
  wire H0_reg_2__FF_INPUT;
  wire H0_reg_30__FF_INPUT;
  wire H0_reg_31__FF_INPUT;
  wire H0_reg_3__FF_INPUT;
  wire H0_reg_4__FF_INPUT;
  wire H0_reg_5__FF_INPUT;
  wire H0_reg_6__FF_INPUT;
  wire H0_reg_7__FF_INPUT;
  wire H0_reg_8__FF_INPUT;
  wire H0_reg_9__FF_INPUT;
  wire H1_reg_0__FF_INPUT;
  wire H1_reg_10__FF_INPUT;
  wire H1_reg_11__FF_INPUT;
  wire H1_reg_12__FF_INPUT;
  wire H1_reg_13__FF_INPUT;
  wire H1_reg_14__FF_INPUT;
  wire H1_reg_15__FF_INPUT;
  wire H1_reg_16__FF_INPUT;
  wire H1_reg_17__FF_INPUT;
  wire H1_reg_18__FF_INPUT;
  wire H1_reg_19__FF_INPUT;
  wire H1_reg_1__FF_INPUT;
  wire H1_reg_20__FF_INPUT;
  wire H1_reg_21__FF_INPUT;
  wire H1_reg_22__FF_INPUT;
  wire H1_reg_23__FF_INPUT;
  wire H1_reg_24__FF_INPUT;
  wire H1_reg_25__FF_INPUT;
  wire H1_reg_26__FF_INPUT;
  wire H1_reg_27__FF_INPUT;
  wire H1_reg_28__FF_INPUT;
  wire H1_reg_29__FF_INPUT;
  wire H1_reg_2__FF_INPUT;
  wire H1_reg_30__FF_INPUT;
  wire H1_reg_31__FF_INPUT;
  wire H1_reg_3__FF_INPUT;
  wire H1_reg_4__FF_INPUT;
  wire H1_reg_5__FF_INPUT;
  wire H1_reg_6__FF_INPUT;
  wire H1_reg_7__FF_INPUT;
  wire H1_reg_8__FF_INPUT;
  wire H1_reg_9__FF_INPUT;
  wire H2_reg_0__FF_INPUT;
  wire H2_reg_10__FF_INPUT;
  wire H2_reg_11__FF_INPUT;
  wire H2_reg_12__FF_INPUT;
  wire H2_reg_13__FF_INPUT;
  wire H2_reg_14__FF_INPUT;
  wire H2_reg_15__FF_INPUT;
  wire H2_reg_16__FF_INPUT;
  wire H2_reg_17__FF_INPUT;
  wire H2_reg_18__FF_INPUT;
  wire H2_reg_19__FF_INPUT;
  wire H2_reg_1__FF_INPUT;
  wire H2_reg_20__FF_INPUT;
  wire H2_reg_21__FF_INPUT;
  wire H2_reg_22__FF_INPUT;
  wire H2_reg_23__FF_INPUT;
  wire H2_reg_24__FF_INPUT;
  wire H2_reg_25__FF_INPUT;
  wire H2_reg_26__FF_INPUT;
  wire H2_reg_27__FF_INPUT;
  wire H2_reg_28__FF_INPUT;
  wire H2_reg_29__FF_INPUT;
  wire H2_reg_2__FF_INPUT;
  wire H2_reg_30__FF_INPUT;
  wire H2_reg_31__FF_INPUT;
  wire H2_reg_3__FF_INPUT;
  wire H2_reg_4__FF_INPUT;
  wire H2_reg_5__FF_INPUT;
  wire H2_reg_6__FF_INPUT;
  wire H2_reg_7__FF_INPUT;
  wire H2_reg_8__FF_INPUT;
  wire H2_reg_9__FF_INPUT;
  wire H3_reg_0__FF_INPUT;
  wire H3_reg_10__FF_INPUT;
  wire H3_reg_11__FF_INPUT;
  wire H3_reg_12__FF_INPUT;
  wire H3_reg_13__FF_INPUT;
  wire H3_reg_14__FF_INPUT;
  wire H3_reg_15__FF_INPUT;
  wire H3_reg_16__FF_INPUT;
  wire H3_reg_17__FF_INPUT;
  wire H3_reg_18__FF_INPUT;
  wire H3_reg_19__FF_INPUT;
  wire H3_reg_1__FF_INPUT;
  wire H3_reg_20__FF_INPUT;
  wire H3_reg_21__FF_INPUT;
  wire H3_reg_22__FF_INPUT;
  wire H3_reg_23__FF_INPUT;
  wire H3_reg_24__FF_INPUT;
  wire H3_reg_25__FF_INPUT;
  wire H3_reg_26__FF_INPUT;
  wire H3_reg_27__FF_INPUT;
  wire H3_reg_28__FF_INPUT;
  wire H3_reg_29__FF_INPUT;
  wire H3_reg_2__FF_INPUT;
  wire H3_reg_30__FF_INPUT;
  wire H3_reg_31__FF_INPUT;
  wire H3_reg_3__FF_INPUT;
  wire H3_reg_4__FF_INPUT;
  wire H3_reg_5__FF_INPUT;
  wire H3_reg_6__FF_INPUT;
  wire H3_reg_7__FF_INPUT;
  wire H3_reg_8__FF_INPUT;
  wire H3_reg_9__FF_INPUT;
  wire H4_reg_0__FF_INPUT;
  wire H4_reg_10__FF_INPUT;
  wire H4_reg_11__FF_INPUT;
  wire H4_reg_12__FF_INPUT;
  wire H4_reg_13__FF_INPUT;
  wire H4_reg_14__FF_INPUT;
  wire H4_reg_15__FF_INPUT;
  wire H4_reg_16__FF_INPUT;
  wire H4_reg_17__FF_INPUT;
  wire H4_reg_18__FF_INPUT;
  wire H4_reg_19__FF_INPUT;
  wire H4_reg_1__FF_INPUT;
  wire H4_reg_20__FF_INPUT;
  wire H4_reg_21__FF_INPUT;
  wire H4_reg_22__FF_INPUT;
  wire H4_reg_23__FF_INPUT;
  wire H4_reg_24__FF_INPUT;
  wire H4_reg_25__FF_INPUT;
  wire H4_reg_26__FF_INPUT;
  wire H4_reg_27__FF_INPUT;
  wire H4_reg_28__FF_INPUT;
  wire H4_reg_29__FF_INPUT;
  wire H4_reg_2__FF_INPUT;
  wire H4_reg_30__FF_INPUT;
  wire H4_reg_31__FF_INPUT;
  wire H4_reg_3__FF_INPUT;
  wire H4_reg_4__FF_INPUT;
  wire H4_reg_5__FF_INPUT;
  wire H4_reg_6__FF_INPUT;
  wire H4_reg_7__FF_INPUT;
  wire H4_reg_8__FF_INPUT;
  wire H4_reg_9__FF_INPUT;
  wire _abc_15724_n1000;
  wire _abc_15724_n1001;
  wire _abc_15724_n1002;
  wire _abc_15724_n1003;
  wire _abc_15724_n1004;
  wire _abc_15724_n1005;
  wire _abc_15724_n1006;
  wire _abc_15724_n1008;
  wire _abc_15724_n1009;
  wire _abc_15724_n1010;
  wire _abc_15724_n1011;
  wire _abc_15724_n1012;
  wire _abc_15724_n1013;
  wire _abc_15724_n1014;
  wire _abc_15724_n1015_1;
  wire _abc_15724_n1016_1;
  wire _abc_15724_n1017;
  wire _abc_15724_n1018_1;
  wire _abc_15724_n1019;
  wire _abc_15724_n1020;
  wire _abc_15724_n1021;
  wire _abc_15724_n1023;
  wire _abc_15724_n1024_1;
  wire _abc_15724_n1025_1;
  wire _abc_15724_n1026_1;
  wire _abc_15724_n1027;
  wire _abc_15724_n1028;
  wire _abc_15724_n1029;
  wire _abc_15724_n1030;
  wire _abc_15724_n1031;
  wire _abc_15724_n1032;
  wire _abc_15724_n1033;
  wire _abc_15724_n1034;
  wire _abc_15724_n1035;
  wire _abc_15724_n1036;
  wire _abc_15724_n1038_1;
  wire _abc_15724_n1039_1;
  wire _abc_15724_n1040;
  wire _abc_15724_n1041;
  wire _abc_15724_n1042;
  wire _abc_15724_n1043;
  wire _abc_15724_n1044;
  wire _abc_15724_n1045;
  wire _abc_15724_n1046;
  wire _abc_15724_n1047_1;
  wire _abc_15724_n1048_1;
  wire _abc_15724_n1049;
  wire _abc_15724_n1050_1;
  wire _abc_15724_n1052;
  wire _abc_15724_n1053;
  wire _abc_15724_n1054;
  wire _abc_15724_n1055;
  wire _abc_15724_n1056;
  wire _abc_15724_n1057;
  wire _abc_15724_n1058;
  wire _abc_15724_n1059;
  wire _abc_15724_n1060_1;
  wire _abc_15724_n1061_1;
  wire _abc_15724_n1062;
  wire _abc_15724_n1063_1;
  wire _abc_15724_n1064;
  wire _abc_15724_n1065;
  wire _abc_15724_n1066;
  wire _abc_15724_n1067;
  wire _abc_15724_n1069_1;
  wire _abc_15724_n1070_1;
  wire _abc_15724_n1071_1;
  wire _abc_15724_n1072;
  wire _abc_15724_n1073;
  wire _abc_15724_n1074;
  wire _abc_15724_n1075;
  wire _abc_15724_n1076;
  wire _abc_15724_n1077;
  wire _abc_15724_n1078;
  wire _abc_15724_n1079;
  wire _abc_15724_n1080;
  wire _abc_15724_n1081;
  wire _abc_15724_n1082_1;
  wire _abc_15724_n1084_1;
  wire _abc_15724_n1085;
  wire _abc_15724_n1086;
  wire _abc_15724_n1087;
  wire _abc_15724_n1088;
  wire _abc_15724_n1089;
  wire _abc_15724_n1090_1;
  wire _abc_15724_n1091_1;
  wire _abc_15724_n1092_1;
  wire _abc_15724_n1093;
  wire _abc_15724_n1094;
  wire _abc_15724_n1095;
  wire _abc_15724_n1096;
  wire _abc_15724_n1097;
  wire _abc_15724_n1099;
  wire _abc_15724_n1100;
  wire _abc_15724_n1101;
  wire _abc_15724_n1102;
  wire _abc_15724_n1103;
  wire _abc_15724_n1104;
  wire _abc_15724_n1105;
  wire _abc_15724_n1106;
  wire _abc_15724_n1107;
  wire _abc_15724_n1108;
  wire _abc_15724_n1109_1;
  wire _abc_15724_n1110_1;
  wire _abc_15724_n1111_1;
  wire _abc_15724_n1113;
  wire _abc_15724_n1114;
  wire _abc_15724_n1115;
  wire _abc_15724_n1116;
  wire _abc_15724_n1117;
  wire _abc_15724_n1118;
  wire _abc_15724_n1119_1;
  wire _abc_15724_n1120_1;
  wire _abc_15724_n1121_1;
  wire _abc_15724_n1122;
  wire _abc_15724_n1123;
  wire _abc_15724_n1124;
  wire _abc_15724_n1126;
  wire _abc_15724_n1127;
  wire _abc_15724_n1128;
  wire _abc_15724_n1129;
  wire _abc_15724_n1130;
  wire _abc_15724_n1131_1;
  wire _abc_15724_n1132_1;
  wire _abc_15724_n1133_1;
  wire _abc_15724_n1134;
  wire _abc_15724_n1135;
  wire _abc_15724_n1136;
  wire _abc_15724_n1137;
  wire _abc_15724_n1139;
  wire _abc_15724_n1140;
  wire _abc_15724_n1141_1;
  wire _abc_15724_n1142_1;
  wire _abc_15724_n1143;
  wire _abc_15724_n1144_1;
  wire _abc_15724_n1145;
  wire _abc_15724_n1146;
  wire _abc_15724_n1147;
  wire _abc_15724_n1148;
  wire _abc_15724_n1149;
  wire _abc_15724_n1150;
  wire _abc_15724_n1151;
  wire _abc_15724_n1153;
  wire _abc_15724_n1154;
  wire _abc_15724_n1155_1;
  wire _abc_15724_n1156_1;
  wire _abc_15724_n1157_1;
  wire _abc_15724_n1158;
  wire _abc_15724_n1159;
  wire _abc_15724_n1160;
  wire _abc_15724_n1161;
  wire _abc_15724_n1162;
  wire _abc_15724_n1163;
  wire _abc_15724_n1164;
  wire _abc_15724_n1166_1;
  wire _abc_15724_n1167_1;
  wire _abc_15724_n1168;
  wire _abc_15724_n1169;
  wire _abc_15724_n1170;
  wire _abc_15724_n1171;
  wire _abc_15724_n1172;
  wire _abc_15724_n1173;
  wire _abc_15724_n1174;
  wire _abc_15724_n1175;
  wire _abc_15724_n1176;
  wire _abc_15724_n1177_1;
  wire _abc_15724_n1178_1;
  wire _abc_15724_n1179_1;
  wire _abc_15724_n1180;
  wire _abc_15724_n1181;
  wire _abc_15724_n1182;
  wire _abc_15724_n1183;
  wire _abc_15724_n1184;
  wire _abc_15724_n1185_1;
  wire _abc_15724_n1186_1;
  wire _abc_15724_n1187_1;
  wire _abc_15724_n1189;
  wire _abc_15724_n1190_1;
  wire _abc_15724_n1191_1;
  wire _abc_15724_n1192;
  wire _abc_15724_n1193_1;
  wire _abc_15724_n1194;
  wire _abc_15724_n1195;
  wire _abc_15724_n1196;
  wire _abc_15724_n1197_1;
  wire _abc_15724_n1198_1;
  wire _abc_15724_n1199;
  wire _abc_15724_n1200_1;
  wire _abc_15724_n1201;
  wire _abc_15724_n1202;
  wire _abc_15724_n1204;
  wire _abc_15724_n1205;
  wire _abc_15724_n1206_1;
  wire _abc_15724_n1207_1;
  wire _abc_15724_n1208;
  wire _abc_15724_n1209_1;
  wire _abc_15724_n1210;
  wire _abc_15724_n1211;
  wire _abc_15724_n1212;
  wire _abc_15724_n1213;
  wire _abc_15724_n1214;
  wire _abc_15724_n1215_1;
  wire _abc_15724_n1216_1;
  wire _abc_15724_n1218_1;
  wire _abc_15724_n1219;
  wire _abc_15724_n1220;
  wire _abc_15724_n1221;
  wire _abc_15724_n1222;
  wire _abc_15724_n1223;
  wire _abc_15724_n1224;
  wire _abc_15724_n1225;
  wire _abc_15724_n1226;
  wire _abc_15724_n1227;
  wire _abc_15724_n1228_1;
  wire _abc_15724_n1229_1;
  wire _abc_15724_n1231_1;
  wire _abc_15724_n1232;
  wire _abc_15724_n1233;
  wire _abc_15724_n1234;
  wire _abc_15724_n1235;
  wire _abc_15724_n1236;
  wire _abc_15724_n1237_1;
  wire _abc_15724_n1238_1;
  wire _abc_15724_n1239;
  wire _abc_15724_n1240_1;
  wire _abc_15724_n1241;
  wire _abc_15724_n1242;
  wire _abc_15724_n1243;
  wire _abc_15724_n1244;
  wire _abc_15724_n1245;
  wire _abc_15724_n1246;
  wire _abc_15724_n1247;
  wire _abc_15724_n1248;
  wire _abc_15724_n1249;
  wire _abc_15724_n1250_1;
  wire _abc_15724_n1251_1;
  wire _abc_15724_n1252;
  wire _abc_15724_n1254;
  wire _abc_15724_n1255;
  wire _abc_15724_n1256;
  wire _abc_15724_n1257;
  wire _abc_15724_n1258;
  wire _abc_15724_n1259_1;
  wire _abc_15724_n1260_1;
  wire _abc_15724_n1261_1;
  wire _abc_15724_n1262;
  wire _abc_15724_n1263;
  wire _abc_15724_n1264;
  wire _abc_15724_n1265;
  wire _abc_15724_n1266;
  wire _abc_15724_n1268;
  wire _abc_15724_n1269;
  wire _abc_15724_n1270;
  wire _abc_15724_n1271;
  wire _abc_15724_n1272;
  wire _abc_15724_n1273;
  wire _abc_15724_n1274_1;
  wire _abc_15724_n1275_1;
  wire _abc_15724_n1276_1;
  wire _abc_15724_n1277;
  wire _abc_15724_n1278;
  wire _abc_15724_n1279;
  wire _abc_15724_n1280;
  wire _abc_15724_n1281;
  wire _abc_15724_n1282;
  wire _abc_15724_n1284_1;
  wire _abc_15724_n1285_1;
  wire _abc_15724_n1286;
  wire _abc_15724_n1287_1;
  wire _abc_15724_n1288;
  wire _abc_15724_n1289;
  wire _abc_15724_n1290;
  wire _abc_15724_n1291;
  wire _abc_15724_n1292;
  wire _abc_15724_n1293;
  wire _abc_15724_n1294;
  wire _abc_15724_n1295;
  wire _abc_15724_n1297_1;
  wire _abc_15724_n1298;
  wire _abc_15724_n1299_1;
  wire _abc_15724_n1300;
  wire _abc_15724_n1301;
  wire _abc_15724_n1302;
  wire _abc_15724_n1303;
  wire _abc_15724_n1304;
  wire _abc_15724_n1305_1;
  wire _abc_15724_n1306_1;
  wire _abc_15724_n1307;
  wire _abc_15724_n1308_1;
  wire _abc_15724_n1309;
  wire _abc_15724_n1310;
  wire _abc_15724_n1311;
  wire _abc_15724_n1312;
  wire _abc_15724_n1313;
  wire _abc_15724_n1314;
  wire _abc_15724_n1315;
  wire _abc_15724_n1316;
  wire _abc_15724_n1317;
  wire _abc_15724_n1318;
  wire _abc_15724_n1319_1;
  wire _abc_15724_n1320_1;
  wire _abc_15724_n1322;
  wire _abc_15724_n1323;
  wire _abc_15724_n1324;
  wire _abc_15724_n1325;
  wire _abc_15724_n1326;
  wire _abc_15724_n1327;
  wire _abc_15724_n1328;
  wire _abc_15724_n1329_1;
  wire _abc_15724_n1330_1;
  wire _abc_15724_n1331;
  wire _abc_15724_n1332_1;
  wire _abc_15724_n1333;
  wire _abc_15724_n1334;
  wire _abc_15724_n1336;
  wire _abc_15724_n1337;
  wire _abc_15724_n1338;
  wire _abc_15724_n1339;
  wire _abc_15724_n1340_1;
  wire _abc_15724_n1341_1;
  wire _abc_15724_n1342;
  wire _abc_15724_n1343_1;
  wire _abc_15724_n1344;
  wire _abc_15724_n1345;
  wire _abc_15724_n1346;
  wire _abc_15724_n1347;
  wire _abc_15724_n1348;
  wire _abc_15724_n1349;
  wire _abc_15724_n1350_1;
  wire _abc_15724_n1352_1;
  wire _abc_15724_n1353;
  wire _abc_15724_n1354;
  wire _abc_15724_n1355;
  wire _abc_15724_n1356;
  wire _abc_15724_n1357;
  wire _abc_15724_n1358;
  wire _abc_15724_n1359;
  wire _abc_15724_n1360;
  wire _abc_15724_n1361;
  wire _abc_15724_n1362;
  wire _abc_15724_n1363;
  wire _abc_15724_n1365;
  wire _abc_15724_n1366;
  wire _abc_15724_n1367;
  wire _abc_15724_n1368_1;
  wire _abc_15724_n1369_1;
  wire _abc_15724_n1370;
  wire _abc_15724_n1371_1;
  wire _abc_15724_n1372;
  wire _abc_15724_n1373;
  wire _abc_15724_n1374;
  wire _abc_15724_n1375;
  wire _abc_15724_n1376;
  wire _abc_15724_n1377_1;
  wire _abc_15724_n1378_1;
  wire _abc_15724_n1379_1;
  wire _abc_15724_n1380;
  wire _abc_15724_n1381;
  wire _abc_15724_n1382;
  wire _abc_15724_n1383;
  wire _abc_15724_n1384;
  wire _abc_15724_n1385;
  wire _abc_15724_n1386;
  wire _abc_15724_n1387;
  wire _abc_15724_n1388;
  wire _abc_15724_n1390_1;
  wire _abc_15724_n1391_1;
  wire _abc_15724_n1392;
  wire _abc_15724_n1393_1;
  wire _abc_15724_n1394;
  wire _abc_15724_n1395;
  wire _abc_15724_n1396;
  wire _abc_15724_n1397;
  wire _abc_15724_n1398;
  wire _abc_15724_n1399_1;
  wire _abc_15724_n1400_1;
  wire _abc_15724_n1401;
  wire _abc_15724_n1402_1;
  wire _abc_15724_n1403;
  wire _abc_15724_n1404;
  wire _abc_15724_n1405;
  wire _abc_15724_n1406;
  wire _abc_15724_n1407;
  wire _abc_15724_n1408;
  wire _abc_15724_n1409;
  wire _abc_15724_n1410;
  wire _abc_15724_n1411;
  wire _abc_15724_n1412;
  wire _abc_15724_n1413_1;
  wire _abc_15724_n1415;
  wire _abc_15724_n1416_1;
  wire _abc_15724_n1417;
  wire _abc_15724_n1418;
  wire _abc_15724_n1419;
  wire _abc_15724_n1420;
  wire _abc_15724_n1421;
  wire _abc_15724_n1422_1;
  wire _abc_15724_n1423_1;
  wire _abc_15724_n1424_1;
  wire _abc_15724_n1425;
  wire _abc_15724_n1426;
  wire _abc_15724_n1427;
  wire _abc_15724_n1428;
  wire _abc_15724_n1430;
  wire _abc_15724_n1431;
  wire _abc_15724_n1432;
  wire _abc_15724_n1433;
  wire _abc_15724_n1434;
  wire _abc_15724_n1435_1;
  wire _abc_15724_n1436_1;
  wire _abc_15724_n1437;
  wire _abc_15724_n1438_1;
  wire _abc_15724_n1439;
  wire _abc_15724_n1440;
  wire _abc_15724_n1441;
  wire _abc_15724_n1442;
  wire _abc_15724_n1443;
  wire _abc_15724_n1444_1;
  wire _abc_15724_n1445_1;
  wire _abc_15724_n1447;
  wire _abc_15724_n1448;
  wire _abc_15724_n1449;
  wire _abc_15724_n1450;
  wire _abc_15724_n1451;
  wire _abc_15724_n1452;
  wire _abc_15724_n1453;
  wire _abc_15724_n1454;
  wire _abc_15724_n1455;
  wire _abc_15724_n1456;
  wire _abc_15724_n1457;
  wire _abc_15724_n1458;
  wire _abc_15724_n1459;
  wire _abc_15724_n1460;
  wire _abc_15724_n1461;
  wire _abc_15724_n1462_1;
  wire _abc_15724_n1464_1;
  wire _abc_15724_n1465;
  wire _abc_15724_n1466;
  wire _abc_15724_n1467;
  wire _abc_15724_n1468;
  wire _abc_15724_n1469;
  wire _abc_15724_n1470;
  wire _abc_15724_n1471;
  wire _abc_15724_n1472_1;
  wire _abc_15724_n1473_1;
  wire _abc_15724_n1474_1;
  wire _abc_15724_n1475;
  wire _abc_15724_n1476;
  wire _abc_15724_n1477;
  wire _abc_15724_n1479;
  wire _abc_15724_n1480;
  wire _abc_15724_n1481;
  wire _abc_15724_n1482;
  wire _abc_15724_n1483;
  wire _abc_15724_n1484_1;
  wire _abc_15724_n1485_1;
  wire _abc_15724_n1486;
  wire _abc_15724_n1487_1;
  wire _abc_15724_n1488;
  wire _abc_15724_n1489;
  wire _abc_15724_n1490;
  wire _abc_15724_n1491;
  wire _abc_15724_n1492;
  wire _abc_15724_n1493_1;
  wire _abc_15724_n1495;
  wire _abc_15724_n1496_1;
  wire _abc_15724_n1497;
  wire _abc_15724_n1498;
  wire _abc_15724_n1499;
  wire _abc_15724_n1500;
  wire _abc_15724_n1501;
  wire _abc_15724_n1502;
  wire _abc_15724_n1503;
  wire _abc_15724_n1504;
  wire _abc_15724_n1505;
  wire _abc_15724_n1506;
  wire _abc_15724_n1507;
  wire _abc_15724_n1509_1;
  wire _abc_15724_n1510_1;
  wire _abc_15724_n1511;
  wire _abc_15724_n1512;
  wire _abc_15724_n1513;
  wire _abc_15724_n1514;
  wire _abc_15724_n1515;
  wire _abc_15724_n1517;
  wire _abc_15724_n1518_1;
  wire _abc_15724_n1519_1;
  wire _abc_15724_n1520_1;
  wire _abc_15724_n1521;
  wire _abc_15724_n1522;
  wire _abc_15724_n1523;
  wire _abc_15724_n1524;
  wire _abc_15724_n1525;
  wire _abc_15724_n1526;
  wire _abc_15724_n1527;
  wire _abc_15724_n1529;
  wire _abc_15724_n1530_1;
  wire _abc_15724_n1531_1;
  wire _abc_15724_n1532;
  wire _abc_15724_n1533_1;
  wire _abc_15724_n1534;
  wire _abc_15724_n1535;
  wire _abc_15724_n1536;
  wire _abc_15724_n1537;
  wire _abc_15724_n1538_1;
  wire _abc_15724_n1539;
  wire _abc_15724_n1540_1;
  wire _abc_15724_n1541;
  wire _abc_15724_n1543_1;
  wire _abc_15724_n1544;
  wire _abc_15724_n1545;
  wire _abc_15724_n1546;
  wire _abc_15724_n1547;
  wire _abc_15724_n1548_1;
  wire _abc_15724_n1549;
  wire _abc_15724_n1550_1;
  wire _abc_15724_n1551;
  wire _abc_15724_n1552;
  wire _abc_15724_n1553;
  wire _abc_15724_n1554;
  wire _abc_15724_n1555;
  wire _abc_15724_n1557_1;
  wire _abc_15724_n1558;
  wire _abc_15724_n1559;
  wire _abc_15724_n1560;
  wire _abc_15724_n1561;
  wire _abc_15724_n1562;
  wire _abc_15724_n1563_1;
  wire _abc_15724_n1564_1;
  wire _abc_15724_n1565;
  wire _abc_15724_n1566;
  wire _abc_15724_n1567;
  wire _abc_15724_n1568;
  wire _abc_15724_n1569;
  wire _abc_15724_n1570_1;
  wire _abc_15724_n1571_1;
  wire _abc_15724_n1573_1;
  wire _abc_15724_n1574;
  wire _abc_15724_n1575;
  wire _abc_15724_n1576;
  wire _abc_15724_n1577;
  wire _abc_15724_n1578_1;
  wire _abc_15724_n1579_1;
  wire _abc_15724_n1580;
  wire _abc_15724_n1581_1;
  wire _abc_15724_n1582;
  wire _abc_15724_n1583;
  wire _abc_15724_n1584_1;
  wire _abc_15724_n1585_1;
  wire _abc_15724_n1587_1;
  wire _abc_15724_n1588;
  wire _abc_15724_n1589;
  wire _abc_15724_n1590_1;
  wire _abc_15724_n1591_1;
  wire _abc_15724_n1592;
  wire _abc_15724_n1593_1;
  wire _abc_15724_n1594;
  wire _abc_15724_n1595;
  wire _abc_15724_n1596_1;
  wire _abc_15724_n1597_1;
  wire _abc_15724_n1598;
  wire _abc_15724_n1599_1;
  wire _abc_15724_n1601;
  wire _abc_15724_n1602_1;
  wire _abc_15724_n1603_1;
  wire _abc_15724_n1604;
  wire _abc_15724_n1605;
  wire _abc_15724_n1606;
  wire _abc_15724_n1607;
  wire _abc_15724_n1608;
  wire _abc_15724_n1609_1;
  wire _abc_15724_n1610_1;
  wire _abc_15724_n1611;
  wire _abc_15724_n1612;
  wire _abc_15724_n1613;
  wire _abc_15724_n1615;
  wire _abc_15724_n1616_1;
  wire _abc_15724_n1617_1;
  wire _abc_15724_n1618;
  wire _abc_15724_n1619;
  wire _abc_15724_n1620;
  wire _abc_15724_n1621;
  wire _abc_15724_n1622;
  wire _abc_15724_n1623_1;
  wire _abc_15724_n1624_1;
  wire _abc_15724_n1625;
  wire _abc_15724_n1626;
  wire _abc_15724_n1627;
  wire _abc_15724_n1628;
  wire _abc_15724_n1629;
  wire _abc_15724_n1631_1;
  wire _abc_15724_n1632;
  wire _abc_15724_n1633_1;
  wire _abc_15724_n1634;
  wire _abc_15724_n1635;
  wire _abc_15724_n1636_1;
  wire _abc_15724_n1637_1;
  wire _abc_15724_n1638;
  wire _abc_15724_n1639_1;
  wire _abc_15724_n1640;
  wire _abc_15724_n1641;
  wire _abc_15724_n1642_1;
  wire _abc_15724_n1644;
  wire _abc_15724_n1645_1;
  wire _abc_15724_n1646;
  wire _abc_15724_n1647;
  wire _abc_15724_n1648_1;
  wire _abc_15724_n1649_1;
  wire _abc_15724_n1650;
  wire _abc_15724_n1651;
  wire _abc_15724_n1652;
  wire _abc_15724_n1653;
  wire _abc_15724_n1654;
  wire _abc_15724_n1655_1;
  wire _abc_15724_n1656_1;
  wire _abc_15724_n1658_1;
  wire _abc_15724_n1659;
  wire _abc_15724_n1660;
  wire _abc_15724_n1661_1;
  wire _abc_15724_n1662_1;
  wire _abc_15724_n1663;
  wire _abc_15724_n1664;
  wire _abc_15724_n1665;
  wire _abc_15724_n1666;
  wire _abc_15724_n1667;
  wire _abc_15724_n1668_1;
  wire _abc_15724_n1669_1;
  wire _abc_15724_n1670;
  wire _abc_15724_n1672;
  wire _abc_15724_n1673;
  wire _abc_15724_n1674;
  wire _abc_15724_n1675_1;
  wire _abc_15724_n1676_1;
  wire _abc_15724_n1677;
  wire _abc_15724_n1678_1;
  wire _abc_15724_n1679;
  wire _abc_15724_n1680;
  wire _abc_15724_n1681_1;
  wire _abc_15724_n1682_1;
  wire _abc_15724_n1683;
  wire _abc_15724_n1684;
  wire _abc_15724_n1685;
  wire _abc_15724_n1686;
  wire _abc_15724_n1687;
  wire _abc_15724_n1688_1;
  wire _abc_15724_n1689;
  wire _abc_15724_n1690;
  wire _abc_15724_n1691;
  wire _abc_15724_n1692_1;
  wire _abc_15724_n1693;
  wire _abc_15724_n1694;
  wire _abc_15724_n1695;
  wire _abc_15724_n1696_1;
  wire _abc_15724_n1698;
  wire _abc_15724_n1699;
  wire _abc_15724_n1700_1;
  wire _abc_15724_n1701;
  wire _abc_15724_n1702;
  wire _abc_15724_n1703;
  wire _abc_15724_n1704_1;
  wire _abc_15724_n1705;
  wire _abc_15724_n1706;
  wire _abc_15724_n1707;
  wire _abc_15724_n1708;
  wire _abc_15724_n1709_1;
  wire _abc_15724_n1711;
  wire _abc_15724_n1712;
  wire _abc_15724_n1713;
  wire _abc_15724_n1714_1;
  wire _abc_15724_n1715;
  wire _abc_15724_n1716;
  wire _abc_15724_n1717;
  wire _abc_15724_n1718;
  wire _abc_15724_n1719_1;
  wire _abc_15724_n1720;
  wire _abc_15724_n1721;
  wire _abc_15724_n1722;
  wire _abc_15724_n1723;
  wire _abc_15724_n1725;
  wire _abc_15724_n1726;
  wire _abc_15724_n1727;
  wire _abc_15724_n1728_1;
  wire _abc_15724_n1729;
  wire _abc_15724_n1730;
  wire _abc_15724_n1731;
  wire _abc_15724_n1732_1;
  wire _abc_15724_n1733;
  wire _abc_15724_n1734;
  wire _abc_15724_n1735;
  wire _abc_15724_n1736;
  wire _abc_15724_n1737_1;
  wire _abc_15724_n1739;
  wire _abc_15724_n1740;
  wire _abc_15724_n1741_1;
  wire _abc_15724_n1742;
  wire _abc_15724_n1743;
  wire _abc_15724_n1744;
  wire _abc_15724_n1745_1;
  wire _abc_15724_n1746;
  wire _abc_15724_n1747;
  wire _abc_15724_n1748;
  wire _abc_15724_n1749;
  wire _abc_15724_n1750_1;
  wire _abc_15724_n1751;
  wire _abc_15724_n1752;
  wire _abc_15724_n1753;
  wire _abc_15724_n1754_1;
  wire _abc_15724_n1755;
  wire _abc_15724_n1756;
  wire _abc_15724_n1757;
  wire _abc_15724_n1758_1;
  wire _abc_15724_n1759;
  wire _abc_15724_n1760;
  wire _abc_15724_n1761;
  wire _abc_15724_n1762_1;
  wire _abc_15724_n1764;
  wire _abc_15724_n1765;
  wire _abc_15724_n1766;
  wire _abc_15724_n1767_1;
  wire _abc_15724_n1768;
  wire _abc_15724_n1769;
  wire _abc_15724_n1770;
  wire _abc_15724_n1771;
  wire _abc_15724_n1772_1;
  wire _abc_15724_n1773;
  wire _abc_15724_n1774;
  wire _abc_15724_n1775;
  wire _abc_15724_n1776;
  wire _abc_15724_n1778;
  wire _abc_15724_n1779;
  wire _abc_15724_n1780;
  wire _abc_15724_n1781_1;
  wire _abc_15724_n1782;
  wire _abc_15724_n1783;
  wire _abc_15724_n1784;
  wire _abc_15724_n1785;
  wire _abc_15724_n1786_1;
  wire _abc_15724_n1787;
  wire _abc_15724_n1788;
  wire _abc_15724_n1789;
  wire _abc_15724_n1790_1;
  wire _abc_15724_n1791;
  wire _abc_15724_n1792;
  wire _abc_15724_n1793;
  wire _abc_15724_n1795_1;
  wire _abc_15724_n1796;
  wire _abc_15724_n1797;
  wire _abc_15724_n1798;
  wire _abc_15724_n1799_1;
  wire _abc_15724_n1800;
  wire _abc_15724_n1801;
  wire _abc_15724_n1802;
  wire _abc_15724_n1803;
  wire _abc_15724_n1804_1;
  wire _abc_15724_n1805;
  wire _abc_15724_n1806;
  wire _abc_15724_n1807;
  wire _abc_15724_n1809_1;
  wire _abc_15724_n1810;
  wire _abc_15724_n1811;
  wire _abc_15724_n1812;
  wire _abc_15724_n1813_1;
  wire _abc_15724_n1814;
  wire _abc_15724_n1815;
  wire _abc_15724_n1816;
  wire _abc_15724_n1817;
  wire _abc_15724_n1818_1;
  wire _abc_15724_n1819;
  wire _abc_15724_n1820;
  wire _abc_15724_n1821;
  wire _abc_15724_n1822;
  wire _abc_15724_n1823_1;
  wire _abc_15724_n1824;
  wire _abc_15724_n1825;
  wire _abc_15724_n1826;
  wire _abc_15724_n1827_1;
  wire _abc_15724_n1828;
  wire _abc_15724_n1829;
  wire _abc_15724_n1830;
  wire _abc_15724_n1832;
  wire _abc_15724_n1833;
  wire _abc_15724_n1834;
  wire _abc_15724_n1835;
  wire _abc_15724_n1836_1;
  wire _abc_15724_n1837;
  wire _abc_15724_n1838;
  wire _abc_15724_n1839;
  wire _abc_15724_n1840;
  wire _abc_15724_n1841_1;
  wire _abc_15724_n1842;
  wire _abc_15724_n1843;
  wire _abc_15724_n1844;
  wire _abc_15724_n1846_1;
  wire _abc_15724_n1847;
  wire _abc_15724_n1848;
  wire _abc_15724_n1849;
  wire _abc_15724_n1850;
  wire _abc_15724_n1851_1;
  wire _abc_15724_n1852;
  wire _abc_15724_n1853;
  wire _abc_15724_n1854;
  wire _abc_15724_n1855;
  wire _abc_15724_n1856_1;
  wire _abc_15724_n1857;
  wire _abc_15724_n1858;
  wire _abc_15724_n1859;
  wire _abc_15724_n1860;
  wire _abc_15724_n1861_1;
  wire _abc_15724_n1863;
  wire _abc_15724_n1864;
  wire _abc_15724_n1865_1;
  wire _abc_15724_n1866;
  wire _abc_15724_n1867;
  wire _abc_15724_n1868;
  wire _abc_15724_n1869;
  wire _abc_15724_n1870_1;
  wire _abc_15724_n1871;
  wire _abc_15724_n1872;
  wire _abc_15724_n1873;
  wire _abc_15724_n1874;
  wire _abc_15724_n1875_1;
  wire _abc_15724_n1877;
  wire _abc_15724_n1878;
  wire _abc_15724_n1879;
  wire _abc_15724_n1880_1;
  wire _abc_15724_n1881;
  wire _abc_15724_n1882;
  wire _abc_15724_n1883;
  wire _abc_15724_n1884;
  wire _abc_15724_n1885_1;
  wire _abc_15724_n1886;
  wire _abc_15724_n1887;
  wire _abc_15724_n1888;
  wire _abc_15724_n1889_1;
  wire _abc_15724_n1890;
  wire _abc_15724_n1891;
  wire _abc_15724_n1892;
  wire _abc_15724_n1893_1;
  wire _abc_15724_n1894;
  wire _abc_15724_n1895;
  wire _abc_15724_n1896;
  wire _abc_15724_n1897_1;
  wire _abc_15724_n1899;
  wire _abc_15724_n1900;
  wire _abc_15724_n1901_1;
  wire _abc_15724_n1902;
  wire _abc_15724_n1903;
  wire _abc_15724_n1904;
  wire _abc_15724_n1905_1;
  wire _abc_15724_n1906;
  wire _abc_15724_n1907;
  wire _abc_15724_n1908;
  wire _abc_15724_n1909_1;
  wire _abc_15724_n1910;
  wire _abc_15724_n1911;
  wire _abc_15724_n1912;
  wire _abc_15724_n1913_1;
  wire _abc_15724_n1915;
  wire _abc_15724_n1916;
  wire _abc_15724_n1917;
  wire _abc_15724_n1918_1;
  wire _abc_15724_n1919;
  wire _abc_15724_n1920;
  wire _abc_15724_n1921;
  wire _abc_15724_n1922;
  wire _abc_15724_n1923_1;
  wire _abc_15724_n1924;
  wire _abc_15724_n1925;
  wire _abc_15724_n1926;
  wire _abc_15724_n1927_1;
  wire _abc_15724_n1929;
  wire _abc_15724_n1930;
  wire _abc_15724_n1931_1;
  wire _abc_15724_n1932;
  wire _abc_15724_n1933;
  wire _abc_15724_n1934;
  wire _abc_15724_n1935_1;
  wire _abc_15724_n1936;
  wire _abc_15724_n1937;
  wire _abc_15724_n1938;
  wire _abc_15724_n1939;
  wire _abc_15724_n1940_1;
  wire _abc_15724_n1941;
  wire _abc_15724_n1943;
  wire _abc_15724_n1944_1;
  wire _abc_15724_n1945;
  wire _abc_15724_n1946;
  wire _abc_15724_n1947;
  wire _abc_15724_n1948_1;
  wire _abc_15724_n1949;
  wire _abc_15724_n1950;
  wire _abc_15724_n1951;
  wire _abc_15724_n1952;
  wire _abc_15724_n1953_1;
  wire _abc_15724_n1954;
  wire _abc_15724_n1955;
  wire _abc_15724_n1956;
  wire _abc_15724_n1957_1;
  wire _abc_15724_n1958;
  wire _abc_15724_n1959;
  wire _abc_15724_n1960;
  wire _abc_15724_n1961;
  wire _abc_15724_n1962_1;
  wire _abc_15724_n1963;
  wire _abc_15724_n1964;
  wire _abc_15724_n1965;
  wire _abc_15724_n1967;
  wire _abc_15724_n1968;
  wire _abc_15724_n1969;
  wire _abc_15724_n1970_1;
  wire _abc_15724_n1971;
  wire _abc_15724_n1972;
  wire _abc_15724_n1973;
  wire _abc_15724_n1974_1;
  wire _abc_15724_n1975;
  wire _abc_15724_n1976;
  wire _abc_15724_n1977;
  wire _abc_15724_n1978;
  wire _abc_15724_n1980;
  wire _abc_15724_n1981;
  wire _abc_15724_n1982;
  wire _abc_15724_n1983_1;
  wire _abc_15724_n1984;
  wire _abc_15724_n1985;
  wire _abc_15724_n1986;
  wire _abc_15724_n1987;
  wire _abc_15724_n1988_1;
  wire _abc_15724_n1989;
  wire _abc_15724_n1990;
  wire _abc_15724_n1991;
  wire _abc_15724_n1992;
  wire _abc_15724_n1993_1;
  wire _abc_15724_n1994;
  wire _abc_15724_n1995;
  wire _abc_15724_n1996;
  wire _abc_15724_n1997;
  wire _abc_15724_n1999;
  wire _abc_15724_n2000;
  wire _abc_15724_n2001;
  wire _abc_15724_n2002_1;
  wire _abc_15724_n2003;
  wire _abc_15724_n2004;
  wire _abc_15724_n2005;
  wire _abc_15724_n2006_1;
  wire _abc_15724_n2007;
  wire _abc_15724_n2008;
  wire _abc_15724_n2009;
  wire _abc_15724_n2010;
  wire _abc_15724_n2011_1;
  wire _abc_15724_n2012;
  wire _abc_15724_n2014;
  wire _abc_15724_n2015;
  wire _abc_15724_n2016_1;
  wire _abc_15724_n2017;
  wire _abc_15724_n2018;
  wire _abc_15724_n2019;
  wire _abc_15724_n2020_1;
  wire _abc_15724_n2022;
  wire _abc_15724_n2023;
  wire _abc_15724_n2024_1;
  wire _abc_15724_n2025;
  wire _abc_15724_n2026;
  wire _abc_15724_n2027;
  wire _abc_15724_n2028;
  wire _abc_15724_n2029_1;
  wire _abc_15724_n2030;
  wire _abc_15724_n2031;
  wire _abc_15724_n2033;
  wire _abc_15724_n2034_1;
  wire _abc_15724_n2035;
  wire _abc_15724_n2036;
  wire _abc_15724_n2037;
  wire _abc_15724_n2038_1;
  wire _abc_15724_n2039;
  wire _abc_15724_n2040;
  wire _abc_15724_n2041;
  wire _abc_15724_n2042;
  wire _abc_15724_n2043_1;
  wire _abc_15724_n2044;
  wire _abc_15724_n2046;
  wire _abc_15724_n2047;
  wire _abc_15724_n2048_1;
  wire _abc_15724_n2049;
  wire _abc_15724_n2050;
  wire _abc_15724_n2051;
  wire _abc_15724_n2052;
  wire _abc_15724_n2053_1;
  wire _abc_15724_n2054;
  wire _abc_15724_n2055;
  wire _abc_15724_n2056;
  wire _abc_15724_n2057_1;
  wire _abc_15724_n2058;
  wire _abc_15724_n2060;
  wire _abc_15724_n2061_1;
  wire _abc_15724_n2062;
  wire _abc_15724_n2063;
  wire _abc_15724_n2064;
  wire _abc_15724_n2065_1;
  wire _abc_15724_n2066;
  wire _abc_15724_n2067;
  wire _abc_15724_n2068;
  wire _abc_15724_n2069;
  wire _abc_15724_n2070_1;
  wire _abc_15724_n2071;
  wire _abc_15724_n2073;
  wire _abc_15724_n2074_1;
  wire _abc_15724_n2075;
  wire _abc_15724_n2076;
  wire _abc_15724_n2077;
  wire _abc_15724_n2078;
  wire _abc_15724_n2079_1;
  wire _abc_15724_n2080;
  wire _abc_15724_n2081;
  wire _abc_15724_n2082;
  wire _abc_15724_n2083_1;
  wire _abc_15724_n2085;
  wire _abc_15724_n2086;
  wire _abc_15724_n2087;
  wire _abc_15724_n2088_1;
  wire _abc_15724_n2089;
  wire _abc_15724_n2090;
  wire _abc_15724_n2091;
  wire _abc_15724_n2092_1;
  wire _abc_15724_n2093;
  wire _abc_15724_n2094;
  wire _abc_15724_n2095;
  wire _abc_15724_n2097;
  wire _abc_15724_n2098;
  wire _abc_15724_n2099;
  wire _abc_15724_n2100;
  wire _abc_15724_n2101_1;
  wire _abc_15724_n2102;
  wire _abc_15724_n2103;
  wire _abc_15724_n2104;
  wire _abc_15724_n2105_1;
  wire _abc_15724_n2106;
  wire _abc_15724_n2107;
  wire _abc_15724_n2108;
  wire _abc_15724_n2109_1;
  wire _abc_15724_n2111;
  wire _abc_15724_n2112;
  wire _abc_15724_n2113;
  wire _abc_15724_n2114_1;
  wire _abc_15724_n2115;
  wire _abc_15724_n2116;
  wire _abc_15724_n2117;
  wire _abc_15724_n2118;
  wire _abc_15724_n2119_1;
  wire _abc_15724_n2120;
  wire _abc_15724_n2121;
  wire _abc_15724_n2122;
  wire _abc_15724_n2123_1;
  wire _abc_15724_n2125;
  wire _abc_15724_n2126;
  wire _abc_15724_n2127_1;
  wire _abc_15724_n2128;
  wire _abc_15724_n2129;
  wire _abc_15724_n2130;
  wire _abc_15724_n2131_1;
  wire _abc_15724_n2132;
  wire _abc_15724_n2133;
  wire _abc_15724_n2134;
  wire _abc_15724_n2135_1;
  wire _abc_15724_n2136;
  wire _abc_15724_n2137;
  wire _abc_15724_n2139_1;
  wire _abc_15724_n2140;
  wire _abc_15724_n2141;
  wire _abc_15724_n2142;
  wire _abc_15724_n2143_1;
  wire _abc_15724_n2144;
  wire _abc_15724_n2145;
  wire _abc_15724_n2146;
  wire _abc_15724_n2147;
  wire _abc_15724_n2148_1;
  wire _abc_15724_n2149;
  wire _abc_15724_n2150;
  wire _abc_15724_n2151;
  wire _abc_15724_n2152_1;
  wire _abc_15724_n2153;
  wire _abc_15724_n2154;
  wire _abc_15724_n2156_1;
  wire _abc_15724_n2157;
  wire _abc_15724_n2158;
  wire _abc_15724_n2159;
  wire _abc_15724_n2160_1;
  wire _abc_15724_n2161;
  wire _abc_15724_n2162;
  wire _abc_15724_n2163_1;
  wire _abc_15724_n2164;
  wire _abc_15724_n2165;
  wire _abc_15724_n2166;
  wire _abc_15724_n2167;
  wire _abc_15724_n2168_1;
  wire _abc_15724_n2170;
  wire _abc_15724_n2171_1;
  wire _abc_15724_n2172_1;
  wire _abc_15724_n2173;
  wire _abc_15724_n2174;
  wire _abc_15724_n2175;
  wire _abc_15724_n2176;
  wire _abc_15724_n2177;
  wire _abc_15724_n2178;
  wire _abc_15724_n2179;
  wire _abc_15724_n2180_1;
  wire _abc_15724_n2181;
  wire _abc_15724_n2182_1;
  wire _abc_15724_n2183;
  wire _abc_15724_n2184;
  wire _abc_15724_n2185;
  wire _abc_15724_n2186;
  wire _abc_15724_n2187;
  wire _abc_15724_n2189;
  wire _abc_15724_n2190;
  wire _abc_15724_n2191;
  wire _abc_15724_n2192;
  wire _abc_15724_n2193;
  wire _abc_15724_n2194;
  wire _abc_15724_n2195_1;
  wire _abc_15724_n2196;
  wire _abc_15724_n2197;
  wire _abc_15724_n2198;
  wire _abc_15724_n2199;
  wire _abc_15724_n2200;
  wire _abc_15724_n2201;
  wire _abc_15724_n2203;
  wire _abc_15724_n2204;
  wire _abc_15724_n2205;
  wire _abc_15724_n2206;
  wire _abc_15724_n2207;
  wire _abc_15724_n2208;
  wire _abc_15724_n2209;
  wire _abc_15724_n2210;
  wire _abc_15724_n2211;
  wire _abc_15724_n2212;
  wire _abc_15724_n2213;
  wire _abc_15724_n2214;
  wire _abc_15724_n2215;
  wire _abc_15724_n2216;
  wire _abc_15724_n2217;
  wire _abc_15724_n2218;
  wire _abc_15724_n2220;
  wire _abc_15724_n2221;
  wire _abc_15724_n2222;
  wire _abc_15724_n2223;
  wire _abc_15724_n2224;
  wire _abc_15724_n2225;
  wire _abc_15724_n2226;
  wire _abc_15724_n2227;
  wire _abc_15724_n2228;
  wire _abc_15724_n2229;
  wire _abc_15724_n2230;
  wire _abc_15724_n2231;
  wire _abc_15724_n2232;
  wire _abc_15724_n2234;
  wire _abc_15724_n2235;
  wire _abc_15724_n2236;
  wire _abc_15724_n2237;
  wire _abc_15724_n2238;
  wire _abc_15724_n2239;
  wire _abc_15724_n2240;
  wire _abc_15724_n2241;
  wire _abc_15724_n2242;
  wire _abc_15724_n2243;
  wire _abc_15724_n2244;
  wire _abc_15724_n2245;
  wire _abc_15724_n2246_1;
  wire _abc_15724_n2247;
  wire _abc_15724_n2248;
  wire _abc_15724_n2249;
  wire _abc_15724_n2250_1;
  wire _abc_15724_n2251;
  wire _abc_15724_n2252;
  wire _abc_15724_n2254;
  wire _abc_15724_n2255;
  wire _abc_15724_n2256;
  wire _abc_15724_n2257;
  wire _abc_15724_n2258;
  wire _abc_15724_n2259;
  wire _abc_15724_n2260;
  wire _abc_15724_n2261;
  wire _abc_15724_n2262;
  wire _abc_15724_n2263;
  wire _abc_15724_n2264;
  wire _abc_15724_n2265;
  wire _abc_15724_n2267;
  wire _abc_15724_n2268;
  wire _abc_15724_n2269;
  wire _abc_15724_n2270;
  wire _abc_15724_n2271;
  wire _abc_15724_n2272;
  wire _abc_15724_n2273;
  wire _abc_15724_n2274;
  wire _abc_15724_n2275;
  wire _abc_15724_n2276;
  wire _abc_15724_n2277;
  wire _abc_15724_n2278;
  wire _abc_15724_n2279;
  wire _abc_15724_n2281;
  wire _abc_15724_n2282;
  wire _abc_15724_n2283;
  wire _abc_15724_n2284;
  wire _abc_15724_n2285;
  wire _abc_15724_n2286;
  wire _abc_15724_n2287_1;
  wire _abc_15724_n2288;
  wire _abc_15724_n2289;
  wire _abc_15724_n2290;
  wire _abc_15724_n2291_1;
  wire _abc_15724_n2292;
  wire _abc_15724_n2293;
  wire _abc_15724_n2295;
  wire _abc_15724_n2296;
  wire _abc_15724_n2297;
  wire _abc_15724_n2298;
  wire _abc_15724_n2299;
  wire _abc_15724_n2300;
  wire _abc_15724_n2301;
  wire _abc_15724_n2302;
  wire _abc_15724_n2303;
  wire _abc_15724_n2304;
  wire _abc_15724_n2305;
  wire _abc_15724_n2306;
  wire _abc_15724_n2307;
  wire _abc_15724_n2308;
  wire _abc_15724_n2309;
  wire _abc_15724_n2310;
  wire _abc_15724_n2311;
  wire _abc_15724_n2312;
  wire _abc_15724_n2313;
  wire _abc_15724_n2314;
  wire _abc_15724_n2315;
  wire _abc_15724_n2317;
  wire _abc_15724_n2318;
  wire _abc_15724_n2319;
  wire _abc_15724_n2320;
  wire _abc_15724_n2321;
  wire _abc_15724_n2322;
  wire _abc_15724_n2323;
  wire _abc_15724_n2324;
  wire _abc_15724_n2325;
  wire _abc_15724_n2326_1;
  wire _abc_15724_n2327;
  wire _abc_15724_n2329;
  wire _abc_15724_n2330_1;
  wire _abc_15724_n2331;
  wire _abc_15724_n2332;
  wire _abc_15724_n2333;
  wire _abc_15724_n2334;
  wire _abc_15724_n2335;
  wire _abc_15724_n2336;
  wire _abc_15724_n2337;
  wire _abc_15724_n2338;
  wire _abc_15724_n2339;
  wire _abc_15724_n2340;
  wire _abc_15724_n2342;
  wire _abc_15724_n2343;
  wire _abc_15724_n2344;
  wire _abc_15724_n2345;
  wire _abc_15724_n2346;
  wire _abc_15724_n2347;
  wire _abc_15724_n2348;
  wire _abc_15724_n2349;
  wire _abc_15724_n2350;
  wire _abc_15724_n2351;
  wire _abc_15724_n2352;
  wire _abc_15724_n2353;
  wire _abc_15724_n2354;
  wire _abc_15724_n2356;
  wire _abc_15724_n2357;
  wire _abc_15724_n2358;
  wire _abc_15724_n2359;
  wire _abc_15724_n2360;
  wire _abc_15724_n2361;
  wire _abc_15724_n2362;
  wire _abc_15724_n2363;
  wire _abc_15724_n2364;
  wire _abc_15724_n2365;
  wire _abc_15724_n2366_1;
  wire _abc_15724_n2367;
  wire _abc_15724_n2368;
  wire _abc_15724_n2369;
  wire _abc_15724_n2370_1;
  wire _abc_15724_n2371;
  wire _abc_15724_n2372;
  wire _abc_15724_n2373;
  wire _abc_15724_n2374;
  wire _abc_15724_n2375;
  wire _abc_15724_n2376;
  wire _abc_15724_n2377;
  wire _abc_15724_n2378;
  wire _abc_15724_n2379;
  wire _abc_15724_n2380;
  wire _abc_15724_n2382;
  wire _abc_15724_n2383;
  wire _abc_15724_n2384;
  wire _abc_15724_n2385;
  wire _abc_15724_n2386;
  wire _abc_15724_n2387;
  wire _abc_15724_n2388;
  wire _abc_15724_n2389;
  wire _abc_15724_n2390;
  wire _abc_15724_n2391;
  wire _abc_15724_n2392;
  wire _abc_15724_n2393;
  wire _abc_15724_n2394;
  wire _abc_15724_n2396;
  wire _abc_15724_n2397;
  wire _abc_15724_n2398;
  wire _abc_15724_n2399;
  wire _abc_15724_n2400;
  wire _abc_15724_n2401;
  wire _abc_15724_n2402;
  wire _abc_15724_n2403;
  wire _abc_15724_n2404;
  wire _abc_15724_n2405;
  wire _abc_15724_n2406_1;
  wire _abc_15724_n2407;
  wire _abc_15724_n2408;
  wire _abc_15724_n2409;
  wire _abc_15724_n2410;
  wire _abc_15724_n2411;
  wire _abc_15724_n2413;
  wire _abc_15724_n2414;
  wire _abc_15724_n2415;
  wire _abc_15724_n2416;
  wire _abc_15724_n2417;
  wire _abc_15724_n2418;
  wire _abc_15724_n2419;
  wire _abc_15724_n2420;
  wire _abc_15724_n2421;
  wire _abc_15724_n2422;
  wire _abc_15724_n2423;
  wire _abc_15724_n2424;
  wire _abc_15724_n2425;
  wire _abc_15724_n2427;
  wire _abc_15724_n2428;
  wire _abc_15724_n2429;
  wire _abc_15724_n2430;
  wire _abc_15724_n2431;
  wire _abc_15724_n2432;
  wire _abc_15724_n2433;
  wire _abc_15724_n2434;
  wire _abc_15724_n2435;
  wire _abc_15724_n2436;
  wire _abc_15724_n2437;
  wire _abc_15724_n2438;
  wire _abc_15724_n2439;
  wire _abc_15724_n2440;
  wire _abc_15724_n2441;
  wire _abc_15724_n2442;
  wire _abc_15724_n2443;
  wire _abc_15724_n2444;
  wire _abc_15724_n2446;
  wire _abc_15724_n2447;
  wire _abc_15724_n2448;
  wire _abc_15724_n2449_1;
  wire _abc_15724_n2450;
  wire _abc_15724_n2451;
  wire _abc_15724_n2452;
  wire _abc_15724_n2453;
  wire _abc_15724_n2454;
  wire _abc_15724_n2455;
  wire _abc_15724_n2456;
  wire _abc_15724_n2457;
  wire _abc_15724_n2458;
  wire _abc_15724_n2460;
  wire _abc_15724_n2461;
  wire _abc_15724_n2462;
  wire _abc_15724_n2463;
  wire _abc_15724_n2464;
  wire _abc_15724_n2465;
  wire _abc_15724_n2466;
  wire _abc_15724_n2467;
  wire _abc_15724_n2468;
  wire _abc_15724_n2469;
  wire _abc_15724_n2470;
  wire _abc_15724_n2471;
  wire _abc_15724_n2472;
  wire _abc_15724_n2473;
  wire _abc_15724_n2474;
  wire _abc_15724_n2475;
  wire _abc_15724_n2477;
  wire _abc_15724_n2478;
  wire _abc_15724_n2479;
  wire _abc_15724_n2480;
  wire _abc_15724_n2481;
  wire _abc_15724_n2482;
  wire _abc_15724_n2483;
  wire _abc_15724_n2484_1;
  wire _abc_15724_n2485;
  wire _abc_15724_n2486;
  wire _abc_15724_n2487;
  wire _abc_15724_n2488_1;
  wire _abc_15724_n2489;
  wire _abc_15724_n2490;
  wire _abc_15724_n2492;
  wire _abc_15724_n2493;
  wire _abc_15724_n2494;
  wire _abc_15724_n2495;
  wire _abc_15724_n2496;
  wire _abc_15724_n2497;
  wire _abc_15724_n2498;
  wire _abc_15724_n2500;
  wire _abc_15724_n2501;
  wire _abc_15724_n2502;
  wire _abc_15724_n2503;
  wire _abc_15724_n2504;
  wire _abc_15724_n2505;
  wire _abc_15724_n2506;
  wire _abc_15724_n2507;
  wire _abc_15724_n2508;
  wire _abc_15724_n2509;
  wire _abc_15724_n2511;
  wire _abc_15724_n2512;
  wire _abc_15724_n2513;
  wire _abc_15724_n2514;
  wire _abc_15724_n2515;
  wire _abc_15724_n2516;
  wire _abc_15724_n2517;
  wire _abc_15724_n2518;
  wire _abc_15724_n2519;
  wire _abc_15724_n2520;
  wire _abc_15724_n2521;
  wire _abc_15724_n2522;
  wire _abc_15724_n2524_1;
  wire _abc_15724_n2525;
  wire _abc_15724_n2526;
  wire _abc_15724_n2527_1;
  wire _abc_15724_n2528;
  wire _abc_15724_n2529;
  wire _abc_15724_n2530;
  wire _abc_15724_n2531;
  wire _abc_15724_n2532;
  wire _abc_15724_n2533;
  wire _abc_15724_n2534;
  wire _abc_15724_n2535;
  wire _abc_15724_n2537;
  wire _abc_15724_n2538;
  wire _abc_15724_n2539;
  wire _abc_15724_n2540;
  wire _abc_15724_n2541;
  wire _abc_15724_n2542;
  wire _abc_15724_n2543;
  wire _abc_15724_n2544;
  wire _abc_15724_n2545;
  wire _abc_15724_n2546;
  wire _abc_15724_n2547;
  wire _abc_15724_n2548;
  wire _abc_15724_n2549;
  wire _abc_15724_n2550;
  wire _abc_15724_n2552;
  wire _abc_15724_n2553;
  wire _abc_15724_n2554;
  wire _abc_15724_n2555;
  wire _abc_15724_n2556;
  wire _abc_15724_n2557;
  wire _abc_15724_n2558;
  wire _abc_15724_n2559;
  wire _abc_15724_n2560;
  wire _abc_15724_n2561;
  wire _abc_15724_n2562;
  wire _abc_15724_n2563;
  wire _abc_15724_n2565;
  wire _abc_15724_n2566;
  wire _abc_15724_n2567;
  wire _abc_15724_n2568;
  wire _abc_15724_n2569;
  wire _abc_15724_n2570_1;
  wire _abc_15724_n2571;
  wire _abc_15724_n2572;
  wire _abc_15724_n2573_1;
  wire _abc_15724_n2574;
  wire _abc_15724_n2575;
  wire _abc_15724_n2576;
  wire _abc_15724_n2578;
  wire _abc_15724_n2579;
  wire _abc_15724_n2580;
  wire _abc_15724_n2581;
  wire _abc_15724_n2582;
  wire _abc_15724_n2583;
  wire _abc_15724_n2584;
  wire _abc_15724_n2585;
  wire _abc_15724_n2586;
  wire _abc_15724_n2587;
  wire _abc_15724_n2588;
  wire _abc_15724_n2589;
  wire _abc_15724_n2590;
  wire _abc_15724_n2591;
  wire _abc_15724_n2592;
  wire _abc_15724_n2594;
  wire _abc_15724_n2595;
  wire _abc_15724_n2596;
  wire _abc_15724_n2597;
  wire _abc_15724_n2598;
  wire _abc_15724_n2599;
  wire _abc_15724_n2600;
  wire _abc_15724_n2601;
  wire _abc_15724_n2602;
  wire _abc_15724_n2603;
  wire _abc_15724_n2604;
  wire _abc_15724_n2605;
  wire _abc_15724_n2606;
  wire _abc_15724_n2607_1;
  wire _abc_15724_n2609;
  wire _abc_15724_n2610;
  wire _abc_15724_n2611;
  wire _abc_15724_n2612_1;
  wire _abc_15724_n2613;
  wire _abc_15724_n2614;
  wire _abc_15724_n2615;
  wire _abc_15724_n2616;
  wire _abc_15724_n2617;
  wire _abc_15724_n2618;
  wire _abc_15724_n2619;
  wire _abc_15724_n2620;
  wire _abc_15724_n2621;
  wire _abc_15724_n2623;
  wire _abc_15724_n2624;
  wire _abc_15724_n2625;
  wire _abc_15724_n2626;
  wire _abc_15724_n2627;
  wire _abc_15724_n2628;
  wire _abc_15724_n2629;
  wire _abc_15724_n2630;
  wire _abc_15724_n2631;
  wire _abc_15724_n2632;
  wire _abc_15724_n2633;
  wire _abc_15724_n2634;
  wire _abc_15724_n2635;
  wire _abc_15724_n2636;
  wire _abc_15724_n2637;
  wire _abc_15724_n2638;
  wire _abc_15724_n2640;
  wire _abc_15724_n2641;
  wire _abc_15724_n2642;
  wire _abc_15724_n2643;
  wire _abc_15724_n2644;
  wire _abc_15724_n2645;
  wire _abc_15724_n2646;
  wire _abc_15724_n2647;
  wire _abc_15724_n2648_1;
  wire _abc_15724_n2649;
  wire _abc_15724_n2650;
  wire _abc_15724_n2651;
  wire _abc_15724_n2653;
  wire _abc_15724_n2654;
  wire _abc_15724_n2655;
  wire _abc_15724_n2656;
  wire _abc_15724_n2657;
  wire _abc_15724_n2658;
  wire _abc_15724_n2659;
  wire _abc_15724_n2660;
  wire _abc_15724_n2661;
  wire _abc_15724_n2662;
  wire _abc_15724_n2663;
  wire _abc_15724_n2664;
  wire _abc_15724_n2665;
  wire _abc_15724_n2666;
  wire _abc_15724_n2667;
  wire _abc_15724_n2668;
  wire _abc_15724_n2669;
  wire _abc_15724_n2670;
  wire _abc_15724_n2671;
  wire _abc_15724_n2672;
  wire _abc_15724_n2673;
  wire _abc_15724_n2675;
  wire _abc_15724_n2676;
  wire _abc_15724_n2677;
  wire _abc_15724_n2678;
  wire _abc_15724_n2679;
  wire _abc_15724_n2680;
  wire _abc_15724_n2681;
  wire _abc_15724_n2682;
  wire _abc_15724_n2683;
  wire _abc_15724_n2684;
  wire _abc_15724_n2685;
  wire _abc_15724_n2686;
  wire _abc_15724_n2687_1;
  wire _abc_15724_n2689;
  wire _abc_15724_n2690;
  wire _abc_15724_n2691_1;
  wire _abc_15724_n2692;
  wire _abc_15724_n2693;
  wire _abc_15724_n2694;
  wire _abc_15724_n2695;
  wire _abc_15724_n2696;
  wire _abc_15724_n2697;
  wire _abc_15724_n2698;
  wire _abc_15724_n2699;
  wire _abc_15724_n2700;
  wire _abc_15724_n2701;
  wire _abc_15724_n2702;
  wire _abc_15724_n2703;
  wire _abc_15724_n2705;
  wire _abc_15724_n2706;
  wire _abc_15724_n2707;
  wire _abc_15724_n2708;
  wire _abc_15724_n2709;
  wire _abc_15724_n2710;
  wire _abc_15724_n2711;
  wire _abc_15724_n2712;
  wire _abc_15724_n2713;
  wire _abc_15724_n2714;
  wire _abc_15724_n2715;
  wire _abc_15724_n2716;
  wire _abc_15724_n2718;
  wire _abc_15724_n2719;
  wire _abc_15724_n2720;
  wire _abc_15724_n2721;
  wire _abc_15724_n2722;
  wire _abc_15724_n2723;
  wire _abc_15724_n2724;
  wire _abc_15724_n2725;
  wire _abc_15724_n2726;
  wire _abc_15724_n2727;
  wire _abc_15724_n2728;
  wire _abc_15724_n2729;
  wire _abc_15724_n2730;
  wire _abc_15724_n2731_1;
  wire _abc_15724_n2732;
  wire _abc_15724_n2733;
  wire _abc_15724_n2734_1;
  wire _abc_15724_n2735;
  wire _abc_15724_n2736;
  wire _abc_15724_n2737;
  wire _abc_15724_n2738;
  wire _abc_15724_n2739;
  wire _abc_15724_n2740;
  wire _abc_15724_n2741;
  wire _abc_15724_n2742;
  wire _abc_15724_n2744;
  wire _abc_15724_n2745;
  wire _abc_15724_n2746;
  wire _abc_15724_n2747;
  wire _abc_15724_n2748;
  wire _abc_15724_n2749;
  wire _abc_15724_n2750;
  wire _abc_15724_n2751;
  wire _abc_15724_n2752;
  wire _abc_15724_n2753;
  wire _abc_15724_n2754;
  wire _abc_15724_n2755;
  wire _abc_15724_n2757;
  wire _abc_15724_n2758;
  wire _abc_15724_n2759;
  wire _abc_15724_n2760;
  wire _abc_15724_n2761;
  wire _abc_15724_n2762;
  wire _abc_15724_n2763;
  wire _abc_15724_n2764;
  wire _abc_15724_n2765;
  wire _abc_15724_n2766;
  wire _abc_15724_n2767;
  wire _abc_15724_n2768_1;
  wire _abc_15724_n2769;
  wire _abc_15724_n2771;
  wire _abc_15724_n2772_1;
  wire _abc_15724_n2773;
  wire _abc_15724_n2774;
  wire _abc_15724_n2775;
  wire _abc_15724_n2776;
  wire _abc_15724_n2777;
  wire _abc_15724_n2778;
  wire _abc_15724_n2779;
  wire _abc_15724_n2780;
  wire _abc_15724_n2781;
  wire _abc_15724_n2782;
  wire _abc_15724_n2784;
  wire _abc_15724_n2785;
  wire _abc_15724_n2786;
  wire _abc_15724_n2787;
  wire _abc_15724_n2788;
  wire _abc_15724_n2789;
  wire _abc_15724_n2790;
  wire _abc_15724_n2791;
  wire _abc_15724_n2792;
  wire _abc_15724_n2793;
  wire _abc_15724_n2794;
  wire _abc_15724_n2795;
  wire _abc_15724_n2796;
  wire _abc_15724_n2797;
  wire _abc_15724_n2798;
  wire _abc_15724_n2799;
  wire _abc_15724_n2800;
  wire _abc_15724_n2801;
  wire _abc_15724_n2802;
  wire _abc_15724_n2803;
  wire _abc_15724_n2804;
  wire _abc_15724_n2805;
  wire _abc_15724_n2806;
  wire _abc_15724_n2807;
  wire _abc_15724_n2809;
  wire _abc_15724_n2810;
  wire _abc_15724_n2811;
  wire _abc_15724_n2812_1;
  wire _abc_15724_n2813;
  wire _abc_15724_n2814;
  wire _abc_15724_n2815;
  wire _abc_15724_n2816;
  wire _abc_15724_n2817;
  wire _abc_15724_n2818;
  wire _abc_15724_n2819;
  wire _abc_15724_n2820;
  wire _abc_15724_n2822;
  wire _abc_15724_n2823;
  wire _abc_15724_n2824;
  wire _abc_15724_n2825;
  wire _abc_15724_n2826;
  wire _abc_15724_n2827;
  wire _abc_15724_n2828;
  wire _abc_15724_n2829;
  wire _abc_15724_n2830;
  wire _abc_15724_n2831;
  wire _abc_15724_n2832;
  wire _abc_15724_n2833;
  wire _abc_15724_n2835;
  wire _abc_15724_n2836;
  wire _abc_15724_n2837;
  wire _abc_15724_n2838;
  wire _abc_15724_n2839;
  wire _abc_15724_n2840;
  wire _abc_15724_n2841;
  wire _abc_15724_n2842;
  wire _abc_15724_n2843;
  wire _abc_15724_n2844;
  wire _abc_15724_n2845_1;
  wire _abc_15724_n2846;
  wire _abc_15724_n2848_1;
  wire _abc_15724_n2849;
  wire _abc_15724_n2850;
  wire _abc_15724_n2851;
  wire _abc_15724_n2852;
  wire _abc_15724_n2853;
  wire _abc_15724_n2854;
  wire _abc_15724_n2855;
  wire _abc_15724_n2856;
  wire _abc_15724_n2857;
  wire _abc_15724_n2858;
  wire _abc_15724_n2859;
  wire _abc_15724_n2860;
  wire _abc_15724_n2861;
  wire _abc_15724_n2862;
  wire _abc_15724_n2863;
  wire _abc_15724_n2864;
  wire _abc_15724_n2865;
  wire _abc_15724_n2866;
  wire _abc_15724_n2867;
  wire _abc_15724_n2868;
  wire _abc_15724_n2869;
  wire _abc_15724_n2870;
  wire _abc_15724_n2871;
  wire _abc_15724_n2872;
  wire _abc_15724_n2874;
  wire _abc_15724_n2875;
  wire _abc_15724_n2876;
  wire _abc_15724_n2877;
  wire _abc_15724_n2878;
  wire _abc_15724_n2879;
  wire _abc_15724_n2880;
  wire _abc_15724_n2881;
  wire _abc_15724_n2882;
  wire _abc_15724_n2883;
  wire _abc_15724_n2884;
  wire _abc_15724_n2885;
  wire _abc_15724_n2886;
  wire _abc_15724_n2888;
  wire _abc_15724_n2889;
  wire _abc_15724_n2890_1;
  wire _abc_15724_n2891;
  wire _abc_15724_n2892;
  wire _abc_15724_n2893;
  wire _abc_15724_n2894_1;
  wire _abc_15724_n2895;
  wire _abc_15724_n2896;
  wire _abc_15724_n2897;
  wire _abc_15724_n2898;
  wire _abc_15724_n2899;
  wire _abc_15724_n2900;
  wire _abc_15724_n2901;
  wire _abc_15724_n2902;
  wire _abc_15724_n2903;
  wire _abc_15724_n2905;
  wire _abc_15724_n2906;
  wire _abc_15724_n2907;
  wire _abc_15724_n2908;
  wire _abc_15724_n2909;
  wire _abc_15724_n2910;
  wire _abc_15724_n2911;
  wire _abc_15724_n2912;
  wire _abc_15724_n2913;
  wire _abc_15724_n2914;
  wire _abc_15724_n2915;
  wire _abc_15724_n2916;
  wire _abc_15724_n2918;
  wire _abc_15724_n2919;
  wire _abc_15724_n2920;
  wire _abc_15724_n2921;
  wire _abc_15724_n2922;
  wire _abc_15724_n2923;
  wire _abc_15724_n2924;
  wire _abc_15724_n2925;
  wire _abc_15724_n2926;
  wire _abc_15724_n2927_1;
  wire _abc_15724_n2928;
  wire _abc_15724_n2929;
  wire _abc_15724_n2930_1;
  wire _abc_15724_n2931;
  wire _abc_15724_n2932;
  wire _abc_15724_n2933;
  wire _abc_15724_n2934;
  wire _abc_15724_n2935;
  wire _abc_15724_n2936;
  wire _abc_15724_n2937;
  wire _abc_15724_n2938;
  wire _abc_15724_n2939;
  wire _abc_15724_n2941;
  wire _abc_15724_n2942;
  wire _abc_15724_n2943;
  wire _abc_15724_n2944;
  wire _abc_15724_n2945;
  wire _abc_15724_n2946;
  wire _abc_15724_n2947;
  wire _abc_15724_n2948;
  wire _abc_15724_n2949;
  wire _abc_15724_n2950;
  wire _abc_15724_n2951;
  wire _abc_15724_n2952;
  wire _abc_15724_n2953;
  wire _abc_15724_n2955;
  wire _abc_15724_n2956;
  wire _abc_15724_n2957;
  wire _abc_15724_n2958;
  wire _abc_15724_n2959;
  wire _abc_15724_n2960;
  wire _abc_15724_n2961;
  wire _abc_15724_n2962;
  wire _abc_15724_n2963;
  wire _abc_15724_n2964_1;
  wire _abc_15724_n2965;
  wire _abc_15724_n2966;
  wire _abc_15724_n2967;
  wire _abc_15724_n2968_1;
  wire _abc_15724_n2969;
  wire _abc_15724_n2970;
  wire _abc_15724_n2971;
  wire _abc_15724_n2972;
  wire _abc_15724_n2973;
  wire _abc_15724_n2975;
  wire _abc_15724_n2976;
  wire _abc_15724_n2977;
  wire _abc_15724_n2978;
  wire _abc_15724_n2979;
  wire _abc_15724_n2980;
  wire _abc_15724_n2981;
  wire _abc_15724_n2982;
  wire _abc_15724_n2983;
  wire _abc_15724_n2984;
  wire _abc_15724_n2985;
  wire _abc_15724_n2986;
  wire _abc_15724_n2988;
  wire _abc_15724_n2990;
  wire _abc_15724_n2991;
  wire _abc_15724_n2992;
  wire _abc_15724_n2992_bF_buf0;
  wire _abc_15724_n2992_bF_buf1;
  wire _abc_15724_n2992_bF_buf10;
  wire _abc_15724_n2992_bF_buf11;
  wire _abc_15724_n2992_bF_buf2;
  wire _abc_15724_n2992_bF_buf3;
  wire _abc_15724_n2992_bF_buf4;
  wire _abc_15724_n2992_bF_buf5;
  wire _abc_15724_n2992_bF_buf6;
  wire _abc_15724_n2992_bF_buf7;
  wire _abc_15724_n2992_bF_buf8;
  wire _abc_15724_n2992_bF_buf9;
  wire _abc_15724_n2993;
  wire _abc_15724_n2994;
  wire _abc_15724_n2994_bF_buf0;
  wire _abc_15724_n2994_bF_buf1;
  wire _abc_15724_n2994_bF_buf10;
  wire _abc_15724_n2994_bF_buf11;
  wire _abc_15724_n2994_bF_buf2;
  wire _abc_15724_n2994_bF_buf3;
  wire _abc_15724_n2994_bF_buf4;
  wire _abc_15724_n2994_bF_buf5;
  wire _abc_15724_n2994_bF_buf6;
  wire _abc_15724_n2994_bF_buf7;
  wire _abc_15724_n2994_bF_buf8;
  wire _abc_15724_n2994_bF_buf9;
  wire _abc_15724_n2995;
  wire _abc_15724_n2996;
  wire _abc_15724_n2997;
  wire _abc_15724_n2998;
  wire _abc_15724_n3000;
  wire _abc_15724_n3001;
  wire _abc_15724_n3002;
  wire _abc_15724_n3003_1;
  wire _abc_15724_n3004;
  wire _abc_15724_n3006;
  wire _abc_15724_n3007;
  wire _abc_15724_n3008;
  wire _abc_15724_n3009;
  wire _abc_15724_n3010;
  wire _abc_15724_n3012;
  wire _abc_15724_n3013;
  wire _abc_15724_n3014;
  wire _abc_15724_n3015;
  wire _abc_15724_n3016;
  wire _abc_15724_n3018;
  wire _abc_15724_n3019;
  wire _abc_15724_n3020;
  wire _abc_15724_n3021;
  wire _abc_15724_n3022;
  wire _abc_15724_n3024;
  wire _abc_15724_n3025;
  wire _abc_15724_n3026;
  wire _abc_15724_n3027;
  wire _abc_15724_n3028;
  wire _abc_15724_n3030;
  wire _abc_15724_n3031;
  wire _abc_15724_n3032;
  wire _abc_15724_n3033;
  wire _abc_15724_n3034;
  wire _abc_15724_n3036;
  wire _abc_15724_n3037;
  wire _abc_15724_n3038;
  wire _abc_15724_n3039;
  wire _abc_15724_n3040_1;
  wire _abc_15724_n3042;
  wire _abc_15724_n3043;
  wire _abc_15724_n3044_1;
  wire _abc_15724_n3045;
  wire _abc_15724_n3046;
  wire _abc_15724_n3048;
  wire _abc_15724_n3049;
  wire _abc_15724_n3050;
  wire _abc_15724_n3051;
  wire _abc_15724_n3052;
  wire _abc_15724_n3054;
  wire _abc_15724_n3055;
  wire _abc_15724_n3056;
  wire _abc_15724_n3057;
  wire _abc_15724_n3058;
  wire _abc_15724_n3060;
  wire _abc_15724_n3061;
  wire _abc_15724_n3062;
  wire _abc_15724_n3063;
  wire _abc_15724_n3064;
  wire _abc_15724_n3066;
  wire _abc_15724_n3067;
  wire _abc_15724_n3068;
  wire _abc_15724_n3069;
  wire _abc_15724_n3070;
  wire _abc_15724_n3072;
  wire _abc_15724_n3073;
  wire _abc_15724_n3074;
  wire _abc_15724_n3075;
  wire _abc_15724_n3076_1;
  wire _abc_15724_n3078;
  wire _abc_15724_n3079_1;
  wire _abc_15724_n3080;
  wire _abc_15724_n3081;
  wire _abc_15724_n3082;
  wire _abc_15724_n3084;
  wire _abc_15724_n3085;
  wire _abc_15724_n3086;
  wire _abc_15724_n3087;
  wire _abc_15724_n3088;
  wire _abc_15724_n3090;
  wire _abc_15724_n3091;
  wire _abc_15724_n3092;
  wire _abc_15724_n3093;
  wire _abc_15724_n3094;
  wire _abc_15724_n3096;
  wire _abc_15724_n3097;
  wire _abc_15724_n3098;
  wire _abc_15724_n3099;
  wire _abc_15724_n3100;
  wire _abc_15724_n3102;
  wire _abc_15724_n3103;
  wire _abc_15724_n3104;
  wire _abc_15724_n3105;
  wire _abc_15724_n3106;
  wire _abc_15724_n3108;
  wire _abc_15724_n3109;
  wire _abc_15724_n3110;
  wire _abc_15724_n3111;
  wire _abc_15724_n3112;
  wire _abc_15724_n3114_1;
  wire _abc_15724_n3115;
  wire _abc_15724_n3116;
  wire _abc_15724_n3117;
  wire _abc_15724_n3118_1;
  wire _abc_15724_n3120;
  wire _abc_15724_n3121;
  wire _abc_15724_n3122;
  wire _abc_15724_n3123;
  wire _abc_15724_n3124;
  wire _abc_15724_n3126;
  wire _abc_15724_n3127;
  wire _abc_15724_n3128;
  wire _abc_15724_n3129;
  wire _abc_15724_n3131;
  wire _abc_15724_n3132;
  wire _abc_15724_n3133;
  wire _abc_15724_n3134;
  wire _abc_15724_n3136;
  wire _abc_15724_n3137;
  wire _abc_15724_n3138;
  wire _abc_15724_n3139;
  wire _abc_15724_n3141;
  wire _abc_15724_n3142;
  wire _abc_15724_n3143;
  wire _abc_15724_n3144;
  wire _abc_15724_n3146;
  wire _abc_15724_n3147;
  wire _abc_15724_n3148;
  wire _abc_15724_n3149;
  wire _abc_15724_n3150_1;
  wire _abc_15724_n3152;
  wire _abc_15724_n3153_1;
  wire _abc_15724_n3154;
  wire _abc_15724_n3155;
  wire _abc_15724_n3156;
  wire _abc_15724_n3158;
  wire _abc_15724_n3159;
  wire _abc_15724_n3160;
  wire _abc_15724_n3161;
  wire _abc_15724_n3162;
  wire _abc_15724_n3164;
  wire _abc_15724_n3165;
  wire _abc_15724_n3166;
  wire _abc_15724_n3167;
  wire _abc_15724_n3169;
  wire _abc_15724_n3170;
  wire _abc_15724_n3171;
  wire _abc_15724_n3172;
  wire _abc_15724_n3174;
  wire _abc_15724_n3175;
  wire _abc_15724_n3176;
  wire _abc_15724_n3177;
  wire _abc_15724_n3179;
  wire _abc_15724_n3180;
  wire _abc_15724_n3181;
  wire _abc_15724_n3182;
  wire _abc_15724_n3184;
  wire _abc_15724_n3185;
  wire _abc_15724_n3186;
  wire _abc_15724_n3187;
  wire _abc_15724_n3189;
  wire _abc_15724_n3190;
  wire _abc_15724_n3191;
  wire _abc_15724_n3192;
  wire _abc_15724_n3194;
  wire _abc_15724_n3195_1;
  wire _abc_15724_n3196;
  wire _abc_15724_n3197;
  wire _abc_15724_n3198_1;
  wire _abc_15724_n3200;
  wire _abc_15724_n3201;
  wire _abc_15724_n3202;
  wire _abc_15724_n3203;
  wire _abc_15724_n3205;
  wire _abc_15724_n3206;
  wire _abc_15724_n3207;
  wire _abc_15724_n3208;
  wire _abc_15724_n3210;
  wire _abc_15724_n3211;
  wire _abc_15724_n3212;
  wire _abc_15724_n3213;
  wire _abc_15724_n3215;
  wire _abc_15724_n3216;
  wire _abc_15724_n3217;
  wire _abc_15724_n3218;
  wire _abc_15724_n3219;
  wire _abc_15724_n3221;
  wire _abc_15724_n3222;
  wire _abc_15724_n3223;
  wire _abc_15724_n3224;
  wire _abc_15724_n3225;
  wire _abc_15724_n3227;
  wire _abc_15724_n3228;
  wire _abc_15724_n3229;
  wire _abc_15724_n3230_1;
  wire _abc_15724_n3231;
  wire _abc_15724_n3233_1;
  wire _abc_15724_n3234;
  wire _abc_15724_n3235;
  wire _abc_15724_n3236;
  wire _abc_15724_n3238;
  wire _abc_15724_n3239;
  wire _abc_15724_n3240;
  wire _abc_15724_n3241;
  wire _abc_15724_n3242;
  wire _abc_15724_n3244;
  wire _abc_15724_n3245;
  wire _abc_15724_n3246;
  wire _abc_15724_n3247;
  wire _abc_15724_n3249;
  wire _abc_15724_n3250;
  wire _abc_15724_n3251;
  wire _abc_15724_n3252;
  wire _abc_15724_n3253;
  wire _abc_15724_n3255;
  wire _abc_15724_n3256;
  wire _abc_15724_n3257;
  wire _abc_15724_n3258;
  wire _abc_15724_n3260;
  wire _abc_15724_n3261;
  wire _abc_15724_n3262;
  wire _abc_15724_n3263;
  wire _abc_15724_n3264;
  wire _abc_15724_n3266;
  wire _abc_15724_n3267;
  wire _abc_15724_n3268;
  wire _abc_15724_n3269;
  wire _abc_15724_n3270_1;
  wire _abc_15724_n3272;
  wire _abc_15724_n3273;
  wire _abc_15724_n3274_1;
  wire _abc_15724_n3275;
  wire _abc_15724_n3277;
  wire _abc_15724_n3278;
  wire _abc_15724_n3279;
  wire _abc_15724_n3280;
  wire _abc_15724_n3281;
  wire _abc_15724_n3283;
  wire _abc_15724_n3284;
  wire _abc_15724_n3285;
  wire _abc_15724_n3286;
  wire _abc_15724_n3287;
  wire _abc_15724_n3289;
  wire _abc_15724_n3290;
  wire _abc_15724_n3291;
  wire _abc_15724_n3292;
  wire _abc_15724_n3294;
  wire _abc_15724_n3295;
  wire _abc_15724_n3296;
  wire _abc_15724_n3297;
  wire _abc_15724_n3299;
  wire _abc_15724_n3300;
  wire _abc_15724_n3301;
  wire _abc_15724_n3302;
  wire _abc_15724_n3303;
  wire _abc_15724_n3305;
  wire _abc_15724_n3306;
  wire _abc_15724_n3307_1;
  wire _abc_15724_n3308;
  wire _abc_15724_n3309;
  wire _abc_15724_n3311_1;
  wire _abc_15724_n3312;
  wire _abc_15724_n3313;
  wire _abc_15724_n3314;
  wire _abc_15724_n3315;
  wire _abc_15724_n3317;
  wire _abc_15724_n3318;
  wire _abc_15724_n3319;
  wire _abc_15724_n3320;
  wire _abc_15724_n3321;
  wire _abc_15724_n3323;
  wire _abc_15724_n3324;
  wire _abc_15724_n3325;
  wire _abc_15724_n3326;
  wire _abc_15724_n3327;
  wire _abc_15724_n3329;
  wire _abc_15724_n3330;
  wire _abc_15724_n3331;
  wire _abc_15724_n3332;
  wire _abc_15724_n3333;
  wire _abc_15724_n3335;
  wire _abc_15724_n3336;
  wire _abc_15724_n3337;
  wire _abc_15724_n3338;
  wire _abc_15724_n3340;
  wire _abc_15724_n3341;
  wire _abc_15724_n3342;
  wire _abc_15724_n3343;
  wire _abc_15724_n3345;
  wire _abc_15724_n3346;
  wire _abc_15724_n3347;
  wire _abc_15724_n3348;
  wire _abc_15724_n3349_1;
  wire _abc_15724_n3351;
  wire _abc_15724_n3352_1;
  wire _abc_15724_n3353;
  wire _abc_15724_n3354;
  wire _abc_15724_n3355;
  wire _abc_15724_n3357;
  wire _abc_15724_n3358;
  wire _abc_15724_n3359;
  wire _abc_15724_n3360;
  wire _abc_15724_n3362;
  wire _abc_15724_n3363;
  wire _abc_15724_n3364;
  wire _abc_15724_n3365;
  wire _abc_15724_n3367;
  wire _abc_15724_n3368;
  wire _abc_15724_n3369;
  wire _abc_15724_n3370;
  wire _abc_15724_n3372;
  wire _abc_15724_n3373;
  wire _abc_15724_n3374;
  wire _abc_15724_n3375;
  wire _abc_15724_n3377;
  wire _abc_15724_n3378;
  wire _abc_15724_n3379;
  wire _abc_15724_n3380;
  wire _abc_15724_n3382;
  wire _abc_15724_n3383;
  wire _abc_15724_n3384;
  wire _abc_15724_n3385;
  wire _abc_15724_n3387;
  wire _abc_15724_n3388;
  wire _abc_15724_n3389_1;
  wire _abc_15724_n3390;
  wire _abc_15724_n3392;
  wire _abc_15724_n3393;
  wire _abc_15724_n3394;
  wire _abc_15724_n3395;
  wire _abc_15724_n3397;
  wire _abc_15724_n3398;
  wire _abc_15724_n3399;
  wire _abc_15724_n3400;
  wire _abc_15724_n3401;
  wire _abc_15724_n3403;
  wire _abc_15724_n3404;
  wire _abc_15724_n3405;
  wire _abc_15724_n3406;
  wire _abc_15724_n3407;
  wire _abc_15724_n3409;
  wire _abc_15724_n3410;
  wire _abc_15724_n3411;
  wire _abc_15724_n3412;
  wire _abc_15724_n3414;
  wire _abc_15724_n3415;
  wire _abc_15724_n3416;
  wire _abc_15724_n3417;
  wire _abc_15724_n3419;
  wire _abc_15724_n3420;
  wire _abc_15724_n3421;
  wire _abc_15724_n3422;
  wire _abc_15724_n3424;
  wire _abc_15724_n3425_1;
  wire _abc_15724_n3426;
  wire _abc_15724_n3427;
  wire _abc_15724_n3428;
  wire _abc_15724_n3430;
  wire _abc_15724_n3431;
  wire _abc_15724_n3432;
  wire _abc_15724_n3433;
  wire _abc_15724_n3435;
  wire _abc_15724_n3436;
  wire _abc_15724_n3437;
  wire _abc_15724_n3438;
  wire _abc_15724_n3440;
  wire _abc_15724_n3441;
  wire _abc_15724_n3442;
  wire _abc_15724_n3443;
  wire _abc_15724_n3444;
  wire _abc_15724_n3446;
  wire _abc_15724_n3447;
  wire _abc_15724_n3448;
  wire _abc_15724_n3449;
  wire _abc_15724_n3451;
  wire _abc_15724_n3452;
  wire _abc_15724_n3453;
  wire _abc_15724_n3454;
  wire _abc_15724_n3455;
  wire _abc_15724_n3457;
  wire _abc_15724_n3458;
  wire _abc_15724_n3459;
  wire _abc_15724_n3460;
  wire _abc_15724_n3462;
  wire _abc_15724_n3463;
  wire _abc_15724_n3464;
  wire _abc_15724_n3465;
  wire _abc_15724_n3465_1;
  wire _abc_15724_n3467;
  wire _abc_15724_n3468_1;
  wire _abc_15724_n3469_1;
  wire _abc_15724_n3470;
  wire _abc_15724_n3472;
  wire _abc_15724_n3473;
  wire _abc_15724_n3474;
  wire _abc_15724_n3475;
  wire _abc_15724_n3476;
  wire _abc_15724_n3478;
  wire _abc_15724_n3479;
  wire _abc_15724_n3480;
  wire _abc_15724_n3481;
  wire _abc_15724_n3483;
  wire _abc_15724_n3483_1;
  wire _abc_15724_n3484;
  wire _abc_15724_n3485;
  wire _abc_15724_n3486;
  wire _abc_15724_n3487;
  wire _abc_15724_n3489;
  wire _abc_15724_n3489_1;
  wire _abc_15724_n3490;
  wire _abc_15724_n3491_1;
  wire _abc_15724_n3492_1;
  wire _abc_15724_n3493;
  wire _abc_15724_n3495;
  wire _abc_15724_n3496;
  wire _abc_15724_n3497_1;
  wire _abc_15724_n3498;
  wire _abc_15724_n3499;
  wire _abc_15724_n3501_1;
  wire _abc_15724_n3502;
  wire _abc_15724_n3503;
  wire _abc_15724_n3504;
  wire _abc_15724_n3506;
  wire _abc_15724_n3507_1;
  wire _abc_15724_n3508;
  wire _abc_15724_n3509;
  wire _abc_15724_n3511;
  wire _abc_15724_n3512;
  wire _abc_15724_n3513_1;
  wire _abc_15724_n3514_1;
  wire _abc_15724_n3515;
  wire _abc_15724_n3517_1;
  wire _abc_15724_n3518;
  wire _abc_15724_n3519;
  wire _abc_15724_n3520;
  wire _abc_15724_n3521_1;
  wire _abc_15724_n3523;
  wire _abc_15724_n3524;
  wire _abc_15724_n3525;
  wire _abc_15724_n3526;
  wire _abc_15724_n3528_1;
  wire _abc_15724_n3529_1;
  wire _abc_15724_n3530;
  wire _abc_15724_n3531;
  wire _abc_15724_n3533;
  wire _abc_15724_n3534;
  wire _abc_15724_n3535_1;
  wire _abc_15724_n3536;
  wire _abc_15724_n3537;
  wire _abc_15724_n3539;
  wire _abc_15724_n3540;
  wire _abc_15724_n3541;
  wire _abc_15724_n3542;
  wire _abc_15724_n3543;
  wire _abc_15724_n3545;
  wire _abc_15724_n3546_1;
  wire _abc_15724_n3547;
  wire _abc_15724_n3548;
  wire _abc_15724_n3550;
  wire _abc_15724_n3551;
  wire _abc_15724_n3552;
  wire _abc_15724_n3553;
  wire _abc_15724_n3554_1;
  wire _abc_15724_n3556;
  wire _abc_15724_n3557;
  wire _abc_15724_n3558;
  wire _abc_15724_n3559;
  wire _abc_15724_n3560;
  wire _abc_15724_n3562;
  wire _abc_15724_n3563;
  wire _abc_15724_n3564_1;
  wire _abc_15724_n3565;
  wire _abc_15724_n3566;
  wire _abc_15724_n3568;
  wire _abc_15724_n3569;
  wire _abc_15724_n3570;
  wire _abc_15724_n3571;
  wire _abc_15724_n3573;
  wire _abc_15724_n3574;
  wire _abc_15724_n3575;
  wire _abc_15724_n3576;
  wire _abc_15724_n3578;
  wire _abc_15724_n3579;
  wire _abc_15724_n3580;
  wire _abc_15724_n3581;
  wire _abc_15724_n3583;
  wire _abc_15724_n3584_1;
  wire _abc_15724_n3585_1;
  wire _abc_15724_n3586;
  wire _abc_15724_n3587;
  wire _abc_15724_n3589;
  wire _abc_15724_n3590;
  wire _abc_15724_n3591_1;
  wire _abc_15724_n3592_1;
  wire _abc_15724_n3594;
  wire _abc_15724_n3595;
  wire _abc_15724_n3596;
  wire _abc_15724_n3597;
  wire _abc_15724_n3598;
  wire _abc_15724_n3600;
  wire _abc_15724_n3601;
  wire _abc_15724_n3602_1;
  wire _abc_15724_n3603_1;
  wire _abc_15724_n3605;
  wire _abc_15724_n3606;
  wire _abc_15724_n3607;
  wire _abc_15724_n3608;
  wire _abc_15724_n3609_1;
  wire _abc_15724_n3611;
  wire _abc_15724_n3612;
  wire _abc_15724_n3613;
  wire _abc_15724_n3614;
  wire _abc_15724_n3616;
  wire _abc_15724_n3617;
  wire _abc_15724_n3618;
  wire _abc_15724_n3619;
  wire _abc_15724_n3621_1;
  wire _abc_15724_n3622;
  wire _abc_15724_n3623;
  wire _abc_15724_n3624;
  wire _abc_15724_n3625;
  wire _abc_15724_n3627;
  wire _abc_15724_n3628;
  wire _abc_15724_n3629_1;
  wire _abc_15724_n3630;
  wire _abc_15724_n3632;
  wire _abc_15724_n3633;
  wire _abc_15724_n3634;
  wire _abc_15724_n3635;
  wire _abc_15724_n3637;
  wire _abc_15724_n3638;
  wire _abc_15724_n3639_1;
  wire _abc_15724_n3640;
  wire _abc_15724_n3641;
  wire _abc_15724_n3643;
  wire _abc_15724_n3644;
  wire _abc_15724_n3645_1;
  wire _abc_15724_n3646_1;
  wire _abc_15724_n3647;
  wire _abc_15724_n3649;
  wire _abc_15724_n3650;
  wire _abc_15724_n3651;
  wire _abc_15724_n3652;
  wire _abc_15724_n3654;
  wire _abc_15724_n3655;
  wire _abc_15724_n3656;
  wire _abc_15724_n3657;
  wire _abc_15724_n3659;
  wire _abc_15724_n3660;
  wire _abc_15724_n3661;
  wire _abc_15724_n3662_1;
  wire _abc_15724_n3664;
  wire _abc_15724_n3665;
  wire _abc_15724_n3666;
  wire _abc_15724_n3667;
  wire _abc_15724_n3669;
  wire _abc_15724_n3670_1;
  wire _abc_15724_n3671_1;
  wire _abc_15724_n3672;
  wire _abc_15724_n3674;
  wire _abc_15724_n3675;
  wire _abc_15724_n3676;
  wire _abc_15724_n3677;
  wire _abc_15724_n3679_1;
  wire _abc_15724_n3680_1;
  wire _abc_15724_n3681;
  wire _abc_15724_n3682;
  wire _abc_15724_n3683;
  wire _abc_15724_n3685;
  wire _abc_15724_n3686_1;
  wire _abc_15724_n3687;
  wire _abc_15724_n3688;
  wire _abc_15724_n3690;
  wire _abc_15724_n3691;
  wire _abc_15724_n3692;
  wire _abc_15724_n3693;
  wire _abc_15724_n3695;
  wire _abc_15724_n3696;
  wire _abc_15724_n3697;
  wire _abc_15724_n3698_1;
  wire _abc_15724_n3700;
  wire _abc_15724_n3701;
  wire _abc_15724_n3702;
  wire _abc_15724_n3703;
  wire _abc_15724_n3704;
  wire _abc_15724_n3705;
  wire _abc_15724_n3706;
  wire _abc_15724_n3707;
  wire _abc_15724_n3708;
  wire _abc_15724_n3709;
  wire _abc_15724_n3710;
  wire _abc_15724_n3711;
  wire _abc_15724_n3712;
  wire _abc_15724_n3713;
  wire _abc_15724_n3714;
  wire _abc_15724_n3715;
  wire _abc_15724_n3716;
  wire _abc_15724_n3717;
  wire _abc_15724_n3718;
  wire _abc_15724_n3719;
  wire _abc_15724_n3720;
  wire _abc_15724_n3721;
  wire _abc_15724_n3721_bF_buf0;
  wire _abc_15724_n3721_bF_buf1;
  wire _abc_15724_n3721_bF_buf2;
  wire _abc_15724_n3721_bF_buf3;
  wire _abc_15724_n3721_bF_buf4;
  wire _abc_15724_n3722;
  wire _abc_15724_n3723;
  wire _abc_15724_n3724;
  wire _abc_15724_n3725;
  wire _abc_15724_n3725_bF_buf0;
  wire _abc_15724_n3725_bF_buf1;
  wire _abc_15724_n3725_bF_buf2;
  wire _abc_15724_n3725_bF_buf3;
  wire _abc_15724_n3726;
  wire _abc_15724_n3726_bF_buf0;
  wire _abc_15724_n3726_bF_buf1;
  wire _abc_15724_n3726_bF_buf2;
  wire _abc_15724_n3726_bF_buf3;
  wire _abc_15724_n3726_bF_buf4;
  wire _abc_15724_n3727;
  wire _abc_15724_n3728;
  wire _abc_15724_n3729;
  wire _abc_15724_n3730;
  wire _abc_15724_n3731;
  wire _abc_15724_n3732;
  wire _abc_15724_n3733;
  wire _abc_15724_n3734;
  wire _abc_15724_n3735;
  wire _abc_15724_n3736;
  wire _abc_15724_n3737;
  wire _abc_15724_n3737_bF_buf0;
  wire _abc_15724_n3737_bF_buf1;
  wire _abc_15724_n3737_bF_buf2;
  wire _abc_15724_n3737_bF_buf3;
  wire _abc_15724_n3737_bF_buf4;
  wire _abc_15724_n3738;
  wire _abc_15724_n3739;
  wire _abc_15724_n3740;
  wire _abc_15724_n3741;
  wire _abc_15724_n3742;
  wire _abc_15724_n3743;
  wire _abc_15724_n3744;
  wire _abc_15724_n3745;
  wire _abc_15724_n3746;
  wire _abc_15724_n3747;
  wire _abc_15724_n3748;
  wire _abc_15724_n3749;
  wire _abc_15724_n3750;
  wire _abc_15724_n3751;
  wire _abc_15724_n3752;
  wire _abc_15724_n3753;
  wire _abc_15724_n3754;
  wire _abc_15724_n3755;
  wire _abc_15724_n3756;
  wire _abc_15724_n3757;
  wire _abc_15724_n3758;
  wire _abc_15724_n3759;
  wire _abc_15724_n3760;
  wire _abc_15724_n3761;
  wire _abc_15724_n3762;
  wire _abc_15724_n3763;
  wire _abc_15724_n3764;
  wire _abc_15724_n3765;
  wire _abc_15724_n3766;
  wire _abc_15724_n3767;
  wire _abc_15724_n3769;
  wire _abc_15724_n3770;
  wire _abc_15724_n3771;
  wire _abc_15724_n3772;
  wire _abc_15724_n3773;
  wire _abc_15724_n3774;
  wire _abc_15724_n3775;
  wire _abc_15724_n3776;
  wire _abc_15724_n3777;
  wire _abc_15724_n3778;
  wire _abc_15724_n3779;
  wire _abc_15724_n3780;
  wire _abc_15724_n3781;
  wire _abc_15724_n3782;
  wire _abc_15724_n3783;
  wire _abc_15724_n3784;
  wire _abc_15724_n3785;
  wire _abc_15724_n3786;
  wire _abc_15724_n3787;
  wire _abc_15724_n3788;
  wire _abc_15724_n3789;
  wire _abc_15724_n3790;
  wire _abc_15724_n3791;
  wire _abc_15724_n3792;
  wire _abc_15724_n3793;
  wire _abc_15724_n3794;
  wire _abc_15724_n3795;
  wire _abc_15724_n3796;
  wire _abc_15724_n3797;
  wire _abc_15724_n3798;
  wire _abc_15724_n3799;
  wire _abc_15724_n3800;
  wire _abc_15724_n3801;
  wire _abc_15724_n3802;
  wire _abc_15724_n3803;
  wire _abc_15724_n3804;
  wire _abc_15724_n3805;
  wire _abc_15724_n3805_bF_buf0;
  wire _abc_15724_n3805_bF_buf1;
  wire _abc_15724_n3805_bF_buf2;
  wire _abc_15724_n3805_bF_buf3;
  wire _abc_15724_n3805_bF_buf4;
  wire _abc_15724_n3806;
  wire _abc_15724_n3806_bF_buf0;
  wire _abc_15724_n3806_bF_buf1;
  wire _abc_15724_n3806_bF_buf2;
  wire _abc_15724_n3806_bF_buf3;
  wire _abc_15724_n3807;
  wire _abc_15724_n3808;
  wire _abc_15724_n3809;
  wire _abc_15724_n3810;
  wire _abc_15724_n3811;
  wire _abc_15724_n3812;
  wire _abc_15724_n3813;
  wire _abc_15724_n3814;
  wire _abc_15724_n3815;
  wire _abc_15724_n3816;
  wire _abc_15724_n3817;
  wire _abc_15724_n3818;
  wire _abc_15724_n3819;
  wire _abc_15724_n3820;
  wire _abc_15724_n3821;
  wire _abc_15724_n3822;
  wire _abc_15724_n3823;
  wire _abc_15724_n3824;
  wire _abc_15724_n3825;
  wire _abc_15724_n3826;
  wire _abc_15724_n3827;
  wire _abc_15724_n3828;
  wire _abc_15724_n3829;
  wire _abc_15724_n3830;
  wire _abc_15724_n3831;
  wire _abc_15724_n3832;
  wire _abc_15724_n3833;
  wire _abc_15724_n3834;
  wire _abc_15724_n3835;
  wire _abc_15724_n3836;
  wire _abc_15724_n3837;
  wire _abc_15724_n3838;
  wire _abc_15724_n3839;
  wire _abc_15724_n3840;
  wire _abc_15724_n3841;
  wire _abc_15724_n3843;
  wire _abc_15724_n3844;
  wire _abc_15724_n3845;
  wire _abc_15724_n3846;
  wire _abc_15724_n3847;
  wire _abc_15724_n3848;
  wire _abc_15724_n3849;
  wire _abc_15724_n3850;
  wire _abc_15724_n3851;
  wire _abc_15724_n3852;
  wire _abc_15724_n3853;
  wire _abc_15724_n3854;
  wire _abc_15724_n3855;
  wire _abc_15724_n3856;
  wire _abc_15724_n3857;
  wire _abc_15724_n3858;
  wire _abc_15724_n3859;
  wire _abc_15724_n3860;
  wire _abc_15724_n3861;
  wire _abc_15724_n3862;
  wire _abc_15724_n3863;
  wire _abc_15724_n3864;
  wire _abc_15724_n3865;
  wire _abc_15724_n3866;
  wire _abc_15724_n3867;
  wire _abc_15724_n3868;
  wire _abc_15724_n3869;
  wire _abc_15724_n3870;
  wire _abc_15724_n3871;
  wire _abc_15724_n3872;
  wire _abc_15724_n3873;
  wire _abc_15724_n3874;
  wire _abc_15724_n3875;
  wire _abc_15724_n3876;
  wire _abc_15724_n3877;
  wire _abc_15724_n3878;
  wire _abc_15724_n3879;
  wire _abc_15724_n3880;
  wire _abc_15724_n3881;
  wire _abc_15724_n3882;
  wire _abc_15724_n3883;
  wire _abc_15724_n3884;
  wire _abc_15724_n3885;
  wire _abc_15724_n3886;
  wire _abc_15724_n3887;
  wire _abc_15724_n3888;
  wire _abc_15724_n3889;
  wire _abc_15724_n3890;
  wire _abc_15724_n3891;
  wire _abc_15724_n3892;
  wire _abc_15724_n3893;
  wire _abc_15724_n3894;
  wire _abc_15724_n3895;
  wire _abc_15724_n3896;
  wire _abc_15724_n3897;
  wire _abc_15724_n3898;
  wire _abc_15724_n3899;
  wire _abc_15724_n3900;
  wire _abc_15724_n3901;
  wire _abc_15724_n3902;
  wire _abc_15724_n3903;
  wire _abc_15724_n3904;
  wire _abc_15724_n3905;
  wire _abc_15724_n3906;
  wire _abc_15724_n3907;
  wire _abc_15724_n3908;
  wire _abc_15724_n3909;
  wire _abc_15724_n3910;
  wire _abc_15724_n3911;
  wire _abc_15724_n3912;
  wire _abc_15724_n3913;
  wire _abc_15724_n3914;
  wire _abc_15724_n3915;
  wire _abc_15724_n3916;
  wire _abc_15724_n3917;
  wire _abc_15724_n3918;
  wire _abc_15724_n3919;
  wire _abc_15724_n3920;
  wire _abc_15724_n3921;
  wire _abc_15724_n3922;
  wire _abc_15724_n3923;
  wire _abc_15724_n3924;
  wire _abc_15724_n3925;
  wire _abc_15724_n3926;
  wire _abc_15724_n3928;
  wire _abc_15724_n3929;
  wire _abc_15724_n3930;
  wire _abc_15724_n3931;
  wire _abc_15724_n3932;
  wire _abc_15724_n3933;
  wire _abc_15724_n3934;
  wire _abc_15724_n3935;
  wire _abc_15724_n3936;
  wire _abc_15724_n3937;
  wire _abc_15724_n3938;
  wire _abc_15724_n3939;
  wire _abc_15724_n3940;
  wire _abc_15724_n3941;
  wire _abc_15724_n3942;
  wire _abc_15724_n3943;
  wire _abc_15724_n3944;
  wire _abc_15724_n3945;
  wire _abc_15724_n3946;
  wire _abc_15724_n3947;
  wire _abc_15724_n3948;
  wire _abc_15724_n3949;
  wire _abc_15724_n3950;
  wire _abc_15724_n3951;
  wire _abc_15724_n3952;
  wire _abc_15724_n3953;
  wire _abc_15724_n3954;
  wire _abc_15724_n3955;
  wire _abc_15724_n3956;
  wire _abc_15724_n3957;
  wire _abc_15724_n3958;
  wire _abc_15724_n3959;
  wire _abc_15724_n3960;
  wire _abc_15724_n3961;
  wire _abc_15724_n3962;
  wire _abc_15724_n3963;
  wire _abc_15724_n3964;
  wire _abc_15724_n3965;
  wire _abc_15724_n3966;
  wire _abc_15724_n3967;
  wire _abc_15724_n3968;
  wire _abc_15724_n3969;
  wire _abc_15724_n3970;
  wire _abc_15724_n3971;
  wire _abc_15724_n3972;
  wire _abc_15724_n3973;
  wire _abc_15724_n3974;
  wire _abc_15724_n3975;
  wire _abc_15724_n3976;
  wire _abc_15724_n3977;
  wire _abc_15724_n3978;
  wire _abc_15724_n3979;
  wire _abc_15724_n3980;
  wire _abc_15724_n3981;
  wire _abc_15724_n3982;
  wire _abc_15724_n3983;
  wire _abc_15724_n3984;
  wire _abc_15724_n3985;
  wire _abc_15724_n3986;
  wire _abc_15724_n3987;
  wire _abc_15724_n3988;
  wire _abc_15724_n3989;
  wire _abc_15724_n3990;
  wire _abc_15724_n3991;
  wire _abc_15724_n3992;
  wire _abc_15724_n3993;
  wire _abc_15724_n3994;
  wire _abc_15724_n3995;
  wire _abc_15724_n3996;
  wire _abc_15724_n3997;
  wire _abc_15724_n3998;
  wire _abc_15724_n3999;
  wire _abc_15724_n4000;
  wire _abc_15724_n4001;
  wire _abc_15724_n4002;
  wire _abc_15724_n4003;
  wire _abc_15724_n4004;
  wire _abc_15724_n4005;
  wire _abc_15724_n4006;
  wire _abc_15724_n4007;
  wire _abc_15724_n4008;
  wire _abc_15724_n4009;
  wire _abc_15724_n4010;
  wire _abc_15724_n4011;
  wire _abc_15724_n4012;
  wire _abc_15724_n4013;
  wire _abc_15724_n4014;
  wire _abc_15724_n4016;
  wire _abc_15724_n4017;
  wire _abc_15724_n4018;
  wire _abc_15724_n4019;
  wire _abc_15724_n4020;
  wire _abc_15724_n4021;
  wire _abc_15724_n4022;
  wire _abc_15724_n4023;
  wire _abc_15724_n4024;
  wire _abc_15724_n4025;
  wire _abc_15724_n4026;
  wire _abc_15724_n4027;
  wire _abc_15724_n4028;
  wire _abc_15724_n4029;
  wire _abc_15724_n4030;
  wire _abc_15724_n4031;
  wire _abc_15724_n4032;
  wire _abc_15724_n4033;
  wire _abc_15724_n4034;
  wire _abc_15724_n4035;
  wire _abc_15724_n4036;
  wire _abc_15724_n4037;
  wire _abc_15724_n4038;
  wire _abc_15724_n4039;
  wire _abc_15724_n4040;
  wire _abc_15724_n4041;
  wire _abc_15724_n4042;
  wire _abc_15724_n4043;
  wire _abc_15724_n4044;
  wire _abc_15724_n4045;
  wire _abc_15724_n4046;
  wire _abc_15724_n4047;
  wire _abc_15724_n4048;
  wire _abc_15724_n4049;
  wire _abc_15724_n4050;
  wire _abc_15724_n4051;
  wire _abc_15724_n4052;
  wire _abc_15724_n4053;
  wire _abc_15724_n4054;
  wire _abc_15724_n4055;
  wire _abc_15724_n4056;
  wire _abc_15724_n4057;
  wire _abc_15724_n4058;
  wire _abc_15724_n4059;
  wire _abc_15724_n4060;
  wire _abc_15724_n4061;
  wire _abc_15724_n4062;
  wire _abc_15724_n4063;
  wire _abc_15724_n4064;
  wire _abc_15724_n4065;
  wire _abc_15724_n4066;
  wire _abc_15724_n4067;
  wire _abc_15724_n4068;
  wire _abc_15724_n4069;
  wire _abc_15724_n4070;
  wire _abc_15724_n4071;
  wire _abc_15724_n4072;
  wire _abc_15724_n4073;
  wire _abc_15724_n4074;
  wire _abc_15724_n4075;
  wire _abc_15724_n4076;
  wire _abc_15724_n4077;
  wire _abc_15724_n4078;
  wire _abc_15724_n4079;
  wire _abc_15724_n4080;
  wire _abc_15724_n4081;
  wire _abc_15724_n4082;
  wire _abc_15724_n4083;
  wire _abc_15724_n4084;
  wire _abc_15724_n4085;
  wire _abc_15724_n4086;
  wire _abc_15724_n4087;
  wire _abc_15724_n4088;
  wire _abc_15724_n4089;
  wire _abc_15724_n4090;
  wire _abc_15724_n4091;
  wire _abc_15724_n4092;
  wire _abc_15724_n4093;
  wire _abc_15724_n4094;
  wire _abc_15724_n4095;
  wire _abc_15724_n4096;
  wire _abc_15724_n4097;
  wire _abc_15724_n4098;
  wire _abc_15724_n4099;
  wire _abc_15724_n4101;
  wire _abc_15724_n4102;
  wire _abc_15724_n4103;
  wire _abc_15724_n4104;
  wire _abc_15724_n4105;
  wire _abc_15724_n4106;
  wire _abc_15724_n4107;
  wire _abc_15724_n4108;
  wire _abc_15724_n4109;
  wire _abc_15724_n4110;
  wire _abc_15724_n4111;
  wire _abc_15724_n4112;
  wire _abc_15724_n4113;
  wire _abc_15724_n4114;
  wire _abc_15724_n4115;
  wire _abc_15724_n4116;
  wire _abc_15724_n4117;
  wire _abc_15724_n4118;
  wire _abc_15724_n4119;
  wire _abc_15724_n4120;
  wire _abc_15724_n4121;
  wire _abc_15724_n4122;
  wire _abc_15724_n4123;
  wire _abc_15724_n4124;
  wire _abc_15724_n4125;
  wire _abc_15724_n4126;
  wire _abc_15724_n4127;
  wire _abc_15724_n4128;
  wire _abc_15724_n4129;
  wire _abc_15724_n4130;
  wire _abc_15724_n4131;
  wire _abc_15724_n4132;
  wire _abc_15724_n4133;
  wire _abc_15724_n4134;
  wire _abc_15724_n4135;
  wire _abc_15724_n4136;
  wire _abc_15724_n4137;
  wire _abc_15724_n4138;
  wire _abc_15724_n4139;
  wire _abc_15724_n4140;
  wire _abc_15724_n4141;
  wire _abc_15724_n4142;
  wire _abc_15724_n4143;
  wire _abc_15724_n4144;
  wire _abc_15724_n4145;
  wire _abc_15724_n4146;
  wire _abc_15724_n4147;
  wire _abc_15724_n4148;
  wire _abc_15724_n4149;
  wire _abc_15724_n4150;
  wire _abc_15724_n4151;
  wire _abc_15724_n4152;
  wire _abc_15724_n4153;
  wire _abc_15724_n4154;
  wire _abc_15724_n4155;
  wire _abc_15724_n4156;
  wire _abc_15724_n4157;
  wire _abc_15724_n4158;
  wire _abc_15724_n4159;
  wire _abc_15724_n4160;
  wire _abc_15724_n4161;
  wire _abc_15724_n4162;
  wire _abc_15724_n4163;
  wire _abc_15724_n4164;
  wire _abc_15724_n4165;
  wire _abc_15724_n4166;
  wire _abc_15724_n4167;
  wire _abc_15724_n4168;
  wire _abc_15724_n4169;
  wire _abc_15724_n4170;
  wire _abc_15724_n4171;
  wire _abc_15724_n4172;
  wire _abc_15724_n4173;
  wire _abc_15724_n4174;
  wire _abc_15724_n4175;
  wire _abc_15724_n4176;
  wire _abc_15724_n4177;
  wire _abc_15724_n4178;
  wire _abc_15724_n4179;
  wire _abc_15724_n4180;
  wire _abc_15724_n4181;
  wire _abc_15724_n4182;
  wire _abc_15724_n4183;
  wire _abc_15724_n4184;
  wire _abc_15724_n4185;
  wire _abc_15724_n4186;
  wire _abc_15724_n4187;
  wire _abc_15724_n4189;
  wire _abc_15724_n4190;
  wire _abc_15724_n4191;
  wire _abc_15724_n4192;
  wire _abc_15724_n4193;
  wire _abc_15724_n4194;
  wire _abc_15724_n4195;
  wire _abc_15724_n4196;
  wire _abc_15724_n4197;
  wire _abc_15724_n4198;
  wire _abc_15724_n4199;
  wire _abc_15724_n4200;
  wire _abc_15724_n4201;
  wire _abc_15724_n4202;
  wire _abc_15724_n4203;
  wire _abc_15724_n4204;
  wire _abc_15724_n4205;
  wire _abc_15724_n4206;
  wire _abc_15724_n4207;
  wire _abc_15724_n4208;
  wire _abc_15724_n4209;
  wire _abc_15724_n4210;
  wire _abc_15724_n4211;
  wire _abc_15724_n4212;
  wire _abc_15724_n4213;
  wire _abc_15724_n4214;
  wire _abc_15724_n4215;
  wire _abc_15724_n4216;
  wire _abc_15724_n4217;
  wire _abc_15724_n4218;
  wire _abc_15724_n4219;
  wire _abc_15724_n4220;
  wire _abc_15724_n4221;
  wire _abc_15724_n4222;
  wire _abc_15724_n4223;
  wire _abc_15724_n4224;
  wire _abc_15724_n4225;
  wire _abc_15724_n4226;
  wire _abc_15724_n4227;
  wire _abc_15724_n4228;
  wire _abc_15724_n4229;
  wire _abc_15724_n4230;
  wire _abc_15724_n4231;
  wire _abc_15724_n4232;
  wire _abc_15724_n4233;
  wire _abc_15724_n4234;
  wire _abc_15724_n4235;
  wire _abc_15724_n4236;
  wire _abc_15724_n4237;
  wire _abc_15724_n4238;
  wire _abc_15724_n4239;
  wire _abc_15724_n4240;
  wire _abc_15724_n4241;
  wire _abc_15724_n4242;
  wire _abc_15724_n4243;
  wire _abc_15724_n4244;
  wire _abc_15724_n4245;
  wire _abc_15724_n4246;
  wire _abc_15724_n4247;
  wire _abc_15724_n4248;
  wire _abc_15724_n4249;
  wire _abc_15724_n4250;
  wire _abc_15724_n4251;
  wire _abc_15724_n4252;
  wire _abc_15724_n4253;
  wire _abc_15724_n4254;
  wire _abc_15724_n4255;
  wire _abc_15724_n4256;
  wire _abc_15724_n4257;
  wire _abc_15724_n4258;
  wire _abc_15724_n4259;
  wire _abc_15724_n4260;
  wire _abc_15724_n4261;
  wire _abc_15724_n4262;
  wire _abc_15724_n4263;
  wire _abc_15724_n4264;
  wire _abc_15724_n4265;
  wire _abc_15724_n4266;
  wire _abc_15724_n4267;
  wire _abc_15724_n4268;
  wire _abc_15724_n4270;
  wire _abc_15724_n4271;
  wire _abc_15724_n4272;
  wire _abc_15724_n4273;
  wire _abc_15724_n4274;
  wire _abc_15724_n4275;
  wire _abc_15724_n4276;
  wire _abc_15724_n4277;
  wire _abc_15724_n4278;
  wire _abc_15724_n4279;
  wire _abc_15724_n4280;
  wire _abc_15724_n4281;
  wire _abc_15724_n4282;
  wire _abc_15724_n4283;
  wire _abc_15724_n4284;
  wire _abc_15724_n4285;
  wire _abc_15724_n4286;
  wire _abc_15724_n4287;
  wire _abc_15724_n4288;
  wire _abc_15724_n4289;
  wire _abc_15724_n4290;
  wire _abc_15724_n4291;
  wire _abc_15724_n4292;
  wire _abc_15724_n4293;
  wire _abc_15724_n4294;
  wire _abc_15724_n4295;
  wire _abc_15724_n4296;
  wire _abc_15724_n4297;
  wire _abc_15724_n4298;
  wire _abc_15724_n4299;
  wire _abc_15724_n4300;
  wire _abc_15724_n4301;
  wire _abc_15724_n4302;
  wire _abc_15724_n4303;
  wire _abc_15724_n4304;
  wire _abc_15724_n4305;
  wire _abc_15724_n4306;
  wire _abc_15724_n4307;
  wire _abc_15724_n4308;
  wire _abc_15724_n4309;
  wire _abc_15724_n4310;
  wire _abc_15724_n4311;
  wire _abc_15724_n4312;
  wire _abc_15724_n4313;
  wire _abc_15724_n4314;
  wire _abc_15724_n4315;
  wire _abc_15724_n4316;
  wire _abc_15724_n4317;
  wire _abc_15724_n4318;
  wire _abc_15724_n4319;
  wire _abc_15724_n4320;
  wire _abc_15724_n4321;
  wire _abc_15724_n4322;
  wire _abc_15724_n4323;
  wire _abc_15724_n4324;
  wire _abc_15724_n4325;
  wire _abc_15724_n4326;
  wire _abc_15724_n4327;
  wire _abc_15724_n4328;
  wire _abc_15724_n4329;
  wire _abc_15724_n4330;
  wire _abc_15724_n4331;
  wire _abc_15724_n4332;
  wire _abc_15724_n4333;
  wire _abc_15724_n4334;
  wire _abc_15724_n4335;
  wire _abc_15724_n4336;
  wire _abc_15724_n4337;
  wire _abc_15724_n4338;
  wire _abc_15724_n4339;
  wire _abc_15724_n4340;
  wire _abc_15724_n4341;
  wire _abc_15724_n4342;
  wire _abc_15724_n4344;
  wire _abc_15724_n4345;
  wire _abc_15724_n4346;
  wire _abc_15724_n4347;
  wire _abc_15724_n4348;
  wire _abc_15724_n4349;
  wire _abc_15724_n4350;
  wire _abc_15724_n4351;
  wire _abc_15724_n4352;
  wire _abc_15724_n4353;
  wire _abc_15724_n4354;
  wire _abc_15724_n4355;
  wire _abc_15724_n4356;
  wire _abc_15724_n4357;
  wire _abc_15724_n4358;
  wire _abc_15724_n4359;
  wire _abc_15724_n4360;
  wire _abc_15724_n4361;
  wire _abc_15724_n4362;
  wire _abc_15724_n4363;
  wire _abc_15724_n4364;
  wire _abc_15724_n4365;
  wire _abc_15724_n4366;
  wire _abc_15724_n4367;
  wire _abc_15724_n4368;
  wire _abc_15724_n4369;
  wire _abc_15724_n4370;
  wire _abc_15724_n4371;
  wire _abc_15724_n4372;
  wire _abc_15724_n4373;
  wire _abc_15724_n4374;
  wire _abc_15724_n4375;
  wire _abc_15724_n4376;
  wire _abc_15724_n4377;
  wire _abc_15724_n4378;
  wire _abc_15724_n4379;
  wire _abc_15724_n4380;
  wire _abc_15724_n4381;
  wire _abc_15724_n4382;
  wire _abc_15724_n4383;
  wire _abc_15724_n4384;
  wire _abc_15724_n4385;
  wire _abc_15724_n4386;
  wire _abc_15724_n4387;
  wire _abc_15724_n4388;
  wire _abc_15724_n4389;
  wire _abc_15724_n4390;
  wire _abc_15724_n4391;
  wire _abc_15724_n4392;
  wire _abc_15724_n4393;
  wire _abc_15724_n4394;
  wire _abc_15724_n4395;
  wire _abc_15724_n4396;
  wire _abc_15724_n4397;
  wire _abc_15724_n4398;
  wire _abc_15724_n4399;
  wire _abc_15724_n4400;
  wire _abc_15724_n4401;
  wire _abc_15724_n4402;
  wire _abc_15724_n4403;
  wire _abc_15724_n4404;
  wire _abc_15724_n4405;
  wire _abc_15724_n4406;
  wire _abc_15724_n4407;
  wire _abc_15724_n4408;
  wire _abc_15724_n4409;
  wire _abc_15724_n4410;
  wire _abc_15724_n4411;
  wire _abc_15724_n4412;
  wire _abc_15724_n4413;
  wire _abc_15724_n4414;
  wire _abc_15724_n4415;
  wire _abc_15724_n4416;
  wire _abc_15724_n4417;
  wire _abc_15724_n4418;
  wire _abc_15724_n4419;
  wire _abc_15724_n4420;
  wire _abc_15724_n4421;
  wire _abc_15724_n4422;
  wire _abc_15724_n4423;
  wire _abc_15724_n4424;
  wire _abc_15724_n4425;
  wire _abc_15724_n4426;
  wire _abc_15724_n4427;
  wire _abc_15724_n4428;
  wire _abc_15724_n4429;
  wire _abc_15724_n4430;
  wire _abc_15724_n4432;
  wire _abc_15724_n4433;
  wire _abc_15724_n4434;
  wire _abc_15724_n4435;
  wire _abc_15724_n4436;
  wire _abc_15724_n4437;
  wire _abc_15724_n4438;
  wire _abc_15724_n4439;
  wire _abc_15724_n4440;
  wire _abc_15724_n4441;
  wire _abc_15724_n4442;
  wire _abc_15724_n4443;
  wire _abc_15724_n4444;
  wire _abc_15724_n4445;
  wire _abc_15724_n4446;
  wire _abc_15724_n4447;
  wire _abc_15724_n4448;
  wire _abc_15724_n4449;
  wire _abc_15724_n4450;
  wire _abc_15724_n4451;
  wire _abc_15724_n4452;
  wire _abc_15724_n4453;
  wire _abc_15724_n4454;
  wire _abc_15724_n4455;
  wire _abc_15724_n4456;
  wire _abc_15724_n4457;
  wire _abc_15724_n4458;
  wire _abc_15724_n4459;
  wire _abc_15724_n4460;
  wire _abc_15724_n4461;
  wire _abc_15724_n4462;
  wire _abc_15724_n4463;
  wire _abc_15724_n4464;
  wire _abc_15724_n4465;
  wire _abc_15724_n4466;
  wire _abc_15724_n4467;
  wire _abc_15724_n4468;
  wire _abc_15724_n4469;
  wire _abc_15724_n4470;
  wire _abc_15724_n4471;
  wire _abc_15724_n4472;
  wire _abc_15724_n4473;
  wire _abc_15724_n4474;
  wire _abc_15724_n4475;
  wire _abc_15724_n4476;
  wire _abc_15724_n4477;
  wire _abc_15724_n4478;
  wire _abc_15724_n4479;
  wire _abc_15724_n4480;
  wire _abc_15724_n4481;
  wire _abc_15724_n4482;
  wire _abc_15724_n4483;
  wire _abc_15724_n4484;
  wire _abc_15724_n4485;
  wire _abc_15724_n4486;
  wire _abc_15724_n4487;
  wire _abc_15724_n4488;
  wire _abc_15724_n4489;
  wire _abc_15724_n4490;
  wire _abc_15724_n4491;
  wire _abc_15724_n4492;
  wire _abc_15724_n4493;
  wire _abc_15724_n4494;
  wire _abc_15724_n4495;
  wire _abc_15724_n4496;
  wire _abc_15724_n4497;
  wire _abc_15724_n4498;
  wire _abc_15724_n4499;
  wire _abc_15724_n4500;
  wire _abc_15724_n4501;
  wire _abc_15724_n4502;
  wire _abc_15724_n4503;
  wire _abc_15724_n4504;
  wire _abc_15724_n4505;
  wire _abc_15724_n4506;
  wire _abc_15724_n4507;
  wire _abc_15724_n4508;
  wire _abc_15724_n4509;
  wire _abc_15724_n4510;
  wire _abc_15724_n4511;
  wire _abc_15724_n4512;
  wire _abc_15724_n4513;
  wire _abc_15724_n4514;
  wire _abc_15724_n4515;
  wire _abc_15724_n4517;
  wire _abc_15724_n4518;
  wire _abc_15724_n4519;
  wire _abc_15724_n4520;
  wire _abc_15724_n4521;
  wire _abc_15724_n4522;
  wire _abc_15724_n4523;
  wire _abc_15724_n4524;
  wire _abc_15724_n4525;
  wire _abc_15724_n4526;
  wire _abc_15724_n4527;
  wire _abc_15724_n4528;
  wire _abc_15724_n4529;
  wire _abc_15724_n4530;
  wire _abc_15724_n4531;
  wire _abc_15724_n4532;
  wire _abc_15724_n4533;
  wire _abc_15724_n4534;
  wire _abc_15724_n4535;
  wire _abc_15724_n4536;
  wire _abc_15724_n4537;
  wire _abc_15724_n4538;
  wire _abc_15724_n4539;
  wire _abc_15724_n4540;
  wire _abc_15724_n4541;
  wire _abc_15724_n4542;
  wire _abc_15724_n4543;
  wire _abc_15724_n4544;
  wire _abc_15724_n4545;
  wire _abc_15724_n4546;
  wire _abc_15724_n4547;
  wire _abc_15724_n4548;
  wire _abc_15724_n4549;
  wire _abc_15724_n4550;
  wire _abc_15724_n4551;
  wire _abc_15724_n4552;
  wire _abc_15724_n4553;
  wire _abc_15724_n4554;
  wire _abc_15724_n4555;
  wire _abc_15724_n4556;
  wire _abc_15724_n4557;
  wire _abc_15724_n4558;
  wire _abc_15724_n4559;
  wire _abc_15724_n4560;
  wire _abc_15724_n4561;
  wire _abc_15724_n4562;
  wire _abc_15724_n4563;
  wire _abc_15724_n4564;
  wire _abc_15724_n4565;
  wire _abc_15724_n4566;
  wire _abc_15724_n4567;
  wire _abc_15724_n4568;
  wire _abc_15724_n4569;
  wire _abc_15724_n4570;
  wire _abc_15724_n4571;
  wire _abc_15724_n4572;
  wire _abc_15724_n4573;
  wire _abc_15724_n4574;
  wire _abc_15724_n4575;
  wire _abc_15724_n4576;
  wire _abc_15724_n4577;
  wire _abc_15724_n4578;
  wire _abc_15724_n4579;
  wire _abc_15724_n4580;
  wire _abc_15724_n4581;
  wire _abc_15724_n4582;
  wire _abc_15724_n4583;
  wire _abc_15724_n4584;
  wire _abc_15724_n4585;
  wire _abc_15724_n4586;
  wire _abc_15724_n4587;
  wire _abc_15724_n4588;
  wire _abc_15724_n4589;
  wire _abc_15724_n4590;
  wire _abc_15724_n4591;
  wire _abc_15724_n4592;
  wire _abc_15724_n4593;
  wire _abc_15724_n4594;
  wire _abc_15724_n4595;
  wire _abc_15724_n4597;
  wire _abc_15724_n4598;
  wire _abc_15724_n4599;
  wire _abc_15724_n4600;
  wire _abc_15724_n4601;
  wire _abc_15724_n4602;
  wire _abc_15724_n4603;
  wire _abc_15724_n4604;
  wire _abc_15724_n4605;
  wire _abc_15724_n4606;
  wire _abc_15724_n4607;
  wire _abc_15724_n4608;
  wire _abc_15724_n4609;
  wire _abc_15724_n4610;
  wire _abc_15724_n4611;
  wire _abc_15724_n4612;
  wire _abc_15724_n4613;
  wire _abc_15724_n4614;
  wire _abc_15724_n4615;
  wire _abc_15724_n4616;
  wire _abc_15724_n4617;
  wire _abc_15724_n4618;
  wire _abc_15724_n4619;
  wire _abc_15724_n4620;
  wire _abc_15724_n4621;
  wire _abc_15724_n4622;
  wire _abc_15724_n4623;
  wire _abc_15724_n4624;
  wire _abc_15724_n4625;
  wire _abc_15724_n4626;
  wire _abc_15724_n4627;
  wire _abc_15724_n4628;
  wire _abc_15724_n4629;
  wire _abc_15724_n4630;
  wire _abc_15724_n4631;
  wire _abc_15724_n4632;
  wire _abc_15724_n4633;
  wire _abc_15724_n4634;
  wire _abc_15724_n4635;
  wire _abc_15724_n4636;
  wire _abc_15724_n4637;
  wire _abc_15724_n4638;
  wire _abc_15724_n4639;
  wire _abc_15724_n4640;
  wire _abc_15724_n4641;
  wire _abc_15724_n4642;
  wire _abc_15724_n4643;
  wire _abc_15724_n4644;
  wire _abc_15724_n4645;
  wire _abc_15724_n4646;
  wire _abc_15724_n4647;
  wire _abc_15724_n4648;
  wire _abc_15724_n4649;
  wire _abc_15724_n4650;
  wire _abc_15724_n4651;
  wire _abc_15724_n4652;
  wire _abc_15724_n4653;
  wire _abc_15724_n4654;
  wire _abc_15724_n4655;
  wire _abc_15724_n4656;
  wire _abc_15724_n4657;
  wire _abc_15724_n4658;
  wire _abc_15724_n4659;
  wire _abc_15724_n4660;
  wire _abc_15724_n4661;
  wire _abc_15724_n4662;
  wire _abc_15724_n4663;
  wire _abc_15724_n4664;
  wire _abc_15724_n4665;
  wire _abc_15724_n4666;
  wire _abc_15724_n4667;
  wire _abc_15724_n4668;
  wire _abc_15724_n4669;
  wire _abc_15724_n4670;
  wire _abc_15724_n4671;
  wire _abc_15724_n4672;
  wire _abc_15724_n4673;
  wire _abc_15724_n4675;
  wire _abc_15724_n4676;
  wire _abc_15724_n4677;
  wire _abc_15724_n4678;
  wire _abc_15724_n4679;
  wire _abc_15724_n4680;
  wire _abc_15724_n4681;
  wire _abc_15724_n4682;
  wire _abc_15724_n4683;
  wire _abc_15724_n4684;
  wire _abc_15724_n4685;
  wire _abc_15724_n4686;
  wire _abc_15724_n4687;
  wire _abc_15724_n4688;
  wire _abc_15724_n4689;
  wire _abc_15724_n4690;
  wire _abc_15724_n4691;
  wire _abc_15724_n4692;
  wire _abc_15724_n4693;
  wire _abc_15724_n4694;
  wire _abc_15724_n4695;
  wire _abc_15724_n4696;
  wire _abc_15724_n4697;
  wire _abc_15724_n4698;
  wire _abc_15724_n4699;
  wire _abc_15724_n4700;
  wire _abc_15724_n4701;
  wire _abc_15724_n4702;
  wire _abc_15724_n4703;
  wire _abc_15724_n4704;
  wire _abc_15724_n4705;
  wire _abc_15724_n4706;
  wire _abc_15724_n4707;
  wire _abc_15724_n4708;
  wire _abc_15724_n4709;
  wire _abc_15724_n4710;
  wire _abc_15724_n4711;
  wire _abc_15724_n4712;
  wire _abc_15724_n4713;
  wire _abc_15724_n4714;
  wire _abc_15724_n4715;
  wire _abc_15724_n4716;
  wire _abc_15724_n4717;
  wire _abc_15724_n4718;
  wire _abc_15724_n4719;
  wire _abc_15724_n4720;
  wire _abc_15724_n4721;
  wire _abc_15724_n4722;
  wire _abc_15724_n4723;
  wire _abc_15724_n4724;
  wire _abc_15724_n4725;
  wire _abc_15724_n4726;
  wire _abc_15724_n4727;
  wire _abc_15724_n4728;
  wire _abc_15724_n4729;
  wire _abc_15724_n4730;
  wire _abc_15724_n4731;
  wire _abc_15724_n4732;
  wire _abc_15724_n4733;
  wire _abc_15724_n4734;
  wire _abc_15724_n4735;
  wire _abc_15724_n4736;
  wire _abc_15724_n4737;
  wire _abc_15724_n4738;
  wire _abc_15724_n4739;
  wire _abc_15724_n4740;
  wire _abc_15724_n4741;
  wire _abc_15724_n4742;
  wire _abc_15724_n4743;
  wire _abc_15724_n4744;
  wire _abc_15724_n4745;
  wire _abc_15724_n4746;
  wire _abc_15724_n4747;
  wire _abc_15724_n4748;
  wire _abc_15724_n4749;
  wire _abc_15724_n4750;
  wire _abc_15724_n4751;
  wire _abc_15724_n4752;
  wire _abc_15724_n4753;
  wire _abc_15724_n4754;
  wire _abc_15724_n4755;
  wire _abc_15724_n4756;
  wire _abc_15724_n4758;
  wire _abc_15724_n4759;
  wire _abc_15724_n4760;
  wire _abc_15724_n4761;
  wire _abc_15724_n4762;
  wire _abc_15724_n4763;
  wire _abc_15724_n4764;
  wire _abc_15724_n4765;
  wire _abc_15724_n4766;
  wire _abc_15724_n4767;
  wire _abc_15724_n4768;
  wire _abc_15724_n4769;
  wire _abc_15724_n4770;
  wire _abc_15724_n4771;
  wire _abc_15724_n4772;
  wire _abc_15724_n4773;
  wire _abc_15724_n4774;
  wire _abc_15724_n4775;
  wire _abc_15724_n4776;
  wire _abc_15724_n4777;
  wire _abc_15724_n4778;
  wire _abc_15724_n4779;
  wire _abc_15724_n4780;
  wire _abc_15724_n4781;
  wire _abc_15724_n4782;
  wire _abc_15724_n4783;
  wire _abc_15724_n4784;
  wire _abc_15724_n4785;
  wire _abc_15724_n4786;
  wire _abc_15724_n4787;
  wire _abc_15724_n4788;
  wire _abc_15724_n4789;
  wire _abc_15724_n4790;
  wire _abc_15724_n4791;
  wire _abc_15724_n4792;
  wire _abc_15724_n4793;
  wire _abc_15724_n4794;
  wire _abc_15724_n4795;
  wire _abc_15724_n4796;
  wire _abc_15724_n4797;
  wire _abc_15724_n4798;
  wire _abc_15724_n4799;
  wire _abc_15724_n4800;
  wire _abc_15724_n4801;
  wire _abc_15724_n4802;
  wire _abc_15724_n4803;
  wire _abc_15724_n4804;
  wire _abc_15724_n4805;
  wire _abc_15724_n4806;
  wire _abc_15724_n4807;
  wire _abc_15724_n4808;
  wire _abc_15724_n4809;
  wire _abc_15724_n4810;
  wire _abc_15724_n4811;
  wire _abc_15724_n4812;
  wire _abc_15724_n4813;
  wire _abc_15724_n4814;
  wire _abc_15724_n4815;
  wire _abc_15724_n4816;
  wire _abc_15724_n4817;
  wire _abc_15724_n4818;
  wire _abc_15724_n4819;
  wire _abc_15724_n4820;
  wire _abc_15724_n4821;
  wire _abc_15724_n4822;
  wire _abc_15724_n4823;
  wire _abc_15724_n4824;
  wire _abc_15724_n4825;
  wire _abc_15724_n4826;
  wire _abc_15724_n4827;
  wire _abc_15724_n4828;
  wire _abc_15724_n4829;
  wire _abc_15724_n4830;
  wire _abc_15724_n4831;
  wire _abc_15724_n4832;
  wire _abc_15724_n4833;
  wire _abc_15724_n4834;
  wire _abc_15724_n4835;
  wire _abc_15724_n4836;
  wire _abc_15724_n4838;
  wire _abc_15724_n4839;
  wire _abc_15724_n4840;
  wire _abc_15724_n4841;
  wire _abc_15724_n4842;
  wire _abc_15724_n4843;
  wire _abc_15724_n4844;
  wire _abc_15724_n4845;
  wire _abc_15724_n4846;
  wire _abc_15724_n4847;
  wire _abc_15724_n4848;
  wire _abc_15724_n4849;
  wire _abc_15724_n4850;
  wire _abc_15724_n4851;
  wire _abc_15724_n4852;
  wire _abc_15724_n4853;
  wire _abc_15724_n4854;
  wire _abc_15724_n4855;
  wire _abc_15724_n4856;
  wire _abc_15724_n4857;
  wire _abc_15724_n4858;
  wire _abc_15724_n4859;
  wire _abc_15724_n4860;
  wire _abc_15724_n4861;
  wire _abc_15724_n4862;
  wire _abc_15724_n4863;
  wire _abc_15724_n4864;
  wire _abc_15724_n4865;
  wire _abc_15724_n4866;
  wire _abc_15724_n4867;
  wire _abc_15724_n4868;
  wire _abc_15724_n4869;
  wire _abc_15724_n4870;
  wire _abc_15724_n4871;
  wire _abc_15724_n4872;
  wire _abc_15724_n4873;
  wire _abc_15724_n4874;
  wire _abc_15724_n4875;
  wire _abc_15724_n4876;
  wire _abc_15724_n4877;
  wire _abc_15724_n4878;
  wire _abc_15724_n4879;
  wire _abc_15724_n4880;
  wire _abc_15724_n4881;
  wire _abc_15724_n4882;
  wire _abc_15724_n4883;
  wire _abc_15724_n4884;
  wire _abc_15724_n4885;
  wire _abc_15724_n4886;
  wire _abc_15724_n4887;
  wire _abc_15724_n4888;
  wire _abc_15724_n4889;
  wire _abc_15724_n4890;
  wire _abc_15724_n4891;
  wire _abc_15724_n4892;
  wire _abc_15724_n4893;
  wire _abc_15724_n4894;
  wire _abc_15724_n4895;
  wire _abc_15724_n4896;
  wire _abc_15724_n4897;
  wire _abc_15724_n4898;
  wire _abc_15724_n4899;
  wire _abc_15724_n4900;
  wire _abc_15724_n4901;
  wire _abc_15724_n4902;
  wire _abc_15724_n4903;
  wire _abc_15724_n4904;
  wire _abc_15724_n4905;
  wire _abc_15724_n4906;
  wire _abc_15724_n4907;
  wire _abc_15724_n4908;
  wire _abc_15724_n4909;
  wire _abc_15724_n4910;
  wire _abc_15724_n4911;
  wire _abc_15724_n4912;
  wire _abc_15724_n4914;
  wire _abc_15724_n4915;
  wire _abc_15724_n4916;
  wire _abc_15724_n4917;
  wire _abc_15724_n4918;
  wire _abc_15724_n4919;
  wire _abc_15724_n4920;
  wire _abc_15724_n4921;
  wire _abc_15724_n4922;
  wire _abc_15724_n4923;
  wire _abc_15724_n4924;
  wire _abc_15724_n4925;
  wire _abc_15724_n4926;
  wire _abc_15724_n4927;
  wire _abc_15724_n4928;
  wire _abc_15724_n4929;
  wire _abc_15724_n4930;
  wire _abc_15724_n4931;
  wire _abc_15724_n4932;
  wire _abc_15724_n4933;
  wire _abc_15724_n4934;
  wire _abc_15724_n4935;
  wire _abc_15724_n4936;
  wire _abc_15724_n4937;
  wire _abc_15724_n4938;
  wire _abc_15724_n4939;
  wire _abc_15724_n4940;
  wire _abc_15724_n4941;
  wire _abc_15724_n4942;
  wire _abc_15724_n4943;
  wire _abc_15724_n4944;
  wire _abc_15724_n4945;
  wire _abc_15724_n4946;
  wire _abc_15724_n4947;
  wire _abc_15724_n4948;
  wire _abc_15724_n4949;
  wire _abc_15724_n4950;
  wire _abc_15724_n4951;
  wire _abc_15724_n4952;
  wire _abc_15724_n4953;
  wire _abc_15724_n4954;
  wire _abc_15724_n4955;
  wire _abc_15724_n4956;
  wire _abc_15724_n4957;
  wire _abc_15724_n4958;
  wire _abc_15724_n4959;
  wire _abc_15724_n4960;
  wire _abc_15724_n4961;
  wire _abc_15724_n4962;
  wire _abc_15724_n4963;
  wire _abc_15724_n4964;
  wire _abc_15724_n4965;
  wire _abc_15724_n4966;
  wire _abc_15724_n4967;
  wire _abc_15724_n4968;
  wire _abc_15724_n4969;
  wire _abc_15724_n4970;
  wire _abc_15724_n4971;
  wire _abc_15724_n4972;
  wire _abc_15724_n4973;
  wire _abc_15724_n4974;
  wire _abc_15724_n4975;
  wire _abc_15724_n4976;
  wire _abc_15724_n4977;
  wire _abc_15724_n4978;
  wire _abc_15724_n4979;
  wire _abc_15724_n4980;
  wire _abc_15724_n4981;
  wire _abc_15724_n4982;
  wire _abc_15724_n4983;
  wire _abc_15724_n4984;
  wire _abc_15724_n4985;
  wire _abc_15724_n4986;
  wire _abc_15724_n4987;
  wire _abc_15724_n4988;
  wire _abc_15724_n4989;
  wire _abc_15724_n4991;
  wire _abc_15724_n4992;
  wire _abc_15724_n4993;
  wire _abc_15724_n4994;
  wire _abc_15724_n4995;
  wire _abc_15724_n4996;
  wire _abc_15724_n4997;
  wire _abc_15724_n4998;
  wire _abc_15724_n4999;
  wire _abc_15724_n5000;
  wire _abc_15724_n5001;
  wire _abc_15724_n5002;
  wire _abc_15724_n5003;
  wire _abc_15724_n5004;
  wire _abc_15724_n5005;
  wire _abc_15724_n5006;
  wire _abc_15724_n5007;
  wire _abc_15724_n5008;
  wire _abc_15724_n5009;
  wire _abc_15724_n5010;
  wire _abc_15724_n5011;
  wire _abc_15724_n5012;
  wire _abc_15724_n5013;
  wire _abc_15724_n5014;
  wire _abc_15724_n5015;
  wire _abc_15724_n5016;
  wire _abc_15724_n5017;
  wire _abc_15724_n5018;
  wire _abc_15724_n5019;
  wire _abc_15724_n5020;
  wire _abc_15724_n5021;
  wire _abc_15724_n5022;
  wire _abc_15724_n5023;
  wire _abc_15724_n5024;
  wire _abc_15724_n5025;
  wire _abc_15724_n5026;
  wire _abc_15724_n5027;
  wire _abc_15724_n5028;
  wire _abc_15724_n5029;
  wire _abc_15724_n5030;
  wire _abc_15724_n5031;
  wire _abc_15724_n5032;
  wire _abc_15724_n5033;
  wire _abc_15724_n5034;
  wire _abc_15724_n5035;
  wire _abc_15724_n5036;
  wire _abc_15724_n5037;
  wire _abc_15724_n5038;
  wire _abc_15724_n5039;
  wire _abc_15724_n5040;
  wire _abc_15724_n5041;
  wire _abc_15724_n5042;
  wire _abc_15724_n5043;
  wire _abc_15724_n5044;
  wire _abc_15724_n5045;
  wire _abc_15724_n5046;
  wire _abc_15724_n5047;
  wire _abc_15724_n5048;
  wire _abc_15724_n5049;
  wire _abc_15724_n5050;
  wire _abc_15724_n5051;
  wire _abc_15724_n5052;
  wire _abc_15724_n5053;
  wire _abc_15724_n5054;
  wire _abc_15724_n5055;
  wire _abc_15724_n5056;
  wire _abc_15724_n5057;
  wire _abc_15724_n5058;
  wire _abc_15724_n5059;
  wire _abc_15724_n5060;
  wire _abc_15724_n5061;
  wire _abc_15724_n5062;
  wire _abc_15724_n5063;
  wire _abc_15724_n5064;
  wire _abc_15724_n5065;
  wire _abc_15724_n5066;
  wire _abc_15724_n5067;
  wire _abc_15724_n5068;
  wire _abc_15724_n5069;
  wire _abc_15724_n5070;
  wire _abc_15724_n5071;
  wire _abc_15724_n5072;
  wire _abc_15724_n5074;
  wire _abc_15724_n5075;
  wire _abc_15724_n5076;
  wire _abc_15724_n5077;
  wire _abc_15724_n5078;
  wire _abc_15724_n5079;
  wire _abc_15724_n5080;
  wire _abc_15724_n5081;
  wire _abc_15724_n5082;
  wire _abc_15724_n5083;
  wire _abc_15724_n5084;
  wire _abc_15724_n5085;
  wire _abc_15724_n5086;
  wire _abc_15724_n5087;
  wire _abc_15724_n5088;
  wire _abc_15724_n5089;
  wire _abc_15724_n5090;
  wire _abc_15724_n5091;
  wire _abc_15724_n5092;
  wire _abc_15724_n5093;
  wire _abc_15724_n5094;
  wire _abc_15724_n5095;
  wire _abc_15724_n5096;
  wire _abc_15724_n5097;
  wire _abc_15724_n5098;
  wire _abc_15724_n5099;
  wire _abc_15724_n5100;
  wire _abc_15724_n5101;
  wire _abc_15724_n5102;
  wire _abc_15724_n5103;
  wire _abc_15724_n5104;
  wire _abc_15724_n5105;
  wire _abc_15724_n5106;
  wire _abc_15724_n5107;
  wire _abc_15724_n5108;
  wire _abc_15724_n5109;
  wire _abc_15724_n5110;
  wire _abc_15724_n5111;
  wire _abc_15724_n5112;
  wire _abc_15724_n5113;
  wire _abc_15724_n5114;
  wire _abc_15724_n5115;
  wire _abc_15724_n5116;
  wire _abc_15724_n5117;
  wire _abc_15724_n5118;
  wire _abc_15724_n5119;
  wire _abc_15724_n5120;
  wire _abc_15724_n5121;
  wire _abc_15724_n5122;
  wire _abc_15724_n5123;
  wire _abc_15724_n5124;
  wire _abc_15724_n5125;
  wire _abc_15724_n5126;
  wire _abc_15724_n5127;
  wire _abc_15724_n5128;
  wire _abc_15724_n5129;
  wire _abc_15724_n5130;
  wire _abc_15724_n5131;
  wire _abc_15724_n5132;
  wire _abc_15724_n5133;
  wire _abc_15724_n5134;
  wire _abc_15724_n5135;
  wire _abc_15724_n5136;
  wire _abc_15724_n5137;
  wire _abc_15724_n5138;
  wire _abc_15724_n5140;
  wire _abc_15724_n5141;
  wire _abc_15724_n5142;
  wire _abc_15724_n5143;
  wire _abc_15724_n5144;
  wire _abc_15724_n5145;
  wire _abc_15724_n5146;
  wire _abc_15724_n5147;
  wire _abc_15724_n5148;
  wire _abc_15724_n5149;
  wire _abc_15724_n5150;
  wire _abc_15724_n5151;
  wire _abc_15724_n5152;
  wire _abc_15724_n5153;
  wire _abc_15724_n5154;
  wire _abc_15724_n5155;
  wire _abc_15724_n5156;
  wire _abc_15724_n5157;
  wire _abc_15724_n5158;
  wire _abc_15724_n5159;
  wire _abc_15724_n5160;
  wire _abc_15724_n5161;
  wire _abc_15724_n5162;
  wire _abc_15724_n5163;
  wire _abc_15724_n5164;
  wire _abc_15724_n5165;
  wire _abc_15724_n5166;
  wire _abc_15724_n5167;
  wire _abc_15724_n5168;
  wire _abc_15724_n5169;
  wire _abc_15724_n5170;
  wire _abc_15724_n5171;
  wire _abc_15724_n5172;
  wire _abc_15724_n5173;
  wire _abc_15724_n5174;
  wire _abc_15724_n5175;
  wire _abc_15724_n5176;
  wire _abc_15724_n5177;
  wire _abc_15724_n5178;
  wire _abc_15724_n5179;
  wire _abc_15724_n5180;
  wire _abc_15724_n5181;
  wire _abc_15724_n5182;
  wire _abc_15724_n5183;
  wire _abc_15724_n5184;
  wire _abc_15724_n5185;
  wire _abc_15724_n5186;
  wire _abc_15724_n5187;
  wire _abc_15724_n5188;
  wire _abc_15724_n5189;
  wire _abc_15724_n5190;
  wire _abc_15724_n5191;
  wire _abc_15724_n5192;
  wire _abc_15724_n5193;
  wire _abc_15724_n5194;
  wire _abc_15724_n5195;
  wire _abc_15724_n5196;
  wire _abc_15724_n5197;
  wire _abc_15724_n5198;
  wire _abc_15724_n5199;
  wire _abc_15724_n5200;
  wire _abc_15724_n5201;
  wire _abc_15724_n5203;
  wire _abc_15724_n5204;
  wire _abc_15724_n5205;
  wire _abc_15724_n5206;
  wire _abc_15724_n5207;
  wire _abc_15724_n5208;
  wire _abc_15724_n5209;
  wire _abc_15724_n5210;
  wire _abc_15724_n5211;
  wire _abc_15724_n5212;
  wire _abc_15724_n5213;
  wire _abc_15724_n5214;
  wire _abc_15724_n5215;
  wire _abc_15724_n5216;
  wire _abc_15724_n5217;
  wire _abc_15724_n5218;
  wire _abc_15724_n5219;
  wire _abc_15724_n5220;
  wire _abc_15724_n5221;
  wire _abc_15724_n5222;
  wire _abc_15724_n5223;
  wire _abc_15724_n5224;
  wire _abc_15724_n5225;
  wire _abc_15724_n5226;
  wire _abc_15724_n5227;
  wire _abc_15724_n5228;
  wire _abc_15724_n5229;
  wire _abc_15724_n5230;
  wire _abc_15724_n5231;
  wire _abc_15724_n5232;
  wire _abc_15724_n5233;
  wire _abc_15724_n5234;
  wire _abc_15724_n5235;
  wire _abc_15724_n5236;
  wire _abc_15724_n5237;
  wire _abc_15724_n5238;
  wire _abc_15724_n5239;
  wire _abc_15724_n5240;
  wire _abc_15724_n5241;
  wire _abc_15724_n5242;
  wire _abc_15724_n5243;
  wire _abc_15724_n5244;
  wire _abc_15724_n5245;
  wire _abc_15724_n5246;
  wire _abc_15724_n5247;
  wire _abc_15724_n5248;
  wire _abc_15724_n5249;
  wire _abc_15724_n5250;
  wire _abc_15724_n5251;
  wire _abc_15724_n5252;
  wire _abc_15724_n5253;
  wire _abc_15724_n5254;
  wire _abc_15724_n5255;
  wire _abc_15724_n5256;
  wire _abc_15724_n5257;
  wire _abc_15724_n5258;
  wire _abc_15724_n5259;
  wire _abc_15724_n5260;
  wire _abc_15724_n5261;
  wire _abc_15724_n5262;
  wire _abc_15724_n5263;
  wire _abc_15724_n5264;
  wire _abc_15724_n5265;
  wire _abc_15724_n5266;
  wire _abc_15724_n5267;
  wire _abc_15724_n5268;
  wire _abc_15724_n5269;
  wire _abc_15724_n5271;
  wire _abc_15724_n5272;
  wire _abc_15724_n5273;
  wire _abc_15724_n5274;
  wire _abc_15724_n5275;
  wire _abc_15724_n5276;
  wire _abc_15724_n5277;
  wire _abc_15724_n5278;
  wire _abc_15724_n5279;
  wire _abc_15724_n5280;
  wire _abc_15724_n5281;
  wire _abc_15724_n5282;
  wire _abc_15724_n5283;
  wire _abc_15724_n5284;
  wire _abc_15724_n5285;
  wire _abc_15724_n5286;
  wire _abc_15724_n5287;
  wire _abc_15724_n5288;
  wire _abc_15724_n5289;
  wire _abc_15724_n5290;
  wire _abc_15724_n5291;
  wire _abc_15724_n5292;
  wire _abc_15724_n5293;
  wire _abc_15724_n5294;
  wire _abc_15724_n5295;
  wire _abc_15724_n5296;
  wire _abc_15724_n5297;
  wire _abc_15724_n5298;
  wire _abc_15724_n5299;
  wire _abc_15724_n5300;
  wire _abc_15724_n5301;
  wire _abc_15724_n5302;
  wire _abc_15724_n5303;
  wire _abc_15724_n5304;
  wire _abc_15724_n5305;
  wire _abc_15724_n5306;
  wire _abc_15724_n5307;
  wire _abc_15724_n5308;
  wire _abc_15724_n5309;
  wire _abc_15724_n5310;
  wire _abc_15724_n5311;
  wire _abc_15724_n5312;
  wire _abc_15724_n5313;
  wire _abc_15724_n5314;
  wire _abc_15724_n5315;
  wire _abc_15724_n5316;
  wire _abc_15724_n5317;
  wire _abc_15724_n5318;
  wire _abc_15724_n5319;
  wire _abc_15724_n5320;
  wire _abc_15724_n5321;
  wire _abc_15724_n5322;
  wire _abc_15724_n5323;
  wire _abc_15724_n5324;
  wire _abc_15724_n5325;
  wire _abc_15724_n5326;
  wire _abc_15724_n5327;
  wire _abc_15724_n5328;
  wire _abc_15724_n5329;
  wire _abc_15724_n5330;
  wire _abc_15724_n5331;
  wire _abc_15724_n5332;
  wire _abc_15724_n5333;
  wire _abc_15724_n5334;
  wire _abc_15724_n5335;
  wire _abc_15724_n5336;
  wire _abc_15724_n5337;
  wire _abc_15724_n5338;
  wire _abc_15724_n5339;
  wire _abc_15724_n5340;
  wire _abc_15724_n5341;
  wire _abc_15724_n5342;
  wire _abc_15724_n5343;
  wire _abc_15724_n5344;
  wire _abc_15724_n5345;
  wire _abc_15724_n5346;
  wire _abc_15724_n5347;
  wire _abc_15724_n5348;
  wire _abc_15724_n5349;
  wire _abc_15724_n5350;
  wire _abc_15724_n5352;
  wire _abc_15724_n5353;
  wire _abc_15724_n5354;
  wire _abc_15724_n5355;
  wire _abc_15724_n5356;
  wire _abc_15724_n5357;
  wire _abc_15724_n5358;
  wire _abc_15724_n5359;
  wire _abc_15724_n5360;
  wire _abc_15724_n5361;
  wire _abc_15724_n5362;
  wire _abc_15724_n5363;
  wire _abc_15724_n5364;
  wire _abc_15724_n5365;
  wire _abc_15724_n5366;
  wire _abc_15724_n5367;
  wire _abc_15724_n5368;
  wire _abc_15724_n5369;
  wire _abc_15724_n5370;
  wire _abc_15724_n5371;
  wire _abc_15724_n5372;
  wire _abc_15724_n5373;
  wire _abc_15724_n5374;
  wire _abc_15724_n5375;
  wire _abc_15724_n5376;
  wire _abc_15724_n5377;
  wire _abc_15724_n5378;
  wire _abc_15724_n5379;
  wire _abc_15724_n5380;
  wire _abc_15724_n5381;
  wire _abc_15724_n5382;
  wire _abc_15724_n5383;
  wire _abc_15724_n5384;
  wire _abc_15724_n5385;
  wire _abc_15724_n5386;
  wire _abc_15724_n5387;
  wire _abc_15724_n5388;
  wire _abc_15724_n5389;
  wire _abc_15724_n5390;
  wire _abc_15724_n5391;
  wire _abc_15724_n5392;
  wire _abc_15724_n5393;
  wire _abc_15724_n5394;
  wire _abc_15724_n5395;
  wire _abc_15724_n5396;
  wire _abc_15724_n5397;
  wire _abc_15724_n5398;
  wire _abc_15724_n5399;
  wire _abc_15724_n5400;
  wire _abc_15724_n5401;
  wire _abc_15724_n5402;
  wire _abc_15724_n5403;
  wire _abc_15724_n5404;
  wire _abc_15724_n5405;
  wire _abc_15724_n5406;
  wire _abc_15724_n5407;
  wire _abc_15724_n5408;
  wire _abc_15724_n5409;
  wire _abc_15724_n5410;
  wire _abc_15724_n5411;
  wire _abc_15724_n5412;
  wire _abc_15724_n5413;
  wire _abc_15724_n5414;
  wire _abc_15724_n5415;
  wire _abc_15724_n5416;
  wire _abc_15724_n5417;
  wire _abc_15724_n5418;
  wire _abc_15724_n5419;
  wire _abc_15724_n5420;
  wire _abc_15724_n5421;
  wire _abc_15724_n5422;
  wire _abc_15724_n5423;
  wire _abc_15724_n5425;
  wire _abc_15724_n5426;
  wire _abc_15724_n5427;
  wire _abc_15724_n5428;
  wire _abc_15724_n5429;
  wire _abc_15724_n5430;
  wire _abc_15724_n5431;
  wire _abc_15724_n5432;
  wire _abc_15724_n5433;
  wire _abc_15724_n5434;
  wire _abc_15724_n5435;
  wire _abc_15724_n5436;
  wire _abc_15724_n5437;
  wire _abc_15724_n5438;
  wire _abc_15724_n5439;
  wire _abc_15724_n5440;
  wire _abc_15724_n5441;
  wire _abc_15724_n5442;
  wire _abc_15724_n5443;
  wire _abc_15724_n5444;
  wire _abc_15724_n5445;
  wire _abc_15724_n5446;
  wire _abc_15724_n5447;
  wire _abc_15724_n5448;
  wire _abc_15724_n5449;
  wire _abc_15724_n5450;
  wire _abc_15724_n5451;
  wire _abc_15724_n5452;
  wire _abc_15724_n5453;
  wire _abc_15724_n5454;
  wire _abc_15724_n5455;
  wire _abc_15724_n5456;
  wire _abc_15724_n5457;
  wire _abc_15724_n5458;
  wire _abc_15724_n5459;
  wire _abc_15724_n5460;
  wire _abc_15724_n5461;
  wire _abc_15724_n5462;
  wire _abc_15724_n5463;
  wire _abc_15724_n5464;
  wire _abc_15724_n5465;
  wire _abc_15724_n5466;
  wire _abc_15724_n5467;
  wire _abc_15724_n5468;
  wire _abc_15724_n5469;
  wire _abc_15724_n5470;
  wire _abc_15724_n5471;
  wire _abc_15724_n5472;
  wire _abc_15724_n5473;
  wire _abc_15724_n5474;
  wire _abc_15724_n5475;
  wire _abc_15724_n5476;
  wire _abc_15724_n5477;
  wire _abc_15724_n5478;
  wire _abc_15724_n5479;
  wire _abc_15724_n5480;
  wire _abc_15724_n5481;
  wire _abc_15724_n5482;
  wire _abc_15724_n5483;
  wire _abc_15724_n5484;
  wire _abc_15724_n5485;
  wire _abc_15724_n5486;
  wire _abc_15724_n5487;
  wire _abc_15724_n5488;
  wire _abc_15724_n5489;
  wire _abc_15724_n5490;
  wire _abc_15724_n5491;
  wire _abc_15724_n5492;
  wire _abc_15724_n5493;
  wire _abc_15724_n5495;
  wire _abc_15724_n5496;
  wire _abc_15724_n5497;
  wire _abc_15724_n5498;
  wire _abc_15724_n5499;
  wire _abc_15724_n5500;
  wire _abc_15724_n5501;
  wire _abc_15724_n5502;
  wire _abc_15724_n5503;
  wire _abc_15724_n5504;
  wire _abc_15724_n5505;
  wire _abc_15724_n5506;
  wire _abc_15724_n5507;
  wire _abc_15724_n5508;
  wire _abc_15724_n5509;
  wire _abc_15724_n5510;
  wire _abc_15724_n5511;
  wire _abc_15724_n5512;
  wire _abc_15724_n5513;
  wire _abc_15724_n5514;
  wire _abc_15724_n5515;
  wire _abc_15724_n5516;
  wire _abc_15724_n5517;
  wire _abc_15724_n5518;
  wire _abc_15724_n5519;
  wire _abc_15724_n5520;
  wire _abc_15724_n5521;
  wire _abc_15724_n5522;
  wire _abc_15724_n5523;
  wire _abc_15724_n5524;
  wire _abc_15724_n5525;
  wire _abc_15724_n5526;
  wire _abc_15724_n5527;
  wire _abc_15724_n5528;
  wire _abc_15724_n5529;
  wire _abc_15724_n5530;
  wire _abc_15724_n5531;
  wire _abc_15724_n5532;
  wire _abc_15724_n5533;
  wire _abc_15724_n5534;
  wire _abc_15724_n5535;
  wire _abc_15724_n5536;
  wire _abc_15724_n5537;
  wire _abc_15724_n5538;
  wire _abc_15724_n5539;
  wire _abc_15724_n5540;
  wire _abc_15724_n5541;
  wire _abc_15724_n5542;
  wire _abc_15724_n5543;
  wire _abc_15724_n5544;
  wire _abc_15724_n5545;
  wire _abc_15724_n5546;
  wire _abc_15724_n5547;
  wire _abc_15724_n5548;
  wire _abc_15724_n5549;
  wire _abc_15724_n5550;
  wire _abc_15724_n5551;
  wire _abc_15724_n5552;
  wire _abc_15724_n5553;
  wire _abc_15724_n5554;
  wire _abc_15724_n5555;
  wire _abc_15724_n5556;
  wire _abc_15724_n5557;
  wire _abc_15724_n5558;
  wire _abc_15724_n5559;
  wire _abc_15724_n5560;
  wire _abc_15724_n5562;
  wire _abc_15724_n5563;
  wire _abc_15724_n5564;
  wire _abc_15724_n5565;
  wire _abc_15724_n5566;
  wire _abc_15724_n5567;
  wire _abc_15724_n5568;
  wire _abc_15724_n5569;
  wire _abc_15724_n5570;
  wire _abc_15724_n5571;
  wire _abc_15724_n5572;
  wire _abc_15724_n5573;
  wire _abc_15724_n5574;
  wire _abc_15724_n5575;
  wire _abc_15724_n5576;
  wire _abc_15724_n5577;
  wire _abc_15724_n5578;
  wire _abc_15724_n5579;
  wire _abc_15724_n5580;
  wire _abc_15724_n5581;
  wire _abc_15724_n5582;
  wire _abc_15724_n5583;
  wire _abc_15724_n5584;
  wire _abc_15724_n5585;
  wire _abc_15724_n5586;
  wire _abc_15724_n5587;
  wire _abc_15724_n5588;
  wire _abc_15724_n5589;
  wire _abc_15724_n5590;
  wire _abc_15724_n5591;
  wire _abc_15724_n5592;
  wire _abc_15724_n5593;
  wire _abc_15724_n5594;
  wire _abc_15724_n5595;
  wire _abc_15724_n5596;
  wire _abc_15724_n5597;
  wire _abc_15724_n5598;
  wire _abc_15724_n5599;
  wire _abc_15724_n5600;
  wire _abc_15724_n5601;
  wire _abc_15724_n5602;
  wire _abc_15724_n5603;
  wire _abc_15724_n5604;
  wire _abc_15724_n5605;
  wire _abc_15724_n5606;
  wire _abc_15724_n5607;
  wire _abc_15724_n5608;
  wire _abc_15724_n5609;
  wire _abc_15724_n5610;
  wire _abc_15724_n5611;
  wire _abc_15724_n5612;
  wire _abc_15724_n5613;
  wire _abc_15724_n5614;
  wire _abc_15724_n5615;
  wire _abc_15724_n5616;
  wire _abc_15724_n5617;
  wire _abc_15724_n5618;
  wire _abc_15724_n5619;
  wire _abc_15724_n5620;
  wire _abc_15724_n5621;
  wire _abc_15724_n5622;
  wire _abc_15724_n5623;
  wire _abc_15724_n5624;
  wire _abc_15724_n5625;
  wire _abc_15724_n5626;
  wire _abc_15724_n5627;
  wire _abc_15724_n5628;
  wire _abc_15724_n5629;
  wire _abc_15724_n5630;
  wire _abc_15724_n5631;
  wire _abc_15724_n5632;
  wire _abc_15724_n5633;
  wire _abc_15724_n5634;
  wire _abc_15724_n5635;
  wire _abc_15724_n5636;
  wire _abc_15724_n5637;
  wire _abc_15724_n5638;
  wire _abc_15724_n5639;
  wire _abc_15724_n5641;
  wire _abc_15724_n5642;
  wire _abc_15724_n5643;
  wire _abc_15724_n5644;
  wire _abc_15724_n5645;
  wire _abc_15724_n5646;
  wire _abc_15724_n5647;
  wire _abc_15724_n5648;
  wire _abc_15724_n5649;
  wire _abc_15724_n5650;
  wire _abc_15724_n5651;
  wire _abc_15724_n5652;
  wire _abc_15724_n5653;
  wire _abc_15724_n5654;
  wire _abc_15724_n5655;
  wire _abc_15724_n5656;
  wire _abc_15724_n5657;
  wire _abc_15724_n5658;
  wire _abc_15724_n5659;
  wire _abc_15724_n5660;
  wire _abc_15724_n5661;
  wire _abc_15724_n5662;
  wire _abc_15724_n5663;
  wire _abc_15724_n5664;
  wire _abc_15724_n5665;
  wire _abc_15724_n5666;
  wire _abc_15724_n5667;
  wire _abc_15724_n5668;
  wire _abc_15724_n5669;
  wire _abc_15724_n5670;
  wire _abc_15724_n5671;
  wire _abc_15724_n5672;
  wire _abc_15724_n5673;
  wire _abc_15724_n5674;
  wire _abc_15724_n5675;
  wire _abc_15724_n5676;
  wire _abc_15724_n5677;
  wire _abc_15724_n5678;
  wire _abc_15724_n5679;
  wire _abc_15724_n5680;
  wire _abc_15724_n5681;
  wire _abc_15724_n5682;
  wire _abc_15724_n5683;
  wire _abc_15724_n5684;
  wire _abc_15724_n5685;
  wire _abc_15724_n5686;
  wire _abc_15724_n5687;
  wire _abc_15724_n5688;
  wire _abc_15724_n5689;
  wire _abc_15724_n5690;
  wire _abc_15724_n5691;
  wire _abc_15724_n5692;
  wire _abc_15724_n5693;
  wire _abc_15724_n5694;
  wire _abc_15724_n5695;
  wire _abc_15724_n5696;
  wire _abc_15724_n5697;
  wire _abc_15724_n5698;
  wire _abc_15724_n5699;
  wire _abc_15724_n5700;
  wire _abc_15724_n5701;
  wire _abc_15724_n5702;
  wire _abc_15724_n5703;
  wire _abc_15724_n5704;
  wire _abc_15724_n5706;
  wire _abc_15724_n5707;
  wire _abc_15724_n5708;
  wire _abc_15724_n5709;
  wire _abc_15724_n5710;
  wire _abc_15724_n5711;
  wire _abc_15724_n5712;
  wire _abc_15724_n5713;
  wire _abc_15724_n5714;
  wire _abc_15724_n5715;
  wire _abc_15724_n5716;
  wire _abc_15724_n5717;
  wire _abc_15724_n5718;
  wire _abc_15724_n5719;
  wire _abc_15724_n5720;
  wire _abc_15724_n5721;
  wire _abc_15724_n5722;
  wire _abc_15724_n5723;
  wire _abc_15724_n5724;
  wire _abc_15724_n5725;
  wire _abc_15724_n5726;
  wire _abc_15724_n5727;
  wire _abc_15724_n5728;
  wire _abc_15724_n5729;
  wire _abc_15724_n5730;
  wire _abc_15724_n5731;
  wire _abc_15724_n5732;
  wire _abc_15724_n5733;
  wire _abc_15724_n5734;
  wire _abc_15724_n5735;
  wire _abc_15724_n5736;
  wire _abc_15724_n5737;
  wire _abc_15724_n5738;
  wire _abc_15724_n5739;
  wire _abc_15724_n5740;
  wire _abc_15724_n5741;
  wire _abc_15724_n5742;
  wire _abc_15724_n5743;
  wire _abc_15724_n5744;
  wire _abc_15724_n5745;
  wire _abc_15724_n5746;
  wire _abc_15724_n5747;
  wire _abc_15724_n5748;
  wire _abc_15724_n5749;
  wire _abc_15724_n5750;
  wire _abc_15724_n5751;
  wire _abc_15724_n5752;
  wire _abc_15724_n5753;
  wire _abc_15724_n5754;
  wire _abc_15724_n5755;
  wire _abc_15724_n5756;
  wire _abc_15724_n5757;
  wire _abc_15724_n5758;
  wire _abc_15724_n5759;
  wire _abc_15724_n5760;
  wire _abc_15724_n5761;
  wire _abc_15724_n5762;
  wire _abc_15724_n5763;
  wire _abc_15724_n5764;
  wire _abc_15724_n5765;
  wire _abc_15724_n5766;
  wire _abc_15724_n5767;
  wire _abc_15724_n5768;
  wire _abc_15724_n5769;
  wire _abc_15724_n5770;
  wire _abc_15724_n5772;
  wire _abc_15724_n5773;
  wire _abc_15724_n5774;
  wire _abc_15724_n5775;
  wire _abc_15724_n5776;
  wire _abc_15724_n5777;
  wire _abc_15724_n5778;
  wire _abc_15724_n5779;
  wire _abc_15724_n5780;
  wire _abc_15724_n5781;
  wire _abc_15724_n5782;
  wire _abc_15724_n5783;
  wire _abc_15724_n5784;
  wire _abc_15724_n5785;
  wire _abc_15724_n5786;
  wire _abc_15724_n5787;
  wire _abc_15724_n5788;
  wire _abc_15724_n5789;
  wire _abc_15724_n5790;
  wire _abc_15724_n5791;
  wire _abc_15724_n5792;
  wire _abc_15724_n5793;
  wire _abc_15724_n5794;
  wire _abc_15724_n5795;
  wire _abc_15724_n5796;
  wire _abc_15724_n5797;
  wire _abc_15724_n5798;
  wire _abc_15724_n5799;
  wire _abc_15724_n5800;
  wire _abc_15724_n5801;
  wire _abc_15724_n5802;
  wire _abc_15724_n5803;
  wire _abc_15724_n5804;
  wire _abc_15724_n5805;
  wire _abc_15724_n5806;
  wire _abc_15724_n5807;
  wire _abc_15724_n5808;
  wire _abc_15724_n5809;
  wire _abc_15724_n5810;
  wire _abc_15724_n5811;
  wire _abc_15724_n5812;
  wire _abc_15724_n5813;
  wire _abc_15724_n5814;
  wire _abc_15724_n5815;
  wire _abc_15724_n5816;
  wire _abc_15724_n5817;
  wire _abc_15724_n5818;
  wire _abc_15724_n5819;
  wire _abc_15724_n5820;
  wire _abc_15724_n5821;
  wire _abc_15724_n5822;
  wire _abc_15724_n5823;
  wire _abc_15724_n5824;
  wire _abc_15724_n5825;
  wire _abc_15724_n5826;
  wire _abc_15724_n5827;
  wire _abc_15724_n5828;
  wire _abc_15724_n5829;
  wire _abc_15724_n5830;
  wire _abc_15724_n5831;
  wire _abc_15724_n5832;
  wire _abc_15724_n5833;
  wire _abc_15724_n5834;
  wire _abc_15724_n5836;
  wire _abc_15724_n5837;
  wire _abc_15724_n5838;
  wire _abc_15724_n5839;
  wire _abc_15724_n5840;
  wire _abc_15724_n5841;
  wire _abc_15724_n5842;
  wire _abc_15724_n5843;
  wire _abc_15724_n5844;
  wire _abc_15724_n5845;
  wire _abc_15724_n5846;
  wire _abc_15724_n5847;
  wire _abc_15724_n5848;
  wire _abc_15724_n5849;
  wire _abc_15724_n5850;
  wire _abc_15724_n5851;
  wire _abc_15724_n5852;
  wire _abc_15724_n5853;
  wire _abc_15724_n5854;
  wire _abc_15724_n5855;
  wire _abc_15724_n5856;
  wire _abc_15724_n5857;
  wire _abc_15724_n5858;
  wire _abc_15724_n5859;
  wire _abc_15724_n5860;
  wire _abc_15724_n5861;
  wire _abc_15724_n5862;
  wire _abc_15724_n5863;
  wire _abc_15724_n5864;
  wire _abc_15724_n5865;
  wire _abc_15724_n5866;
  wire _abc_15724_n5867;
  wire _abc_15724_n5868;
  wire _abc_15724_n5869;
  wire _abc_15724_n5870;
  wire _abc_15724_n5871;
  wire _abc_15724_n5872;
  wire _abc_15724_n5873;
  wire _abc_15724_n5874;
  wire _abc_15724_n5875;
  wire _abc_15724_n5876;
  wire _abc_15724_n5877;
  wire _abc_15724_n5878;
  wire _abc_15724_n5879;
  wire _abc_15724_n5880;
  wire _abc_15724_n5881;
  wire _abc_15724_n5882;
  wire _abc_15724_n5883;
  wire _abc_15724_n5884;
  wire _abc_15724_n5885;
  wire _abc_15724_n5886;
  wire _abc_15724_n5887;
  wire _abc_15724_n5888;
  wire _abc_15724_n5889;
  wire _abc_15724_n5890;
  wire _abc_15724_n5891;
  wire _abc_15724_n5892;
  wire _abc_15724_n5893;
  wire _abc_15724_n5894;
  wire _abc_15724_n5895;
  wire _abc_15724_n5896;
  wire _abc_15724_n5897;
  wire _abc_15724_n5898;
  wire _abc_15724_n5899;
  wire _abc_15724_n5900;
  wire _abc_15724_n5901;
  wire _abc_15724_n5902;
  wire _abc_15724_n5903;
  wire _abc_15724_n5904;
  wire _abc_15724_n5905;
  wire _abc_15724_n5906;
  wire _abc_15724_n5907;
  wire _abc_15724_n5908;
  wire _abc_15724_n5909;
  wire _abc_15724_n5910;
  wire _abc_15724_n5912;
  wire _abc_15724_n5913;
  wire _abc_15724_n5914;
  wire _abc_15724_n5915;
  wire _abc_15724_n5916;
  wire _abc_15724_n5917;
  wire _abc_15724_n5918;
  wire _abc_15724_n5919;
  wire _abc_15724_n5920;
  wire _abc_15724_n5921;
  wire _abc_15724_n5922;
  wire _abc_15724_n5923;
  wire _abc_15724_n5924;
  wire _abc_15724_n5925;
  wire _abc_15724_n5926;
  wire _abc_15724_n5927;
  wire _abc_15724_n5928;
  wire _abc_15724_n5929;
  wire _abc_15724_n5930;
  wire _abc_15724_n5931;
  wire _abc_15724_n5932;
  wire _abc_15724_n5933;
  wire _abc_15724_n5934;
  wire _abc_15724_n5935;
  wire _abc_15724_n5936;
  wire _abc_15724_n5937;
  wire _abc_15724_n5938;
  wire _abc_15724_n5939;
  wire _abc_15724_n5940;
  wire _abc_15724_n5941;
  wire _abc_15724_n5942;
  wire _abc_15724_n5943;
  wire _abc_15724_n5944;
  wire _abc_15724_n5945;
  wire _abc_15724_n5946;
  wire _abc_15724_n5947;
  wire _abc_15724_n5948;
  wire _abc_15724_n5949;
  wire _abc_15724_n5950;
  wire _abc_15724_n5951;
  wire _abc_15724_n5952;
  wire _abc_15724_n5953;
  wire _abc_15724_n5954;
  wire _abc_15724_n5955;
  wire _abc_15724_n5956;
  wire _abc_15724_n5957;
  wire _abc_15724_n5958;
  wire _abc_15724_n5959;
  wire _abc_15724_n5960;
  wire _abc_15724_n5961;
  wire _abc_15724_n5962;
  wire _abc_15724_n5963;
  wire _abc_15724_n5964;
  wire _abc_15724_n5965;
  wire _abc_15724_n5966;
  wire _abc_15724_n5967;
  wire _abc_15724_n5968;
  wire _abc_15724_n5969;
  wire _abc_15724_n5970;
  wire _abc_15724_n5971;
  wire _abc_15724_n5972;
  wire _abc_15724_n5973;
  wire _abc_15724_n5974;
  wire _abc_15724_n5975;
  wire _abc_15724_n5976;
  wire _abc_15724_n5977;
  wire _abc_15724_n5978;
  wire _abc_15724_n5979;
  wire _abc_15724_n5980;
  wire _abc_15724_n5982;
  wire _abc_15724_n5983;
  wire _abc_15724_n5984;
  wire _abc_15724_n5985;
  wire _abc_15724_n5986;
  wire _abc_15724_n5987;
  wire _abc_15724_n5988;
  wire _abc_15724_n5989;
  wire _abc_15724_n5990;
  wire _abc_15724_n5991;
  wire _abc_15724_n5992;
  wire _abc_15724_n5993;
  wire _abc_15724_n5994;
  wire _abc_15724_n5995;
  wire _abc_15724_n5996;
  wire _abc_15724_n5997;
  wire _abc_15724_n5998;
  wire _abc_15724_n5999;
  wire _abc_15724_n6000;
  wire _abc_15724_n6001;
  wire _abc_15724_n6002;
  wire _abc_15724_n6003;
  wire _abc_15724_n6004;
  wire _abc_15724_n6005;
  wire _abc_15724_n6006;
  wire _abc_15724_n6007;
  wire _abc_15724_n6008;
  wire _abc_15724_n6009;
  wire _abc_15724_n6010;
  wire _abc_15724_n6011;
  wire _abc_15724_n6012;
  wire _abc_15724_n6013;
  wire _abc_15724_n6014;
  wire _abc_15724_n6015;
  wire _abc_15724_n6016;
  wire _abc_15724_n6017;
  wire _abc_15724_n6018;
  wire _abc_15724_n6019;
  wire _abc_15724_n6020;
  wire _abc_15724_n6021;
  wire _abc_15724_n6022;
  wire _abc_15724_n6023;
  wire _abc_15724_n6024;
  wire _abc_15724_n6025;
  wire _abc_15724_n6026;
  wire _abc_15724_n6027;
  wire _abc_15724_n6028;
  wire _abc_15724_n6029;
  wire _abc_15724_n6030;
  wire _abc_15724_n6031;
  wire _abc_15724_n6032;
  wire _abc_15724_n6033;
  wire _abc_15724_n6034;
  wire _abc_15724_n6035;
  wire _abc_15724_n6036;
  wire _abc_15724_n6037;
  wire _abc_15724_n6038;
  wire _abc_15724_n6039;
  wire _abc_15724_n6040;
  wire _abc_15724_n6041;
  wire _abc_15724_n6042;
  wire _abc_15724_n6043;
  wire _abc_15724_n6044;
  wire _abc_15724_n6045;
  wire _abc_15724_n6046;
  wire _abc_15724_n6047;
  wire _abc_15724_n6048;
  wire _abc_15724_n6050;
  wire _abc_15724_n6051;
  wire _abc_15724_n6052;
  wire _abc_15724_n6053;
  wire _abc_15724_n6054;
  wire _abc_15724_n6055;
  wire _abc_15724_n6056;
  wire _abc_15724_n6057;
  wire _abc_15724_n6058;
  wire _abc_15724_n6059;
  wire _abc_15724_n6060;
  wire _abc_15724_n6061;
  wire _abc_15724_n6062;
  wire _abc_15724_n6063;
  wire _abc_15724_n6064;
  wire _abc_15724_n6065;
  wire _abc_15724_n6066;
  wire _abc_15724_n6067;
  wire _abc_15724_n6068;
  wire _abc_15724_n6069;
  wire _abc_15724_n6070;
  wire _abc_15724_n6071;
  wire _abc_15724_n6072;
  wire _abc_15724_n6073;
  wire _abc_15724_n6074;
  wire _abc_15724_n6075;
  wire _abc_15724_n6076;
  wire _abc_15724_n6077;
  wire _abc_15724_n6078;
  wire _abc_15724_n6079;
  wire _abc_15724_n6080;
  wire _abc_15724_n6081;
  wire _abc_15724_n6082;
  wire _abc_15724_n6083;
  wire _abc_15724_n6084;
  wire _abc_15724_n6085;
  wire _abc_15724_n6086;
  wire _abc_15724_n6087;
  wire _abc_15724_n6088;
  wire _abc_15724_n6089;
  wire _abc_15724_n6090;
  wire _abc_15724_n6091;
  wire _abc_15724_n6092;
  wire _abc_15724_n6093;
  wire _abc_15724_n6094;
  wire _abc_15724_n6095;
  wire _abc_15724_n6096;
  wire _abc_15724_n6097;
  wire _abc_15724_n6098;
  wire _abc_15724_n6099;
  wire _abc_15724_n6100;
  wire _abc_15724_n6101;
  wire _abc_15724_n6102;
  wire _abc_15724_n6103;
  wire _abc_15724_n6104;
  wire _abc_15724_n6105;
  wire _abc_15724_n6106;
  wire _abc_15724_n6107;
  wire _abc_15724_n6108;
  wire _abc_15724_n6109;
  wire _abc_15724_n6110;
  wire _abc_15724_n6111;
  wire _abc_15724_n6112;
  wire _abc_15724_n6113;
  wire _abc_15724_n6114;
  wire _abc_15724_n6116;
  wire _abc_15724_n6117;
  wire _abc_15724_n6118;
  wire _abc_15724_n6119;
  wire _abc_15724_n6120;
  wire _abc_15724_n6121;
  wire _abc_15724_n6123;
  wire _abc_15724_n6124;
  wire _abc_15724_n6125;
  wire _abc_15724_n6126;
  wire _abc_15724_n6128;
  wire _abc_15724_n6129;
  wire _abc_15724_n6130;
  wire _abc_15724_n6132;
  wire _abc_15724_n6134;
  wire _abc_15724_n6135;
  wire _abc_15724_n6136;
  wire _abc_15724_n6138;
  wire _abc_15724_n6139;
  wire _abc_15724_n6140;
  wire _abc_15724_n6141;
  wire _abc_15724_n6142;
  wire _abc_15724_n6144;
  wire _abc_15724_n6145;
  wire _abc_15724_n6146;
  wire _abc_15724_n6147;
  wire _abc_15724_n6148;
  wire _abc_15724_n6149;
  wire _abc_15724_n6151;
  wire _abc_15724_n6152;
  wire _abc_15724_n6153;
  wire _abc_15724_n6154;
  wire _abc_15724_n6156;
  wire _abc_15724_n6157;
  wire _abc_15724_n6158;
  wire _abc_15724_n6159;
  wire _abc_15724_n6160;
  wire _abc_15724_n6162;
  wire _abc_15724_n6163;
  wire _abc_15724_n6164;
  wire _abc_15724_n6165;
  wire _abc_15724_n6166;
  wire _abc_15724_n6167;
  wire _abc_15724_n6169;
  wire _abc_15724_n6170;
  wire _abc_15724_n6171;
  wire _abc_15724_n6172;
  wire _abc_15724_n6173;
  wire _abc_15724_n6175;
  wire _abc_15724_n6176;
  wire _abc_15724_n6177;
  wire _abc_15724_n6178;
  wire _abc_15724_n6179;
  wire _abc_15724_n6181;
  wire _abc_15724_n6182;
  wire _abc_15724_n6183;
  wire _abc_15724_n6184;
  wire _abc_15724_n6186;
  wire _abc_15724_n6187;
  wire _abc_15724_n6188;
  wire _abc_15724_n6189;
  wire _abc_15724_n6190;
  wire _abc_15724_n6192;
  wire _abc_15724_n6193;
  wire _abc_15724_n6194;
  wire _abc_15724_n6195;
  wire _abc_15724_n6196;
  wire _abc_15724_n6197;
  wire _abc_15724_n6198;
  wire _abc_15724_n6199;
  wire _abc_15724_n6200;
  wire _abc_15724_n6202;
  wire _abc_15724_n6203;
  wire _abc_15724_n6204;
  wire _abc_15724_n6205;
  wire _abc_15724_n6206;
  wire _abc_15724_n6208;
  wire _abc_15724_n6209;
  wire _abc_15724_n6210;
  wire _abc_15724_n6211;
  wire _abc_15724_n6212;
  wire _abc_15724_n6213;
  wire _abc_15724_n6214;
  wire _abc_15724_n6215;
  wire _abc_15724_n6216;
  wire _abc_15724_n6218;
  wire _abc_15724_n6219;
  wire _abc_15724_n6220;
  wire _abc_15724_n6221;
  wire _abc_15724_n6222;
  wire _abc_15724_n6223;
  wire _abc_15724_n6225;
  wire _abc_15724_n6226;
  wire _abc_15724_n6227;
  wire _abc_15724_n6228;
  wire _abc_15724_n6229;
  wire _abc_15724_n6230;
  wire _abc_15724_n6231;
  wire _abc_15724_n6232;
  wire _abc_15724_n6234;
  wire _abc_15724_n6235;
  wire _abc_15724_n6236;
  wire _abc_15724_n6237;
  wire _abc_15724_n6238;
  wire _abc_15724_n6239;
  wire _abc_15724_n6241;
  wire _abc_15724_n6242;
  wire _abc_15724_n6243;
  wire _abc_15724_n6244;
  wire _abc_15724_n6245;
  wire _abc_15724_n6246;
  wire _abc_15724_n6247;
  wire _abc_15724_n6248;
  wire _abc_15724_n6250;
  wire _abc_15724_n6251;
  wire _abc_15724_n6252;
  wire _abc_15724_n6253;
  wire _abc_15724_n6254;
  wire _abc_15724_n6255;
  wire _abc_15724_n6256;
  wire _abc_15724_n6257;
  wire _abc_15724_n6259;
  wire _abc_15724_n6260;
  wire _abc_15724_n6261;
  wire _abc_15724_n6262;
  wire _abc_15724_n6263;
  wire _abc_15724_n6264;
  wire _abc_15724_n6265;
  wire _abc_15724_n6266;
  wire _abc_15724_n6268;
  wire _abc_15724_n6269;
  wire _abc_15724_n6270;
  wire _abc_15724_n6271;
  wire _abc_15724_n6272;
  wire _abc_15724_n6273;
  wire _abc_15724_n6275;
  wire _abc_15724_n6276;
  wire _abc_15724_n6277;
  wire _abc_15724_n6278;
  wire _abc_15724_n6279;
  wire _abc_15724_n6280;
  wire _abc_15724_n6281;
  wire _abc_15724_n6282;
  wire _abc_15724_n6284;
  wire _abc_15724_n6285;
  wire _abc_15724_n6286;
  wire _abc_15724_n6287;
  wire _abc_15724_n6288;
  wire _abc_15724_n6289;
  wire _abc_15724_n6290;
  wire _abc_15724_n6291;
  wire _abc_15724_n6293;
  wire _abc_15724_n6294;
  wire _abc_15724_n6295;
  wire _abc_15724_n6296;
  wire _abc_15724_n6297;
  wire _abc_15724_n6298;
  wire _abc_15724_n6299;
  wire _abc_15724_n6300;
  wire _abc_15724_n6302;
  wire _abc_15724_n6303;
  wire _abc_15724_n6304;
  wire _abc_15724_n6305;
  wire _abc_15724_n6306;
  wire _abc_15724_n6307;
  wire _abc_15724_n6309;
  wire _abc_15724_n6310;
  wire _abc_15724_n6311;
  wire _abc_15724_n6312;
  wire _abc_15724_n6313;
  wire _abc_15724_n6314;
  wire _abc_15724_n6315;
  wire _abc_15724_n6317;
  wire _abc_15724_n6318;
  wire _abc_15724_n6319;
  wire _abc_15724_n6320;
  wire _abc_15724_n6321;
  wire _abc_15724_n6322;
  wire _abc_15724_n6323;
  wire _abc_15724_n6324;
  wire _abc_15724_n6326;
  wire _abc_15724_n6327;
  wire _abc_15724_n6328;
  wire _abc_15724_n6329;
  wire _abc_15724_n6330;
  wire _abc_15724_n6331;
  wire _abc_15724_n6332;
  wire _abc_15724_n6333;
  wire _abc_15724_n6335;
  wire _abc_15724_n6336;
  wire _abc_15724_n6337;
  wire _abc_15724_n6338;
  wire _abc_15724_n6339;
  wire _abc_15724_n6340;
  wire _abc_15724_n6342;
  wire _abc_15724_n6343;
  wire _abc_15724_n6344;
  wire _abc_15724_n6345;
  wire _abc_15724_n6346;
  wire _abc_15724_n6347;
  wire _abc_15724_n6348;
  wire _abc_15724_n6349;
  wire _abc_15724_n698;
  wire _abc_15724_n699;
  wire _abc_15724_n700;
  wire _abc_15724_n701;
  wire _abc_15724_n702;
  wire _abc_15724_n703;
  wire _abc_15724_n704;
  wire _abc_15724_n705;
  wire _abc_15724_n706;
  wire _abc_15724_n707;
  wire _abc_15724_n708_1;
  wire _abc_15724_n709_1;
  wire _abc_15724_n710_1;
  wire _abc_15724_n711;
  wire _abc_15724_n712;
  wire _abc_15724_n713;
  wire _abc_15724_n714;
  wire _abc_15724_n715;
  wire _abc_15724_n716;
  wire _abc_15724_n717;
  wire _abc_15724_n718_1;
  wire _abc_15724_n719_1;
  wire _abc_15724_n720;
  wire _abc_15724_n721_1;
  wire _abc_15724_n722;
  wire _abc_15724_n723;
  wire _abc_15724_n724;
  wire _abc_15724_n725;
  wire _abc_15724_n726;
  wire _abc_15724_n727;
  wire _abc_15724_n728;
  wire _abc_15724_n729_1;
  wire _abc_15724_n730_1;
  wire _abc_15724_n731_1;
  wire _abc_15724_n732;
  wire _abc_15724_n733;
  wire _abc_15724_n734;
  wire _abc_15724_n735;
  wire _abc_15724_n736;
  wire _abc_15724_n737;
  wire _abc_15724_n738_1;
  wire _abc_15724_n739_1;
  wire _abc_15724_n740;
  wire _abc_15724_n741_1;
  wire _abc_15724_n742;
  wire _abc_15724_n743;
  wire _abc_15724_n744;
  wire _abc_15724_n745;
  wire _abc_15724_n746;
  wire _abc_15724_n747;
  wire _abc_15724_n748;
  wire _abc_15724_n749;
  wire _abc_15724_n750;
  wire _abc_15724_n751;
  wire _abc_15724_n752;
  wire _abc_15724_n753;
  wire _abc_15724_n754;
  wire _abc_15724_n755;
  wire _abc_15724_n756;
  wire _abc_15724_n757_1;
  wire _abc_15724_n758_1;
  wire _abc_15724_n759;
  wire _abc_15724_n760_1;
  wire _abc_15724_n761;
  wire _abc_15724_n762;
  wire _abc_15724_n763;
  wire _abc_15724_n764;
  wire _abc_15724_n765;
  wire _abc_15724_n766_1;
  wire _abc_15724_n767_1;
  wire _abc_15724_n768;
  wire _abc_15724_n769_1;
  wire _abc_15724_n770;
  wire _abc_15724_n771;
  wire _abc_15724_n772;
  wire _abc_15724_n773;
  wire _abc_15724_n774;
  wire _abc_15724_n775;
  wire _abc_15724_n776;
  wire _abc_15724_n777;
  wire _abc_15724_n778;
  wire _abc_15724_n779_1;
  wire _abc_15724_n780_1;
  wire _abc_15724_n781_1;
  wire _abc_15724_n782;
  wire _abc_15724_n783;
  wire _abc_15724_n784;
  wire _abc_15724_n785;
  wire _abc_15724_n786;
  wire _abc_15724_n787;
  wire _abc_15724_n788;
  wire _abc_15724_n789_1;
  wire _abc_15724_n790_1;
  wire _abc_15724_n791_1;
  wire _abc_15724_n792;
  wire _abc_15724_n793;
  wire _abc_15724_n794;
  wire _abc_15724_n795;
  wire _abc_15724_n796;
  wire _abc_15724_n797;
  wire _abc_15724_n798;
  wire _abc_15724_n799;
  wire _abc_15724_n800;
  wire _abc_15724_n801;
  wire _abc_15724_n802;
  wire _abc_15724_n803_1;
  wire _abc_15724_n804_1;
  wire _abc_15724_n805;
  wire _abc_15724_n806_1;
  wire _abc_15724_n807;
  wire _abc_15724_n808;
  wire _abc_15724_n809;
  wire _abc_15724_n810;
  wire _abc_15724_n811;
  wire _abc_15724_n812_1;
  wire _abc_15724_n813_1;
  wire _abc_15724_n814;
  wire _abc_15724_n815_1;
  wire _abc_15724_n816;
  wire _abc_15724_n817;
  wire _abc_15724_n818;
  wire _abc_15724_n819;
  wire _abc_15724_n820;
  wire _abc_15724_n821;
  wire _abc_15724_n822;
  wire _abc_15724_n823;
  wire _abc_15724_n824_1;
  wire _abc_15724_n825_1;
  wire _abc_15724_n826_1;
  wire _abc_15724_n827;
  wire _abc_15724_n828;
  wire _abc_15724_n829;
  wire _abc_15724_n830;
  wire _abc_15724_n831;
  wire _abc_15724_n832_1;
  wire _abc_15724_n833_1;
  wire _abc_15724_n834_1;
  wire _abc_15724_n835;
  wire _abc_15724_n836;
  wire _abc_15724_n837_1;
  wire _abc_15724_n838_1;
  wire _abc_15724_n839;
  wire _abc_15724_n840_1;
  wire _abc_15724_n841;
  wire _abc_15724_n842;
  wire _abc_15724_n843;
  wire _abc_15724_n844_1;
  wire _abc_15724_n845_1;
  wire _abc_15724_n846;
  wire _abc_15724_n847_1;
  wire _abc_15724_n848;
  wire _abc_15724_n849;
  wire _abc_15724_n850;
  wire _abc_15724_n850_bF_buf0;
  wire _abc_15724_n850_bF_buf1;
  wire _abc_15724_n850_bF_buf2;
  wire _abc_15724_n850_bF_buf3;
  wire _abc_15724_n850_bF_buf4;
  wire _abc_15724_n850_bF_buf5;
  wire _abc_15724_n850_bF_buf6;
  wire _abc_15724_n850_bF_buf7;
  wire _abc_15724_n850_bF_buf8;
  wire _abc_15724_n851;
  wire _abc_15724_n851_bF_buf0;
  wire _abc_15724_n851_bF_buf1;
  wire _abc_15724_n851_bF_buf2;
  wire _abc_15724_n851_bF_buf3;
  wire _abc_15724_n851_bF_buf4;
  wire _abc_15724_n851_bF_buf5;
  wire _abc_15724_n851_bF_buf6;
  wire _abc_15724_n851_bF_buf7;
  wire _abc_15724_n851_bF_buf8;
  wire _abc_15724_n852;
  wire _abc_15724_n853_1;
  wire _abc_15724_n855_1;
  wire _abc_15724_n856;
  wire _abc_15724_n857;
  wire _abc_15724_n858;
  wire _abc_15724_n859;
  wire _abc_15724_n860;
  wire _abc_15724_n861;
  wire _abc_15724_n862;
  wire _abc_15724_n863_1;
  wire _abc_15724_n864_1;
  wire _abc_15724_n865;
  wire _abc_15724_n866_1;
  wire _abc_15724_n867;
  wire _abc_15724_n869;
  wire _abc_15724_n870;
  wire _abc_15724_n871;
  wire _abc_15724_n872;
  wire _abc_15724_n873;
  wire _abc_15724_n874;
  wire _abc_15724_n875_1;
  wire _abc_15724_n876_1;
  wire _abc_15724_n877;
  wire _abc_15724_n878_1;
  wire _abc_15724_n879;
  wire _abc_15724_n880;
  wire _abc_15724_n881;
  wire _abc_15724_n882;
  wire _abc_15724_n883;
  wire _abc_15724_n884_1;
  wire _abc_15724_n885_1;
  wire _abc_15724_n886;
  wire _abc_15724_n887_1;
  wire _abc_15724_n888;
  wire _abc_15724_n889;
  wire _abc_15724_n890;
  wire _abc_15724_n892;
  wire _abc_15724_n893;
  wire _abc_15724_n894;
  wire _abc_15724_n895;
  wire _abc_15724_n896;
  wire _abc_15724_n897_1;
  wire _abc_15724_n898_1;
  wire _abc_15724_n899_1;
  wire _abc_15724_n900;
  wire _abc_15724_n901;
  wire _abc_15724_n902;
  wire _abc_15724_n903;
  wire _abc_15724_n904;
  wire _abc_15724_n906;
  wire _abc_15724_n906_bF_buf0;
  wire _abc_15724_n906_bF_buf1;
  wire _abc_15724_n906_bF_buf2;
  wire _abc_15724_n906_bF_buf3;
  wire _abc_15724_n906_bF_buf4;
  wire _abc_15724_n906_bF_buf5;
  wire _abc_15724_n906_bF_buf6;
  wire _abc_15724_n906_bF_buf7;
  wire _abc_15724_n906_bF_buf8;
  wire _abc_15724_n907_1;
  wire _abc_15724_n907_1_bF_buf0;
  wire _abc_15724_n907_1_bF_buf1;
  wire _abc_15724_n907_1_bF_buf2;
  wire _abc_15724_n907_1_bF_buf3;
  wire _abc_15724_n907_1_bF_buf4;
  wire _abc_15724_n907_1_bF_buf5;
  wire _abc_15724_n907_1_bF_buf6;
  wire _abc_15724_n907_1_bF_buf7;
  wire _abc_15724_n908_1;
  wire _abc_15724_n909_1;
  wire _abc_15724_n910;
  wire _abc_15724_n911;
  wire _abc_15724_n912;
  wire _abc_15724_n913;
  wire _abc_15724_n914;
  wire _abc_15724_n915;
  wire _abc_15724_n916;
  wire _abc_15724_n917;
  wire _abc_15724_n918;
  wire _abc_15724_n919;
  wire _abc_15724_n920;
  wire _abc_15724_n921_1;
  wire _abc_15724_n922_1;
  wire _abc_15724_n924;
  wire _abc_15724_n925;
  wire _abc_15724_n926;
  wire _abc_15724_n927;
  wire _abc_15724_n928;
  wire _abc_15724_n929;
  wire _abc_15724_n930;
  wire _abc_15724_n931_1;
  wire _abc_15724_n932_1;
  wire _abc_15724_n933;
  wire _abc_15724_n934_1;
  wire _abc_15724_n935;
  wire _abc_15724_n936;
  wire _abc_15724_n937;
  wire _abc_15724_n938;
  wire _abc_15724_n940;
  wire _abc_15724_n941;
  wire _abc_15724_n942;
  wire _abc_15724_n943_1;
  wire _abc_15724_n944_1;
  wire _abc_15724_n945_1;
  wire _abc_15724_n946;
  wire _abc_15724_n947;
  wire _abc_15724_n948;
  wire _abc_15724_n949;
  wire _abc_15724_n950;
  wire _abc_15724_n951;
  wire _abc_15724_n952;
  wire _abc_15724_n954_1;
  wire _abc_15724_n955;
  wire _abc_15724_n956_1;
  wire _abc_15724_n957;
  wire _abc_15724_n958;
  wire _abc_15724_n959;
  wire _abc_15724_n960;
  wire _abc_15724_n961;
  wire _abc_15724_n962;
  wire _abc_15724_n963;
  wire _abc_15724_n964;
  wire _abc_15724_n965;
  wire _abc_15724_n966_1;
  wire _abc_15724_n968_1;
  wire _abc_15724_n969;
  wire _abc_15724_n970;
  wire _abc_15724_n971;
  wire _abc_15724_n972;
  wire _abc_15724_n973;
  wire _abc_15724_n974;
  wire _abc_15724_n975;
  wire _abc_15724_n976_1;
  wire _abc_15724_n977_1;
  wire _abc_15724_n978;
  wire _abc_15724_n979_1;
  wire _abc_15724_n980;
  wire _abc_15724_n981;
  wire _abc_15724_n982;
  wire _abc_15724_n983;
  wire _abc_15724_n985;
  wire _abc_15724_n986;
  wire _abc_15724_n987_1;
  wire _abc_15724_n988_1;
  wire _abc_15724_n989_1;
  wire _abc_15724_n990;
  wire _abc_15724_n991;
  wire _abc_15724_n992;
  wire _abc_15724_n993;
  wire _abc_15724_n994;
  wire _abc_15724_n995;
  wire _abc_15724_n996_1;
  wire _abc_15724_n997_1;
  wire _abc_15724_n998_1;
  wire _auto_iopadmap_cc_313_execute_26059_0_;
  wire _auto_iopadmap_cc_313_execute_26059_100_;
  wire _auto_iopadmap_cc_313_execute_26059_101_;
  wire _auto_iopadmap_cc_313_execute_26059_102_;
  wire _auto_iopadmap_cc_313_execute_26059_103_;
  wire _auto_iopadmap_cc_313_execute_26059_104_;
  wire _auto_iopadmap_cc_313_execute_26059_105_;
  wire _auto_iopadmap_cc_313_execute_26059_106_;
  wire _auto_iopadmap_cc_313_execute_26059_107_;
  wire _auto_iopadmap_cc_313_execute_26059_108_;
  wire _auto_iopadmap_cc_313_execute_26059_109_;
  wire _auto_iopadmap_cc_313_execute_26059_10_;
  wire _auto_iopadmap_cc_313_execute_26059_110_;
  wire _auto_iopadmap_cc_313_execute_26059_111_;
  wire _auto_iopadmap_cc_313_execute_26059_112_;
  wire _auto_iopadmap_cc_313_execute_26059_113_;
  wire _auto_iopadmap_cc_313_execute_26059_114_;
  wire _auto_iopadmap_cc_313_execute_26059_115_;
  wire _auto_iopadmap_cc_313_execute_26059_116_;
  wire _auto_iopadmap_cc_313_execute_26059_117_;
  wire _auto_iopadmap_cc_313_execute_26059_118_;
  wire _auto_iopadmap_cc_313_execute_26059_119_;
  wire _auto_iopadmap_cc_313_execute_26059_11_;
  wire _auto_iopadmap_cc_313_execute_26059_120_;
  wire _auto_iopadmap_cc_313_execute_26059_121_;
  wire _auto_iopadmap_cc_313_execute_26059_122_;
  wire _auto_iopadmap_cc_313_execute_26059_123_;
  wire _auto_iopadmap_cc_313_execute_26059_124_;
  wire _auto_iopadmap_cc_313_execute_26059_125_;
  wire _auto_iopadmap_cc_313_execute_26059_126_;
  wire _auto_iopadmap_cc_313_execute_26059_127_;
  wire _auto_iopadmap_cc_313_execute_26059_128_;
  wire _auto_iopadmap_cc_313_execute_26059_129_;
  wire _auto_iopadmap_cc_313_execute_26059_12_;
  wire _auto_iopadmap_cc_313_execute_26059_130_;
  wire _auto_iopadmap_cc_313_execute_26059_131_;
  wire _auto_iopadmap_cc_313_execute_26059_132_;
  wire _auto_iopadmap_cc_313_execute_26059_133_;
  wire _auto_iopadmap_cc_313_execute_26059_134_;
  wire _auto_iopadmap_cc_313_execute_26059_135_;
  wire _auto_iopadmap_cc_313_execute_26059_136_;
  wire _auto_iopadmap_cc_313_execute_26059_137_;
  wire _auto_iopadmap_cc_313_execute_26059_138_;
  wire _auto_iopadmap_cc_313_execute_26059_139_;
  wire _auto_iopadmap_cc_313_execute_26059_13_;
  wire _auto_iopadmap_cc_313_execute_26059_140_;
  wire _auto_iopadmap_cc_313_execute_26059_141_;
  wire _auto_iopadmap_cc_313_execute_26059_142_;
  wire _auto_iopadmap_cc_313_execute_26059_143_;
  wire _auto_iopadmap_cc_313_execute_26059_144_;
  wire _auto_iopadmap_cc_313_execute_26059_145_;
  wire _auto_iopadmap_cc_313_execute_26059_146_;
  wire _auto_iopadmap_cc_313_execute_26059_147_;
  wire _auto_iopadmap_cc_313_execute_26059_148_;
  wire _auto_iopadmap_cc_313_execute_26059_149_;
  wire _auto_iopadmap_cc_313_execute_26059_14_;
  wire _auto_iopadmap_cc_313_execute_26059_150_;
  wire _auto_iopadmap_cc_313_execute_26059_151_;
  wire _auto_iopadmap_cc_313_execute_26059_152_;
  wire _auto_iopadmap_cc_313_execute_26059_153_;
  wire _auto_iopadmap_cc_313_execute_26059_154_;
  wire _auto_iopadmap_cc_313_execute_26059_155_;
  wire _auto_iopadmap_cc_313_execute_26059_156_;
  wire _auto_iopadmap_cc_313_execute_26059_157_;
  wire _auto_iopadmap_cc_313_execute_26059_158_;
  wire _auto_iopadmap_cc_313_execute_26059_159_;
  wire _auto_iopadmap_cc_313_execute_26059_15_;
  wire _auto_iopadmap_cc_313_execute_26059_16_;
  wire _auto_iopadmap_cc_313_execute_26059_17_;
  wire _auto_iopadmap_cc_313_execute_26059_18_;
  wire _auto_iopadmap_cc_313_execute_26059_19_;
  wire _auto_iopadmap_cc_313_execute_26059_1_;
  wire _auto_iopadmap_cc_313_execute_26059_20_;
  wire _auto_iopadmap_cc_313_execute_26059_21_;
  wire _auto_iopadmap_cc_313_execute_26059_22_;
  wire _auto_iopadmap_cc_313_execute_26059_23_;
  wire _auto_iopadmap_cc_313_execute_26059_24_;
  wire _auto_iopadmap_cc_313_execute_26059_25_;
  wire _auto_iopadmap_cc_313_execute_26059_26_;
  wire _auto_iopadmap_cc_313_execute_26059_27_;
  wire _auto_iopadmap_cc_313_execute_26059_28_;
  wire _auto_iopadmap_cc_313_execute_26059_29_;
  wire _auto_iopadmap_cc_313_execute_26059_2_;
  wire _auto_iopadmap_cc_313_execute_26059_30_;
  wire _auto_iopadmap_cc_313_execute_26059_31_;
  wire _auto_iopadmap_cc_313_execute_26059_32_;
  wire _auto_iopadmap_cc_313_execute_26059_33_;
  wire _auto_iopadmap_cc_313_execute_26059_34_;
  wire _auto_iopadmap_cc_313_execute_26059_35_;
  wire _auto_iopadmap_cc_313_execute_26059_36_;
  wire _auto_iopadmap_cc_313_execute_26059_37_;
  wire _auto_iopadmap_cc_313_execute_26059_38_;
  wire _auto_iopadmap_cc_313_execute_26059_39_;
  wire _auto_iopadmap_cc_313_execute_26059_3_;
  wire _auto_iopadmap_cc_313_execute_26059_40_;
  wire _auto_iopadmap_cc_313_execute_26059_41_;
  wire _auto_iopadmap_cc_313_execute_26059_42_;
  wire _auto_iopadmap_cc_313_execute_26059_43_;
  wire _auto_iopadmap_cc_313_execute_26059_44_;
  wire _auto_iopadmap_cc_313_execute_26059_45_;
  wire _auto_iopadmap_cc_313_execute_26059_46_;
  wire _auto_iopadmap_cc_313_execute_26059_47_;
  wire _auto_iopadmap_cc_313_execute_26059_48_;
  wire _auto_iopadmap_cc_313_execute_26059_49_;
  wire _auto_iopadmap_cc_313_execute_26059_4_;
  wire _auto_iopadmap_cc_313_execute_26059_50_;
  wire _auto_iopadmap_cc_313_execute_26059_51_;
  wire _auto_iopadmap_cc_313_execute_26059_52_;
  wire _auto_iopadmap_cc_313_execute_26059_53_;
  wire _auto_iopadmap_cc_313_execute_26059_54_;
  wire _auto_iopadmap_cc_313_execute_26059_55_;
  wire _auto_iopadmap_cc_313_execute_26059_56_;
  wire _auto_iopadmap_cc_313_execute_26059_57_;
  wire _auto_iopadmap_cc_313_execute_26059_58_;
  wire _auto_iopadmap_cc_313_execute_26059_59_;
  wire _auto_iopadmap_cc_313_execute_26059_5_;
  wire _auto_iopadmap_cc_313_execute_26059_60_;
  wire _auto_iopadmap_cc_313_execute_26059_61_;
  wire _auto_iopadmap_cc_313_execute_26059_62_;
  wire _auto_iopadmap_cc_313_execute_26059_63_;
  wire _auto_iopadmap_cc_313_execute_26059_64_;
  wire _auto_iopadmap_cc_313_execute_26059_65_;
  wire _auto_iopadmap_cc_313_execute_26059_66_;
  wire _auto_iopadmap_cc_313_execute_26059_67_;
  wire _auto_iopadmap_cc_313_execute_26059_68_;
  wire _auto_iopadmap_cc_313_execute_26059_69_;
  wire _auto_iopadmap_cc_313_execute_26059_6_;
  wire _auto_iopadmap_cc_313_execute_26059_70_;
  wire _auto_iopadmap_cc_313_execute_26059_71_;
  wire _auto_iopadmap_cc_313_execute_26059_72_;
  wire _auto_iopadmap_cc_313_execute_26059_73_;
  wire _auto_iopadmap_cc_313_execute_26059_74_;
  wire _auto_iopadmap_cc_313_execute_26059_75_;
  wire _auto_iopadmap_cc_313_execute_26059_76_;
  wire _auto_iopadmap_cc_313_execute_26059_77_;
  wire _auto_iopadmap_cc_313_execute_26059_78_;
  wire _auto_iopadmap_cc_313_execute_26059_79_;
  wire _auto_iopadmap_cc_313_execute_26059_7_;
  wire _auto_iopadmap_cc_313_execute_26059_80_;
  wire _auto_iopadmap_cc_313_execute_26059_81_;
  wire _auto_iopadmap_cc_313_execute_26059_82_;
  wire _auto_iopadmap_cc_313_execute_26059_83_;
  wire _auto_iopadmap_cc_313_execute_26059_84_;
  wire _auto_iopadmap_cc_313_execute_26059_85_;
  wire _auto_iopadmap_cc_313_execute_26059_86_;
  wire _auto_iopadmap_cc_313_execute_26059_87_;
  wire _auto_iopadmap_cc_313_execute_26059_88_;
  wire _auto_iopadmap_cc_313_execute_26059_89_;
  wire _auto_iopadmap_cc_313_execute_26059_8_;
  wire _auto_iopadmap_cc_313_execute_26059_90_;
  wire _auto_iopadmap_cc_313_execute_26059_91_;
  wire _auto_iopadmap_cc_313_execute_26059_92_;
  wire _auto_iopadmap_cc_313_execute_26059_93_;
  wire _auto_iopadmap_cc_313_execute_26059_94_;
  wire _auto_iopadmap_cc_313_execute_26059_95_;
  wire _auto_iopadmap_cc_313_execute_26059_96_;
  wire _auto_iopadmap_cc_313_execute_26059_97_;
  wire _auto_iopadmap_cc_313_execute_26059_98_;
  wire _auto_iopadmap_cc_313_execute_26059_99_;
  wire _auto_iopadmap_cc_313_execute_26059_9_;
  wire _auto_iopadmap_cc_313_execute_26220;
  wire _auto_iopadmap_cc_313_execute_26222;
  wire a_reg_0_;
  wire a_reg_0__FF_INPUT;
  wire a_reg_10_;
  wire a_reg_10__FF_INPUT;
  wire a_reg_11_;
  wire a_reg_11__FF_INPUT;
  wire a_reg_12_;
  wire a_reg_12__FF_INPUT;
  wire a_reg_13_;
  wire a_reg_13__FF_INPUT;
  wire a_reg_14_;
  wire a_reg_14__FF_INPUT;
  wire a_reg_15_;
  wire a_reg_15__FF_INPUT;
  wire a_reg_16_;
  wire a_reg_16__FF_INPUT;
  wire a_reg_17_;
  wire a_reg_17__FF_INPUT;
  wire a_reg_18_;
  wire a_reg_18__FF_INPUT;
  wire a_reg_19_;
  wire a_reg_19__FF_INPUT;
  wire a_reg_1_;
  wire a_reg_1__FF_INPUT;
  wire a_reg_20_;
  wire a_reg_20__FF_INPUT;
  wire a_reg_21_;
  wire a_reg_21__FF_INPUT;
  wire a_reg_22_;
  wire a_reg_22__FF_INPUT;
  wire a_reg_23_;
  wire a_reg_23__FF_INPUT;
  wire a_reg_24_;
  wire a_reg_24__FF_INPUT;
  wire a_reg_25_;
  wire a_reg_25__FF_INPUT;
  wire a_reg_26_;
  wire a_reg_26__FF_INPUT;
  wire a_reg_27_;
  wire a_reg_27__FF_INPUT;
  wire a_reg_28_;
  wire a_reg_28__FF_INPUT;
  wire a_reg_29_;
  wire a_reg_29__FF_INPUT;
  wire a_reg_2_;
  wire a_reg_2__FF_INPUT;
  wire a_reg_30_;
  wire a_reg_30__FF_INPUT;
  wire a_reg_31_;
  wire a_reg_31__FF_INPUT;
  wire a_reg_3_;
  wire a_reg_3__FF_INPUT;
  wire a_reg_4_;
  wire a_reg_4__FF_INPUT;
  wire a_reg_5_;
  wire a_reg_5__FF_INPUT;
  wire a_reg_6_;
  wire a_reg_6__FF_INPUT;
  wire a_reg_7_;
  wire a_reg_7__FF_INPUT;
  wire a_reg_8_;
  wire a_reg_8__FF_INPUT;
  wire a_reg_9_;
  wire a_reg_9__FF_INPUT;
  wire b_reg_0_;
  wire b_reg_0__FF_INPUT;
  wire b_reg_10_;
  wire b_reg_10__FF_INPUT;
  wire b_reg_11_;
  wire b_reg_11__FF_INPUT;
  wire b_reg_12_;
  wire b_reg_12__FF_INPUT;
  wire b_reg_13_;
  wire b_reg_13__FF_INPUT;
  wire b_reg_14_;
  wire b_reg_14__FF_INPUT;
  wire b_reg_15_;
  wire b_reg_15__FF_INPUT;
  wire b_reg_16_;
  wire b_reg_16__FF_INPUT;
  wire b_reg_17_;
  wire b_reg_17__FF_INPUT;
  wire b_reg_18_;
  wire b_reg_18__FF_INPUT;
  wire b_reg_19_;
  wire b_reg_19__FF_INPUT;
  wire b_reg_1_;
  wire b_reg_1__FF_INPUT;
  wire b_reg_20_;
  wire b_reg_20__FF_INPUT;
  wire b_reg_21_;
  wire b_reg_21__FF_INPUT;
  wire b_reg_22_;
  wire b_reg_22__FF_INPUT;
  wire b_reg_23_;
  wire b_reg_23__FF_INPUT;
  wire b_reg_24_;
  wire b_reg_24__FF_INPUT;
  wire b_reg_25_;
  wire b_reg_25__FF_INPUT;
  wire b_reg_26_;
  wire b_reg_26__FF_INPUT;
  wire b_reg_27_;
  wire b_reg_27__FF_INPUT;
  wire b_reg_28_;
  wire b_reg_28__FF_INPUT;
  wire b_reg_29_;
  wire b_reg_29__FF_INPUT;
  wire b_reg_2_;
  wire b_reg_2__FF_INPUT;
  wire b_reg_30_;
  wire b_reg_30__FF_INPUT;
  wire b_reg_31_;
  wire b_reg_31__FF_INPUT;
  wire b_reg_3_;
  wire b_reg_3__FF_INPUT;
  wire b_reg_4_;
  wire b_reg_4__FF_INPUT;
  wire b_reg_5_;
  wire b_reg_5__FF_INPUT;
  wire b_reg_6_;
  wire b_reg_6__FF_INPUT;
  wire b_reg_7_;
  wire b_reg_7__FF_INPUT;
  wire b_reg_8_;
  wire b_reg_8__FF_INPUT;
  wire b_reg_9_;
  wire b_reg_9__FF_INPUT;
  input \block[0] ;
  input \block[100] ;
  input \block[101] ;
  input \block[102] ;
  input \block[103] ;
  input \block[104] ;
  input \block[105] ;
  input \block[106] ;
  input \block[107] ;
  input \block[108] ;
  input \block[109] ;
  input \block[10] ;
  input \block[110] ;
  input \block[111] ;
  input \block[112] ;
  input \block[113] ;
  input \block[114] ;
  input \block[115] ;
  input \block[116] ;
  input \block[117] ;
  input \block[118] ;
  input \block[119] ;
  input \block[11] ;
  input \block[120] ;
  input \block[121] ;
  input \block[122] ;
  input \block[123] ;
  input \block[124] ;
  input \block[125] ;
  input \block[126] ;
  input \block[127] ;
  input \block[128] ;
  input \block[129] ;
  input \block[12] ;
  input \block[130] ;
  input \block[131] ;
  input \block[132] ;
  input \block[133] ;
  input \block[134] ;
  input \block[135] ;
  input \block[136] ;
  input \block[137] ;
  input \block[138] ;
  input \block[139] ;
  input \block[13] ;
  input \block[140] ;
  input \block[141] ;
  input \block[142] ;
  input \block[143] ;
  input \block[144] ;
  input \block[145] ;
  input \block[146] ;
  input \block[147] ;
  input \block[148] ;
  input \block[149] ;
  input \block[14] ;
  input \block[150] ;
  input \block[151] ;
  input \block[152] ;
  input \block[153] ;
  input \block[154] ;
  input \block[155] ;
  input \block[156] ;
  input \block[157] ;
  input \block[158] ;
  input \block[159] ;
  input \block[15] ;
  input \block[160] ;
  input \block[161] ;
  input \block[162] ;
  input \block[163] ;
  input \block[164] ;
  input \block[165] ;
  input \block[166] ;
  input \block[167] ;
  input \block[168] ;
  input \block[169] ;
  input \block[16] ;
  input \block[170] ;
  input \block[171] ;
  input \block[172] ;
  input \block[173] ;
  input \block[174] ;
  input \block[175] ;
  input \block[176] ;
  input \block[177] ;
  input \block[178] ;
  input \block[179] ;
  input \block[17] ;
  input \block[180] ;
  input \block[181] ;
  input \block[182] ;
  input \block[183] ;
  input \block[184] ;
  input \block[185] ;
  input \block[186] ;
  input \block[187] ;
  input \block[188] ;
  input \block[189] ;
  input \block[18] ;
  input \block[190] ;
  input \block[191] ;
  input \block[192] ;
  input \block[193] ;
  input \block[194] ;
  input \block[195] ;
  input \block[196] ;
  input \block[197] ;
  input \block[198] ;
  input \block[199] ;
  input \block[19] ;
  input \block[1] ;
  input \block[200] ;
  input \block[201] ;
  input \block[202] ;
  input \block[203] ;
  input \block[204] ;
  input \block[205] ;
  input \block[206] ;
  input \block[207] ;
  input \block[208] ;
  input \block[209] ;
  input \block[20] ;
  input \block[210] ;
  input \block[211] ;
  input \block[212] ;
  input \block[213] ;
  input \block[214] ;
  input \block[215] ;
  input \block[216] ;
  input \block[217] ;
  input \block[218] ;
  input \block[219] ;
  input \block[21] ;
  input \block[220] ;
  input \block[221] ;
  input \block[222] ;
  input \block[223] ;
  input \block[224] ;
  input \block[225] ;
  input \block[226] ;
  input \block[227] ;
  input \block[228] ;
  input \block[229] ;
  input \block[22] ;
  input \block[230] ;
  input \block[231] ;
  input \block[232] ;
  input \block[233] ;
  input \block[234] ;
  input \block[235] ;
  input \block[236] ;
  input \block[237] ;
  input \block[238] ;
  input \block[239] ;
  input \block[23] ;
  input \block[240] ;
  input \block[241] ;
  input \block[242] ;
  input \block[243] ;
  input \block[244] ;
  input \block[245] ;
  input \block[246] ;
  input \block[247] ;
  input \block[248] ;
  input \block[249] ;
  input \block[24] ;
  input \block[250] ;
  input \block[251] ;
  input \block[252] ;
  input \block[253] ;
  input \block[254] ;
  input \block[255] ;
  input \block[256] ;
  input \block[257] ;
  input \block[258] ;
  input \block[259] ;
  input \block[25] ;
  input \block[260] ;
  input \block[261] ;
  input \block[262] ;
  input \block[263] ;
  input \block[264] ;
  input \block[265] ;
  input \block[266] ;
  input \block[267] ;
  input \block[268] ;
  input \block[269] ;
  input \block[26] ;
  input \block[270] ;
  input \block[271] ;
  input \block[272] ;
  input \block[273] ;
  input \block[274] ;
  input \block[275] ;
  input \block[276] ;
  input \block[277] ;
  input \block[278] ;
  input \block[279] ;
  input \block[27] ;
  input \block[280] ;
  input \block[281] ;
  input \block[282] ;
  input \block[283] ;
  input \block[284] ;
  input \block[285] ;
  input \block[286] ;
  input \block[287] ;
  input \block[288] ;
  input \block[289] ;
  input \block[28] ;
  input \block[290] ;
  input \block[291] ;
  input \block[292] ;
  input \block[293] ;
  input \block[294] ;
  input \block[295] ;
  input \block[296] ;
  input \block[297] ;
  input \block[298] ;
  input \block[299] ;
  input \block[29] ;
  input \block[2] ;
  input \block[300] ;
  input \block[301] ;
  input \block[302] ;
  input \block[303] ;
  input \block[304] ;
  input \block[305] ;
  input \block[306] ;
  input \block[307] ;
  input \block[308] ;
  input \block[309] ;
  input \block[30] ;
  input \block[310] ;
  input \block[311] ;
  input \block[312] ;
  input \block[313] ;
  input \block[314] ;
  input \block[315] ;
  input \block[316] ;
  input \block[317] ;
  input \block[318] ;
  input \block[319] ;
  input \block[31] ;
  input \block[320] ;
  input \block[321] ;
  input \block[322] ;
  input \block[323] ;
  input \block[324] ;
  input \block[325] ;
  input \block[326] ;
  input \block[327] ;
  input \block[328] ;
  input \block[329] ;
  input \block[32] ;
  input \block[330] ;
  input \block[331] ;
  input \block[332] ;
  input \block[333] ;
  input \block[334] ;
  input \block[335] ;
  input \block[336] ;
  input \block[337] ;
  input \block[338] ;
  input \block[339] ;
  input \block[33] ;
  input \block[340] ;
  input \block[341] ;
  input \block[342] ;
  input \block[343] ;
  input \block[344] ;
  input \block[345] ;
  input \block[346] ;
  input \block[347] ;
  input \block[348] ;
  input \block[349] ;
  input \block[34] ;
  input \block[350] ;
  input \block[351] ;
  input \block[352] ;
  input \block[353] ;
  input \block[354] ;
  input \block[355] ;
  input \block[356] ;
  input \block[357] ;
  input \block[358] ;
  input \block[359] ;
  input \block[35] ;
  input \block[360] ;
  input \block[361] ;
  input \block[362] ;
  input \block[363] ;
  input \block[364] ;
  input \block[365] ;
  input \block[366] ;
  input \block[367] ;
  input \block[368] ;
  input \block[369] ;
  input \block[36] ;
  input \block[370] ;
  input \block[371] ;
  input \block[372] ;
  input \block[373] ;
  input \block[374] ;
  input \block[375] ;
  input \block[376] ;
  input \block[377] ;
  input \block[378] ;
  input \block[379] ;
  input \block[37] ;
  input \block[380] ;
  input \block[381] ;
  input \block[382] ;
  input \block[383] ;
  input \block[384] ;
  input \block[385] ;
  input \block[386] ;
  input \block[387] ;
  input \block[388] ;
  input \block[389] ;
  input \block[38] ;
  input \block[390] ;
  input \block[391] ;
  input \block[392] ;
  input \block[393] ;
  input \block[394] ;
  input \block[395] ;
  input \block[396] ;
  input \block[397] ;
  input \block[398] ;
  input \block[399] ;
  input \block[39] ;
  input \block[3] ;
  input \block[400] ;
  input \block[401] ;
  input \block[402] ;
  input \block[403] ;
  input \block[404] ;
  input \block[405] ;
  input \block[406] ;
  input \block[407] ;
  input \block[408] ;
  input \block[409] ;
  input \block[40] ;
  input \block[410] ;
  input \block[411] ;
  input \block[412] ;
  input \block[413] ;
  input \block[414] ;
  input \block[415] ;
  input \block[416] ;
  input \block[417] ;
  input \block[418] ;
  input \block[419] ;
  input \block[41] ;
  input \block[420] ;
  input \block[421] ;
  input \block[422] ;
  input \block[423] ;
  input \block[424] ;
  input \block[425] ;
  input \block[426] ;
  input \block[427] ;
  input \block[428] ;
  input \block[429] ;
  input \block[42] ;
  input \block[430] ;
  input \block[431] ;
  input \block[432] ;
  input \block[433] ;
  input \block[434] ;
  input \block[435] ;
  input \block[436] ;
  input \block[437] ;
  input \block[438] ;
  input \block[439] ;
  input \block[43] ;
  input \block[440] ;
  input \block[441] ;
  input \block[442] ;
  input \block[443] ;
  input \block[444] ;
  input \block[445] ;
  input \block[446] ;
  input \block[447] ;
  input \block[448] ;
  input \block[449] ;
  input \block[44] ;
  input \block[450] ;
  input \block[451] ;
  input \block[452] ;
  input \block[453] ;
  input \block[454] ;
  input \block[455] ;
  input \block[456] ;
  input \block[457] ;
  input \block[458] ;
  input \block[459] ;
  input \block[45] ;
  input \block[460] ;
  input \block[461] ;
  input \block[462] ;
  input \block[463] ;
  input \block[464] ;
  input \block[465] ;
  input \block[466] ;
  input \block[467] ;
  input \block[468] ;
  input \block[469] ;
  input \block[46] ;
  input \block[470] ;
  input \block[471] ;
  input \block[472] ;
  input \block[473] ;
  input \block[474] ;
  input \block[475] ;
  input \block[476] ;
  input \block[477] ;
  input \block[478] ;
  input \block[479] ;
  input \block[47] ;
  input \block[480] ;
  input \block[481] ;
  input \block[482] ;
  input \block[483] ;
  input \block[484] ;
  input \block[485] ;
  input \block[486] ;
  input \block[487] ;
  input \block[488] ;
  input \block[489] ;
  input \block[48] ;
  input \block[490] ;
  input \block[491] ;
  input \block[492] ;
  input \block[493] ;
  input \block[494] ;
  input \block[495] ;
  input \block[496] ;
  input \block[497] ;
  input \block[498] ;
  input \block[499] ;
  input \block[49] ;
  input \block[4] ;
  input \block[500] ;
  input \block[501] ;
  input \block[502] ;
  input \block[503] ;
  input \block[504] ;
  input \block[505] ;
  input \block[506] ;
  input \block[507] ;
  input \block[508] ;
  input \block[509] ;
  input \block[50] ;
  input \block[510] ;
  input \block[511] ;
  input \block[51] ;
  input \block[52] ;
  input \block[53] ;
  input \block[54] ;
  input \block[55] ;
  input \block[56] ;
  input \block[57] ;
  input \block[58] ;
  input \block[59] ;
  input \block[5] ;
  input \block[60] ;
  input \block[61] ;
  input \block[62] ;
  input \block[63] ;
  input \block[64] ;
  input \block[65] ;
  input \block[66] ;
  input \block[67] ;
  input \block[68] ;
  input \block[69] ;
  input \block[6] ;
  input \block[70] ;
  input \block[71] ;
  input \block[72] ;
  input \block[73] ;
  input \block[74] ;
  input \block[75] ;
  input \block[76] ;
  input \block[77] ;
  input \block[78] ;
  input \block[79] ;
  input \block[7] ;
  input \block[80] ;
  input \block[81] ;
  input \block[82] ;
  input \block[83] ;
  input \block[84] ;
  input \block[85] ;
  input \block[86] ;
  input \block[87] ;
  input \block[88] ;
  input \block[89] ;
  input \block[8] ;
  input \block[90] ;
  input \block[91] ;
  input \block[92] ;
  input \block[93] ;
  input \block[94] ;
  input \block[95] ;
  input \block[96] ;
  input \block[97] ;
  input \block[98] ;
  input \block[99] ;
  input \block[9] ;
  wire c_reg_0_;
  wire c_reg_0__FF_INPUT;
  wire c_reg_10_;
  wire c_reg_10__FF_INPUT;
  wire c_reg_11_;
  wire c_reg_11__FF_INPUT;
  wire c_reg_12_;
  wire c_reg_12__FF_INPUT;
  wire c_reg_13_;
  wire c_reg_13__FF_INPUT;
  wire c_reg_14_;
  wire c_reg_14__FF_INPUT;
  wire c_reg_15_;
  wire c_reg_15__FF_INPUT;
  wire c_reg_16_;
  wire c_reg_16__FF_INPUT;
  wire c_reg_17_;
  wire c_reg_17__FF_INPUT;
  wire c_reg_18_;
  wire c_reg_18__FF_INPUT;
  wire c_reg_19_;
  wire c_reg_19__FF_INPUT;
  wire c_reg_1_;
  wire c_reg_1__FF_INPUT;
  wire c_reg_20_;
  wire c_reg_20__FF_INPUT;
  wire c_reg_21_;
  wire c_reg_21__FF_INPUT;
  wire c_reg_22_;
  wire c_reg_22__FF_INPUT;
  wire c_reg_23_;
  wire c_reg_23__FF_INPUT;
  wire c_reg_24_;
  wire c_reg_24__FF_INPUT;
  wire c_reg_25_;
  wire c_reg_25__FF_INPUT;
  wire c_reg_26_;
  wire c_reg_26__FF_INPUT;
  wire c_reg_27_;
  wire c_reg_27__FF_INPUT;
  wire c_reg_28_;
  wire c_reg_28__FF_INPUT;
  wire c_reg_29_;
  wire c_reg_29__FF_INPUT;
  wire c_reg_2_;
  wire c_reg_2__FF_INPUT;
  wire c_reg_30_;
  wire c_reg_30__FF_INPUT;
  wire c_reg_31_;
  wire c_reg_31__FF_INPUT;
  wire c_reg_3_;
  wire c_reg_3__FF_INPUT;
  wire c_reg_4_;
  wire c_reg_4__FF_INPUT;
  wire c_reg_5_;
  wire c_reg_5__FF_INPUT;
  wire c_reg_6_;
  wire c_reg_6__FF_INPUT;
  wire c_reg_7_;
  wire c_reg_7__FF_INPUT;
  wire c_reg_8_;
  wire c_reg_8__FF_INPUT;
  wire c_reg_9_;
  wire c_reg_9__FF_INPUT;
  input clk;
  wire clk_bF_buf0;
  wire clk_bF_buf1;
  wire clk_bF_buf10;
  wire clk_bF_buf11;
  wire clk_bF_buf12;
  wire clk_bF_buf13;
  wire clk_bF_buf14;
  wire clk_bF_buf15;
  wire clk_bF_buf16;
  wire clk_bF_buf17;
  wire clk_bF_buf18;
  wire clk_bF_buf19;
  wire clk_bF_buf2;
  wire clk_bF_buf20;
  wire clk_bF_buf21;
  wire clk_bF_buf22;
  wire clk_bF_buf23;
  wire clk_bF_buf24;
  wire clk_bF_buf25;
  wire clk_bF_buf26;
  wire clk_bF_buf27;
  wire clk_bF_buf28;
  wire clk_bF_buf29;
  wire clk_bF_buf3;
  wire clk_bF_buf30;
  wire clk_bF_buf31;
  wire clk_bF_buf32;
  wire clk_bF_buf33;
  wire clk_bF_buf34;
  wire clk_bF_buf35;
  wire clk_bF_buf36;
  wire clk_bF_buf37;
  wire clk_bF_buf38;
  wire clk_bF_buf39;
  wire clk_bF_buf4;
  wire clk_bF_buf40;
  wire clk_bF_buf41;
  wire clk_bF_buf42;
  wire clk_bF_buf43;
  wire clk_bF_buf44;
  wire clk_bF_buf45;
  wire clk_bF_buf46;
  wire clk_bF_buf47;
  wire clk_bF_buf48;
  wire clk_bF_buf49;
  wire clk_bF_buf5;
  wire clk_bF_buf50;
  wire clk_bF_buf51;
  wire clk_bF_buf52;
  wire clk_bF_buf53;
  wire clk_bF_buf54;
  wire clk_bF_buf55;
  wire clk_bF_buf56;
  wire clk_bF_buf57;
  wire clk_bF_buf58;
  wire clk_bF_buf59;
  wire clk_bF_buf6;
  wire clk_bF_buf60;
  wire clk_bF_buf61;
  wire clk_bF_buf62;
  wire clk_bF_buf63;
  wire clk_bF_buf64;
  wire clk_bF_buf65;
  wire clk_bF_buf66;
  wire clk_bF_buf67;
  wire clk_bF_buf68;
  wire clk_bF_buf69;
  wire clk_bF_buf7;
  wire clk_bF_buf70;
  wire clk_bF_buf71;
  wire clk_bF_buf72;
  wire clk_bF_buf73;
  wire clk_bF_buf74;
  wire clk_bF_buf75;
  wire clk_bF_buf76;
  wire clk_bF_buf77;
  wire clk_bF_buf78;
  wire clk_bF_buf79;
  wire clk_bF_buf8;
  wire clk_bF_buf80;
  wire clk_bF_buf81;
  wire clk_bF_buf82;
  wire clk_bF_buf83;
  wire clk_bF_buf84;
  wire clk_bF_buf85;
  wire clk_bF_buf86;
  wire clk_bF_buf87;
  wire clk_bF_buf88;
  wire clk_bF_buf9;
  wire clk_hier0_bF_buf0;
  wire clk_hier0_bF_buf1;
  wire clk_hier0_bF_buf2;
  wire clk_hier0_bF_buf3;
  wire clk_hier0_bF_buf4;
  wire clk_hier0_bF_buf5;
  wire clk_hier0_bF_buf6;
  wire clk_hier0_bF_buf7;
  wire clk_hier0_bF_buf8;
  wire d_reg_0_;
  wire d_reg_0__FF_INPUT;
  wire d_reg_10_;
  wire d_reg_10__FF_INPUT;
  wire d_reg_11_;
  wire d_reg_11__FF_INPUT;
  wire d_reg_12_;
  wire d_reg_12__FF_INPUT;
  wire d_reg_13_;
  wire d_reg_13__FF_INPUT;
  wire d_reg_14_;
  wire d_reg_14__FF_INPUT;
  wire d_reg_15_;
  wire d_reg_15__FF_INPUT;
  wire d_reg_16_;
  wire d_reg_16__FF_INPUT;
  wire d_reg_17_;
  wire d_reg_17__FF_INPUT;
  wire d_reg_18_;
  wire d_reg_18__FF_INPUT;
  wire d_reg_19_;
  wire d_reg_19__FF_INPUT;
  wire d_reg_1_;
  wire d_reg_1__FF_INPUT;
  wire d_reg_20_;
  wire d_reg_20__FF_INPUT;
  wire d_reg_21_;
  wire d_reg_21__FF_INPUT;
  wire d_reg_22_;
  wire d_reg_22__FF_INPUT;
  wire d_reg_23_;
  wire d_reg_23__FF_INPUT;
  wire d_reg_24_;
  wire d_reg_24__FF_INPUT;
  wire d_reg_25_;
  wire d_reg_25__FF_INPUT;
  wire d_reg_26_;
  wire d_reg_26__FF_INPUT;
  wire d_reg_27_;
  wire d_reg_27__FF_INPUT;
  wire d_reg_28_;
  wire d_reg_28__FF_INPUT;
  wire d_reg_29_;
  wire d_reg_29__FF_INPUT;
  wire d_reg_2_;
  wire d_reg_2__FF_INPUT;
  wire d_reg_30_;
  wire d_reg_30__FF_INPUT;
  wire d_reg_31_;
  wire d_reg_31__FF_INPUT;
  wire d_reg_3_;
  wire d_reg_3__FF_INPUT;
  wire d_reg_4_;
  wire d_reg_4__FF_INPUT;
  wire d_reg_5_;
  wire d_reg_5__FF_INPUT;
  wire d_reg_6_;
  wire d_reg_6__FF_INPUT;
  wire d_reg_7_;
  wire d_reg_7__FF_INPUT;
  wire d_reg_8_;
  wire d_reg_8__FF_INPUT;
  wire d_reg_9_;
  wire d_reg_9__FF_INPUT;
  output \digest[0] ;
  output \digest[100] ;
  output \digest[101] ;
  output \digest[102] ;
  output \digest[103] ;
  output \digest[104] ;
  output \digest[105] ;
  output \digest[106] ;
  output \digest[107] ;
  output \digest[108] ;
  output \digest[109] ;
  output \digest[10] ;
  output \digest[110] ;
  output \digest[111] ;
  output \digest[112] ;
  output \digest[113] ;
  output \digest[114] ;
  output \digest[115] ;
  output \digest[116] ;
  output \digest[117] ;
  output \digest[118] ;
  output \digest[119] ;
  output \digest[11] ;
  output \digest[120] ;
  output \digest[121] ;
  output \digest[122] ;
  output \digest[123] ;
  output \digest[124] ;
  output \digest[125] ;
  output \digest[126] ;
  output \digest[127] ;
  output \digest[128] ;
  output \digest[129] ;
  output \digest[12] ;
  output \digest[130] ;
  output \digest[131] ;
  output \digest[132] ;
  output \digest[133] ;
  output \digest[134] ;
  output \digest[135] ;
  output \digest[136] ;
  output \digest[137] ;
  output \digest[138] ;
  output \digest[139] ;
  output \digest[13] ;
  output \digest[140] ;
  output \digest[141] ;
  output \digest[142] ;
  output \digest[143] ;
  output \digest[144] ;
  output \digest[145] ;
  output \digest[146] ;
  output \digest[147] ;
  output \digest[148] ;
  output \digest[149] ;
  output \digest[14] ;
  output \digest[150] ;
  output \digest[151] ;
  output \digest[152] ;
  output \digest[153] ;
  output \digest[154] ;
  output \digest[155] ;
  output \digest[156] ;
  output \digest[157] ;
  output \digest[158] ;
  output \digest[159] ;
  output \digest[15] ;
  output \digest[16] ;
  output \digest[17] ;
  output \digest[18] ;
  output \digest[19] ;
  output \digest[1] ;
  output \digest[20] ;
  output \digest[21] ;
  output \digest[22] ;
  output \digest[23] ;
  output \digest[24] ;
  output \digest[25] ;
  output \digest[26] ;
  output \digest[27] ;
  output \digest[28] ;
  output \digest[29] ;
  output \digest[2] ;
  output \digest[30] ;
  output \digest[31] ;
  output \digest[32] ;
  output \digest[33] ;
  output \digest[34] ;
  output \digest[35] ;
  output \digest[36] ;
  output \digest[37] ;
  output \digest[38] ;
  output \digest[39] ;
  output \digest[3] ;
  output \digest[40] ;
  output \digest[41] ;
  output \digest[42] ;
  output \digest[43] ;
  output \digest[44] ;
  output \digest[45] ;
  output \digest[46] ;
  output \digest[47] ;
  output \digest[48] ;
  output \digest[49] ;
  output \digest[4] ;
  output \digest[50] ;
  output \digest[51] ;
  output \digest[52] ;
  output \digest[53] ;
  output \digest[54] ;
  output \digest[55] ;
  output \digest[56] ;
  output \digest[57] ;
  output \digest[58] ;
  output \digest[59] ;
  output \digest[5] ;
  output \digest[60] ;
  output \digest[61] ;
  output \digest[62] ;
  output \digest[63] ;
  output \digest[64] ;
  output \digest[65] ;
  output \digest[66] ;
  output \digest[67] ;
  output \digest[68] ;
  output \digest[69] ;
  output \digest[6] ;
  output \digest[70] ;
  output \digest[71] ;
  output \digest[72] ;
  output \digest[73] ;
  output \digest[74] ;
  output \digest[75] ;
  output \digest[76] ;
  output \digest[77] ;
  output \digest[78] ;
  output \digest[79] ;
  output \digest[7] ;
  output \digest[80] ;
  output \digest[81] ;
  output \digest[82] ;
  output \digest[83] ;
  output \digest[84] ;
  output \digest[85] ;
  output \digest[86] ;
  output \digest[87] ;
  output \digest[88] ;
  output \digest[89] ;
  output \digest[8] ;
  output \digest[90] ;
  output \digest[91] ;
  output \digest[92] ;
  output \digest[93] ;
  output \digest[94] ;
  output \digest[95] ;
  output \digest[96] ;
  output \digest[97] ;
  output \digest[98] ;
  output \digest[99] ;
  output \digest[9] ;
  wire digest_update;
  wire digest_update_bF_buf0;
  wire digest_update_bF_buf1;
  wire digest_update_bF_buf10;
  wire digest_update_bF_buf11;
  wire digest_update_bF_buf2;
  wire digest_update_bF_buf3;
  wire digest_update_bF_buf4;
  wire digest_update_bF_buf5;
  wire digest_update_bF_buf6;
  wire digest_update_bF_buf7;
  wire digest_update_bF_buf8;
  wire digest_update_bF_buf9;
  output digest_valid;
  wire digest_valid_reg_FF_INPUT;
  wire e_reg_0_;
  wire e_reg_0__FF_INPUT;
  wire e_reg_10_;
  wire e_reg_10__FF_INPUT;
  wire e_reg_11_;
  wire e_reg_11__FF_INPUT;
  wire e_reg_12_;
  wire e_reg_12__FF_INPUT;
  wire e_reg_13_;
  wire e_reg_13__FF_INPUT;
  wire e_reg_14_;
  wire e_reg_14__FF_INPUT;
  wire e_reg_15_;
  wire e_reg_15__FF_INPUT;
  wire e_reg_16_;
  wire e_reg_16__FF_INPUT;
  wire e_reg_17_;
  wire e_reg_17__FF_INPUT;
  wire e_reg_18_;
  wire e_reg_18__FF_INPUT;
  wire e_reg_19_;
  wire e_reg_19__FF_INPUT;
  wire e_reg_1_;
  wire e_reg_1__FF_INPUT;
  wire e_reg_20_;
  wire e_reg_20__FF_INPUT;
  wire e_reg_21_;
  wire e_reg_21__FF_INPUT;
  wire e_reg_22_;
  wire e_reg_22__FF_INPUT;
  wire e_reg_23_;
  wire e_reg_23__FF_INPUT;
  wire e_reg_24_;
  wire e_reg_24__FF_INPUT;
  wire e_reg_25_;
  wire e_reg_25__FF_INPUT;
  wire e_reg_26_;
  wire e_reg_26__FF_INPUT;
  wire e_reg_27_;
  wire e_reg_27__FF_INPUT;
  wire e_reg_28_;
  wire e_reg_28__FF_INPUT;
  wire e_reg_29_;
  wire e_reg_29__FF_INPUT;
  wire e_reg_2_;
  wire e_reg_2__FF_INPUT;
  wire e_reg_30_;
  wire e_reg_30__FF_INPUT;
  wire e_reg_31_;
  wire e_reg_31__FF_INPUT;
  wire e_reg_3_;
  wire e_reg_3__FF_INPUT;
  wire e_reg_4_;
  wire e_reg_4__FF_INPUT;
  wire e_reg_5_;
  wire e_reg_5__FF_INPUT;
  wire e_reg_6_;
  wire e_reg_6__FF_INPUT;
  wire e_reg_7_;
  wire e_reg_7__FF_INPUT;
  wire e_reg_8_;
  wire e_reg_8__FF_INPUT;
  wire e_reg_9_;
  wire e_reg_9__FF_INPUT;
  input init;
  input next;
  output ready;
  input reset_n;
  wire reset_n_bF_buf0;
  wire reset_n_bF_buf1;
  wire reset_n_bF_buf10;
  wire reset_n_bF_buf11;
  wire reset_n_bF_buf12;
  wire reset_n_bF_buf13;
  wire reset_n_bF_buf14;
  wire reset_n_bF_buf15;
  wire reset_n_bF_buf16;
  wire reset_n_bF_buf17;
  wire reset_n_bF_buf18;
  wire reset_n_bF_buf19;
  wire reset_n_bF_buf2;
  wire reset_n_bF_buf20;
  wire reset_n_bF_buf21;
  wire reset_n_bF_buf22;
  wire reset_n_bF_buf23;
  wire reset_n_bF_buf24;
  wire reset_n_bF_buf25;
  wire reset_n_bF_buf26;
  wire reset_n_bF_buf27;
  wire reset_n_bF_buf28;
  wire reset_n_bF_buf29;
  wire reset_n_bF_buf3;
  wire reset_n_bF_buf30;
  wire reset_n_bF_buf31;
  wire reset_n_bF_buf32;
  wire reset_n_bF_buf33;
  wire reset_n_bF_buf34;
  wire reset_n_bF_buf35;
  wire reset_n_bF_buf36;
  wire reset_n_bF_buf37;
  wire reset_n_bF_buf38;
  wire reset_n_bF_buf39;
  wire reset_n_bF_buf4;
  wire reset_n_bF_buf40;
  wire reset_n_bF_buf41;
  wire reset_n_bF_buf42;
  wire reset_n_bF_buf43;
  wire reset_n_bF_buf44;
  wire reset_n_bF_buf45;
  wire reset_n_bF_buf46;
  wire reset_n_bF_buf47;
  wire reset_n_bF_buf48;
  wire reset_n_bF_buf49;
  wire reset_n_bF_buf5;
  wire reset_n_bF_buf50;
  wire reset_n_bF_buf51;
  wire reset_n_bF_buf52;
  wire reset_n_bF_buf53;
  wire reset_n_bF_buf54;
  wire reset_n_bF_buf55;
  wire reset_n_bF_buf56;
  wire reset_n_bF_buf57;
  wire reset_n_bF_buf58;
  wire reset_n_bF_buf59;
  wire reset_n_bF_buf6;
  wire reset_n_bF_buf60;
  wire reset_n_bF_buf61;
  wire reset_n_bF_buf62;
  wire reset_n_bF_buf63;
  wire reset_n_bF_buf64;
  wire reset_n_bF_buf65;
  wire reset_n_bF_buf66;
  wire reset_n_bF_buf67;
  wire reset_n_bF_buf68;
  wire reset_n_bF_buf69;
  wire reset_n_bF_buf7;
  wire reset_n_bF_buf70;
  wire reset_n_bF_buf71;
  wire reset_n_bF_buf72;
  wire reset_n_bF_buf73;
  wire reset_n_bF_buf74;
  wire reset_n_bF_buf75;
  wire reset_n_bF_buf76;
  wire reset_n_bF_buf77;
  wire reset_n_bF_buf78;
  wire reset_n_bF_buf79;
  wire reset_n_bF_buf8;
  wire reset_n_bF_buf80;
  wire reset_n_bF_buf81;
  wire reset_n_bF_buf82;
  wire reset_n_bF_buf83;
  wire reset_n_bF_buf84;
  wire reset_n_bF_buf85;
  wire reset_n_bF_buf86;
  wire reset_n_bF_buf87;
  wire reset_n_bF_buf88;
  wire reset_n_bF_buf9;
  wire reset_n_hier0_bF_buf0;
  wire reset_n_hier0_bF_buf1;
  wire reset_n_hier0_bF_buf2;
  wire reset_n_hier0_bF_buf3;
  wire reset_n_hier0_bF_buf4;
  wire reset_n_hier0_bF_buf5;
  wire reset_n_hier0_bF_buf6;
  wire reset_n_hier0_bF_buf7;
  wire reset_n_hier0_bF_buf8;
  wire round_ctr_inc;
  wire round_ctr_inc_bF_buf0;
  wire round_ctr_inc_bF_buf1;
  wire round_ctr_inc_bF_buf10;
  wire round_ctr_inc_bF_buf11;
  wire round_ctr_inc_bF_buf12;
  wire round_ctr_inc_bF_buf2;
  wire round_ctr_inc_bF_buf3;
  wire round_ctr_inc_bF_buf4;
  wire round_ctr_inc_bF_buf5;
  wire round_ctr_inc_bF_buf6;
  wire round_ctr_inc_bF_buf7;
  wire round_ctr_inc_bF_buf8;
  wire round_ctr_inc_bF_buf9;
  wire round_ctr_reg_0_;
  wire round_ctr_reg_0__FF_INPUT;
  wire round_ctr_reg_1_;
  wire round_ctr_reg_1__FF_INPUT;
  wire round_ctr_reg_2_;
  wire round_ctr_reg_2__FF_INPUT;
  wire round_ctr_reg_3_;
  wire round_ctr_reg_3__FF_INPUT;
  wire round_ctr_reg_4_;
  wire round_ctr_reg_4__FF_INPUT;
  wire round_ctr_reg_5_;
  wire round_ctr_reg_5__FF_INPUT;
  wire round_ctr_reg_6_;
  wire round_ctr_reg_6__FF_INPUT;
  wire round_ctr_rst;
  wire round_ctr_rst_bF_buf0;
  wire round_ctr_rst_bF_buf1;
  wire round_ctr_rst_bF_buf10;
  wire round_ctr_rst_bF_buf11;
  wire round_ctr_rst_bF_buf12;
  wire round_ctr_rst_bF_buf13;
  wire round_ctr_rst_bF_buf14;
  wire round_ctr_rst_bF_buf15;
  wire round_ctr_rst_bF_buf16;
  wire round_ctr_rst_bF_buf17;
  wire round_ctr_rst_bF_buf18;
  wire round_ctr_rst_bF_buf19;
  wire round_ctr_rst_bF_buf2;
  wire round_ctr_rst_bF_buf20;
  wire round_ctr_rst_bF_buf21;
  wire round_ctr_rst_bF_buf22;
  wire round_ctr_rst_bF_buf23;
  wire round_ctr_rst_bF_buf24;
  wire round_ctr_rst_bF_buf25;
  wire round_ctr_rst_bF_buf26;
  wire round_ctr_rst_bF_buf27;
  wire round_ctr_rst_bF_buf28;
  wire round_ctr_rst_bF_buf29;
  wire round_ctr_rst_bF_buf3;
  wire round_ctr_rst_bF_buf30;
  wire round_ctr_rst_bF_buf31;
  wire round_ctr_rst_bF_buf32;
  wire round_ctr_rst_bF_buf33;
  wire round_ctr_rst_bF_buf34;
  wire round_ctr_rst_bF_buf35;
  wire round_ctr_rst_bF_buf36;
  wire round_ctr_rst_bF_buf37;
  wire round_ctr_rst_bF_buf38;
  wire round_ctr_rst_bF_buf39;
  wire round_ctr_rst_bF_buf4;
  wire round_ctr_rst_bF_buf40;
  wire round_ctr_rst_bF_buf41;
  wire round_ctr_rst_bF_buf42;
  wire round_ctr_rst_bF_buf43;
  wire round_ctr_rst_bF_buf44;
  wire round_ctr_rst_bF_buf45;
  wire round_ctr_rst_bF_buf46;
  wire round_ctr_rst_bF_buf47;
  wire round_ctr_rst_bF_buf48;
  wire round_ctr_rst_bF_buf49;
  wire round_ctr_rst_bF_buf5;
  wire round_ctr_rst_bF_buf50;
  wire round_ctr_rst_bF_buf51;
  wire round_ctr_rst_bF_buf52;
  wire round_ctr_rst_bF_buf53;
  wire round_ctr_rst_bF_buf54;
  wire round_ctr_rst_bF_buf55;
  wire round_ctr_rst_bF_buf56;
  wire round_ctr_rst_bF_buf57;
  wire round_ctr_rst_bF_buf58;
  wire round_ctr_rst_bF_buf59;
  wire round_ctr_rst_bF_buf6;
  wire round_ctr_rst_bF_buf60;
  wire round_ctr_rst_bF_buf61;
  wire round_ctr_rst_bF_buf62;
  wire round_ctr_rst_bF_buf63;
  wire round_ctr_rst_bF_buf7;
  wire round_ctr_rst_bF_buf8;
  wire round_ctr_rst_bF_buf9;
  wire round_ctr_rst_hier0_bF_buf0;
  wire round_ctr_rst_hier0_bF_buf1;
  wire round_ctr_rst_hier0_bF_buf2;
  wire round_ctr_rst_hier0_bF_buf3;
  wire round_ctr_rst_hier0_bF_buf4;
  wire round_ctr_rst_hier0_bF_buf5;
  wire round_ctr_rst_hier0_bF_buf6;
  wire round_ctr_rst_hier0_bF_buf7;
  wire w_0_;
  wire w_10_;
  wire w_11_;
  wire w_12_;
  wire w_13_;
  wire w_14_;
  wire w_15_;
  wire w_16_;
  wire w_17_;
  wire w_18_;
  wire w_19_;
  wire w_1_;
  wire w_20_;
  wire w_21_;
  wire w_22_;
  wire w_23_;
  wire w_24_;
  wire w_25_;
  wire w_26_;
  wire w_27_;
  wire w_28_;
  wire w_29_;
  wire w_2_;
  wire w_30_;
  wire w_31_;
  wire w_3_;
  wire w_4_;
  wire w_5_;
  wire w_6_;
  wire w_7_;
  wire w_8_;
  wire w_9_;
  wire w_mem_inst__0w_mem_0__31_0__0_;
  wire w_mem_inst__0w_mem_0__31_0__10_;
  wire w_mem_inst__0w_mem_0__31_0__11_;
  wire w_mem_inst__0w_mem_0__31_0__12_;
  wire w_mem_inst__0w_mem_0__31_0__13_;
  wire w_mem_inst__0w_mem_0__31_0__14_;
  wire w_mem_inst__0w_mem_0__31_0__15_;
  wire w_mem_inst__0w_mem_0__31_0__16_;
  wire w_mem_inst__0w_mem_0__31_0__17_;
  wire w_mem_inst__0w_mem_0__31_0__18_;
  wire w_mem_inst__0w_mem_0__31_0__19_;
  wire w_mem_inst__0w_mem_0__31_0__1_;
  wire w_mem_inst__0w_mem_0__31_0__20_;
  wire w_mem_inst__0w_mem_0__31_0__21_;
  wire w_mem_inst__0w_mem_0__31_0__22_;
  wire w_mem_inst__0w_mem_0__31_0__23_;
  wire w_mem_inst__0w_mem_0__31_0__24_;
  wire w_mem_inst__0w_mem_0__31_0__25_;
  wire w_mem_inst__0w_mem_0__31_0__26_;
  wire w_mem_inst__0w_mem_0__31_0__27_;
  wire w_mem_inst__0w_mem_0__31_0__28_;
  wire w_mem_inst__0w_mem_0__31_0__29_;
  wire w_mem_inst__0w_mem_0__31_0__2_;
  wire w_mem_inst__0w_mem_0__31_0__30_;
  wire w_mem_inst__0w_mem_0__31_0__31_;
  wire w_mem_inst__0w_mem_0__31_0__3_;
  wire w_mem_inst__0w_mem_0__31_0__4_;
  wire w_mem_inst__0w_mem_0__31_0__5_;
  wire w_mem_inst__0w_mem_0__31_0__6_;
  wire w_mem_inst__0w_mem_0__31_0__7_;
  wire w_mem_inst__0w_mem_0__31_0__8_;
  wire w_mem_inst__0w_mem_0__31_0__9_;
  wire w_mem_inst__0w_mem_10__31_0__0_;
  wire w_mem_inst__0w_mem_10__31_0__10_;
  wire w_mem_inst__0w_mem_10__31_0__11_;
  wire w_mem_inst__0w_mem_10__31_0__12_;
  wire w_mem_inst__0w_mem_10__31_0__13_;
  wire w_mem_inst__0w_mem_10__31_0__14_;
  wire w_mem_inst__0w_mem_10__31_0__15_;
  wire w_mem_inst__0w_mem_10__31_0__16_;
  wire w_mem_inst__0w_mem_10__31_0__17_;
  wire w_mem_inst__0w_mem_10__31_0__18_;
  wire w_mem_inst__0w_mem_10__31_0__19_;
  wire w_mem_inst__0w_mem_10__31_0__1_;
  wire w_mem_inst__0w_mem_10__31_0__20_;
  wire w_mem_inst__0w_mem_10__31_0__21_;
  wire w_mem_inst__0w_mem_10__31_0__22_;
  wire w_mem_inst__0w_mem_10__31_0__23_;
  wire w_mem_inst__0w_mem_10__31_0__24_;
  wire w_mem_inst__0w_mem_10__31_0__25_;
  wire w_mem_inst__0w_mem_10__31_0__26_;
  wire w_mem_inst__0w_mem_10__31_0__27_;
  wire w_mem_inst__0w_mem_10__31_0__28_;
  wire w_mem_inst__0w_mem_10__31_0__29_;
  wire w_mem_inst__0w_mem_10__31_0__2_;
  wire w_mem_inst__0w_mem_10__31_0__30_;
  wire w_mem_inst__0w_mem_10__31_0__31_;
  wire w_mem_inst__0w_mem_10__31_0__3_;
  wire w_mem_inst__0w_mem_10__31_0__4_;
  wire w_mem_inst__0w_mem_10__31_0__5_;
  wire w_mem_inst__0w_mem_10__31_0__6_;
  wire w_mem_inst__0w_mem_10__31_0__7_;
  wire w_mem_inst__0w_mem_10__31_0__8_;
  wire w_mem_inst__0w_mem_10__31_0__9_;
  wire w_mem_inst__0w_mem_11__31_0__0_;
  wire w_mem_inst__0w_mem_11__31_0__10_;
  wire w_mem_inst__0w_mem_11__31_0__11_;
  wire w_mem_inst__0w_mem_11__31_0__12_;
  wire w_mem_inst__0w_mem_11__31_0__13_;
  wire w_mem_inst__0w_mem_11__31_0__14_;
  wire w_mem_inst__0w_mem_11__31_0__15_;
  wire w_mem_inst__0w_mem_11__31_0__16_;
  wire w_mem_inst__0w_mem_11__31_0__17_;
  wire w_mem_inst__0w_mem_11__31_0__18_;
  wire w_mem_inst__0w_mem_11__31_0__19_;
  wire w_mem_inst__0w_mem_11__31_0__1_;
  wire w_mem_inst__0w_mem_11__31_0__20_;
  wire w_mem_inst__0w_mem_11__31_0__21_;
  wire w_mem_inst__0w_mem_11__31_0__22_;
  wire w_mem_inst__0w_mem_11__31_0__23_;
  wire w_mem_inst__0w_mem_11__31_0__24_;
  wire w_mem_inst__0w_mem_11__31_0__25_;
  wire w_mem_inst__0w_mem_11__31_0__26_;
  wire w_mem_inst__0w_mem_11__31_0__27_;
  wire w_mem_inst__0w_mem_11__31_0__28_;
  wire w_mem_inst__0w_mem_11__31_0__29_;
  wire w_mem_inst__0w_mem_11__31_0__2_;
  wire w_mem_inst__0w_mem_11__31_0__30_;
  wire w_mem_inst__0w_mem_11__31_0__31_;
  wire w_mem_inst__0w_mem_11__31_0__3_;
  wire w_mem_inst__0w_mem_11__31_0__4_;
  wire w_mem_inst__0w_mem_11__31_0__5_;
  wire w_mem_inst__0w_mem_11__31_0__6_;
  wire w_mem_inst__0w_mem_11__31_0__7_;
  wire w_mem_inst__0w_mem_11__31_0__8_;
  wire w_mem_inst__0w_mem_11__31_0__9_;
  wire w_mem_inst__0w_mem_12__31_0__0_;
  wire w_mem_inst__0w_mem_12__31_0__10_;
  wire w_mem_inst__0w_mem_12__31_0__11_;
  wire w_mem_inst__0w_mem_12__31_0__12_;
  wire w_mem_inst__0w_mem_12__31_0__13_;
  wire w_mem_inst__0w_mem_12__31_0__14_;
  wire w_mem_inst__0w_mem_12__31_0__15_;
  wire w_mem_inst__0w_mem_12__31_0__16_;
  wire w_mem_inst__0w_mem_12__31_0__17_;
  wire w_mem_inst__0w_mem_12__31_0__18_;
  wire w_mem_inst__0w_mem_12__31_0__19_;
  wire w_mem_inst__0w_mem_12__31_0__1_;
  wire w_mem_inst__0w_mem_12__31_0__20_;
  wire w_mem_inst__0w_mem_12__31_0__21_;
  wire w_mem_inst__0w_mem_12__31_0__22_;
  wire w_mem_inst__0w_mem_12__31_0__23_;
  wire w_mem_inst__0w_mem_12__31_0__24_;
  wire w_mem_inst__0w_mem_12__31_0__25_;
  wire w_mem_inst__0w_mem_12__31_0__26_;
  wire w_mem_inst__0w_mem_12__31_0__27_;
  wire w_mem_inst__0w_mem_12__31_0__28_;
  wire w_mem_inst__0w_mem_12__31_0__29_;
  wire w_mem_inst__0w_mem_12__31_0__2_;
  wire w_mem_inst__0w_mem_12__31_0__30_;
  wire w_mem_inst__0w_mem_12__31_0__31_;
  wire w_mem_inst__0w_mem_12__31_0__3_;
  wire w_mem_inst__0w_mem_12__31_0__4_;
  wire w_mem_inst__0w_mem_12__31_0__5_;
  wire w_mem_inst__0w_mem_12__31_0__6_;
  wire w_mem_inst__0w_mem_12__31_0__7_;
  wire w_mem_inst__0w_mem_12__31_0__8_;
  wire w_mem_inst__0w_mem_12__31_0__9_;
  wire w_mem_inst__0w_mem_13__31_0__0_;
  wire w_mem_inst__0w_mem_13__31_0__10_;
  wire w_mem_inst__0w_mem_13__31_0__11_;
  wire w_mem_inst__0w_mem_13__31_0__12_;
  wire w_mem_inst__0w_mem_13__31_0__13_;
  wire w_mem_inst__0w_mem_13__31_0__14_;
  wire w_mem_inst__0w_mem_13__31_0__15_;
  wire w_mem_inst__0w_mem_13__31_0__16_;
  wire w_mem_inst__0w_mem_13__31_0__17_;
  wire w_mem_inst__0w_mem_13__31_0__18_;
  wire w_mem_inst__0w_mem_13__31_0__19_;
  wire w_mem_inst__0w_mem_13__31_0__1_;
  wire w_mem_inst__0w_mem_13__31_0__20_;
  wire w_mem_inst__0w_mem_13__31_0__21_;
  wire w_mem_inst__0w_mem_13__31_0__22_;
  wire w_mem_inst__0w_mem_13__31_0__23_;
  wire w_mem_inst__0w_mem_13__31_0__24_;
  wire w_mem_inst__0w_mem_13__31_0__25_;
  wire w_mem_inst__0w_mem_13__31_0__26_;
  wire w_mem_inst__0w_mem_13__31_0__27_;
  wire w_mem_inst__0w_mem_13__31_0__28_;
  wire w_mem_inst__0w_mem_13__31_0__29_;
  wire w_mem_inst__0w_mem_13__31_0__2_;
  wire w_mem_inst__0w_mem_13__31_0__30_;
  wire w_mem_inst__0w_mem_13__31_0__31_;
  wire w_mem_inst__0w_mem_13__31_0__3_;
  wire w_mem_inst__0w_mem_13__31_0__4_;
  wire w_mem_inst__0w_mem_13__31_0__5_;
  wire w_mem_inst__0w_mem_13__31_0__6_;
  wire w_mem_inst__0w_mem_13__31_0__7_;
  wire w_mem_inst__0w_mem_13__31_0__8_;
  wire w_mem_inst__0w_mem_13__31_0__9_;
  wire w_mem_inst__0w_mem_14__31_0__0_;
  wire w_mem_inst__0w_mem_14__31_0__10_;
  wire w_mem_inst__0w_mem_14__31_0__11_;
  wire w_mem_inst__0w_mem_14__31_0__12_;
  wire w_mem_inst__0w_mem_14__31_0__13_;
  wire w_mem_inst__0w_mem_14__31_0__14_;
  wire w_mem_inst__0w_mem_14__31_0__15_;
  wire w_mem_inst__0w_mem_14__31_0__16_;
  wire w_mem_inst__0w_mem_14__31_0__17_;
  wire w_mem_inst__0w_mem_14__31_0__18_;
  wire w_mem_inst__0w_mem_14__31_0__19_;
  wire w_mem_inst__0w_mem_14__31_0__1_;
  wire w_mem_inst__0w_mem_14__31_0__20_;
  wire w_mem_inst__0w_mem_14__31_0__21_;
  wire w_mem_inst__0w_mem_14__31_0__22_;
  wire w_mem_inst__0w_mem_14__31_0__23_;
  wire w_mem_inst__0w_mem_14__31_0__24_;
  wire w_mem_inst__0w_mem_14__31_0__25_;
  wire w_mem_inst__0w_mem_14__31_0__26_;
  wire w_mem_inst__0w_mem_14__31_0__27_;
  wire w_mem_inst__0w_mem_14__31_0__28_;
  wire w_mem_inst__0w_mem_14__31_0__29_;
  wire w_mem_inst__0w_mem_14__31_0__2_;
  wire w_mem_inst__0w_mem_14__31_0__30_;
  wire w_mem_inst__0w_mem_14__31_0__31_;
  wire w_mem_inst__0w_mem_14__31_0__3_;
  wire w_mem_inst__0w_mem_14__31_0__4_;
  wire w_mem_inst__0w_mem_14__31_0__5_;
  wire w_mem_inst__0w_mem_14__31_0__6_;
  wire w_mem_inst__0w_mem_14__31_0__7_;
  wire w_mem_inst__0w_mem_14__31_0__8_;
  wire w_mem_inst__0w_mem_14__31_0__9_;
  wire w_mem_inst__0w_mem_15__31_0__0_;
  wire w_mem_inst__0w_mem_15__31_0__10_;
  wire w_mem_inst__0w_mem_15__31_0__11_;
  wire w_mem_inst__0w_mem_15__31_0__12_;
  wire w_mem_inst__0w_mem_15__31_0__13_;
  wire w_mem_inst__0w_mem_15__31_0__14_;
  wire w_mem_inst__0w_mem_15__31_0__15_;
  wire w_mem_inst__0w_mem_15__31_0__16_;
  wire w_mem_inst__0w_mem_15__31_0__17_;
  wire w_mem_inst__0w_mem_15__31_0__18_;
  wire w_mem_inst__0w_mem_15__31_0__19_;
  wire w_mem_inst__0w_mem_15__31_0__1_;
  wire w_mem_inst__0w_mem_15__31_0__20_;
  wire w_mem_inst__0w_mem_15__31_0__21_;
  wire w_mem_inst__0w_mem_15__31_0__22_;
  wire w_mem_inst__0w_mem_15__31_0__23_;
  wire w_mem_inst__0w_mem_15__31_0__24_;
  wire w_mem_inst__0w_mem_15__31_0__25_;
  wire w_mem_inst__0w_mem_15__31_0__26_;
  wire w_mem_inst__0w_mem_15__31_0__27_;
  wire w_mem_inst__0w_mem_15__31_0__28_;
  wire w_mem_inst__0w_mem_15__31_0__29_;
  wire w_mem_inst__0w_mem_15__31_0__2_;
  wire w_mem_inst__0w_mem_15__31_0__30_;
  wire w_mem_inst__0w_mem_15__31_0__31_;
  wire w_mem_inst__0w_mem_15__31_0__3_;
  wire w_mem_inst__0w_mem_15__31_0__4_;
  wire w_mem_inst__0w_mem_15__31_0__5_;
  wire w_mem_inst__0w_mem_15__31_0__6_;
  wire w_mem_inst__0w_mem_15__31_0__7_;
  wire w_mem_inst__0w_mem_15__31_0__8_;
  wire w_mem_inst__0w_mem_15__31_0__9_;
  wire w_mem_inst__0w_mem_1__31_0__0_;
  wire w_mem_inst__0w_mem_1__31_0__10_;
  wire w_mem_inst__0w_mem_1__31_0__11_;
  wire w_mem_inst__0w_mem_1__31_0__12_;
  wire w_mem_inst__0w_mem_1__31_0__13_;
  wire w_mem_inst__0w_mem_1__31_0__14_;
  wire w_mem_inst__0w_mem_1__31_0__15_;
  wire w_mem_inst__0w_mem_1__31_0__16_;
  wire w_mem_inst__0w_mem_1__31_0__17_;
  wire w_mem_inst__0w_mem_1__31_0__18_;
  wire w_mem_inst__0w_mem_1__31_0__19_;
  wire w_mem_inst__0w_mem_1__31_0__1_;
  wire w_mem_inst__0w_mem_1__31_0__20_;
  wire w_mem_inst__0w_mem_1__31_0__21_;
  wire w_mem_inst__0w_mem_1__31_0__22_;
  wire w_mem_inst__0w_mem_1__31_0__23_;
  wire w_mem_inst__0w_mem_1__31_0__24_;
  wire w_mem_inst__0w_mem_1__31_0__25_;
  wire w_mem_inst__0w_mem_1__31_0__26_;
  wire w_mem_inst__0w_mem_1__31_0__27_;
  wire w_mem_inst__0w_mem_1__31_0__28_;
  wire w_mem_inst__0w_mem_1__31_0__29_;
  wire w_mem_inst__0w_mem_1__31_0__2_;
  wire w_mem_inst__0w_mem_1__31_0__30_;
  wire w_mem_inst__0w_mem_1__31_0__31_;
  wire w_mem_inst__0w_mem_1__31_0__3_;
  wire w_mem_inst__0w_mem_1__31_0__4_;
  wire w_mem_inst__0w_mem_1__31_0__5_;
  wire w_mem_inst__0w_mem_1__31_0__6_;
  wire w_mem_inst__0w_mem_1__31_0__7_;
  wire w_mem_inst__0w_mem_1__31_0__8_;
  wire w_mem_inst__0w_mem_1__31_0__9_;
  wire w_mem_inst__0w_mem_2__31_0__0_;
  wire w_mem_inst__0w_mem_2__31_0__10_;
  wire w_mem_inst__0w_mem_2__31_0__11_;
  wire w_mem_inst__0w_mem_2__31_0__12_;
  wire w_mem_inst__0w_mem_2__31_0__13_;
  wire w_mem_inst__0w_mem_2__31_0__14_;
  wire w_mem_inst__0w_mem_2__31_0__15_;
  wire w_mem_inst__0w_mem_2__31_0__16_;
  wire w_mem_inst__0w_mem_2__31_0__17_;
  wire w_mem_inst__0w_mem_2__31_0__18_;
  wire w_mem_inst__0w_mem_2__31_0__19_;
  wire w_mem_inst__0w_mem_2__31_0__1_;
  wire w_mem_inst__0w_mem_2__31_0__20_;
  wire w_mem_inst__0w_mem_2__31_0__21_;
  wire w_mem_inst__0w_mem_2__31_0__22_;
  wire w_mem_inst__0w_mem_2__31_0__23_;
  wire w_mem_inst__0w_mem_2__31_0__24_;
  wire w_mem_inst__0w_mem_2__31_0__25_;
  wire w_mem_inst__0w_mem_2__31_0__26_;
  wire w_mem_inst__0w_mem_2__31_0__27_;
  wire w_mem_inst__0w_mem_2__31_0__28_;
  wire w_mem_inst__0w_mem_2__31_0__29_;
  wire w_mem_inst__0w_mem_2__31_0__2_;
  wire w_mem_inst__0w_mem_2__31_0__30_;
  wire w_mem_inst__0w_mem_2__31_0__31_;
  wire w_mem_inst__0w_mem_2__31_0__3_;
  wire w_mem_inst__0w_mem_2__31_0__4_;
  wire w_mem_inst__0w_mem_2__31_0__5_;
  wire w_mem_inst__0w_mem_2__31_0__6_;
  wire w_mem_inst__0w_mem_2__31_0__7_;
  wire w_mem_inst__0w_mem_2__31_0__8_;
  wire w_mem_inst__0w_mem_2__31_0__9_;
  wire w_mem_inst__0w_mem_3__31_0__0_;
  wire w_mem_inst__0w_mem_3__31_0__10_;
  wire w_mem_inst__0w_mem_3__31_0__11_;
  wire w_mem_inst__0w_mem_3__31_0__12_;
  wire w_mem_inst__0w_mem_3__31_0__13_;
  wire w_mem_inst__0w_mem_3__31_0__14_;
  wire w_mem_inst__0w_mem_3__31_0__15_;
  wire w_mem_inst__0w_mem_3__31_0__16_;
  wire w_mem_inst__0w_mem_3__31_0__17_;
  wire w_mem_inst__0w_mem_3__31_0__18_;
  wire w_mem_inst__0w_mem_3__31_0__19_;
  wire w_mem_inst__0w_mem_3__31_0__1_;
  wire w_mem_inst__0w_mem_3__31_0__20_;
  wire w_mem_inst__0w_mem_3__31_0__21_;
  wire w_mem_inst__0w_mem_3__31_0__22_;
  wire w_mem_inst__0w_mem_3__31_0__23_;
  wire w_mem_inst__0w_mem_3__31_0__24_;
  wire w_mem_inst__0w_mem_3__31_0__25_;
  wire w_mem_inst__0w_mem_3__31_0__26_;
  wire w_mem_inst__0w_mem_3__31_0__27_;
  wire w_mem_inst__0w_mem_3__31_0__28_;
  wire w_mem_inst__0w_mem_3__31_0__29_;
  wire w_mem_inst__0w_mem_3__31_0__2_;
  wire w_mem_inst__0w_mem_3__31_0__30_;
  wire w_mem_inst__0w_mem_3__31_0__31_;
  wire w_mem_inst__0w_mem_3__31_0__3_;
  wire w_mem_inst__0w_mem_3__31_0__4_;
  wire w_mem_inst__0w_mem_3__31_0__5_;
  wire w_mem_inst__0w_mem_3__31_0__6_;
  wire w_mem_inst__0w_mem_3__31_0__7_;
  wire w_mem_inst__0w_mem_3__31_0__8_;
  wire w_mem_inst__0w_mem_3__31_0__9_;
  wire w_mem_inst__0w_mem_4__31_0__0_;
  wire w_mem_inst__0w_mem_4__31_0__10_;
  wire w_mem_inst__0w_mem_4__31_0__11_;
  wire w_mem_inst__0w_mem_4__31_0__12_;
  wire w_mem_inst__0w_mem_4__31_0__13_;
  wire w_mem_inst__0w_mem_4__31_0__14_;
  wire w_mem_inst__0w_mem_4__31_0__15_;
  wire w_mem_inst__0w_mem_4__31_0__16_;
  wire w_mem_inst__0w_mem_4__31_0__17_;
  wire w_mem_inst__0w_mem_4__31_0__18_;
  wire w_mem_inst__0w_mem_4__31_0__19_;
  wire w_mem_inst__0w_mem_4__31_0__1_;
  wire w_mem_inst__0w_mem_4__31_0__20_;
  wire w_mem_inst__0w_mem_4__31_0__21_;
  wire w_mem_inst__0w_mem_4__31_0__22_;
  wire w_mem_inst__0w_mem_4__31_0__23_;
  wire w_mem_inst__0w_mem_4__31_0__24_;
  wire w_mem_inst__0w_mem_4__31_0__25_;
  wire w_mem_inst__0w_mem_4__31_0__26_;
  wire w_mem_inst__0w_mem_4__31_0__27_;
  wire w_mem_inst__0w_mem_4__31_0__28_;
  wire w_mem_inst__0w_mem_4__31_0__29_;
  wire w_mem_inst__0w_mem_4__31_0__2_;
  wire w_mem_inst__0w_mem_4__31_0__30_;
  wire w_mem_inst__0w_mem_4__31_0__31_;
  wire w_mem_inst__0w_mem_4__31_0__3_;
  wire w_mem_inst__0w_mem_4__31_0__4_;
  wire w_mem_inst__0w_mem_4__31_0__5_;
  wire w_mem_inst__0w_mem_4__31_0__6_;
  wire w_mem_inst__0w_mem_4__31_0__7_;
  wire w_mem_inst__0w_mem_4__31_0__8_;
  wire w_mem_inst__0w_mem_4__31_0__9_;
  wire w_mem_inst__0w_mem_5__31_0__0_;
  wire w_mem_inst__0w_mem_5__31_0__10_;
  wire w_mem_inst__0w_mem_5__31_0__11_;
  wire w_mem_inst__0w_mem_5__31_0__12_;
  wire w_mem_inst__0w_mem_5__31_0__13_;
  wire w_mem_inst__0w_mem_5__31_0__14_;
  wire w_mem_inst__0w_mem_5__31_0__15_;
  wire w_mem_inst__0w_mem_5__31_0__16_;
  wire w_mem_inst__0w_mem_5__31_0__17_;
  wire w_mem_inst__0w_mem_5__31_0__18_;
  wire w_mem_inst__0w_mem_5__31_0__19_;
  wire w_mem_inst__0w_mem_5__31_0__1_;
  wire w_mem_inst__0w_mem_5__31_0__20_;
  wire w_mem_inst__0w_mem_5__31_0__21_;
  wire w_mem_inst__0w_mem_5__31_0__22_;
  wire w_mem_inst__0w_mem_5__31_0__23_;
  wire w_mem_inst__0w_mem_5__31_0__24_;
  wire w_mem_inst__0w_mem_5__31_0__25_;
  wire w_mem_inst__0w_mem_5__31_0__26_;
  wire w_mem_inst__0w_mem_5__31_0__27_;
  wire w_mem_inst__0w_mem_5__31_0__28_;
  wire w_mem_inst__0w_mem_5__31_0__29_;
  wire w_mem_inst__0w_mem_5__31_0__2_;
  wire w_mem_inst__0w_mem_5__31_0__30_;
  wire w_mem_inst__0w_mem_5__31_0__31_;
  wire w_mem_inst__0w_mem_5__31_0__3_;
  wire w_mem_inst__0w_mem_5__31_0__4_;
  wire w_mem_inst__0w_mem_5__31_0__5_;
  wire w_mem_inst__0w_mem_5__31_0__6_;
  wire w_mem_inst__0w_mem_5__31_0__7_;
  wire w_mem_inst__0w_mem_5__31_0__8_;
  wire w_mem_inst__0w_mem_5__31_0__9_;
  wire w_mem_inst__0w_mem_6__31_0__0_;
  wire w_mem_inst__0w_mem_6__31_0__10_;
  wire w_mem_inst__0w_mem_6__31_0__11_;
  wire w_mem_inst__0w_mem_6__31_0__12_;
  wire w_mem_inst__0w_mem_6__31_0__13_;
  wire w_mem_inst__0w_mem_6__31_0__14_;
  wire w_mem_inst__0w_mem_6__31_0__15_;
  wire w_mem_inst__0w_mem_6__31_0__16_;
  wire w_mem_inst__0w_mem_6__31_0__17_;
  wire w_mem_inst__0w_mem_6__31_0__18_;
  wire w_mem_inst__0w_mem_6__31_0__19_;
  wire w_mem_inst__0w_mem_6__31_0__1_;
  wire w_mem_inst__0w_mem_6__31_0__20_;
  wire w_mem_inst__0w_mem_6__31_0__21_;
  wire w_mem_inst__0w_mem_6__31_0__22_;
  wire w_mem_inst__0w_mem_6__31_0__23_;
  wire w_mem_inst__0w_mem_6__31_0__24_;
  wire w_mem_inst__0w_mem_6__31_0__25_;
  wire w_mem_inst__0w_mem_6__31_0__26_;
  wire w_mem_inst__0w_mem_6__31_0__27_;
  wire w_mem_inst__0w_mem_6__31_0__28_;
  wire w_mem_inst__0w_mem_6__31_0__29_;
  wire w_mem_inst__0w_mem_6__31_0__2_;
  wire w_mem_inst__0w_mem_6__31_0__30_;
  wire w_mem_inst__0w_mem_6__31_0__31_;
  wire w_mem_inst__0w_mem_6__31_0__3_;
  wire w_mem_inst__0w_mem_6__31_0__4_;
  wire w_mem_inst__0w_mem_6__31_0__5_;
  wire w_mem_inst__0w_mem_6__31_0__6_;
  wire w_mem_inst__0w_mem_6__31_0__7_;
  wire w_mem_inst__0w_mem_6__31_0__8_;
  wire w_mem_inst__0w_mem_6__31_0__9_;
  wire w_mem_inst__0w_mem_7__31_0__0_;
  wire w_mem_inst__0w_mem_7__31_0__10_;
  wire w_mem_inst__0w_mem_7__31_0__11_;
  wire w_mem_inst__0w_mem_7__31_0__12_;
  wire w_mem_inst__0w_mem_7__31_0__13_;
  wire w_mem_inst__0w_mem_7__31_0__14_;
  wire w_mem_inst__0w_mem_7__31_0__15_;
  wire w_mem_inst__0w_mem_7__31_0__16_;
  wire w_mem_inst__0w_mem_7__31_0__17_;
  wire w_mem_inst__0w_mem_7__31_0__18_;
  wire w_mem_inst__0w_mem_7__31_0__19_;
  wire w_mem_inst__0w_mem_7__31_0__1_;
  wire w_mem_inst__0w_mem_7__31_0__20_;
  wire w_mem_inst__0w_mem_7__31_0__21_;
  wire w_mem_inst__0w_mem_7__31_0__22_;
  wire w_mem_inst__0w_mem_7__31_0__23_;
  wire w_mem_inst__0w_mem_7__31_0__24_;
  wire w_mem_inst__0w_mem_7__31_0__25_;
  wire w_mem_inst__0w_mem_7__31_0__26_;
  wire w_mem_inst__0w_mem_7__31_0__27_;
  wire w_mem_inst__0w_mem_7__31_0__28_;
  wire w_mem_inst__0w_mem_7__31_0__29_;
  wire w_mem_inst__0w_mem_7__31_0__2_;
  wire w_mem_inst__0w_mem_7__31_0__30_;
  wire w_mem_inst__0w_mem_7__31_0__31_;
  wire w_mem_inst__0w_mem_7__31_0__3_;
  wire w_mem_inst__0w_mem_7__31_0__4_;
  wire w_mem_inst__0w_mem_7__31_0__5_;
  wire w_mem_inst__0w_mem_7__31_0__6_;
  wire w_mem_inst__0w_mem_7__31_0__7_;
  wire w_mem_inst__0w_mem_7__31_0__8_;
  wire w_mem_inst__0w_mem_7__31_0__9_;
  wire w_mem_inst__0w_mem_8__31_0__0_;
  wire w_mem_inst__0w_mem_8__31_0__10_;
  wire w_mem_inst__0w_mem_8__31_0__11_;
  wire w_mem_inst__0w_mem_8__31_0__12_;
  wire w_mem_inst__0w_mem_8__31_0__13_;
  wire w_mem_inst__0w_mem_8__31_0__14_;
  wire w_mem_inst__0w_mem_8__31_0__15_;
  wire w_mem_inst__0w_mem_8__31_0__16_;
  wire w_mem_inst__0w_mem_8__31_0__17_;
  wire w_mem_inst__0w_mem_8__31_0__18_;
  wire w_mem_inst__0w_mem_8__31_0__19_;
  wire w_mem_inst__0w_mem_8__31_0__1_;
  wire w_mem_inst__0w_mem_8__31_0__20_;
  wire w_mem_inst__0w_mem_8__31_0__21_;
  wire w_mem_inst__0w_mem_8__31_0__22_;
  wire w_mem_inst__0w_mem_8__31_0__23_;
  wire w_mem_inst__0w_mem_8__31_0__24_;
  wire w_mem_inst__0w_mem_8__31_0__25_;
  wire w_mem_inst__0w_mem_8__31_0__26_;
  wire w_mem_inst__0w_mem_8__31_0__27_;
  wire w_mem_inst__0w_mem_8__31_0__28_;
  wire w_mem_inst__0w_mem_8__31_0__29_;
  wire w_mem_inst__0w_mem_8__31_0__2_;
  wire w_mem_inst__0w_mem_8__31_0__30_;
  wire w_mem_inst__0w_mem_8__31_0__31_;
  wire w_mem_inst__0w_mem_8__31_0__3_;
  wire w_mem_inst__0w_mem_8__31_0__4_;
  wire w_mem_inst__0w_mem_8__31_0__5_;
  wire w_mem_inst__0w_mem_8__31_0__6_;
  wire w_mem_inst__0w_mem_8__31_0__7_;
  wire w_mem_inst__0w_mem_8__31_0__8_;
  wire w_mem_inst__0w_mem_8__31_0__9_;
  wire w_mem_inst__0w_mem_9__31_0__0_;
  wire w_mem_inst__0w_mem_9__31_0__10_;
  wire w_mem_inst__0w_mem_9__31_0__11_;
  wire w_mem_inst__0w_mem_9__31_0__12_;
  wire w_mem_inst__0w_mem_9__31_0__13_;
  wire w_mem_inst__0w_mem_9__31_0__14_;
  wire w_mem_inst__0w_mem_9__31_0__15_;
  wire w_mem_inst__0w_mem_9__31_0__16_;
  wire w_mem_inst__0w_mem_9__31_0__17_;
  wire w_mem_inst__0w_mem_9__31_0__18_;
  wire w_mem_inst__0w_mem_9__31_0__19_;
  wire w_mem_inst__0w_mem_9__31_0__1_;
  wire w_mem_inst__0w_mem_9__31_0__20_;
  wire w_mem_inst__0w_mem_9__31_0__21_;
  wire w_mem_inst__0w_mem_9__31_0__22_;
  wire w_mem_inst__0w_mem_9__31_0__23_;
  wire w_mem_inst__0w_mem_9__31_0__24_;
  wire w_mem_inst__0w_mem_9__31_0__25_;
  wire w_mem_inst__0w_mem_9__31_0__26_;
  wire w_mem_inst__0w_mem_9__31_0__27_;
  wire w_mem_inst__0w_mem_9__31_0__28_;
  wire w_mem_inst__0w_mem_9__31_0__29_;
  wire w_mem_inst__0w_mem_9__31_0__2_;
  wire w_mem_inst__0w_mem_9__31_0__30_;
  wire w_mem_inst__0w_mem_9__31_0__31_;
  wire w_mem_inst__0w_mem_9__31_0__3_;
  wire w_mem_inst__0w_mem_9__31_0__4_;
  wire w_mem_inst__0w_mem_9__31_0__5_;
  wire w_mem_inst__0w_mem_9__31_0__6_;
  wire w_mem_inst__0w_mem_9__31_0__7_;
  wire w_mem_inst__0w_mem_9__31_0__8_;
  wire w_mem_inst__0w_mem_9__31_0__9_;
  wire w_mem_inst__abc_21378_n1585;
  wire w_mem_inst__abc_21378_n1586;
  wire w_mem_inst__abc_21378_n1586_bF_buf0;
  wire w_mem_inst__abc_21378_n1586_bF_buf1;
  wire w_mem_inst__abc_21378_n1586_bF_buf2;
  wire w_mem_inst__abc_21378_n1586_bF_buf3;
  wire w_mem_inst__abc_21378_n1586_bF_buf4;
  wire w_mem_inst__abc_21378_n1587;
  wire w_mem_inst__abc_21378_n1587_bF_buf0;
  wire w_mem_inst__abc_21378_n1587_bF_buf1;
  wire w_mem_inst__abc_21378_n1587_bF_buf2;
  wire w_mem_inst__abc_21378_n1587_bF_buf3;
  wire w_mem_inst__abc_21378_n1587_bF_buf4;
  wire w_mem_inst__abc_21378_n1588;
  wire w_mem_inst__abc_21378_n1589;
  wire w_mem_inst__abc_21378_n1590;
  wire w_mem_inst__abc_21378_n1591;
  wire w_mem_inst__abc_21378_n1592;
  wire w_mem_inst__abc_21378_n1593;
  wire w_mem_inst__abc_21378_n1594_1;
  wire w_mem_inst__abc_21378_n1595;
  wire w_mem_inst__abc_21378_n1596;
  wire w_mem_inst__abc_21378_n1597;
  wire w_mem_inst__abc_21378_n1598;
  wire w_mem_inst__abc_21378_n1599_1;
  wire w_mem_inst__abc_21378_n1600;
  wire w_mem_inst__abc_21378_n1601_1;
  wire w_mem_inst__abc_21378_n1602;
  wire w_mem_inst__abc_21378_n1603_1;
  wire w_mem_inst__abc_21378_n1604;
  wire w_mem_inst__abc_21378_n1605;
  wire w_mem_inst__abc_21378_n1605_bF_buf0;
  wire w_mem_inst__abc_21378_n1605_bF_buf1;
  wire w_mem_inst__abc_21378_n1605_bF_buf2;
  wire w_mem_inst__abc_21378_n1605_bF_buf3;
  wire w_mem_inst__abc_21378_n1605_bF_buf4;
  wire w_mem_inst__abc_21378_n1606_1;
  wire w_mem_inst__abc_21378_n1607_1;
  wire w_mem_inst__abc_21378_n1608;
  wire w_mem_inst__abc_21378_n1609;
  wire w_mem_inst__abc_21378_n1610_1;
  wire w_mem_inst__abc_21378_n1610_1_bF_buf0;
  wire w_mem_inst__abc_21378_n1610_1_bF_buf1;
  wire w_mem_inst__abc_21378_n1610_1_bF_buf2;
  wire w_mem_inst__abc_21378_n1610_1_bF_buf3;
  wire w_mem_inst__abc_21378_n1610_1_bF_buf4;
  wire w_mem_inst__abc_21378_n1611_1;
  wire w_mem_inst__abc_21378_n1612;
  wire w_mem_inst__abc_21378_n1613;
  wire w_mem_inst__abc_21378_n1614_1;
  wire w_mem_inst__abc_21378_n1615_1;
  wire w_mem_inst__abc_21378_n1616;
  wire w_mem_inst__abc_21378_n1616_bF_buf0;
  wire w_mem_inst__abc_21378_n1616_bF_buf1;
  wire w_mem_inst__abc_21378_n1616_bF_buf2;
  wire w_mem_inst__abc_21378_n1616_bF_buf3;
  wire w_mem_inst__abc_21378_n1616_bF_buf4;
  wire w_mem_inst__abc_21378_n1617;
  wire w_mem_inst__abc_21378_n1618_1;
  wire w_mem_inst__abc_21378_n1618_1_bF_buf0;
  wire w_mem_inst__abc_21378_n1618_1_bF_buf1;
  wire w_mem_inst__abc_21378_n1618_1_bF_buf2;
  wire w_mem_inst__abc_21378_n1618_1_bF_buf3;
  wire w_mem_inst__abc_21378_n1618_1_bF_buf4;
  wire w_mem_inst__abc_21378_n1619_1;
  wire w_mem_inst__abc_21378_n1620;
  wire w_mem_inst__abc_21378_n1621;
  wire w_mem_inst__abc_21378_n1622_1;
  wire w_mem_inst__abc_21378_n1623_1;
  wire w_mem_inst__abc_21378_n1624;
  wire w_mem_inst__abc_21378_n1625;
  wire w_mem_inst__abc_21378_n1625_bF_buf0;
  wire w_mem_inst__abc_21378_n1625_bF_buf1;
  wire w_mem_inst__abc_21378_n1625_bF_buf2;
  wire w_mem_inst__abc_21378_n1625_bF_buf3;
  wire w_mem_inst__abc_21378_n1625_bF_buf4;
  wire w_mem_inst__abc_21378_n1626_1;
  wire w_mem_inst__abc_21378_n1627_1;
  wire w_mem_inst__abc_21378_n1627_1_bF_buf0;
  wire w_mem_inst__abc_21378_n1627_1_bF_buf1;
  wire w_mem_inst__abc_21378_n1627_1_bF_buf2;
  wire w_mem_inst__abc_21378_n1627_1_bF_buf3;
  wire w_mem_inst__abc_21378_n1627_1_bF_buf4;
  wire w_mem_inst__abc_21378_n1628;
  wire w_mem_inst__abc_21378_n1629;
  wire w_mem_inst__abc_21378_n1630_1;
  wire w_mem_inst__abc_21378_n1630_1_bF_buf0;
  wire w_mem_inst__abc_21378_n1630_1_bF_buf1;
  wire w_mem_inst__abc_21378_n1630_1_bF_buf2;
  wire w_mem_inst__abc_21378_n1630_1_bF_buf3;
  wire w_mem_inst__abc_21378_n1630_1_bF_buf4;
  wire w_mem_inst__abc_21378_n1631_1;
  wire w_mem_inst__abc_21378_n1632;
  wire w_mem_inst__abc_21378_n1633;
  wire w_mem_inst__abc_21378_n1634_1;
  wire w_mem_inst__abc_21378_n1634_1_bF_buf0;
  wire w_mem_inst__abc_21378_n1634_1_bF_buf1;
  wire w_mem_inst__abc_21378_n1634_1_bF_buf2;
  wire w_mem_inst__abc_21378_n1634_1_bF_buf3;
  wire w_mem_inst__abc_21378_n1634_1_bF_buf4;
  wire w_mem_inst__abc_21378_n1635_1;
  wire w_mem_inst__abc_21378_n1636;
  wire w_mem_inst__abc_21378_n1637;
  wire w_mem_inst__abc_21378_n1638_1;
  wire w_mem_inst__abc_21378_n1638_1_bF_buf0;
  wire w_mem_inst__abc_21378_n1638_1_bF_buf1;
  wire w_mem_inst__abc_21378_n1638_1_bF_buf2;
  wire w_mem_inst__abc_21378_n1638_1_bF_buf3;
  wire w_mem_inst__abc_21378_n1638_1_bF_buf4;
  wire w_mem_inst__abc_21378_n1639_1;
  wire w_mem_inst__abc_21378_n1640;
  wire w_mem_inst__abc_21378_n1640_bF_buf0;
  wire w_mem_inst__abc_21378_n1640_bF_buf1;
  wire w_mem_inst__abc_21378_n1640_bF_buf2;
  wire w_mem_inst__abc_21378_n1640_bF_buf3;
  wire w_mem_inst__abc_21378_n1640_bF_buf4;
  wire w_mem_inst__abc_21378_n1641;
  wire w_mem_inst__abc_21378_n1642_1;
  wire w_mem_inst__abc_21378_n1643_1;
  wire w_mem_inst__abc_21378_n1643_1_bF_buf0;
  wire w_mem_inst__abc_21378_n1643_1_bF_buf1;
  wire w_mem_inst__abc_21378_n1643_1_bF_buf2;
  wire w_mem_inst__abc_21378_n1643_1_bF_buf3;
  wire w_mem_inst__abc_21378_n1643_1_bF_buf4;
  wire w_mem_inst__abc_21378_n1644;
  wire w_mem_inst__abc_21378_n1645;
  wire w_mem_inst__abc_21378_n1645_bF_buf0;
  wire w_mem_inst__abc_21378_n1645_bF_buf1;
  wire w_mem_inst__abc_21378_n1645_bF_buf2;
  wire w_mem_inst__abc_21378_n1645_bF_buf3;
  wire w_mem_inst__abc_21378_n1645_bF_buf4;
  wire w_mem_inst__abc_21378_n1646_1;
  wire w_mem_inst__abc_21378_n1647_1;
  wire w_mem_inst__abc_21378_n1648;
  wire w_mem_inst__abc_21378_n1649;
  wire w_mem_inst__abc_21378_n1649_bF_buf0;
  wire w_mem_inst__abc_21378_n1649_bF_buf1;
  wire w_mem_inst__abc_21378_n1649_bF_buf2;
  wire w_mem_inst__abc_21378_n1649_bF_buf3;
  wire w_mem_inst__abc_21378_n1649_bF_buf4;
  wire w_mem_inst__abc_21378_n1650_1;
  wire w_mem_inst__abc_21378_n1651_1;
  wire w_mem_inst__abc_21378_n1651_1_bF_buf0;
  wire w_mem_inst__abc_21378_n1651_1_bF_buf1;
  wire w_mem_inst__abc_21378_n1651_1_bF_buf2;
  wire w_mem_inst__abc_21378_n1651_1_bF_buf3;
  wire w_mem_inst__abc_21378_n1651_1_bF_buf4;
  wire w_mem_inst__abc_21378_n1652;
  wire w_mem_inst__abc_21378_n1653;
  wire w_mem_inst__abc_21378_n1654_1;
  wire w_mem_inst__abc_21378_n1654_1_bF_buf0;
  wire w_mem_inst__abc_21378_n1654_1_bF_buf1;
  wire w_mem_inst__abc_21378_n1654_1_bF_buf2;
  wire w_mem_inst__abc_21378_n1654_1_bF_buf3;
  wire w_mem_inst__abc_21378_n1654_1_bF_buf4;
  wire w_mem_inst__abc_21378_n1655_1;
  wire w_mem_inst__abc_21378_n1656;
  wire w_mem_inst__abc_21378_n1656_bF_buf0;
  wire w_mem_inst__abc_21378_n1656_bF_buf1;
  wire w_mem_inst__abc_21378_n1656_bF_buf2;
  wire w_mem_inst__abc_21378_n1656_bF_buf3;
  wire w_mem_inst__abc_21378_n1656_bF_buf4;
  wire w_mem_inst__abc_21378_n1657;
  wire w_mem_inst__abc_21378_n1658_1;
  wire w_mem_inst__abc_21378_n1659_1;
  wire w_mem_inst__abc_21378_n1660;
  wire w_mem_inst__abc_21378_n1661;
  wire w_mem_inst__abc_21378_n1662_1;
  wire w_mem_inst__abc_21378_n1664;
  wire w_mem_inst__abc_21378_n1665;
  wire w_mem_inst__abc_21378_n1666_1;
  wire w_mem_inst__abc_21378_n1667_1;
  wire w_mem_inst__abc_21378_n1668;
  wire w_mem_inst__abc_21378_n1669;
  wire w_mem_inst__abc_21378_n1670_1;
  wire w_mem_inst__abc_21378_n1671_1;
  wire w_mem_inst__abc_21378_n1672;
  wire w_mem_inst__abc_21378_n1673;
  wire w_mem_inst__abc_21378_n1674_1;
  wire w_mem_inst__abc_21378_n1675_1;
  wire w_mem_inst__abc_21378_n1676;
  wire w_mem_inst__abc_21378_n1677;
  wire w_mem_inst__abc_21378_n1678_1;
  wire w_mem_inst__abc_21378_n1679_1;
  wire w_mem_inst__abc_21378_n1680;
  wire w_mem_inst__abc_21378_n1681;
  wire w_mem_inst__abc_21378_n1682_1;
  wire w_mem_inst__abc_21378_n1683_1;
  wire w_mem_inst__abc_21378_n1684;
  wire w_mem_inst__abc_21378_n1685;
  wire w_mem_inst__abc_21378_n1686_1;
  wire w_mem_inst__abc_21378_n1687_1;
  wire w_mem_inst__abc_21378_n1688;
  wire w_mem_inst__abc_21378_n1689;
  wire w_mem_inst__abc_21378_n1690_1;
  wire w_mem_inst__abc_21378_n1691_1;
  wire w_mem_inst__abc_21378_n1692;
  wire w_mem_inst__abc_21378_n1693;
  wire w_mem_inst__abc_21378_n1694_1;
  wire w_mem_inst__abc_21378_n1695_1;
  wire w_mem_inst__abc_21378_n1696;
  wire w_mem_inst__abc_21378_n1697;
  wire w_mem_inst__abc_21378_n1698_1;
  wire w_mem_inst__abc_21378_n1699_1;
  wire w_mem_inst__abc_21378_n1700;
  wire w_mem_inst__abc_21378_n1701;
  wire w_mem_inst__abc_21378_n1702_1;
  wire w_mem_inst__abc_21378_n1703_1;
  wire w_mem_inst__abc_21378_n1704;
  wire w_mem_inst__abc_21378_n1705;
  wire w_mem_inst__abc_21378_n1706_1;
  wire w_mem_inst__abc_21378_n1707_1;
  wire w_mem_inst__abc_21378_n1708;
  wire w_mem_inst__abc_21378_n1709;
  wire w_mem_inst__abc_21378_n1710_1;
  wire w_mem_inst__abc_21378_n1712;
  wire w_mem_inst__abc_21378_n1713;
  wire w_mem_inst__abc_21378_n1714_1;
  wire w_mem_inst__abc_21378_n1715_1;
  wire w_mem_inst__abc_21378_n1716;
  wire w_mem_inst__abc_21378_n1717;
  wire w_mem_inst__abc_21378_n1718_1;
  wire w_mem_inst__abc_21378_n1719_1;
  wire w_mem_inst__abc_21378_n1720;
  wire w_mem_inst__abc_21378_n1721;
  wire w_mem_inst__abc_21378_n1722_1;
  wire w_mem_inst__abc_21378_n1723_1;
  wire w_mem_inst__abc_21378_n1724;
  wire w_mem_inst__abc_21378_n1725;
  wire w_mem_inst__abc_21378_n1726_1;
  wire w_mem_inst__abc_21378_n1727_1;
  wire w_mem_inst__abc_21378_n1728;
  wire w_mem_inst__abc_21378_n1729;
  wire w_mem_inst__abc_21378_n1730_1;
  wire w_mem_inst__abc_21378_n1731_1;
  wire w_mem_inst__abc_21378_n1732;
  wire w_mem_inst__abc_21378_n1733;
  wire w_mem_inst__abc_21378_n1734_1;
  wire w_mem_inst__abc_21378_n1735_1;
  wire w_mem_inst__abc_21378_n1736;
  wire w_mem_inst__abc_21378_n1737;
  wire w_mem_inst__abc_21378_n1738_1;
  wire w_mem_inst__abc_21378_n1739_1;
  wire w_mem_inst__abc_21378_n1740;
  wire w_mem_inst__abc_21378_n1741;
  wire w_mem_inst__abc_21378_n1742_1;
  wire w_mem_inst__abc_21378_n1743_1;
  wire w_mem_inst__abc_21378_n1744;
  wire w_mem_inst__abc_21378_n1745;
  wire w_mem_inst__abc_21378_n1746_1;
  wire w_mem_inst__abc_21378_n1747_1;
  wire w_mem_inst__abc_21378_n1748;
  wire w_mem_inst__abc_21378_n1749;
  wire w_mem_inst__abc_21378_n1750_1;
  wire w_mem_inst__abc_21378_n1751_1;
  wire w_mem_inst__abc_21378_n1752;
  wire w_mem_inst__abc_21378_n1753;
  wire w_mem_inst__abc_21378_n1754_1;
  wire w_mem_inst__abc_21378_n1755_1;
  wire w_mem_inst__abc_21378_n1756;
  wire w_mem_inst__abc_21378_n1757;
  wire w_mem_inst__abc_21378_n1758_1;
  wire w_mem_inst__abc_21378_n1760;
  wire w_mem_inst__abc_21378_n1761;
  wire w_mem_inst__abc_21378_n1762_1;
  wire w_mem_inst__abc_21378_n1763_1;
  wire w_mem_inst__abc_21378_n1764;
  wire w_mem_inst__abc_21378_n1765;
  wire w_mem_inst__abc_21378_n1766_1;
  wire w_mem_inst__abc_21378_n1767_1;
  wire w_mem_inst__abc_21378_n1768;
  wire w_mem_inst__abc_21378_n1769;
  wire w_mem_inst__abc_21378_n1770_1;
  wire w_mem_inst__abc_21378_n1771_1;
  wire w_mem_inst__abc_21378_n1772;
  wire w_mem_inst__abc_21378_n1773;
  wire w_mem_inst__abc_21378_n1774_1;
  wire w_mem_inst__abc_21378_n1775_1;
  wire w_mem_inst__abc_21378_n1776;
  wire w_mem_inst__abc_21378_n1777;
  wire w_mem_inst__abc_21378_n1778_1;
  wire w_mem_inst__abc_21378_n1779_1;
  wire w_mem_inst__abc_21378_n1780;
  wire w_mem_inst__abc_21378_n1781;
  wire w_mem_inst__abc_21378_n1782_1;
  wire w_mem_inst__abc_21378_n1783_1;
  wire w_mem_inst__abc_21378_n1784;
  wire w_mem_inst__abc_21378_n1785;
  wire w_mem_inst__abc_21378_n1786_1;
  wire w_mem_inst__abc_21378_n1787_1;
  wire w_mem_inst__abc_21378_n1788;
  wire w_mem_inst__abc_21378_n1789;
  wire w_mem_inst__abc_21378_n1790_1;
  wire w_mem_inst__abc_21378_n1791_1;
  wire w_mem_inst__abc_21378_n1792;
  wire w_mem_inst__abc_21378_n1793;
  wire w_mem_inst__abc_21378_n1794_1;
  wire w_mem_inst__abc_21378_n1795_1;
  wire w_mem_inst__abc_21378_n1796;
  wire w_mem_inst__abc_21378_n1797;
  wire w_mem_inst__abc_21378_n1798_1;
  wire w_mem_inst__abc_21378_n1799_1;
  wire w_mem_inst__abc_21378_n1800;
  wire w_mem_inst__abc_21378_n1801;
  wire w_mem_inst__abc_21378_n1802_1;
  wire w_mem_inst__abc_21378_n1803_1;
  wire w_mem_inst__abc_21378_n1804;
  wire w_mem_inst__abc_21378_n1805;
  wire w_mem_inst__abc_21378_n1806_1;
  wire w_mem_inst__abc_21378_n1808;
  wire w_mem_inst__abc_21378_n1809;
  wire w_mem_inst__abc_21378_n1810_1;
  wire w_mem_inst__abc_21378_n1811_1;
  wire w_mem_inst__abc_21378_n1812;
  wire w_mem_inst__abc_21378_n1813;
  wire w_mem_inst__abc_21378_n1814_1;
  wire w_mem_inst__abc_21378_n1815_1;
  wire w_mem_inst__abc_21378_n1816;
  wire w_mem_inst__abc_21378_n1817;
  wire w_mem_inst__abc_21378_n1818_1;
  wire w_mem_inst__abc_21378_n1819_1;
  wire w_mem_inst__abc_21378_n1820;
  wire w_mem_inst__abc_21378_n1821;
  wire w_mem_inst__abc_21378_n1822_1;
  wire w_mem_inst__abc_21378_n1823_1;
  wire w_mem_inst__abc_21378_n1824;
  wire w_mem_inst__abc_21378_n1825;
  wire w_mem_inst__abc_21378_n1826_1;
  wire w_mem_inst__abc_21378_n1827_1;
  wire w_mem_inst__abc_21378_n1828;
  wire w_mem_inst__abc_21378_n1829;
  wire w_mem_inst__abc_21378_n1830_1;
  wire w_mem_inst__abc_21378_n1831_1;
  wire w_mem_inst__abc_21378_n1832;
  wire w_mem_inst__abc_21378_n1833;
  wire w_mem_inst__abc_21378_n1834_1;
  wire w_mem_inst__abc_21378_n1835_1;
  wire w_mem_inst__abc_21378_n1836;
  wire w_mem_inst__abc_21378_n1837;
  wire w_mem_inst__abc_21378_n1838_1;
  wire w_mem_inst__abc_21378_n1839_1;
  wire w_mem_inst__abc_21378_n1840;
  wire w_mem_inst__abc_21378_n1841;
  wire w_mem_inst__abc_21378_n1842_1;
  wire w_mem_inst__abc_21378_n1843_1;
  wire w_mem_inst__abc_21378_n1844;
  wire w_mem_inst__abc_21378_n1845;
  wire w_mem_inst__abc_21378_n1846_1;
  wire w_mem_inst__abc_21378_n1847_1;
  wire w_mem_inst__abc_21378_n1848;
  wire w_mem_inst__abc_21378_n1849;
  wire w_mem_inst__abc_21378_n1850_1;
  wire w_mem_inst__abc_21378_n1851_1;
  wire w_mem_inst__abc_21378_n1852;
  wire w_mem_inst__abc_21378_n1853;
  wire w_mem_inst__abc_21378_n1854_1;
  wire w_mem_inst__abc_21378_n1856;
  wire w_mem_inst__abc_21378_n1857;
  wire w_mem_inst__abc_21378_n1858_1;
  wire w_mem_inst__abc_21378_n1859_1;
  wire w_mem_inst__abc_21378_n1860;
  wire w_mem_inst__abc_21378_n1861;
  wire w_mem_inst__abc_21378_n1862_1;
  wire w_mem_inst__abc_21378_n1863_1;
  wire w_mem_inst__abc_21378_n1864;
  wire w_mem_inst__abc_21378_n1865;
  wire w_mem_inst__abc_21378_n1866_1;
  wire w_mem_inst__abc_21378_n1867_1;
  wire w_mem_inst__abc_21378_n1868;
  wire w_mem_inst__abc_21378_n1869;
  wire w_mem_inst__abc_21378_n1870_1;
  wire w_mem_inst__abc_21378_n1871_1;
  wire w_mem_inst__abc_21378_n1872;
  wire w_mem_inst__abc_21378_n1873;
  wire w_mem_inst__abc_21378_n1874_1;
  wire w_mem_inst__abc_21378_n1875_1;
  wire w_mem_inst__abc_21378_n1876;
  wire w_mem_inst__abc_21378_n1877;
  wire w_mem_inst__abc_21378_n1878_1;
  wire w_mem_inst__abc_21378_n1879_1;
  wire w_mem_inst__abc_21378_n1880;
  wire w_mem_inst__abc_21378_n1881;
  wire w_mem_inst__abc_21378_n1882_1;
  wire w_mem_inst__abc_21378_n1883_1;
  wire w_mem_inst__abc_21378_n1884;
  wire w_mem_inst__abc_21378_n1885;
  wire w_mem_inst__abc_21378_n1886_1;
  wire w_mem_inst__abc_21378_n1887_1;
  wire w_mem_inst__abc_21378_n1888;
  wire w_mem_inst__abc_21378_n1889;
  wire w_mem_inst__abc_21378_n1890_1;
  wire w_mem_inst__abc_21378_n1891_1;
  wire w_mem_inst__abc_21378_n1892;
  wire w_mem_inst__abc_21378_n1893;
  wire w_mem_inst__abc_21378_n1894_1;
  wire w_mem_inst__abc_21378_n1895_1;
  wire w_mem_inst__abc_21378_n1896;
  wire w_mem_inst__abc_21378_n1897;
  wire w_mem_inst__abc_21378_n1898_1;
  wire w_mem_inst__abc_21378_n1899_1;
  wire w_mem_inst__abc_21378_n1900;
  wire w_mem_inst__abc_21378_n1901;
  wire w_mem_inst__abc_21378_n1902_1;
  wire w_mem_inst__abc_21378_n1904;
  wire w_mem_inst__abc_21378_n1905;
  wire w_mem_inst__abc_21378_n1906_1;
  wire w_mem_inst__abc_21378_n1907_1;
  wire w_mem_inst__abc_21378_n1908;
  wire w_mem_inst__abc_21378_n1909;
  wire w_mem_inst__abc_21378_n1910_1;
  wire w_mem_inst__abc_21378_n1911_1;
  wire w_mem_inst__abc_21378_n1912;
  wire w_mem_inst__abc_21378_n1913;
  wire w_mem_inst__abc_21378_n1914_1;
  wire w_mem_inst__abc_21378_n1915_1;
  wire w_mem_inst__abc_21378_n1916;
  wire w_mem_inst__abc_21378_n1917;
  wire w_mem_inst__abc_21378_n1918_1;
  wire w_mem_inst__abc_21378_n1919_1;
  wire w_mem_inst__abc_21378_n1920;
  wire w_mem_inst__abc_21378_n1921;
  wire w_mem_inst__abc_21378_n1922_1;
  wire w_mem_inst__abc_21378_n1923_1;
  wire w_mem_inst__abc_21378_n1924;
  wire w_mem_inst__abc_21378_n1925;
  wire w_mem_inst__abc_21378_n1926_1;
  wire w_mem_inst__abc_21378_n1927_1;
  wire w_mem_inst__abc_21378_n1928;
  wire w_mem_inst__abc_21378_n1929;
  wire w_mem_inst__abc_21378_n1930_1;
  wire w_mem_inst__abc_21378_n1931_1;
  wire w_mem_inst__abc_21378_n1932;
  wire w_mem_inst__abc_21378_n1933;
  wire w_mem_inst__abc_21378_n1934_1;
  wire w_mem_inst__abc_21378_n1935_1;
  wire w_mem_inst__abc_21378_n1936;
  wire w_mem_inst__abc_21378_n1937;
  wire w_mem_inst__abc_21378_n1938_1;
  wire w_mem_inst__abc_21378_n1939_1;
  wire w_mem_inst__abc_21378_n1940;
  wire w_mem_inst__abc_21378_n1941;
  wire w_mem_inst__abc_21378_n1942_1;
  wire w_mem_inst__abc_21378_n1943_1;
  wire w_mem_inst__abc_21378_n1944;
  wire w_mem_inst__abc_21378_n1945;
  wire w_mem_inst__abc_21378_n1946_1;
  wire w_mem_inst__abc_21378_n1947_1;
  wire w_mem_inst__abc_21378_n1948;
  wire w_mem_inst__abc_21378_n1949;
  wire w_mem_inst__abc_21378_n1950_1;
  wire w_mem_inst__abc_21378_n1952;
  wire w_mem_inst__abc_21378_n1953;
  wire w_mem_inst__abc_21378_n1954_1;
  wire w_mem_inst__abc_21378_n1955_1;
  wire w_mem_inst__abc_21378_n1956;
  wire w_mem_inst__abc_21378_n1957;
  wire w_mem_inst__abc_21378_n1958_1;
  wire w_mem_inst__abc_21378_n1959_1;
  wire w_mem_inst__abc_21378_n1960;
  wire w_mem_inst__abc_21378_n1961;
  wire w_mem_inst__abc_21378_n1962_1;
  wire w_mem_inst__abc_21378_n1963_1;
  wire w_mem_inst__abc_21378_n1964;
  wire w_mem_inst__abc_21378_n1965;
  wire w_mem_inst__abc_21378_n1966_1;
  wire w_mem_inst__abc_21378_n1967_1;
  wire w_mem_inst__abc_21378_n1968;
  wire w_mem_inst__abc_21378_n1969;
  wire w_mem_inst__abc_21378_n1970_1;
  wire w_mem_inst__abc_21378_n1971_1;
  wire w_mem_inst__abc_21378_n1972;
  wire w_mem_inst__abc_21378_n1973;
  wire w_mem_inst__abc_21378_n1974_1;
  wire w_mem_inst__abc_21378_n1975_1;
  wire w_mem_inst__abc_21378_n1976;
  wire w_mem_inst__abc_21378_n1977;
  wire w_mem_inst__abc_21378_n1978_1;
  wire w_mem_inst__abc_21378_n1979_1;
  wire w_mem_inst__abc_21378_n1980;
  wire w_mem_inst__abc_21378_n1981;
  wire w_mem_inst__abc_21378_n1982_1;
  wire w_mem_inst__abc_21378_n1983_1;
  wire w_mem_inst__abc_21378_n1984;
  wire w_mem_inst__abc_21378_n1985;
  wire w_mem_inst__abc_21378_n1986_1;
  wire w_mem_inst__abc_21378_n1987_1;
  wire w_mem_inst__abc_21378_n1988;
  wire w_mem_inst__abc_21378_n1989;
  wire w_mem_inst__abc_21378_n1990_1;
  wire w_mem_inst__abc_21378_n1991_1;
  wire w_mem_inst__abc_21378_n1992;
  wire w_mem_inst__abc_21378_n1993;
  wire w_mem_inst__abc_21378_n1994_1;
  wire w_mem_inst__abc_21378_n1995_1;
  wire w_mem_inst__abc_21378_n1996;
  wire w_mem_inst__abc_21378_n1997;
  wire w_mem_inst__abc_21378_n1998_1;
  wire w_mem_inst__abc_21378_n2000;
  wire w_mem_inst__abc_21378_n2001;
  wire w_mem_inst__abc_21378_n2002_1;
  wire w_mem_inst__abc_21378_n2003_1;
  wire w_mem_inst__abc_21378_n2004;
  wire w_mem_inst__abc_21378_n2005;
  wire w_mem_inst__abc_21378_n2006_1;
  wire w_mem_inst__abc_21378_n2007_1;
  wire w_mem_inst__abc_21378_n2008;
  wire w_mem_inst__abc_21378_n2009;
  wire w_mem_inst__abc_21378_n2010_1;
  wire w_mem_inst__abc_21378_n2011_1;
  wire w_mem_inst__abc_21378_n2012;
  wire w_mem_inst__abc_21378_n2013;
  wire w_mem_inst__abc_21378_n2014_1;
  wire w_mem_inst__abc_21378_n2015_1;
  wire w_mem_inst__abc_21378_n2016;
  wire w_mem_inst__abc_21378_n2017;
  wire w_mem_inst__abc_21378_n2018_1;
  wire w_mem_inst__abc_21378_n2019_1;
  wire w_mem_inst__abc_21378_n2020;
  wire w_mem_inst__abc_21378_n2021;
  wire w_mem_inst__abc_21378_n2022_1;
  wire w_mem_inst__abc_21378_n2023_1;
  wire w_mem_inst__abc_21378_n2024;
  wire w_mem_inst__abc_21378_n2025;
  wire w_mem_inst__abc_21378_n2026_1;
  wire w_mem_inst__abc_21378_n2027_1;
  wire w_mem_inst__abc_21378_n2028;
  wire w_mem_inst__abc_21378_n2029;
  wire w_mem_inst__abc_21378_n2030_1;
  wire w_mem_inst__abc_21378_n2031_1;
  wire w_mem_inst__abc_21378_n2032;
  wire w_mem_inst__abc_21378_n2033;
  wire w_mem_inst__abc_21378_n2034_1;
  wire w_mem_inst__abc_21378_n2035_1;
  wire w_mem_inst__abc_21378_n2036;
  wire w_mem_inst__abc_21378_n2037;
  wire w_mem_inst__abc_21378_n2038_1;
  wire w_mem_inst__abc_21378_n2039_1;
  wire w_mem_inst__abc_21378_n2040;
  wire w_mem_inst__abc_21378_n2041;
  wire w_mem_inst__abc_21378_n2042_1;
  wire w_mem_inst__abc_21378_n2043_1;
  wire w_mem_inst__abc_21378_n2044;
  wire w_mem_inst__abc_21378_n2045;
  wire w_mem_inst__abc_21378_n2046_1;
  wire w_mem_inst__abc_21378_n2048;
  wire w_mem_inst__abc_21378_n2049;
  wire w_mem_inst__abc_21378_n2050_1;
  wire w_mem_inst__abc_21378_n2051_1;
  wire w_mem_inst__abc_21378_n2052;
  wire w_mem_inst__abc_21378_n2053;
  wire w_mem_inst__abc_21378_n2054_1;
  wire w_mem_inst__abc_21378_n2055_1;
  wire w_mem_inst__abc_21378_n2056;
  wire w_mem_inst__abc_21378_n2057;
  wire w_mem_inst__abc_21378_n2058_1;
  wire w_mem_inst__abc_21378_n2059_1;
  wire w_mem_inst__abc_21378_n2060;
  wire w_mem_inst__abc_21378_n2061;
  wire w_mem_inst__abc_21378_n2062_1;
  wire w_mem_inst__abc_21378_n2063_1;
  wire w_mem_inst__abc_21378_n2064;
  wire w_mem_inst__abc_21378_n2065;
  wire w_mem_inst__abc_21378_n2066_1;
  wire w_mem_inst__abc_21378_n2067_1;
  wire w_mem_inst__abc_21378_n2068;
  wire w_mem_inst__abc_21378_n2069;
  wire w_mem_inst__abc_21378_n2070_1;
  wire w_mem_inst__abc_21378_n2071_1;
  wire w_mem_inst__abc_21378_n2072;
  wire w_mem_inst__abc_21378_n2073;
  wire w_mem_inst__abc_21378_n2074_1;
  wire w_mem_inst__abc_21378_n2075_1;
  wire w_mem_inst__abc_21378_n2076;
  wire w_mem_inst__abc_21378_n2077;
  wire w_mem_inst__abc_21378_n2078_1;
  wire w_mem_inst__abc_21378_n2079_1;
  wire w_mem_inst__abc_21378_n2080;
  wire w_mem_inst__abc_21378_n2081;
  wire w_mem_inst__abc_21378_n2082_1;
  wire w_mem_inst__abc_21378_n2083_1;
  wire w_mem_inst__abc_21378_n2084;
  wire w_mem_inst__abc_21378_n2085;
  wire w_mem_inst__abc_21378_n2086_1;
  wire w_mem_inst__abc_21378_n2087_1;
  wire w_mem_inst__abc_21378_n2088;
  wire w_mem_inst__abc_21378_n2089;
  wire w_mem_inst__abc_21378_n2090_1;
  wire w_mem_inst__abc_21378_n2091_1;
  wire w_mem_inst__abc_21378_n2092;
  wire w_mem_inst__abc_21378_n2093;
  wire w_mem_inst__abc_21378_n2094_1;
  wire w_mem_inst__abc_21378_n2096;
  wire w_mem_inst__abc_21378_n2097;
  wire w_mem_inst__abc_21378_n2098_1;
  wire w_mem_inst__abc_21378_n2099_1;
  wire w_mem_inst__abc_21378_n2100;
  wire w_mem_inst__abc_21378_n2101;
  wire w_mem_inst__abc_21378_n2102_1;
  wire w_mem_inst__abc_21378_n2103_1;
  wire w_mem_inst__abc_21378_n2104;
  wire w_mem_inst__abc_21378_n2105;
  wire w_mem_inst__abc_21378_n2106_1;
  wire w_mem_inst__abc_21378_n2107_1;
  wire w_mem_inst__abc_21378_n2108;
  wire w_mem_inst__abc_21378_n2109;
  wire w_mem_inst__abc_21378_n2110_1;
  wire w_mem_inst__abc_21378_n2111_1;
  wire w_mem_inst__abc_21378_n2112;
  wire w_mem_inst__abc_21378_n2113;
  wire w_mem_inst__abc_21378_n2114_1;
  wire w_mem_inst__abc_21378_n2115_1;
  wire w_mem_inst__abc_21378_n2116;
  wire w_mem_inst__abc_21378_n2117;
  wire w_mem_inst__abc_21378_n2118_1;
  wire w_mem_inst__abc_21378_n2119_1;
  wire w_mem_inst__abc_21378_n2120;
  wire w_mem_inst__abc_21378_n2121;
  wire w_mem_inst__abc_21378_n2122_1;
  wire w_mem_inst__abc_21378_n2123_1;
  wire w_mem_inst__abc_21378_n2124;
  wire w_mem_inst__abc_21378_n2125;
  wire w_mem_inst__abc_21378_n2126_1;
  wire w_mem_inst__abc_21378_n2127_1;
  wire w_mem_inst__abc_21378_n2128;
  wire w_mem_inst__abc_21378_n2129;
  wire w_mem_inst__abc_21378_n2130_1;
  wire w_mem_inst__abc_21378_n2131_1;
  wire w_mem_inst__abc_21378_n2132;
  wire w_mem_inst__abc_21378_n2133;
  wire w_mem_inst__abc_21378_n2134_1;
  wire w_mem_inst__abc_21378_n2135_1;
  wire w_mem_inst__abc_21378_n2136;
  wire w_mem_inst__abc_21378_n2137;
  wire w_mem_inst__abc_21378_n2138_1;
  wire w_mem_inst__abc_21378_n2139_1;
  wire w_mem_inst__abc_21378_n2140;
  wire w_mem_inst__abc_21378_n2141;
  wire w_mem_inst__abc_21378_n2142_1;
  wire w_mem_inst__abc_21378_n2144;
  wire w_mem_inst__abc_21378_n2145;
  wire w_mem_inst__abc_21378_n2146_1;
  wire w_mem_inst__abc_21378_n2147_1;
  wire w_mem_inst__abc_21378_n2148;
  wire w_mem_inst__abc_21378_n2149;
  wire w_mem_inst__abc_21378_n2150_1;
  wire w_mem_inst__abc_21378_n2151_1;
  wire w_mem_inst__abc_21378_n2152;
  wire w_mem_inst__abc_21378_n2153;
  wire w_mem_inst__abc_21378_n2154_1;
  wire w_mem_inst__abc_21378_n2155_1;
  wire w_mem_inst__abc_21378_n2156;
  wire w_mem_inst__abc_21378_n2157;
  wire w_mem_inst__abc_21378_n2158_1;
  wire w_mem_inst__abc_21378_n2159_1;
  wire w_mem_inst__abc_21378_n2160;
  wire w_mem_inst__abc_21378_n2161;
  wire w_mem_inst__abc_21378_n2162_1;
  wire w_mem_inst__abc_21378_n2163_1;
  wire w_mem_inst__abc_21378_n2164;
  wire w_mem_inst__abc_21378_n2165;
  wire w_mem_inst__abc_21378_n2166_1;
  wire w_mem_inst__abc_21378_n2167_1;
  wire w_mem_inst__abc_21378_n2168;
  wire w_mem_inst__abc_21378_n2169;
  wire w_mem_inst__abc_21378_n2170_1;
  wire w_mem_inst__abc_21378_n2171_1;
  wire w_mem_inst__abc_21378_n2172;
  wire w_mem_inst__abc_21378_n2173;
  wire w_mem_inst__abc_21378_n2174_1;
  wire w_mem_inst__abc_21378_n2175_1;
  wire w_mem_inst__abc_21378_n2176;
  wire w_mem_inst__abc_21378_n2177;
  wire w_mem_inst__abc_21378_n2178_1;
  wire w_mem_inst__abc_21378_n2179_1;
  wire w_mem_inst__abc_21378_n2180;
  wire w_mem_inst__abc_21378_n2181;
  wire w_mem_inst__abc_21378_n2182_1;
  wire w_mem_inst__abc_21378_n2183_1;
  wire w_mem_inst__abc_21378_n2184;
  wire w_mem_inst__abc_21378_n2185;
  wire w_mem_inst__abc_21378_n2186_1;
  wire w_mem_inst__abc_21378_n2187_1;
  wire w_mem_inst__abc_21378_n2188;
  wire w_mem_inst__abc_21378_n2189;
  wire w_mem_inst__abc_21378_n2190_1;
  wire w_mem_inst__abc_21378_n2192;
  wire w_mem_inst__abc_21378_n2193;
  wire w_mem_inst__abc_21378_n2194_1;
  wire w_mem_inst__abc_21378_n2195_1;
  wire w_mem_inst__abc_21378_n2196;
  wire w_mem_inst__abc_21378_n2197;
  wire w_mem_inst__abc_21378_n2198_1;
  wire w_mem_inst__abc_21378_n2199_1;
  wire w_mem_inst__abc_21378_n2200;
  wire w_mem_inst__abc_21378_n2201;
  wire w_mem_inst__abc_21378_n2202_1;
  wire w_mem_inst__abc_21378_n2203_1;
  wire w_mem_inst__abc_21378_n2204;
  wire w_mem_inst__abc_21378_n2205;
  wire w_mem_inst__abc_21378_n2206_1;
  wire w_mem_inst__abc_21378_n2207_1;
  wire w_mem_inst__abc_21378_n2208;
  wire w_mem_inst__abc_21378_n2209;
  wire w_mem_inst__abc_21378_n2210_1;
  wire w_mem_inst__abc_21378_n2211_1;
  wire w_mem_inst__abc_21378_n2212;
  wire w_mem_inst__abc_21378_n2213;
  wire w_mem_inst__abc_21378_n2214_1;
  wire w_mem_inst__abc_21378_n2215_1;
  wire w_mem_inst__abc_21378_n2216;
  wire w_mem_inst__abc_21378_n2217;
  wire w_mem_inst__abc_21378_n2218_1;
  wire w_mem_inst__abc_21378_n2219_1;
  wire w_mem_inst__abc_21378_n2220;
  wire w_mem_inst__abc_21378_n2221;
  wire w_mem_inst__abc_21378_n2222_1;
  wire w_mem_inst__abc_21378_n2223_1;
  wire w_mem_inst__abc_21378_n2224;
  wire w_mem_inst__abc_21378_n2225;
  wire w_mem_inst__abc_21378_n2226_1;
  wire w_mem_inst__abc_21378_n2227_1;
  wire w_mem_inst__abc_21378_n2228;
  wire w_mem_inst__abc_21378_n2229;
  wire w_mem_inst__abc_21378_n2230_1;
  wire w_mem_inst__abc_21378_n2231_1;
  wire w_mem_inst__abc_21378_n2232;
  wire w_mem_inst__abc_21378_n2233;
  wire w_mem_inst__abc_21378_n2234_1;
  wire w_mem_inst__abc_21378_n2235_1;
  wire w_mem_inst__abc_21378_n2236;
  wire w_mem_inst__abc_21378_n2237;
  wire w_mem_inst__abc_21378_n2238_1;
  wire w_mem_inst__abc_21378_n2240;
  wire w_mem_inst__abc_21378_n2241;
  wire w_mem_inst__abc_21378_n2242_1;
  wire w_mem_inst__abc_21378_n2243_1;
  wire w_mem_inst__abc_21378_n2244;
  wire w_mem_inst__abc_21378_n2245;
  wire w_mem_inst__abc_21378_n2246_1;
  wire w_mem_inst__abc_21378_n2247_1;
  wire w_mem_inst__abc_21378_n2248;
  wire w_mem_inst__abc_21378_n2249;
  wire w_mem_inst__abc_21378_n2250_1;
  wire w_mem_inst__abc_21378_n2251_1;
  wire w_mem_inst__abc_21378_n2252;
  wire w_mem_inst__abc_21378_n2253;
  wire w_mem_inst__abc_21378_n2254_1;
  wire w_mem_inst__abc_21378_n2255_1;
  wire w_mem_inst__abc_21378_n2256;
  wire w_mem_inst__abc_21378_n2257;
  wire w_mem_inst__abc_21378_n2258_1;
  wire w_mem_inst__abc_21378_n2259_1;
  wire w_mem_inst__abc_21378_n2260;
  wire w_mem_inst__abc_21378_n2261;
  wire w_mem_inst__abc_21378_n2262_1;
  wire w_mem_inst__abc_21378_n2263_1;
  wire w_mem_inst__abc_21378_n2264;
  wire w_mem_inst__abc_21378_n2265;
  wire w_mem_inst__abc_21378_n2266_1;
  wire w_mem_inst__abc_21378_n2267_1;
  wire w_mem_inst__abc_21378_n2268;
  wire w_mem_inst__abc_21378_n2269;
  wire w_mem_inst__abc_21378_n2270_1;
  wire w_mem_inst__abc_21378_n2271_1;
  wire w_mem_inst__abc_21378_n2272;
  wire w_mem_inst__abc_21378_n2273;
  wire w_mem_inst__abc_21378_n2274_1;
  wire w_mem_inst__abc_21378_n2275_1;
  wire w_mem_inst__abc_21378_n2276;
  wire w_mem_inst__abc_21378_n2277;
  wire w_mem_inst__abc_21378_n2278_1;
  wire w_mem_inst__abc_21378_n2279_1;
  wire w_mem_inst__abc_21378_n2280;
  wire w_mem_inst__abc_21378_n2281;
  wire w_mem_inst__abc_21378_n2282_1;
  wire w_mem_inst__abc_21378_n2283_1;
  wire w_mem_inst__abc_21378_n2284;
  wire w_mem_inst__abc_21378_n2285;
  wire w_mem_inst__abc_21378_n2286_1;
  wire w_mem_inst__abc_21378_n2288;
  wire w_mem_inst__abc_21378_n2289;
  wire w_mem_inst__abc_21378_n2290_1;
  wire w_mem_inst__abc_21378_n2291_1;
  wire w_mem_inst__abc_21378_n2292;
  wire w_mem_inst__abc_21378_n2293;
  wire w_mem_inst__abc_21378_n2294_1;
  wire w_mem_inst__abc_21378_n2295_1;
  wire w_mem_inst__abc_21378_n2296;
  wire w_mem_inst__abc_21378_n2297;
  wire w_mem_inst__abc_21378_n2298_1;
  wire w_mem_inst__abc_21378_n2299_1;
  wire w_mem_inst__abc_21378_n2300;
  wire w_mem_inst__abc_21378_n2301;
  wire w_mem_inst__abc_21378_n2302_1;
  wire w_mem_inst__abc_21378_n2303_1;
  wire w_mem_inst__abc_21378_n2304;
  wire w_mem_inst__abc_21378_n2305;
  wire w_mem_inst__abc_21378_n2306_1;
  wire w_mem_inst__abc_21378_n2307_1;
  wire w_mem_inst__abc_21378_n2308;
  wire w_mem_inst__abc_21378_n2309;
  wire w_mem_inst__abc_21378_n2310_1;
  wire w_mem_inst__abc_21378_n2311_1;
  wire w_mem_inst__abc_21378_n2312;
  wire w_mem_inst__abc_21378_n2313;
  wire w_mem_inst__abc_21378_n2314_1;
  wire w_mem_inst__abc_21378_n2315_1;
  wire w_mem_inst__abc_21378_n2316;
  wire w_mem_inst__abc_21378_n2317;
  wire w_mem_inst__abc_21378_n2318_1;
  wire w_mem_inst__abc_21378_n2319_1;
  wire w_mem_inst__abc_21378_n2320;
  wire w_mem_inst__abc_21378_n2321;
  wire w_mem_inst__abc_21378_n2322_1;
  wire w_mem_inst__abc_21378_n2323_1;
  wire w_mem_inst__abc_21378_n2324;
  wire w_mem_inst__abc_21378_n2325;
  wire w_mem_inst__abc_21378_n2326_1;
  wire w_mem_inst__abc_21378_n2327_1;
  wire w_mem_inst__abc_21378_n2328;
  wire w_mem_inst__abc_21378_n2329;
  wire w_mem_inst__abc_21378_n2330_1;
  wire w_mem_inst__abc_21378_n2331_1;
  wire w_mem_inst__abc_21378_n2332;
  wire w_mem_inst__abc_21378_n2333;
  wire w_mem_inst__abc_21378_n2334_1;
  wire w_mem_inst__abc_21378_n2336;
  wire w_mem_inst__abc_21378_n2337;
  wire w_mem_inst__abc_21378_n2338_1;
  wire w_mem_inst__abc_21378_n2339_1;
  wire w_mem_inst__abc_21378_n2340;
  wire w_mem_inst__abc_21378_n2341;
  wire w_mem_inst__abc_21378_n2342_1;
  wire w_mem_inst__abc_21378_n2343_1;
  wire w_mem_inst__abc_21378_n2344;
  wire w_mem_inst__abc_21378_n2345;
  wire w_mem_inst__abc_21378_n2346_1;
  wire w_mem_inst__abc_21378_n2347_1;
  wire w_mem_inst__abc_21378_n2348;
  wire w_mem_inst__abc_21378_n2349;
  wire w_mem_inst__abc_21378_n2350_1;
  wire w_mem_inst__abc_21378_n2351_1;
  wire w_mem_inst__abc_21378_n2352;
  wire w_mem_inst__abc_21378_n2353;
  wire w_mem_inst__abc_21378_n2354_1;
  wire w_mem_inst__abc_21378_n2355_1;
  wire w_mem_inst__abc_21378_n2356;
  wire w_mem_inst__abc_21378_n2357;
  wire w_mem_inst__abc_21378_n2358_1;
  wire w_mem_inst__abc_21378_n2359_1;
  wire w_mem_inst__abc_21378_n2360;
  wire w_mem_inst__abc_21378_n2361;
  wire w_mem_inst__abc_21378_n2362_1;
  wire w_mem_inst__abc_21378_n2363_1;
  wire w_mem_inst__abc_21378_n2364;
  wire w_mem_inst__abc_21378_n2365;
  wire w_mem_inst__abc_21378_n2366_1;
  wire w_mem_inst__abc_21378_n2367_1;
  wire w_mem_inst__abc_21378_n2368;
  wire w_mem_inst__abc_21378_n2369;
  wire w_mem_inst__abc_21378_n2370_1;
  wire w_mem_inst__abc_21378_n2371_1;
  wire w_mem_inst__abc_21378_n2372;
  wire w_mem_inst__abc_21378_n2373;
  wire w_mem_inst__abc_21378_n2374_1;
  wire w_mem_inst__abc_21378_n2375_1;
  wire w_mem_inst__abc_21378_n2376;
  wire w_mem_inst__abc_21378_n2377;
  wire w_mem_inst__abc_21378_n2378_1;
  wire w_mem_inst__abc_21378_n2379_1;
  wire w_mem_inst__abc_21378_n2380;
  wire w_mem_inst__abc_21378_n2381;
  wire w_mem_inst__abc_21378_n2382_1;
  wire w_mem_inst__abc_21378_n2384;
  wire w_mem_inst__abc_21378_n2385;
  wire w_mem_inst__abc_21378_n2386_1;
  wire w_mem_inst__abc_21378_n2387_1;
  wire w_mem_inst__abc_21378_n2388;
  wire w_mem_inst__abc_21378_n2389;
  wire w_mem_inst__abc_21378_n2390_1;
  wire w_mem_inst__abc_21378_n2391_1;
  wire w_mem_inst__abc_21378_n2392;
  wire w_mem_inst__abc_21378_n2393;
  wire w_mem_inst__abc_21378_n2394_1;
  wire w_mem_inst__abc_21378_n2395_1;
  wire w_mem_inst__abc_21378_n2396;
  wire w_mem_inst__abc_21378_n2397;
  wire w_mem_inst__abc_21378_n2398_1;
  wire w_mem_inst__abc_21378_n2399_1;
  wire w_mem_inst__abc_21378_n2400;
  wire w_mem_inst__abc_21378_n2401;
  wire w_mem_inst__abc_21378_n2402_1;
  wire w_mem_inst__abc_21378_n2403_1;
  wire w_mem_inst__abc_21378_n2404;
  wire w_mem_inst__abc_21378_n2405;
  wire w_mem_inst__abc_21378_n2406_1;
  wire w_mem_inst__abc_21378_n2407_1;
  wire w_mem_inst__abc_21378_n2408;
  wire w_mem_inst__abc_21378_n2409;
  wire w_mem_inst__abc_21378_n2410_1;
  wire w_mem_inst__abc_21378_n2411_1;
  wire w_mem_inst__abc_21378_n2412;
  wire w_mem_inst__abc_21378_n2413;
  wire w_mem_inst__abc_21378_n2414_1;
  wire w_mem_inst__abc_21378_n2415_1;
  wire w_mem_inst__abc_21378_n2416;
  wire w_mem_inst__abc_21378_n2417;
  wire w_mem_inst__abc_21378_n2418_1;
  wire w_mem_inst__abc_21378_n2419_1;
  wire w_mem_inst__abc_21378_n2420;
  wire w_mem_inst__abc_21378_n2421;
  wire w_mem_inst__abc_21378_n2422_1;
  wire w_mem_inst__abc_21378_n2423_1;
  wire w_mem_inst__abc_21378_n2424;
  wire w_mem_inst__abc_21378_n2425;
  wire w_mem_inst__abc_21378_n2426_1;
  wire w_mem_inst__abc_21378_n2427_1;
  wire w_mem_inst__abc_21378_n2428;
  wire w_mem_inst__abc_21378_n2429;
  wire w_mem_inst__abc_21378_n2430_1;
  wire w_mem_inst__abc_21378_n2432;
  wire w_mem_inst__abc_21378_n2433;
  wire w_mem_inst__abc_21378_n2434_1;
  wire w_mem_inst__abc_21378_n2435_1;
  wire w_mem_inst__abc_21378_n2436;
  wire w_mem_inst__abc_21378_n2437;
  wire w_mem_inst__abc_21378_n2438_1;
  wire w_mem_inst__abc_21378_n2439_1;
  wire w_mem_inst__abc_21378_n2440;
  wire w_mem_inst__abc_21378_n2441;
  wire w_mem_inst__abc_21378_n2442_1;
  wire w_mem_inst__abc_21378_n2443_1;
  wire w_mem_inst__abc_21378_n2444;
  wire w_mem_inst__abc_21378_n2445;
  wire w_mem_inst__abc_21378_n2446_1;
  wire w_mem_inst__abc_21378_n2447_1;
  wire w_mem_inst__abc_21378_n2448;
  wire w_mem_inst__abc_21378_n2449;
  wire w_mem_inst__abc_21378_n2450_1;
  wire w_mem_inst__abc_21378_n2451_1;
  wire w_mem_inst__abc_21378_n2452;
  wire w_mem_inst__abc_21378_n2453;
  wire w_mem_inst__abc_21378_n2454_1;
  wire w_mem_inst__abc_21378_n2455_1;
  wire w_mem_inst__abc_21378_n2456;
  wire w_mem_inst__abc_21378_n2457;
  wire w_mem_inst__abc_21378_n2458_1;
  wire w_mem_inst__abc_21378_n2459_1;
  wire w_mem_inst__abc_21378_n2460;
  wire w_mem_inst__abc_21378_n2461;
  wire w_mem_inst__abc_21378_n2462_1;
  wire w_mem_inst__abc_21378_n2463_1;
  wire w_mem_inst__abc_21378_n2464;
  wire w_mem_inst__abc_21378_n2465;
  wire w_mem_inst__abc_21378_n2466_1;
  wire w_mem_inst__abc_21378_n2467_1;
  wire w_mem_inst__abc_21378_n2468;
  wire w_mem_inst__abc_21378_n2469;
  wire w_mem_inst__abc_21378_n2470_1;
  wire w_mem_inst__abc_21378_n2471_1;
  wire w_mem_inst__abc_21378_n2472;
  wire w_mem_inst__abc_21378_n2473;
  wire w_mem_inst__abc_21378_n2474_1;
  wire w_mem_inst__abc_21378_n2475_1;
  wire w_mem_inst__abc_21378_n2476;
  wire w_mem_inst__abc_21378_n2477;
  wire w_mem_inst__abc_21378_n2478_1;
  wire w_mem_inst__abc_21378_n2480;
  wire w_mem_inst__abc_21378_n2481;
  wire w_mem_inst__abc_21378_n2482_1;
  wire w_mem_inst__abc_21378_n2483_1;
  wire w_mem_inst__abc_21378_n2484;
  wire w_mem_inst__abc_21378_n2485;
  wire w_mem_inst__abc_21378_n2486_1;
  wire w_mem_inst__abc_21378_n2487_1;
  wire w_mem_inst__abc_21378_n2488;
  wire w_mem_inst__abc_21378_n2489;
  wire w_mem_inst__abc_21378_n2490_1;
  wire w_mem_inst__abc_21378_n2491_1;
  wire w_mem_inst__abc_21378_n2492;
  wire w_mem_inst__abc_21378_n2493;
  wire w_mem_inst__abc_21378_n2494_1;
  wire w_mem_inst__abc_21378_n2495_1;
  wire w_mem_inst__abc_21378_n2496;
  wire w_mem_inst__abc_21378_n2497;
  wire w_mem_inst__abc_21378_n2498_1;
  wire w_mem_inst__abc_21378_n2499_1;
  wire w_mem_inst__abc_21378_n2500;
  wire w_mem_inst__abc_21378_n2501;
  wire w_mem_inst__abc_21378_n2502_1;
  wire w_mem_inst__abc_21378_n2503_1;
  wire w_mem_inst__abc_21378_n2504;
  wire w_mem_inst__abc_21378_n2505;
  wire w_mem_inst__abc_21378_n2506_1;
  wire w_mem_inst__abc_21378_n2507_1;
  wire w_mem_inst__abc_21378_n2508;
  wire w_mem_inst__abc_21378_n2509;
  wire w_mem_inst__abc_21378_n2510_1;
  wire w_mem_inst__abc_21378_n2511_1;
  wire w_mem_inst__abc_21378_n2512;
  wire w_mem_inst__abc_21378_n2513;
  wire w_mem_inst__abc_21378_n2514_1;
  wire w_mem_inst__abc_21378_n2515_1;
  wire w_mem_inst__abc_21378_n2516;
  wire w_mem_inst__abc_21378_n2517;
  wire w_mem_inst__abc_21378_n2518_1;
  wire w_mem_inst__abc_21378_n2519_1;
  wire w_mem_inst__abc_21378_n2520;
  wire w_mem_inst__abc_21378_n2521;
  wire w_mem_inst__abc_21378_n2522_1;
  wire w_mem_inst__abc_21378_n2523_1;
  wire w_mem_inst__abc_21378_n2524;
  wire w_mem_inst__abc_21378_n2525;
  wire w_mem_inst__abc_21378_n2526_1;
  wire w_mem_inst__abc_21378_n2528;
  wire w_mem_inst__abc_21378_n2529;
  wire w_mem_inst__abc_21378_n2530_1;
  wire w_mem_inst__abc_21378_n2531_1;
  wire w_mem_inst__abc_21378_n2532;
  wire w_mem_inst__abc_21378_n2533;
  wire w_mem_inst__abc_21378_n2534_1;
  wire w_mem_inst__abc_21378_n2535_1;
  wire w_mem_inst__abc_21378_n2536;
  wire w_mem_inst__abc_21378_n2537;
  wire w_mem_inst__abc_21378_n2538_1;
  wire w_mem_inst__abc_21378_n2539_1;
  wire w_mem_inst__abc_21378_n2540;
  wire w_mem_inst__abc_21378_n2541;
  wire w_mem_inst__abc_21378_n2542_1;
  wire w_mem_inst__abc_21378_n2543_1;
  wire w_mem_inst__abc_21378_n2544;
  wire w_mem_inst__abc_21378_n2545;
  wire w_mem_inst__abc_21378_n2546_1;
  wire w_mem_inst__abc_21378_n2547_1;
  wire w_mem_inst__abc_21378_n2548;
  wire w_mem_inst__abc_21378_n2549;
  wire w_mem_inst__abc_21378_n2550_1;
  wire w_mem_inst__abc_21378_n2551_1;
  wire w_mem_inst__abc_21378_n2552;
  wire w_mem_inst__abc_21378_n2553;
  wire w_mem_inst__abc_21378_n2554_1;
  wire w_mem_inst__abc_21378_n2555_1;
  wire w_mem_inst__abc_21378_n2556;
  wire w_mem_inst__abc_21378_n2557;
  wire w_mem_inst__abc_21378_n2558_1;
  wire w_mem_inst__abc_21378_n2559_1;
  wire w_mem_inst__abc_21378_n2560;
  wire w_mem_inst__abc_21378_n2561;
  wire w_mem_inst__abc_21378_n2562_1;
  wire w_mem_inst__abc_21378_n2563_1;
  wire w_mem_inst__abc_21378_n2564;
  wire w_mem_inst__abc_21378_n2565;
  wire w_mem_inst__abc_21378_n2566_1;
  wire w_mem_inst__abc_21378_n2567_1;
  wire w_mem_inst__abc_21378_n2568;
  wire w_mem_inst__abc_21378_n2569;
  wire w_mem_inst__abc_21378_n2570_1;
  wire w_mem_inst__abc_21378_n2571_1;
  wire w_mem_inst__abc_21378_n2572;
  wire w_mem_inst__abc_21378_n2573;
  wire w_mem_inst__abc_21378_n2574_1;
  wire w_mem_inst__abc_21378_n2576;
  wire w_mem_inst__abc_21378_n2577;
  wire w_mem_inst__abc_21378_n2578_1;
  wire w_mem_inst__abc_21378_n2579_1;
  wire w_mem_inst__abc_21378_n2580;
  wire w_mem_inst__abc_21378_n2581;
  wire w_mem_inst__abc_21378_n2582_1;
  wire w_mem_inst__abc_21378_n2583_1;
  wire w_mem_inst__abc_21378_n2584;
  wire w_mem_inst__abc_21378_n2585;
  wire w_mem_inst__abc_21378_n2586_1;
  wire w_mem_inst__abc_21378_n2587_1;
  wire w_mem_inst__abc_21378_n2588;
  wire w_mem_inst__abc_21378_n2589;
  wire w_mem_inst__abc_21378_n2590_1;
  wire w_mem_inst__abc_21378_n2591_1;
  wire w_mem_inst__abc_21378_n2592;
  wire w_mem_inst__abc_21378_n2593;
  wire w_mem_inst__abc_21378_n2594_1;
  wire w_mem_inst__abc_21378_n2595_1;
  wire w_mem_inst__abc_21378_n2596;
  wire w_mem_inst__abc_21378_n2597;
  wire w_mem_inst__abc_21378_n2598_1;
  wire w_mem_inst__abc_21378_n2599_1;
  wire w_mem_inst__abc_21378_n2600;
  wire w_mem_inst__abc_21378_n2601;
  wire w_mem_inst__abc_21378_n2602_1;
  wire w_mem_inst__abc_21378_n2603_1;
  wire w_mem_inst__abc_21378_n2604;
  wire w_mem_inst__abc_21378_n2605;
  wire w_mem_inst__abc_21378_n2606_1;
  wire w_mem_inst__abc_21378_n2607_1;
  wire w_mem_inst__abc_21378_n2608;
  wire w_mem_inst__abc_21378_n2609;
  wire w_mem_inst__abc_21378_n2610_1;
  wire w_mem_inst__abc_21378_n2611_1;
  wire w_mem_inst__abc_21378_n2612;
  wire w_mem_inst__abc_21378_n2613;
  wire w_mem_inst__abc_21378_n2614_1;
  wire w_mem_inst__abc_21378_n2615_1;
  wire w_mem_inst__abc_21378_n2616;
  wire w_mem_inst__abc_21378_n2617;
  wire w_mem_inst__abc_21378_n2618_1;
  wire w_mem_inst__abc_21378_n2619_1;
  wire w_mem_inst__abc_21378_n2620;
  wire w_mem_inst__abc_21378_n2621;
  wire w_mem_inst__abc_21378_n2622_1;
  wire w_mem_inst__abc_21378_n2624;
  wire w_mem_inst__abc_21378_n2625;
  wire w_mem_inst__abc_21378_n2626_1;
  wire w_mem_inst__abc_21378_n2627_1;
  wire w_mem_inst__abc_21378_n2628;
  wire w_mem_inst__abc_21378_n2629;
  wire w_mem_inst__abc_21378_n2630_1;
  wire w_mem_inst__abc_21378_n2631_1;
  wire w_mem_inst__abc_21378_n2632;
  wire w_mem_inst__abc_21378_n2633;
  wire w_mem_inst__abc_21378_n2634_1;
  wire w_mem_inst__abc_21378_n2635_1;
  wire w_mem_inst__abc_21378_n2636;
  wire w_mem_inst__abc_21378_n2637;
  wire w_mem_inst__abc_21378_n2638_1;
  wire w_mem_inst__abc_21378_n2639_1;
  wire w_mem_inst__abc_21378_n2640;
  wire w_mem_inst__abc_21378_n2641;
  wire w_mem_inst__abc_21378_n2642_1;
  wire w_mem_inst__abc_21378_n2643_1;
  wire w_mem_inst__abc_21378_n2644;
  wire w_mem_inst__abc_21378_n2645;
  wire w_mem_inst__abc_21378_n2646_1;
  wire w_mem_inst__abc_21378_n2647_1;
  wire w_mem_inst__abc_21378_n2648;
  wire w_mem_inst__abc_21378_n2649;
  wire w_mem_inst__abc_21378_n2650_1;
  wire w_mem_inst__abc_21378_n2651_1;
  wire w_mem_inst__abc_21378_n2652;
  wire w_mem_inst__abc_21378_n2653;
  wire w_mem_inst__abc_21378_n2654_1;
  wire w_mem_inst__abc_21378_n2655_1;
  wire w_mem_inst__abc_21378_n2656;
  wire w_mem_inst__abc_21378_n2657;
  wire w_mem_inst__abc_21378_n2658_1;
  wire w_mem_inst__abc_21378_n2659_1;
  wire w_mem_inst__abc_21378_n2660;
  wire w_mem_inst__abc_21378_n2661;
  wire w_mem_inst__abc_21378_n2662_1;
  wire w_mem_inst__abc_21378_n2663_1;
  wire w_mem_inst__abc_21378_n2664;
  wire w_mem_inst__abc_21378_n2665;
  wire w_mem_inst__abc_21378_n2666_1;
  wire w_mem_inst__abc_21378_n2667_1;
  wire w_mem_inst__abc_21378_n2668;
  wire w_mem_inst__abc_21378_n2669;
  wire w_mem_inst__abc_21378_n2670_1;
  wire w_mem_inst__abc_21378_n2672;
  wire w_mem_inst__abc_21378_n2673;
  wire w_mem_inst__abc_21378_n2674_1;
  wire w_mem_inst__abc_21378_n2675_1;
  wire w_mem_inst__abc_21378_n2676;
  wire w_mem_inst__abc_21378_n2677;
  wire w_mem_inst__abc_21378_n2678_1;
  wire w_mem_inst__abc_21378_n2679_1;
  wire w_mem_inst__abc_21378_n2680;
  wire w_mem_inst__abc_21378_n2681;
  wire w_mem_inst__abc_21378_n2682_1;
  wire w_mem_inst__abc_21378_n2683_1;
  wire w_mem_inst__abc_21378_n2684;
  wire w_mem_inst__abc_21378_n2685;
  wire w_mem_inst__abc_21378_n2686_1;
  wire w_mem_inst__abc_21378_n2687_1;
  wire w_mem_inst__abc_21378_n2688;
  wire w_mem_inst__abc_21378_n2689;
  wire w_mem_inst__abc_21378_n2690_1;
  wire w_mem_inst__abc_21378_n2691_1;
  wire w_mem_inst__abc_21378_n2692;
  wire w_mem_inst__abc_21378_n2693;
  wire w_mem_inst__abc_21378_n2694_1;
  wire w_mem_inst__abc_21378_n2695_1;
  wire w_mem_inst__abc_21378_n2696;
  wire w_mem_inst__abc_21378_n2697;
  wire w_mem_inst__abc_21378_n2698_1;
  wire w_mem_inst__abc_21378_n2699_1;
  wire w_mem_inst__abc_21378_n2700;
  wire w_mem_inst__abc_21378_n2701;
  wire w_mem_inst__abc_21378_n2702_1;
  wire w_mem_inst__abc_21378_n2703_1;
  wire w_mem_inst__abc_21378_n2704;
  wire w_mem_inst__abc_21378_n2705;
  wire w_mem_inst__abc_21378_n2706_1;
  wire w_mem_inst__abc_21378_n2707_1;
  wire w_mem_inst__abc_21378_n2708;
  wire w_mem_inst__abc_21378_n2709;
  wire w_mem_inst__abc_21378_n2710_1;
  wire w_mem_inst__abc_21378_n2711_1;
  wire w_mem_inst__abc_21378_n2712;
  wire w_mem_inst__abc_21378_n2713;
  wire w_mem_inst__abc_21378_n2714_1;
  wire w_mem_inst__abc_21378_n2715_1;
  wire w_mem_inst__abc_21378_n2716;
  wire w_mem_inst__abc_21378_n2717;
  wire w_mem_inst__abc_21378_n2718_1;
  wire w_mem_inst__abc_21378_n2720;
  wire w_mem_inst__abc_21378_n2721;
  wire w_mem_inst__abc_21378_n2722_1;
  wire w_mem_inst__abc_21378_n2723_1;
  wire w_mem_inst__abc_21378_n2724;
  wire w_mem_inst__abc_21378_n2725;
  wire w_mem_inst__abc_21378_n2726_1;
  wire w_mem_inst__abc_21378_n2727_1;
  wire w_mem_inst__abc_21378_n2728;
  wire w_mem_inst__abc_21378_n2729;
  wire w_mem_inst__abc_21378_n2730_1;
  wire w_mem_inst__abc_21378_n2731_1;
  wire w_mem_inst__abc_21378_n2732;
  wire w_mem_inst__abc_21378_n2733;
  wire w_mem_inst__abc_21378_n2734_1;
  wire w_mem_inst__abc_21378_n2735_1;
  wire w_mem_inst__abc_21378_n2736;
  wire w_mem_inst__abc_21378_n2737;
  wire w_mem_inst__abc_21378_n2738_1;
  wire w_mem_inst__abc_21378_n2739_1;
  wire w_mem_inst__abc_21378_n2740;
  wire w_mem_inst__abc_21378_n2741;
  wire w_mem_inst__abc_21378_n2742_1;
  wire w_mem_inst__abc_21378_n2743_1;
  wire w_mem_inst__abc_21378_n2744;
  wire w_mem_inst__abc_21378_n2745;
  wire w_mem_inst__abc_21378_n2746_1;
  wire w_mem_inst__abc_21378_n2747_1;
  wire w_mem_inst__abc_21378_n2748;
  wire w_mem_inst__abc_21378_n2749;
  wire w_mem_inst__abc_21378_n2750_1;
  wire w_mem_inst__abc_21378_n2751_1;
  wire w_mem_inst__abc_21378_n2752;
  wire w_mem_inst__abc_21378_n2753;
  wire w_mem_inst__abc_21378_n2754_1;
  wire w_mem_inst__abc_21378_n2755_1;
  wire w_mem_inst__abc_21378_n2756;
  wire w_mem_inst__abc_21378_n2757;
  wire w_mem_inst__abc_21378_n2758_1;
  wire w_mem_inst__abc_21378_n2759_1;
  wire w_mem_inst__abc_21378_n2760;
  wire w_mem_inst__abc_21378_n2761;
  wire w_mem_inst__abc_21378_n2762_1;
  wire w_mem_inst__abc_21378_n2763_1;
  wire w_mem_inst__abc_21378_n2764;
  wire w_mem_inst__abc_21378_n2765;
  wire w_mem_inst__abc_21378_n2766_1;
  wire w_mem_inst__abc_21378_n2768;
  wire w_mem_inst__abc_21378_n2769;
  wire w_mem_inst__abc_21378_n2770_1;
  wire w_mem_inst__abc_21378_n2771_1;
  wire w_mem_inst__abc_21378_n2772;
  wire w_mem_inst__abc_21378_n2773;
  wire w_mem_inst__abc_21378_n2774_1;
  wire w_mem_inst__abc_21378_n2775_1;
  wire w_mem_inst__abc_21378_n2776;
  wire w_mem_inst__abc_21378_n2777;
  wire w_mem_inst__abc_21378_n2778_1;
  wire w_mem_inst__abc_21378_n2779_1;
  wire w_mem_inst__abc_21378_n2780;
  wire w_mem_inst__abc_21378_n2781;
  wire w_mem_inst__abc_21378_n2782_1;
  wire w_mem_inst__abc_21378_n2783_1;
  wire w_mem_inst__abc_21378_n2784;
  wire w_mem_inst__abc_21378_n2785;
  wire w_mem_inst__abc_21378_n2786_1;
  wire w_mem_inst__abc_21378_n2787_1;
  wire w_mem_inst__abc_21378_n2788;
  wire w_mem_inst__abc_21378_n2789;
  wire w_mem_inst__abc_21378_n2790_1;
  wire w_mem_inst__abc_21378_n2791_1;
  wire w_mem_inst__abc_21378_n2792;
  wire w_mem_inst__abc_21378_n2793;
  wire w_mem_inst__abc_21378_n2794_1;
  wire w_mem_inst__abc_21378_n2795_1;
  wire w_mem_inst__abc_21378_n2796;
  wire w_mem_inst__abc_21378_n2797;
  wire w_mem_inst__abc_21378_n2798_1;
  wire w_mem_inst__abc_21378_n2799_1;
  wire w_mem_inst__abc_21378_n2800;
  wire w_mem_inst__abc_21378_n2801;
  wire w_mem_inst__abc_21378_n2802_1;
  wire w_mem_inst__abc_21378_n2803_1;
  wire w_mem_inst__abc_21378_n2804;
  wire w_mem_inst__abc_21378_n2805;
  wire w_mem_inst__abc_21378_n2806_1;
  wire w_mem_inst__abc_21378_n2807_1;
  wire w_mem_inst__abc_21378_n2808;
  wire w_mem_inst__abc_21378_n2809;
  wire w_mem_inst__abc_21378_n2810_1;
  wire w_mem_inst__abc_21378_n2811_1;
  wire w_mem_inst__abc_21378_n2812;
  wire w_mem_inst__abc_21378_n2813;
  wire w_mem_inst__abc_21378_n2814_1;
  wire w_mem_inst__abc_21378_n2816;
  wire w_mem_inst__abc_21378_n2817;
  wire w_mem_inst__abc_21378_n2818_1;
  wire w_mem_inst__abc_21378_n2819_1;
  wire w_mem_inst__abc_21378_n2820;
  wire w_mem_inst__abc_21378_n2821;
  wire w_mem_inst__abc_21378_n2822_1;
  wire w_mem_inst__abc_21378_n2823_1;
  wire w_mem_inst__abc_21378_n2824;
  wire w_mem_inst__abc_21378_n2825;
  wire w_mem_inst__abc_21378_n2826_1;
  wire w_mem_inst__abc_21378_n2827_1;
  wire w_mem_inst__abc_21378_n2828;
  wire w_mem_inst__abc_21378_n2829;
  wire w_mem_inst__abc_21378_n2830_1;
  wire w_mem_inst__abc_21378_n2831_1;
  wire w_mem_inst__abc_21378_n2832;
  wire w_mem_inst__abc_21378_n2833;
  wire w_mem_inst__abc_21378_n2834_1;
  wire w_mem_inst__abc_21378_n2835_1;
  wire w_mem_inst__abc_21378_n2836;
  wire w_mem_inst__abc_21378_n2837;
  wire w_mem_inst__abc_21378_n2838_1;
  wire w_mem_inst__abc_21378_n2839_1;
  wire w_mem_inst__abc_21378_n2840;
  wire w_mem_inst__abc_21378_n2841;
  wire w_mem_inst__abc_21378_n2842_1;
  wire w_mem_inst__abc_21378_n2843_1;
  wire w_mem_inst__abc_21378_n2844;
  wire w_mem_inst__abc_21378_n2845;
  wire w_mem_inst__abc_21378_n2846_1;
  wire w_mem_inst__abc_21378_n2847_1;
  wire w_mem_inst__abc_21378_n2848;
  wire w_mem_inst__abc_21378_n2849;
  wire w_mem_inst__abc_21378_n2850_1;
  wire w_mem_inst__abc_21378_n2851_1;
  wire w_mem_inst__abc_21378_n2852;
  wire w_mem_inst__abc_21378_n2853;
  wire w_mem_inst__abc_21378_n2854_1;
  wire w_mem_inst__abc_21378_n2855_1;
  wire w_mem_inst__abc_21378_n2856;
  wire w_mem_inst__abc_21378_n2857;
  wire w_mem_inst__abc_21378_n2858_1;
  wire w_mem_inst__abc_21378_n2859_1;
  wire w_mem_inst__abc_21378_n2860;
  wire w_mem_inst__abc_21378_n2861;
  wire w_mem_inst__abc_21378_n2862_1;
  wire w_mem_inst__abc_21378_n2864;
  wire w_mem_inst__abc_21378_n2865;
  wire w_mem_inst__abc_21378_n2866_1;
  wire w_mem_inst__abc_21378_n2867_1;
  wire w_mem_inst__abc_21378_n2868;
  wire w_mem_inst__abc_21378_n2869;
  wire w_mem_inst__abc_21378_n2870_1;
  wire w_mem_inst__abc_21378_n2871_1;
  wire w_mem_inst__abc_21378_n2872;
  wire w_mem_inst__abc_21378_n2873;
  wire w_mem_inst__abc_21378_n2874_1;
  wire w_mem_inst__abc_21378_n2875_1;
  wire w_mem_inst__abc_21378_n2876;
  wire w_mem_inst__abc_21378_n2877;
  wire w_mem_inst__abc_21378_n2878_1;
  wire w_mem_inst__abc_21378_n2879_1;
  wire w_mem_inst__abc_21378_n2880;
  wire w_mem_inst__abc_21378_n2881;
  wire w_mem_inst__abc_21378_n2882_1;
  wire w_mem_inst__abc_21378_n2883_1;
  wire w_mem_inst__abc_21378_n2884;
  wire w_mem_inst__abc_21378_n2885;
  wire w_mem_inst__abc_21378_n2886_1;
  wire w_mem_inst__abc_21378_n2887_1;
  wire w_mem_inst__abc_21378_n2888;
  wire w_mem_inst__abc_21378_n2889;
  wire w_mem_inst__abc_21378_n2890_1;
  wire w_mem_inst__abc_21378_n2891_1;
  wire w_mem_inst__abc_21378_n2892;
  wire w_mem_inst__abc_21378_n2893;
  wire w_mem_inst__abc_21378_n2894_1;
  wire w_mem_inst__abc_21378_n2895_1;
  wire w_mem_inst__abc_21378_n2896;
  wire w_mem_inst__abc_21378_n2897;
  wire w_mem_inst__abc_21378_n2898_1;
  wire w_mem_inst__abc_21378_n2899_1;
  wire w_mem_inst__abc_21378_n2900;
  wire w_mem_inst__abc_21378_n2901;
  wire w_mem_inst__abc_21378_n2902_1;
  wire w_mem_inst__abc_21378_n2903_1;
  wire w_mem_inst__abc_21378_n2904;
  wire w_mem_inst__abc_21378_n2905;
  wire w_mem_inst__abc_21378_n2906_1;
  wire w_mem_inst__abc_21378_n2907_1;
  wire w_mem_inst__abc_21378_n2908;
  wire w_mem_inst__abc_21378_n2909;
  wire w_mem_inst__abc_21378_n2910_1;
  wire w_mem_inst__abc_21378_n2912;
  wire w_mem_inst__abc_21378_n2913;
  wire w_mem_inst__abc_21378_n2914_1;
  wire w_mem_inst__abc_21378_n2915_1;
  wire w_mem_inst__abc_21378_n2916;
  wire w_mem_inst__abc_21378_n2917;
  wire w_mem_inst__abc_21378_n2918_1;
  wire w_mem_inst__abc_21378_n2919_1;
  wire w_mem_inst__abc_21378_n2920;
  wire w_mem_inst__abc_21378_n2921;
  wire w_mem_inst__abc_21378_n2922_1;
  wire w_mem_inst__abc_21378_n2923_1;
  wire w_mem_inst__abc_21378_n2924;
  wire w_mem_inst__abc_21378_n2925;
  wire w_mem_inst__abc_21378_n2926_1;
  wire w_mem_inst__abc_21378_n2927_1;
  wire w_mem_inst__abc_21378_n2928;
  wire w_mem_inst__abc_21378_n2929;
  wire w_mem_inst__abc_21378_n2930_1;
  wire w_mem_inst__abc_21378_n2931_1;
  wire w_mem_inst__abc_21378_n2932;
  wire w_mem_inst__abc_21378_n2933;
  wire w_mem_inst__abc_21378_n2934_1;
  wire w_mem_inst__abc_21378_n2935_1;
  wire w_mem_inst__abc_21378_n2936;
  wire w_mem_inst__abc_21378_n2937;
  wire w_mem_inst__abc_21378_n2938_1;
  wire w_mem_inst__abc_21378_n2939_1;
  wire w_mem_inst__abc_21378_n2940;
  wire w_mem_inst__abc_21378_n2941;
  wire w_mem_inst__abc_21378_n2942_1;
  wire w_mem_inst__abc_21378_n2943_1;
  wire w_mem_inst__abc_21378_n2944;
  wire w_mem_inst__abc_21378_n2945;
  wire w_mem_inst__abc_21378_n2946_1;
  wire w_mem_inst__abc_21378_n2947_1;
  wire w_mem_inst__abc_21378_n2948;
  wire w_mem_inst__abc_21378_n2949;
  wire w_mem_inst__abc_21378_n2950_1;
  wire w_mem_inst__abc_21378_n2951_1;
  wire w_mem_inst__abc_21378_n2952;
  wire w_mem_inst__abc_21378_n2953;
  wire w_mem_inst__abc_21378_n2954_1;
  wire w_mem_inst__abc_21378_n2955_1;
  wire w_mem_inst__abc_21378_n2956;
  wire w_mem_inst__abc_21378_n2957;
  wire w_mem_inst__abc_21378_n2958_1;
  wire w_mem_inst__abc_21378_n2960;
  wire w_mem_inst__abc_21378_n2961;
  wire w_mem_inst__abc_21378_n2962_1;
  wire w_mem_inst__abc_21378_n2963_1;
  wire w_mem_inst__abc_21378_n2964;
  wire w_mem_inst__abc_21378_n2965;
  wire w_mem_inst__abc_21378_n2966_1;
  wire w_mem_inst__abc_21378_n2967_1;
  wire w_mem_inst__abc_21378_n2968;
  wire w_mem_inst__abc_21378_n2969;
  wire w_mem_inst__abc_21378_n2970_1;
  wire w_mem_inst__abc_21378_n2971_1;
  wire w_mem_inst__abc_21378_n2972;
  wire w_mem_inst__abc_21378_n2973;
  wire w_mem_inst__abc_21378_n2974_1;
  wire w_mem_inst__abc_21378_n2975_1;
  wire w_mem_inst__abc_21378_n2976;
  wire w_mem_inst__abc_21378_n2977;
  wire w_mem_inst__abc_21378_n2978_1;
  wire w_mem_inst__abc_21378_n2979_1;
  wire w_mem_inst__abc_21378_n2980;
  wire w_mem_inst__abc_21378_n2981;
  wire w_mem_inst__abc_21378_n2982_1;
  wire w_mem_inst__abc_21378_n2983_1;
  wire w_mem_inst__abc_21378_n2984;
  wire w_mem_inst__abc_21378_n2985;
  wire w_mem_inst__abc_21378_n2986_1;
  wire w_mem_inst__abc_21378_n2987_1;
  wire w_mem_inst__abc_21378_n2988;
  wire w_mem_inst__abc_21378_n2989;
  wire w_mem_inst__abc_21378_n2990_1;
  wire w_mem_inst__abc_21378_n2991_1;
  wire w_mem_inst__abc_21378_n2992;
  wire w_mem_inst__abc_21378_n2993;
  wire w_mem_inst__abc_21378_n2994_1;
  wire w_mem_inst__abc_21378_n2995_1;
  wire w_mem_inst__abc_21378_n2996;
  wire w_mem_inst__abc_21378_n2997;
  wire w_mem_inst__abc_21378_n2998_1;
  wire w_mem_inst__abc_21378_n2999_1;
  wire w_mem_inst__abc_21378_n3000;
  wire w_mem_inst__abc_21378_n3001;
  wire w_mem_inst__abc_21378_n3002_1;
  wire w_mem_inst__abc_21378_n3003_1;
  wire w_mem_inst__abc_21378_n3004;
  wire w_mem_inst__abc_21378_n3005;
  wire w_mem_inst__abc_21378_n3006_1;
  wire w_mem_inst__abc_21378_n3008;
  wire w_mem_inst__abc_21378_n3009;
  wire w_mem_inst__abc_21378_n3010_1;
  wire w_mem_inst__abc_21378_n3011_1;
  wire w_mem_inst__abc_21378_n3012;
  wire w_mem_inst__abc_21378_n3013;
  wire w_mem_inst__abc_21378_n3014_1;
  wire w_mem_inst__abc_21378_n3015_1;
  wire w_mem_inst__abc_21378_n3016;
  wire w_mem_inst__abc_21378_n3017;
  wire w_mem_inst__abc_21378_n3018_1;
  wire w_mem_inst__abc_21378_n3019_1;
  wire w_mem_inst__abc_21378_n3020;
  wire w_mem_inst__abc_21378_n3021;
  wire w_mem_inst__abc_21378_n3022_1;
  wire w_mem_inst__abc_21378_n3023_1;
  wire w_mem_inst__abc_21378_n3024;
  wire w_mem_inst__abc_21378_n3025;
  wire w_mem_inst__abc_21378_n3026_1;
  wire w_mem_inst__abc_21378_n3027_1;
  wire w_mem_inst__abc_21378_n3028;
  wire w_mem_inst__abc_21378_n3029;
  wire w_mem_inst__abc_21378_n3030_1;
  wire w_mem_inst__abc_21378_n3031_1;
  wire w_mem_inst__abc_21378_n3032;
  wire w_mem_inst__abc_21378_n3033;
  wire w_mem_inst__abc_21378_n3034_1;
  wire w_mem_inst__abc_21378_n3035_1;
  wire w_mem_inst__abc_21378_n3036;
  wire w_mem_inst__abc_21378_n3037;
  wire w_mem_inst__abc_21378_n3038_1;
  wire w_mem_inst__abc_21378_n3039_1;
  wire w_mem_inst__abc_21378_n3040;
  wire w_mem_inst__abc_21378_n3041;
  wire w_mem_inst__abc_21378_n3042_1;
  wire w_mem_inst__abc_21378_n3043_1;
  wire w_mem_inst__abc_21378_n3044;
  wire w_mem_inst__abc_21378_n3045;
  wire w_mem_inst__abc_21378_n3046_1;
  wire w_mem_inst__abc_21378_n3047_1;
  wire w_mem_inst__abc_21378_n3048;
  wire w_mem_inst__abc_21378_n3049;
  wire w_mem_inst__abc_21378_n3050_1;
  wire w_mem_inst__abc_21378_n3051_1;
  wire w_mem_inst__abc_21378_n3052;
  wire w_mem_inst__abc_21378_n3053;
  wire w_mem_inst__abc_21378_n3054_1;
  wire w_mem_inst__abc_21378_n3056;
  wire w_mem_inst__abc_21378_n3057;
  wire w_mem_inst__abc_21378_n3058_1;
  wire w_mem_inst__abc_21378_n3059_1;
  wire w_mem_inst__abc_21378_n3060;
  wire w_mem_inst__abc_21378_n3061;
  wire w_mem_inst__abc_21378_n3062_1;
  wire w_mem_inst__abc_21378_n3063_1;
  wire w_mem_inst__abc_21378_n3064;
  wire w_mem_inst__abc_21378_n3065;
  wire w_mem_inst__abc_21378_n3066_1;
  wire w_mem_inst__abc_21378_n3067_1;
  wire w_mem_inst__abc_21378_n3068;
  wire w_mem_inst__abc_21378_n3069;
  wire w_mem_inst__abc_21378_n3070_1;
  wire w_mem_inst__abc_21378_n3071_1;
  wire w_mem_inst__abc_21378_n3072;
  wire w_mem_inst__abc_21378_n3073;
  wire w_mem_inst__abc_21378_n3074_1;
  wire w_mem_inst__abc_21378_n3075_1;
  wire w_mem_inst__abc_21378_n3076;
  wire w_mem_inst__abc_21378_n3077;
  wire w_mem_inst__abc_21378_n3078_1;
  wire w_mem_inst__abc_21378_n3079_1;
  wire w_mem_inst__abc_21378_n3080;
  wire w_mem_inst__abc_21378_n3081;
  wire w_mem_inst__abc_21378_n3082_1;
  wire w_mem_inst__abc_21378_n3083_1;
  wire w_mem_inst__abc_21378_n3084;
  wire w_mem_inst__abc_21378_n3085;
  wire w_mem_inst__abc_21378_n3086_1;
  wire w_mem_inst__abc_21378_n3087_1;
  wire w_mem_inst__abc_21378_n3088;
  wire w_mem_inst__abc_21378_n3089;
  wire w_mem_inst__abc_21378_n3090_1;
  wire w_mem_inst__abc_21378_n3091_1;
  wire w_mem_inst__abc_21378_n3092;
  wire w_mem_inst__abc_21378_n3093;
  wire w_mem_inst__abc_21378_n3094_1;
  wire w_mem_inst__abc_21378_n3095_1;
  wire w_mem_inst__abc_21378_n3096;
  wire w_mem_inst__abc_21378_n3097;
  wire w_mem_inst__abc_21378_n3098_1;
  wire w_mem_inst__abc_21378_n3099_1;
  wire w_mem_inst__abc_21378_n3100;
  wire w_mem_inst__abc_21378_n3101;
  wire w_mem_inst__abc_21378_n3102_1;
  wire w_mem_inst__abc_21378_n3104;
  wire w_mem_inst__abc_21378_n3105;
  wire w_mem_inst__abc_21378_n3106_1;
  wire w_mem_inst__abc_21378_n3107_1;
  wire w_mem_inst__abc_21378_n3108;
  wire w_mem_inst__abc_21378_n3109;
  wire w_mem_inst__abc_21378_n3110_1;
  wire w_mem_inst__abc_21378_n3111_1;
  wire w_mem_inst__abc_21378_n3112;
  wire w_mem_inst__abc_21378_n3113;
  wire w_mem_inst__abc_21378_n3114_1;
  wire w_mem_inst__abc_21378_n3115_1;
  wire w_mem_inst__abc_21378_n3116;
  wire w_mem_inst__abc_21378_n3117;
  wire w_mem_inst__abc_21378_n3118_1;
  wire w_mem_inst__abc_21378_n3119_1;
  wire w_mem_inst__abc_21378_n3120;
  wire w_mem_inst__abc_21378_n3121;
  wire w_mem_inst__abc_21378_n3122_1;
  wire w_mem_inst__abc_21378_n3123_1;
  wire w_mem_inst__abc_21378_n3124;
  wire w_mem_inst__abc_21378_n3125;
  wire w_mem_inst__abc_21378_n3126_1;
  wire w_mem_inst__abc_21378_n3127_1;
  wire w_mem_inst__abc_21378_n3128;
  wire w_mem_inst__abc_21378_n3129;
  wire w_mem_inst__abc_21378_n3130_1;
  wire w_mem_inst__abc_21378_n3131_1;
  wire w_mem_inst__abc_21378_n3132;
  wire w_mem_inst__abc_21378_n3133;
  wire w_mem_inst__abc_21378_n3134_1;
  wire w_mem_inst__abc_21378_n3135_1;
  wire w_mem_inst__abc_21378_n3136;
  wire w_mem_inst__abc_21378_n3137;
  wire w_mem_inst__abc_21378_n3138_1;
  wire w_mem_inst__abc_21378_n3139_1;
  wire w_mem_inst__abc_21378_n3140;
  wire w_mem_inst__abc_21378_n3141;
  wire w_mem_inst__abc_21378_n3142_1;
  wire w_mem_inst__abc_21378_n3143_1;
  wire w_mem_inst__abc_21378_n3144;
  wire w_mem_inst__abc_21378_n3145;
  wire w_mem_inst__abc_21378_n3146_1;
  wire w_mem_inst__abc_21378_n3147_1;
  wire w_mem_inst__abc_21378_n3148;
  wire w_mem_inst__abc_21378_n3149;
  wire w_mem_inst__abc_21378_n3150_1;
  wire w_mem_inst__abc_21378_n3152;
  wire w_mem_inst__abc_21378_n3152_bF_buf0;
  wire w_mem_inst__abc_21378_n3152_bF_buf1;
  wire w_mem_inst__abc_21378_n3152_bF_buf10;
  wire w_mem_inst__abc_21378_n3152_bF_buf11;
  wire w_mem_inst__abc_21378_n3152_bF_buf12;
  wire w_mem_inst__abc_21378_n3152_bF_buf13;
  wire w_mem_inst__abc_21378_n3152_bF_buf14;
  wire w_mem_inst__abc_21378_n3152_bF_buf15;
  wire w_mem_inst__abc_21378_n3152_bF_buf16;
  wire w_mem_inst__abc_21378_n3152_bF_buf17;
  wire w_mem_inst__abc_21378_n3152_bF_buf18;
  wire w_mem_inst__abc_21378_n3152_bF_buf19;
  wire w_mem_inst__abc_21378_n3152_bF_buf2;
  wire w_mem_inst__abc_21378_n3152_bF_buf20;
  wire w_mem_inst__abc_21378_n3152_bF_buf21;
  wire w_mem_inst__abc_21378_n3152_bF_buf22;
  wire w_mem_inst__abc_21378_n3152_bF_buf23;
  wire w_mem_inst__abc_21378_n3152_bF_buf24;
  wire w_mem_inst__abc_21378_n3152_bF_buf25;
  wire w_mem_inst__abc_21378_n3152_bF_buf26;
  wire w_mem_inst__abc_21378_n3152_bF_buf27;
  wire w_mem_inst__abc_21378_n3152_bF_buf28;
  wire w_mem_inst__abc_21378_n3152_bF_buf29;
  wire w_mem_inst__abc_21378_n3152_bF_buf3;
  wire w_mem_inst__abc_21378_n3152_bF_buf30;
  wire w_mem_inst__abc_21378_n3152_bF_buf31;
  wire w_mem_inst__abc_21378_n3152_bF_buf32;
  wire w_mem_inst__abc_21378_n3152_bF_buf33;
  wire w_mem_inst__abc_21378_n3152_bF_buf34;
  wire w_mem_inst__abc_21378_n3152_bF_buf35;
  wire w_mem_inst__abc_21378_n3152_bF_buf36;
  wire w_mem_inst__abc_21378_n3152_bF_buf37;
  wire w_mem_inst__abc_21378_n3152_bF_buf38;
  wire w_mem_inst__abc_21378_n3152_bF_buf39;
  wire w_mem_inst__abc_21378_n3152_bF_buf4;
  wire w_mem_inst__abc_21378_n3152_bF_buf40;
  wire w_mem_inst__abc_21378_n3152_bF_buf41;
  wire w_mem_inst__abc_21378_n3152_bF_buf42;
  wire w_mem_inst__abc_21378_n3152_bF_buf43;
  wire w_mem_inst__abc_21378_n3152_bF_buf44;
  wire w_mem_inst__abc_21378_n3152_bF_buf45;
  wire w_mem_inst__abc_21378_n3152_bF_buf46;
  wire w_mem_inst__abc_21378_n3152_bF_buf47;
  wire w_mem_inst__abc_21378_n3152_bF_buf48;
  wire w_mem_inst__abc_21378_n3152_bF_buf49;
  wire w_mem_inst__abc_21378_n3152_bF_buf5;
  wire w_mem_inst__abc_21378_n3152_bF_buf50;
  wire w_mem_inst__abc_21378_n3152_bF_buf51;
  wire w_mem_inst__abc_21378_n3152_bF_buf52;
  wire w_mem_inst__abc_21378_n3152_bF_buf53;
  wire w_mem_inst__abc_21378_n3152_bF_buf54;
  wire w_mem_inst__abc_21378_n3152_bF_buf55;
  wire w_mem_inst__abc_21378_n3152_bF_buf56;
  wire w_mem_inst__abc_21378_n3152_bF_buf57;
  wire w_mem_inst__abc_21378_n3152_bF_buf58;
  wire w_mem_inst__abc_21378_n3152_bF_buf59;
  wire w_mem_inst__abc_21378_n3152_bF_buf6;
  wire w_mem_inst__abc_21378_n3152_bF_buf60;
  wire w_mem_inst__abc_21378_n3152_bF_buf61;
  wire w_mem_inst__abc_21378_n3152_bF_buf62;
  wire w_mem_inst__abc_21378_n3152_bF_buf63;
  wire w_mem_inst__abc_21378_n3152_bF_buf7;
  wire w_mem_inst__abc_21378_n3152_bF_buf8;
  wire w_mem_inst__abc_21378_n3152_bF_buf9;
  wire w_mem_inst__abc_21378_n3152_hier0_bF_buf0;
  wire w_mem_inst__abc_21378_n3152_hier0_bF_buf1;
  wire w_mem_inst__abc_21378_n3152_hier0_bF_buf2;
  wire w_mem_inst__abc_21378_n3152_hier0_bF_buf3;
  wire w_mem_inst__abc_21378_n3152_hier0_bF_buf4;
  wire w_mem_inst__abc_21378_n3152_hier0_bF_buf5;
  wire w_mem_inst__abc_21378_n3152_hier0_bF_buf6;
  wire w_mem_inst__abc_21378_n3152_hier0_bF_buf7;
  wire w_mem_inst__abc_21378_n3153;
  wire w_mem_inst__abc_21378_n3154_1;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf0;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf1;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf10;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf11;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf12;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf13;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf14;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf15;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf16;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf17;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf18;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf19;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf2;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf20;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf21;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf22;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf23;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf24;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf25;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf26;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf27;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf28;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf29;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf3;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf30;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf31;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf32;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf33;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf34;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf35;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf36;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf37;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf38;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf39;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf4;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf40;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf41;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf42;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf43;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf44;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf45;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf46;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf47;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf48;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf49;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf5;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf50;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf51;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf52;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf53;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf54;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf55;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf56;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf57;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf58;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf59;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf6;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf60;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf61;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf62;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf63;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf7;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf8;
  wire w_mem_inst__abc_21378_n3154_1_bF_buf9;
  wire w_mem_inst__abc_21378_n3154_1_hier0_bF_buf0;
  wire w_mem_inst__abc_21378_n3154_1_hier0_bF_buf1;
  wire w_mem_inst__abc_21378_n3154_1_hier0_bF_buf2;
  wire w_mem_inst__abc_21378_n3154_1_hier0_bF_buf3;
  wire w_mem_inst__abc_21378_n3154_1_hier0_bF_buf4;
  wire w_mem_inst__abc_21378_n3154_1_hier0_bF_buf5;
  wire w_mem_inst__abc_21378_n3154_1_hier0_bF_buf6;
  wire w_mem_inst__abc_21378_n3154_1_hier0_bF_buf7;
  wire w_mem_inst__abc_21378_n3155_1;
  wire w_mem_inst__abc_21378_n3156;
  wire w_mem_inst__abc_21378_n3156_bF_buf0;
  wire w_mem_inst__abc_21378_n3156_bF_buf1;
  wire w_mem_inst__abc_21378_n3156_bF_buf2;
  wire w_mem_inst__abc_21378_n3156_bF_buf3;
  wire w_mem_inst__abc_21378_n3156_bF_buf4;
  wire w_mem_inst__abc_21378_n3157;
  wire w_mem_inst__abc_21378_n3158_1;
  wire w_mem_inst__abc_21378_n3159_1;
  wire w_mem_inst__abc_21378_n3161;
  wire w_mem_inst__abc_21378_n3162_1;
  wire w_mem_inst__abc_21378_n3163_1;
  wire w_mem_inst__abc_21378_n3164;
  wire w_mem_inst__abc_21378_n3165;
  wire w_mem_inst__abc_21378_n3167_1;
  wire w_mem_inst__abc_21378_n3168;
  wire w_mem_inst__abc_21378_n3169;
  wire w_mem_inst__abc_21378_n3170_1;
  wire w_mem_inst__abc_21378_n3171_1;
  wire w_mem_inst__abc_21378_n3173;
  wire w_mem_inst__abc_21378_n3174_1;
  wire w_mem_inst__abc_21378_n3175_1;
  wire w_mem_inst__abc_21378_n3176;
  wire w_mem_inst__abc_21378_n3177;
  wire w_mem_inst__abc_21378_n3179_1;
  wire w_mem_inst__abc_21378_n3180;
  wire w_mem_inst__abc_21378_n3181;
  wire w_mem_inst__abc_21378_n3182_1;
  wire w_mem_inst__abc_21378_n3183_1;
  wire w_mem_inst__abc_21378_n3185;
  wire w_mem_inst__abc_21378_n3186_1;
  wire w_mem_inst__abc_21378_n3187_1;
  wire w_mem_inst__abc_21378_n3188;
  wire w_mem_inst__abc_21378_n3189;
  wire w_mem_inst__abc_21378_n3191_1;
  wire w_mem_inst__abc_21378_n3192;
  wire w_mem_inst__abc_21378_n3193;
  wire w_mem_inst__abc_21378_n3194_1;
  wire w_mem_inst__abc_21378_n3195_1;
  wire w_mem_inst__abc_21378_n3197;
  wire w_mem_inst__abc_21378_n3198_1;
  wire w_mem_inst__abc_21378_n3199_1;
  wire w_mem_inst__abc_21378_n3200;
  wire w_mem_inst__abc_21378_n3201;
  wire w_mem_inst__abc_21378_n3203_1;
  wire w_mem_inst__abc_21378_n3204;
  wire w_mem_inst__abc_21378_n3205;
  wire w_mem_inst__abc_21378_n3206_1;
  wire w_mem_inst__abc_21378_n3207_1;
  wire w_mem_inst__abc_21378_n3209;
  wire w_mem_inst__abc_21378_n3210_1;
  wire w_mem_inst__abc_21378_n3211_1;
  wire w_mem_inst__abc_21378_n3212;
  wire w_mem_inst__abc_21378_n3213;
  wire w_mem_inst__abc_21378_n3215_1;
  wire w_mem_inst__abc_21378_n3216;
  wire w_mem_inst__abc_21378_n3217;
  wire w_mem_inst__abc_21378_n3218_1;
  wire w_mem_inst__abc_21378_n3219_1;
  wire w_mem_inst__abc_21378_n3221;
  wire w_mem_inst__abc_21378_n3222_1;
  wire w_mem_inst__abc_21378_n3223_1;
  wire w_mem_inst__abc_21378_n3224;
  wire w_mem_inst__abc_21378_n3225;
  wire w_mem_inst__abc_21378_n3227_1;
  wire w_mem_inst__abc_21378_n3228;
  wire w_mem_inst__abc_21378_n3229;
  wire w_mem_inst__abc_21378_n3230_1;
  wire w_mem_inst__abc_21378_n3231_1;
  wire w_mem_inst__abc_21378_n3233;
  wire w_mem_inst__abc_21378_n3234_1;
  wire w_mem_inst__abc_21378_n3235_1;
  wire w_mem_inst__abc_21378_n3236;
  wire w_mem_inst__abc_21378_n3237;
  wire w_mem_inst__abc_21378_n3239_1;
  wire w_mem_inst__abc_21378_n3240;
  wire w_mem_inst__abc_21378_n3241;
  wire w_mem_inst__abc_21378_n3242_1;
  wire w_mem_inst__abc_21378_n3243_1;
  wire w_mem_inst__abc_21378_n3245;
  wire w_mem_inst__abc_21378_n3246_1;
  wire w_mem_inst__abc_21378_n3247_1;
  wire w_mem_inst__abc_21378_n3248;
  wire w_mem_inst__abc_21378_n3249;
  wire w_mem_inst__abc_21378_n3251_1;
  wire w_mem_inst__abc_21378_n3252;
  wire w_mem_inst__abc_21378_n3253;
  wire w_mem_inst__abc_21378_n3254_1;
  wire w_mem_inst__abc_21378_n3255_1;
  wire w_mem_inst__abc_21378_n3257;
  wire w_mem_inst__abc_21378_n3258_1;
  wire w_mem_inst__abc_21378_n3259_1;
  wire w_mem_inst__abc_21378_n3260;
  wire w_mem_inst__abc_21378_n3261;
  wire w_mem_inst__abc_21378_n3263_1;
  wire w_mem_inst__abc_21378_n3264;
  wire w_mem_inst__abc_21378_n3265;
  wire w_mem_inst__abc_21378_n3266_1;
  wire w_mem_inst__abc_21378_n3267_1;
  wire w_mem_inst__abc_21378_n3269;
  wire w_mem_inst__abc_21378_n3270_1;
  wire w_mem_inst__abc_21378_n3271_1;
  wire w_mem_inst__abc_21378_n3272;
  wire w_mem_inst__abc_21378_n3273;
  wire w_mem_inst__abc_21378_n3275_1;
  wire w_mem_inst__abc_21378_n3276;
  wire w_mem_inst__abc_21378_n3277;
  wire w_mem_inst__abc_21378_n3278_1;
  wire w_mem_inst__abc_21378_n3279_1;
  wire w_mem_inst__abc_21378_n3281;
  wire w_mem_inst__abc_21378_n3282_1;
  wire w_mem_inst__abc_21378_n3283_1;
  wire w_mem_inst__abc_21378_n3284;
  wire w_mem_inst__abc_21378_n3285;
  wire w_mem_inst__abc_21378_n3287_1;
  wire w_mem_inst__abc_21378_n3288;
  wire w_mem_inst__abc_21378_n3289;
  wire w_mem_inst__abc_21378_n3290_1;
  wire w_mem_inst__abc_21378_n3291_1;
  wire w_mem_inst__abc_21378_n3293;
  wire w_mem_inst__abc_21378_n3294_1;
  wire w_mem_inst__abc_21378_n3295_1;
  wire w_mem_inst__abc_21378_n3296;
  wire w_mem_inst__abc_21378_n3297;
  wire w_mem_inst__abc_21378_n3299_1;
  wire w_mem_inst__abc_21378_n3300;
  wire w_mem_inst__abc_21378_n3301;
  wire w_mem_inst__abc_21378_n3302_1;
  wire w_mem_inst__abc_21378_n3303_1;
  wire w_mem_inst__abc_21378_n3305;
  wire w_mem_inst__abc_21378_n3306_1;
  wire w_mem_inst__abc_21378_n3307_1;
  wire w_mem_inst__abc_21378_n3308;
  wire w_mem_inst__abc_21378_n3309;
  wire w_mem_inst__abc_21378_n3311_1;
  wire w_mem_inst__abc_21378_n3312;
  wire w_mem_inst__abc_21378_n3313;
  wire w_mem_inst__abc_21378_n3314_1;
  wire w_mem_inst__abc_21378_n3315_1;
  wire w_mem_inst__abc_21378_n3317;
  wire w_mem_inst__abc_21378_n3318_1;
  wire w_mem_inst__abc_21378_n3319_1;
  wire w_mem_inst__abc_21378_n3320;
  wire w_mem_inst__abc_21378_n3321;
  wire w_mem_inst__abc_21378_n3323_1;
  wire w_mem_inst__abc_21378_n3324;
  wire w_mem_inst__abc_21378_n3325;
  wire w_mem_inst__abc_21378_n3326_1;
  wire w_mem_inst__abc_21378_n3327_1;
  wire w_mem_inst__abc_21378_n3329;
  wire w_mem_inst__abc_21378_n3330_1;
  wire w_mem_inst__abc_21378_n3331_1;
  wire w_mem_inst__abc_21378_n3332;
  wire w_mem_inst__abc_21378_n3333;
  wire w_mem_inst__abc_21378_n3335_1;
  wire w_mem_inst__abc_21378_n3336;
  wire w_mem_inst__abc_21378_n3337;
  wire w_mem_inst__abc_21378_n3338_1;
  wire w_mem_inst__abc_21378_n3339_1;
  wire w_mem_inst__abc_21378_n3341;
  wire w_mem_inst__abc_21378_n3342_1;
  wire w_mem_inst__abc_21378_n3343_1;
  wire w_mem_inst__abc_21378_n3344;
  wire w_mem_inst__abc_21378_n3345;
  wire w_mem_inst__abc_21378_n3347_1;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf0;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf1;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf10;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf11;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf12;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf13;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf14;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf15;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf16;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf17;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf18;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf19;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf2;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf20;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf21;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf22;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf23;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf24;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf25;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf26;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf27;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf28;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf29;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf3;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf30;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf31;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf32;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf33;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf34;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf35;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf36;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf37;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf38;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf39;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf4;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf40;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf41;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf42;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf43;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf44;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf45;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf46;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf47;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf48;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf49;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf5;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf50;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf51;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf52;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf53;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf54;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf55;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf56;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf57;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf58;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf59;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf6;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf60;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf7;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf8;
  wire w_mem_inst__abc_21378_n3347_1_bF_buf9;
  wire w_mem_inst__abc_21378_n3347_1_hier0_bF_buf0;
  wire w_mem_inst__abc_21378_n3347_1_hier0_bF_buf1;
  wire w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2;
  wire w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3;
  wire w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4;
  wire w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5;
  wire w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6;
  wire w_mem_inst__abc_21378_n3348;
  wire w_mem_inst__abc_21378_n3349;
  wire w_mem_inst__abc_21378_n3350_1;
  wire w_mem_inst__abc_21378_n3351_1;
  wire w_mem_inst__abc_21378_n3352;
  wire w_mem_inst__abc_21378_n3354_1;
  wire w_mem_inst__abc_21378_n3355_1;
  wire w_mem_inst__abc_21378_n3356;
  wire w_mem_inst__abc_21378_n3357;
  wire w_mem_inst__abc_21378_n3358_1;
  wire w_mem_inst__abc_21378_n3360;
  wire w_mem_inst__abc_21378_n3361;
  wire w_mem_inst__abc_21378_n3362_1;
  wire w_mem_inst__abc_21378_n3363_1;
  wire w_mem_inst__abc_21378_n3364;
  wire w_mem_inst__abc_21378_n3366_1;
  wire w_mem_inst__abc_21378_n3367_1;
  wire w_mem_inst__abc_21378_n3368;
  wire w_mem_inst__abc_21378_n3369;
  wire w_mem_inst__abc_21378_n3370_1;
  wire w_mem_inst__abc_21378_n3372;
  wire w_mem_inst__abc_21378_n3373;
  wire w_mem_inst__abc_21378_n3374_1;
  wire w_mem_inst__abc_21378_n3375_1;
  wire w_mem_inst__abc_21378_n3376;
  wire w_mem_inst__abc_21378_n3378_1;
  wire w_mem_inst__abc_21378_n3379_1;
  wire w_mem_inst__abc_21378_n3380;
  wire w_mem_inst__abc_21378_n3381;
  wire w_mem_inst__abc_21378_n3382_1;
  wire w_mem_inst__abc_21378_n3384;
  wire w_mem_inst__abc_21378_n3385;
  wire w_mem_inst__abc_21378_n3386_1;
  wire w_mem_inst__abc_21378_n3387_1;
  wire w_mem_inst__abc_21378_n3388;
  wire w_mem_inst__abc_21378_n3390_1;
  wire w_mem_inst__abc_21378_n3391_1;
  wire w_mem_inst__abc_21378_n3392;
  wire w_mem_inst__abc_21378_n3393;
  wire w_mem_inst__abc_21378_n3394_1;
  wire w_mem_inst__abc_21378_n3396;
  wire w_mem_inst__abc_21378_n3397;
  wire w_mem_inst__abc_21378_n3398_1;
  wire w_mem_inst__abc_21378_n3399_1;
  wire w_mem_inst__abc_21378_n3400;
  wire w_mem_inst__abc_21378_n3402_1;
  wire w_mem_inst__abc_21378_n3403_1;
  wire w_mem_inst__abc_21378_n3404;
  wire w_mem_inst__abc_21378_n3405;
  wire w_mem_inst__abc_21378_n3406_1;
  wire w_mem_inst__abc_21378_n3408;
  wire w_mem_inst__abc_21378_n3409;
  wire w_mem_inst__abc_21378_n3410_1;
  wire w_mem_inst__abc_21378_n3411_1;
  wire w_mem_inst__abc_21378_n3412;
  wire w_mem_inst__abc_21378_n3414_1;
  wire w_mem_inst__abc_21378_n3415_1;
  wire w_mem_inst__abc_21378_n3416;
  wire w_mem_inst__abc_21378_n3417;
  wire w_mem_inst__abc_21378_n3418_1;
  wire w_mem_inst__abc_21378_n3420;
  wire w_mem_inst__abc_21378_n3421;
  wire w_mem_inst__abc_21378_n3422_1;
  wire w_mem_inst__abc_21378_n3423_1;
  wire w_mem_inst__abc_21378_n3424;
  wire w_mem_inst__abc_21378_n3426_1;
  wire w_mem_inst__abc_21378_n3427_1;
  wire w_mem_inst__abc_21378_n3428;
  wire w_mem_inst__abc_21378_n3429;
  wire w_mem_inst__abc_21378_n3430_1;
  wire w_mem_inst__abc_21378_n3432;
  wire w_mem_inst__abc_21378_n3433;
  wire w_mem_inst__abc_21378_n3434_1;
  wire w_mem_inst__abc_21378_n3435_1;
  wire w_mem_inst__abc_21378_n3436;
  wire w_mem_inst__abc_21378_n3438_1;
  wire w_mem_inst__abc_21378_n3439_1;
  wire w_mem_inst__abc_21378_n3440;
  wire w_mem_inst__abc_21378_n3441;
  wire w_mem_inst__abc_21378_n3442_1;
  wire w_mem_inst__abc_21378_n3444;
  wire w_mem_inst__abc_21378_n3445;
  wire w_mem_inst__abc_21378_n3446_1;
  wire w_mem_inst__abc_21378_n3447_1;
  wire w_mem_inst__abc_21378_n3448;
  wire w_mem_inst__abc_21378_n3450_1;
  wire w_mem_inst__abc_21378_n3451_1;
  wire w_mem_inst__abc_21378_n3452;
  wire w_mem_inst__abc_21378_n3453;
  wire w_mem_inst__abc_21378_n3454_1;
  wire w_mem_inst__abc_21378_n3456;
  wire w_mem_inst__abc_21378_n3457;
  wire w_mem_inst__abc_21378_n3458_1;
  wire w_mem_inst__abc_21378_n3459_1;
  wire w_mem_inst__abc_21378_n3460;
  wire w_mem_inst__abc_21378_n3462_1;
  wire w_mem_inst__abc_21378_n3463_1;
  wire w_mem_inst__abc_21378_n3464;
  wire w_mem_inst__abc_21378_n3465;
  wire w_mem_inst__abc_21378_n3466_1;
  wire w_mem_inst__abc_21378_n3468;
  wire w_mem_inst__abc_21378_n3469;
  wire w_mem_inst__abc_21378_n3470_1;
  wire w_mem_inst__abc_21378_n3471_1;
  wire w_mem_inst__abc_21378_n3472;
  wire w_mem_inst__abc_21378_n3474_1;
  wire w_mem_inst__abc_21378_n3475_1;
  wire w_mem_inst__abc_21378_n3476;
  wire w_mem_inst__abc_21378_n3477;
  wire w_mem_inst__abc_21378_n3478_1;
  wire w_mem_inst__abc_21378_n3480;
  wire w_mem_inst__abc_21378_n3481;
  wire w_mem_inst__abc_21378_n3482_1;
  wire w_mem_inst__abc_21378_n3483_1;
  wire w_mem_inst__abc_21378_n3484;
  wire w_mem_inst__abc_21378_n3486_1;
  wire w_mem_inst__abc_21378_n3487_1;
  wire w_mem_inst__abc_21378_n3488;
  wire w_mem_inst__abc_21378_n3489;
  wire w_mem_inst__abc_21378_n3490_1;
  wire w_mem_inst__abc_21378_n3492;
  wire w_mem_inst__abc_21378_n3493;
  wire w_mem_inst__abc_21378_n3494_1;
  wire w_mem_inst__abc_21378_n3495_1;
  wire w_mem_inst__abc_21378_n3496;
  wire w_mem_inst__abc_21378_n3498_1;
  wire w_mem_inst__abc_21378_n3499_1;
  wire w_mem_inst__abc_21378_n3500;
  wire w_mem_inst__abc_21378_n3501;
  wire w_mem_inst__abc_21378_n3502_1;
  wire w_mem_inst__abc_21378_n3504;
  wire w_mem_inst__abc_21378_n3505;
  wire w_mem_inst__abc_21378_n3506_1;
  wire w_mem_inst__abc_21378_n3507_1;
  wire w_mem_inst__abc_21378_n3508;
  wire w_mem_inst__abc_21378_n3510_1;
  wire w_mem_inst__abc_21378_n3511_1;
  wire w_mem_inst__abc_21378_n3512;
  wire w_mem_inst__abc_21378_n3513;
  wire w_mem_inst__abc_21378_n3514_1;
  wire w_mem_inst__abc_21378_n3516;
  wire w_mem_inst__abc_21378_n3517;
  wire w_mem_inst__abc_21378_n3518_1;
  wire w_mem_inst__abc_21378_n3519_1;
  wire w_mem_inst__abc_21378_n3520;
  wire w_mem_inst__abc_21378_n3522_1;
  wire w_mem_inst__abc_21378_n3523_1;
  wire w_mem_inst__abc_21378_n3524;
  wire w_mem_inst__abc_21378_n3525;
  wire w_mem_inst__abc_21378_n3526_1;
  wire w_mem_inst__abc_21378_n3528;
  wire w_mem_inst__abc_21378_n3529;
  wire w_mem_inst__abc_21378_n3530_1;
  wire w_mem_inst__abc_21378_n3531_1;
  wire w_mem_inst__abc_21378_n3532;
  wire w_mem_inst__abc_21378_n3534_1;
  wire w_mem_inst__abc_21378_n3535_1;
  wire w_mem_inst__abc_21378_n3536;
  wire w_mem_inst__abc_21378_n3537;
  wire w_mem_inst__abc_21378_n3538_1;
  wire w_mem_inst__abc_21378_n3540;
  wire w_mem_inst__abc_21378_n3541;
  wire w_mem_inst__abc_21378_n3542_1;
  wire w_mem_inst__abc_21378_n3543_1;
  wire w_mem_inst__abc_21378_n3544;
  wire w_mem_inst__abc_21378_n3546_1;
  wire w_mem_inst__abc_21378_n3547_1;
  wire w_mem_inst__abc_21378_n3548;
  wire w_mem_inst__abc_21378_n3549;
  wire w_mem_inst__abc_21378_n3550_1;
  wire w_mem_inst__abc_21378_n3552;
  wire w_mem_inst__abc_21378_n3553;
  wire w_mem_inst__abc_21378_n3554_1;
  wire w_mem_inst__abc_21378_n3555_1;
  wire w_mem_inst__abc_21378_n3556;
  wire w_mem_inst__abc_21378_n3558_1;
  wire w_mem_inst__abc_21378_n3559_1;
  wire w_mem_inst__abc_21378_n3560;
  wire w_mem_inst__abc_21378_n3561;
  wire w_mem_inst__abc_21378_n3562_1;
  wire w_mem_inst__abc_21378_n3564;
  wire w_mem_inst__abc_21378_n3565;
  wire w_mem_inst__abc_21378_n3566_1;
  wire w_mem_inst__abc_21378_n3567_1;
  wire w_mem_inst__abc_21378_n3568;
  wire w_mem_inst__abc_21378_n3570_1;
  wire w_mem_inst__abc_21378_n3571_1;
  wire w_mem_inst__abc_21378_n3572;
  wire w_mem_inst__abc_21378_n3573;
  wire w_mem_inst__abc_21378_n3574_1;
  wire w_mem_inst__abc_21378_n3576;
  wire w_mem_inst__abc_21378_n3577;
  wire w_mem_inst__abc_21378_n3578_1;
  wire w_mem_inst__abc_21378_n3579_1;
  wire w_mem_inst__abc_21378_n3580;
  wire w_mem_inst__abc_21378_n3582_1;
  wire w_mem_inst__abc_21378_n3583_1;
  wire w_mem_inst__abc_21378_n3584;
  wire w_mem_inst__abc_21378_n3585;
  wire w_mem_inst__abc_21378_n3586_1;
  wire w_mem_inst__abc_21378_n3588;
  wire w_mem_inst__abc_21378_n3589;
  wire w_mem_inst__abc_21378_n3590_1;
  wire w_mem_inst__abc_21378_n3591_1;
  wire w_mem_inst__abc_21378_n3592;
  wire w_mem_inst__abc_21378_n3594_1;
  wire w_mem_inst__abc_21378_n3595_1;
  wire w_mem_inst__abc_21378_n3596;
  wire w_mem_inst__abc_21378_n3597;
  wire w_mem_inst__abc_21378_n3598_1;
  wire w_mem_inst__abc_21378_n3600;
  wire w_mem_inst__abc_21378_n3601;
  wire w_mem_inst__abc_21378_n3602_1;
  wire w_mem_inst__abc_21378_n3603_1;
  wire w_mem_inst__abc_21378_n3604;
  wire w_mem_inst__abc_21378_n3606_1;
  wire w_mem_inst__abc_21378_n3607_1;
  wire w_mem_inst__abc_21378_n3608;
  wire w_mem_inst__abc_21378_n3609;
  wire w_mem_inst__abc_21378_n3610_1;
  wire w_mem_inst__abc_21378_n3612;
  wire w_mem_inst__abc_21378_n3613;
  wire w_mem_inst__abc_21378_n3614_1;
  wire w_mem_inst__abc_21378_n3615_1;
  wire w_mem_inst__abc_21378_n3616;
  wire w_mem_inst__abc_21378_n3618_1;
  wire w_mem_inst__abc_21378_n3619_1;
  wire w_mem_inst__abc_21378_n3620;
  wire w_mem_inst__abc_21378_n3621;
  wire w_mem_inst__abc_21378_n3622_1;
  wire w_mem_inst__abc_21378_n3624;
  wire w_mem_inst__abc_21378_n3625;
  wire w_mem_inst__abc_21378_n3626_1;
  wire w_mem_inst__abc_21378_n3627_1;
  wire w_mem_inst__abc_21378_n3628;
  wire w_mem_inst__abc_21378_n3630_1;
  wire w_mem_inst__abc_21378_n3631_1;
  wire w_mem_inst__abc_21378_n3632;
  wire w_mem_inst__abc_21378_n3633;
  wire w_mem_inst__abc_21378_n3634_1;
  wire w_mem_inst__abc_21378_n3636;
  wire w_mem_inst__abc_21378_n3637;
  wire w_mem_inst__abc_21378_n3638_1;
  wire w_mem_inst__abc_21378_n3639_1;
  wire w_mem_inst__abc_21378_n3640;
  wire w_mem_inst__abc_21378_n3642_1;
  wire w_mem_inst__abc_21378_n3643_1;
  wire w_mem_inst__abc_21378_n3644;
  wire w_mem_inst__abc_21378_n3645;
  wire w_mem_inst__abc_21378_n3646_1;
  wire w_mem_inst__abc_21378_n3648;
  wire w_mem_inst__abc_21378_n3649;
  wire w_mem_inst__abc_21378_n3650_1;
  wire w_mem_inst__abc_21378_n3651;
  wire w_mem_inst__abc_21378_n3652;
  wire w_mem_inst__abc_21378_n3654;
  wire w_mem_inst__abc_21378_n3655;
  wire w_mem_inst__abc_21378_n3656;
  wire w_mem_inst__abc_21378_n3657_1;
  wire w_mem_inst__abc_21378_n3658;
  wire w_mem_inst__abc_21378_n3660;
  wire w_mem_inst__abc_21378_n3661;
  wire w_mem_inst__abc_21378_n3662_1;
  wire w_mem_inst__abc_21378_n3663;
  wire w_mem_inst__abc_21378_n3664;
  wire w_mem_inst__abc_21378_n3666;
  wire w_mem_inst__abc_21378_n3667;
  wire w_mem_inst__abc_21378_n3668;
  wire w_mem_inst__abc_21378_n3669_1;
  wire w_mem_inst__abc_21378_n3670;
  wire w_mem_inst__abc_21378_n3672;
  wire w_mem_inst__abc_21378_n3673_1;
  wire w_mem_inst__abc_21378_n3674;
  wire w_mem_inst__abc_21378_n3675;
  wire w_mem_inst__abc_21378_n3676;
  wire w_mem_inst__abc_21378_n3678;
  wire w_mem_inst__abc_21378_n3679;
  wire w_mem_inst__abc_21378_n3680;
  wire w_mem_inst__abc_21378_n3681;
  wire w_mem_inst__abc_21378_n3682;
  wire w_mem_inst__abc_21378_n3684;
  wire w_mem_inst__abc_21378_n3685;
  wire w_mem_inst__abc_21378_n3686;
  wire w_mem_inst__abc_21378_n3687;
  wire w_mem_inst__abc_21378_n3688;
  wire w_mem_inst__abc_21378_n3690;
  wire w_mem_inst__abc_21378_n3691;
  wire w_mem_inst__abc_21378_n3692;
  wire w_mem_inst__abc_21378_n3693;
  wire w_mem_inst__abc_21378_n3694;
  wire w_mem_inst__abc_21378_n3696;
  wire w_mem_inst__abc_21378_n3697;
  wire w_mem_inst__abc_21378_n3698;
  wire w_mem_inst__abc_21378_n3699;
  wire w_mem_inst__abc_21378_n3700;
  wire w_mem_inst__abc_21378_n3702;
  wire w_mem_inst__abc_21378_n3703;
  wire w_mem_inst__abc_21378_n3704;
  wire w_mem_inst__abc_21378_n3705;
  wire w_mem_inst__abc_21378_n3706;
  wire w_mem_inst__abc_21378_n3708;
  wire w_mem_inst__abc_21378_n3709;
  wire w_mem_inst__abc_21378_n3710;
  wire w_mem_inst__abc_21378_n3711;
  wire w_mem_inst__abc_21378_n3712;
  wire w_mem_inst__abc_21378_n3714;
  wire w_mem_inst__abc_21378_n3715;
  wire w_mem_inst__abc_21378_n3716;
  wire w_mem_inst__abc_21378_n3717;
  wire w_mem_inst__abc_21378_n3718;
  wire w_mem_inst__abc_21378_n3720;
  wire w_mem_inst__abc_21378_n3721;
  wire w_mem_inst__abc_21378_n3722;
  wire w_mem_inst__abc_21378_n3723;
  wire w_mem_inst__abc_21378_n3724;
  wire w_mem_inst__abc_21378_n3726;
  wire w_mem_inst__abc_21378_n3727;
  wire w_mem_inst__abc_21378_n3728;
  wire w_mem_inst__abc_21378_n3729;
  wire w_mem_inst__abc_21378_n3730;
  wire w_mem_inst__abc_21378_n3732;
  wire w_mem_inst__abc_21378_n3733;
  wire w_mem_inst__abc_21378_n3734;
  wire w_mem_inst__abc_21378_n3735;
  wire w_mem_inst__abc_21378_n3736;
  wire w_mem_inst__abc_21378_n3738;
  wire w_mem_inst__abc_21378_n3739;
  wire w_mem_inst__abc_21378_n3740;
  wire w_mem_inst__abc_21378_n3741;
  wire w_mem_inst__abc_21378_n3742;
  wire w_mem_inst__abc_21378_n3744;
  wire w_mem_inst__abc_21378_n3745;
  wire w_mem_inst__abc_21378_n3746;
  wire w_mem_inst__abc_21378_n3747;
  wire w_mem_inst__abc_21378_n3748;
  wire w_mem_inst__abc_21378_n3750;
  wire w_mem_inst__abc_21378_n3751;
  wire w_mem_inst__abc_21378_n3752;
  wire w_mem_inst__abc_21378_n3753;
  wire w_mem_inst__abc_21378_n3754;
  wire w_mem_inst__abc_21378_n3756;
  wire w_mem_inst__abc_21378_n3757;
  wire w_mem_inst__abc_21378_n3758;
  wire w_mem_inst__abc_21378_n3759;
  wire w_mem_inst__abc_21378_n3760;
  wire w_mem_inst__abc_21378_n3762;
  wire w_mem_inst__abc_21378_n3763;
  wire w_mem_inst__abc_21378_n3764;
  wire w_mem_inst__abc_21378_n3765;
  wire w_mem_inst__abc_21378_n3766;
  wire w_mem_inst__abc_21378_n3768;
  wire w_mem_inst__abc_21378_n3769;
  wire w_mem_inst__abc_21378_n3770;
  wire w_mem_inst__abc_21378_n3771;
  wire w_mem_inst__abc_21378_n3772;
  wire w_mem_inst__abc_21378_n3774;
  wire w_mem_inst__abc_21378_n3775;
  wire w_mem_inst__abc_21378_n3776;
  wire w_mem_inst__abc_21378_n3777;
  wire w_mem_inst__abc_21378_n3778;
  wire w_mem_inst__abc_21378_n3780;
  wire w_mem_inst__abc_21378_n3781;
  wire w_mem_inst__abc_21378_n3782;
  wire w_mem_inst__abc_21378_n3783;
  wire w_mem_inst__abc_21378_n3784;
  wire w_mem_inst__abc_21378_n3786;
  wire w_mem_inst__abc_21378_n3787;
  wire w_mem_inst__abc_21378_n3788;
  wire w_mem_inst__abc_21378_n3789;
  wire w_mem_inst__abc_21378_n3790;
  wire w_mem_inst__abc_21378_n3792;
  wire w_mem_inst__abc_21378_n3793;
  wire w_mem_inst__abc_21378_n3794;
  wire w_mem_inst__abc_21378_n3795;
  wire w_mem_inst__abc_21378_n3796;
  wire w_mem_inst__abc_21378_n3798;
  wire w_mem_inst__abc_21378_n3799;
  wire w_mem_inst__abc_21378_n3800;
  wire w_mem_inst__abc_21378_n3801;
  wire w_mem_inst__abc_21378_n3802;
  wire w_mem_inst__abc_21378_n3804;
  wire w_mem_inst__abc_21378_n3805;
  wire w_mem_inst__abc_21378_n3806;
  wire w_mem_inst__abc_21378_n3807;
  wire w_mem_inst__abc_21378_n3808;
  wire w_mem_inst__abc_21378_n3810;
  wire w_mem_inst__abc_21378_n3811;
  wire w_mem_inst__abc_21378_n3812;
  wire w_mem_inst__abc_21378_n3813;
  wire w_mem_inst__abc_21378_n3814;
  wire w_mem_inst__abc_21378_n3816;
  wire w_mem_inst__abc_21378_n3817;
  wire w_mem_inst__abc_21378_n3818;
  wire w_mem_inst__abc_21378_n3819;
  wire w_mem_inst__abc_21378_n3820;
  wire w_mem_inst__abc_21378_n3822;
  wire w_mem_inst__abc_21378_n3823;
  wire w_mem_inst__abc_21378_n3824;
  wire w_mem_inst__abc_21378_n3825;
  wire w_mem_inst__abc_21378_n3826;
  wire w_mem_inst__abc_21378_n3828;
  wire w_mem_inst__abc_21378_n3829;
  wire w_mem_inst__abc_21378_n3830;
  wire w_mem_inst__abc_21378_n3831;
  wire w_mem_inst__abc_21378_n3832;
  wire w_mem_inst__abc_21378_n3834;
  wire w_mem_inst__abc_21378_n3835;
  wire w_mem_inst__abc_21378_n3836;
  wire w_mem_inst__abc_21378_n3837;
  wire w_mem_inst__abc_21378_n3838;
  wire w_mem_inst__abc_21378_n3840;
  wire w_mem_inst__abc_21378_n3841;
  wire w_mem_inst__abc_21378_n3842;
  wire w_mem_inst__abc_21378_n3843;
  wire w_mem_inst__abc_21378_n3844;
  wire w_mem_inst__abc_21378_n3846;
  wire w_mem_inst__abc_21378_n3847;
  wire w_mem_inst__abc_21378_n3848;
  wire w_mem_inst__abc_21378_n3849;
  wire w_mem_inst__abc_21378_n3850;
  wire w_mem_inst__abc_21378_n3852;
  wire w_mem_inst__abc_21378_n3853;
  wire w_mem_inst__abc_21378_n3854;
  wire w_mem_inst__abc_21378_n3855;
  wire w_mem_inst__abc_21378_n3856;
  wire w_mem_inst__abc_21378_n3858;
  wire w_mem_inst__abc_21378_n3859;
  wire w_mem_inst__abc_21378_n3860;
  wire w_mem_inst__abc_21378_n3861;
  wire w_mem_inst__abc_21378_n3862;
  wire w_mem_inst__abc_21378_n3864;
  wire w_mem_inst__abc_21378_n3865;
  wire w_mem_inst__abc_21378_n3866;
  wire w_mem_inst__abc_21378_n3867;
  wire w_mem_inst__abc_21378_n3868;
  wire w_mem_inst__abc_21378_n3870;
  wire w_mem_inst__abc_21378_n3871;
  wire w_mem_inst__abc_21378_n3872;
  wire w_mem_inst__abc_21378_n3873;
  wire w_mem_inst__abc_21378_n3874;
  wire w_mem_inst__abc_21378_n3876;
  wire w_mem_inst__abc_21378_n3877;
  wire w_mem_inst__abc_21378_n3878;
  wire w_mem_inst__abc_21378_n3879;
  wire w_mem_inst__abc_21378_n3880;
  wire w_mem_inst__abc_21378_n3882;
  wire w_mem_inst__abc_21378_n3883;
  wire w_mem_inst__abc_21378_n3884;
  wire w_mem_inst__abc_21378_n3885;
  wire w_mem_inst__abc_21378_n3886;
  wire w_mem_inst__abc_21378_n3888;
  wire w_mem_inst__abc_21378_n3889;
  wire w_mem_inst__abc_21378_n3890;
  wire w_mem_inst__abc_21378_n3891;
  wire w_mem_inst__abc_21378_n3892;
  wire w_mem_inst__abc_21378_n3894;
  wire w_mem_inst__abc_21378_n3895;
  wire w_mem_inst__abc_21378_n3896;
  wire w_mem_inst__abc_21378_n3897;
  wire w_mem_inst__abc_21378_n3898;
  wire w_mem_inst__abc_21378_n3900;
  wire w_mem_inst__abc_21378_n3901;
  wire w_mem_inst__abc_21378_n3902;
  wire w_mem_inst__abc_21378_n3903;
  wire w_mem_inst__abc_21378_n3904;
  wire w_mem_inst__abc_21378_n3906;
  wire w_mem_inst__abc_21378_n3907;
  wire w_mem_inst__abc_21378_n3908;
  wire w_mem_inst__abc_21378_n3909;
  wire w_mem_inst__abc_21378_n3910;
  wire w_mem_inst__abc_21378_n3912;
  wire w_mem_inst__abc_21378_n3913;
  wire w_mem_inst__abc_21378_n3914;
  wire w_mem_inst__abc_21378_n3915;
  wire w_mem_inst__abc_21378_n3916;
  wire w_mem_inst__abc_21378_n3918;
  wire w_mem_inst__abc_21378_n3919;
  wire w_mem_inst__abc_21378_n3920;
  wire w_mem_inst__abc_21378_n3921;
  wire w_mem_inst__abc_21378_n3922;
  wire w_mem_inst__abc_21378_n3924;
  wire w_mem_inst__abc_21378_n3925;
  wire w_mem_inst__abc_21378_n3926;
  wire w_mem_inst__abc_21378_n3927;
  wire w_mem_inst__abc_21378_n3928;
  wire w_mem_inst__abc_21378_n3930;
  wire w_mem_inst__abc_21378_n3931;
  wire w_mem_inst__abc_21378_n3932;
  wire w_mem_inst__abc_21378_n3933;
  wire w_mem_inst__abc_21378_n3934;
  wire w_mem_inst__abc_21378_n3936;
  wire w_mem_inst__abc_21378_n3937;
  wire w_mem_inst__abc_21378_n3938;
  wire w_mem_inst__abc_21378_n3939;
  wire w_mem_inst__abc_21378_n3940;
  wire w_mem_inst__abc_21378_n3942;
  wire w_mem_inst__abc_21378_n3943;
  wire w_mem_inst__abc_21378_n3944;
  wire w_mem_inst__abc_21378_n3945;
  wire w_mem_inst__abc_21378_n3946;
  wire w_mem_inst__abc_21378_n3948;
  wire w_mem_inst__abc_21378_n3949;
  wire w_mem_inst__abc_21378_n3950;
  wire w_mem_inst__abc_21378_n3951;
  wire w_mem_inst__abc_21378_n3952;
  wire w_mem_inst__abc_21378_n3954;
  wire w_mem_inst__abc_21378_n3955;
  wire w_mem_inst__abc_21378_n3956;
  wire w_mem_inst__abc_21378_n3957;
  wire w_mem_inst__abc_21378_n3958;
  wire w_mem_inst__abc_21378_n3960;
  wire w_mem_inst__abc_21378_n3961;
  wire w_mem_inst__abc_21378_n3962;
  wire w_mem_inst__abc_21378_n3963;
  wire w_mem_inst__abc_21378_n3964;
  wire w_mem_inst__abc_21378_n3966;
  wire w_mem_inst__abc_21378_n3967;
  wire w_mem_inst__abc_21378_n3968;
  wire w_mem_inst__abc_21378_n3969;
  wire w_mem_inst__abc_21378_n3970;
  wire w_mem_inst__abc_21378_n3972;
  wire w_mem_inst__abc_21378_n3973;
  wire w_mem_inst__abc_21378_n3974;
  wire w_mem_inst__abc_21378_n3975;
  wire w_mem_inst__abc_21378_n3976;
  wire w_mem_inst__abc_21378_n3978;
  wire w_mem_inst__abc_21378_n3979;
  wire w_mem_inst__abc_21378_n3980;
  wire w_mem_inst__abc_21378_n3981;
  wire w_mem_inst__abc_21378_n3982;
  wire w_mem_inst__abc_21378_n3984;
  wire w_mem_inst__abc_21378_n3985;
  wire w_mem_inst__abc_21378_n3986;
  wire w_mem_inst__abc_21378_n3987;
  wire w_mem_inst__abc_21378_n3988;
  wire w_mem_inst__abc_21378_n3990;
  wire w_mem_inst__abc_21378_n3991;
  wire w_mem_inst__abc_21378_n3992;
  wire w_mem_inst__abc_21378_n3993;
  wire w_mem_inst__abc_21378_n3994;
  wire w_mem_inst__abc_21378_n3996;
  wire w_mem_inst__abc_21378_n3997;
  wire w_mem_inst__abc_21378_n3998;
  wire w_mem_inst__abc_21378_n3999;
  wire w_mem_inst__abc_21378_n4000;
  wire w_mem_inst__abc_21378_n4002;
  wire w_mem_inst__abc_21378_n4003;
  wire w_mem_inst__abc_21378_n4004;
  wire w_mem_inst__abc_21378_n4005;
  wire w_mem_inst__abc_21378_n4006;
  wire w_mem_inst__abc_21378_n4008;
  wire w_mem_inst__abc_21378_n4009;
  wire w_mem_inst__abc_21378_n4010;
  wire w_mem_inst__abc_21378_n4011;
  wire w_mem_inst__abc_21378_n4012;
  wire w_mem_inst__abc_21378_n4014;
  wire w_mem_inst__abc_21378_n4015;
  wire w_mem_inst__abc_21378_n4016;
  wire w_mem_inst__abc_21378_n4017;
  wire w_mem_inst__abc_21378_n4018;
  wire w_mem_inst__abc_21378_n4020;
  wire w_mem_inst__abc_21378_n4021;
  wire w_mem_inst__abc_21378_n4022;
  wire w_mem_inst__abc_21378_n4023;
  wire w_mem_inst__abc_21378_n4024;
  wire w_mem_inst__abc_21378_n4026;
  wire w_mem_inst__abc_21378_n4027;
  wire w_mem_inst__abc_21378_n4028;
  wire w_mem_inst__abc_21378_n4029;
  wire w_mem_inst__abc_21378_n4030;
  wire w_mem_inst__abc_21378_n4032;
  wire w_mem_inst__abc_21378_n4033;
  wire w_mem_inst__abc_21378_n4034;
  wire w_mem_inst__abc_21378_n4035;
  wire w_mem_inst__abc_21378_n4036;
  wire w_mem_inst__abc_21378_n4038;
  wire w_mem_inst__abc_21378_n4039;
  wire w_mem_inst__abc_21378_n4040;
  wire w_mem_inst__abc_21378_n4041;
  wire w_mem_inst__abc_21378_n4042;
  wire w_mem_inst__abc_21378_n4044;
  wire w_mem_inst__abc_21378_n4045;
  wire w_mem_inst__abc_21378_n4046;
  wire w_mem_inst__abc_21378_n4047;
  wire w_mem_inst__abc_21378_n4048;
  wire w_mem_inst__abc_21378_n4050;
  wire w_mem_inst__abc_21378_n4051;
  wire w_mem_inst__abc_21378_n4052;
  wire w_mem_inst__abc_21378_n4053;
  wire w_mem_inst__abc_21378_n4054;
  wire w_mem_inst__abc_21378_n4056;
  wire w_mem_inst__abc_21378_n4057;
  wire w_mem_inst__abc_21378_n4058;
  wire w_mem_inst__abc_21378_n4059;
  wire w_mem_inst__abc_21378_n4060;
  wire w_mem_inst__abc_21378_n4062;
  wire w_mem_inst__abc_21378_n4063;
  wire w_mem_inst__abc_21378_n4064;
  wire w_mem_inst__abc_21378_n4065;
  wire w_mem_inst__abc_21378_n4066;
  wire w_mem_inst__abc_21378_n4068;
  wire w_mem_inst__abc_21378_n4069;
  wire w_mem_inst__abc_21378_n4070;
  wire w_mem_inst__abc_21378_n4071;
  wire w_mem_inst__abc_21378_n4072;
  wire w_mem_inst__abc_21378_n4074;
  wire w_mem_inst__abc_21378_n4075;
  wire w_mem_inst__abc_21378_n4076;
  wire w_mem_inst__abc_21378_n4077;
  wire w_mem_inst__abc_21378_n4078;
  wire w_mem_inst__abc_21378_n4080;
  wire w_mem_inst__abc_21378_n4081;
  wire w_mem_inst__abc_21378_n4082;
  wire w_mem_inst__abc_21378_n4083;
  wire w_mem_inst__abc_21378_n4084;
  wire w_mem_inst__abc_21378_n4086;
  wire w_mem_inst__abc_21378_n4087;
  wire w_mem_inst__abc_21378_n4088;
  wire w_mem_inst__abc_21378_n4089;
  wire w_mem_inst__abc_21378_n4090;
  wire w_mem_inst__abc_21378_n4092;
  wire w_mem_inst__abc_21378_n4093;
  wire w_mem_inst__abc_21378_n4094;
  wire w_mem_inst__abc_21378_n4095;
  wire w_mem_inst__abc_21378_n4096;
  wire w_mem_inst__abc_21378_n4098;
  wire w_mem_inst__abc_21378_n4099;
  wire w_mem_inst__abc_21378_n4100;
  wire w_mem_inst__abc_21378_n4101;
  wire w_mem_inst__abc_21378_n4102;
  wire w_mem_inst__abc_21378_n4104;
  wire w_mem_inst__abc_21378_n4105;
  wire w_mem_inst__abc_21378_n4106;
  wire w_mem_inst__abc_21378_n4107;
  wire w_mem_inst__abc_21378_n4108;
  wire w_mem_inst__abc_21378_n4110;
  wire w_mem_inst__abc_21378_n4111;
  wire w_mem_inst__abc_21378_n4112;
  wire w_mem_inst__abc_21378_n4113;
  wire w_mem_inst__abc_21378_n4114;
  wire w_mem_inst__abc_21378_n4116;
  wire w_mem_inst__abc_21378_n4117;
  wire w_mem_inst__abc_21378_n4118;
  wire w_mem_inst__abc_21378_n4119;
  wire w_mem_inst__abc_21378_n4120;
  wire w_mem_inst__abc_21378_n4122;
  wire w_mem_inst__abc_21378_n4123;
  wire w_mem_inst__abc_21378_n4124;
  wire w_mem_inst__abc_21378_n4125;
  wire w_mem_inst__abc_21378_n4126;
  wire w_mem_inst__abc_21378_n4128;
  wire w_mem_inst__abc_21378_n4129;
  wire w_mem_inst__abc_21378_n4130;
  wire w_mem_inst__abc_21378_n4131;
  wire w_mem_inst__abc_21378_n4132;
  wire w_mem_inst__abc_21378_n4134;
  wire w_mem_inst__abc_21378_n4135;
  wire w_mem_inst__abc_21378_n4136;
  wire w_mem_inst__abc_21378_n4137;
  wire w_mem_inst__abc_21378_n4138;
  wire w_mem_inst__abc_21378_n4140;
  wire w_mem_inst__abc_21378_n4141;
  wire w_mem_inst__abc_21378_n4142;
  wire w_mem_inst__abc_21378_n4143;
  wire w_mem_inst__abc_21378_n4144;
  wire w_mem_inst__abc_21378_n4146;
  wire w_mem_inst__abc_21378_n4147;
  wire w_mem_inst__abc_21378_n4148;
  wire w_mem_inst__abc_21378_n4149;
  wire w_mem_inst__abc_21378_n4150;
  wire w_mem_inst__abc_21378_n4152;
  wire w_mem_inst__abc_21378_n4153;
  wire w_mem_inst__abc_21378_n4154;
  wire w_mem_inst__abc_21378_n4155;
  wire w_mem_inst__abc_21378_n4156;
  wire w_mem_inst__abc_21378_n4158;
  wire w_mem_inst__abc_21378_n4159;
  wire w_mem_inst__abc_21378_n4160;
  wire w_mem_inst__abc_21378_n4161;
  wire w_mem_inst__abc_21378_n4162;
  wire w_mem_inst__abc_21378_n4164;
  wire w_mem_inst__abc_21378_n4165;
  wire w_mem_inst__abc_21378_n4166;
  wire w_mem_inst__abc_21378_n4167;
  wire w_mem_inst__abc_21378_n4168;
  wire w_mem_inst__abc_21378_n4170;
  wire w_mem_inst__abc_21378_n4171;
  wire w_mem_inst__abc_21378_n4172;
  wire w_mem_inst__abc_21378_n4173;
  wire w_mem_inst__abc_21378_n4174;
  wire w_mem_inst__abc_21378_n4176;
  wire w_mem_inst__abc_21378_n4177;
  wire w_mem_inst__abc_21378_n4178;
  wire w_mem_inst__abc_21378_n4179;
  wire w_mem_inst__abc_21378_n4180;
  wire w_mem_inst__abc_21378_n4182;
  wire w_mem_inst__abc_21378_n4183;
  wire w_mem_inst__abc_21378_n4184;
  wire w_mem_inst__abc_21378_n4185;
  wire w_mem_inst__abc_21378_n4186;
  wire w_mem_inst__abc_21378_n4188;
  wire w_mem_inst__abc_21378_n4189;
  wire w_mem_inst__abc_21378_n4190;
  wire w_mem_inst__abc_21378_n4191;
  wire w_mem_inst__abc_21378_n4192;
  wire w_mem_inst__abc_21378_n4194;
  wire w_mem_inst__abc_21378_n4195;
  wire w_mem_inst__abc_21378_n4196;
  wire w_mem_inst__abc_21378_n4197;
  wire w_mem_inst__abc_21378_n4198;
  wire w_mem_inst__abc_21378_n4200;
  wire w_mem_inst__abc_21378_n4201;
  wire w_mem_inst__abc_21378_n4202;
  wire w_mem_inst__abc_21378_n4203;
  wire w_mem_inst__abc_21378_n4204;
  wire w_mem_inst__abc_21378_n4206;
  wire w_mem_inst__abc_21378_n4207;
  wire w_mem_inst__abc_21378_n4208;
  wire w_mem_inst__abc_21378_n4209;
  wire w_mem_inst__abc_21378_n4210;
  wire w_mem_inst__abc_21378_n4212;
  wire w_mem_inst__abc_21378_n4213;
  wire w_mem_inst__abc_21378_n4214;
  wire w_mem_inst__abc_21378_n4215;
  wire w_mem_inst__abc_21378_n4216;
  wire w_mem_inst__abc_21378_n4218;
  wire w_mem_inst__abc_21378_n4219;
  wire w_mem_inst__abc_21378_n4220;
  wire w_mem_inst__abc_21378_n4221;
  wire w_mem_inst__abc_21378_n4222;
  wire w_mem_inst__abc_21378_n4224;
  wire w_mem_inst__abc_21378_n4225;
  wire w_mem_inst__abc_21378_n4226;
  wire w_mem_inst__abc_21378_n4227;
  wire w_mem_inst__abc_21378_n4228;
  wire w_mem_inst__abc_21378_n4230;
  wire w_mem_inst__abc_21378_n4231;
  wire w_mem_inst__abc_21378_n4232;
  wire w_mem_inst__abc_21378_n4233;
  wire w_mem_inst__abc_21378_n4234;
  wire w_mem_inst__abc_21378_n4236;
  wire w_mem_inst__abc_21378_n4237;
  wire w_mem_inst__abc_21378_n4238;
  wire w_mem_inst__abc_21378_n4239;
  wire w_mem_inst__abc_21378_n4240;
  wire w_mem_inst__abc_21378_n4242;
  wire w_mem_inst__abc_21378_n4243;
  wire w_mem_inst__abc_21378_n4244;
  wire w_mem_inst__abc_21378_n4245;
  wire w_mem_inst__abc_21378_n4246;
  wire w_mem_inst__abc_21378_n4248;
  wire w_mem_inst__abc_21378_n4249;
  wire w_mem_inst__abc_21378_n4250;
  wire w_mem_inst__abc_21378_n4251;
  wire w_mem_inst__abc_21378_n4252;
  wire w_mem_inst__abc_21378_n4254;
  wire w_mem_inst__abc_21378_n4255;
  wire w_mem_inst__abc_21378_n4256;
  wire w_mem_inst__abc_21378_n4257;
  wire w_mem_inst__abc_21378_n4258;
  wire w_mem_inst__abc_21378_n4260;
  wire w_mem_inst__abc_21378_n4261;
  wire w_mem_inst__abc_21378_n4262;
  wire w_mem_inst__abc_21378_n4263;
  wire w_mem_inst__abc_21378_n4264;
  wire w_mem_inst__abc_21378_n4266;
  wire w_mem_inst__abc_21378_n4267;
  wire w_mem_inst__abc_21378_n4268;
  wire w_mem_inst__abc_21378_n4269;
  wire w_mem_inst__abc_21378_n4270;
  wire w_mem_inst__abc_21378_n4272;
  wire w_mem_inst__abc_21378_n4273;
  wire w_mem_inst__abc_21378_n4274;
  wire w_mem_inst__abc_21378_n4275;
  wire w_mem_inst__abc_21378_n4276;
  wire w_mem_inst__abc_21378_n4278;
  wire w_mem_inst__abc_21378_n4279;
  wire w_mem_inst__abc_21378_n4280;
  wire w_mem_inst__abc_21378_n4281;
  wire w_mem_inst__abc_21378_n4282;
  wire w_mem_inst__abc_21378_n4284;
  wire w_mem_inst__abc_21378_n4285;
  wire w_mem_inst__abc_21378_n4286;
  wire w_mem_inst__abc_21378_n4287;
  wire w_mem_inst__abc_21378_n4288;
  wire w_mem_inst__abc_21378_n4290;
  wire w_mem_inst__abc_21378_n4291;
  wire w_mem_inst__abc_21378_n4292;
  wire w_mem_inst__abc_21378_n4293;
  wire w_mem_inst__abc_21378_n4294;
  wire w_mem_inst__abc_21378_n4296;
  wire w_mem_inst__abc_21378_n4297;
  wire w_mem_inst__abc_21378_n4298;
  wire w_mem_inst__abc_21378_n4299;
  wire w_mem_inst__abc_21378_n4300;
  wire w_mem_inst__abc_21378_n4302;
  wire w_mem_inst__abc_21378_n4303;
  wire w_mem_inst__abc_21378_n4304;
  wire w_mem_inst__abc_21378_n4305;
  wire w_mem_inst__abc_21378_n4306;
  wire w_mem_inst__abc_21378_n4308;
  wire w_mem_inst__abc_21378_n4309;
  wire w_mem_inst__abc_21378_n4310;
  wire w_mem_inst__abc_21378_n4311;
  wire w_mem_inst__abc_21378_n4312;
  wire w_mem_inst__abc_21378_n4314;
  wire w_mem_inst__abc_21378_n4315;
  wire w_mem_inst__abc_21378_n4316;
  wire w_mem_inst__abc_21378_n4317;
  wire w_mem_inst__abc_21378_n4318;
  wire w_mem_inst__abc_21378_n4320;
  wire w_mem_inst__abc_21378_n4321;
  wire w_mem_inst__abc_21378_n4322;
  wire w_mem_inst__abc_21378_n4323;
  wire w_mem_inst__abc_21378_n4324;
  wire w_mem_inst__abc_21378_n4326;
  wire w_mem_inst__abc_21378_n4327;
  wire w_mem_inst__abc_21378_n4328;
  wire w_mem_inst__abc_21378_n4329;
  wire w_mem_inst__abc_21378_n4330;
  wire w_mem_inst__abc_21378_n4332;
  wire w_mem_inst__abc_21378_n4333;
  wire w_mem_inst__abc_21378_n4334;
  wire w_mem_inst__abc_21378_n4335;
  wire w_mem_inst__abc_21378_n4336;
  wire w_mem_inst__abc_21378_n4338;
  wire w_mem_inst__abc_21378_n4339;
  wire w_mem_inst__abc_21378_n4340;
  wire w_mem_inst__abc_21378_n4341;
  wire w_mem_inst__abc_21378_n4342;
  wire w_mem_inst__abc_21378_n4344;
  wire w_mem_inst__abc_21378_n4345;
  wire w_mem_inst__abc_21378_n4346;
  wire w_mem_inst__abc_21378_n4347;
  wire w_mem_inst__abc_21378_n4348;
  wire w_mem_inst__abc_21378_n4350;
  wire w_mem_inst__abc_21378_n4351;
  wire w_mem_inst__abc_21378_n4352;
  wire w_mem_inst__abc_21378_n4353;
  wire w_mem_inst__abc_21378_n4354;
  wire w_mem_inst__abc_21378_n4356;
  wire w_mem_inst__abc_21378_n4357;
  wire w_mem_inst__abc_21378_n4358;
  wire w_mem_inst__abc_21378_n4359;
  wire w_mem_inst__abc_21378_n4360;
  wire w_mem_inst__abc_21378_n4362;
  wire w_mem_inst__abc_21378_n4363;
  wire w_mem_inst__abc_21378_n4364;
  wire w_mem_inst__abc_21378_n4365;
  wire w_mem_inst__abc_21378_n4366;
  wire w_mem_inst__abc_21378_n4368;
  wire w_mem_inst__abc_21378_n4369;
  wire w_mem_inst__abc_21378_n4370;
  wire w_mem_inst__abc_21378_n4371;
  wire w_mem_inst__abc_21378_n4372;
  wire w_mem_inst__abc_21378_n4374;
  wire w_mem_inst__abc_21378_n4375;
  wire w_mem_inst__abc_21378_n4376;
  wire w_mem_inst__abc_21378_n4377;
  wire w_mem_inst__abc_21378_n4378;
  wire w_mem_inst__abc_21378_n4380;
  wire w_mem_inst__abc_21378_n4381;
  wire w_mem_inst__abc_21378_n4382;
  wire w_mem_inst__abc_21378_n4383;
  wire w_mem_inst__abc_21378_n4384;
  wire w_mem_inst__abc_21378_n4386;
  wire w_mem_inst__abc_21378_n4387;
  wire w_mem_inst__abc_21378_n4388;
  wire w_mem_inst__abc_21378_n4389;
  wire w_mem_inst__abc_21378_n4390;
  wire w_mem_inst__abc_21378_n4392;
  wire w_mem_inst__abc_21378_n4393;
  wire w_mem_inst__abc_21378_n4394;
  wire w_mem_inst__abc_21378_n4395;
  wire w_mem_inst__abc_21378_n4396;
  wire w_mem_inst__abc_21378_n4398;
  wire w_mem_inst__abc_21378_n4399;
  wire w_mem_inst__abc_21378_n4400;
  wire w_mem_inst__abc_21378_n4401;
  wire w_mem_inst__abc_21378_n4402;
  wire w_mem_inst__abc_21378_n4404;
  wire w_mem_inst__abc_21378_n4405;
  wire w_mem_inst__abc_21378_n4406;
  wire w_mem_inst__abc_21378_n4407;
  wire w_mem_inst__abc_21378_n4408;
  wire w_mem_inst__abc_21378_n4410;
  wire w_mem_inst__abc_21378_n4411;
  wire w_mem_inst__abc_21378_n4412;
  wire w_mem_inst__abc_21378_n4413;
  wire w_mem_inst__abc_21378_n4414;
  wire w_mem_inst__abc_21378_n4416;
  wire w_mem_inst__abc_21378_n4417;
  wire w_mem_inst__abc_21378_n4418;
  wire w_mem_inst__abc_21378_n4419;
  wire w_mem_inst__abc_21378_n4420;
  wire w_mem_inst__abc_21378_n4422;
  wire w_mem_inst__abc_21378_n4423;
  wire w_mem_inst__abc_21378_n4424;
  wire w_mem_inst__abc_21378_n4425;
  wire w_mem_inst__abc_21378_n4426;
  wire w_mem_inst__abc_21378_n4428;
  wire w_mem_inst__abc_21378_n4429;
  wire w_mem_inst__abc_21378_n4430;
  wire w_mem_inst__abc_21378_n4431;
  wire w_mem_inst__abc_21378_n4432;
  wire w_mem_inst__abc_21378_n4434;
  wire w_mem_inst__abc_21378_n4435;
  wire w_mem_inst__abc_21378_n4436;
  wire w_mem_inst__abc_21378_n4437;
  wire w_mem_inst__abc_21378_n4438;
  wire w_mem_inst__abc_21378_n4440;
  wire w_mem_inst__abc_21378_n4441;
  wire w_mem_inst__abc_21378_n4442;
  wire w_mem_inst__abc_21378_n4443;
  wire w_mem_inst__abc_21378_n4444;
  wire w_mem_inst__abc_21378_n4446;
  wire w_mem_inst__abc_21378_n4447;
  wire w_mem_inst__abc_21378_n4448;
  wire w_mem_inst__abc_21378_n4449;
  wire w_mem_inst__abc_21378_n4450;
  wire w_mem_inst__abc_21378_n4452;
  wire w_mem_inst__abc_21378_n4453;
  wire w_mem_inst__abc_21378_n4454;
  wire w_mem_inst__abc_21378_n4455;
  wire w_mem_inst__abc_21378_n4456;
  wire w_mem_inst__abc_21378_n4458;
  wire w_mem_inst__abc_21378_n4459;
  wire w_mem_inst__abc_21378_n4460;
  wire w_mem_inst__abc_21378_n4461;
  wire w_mem_inst__abc_21378_n4462;
  wire w_mem_inst__abc_21378_n4464;
  wire w_mem_inst__abc_21378_n4465;
  wire w_mem_inst__abc_21378_n4466;
  wire w_mem_inst__abc_21378_n4467;
  wire w_mem_inst__abc_21378_n4468;
  wire w_mem_inst__abc_21378_n4470;
  wire w_mem_inst__abc_21378_n4471;
  wire w_mem_inst__abc_21378_n4472;
  wire w_mem_inst__abc_21378_n4473;
  wire w_mem_inst__abc_21378_n4474;
  wire w_mem_inst__abc_21378_n4476;
  wire w_mem_inst__abc_21378_n4477;
  wire w_mem_inst__abc_21378_n4478;
  wire w_mem_inst__abc_21378_n4479;
  wire w_mem_inst__abc_21378_n4480;
  wire w_mem_inst__abc_21378_n4482;
  wire w_mem_inst__abc_21378_n4483;
  wire w_mem_inst__abc_21378_n4484;
  wire w_mem_inst__abc_21378_n4485;
  wire w_mem_inst__abc_21378_n4486;
  wire w_mem_inst__abc_21378_n4488;
  wire w_mem_inst__abc_21378_n4489;
  wire w_mem_inst__abc_21378_n4490;
  wire w_mem_inst__abc_21378_n4491;
  wire w_mem_inst__abc_21378_n4492;
  wire w_mem_inst__abc_21378_n4494;
  wire w_mem_inst__abc_21378_n4495;
  wire w_mem_inst__abc_21378_n4496;
  wire w_mem_inst__abc_21378_n4497;
  wire w_mem_inst__abc_21378_n4498;
  wire w_mem_inst__abc_21378_n4500;
  wire w_mem_inst__abc_21378_n4501;
  wire w_mem_inst__abc_21378_n4502;
  wire w_mem_inst__abc_21378_n4503;
  wire w_mem_inst__abc_21378_n4504;
  wire w_mem_inst__abc_21378_n4506;
  wire w_mem_inst__abc_21378_n4507;
  wire w_mem_inst__abc_21378_n4508;
  wire w_mem_inst__abc_21378_n4509;
  wire w_mem_inst__abc_21378_n4510;
  wire w_mem_inst__abc_21378_n4512;
  wire w_mem_inst__abc_21378_n4513;
  wire w_mem_inst__abc_21378_n4514;
  wire w_mem_inst__abc_21378_n4515;
  wire w_mem_inst__abc_21378_n4516;
  wire w_mem_inst__abc_21378_n4518;
  wire w_mem_inst__abc_21378_n4519;
  wire w_mem_inst__abc_21378_n4520;
  wire w_mem_inst__abc_21378_n4521;
  wire w_mem_inst__abc_21378_n4522;
  wire w_mem_inst__abc_21378_n4524;
  wire w_mem_inst__abc_21378_n4525;
  wire w_mem_inst__abc_21378_n4526;
  wire w_mem_inst__abc_21378_n4527;
  wire w_mem_inst__abc_21378_n4528;
  wire w_mem_inst__abc_21378_n4530;
  wire w_mem_inst__abc_21378_n4531;
  wire w_mem_inst__abc_21378_n4532;
  wire w_mem_inst__abc_21378_n4533;
  wire w_mem_inst__abc_21378_n4534;
  wire w_mem_inst__abc_21378_n4536;
  wire w_mem_inst__abc_21378_n4537;
  wire w_mem_inst__abc_21378_n4538;
  wire w_mem_inst__abc_21378_n4539;
  wire w_mem_inst__abc_21378_n4540;
  wire w_mem_inst__abc_21378_n4542;
  wire w_mem_inst__abc_21378_n4543;
  wire w_mem_inst__abc_21378_n4544;
  wire w_mem_inst__abc_21378_n4545;
  wire w_mem_inst__abc_21378_n4546;
  wire w_mem_inst__abc_21378_n4548;
  wire w_mem_inst__abc_21378_n4549;
  wire w_mem_inst__abc_21378_n4550;
  wire w_mem_inst__abc_21378_n4551;
  wire w_mem_inst__abc_21378_n4552;
  wire w_mem_inst__abc_21378_n4554;
  wire w_mem_inst__abc_21378_n4555;
  wire w_mem_inst__abc_21378_n4556;
  wire w_mem_inst__abc_21378_n4557;
  wire w_mem_inst__abc_21378_n4558;
  wire w_mem_inst__abc_21378_n4560;
  wire w_mem_inst__abc_21378_n4561;
  wire w_mem_inst__abc_21378_n4562;
  wire w_mem_inst__abc_21378_n4563;
  wire w_mem_inst__abc_21378_n4564;
  wire w_mem_inst__abc_21378_n4566;
  wire w_mem_inst__abc_21378_n4567;
  wire w_mem_inst__abc_21378_n4568;
  wire w_mem_inst__abc_21378_n4569;
  wire w_mem_inst__abc_21378_n4570;
  wire w_mem_inst__abc_21378_n4572;
  wire w_mem_inst__abc_21378_n4573;
  wire w_mem_inst__abc_21378_n4574;
  wire w_mem_inst__abc_21378_n4575;
  wire w_mem_inst__abc_21378_n4576;
  wire w_mem_inst__abc_21378_n4578;
  wire w_mem_inst__abc_21378_n4579;
  wire w_mem_inst__abc_21378_n4580;
  wire w_mem_inst__abc_21378_n4581;
  wire w_mem_inst__abc_21378_n4582;
  wire w_mem_inst__abc_21378_n4584;
  wire w_mem_inst__abc_21378_n4585;
  wire w_mem_inst__abc_21378_n4586;
  wire w_mem_inst__abc_21378_n4587;
  wire w_mem_inst__abc_21378_n4588;
  wire w_mem_inst__abc_21378_n4590;
  wire w_mem_inst__abc_21378_n4591;
  wire w_mem_inst__abc_21378_n4592;
  wire w_mem_inst__abc_21378_n4593;
  wire w_mem_inst__abc_21378_n4594;
  wire w_mem_inst__abc_21378_n4596;
  wire w_mem_inst__abc_21378_n4597;
  wire w_mem_inst__abc_21378_n4598;
  wire w_mem_inst__abc_21378_n4599;
  wire w_mem_inst__abc_21378_n4600;
  wire w_mem_inst__abc_21378_n4602;
  wire w_mem_inst__abc_21378_n4603;
  wire w_mem_inst__abc_21378_n4604;
  wire w_mem_inst__abc_21378_n4605;
  wire w_mem_inst__abc_21378_n4606;
  wire w_mem_inst__abc_21378_n4608;
  wire w_mem_inst__abc_21378_n4609;
  wire w_mem_inst__abc_21378_n4610;
  wire w_mem_inst__abc_21378_n4611;
  wire w_mem_inst__abc_21378_n4612;
  wire w_mem_inst__abc_21378_n4614;
  wire w_mem_inst__abc_21378_n4615;
  wire w_mem_inst__abc_21378_n4616;
  wire w_mem_inst__abc_21378_n4617;
  wire w_mem_inst__abc_21378_n4618;
  wire w_mem_inst__abc_21378_n4620;
  wire w_mem_inst__abc_21378_n4621;
  wire w_mem_inst__abc_21378_n4622;
  wire w_mem_inst__abc_21378_n4623;
  wire w_mem_inst__abc_21378_n4624;
  wire w_mem_inst__abc_21378_n4626;
  wire w_mem_inst__abc_21378_n4627;
  wire w_mem_inst__abc_21378_n4628;
  wire w_mem_inst__abc_21378_n4629;
  wire w_mem_inst__abc_21378_n4630;
  wire w_mem_inst__abc_21378_n4632;
  wire w_mem_inst__abc_21378_n4633;
  wire w_mem_inst__abc_21378_n4634;
  wire w_mem_inst__abc_21378_n4635;
  wire w_mem_inst__abc_21378_n4636;
  wire w_mem_inst__abc_21378_n4638;
  wire w_mem_inst__abc_21378_n4639;
  wire w_mem_inst__abc_21378_n4640;
  wire w_mem_inst__abc_21378_n4641;
  wire w_mem_inst__abc_21378_n4642;
  wire w_mem_inst__abc_21378_n4644;
  wire w_mem_inst__abc_21378_n4645;
  wire w_mem_inst__abc_21378_n4646;
  wire w_mem_inst__abc_21378_n4647;
  wire w_mem_inst__abc_21378_n4648;
  wire w_mem_inst__abc_21378_n4650;
  wire w_mem_inst__abc_21378_n4651;
  wire w_mem_inst__abc_21378_n4652;
  wire w_mem_inst__abc_21378_n4653;
  wire w_mem_inst__abc_21378_n4654;
  wire w_mem_inst__abc_21378_n4656;
  wire w_mem_inst__abc_21378_n4657;
  wire w_mem_inst__abc_21378_n4658;
  wire w_mem_inst__abc_21378_n4659;
  wire w_mem_inst__abc_21378_n4660;
  wire w_mem_inst__abc_21378_n4662;
  wire w_mem_inst__abc_21378_n4663;
  wire w_mem_inst__abc_21378_n4664;
  wire w_mem_inst__abc_21378_n4665;
  wire w_mem_inst__abc_21378_n4666;
  wire w_mem_inst__abc_21378_n4668;
  wire w_mem_inst__abc_21378_n4669;
  wire w_mem_inst__abc_21378_n4670;
  wire w_mem_inst__abc_21378_n4671;
  wire w_mem_inst__abc_21378_n4672;
  wire w_mem_inst__abc_21378_n4674;
  wire w_mem_inst__abc_21378_n4675;
  wire w_mem_inst__abc_21378_n4676;
  wire w_mem_inst__abc_21378_n4677;
  wire w_mem_inst__abc_21378_n4678;
  wire w_mem_inst__abc_21378_n4680;
  wire w_mem_inst__abc_21378_n4681;
  wire w_mem_inst__abc_21378_n4682;
  wire w_mem_inst__abc_21378_n4683;
  wire w_mem_inst__abc_21378_n4684;
  wire w_mem_inst__abc_21378_n4686;
  wire w_mem_inst__abc_21378_n4687;
  wire w_mem_inst__abc_21378_n4688;
  wire w_mem_inst__abc_21378_n4689;
  wire w_mem_inst__abc_21378_n4690;
  wire w_mem_inst__abc_21378_n4692;
  wire w_mem_inst__abc_21378_n4693;
  wire w_mem_inst__abc_21378_n4694;
  wire w_mem_inst__abc_21378_n4695;
  wire w_mem_inst__abc_21378_n4696;
  wire w_mem_inst__abc_21378_n4698;
  wire w_mem_inst__abc_21378_n4699;
  wire w_mem_inst__abc_21378_n4700;
  wire w_mem_inst__abc_21378_n4701;
  wire w_mem_inst__abc_21378_n4702;
  wire w_mem_inst__abc_21378_n4704;
  wire w_mem_inst__abc_21378_n4705;
  wire w_mem_inst__abc_21378_n4706;
  wire w_mem_inst__abc_21378_n4707;
  wire w_mem_inst__abc_21378_n4708;
  wire w_mem_inst__abc_21378_n4710;
  wire w_mem_inst__abc_21378_n4711;
  wire w_mem_inst__abc_21378_n4712;
  wire w_mem_inst__abc_21378_n4713;
  wire w_mem_inst__abc_21378_n4714;
  wire w_mem_inst__abc_21378_n4716;
  wire w_mem_inst__abc_21378_n4717;
  wire w_mem_inst__abc_21378_n4718;
  wire w_mem_inst__abc_21378_n4719;
  wire w_mem_inst__abc_21378_n4720;
  wire w_mem_inst__abc_21378_n4722;
  wire w_mem_inst__abc_21378_n4723;
  wire w_mem_inst__abc_21378_n4724;
  wire w_mem_inst__abc_21378_n4725;
  wire w_mem_inst__abc_21378_n4726;
  wire w_mem_inst__abc_21378_n4728;
  wire w_mem_inst__abc_21378_n4729;
  wire w_mem_inst__abc_21378_n4730;
  wire w_mem_inst__abc_21378_n4731;
  wire w_mem_inst__abc_21378_n4732;
  wire w_mem_inst__abc_21378_n4734;
  wire w_mem_inst__abc_21378_n4735;
  wire w_mem_inst__abc_21378_n4736;
  wire w_mem_inst__abc_21378_n4737;
  wire w_mem_inst__abc_21378_n4738;
  wire w_mem_inst__abc_21378_n4740;
  wire w_mem_inst__abc_21378_n4741;
  wire w_mem_inst__abc_21378_n4742;
  wire w_mem_inst__abc_21378_n4743;
  wire w_mem_inst__abc_21378_n4744;
  wire w_mem_inst__abc_21378_n4746;
  wire w_mem_inst__abc_21378_n4747;
  wire w_mem_inst__abc_21378_n4748;
  wire w_mem_inst__abc_21378_n4749;
  wire w_mem_inst__abc_21378_n4750;
  wire w_mem_inst__abc_21378_n4752;
  wire w_mem_inst__abc_21378_n4753;
  wire w_mem_inst__abc_21378_n4754;
  wire w_mem_inst__abc_21378_n4755;
  wire w_mem_inst__abc_21378_n4756;
  wire w_mem_inst__abc_21378_n4758;
  wire w_mem_inst__abc_21378_n4759;
  wire w_mem_inst__abc_21378_n4760;
  wire w_mem_inst__abc_21378_n4761;
  wire w_mem_inst__abc_21378_n4762;
  wire w_mem_inst__abc_21378_n4764;
  wire w_mem_inst__abc_21378_n4765;
  wire w_mem_inst__abc_21378_n4766;
  wire w_mem_inst__abc_21378_n4767;
  wire w_mem_inst__abc_21378_n4768;
  wire w_mem_inst__abc_21378_n4770;
  wire w_mem_inst__abc_21378_n4771;
  wire w_mem_inst__abc_21378_n4772;
  wire w_mem_inst__abc_21378_n4773;
  wire w_mem_inst__abc_21378_n4774;
  wire w_mem_inst__abc_21378_n4776;
  wire w_mem_inst__abc_21378_n4777;
  wire w_mem_inst__abc_21378_n4778;
  wire w_mem_inst__abc_21378_n4779;
  wire w_mem_inst__abc_21378_n4780;
  wire w_mem_inst__abc_21378_n4782;
  wire w_mem_inst__abc_21378_n4783;
  wire w_mem_inst__abc_21378_n4784;
  wire w_mem_inst__abc_21378_n4785;
  wire w_mem_inst__abc_21378_n4786;
  wire w_mem_inst__abc_21378_n4788;
  wire w_mem_inst__abc_21378_n4789;
  wire w_mem_inst__abc_21378_n4790;
  wire w_mem_inst__abc_21378_n4791;
  wire w_mem_inst__abc_21378_n4792;
  wire w_mem_inst__abc_21378_n4794;
  wire w_mem_inst__abc_21378_n4795;
  wire w_mem_inst__abc_21378_n4796;
  wire w_mem_inst__abc_21378_n4797;
  wire w_mem_inst__abc_21378_n4798;
  wire w_mem_inst__abc_21378_n4800;
  wire w_mem_inst__abc_21378_n4801;
  wire w_mem_inst__abc_21378_n4802;
  wire w_mem_inst__abc_21378_n4803;
  wire w_mem_inst__abc_21378_n4804;
  wire w_mem_inst__abc_21378_n4806;
  wire w_mem_inst__abc_21378_n4807;
  wire w_mem_inst__abc_21378_n4808;
  wire w_mem_inst__abc_21378_n4809;
  wire w_mem_inst__abc_21378_n4810;
  wire w_mem_inst__abc_21378_n4812;
  wire w_mem_inst__abc_21378_n4813;
  wire w_mem_inst__abc_21378_n4814;
  wire w_mem_inst__abc_21378_n4815;
  wire w_mem_inst__abc_21378_n4816;
  wire w_mem_inst__abc_21378_n4818;
  wire w_mem_inst__abc_21378_n4819;
  wire w_mem_inst__abc_21378_n4820;
  wire w_mem_inst__abc_21378_n4821;
  wire w_mem_inst__abc_21378_n4822;
  wire w_mem_inst__abc_21378_n4824;
  wire w_mem_inst__abc_21378_n4825;
  wire w_mem_inst__abc_21378_n4826;
  wire w_mem_inst__abc_21378_n4827;
  wire w_mem_inst__abc_21378_n4828;
  wire w_mem_inst__abc_21378_n4830;
  wire w_mem_inst__abc_21378_n4831;
  wire w_mem_inst__abc_21378_n4832;
  wire w_mem_inst__abc_21378_n4833;
  wire w_mem_inst__abc_21378_n4834;
  wire w_mem_inst__abc_21378_n4836;
  wire w_mem_inst__abc_21378_n4837;
  wire w_mem_inst__abc_21378_n4838;
  wire w_mem_inst__abc_21378_n4839;
  wire w_mem_inst__abc_21378_n4840;
  wire w_mem_inst__abc_21378_n4842;
  wire w_mem_inst__abc_21378_n4843;
  wire w_mem_inst__abc_21378_n4844;
  wire w_mem_inst__abc_21378_n4845;
  wire w_mem_inst__abc_21378_n4846;
  wire w_mem_inst__abc_21378_n4848;
  wire w_mem_inst__abc_21378_n4849;
  wire w_mem_inst__abc_21378_n4850;
  wire w_mem_inst__abc_21378_n4851;
  wire w_mem_inst__abc_21378_n4852;
  wire w_mem_inst__abc_21378_n4854;
  wire w_mem_inst__abc_21378_n4855;
  wire w_mem_inst__abc_21378_n4856;
  wire w_mem_inst__abc_21378_n4857;
  wire w_mem_inst__abc_21378_n4858;
  wire w_mem_inst__abc_21378_n4860;
  wire w_mem_inst__abc_21378_n4861;
  wire w_mem_inst__abc_21378_n4862;
  wire w_mem_inst__abc_21378_n4863;
  wire w_mem_inst__abc_21378_n4864;
  wire w_mem_inst__abc_21378_n4866;
  wire w_mem_inst__abc_21378_n4867;
  wire w_mem_inst__abc_21378_n4868;
  wire w_mem_inst__abc_21378_n4869;
  wire w_mem_inst__abc_21378_n4870;
  wire w_mem_inst__abc_21378_n4872;
  wire w_mem_inst__abc_21378_n4873;
  wire w_mem_inst__abc_21378_n4874;
  wire w_mem_inst__abc_21378_n4875;
  wire w_mem_inst__abc_21378_n4876;
  wire w_mem_inst__abc_21378_n4878;
  wire w_mem_inst__abc_21378_n4879;
  wire w_mem_inst__abc_21378_n4880;
  wire w_mem_inst__abc_21378_n4881;
  wire w_mem_inst__abc_21378_n4882;
  wire w_mem_inst__abc_21378_n4884;
  wire w_mem_inst__abc_21378_n4885;
  wire w_mem_inst__abc_21378_n4886;
  wire w_mem_inst__abc_21378_n4887;
  wire w_mem_inst__abc_21378_n4888;
  wire w_mem_inst__abc_21378_n4890;
  wire w_mem_inst__abc_21378_n4891;
  wire w_mem_inst__abc_21378_n4892;
  wire w_mem_inst__abc_21378_n4893;
  wire w_mem_inst__abc_21378_n4894;
  wire w_mem_inst__abc_21378_n4896;
  wire w_mem_inst__abc_21378_n4897;
  wire w_mem_inst__abc_21378_n4898;
  wire w_mem_inst__abc_21378_n4899;
  wire w_mem_inst__abc_21378_n4900;
  wire w_mem_inst__abc_21378_n4902;
  wire w_mem_inst__abc_21378_n4903;
  wire w_mem_inst__abc_21378_n4904;
  wire w_mem_inst__abc_21378_n4905;
  wire w_mem_inst__abc_21378_n4906;
  wire w_mem_inst__abc_21378_n4908;
  wire w_mem_inst__abc_21378_n4909;
  wire w_mem_inst__abc_21378_n4910;
  wire w_mem_inst__abc_21378_n4911;
  wire w_mem_inst__abc_21378_n4912;
  wire w_mem_inst__abc_21378_n4914;
  wire w_mem_inst__abc_21378_n4915;
  wire w_mem_inst__abc_21378_n4916;
  wire w_mem_inst__abc_21378_n4917;
  wire w_mem_inst__abc_21378_n4918;
  wire w_mem_inst__abc_21378_n4920;
  wire w_mem_inst__abc_21378_n4921;
  wire w_mem_inst__abc_21378_n4922;
  wire w_mem_inst__abc_21378_n4923;
  wire w_mem_inst__abc_21378_n4924;
  wire w_mem_inst__abc_21378_n4926;
  wire w_mem_inst__abc_21378_n4927;
  wire w_mem_inst__abc_21378_n4928;
  wire w_mem_inst__abc_21378_n4929;
  wire w_mem_inst__abc_21378_n4930;
  wire w_mem_inst__abc_21378_n4932;
  wire w_mem_inst__abc_21378_n4933;
  wire w_mem_inst__abc_21378_n4934;
  wire w_mem_inst__abc_21378_n4935;
  wire w_mem_inst__abc_21378_n4936;
  wire w_mem_inst__abc_21378_n4938;
  wire w_mem_inst__abc_21378_n4939;
  wire w_mem_inst__abc_21378_n4940;
  wire w_mem_inst__abc_21378_n4941;
  wire w_mem_inst__abc_21378_n4942;
  wire w_mem_inst__abc_21378_n4944;
  wire w_mem_inst__abc_21378_n4945;
  wire w_mem_inst__abc_21378_n4946;
  wire w_mem_inst__abc_21378_n4947;
  wire w_mem_inst__abc_21378_n4948;
  wire w_mem_inst__abc_21378_n4950;
  wire w_mem_inst__abc_21378_n4951;
  wire w_mem_inst__abc_21378_n4952;
  wire w_mem_inst__abc_21378_n4953;
  wire w_mem_inst__abc_21378_n4954;
  wire w_mem_inst__abc_21378_n4956;
  wire w_mem_inst__abc_21378_n4957;
  wire w_mem_inst__abc_21378_n4958;
  wire w_mem_inst__abc_21378_n4959;
  wire w_mem_inst__abc_21378_n4960;
  wire w_mem_inst__abc_21378_n4962;
  wire w_mem_inst__abc_21378_n4963;
  wire w_mem_inst__abc_21378_n4964;
  wire w_mem_inst__abc_21378_n4965;
  wire w_mem_inst__abc_21378_n4966;
  wire w_mem_inst__abc_21378_n4968;
  wire w_mem_inst__abc_21378_n4969;
  wire w_mem_inst__abc_21378_n4970;
  wire w_mem_inst__abc_21378_n4971;
  wire w_mem_inst__abc_21378_n4972;
  wire w_mem_inst__abc_21378_n4974;
  wire w_mem_inst__abc_21378_n4975;
  wire w_mem_inst__abc_21378_n4976;
  wire w_mem_inst__abc_21378_n4977;
  wire w_mem_inst__abc_21378_n4978;
  wire w_mem_inst__abc_21378_n4980;
  wire w_mem_inst__abc_21378_n4981;
  wire w_mem_inst__abc_21378_n4982;
  wire w_mem_inst__abc_21378_n4983;
  wire w_mem_inst__abc_21378_n4984;
  wire w_mem_inst__abc_21378_n4986;
  wire w_mem_inst__abc_21378_n4987;
  wire w_mem_inst__abc_21378_n4988;
  wire w_mem_inst__abc_21378_n4989;
  wire w_mem_inst__abc_21378_n4990;
  wire w_mem_inst__abc_21378_n4992;
  wire w_mem_inst__abc_21378_n4993;
  wire w_mem_inst__abc_21378_n4994;
  wire w_mem_inst__abc_21378_n4995;
  wire w_mem_inst__abc_21378_n4996;
  wire w_mem_inst__abc_21378_n4998;
  wire w_mem_inst__abc_21378_n4999;
  wire w_mem_inst__abc_21378_n5000;
  wire w_mem_inst__abc_21378_n5001;
  wire w_mem_inst__abc_21378_n5002;
  wire w_mem_inst__abc_21378_n5004;
  wire w_mem_inst__abc_21378_n5005;
  wire w_mem_inst__abc_21378_n5006;
  wire w_mem_inst__abc_21378_n5007;
  wire w_mem_inst__abc_21378_n5008;
  wire w_mem_inst__abc_21378_n5010;
  wire w_mem_inst__abc_21378_n5011;
  wire w_mem_inst__abc_21378_n5012;
  wire w_mem_inst__abc_21378_n5013;
  wire w_mem_inst__abc_21378_n5014;
  wire w_mem_inst__abc_21378_n5016;
  wire w_mem_inst__abc_21378_n5017;
  wire w_mem_inst__abc_21378_n5018;
  wire w_mem_inst__abc_21378_n5019;
  wire w_mem_inst__abc_21378_n5020;
  wire w_mem_inst__abc_21378_n5022;
  wire w_mem_inst__abc_21378_n5023;
  wire w_mem_inst__abc_21378_n5024;
  wire w_mem_inst__abc_21378_n5025;
  wire w_mem_inst__abc_21378_n5026;
  wire w_mem_inst__abc_21378_n5028;
  wire w_mem_inst__abc_21378_n5029;
  wire w_mem_inst__abc_21378_n5030;
  wire w_mem_inst__abc_21378_n5031;
  wire w_mem_inst__abc_21378_n5032;
  wire w_mem_inst__abc_21378_n5034;
  wire w_mem_inst__abc_21378_n5035;
  wire w_mem_inst__abc_21378_n5036;
  wire w_mem_inst__abc_21378_n5037;
  wire w_mem_inst__abc_21378_n5038;
  wire w_mem_inst__abc_21378_n5040;
  wire w_mem_inst__abc_21378_n5041;
  wire w_mem_inst__abc_21378_n5042;
  wire w_mem_inst__abc_21378_n5043;
  wire w_mem_inst__abc_21378_n5044;
  wire w_mem_inst__abc_21378_n5046;
  wire w_mem_inst__abc_21378_n5047;
  wire w_mem_inst__abc_21378_n5048;
  wire w_mem_inst__abc_21378_n5049;
  wire w_mem_inst__abc_21378_n5050;
  wire w_mem_inst__abc_21378_n5052;
  wire w_mem_inst__abc_21378_n5053;
  wire w_mem_inst__abc_21378_n5054;
  wire w_mem_inst__abc_21378_n5055;
  wire w_mem_inst__abc_21378_n5056;
  wire w_mem_inst__abc_21378_n5058;
  wire w_mem_inst__abc_21378_n5059;
  wire w_mem_inst__abc_21378_n5060;
  wire w_mem_inst__abc_21378_n5061;
  wire w_mem_inst__abc_21378_n5062;
  wire w_mem_inst__abc_21378_n5064;
  wire w_mem_inst__abc_21378_n5065;
  wire w_mem_inst__abc_21378_n5066;
  wire w_mem_inst__abc_21378_n5067;
  wire w_mem_inst__abc_21378_n5068;
  wire w_mem_inst__abc_21378_n5070;
  wire w_mem_inst__abc_21378_n5071;
  wire w_mem_inst__abc_21378_n5072;
  wire w_mem_inst__abc_21378_n5073;
  wire w_mem_inst__abc_21378_n5074;
  wire w_mem_inst__abc_21378_n5076;
  wire w_mem_inst__abc_21378_n5077;
  wire w_mem_inst__abc_21378_n5078;
  wire w_mem_inst__abc_21378_n5079;
  wire w_mem_inst__abc_21378_n5080;
  wire w_mem_inst__abc_21378_n5082;
  wire w_mem_inst__abc_21378_n5083;
  wire w_mem_inst__abc_21378_n5084;
  wire w_mem_inst__abc_21378_n5085;
  wire w_mem_inst__abc_21378_n5086;
  wire w_mem_inst__abc_21378_n5088;
  wire w_mem_inst__abc_21378_n5089;
  wire w_mem_inst__abc_21378_n5090;
  wire w_mem_inst__abc_21378_n5091;
  wire w_mem_inst__abc_21378_n5092;
  wire w_mem_inst__abc_21378_n5094;
  wire w_mem_inst__abc_21378_n5095;
  wire w_mem_inst__abc_21378_n5096;
  wire w_mem_inst__abc_21378_n5097;
  wire w_mem_inst__abc_21378_n5098;
  wire w_mem_inst__abc_21378_n5100;
  wire w_mem_inst__abc_21378_n5101;
  wire w_mem_inst__abc_21378_n5102;
  wire w_mem_inst__abc_21378_n5103;
  wire w_mem_inst__abc_21378_n5104;
  wire w_mem_inst__abc_21378_n5106;
  wire w_mem_inst__abc_21378_n5107;
  wire w_mem_inst__abc_21378_n5108;
  wire w_mem_inst__abc_21378_n5109;
  wire w_mem_inst__abc_21378_n5110;
  wire w_mem_inst__abc_21378_n5112;
  wire w_mem_inst__abc_21378_n5113;
  wire w_mem_inst__abc_21378_n5114;
  wire w_mem_inst__abc_21378_n5115;
  wire w_mem_inst__abc_21378_n5116;
  wire w_mem_inst__abc_21378_n5118;
  wire w_mem_inst__abc_21378_n5119;
  wire w_mem_inst__abc_21378_n5120;
  wire w_mem_inst__abc_21378_n5121;
  wire w_mem_inst__abc_21378_n5122;
  wire w_mem_inst__abc_21378_n5124;
  wire w_mem_inst__abc_21378_n5125;
  wire w_mem_inst__abc_21378_n5126;
  wire w_mem_inst__abc_21378_n5127;
  wire w_mem_inst__abc_21378_n5128;
  wire w_mem_inst__abc_21378_n5130;
  wire w_mem_inst__abc_21378_n5131;
  wire w_mem_inst__abc_21378_n5132;
  wire w_mem_inst__abc_21378_n5133;
  wire w_mem_inst__abc_21378_n5134;
  wire w_mem_inst__abc_21378_n5136;
  wire w_mem_inst__abc_21378_n5137;
  wire w_mem_inst__abc_21378_n5138;
  wire w_mem_inst__abc_21378_n5139;
  wire w_mem_inst__abc_21378_n5140;
  wire w_mem_inst__abc_21378_n5142;
  wire w_mem_inst__abc_21378_n5143;
  wire w_mem_inst__abc_21378_n5144;
  wire w_mem_inst__abc_21378_n5145;
  wire w_mem_inst__abc_21378_n5146;
  wire w_mem_inst__abc_21378_n5148;
  wire w_mem_inst__abc_21378_n5149;
  wire w_mem_inst__abc_21378_n5150;
  wire w_mem_inst__abc_21378_n5151;
  wire w_mem_inst__abc_21378_n5152;
  wire w_mem_inst__abc_21378_n5154;
  wire w_mem_inst__abc_21378_n5155;
  wire w_mem_inst__abc_21378_n5156;
  wire w_mem_inst__abc_21378_n5157;
  wire w_mem_inst__abc_21378_n5158;
  wire w_mem_inst__abc_21378_n5160;
  wire w_mem_inst__abc_21378_n5161;
  wire w_mem_inst__abc_21378_n5162;
  wire w_mem_inst__abc_21378_n5163;
  wire w_mem_inst__abc_21378_n5164;
  wire w_mem_inst__abc_21378_n5166;
  wire w_mem_inst__abc_21378_n5167;
  wire w_mem_inst__abc_21378_n5168;
  wire w_mem_inst__abc_21378_n5169;
  wire w_mem_inst__abc_21378_n5170;
  wire w_mem_inst__abc_21378_n5172;
  wire w_mem_inst__abc_21378_n5173;
  wire w_mem_inst__abc_21378_n5174;
  wire w_mem_inst__abc_21378_n5175;
  wire w_mem_inst__abc_21378_n5176;
  wire w_mem_inst__abc_21378_n5178;
  wire w_mem_inst__abc_21378_n5179;
  wire w_mem_inst__abc_21378_n5180;
  wire w_mem_inst__abc_21378_n5181;
  wire w_mem_inst__abc_21378_n5182;
  wire w_mem_inst__abc_21378_n5184;
  wire w_mem_inst__abc_21378_n5185;
  wire w_mem_inst__abc_21378_n5186;
  wire w_mem_inst__abc_21378_n5187;
  wire w_mem_inst__abc_21378_n5188;
  wire w_mem_inst__abc_21378_n5190;
  wire w_mem_inst__abc_21378_n5191;
  wire w_mem_inst__abc_21378_n5192;
  wire w_mem_inst__abc_21378_n5193;
  wire w_mem_inst__abc_21378_n5194;
  wire w_mem_inst__abc_21378_n5196;
  wire w_mem_inst__abc_21378_n5197;
  wire w_mem_inst__abc_21378_n5198;
  wire w_mem_inst__abc_21378_n5199;
  wire w_mem_inst__abc_21378_n5200;
  wire w_mem_inst__abc_21378_n5202;
  wire w_mem_inst__abc_21378_n5203;
  wire w_mem_inst__abc_21378_n5204;
  wire w_mem_inst__abc_21378_n5205;
  wire w_mem_inst__abc_21378_n5206;
  wire w_mem_inst__abc_21378_n5208;
  wire w_mem_inst__abc_21378_n5209;
  wire w_mem_inst__abc_21378_n5210;
  wire w_mem_inst__abc_21378_n5211;
  wire w_mem_inst__abc_21378_n5212;
  wire w_mem_inst__abc_21378_n5214;
  wire w_mem_inst__abc_21378_n5215;
  wire w_mem_inst__abc_21378_n5216;
  wire w_mem_inst__abc_21378_n5217;
  wire w_mem_inst__abc_21378_n5218;
  wire w_mem_inst__abc_21378_n5220;
  wire w_mem_inst__abc_21378_n5221;
  wire w_mem_inst__abc_21378_n5222;
  wire w_mem_inst__abc_21378_n5223;
  wire w_mem_inst__abc_21378_n5224;
  wire w_mem_inst__abc_21378_n5226;
  wire w_mem_inst__abc_21378_n5227;
  wire w_mem_inst__abc_21378_n5228;
  wire w_mem_inst__abc_21378_n5229;
  wire w_mem_inst__abc_21378_n5230;
  wire w_mem_inst__abc_21378_n5232;
  wire w_mem_inst__abc_21378_n5233;
  wire w_mem_inst__abc_21378_n5234;
  wire w_mem_inst__abc_21378_n5235;
  wire w_mem_inst__abc_21378_n5236;
  wire w_mem_inst__abc_21378_n5238;
  wire w_mem_inst__abc_21378_n5239;
  wire w_mem_inst__abc_21378_n5240;
  wire w_mem_inst__abc_21378_n5241;
  wire w_mem_inst__abc_21378_n5242;
  wire w_mem_inst__abc_21378_n5244;
  wire w_mem_inst__abc_21378_n5245;
  wire w_mem_inst__abc_21378_n5246;
  wire w_mem_inst__abc_21378_n5247;
  wire w_mem_inst__abc_21378_n5248;
  wire w_mem_inst__abc_21378_n5250;
  wire w_mem_inst__abc_21378_n5251;
  wire w_mem_inst__abc_21378_n5252;
  wire w_mem_inst__abc_21378_n5253;
  wire w_mem_inst__abc_21378_n5254;
  wire w_mem_inst__abc_21378_n5256;
  wire w_mem_inst__abc_21378_n5257;
  wire w_mem_inst__abc_21378_n5258;
  wire w_mem_inst__abc_21378_n5259;
  wire w_mem_inst__abc_21378_n5260;
  wire w_mem_inst__abc_21378_n5262;
  wire w_mem_inst__abc_21378_n5263;
  wire w_mem_inst__abc_21378_n5264;
  wire w_mem_inst__abc_21378_n5265;
  wire w_mem_inst__abc_21378_n5266;
  wire w_mem_inst__abc_21378_n5268;
  wire w_mem_inst__abc_21378_n5269;
  wire w_mem_inst__abc_21378_n5270;
  wire w_mem_inst__abc_21378_n5271;
  wire w_mem_inst__abc_21378_n5272;
  wire w_mem_inst__abc_21378_n5274;
  wire w_mem_inst__abc_21378_n5275;
  wire w_mem_inst__abc_21378_n5276;
  wire w_mem_inst__abc_21378_n5277;
  wire w_mem_inst__abc_21378_n5278;
  wire w_mem_inst__abc_21378_n5280;
  wire w_mem_inst__abc_21378_n5281;
  wire w_mem_inst__abc_21378_n5282;
  wire w_mem_inst__abc_21378_n5283;
  wire w_mem_inst__abc_21378_n5284;
  wire w_mem_inst__abc_21378_n5286;
  wire w_mem_inst__abc_21378_n5287;
  wire w_mem_inst__abc_21378_n5288;
  wire w_mem_inst__abc_21378_n5289;
  wire w_mem_inst__abc_21378_n5290;
  wire w_mem_inst__abc_21378_n5292;
  wire w_mem_inst__abc_21378_n5293;
  wire w_mem_inst__abc_21378_n5294;
  wire w_mem_inst__abc_21378_n5295;
  wire w_mem_inst__abc_21378_n5296;
  wire w_mem_inst__abc_21378_n5298;
  wire w_mem_inst__abc_21378_n5299;
  wire w_mem_inst__abc_21378_n5300;
  wire w_mem_inst__abc_21378_n5301;
  wire w_mem_inst__abc_21378_n5302;
  wire w_mem_inst__abc_21378_n5304;
  wire w_mem_inst__abc_21378_n5305;
  wire w_mem_inst__abc_21378_n5306;
  wire w_mem_inst__abc_21378_n5307;
  wire w_mem_inst__abc_21378_n5308;
  wire w_mem_inst__abc_21378_n5310;
  wire w_mem_inst__abc_21378_n5311;
  wire w_mem_inst__abc_21378_n5312;
  wire w_mem_inst__abc_21378_n5313;
  wire w_mem_inst__abc_21378_n5314;
  wire w_mem_inst__abc_21378_n5316;
  wire w_mem_inst__abc_21378_n5317;
  wire w_mem_inst__abc_21378_n5318;
  wire w_mem_inst__abc_21378_n5319;
  wire w_mem_inst__abc_21378_n5320;
  wire w_mem_inst__abc_21378_n5322;
  wire w_mem_inst__abc_21378_n5323;
  wire w_mem_inst__abc_21378_n5324;
  wire w_mem_inst__abc_21378_n5325;
  wire w_mem_inst__abc_21378_n5326;
  wire w_mem_inst__abc_21378_n5328;
  wire w_mem_inst__abc_21378_n5329;
  wire w_mem_inst__abc_21378_n5330;
  wire w_mem_inst__abc_21378_n5331;
  wire w_mem_inst__abc_21378_n5332;
  wire w_mem_inst__abc_21378_n5334;
  wire w_mem_inst__abc_21378_n5335;
  wire w_mem_inst__abc_21378_n5336;
  wire w_mem_inst__abc_21378_n5337;
  wire w_mem_inst__abc_21378_n5338;
  wire w_mem_inst__abc_21378_n5340;
  wire w_mem_inst__abc_21378_n5341;
  wire w_mem_inst__abc_21378_n5342;
  wire w_mem_inst__abc_21378_n5343;
  wire w_mem_inst__abc_21378_n5344;
  wire w_mem_inst__abc_21378_n5346;
  wire w_mem_inst__abc_21378_n5347;
  wire w_mem_inst__abc_21378_n5348;
  wire w_mem_inst__abc_21378_n5349;
  wire w_mem_inst__abc_21378_n5350;
  wire w_mem_inst__abc_21378_n5352;
  wire w_mem_inst__abc_21378_n5353;
  wire w_mem_inst__abc_21378_n5354;
  wire w_mem_inst__abc_21378_n5355;
  wire w_mem_inst__abc_21378_n5356;
  wire w_mem_inst__abc_21378_n5358;
  wire w_mem_inst__abc_21378_n5359;
  wire w_mem_inst__abc_21378_n5360;
  wire w_mem_inst__abc_21378_n5361;
  wire w_mem_inst__abc_21378_n5362;
  wire w_mem_inst__abc_21378_n5364;
  wire w_mem_inst__abc_21378_n5365;
  wire w_mem_inst__abc_21378_n5366;
  wire w_mem_inst__abc_21378_n5367;
  wire w_mem_inst__abc_21378_n5368;
  wire w_mem_inst__abc_21378_n5370;
  wire w_mem_inst__abc_21378_n5371;
  wire w_mem_inst__abc_21378_n5372;
  wire w_mem_inst__abc_21378_n5373;
  wire w_mem_inst__abc_21378_n5374;
  wire w_mem_inst__abc_21378_n5376;
  wire w_mem_inst__abc_21378_n5377;
  wire w_mem_inst__abc_21378_n5378;
  wire w_mem_inst__abc_21378_n5379;
  wire w_mem_inst__abc_21378_n5380;
  wire w_mem_inst__abc_21378_n5382;
  wire w_mem_inst__abc_21378_n5383;
  wire w_mem_inst__abc_21378_n5384;
  wire w_mem_inst__abc_21378_n5385;
  wire w_mem_inst__abc_21378_n5386;
  wire w_mem_inst__abc_21378_n5388;
  wire w_mem_inst__abc_21378_n5389;
  wire w_mem_inst__abc_21378_n5390;
  wire w_mem_inst__abc_21378_n5391;
  wire w_mem_inst__abc_21378_n5392;
  wire w_mem_inst__abc_21378_n5394;
  wire w_mem_inst__abc_21378_n5395;
  wire w_mem_inst__abc_21378_n5396;
  wire w_mem_inst__abc_21378_n5397;
  wire w_mem_inst__abc_21378_n5398;
  wire w_mem_inst__abc_21378_n5400;
  wire w_mem_inst__abc_21378_n5401;
  wire w_mem_inst__abc_21378_n5402;
  wire w_mem_inst__abc_21378_n5403;
  wire w_mem_inst__abc_21378_n5404;
  wire w_mem_inst__abc_21378_n5406;
  wire w_mem_inst__abc_21378_n5407;
  wire w_mem_inst__abc_21378_n5408;
  wire w_mem_inst__abc_21378_n5409;
  wire w_mem_inst__abc_21378_n5410;
  wire w_mem_inst__abc_21378_n5412;
  wire w_mem_inst__abc_21378_n5413;
  wire w_mem_inst__abc_21378_n5414;
  wire w_mem_inst__abc_21378_n5415;
  wire w_mem_inst__abc_21378_n5416;
  wire w_mem_inst__abc_21378_n5418;
  wire w_mem_inst__abc_21378_n5419;
  wire w_mem_inst__abc_21378_n5420;
  wire w_mem_inst__abc_21378_n5421;
  wire w_mem_inst__abc_21378_n5422;
  wire w_mem_inst__abc_21378_n5424;
  wire w_mem_inst__abc_21378_n5425;
  wire w_mem_inst__abc_21378_n5426;
  wire w_mem_inst__abc_21378_n5427;
  wire w_mem_inst__abc_21378_n5428;
  wire w_mem_inst__abc_21378_n5430;
  wire w_mem_inst__abc_21378_n5431;
  wire w_mem_inst__abc_21378_n5432;
  wire w_mem_inst__abc_21378_n5433;
  wire w_mem_inst__abc_21378_n5434;
  wire w_mem_inst__abc_21378_n5436;
  wire w_mem_inst__abc_21378_n5437;
  wire w_mem_inst__abc_21378_n5438;
  wire w_mem_inst__abc_21378_n5439;
  wire w_mem_inst__abc_21378_n5440;
  wire w_mem_inst__abc_21378_n5442;
  wire w_mem_inst__abc_21378_n5443;
  wire w_mem_inst__abc_21378_n5444;
  wire w_mem_inst__abc_21378_n5445;
  wire w_mem_inst__abc_21378_n5446;
  wire w_mem_inst__abc_21378_n5448;
  wire w_mem_inst__abc_21378_n5449;
  wire w_mem_inst__abc_21378_n5450;
  wire w_mem_inst__abc_21378_n5451;
  wire w_mem_inst__abc_21378_n5452;
  wire w_mem_inst__abc_21378_n5454;
  wire w_mem_inst__abc_21378_n5455;
  wire w_mem_inst__abc_21378_n5456;
  wire w_mem_inst__abc_21378_n5457;
  wire w_mem_inst__abc_21378_n5458;
  wire w_mem_inst__abc_21378_n5460;
  wire w_mem_inst__abc_21378_n5461;
  wire w_mem_inst__abc_21378_n5462;
  wire w_mem_inst__abc_21378_n5463;
  wire w_mem_inst__abc_21378_n5464;
  wire w_mem_inst__abc_21378_n5466;
  wire w_mem_inst__abc_21378_n5467;
  wire w_mem_inst__abc_21378_n5468;
  wire w_mem_inst__abc_21378_n5469;
  wire w_mem_inst__abc_21378_n5470;
  wire w_mem_inst__abc_21378_n5472;
  wire w_mem_inst__abc_21378_n5473;
  wire w_mem_inst__abc_21378_n5474;
  wire w_mem_inst__abc_21378_n5475;
  wire w_mem_inst__abc_21378_n5476;
  wire w_mem_inst__abc_21378_n5478;
  wire w_mem_inst__abc_21378_n5479;
  wire w_mem_inst__abc_21378_n5480;
  wire w_mem_inst__abc_21378_n5481;
  wire w_mem_inst__abc_21378_n5482;
  wire w_mem_inst__abc_21378_n5484;
  wire w_mem_inst__abc_21378_n5485;
  wire w_mem_inst__abc_21378_n5486;
  wire w_mem_inst__abc_21378_n5487;
  wire w_mem_inst__abc_21378_n5488;
  wire w_mem_inst__abc_21378_n5490;
  wire w_mem_inst__abc_21378_n5491;
  wire w_mem_inst__abc_21378_n5492;
  wire w_mem_inst__abc_21378_n5493;
  wire w_mem_inst__abc_21378_n5494;
  wire w_mem_inst__abc_21378_n5496;
  wire w_mem_inst__abc_21378_n5497;
  wire w_mem_inst__abc_21378_n5498;
  wire w_mem_inst__abc_21378_n5499;
  wire w_mem_inst__abc_21378_n5500;
  wire w_mem_inst__abc_21378_n5502;
  wire w_mem_inst__abc_21378_n5503;
  wire w_mem_inst__abc_21378_n5504;
  wire w_mem_inst__abc_21378_n5505;
  wire w_mem_inst__abc_21378_n5506;
  wire w_mem_inst__abc_21378_n5508;
  wire w_mem_inst__abc_21378_n5509;
  wire w_mem_inst__abc_21378_n5510;
  wire w_mem_inst__abc_21378_n5511;
  wire w_mem_inst__abc_21378_n5512;
  wire w_mem_inst__abc_21378_n5514;
  wire w_mem_inst__abc_21378_n5515;
  wire w_mem_inst__abc_21378_n5516;
  wire w_mem_inst__abc_21378_n5517;
  wire w_mem_inst__abc_21378_n5518;
  wire w_mem_inst__abc_21378_n5520;
  wire w_mem_inst__abc_21378_n5521;
  wire w_mem_inst__abc_21378_n5522;
  wire w_mem_inst__abc_21378_n5523;
  wire w_mem_inst__abc_21378_n5524;
  wire w_mem_inst__abc_21378_n5526;
  wire w_mem_inst__abc_21378_n5527;
  wire w_mem_inst__abc_21378_n5528;
  wire w_mem_inst__abc_21378_n5529;
  wire w_mem_inst__abc_21378_n5530;
  wire w_mem_inst__abc_21378_n5532;
  wire w_mem_inst__abc_21378_n5533;
  wire w_mem_inst__abc_21378_n5534;
  wire w_mem_inst__abc_21378_n5535;
  wire w_mem_inst__abc_21378_n5536;
  wire w_mem_inst__abc_21378_n5538;
  wire w_mem_inst__abc_21378_n5539;
  wire w_mem_inst__abc_21378_n5540;
  wire w_mem_inst__abc_21378_n5541;
  wire w_mem_inst__abc_21378_n5542;
  wire w_mem_inst__abc_21378_n5544;
  wire w_mem_inst__abc_21378_n5545;
  wire w_mem_inst__abc_21378_n5546;
  wire w_mem_inst__abc_21378_n5547;
  wire w_mem_inst__abc_21378_n5548;
  wire w_mem_inst__abc_21378_n5550;
  wire w_mem_inst__abc_21378_n5551;
  wire w_mem_inst__abc_21378_n5552;
  wire w_mem_inst__abc_21378_n5553;
  wire w_mem_inst__abc_21378_n5554;
  wire w_mem_inst__abc_21378_n5556;
  wire w_mem_inst__abc_21378_n5557;
  wire w_mem_inst__abc_21378_n5558;
  wire w_mem_inst__abc_21378_n5559;
  wire w_mem_inst__abc_21378_n5560;
  wire w_mem_inst__abc_21378_n5562;
  wire w_mem_inst__abc_21378_n5563;
  wire w_mem_inst__abc_21378_n5564;
  wire w_mem_inst__abc_21378_n5565;
  wire w_mem_inst__abc_21378_n5566;
  wire w_mem_inst__abc_21378_n5568;
  wire w_mem_inst__abc_21378_n5569;
  wire w_mem_inst__abc_21378_n5570;
  wire w_mem_inst__abc_21378_n5571;
  wire w_mem_inst__abc_21378_n5572;
  wire w_mem_inst__abc_21378_n5574;
  wire w_mem_inst__abc_21378_n5575;
  wire w_mem_inst__abc_21378_n5576;
  wire w_mem_inst__abc_21378_n5577;
  wire w_mem_inst__abc_21378_n5578;
  wire w_mem_inst__abc_21378_n5580;
  wire w_mem_inst__abc_21378_n5581;
  wire w_mem_inst__abc_21378_n5582;
  wire w_mem_inst__abc_21378_n5583;
  wire w_mem_inst__abc_21378_n5584;
  wire w_mem_inst__abc_21378_n5586;
  wire w_mem_inst__abc_21378_n5587;
  wire w_mem_inst__abc_21378_n5588;
  wire w_mem_inst__abc_21378_n5589;
  wire w_mem_inst__abc_21378_n5590;
  wire w_mem_inst__abc_21378_n5592;
  wire w_mem_inst__abc_21378_n5593;
  wire w_mem_inst__abc_21378_n5594;
  wire w_mem_inst__abc_21378_n5595;
  wire w_mem_inst__abc_21378_n5596;
  wire w_mem_inst__abc_21378_n5598;
  wire w_mem_inst__abc_21378_n5599;
  wire w_mem_inst__abc_21378_n5600;
  wire w_mem_inst__abc_21378_n5601;
  wire w_mem_inst__abc_21378_n5602;
  wire w_mem_inst__abc_21378_n5604;
  wire w_mem_inst__abc_21378_n5605;
  wire w_mem_inst__abc_21378_n5606;
  wire w_mem_inst__abc_21378_n5607;
  wire w_mem_inst__abc_21378_n5608;
  wire w_mem_inst__abc_21378_n5610;
  wire w_mem_inst__abc_21378_n5611;
  wire w_mem_inst__abc_21378_n5612;
  wire w_mem_inst__abc_21378_n5613;
  wire w_mem_inst__abc_21378_n5614;
  wire w_mem_inst__abc_21378_n5616;
  wire w_mem_inst__abc_21378_n5617;
  wire w_mem_inst__abc_21378_n5618;
  wire w_mem_inst__abc_21378_n5619;
  wire w_mem_inst__abc_21378_n5620;
  wire w_mem_inst__abc_21378_n5622;
  wire w_mem_inst__abc_21378_n5623;
  wire w_mem_inst__abc_21378_n5624;
  wire w_mem_inst__abc_21378_n5625;
  wire w_mem_inst__abc_21378_n5626;
  wire w_mem_inst__abc_21378_n5628;
  wire w_mem_inst__abc_21378_n5629;
  wire w_mem_inst__abc_21378_n5630;
  wire w_mem_inst__abc_21378_n5631;
  wire w_mem_inst__abc_21378_n5632;
  wire w_mem_inst__abc_21378_n5634;
  wire w_mem_inst__abc_21378_n5635;
  wire w_mem_inst__abc_21378_n5636;
  wire w_mem_inst__abc_21378_n5637;
  wire w_mem_inst__abc_21378_n5638;
  wire w_mem_inst__abc_21378_n5640;
  wire w_mem_inst__abc_21378_n5641;
  wire w_mem_inst__abc_21378_n5642;
  wire w_mem_inst__abc_21378_n5643;
  wire w_mem_inst__abc_21378_n5644;
  wire w_mem_inst__abc_21378_n5646;
  wire w_mem_inst__abc_21378_n5647;
  wire w_mem_inst__abc_21378_n5648;
  wire w_mem_inst__abc_21378_n5649;
  wire w_mem_inst__abc_21378_n5650;
  wire w_mem_inst__abc_21378_n5652;
  wire w_mem_inst__abc_21378_n5653;
  wire w_mem_inst__abc_21378_n5654;
  wire w_mem_inst__abc_21378_n5655;
  wire w_mem_inst__abc_21378_n5656;
  wire w_mem_inst__abc_21378_n5658;
  wire w_mem_inst__abc_21378_n5659;
  wire w_mem_inst__abc_21378_n5660;
  wire w_mem_inst__abc_21378_n5661;
  wire w_mem_inst__abc_21378_n5662;
  wire w_mem_inst__abc_21378_n5664;
  wire w_mem_inst__abc_21378_n5665;
  wire w_mem_inst__abc_21378_n5666;
  wire w_mem_inst__abc_21378_n5667;
  wire w_mem_inst__abc_21378_n5668;
  wire w_mem_inst__abc_21378_n5670;
  wire w_mem_inst__abc_21378_n5671;
  wire w_mem_inst__abc_21378_n5672;
  wire w_mem_inst__abc_21378_n5673;
  wire w_mem_inst__abc_21378_n5674;
  wire w_mem_inst__abc_21378_n5676;
  wire w_mem_inst__abc_21378_n5677;
  wire w_mem_inst__abc_21378_n5678;
  wire w_mem_inst__abc_21378_n5679;
  wire w_mem_inst__abc_21378_n5680;
  wire w_mem_inst__abc_21378_n5682;
  wire w_mem_inst__abc_21378_n5683;
  wire w_mem_inst__abc_21378_n5684;
  wire w_mem_inst__abc_21378_n5685;
  wire w_mem_inst__abc_21378_n5686;
  wire w_mem_inst__abc_21378_n5688;
  wire w_mem_inst__abc_21378_n5689;
  wire w_mem_inst__abc_21378_n5690;
  wire w_mem_inst__abc_21378_n5691;
  wire w_mem_inst__abc_21378_n5692;
  wire w_mem_inst__abc_21378_n5694;
  wire w_mem_inst__abc_21378_n5695;
  wire w_mem_inst__abc_21378_n5696;
  wire w_mem_inst__abc_21378_n5697;
  wire w_mem_inst__abc_21378_n5698;
  wire w_mem_inst__abc_21378_n5700;
  wire w_mem_inst__abc_21378_n5701;
  wire w_mem_inst__abc_21378_n5702;
  wire w_mem_inst__abc_21378_n5703;
  wire w_mem_inst__abc_21378_n5704;
  wire w_mem_inst__abc_21378_n5706;
  wire w_mem_inst__abc_21378_n5707;
  wire w_mem_inst__abc_21378_n5708;
  wire w_mem_inst__abc_21378_n5709;
  wire w_mem_inst__abc_21378_n5710;
  wire w_mem_inst__abc_21378_n5712;
  wire w_mem_inst__abc_21378_n5713;
  wire w_mem_inst__abc_21378_n5714;
  wire w_mem_inst__abc_21378_n5715;
  wire w_mem_inst__abc_21378_n5716;
  wire w_mem_inst__abc_21378_n5718;
  wire w_mem_inst__abc_21378_n5719;
  wire w_mem_inst__abc_21378_n5720;
  wire w_mem_inst__abc_21378_n5721;
  wire w_mem_inst__abc_21378_n5722;
  wire w_mem_inst__abc_21378_n5724;
  wire w_mem_inst__abc_21378_n5725;
  wire w_mem_inst__abc_21378_n5726;
  wire w_mem_inst__abc_21378_n5727;
  wire w_mem_inst__abc_21378_n5728;
  wire w_mem_inst__abc_21378_n5730;
  wire w_mem_inst__abc_21378_n5731;
  wire w_mem_inst__abc_21378_n5732;
  wire w_mem_inst__abc_21378_n5733;
  wire w_mem_inst__abc_21378_n5734;
  wire w_mem_inst__abc_21378_n5736;
  wire w_mem_inst__abc_21378_n5737;
  wire w_mem_inst__abc_21378_n5738;
  wire w_mem_inst__abc_21378_n5739;
  wire w_mem_inst__abc_21378_n5740;
  wire w_mem_inst__abc_21378_n5742;
  wire w_mem_inst__abc_21378_n5743;
  wire w_mem_inst__abc_21378_n5744;
  wire w_mem_inst__abc_21378_n5745;
  wire w_mem_inst__abc_21378_n5746;
  wire w_mem_inst__abc_21378_n5748;
  wire w_mem_inst__abc_21378_n5749;
  wire w_mem_inst__abc_21378_n5750;
  wire w_mem_inst__abc_21378_n5751;
  wire w_mem_inst__abc_21378_n5752;
  wire w_mem_inst__abc_21378_n5754;
  wire w_mem_inst__abc_21378_n5755;
  wire w_mem_inst__abc_21378_n5756;
  wire w_mem_inst__abc_21378_n5757;
  wire w_mem_inst__abc_21378_n5758;
  wire w_mem_inst__abc_21378_n5760;
  wire w_mem_inst__abc_21378_n5761;
  wire w_mem_inst__abc_21378_n5762;
  wire w_mem_inst__abc_21378_n5763;
  wire w_mem_inst__abc_21378_n5764;
  wire w_mem_inst__abc_21378_n5766;
  wire w_mem_inst__abc_21378_n5767;
  wire w_mem_inst__abc_21378_n5768;
  wire w_mem_inst__abc_21378_n5769;
  wire w_mem_inst__abc_21378_n5770;
  wire w_mem_inst__abc_21378_n5772;
  wire w_mem_inst__abc_21378_n5773;
  wire w_mem_inst__abc_21378_n5774;
  wire w_mem_inst__abc_21378_n5775;
  wire w_mem_inst__abc_21378_n5776;
  wire w_mem_inst__abc_21378_n5778;
  wire w_mem_inst__abc_21378_n5779;
  wire w_mem_inst__abc_21378_n5780;
  wire w_mem_inst__abc_21378_n5781;
  wire w_mem_inst__abc_21378_n5782;
  wire w_mem_inst__abc_21378_n5784;
  wire w_mem_inst__abc_21378_n5785;
  wire w_mem_inst__abc_21378_n5786;
  wire w_mem_inst__abc_21378_n5787;
  wire w_mem_inst__abc_21378_n5788;
  wire w_mem_inst__abc_21378_n5790;
  wire w_mem_inst__abc_21378_n5791;
  wire w_mem_inst__abc_21378_n5792;
  wire w_mem_inst__abc_21378_n5793;
  wire w_mem_inst__abc_21378_n5794;
  wire w_mem_inst__abc_21378_n5796;
  wire w_mem_inst__abc_21378_n5797;
  wire w_mem_inst__abc_21378_n5798;
  wire w_mem_inst__abc_21378_n5799;
  wire w_mem_inst__abc_21378_n5800;
  wire w_mem_inst__abc_21378_n5802;
  wire w_mem_inst__abc_21378_n5803;
  wire w_mem_inst__abc_21378_n5804;
  wire w_mem_inst__abc_21378_n5805;
  wire w_mem_inst__abc_21378_n5806;
  wire w_mem_inst__abc_21378_n5808;
  wire w_mem_inst__abc_21378_n5809;
  wire w_mem_inst__abc_21378_n5810;
  wire w_mem_inst__abc_21378_n5811;
  wire w_mem_inst__abc_21378_n5812;
  wire w_mem_inst__abc_21378_n5814;
  wire w_mem_inst__abc_21378_n5815;
  wire w_mem_inst__abc_21378_n5816;
  wire w_mem_inst__abc_21378_n5817;
  wire w_mem_inst__abc_21378_n5818;
  wire w_mem_inst__abc_21378_n5820;
  wire w_mem_inst__abc_21378_n5821;
  wire w_mem_inst__abc_21378_n5822;
  wire w_mem_inst__abc_21378_n5823;
  wire w_mem_inst__abc_21378_n5824;
  wire w_mem_inst__abc_21378_n5826;
  wire w_mem_inst__abc_21378_n5827;
  wire w_mem_inst__abc_21378_n5828;
  wire w_mem_inst__abc_21378_n5829;
  wire w_mem_inst__abc_21378_n5830;
  wire w_mem_inst__abc_21378_n5832;
  wire w_mem_inst__abc_21378_n5833;
  wire w_mem_inst__abc_21378_n5834;
  wire w_mem_inst__abc_21378_n5835;
  wire w_mem_inst__abc_21378_n5836;
  wire w_mem_inst__abc_21378_n5838;
  wire w_mem_inst__abc_21378_n5839;
  wire w_mem_inst__abc_21378_n5840;
  wire w_mem_inst__abc_21378_n5841;
  wire w_mem_inst__abc_21378_n5842;
  wire w_mem_inst__abc_21378_n5844;
  wire w_mem_inst__abc_21378_n5845;
  wire w_mem_inst__abc_21378_n5846;
  wire w_mem_inst__abc_21378_n5847;
  wire w_mem_inst__abc_21378_n5848;
  wire w_mem_inst__abc_21378_n5850;
  wire w_mem_inst__abc_21378_n5851;
  wire w_mem_inst__abc_21378_n5852;
  wire w_mem_inst__abc_21378_n5853;
  wire w_mem_inst__abc_21378_n5854;
  wire w_mem_inst__abc_21378_n5856;
  wire w_mem_inst__abc_21378_n5857;
  wire w_mem_inst__abc_21378_n5858;
  wire w_mem_inst__abc_21378_n5859;
  wire w_mem_inst__abc_21378_n5860;
  wire w_mem_inst__abc_21378_n5862;
  wire w_mem_inst__abc_21378_n5863;
  wire w_mem_inst__abc_21378_n5864;
  wire w_mem_inst__abc_21378_n5865;
  wire w_mem_inst__abc_21378_n5866;
  wire w_mem_inst__abc_21378_n5868;
  wire w_mem_inst__abc_21378_n5869;
  wire w_mem_inst__abc_21378_n5870;
  wire w_mem_inst__abc_21378_n5871;
  wire w_mem_inst__abc_21378_n5872;
  wire w_mem_inst__abc_21378_n5874;
  wire w_mem_inst__abc_21378_n5875;
  wire w_mem_inst__abc_21378_n5876;
  wire w_mem_inst__abc_21378_n5877;
  wire w_mem_inst__abc_21378_n5878;
  wire w_mem_inst__abc_21378_n5880;
  wire w_mem_inst__abc_21378_n5881;
  wire w_mem_inst__abc_21378_n5882;
  wire w_mem_inst__abc_21378_n5883;
  wire w_mem_inst__abc_21378_n5884;
  wire w_mem_inst__abc_21378_n5886;
  wire w_mem_inst__abc_21378_n5887;
  wire w_mem_inst__abc_21378_n5888;
  wire w_mem_inst__abc_21378_n5889;
  wire w_mem_inst__abc_21378_n5890;
  wire w_mem_inst__abc_21378_n5892;
  wire w_mem_inst__abc_21378_n5893;
  wire w_mem_inst__abc_21378_n5894;
  wire w_mem_inst__abc_21378_n5895;
  wire w_mem_inst__abc_21378_n5896;
  wire w_mem_inst__abc_21378_n5898;
  wire w_mem_inst__abc_21378_n5899;
  wire w_mem_inst__abc_21378_n5900;
  wire w_mem_inst__abc_21378_n5901;
  wire w_mem_inst__abc_21378_n5902;
  wire w_mem_inst__abc_21378_n5904;
  wire w_mem_inst__abc_21378_n5905;
  wire w_mem_inst__abc_21378_n5906;
  wire w_mem_inst__abc_21378_n5907;
  wire w_mem_inst__abc_21378_n5908;
  wire w_mem_inst__abc_21378_n5910;
  wire w_mem_inst__abc_21378_n5911;
  wire w_mem_inst__abc_21378_n5912;
  wire w_mem_inst__abc_21378_n5913;
  wire w_mem_inst__abc_21378_n5914;
  wire w_mem_inst__abc_21378_n5916;
  wire w_mem_inst__abc_21378_n5917;
  wire w_mem_inst__abc_21378_n5918;
  wire w_mem_inst__abc_21378_n5919;
  wire w_mem_inst__abc_21378_n5920;
  wire w_mem_inst__abc_21378_n5922;
  wire w_mem_inst__abc_21378_n5923;
  wire w_mem_inst__abc_21378_n5924;
  wire w_mem_inst__abc_21378_n5925;
  wire w_mem_inst__abc_21378_n5926;
  wire w_mem_inst__abc_21378_n5928;
  wire w_mem_inst__abc_21378_n5929;
  wire w_mem_inst__abc_21378_n5930;
  wire w_mem_inst__abc_21378_n5931;
  wire w_mem_inst__abc_21378_n5932;
  wire w_mem_inst__abc_21378_n5934;
  wire w_mem_inst__abc_21378_n5935;
  wire w_mem_inst__abc_21378_n5936;
  wire w_mem_inst__abc_21378_n5937;
  wire w_mem_inst__abc_21378_n5938;
  wire w_mem_inst__abc_21378_n5940;
  wire w_mem_inst__abc_21378_n5941;
  wire w_mem_inst__abc_21378_n5942;
  wire w_mem_inst__abc_21378_n5943;
  wire w_mem_inst__abc_21378_n5944;
  wire w_mem_inst__abc_21378_n5946;
  wire w_mem_inst__abc_21378_n5947;
  wire w_mem_inst__abc_21378_n5948;
  wire w_mem_inst__abc_21378_n5949;
  wire w_mem_inst__abc_21378_n5950;
  wire w_mem_inst__abc_21378_n5952;
  wire w_mem_inst__abc_21378_n5953;
  wire w_mem_inst__abc_21378_n5954;
  wire w_mem_inst__abc_21378_n5955;
  wire w_mem_inst__abc_21378_n5956;
  wire w_mem_inst__abc_21378_n5958;
  wire w_mem_inst__abc_21378_n5959;
  wire w_mem_inst__abc_21378_n5960;
  wire w_mem_inst__abc_21378_n5961;
  wire w_mem_inst__abc_21378_n5962;
  wire w_mem_inst__abc_21378_n5964;
  wire w_mem_inst__abc_21378_n5965;
  wire w_mem_inst__abc_21378_n5966;
  wire w_mem_inst__abc_21378_n5967;
  wire w_mem_inst__abc_21378_n5968;
  wire w_mem_inst__abc_21378_n5970;
  wire w_mem_inst__abc_21378_n5971;
  wire w_mem_inst__abc_21378_n5972;
  wire w_mem_inst__abc_21378_n5973;
  wire w_mem_inst__abc_21378_n5974;
  wire w_mem_inst__abc_21378_n5976;
  wire w_mem_inst__abc_21378_n5977;
  wire w_mem_inst__abc_21378_n5978;
  wire w_mem_inst__abc_21378_n5979;
  wire w_mem_inst__abc_21378_n5980;
  wire w_mem_inst__abc_21378_n5982;
  wire w_mem_inst__abc_21378_n5983;
  wire w_mem_inst__abc_21378_n5984;
  wire w_mem_inst__abc_21378_n5985;
  wire w_mem_inst__abc_21378_n5986;
  wire w_mem_inst__abc_21378_n5988;
  wire w_mem_inst__abc_21378_n5989;
  wire w_mem_inst__abc_21378_n5990;
  wire w_mem_inst__abc_21378_n5991;
  wire w_mem_inst__abc_21378_n5992;
  wire w_mem_inst__abc_21378_n5994;
  wire w_mem_inst__abc_21378_n5995;
  wire w_mem_inst__abc_21378_n5996;
  wire w_mem_inst__abc_21378_n5997;
  wire w_mem_inst__abc_21378_n5998;
  wire w_mem_inst__abc_21378_n6000;
  wire w_mem_inst__abc_21378_n6001;
  wire w_mem_inst__abc_21378_n6002;
  wire w_mem_inst__abc_21378_n6003;
  wire w_mem_inst__abc_21378_n6004;
  wire w_mem_inst__abc_21378_n6006;
  wire w_mem_inst__abc_21378_n6007;
  wire w_mem_inst__abc_21378_n6008;
  wire w_mem_inst__abc_21378_n6009;
  wire w_mem_inst__abc_21378_n6010;
  wire w_mem_inst__abc_21378_n6012;
  wire w_mem_inst__abc_21378_n6013;
  wire w_mem_inst__abc_21378_n6014;
  wire w_mem_inst__abc_21378_n6015;
  wire w_mem_inst__abc_21378_n6016;
  wire w_mem_inst__abc_21378_n6018;
  wire w_mem_inst__abc_21378_n6019;
  wire w_mem_inst__abc_21378_n6020;
  wire w_mem_inst__abc_21378_n6021;
  wire w_mem_inst__abc_21378_n6022;
  wire w_mem_inst__abc_21378_n6024;
  wire w_mem_inst__abc_21378_n6025;
  wire w_mem_inst__abc_21378_n6026;
  wire w_mem_inst__abc_21378_n6027;
  wire w_mem_inst__abc_21378_n6028;
  wire w_mem_inst__abc_21378_n6030;
  wire w_mem_inst__abc_21378_n6031;
  wire w_mem_inst__abc_21378_n6032;
  wire w_mem_inst__abc_21378_n6033;
  wire w_mem_inst__abc_21378_n6034;
  wire w_mem_inst__abc_21378_n6036;
  wire w_mem_inst__abc_21378_n6037;
  wire w_mem_inst__abc_21378_n6038;
  wire w_mem_inst__abc_21378_n6039;
  wire w_mem_inst__abc_21378_n6040;
  wire w_mem_inst__abc_21378_n6042;
  wire w_mem_inst__abc_21378_n6043;
  wire w_mem_inst__abc_21378_n6044;
  wire w_mem_inst__abc_21378_n6045;
  wire w_mem_inst__abc_21378_n6046;
  wire w_mem_inst__abc_21378_n6048;
  wire w_mem_inst__abc_21378_n6049;
  wire w_mem_inst__abc_21378_n6050;
  wire w_mem_inst__abc_21378_n6051;
  wire w_mem_inst__abc_21378_n6052;
  wire w_mem_inst__abc_21378_n6054;
  wire w_mem_inst__abc_21378_n6055;
  wire w_mem_inst__abc_21378_n6056;
  wire w_mem_inst__abc_21378_n6057;
  wire w_mem_inst__abc_21378_n6058;
  wire w_mem_inst__abc_21378_n6060;
  wire w_mem_inst__abc_21378_n6061;
  wire w_mem_inst__abc_21378_n6062;
  wire w_mem_inst__abc_21378_n6063;
  wire w_mem_inst__abc_21378_n6064;
  wire w_mem_inst__abc_21378_n6066;
  wire w_mem_inst__abc_21378_n6067;
  wire w_mem_inst__abc_21378_n6068;
  wire w_mem_inst__abc_21378_n6069;
  wire w_mem_inst__abc_21378_n6070;
  wire w_mem_inst__abc_21378_n6072;
  wire w_mem_inst__abc_21378_n6073;
  wire w_mem_inst__abc_21378_n6074;
  wire w_mem_inst__abc_21378_n6075;
  wire w_mem_inst__abc_21378_n6076;
  wire w_mem_inst__abc_21378_n6078;
  wire w_mem_inst__abc_21378_n6079;
  wire w_mem_inst__abc_21378_n6080;
  wire w_mem_inst__abc_21378_n6081;
  wire w_mem_inst__abc_21378_n6082;
  wire w_mem_inst__abc_21378_n6084;
  wire w_mem_inst__abc_21378_n6085;
  wire w_mem_inst__abc_21378_n6086;
  wire w_mem_inst__abc_21378_n6087;
  wire w_mem_inst__abc_21378_n6088;
  wire w_mem_inst__abc_21378_n6090;
  wire w_mem_inst__abc_21378_n6091;
  wire w_mem_inst__abc_21378_n6092;
  wire w_mem_inst__abc_21378_n6093;
  wire w_mem_inst__abc_21378_n6094;
  wire w_mem_inst__abc_21378_n6096;
  wire w_mem_inst__abc_21378_n6097;
  wire w_mem_inst__abc_21378_n6098;
  wire w_mem_inst__abc_21378_n6099;
  wire w_mem_inst__abc_21378_n6100;
  wire w_mem_inst__abc_21378_n6102;
  wire w_mem_inst__abc_21378_n6103;
  wire w_mem_inst__abc_21378_n6104;
  wire w_mem_inst__abc_21378_n6105;
  wire w_mem_inst__abc_21378_n6106;
  wire w_mem_inst__abc_21378_n6108;
  wire w_mem_inst__abc_21378_n6109;
  wire w_mem_inst__abc_21378_n6110;
  wire w_mem_inst__abc_21378_n6111;
  wire w_mem_inst__abc_21378_n6112;
  wire w_mem_inst__abc_21378_n6114;
  wire w_mem_inst__abc_21378_n6115;
  wire w_mem_inst__abc_21378_n6116;
  wire w_mem_inst__abc_21378_n6117;
  wire w_mem_inst__abc_21378_n6118;
  wire w_mem_inst__abc_21378_n6120;
  wire w_mem_inst__abc_21378_n6121;
  wire w_mem_inst__abc_21378_n6122;
  wire w_mem_inst__abc_21378_n6123;
  wire w_mem_inst__abc_21378_n6124;
  wire w_mem_inst__abc_21378_n6126;
  wire w_mem_inst__abc_21378_n6127;
  wire w_mem_inst__abc_21378_n6128;
  wire w_mem_inst__abc_21378_n6129;
  wire w_mem_inst__abc_21378_n6130;
  wire w_mem_inst__abc_21378_n6132;
  wire w_mem_inst__abc_21378_n6133;
  wire w_mem_inst__abc_21378_n6134;
  wire w_mem_inst__abc_21378_n6135;
  wire w_mem_inst__abc_21378_n6136;
  wire w_mem_inst__abc_21378_n6138;
  wire w_mem_inst__abc_21378_n6139;
  wire w_mem_inst__abc_21378_n6140;
  wire w_mem_inst__abc_21378_n6141;
  wire w_mem_inst__abc_21378_n6142;
  wire w_mem_inst__abc_21378_n6144;
  wire w_mem_inst__abc_21378_n6145;
  wire w_mem_inst__abc_21378_n6146;
  wire w_mem_inst__abc_21378_n6147;
  wire w_mem_inst__abc_21378_n6148;
  wire w_mem_inst__abc_21378_n6150;
  wire w_mem_inst__abc_21378_n6151;
  wire w_mem_inst__abc_21378_n6152;
  wire w_mem_inst__abc_21378_n6153;
  wire w_mem_inst__abc_21378_n6154;
  wire w_mem_inst__abc_21378_n6156;
  wire w_mem_inst__abc_21378_n6157;
  wire w_mem_inst__abc_21378_n6158;
  wire w_mem_inst__abc_21378_n6159;
  wire w_mem_inst__abc_21378_n6160;
  wire w_mem_inst__abc_21378_n6162;
  wire w_mem_inst__abc_21378_n6163;
  wire w_mem_inst__abc_21378_n6164;
  wire w_mem_inst__abc_21378_n6165;
  wire w_mem_inst__abc_21378_n6166;
  wire w_mem_inst__abc_21378_n6168;
  wire w_mem_inst__abc_21378_n6169;
  wire w_mem_inst__abc_21378_n6170;
  wire w_mem_inst__abc_21378_n6171;
  wire w_mem_inst__abc_21378_n6172;
  wire w_mem_inst__abc_21378_n6174;
  wire w_mem_inst__abc_21378_n6175;
  wire w_mem_inst__abc_21378_n6176;
  wire w_mem_inst__abc_21378_n6177;
  wire w_mem_inst__abc_21378_n6178;
  wire w_mem_inst__abc_21378_n6180;
  wire w_mem_inst__abc_21378_n6181;
  wire w_mem_inst__abc_21378_n6182;
  wire w_mem_inst__abc_21378_n6183;
  wire w_mem_inst__abc_21378_n6184;
  wire w_mem_inst__abc_21378_n6186;
  wire w_mem_inst__abc_21378_n6187;
  wire w_mem_inst__abc_21378_n6188;
  wire w_mem_inst__abc_21378_n6189;
  wire w_mem_inst__abc_21378_n6190;
  wire w_mem_inst__abc_21378_n6192;
  wire w_mem_inst__abc_21378_n6193;
  wire w_mem_inst__abc_21378_n6194;
  wire w_mem_inst__abc_21378_n6195;
  wire w_mem_inst__abc_21378_n6196;
  wire w_mem_inst__abc_21378_n6198;
  wire w_mem_inst__abc_21378_n6199;
  wire w_mem_inst__abc_21378_n6200;
  wire w_mem_inst__abc_21378_n6201;
  wire w_mem_inst__abc_21378_n6202;
  wire w_mem_inst__abc_21378_n6204;
  wire w_mem_inst__abc_21378_n6205;
  wire w_mem_inst__abc_21378_n6206;
  wire w_mem_inst__abc_21378_n6207;
  wire w_mem_inst__abc_21378_n6208;
  wire w_mem_inst__abc_21378_n6210;
  wire w_mem_inst__abc_21378_n6211;
  wire w_mem_inst__abc_21378_n6212;
  wire w_mem_inst__abc_21378_n6213;
  wire w_mem_inst__abc_21378_n6214;
  wire w_mem_inst__abc_21378_n6216;
  wire w_mem_inst__abc_21378_n6217;
  wire w_mem_inst__abc_21378_n6218;
  wire w_mem_inst__abc_21378_n6219;
  wire w_mem_inst__abc_21378_n6220;
  wire w_mem_inst__abc_21378_n6222;
  wire w_mem_inst__abc_21378_n6223;
  wire w_mem_inst__abc_21378_n6224;
  wire w_mem_inst__abc_21378_n6225;
  wire w_mem_inst__abc_21378_n6226;
  wire w_mem_inst__abc_21378_n6228;
  wire w_mem_inst__abc_21378_n6229;
  wire w_mem_inst__abc_21378_n6230;
  wire w_mem_inst__abc_21378_n6231;
  wire w_mem_inst__abc_21378_n6233;
  wire w_mem_inst__abc_21378_n6234;
  wire w_mem_inst__abc_21378_n6235;
  wire w_mem_inst__abc_21378_n6237;
  wire w_mem_inst__abc_21378_n6238;
  wire w_mem_inst__abc_21378_n6239;
  wire w_mem_inst__abc_21378_n6240;
  wire w_mem_inst__abc_21378_n6241;
  wire w_mem_inst__abc_21378_n6242;
  wire w_mem_inst__abc_21378_n6243;
  wire w_mem_inst__abc_21378_n6245;
  wire w_mem_inst__abc_21378_n6246;
  wire w_mem_inst__abc_21378_n6247;
  wire w_mem_inst__abc_21378_n6248;
  wire w_mem_inst__abc_21378_n6250;
  wire w_mem_inst__abc_21378_n6251;
  wire w_mem_inst__abc_21378_n6252;
  wire w_mem_inst__abc_21378_n6253;
  wire w_mem_inst__abc_21378_n6255;
  wire w_mem_inst__abc_21378_n6256;
  wire w_mem_inst__abc_21378_n6257;
  wire w_mem_inst__abc_21378_n6258;
  wire w_mem_inst__abc_21378_n6260;
  wire w_mem_inst__abc_21378_n6261;
  wire w_mem_inst__abc_21378_n6262;
  wire w_mem_inst__abc_21378_n6263;
  wire w_mem_inst_w_ctr_reg_0_;
  wire w_mem_inst_w_ctr_reg_0__FF_INPUT;
  wire w_mem_inst_w_ctr_reg_1_;
  wire w_mem_inst_w_ctr_reg_1__FF_INPUT;
  wire w_mem_inst_w_ctr_reg_2_;
  wire w_mem_inst_w_ctr_reg_2__FF_INPUT;
  wire w_mem_inst_w_ctr_reg_3_;
  wire w_mem_inst_w_ctr_reg_3__FF_INPUT;
  wire w_mem_inst_w_ctr_reg_4_;
  wire w_mem_inst_w_ctr_reg_4__FF_INPUT;
  wire w_mem_inst_w_ctr_reg_5_;
  wire w_mem_inst_w_ctr_reg_5__FF_INPUT;
  wire w_mem_inst_w_ctr_reg_6_;
  wire w_mem_inst_w_ctr_reg_6__FF_INPUT;
  wire w_mem_inst_w_mem_0__0_;
  wire w_mem_inst_w_mem_0__10_;
  wire w_mem_inst_w_mem_0__11_;
  wire w_mem_inst_w_mem_0__12_;
  wire w_mem_inst_w_mem_0__13_;
  wire w_mem_inst_w_mem_0__14_;
  wire w_mem_inst_w_mem_0__15_;
  wire w_mem_inst_w_mem_0__16_;
  wire w_mem_inst_w_mem_0__17_;
  wire w_mem_inst_w_mem_0__18_;
  wire w_mem_inst_w_mem_0__19_;
  wire w_mem_inst_w_mem_0__1_;
  wire w_mem_inst_w_mem_0__20_;
  wire w_mem_inst_w_mem_0__21_;
  wire w_mem_inst_w_mem_0__22_;
  wire w_mem_inst_w_mem_0__23_;
  wire w_mem_inst_w_mem_0__24_;
  wire w_mem_inst_w_mem_0__25_;
  wire w_mem_inst_w_mem_0__26_;
  wire w_mem_inst_w_mem_0__27_;
  wire w_mem_inst_w_mem_0__28_;
  wire w_mem_inst_w_mem_0__29_;
  wire w_mem_inst_w_mem_0__2_;
  wire w_mem_inst_w_mem_0__30_;
  wire w_mem_inst_w_mem_0__31_;
  wire w_mem_inst_w_mem_0__3_;
  wire w_mem_inst_w_mem_0__4_;
  wire w_mem_inst_w_mem_0__5_;
  wire w_mem_inst_w_mem_0__6_;
  wire w_mem_inst_w_mem_0__7_;
  wire w_mem_inst_w_mem_0__8_;
  wire w_mem_inst_w_mem_0__9_;
  wire w_mem_inst_w_mem_10__0_;
  wire w_mem_inst_w_mem_10__10_;
  wire w_mem_inst_w_mem_10__11_;
  wire w_mem_inst_w_mem_10__12_;
  wire w_mem_inst_w_mem_10__13_;
  wire w_mem_inst_w_mem_10__14_;
  wire w_mem_inst_w_mem_10__15_;
  wire w_mem_inst_w_mem_10__16_;
  wire w_mem_inst_w_mem_10__17_;
  wire w_mem_inst_w_mem_10__18_;
  wire w_mem_inst_w_mem_10__19_;
  wire w_mem_inst_w_mem_10__1_;
  wire w_mem_inst_w_mem_10__20_;
  wire w_mem_inst_w_mem_10__21_;
  wire w_mem_inst_w_mem_10__22_;
  wire w_mem_inst_w_mem_10__23_;
  wire w_mem_inst_w_mem_10__24_;
  wire w_mem_inst_w_mem_10__25_;
  wire w_mem_inst_w_mem_10__26_;
  wire w_mem_inst_w_mem_10__27_;
  wire w_mem_inst_w_mem_10__28_;
  wire w_mem_inst_w_mem_10__29_;
  wire w_mem_inst_w_mem_10__2_;
  wire w_mem_inst_w_mem_10__30_;
  wire w_mem_inst_w_mem_10__31_;
  wire w_mem_inst_w_mem_10__3_;
  wire w_mem_inst_w_mem_10__4_;
  wire w_mem_inst_w_mem_10__5_;
  wire w_mem_inst_w_mem_10__6_;
  wire w_mem_inst_w_mem_10__7_;
  wire w_mem_inst_w_mem_10__8_;
  wire w_mem_inst_w_mem_10__9_;
  wire w_mem_inst_w_mem_11__0_;
  wire w_mem_inst_w_mem_11__10_;
  wire w_mem_inst_w_mem_11__11_;
  wire w_mem_inst_w_mem_11__12_;
  wire w_mem_inst_w_mem_11__13_;
  wire w_mem_inst_w_mem_11__14_;
  wire w_mem_inst_w_mem_11__15_;
  wire w_mem_inst_w_mem_11__16_;
  wire w_mem_inst_w_mem_11__17_;
  wire w_mem_inst_w_mem_11__18_;
  wire w_mem_inst_w_mem_11__19_;
  wire w_mem_inst_w_mem_11__1_;
  wire w_mem_inst_w_mem_11__20_;
  wire w_mem_inst_w_mem_11__21_;
  wire w_mem_inst_w_mem_11__22_;
  wire w_mem_inst_w_mem_11__23_;
  wire w_mem_inst_w_mem_11__24_;
  wire w_mem_inst_w_mem_11__25_;
  wire w_mem_inst_w_mem_11__26_;
  wire w_mem_inst_w_mem_11__27_;
  wire w_mem_inst_w_mem_11__28_;
  wire w_mem_inst_w_mem_11__29_;
  wire w_mem_inst_w_mem_11__2_;
  wire w_mem_inst_w_mem_11__30_;
  wire w_mem_inst_w_mem_11__31_;
  wire w_mem_inst_w_mem_11__3_;
  wire w_mem_inst_w_mem_11__4_;
  wire w_mem_inst_w_mem_11__5_;
  wire w_mem_inst_w_mem_11__6_;
  wire w_mem_inst_w_mem_11__7_;
  wire w_mem_inst_w_mem_11__8_;
  wire w_mem_inst_w_mem_11__9_;
  wire w_mem_inst_w_mem_12__0_;
  wire w_mem_inst_w_mem_12__10_;
  wire w_mem_inst_w_mem_12__11_;
  wire w_mem_inst_w_mem_12__12_;
  wire w_mem_inst_w_mem_12__13_;
  wire w_mem_inst_w_mem_12__14_;
  wire w_mem_inst_w_mem_12__15_;
  wire w_mem_inst_w_mem_12__16_;
  wire w_mem_inst_w_mem_12__17_;
  wire w_mem_inst_w_mem_12__18_;
  wire w_mem_inst_w_mem_12__19_;
  wire w_mem_inst_w_mem_12__1_;
  wire w_mem_inst_w_mem_12__20_;
  wire w_mem_inst_w_mem_12__21_;
  wire w_mem_inst_w_mem_12__22_;
  wire w_mem_inst_w_mem_12__23_;
  wire w_mem_inst_w_mem_12__24_;
  wire w_mem_inst_w_mem_12__25_;
  wire w_mem_inst_w_mem_12__26_;
  wire w_mem_inst_w_mem_12__27_;
  wire w_mem_inst_w_mem_12__28_;
  wire w_mem_inst_w_mem_12__29_;
  wire w_mem_inst_w_mem_12__2_;
  wire w_mem_inst_w_mem_12__30_;
  wire w_mem_inst_w_mem_12__31_;
  wire w_mem_inst_w_mem_12__3_;
  wire w_mem_inst_w_mem_12__4_;
  wire w_mem_inst_w_mem_12__5_;
  wire w_mem_inst_w_mem_12__6_;
  wire w_mem_inst_w_mem_12__7_;
  wire w_mem_inst_w_mem_12__8_;
  wire w_mem_inst_w_mem_12__9_;
  wire w_mem_inst_w_mem_13__0_;
  wire w_mem_inst_w_mem_13__10_;
  wire w_mem_inst_w_mem_13__11_;
  wire w_mem_inst_w_mem_13__12_;
  wire w_mem_inst_w_mem_13__13_;
  wire w_mem_inst_w_mem_13__14_;
  wire w_mem_inst_w_mem_13__15_;
  wire w_mem_inst_w_mem_13__16_;
  wire w_mem_inst_w_mem_13__17_;
  wire w_mem_inst_w_mem_13__18_;
  wire w_mem_inst_w_mem_13__19_;
  wire w_mem_inst_w_mem_13__1_;
  wire w_mem_inst_w_mem_13__20_;
  wire w_mem_inst_w_mem_13__21_;
  wire w_mem_inst_w_mem_13__22_;
  wire w_mem_inst_w_mem_13__23_;
  wire w_mem_inst_w_mem_13__24_;
  wire w_mem_inst_w_mem_13__25_;
  wire w_mem_inst_w_mem_13__26_;
  wire w_mem_inst_w_mem_13__27_;
  wire w_mem_inst_w_mem_13__28_;
  wire w_mem_inst_w_mem_13__29_;
  wire w_mem_inst_w_mem_13__2_;
  wire w_mem_inst_w_mem_13__30_;
  wire w_mem_inst_w_mem_13__31_;
  wire w_mem_inst_w_mem_13__3_;
  wire w_mem_inst_w_mem_13__4_;
  wire w_mem_inst_w_mem_13__5_;
  wire w_mem_inst_w_mem_13__6_;
  wire w_mem_inst_w_mem_13__7_;
  wire w_mem_inst_w_mem_13__8_;
  wire w_mem_inst_w_mem_13__9_;
  wire w_mem_inst_w_mem_14__0_;
  wire w_mem_inst_w_mem_14__10_;
  wire w_mem_inst_w_mem_14__11_;
  wire w_mem_inst_w_mem_14__12_;
  wire w_mem_inst_w_mem_14__13_;
  wire w_mem_inst_w_mem_14__14_;
  wire w_mem_inst_w_mem_14__15_;
  wire w_mem_inst_w_mem_14__16_;
  wire w_mem_inst_w_mem_14__17_;
  wire w_mem_inst_w_mem_14__18_;
  wire w_mem_inst_w_mem_14__19_;
  wire w_mem_inst_w_mem_14__1_;
  wire w_mem_inst_w_mem_14__20_;
  wire w_mem_inst_w_mem_14__21_;
  wire w_mem_inst_w_mem_14__22_;
  wire w_mem_inst_w_mem_14__23_;
  wire w_mem_inst_w_mem_14__24_;
  wire w_mem_inst_w_mem_14__25_;
  wire w_mem_inst_w_mem_14__26_;
  wire w_mem_inst_w_mem_14__27_;
  wire w_mem_inst_w_mem_14__28_;
  wire w_mem_inst_w_mem_14__29_;
  wire w_mem_inst_w_mem_14__2_;
  wire w_mem_inst_w_mem_14__30_;
  wire w_mem_inst_w_mem_14__31_;
  wire w_mem_inst_w_mem_14__3_;
  wire w_mem_inst_w_mem_14__4_;
  wire w_mem_inst_w_mem_14__5_;
  wire w_mem_inst_w_mem_14__6_;
  wire w_mem_inst_w_mem_14__7_;
  wire w_mem_inst_w_mem_14__8_;
  wire w_mem_inst_w_mem_14__9_;
  wire w_mem_inst_w_mem_15__0_;
  wire w_mem_inst_w_mem_15__10_;
  wire w_mem_inst_w_mem_15__11_;
  wire w_mem_inst_w_mem_15__12_;
  wire w_mem_inst_w_mem_15__13_;
  wire w_mem_inst_w_mem_15__14_;
  wire w_mem_inst_w_mem_15__15_;
  wire w_mem_inst_w_mem_15__16_;
  wire w_mem_inst_w_mem_15__17_;
  wire w_mem_inst_w_mem_15__18_;
  wire w_mem_inst_w_mem_15__19_;
  wire w_mem_inst_w_mem_15__1_;
  wire w_mem_inst_w_mem_15__20_;
  wire w_mem_inst_w_mem_15__21_;
  wire w_mem_inst_w_mem_15__22_;
  wire w_mem_inst_w_mem_15__23_;
  wire w_mem_inst_w_mem_15__24_;
  wire w_mem_inst_w_mem_15__25_;
  wire w_mem_inst_w_mem_15__26_;
  wire w_mem_inst_w_mem_15__27_;
  wire w_mem_inst_w_mem_15__28_;
  wire w_mem_inst_w_mem_15__29_;
  wire w_mem_inst_w_mem_15__2_;
  wire w_mem_inst_w_mem_15__30_;
  wire w_mem_inst_w_mem_15__31_;
  wire w_mem_inst_w_mem_15__3_;
  wire w_mem_inst_w_mem_15__4_;
  wire w_mem_inst_w_mem_15__5_;
  wire w_mem_inst_w_mem_15__6_;
  wire w_mem_inst_w_mem_15__7_;
  wire w_mem_inst_w_mem_15__8_;
  wire w_mem_inst_w_mem_15__9_;
  wire w_mem_inst_w_mem_1__0_;
  wire w_mem_inst_w_mem_1__10_;
  wire w_mem_inst_w_mem_1__11_;
  wire w_mem_inst_w_mem_1__12_;
  wire w_mem_inst_w_mem_1__13_;
  wire w_mem_inst_w_mem_1__14_;
  wire w_mem_inst_w_mem_1__15_;
  wire w_mem_inst_w_mem_1__16_;
  wire w_mem_inst_w_mem_1__17_;
  wire w_mem_inst_w_mem_1__18_;
  wire w_mem_inst_w_mem_1__19_;
  wire w_mem_inst_w_mem_1__1_;
  wire w_mem_inst_w_mem_1__20_;
  wire w_mem_inst_w_mem_1__21_;
  wire w_mem_inst_w_mem_1__22_;
  wire w_mem_inst_w_mem_1__23_;
  wire w_mem_inst_w_mem_1__24_;
  wire w_mem_inst_w_mem_1__25_;
  wire w_mem_inst_w_mem_1__26_;
  wire w_mem_inst_w_mem_1__27_;
  wire w_mem_inst_w_mem_1__28_;
  wire w_mem_inst_w_mem_1__29_;
  wire w_mem_inst_w_mem_1__2_;
  wire w_mem_inst_w_mem_1__30_;
  wire w_mem_inst_w_mem_1__31_;
  wire w_mem_inst_w_mem_1__3_;
  wire w_mem_inst_w_mem_1__4_;
  wire w_mem_inst_w_mem_1__5_;
  wire w_mem_inst_w_mem_1__6_;
  wire w_mem_inst_w_mem_1__7_;
  wire w_mem_inst_w_mem_1__8_;
  wire w_mem_inst_w_mem_1__9_;
  wire w_mem_inst_w_mem_2__0_;
  wire w_mem_inst_w_mem_2__10_;
  wire w_mem_inst_w_mem_2__11_;
  wire w_mem_inst_w_mem_2__12_;
  wire w_mem_inst_w_mem_2__13_;
  wire w_mem_inst_w_mem_2__14_;
  wire w_mem_inst_w_mem_2__15_;
  wire w_mem_inst_w_mem_2__16_;
  wire w_mem_inst_w_mem_2__17_;
  wire w_mem_inst_w_mem_2__18_;
  wire w_mem_inst_w_mem_2__19_;
  wire w_mem_inst_w_mem_2__1_;
  wire w_mem_inst_w_mem_2__20_;
  wire w_mem_inst_w_mem_2__21_;
  wire w_mem_inst_w_mem_2__22_;
  wire w_mem_inst_w_mem_2__23_;
  wire w_mem_inst_w_mem_2__24_;
  wire w_mem_inst_w_mem_2__25_;
  wire w_mem_inst_w_mem_2__26_;
  wire w_mem_inst_w_mem_2__27_;
  wire w_mem_inst_w_mem_2__28_;
  wire w_mem_inst_w_mem_2__29_;
  wire w_mem_inst_w_mem_2__2_;
  wire w_mem_inst_w_mem_2__30_;
  wire w_mem_inst_w_mem_2__31_;
  wire w_mem_inst_w_mem_2__3_;
  wire w_mem_inst_w_mem_2__4_;
  wire w_mem_inst_w_mem_2__5_;
  wire w_mem_inst_w_mem_2__6_;
  wire w_mem_inst_w_mem_2__7_;
  wire w_mem_inst_w_mem_2__8_;
  wire w_mem_inst_w_mem_2__9_;
  wire w_mem_inst_w_mem_3__0_;
  wire w_mem_inst_w_mem_3__10_;
  wire w_mem_inst_w_mem_3__11_;
  wire w_mem_inst_w_mem_3__12_;
  wire w_mem_inst_w_mem_3__13_;
  wire w_mem_inst_w_mem_3__14_;
  wire w_mem_inst_w_mem_3__15_;
  wire w_mem_inst_w_mem_3__16_;
  wire w_mem_inst_w_mem_3__17_;
  wire w_mem_inst_w_mem_3__18_;
  wire w_mem_inst_w_mem_3__19_;
  wire w_mem_inst_w_mem_3__1_;
  wire w_mem_inst_w_mem_3__20_;
  wire w_mem_inst_w_mem_3__21_;
  wire w_mem_inst_w_mem_3__22_;
  wire w_mem_inst_w_mem_3__23_;
  wire w_mem_inst_w_mem_3__24_;
  wire w_mem_inst_w_mem_3__25_;
  wire w_mem_inst_w_mem_3__26_;
  wire w_mem_inst_w_mem_3__27_;
  wire w_mem_inst_w_mem_3__28_;
  wire w_mem_inst_w_mem_3__29_;
  wire w_mem_inst_w_mem_3__2_;
  wire w_mem_inst_w_mem_3__30_;
  wire w_mem_inst_w_mem_3__31_;
  wire w_mem_inst_w_mem_3__3_;
  wire w_mem_inst_w_mem_3__4_;
  wire w_mem_inst_w_mem_3__5_;
  wire w_mem_inst_w_mem_3__6_;
  wire w_mem_inst_w_mem_3__7_;
  wire w_mem_inst_w_mem_3__8_;
  wire w_mem_inst_w_mem_3__9_;
  wire w_mem_inst_w_mem_4__0_;
  wire w_mem_inst_w_mem_4__10_;
  wire w_mem_inst_w_mem_4__11_;
  wire w_mem_inst_w_mem_4__12_;
  wire w_mem_inst_w_mem_4__13_;
  wire w_mem_inst_w_mem_4__14_;
  wire w_mem_inst_w_mem_4__15_;
  wire w_mem_inst_w_mem_4__16_;
  wire w_mem_inst_w_mem_4__17_;
  wire w_mem_inst_w_mem_4__18_;
  wire w_mem_inst_w_mem_4__19_;
  wire w_mem_inst_w_mem_4__1_;
  wire w_mem_inst_w_mem_4__20_;
  wire w_mem_inst_w_mem_4__21_;
  wire w_mem_inst_w_mem_4__22_;
  wire w_mem_inst_w_mem_4__23_;
  wire w_mem_inst_w_mem_4__24_;
  wire w_mem_inst_w_mem_4__25_;
  wire w_mem_inst_w_mem_4__26_;
  wire w_mem_inst_w_mem_4__27_;
  wire w_mem_inst_w_mem_4__28_;
  wire w_mem_inst_w_mem_4__29_;
  wire w_mem_inst_w_mem_4__2_;
  wire w_mem_inst_w_mem_4__30_;
  wire w_mem_inst_w_mem_4__31_;
  wire w_mem_inst_w_mem_4__3_;
  wire w_mem_inst_w_mem_4__4_;
  wire w_mem_inst_w_mem_4__5_;
  wire w_mem_inst_w_mem_4__6_;
  wire w_mem_inst_w_mem_4__7_;
  wire w_mem_inst_w_mem_4__8_;
  wire w_mem_inst_w_mem_4__9_;
  wire w_mem_inst_w_mem_5__0_;
  wire w_mem_inst_w_mem_5__10_;
  wire w_mem_inst_w_mem_5__11_;
  wire w_mem_inst_w_mem_5__12_;
  wire w_mem_inst_w_mem_5__13_;
  wire w_mem_inst_w_mem_5__14_;
  wire w_mem_inst_w_mem_5__15_;
  wire w_mem_inst_w_mem_5__16_;
  wire w_mem_inst_w_mem_5__17_;
  wire w_mem_inst_w_mem_5__18_;
  wire w_mem_inst_w_mem_5__19_;
  wire w_mem_inst_w_mem_5__1_;
  wire w_mem_inst_w_mem_5__20_;
  wire w_mem_inst_w_mem_5__21_;
  wire w_mem_inst_w_mem_5__22_;
  wire w_mem_inst_w_mem_5__23_;
  wire w_mem_inst_w_mem_5__24_;
  wire w_mem_inst_w_mem_5__25_;
  wire w_mem_inst_w_mem_5__26_;
  wire w_mem_inst_w_mem_5__27_;
  wire w_mem_inst_w_mem_5__28_;
  wire w_mem_inst_w_mem_5__29_;
  wire w_mem_inst_w_mem_5__2_;
  wire w_mem_inst_w_mem_5__30_;
  wire w_mem_inst_w_mem_5__31_;
  wire w_mem_inst_w_mem_5__3_;
  wire w_mem_inst_w_mem_5__4_;
  wire w_mem_inst_w_mem_5__5_;
  wire w_mem_inst_w_mem_5__6_;
  wire w_mem_inst_w_mem_5__7_;
  wire w_mem_inst_w_mem_5__8_;
  wire w_mem_inst_w_mem_5__9_;
  wire w_mem_inst_w_mem_6__0_;
  wire w_mem_inst_w_mem_6__10_;
  wire w_mem_inst_w_mem_6__11_;
  wire w_mem_inst_w_mem_6__12_;
  wire w_mem_inst_w_mem_6__13_;
  wire w_mem_inst_w_mem_6__14_;
  wire w_mem_inst_w_mem_6__15_;
  wire w_mem_inst_w_mem_6__16_;
  wire w_mem_inst_w_mem_6__17_;
  wire w_mem_inst_w_mem_6__18_;
  wire w_mem_inst_w_mem_6__19_;
  wire w_mem_inst_w_mem_6__1_;
  wire w_mem_inst_w_mem_6__20_;
  wire w_mem_inst_w_mem_6__21_;
  wire w_mem_inst_w_mem_6__22_;
  wire w_mem_inst_w_mem_6__23_;
  wire w_mem_inst_w_mem_6__24_;
  wire w_mem_inst_w_mem_6__25_;
  wire w_mem_inst_w_mem_6__26_;
  wire w_mem_inst_w_mem_6__27_;
  wire w_mem_inst_w_mem_6__28_;
  wire w_mem_inst_w_mem_6__29_;
  wire w_mem_inst_w_mem_6__2_;
  wire w_mem_inst_w_mem_6__30_;
  wire w_mem_inst_w_mem_6__31_;
  wire w_mem_inst_w_mem_6__3_;
  wire w_mem_inst_w_mem_6__4_;
  wire w_mem_inst_w_mem_6__5_;
  wire w_mem_inst_w_mem_6__6_;
  wire w_mem_inst_w_mem_6__7_;
  wire w_mem_inst_w_mem_6__8_;
  wire w_mem_inst_w_mem_6__9_;
  wire w_mem_inst_w_mem_7__0_;
  wire w_mem_inst_w_mem_7__10_;
  wire w_mem_inst_w_mem_7__11_;
  wire w_mem_inst_w_mem_7__12_;
  wire w_mem_inst_w_mem_7__13_;
  wire w_mem_inst_w_mem_7__14_;
  wire w_mem_inst_w_mem_7__15_;
  wire w_mem_inst_w_mem_7__16_;
  wire w_mem_inst_w_mem_7__17_;
  wire w_mem_inst_w_mem_7__18_;
  wire w_mem_inst_w_mem_7__19_;
  wire w_mem_inst_w_mem_7__1_;
  wire w_mem_inst_w_mem_7__20_;
  wire w_mem_inst_w_mem_7__21_;
  wire w_mem_inst_w_mem_7__22_;
  wire w_mem_inst_w_mem_7__23_;
  wire w_mem_inst_w_mem_7__24_;
  wire w_mem_inst_w_mem_7__25_;
  wire w_mem_inst_w_mem_7__26_;
  wire w_mem_inst_w_mem_7__27_;
  wire w_mem_inst_w_mem_7__28_;
  wire w_mem_inst_w_mem_7__29_;
  wire w_mem_inst_w_mem_7__2_;
  wire w_mem_inst_w_mem_7__30_;
  wire w_mem_inst_w_mem_7__31_;
  wire w_mem_inst_w_mem_7__3_;
  wire w_mem_inst_w_mem_7__4_;
  wire w_mem_inst_w_mem_7__5_;
  wire w_mem_inst_w_mem_7__6_;
  wire w_mem_inst_w_mem_7__7_;
  wire w_mem_inst_w_mem_7__8_;
  wire w_mem_inst_w_mem_7__9_;
  wire w_mem_inst_w_mem_8__0_;
  wire w_mem_inst_w_mem_8__10_;
  wire w_mem_inst_w_mem_8__11_;
  wire w_mem_inst_w_mem_8__12_;
  wire w_mem_inst_w_mem_8__13_;
  wire w_mem_inst_w_mem_8__14_;
  wire w_mem_inst_w_mem_8__15_;
  wire w_mem_inst_w_mem_8__16_;
  wire w_mem_inst_w_mem_8__17_;
  wire w_mem_inst_w_mem_8__18_;
  wire w_mem_inst_w_mem_8__19_;
  wire w_mem_inst_w_mem_8__1_;
  wire w_mem_inst_w_mem_8__20_;
  wire w_mem_inst_w_mem_8__21_;
  wire w_mem_inst_w_mem_8__22_;
  wire w_mem_inst_w_mem_8__23_;
  wire w_mem_inst_w_mem_8__24_;
  wire w_mem_inst_w_mem_8__25_;
  wire w_mem_inst_w_mem_8__26_;
  wire w_mem_inst_w_mem_8__27_;
  wire w_mem_inst_w_mem_8__28_;
  wire w_mem_inst_w_mem_8__29_;
  wire w_mem_inst_w_mem_8__2_;
  wire w_mem_inst_w_mem_8__30_;
  wire w_mem_inst_w_mem_8__31_;
  wire w_mem_inst_w_mem_8__3_;
  wire w_mem_inst_w_mem_8__4_;
  wire w_mem_inst_w_mem_8__5_;
  wire w_mem_inst_w_mem_8__6_;
  wire w_mem_inst_w_mem_8__7_;
  wire w_mem_inst_w_mem_8__8_;
  wire w_mem_inst_w_mem_8__9_;
  wire w_mem_inst_w_mem_9__0_;
  wire w_mem_inst_w_mem_9__10_;
  wire w_mem_inst_w_mem_9__11_;
  wire w_mem_inst_w_mem_9__12_;
  wire w_mem_inst_w_mem_9__13_;
  wire w_mem_inst_w_mem_9__14_;
  wire w_mem_inst_w_mem_9__15_;
  wire w_mem_inst_w_mem_9__16_;
  wire w_mem_inst_w_mem_9__17_;
  wire w_mem_inst_w_mem_9__18_;
  wire w_mem_inst_w_mem_9__19_;
  wire w_mem_inst_w_mem_9__1_;
  wire w_mem_inst_w_mem_9__20_;
  wire w_mem_inst_w_mem_9__21_;
  wire w_mem_inst_w_mem_9__22_;
  wire w_mem_inst_w_mem_9__23_;
  wire w_mem_inst_w_mem_9__24_;
  wire w_mem_inst_w_mem_9__25_;
  wire w_mem_inst_w_mem_9__26_;
  wire w_mem_inst_w_mem_9__27_;
  wire w_mem_inst_w_mem_9__28_;
  wire w_mem_inst_w_mem_9__29_;
  wire w_mem_inst_w_mem_9__2_;
  wire w_mem_inst_w_mem_9__30_;
  wire w_mem_inst_w_mem_9__31_;
  wire w_mem_inst_w_mem_9__3_;
  wire w_mem_inst_w_mem_9__4_;
  wire w_mem_inst_w_mem_9__5_;
  wire w_mem_inst_w_mem_9__6_;
  wire w_mem_inst_w_mem_9__7_;
  wire w_mem_inst_w_mem_9__8_;
  wire w_mem_inst_w_mem_9__9_;
  AND2X2 AND2X2_1 ( .A(e_reg_21_), .B(_auto_iopadmap_cc_313_execute_26059_21_), .Y(_abc_15724_n698) );
  AND2X2 AND2X2_10 ( .A(_auto_iopadmap_cc_313_execute_26059_17_), .B(e_reg_17_), .Y(_abc_15724_n714) );
  AND2X2 AND2X2_100 ( .A(_abc_15724_n889), .B(_abc_15724_n850_bF_buf6), .Y(_abc_15724_n890) );
  AND2X2 AND2X2_1000 ( .A(_abc_15724_n2752), .B(_abc_15724_n2746), .Y(_abc_15724_n2757) );
  AND2X2 AND2X2_1001 ( .A(_auto_iopadmap_cc_313_execute_26059_146_), .B(a_reg_18_), .Y(_abc_15724_n2760) );
  AND2X2 AND2X2_1002 ( .A(_abc_15724_n2761), .B(_abc_15724_n2759), .Y(_abc_15724_n2762) );
  AND2X2 AND2X2_1003 ( .A(_abc_15724_n2758), .B(_abc_15724_n2762), .Y(_abc_15724_n2764) );
  AND2X2 AND2X2_1004 ( .A(_abc_15724_n2765), .B(_abc_15724_n2763), .Y(_abc_15724_n2766) );
  AND2X2 AND2X2_1005 ( .A(_abc_15724_n2766), .B(digest_update_bF_buf6), .Y(_abc_15724_n2767) );
  AND2X2 AND2X2_1006 ( .A(_abc_15724_n2768_1), .B(_abc_15724_n850_bF_buf3), .Y(_abc_15724_n2769) );
  AND2X2 AND2X2_1007 ( .A(_abc_15724_n2765), .B(_abc_15724_n2761), .Y(_abc_15724_n2771) );
  AND2X2 AND2X2_1008 ( .A(_auto_iopadmap_cc_313_execute_26059_147_), .B(a_reg_19_), .Y(_abc_15724_n2773) );
  AND2X2 AND2X2_1009 ( .A(_abc_15724_n2774), .B(_abc_15724_n2772_1), .Y(_abc_15724_n2775) );
  AND2X2 AND2X2_101 ( .A(_abc_15724_n886), .B(_abc_15724_n882), .Y(_abc_15724_n892) );
  AND2X2 AND2X2_1010 ( .A(_abc_15724_n2771), .B(_abc_15724_n2775), .Y(_abc_15724_n2776) );
  AND2X2 AND2X2_1011 ( .A(_abc_15724_n2777), .B(_abc_15724_n2778), .Y(_abc_15724_n2779) );
  AND2X2 AND2X2_1012 ( .A(_abc_15724_n2780), .B(digest_update_bF_buf5), .Y(_abc_15724_n2781) );
  AND2X2 AND2X2_1013 ( .A(_abc_15724_n907_1_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_147_), .Y(_abc_15724_n2782) );
  AND2X2 AND2X2_1014 ( .A(_abc_15724_n907_1_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_148_), .Y(_abc_15724_n2784) );
  AND2X2 AND2X2_1015 ( .A(_abc_15724_n2735), .B(_abc_15724_n2747), .Y(_abc_15724_n2785) );
  AND2X2 AND2X2_1016 ( .A(_abc_15724_n2762), .B(_abc_15724_n2775), .Y(_abc_15724_n2786) );
  AND2X2 AND2X2_1017 ( .A(_abc_15724_n2785), .B(_abc_15724_n2786), .Y(_abc_15724_n2787) );
  AND2X2 AND2X2_1018 ( .A(_abc_15724_n2744), .B(_abc_15724_n2733), .Y(_abc_15724_n2790) );
  AND2X2 AND2X2_1019 ( .A(_abc_15724_n2786), .B(_abc_15724_n2791), .Y(_abc_15724_n2792) );
  AND2X2 AND2X2_102 ( .A(e_reg_25_), .B(_auto_iopadmap_cc_313_execute_26059_25_), .Y(_abc_15724_n895) );
  AND2X2 AND2X2_1020 ( .A(_abc_15724_n2772_1), .B(_abc_15724_n2760), .Y(_abc_15724_n2793) );
  AND2X2 AND2X2_1021 ( .A(_abc_15724_n2789), .B(_abc_15724_n2796), .Y(_abc_15724_n2797) );
  AND2X2 AND2X2_1022 ( .A(_auto_iopadmap_cc_313_execute_26059_148_), .B(a_reg_20_), .Y(_abc_15724_n2800) );
  AND2X2 AND2X2_1023 ( .A(_abc_15724_n2801), .B(_abc_15724_n2799), .Y(_abc_15724_n2802) );
  AND2X2 AND2X2_1024 ( .A(_abc_15724_n2798), .B(_abc_15724_n2802), .Y(_abc_15724_n2804) );
  AND2X2 AND2X2_1025 ( .A(_abc_15724_n2805), .B(_abc_15724_n2803), .Y(_abc_15724_n2806) );
  AND2X2 AND2X2_1026 ( .A(_abc_15724_n2806), .B(digest_update_bF_buf4), .Y(_abc_15724_n2807) );
  AND2X2 AND2X2_1027 ( .A(_auto_iopadmap_cc_313_execute_26059_149_), .B(a_reg_21_), .Y(_abc_15724_n2810) );
  AND2X2 AND2X2_1028 ( .A(_abc_15724_n2811), .B(_abc_15724_n2809), .Y(_abc_15724_n2812_1) );
  AND2X2 AND2X2_1029 ( .A(_abc_15724_n2805), .B(_abc_15724_n2801), .Y(_abc_15724_n2813) );
  AND2X2 AND2X2_103 ( .A(_abc_15724_n896), .B(_abc_15724_n894), .Y(_abc_15724_n897_1) );
  AND2X2 AND2X2_1030 ( .A(_abc_15724_n2814), .B(_abc_15724_n2812_1), .Y(_abc_15724_n2816) );
  AND2X2 AND2X2_1031 ( .A(_abc_15724_n2817), .B(_abc_15724_n2815), .Y(_abc_15724_n2818) );
  AND2X2 AND2X2_1032 ( .A(_abc_15724_n2818), .B(digest_update_bF_buf3), .Y(_abc_15724_n2819) );
  AND2X2 AND2X2_1033 ( .A(_abc_15724_n907_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_149_), .Y(_abc_15724_n2820) );
  AND2X2 AND2X2_1034 ( .A(_auto_iopadmap_cc_313_execute_26059_150_), .B(a_reg_22_), .Y(_abc_15724_n2824) );
  AND2X2 AND2X2_1035 ( .A(_abc_15724_n2825), .B(_abc_15724_n2823), .Y(_abc_15724_n2826) );
  AND2X2 AND2X2_1036 ( .A(_abc_15724_n2822), .B(_abc_15724_n2826), .Y(_abc_15724_n2828) );
  AND2X2 AND2X2_1037 ( .A(_abc_15724_n2829), .B(_abc_15724_n2827), .Y(_abc_15724_n2830) );
  AND2X2 AND2X2_1038 ( .A(_abc_15724_n2830), .B(digest_update_bF_buf2), .Y(_abc_15724_n2831) );
  AND2X2 AND2X2_1039 ( .A(_abc_15724_n2832), .B(_abc_15724_n850_bF_buf2), .Y(_abc_15724_n2833) );
  AND2X2 AND2X2_104 ( .A(_abc_15724_n898_1), .B(_abc_15724_n900), .Y(_abc_15724_n901) );
  AND2X2 AND2X2_1040 ( .A(_auto_iopadmap_cc_313_execute_26059_151_), .B(a_reg_23_), .Y(_abc_15724_n2838) );
  AND2X2 AND2X2_1041 ( .A(_abc_15724_n2839), .B(_abc_15724_n2837), .Y(_abc_15724_n2840) );
  AND2X2 AND2X2_1042 ( .A(_abc_15724_n2836), .B(_abc_15724_n2840), .Y(_abc_15724_n2841) );
  AND2X2 AND2X2_1043 ( .A(_abc_15724_n2835), .B(_abc_15724_n2842), .Y(_abc_15724_n2843) );
  AND2X2 AND2X2_1044 ( .A(_abc_15724_n2844), .B(digest_update_bF_buf1), .Y(_abc_15724_n2845_1) );
  AND2X2 AND2X2_1045 ( .A(_abc_15724_n907_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_151_), .Y(_abc_15724_n2846) );
  AND2X2 AND2X2_1046 ( .A(_abc_15724_n2809), .B(_abc_15724_n2800), .Y(_abc_15724_n2848_1) );
  AND2X2 AND2X2_1047 ( .A(_abc_15724_n2826), .B(_abc_15724_n2840), .Y(_abc_15724_n2850) );
  AND2X2 AND2X2_1048 ( .A(_abc_15724_n2850), .B(_abc_15724_n2849), .Y(_abc_15724_n2851) );
  AND2X2 AND2X2_1049 ( .A(_abc_15724_n2837), .B(_abc_15724_n2824), .Y(_abc_15724_n2852) );
  AND2X2 AND2X2_105 ( .A(_abc_15724_n901), .B(digest_update_bF_buf7), .Y(_abc_15724_n902) );
  AND2X2 AND2X2_1050 ( .A(_abc_15724_n2802), .B(_abc_15724_n2812_1), .Y(_abc_15724_n2856) );
  AND2X2 AND2X2_1051 ( .A(_abc_15724_n2856), .B(_abc_15724_n2850), .Y(_abc_15724_n2857) );
  AND2X2 AND2X2_1052 ( .A(_abc_15724_n2859), .B(_abc_15724_n2855), .Y(_abc_15724_n2860) );
  AND2X2 AND2X2_1053 ( .A(_auto_iopadmap_cc_313_execute_26059_152_), .B(a_reg_24_), .Y(_abc_15724_n2863) );
  AND2X2 AND2X2_1054 ( .A(_abc_15724_n2864), .B(_abc_15724_n2862), .Y(_abc_15724_n2865) );
  AND2X2 AND2X2_1055 ( .A(_abc_15724_n2861), .B(_abc_15724_n2865), .Y(_abc_15724_n2867) );
  AND2X2 AND2X2_1056 ( .A(_abc_15724_n2868), .B(_abc_15724_n2866), .Y(_abc_15724_n2869) );
  AND2X2 AND2X2_1057 ( .A(_abc_15724_n2869), .B(digest_update_bF_buf0), .Y(_abc_15724_n2870) );
  AND2X2 AND2X2_1058 ( .A(_abc_15724_n2871), .B(_abc_15724_n850_bF_buf1), .Y(_abc_15724_n2872) );
  AND2X2 AND2X2_1059 ( .A(_abc_15724_n2868), .B(_abc_15724_n2864), .Y(_abc_15724_n2874) );
  AND2X2 AND2X2_106 ( .A(_abc_15724_n903), .B(_abc_15724_n850_bF_buf5), .Y(_abc_15724_n904) );
  AND2X2 AND2X2_1060 ( .A(_auto_iopadmap_cc_313_execute_26059_153_), .B(a_reg_25_), .Y(_abc_15724_n2877) );
  AND2X2 AND2X2_1061 ( .A(_abc_15724_n2878), .B(_abc_15724_n2876), .Y(_abc_15724_n2879) );
  AND2X2 AND2X2_1062 ( .A(_abc_15724_n2880), .B(_abc_15724_n2882), .Y(_abc_15724_n2883) );
  AND2X2 AND2X2_1063 ( .A(_abc_15724_n2883), .B(digest_update_bF_buf11), .Y(_abc_15724_n2884) );
  AND2X2 AND2X2_1064 ( .A(_abc_15724_n2885), .B(_abc_15724_n850_bF_buf0), .Y(_abc_15724_n2886) );
  AND2X2 AND2X2_1065 ( .A(_abc_15724_n2865), .B(_abc_15724_n2879), .Y(_abc_15724_n2888) );
  AND2X2 AND2X2_1066 ( .A(_abc_15724_n2861), .B(_abc_15724_n2888), .Y(_abc_15724_n2889) );
  AND2X2 AND2X2_1067 ( .A(_abc_15724_n2876), .B(_abc_15724_n2863), .Y(_abc_15724_n2890_1) );
  AND2X2 AND2X2_1068 ( .A(_auto_iopadmap_cc_313_execute_26059_154_), .B(a_reg_26_), .Y(_abc_15724_n2894_1) );
  AND2X2 AND2X2_1069 ( .A(_abc_15724_n2895), .B(_abc_15724_n2893), .Y(_abc_15724_n2896) );
  AND2X2 AND2X2_107 ( .A(_abc_15724_n906_bF_buf8), .B(_abc_15724_n850_bF_buf4), .Y(_abc_15724_n907_1) );
  AND2X2 AND2X2_1070 ( .A(_abc_15724_n2892), .B(_abc_15724_n2896), .Y(_abc_15724_n2898) );
  AND2X2 AND2X2_1071 ( .A(_abc_15724_n2899), .B(_abc_15724_n2897), .Y(_abc_15724_n2900) );
  AND2X2 AND2X2_1072 ( .A(_abc_15724_n2900), .B(digest_update_bF_buf10), .Y(_abc_15724_n2901) );
  AND2X2 AND2X2_1073 ( .A(_abc_15724_n2902), .B(_abc_15724_n850_bF_buf8), .Y(_abc_15724_n2903) );
  AND2X2 AND2X2_1074 ( .A(_abc_15724_n907_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_155_), .Y(_abc_15724_n2905) );
  AND2X2 AND2X2_1075 ( .A(_auto_iopadmap_cc_313_execute_26059_155_), .B(a_reg_27_), .Y(_abc_15724_n2907) );
  AND2X2 AND2X2_1076 ( .A(_abc_15724_n2908), .B(_abc_15724_n2906), .Y(_abc_15724_n2909) );
  AND2X2 AND2X2_1077 ( .A(_abc_15724_n2899), .B(_abc_15724_n2895), .Y(_abc_15724_n2913) );
  AND2X2 AND2X2_1078 ( .A(_abc_15724_n2914), .B(_abc_15724_n2911), .Y(_abc_15724_n2915) );
  AND2X2 AND2X2_1079 ( .A(_abc_15724_n2915), .B(digest_update_bF_buf9), .Y(_abc_15724_n2916) );
  AND2X2 AND2X2_108 ( .A(_abc_15724_n907_1_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_26_), .Y(_abc_15724_n908_1) );
  AND2X2 AND2X2_1080 ( .A(_abc_15724_n907_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_156_), .Y(_abc_15724_n2918) );
  AND2X2 AND2X2_1081 ( .A(_abc_15724_n2909), .B(_abc_15724_n2894_1), .Y(_abc_15724_n2919) );
  AND2X2 AND2X2_1082 ( .A(_abc_15724_n2920), .B(_abc_15724_n2908), .Y(_abc_15724_n2921) );
  AND2X2 AND2X2_1083 ( .A(_abc_15724_n2896), .B(_abc_15724_n2909), .Y(_abc_15724_n2922) );
  AND2X2 AND2X2_1084 ( .A(_abc_15724_n2922), .B(_abc_15724_n2891), .Y(_abc_15724_n2923) );
  AND2X2 AND2X2_1085 ( .A(_abc_15724_n2924), .B(_abc_15724_n2921), .Y(_abc_15724_n2925) );
  AND2X2 AND2X2_1086 ( .A(_abc_15724_n2888), .B(_abc_15724_n2922), .Y(_abc_15724_n2926) );
  AND2X2 AND2X2_1087 ( .A(_abc_15724_n2928), .B(_abc_15724_n2925), .Y(_abc_15724_n2929) );
  AND2X2 AND2X2_1088 ( .A(_auto_iopadmap_cc_313_execute_26059_156_), .B(a_reg_28_), .Y(_abc_15724_n2932) );
  AND2X2 AND2X2_1089 ( .A(_abc_15724_n2933), .B(_abc_15724_n2931), .Y(_abc_15724_n2934) );
  AND2X2 AND2X2_109 ( .A(_abc_15724_n883), .B(_abc_15724_n897_1), .Y(_abc_15724_n909_1) );
  AND2X2 AND2X2_1090 ( .A(_abc_15724_n2930_1), .B(_abc_15724_n2934), .Y(_abc_15724_n2936) );
  AND2X2 AND2X2_1091 ( .A(_abc_15724_n2937), .B(_abc_15724_n2935), .Y(_abc_15724_n2938) );
  AND2X2 AND2X2_1092 ( .A(_abc_15724_n2938), .B(digest_update_bF_buf8), .Y(_abc_15724_n2939) );
  AND2X2 AND2X2_1093 ( .A(_abc_15724_n2937), .B(_abc_15724_n2933), .Y(_abc_15724_n2941) );
  AND2X2 AND2X2_1094 ( .A(_auto_iopadmap_cc_313_execute_26059_157_), .B(a_reg_29_), .Y(_abc_15724_n2943) );
  AND2X2 AND2X2_1095 ( .A(_abc_15724_n2944), .B(_abc_15724_n2942), .Y(_abc_15724_n2945) );
  AND2X2 AND2X2_1096 ( .A(_abc_15724_n2949), .B(digest_update_bF_buf7), .Y(_abc_15724_n2950) );
  AND2X2 AND2X2_1097 ( .A(_abc_15724_n2950), .B(_abc_15724_n2947), .Y(_abc_15724_n2951) );
  AND2X2 AND2X2_1098 ( .A(_abc_15724_n2952), .B(_abc_15724_n850_bF_buf7), .Y(_abc_15724_n2953) );
  AND2X2 AND2X2_1099 ( .A(_auto_iopadmap_cc_313_execute_26059_158_), .B(a_reg_30_), .Y(_abc_15724_n2956) );
  AND2X2 AND2X2_11 ( .A(e_reg_16_), .B(_auto_iopadmap_cc_313_execute_26059_16_), .Y(_abc_15724_n716) );
  AND2X2 AND2X2_110 ( .A(_abc_15724_n879), .B(_abc_15724_n909_1), .Y(_abc_15724_n910) );
  AND2X2 AND2X2_1100 ( .A(_abc_15724_n2957), .B(_abc_15724_n2955), .Y(_abc_15724_n2958) );
  AND2X2 AND2X2_1101 ( .A(_abc_15724_n2945), .B(_abc_15724_n2932), .Y(_abc_15724_n2959) );
  AND2X2 AND2X2_1102 ( .A(_abc_15724_n2934), .B(_abc_15724_n2945), .Y(_abc_15724_n2962) );
  AND2X2 AND2X2_1103 ( .A(_abc_15724_n2964_1), .B(_abc_15724_n2961), .Y(_abc_15724_n2965) );
  AND2X2 AND2X2_1104 ( .A(_abc_15724_n2969), .B(digest_update_bF_buf6), .Y(_abc_15724_n2970) );
  AND2X2 AND2X2_1105 ( .A(_abc_15724_n2970), .B(_abc_15724_n2967), .Y(_abc_15724_n2971) );
  AND2X2 AND2X2_1106 ( .A(_abc_15724_n2972), .B(_abc_15724_n850_bF_buf6), .Y(_abc_15724_n2973) );
  AND2X2 AND2X2_1107 ( .A(_abc_15724_n2969), .B(_abc_15724_n2957), .Y(_abc_15724_n2975) );
  AND2X2 AND2X2_1108 ( .A(_auto_iopadmap_cc_313_execute_26059_159_), .B(a_reg_31_), .Y(_abc_15724_n2977) );
  AND2X2 AND2X2_1109 ( .A(_abc_15724_n2978), .B(_abc_15724_n2976), .Y(_abc_15724_n2979) );
  AND2X2 AND2X2_111 ( .A(_abc_15724_n894), .B(_abc_15724_n881), .Y(_abc_15724_n911) );
  AND2X2 AND2X2_1110 ( .A(_abc_15724_n2975), .B(_abc_15724_n2979), .Y(_abc_15724_n2980) );
  AND2X2 AND2X2_1111 ( .A(_abc_15724_n2981), .B(_abc_15724_n2982), .Y(_abc_15724_n2983) );
  AND2X2 AND2X2_1112 ( .A(_abc_15724_n2984), .B(digest_update_bF_buf5), .Y(_abc_15724_n2985) );
  AND2X2 AND2X2_1113 ( .A(_abc_15724_n907_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_159_), .Y(_abc_15724_n2986) );
  AND2X2 AND2X2_1114 ( .A(_abc_15724_n2988), .B(_auto_iopadmap_cc_313_execute_26222), .Y(round_ctr_rst) );
  AND2X2 AND2X2_1115 ( .A(_abc_15724_n2991), .B(_abc_15724_n2990), .Y(_abc_15724_n2992) );
  AND2X2 AND2X2_1116 ( .A(_abc_15724_n2992_bF_buf11), .B(e_reg_0_), .Y(_abc_15724_n2993) );
  AND2X2 AND2X2_1117 ( .A(round_ctr_rst_bF_buf62), .B(_abc_15724_n2990), .Y(_abc_15724_n2994) );
  AND2X2 AND2X2_1118 ( .A(_abc_15724_n906_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_0_), .Y(_abc_15724_n2995) );
  AND2X2 AND2X2_1119 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n2995), .Y(_abc_15724_n2996) );
  AND2X2 AND2X2_112 ( .A(_auto_iopadmap_cc_313_execute_26059_26_), .B(e_reg_26_), .Y(_abc_15724_n915) );
  AND2X2 AND2X2_1120 ( .A(d_reg_0_), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n2997) );
  AND2X2 AND2X2_1121 ( .A(_abc_15724_n2992_bF_buf10), .B(e_reg_1_), .Y(_abc_15724_n3000) );
  AND2X2 AND2X2_1122 ( .A(_abc_15724_n906_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_1_), .Y(_abc_15724_n3001) );
  AND2X2 AND2X2_1123 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n3001), .Y(_abc_15724_n3002) );
  AND2X2 AND2X2_1124 ( .A(d_reg_1_), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n3003_1) );
  AND2X2 AND2X2_1125 ( .A(_abc_15724_n2992_bF_buf9), .B(e_reg_2_), .Y(_abc_15724_n3006) );
  AND2X2 AND2X2_1126 ( .A(_abc_15724_n906_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_2_), .Y(_abc_15724_n3007) );
  AND2X2 AND2X2_1127 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n3007), .Y(_abc_15724_n3008) );
  AND2X2 AND2X2_1128 ( .A(d_reg_2_), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n3009) );
  AND2X2 AND2X2_1129 ( .A(_abc_15724_n2992_bF_buf8), .B(e_reg_3_), .Y(_abc_15724_n3012) );
  AND2X2 AND2X2_113 ( .A(_abc_15724_n916), .B(_abc_15724_n914), .Y(_abc_15724_n917) );
  AND2X2 AND2X2_1130 ( .A(_abc_15724_n906_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_3_), .Y(_abc_15724_n3013) );
  AND2X2 AND2X2_1131 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n3013), .Y(_abc_15724_n3014) );
  AND2X2 AND2X2_1132 ( .A(d_reg_3_), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n3015) );
  AND2X2 AND2X2_1133 ( .A(_abc_15724_n2992_bF_buf7), .B(e_reg_4_), .Y(_abc_15724_n3018) );
  AND2X2 AND2X2_1134 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n3019), .Y(_abc_15724_n3020) );
  AND2X2 AND2X2_1135 ( .A(d_reg_4_), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n3021) );
  AND2X2 AND2X2_1136 ( .A(_abc_15724_n2992_bF_buf6), .B(e_reg_5_), .Y(_abc_15724_n3024) );
  AND2X2 AND2X2_1137 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n3025), .Y(_abc_15724_n3026) );
  AND2X2 AND2X2_1138 ( .A(d_reg_5_), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n3027) );
  AND2X2 AND2X2_1139 ( .A(_abc_15724_n2992_bF_buf5), .B(e_reg_6_), .Y(_abc_15724_n3030) );
  AND2X2 AND2X2_114 ( .A(_abc_15724_n913), .B(_abc_15724_n917), .Y(_abc_15724_n919) );
  AND2X2 AND2X2_1140 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n3031), .Y(_abc_15724_n3032) );
  AND2X2 AND2X2_1141 ( .A(d_reg_6_), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n3033) );
  AND2X2 AND2X2_1142 ( .A(_abc_15724_n2992_bF_buf4), .B(e_reg_7_), .Y(_abc_15724_n3036) );
  AND2X2 AND2X2_1143 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n3037), .Y(_abc_15724_n3038) );
  AND2X2 AND2X2_1144 ( .A(d_reg_7_), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n3039) );
  AND2X2 AND2X2_1145 ( .A(_abc_15724_n2992_bF_buf3), .B(e_reg_8_), .Y(_abc_15724_n3042) );
  AND2X2 AND2X2_1146 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n3043), .Y(_abc_15724_n3044_1) );
  AND2X2 AND2X2_1147 ( .A(d_reg_8_), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n3045) );
  AND2X2 AND2X2_1148 ( .A(_abc_15724_n2992_bF_buf2), .B(e_reg_9_), .Y(_abc_15724_n3048) );
  AND2X2 AND2X2_1149 ( .A(_abc_15724_n906_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_9_), .Y(_abc_15724_n3049) );
  AND2X2 AND2X2_115 ( .A(_abc_15724_n920), .B(_abc_15724_n918), .Y(_abc_15724_n921_1) );
  AND2X2 AND2X2_1150 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n3049), .Y(_abc_15724_n3050) );
  AND2X2 AND2X2_1151 ( .A(d_reg_9_), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n3051) );
  AND2X2 AND2X2_1152 ( .A(_abc_15724_n2992_bF_buf1), .B(e_reg_10_), .Y(_abc_15724_n3054) );
  AND2X2 AND2X2_1153 ( .A(_abc_15724_n906_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_10_), .Y(_abc_15724_n3055) );
  AND2X2 AND2X2_1154 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n3055), .Y(_abc_15724_n3056) );
  AND2X2 AND2X2_1155 ( .A(d_reg_10_), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n3057) );
  AND2X2 AND2X2_1156 ( .A(_abc_15724_n2992_bF_buf0), .B(e_reg_11_), .Y(_abc_15724_n3060) );
  AND2X2 AND2X2_1157 ( .A(_abc_15724_n906_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_11_), .Y(_abc_15724_n3061) );
  AND2X2 AND2X2_1158 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n3061), .Y(_abc_15724_n3062) );
  AND2X2 AND2X2_1159 ( .A(d_reg_11_), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n3063) );
  AND2X2 AND2X2_116 ( .A(_abc_15724_n921_1), .B(digest_update_bF_buf6), .Y(_abc_15724_n922_1) );
  AND2X2 AND2X2_1160 ( .A(_abc_15724_n2992_bF_buf11), .B(e_reg_12_), .Y(_abc_15724_n3066) );
  AND2X2 AND2X2_1161 ( .A(_abc_15724_n906_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_12_), .Y(_abc_15724_n3067) );
  AND2X2 AND2X2_1162 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n3067), .Y(_abc_15724_n3068) );
  AND2X2 AND2X2_1163 ( .A(d_reg_12_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n3069) );
  AND2X2 AND2X2_1164 ( .A(_abc_15724_n2992_bF_buf10), .B(e_reg_13_), .Y(_abc_15724_n3072) );
  AND2X2 AND2X2_1165 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n3073), .Y(_abc_15724_n3074) );
  AND2X2 AND2X2_1166 ( .A(d_reg_13_), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n3075) );
  AND2X2 AND2X2_1167 ( .A(_abc_15724_n2992_bF_buf9), .B(e_reg_14_), .Y(_abc_15724_n3078) );
  AND2X2 AND2X2_1168 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n3079_1), .Y(_abc_15724_n3080) );
  AND2X2 AND2X2_1169 ( .A(d_reg_14_), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n3081) );
  AND2X2 AND2X2_117 ( .A(_abc_15724_n907_1_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_27_), .Y(_abc_15724_n924) );
  AND2X2 AND2X2_1170 ( .A(_abc_15724_n2992_bF_buf8), .B(e_reg_15_), .Y(_abc_15724_n3084) );
  AND2X2 AND2X2_1171 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n3085), .Y(_abc_15724_n3086) );
  AND2X2 AND2X2_1172 ( .A(d_reg_15_), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n3087) );
  AND2X2 AND2X2_1173 ( .A(_abc_15724_n2992_bF_buf7), .B(e_reg_16_), .Y(_abc_15724_n3090) );
  AND2X2 AND2X2_1174 ( .A(_abc_15724_n906_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_16_), .Y(_abc_15724_n3091) );
  AND2X2 AND2X2_1175 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n3091), .Y(_abc_15724_n3092) );
  AND2X2 AND2X2_1176 ( .A(d_reg_16_), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n3093) );
  AND2X2 AND2X2_1177 ( .A(_abc_15724_n2992_bF_buf6), .B(e_reg_17_), .Y(_abc_15724_n3096) );
  AND2X2 AND2X2_1178 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n3097), .Y(_abc_15724_n3098) );
  AND2X2 AND2X2_1179 ( .A(d_reg_17_), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n3099) );
  AND2X2 AND2X2_118 ( .A(_auto_iopadmap_cc_313_execute_26059_27_), .B(e_reg_27_), .Y(_abc_15724_n926) );
  AND2X2 AND2X2_1180 ( .A(_abc_15724_n2992_bF_buf5), .B(e_reg_18_), .Y(_abc_15724_n3102) );
  AND2X2 AND2X2_1181 ( .A(_abc_15724_n906_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_18_), .Y(_abc_15724_n3103) );
  AND2X2 AND2X2_1182 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n3103), .Y(_abc_15724_n3104) );
  AND2X2 AND2X2_1183 ( .A(d_reg_18_), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n3105) );
  AND2X2 AND2X2_1184 ( .A(_abc_15724_n2992_bF_buf4), .B(e_reg_19_), .Y(_abc_15724_n3108) );
  AND2X2 AND2X2_1185 ( .A(_abc_15724_n906_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_19_), .Y(_abc_15724_n3109) );
  AND2X2 AND2X2_1186 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n3109), .Y(_abc_15724_n3110) );
  AND2X2 AND2X2_1187 ( .A(d_reg_19_), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n3111) );
  AND2X2 AND2X2_1188 ( .A(_abc_15724_n2992_bF_buf3), .B(e_reg_20_), .Y(_abc_15724_n3114_1) );
  AND2X2 AND2X2_1189 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n3115), .Y(_abc_15724_n3116) );
  AND2X2 AND2X2_119 ( .A(_abc_15724_n927), .B(_abc_15724_n925), .Y(_abc_15724_n928) );
  AND2X2 AND2X2_1190 ( .A(d_reg_20_), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n3117) );
  AND2X2 AND2X2_1191 ( .A(_abc_15724_n2992_bF_buf2), .B(e_reg_21_), .Y(_abc_15724_n3120) );
  AND2X2 AND2X2_1192 ( .A(_abc_15724_n906_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_21_), .Y(_abc_15724_n3121) );
  AND2X2 AND2X2_1193 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n3121), .Y(_abc_15724_n3122) );
  AND2X2 AND2X2_1194 ( .A(d_reg_21_), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n3123) );
  AND2X2 AND2X2_1195 ( .A(_abc_15724_n2992_bF_buf1), .B(e_reg_22_), .Y(_abc_15724_n3126) );
  AND2X2 AND2X2_1196 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n852), .Y(_abc_15724_n3127) );
  AND2X2 AND2X2_1197 ( .A(d_reg_22_), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n3128) );
  AND2X2 AND2X2_1198 ( .A(_abc_15724_n2992_bF_buf0), .B(e_reg_23_), .Y(_abc_15724_n3131) );
  AND2X2 AND2X2_1199 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n866_1), .Y(_abc_15724_n3132) );
  AND2X2 AND2X2_12 ( .A(_abc_15724_n715), .B(_abc_15724_n718_1), .Y(_abc_15724_n719_1) );
  AND2X2 AND2X2_120 ( .A(_abc_15724_n917), .B(_abc_15724_n928), .Y(_abc_15724_n931_1) );
  AND2X2 AND2X2_1200 ( .A(d_reg_23_), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n3133) );
  AND2X2 AND2X2_1201 ( .A(_abc_15724_n2992_bF_buf11), .B(e_reg_24_), .Y(_abc_15724_n3136) );
  AND2X2 AND2X2_1202 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n889), .Y(_abc_15724_n3137) );
  AND2X2 AND2X2_1203 ( .A(d_reg_24_), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n3138) );
  AND2X2 AND2X2_1204 ( .A(_abc_15724_n2992_bF_buf10), .B(e_reg_25_), .Y(_abc_15724_n3141) );
  AND2X2 AND2X2_1205 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n903), .Y(_abc_15724_n3142) );
  AND2X2 AND2X2_1206 ( .A(d_reg_25_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n3143) );
  AND2X2 AND2X2_1207 ( .A(_abc_15724_n2992_bF_buf9), .B(e_reg_26_), .Y(_abc_15724_n3146) );
  AND2X2 AND2X2_1208 ( .A(_abc_15724_n906_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_26_), .Y(_abc_15724_n3147) );
  AND2X2 AND2X2_1209 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n3147), .Y(_abc_15724_n3148) );
  AND2X2 AND2X2_121 ( .A(_abc_15724_n913), .B(_abc_15724_n931_1), .Y(_abc_15724_n932_1) );
  AND2X2 AND2X2_1210 ( .A(d_reg_26_), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n3149) );
  AND2X2 AND2X2_1211 ( .A(_abc_15724_n2992_bF_buf8), .B(e_reg_27_), .Y(_abc_15724_n3152) );
  AND2X2 AND2X2_1212 ( .A(_abc_15724_n906_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_27_), .Y(_abc_15724_n3153_1) );
  AND2X2 AND2X2_1213 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n3153_1), .Y(_abc_15724_n3154) );
  AND2X2 AND2X2_1214 ( .A(d_reg_27_), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n3155) );
  AND2X2 AND2X2_1215 ( .A(_abc_15724_n2992_bF_buf7), .B(e_reg_28_), .Y(_abc_15724_n3158) );
  AND2X2 AND2X2_1216 ( .A(_abc_15724_n906_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_28_), .Y(_abc_15724_n3159) );
  AND2X2 AND2X2_1217 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n3159), .Y(_abc_15724_n3160) );
  AND2X2 AND2X2_1218 ( .A(d_reg_28_), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n3161) );
  AND2X2 AND2X2_1219 ( .A(_abc_15724_n2992_bF_buf6), .B(e_reg_29_), .Y(_abc_15724_n3164) );
  AND2X2 AND2X2_122 ( .A(_abc_15724_n928), .B(_abc_15724_n915), .Y(_abc_15724_n934_1) );
  AND2X2 AND2X2_1220 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n954_1), .Y(_abc_15724_n3165) );
  AND2X2 AND2X2_1221 ( .A(d_reg_29_), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n3166) );
  AND2X2 AND2X2_1222 ( .A(_abc_15724_n2992_bF_buf5), .B(e_reg_30_), .Y(_abc_15724_n3169) );
  AND2X2 AND2X2_1223 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n982), .Y(_abc_15724_n3170) );
  AND2X2 AND2X2_1224 ( .A(d_reg_30_), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n3171) );
  AND2X2 AND2X2_1225 ( .A(_abc_15724_n2992_bF_buf4), .B(e_reg_31_), .Y(_abc_15724_n3174) );
  AND2X2 AND2X2_1226 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n997_1), .Y(_abc_15724_n3175) );
  AND2X2 AND2X2_1227 ( .A(d_reg_31_), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n3176) );
  AND2X2 AND2X2_1228 ( .A(_abc_15724_n2992_bF_buf3), .B(d_reg_0_), .Y(_abc_15724_n3179) );
  AND2X2 AND2X2_1229 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n1005), .Y(_abc_15724_n3180) );
  AND2X2 AND2X2_123 ( .A(_abc_15724_n935), .B(digest_update_bF_buf5), .Y(_abc_15724_n936) );
  AND2X2 AND2X2_1230 ( .A(c_reg_0_), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n3181) );
  AND2X2 AND2X2_1231 ( .A(_abc_15724_n2992_bF_buf2), .B(d_reg_1_), .Y(_abc_15724_n3184) );
  AND2X2 AND2X2_1232 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n1020), .Y(_abc_15724_n3185) );
  AND2X2 AND2X2_1233 ( .A(c_reg_1_), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n3186) );
  AND2X2 AND2X2_1234 ( .A(_abc_15724_n2992_bF_buf1), .B(d_reg_2_), .Y(_abc_15724_n3189) );
  AND2X2 AND2X2_1235 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n1035), .Y(_abc_15724_n3190) );
  AND2X2 AND2X2_1236 ( .A(c_reg_2_), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n3191) );
  AND2X2 AND2X2_1237 ( .A(_abc_15724_n2992_bF_buf0), .B(d_reg_3_), .Y(_abc_15724_n3194) );
  AND2X2 AND2X2_1238 ( .A(_abc_15724_n906_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_35_), .Y(_abc_15724_n3195_1) );
  AND2X2 AND2X2_1239 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n3195_1), .Y(_abc_15724_n3196) );
  AND2X2 AND2X2_124 ( .A(_abc_15724_n933), .B(_abc_15724_n936), .Y(_abc_15724_n937) );
  AND2X2 AND2X2_1240 ( .A(c_reg_3_), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n3197) );
  AND2X2 AND2X2_1241 ( .A(_abc_15724_n2992_bF_buf11), .B(d_reg_4_), .Y(_abc_15724_n3200) );
  AND2X2 AND2X2_1242 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n1066), .Y(_abc_15724_n3201) );
  AND2X2 AND2X2_1243 ( .A(c_reg_4_), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n3202) );
  AND2X2 AND2X2_1244 ( .A(_abc_15724_n2992_bF_buf10), .B(d_reg_5_), .Y(_abc_15724_n3205) );
  AND2X2 AND2X2_1245 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n1081), .Y(_abc_15724_n3206) );
  AND2X2 AND2X2_1246 ( .A(c_reg_5_), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n3207) );
  AND2X2 AND2X2_1247 ( .A(_abc_15724_n2992_bF_buf9), .B(d_reg_6_), .Y(_abc_15724_n3210) );
  AND2X2 AND2X2_1248 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n1096), .Y(_abc_15724_n3211) );
  AND2X2 AND2X2_1249 ( .A(c_reg_6_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n3212) );
  AND2X2 AND2X2_125 ( .A(_abc_15724_n937), .B(_abc_15724_n930), .Y(_abc_15724_n938) );
  AND2X2 AND2X2_1250 ( .A(_abc_15724_n2992_bF_buf8), .B(d_reg_7_), .Y(_abc_15724_n3215) );
  AND2X2 AND2X2_1251 ( .A(_abc_15724_n906_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_39_), .Y(_abc_15724_n3216) );
  AND2X2 AND2X2_1252 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n3216), .Y(_abc_15724_n3217) );
  AND2X2 AND2X2_1253 ( .A(c_reg_7_), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n3218) );
  AND2X2 AND2X2_1254 ( .A(_abc_15724_n2992_bF_buf7), .B(d_reg_8_), .Y(_abc_15724_n3221) );
  AND2X2 AND2X2_1255 ( .A(_abc_15724_n906_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_40_), .Y(_abc_15724_n3222) );
  AND2X2 AND2X2_1256 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n3222), .Y(_abc_15724_n3223) );
  AND2X2 AND2X2_1257 ( .A(c_reg_8_), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n3224) );
  AND2X2 AND2X2_1258 ( .A(_abc_15724_n2992_bF_buf6), .B(d_reg_9_), .Y(_abc_15724_n3227) );
  AND2X2 AND2X2_1259 ( .A(_abc_15724_n906_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_41_), .Y(_abc_15724_n3228) );
  AND2X2 AND2X2_126 ( .A(_abc_15724_n907_1_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_28_), .Y(_abc_15724_n940) );
  AND2X2 AND2X2_1260 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n3228), .Y(_abc_15724_n3229) );
  AND2X2 AND2X2_1261 ( .A(c_reg_9_), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n3230_1) );
  AND2X2 AND2X2_1262 ( .A(_abc_15724_n2992_bF_buf5), .B(d_reg_10_), .Y(_abc_15724_n3233_1) );
  AND2X2 AND2X2_1263 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n1150), .Y(_abc_15724_n3234) );
  AND2X2 AND2X2_1264 ( .A(c_reg_10_), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n3235) );
  AND2X2 AND2X2_1265 ( .A(_abc_15724_n2992_bF_buf4), .B(d_reg_11_), .Y(_abc_15724_n3238) );
  AND2X2 AND2X2_1266 ( .A(_abc_15724_n906_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_43_), .Y(_abc_15724_n3239) );
  AND2X2 AND2X2_1267 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n3239), .Y(_abc_15724_n3240) );
  AND2X2 AND2X2_1268 ( .A(c_reg_11_), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n3241) );
  AND2X2 AND2X2_1269 ( .A(_abc_15724_n2992_bF_buf3), .B(d_reg_12_), .Y(_abc_15724_n3244) );
  AND2X2 AND2X2_127 ( .A(_abc_15724_n935), .B(_abc_15724_n927), .Y(_abc_15724_n941) );
  AND2X2 AND2X2_1270 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n1186_1), .Y(_abc_15724_n3245) );
  AND2X2 AND2X2_1271 ( .A(c_reg_12_), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n3246) );
  AND2X2 AND2X2_1272 ( .A(_abc_15724_n2992_bF_buf2), .B(d_reg_13_), .Y(_abc_15724_n3249) );
  AND2X2 AND2X2_1273 ( .A(_abc_15724_n906_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_45_), .Y(_abc_15724_n3250) );
  AND2X2 AND2X2_1274 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n3250), .Y(_abc_15724_n3251) );
  AND2X2 AND2X2_1275 ( .A(c_reg_13_), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n3252) );
  AND2X2 AND2X2_1276 ( .A(_abc_15724_n2992_bF_buf1), .B(d_reg_14_), .Y(_abc_15724_n3255) );
  AND2X2 AND2X2_1277 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n1215_1), .Y(_abc_15724_n3256) );
  AND2X2 AND2X2_1278 ( .A(c_reg_14_), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n3257) );
  AND2X2 AND2X2_1279 ( .A(_abc_15724_n2992_bF_buf0), .B(d_reg_15_), .Y(_abc_15724_n3260) );
  AND2X2 AND2X2_128 ( .A(_auto_iopadmap_cc_313_execute_26059_28_), .B(e_reg_28_), .Y(_abc_15724_n945_1) );
  AND2X2 AND2X2_1280 ( .A(_abc_15724_n906_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_47_), .Y(_abc_15724_n3261) );
  AND2X2 AND2X2_1281 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n3261), .Y(_abc_15724_n3262) );
  AND2X2 AND2X2_1282 ( .A(c_reg_15_), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n3263) );
  AND2X2 AND2X2_1283 ( .A(_abc_15724_n2992_bF_buf11), .B(d_reg_16_), .Y(_abc_15724_n3266) );
  AND2X2 AND2X2_1284 ( .A(_abc_15724_n906_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_48_), .Y(_abc_15724_n3267) );
  AND2X2 AND2X2_1285 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n3267), .Y(_abc_15724_n3268) );
  AND2X2 AND2X2_1286 ( .A(c_reg_16_), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n3269) );
  AND2X2 AND2X2_1287 ( .A(_abc_15724_n2992_bF_buf10), .B(d_reg_17_), .Y(_abc_15724_n3272) );
  AND2X2 AND2X2_1288 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n1265), .Y(_abc_15724_n3273) );
  AND2X2 AND2X2_1289 ( .A(c_reg_17_), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n3274_1) );
  AND2X2 AND2X2_129 ( .A(_abc_15724_n946), .B(_abc_15724_n944_1), .Y(_abc_15724_n947) );
  AND2X2 AND2X2_1290 ( .A(_abc_15724_n2992_bF_buf9), .B(d_reg_18_), .Y(_abc_15724_n3277) );
  AND2X2 AND2X2_1291 ( .A(_abc_15724_n906_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_50_), .Y(_abc_15724_n3278) );
  AND2X2 AND2X2_1292 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n3278), .Y(_abc_15724_n3279) );
  AND2X2 AND2X2_1293 ( .A(c_reg_18_), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n3280) );
  AND2X2 AND2X2_1294 ( .A(_abc_15724_n2992_bF_buf8), .B(d_reg_19_), .Y(_abc_15724_n3283) );
  AND2X2 AND2X2_1295 ( .A(_abc_15724_n906_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_51_), .Y(_abc_15724_n3284) );
  AND2X2 AND2X2_1296 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n3284), .Y(_abc_15724_n3285) );
  AND2X2 AND2X2_1297 ( .A(c_reg_19_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n3286) );
  AND2X2 AND2X2_1298 ( .A(_abc_15724_n2992_bF_buf7), .B(d_reg_20_), .Y(_abc_15724_n3289) );
  AND2X2 AND2X2_1299 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n1319_1), .Y(_abc_15724_n3290) );
  AND2X2 AND2X2_13 ( .A(_abc_15724_n721_1), .B(_abc_15724_n715), .Y(_abc_15724_n722) );
  AND2X2 AND2X2_130 ( .A(_abc_15724_n943_1), .B(_abc_15724_n947), .Y(_abc_15724_n949) );
  AND2X2 AND2X2_1300 ( .A(c_reg_20_), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n3291) );
  AND2X2 AND2X2_1301 ( .A(_abc_15724_n2992_bF_buf6), .B(d_reg_21_), .Y(_abc_15724_n3294) );
  AND2X2 AND2X2_1302 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n1333), .Y(_abc_15724_n3295) );
  AND2X2 AND2X2_1303 ( .A(c_reg_21_), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n3296) );
  AND2X2 AND2X2_1304 ( .A(_abc_15724_n2992_bF_buf5), .B(d_reg_22_), .Y(_abc_15724_n3299) );
  AND2X2 AND2X2_1305 ( .A(_abc_15724_n906_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_54_), .Y(_abc_15724_n3300) );
  AND2X2 AND2X2_1306 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n3300), .Y(_abc_15724_n3301) );
  AND2X2 AND2X2_1307 ( .A(c_reg_22_), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n3302) );
  AND2X2 AND2X2_1308 ( .A(_abc_15724_n2992_bF_buf4), .B(d_reg_23_), .Y(_abc_15724_n3305) );
  AND2X2 AND2X2_1309 ( .A(_abc_15724_n906_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_55_), .Y(_abc_15724_n3306) );
  AND2X2 AND2X2_131 ( .A(_abc_15724_n950), .B(_abc_15724_n948), .Y(_abc_15724_n951) );
  AND2X2 AND2X2_1310 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n3306), .Y(_abc_15724_n3307_1) );
  AND2X2 AND2X2_1311 ( .A(c_reg_23_), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n3308) );
  AND2X2 AND2X2_1312 ( .A(_abc_15724_n2992_bF_buf3), .B(d_reg_24_), .Y(_abc_15724_n3311_1) );
  AND2X2 AND2X2_1313 ( .A(_abc_15724_n906_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_56_), .Y(_abc_15724_n3312) );
  AND2X2 AND2X2_1314 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n3312), .Y(_abc_15724_n3313) );
  AND2X2 AND2X2_1315 ( .A(c_reg_24_), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n3314) );
  AND2X2 AND2X2_1316 ( .A(_abc_15724_n2992_bF_buf2), .B(d_reg_25_), .Y(_abc_15724_n3317) );
  AND2X2 AND2X2_1317 ( .A(_abc_15724_n906_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_57_), .Y(_abc_15724_n3318) );
  AND2X2 AND2X2_1318 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n3318), .Y(_abc_15724_n3319) );
  AND2X2 AND2X2_1319 ( .A(c_reg_25_), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n3320) );
  AND2X2 AND2X2_132 ( .A(_abc_15724_n951), .B(digest_update_bF_buf4), .Y(_abc_15724_n952) );
  AND2X2 AND2X2_1320 ( .A(_abc_15724_n2992_bF_buf1), .B(d_reg_26_), .Y(_abc_15724_n3323) );
  AND2X2 AND2X2_1321 ( .A(_abc_15724_n906_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_58_), .Y(_abc_15724_n3324) );
  AND2X2 AND2X2_1322 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n3324), .Y(_abc_15724_n3325) );
  AND2X2 AND2X2_1323 ( .A(c_reg_26_), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n3326) );
  AND2X2 AND2X2_1324 ( .A(_abc_15724_n2992_bF_buf0), .B(d_reg_27_), .Y(_abc_15724_n3329) );
  AND2X2 AND2X2_1325 ( .A(_abc_15724_n906_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_59_), .Y(_abc_15724_n3330) );
  AND2X2 AND2X2_1326 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n3330), .Y(_abc_15724_n3331) );
  AND2X2 AND2X2_1327 ( .A(c_reg_27_), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n3332) );
  AND2X2 AND2X2_1328 ( .A(_abc_15724_n2992_bF_buf11), .B(d_reg_28_), .Y(_abc_15724_n3335) );
  AND2X2 AND2X2_1329 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n1461), .Y(_abc_15724_n3336) );
  AND2X2 AND2X2_133 ( .A(_abc_15724_n906_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_29_), .Y(_abc_15724_n954_1) );
  AND2X2 AND2X2_1330 ( .A(c_reg_28_), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n3337) );
  AND2X2 AND2X2_1331 ( .A(_abc_15724_n2992_bF_buf10), .B(d_reg_29_), .Y(_abc_15724_n3340) );
  AND2X2 AND2X2_1332 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n1464_1), .Y(_abc_15724_n3341) );
  AND2X2 AND2X2_1333 ( .A(c_reg_29_), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n3342) );
  AND2X2 AND2X2_1334 ( .A(_abc_15724_n2992_bF_buf9), .B(d_reg_30_), .Y(_abc_15724_n3345) );
  AND2X2 AND2X2_1335 ( .A(_abc_15724_n906_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_62_), .Y(_abc_15724_n3346) );
  AND2X2 AND2X2_1336 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n3346), .Y(_abc_15724_n3347) );
  AND2X2 AND2X2_1337 ( .A(c_reg_30_), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n3348) );
  AND2X2 AND2X2_1338 ( .A(_abc_15724_n2992_bF_buf8), .B(d_reg_31_), .Y(_abc_15724_n3351) );
  AND2X2 AND2X2_1339 ( .A(_abc_15724_n906_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_63_), .Y(_abc_15724_n3352_1) );
  AND2X2 AND2X2_134 ( .A(_abc_15724_n950), .B(_abc_15724_n946), .Y(_abc_15724_n956_1) );
  AND2X2 AND2X2_1340 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n3352_1), .Y(_abc_15724_n3353) );
  AND2X2 AND2X2_1341 ( .A(c_reg_31_), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n3354) );
  AND2X2 AND2X2_1342 ( .A(_abc_15724_n2992_bF_buf7), .B(c_reg_0_), .Y(_abc_15724_n3357) );
  AND2X2 AND2X2_1343 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n1514), .Y(_abc_15724_n3358) );
  AND2X2 AND2X2_1344 ( .A(b_reg_2_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n3359) );
  AND2X2 AND2X2_1345 ( .A(_abc_15724_n2992_bF_buf6), .B(c_reg_1_), .Y(_abc_15724_n3362) );
  AND2X2 AND2X2_1346 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n1526), .Y(_abc_15724_n3363) );
  AND2X2 AND2X2_1347 ( .A(b_reg_3_), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n3364) );
  AND2X2 AND2X2_1348 ( .A(_abc_15724_n2992_bF_buf5), .B(c_reg_2_), .Y(_abc_15724_n3367) );
  AND2X2 AND2X2_1349 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n1540_1), .Y(_abc_15724_n3368) );
  AND2X2 AND2X2_135 ( .A(_auto_iopadmap_cc_313_execute_26059_29_), .B(e_reg_29_), .Y(_abc_15724_n959) );
  AND2X2 AND2X2_1350 ( .A(b_reg_4_), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n3369) );
  AND2X2 AND2X2_1351 ( .A(_abc_15724_n2992_bF_buf4), .B(c_reg_3_), .Y(_abc_15724_n3372) );
  AND2X2 AND2X2_1352 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n1554), .Y(_abc_15724_n3373) );
  AND2X2 AND2X2_1353 ( .A(b_reg_5_), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n3374) );
  AND2X2 AND2X2_1354 ( .A(_abc_15724_n2992_bF_buf3), .B(c_reg_4_), .Y(_abc_15724_n3377) );
  AND2X2 AND2X2_1355 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n1570_1), .Y(_abc_15724_n3378) );
  AND2X2 AND2X2_1356 ( .A(b_reg_6_), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n3379) );
  AND2X2 AND2X2_1357 ( .A(_abc_15724_n2992_bF_buf2), .B(c_reg_5_), .Y(_abc_15724_n3382) );
  AND2X2 AND2X2_1358 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n1584_1), .Y(_abc_15724_n3383) );
  AND2X2 AND2X2_1359 ( .A(b_reg_7_), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n3384) );
  AND2X2 AND2X2_136 ( .A(_abc_15724_n960), .B(_abc_15724_n958), .Y(_abc_15724_n961) );
  AND2X2 AND2X2_1360 ( .A(_abc_15724_n2992_bF_buf1), .B(c_reg_6_), .Y(_abc_15724_n3387) );
  AND2X2 AND2X2_1361 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n1598), .Y(_abc_15724_n3388) );
  AND2X2 AND2X2_1362 ( .A(b_reg_8_), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n3389_1) );
  AND2X2 AND2X2_1363 ( .A(_abc_15724_n2992_bF_buf0), .B(c_reg_7_), .Y(_abc_15724_n3392) );
  AND2X2 AND2X2_1364 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n1612), .Y(_abc_15724_n3393) );
  AND2X2 AND2X2_1365 ( .A(b_reg_9_), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n3394) );
  AND2X2 AND2X2_1366 ( .A(_abc_15724_n2992_bF_buf11), .B(c_reg_8_), .Y(_abc_15724_n3397) );
  AND2X2 AND2X2_1367 ( .A(_abc_15724_n906_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_72_), .Y(_abc_15724_n3398) );
  AND2X2 AND2X2_1368 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n3398), .Y(_abc_15724_n3399) );
  AND2X2 AND2X2_1369 ( .A(b_reg_10_), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n3400) );
  AND2X2 AND2X2_137 ( .A(_abc_15724_n962), .B(_abc_15724_n964), .Y(_abc_15724_n965) );
  AND2X2 AND2X2_1370 ( .A(_abc_15724_n2992_bF_buf10), .B(c_reg_9_), .Y(_abc_15724_n3403) );
  AND2X2 AND2X2_1371 ( .A(_abc_15724_n906_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_73_), .Y(_abc_15724_n3404) );
  AND2X2 AND2X2_1372 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n3404), .Y(_abc_15724_n3405) );
  AND2X2 AND2X2_1373 ( .A(b_reg_11_), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n3406) );
  AND2X2 AND2X2_1374 ( .A(_abc_15724_n2992_bF_buf9), .B(c_reg_10_), .Y(_abc_15724_n3409) );
  AND2X2 AND2X2_1375 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n1655_1), .Y(_abc_15724_n3410) );
  AND2X2 AND2X2_1376 ( .A(b_reg_12_), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n3411) );
  AND2X2 AND2X2_1377 ( .A(_abc_15724_n2992_bF_buf8), .B(c_reg_11_), .Y(_abc_15724_n3414) );
  AND2X2 AND2X2_1378 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n1669_1), .Y(_abc_15724_n3415) );
  AND2X2 AND2X2_1379 ( .A(b_reg_13_), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n3416) );
  AND2X2 AND2X2_138 ( .A(_abc_15724_n966_1), .B(_abc_15724_n955), .Y(H4_reg_29__FF_INPUT) );
  AND2X2 AND2X2_1380 ( .A(_abc_15724_n2992_bF_buf7), .B(c_reg_12_), .Y(_abc_15724_n3419) );
  AND2X2 AND2X2_1381 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n1695), .Y(_abc_15724_n3420) );
  AND2X2 AND2X2_1382 ( .A(b_reg_14_), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n3421) );
  AND2X2 AND2X2_1383 ( .A(_abc_15724_n2992_bF_buf6), .B(c_reg_13_), .Y(_abc_15724_n3424) );
  AND2X2 AND2X2_1384 ( .A(_abc_15724_n906_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_77_), .Y(_abc_15724_n3425_1) );
  AND2X2 AND2X2_1385 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n3425_1), .Y(_abc_15724_n3426) );
  AND2X2 AND2X2_1386 ( .A(b_reg_15_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n3427) );
  AND2X2 AND2X2_1387 ( .A(_abc_15724_n2992_bF_buf5), .B(c_reg_14_), .Y(_abc_15724_n3430) );
  AND2X2 AND2X2_1388 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n1722), .Y(_abc_15724_n3431) );
  AND2X2 AND2X2_1389 ( .A(b_reg_16_), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n3432) );
  AND2X2 AND2X2_139 ( .A(e_reg_30_), .B(_auto_iopadmap_cc_313_execute_26059_30_), .Y(_abc_15724_n969) );
  AND2X2 AND2X2_1390 ( .A(_abc_15724_n2992_bF_buf4), .B(c_reg_15_), .Y(_abc_15724_n3435) );
  AND2X2 AND2X2_1391 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n1736), .Y(_abc_15724_n3436) );
  AND2X2 AND2X2_1392 ( .A(b_reg_17_), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n3437) );
  AND2X2 AND2X2_1393 ( .A(_abc_15724_n2992_bF_buf3), .B(c_reg_16_), .Y(_abc_15724_n3440) );
  AND2X2 AND2X2_1394 ( .A(_abc_15724_n906_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_80_), .Y(_abc_15724_n3441) );
  AND2X2 AND2X2_1395 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n3441), .Y(_abc_15724_n3442) );
  AND2X2 AND2X2_1396 ( .A(b_reg_18_), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n3443) );
  AND2X2 AND2X2_1397 ( .A(_abc_15724_n2992_bF_buf2), .B(c_reg_17_), .Y(_abc_15724_n3446) );
  AND2X2 AND2X2_1398 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n1775), .Y(_abc_15724_n3447) );
  AND2X2 AND2X2_1399 ( .A(b_reg_19_), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n3448) );
  AND2X2 AND2X2_14 ( .A(_abc_15724_n723), .B(_abc_15724_n713), .Y(_abc_15724_n724) );
  AND2X2 AND2X2_140 ( .A(_abc_15724_n970), .B(_abc_15724_n968_1), .Y(_abc_15724_n971) );
  AND2X2 AND2X2_1400 ( .A(_abc_15724_n2992_bF_buf1), .B(c_reg_18_), .Y(_abc_15724_n3451) );
  AND2X2 AND2X2_1401 ( .A(_abc_15724_n906_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_82_), .Y(_abc_15724_n3452) );
  AND2X2 AND2X2_1402 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n3452), .Y(_abc_15724_n3453) );
  AND2X2 AND2X2_1403 ( .A(b_reg_20_), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n3454) );
  AND2X2 AND2X2_1404 ( .A(_abc_15724_n2992_bF_buf0), .B(c_reg_19_), .Y(_abc_15724_n3457) );
  AND2X2 AND2X2_1405 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n1806), .Y(_abc_15724_n3458) );
  AND2X2 AND2X2_1406 ( .A(b_reg_21_), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n3459) );
  AND2X2 AND2X2_1407 ( .A(_abc_15724_n2992_bF_buf11), .B(c_reg_20_), .Y(_abc_15724_n3462) );
  AND2X2 AND2X2_1408 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n1829), .Y(_abc_15724_n3463) );
  AND2X2 AND2X2_1409 ( .A(b_reg_22_), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n3464) );
  AND2X2 AND2X2_141 ( .A(_abc_15724_n961), .B(_abc_15724_n945_1), .Y(_abc_15724_n972) );
  AND2X2 AND2X2_1410 ( .A(_abc_15724_n2992_bF_buf10), .B(c_reg_21_), .Y(_abc_15724_n3467) );
  AND2X2 AND2X2_1411 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n1843), .Y(_abc_15724_n3468_1) );
  AND2X2 AND2X2_1412 ( .A(b_reg_23_), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n3469_1) );
  AND2X2 AND2X2_1413 ( .A(_abc_15724_n2992_bF_buf9), .B(c_reg_22_), .Y(_abc_15724_n3472) );
  AND2X2 AND2X2_1414 ( .A(_abc_15724_n906_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_86_), .Y(_abc_15724_n3473) );
  AND2X2 AND2X2_1415 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n3473), .Y(_abc_15724_n3474) );
  AND2X2 AND2X2_1416 ( .A(b_reg_24_), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n3475) );
  AND2X2 AND2X2_1417 ( .A(_abc_15724_n2992_bF_buf8), .B(c_reg_23_), .Y(_abc_15724_n3478) );
  AND2X2 AND2X2_1418 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n1874), .Y(_abc_15724_n3479) );
  AND2X2 AND2X2_1419 ( .A(b_reg_25_), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n3480) );
  AND2X2 AND2X2_142 ( .A(_abc_15724_n947), .B(_abc_15724_n961), .Y(_abc_15724_n974) );
  AND2X2 AND2X2_1420 ( .A(_abc_15724_n2992_bF_buf7), .B(c_reg_24_), .Y(_abc_15724_n3483_1) );
  AND2X2 AND2X2_1421 ( .A(_abc_15724_n906_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_88_), .Y(_abc_15724_n3484) );
  AND2X2 AND2X2_1422 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n3484), .Y(_abc_15724_n3485) );
  AND2X2 AND2X2_1423 ( .A(b_reg_26_), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n3486) );
  AND2X2 AND2X2_1424 ( .A(_abc_15724_n2992_bF_buf6), .B(c_reg_25_), .Y(_abc_15724_n3489_1) );
  AND2X2 AND2X2_1425 ( .A(_abc_15724_n906_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_89_), .Y(_abc_15724_n3490) );
  AND2X2 AND2X2_1426 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n3490), .Y(_abc_15724_n3491_1) );
  AND2X2 AND2X2_1427 ( .A(b_reg_27_), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n3492_1) );
  AND2X2 AND2X2_1428 ( .A(_abc_15724_n2992_bF_buf5), .B(c_reg_26_), .Y(_abc_15724_n3495) );
  AND2X2 AND2X2_1429 ( .A(_abc_15724_n906_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_90_), .Y(_abc_15724_n3496) );
  AND2X2 AND2X2_143 ( .A(_abc_15724_n943_1), .B(_abc_15724_n974), .Y(_abc_15724_n975) );
  AND2X2 AND2X2_1430 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n3496), .Y(_abc_15724_n3497_1) );
  AND2X2 AND2X2_1431 ( .A(b_reg_28_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n3498) );
  AND2X2 AND2X2_1432 ( .A(_abc_15724_n2992_bF_buf4), .B(c_reg_27_), .Y(_abc_15724_n3501_1) );
  AND2X2 AND2X2_1433 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n1940_1), .Y(_abc_15724_n3502) );
  AND2X2 AND2X2_1434 ( .A(b_reg_29_), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n3503) );
  AND2X2 AND2X2_1435 ( .A(_abc_15724_n2992_bF_buf3), .B(c_reg_28_), .Y(_abc_15724_n3506) );
  AND2X2 AND2X2_1436 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n1964), .Y(_abc_15724_n3507_1) );
  AND2X2 AND2X2_1437 ( .A(b_reg_30_), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n3508) );
  AND2X2 AND2X2_1438 ( .A(_abc_15724_n2992_bF_buf2), .B(c_reg_29_), .Y(_abc_15724_n3511) );
  AND2X2 AND2X2_1439 ( .A(_abc_15724_n906_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_93_), .Y(_abc_15724_n3512) );
  AND2X2 AND2X2_144 ( .A(_abc_15724_n976_1), .B(_abc_15724_n971), .Y(_abc_15724_n978) );
  AND2X2 AND2X2_1440 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n3512), .Y(_abc_15724_n3513_1) );
  AND2X2 AND2X2_1441 ( .A(b_reg_31_), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n3514_1) );
  AND2X2 AND2X2_1442 ( .A(_abc_15724_n2992_bF_buf1), .B(c_reg_30_), .Y(_abc_15724_n3517_1) );
  AND2X2 AND2X2_1443 ( .A(_abc_15724_n906_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_94_), .Y(_abc_15724_n3518) );
  AND2X2 AND2X2_1444 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n3518), .Y(_abc_15724_n3519) );
  AND2X2 AND2X2_1445 ( .A(b_reg_0_), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n3520) );
  AND2X2 AND2X2_1446 ( .A(_abc_15724_n2992_bF_buf0), .B(c_reg_31_), .Y(_abc_15724_n3523) );
  AND2X2 AND2X2_1447 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n2011_1), .Y(_abc_15724_n3524) );
  AND2X2 AND2X2_1448 ( .A(b_reg_1_), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n3525) );
  AND2X2 AND2X2_1449 ( .A(_abc_15724_n2992_bF_buf11), .B(b_reg_0_), .Y(_abc_15724_n3528_1) );
  AND2X2 AND2X2_145 ( .A(_abc_15724_n979_1), .B(_abc_15724_n977_1), .Y(_abc_15724_n980) );
  AND2X2 AND2X2_1450 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n2019), .Y(_abc_15724_n3529_1) );
  AND2X2 AND2X2_1451 ( .A(a_reg_0_), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n3530) );
  AND2X2 AND2X2_1452 ( .A(_abc_15724_n2992_bF_buf10), .B(b_reg_1_), .Y(_abc_15724_n3533) );
  AND2X2 AND2X2_1453 ( .A(_abc_15724_n906_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_97_), .Y(_abc_15724_n3534) );
  AND2X2 AND2X2_1454 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n3534), .Y(_abc_15724_n3535_1) );
  AND2X2 AND2X2_1455 ( .A(a_reg_1_), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n3536) );
  AND2X2 AND2X2_1456 ( .A(_abc_15724_n2992_bF_buf9), .B(b_reg_2_), .Y(_abc_15724_n3539) );
  AND2X2 AND2X2_1457 ( .A(_abc_15724_n906_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_98_), .Y(_abc_15724_n3540) );
  AND2X2 AND2X2_1458 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n3540), .Y(_abc_15724_n3541) );
  AND2X2 AND2X2_1459 ( .A(a_reg_2_), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n3542) );
  AND2X2 AND2X2_146 ( .A(_abc_15724_n980), .B(digest_update_bF_buf2), .Y(_abc_15724_n981) );
  AND2X2 AND2X2_1460 ( .A(_abc_15724_n2992_bF_buf8), .B(b_reg_3_), .Y(_abc_15724_n3545) );
  AND2X2 AND2X2_1461 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n2057_1), .Y(_abc_15724_n3546_1) );
  AND2X2 AND2X2_1462 ( .A(a_reg_3_), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n3547) );
  AND2X2 AND2X2_1463 ( .A(_abc_15724_n2992_bF_buf7), .B(b_reg_4_), .Y(_abc_15724_n3550) );
  AND2X2 AND2X2_1464 ( .A(_abc_15724_n906_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_100_), .Y(_abc_15724_n3551) );
  AND2X2 AND2X2_1465 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n3551), .Y(_abc_15724_n3552) );
  AND2X2 AND2X2_1466 ( .A(a_reg_4_), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n3553) );
  AND2X2 AND2X2_1467 ( .A(_abc_15724_n2992_bF_buf6), .B(b_reg_5_), .Y(_abc_15724_n3556) );
  AND2X2 AND2X2_1468 ( .A(_abc_15724_n906_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_101_), .Y(_abc_15724_n3557) );
  AND2X2 AND2X2_1469 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n3557), .Y(_abc_15724_n3558) );
  AND2X2 AND2X2_147 ( .A(_abc_15724_n982), .B(_abc_15724_n850_bF_buf2), .Y(_abc_15724_n983) );
  AND2X2 AND2X2_1470 ( .A(a_reg_5_), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n3559) );
  AND2X2 AND2X2_1471 ( .A(_abc_15724_n2992_bF_buf5), .B(b_reg_6_), .Y(_abc_15724_n3562) );
  AND2X2 AND2X2_1472 ( .A(_abc_15724_n906_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_102_), .Y(_abc_15724_n3563) );
  AND2X2 AND2X2_1473 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n3563), .Y(_abc_15724_n3564_1) );
  AND2X2 AND2X2_1474 ( .A(a_reg_6_), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n3565) );
  AND2X2 AND2X2_1475 ( .A(_abc_15724_n2992_bF_buf4), .B(b_reg_7_), .Y(_abc_15724_n3568) );
  AND2X2 AND2X2_1476 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n2097), .Y(_abc_15724_n3569) );
  AND2X2 AND2X2_1477 ( .A(a_reg_7_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n3570) );
  AND2X2 AND2X2_1478 ( .A(_abc_15724_n2992_bF_buf3), .B(b_reg_8_), .Y(_abc_15724_n3573) );
  AND2X2 AND2X2_1479 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n2122), .Y(_abc_15724_n3574) );
  AND2X2 AND2X2_148 ( .A(_abc_15724_n987_1), .B(_abc_15724_n989_1), .Y(_abc_15724_n990) );
  AND2X2 AND2X2_1480 ( .A(a_reg_8_), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n3575) );
  AND2X2 AND2X2_1481 ( .A(_abc_15724_n2992_bF_buf2), .B(b_reg_9_), .Y(_abc_15724_n3578) );
  AND2X2 AND2X2_1482 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n2136), .Y(_abc_15724_n3579) );
  AND2X2 AND2X2_1483 ( .A(a_reg_9_), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n3580) );
  AND2X2 AND2X2_1484 ( .A(_abc_15724_n2992_bF_buf1), .B(b_reg_10_), .Y(_abc_15724_n3583) );
  AND2X2 AND2X2_1485 ( .A(_abc_15724_n906_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_106_), .Y(_abc_15724_n3584_1) );
  AND2X2 AND2X2_1486 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n3584_1), .Y(_abc_15724_n3585_1) );
  AND2X2 AND2X2_1487 ( .A(a_reg_10_), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n3586) );
  AND2X2 AND2X2_1488 ( .A(_abc_15724_n2992_bF_buf0), .B(b_reg_11_), .Y(_abc_15724_n3589) );
  AND2X2 AND2X2_1489 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n2167), .Y(_abc_15724_n3590) );
  AND2X2 AND2X2_149 ( .A(_abc_15724_n994), .B(_abc_15724_n992), .Y(_abc_15724_n995) );
  AND2X2 AND2X2_1490 ( .A(a_reg_11_), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n3591_1) );
  AND2X2 AND2X2_1491 ( .A(_abc_15724_n2992_bF_buf11), .B(b_reg_12_), .Y(_abc_15724_n3594) );
  AND2X2 AND2X2_1492 ( .A(_abc_15724_n906_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_108_), .Y(_abc_15724_n3595) );
  AND2X2 AND2X2_1493 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n3595), .Y(_abc_15724_n3596) );
  AND2X2 AND2X2_1494 ( .A(a_reg_12_), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n3597) );
  AND2X2 AND2X2_1495 ( .A(_abc_15724_n2992_bF_buf10), .B(b_reg_13_), .Y(_abc_15724_n3600) );
  AND2X2 AND2X2_1496 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n2200), .Y(_abc_15724_n3601) );
  AND2X2 AND2X2_1497 ( .A(a_reg_13_), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n3602_1) );
  AND2X2 AND2X2_1498 ( .A(_abc_15724_n2992_bF_buf9), .B(b_reg_14_), .Y(_abc_15724_n3605) );
  AND2X2 AND2X2_1499 ( .A(_abc_15724_n906_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_110_), .Y(_abc_15724_n3606) );
  AND2X2 AND2X2_15 ( .A(_abc_15724_n707), .B(_abc_15724_n709_1), .Y(_abc_15724_n725) );
  AND2X2 AND2X2_150 ( .A(_abc_15724_n995), .B(digest_update_bF_buf1), .Y(_abc_15724_n996_1) );
  AND2X2 AND2X2_1500 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n3606), .Y(_abc_15724_n3607) );
  AND2X2 AND2X2_1501 ( .A(a_reg_14_), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n3608) );
  AND2X2 AND2X2_1502 ( .A(_abc_15724_n2992_bF_buf8), .B(b_reg_15_), .Y(_abc_15724_n3611) );
  AND2X2 AND2X2_1503 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n2231), .Y(_abc_15724_n3612) );
  AND2X2 AND2X2_1504 ( .A(a_reg_15_), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n3613) );
  AND2X2 AND2X2_1505 ( .A(_abc_15724_n2992_bF_buf7), .B(b_reg_16_), .Y(_abc_15724_n3616) );
  AND2X2 AND2X2_1506 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n2251), .Y(_abc_15724_n3617) );
  AND2X2 AND2X2_1507 ( .A(a_reg_16_), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n3618) );
  AND2X2 AND2X2_1508 ( .A(_abc_15724_n2992_bF_buf6), .B(b_reg_17_), .Y(_abc_15724_n3621_1) );
  AND2X2 AND2X2_1509 ( .A(_abc_15724_n906_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_113_), .Y(_abc_15724_n3622) );
  AND2X2 AND2X2_151 ( .A(_abc_15724_n997_1), .B(_abc_15724_n850_bF_buf1), .Y(_abc_15724_n998_1) );
  AND2X2 AND2X2_1510 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n3622), .Y(_abc_15724_n3623) );
  AND2X2 AND2X2_1511 ( .A(a_reg_17_), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n3624) );
  AND2X2 AND2X2_1512 ( .A(_abc_15724_n2992_bF_buf5), .B(b_reg_18_), .Y(_abc_15724_n3627) );
  AND2X2 AND2X2_1513 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n2278), .Y(_abc_15724_n3628) );
  AND2X2 AND2X2_1514 ( .A(a_reg_18_), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n3629_1) );
  AND2X2 AND2X2_1515 ( .A(_abc_15724_n2992_bF_buf4), .B(b_reg_19_), .Y(_abc_15724_n3632) );
  AND2X2 AND2X2_1516 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n2292), .Y(_abc_15724_n3633) );
  AND2X2 AND2X2_1517 ( .A(a_reg_19_), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n3634) );
  AND2X2 AND2X2_1518 ( .A(_abc_15724_n2992_bF_buf3), .B(b_reg_20_), .Y(_abc_15724_n3637) );
  AND2X2 AND2X2_1519 ( .A(_abc_15724_n906_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_116_), .Y(_abc_15724_n3638) );
  AND2X2 AND2X2_152 ( .A(_auto_iopadmap_cc_313_execute_26059_32_), .B(d_reg_0_), .Y(_abc_15724_n1001) );
  AND2X2 AND2X2_1520 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n3638), .Y(_abc_15724_n3639_1) );
  AND2X2 AND2X2_1521 ( .A(a_reg_20_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n3640) );
  AND2X2 AND2X2_1522 ( .A(_abc_15724_n2992_bF_buf2), .B(b_reg_21_), .Y(_abc_15724_n3643) );
  AND2X2 AND2X2_1523 ( .A(_abc_15724_n906_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_117_), .Y(_abc_15724_n3644) );
  AND2X2 AND2X2_1524 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n3644), .Y(_abc_15724_n3645_1) );
  AND2X2 AND2X2_1525 ( .A(a_reg_21_), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n3646_1) );
  AND2X2 AND2X2_1526 ( .A(_abc_15724_n2992_bF_buf1), .B(b_reg_22_), .Y(_abc_15724_n3649) );
  AND2X2 AND2X2_1527 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n2339), .Y(_abc_15724_n3650) );
  AND2X2 AND2X2_1528 ( .A(a_reg_22_), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n3651) );
  AND2X2 AND2X2_1529 ( .A(_abc_15724_n2992_bF_buf0), .B(b_reg_23_), .Y(_abc_15724_n3654) );
  AND2X2 AND2X2_153 ( .A(_abc_15724_n1002), .B(_abc_15724_n1000), .Y(_abc_15724_n1003) );
  AND2X2 AND2X2_1530 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n2353), .Y(_abc_15724_n3655) );
  AND2X2 AND2X2_1531 ( .A(a_reg_23_), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n3656) );
  AND2X2 AND2X2_1532 ( .A(_abc_15724_n2992_bF_buf11), .B(b_reg_24_), .Y(_abc_15724_n3659) );
  AND2X2 AND2X2_1533 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n2379), .Y(_abc_15724_n3660) );
  AND2X2 AND2X2_1534 ( .A(a_reg_24_), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n3661) );
  AND2X2 AND2X2_1535 ( .A(_abc_15724_n2992_bF_buf10), .B(b_reg_25_), .Y(_abc_15724_n3664) );
  AND2X2 AND2X2_1536 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n2393), .Y(_abc_15724_n3665) );
  AND2X2 AND2X2_1537 ( .A(a_reg_25_), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n3666) );
  AND2X2 AND2X2_1538 ( .A(_abc_15724_n2992_bF_buf9), .B(b_reg_26_), .Y(_abc_15724_n3669) );
  AND2X2 AND2X2_1539 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n2410), .Y(_abc_15724_n3670_1) );
  AND2X2 AND2X2_154 ( .A(_abc_15724_n906_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_32_), .Y(_abc_15724_n1005) );
  AND2X2 AND2X2_1540 ( .A(a_reg_26_), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n3671_1) );
  AND2X2 AND2X2_1541 ( .A(_abc_15724_n2992_bF_buf8), .B(b_reg_27_), .Y(_abc_15724_n3674) );
  AND2X2 AND2X2_1542 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n2424), .Y(_abc_15724_n3675) );
  AND2X2 AND2X2_1543 ( .A(a_reg_27_), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n3676) );
  AND2X2 AND2X2_1544 ( .A(_abc_15724_n2992_bF_buf7), .B(b_reg_28_), .Y(_abc_15724_n3679_1) );
  AND2X2 AND2X2_1545 ( .A(_abc_15724_n906_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_124_), .Y(_abc_15724_n3680_1) );
  AND2X2 AND2X2_1546 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n3680_1), .Y(_abc_15724_n3681) );
  AND2X2 AND2X2_1547 ( .A(a_reg_28_), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n3682) );
  AND2X2 AND2X2_1548 ( .A(_abc_15724_n2992_bF_buf6), .B(b_reg_29_), .Y(_abc_15724_n3685) );
  AND2X2 AND2X2_1549 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n2457), .Y(_abc_15724_n3686_1) );
  AND2X2 AND2X2_155 ( .A(_abc_15724_n1004), .B(_abc_15724_n1006), .Y(H3_reg_0__FF_INPUT) );
  AND2X2 AND2X2_1550 ( .A(a_reg_29_), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n3687) );
  AND2X2 AND2X2_1551 ( .A(_abc_15724_n2992_bF_buf5), .B(b_reg_30_), .Y(_abc_15724_n3690) );
  AND2X2 AND2X2_1552 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n2474), .Y(_abc_15724_n3691) );
  AND2X2 AND2X2_1553 ( .A(a_reg_30_), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n3692) );
  AND2X2 AND2X2_1554 ( .A(_abc_15724_n2992_bF_buf4), .B(b_reg_31_), .Y(_abc_15724_n3695) );
  AND2X2 AND2X2_1555 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n2489), .Y(_abc_15724_n3696) );
  AND2X2 AND2X2_1556 ( .A(a_reg_31_), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n3697) );
  AND2X2 AND2X2_1557 ( .A(round_ctr_reg_5_), .B(round_ctr_reg_4_), .Y(_abc_15724_n3700) );
  AND2X2 AND2X2_1558 ( .A(round_ctr_reg_3_), .B(round_ctr_reg_5_), .Y(_abc_15724_n3703) );
  AND2X2 AND2X2_1559 ( .A(_abc_15724_n3704), .B(_abc_15724_n3702), .Y(_abc_15724_n3705) );
  AND2X2 AND2X2_156 ( .A(_abc_15724_n1008), .B(_abc_15724_n1009), .Y(_abc_15724_n1010) );
  AND2X2 AND2X2_1560 ( .A(_abc_15724_n3705), .B(_abc_15724_n3701), .Y(_abc_15724_n3706) );
  AND2X2 AND2X2_1561 ( .A(c_reg_0_), .B(b_reg_0_), .Y(_abc_15724_n3708) );
  AND2X2 AND2X2_1562 ( .A(_abc_15724_n3709), .B(_abc_15724_n3710), .Y(_abc_15724_n3711) );
  AND2X2 AND2X2_1563 ( .A(_abc_15724_n3713), .B(_abc_15724_n3707), .Y(_abc_15724_n3714) );
  AND2X2 AND2X2_1564 ( .A(_abc_15724_n3712), .B(d_reg_0_), .Y(_abc_15724_n3715) );
  AND2X2 AND2X2_1565 ( .A(round_ctr_reg_2_), .B(round_ctr_reg_4_), .Y(_abc_15724_n3717) );
  AND2X2 AND2X2_1566 ( .A(round_ctr_reg_3_), .B(round_ctr_reg_4_), .Y(_abc_15724_n3719) );
  AND2X2 AND2X2_1567 ( .A(round_ctr_reg_2_), .B(round_ctr_reg_3_), .Y(_abc_15724_n3722) );
  AND2X2 AND2X2_1568 ( .A(_abc_15724_n3700), .B(_abc_15724_n3722), .Y(_abc_15724_n3723) );
  AND2X2 AND2X2_1569 ( .A(_abc_15724_n3725_bF_buf3), .B(_abc_15724_n3721_bF_buf4), .Y(_abc_15724_n3726) );
  AND2X2 AND2X2_157 ( .A(_auto_iopadmap_cc_313_execute_26059_33_), .B(d_reg_1_), .Y(_abc_15724_n1011) );
  AND2X2 AND2X2_1570 ( .A(_abc_15724_n3726_bF_buf4), .B(_abc_15724_n3716), .Y(_abc_15724_n3727) );
  AND2X2 AND2X2_1571 ( .A(_abc_15724_n3709), .B(b_reg_0_), .Y(_abc_15724_n3729) );
  AND2X2 AND2X2_1572 ( .A(_abc_15724_n3707), .B(_abc_15724_n3710), .Y(_abc_15724_n3730) );
  AND2X2 AND2X2_1573 ( .A(_abc_15724_n3735), .B(_abc_15724_n3702), .Y(_abc_15724_n3736) );
  AND2X2 AND2X2_1574 ( .A(_abc_15724_n3736), .B(_abc_15724_n3734), .Y(_abc_15724_n3737) );
  AND2X2 AND2X2_1575 ( .A(_abc_15724_n3738), .B(_abc_15724_n3739), .Y(_abc_15724_n3740) );
  AND2X2 AND2X2_1576 ( .A(_abc_15724_n3737_bF_buf4), .B(_abc_15724_n3740), .Y(_abc_15724_n3741) );
  AND2X2 AND2X2_1577 ( .A(_abc_15724_n3742), .B(_abc_15724_n3732), .Y(_abc_15724_n3743) );
  AND2X2 AND2X2_1578 ( .A(_abc_15724_n3728), .B(_abc_15724_n3743), .Y(_abc_15724_n3744) );
  AND2X2 AND2X2_1579 ( .A(a_reg_27_), .B(e_reg_0_), .Y(_abc_15724_n3747) );
  AND2X2 AND2X2_158 ( .A(_abc_15724_n1015_1), .B(_abc_15724_n1014), .Y(_abc_15724_n1016_1) );
  AND2X2 AND2X2_1580 ( .A(_abc_15724_n3748), .B(_abc_15724_n3746), .Y(_abc_15724_n3749) );
  AND2X2 AND2X2_1581 ( .A(_abc_15724_n3749), .B(w_0_), .Y(_abc_15724_n3750) );
  AND2X2 AND2X2_1582 ( .A(_abc_15724_n3752), .B(_abc_15724_n3751), .Y(_abc_15724_n3753) );
  AND2X2 AND2X2_1583 ( .A(_abc_15724_n3745), .B(_abc_15724_n3755), .Y(_abc_15724_n3756) );
  AND2X2 AND2X2_1584 ( .A(_abc_15724_n3744), .B(_abc_15724_n3754), .Y(_abc_15724_n3757) );
  AND2X2 AND2X2_1585 ( .A(_abc_15724_n3759), .B(_abc_15724_n3706), .Y(_abc_15724_n3761) );
  AND2X2 AND2X2_1586 ( .A(_abc_15724_n3762), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n3763) );
  AND2X2 AND2X2_1587 ( .A(_abc_15724_n3763), .B(_abc_15724_n3760), .Y(_abc_15724_n3764) );
  AND2X2 AND2X2_1588 ( .A(_abc_15724_n2992_bF_buf3), .B(a_reg_0_), .Y(_abc_15724_n3765) );
  AND2X2 AND2X2_1589 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n2497), .Y(_abc_15724_n3766) );
  AND2X2 AND2X2_159 ( .A(_abc_15724_n1013), .B(_abc_15724_n1017), .Y(_abc_15724_n1018_1) );
  AND2X2 AND2X2_1590 ( .A(_abc_15724_n3770), .B(_abc_15724_n3771), .Y(_abc_15724_n3772) );
  AND2X2 AND2X2_1591 ( .A(c_reg_1_), .B(b_reg_1_), .Y(_abc_15724_n3773) );
  AND2X2 AND2X2_1592 ( .A(_abc_15724_n3774), .B(_abc_15724_n1009), .Y(_abc_15724_n3776) );
  AND2X2 AND2X2_1593 ( .A(_abc_15724_n3777), .B(_abc_15724_n3775), .Y(_abc_15724_n3778) );
  AND2X2 AND2X2_1594 ( .A(_abc_15724_n3726_bF_buf3), .B(_abc_15724_n3778), .Y(_abc_15724_n3779) );
  AND2X2 AND2X2_1595 ( .A(_abc_15724_n3780), .B(_abc_15724_n1009), .Y(_abc_15724_n3781) );
  AND2X2 AND2X2_1596 ( .A(_abc_15724_n3770), .B(b_reg_1_), .Y(_abc_15724_n3782) );
  AND2X2 AND2X2_1597 ( .A(_abc_15724_n3737_bF_buf3), .B(_abc_15724_n3787), .Y(_abc_15724_n3788) );
  AND2X2 AND2X2_1598 ( .A(a_reg_28_), .B(e_reg_1_), .Y(_abc_15724_n3793) );
  AND2X2 AND2X2_1599 ( .A(_abc_15724_n3794), .B(_abc_15724_n3792), .Y(_abc_15724_n3795) );
  AND2X2 AND2X2_16 ( .A(_auto_iopadmap_cc_313_execute_26059_15_), .B(e_reg_15_), .Y(_abc_15724_n729_1) );
  AND2X2 AND2X2_160 ( .A(_abc_15724_n1019), .B(_abc_15724_n1021), .Y(H3_reg_1__FF_INPUT) );
  AND2X2 AND2X2_1600 ( .A(_abc_15724_n3795), .B(w_1_), .Y(_abc_15724_n3796) );
  AND2X2 AND2X2_1601 ( .A(_abc_15724_n3797), .B(_abc_15724_n3798), .Y(_abc_15724_n3799) );
  AND2X2 AND2X2_1602 ( .A(_abc_15724_n3799), .B(_abc_15724_n3791), .Y(_abc_15724_n3800) );
  AND2X2 AND2X2_1603 ( .A(_abc_15724_n3801), .B(_abc_15724_n3802), .Y(_abc_15724_n3803) );
  AND2X2 AND2X2_1604 ( .A(_abc_15724_n3790), .B(_abc_15724_n3803), .Y(_abc_15724_n3804) );
  AND2X2 AND2X2_1605 ( .A(_abc_15724_n3807), .B(d_reg_1_), .Y(_abc_15724_n3808) );
  AND2X2 AND2X2_1606 ( .A(_abc_15724_n3811), .B(_abc_15724_n3784), .Y(_abc_15724_n3812) );
  AND2X2 AND2X2_1607 ( .A(_abc_15724_n3810), .B(_abc_15724_n3812), .Y(_abc_15724_n3813) );
  AND2X2 AND2X2_1608 ( .A(_abc_15724_n3816), .B(_abc_15724_n3814), .Y(_abc_15724_n3817) );
  AND2X2 AND2X2_1609 ( .A(_abc_15724_n3813), .B(_abc_15724_n3818), .Y(_abc_15724_n3819) );
  AND2X2 AND2X2_161 ( .A(_abc_15724_n1013), .B(_abc_15724_n1015_1), .Y(_abc_15724_n1023) );
  AND2X2 AND2X2_1610 ( .A(_abc_15724_n3823), .B(_abc_15724_n3822), .Y(_abc_15724_n3824) );
  AND2X2 AND2X2_1611 ( .A(_abc_15724_n3821), .B(_abc_15724_n3825), .Y(_abc_15724_n3826) );
  AND2X2 AND2X2_1612 ( .A(_abc_15724_n3826), .B(_abc_15724_n3724), .Y(_abc_15724_n3827) );
  AND2X2 AND2X2_1613 ( .A(_abc_15724_n3828), .B(_abc_15724_n3829), .Y(_abc_15724_n3830) );
  AND2X2 AND2X2_1614 ( .A(_abc_15724_n3830), .B(_abc_15724_n3736), .Y(_abc_15724_n3831) );
  AND2X2 AND2X2_1615 ( .A(_abc_15724_n3835), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n3836) );
  AND2X2 AND2X2_1616 ( .A(_abc_15724_n3836), .B(_abc_15724_n3833), .Y(_abc_15724_n3837) );
  AND2X2 AND2X2_1617 ( .A(_abc_15724_n2992_bF_buf2), .B(a_reg_1_), .Y(_abc_15724_n3838) );
  AND2X2 AND2X2_1618 ( .A(_abc_15724_n906_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_129_), .Y(_abc_15724_n3839) );
  AND2X2 AND2X2_1619 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n3839), .Y(_abc_15724_n3840) );
  AND2X2 AND2X2_162 ( .A(_auto_iopadmap_cc_313_execute_26059_34_), .B(d_reg_2_), .Y(_abc_15724_n1025_1) );
  AND2X2 AND2X2_1620 ( .A(_abc_15724_n3844), .B(_abc_15724_n3821), .Y(_abc_15724_n3845) );
  AND2X2 AND2X2_1621 ( .A(_abc_15724_n3822), .B(_abc_15724_n3801), .Y(_abc_15724_n3846) );
  AND2X2 AND2X2_1622 ( .A(_abc_15724_n3847), .B(_abc_15724_n3848), .Y(_abc_15724_n3849) );
  AND2X2 AND2X2_1623 ( .A(c_reg_2_), .B(b_reg_2_), .Y(_abc_15724_n3850) );
  AND2X2 AND2X2_1624 ( .A(_abc_15724_n3852), .B(d_reg_2_), .Y(_abc_15724_n3853) );
  AND2X2 AND2X2_1625 ( .A(_abc_15724_n3851), .B(_abc_15724_n3854), .Y(_abc_15724_n3855) );
  AND2X2 AND2X2_1626 ( .A(_abc_15724_n3858), .B(_abc_15724_n3854), .Y(_abc_15724_n3859) );
  AND2X2 AND2X2_1627 ( .A(_abc_15724_n3847), .B(b_reg_2_), .Y(_abc_15724_n3860) );
  AND2X2 AND2X2_1628 ( .A(_abc_15724_n3864), .B(_abc_15724_n3862), .Y(_abc_15724_n3865) );
  AND2X2 AND2X2_1629 ( .A(_abc_15724_n3857), .B(_abc_15724_n3865), .Y(_abc_15724_n3866) );
  AND2X2 AND2X2_163 ( .A(_abc_15724_n1026_1), .B(_abc_15724_n1024_1), .Y(_abc_15724_n1027) );
  AND2X2 AND2X2_1630 ( .A(a_reg_29_), .B(e_reg_2_), .Y(_abc_15724_n3869) );
  AND2X2 AND2X2_1631 ( .A(_abc_15724_n3870), .B(_abc_15724_n3868), .Y(_abc_15724_n3871) );
  AND2X2 AND2X2_1632 ( .A(_abc_15724_n3871), .B(w_2_), .Y(_abc_15724_n3872) );
  AND2X2 AND2X2_1633 ( .A(_abc_15724_n3873), .B(_abc_15724_n3874), .Y(_abc_15724_n3875) );
  AND2X2 AND2X2_1634 ( .A(_abc_15724_n3875), .B(_abc_15724_n3867), .Y(_abc_15724_n3876) );
  AND2X2 AND2X2_1635 ( .A(_abc_15724_n3879), .B(_abc_15724_n3877), .Y(_abc_15724_n3880) );
  AND2X2 AND2X2_1636 ( .A(_abc_15724_n3866), .B(_abc_15724_n3881), .Y(_abc_15724_n3882) );
  AND2X2 AND2X2_1637 ( .A(_abc_15724_n3884), .B(_abc_15724_n3883), .Y(_abc_15724_n3885) );
  AND2X2 AND2X2_1638 ( .A(_abc_15724_n3726_bF_buf2), .B(_abc_15724_n3885), .Y(_abc_15724_n3886) );
  AND2X2 AND2X2_1639 ( .A(_abc_15724_n3737_bF_buf1), .B(_abc_15724_n3888), .Y(_abc_15724_n3889) );
  AND2X2 AND2X2_164 ( .A(_abc_15724_n1016_1), .B(_abc_15724_n1001), .Y(_abc_15724_n1030) );
  AND2X2 AND2X2_1640 ( .A(_abc_15724_n3892), .B(_abc_15724_n3893), .Y(_abc_15724_n3894) );
  AND2X2 AND2X2_1641 ( .A(_abc_15724_n3891), .B(_abc_15724_n3894), .Y(_abc_15724_n3895) );
  AND2X2 AND2X2_1642 ( .A(_abc_15724_n3899), .B(_abc_15724_n3900), .Y(_abc_15724_n3901) );
  AND2X2 AND2X2_1643 ( .A(_abc_15724_n3902), .B(_abc_15724_n3897), .Y(_abc_15724_n3903) );
  AND2X2 AND2X2_1644 ( .A(_abc_15724_n3906), .B(_abc_15724_n3905), .Y(_abc_15724_n3907) );
  AND2X2 AND2X2_1645 ( .A(_abc_15724_n3904), .B(_abc_15724_n3908), .Y(_abc_15724_n3909) );
  AND2X2 AND2X2_1646 ( .A(_abc_15724_n3907), .B(_abc_15724_n3706), .Y(_abc_15724_n3913) );
  AND2X2 AND2X2_1647 ( .A(_abc_15724_n3903), .B(_abc_15724_n3734), .Y(_abc_15724_n3914) );
  AND2X2 AND2X2_1648 ( .A(_abc_15724_n3916), .B(_abc_15724_n3910), .Y(_abc_15724_n3917) );
  AND2X2 AND2X2_1649 ( .A(_abc_15724_n3920), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n3921) );
  AND2X2 AND2X2_165 ( .A(_abc_15724_n1029), .B(_abc_15724_n1032), .Y(_abc_15724_n1033) );
  AND2X2 AND2X2_1650 ( .A(_abc_15724_n3921), .B(_abc_15724_n3919), .Y(_abc_15724_n3922) );
  AND2X2 AND2X2_1651 ( .A(_abc_15724_n2992_bF_buf1), .B(a_reg_2_), .Y(_abc_15724_n3923) );
  AND2X2 AND2X2_1652 ( .A(_abc_15724_n906_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_130_), .Y(_abc_15724_n3924) );
  AND2X2 AND2X2_1653 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n3924), .Y(_abc_15724_n3925) );
  AND2X2 AND2X2_1654 ( .A(_abc_15724_n3909), .B(_abc_15724_n3912), .Y(_abc_15724_n3929) );
  AND2X2 AND2X2_1655 ( .A(_abc_15724_n3934), .B(_abc_15724_n3935), .Y(_abc_15724_n3936) );
  AND2X2 AND2X2_1656 ( .A(c_reg_3_), .B(b_reg_3_), .Y(_abc_15724_n3937) );
  AND2X2 AND2X2_1657 ( .A(_abc_15724_n3938), .B(_abc_15724_n3933), .Y(_abc_15724_n3939) );
  AND2X2 AND2X2_1658 ( .A(_abc_15724_n3940), .B(_abc_15724_n3941), .Y(_abc_15724_n3942) );
  AND2X2 AND2X2_1659 ( .A(_abc_15724_n3726_bF_buf1), .B(_abc_15724_n3942), .Y(_abc_15724_n3943) );
  AND2X2 AND2X2_166 ( .A(_abc_15724_n1034), .B(_abc_15724_n1036), .Y(H3_reg_2__FF_INPUT) );
  AND2X2 AND2X2_1660 ( .A(_abc_15724_n3944), .B(_abc_15724_n3933), .Y(_abc_15724_n3945) );
  AND2X2 AND2X2_1661 ( .A(_abc_15724_n3934), .B(b_reg_3_), .Y(_abc_15724_n3946) );
  AND2X2 AND2X2_1662 ( .A(_abc_15724_n3737_bF_buf0), .B(_abc_15724_n3951), .Y(_abc_15724_n3952) );
  AND2X2 AND2X2_1663 ( .A(a_reg_30_), .B(e_reg_3_), .Y(_abc_15724_n3957) );
  AND2X2 AND2X2_1664 ( .A(_abc_15724_n3958), .B(_abc_15724_n3956), .Y(_abc_15724_n3959) );
  AND2X2 AND2X2_1665 ( .A(_abc_15724_n3959), .B(w_3_), .Y(_abc_15724_n3960) );
  AND2X2 AND2X2_1666 ( .A(_abc_15724_n3961), .B(_abc_15724_n3962), .Y(_abc_15724_n3963) );
  AND2X2 AND2X2_1667 ( .A(_abc_15724_n3963), .B(_abc_15724_n3955), .Y(_abc_15724_n3964) );
  AND2X2 AND2X2_1668 ( .A(_abc_15724_n3965), .B(_abc_15724_n3966), .Y(_abc_15724_n3967) );
  AND2X2 AND2X2_1669 ( .A(_abc_15724_n3972), .B(_abc_15724_n3948), .Y(_abc_15724_n3973) );
  AND2X2 AND2X2_167 ( .A(_abc_15724_n1029), .B(_abc_15724_n1026_1), .Y(_abc_15724_n1038_1) );
  AND2X2 AND2X2_1670 ( .A(_abc_15724_n3971), .B(_abc_15724_n3973), .Y(_abc_15724_n3974) );
  AND2X2 AND2X2_1671 ( .A(_abc_15724_n3977), .B(_abc_15724_n3975), .Y(_abc_15724_n3978) );
  AND2X2 AND2X2_1672 ( .A(_abc_15724_n3968), .B(_abc_15724_n3980), .Y(_abc_15724_n3981) );
  AND2X2 AND2X2_1673 ( .A(_abc_15724_n3932), .B(_abc_15724_n3981), .Y(_abc_15724_n3982) );
  AND2X2 AND2X2_1674 ( .A(_abc_15724_n3900), .B(_abc_15724_n3892), .Y(_abc_15724_n3983) );
  AND2X2 AND2X2_1675 ( .A(_abc_15724_n3974), .B(_abc_15724_n3979), .Y(_abc_15724_n3984) );
  AND2X2 AND2X2_1676 ( .A(_abc_15724_n3954), .B(_abc_15724_n3967), .Y(_abc_15724_n3985) );
  AND2X2 AND2X2_1677 ( .A(_abc_15724_n3986), .B(_abc_15724_n3983), .Y(_abc_15724_n3987) );
  AND2X2 AND2X2_1678 ( .A(_abc_15724_n3991), .B(_abc_15724_n3990), .Y(_abc_15724_n3992) );
  AND2X2 AND2X2_1679 ( .A(_abc_15724_n3989), .B(_abc_15724_n3993), .Y(_abc_15724_n3994) );
  AND2X2 AND2X2_168 ( .A(_auto_iopadmap_cc_313_execute_26059_35_), .B(d_reg_3_), .Y(_abc_15724_n1040) );
  AND2X2 AND2X2_1680 ( .A(_abc_15724_n3994), .B(_abc_15724_n3931), .Y(_abc_15724_n3995) );
  AND2X2 AND2X2_1681 ( .A(_abc_15724_n3908), .B(_abc_15724_n3897), .Y(_abc_15724_n3996) );
  AND2X2 AND2X2_1682 ( .A(_abc_15724_n3992), .B(_abc_15724_n3806_bF_buf3), .Y(_abc_15724_n3997) );
  AND2X2 AND2X2_1683 ( .A(_abc_15724_n3988), .B(_abc_15724_n3726_bF_buf4), .Y(_abc_15724_n3998) );
  AND2X2 AND2X2_1684 ( .A(_abc_15724_n3999), .B(_abc_15724_n3996), .Y(_abc_15724_n4000) );
  AND2X2 AND2X2_1685 ( .A(_abc_15724_n4007), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n4008) );
  AND2X2 AND2X2_1686 ( .A(_abc_15724_n4005), .B(_abc_15724_n4008), .Y(_abc_15724_n4009) );
  AND2X2 AND2X2_1687 ( .A(_abc_15724_n4009), .B(_abc_15724_n4004), .Y(_abc_15724_n4010) );
  AND2X2 AND2X2_1688 ( .A(_abc_15724_n2992_bF_buf0), .B(a_reg_3_), .Y(_abc_15724_n4011) );
  AND2X2 AND2X2_1689 ( .A(_abc_15724_n906_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_131_), .Y(_abc_15724_n4012) );
  AND2X2 AND2X2_169 ( .A(_abc_15724_n1041), .B(_abc_15724_n1039_1), .Y(_abc_15724_n1042) );
  AND2X2 AND2X2_1690 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n4012), .Y(_abc_15724_n4013) );
  AND2X2 AND2X2_1691 ( .A(_abc_15724_n4007), .B(_abc_15724_n4016), .Y(_abc_15724_n4017) );
  AND2X2 AND2X2_1692 ( .A(_abc_15724_n4005), .B(_abc_15724_n4017), .Y(_abc_15724_n4018) );
  AND2X2 AND2X2_1693 ( .A(_abc_15724_n3989), .B(_abc_15724_n3990), .Y(_abc_15724_n4020) );
  AND2X2 AND2X2_1694 ( .A(_abc_15724_n3706), .B(_abc_15724_n3721_bF_buf3), .Y(_abc_15724_n4021) );
  AND2X2 AND2X2_1695 ( .A(_abc_15724_n3980), .B(_abc_15724_n3965), .Y(_abc_15724_n4023) );
  AND2X2 AND2X2_1696 ( .A(_abc_15724_n4025), .B(_abc_15724_n4026), .Y(_abc_15724_n4027) );
  AND2X2 AND2X2_1697 ( .A(c_reg_4_), .B(b_reg_4_), .Y(_abc_15724_n4028) );
  AND2X2 AND2X2_1698 ( .A(_abc_15724_n4029), .B(_abc_15724_n4024), .Y(_abc_15724_n4030) );
  AND2X2 AND2X2_1699 ( .A(_abc_15724_n4035), .B(_abc_15724_n4024), .Y(_abc_15724_n4036) );
  AND2X2 AND2X2_17 ( .A(_abc_15724_n730_1), .B(_abc_15724_n731_1), .Y(_abc_15724_n732) );
  AND2X2 AND2X2_170 ( .A(_abc_15724_n1031), .B(_abc_15724_n1027), .Y(_abc_15724_n1045) );
  AND2X2 AND2X2_1700 ( .A(_abc_15724_n4025), .B(b_reg_4_), .Y(_abc_15724_n4037) );
  AND2X2 AND2X2_1701 ( .A(_abc_15724_n4041), .B(_abc_15724_n4039), .Y(_abc_15724_n4042) );
  AND2X2 AND2X2_1702 ( .A(_abc_15724_n4034), .B(_abc_15724_n4042), .Y(_abc_15724_n4043) );
  AND2X2 AND2X2_1703 ( .A(a_reg_31_), .B(e_reg_4_), .Y(_abc_15724_n4046) );
  AND2X2 AND2X2_1704 ( .A(_abc_15724_n4047), .B(_abc_15724_n4045), .Y(_abc_15724_n4048) );
  AND2X2 AND2X2_1705 ( .A(_abc_15724_n4048), .B(w_4_), .Y(_abc_15724_n4049) );
  AND2X2 AND2X2_1706 ( .A(_abc_15724_n4050), .B(_abc_15724_n4051), .Y(_abc_15724_n4052) );
  AND2X2 AND2X2_1707 ( .A(_abc_15724_n4052), .B(_abc_15724_n4044), .Y(_abc_15724_n4053) );
  AND2X2 AND2X2_1708 ( .A(_abc_15724_n4056), .B(_abc_15724_n4054), .Y(_abc_15724_n4057) );
  AND2X2 AND2X2_1709 ( .A(_abc_15724_n4043), .B(_abc_15724_n4058), .Y(_abc_15724_n4059) );
  AND2X2 AND2X2_171 ( .A(_abc_15724_n1044), .B(_abc_15724_n1047_1), .Y(_abc_15724_n1048_1) );
  AND2X2 AND2X2_1710 ( .A(_abc_15724_n4060), .B(_abc_15724_n4031), .Y(_abc_15724_n4061) );
  AND2X2 AND2X2_1711 ( .A(_abc_15724_n3726_bF_buf3), .B(_abc_15724_n4061), .Y(_abc_15724_n4062) );
  AND2X2 AND2X2_1712 ( .A(_abc_15724_n3737_bF_buf4), .B(_abc_15724_n4064), .Y(_abc_15724_n4065) );
  AND2X2 AND2X2_1713 ( .A(_abc_15724_n4068), .B(_abc_15724_n4069), .Y(_abc_15724_n4070) );
  AND2X2 AND2X2_1714 ( .A(_abc_15724_n4067), .B(_abc_15724_n4070), .Y(_abc_15724_n4071) );
  AND2X2 AND2X2_1715 ( .A(_abc_15724_n4075), .B(_abc_15724_n4076), .Y(_abc_15724_n4077) );
  AND2X2 AND2X2_1716 ( .A(_abc_15724_n4078), .B(_abc_15724_n4073), .Y(_abc_15724_n4079) );
  AND2X2 AND2X2_1717 ( .A(_abc_15724_n4079), .B(_abc_15724_n4022), .Y(_abc_15724_n4080) );
  AND2X2 AND2X2_1718 ( .A(_abc_15724_n4074), .B(_abc_15724_n4077), .Y(_abc_15724_n4081) );
  AND2X2 AND2X2_1719 ( .A(_abc_15724_n4072), .B(_abc_15724_n4023), .Y(_abc_15724_n4082) );
  AND2X2 AND2X2_172 ( .A(_abc_15724_n1048_1), .B(digest_update_bF_buf9), .Y(_abc_15724_n1049) );
  AND2X2 AND2X2_1720 ( .A(_abc_15724_n4083), .B(_abc_15724_n4021), .Y(_abc_15724_n4084) );
  AND2X2 AND2X2_1721 ( .A(_abc_15724_n4085), .B(_abc_15724_n4020), .Y(_abc_15724_n4088) );
  AND2X2 AND2X2_1722 ( .A(_abc_15724_n4019), .B(_abc_15724_n4090), .Y(_abc_15724_n4092) );
  AND2X2 AND2X2_1723 ( .A(_abc_15724_n4093), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n4094) );
  AND2X2 AND2X2_1724 ( .A(_abc_15724_n4094), .B(_abc_15724_n4091), .Y(_abc_15724_n4095) );
  AND2X2 AND2X2_1725 ( .A(_abc_15724_n2992_bF_buf11), .B(a_reg_4_), .Y(_abc_15724_n4096) );
  AND2X2 AND2X2_1726 ( .A(_abc_15724_n906_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_132_), .Y(_abc_15724_n4097) );
  AND2X2 AND2X2_1727 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n4097), .Y(_abc_15724_n4098) );
  AND2X2 AND2X2_1728 ( .A(_abc_15724_n4076), .B(_abc_15724_n4068), .Y(_abc_15724_n4102) );
  AND2X2 AND2X2_1729 ( .A(_abc_15724_n4104), .B(_abc_15724_n4105), .Y(_abc_15724_n4106) );
  AND2X2 AND2X2_173 ( .A(_abc_15724_n907_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_35_), .Y(_abc_15724_n1050_1) );
  AND2X2 AND2X2_1730 ( .A(c_reg_5_), .B(b_reg_5_), .Y(_abc_15724_n4107) );
  AND2X2 AND2X2_1731 ( .A(_abc_15724_n4108), .B(_abc_15724_n4103), .Y(_abc_15724_n4109) );
  AND2X2 AND2X2_1732 ( .A(_abc_15724_n4114), .B(_abc_15724_n4103), .Y(_abc_15724_n4115) );
  AND2X2 AND2X2_1733 ( .A(_abc_15724_n4104), .B(b_reg_5_), .Y(_abc_15724_n4116) );
  AND2X2 AND2X2_1734 ( .A(_abc_15724_n4120), .B(_abc_15724_n4118), .Y(_abc_15724_n4121) );
  AND2X2 AND2X2_1735 ( .A(_abc_15724_n4113), .B(_abc_15724_n4121), .Y(_abc_15724_n4122) );
  AND2X2 AND2X2_1736 ( .A(a_reg_0_), .B(e_reg_5_), .Y(_abc_15724_n4125) );
  AND2X2 AND2X2_1737 ( .A(_abc_15724_n4126), .B(_abc_15724_n4124), .Y(_abc_15724_n4127) );
  AND2X2 AND2X2_1738 ( .A(_abc_15724_n4127), .B(w_5_), .Y(_abc_15724_n4128) );
  AND2X2 AND2X2_1739 ( .A(_abc_15724_n4129), .B(_abc_15724_n4130), .Y(_abc_15724_n4131) );
  AND2X2 AND2X2_174 ( .A(_auto_iopadmap_cc_313_execute_26059_36_), .B(d_reg_4_), .Y(_abc_15724_n1053) );
  AND2X2 AND2X2_1740 ( .A(_abc_15724_n4131), .B(_abc_15724_n4123), .Y(_abc_15724_n4132) );
  AND2X2 AND2X2_1741 ( .A(_abc_15724_n4135), .B(_abc_15724_n4133), .Y(_abc_15724_n4136) );
  AND2X2 AND2X2_1742 ( .A(_abc_15724_n4122), .B(_abc_15724_n4137), .Y(_abc_15724_n4138) );
  AND2X2 AND2X2_1743 ( .A(_abc_15724_n4139), .B(_abc_15724_n4110), .Y(_abc_15724_n4140) );
  AND2X2 AND2X2_1744 ( .A(_abc_15724_n3726_bF_buf2), .B(_abc_15724_n4140), .Y(_abc_15724_n4141) );
  AND2X2 AND2X2_1745 ( .A(_abc_15724_n3737_bF_buf3), .B(_abc_15724_n4143), .Y(_abc_15724_n4144) );
  AND2X2 AND2X2_1746 ( .A(_abc_15724_n4147), .B(_abc_15724_n4148), .Y(_abc_15724_n4149) );
  AND2X2 AND2X2_1747 ( .A(_abc_15724_n4146), .B(_abc_15724_n4149), .Y(_abc_15724_n4150) );
  AND2X2 AND2X2_1748 ( .A(_abc_15724_n4154), .B(_abc_15724_n4155), .Y(_abc_15724_n4156) );
  AND2X2 AND2X2_1749 ( .A(_abc_15724_n4157), .B(_abc_15724_n4152), .Y(_abc_15724_n4158) );
  AND2X2 AND2X2_175 ( .A(_abc_15724_n1054), .B(_abc_15724_n1052), .Y(_abc_15724_n1055) );
  AND2X2 AND2X2_1750 ( .A(_abc_15724_n4153), .B(_abc_15724_n4156), .Y(_abc_15724_n4160) );
  AND2X2 AND2X2_1751 ( .A(_abc_15724_n4151), .B(_abc_15724_n4102), .Y(_abc_15724_n4161) );
  AND2X2 AND2X2_1752 ( .A(_abc_15724_n4163), .B(_abc_15724_n4159), .Y(_abc_15724_n4164) );
  AND2X2 AND2X2_1753 ( .A(_abc_15724_n4164), .B(_abc_15724_n4101), .Y(_abc_15724_n4165) );
  AND2X2 AND2X2_1754 ( .A(_abc_15724_n4166), .B(_abc_15724_n4073), .Y(_abc_15724_n4167) );
  AND2X2 AND2X2_1755 ( .A(_abc_15724_n4162), .B(_abc_15724_n4022), .Y(_abc_15724_n4168) );
  AND2X2 AND2X2_1756 ( .A(_abc_15724_n4158), .B(_abc_15724_n4021), .Y(_abc_15724_n4169) );
  AND2X2 AND2X2_1757 ( .A(_abc_15724_n4170), .B(_abc_15724_n4167), .Y(_abc_15724_n4171) );
  AND2X2 AND2X2_1758 ( .A(_abc_15724_n4019), .B(_abc_15724_n4177), .Y(_abc_15724_n4178) );
  AND2X2 AND2X2_1759 ( .A(_abc_15724_n4180), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n4181) );
  AND2X2 AND2X2_176 ( .A(_abc_15724_n1058), .B(_abc_15724_n1041), .Y(_abc_15724_n1059) );
  AND2X2 AND2X2_1760 ( .A(_abc_15724_n4179), .B(_abc_15724_n4181), .Y(_abc_15724_n4182) );
  AND2X2 AND2X2_1761 ( .A(_abc_15724_n4182), .B(_abc_15724_n4175), .Y(_abc_15724_n4183) );
  AND2X2 AND2X2_1762 ( .A(_abc_15724_n2992_bF_buf10), .B(a_reg_5_), .Y(_abc_15724_n4184) );
  AND2X2 AND2X2_1763 ( .A(_abc_15724_n906_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_133_), .Y(_abc_15724_n4185) );
  AND2X2 AND2X2_1764 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n4185), .Y(_abc_15724_n4186) );
  AND2X2 AND2X2_1765 ( .A(_abc_15724_n4180), .B(_abc_15724_n4189), .Y(_abc_15724_n4190) );
  AND2X2 AND2X2_1766 ( .A(_abc_15724_n4179), .B(_abc_15724_n4190), .Y(_abc_15724_n4191) );
  AND2X2 AND2X2_1767 ( .A(_abc_15724_n4163), .B(_abc_15724_n4152), .Y(_abc_15724_n4193) );
  AND2X2 AND2X2_1768 ( .A(_abc_15724_n4155), .B(_abc_15724_n4147), .Y(_abc_15724_n4195) );
  AND2X2 AND2X2_1769 ( .A(_abc_15724_n4197), .B(_abc_15724_n4198), .Y(_abc_15724_n4199) );
  AND2X2 AND2X2_177 ( .A(_abc_15724_n1046), .B(_abc_15724_n1039_1), .Y(_abc_15724_n1061_1) );
  AND2X2 AND2X2_1770 ( .A(c_reg_6_), .B(b_reg_6_), .Y(_abc_15724_n4200) );
  AND2X2 AND2X2_1771 ( .A(_abc_15724_n4201), .B(_abc_15724_n4196), .Y(_abc_15724_n4202) );
  AND2X2 AND2X2_1772 ( .A(_abc_15724_n4203), .B(_abc_15724_n4204), .Y(_abc_15724_n4205) );
  AND2X2 AND2X2_1773 ( .A(_abc_15724_n3726_bF_buf1), .B(_abc_15724_n4205), .Y(_abc_15724_n4206) );
  AND2X2 AND2X2_1774 ( .A(_abc_15724_n4196), .B(_abc_15724_n4198), .Y(_abc_15724_n4207) );
  AND2X2 AND2X2_1775 ( .A(_abc_15724_n4197), .B(b_reg_6_), .Y(_abc_15724_n4208) );
  AND2X2 AND2X2_1776 ( .A(_abc_15724_n4212), .B(_abc_15724_n4196), .Y(_abc_15724_n4213) );
  AND2X2 AND2X2_1777 ( .A(_abc_15724_n3737_bF_buf2), .B(_abc_15724_n4215), .Y(_abc_15724_n4216) );
  AND2X2 AND2X2_1778 ( .A(_abc_15724_n4129), .B(_abc_15724_n4126), .Y(_abc_15724_n4220) );
  AND2X2 AND2X2_1779 ( .A(a_reg_1_), .B(e_reg_6_), .Y(_abc_15724_n4223) );
  AND2X2 AND2X2_178 ( .A(_abc_15724_n1060_1), .B(_abc_15724_n1063_1), .Y(_abc_15724_n1064) );
  AND2X2 AND2X2_1780 ( .A(_abc_15724_n4224), .B(_abc_15724_n4222), .Y(_abc_15724_n4225) );
  AND2X2 AND2X2_1781 ( .A(_abc_15724_n4225), .B(w_6_), .Y(_abc_15724_n4226) );
  AND2X2 AND2X2_1782 ( .A(_abc_15724_n4227), .B(_abc_15724_n4228), .Y(_abc_15724_n4229) );
  AND2X2 AND2X2_1783 ( .A(_abc_15724_n4221), .B(_abc_15724_n4229), .Y(_abc_15724_n4230) );
  AND2X2 AND2X2_1784 ( .A(_abc_15724_n4231), .B(_abc_15724_n4220), .Y(_abc_15724_n4232) );
  AND2X2 AND2X2_1785 ( .A(_abc_15724_n4219), .B(_abc_15724_n4233), .Y(_abc_15724_n4234) );
  AND2X2 AND2X2_1786 ( .A(_abc_15724_n4235), .B(_abc_15724_n4236), .Y(_abc_15724_n4237) );
  AND2X2 AND2X2_1787 ( .A(_abc_15724_n4237), .B(_abc_15724_n4218), .Y(_abc_15724_n4238) );
  AND2X2 AND2X2_1788 ( .A(_abc_15724_n4243), .B(_abc_15724_n4242), .Y(_abc_15724_n4244) );
  AND2X2 AND2X2_1789 ( .A(_abc_15724_n4245), .B(_abc_15724_n4240), .Y(_abc_15724_n4246) );
  AND2X2 AND2X2_179 ( .A(_abc_15724_n1065), .B(_abc_15724_n1067), .Y(H3_reg_4__FF_INPUT) );
  AND2X2 AND2X2_1790 ( .A(_abc_15724_n4244), .B(_abc_15724_n4241), .Y(_abc_15724_n4248) );
  AND2X2 AND2X2_1791 ( .A(_abc_15724_n4239), .B(_abc_15724_n4195), .Y(_abc_15724_n4249) );
  AND2X2 AND2X2_1792 ( .A(_abc_15724_n4251), .B(_abc_15724_n4247), .Y(_abc_15724_n4252) );
  AND2X2 AND2X2_1793 ( .A(_abc_15724_n4194), .B(_abc_15724_n4252), .Y(_abc_15724_n4253) );
  AND2X2 AND2X2_1794 ( .A(_abc_15724_n4250), .B(_abc_15724_n3706), .Y(_abc_15724_n4254) );
  AND2X2 AND2X2_1795 ( .A(_abc_15724_n4246), .B(_abc_15724_n3734), .Y(_abc_15724_n4255) );
  AND2X2 AND2X2_1796 ( .A(_abc_15724_n4256), .B(_abc_15724_n4193), .Y(_abc_15724_n4257) );
  AND2X2 AND2X2_1797 ( .A(_abc_15724_n4192), .B(_abc_15724_n4259), .Y(_abc_15724_n4260) );
  AND2X2 AND2X2_1798 ( .A(_abc_15724_n4262), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n4263) );
  AND2X2 AND2X2_1799 ( .A(_abc_15724_n4263), .B(_abc_15724_n4261), .Y(_abc_15724_n4264) );
  AND2X2 AND2X2_18 ( .A(_auto_iopadmap_cc_313_execute_26059_14_), .B(e_reg_14_), .Y(_abc_15724_n733) );
  AND2X2 AND2X2_180 ( .A(_abc_15724_n1062), .B(_abc_15724_n1055), .Y(_abc_15724_n1069_1) );
  AND2X2 AND2X2_1800 ( .A(_abc_15724_n2992_bF_buf9), .B(a_reg_6_), .Y(_abc_15724_n4265) );
  AND2X2 AND2X2_1801 ( .A(_abc_15724_n906_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_134_), .Y(_abc_15724_n4266) );
  AND2X2 AND2X2_1802 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n4266), .Y(_abc_15724_n4267) );
  AND2X2 AND2X2_1803 ( .A(_abc_15724_n4261), .B(_abc_15724_n4270), .Y(_abc_15724_n4271) );
  AND2X2 AND2X2_1804 ( .A(_abc_15724_n4243), .B(_abc_15724_n4235), .Y(_abc_15724_n4274) );
  AND2X2 AND2X2_1805 ( .A(_abc_15724_n4277), .B(_abc_15724_n4278), .Y(_abc_15724_n4279) );
  AND2X2 AND2X2_1806 ( .A(c_reg_7_), .B(b_reg_7_), .Y(_abc_15724_n4280) );
  AND2X2 AND2X2_1807 ( .A(_abc_15724_n4281), .B(_abc_15724_n4276), .Y(_abc_15724_n4282) );
  AND2X2 AND2X2_1808 ( .A(_abc_15724_n4287), .B(_abc_15724_n4276), .Y(_abc_15724_n4288) );
  AND2X2 AND2X2_1809 ( .A(_abc_15724_n4277), .B(b_reg_7_), .Y(_abc_15724_n4289) );
  AND2X2 AND2X2_181 ( .A(_auto_iopadmap_cc_313_execute_26059_37_), .B(d_reg_5_), .Y(_abc_15724_n1072) );
  AND2X2 AND2X2_1810 ( .A(_abc_15724_n4293), .B(_abc_15724_n4291), .Y(_abc_15724_n4294) );
  AND2X2 AND2X2_1811 ( .A(_abc_15724_n4286), .B(_abc_15724_n4294), .Y(_abc_15724_n4295) );
  AND2X2 AND2X2_1812 ( .A(a_reg_2_), .B(e_reg_7_), .Y(_abc_15724_n4298) );
  AND2X2 AND2X2_1813 ( .A(_abc_15724_n4299), .B(_abc_15724_n4297), .Y(_abc_15724_n4300) );
  AND2X2 AND2X2_1814 ( .A(_abc_15724_n4300), .B(w_7_), .Y(_abc_15724_n4301) );
  AND2X2 AND2X2_1815 ( .A(_abc_15724_n4302), .B(_abc_15724_n4303), .Y(_abc_15724_n4304) );
  AND2X2 AND2X2_1816 ( .A(_abc_15724_n4304), .B(_abc_15724_n4296), .Y(_abc_15724_n4305) );
  AND2X2 AND2X2_1817 ( .A(_abc_15724_n4308), .B(_abc_15724_n4306), .Y(_abc_15724_n4309) );
  AND2X2 AND2X2_1818 ( .A(_abc_15724_n4295), .B(_abc_15724_n4310), .Y(_abc_15724_n4311) );
  AND2X2 AND2X2_1819 ( .A(_abc_15724_n4312), .B(_abc_15724_n4283), .Y(_abc_15724_n4313) );
  AND2X2 AND2X2_182 ( .A(_abc_15724_n1073), .B(_abc_15724_n1071_1), .Y(_abc_15724_n1074) );
  AND2X2 AND2X2_1820 ( .A(_abc_15724_n3726_bF_buf0), .B(_abc_15724_n4313), .Y(_abc_15724_n4314) );
  AND2X2 AND2X2_1821 ( .A(_abc_15724_n3737_bF_buf1), .B(_abc_15724_n4316), .Y(_abc_15724_n4317) );
  AND2X2 AND2X2_1822 ( .A(_abc_15724_n4320), .B(_abc_15724_n4321), .Y(_abc_15724_n4322) );
  AND2X2 AND2X2_1823 ( .A(_abc_15724_n4319), .B(_abc_15724_n4322), .Y(_abc_15724_n4323) );
  AND2X2 AND2X2_1824 ( .A(_abc_15724_n4275), .B(_abc_15724_n4325), .Y(_abc_15724_n4326) );
  AND2X2 AND2X2_1825 ( .A(_abc_15724_n4274), .B(_abc_15724_n4324), .Y(_abc_15724_n4327) );
  AND2X2 AND2X2_1826 ( .A(_abc_15724_n4273), .B(_abc_15724_n4328), .Y(_abc_15724_n4329) );
  AND2X2 AND2X2_1827 ( .A(_abc_15724_n4251), .B(_abc_15724_n4240), .Y(_abc_15724_n4330) );
  AND2X2 AND2X2_1828 ( .A(_abc_15724_n4330), .B(_abc_15724_n4331), .Y(_abc_15724_n4332) );
  AND2X2 AND2X2_1829 ( .A(_abc_15724_n4336), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n4337) );
  AND2X2 AND2X2_183 ( .A(_abc_15724_n1060_1), .B(_abc_15724_n1054), .Y(_abc_15724_n1076) );
  AND2X2 AND2X2_1830 ( .A(_abc_15724_n4337), .B(_abc_15724_n4335), .Y(_abc_15724_n4338) );
  AND2X2 AND2X2_1831 ( .A(_abc_15724_n2992_bF_buf8), .B(a_reg_7_), .Y(_abc_15724_n4339) );
  AND2X2 AND2X2_1832 ( .A(_abc_15724_n906_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_135_), .Y(_abc_15724_n4340) );
  AND2X2 AND2X2_1833 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n4340), .Y(_abc_15724_n4341) );
  AND2X2 AND2X2_1834 ( .A(_abc_15724_n4270), .B(_abc_15724_n4348), .Y(_abc_15724_n4349) );
  AND2X2 AND2X2_1835 ( .A(_abc_15724_n4347), .B(_abc_15724_n4350), .Y(_abc_15724_n4351) );
  AND2X2 AND2X2_1836 ( .A(_abc_15724_n4346), .B(_abc_15724_n4351), .Y(_abc_15724_n4352) );
  AND2X2 AND2X2_1837 ( .A(_abc_15724_n4354), .B(_abc_15724_n4320), .Y(_abc_15724_n4355) );
  AND2X2 AND2X2_1838 ( .A(_abc_15724_n4357), .B(_abc_15724_n4358), .Y(_abc_15724_n4359) );
  AND2X2 AND2X2_1839 ( .A(c_reg_8_), .B(b_reg_8_), .Y(_abc_15724_n4360) );
  AND2X2 AND2X2_184 ( .A(_abc_15724_n1078), .B(_abc_15724_n1075), .Y(_abc_15724_n1079) );
  AND2X2 AND2X2_1840 ( .A(_abc_15724_n4361), .B(_abc_15724_n4356), .Y(_abc_15724_n4362) );
  AND2X2 AND2X2_1841 ( .A(_abc_15724_n4367), .B(_abc_15724_n4356), .Y(_abc_15724_n4368) );
  AND2X2 AND2X2_1842 ( .A(_abc_15724_n4357), .B(b_reg_8_), .Y(_abc_15724_n4369) );
  AND2X2 AND2X2_1843 ( .A(_abc_15724_n4373), .B(_abc_15724_n4371), .Y(_abc_15724_n4374) );
  AND2X2 AND2X2_1844 ( .A(_abc_15724_n4366), .B(_abc_15724_n4374), .Y(_abc_15724_n4375) );
  AND2X2 AND2X2_1845 ( .A(a_reg_3_), .B(e_reg_8_), .Y(_abc_15724_n4378) );
  AND2X2 AND2X2_1846 ( .A(_abc_15724_n4379), .B(_abc_15724_n4377), .Y(_abc_15724_n4380) );
  AND2X2 AND2X2_1847 ( .A(_abc_15724_n4380), .B(w_8_), .Y(_abc_15724_n4381) );
  AND2X2 AND2X2_1848 ( .A(_abc_15724_n4382), .B(_abc_15724_n4383), .Y(_abc_15724_n4384) );
  AND2X2 AND2X2_1849 ( .A(_abc_15724_n4384), .B(_abc_15724_n4376), .Y(_abc_15724_n4385) );
  AND2X2 AND2X2_185 ( .A(_abc_15724_n1079), .B(digest_update_bF_buf7), .Y(_abc_15724_n1080) );
  AND2X2 AND2X2_1850 ( .A(_abc_15724_n4388), .B(_abc_15724_n4386), .Y(_abc_15724_n4389) );
  AND2X2 AND2X2_1851 ( .A(_abc_15724_n4375), .B(_abc_15724_n4390), .Y(_abc_15724_n4391) );
  AND2X2 AND2X2_1852 ( .A(_abc_15724_n4392), .B(_abc_15724_n4363), .Y(_abc_15724_n4393) );
  AND2X2 AND2X2_1853 ( .A(_abc_15724_n3726_bF_buf4), .B(_abc_15724_n4393), .Y(_abc_15724_n4394) );
  AND2X2 AND2X2_1854 ( .A(_abc_15724_n3737_bF_buf0), .B(_abc_15724_n4396), .Y(_abc_15724_n4397) );
  AND2X2 AND2X2_1855 ( .A(_abc_15724_n4400), .B(_abc_15724_n4401), .Y(_abc_15724_n4402) );
  AND2X2 AND2X2_1856 ( .A(_abc_15724_n4399), .B(_abc_15724_n4402), .Y(_abc_15724_n4403) );
  AND2X2 AND2X2_1857 ( .A(_abc_15724_n4407), .B(_abc_15724_n4408), .Y(_abc_15724_n4409) );
  AND2X2 AND2X2_1858 ( .A(_abc_15724_n4410), .B(_abc_15724_n4405), .Y(_abc_15724_n4411) );
  AND2X2 AND2X2_1859 ( .A(_abc_15724_n4411), .B(_abc_15724_n3725_bF_buf3), .Y(_abc_15724_n4412) );
  AND2X2 AND2X2_186 ( .A(_abc_15724_n1081), .B(_abc_15724_n850_bF_buf5), .Y(_abc_15724_n1082_1) );
  AND2X2 AND2X2_1860 ( .A(_abc_15724_n4406), .B(_abc_15724_n4409), .Y(_abc_15724_n4413) );
  AND2X2 AND2X2_1861 ( .A(_abc_15724_n4404), .B(_abc_15724_n4355), .Y(_abc_15724_n4414) );
  AND2X2 AND2X2_1862 ( .A(_abc_15724_n4415), .B(_abc_15724_n3737_bF_buf4), .Y(_abc_15724_n4416) );
  AND2X2 AND2X2_1863 ( .A(_abc_15724_n4417), .B(_abc_15724_n4327), .Y(_abc_15724_n4420) );
  AND2X2 AND2X2_1864 ( .A(_abc_15724_n4353), .B(_abc_15724_n4422), .Y(_abc_15724_n4423) );
  AND2X2 AND2X2_1865 ( .A(_abc_15724_n4425), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n4426) );
  AND2X2 AND2X2_1866 ( .A(_abc_15724_n4426), .B(_abc_15724_n4424), .Y(_abc_15724_n4427) );
  AND2X2 AND2X2_1867 ( .A(_abc_15724_n2992_bF_buf7), .B(a_reg_8_), .Y(_abc_15724_n4428) );
  AND2X2 AND2X2_1868 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n2606), .Y(_abc_15724_n4429) );
  AND2X2 AND2X2_1869 ( .A(_abc_15724_n4408), .B(_abc_15724_n4400), .Y(_abc_15724_n4433) );
  AND2X2 AND2X2_187 ( .A(_abc_15724_n1070_1), .B(_abc_15724_n1074), .Y(_abc_15724_n1084_1) );
  AND2X2 AND2X2_1870 ( .A(_abc_15724_n4435), .B(_abc_15724_n4436), .Y(_abc_15724_n4437) );
  AND2X2 AND2X2_1871 ( .A(c_reg_9_), .B(b_reg_9_), .Y(_abc_15724_n4438) );
  AND2X2 AND2X2_1872 ( .A(_abc_15724_n4439), .B(_abc_15724_n4434), .Y(_abc_15724_n4440) );
  AND2X2 AND2X2_1873 ( .A(_abc_15724_n4445), .B(_abc_15724_n4434), .Y(_abc_15724_n4446) );
  AND2X2 AND2X2_1874 ( .A(_abc_15724_n4435), .B(b_reg_9_), .Y(_abc_15724_n4447) );
  AND2X2 AND2X2_1875 ( .A(_abc_15724_n4451), .B(_abc_15724_n4449), .Y(_abc_15724_n4452) );
  AND2X2 AND2X2_1876 ( .A(_abc_15724_n4444), .B(_abc_15724_n4452), .Y(_abc_15724_n4453) );
  AND2X2 AND2X2_1877 ( .A(a_reg_4_), .B(e_reg_9_), .Y(_abc_15724_n4456) );
  AND2X2 AND2X2_1878 ( .A(_abc_15724_n4457), .B(_abc_15724_n4455), .Y(_abc_15724_n4458) );
  AND2X2 AND2X2_1879 ( .A(_abc_15724_n4458), .B(w_9_), .Y(_abc_15724_n4459) );
  AND2X2 AND2X2_188 ( .A(_auto_iopadmap_cc_313_execute_26059_38_), .B(d_reg_6_), .Y(_abc_15724_n1087) );
  AND2X2 AND2X2_1880 ( .A(_abc_15724_n4460), .B(_abc_15724_n4461), .Y(_abc_15724_n4462) );
  AND2X2 AND2X2_1881 ( .A(_abc_15724_n4462), .B(_abc_15724_n4454), .Y(_abc_15724_n4463) );
  AND2X2 AND2X2_1882 ( .A(_abc_15724_n4466), .B(_abc_15724_n4464), .Y(_abc_15724_n4467) );
  AND2X2 AND2X2_1883 ( .A(_abc_15724_n4453), .B(_abc_15724_n4468), .Y(_abc_15724_n4469) );
  AND2X2 AND2X2_1884 ( .A(_abc_15724_n4470), .B(_abc_15724_n4441), .Y(_abc_15724_n4471) );
  AND2X2 AND2X2_1885 ( .A(_abc_15724_n3726_bF_buf3), .B(_abc_15724_n4471), .Y(_abc_15724_n4472) );
  AND2X2 AND2X2_1886 ( .A(_abc_15724_n3737_bF_buf3), .B(_abc_15724_n4474), .Y(_abc_15724_n4475) );
  AND2X2 AND2X2_1887 ( .A(_abc_15724_n4478), .B(_abc_15724_n4479), .Y(_abc_15724_n4480) );
  AND2X2 AND2X2_1888 ( .A(_abc_15724_n4477), .B(_abc_15724_n4480), .Y(_abc_15724_n4481) );
  AND2X2 AND2X2_1889 ( .A(_abc_15724_n4485), .B(_abc_15724_n4486), .Y(_abc_15724_n4487) );
  AND2X2 AND2X2_189 ( .A(_abc_15724_n1088), .B(_abc_15724_n1086), .Y(_abc_15724_n1089) );
  AND2X2 AND2X2_1890 ( .A(_abc_15724_n4488), .B(_abc_15724_n4483), .Y(_abc_15724_n4489) );
  AND2X2 AND2X2_1891 ( .A(_abc_15724_n4484), .B(_abc_15724_n4487), .Y(_abc_15724_n4491) );
  AND2X2 AND2X2_1892 ( .A(_abc_15724_n4482), .B(_abc_15724_n4433), .Y(_abc_15724_n4492) );
  AND2X2 AND2X2_1893 ( .A(_abc_15724_n4494), .B(_abc_15724_n4490), .Y(_abc_15724_n4495) );
  AND2X2 AND2X2_1894 ( .A(_abc_15724_n4495), .B(_abc_15724_n4432), .Y(_abc_15724_n4496) );
  AND2X2 AND2X2_1895 ( .A(_abc_15724_n4497), .B(_abc_15724_n4405), .Y(_abc_15724_n4498) );
  AND2X2 AND2X2_1896 ( .A(_abc_15724_n4493), .B(_abc_15724_n4022), .Y(_abc_15724_n4499) );
  AND2X2 AND2X2_1897 ( .A(_abc_15724_n4489), .B(_abc_15724_n4021), .Y(_abc_15724_n4500) );
  AND2X2 AND2X2_1898 ( .A(_abc_15724_n4501), .B(_abc_15724_n4498), .Y(_abc_15724_n4502) );
  AND2X2 AND2X2_1899 ( .A(_abc_15724_n4423), .B(_abc_15724_n4504), .Y(_abc_15724_n4505) );
  AND2X2 AND2X2_19 ( .A(_abc_15724_n734), .B(_abc_15724_n735), .Y(_abc_15724_n736) );
  AND2X2 AND2X2_190 ( .A(_abc_15724_n1078), .B(_abc_15724_n1073), .Y(_abc_15724_n1091_1) );
  AND2X2 AND2X2_1900 ( .A(_abc_15724_n4509), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n4510) );
  AND2X2 AND2X2_1901 ( .A(_abc_15724_n4508), .B(_abc_15724_n4510), .Y(_abc_15724_n4511) );
  AND2X2 AND2X2_1902 ( .A(_abc_15724_n4511), .B(_abc_15724_n4506), .Y(_abc_15724_n4512) );
  AND2X2 AND2X2_1903 ( .A(_abc_15724_n2992_bF_buf6), .B(a_reg_9_), .Y(_abc_15724_n4513) );
  AND2X2 AND2X2_1904 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n2620), .Y(_abc_15724_n4514) );
  AND2X2 AND2X2_1905 ( .A(_abc_15724_n4509), .B(_abc_15724_n4517), .Y(_abc_15724_n4518) );
  AND2X2 AND2X2_1906 ( .A(_abc_15724_n4494), .B(_abc_15724_n4483), .Y(_abc_15724_n4521) );
  AND2X2 AND2X2_1907 ( .A(_abc_15724_n4486), .B(_abc_15724_n4478), .Y(_abc_15724_n4523) );
  AND2X2 AND2X2_1908 ( .A(_abc_15724_n4525), .B(_abc_15724_n4526), .Y(_abc_15724_n4527) );
  AND2X2 AND2X2_1909 ( .A(c_reg_10_), .B(b_reg_10_), .Y(_abc_15724_n4528) );
  AND2X2 AND2X2_191 ( .A(_abc_15724_n1093), .B(_abc_15724_n1090_1), .Y(_abc_15724_n1094) );
  AND2X2 AND2X2_1910 ( .A(_abc_15724_n4529), .B(_abc_15724_n4524), .Y(_abc_15724_n4530) );
  AND2X2 AND2X2_1911 ( .A(_abc_15724_n4531), .B(_abc_15724_n4532), .Y(_abc_15724_n4533) );
  AND2X2 AND2X2_1912 ( .A(_abc_15724_n3726_bF_buf2), .B(_abc_15724_n4533), .Y(_abc_15724_n4534) );
  AND2X2 AND2X2_1913 ( .A(_abc_15724_n4524), .B(_abc_15724_n4526), .Y(_abc_15724_n4536) );
  AND2X2 AND2X2_1914 ( .A(_abc_15724_n4525), .B(b_reg_10_), .Y(_abc_15724_n4537) );
  AND2X2 AND2X2_1915 ( .A(_abc_15724_n4540), .B(_abc_15724_n4524), .Y(_abc_15724_n4541) );
  AND2X2 AND2X2_1916 ( .A(_abc_15724_n4543), .B(_abc_15724_n4539), .Y(_abc_15724_n4544) );
  AND2X2 AND2X2_1917 ( .A(_abc_15724_n4535), .B(_abc_15724_n4544), .Y(_abc_15724_n4545) );
  AND2X2 AND2X2_1918 ( .A(_abc_15724_n4460), .B(_abc_15724_n4457), .Y(_abc_15724_n4546) );
  AND2X2 AND2X2_1919 ( .A(a_reg_5_), .B(e_reg_10_), .Y(_abc_15724_n4549) );
  AND2X2 AND2X2_192 ( .A(_abc_15724_n1094), .B(digest_update_bF_buf6), .Y(_abc_15724_n1095) );
  AND2X2 AND2X2_1920 ( .A(_abc_15724_n4550), .B(_abc_15724_n4548), .Y(_abc_15724_n4551) );
  AND2X2 AND2X2_1921 ( .A(_abc_15724_n4551), .B(w_10_), .Y(_abc_15724_n4552) );
  AND2X2 AND2X2_1922 ( .A(_abc_15724_n4553), .B(_abc_15724_n4554), .Y(_abc_15724_n4555) );
  AND2X2 AND2X2_1923 ( .A(_abc_15724_n4547), .B(_abc_15724_n4555), .Y(_abc_15724_n4556) );
  AND2X2 AND2X2_1924 ( .A(_abc_15724_n4559), .B(_abc_15724_n4545), .Y(_abc_15724_n4560) );
  AND2X2 AND2X2_1925 ( .A(_abc_15724_n4563), .B(_abc_15724_n4557), .Y(_abc_15724_n4564) );
  AND2X2 AND2X2_1926 ( .A(_abc_15724_n4562), .B(_abc_15724_n4564), .Y(_abc_15724_n4565) );
  AND2X2 AND2X2_1927 ( .A(_abc_15724_n4570), .B(_abc_15724_n4569), .Y(_abc_15724_n4571) );
  AND2X2 AND2X2_1928 ( .A(_abc_15724_n4567), .B(_abc_15724_n4572), .Y(_abc_15724_n4573) );
  AND2X2 AND2X2_1929 ( .A(_abc_15724_n4571), .B(_abc_15724_n4568), .Y(_abc_15724_n4575) );
  AND2X2 AND2X2_193 ( .A(_abc_15724_n1096), .B(_abc_15724_n850_bF_buf4), .Y(_abc_15724_n1097) );
  AND2X2 AND2X2_1930 ( .A(_abc_15724_n4566), .B(_abc_15724_n4523), .Y(_abc_15724_n4576) );
  AND2X2 AND2X2_1931 ( .A(_abc_15724_n4578), .B(_abc_15724_n4574), .Y(_abc_15724_n4579) );
  AND2X2 AND2X2_1932 ( .A(_abc_15724_n4579), .B(_abc_15724_n4522), .Y(_abc_15724_n4580) );
  AND2X2 AND2X2_1933 ( .A(_abc_15724_n4577), .B(_abc_15724_n3725_bF_buf3), .Y(_abc_15724_n4581) );
  AND2X2 AND2X2_1934 ( .A(_abc_15724_n4573), .B(_abc_15724_n3737_bF_buf0), .Y(_abc_15724_n4582) );
  AND2X2 AND2X2_1935 ( .A(_abc_15724_n4583), .B(_abc_15724_n4521), .Y(_abc_15724_n4584) );
  AND2X2 AND2X2_1936 ( .A(_abc_15724_n4520), .B(_abc_15724_n4586), .Y(_abc_15724_n4587) );
  AND2X2 AND2X2_1937 ( .A(_abc_15724_n4589), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n4590) );
  AND2X2 AND2X2_1938 ( .A(_abc_15724_n4590), .B(_abc_15724_n4588), .Y(_abc_15724_n4591) );
  AND2X2 AND2X2_1939 ( .A(_abc_15724_n2992_bF_buf5), .B(a_reg_10_), .Y(_abc_15724_n4592) );
  AND2X2 AND2X2_194 ( .A(_abc_15724_n907_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_39_), .Y(_abc_15724_n1099) );
  AND2X2 AND2X2_1940 ( .A(_abc_15724_n906_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_138_), .Y(_abc_15724_n4593) );
  AND2X2 AND2X2_1941 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n4593), .Y(_abc_15724_n4594) );
  AND2X2 AND2X2_1942 ( .A(_abc_15724_n4588), .B(_abc_15724_n4597), .Y(_abc_15724_n4598) );
  AND2X2 AND2X2_1943 ( .A(_abc_15724_n4602), .B(_abc_15724_n4603), .Y(_abc_15724_n4604) );
  AND2X2 AND2X2_1944 ( .A(c_reg_11_), .B(b_reg_11_), .Y(_abc_15724_n4605) );
  AND2X2 AND2X2_1945 ( .A(_abc_15724_n4606), .B(_abc_15724_n4601), .Y(_abc_15724_n4607) );
  AND2X2 AND2X2_1946 ( .A(_abc_15724_n4608), .B(_abc_15724_n4609), .Y(_abc_15724_n4610) );
  AND2X2 AND2X2_1947 ( .A(_abc_15724_n3726_bF_buf1), .B(_abc_15724_n4610), .Y(_abc_15724_n4611) );
  AND2X2 AND2X2_1948 ( .A(_abc_15724_n4601), .B(_abc_15724_n4603), .Y(_abc_15724_n4612) );
  AND2X2 AND2X2_1949 ( .A(_abc_15724_n4602), .B(b_reg_11_), .Y(_abc_15724_n4613) );
  AND2X2 AND2X2_195 ( .A(_auto_iopadmap_cc_313_execute_26059_39_), .B(d_reg_7_), .Y(_abc_15724_n1101) );
  AND2X2 AND2X2_1950 ( .A(_abc_15724_n4616), .B(_abc_15724_n4601), .Y(_abc_15724_n4617) );
  AND2X2 AND2X2_1951 ( .A(_abc_15724_n4619), .B(_abc_15724_n4615), .Y(_abc_15724_n4620) );
  AND2X2 AND2X2_1952 ( .A(_abc_15724_n4553), .B(_abc_15724_n4550), .Y(_abc_15724_n4623) );
  AND2X2 AND2X2_1953 ( .A(a_reg_6_), .B(e_reg_11_), .Y(_abc_15724_n4626) );
  AND2X2 AND2X2_1954 ( .A(_abc_15724_n4627), .B(_abc_15724_n4625), .Y(_abc_15724_n4628) );
  AND2X2 AND2X2_1955 ( .A(_abc_15724_n4628), .B(w_11_), .Y(_abc_15724_n4629) );
  AND2X2 AND2X2_1956 ( .A(_abc_15724_n4630), .B(_abc_15724_n4631), .Y(_abc_15724_n4632) );
  AND2X2 AND2X2_1957 ( .A(_abc_15724_n4624), .B(_abc_15724_n4632), .Y(_abc_15724_n4633) );
  AND2X2 AND2X2_1958 ( .A(_abc_15724_n4634), .B(_abc_15724_n4635), .Y(_abc_15724_n4636) );
  AND2X2 AND2X2_1959 ( .A(_abc_15724_n4638), .B(_abc_15724_n4620), .Y(_abc_15724_n4639) );
  AND2X2 AND2X2_196 ( .A(_abc_15724_n1102), .B(_abc_15724_n1100), .Y(_abc_15724_n1103) );
  AND2X2 AND2X2_1960 ( .A(_abc_15724_n4642), .B(_abc_15724_n4637), .Y(_abc_15724_n4643) );
  AND2X2 AND2X2_1961 ( .A(_abc_15724_n4643), .B(_abc_15724_n4600), .Y(_abc_15724_n4644) );
  AND2X2 AND2X2_1962 ( .A(_abc_15724_n4570), .B(_abc_15724_n4563), .Y(_abc_15724_n4645) );
  AND2X2 AND2X2_1963 ( .A(_abc_15724_n4641), .B(_abc_15724_n4639), .Y(_abc_15724_n4646) );
  AND2X2 AND2X2_1964 ( .A(_abc_15724_n4622), .B(_abc_15724_n4636), .Y(_abc_15724_n4647) );
  AND2X2 AND2X2_1965 ( .A(_abc_15724_n4648), .B(_abc_15724_n4645), .Y(_abc_15724_n4649) );
  AND2X2 AND2X2_1966 ( .A(_abc_15724_n4652), .B(_abc_15724_n4653), .Y(_abc_15724_n4654) );
  AND2X2 AND2X2_1967 ( .A(_abc_15724_n4651), .B(_abc_15724_n4655), .Y(_abc_15724_n4656) );
  AND2X2 AND2X2_1968 ( .A(_abc_15724_n4656), .B(_abc_15724_n4599), .Y(_abc_15724_n4657) );
  AND2X2 AND2X2_1969 ( .A(_abc_15724_n4578), .B(_abc_15724_n4567), .Y(_abc_15724_n4658) );
  AND2X2 AND2X2_197 ( .A(_abc_15724_n1085), .B(_abc_15724_n1089), .Y(_abc_15724_n1104) );
  AND2X2 AND2X2_1970 ( .A(_abc_15724_n4654), .B(_abc_15724_n3736), .Y(_abc_15724_n4659) );
  AND2X2 AND2X2_1971 ( .A(_abc_15724_n4650), .B(_abc_15724_n3724), .Y(_abc_15724_n4660) );
  AND2X2 AND2X2_1972 ( .A(_abc_15724_n4661), .B(_abc_15724_n4658), .Y(_abc_15724_n4662) );
  AND2X2 AND2X2_1973 ( .A(_abc_15724_n4667), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n4668) );
  AND2X2 AND2X2_1974 ( .A(_abc_15724_n4668), .B(_abc_15724_n4664), .Y(_abc_15724_n4669) );
  AND2X2 AND2X2_1975 ( .A(_abc_15724_n2992_bF_buf4), .B(a_reg_11_), .Y(_abc_15724_n4670) );
  AND2X2 AND2X2_1976 ( .A(_abc_15724_n906_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_139_), .Y(_abc_15724_n4671) );
  AND2X2 AND2X2_1977 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n4671), .Y(_abc_15724_n4672) );
  AND2X2 AND2X2_1978 ( .A(_abc_15724_n4680), .B(_abc_15724_n4679), .Y(_abc_15724_n4681) );
  AND2X2 AND2X2_1979 ( .A(_abc_15724_n4682), .B(_abc_15724_n4681), .Y(_abc_15724_n4683) );
  AND2X2 AND2X2_198 ( .A(_abc_15724_n1093), .B(_abc_15724_n1088), .Y(_abc_15724_n1108) );
  AND2X2 AND2X2_1980 ( .A(_abc_15724_n4678), .B(_abc_15724_n4683), .Y(_abc_15724_n4684) );
  AND2X2 AND2X2_1981 ( .A(_abc_15724_n4651), .B(_abc_15724_n4652), .Y(_abc_15724_n4686) );
  AND2X2 AND2X2_1982 ( .A(_abc_15724_n4689), .B(_abc_15724_n4690), .Y(_abc_15724_n4691) );
  AND2X2 AND2X2_1983 ( .A(c_reg_12_), .B(b_reg_12_), .Y(_abc_15724_n4692) );
  AND2X2 AND2X2_1984 ( .A(_abc_15724_n4693), .B(_abc_15724_n4688), .Y(_abc_15724_n4694) );
  AND2X2 AND2X2_1985 ( .A(_abc_15724_n4695), .B(_abc_15724_n4696), .Y(_abc_15724_n4697) );
  AND2X2 AND2X2_1986 ( .A(_abc_15724_n3726_bF_buf0), .B(_abc_15724_n4697), .Y(_abc_15724_n4698) );
  AND2X2 AND2X2_1987 ( .A(_abc_15724_n4688), .B(_abc_15724_n4690), .Y(_abc_15724_n4700) );
  AND2X2 AND2X2_1988 ( .A(_abc_15724_n4689), .B(b_reg_12_), .Y(_abc_15724_n4701) );
  AND2X2 AND2X2_1989 ( .A(_abc_15724_n4704), .B(_abc_15724_n4688), .Y(_abc_15724_n4705) );
  AND2X2 AND2X2_199 ( .A(_abc_15724_n1109_1), .B(_abc_15724_n1106), .Y(_abc_15724_n1110_1) );
  AND2X2 AND2X2_1990 ( .A(_abc_15724_n4707), .B(_abc_15724_n4703), .Y(_abc_15724_n4708) );
  AND2X2 AND2X2_1991 ( .A(_abc_15724_n4699), .B(_abc_15724_n4708), .Y(_abc_15724_n4709) );
  AND2X2 AND2X2_1992 ( .A(_abc_15724_n4630), .B(_abc_15724_n4627), .Y(_abc_15724_n4711) );
  AND2X2 AND2X2_1993 ( .A(a_reg_7_), .B(e_reg_12_), .Y(_abc_15724_n4714) );
  AND2X2 AND2X2_1994 ( .A(_abc_15724_n4715), .B(_abc_15724_n4713), .Y(_abc_15724_n4716) );
  AND2X2 AND2X2_1995 ( .A(_abc_15724_n4716), .B(w_12_), .Y(_abc_15724_n4717) );
  AND2X2 AND2X2_1996 ( .A(_abc_15724_n4718), .B(_abc_15724_n4719), .Y(_abc_15724_n4720) );
  AND2X2 AND2X2_1997 ( .A(_abc_15724_n4712), .B(_abc_15724_n4720), .Y(_abc_15724_n4721) );
  AND2X2 AND2X2_1998 ( .A(_abc_15724_n4722), .B(_abc_15724_n4723), .Y(_abc_15724_n4724) );
  AND2X2 AND2X2_1999 ( .A(_abc_15724_n4725), .B(_abc_15724_n4728), .Y(_abc_15724_n4729) );
  AND2X2 AND2X2_2 ( .A(_auto_iopadmap_cc_313_execute_26059_20_), .B(e_reg_20_), .Y(_abc_15724_n699) );
  AND2X2 AND2X2_20 ( .A(_abc_15724_n732), .B(_abc_15724_n736), .Y(_abc_15724_n737) );
  AND2X2 AND2X2_200 ( .A(_abc_15724_n1110_1), .B(digest_update_bF_buf5), .Y(_abc_15724_n1111_1) );
  AND2X2 AND2X2_2000 ( .A(_abc_15724_n4729), .B(_abc_15724_n4687), .Y(_abc_15724_n4730) );
  AND2X2 AND2X2_2001 ( .A(_abc_15724_n4642), .B(_abc_15724_n4634), .Y(_abc_15724_n4731) );
  AND2X2 AND2X2_2002 ( .A(_abc_15724_n4727), .B(_abc_15724_n4709), .Y(_abc_15724_n4732) );
  AND2X2 AND2X2_2003 ( .A(_abc_15724_n4710), .B(_abc_15724_n4724), .Y(_abc_15724_n4733) );
  AND2X2 AND2X2_2004 ( .A(_abc_15724_n4734), .B(_abc_15724_n4731), .Y(_abc_15724_n4735) );
  AND2X2 AND2X2_2005 ( .A(_abc_15724_n4736), .B(_abc_15724_n3726_bF_buf4), .Y(_abc_15724_n4737) );
  AND2X2 AND2X2_2006 ( .A(_abc_15724_n4739), .B(_abc_15724_n4738), .Y(_abc_15724_n4740) );
  AND2X2 AND2X2_2007 ( .A(_abc_15724_n4740), .B(_abc_15724_n3806_bF_buf1), .Y(_abc_15724_n4741) );
  AND2X2 AND2X2_2008 ( .A(_abc_15724_n4742), .B(_abc_15724_n4686), .Y(_abc_15724_n4745) );
  AND2X2 AND2X2_2009 ( .A(_abc_15724_n4685), .B(_abc_15724_n4747), .Y(_abc_15724_n4749) );
  AND2X2 AND2X2_201 ( .A(_abc_15724_n907_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_40_), .Y(_abc_15724_n1113) );
  AND2X2 AND2X2_2010 ( .A(_abc_15724_n4750), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n4751) );
  AND2X2 AND2X2_2011 ( .A(_abc_15724_n4751), .B(_abc_15724_n4748), .Y(_abc_15724_n4752) );
  AND2X2 AND2X2_2012 ( .A(_abc_15724_n2992_bF_buf3), .B(a_reg_12_), .Y(_abc_15724_n4753) );
  AND2X2 AND2X2_2013 ( .A(_abc_15724_n906_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_140_), .Y(_abc_15724_n4754) );
  AND2X2 AND2X2_2014 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n4754), .Y(_abc_15724_n4755) );
  AND2X2 AND2X2_2015 ( .A(_abc_15724_n4728), .B(_abc_15724_n4722), .Y(_abc_15724_n4759) );
  AND2X2 AND2X2_2016 ( .A(_abc_15724_n4761), .B(_abc_15724_n4762), .Y(_abc_15724_n4763) );
  AND2X2 AND2X2_2017 ( .A(c_reg_13_), .B(b_reg_13_), .Y(_abc_15724_n4764) );
  AND2X2 AND2X2_2018 ( .A(_abc_15724_n4765), .B(_abc_15724_n4760), .Y(_abc_15724_n4766) );
  AND2X2 AND2X2_2019 ( .A(_abc_15724_n4767), .B(_abc_15724_n4768), .Y(_abc_15724_n4769) );
  AND2X2 AND2X2_202 ( .A(_abc_15724_n1105), .B(_abc_15724_n1103), .Y(_abc_15724_n1114) );
  AND2X2 AND2X2_2020 ( .A(_abc_15724_n3726_bF_buf3), .B(_abc_15724_n4769), .Y(_abc_15724_n4770) );
  AND2X2 AND2X2_2021 ( .A(_abc_15724_n4760), .B(_abc_15724_n4762), .Y(_abc_15724_n4772) );
  AND2X2 AND2X2_2022 ( .A(_abc_15724_n4761), .B(b_reg_13_), .Y(_abc_15724_n4773) );
  AND2X2 AND2X2_2023 ( .A(_abc_15724_n4776), .B(_abc_15724_n4760), .Y(_abc_15724_n4777) );
  AND2X2 AND2X2_2024 ( .A(_abc_15724_n4779), .B(_abc_15724_n4775), .Y(_abc_15724_n4780) );
  AND2X2 AND2X2_2025 ( .A(_abc_15724_n4771), .B(_abc_15724_n4780), .Y(_abc_15724_n4781) );
  AND2X2 AND2X2_2026 ( .A(_abc_15724_n4718), .B(_abc_15724_n4715), .Y(_abc_15724_n4782) );
  AND2X2 AND2X2_2027 ( .A(a_reg_8_), .B(e_reg_13_), .Y(_abc_15724_n4785) );
  AND2X2 AND2X2_2028 ( .A(_abc_15724_n4786), .B(_abc_15724_n4784), .Y(_abc_15724_n4787) );
  AND2X2 AND2X2_2029 ( .A(_abc_15724_n4787), .B(w_13_), .Y(_abc_15724_n4788) );
  AND2X2 AND2X2_203 ( .A(_auto_iopadmap_cc_313_execute_26059_40_), .B(d_reg_8_), .Y(_abc_15724_n1117) );
  AND2X2 AND2X2_2030 ( .A(_abc_15724_n4789), .B(_abc_15724_n4790), .Y(_abc_15724_n4791) );
  AND2X2 AND2X2_2031 ( .A(_abc_15724_n4783), .B(_abc_15724_n4791), .Y(_abc_15724_n4792) );
  AND2X2 AND2X2_2032 ( .A(_abc_15724_n4795), .B(_abc_15724_n4781), .Y(_abc_15724_n4796) );
  AND2X2 AND2X2_2033 ( .A(_abc_15724_n4798), .B(_abc_15724_n4793), .Y(_abc_15724_n4799) );
  AND2X2 AND2X2_2034 ( .A(_abc_15724_n4797), .B(_abc_15724_n4799), .Y(_abc_15724_n4800) );
  AND2X2 AND2X2_2035 ( .A(_abc_15724_n4804), .B(_abc_15724_n4805), .Y(_abc_15724_n4806) );
  AND2X2 AND2X2_2036 ( .A(_abc_15724_n4807), .B(_abc_15724_n4802), .Y(_abc_15724_n4808) );
  AND2X2 AND2X2_2037 ( .A(_abc_15724_n4803), .B(_abc_15724_n4806), .Y(_abc_15724_n4810) );
  AND2X2 AND2X2_2038 ( .A(_abc_15724_n4801), .B(_abc_15724_n4759), .Y(_abc_15724_n4811) );
  AND2X2 AND2X2_2039 ( .A(_abc_15724_n4813), .B(_abc_15724_n4809), .Y(_abc_15724_n4814) );
  AND2X2 AND2X2_204 ( .A(_abc_15724_n1118), .B(_abc_15724_n1116), .Y(_abc_15724_n1119_1) );
  AND2X2 AND2X2_2040 ( .A(_abc_15724_n4814), .B(_abc_15724_n4758), .Y(_abc_15724_n4815) );
  AND2X2 AND2X2_2041 ( .A(_abc_15724_n4816), .B(_abc_15724_n4738), .Y(_abc_15724_n4817) );
  AND2X2 AND2X2_2042 ( .A(_abc_15724_n4812), .B(_abc_15724_n3724), .Y(_abc_15724_n4818) );
  AND2X2 AND2X2_2043 ( .A(_abc_15724_n4808), .B(_abc_15724_n3736), .Y(_abc_15724_n4819) );
  AND2X2 AND2X2_2044 ( .A(_abc_15724_n4820), .B(_abc_15724_n4817), .Y(_abc_15724_n4821) );
  AND2X2 AND2X2_2045 ( .A(_abc_15724_n4685), .B(_abc_15724_n4827), .Y(_abc_15724_n4828) );
  AND2X2 AND2X2_2046 ( .A(_abc_15724_n4830), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n4831) );
  AND2X2 AND2X2_2047 ( .A(_abc_15724_n4829), .B(_abc_15724_n4831), .Y(_abc_15724_n4832) );
  AND2X2 AND2X2_2048 ( .A(_abc_15724_n4832), .B(_abc_15724_n4825), .Y(_abc_15724_n4833) );
  AND2X2 AND2X2_2049 ( .A(_abc_15724_n2992_bF_buf2), .B(a_reg_13_), .Y(_abc_15724_n4834) );
  AND2X2 AND2X2_205 ( .A(_abc_15724_n1115), .B(_abc_15724_n1119_1), .Y(_abc_15724_n1121_1) );
  AND2X2 AND2X2_2050 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n2686), .Y(_abc_15724_n4835) );
  AND2X2 AND2X2_2051 ( .A(_abc_15724_n4830), .B(_abc_15724_n4838), .Y(_abc_15724_n4839) );
  AND2X2 AND2X2_2052 ( .A(_abc_15724_n4829), .B(_abc_15724_n4839), .Y(_abc_15724_n4840) );
  AND2X2 AND2X2_2053 ( .A(_abc_15724_n4813), .B(_abc_15724_n4802), .Y(_abc_15724_n4842) );
  AND2X2 AND2X2_2054 ( .A(_abc_15724_n4805), .B(_abc_15724_n4798), .Y(_abc_15724_n4844) );
  AND2X2 AND2X2_2055 ( .A(_abc_15724_n4846), .B(_abc_15724_n4847), .Y(_abc_15724_n4848) );
  AND2X2 AND2X2_2056 ( .A(c_reg_14_), .B(b_reg_14_), .Y(_abc_15724_n4849) );
  AND2X2 AND2X2_2057 ( .A(_abc_15724_n4850), .B(_abc_15724_n4845), .Y(_abc_15724_n4851) );
  AND2X2 AND2X2_2058 ( .A(_abc_15724_n4852), .B(_abc_15724_n4845), .Y(_abc_15724_n4853) );
  AND2X2 AND2X2_2059 ( .A(_abc_15724_n4855), .B(_abc_15724_n4852), .Y(_abc_15724_n4856) );
  AND2X2 AND2X2_206 ( .A(_abc_15724_n1122), .B(_abc_15724_n1120_1), .Y(_abc_15724_n1123) );
  AND2X2 AND2X2_2060 ( .A(_abc_15724_n4846), .B(b_reg_14_), .Y(_abc_15724_n4859) );
  AND2X2 AND2X2_2061 ( .A(_abc_15724_n3737_bF_buf4), .B(_abc_15724_n4855), .Y(_abc_15724_n4862) );
  AND2X2 AND2X2_2062 ( .A(_abc_15724_n4863), .B(_abc_15724_n4861), .Y(_abc_15724_n4864) );
  AND2X2 AND2X2_2063 ( .A(_abc_15724_n4858), .B(_abc_15724_n4864), .Y(_abc_15724_n4865) );
  AND2X2 AND2X2_2064 ( .A(_abc_15724_n4789), .B(_abc_15724_n4786), .Y(_abc_15724_n4866) );
  AND2X2 AND2X2_2065 ( .A(a_reg_9_), .B(e_reg_14_), .Y(_abc_15724_n4869) );
  AND2X2 AND2X2_2066 ( .A(_abc_15724_n4870), .B(_abc_15724_n4868), .Y(_abc_15724_n4871) );
  AND2X2 AND2X2_2067 ( .A(_abc_15724_n4871), .B(w_14_), .Y(_abc_15724_n4872) );
  AND2X2 AND2X2_2068 ( .A(_abc_15724_n4873), .B(_abc_15724_n4874), .Y(_abc_15724_n4875) );
  AND2X2 AND2X2_2069 ( .A(_abc_15724_n4867), .B(_abc_15724_n4875), .Y(_abc_15724_n4876) );
  AND2X2 AND2X2_207 ( .A(_abc_15724_n1123), .B(digest_update_bF_buf4), .Y(_abc_15724_n1124) );
  AND2X2 AND2X2_2070 ( .A(_abc_15724_n4877), .B(_abc_15724_n4878), .Y(_abc_15724_n4879) );
  AND2X2 AND2X2_2071 ( .A(_abc_15724_n4880), .B(_abc_15724_n4865), .Y(_abc_15724_n4881) );
  AND2X2 AND2X2_2072 ( .A(_abc_15724_n4887), .B(_abc_15724_n4882), .Y(_abc_15724_n4888) );
  AND2X2 AND2X2_2073 ( .A(_abc_15724_n4885), .B(_abc_15724_n4889), .Y(_abc_15724_n4890) );
  AND2X2 AND2X2_2074 ( .A(_abc_15724_n4888), .B(_abc_15724_n4886), .Y(_abc_15724_n4892) );
  AND2X2 AND2X2_2075 ( .A(_abc_15724_n4884), .B(_abc_15724_n4844), .Y(_abc_15724_n4893) );
  AND2X2 AND2X2_2076 ( .A(_abc_15724_n4895), .B(_abc_15724_n4891), .Y(_abc_15724_n4896) );
  AND2X2 AND2X2_2077 ( .A(_abc_15724_n4896), .B(_abc_15724_n4843), .Y(_abc_15724_n4897) );
  AND2X2 AND2X2_2078 ( .A(_abc_15724_n4894), .B(_abc_15724_n3737_bF_buf2), .Y(_abc_15724_n4898) );
  AND2X2 AND2X2_2079 ( .A(_abc_15724_n4890), .B(_abc_15724_n3725_bF_buf2), .Y(_abc_15724_n4899) );
  AND2X2 AND2X2_208 ( .A(_auto_iopadmap_cc_313_execute_26059_41_), .B(d_reg_9_), .Y(_abc_15724_n1127) );
  AND2X2 AND2X2_2080 ( .A(_abc_15724_n4900), .B(_abc_15724_n4842), .Y(_abc_15724_n4901) );
  AND2X2 AND2X2_2081 ( .A(_abc_15724_n4841), .B(_abc_15724_n4903), .Y(_abc_15724_n4904) );
  AND2X2 AND2X2_2082 ( .A(_abc_15724_n4906), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n4907) );
  AND2X2 AND2X2_2083 ( .A(_abc_15724_n4907), .B(_abc_15724_n4905), .Y(_abc_15724_n4908) );
  AND2X2 AND2X2_2084 ( .A(_abc_15724_n2992_bF_buf1), .B(a_reg_14_), .Y(_abc_15724_n4909) );
  AND2X2 AND2X2_2085 ( .A(_abc_15724_n906_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_142_), .Y(_abc_15724_n4910) );
  AND2X2 AND2X2_2086 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n4910), .Y(_abc_15724_n4911) );
  AND2X2 AND2X2_2087 ( .A(_abc_15724_n4905), .B(_abc_15724_n4914), .Y(_abc_15724_n4915) );
  AND2X2 AND2X2_2088 ( .A(_abc_15724_n4882), .B(_abc_15724_n4877), .Y(_abc_15724_n4918) );
  AND2X2 AND2X2_2089 ( .A(c_reg_15_), .B(b_reg_15_), .Y(_abc_15724_n4920) );
  AND2X2 AND2X2_209 ( .A(_abc_15724_n1128), .B(_abc_15724_n1126), .Y(_abc_15724_n1129) );
  AND2X2 AND2X2_2090 ( .A(_abc_15724_n4923), .B(_abc_15724_n4921), .Y(_abc_15724_n4924) );
  AND2X2 AND2X2_2091 ( .A(_abc_15724_n3805_bF_buf3), .B(_abc_15724_n4924), .Y(_abc_15724_n4925) );
  AND2X2 AND2X2_2092 ( .A(_abc_15724_n4921), .B(_abc_15724_n4926), .Y(_abc_15724_n4927) );
  AND2X2 AND2X2_2093 ( .A(_abc_15724_n4927), .B(d_reg_15_), .Y(_abc_15724_n4929) );
  AND2X2 AND2X2_2094 ( .A(_abc_15724_n4930), .B(_abc_15724_n4928), .Y(_abc_15724_n4931) );
  AND2X2 AND2X2_2095 ( .A(_abc_15724_n3726_bF_buf1), .B(_abc_15724_n4931), .Y(_abc_15724_n4932) );
  AND2X2 AND2X2_2096 ( .A(_abc_15724_n4921), .B(_abc_15724_n4922), .Y(_abc_15724_n4934) );
  AND2X2 AND2X2_2097 ( .A(_abc_15724_n4937), .B(_abc_15724_n3721_bF_buf1), .Y(_abc_15724_n4938) );
  AND2X2 AND2X2_2098 ( .A(_abc_15724_n4933), .B(_abc_15724_n4938), .Y(_abc_15724_n4939) );
  AND2X2 AND2X2_2099 ( .A(a_reg_10_), .B(e_reg_15_), .Y(_abc_15724_n4943) );
  AND2X2 AND2X2_21 ( .A(_auto_iopadmap_cc_313_execute_26059_13_), .B(e_reg_13_), .Y(_abc_15724_n739_1) );
  AND2X2 AND2X2_210 ( .A(_abc_15724_n1122), .B(_abc_15724_n1118), .Y(_abc_15724_n1130) );
  AND2X2 AND2X2_2100 ( .A(_abc_15724_n4944), .B(_abc_15724_n4942), .Y(_abc_15724_n4945) );
  AND2X2 AND2X2_2101 ( .A(_abc_15724_n4945), .B(w_15_), .Y(_abc_15724_n4946) );
  AND2X2 AND2X2_2102 ( .A(_abc_15724_n4947), .B(_abc_15724_n4948), .Y(_abc_15724_n4949) );
  AND2X2 AND2X2_2103 ( .A(_abc_15724_n4949), .B(_abc_15724_n4941), .Y(_abc_15724_n4950) );
  AND2X2 AND2X2_2104 ( .A(_abc_15724_n4951), .B(_abc_15724_n4952), .Y(_abc_15724_n4953) );
  AND2X2 AND2X2_2105 ( .A(_abc_15724_n4958), .B(_abc_15724_n4956), .Y(_abc_15724_n4959) );
  AND2X2 AND2X2_2106 ( .A(_abc_15724_n4960), .B(_abc_15724_n4955), .Y(_abc_15724_n4961) );
  AND2X2 AND2X2_2107 ( .A(_abc_15724_n4961), .B(_abc_15724_n4919), .Y(_abc_15724_n4962) );
  AND2X2 AND2X2_2108 ( .A(_abc_15724_n4959), .B(_abc_15724_n4953), .Y(_abc_15724_n4963) );
  AND2X2 AND2X2_2109 ( .A(_abc_15724_n4940), .B(_abc_15724_n4954), .Y(_abc_15724_n4964) );
  AND2X2 AND2X2_211 ( .A(_abc_15724_n1131_1), .B(_abc_15724_n1129), .Y(_abc_15724_n1133_1) );
  AND2X2 AND2X2_2110 ( .A(_abc_15724_n4965), .B(_abc_15724_n4918), .Y(_abc_15724_n4966) );
  AND2X2 AND2X2_2111 ( .A(_abc_15724_n4970), .B(_abc_15724_n4969), .Y(_abc_15724_n4971) );
  AND2X2 AND2X2_2112 ( .A(_abc_15724_n4968), .B(_abc_15724_n4972), .Y(_abc_15724_n4973) );
  AND2X2 AND2X2_2113 ( .A(_abc_15724_n4917), .B(_abc_15724_n4973), .Y(_abc_15724_n4974) );
  AND2X2 AND2X2_2114 ( .A(_abc_15724_n4895), .B(_abc_15724_n4885), .Y(_abc_15724_n4975) );
  AND2X2 AND2X2_2115 ( .A(_abc_15724_n4971), .B(_abc_15724_n3721_bF_buf4), .Y(_abc_15724_n4976) );
  AND2X2 AND2X2_2116 ( .A(_abc_15724_n4967), .B(_abc_15724_n3805_bF_buf1), .Y(_abc_15724_n4977) );
  AND2X2 AND2X2_2117 ( .A(_abc_15724_n4978), .B(_abc_15724_n4975), .Y(_abc_15724_n4979) );
  AND2X2 AND2X2_2118 ( .A(_abc_15724_n4983), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n4984) );
  AND2X2 AND2X2_2119 ( .A(_abc_15724_n4984), .B(_abc_15724_n4982), .Y(_abc_15724_n4985) );
  AND2X2 AND2X2_212 ( .A(_abc_15724_n1134), .B(_abc_15724_n1132_1), .Y(_abc_15724_n1135) );
  AND2X2 AND2X2_2120 ( .A(_abc_15724_n2992_bF_buf0), .B(a_reg_15_), .Y(_abc_15724_n4986) );
  AND2X2 AND2X2_2121 ( .A(_abc_15724_n906_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_143_), .Y(_abc_15724_n4987) );
  AND2X2 AND2X2_2122 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n4987), .Y(_abc_15724_n4988) );
  AND2X2 AND2X2_2123 ( .A(_abc_15724_n4996), .B(_abc_15724_n4897), .Y(_abc_15724_n4997) );
  AND2X2 AND2X2_2124 ( .A(_abc_15724_n4995), .B(_abc_15724_n4999), .Y(_abc_15724_n5000) );
  AND2X2 AND2X2_2125 ( .A(_abc_15724_n5001), .B(_abc_15724_n5000), .Y(_abc_15724_n5002) );
  AND2X2 AND2X2_2126 ( .A(_abc_15724_n4994), .B(_abc_15724_n5002), .Y(_abc_15724_n5003) );
  AND2X2 AND2X2_2127 ( .A(_abc_15724_n4968), .B(_abc_15724_n4969), .Y(_abc_15724_n5005) );
  AND2X2 AND2X2_2128 ( .A(_abc_15724_n4022), .B(_abc_15724_n3725_bF_buf0), .Y(_abc_15724_n5006) );
  AND2X2 AND2X2_2129 ( .A(_abc_15724_n4955), .B(_abc_15724_n4951), .Y(_abc_15724_n5007) );
  AND2X2 AND2X2_213 ( .A(_abc_15724_n1135), .B(digest_update_bF_buf3), .Y(_abc_15724_n1136) );
  AND2X2 AND2X2_2130 ( .A(_abc_15724_n5009), .B(_abc_15724_n5010), .Y(_abc_15724_n5011) );
  AND2X2 AND2X2_2131 ( .A(c_reg_16_), .B(b_reg_16_), .Y(_abc_15724_n5013) );
  AND2X2 AND2X2_2132 ( .A(_abc_15724_n5012), .B(_abc_15724_n5014), .Y(_abc_15724_n5015) );
  AND2X2 AND2X2_2133 ( .A(_abc_15724_n5012), .B(_abc_15724_n5017), .Y(_abc_15724_n5018) );
  AND2X2 AND2X2_2134 ( .A(_abc_15724_n5018), .B(_abc_15724_n5014), .Y(_abc_15724_n5019) );
  AND2X2 AND2X2_2135 ( .A(_abc_15724_n5020), .B(_abc_15724_n5016), .Y(_abc_15724_n5021) );
  AND2X2 AND2X2_2136 ( .A(_abc_15724_n5021), .B(_abc_15724_n3726_bF_buf0), .Y(_abc_15724_n5022) );
  AND2X2 AND2X2_2137 ( .A(_abc_15724_n5009), .B(b_reg_16_), .Y(_abc_15724_n5025) );
  AND2X2 AND2X2_2138 ( .A(_abc_15724_n3737_bF_buf1), .B(_abc_15724_n5018), .Y(_abc_15724_n5028) );
  AND2X2 AND2X2_2139 ( .A(_abc_15724_n5029), .B(_abc_15724_n5027), .Y(_abc_15724_n5030) );
  AND2X2 AND2X2_214 ( .A(_abc_15724_n907_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_41_), .Y(_abc_15724_n1137) );
  AND2X2 AND2X2_2140 ( .A(_abc_15724_n5023), .B(_abc_15724_n5030), .Y(_abc_15724_n5031) );
  AND2X2 AND2X2_2141 ( .A(_abc_15724_n4947), .B(_abc_15724_n4944), .Y(_abc_15724_n5032) );
  AND2X2 AND2X2_2142 ( .A(a_reg_11_), .B(e_reg_16_), .Y(_abc_15724_n5035) );
  AND2X2 AND2X2_2143 ( .A(_abc_15724_n5036), .B(_abc_15724_n5034), .Y(_abc_15724_n5037) );
  AND2X2 AND2X2_2144 ( .A(_abc_15724_n5037), .B(w_16_), .Y(_abc_15724_n5038) );
  AND2X2 AND2X2_2145 ( .A(_abc_15724_n5039), .B(_abc_15724_n5040), .Y(_abc_15724_n5041) );
  AND2X2 AND2X2_2146 ( .A(_abc_15724_n5033), .B(_abc_15724_n5041), .Y(_abc_15724_n5042) );
  AND2X2 AND2X2_2147 ( .A(_abc_15724_n5043), .B(_abc_15724_n5044), .Y(_abc_15724_n5045) );
  AND2X2 AND2X2_2148 ( .A(_abc_15724_n5046), .B(_abc_15724_n5031), .Y(_abc_15724_n5047) );
  AND2X2 AND2X2_2149 ( .A(_abc_15724_n5051), .B(_abc_15724_n5008), .Y(_abc_15724_n5052) );
  AND2X2 AND2X2_215 ( .A(_abc_15724_n1134), .B(_abc_15724_n1128), .Y(_abc_15724_n1139) );
  AND2X2 AND2X2_2150 ( .A(_abc_15724_n5050), .B(_abc_15724_n5007), .Y(_abc_15724_n5053) );
  AND2X2 AND2X2_2151 ( .A(_abc_15724_n5054), .B(_abc_15724_n5006), .Y(_abc_15724_n5055) );
  AND2X2 AND2X2_2152 ( .A(_abc_15724_n5057), .B(_abc_15724_n5056), .Y(_abc_15724_n5058) );
  AND2X2 AND2X2_2153 ( .A(_abc_15724_n5059), .B(_abc_15724_n5005), .Y(_abc_15724_n5062) );
  AND2X2 AND2X2_2154 ( .A(_abc_15724_n5004), .B(_abc_15724_n5064), .Y(_abc_15724_n5066) );
  AND2X2 AND2X2_2155 ( .A(_abc_15724_n5067), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n5068) );
  AND2X2 AND2X2_2156 ( .A(_abc_15724_n5068), .B(_abc_15724_n5065), .Y(_abc_15724_n5069) );
  AND2X2 AND2X2_2157 ( .A(_abc_15724_n2992_bF_buf11), .B(a_reg_16_), .Y(_abc_15724_n5070) );
  AND2X2 AND2X2_2158 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n2741), .Y(_abc_15724_n5071) );
  AND2X2 AND2X2_2159 ( .A(_abc_15724_n5075), .B(_abc_15724_n5074), .Y(_abc_15724_n5076) );
  AND2X2 AND2X2_216 ( .A(_auto_iopadmap_cc_313_execute_26059_42_), .B(d_reg_10_), .Y(_abc_15724_n1142_1) );
  AND2X2 AND2X2_2160 ( .A(_abc_15724_n5048), .B(_abc_15724_n5043), .Y(_abc_15724_n5077) );
  AND2X2 AND2X2_2161 ( .A(c_reg_17_), .B(b_reg_17_), .Y(_abc_15724_n5079) );
  AND2X2 AND2X2_2162 ( .A(_abc_15724_n5082), .B(_abc_15724_n5080), .Y(_abc_15724_n5083) );
  AND2X2 AND2X2_2163 ( .A(_abc_15724_n3805_bF_buf0), .B(_abc_15724_n5083), .Y(_abc_15724_n5084) );
  AND2X2 AND2X2_2164 ( .A(_abc_15724_n5080), .B(_abc_15724_n5086), .Y(_abc_15724_n5087) );
  AND2X2 AND2X2_2165 ( .A(_abc_15724_n5087), .B(d_reg_17_), .Y(_abc_15724_n5089) );
  AND2X2 AND2X2_2166 ( .A(_abc_15724_n5090), .B(_abc_15724_n5088), .Y(_abc_15724_n5091) );
  AND2X2 AND2X2_2167 ( .A(_abc_15724_n3726_bF_buf4), .B(_abc_15724_n5091), .Y(_abc_15724_n5092) );
  AND2X2 AND2X2_2168 ( .A(_abc_15724_n5093), .B(_abc_15724_n5086), .Y(_abc_15724_n5094) );
  AND2X2 AND2X2_2169 ( .A(_abc_15724_n3737_bF_buf0), .B(_abc_15724_n5094), .Y(_abc_15724_n5095) );
  AND2X2 AND2X2_217 ( .A(_abc_15724_n1143), .B(_abc_15724_n1141_1), .Y(_abc_15724_n1144_1) );
  AND2X2 AND2X2_2170 ( .A(_abc_15724_n5097), .B(_abc_15724_n5085), .Y(_abc_15724_n5098) );
  AND2X2 AND2X2_2171 ( .A(_abc_15724_n5039), .B(_abc_15724_n5036), .Y(_abc_15724_n5099) );
  AND2X2 AND2X2_2172 ( .A(a_reg_12_), .B(e_reg_17_), .Y(_abc_15724_n5102) );
  AND2X2 AND2X2_2173 ( .A(_abc_15724_n5103), .B(_abc_15724_n5101), .Y(_abc_15724_n5104) );
  AND2X2 AND2X2_2174 ( .A(_abc_15724_n5104), .B(w_17_), .Y(_abc_15724_n5105) );
  AND2X2 AND2X2_2175 ( .A(_abc_15724_n5106), .B(_abc_15724_n5107), .Y(_abc_15724_n5108) );
  AND2X2 AND2X2_2176 ( .A(_abc_15724_n5100), .B(_abc_15724_n5108), .Y(_abc_15724_n5109) );
  AND2X2 AND2X2_2177 ( .A(_abc_15724_n5110), .B(_abc_15724_n5111), .Y(_abc_15724_n5112) );
  AND2X2 AND2X2_2178 ( .A(_abc_15724_n5098), .B(_abc_15724_n5112), .Y(_abc_15724_n5113) );
  AND2X2 AND2X2_2179 ( .A(_abc_15724_n5114), .B(_abc_15724_n5115), .Y(_abc_15724_n5116) );
  AND2X2 AND2X2_218 ( .A(_abc_15724_n1140), .B(_abc_15724_n1144_1), .Y(_abc_15724_n1146) );
  AND2X2 AND2X2_2180 ( .A(_abc_15724_n5078), .B(_abc_15724_n5116), .Y(_abc_15724_n5117) );
  AND2X2 AND2X2_2181 ( .A(_abc_15724_n5118), .B(_abc_15724_n5119), .Y(_abc_15724_n5120) );
  AND2X2 AND2X2_2182 ( .A(_abc_15724_n5121), .B(_abc_15724_n4021), .Y(_abc_15724_n5122) );
  AND2X2 AND2X2_2183 ( .A(_abc_15724_n5120), .B(_abc_15724_n4022), .Y(_abc_15724_n5123) );
  AND2X2 AND2X2_2184 ( .A(_abc_15724_n5124), .B(_abc_15724_n5076), .Y(_abc_15724_n5126) );
  AND2X2 AND2X2_2185 ( .A(_abc_15724_n5127), .B(_abc_15724_n5125), .Y(_abc_15724_n5128) );
  AND2X2 AND2X2_2186 ( .A(_abc_15724_n5129), .B(_abc_15724_n5128), .Y(_abc_15724_n5130) );
  AND2X2 AND2X2_2187 ( .A(_abc_15724_n5132), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n5133) );
  AND2X2 AND2X2_2188 ( .A(_abc_15724_n5133), .B(_abc_15724_n5131), .Y(_abc_15724_n5134) );
  AND2X2 AND2X2_2189 ( .A(_abc_15724_n2992_bF_buf10), .B(a_reg_17_), .Y(_abc_15724_n5135) );
  AND2X2 AND2X2_219 ( .A(_abc_15724_n1147), .B(_abc_15724_n1145), .Y(_abc_15724_n1148) );
  AND2X2 AND2X2_2190 ( .A(_abc_15724_n906_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_145_), .Y(_abc_15724_n5136) );
  AND2X2 AND2X2_2191 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n5136), .Y(_abc_15724_n5137) );
  AND2X2 AND2X2_2192 ( .A(_abc_15724_n5131), .B(_abc_15724_n5125), .Y(_abc_15724_n5140) );
  AND2X2 AND2X2_2193 ( .A(_abc_15724_n5114), .B(_abc_15724_n5110), .Y(_abc_15724_n5143) );
  AND2X2 AND2X2_2194 ( .A(_abc_15724_n5146), .B(_abc_15724_n5147), .Y(_abc_15724_n5148) );
  AND2X2 AND2X2_2195 ( .A(c_reg_18_), .B(b_reg_18_), .Y(_abc_15724_n5149) );
  AND2X2 AND2X2_2196 ( .A(_abc_15724_n5150), .B(_abc_15724_n5145), .Y(_abc_15724_n5151) );
  AND2X2 AND2X2_2197 ( .A(_abc_15724_n5152), .B(_abc_15724_n5145), .Y(_abc_15724_n5153) );
  AND2X2 AND2X2_2198 ( .A(_abc_15724_n5155), .B(_abc_15724_n5152), .Y(_abc_15724_n5156) );
  AND2X2 AND2X2_2199 ( .A(_abc_15724_n5146), .B(b_reg_18_), .Y(_abc_15724_n5159) );
  AND2X2 AND2X2_22 ( .A(e_reg_12_), .B(_auto_iopadmap_cc_313_execute_26059_12_), .Y(_abc_15724_n741_1) );
  AND2X2 AND2X2_220 ( .A(_abc_15724_n1148), .B(digest_update_bF_buf2), .Y(_abc_15724_n1149) );
  AND2X2 AND2X2_2200 ( .A(_abc_15724_n3737_bF_buf4), .B(_abc_15724_n5155), .Y(_abc_15724_n5162) );
  AND2X2 AND2X2_2201 ( .A(_abc_15724_n5163), .B(_abc_15724_n5161), .Y(_abc_15724_n5164) );
  AND2X2 AND2X2_2202 ( .A(_abc_15724_n5158), .B(_abc_15724_n5164), .Y(_abc_15724_n5165) );
  AND2X2 AND2X2_2203 ( .A(_abc_15724_n5106), .B(_abc_15724_n5103), .Y(_abc_15724_n5166) );
  AND2X2 AND2X2_2204 ( .A(a_reg_13_), .B(e_reg_18_), .Y(_abc_15724_n5169) );
  AND2X2 AND2X2_2205 ( .A(_abc_15724_n5170), .B(_abc_15724_n5168), .Y(_abc_15724_n5171) );
  AND2X2 AND2X2_2206 ( .A(_abc_15724_n5171), .B(w_18_), .Y(_abc_15724_n5172) );
  AND2X2 AND2X2_2207 ( .A(_abc_15724_n5173), .B(_abc_15724_n5174), .Y(_abc_15724_n5175) );
  AND2X2 AND2X2_2208 ( .A(_abc_15724_n5167), .B(_abc_15724_n5175), .Y(_abc_15724_n5176) );
  AND2X2 AND2X2_2209 ( .A(_abc_15724_n5177), .B(_abc_15724_n5178), .Y(_abc_15724_n5179) );
  AND2X2 AND2X2_221 ( .A(_abc_15724_n1150), .B(_abc_15724_n850_bF_buf3), .Y(_abc_15724_n1151) );
  AND2X2 AND2X2_2210 ( .A(_abc_15724_n5180), .B(_abc_15724_n5165), .Y(_abc_15724_n5181) );
  AND2X2 AND2X2_2211 ( .A(_abc_15724_n5185), .B(_abc_15724_n5144), .Y(_abc_15724_n5186) );
  AND2X2 AND2X2_2212 ( .A(_abc_15724_n5184), .B(_abc_15724_n5143), .Y(_abc_15724_n5187) );
  AND2X2 AND2X2_2213 ( .A(_abc_15724_n5142), .B(_abc_15724_n5189), .Y(_abc_15724_n5190) );
  AND2X2 AND2X2_2214 ( .A(_abc_15724_n5191), .B(_abc_15724_n5188), .Y(_abc_15724_n5192) );
  AND2X2 AND2X2_2215 ( .A(_abc_15724_n5196), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n5197) );
  AND2X2 AND2X2_2216 ( .A(_abc_15724_n5197), .B(_abc_15724_n5195), .Y(_abc_15724_n5198) );
  AND2X2 AND2X2_2217 ( .A(_abc_15724_n2992_bF_buf9), .B(a_reg_18_), .Y(_abc_15724_n5199) );
  AND2X2 AND2X2_2218 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n2768_1), .Y(_abc_15724_n5200) );
  AND2X2 AND2X2_2219 ( .A(_abc_15724_n5196), .B(_abc_15724_n5203), .Y(_abc_15724_n5204) );
  AND2X2 AND2X2_222 ( .A(_abc_15724_n1147), .B(_abc_15724_n1143), .Y(_abc_15724_n1153) );
  AND2X2 AND2X2_2220 ( .A(_abc_15724_n5182), .B(_abc_15724_n5177), .Y(_abc_15724_n5206) );
  AND2X2 AND2X2_2221 ( .A(_abc_15724_n5209), .B(_abc_15724_n5210), .Y(_abc_15724_n5211) );
  AND2X2 AND2X2_2222 ( .A(c_reg_19_), .B(b_reg_19_), .Y(_abc_15724_n5212) );
  AND2X2 AND2X2_2223 ( .A(_abc_15724_n5213), .B(_abc_15724_n5208), .Y(_abc_15724_n5214) );
  AND2X2 AND2X2_2224 ( .A(_abc_15724_n5215), .B(_abc_15724_n5216), .Y(_abc_15724_n5217) );
  AND2X2 AND2X2_2225 ( .A(_abc_15724_n3726_bF_buf3), .B(_abc_15724_n5217), .Y(_abc_15724_n5218) );
  AND2X2 AND2X2_2226 ( .A(_abc_15724_n5220), .B(_abc_15724_n5208), .Y(_abc_15724_n5221) );
  AND2X2 AND2X2_2227 ( .A(_abc_15724_n5209), .B(b_reg_19_), .Y(_abc_15724_n5222) );
  AND2X2 AND2X2_2228 ( .A(_abc_15724_n5226), .B(_abc_15724_n5224), .Y(_abc_15724_n5227) );
  AND2X2 AND2X2_2229 ( .A(_abc_15724_n5219), .B(_abc_15724_n5227), .Y(_abc_15724_n5228) );
  AND2X2 AND2X2_223 ( .A(_auto_iopadmap_cc_313_execute_26059_43_), .B(d_reg_11_), .Y(_abc_15724_n1155_1) );
  AND2X2 AND2X2_2230 ( .A(_abc_15724_n5173), .B(_abc_15724_n5170), .Y(_abc_15724_n5229) );
  AND2X2 AND2X2_2231 ( .A(a_reg_14_), .B(e_reg_19_), .Y(_abc_15724_n5232) );
  AND2X2 AND2X2_2232 ( .A(_abc_15724_n5233), .B(_abc_15724_n5231), .Y(_abc_15724_n5234) );
  AND2X2 AND2X2_2233 ( .A(_abc_15724_n5234), .B(w_19_), .Y(_abc_15724_n5235) );
  AND2X2 AND2X2_2234 ( .A(_abc_15724_n5236), .B(_abc_15724_n5237), .Y(_abc_15724_n5238) );
  AND2X2 AND2X2_2235 ( .A(_abc_15724_n5230), .B(_abc_15724_n5238), .Y(_abc_15724_n5239) );
  AND2X2 AND2X2_2236 ( .A(_abc_15724_n5240), .B(_abc_15724_n5241), .Y(_abc_15724_n5242) );
  AND2X2 AND2X2_2237 ( .A(_abc_15724_n5243), .B(_abc_15724_n5228), .Y(_abc_15724_n5244) );
  AND2X2 AND2X2_2238 ( .A(_abc_15724_n5245), .B(_abc_15724_n5246), .Y(_abc_15724_n5247) );
  AND2X2 AND2X2_2239 ( .A(_abc_15724_n5207), .B(_abc_15724_n5247), .Y(_abc_15724_n5248) );
  AND2X2 AND2X2_224 ( .A(_abc_15724_n1156_1), .B(_abc_15724_n1154), .Y(_abc_15724_n1157_1) );
  AND2X2 AND2X2_2240 ( .A(_abc_15724_n5249), .B(_abc_15724_n5250), .Y(_abc_15724_n5251) );
  AND2X2 AND2X2_2241 ( .A(_abc_15724_n5251), .B(_abc_15724_n5056), .Y(_abc_15724_n5252) );
  AND2X2 AND2X2_2242 ( .A(_abc_15724_n5253), .B(_abc_15724_n5254), .Y(_abc_15724_n5255) );
  AND2X2 AND2X2_2243 ( .A(_abc_15724_n5255), .B(_abc_15724_n5186), .Y(_abc_15724_n5256) );
  AND2X2 AND2X2_2244 ( .A(_abc_15724_n5258), .B(_abc_15724_n5257), .Y(_abc_15724_n5259) );
  AND2X2 AND2X2_2245 ( .A(_abc_15724_n5263), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n5264) );
  AND2X2 AND2X2_2246 ( .A(_abc_15724_n5264), .B(_abc_15724_n5262), .Y(_abc_15724_n5265) );
  AND2X2 AND2X2_2247 ( .A(_abc_15724_n2992_bF_buf8), .B(a_reg_19_), .Y(_abc_15724_n5266) );
  AND2X2 AND2X2_2248 ( .A(_abc_15724_n906_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_147_), .Y(_abc_15724_n5267) );
  AND2X2 AND2X2_2249 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n5267), .Y(_abc_15724_n5268) );
  AND2X2 AND2X2_225 ( .A(_abc_15724_n1153), .B(_abc_15724_n1157_1), .Y(_abc_15724_n1158) );
  AND2X2 AND2X2_2250 ( .A(_abc_15724_n5271), .B(_abc_15724_n5272), .Y(_abc_15724_n5273) );
  AND2X2 AND2X2_2251 ( .A(_abc_15724_n5060), .B(_abc_15724_n5125), .Y(_abc_15724_n5275) );
  AND2X2 AND2X2_2252 ( .A(_abc_15724_n5278), .B(_abc_15724_n5274), .Y(_abc_15724_n5279) );
  AND2X2 AND2X2_2253 ( .A(_abc_15724_n5283), .B(_abc_15724_n5279), .Y(_abc_15724_n5284) );
  AND2X2 AND2X2_2254 ( .A(_abc_15724_n5253), .B(_abc_15724_n5249), .Y(_abc_15724_n5286) );
  AND2X2 AND2X2_2255 ( .A(_abc_15724_n5246), .B(_abc_15724_n5240), .Y(_abc_15724_n5288) );
  AND2X2 AND2X2_2256 ( .A(_abc_15724_n5291), .B(_abc_15724_n5292), .Y(_abc_15724_n5293) );
  AND2X2 AND2X2_2257 ( .A(c_reg_20_), .B(b_reg_20_), .Y(_abc_15724_n5294) );
  AND2X2 AND2X2_2258 ( .A(_abc_15724_n5295), .B(_abc_15724_n5290), .Y(_abc_15724_n5296) );
  AND2X2 AND2X2_2259 ( .A(_abc_15724_n5297), .B(_abc_15724_n5290), .Y(_abc_15724_n5298) );
  AND2X2 AND2X2_226 ( .A(_abc_15724_n1159), .B(_abc_15724_n1160), .Y(_abc_15724_n1161) );
  AND2X2 AND2X2_2260 ( .A(_abc_15724_n5300), .B(_abc_15724_n5297), .Y(_abc_15724_n5301) );
  AND2X2 AND2X2_2261 ( .A(_abc_15724_n5291), .B(b_reg_20_), .Y(_abc_15724_n5304) );
  AND2X2 AND2X2_2262 ( .A(_abc_15724_n3737_bF_buf3), .B(_abc_15724_n5300), .Y(_abc_15724_n5307) );
  AND2X2 AND2X2_2263 ( .A(_abc_15724_n5308), .B(_abc_15724_n5306), .Y(_abc_15724_n5309) );
  AND2X2 AND2X2_2264 ( .A(_abc_15724_n5303), .B(_abc_15724_n5309), .Y(_abc_15724_n5310) );
  AND2X2 AND2X2_2265 ( .A(_abc_15724_n5236), .B(_abc_15724_n5233), .Y(_abc_15724_n5311) );
  AND2X2 AND2X2_2266 ( .A(a_reg_15_), .B(e_reg_20_), .Y(_abc_15724_n5314) );
  AND2X2 AND2X2_2267 ( .A(_abc_15724_n5315), .B(_abc_15724_n5313), .Y(_abc_15724_n5316) );
  AND2X2 AND2X2_2268 ( .A(_abc_15724_n5316), .B(w_20_), .Y(_abc_15724_n5317) );
  AND2X2 AND2X2_2269 ( .A(_abc_15724_n5318), .B(_abc_15724_n5319), .Y(_abc_15724_n5320) );
  AND2X2 AND2X2_227 ( .A(_abc_15724_n1162), .B(digest_update_bF_buf1), .Y(_abc_15724_n1163) );
  AND2X2 AND2X2_2270 ( .A(_abc_15724_n5312), .B(_abc_15724_n5320), .Y(_abc_15724_n5321) );
  AND2X2 AND2X2_2271 ( .A(_abc_15724_n5322), .B(_abc_15724_n5323), .Y(_abc_15724_n5324) );
  AND2X2 AND2X2_2272 ( .A(_abc_15724_n5325), .B(_abc_15724_n5310), .Y(_abc_15724_n5326) );
  AND2X2 AND2X2_2273 ( .A(_abc_15724_n5330), .B(_abc_15724_n5289), .Y(_abc_15724_n5331) );
  AND2X2 AND2X2_2274 ( .A(_abc_15724_n5329), .B(_abc_15724_n5288), .Y(_abc_15724_n5332) );
  AND2X2 AND2X2_2275 ( .A(_abc_15724_n5333), .B(_abc_15724_n5006), .Y(_abc_15724_n5334) );
  AND2X2 AND2X2_2276 ( .A(_abc_15724_n5338), .B(_abc_15724_n5287), .Y(_abc_15724_n5339) );
  AND2X2 AND2X2_2277 ( .A(_abc_15724_n5337), .B(_abc_15724_n5286), .Y(_abc_15724_n5340) );
  AND2X2 AND2X2_2278 ( .A(_abc_15724_n5344), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n5345) );
  AND2X2 AND2X2_2279 ( .A(_abc_15724_n5345), .B(_abc_15724_n5343), .Y(_abc_15724_n5346) );
  AND2X2 AND2X2_228 ( .A(_abc_15724_n907_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_43_), .Y(_abc_15724_n1164) );
  AND2X2 AND2X2_2280 ( .A(_abc_15724_n2992_bF_buf7), .B(a_reg_20_), .Y(_abc_15724_n5347) );
  AND2X2 AND2X2_2281 ( .A(_abc_15724_n906_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_148_), .Y(_abc_15724_n5348) );
  AND2X2 AND2X2_2282 ( .A(_abc_15724_n2994_bF_buf7), .B(_abc_15724_n5348), .Y(_abc_15724_n5349) );
  AND2X2 AND2X2_2283 ( .A(_abc_15724_n5335), .B(_abc_15724_n5353), .Y(_abc_15724_n5354) );
  AND2X2 AND2X2_2284 ( .A(_abc_15724_n5327), .B(_abc_15724_n5322), .Y(_abc_15724_n5356) );
  AND2X2 AND2X2_2285 ( .A(_abc_15724_n5359), .B(_abc_15724_n5360), .Y(_abc_15724_n5361) );
  AND2X2 AND2X2_2286 ( .A(c_reg_21_), .B(b_reg_21_), .Y(_abc_15724_n5362) );
  AND2X2 AND2X2_2287 ( .A(_abc_15724_n5363), .B(_abc_15724_n5358), .Y(_abc_15724_n5364) );
  AND2X2 AND2X2_2288 ( .A(_abc_15724_n5365), .B(_abc_15724_n5358), .Y(_abc_15724_n5366) );
  AND2X2 AND2X2_2289 ( .A(_abc_15724_n5368), .B(_abc_15724_n5365), .Y(_abc_15724_n5369) );
  AND2X2 AND2X2_229 ( .A(_abc_15724_n1126), .B(_abc_15724_n1117), .Y(_abc_15724_n1166_1) );
  AND2X2 AND2X2_2290 ( .A(_abc_15724_n5359), .B(b_reg_21_), .Y(_abc_15724_n5372) );
  AND2X2 AND2X2_2291 ( .A(_abc_15724_n3737_bF_buf2), .B(_abc_15724_n5368), .Y(_abc_15724_n5375) );
  AND2X2 AND2X2_2292 ( .A(_abc_15724_n5376), .B(_abc_15724_n5374), .Y(_abc_15724_n5377) );
  AND2X2 AND2X2_2293 ( .A(_abc_15724_n5371), .B(_abc_15724_n5377), .Y(_abc_15724_n5378) );
  AND2X2 AND2X2_2294 ( .A(_abc_15724_n5318), .B(_abc_15724_n5315), .Y(_abc_15724_n5379) );
  AND2X2 AND2X2_2295 ( .A(e_reg_21_), .B(a_reg_16_), .Y(_abc_15724_n5382) );
  AND2X2 AND2X2_2296 ( .A(_abc_15724_n5383), .B(_abc_15724_n5381), .Y(_abc_15724_n5384) );
  AND2X2 AND2X2_2297 ( .A(_abc_15724_n5384), .B(w_21_), .Y(_abc_15724_n5385) );
  AND2X2 AND2X2_2298 ( .A(_abc_15724_n5386), .B(_abc_15724_n5387), .Y(_abc_15724_n5388) );
  AND2X2 AND2X2_2299 ( .A(_abc_15724_n5380), .B(_abc_15724_n5388), .Y(_abc_15724_n5389) );
  AND2X2 AND2X2_23 ( .A(_abc_15724_n740), .B(_abc_15724_n742), .Y(_abc_15724_n743) );
  AND2X2 AND2X2_230 ( .A(_abc_15724_n1144_1), .B(_abc_15724_n1157_1), .Y(_abc_15724_n1168) );
  AND2X2 AND2X2_2300 ( .A(_abc_15724_n5390), .B(_abc_15724_n5391), .Y(_abc_15724_n5392) );
  AND2X2 AND2X2_2301 ( .A(_abc_15724_n5393), .B(_abc_15724_n5378), .Y(_abc_15724_n5394) );
  AND2X2 AND2X2_2302 ( .A(_abc_15724_n5395), .B(_abc_15724_n5396), .Y(_abc_15724_n5397) );
  AND2X2 AND2X2_2303 ( .A(_abc_15724_n5357), .B(_abc_15724_n5397), .Y(_abc_15724_n5398) );
  AND2X2 AND2X2_2304 ( .A(_abc_15724_n5399), .B(_abc_15724_n5400), .Y(_abc_15724_n5401) );
  AND2X2 AND2X2_2305 ( .A(_abc_15724_n5402), .B(_abc_15724_n3736), .Y(_abc_15724_n5403) );
  AND2X2 AND2X2_2306 ( .A(_abc_15724_n5401), .B(_abc_15724_n3724), .Y(_abc_15724_n5404) );
  AND2X2 AND2X2_2307 ( .A(_abc_15724_n5406), .B(_abc_15724_n5355), .Y(_abc_15724_n5407) );
  AND2X2 AND2X2_2308 ( .A(_abc_15724_n5405), .B(_abc_15724_n5354), .Y(_abc_15724_n5408) );
  AND2X2 AND2X2_2309 ( .A(_abc_15724_n5414), .B(_abc_15724_n5416), .Y(_abc_15724_n5417) );
  AND2X2 AND2X2_231 ( .A(_abc_15724_n1168), .B(_abc_15724_n1167_1), .Y(_abc_15724_n1169) );
  AND2X2 AND2X2_2310 ( .A(_abc_15724_n5417), .B(round_ctr_inc_bF_buf5), .Y(_abc_15724_n5418) );
  AND2X2 AND2X2_2311 ( .A(_abc_15724_n5418), .B(_abc_15724_n5412), .Y(_abc_15724_n5419) );
  AND2X2 AND2X2_2312 ( .A(_abc_15724_n2992_bF_buf6), .B(a_reg_21_), .Y(_abc_15724_n5420) );
  AND2X2 AND2X2_2313 ( .A(_abc_15724_n906_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_149_), .Y(_abc_15724_n5421) );
  AND2X2 AND2X2_2314 ( .A(_abc_15724_n2994_bF_buf6), .B(_abc_15724_n5421), .Y(_abc_15724_n5422) );
  AND2X2 AND2X2_2315 ( .A(_abc_15724_n5416), .B(_abc_15724_n5425), .Y(_abc_15724_n5426) );
  AND2X2 AND2X2_2316 ( .A(_abc_15724_n5414), .B(_abc_15724_n5426), .Y(_abc_15724_n5427) );
  AND2X2 AND2X2_2317 ( .A(_abc_15724_n5429), .B(_abc_15724_n5399), .Y(_abc_15724_n5430) );
  AND2X2 AND2X2_2318 ( .A(_abc_15724_n5396), .B(_abc_15724_n5390), .Y(_abc_15724_n5432) );
  AND2X2 AND2X2_2319 ( .A(_abc_15724_n5435), .B(_abc_15724_n5436), .Y(_abc_15724_n5437) );
  AND2X2 AND2X2_232 ( .A(_abc_15724_n1154), .B(_abc_15724_n1142_1), .Y(_abc_15724_n1170) );
  AND2X2 AND2X2_2320 ( .A(c_reg_22_), .B(b_reg_22_), .Y(_abc_15724_n5438) );
  AND2X2 AND2X2_2321 ( .A(_abc_15724_n5439), .B(_abc_15724_n5434), .Y(_abc_15724_n5440) );
  AND2X2 AND2X2_2322 ( .A(_abc_15724_n5441), .B(_abc_15724_n5434), .Y(_abc_15724_n5442) );
  AND2X2 AND2X2_2323 ( .A(_abc_15724_n5444), .B(_abc_15724_n5441), .Y(_abc_15724_n5445) );
  AND2X2 AND2X2_2324 ( .A(_abc_15724_n5435), .B(b_reg_22_), .Y(_abc_15724_n5448) );
  AND2X2 AND2X2_2325 ( .A(_abc_15724_n3737_bF_buf1), .B(_abc_15724_n5444), .Y(_abc_15724_n5451) );
  AND2X2 AND2X2_2326 ( .A(_abc_15724_n5452), .B(_abc_15724_n5450), .Y(_abc_15724_n5453) );
  AND2X2 AND2X2_2327 ( .A(_abc_15724_n5447), .B(_abc_15724_n5453), .Y(_abc_15724_n5454) );
  AND2X2 AND2X2_2328 ( .A(_abc_15724_n5386), .B(_abc_15724_n5383), .Y(_abc_15724_n5455) );
  AND2X2 AND2X2_2329 ( .A(e_reg_22_), .B(a_reg_17_), .Y(_abc_15724_n5458) );
  AND2X2 AND2X2_233 ( .A(_abc_15724_n1119_1), .B(_abc_15724_n1129), .Y(_abc_15724_n1173) );
  AND2X2 AND2X2_2330 ( .A(_abc_15724_n5459), .B(_abc_15724_n5457), .Y(_abc_15724_n5460) );
  AND2X2 AND2X2_2331 ( .A(_abc_15724_n5460), .B(w_22_), .Y(_abc_15724_n5461) );
  AND2X2 AND2X2_2332 ( .A(_abc_15724_n5462), .B(_abc_15724_n5463), .Y(_abc_15724_n5464) );
  AND2X2 AND2X2_2333 ( .A(_abc_15724_n5456), .B(_abc_15724_n5464), .Y(_abc_15724_n5465) );
  AND2X2 AND2X2_2334 ( .A(_abc_15724_n5466), .B(_abc_15724_n5467), .Y(_abc_15724_n5468) );
  AND2X2 AND2X2_2335 ( .A(_abc_15724_n5469), .B(_abc_15724_n5454), .Y(_abc_15724_n5470) );
  AND2X2 AND2X2_2336 ( .A(_abc_15724_n5471), .B(_abc_15724_n5472), .Y(_abc_15724_n5473) );
  AND2X2 AND2X2_2337 ( .A(_abc_15724_n5433), .B(_abc_15724_n5473), .Y(_abc_15724_n5474) );
  AND2X2 AND2X2_2338 ( .A(_abc_15724_n5475), .B(_abc_15724_n5476), .Y(_abc_15724_n5477) );
  AND2X2 AND2X2_2339 ( .A(_abc_15724_n5478), .B(_abc_15724_n3806_bF_buf3), .Y(_abc_15724_n5479) );
  AND2X2 AND2X2_234 ( .A(_abc_15724_n1173), .B(_abc_15724_n1168), .Y(_abc_15724_n1174) );
  AND2X2 AND2X2_2340 ( .A(_abc_15724_n5477), .B(_abc_15724_n3726_bF_buf2), .Y(_abc_15724_n5480) );
  AND2X2 AND2X2_2341 ( .A(_abc_15724_n5482), .B(_abc_15724_n5431), .Y(_abc_15724_n5483) );
  AND2X2 AND2X2_2342 ( .A(_abc_15724_n5481), .B(_abc_15724_n5430), .Y(_abc_15724_n5484) );
  AND2X2 AND2X2_2343 ( .A(_abc_15724_n5488), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n5489) );
  AND2X2 AND2X2_2344 ( .A(_abc_15724_n5489), .B(_abc_15724_n5487), .Y(_abc_15724_n5490) );
  AND2X2 AND2X2_2345 ( .A(_abc_15724_n2992_bF_buf5), .B(a_reg_22_), .Y(_abc_15724_n5491) );
  AND2X2 AND2X2_2346 ( .A(_abc_15724_n2994_bF_buf5), .B(_abc_15724_n2832), .Y(_abc_15724_n5492) );
  AND2X2 AND2X2_2347 ( .A(_abc_15724_n5488), .B(_abc_15724_n5495), .Y(_abc_15724_n5496) );
  AND2X2 AND2X2_2348 ( .A(_abc_15724_n5472), .B(_abc_15724_n5466), .Y(_abc_15724_n5499) );
  AND2X2 AND2X2_2349 ( .A(c_reg_23_), .B(b_reg_23_), .Y(_abc_15724_n5501) );
  AND2X2 AND2X2_235 ( .A(_abc_15724_n1115), .B(_abc_15724_n1174), .Y(_abc_15724_n1175) );
  AND2X2 AND2X2_2350 ( .A(_abc_15724_n5504), .B(_abc_15724_n5502), .Y(_abc_15724_n5505) );
  AND2X2 AND2X2_2351 ( .A(_abc_15724_n3805_bF_buf3), .B(_abc_15724_n5505), .Y(_abc_15724_n5506) );
  AND2X2 AND2X2_2352 ( .A(_abc_15724_n5502), .B(_abc_15724_n5508), .Y(_abc_15724_n5509) );
  AND2X2 AND2X2_2353 ( .A(_abc_15724_n5509), .B(d_reg_23_), .Y(_abc_15724_n5511) );
  AND2X2 AND2X2_2354 ( .A(_abc_15724_n5512), .B(_abc_15724_n5510), .Y(_abc_15724_n5513) );
  AND2X2 AND2X2_2355 ( .A(_abc_15724_n3726_bF_buf1), .B(_abc_15724_n5513), .Y(_abc_15724_n5514) );
  AND2X2 AND2X2_2356 ( .A(_abc_15724_n5515), .B(_abc_15724_n5508), .Y(_abc_15724_n5516) );
  AND2X2 AND2X2_2357 ( .A(_abc_15724_n3737_bF_buf0), .B(_abc_15724_n5516), .Y(_abc_15724_n5517) );
  AND2X2 AND2X2_2358 ( .A(_abc_15724_n5519), .B(_abc_15724_n5507), .Y(_abc_15724_n5520) );
  AND2X2 AND2X2_2359 ( .A(_abc_15724_n5462), .B(_abc_15724_n5459), .Y(_abc_15724_n5521) );
  AND2X2 AND2X2_236 ( .A(_auto_iopadmap_cc_313_execute_26059_44_), .B(d_reg_12_), .Y(_abc_15724_n1178_1) );
  AND2X2 AND2X2_2360 ( .A(e_reg_23_), .B(a_reg_18_), .Y(_abc_15724_n5524) );
  AND2X2 AND2X2_2361 ( .A(_abc_15724_n5525), .B(_abc_15724_n5523), .Y(_abc_15724_n5526) );
  AND2X2 AND2X2_2362 ( .A(_abc_15724_n5526), .B(w_23_), .Y(_abc_15724_n5527) );
  AND2X2 AND2X2_2363 ( .A(_abc_15724_n5528), .B(_abc_15724_n5529), .Y(_abc_15724_n5530) );
  AND2X2 AND2X2_2364 ( .A(_abc_15724_n5522), .B(_abc_15724_n5530), .Y(_abc_15724_n5531) );
  AND2X2 AND2X2_2365 ( .A(_abc_15724_n5532), .B(_abc_15724_n5533), .Y(_abc_15724_n5534) );
  AND2X2 AND2X2_2366 ( .A(_abc_15724_n5520), .B(_abc_15724_n5534), .Y(_abc_15724_n5535) );
  AND2X2 AND2X2_2367 ( .A(_abc_15724_n5536), .B(_abc_15724_n5537), .Y(_abc_15724_n5538) );
  AND2X2 AND2X2_2368 ( .A(_abc_15724_n5500), .B(_abc_15724_n5538), .Y(_abc_15724_n5539) );
  AND2X2 AND2X2_2369 ( .A(_abc_15724_n5540), .B(_abc_15724_n5541), .Y(_abc_15724_n5542) );
  AND2X2 AND2X2_237 ( .A(_abc_15724_n1179_1), .B(_abc_15724_n1177_1), .Y(_abc_15724_n1180) );
  AND2X2 AND2X2_2370 ( .A(_abc_15724_n5542), .B(_abc_15724_n3706), .Y(_abc_15724_n5543) );
  AND2X2 AND2X2_2371 ( .A(_abc_15724_n5544), .B(_abc_15724_n5545), .Y(_abc_15724_n5546) );
  AND2X2 AND2X2_2372 ( .A(_abc_15724_n5546), .B(_abc_15724_n5498), .Y(_abc_15724_n5547) );
  AND2X2 AND2X2_2373 ( .A(_abc_15724_n5549), .B(_abc_15724_n5548), .Y(_abc_15724_n5550) );
  AND2X2 AND2X2_2374 ( .A(_abc_15724_n5554), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n5555) );
  AND2X2 AND2X2_2375 ( .A(_abc_15724_n5555), .B(_abc_15724_n5553), .Y(_abc_15724_n5556) );
  AND2X2 AND2X2_2376 ( .A(_abc_15724_n2992_bF_buf4), .B(a_reg_23_), .Y(_abc_15724_n5557) );
  AND2X2 AND2X2_2377 ( .A(_abc_15724_n906_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_151_), .Y(_abc_15724_n5558) );
  AND2X2 AND2X2_2378 ( .A(_abc_15724_n2994_bF_buf4), .B(_abc_15724_n5558), .Y(_abc_15724_n5559) );
  AND2X2 AND2X2_2379 ( .A(_abc_15724_n5567), .B(_abc_15724_n5566), .Y(_abc_15724_n5568) );
  AND2X2 AND2X2_238 ( .A(_abc_15724_n1176), .B(_abc_15724_n1180), .Y(_abc_15724_n1182) );
  AND2X2 AND2X2_2380 ( .A(_abc_15724_n5565), .B(_abc_15724_n5568), .Y(_abc_15724_n5569) );
  AND2X2 AND2X2_2381 ( .A(_abc_15724_n5569), .B(_abc_15724_n5564), .Y(_abc_15724_n5570) );
  AND2X2 AND2X2_2382 ( .A(_abc_15724_n5572), .B(_abc_15724_n5570), .Y(_abc_15724_n5573) );
  AND2X2 AND2X2_2383 ( .A(_abc_15724_n5544), .B(_abc_15724_n5540), .Y(_abc_15724_n5575) );
  AND2X2 AND2X2_2384 ( .A(_abc_15724_n5536), .B(_abc_15724_n5532), .Y(_abc_15724_n5577) );
  AND2X2 AND2X2_2385 ( .A(c_reg_24_), .B(b_reg_24_), .Y(_abc_15724_n5579) );
  AND2X2 AND2X2_2386 ( .A(_abc_15724_n5582), .B(_abc_15724_n5580), .Y(_abc_15724_n5583) );
  AND2X2 AND2X2_2387 ( .A(_abc_15724_n3805_bF_buf1), .B(_abc_15724_n5583), .Y(_abc_15724_n5584) );
  AND2X2 AND2X2_2388 ( .A(_abc_15724_n5580), .B(_abc_15724_n5586), .Y(_abc_15724_n5587) );
  AND2X2 AND2X2_2389 ( .A(_abc_15724_n5587), .B(d_reg_24_), .Y(_abc_15724_n5589) );
  AND2X2 AND2X2_239 ( .A(_abc_15724_n1183), .B(_abc_15724_n1181), .Y(_abc_15724_n1184) );
  AND2X2 AND2X2_2390 ( .A(_abc_15724_n5590), .B(_abc_15724_n5588), .Y(_abc_15724_n5591) );
  AND2X2 AND2X2_2391 ( .A(_abc_15724_n3726_bF_buf0), .B(_abc_15724_n5591), .Y(_abc_15724_n5592) );
  AND2X2 AND2X2_2392 ( .A(_abc_15724_n5580), .B(_abc_15724_n5581), .Y(_abc_15724_n5593) );
  AND2X2 AND2X2_2393 ( .A(_abc_15724_n3737_bF_buf4), .B(_abc_15724_n5596), .Y(_abc_15724_n5597) );
  AND2X2 AND2X2_2394 ( .A(_abc_15724_n5599), .B(_abc_15724_n5585), .Y(_abc_15724_n5600) );
  AND2X2 AND2X2_2395 ( .A(_abc_15724_n5528), .B(_abc_15724_n5525), .Y(_abc_15724_n5601) );
  AND2X2 AND2X2_2396 ( .A(e_reg_24_), .B(a_reg_19_), .Y(_abc_15724_n5604) );
  AND2X2 AND2X2_2397 ( .A(_abc_15724_n5605), .B(_abc_15724_n5603), .Y(_abc_15724_n5606) );
  AND2X2 AND2X2_2398 ( .A(_abc_15724_n5606), .B(w_24_), .Y(_abc_15724_n5607) );
  AND2X2 AND2X2_2399 ( .A(_abc_15724_n5608), .B(_abc_15724_n5609), .Y(_abc_15724_n5610) );
  AND2X2 AND2X2_24 ( .A(_abc_15724_n744), .B(_abc_15724_n738_1), .Y(_abc_15724_n745) );
  AND2X2 AND2X2_240 ( .A(_abc_15724_n1184), .B(digest_update_bF_buf0), .Y(_abc_15724_n1185_1) );
  AND2X2 AND2X2_2400 ( .A(_abc_15724_n5602), .B(_abc_15724_n5610), .Y(_abc_15724_n5611) );
  AND2X2 AND2X2_2401 ( .A(_abc_15724_n5612), .B(_abc_15724_n5613), .Y(_abc_15724_n5614) );
  AND2X2 AND2X2_2402 ( .A(_abc_15724_n5600), .B(_abc_15724_n5614), .Y(_abc_15724_n5615) );
  AND2X2 AND2X2_2403 ( .A(_abc_15724_n5616), .B(_abc_15724_n5617), .Y(_abc_15724_n5618) );
  AND2X2 AND2X2_2404 ( .A(_abc_15724_n5578), .B(_abc_15724_n5618), .Y(_abc_15724_n5619) );
  AND2X2 AND2X2_2405 ( .A(_abc_15724_n5620), .B(_abc_15724_n5621), .Y(_abc_15724_n5622) );
  AND2X2 AND2X2_2406 ( .A(_abc_15724_n5623), .B(_abc_15724_n3725_bF_buf2), .Y(_abc_15724_n5624) );
  AND2X2 AND2X2_2407 ( .A(_abc_15724_n5622), .B(_abc_15724_n3737_bF_buf3), .Y(_abc_15724_n5625) );
  AND2X2 AND2X2_2408 ( .A(_abc_15724_n5627), .B(_abc_15724_n5576), .Y(_abc_15724_n5628) );
  AND2X2 AND2X2_2409 ( .A(_abc_15724_n5626), .B(_abc_15724_n5575), .Y(_abc_15724_n5629) );
  AND2X2 AND2X2_241 ( .A(_abc_15724_n1186_1), .B(_abc_15724_n850_bF_buf2), .Y(_abc_15724_n1187_1) );
  AND2X2 AND2X2_2410 ( .A(_abc_15724_n5574), .B(_abc_15724_n5631), .Y(_abc_15724_n5632) );
  AND2X2 AND2X2_2411 ( .A(_abc_15724_n5634), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n5635) );
  AND2X2 AND2X2_2412 ( .A(_abc_15724_n5635), .B(_abc_15724_n5633), .Y(_abc_15724_n5636) );
  AND2X2 AND2X2_2413 ( .A(_abc_15724_n2992_bF_buf3), .B(a_reg_24_), .Y(_abc_15724_n5637) );
  AND2X2 AND2X2_2414 ( .A(_abc_15724_n2994_bF_buf3), .B(_abc_15724_n2871), .Y(_abc_15724_n5638) );
  AND2X2 AND2X2_2415 ( .A(_abc_15724_n5616), .B(_abc_15724_n5612), .Y(_abc_15724_n5642) );
  AND2X2 AND2X2_2416 ( .A(c_reg_25_), .B(b_reg_25_), .Y(_abc_15724_n5644) );
  AND2X2 AND2X2_2417 ( .A(_abc_15724_n5647), .B(_abc_15724_n5645), .Y(_abc_15724_n5648) );
  AND2X2 AND2X2_2418 ( .A(_abc_15724_n3805_bF_buf4), .B(_abc_15724_n5648), .Y(_abc_15724_n5649) );
  AND2X2 AND2X2_2419 ( .A(_abc_15724_n5645), .B(_abc_15724_n5651), .Y(_abc_15724_n5652) );
  AND2X2 AND2X2_242 ( .A(_abc_15724_n907_1_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_45_), .Y(_abc_15724_n1189) );
  AND2X2 AND2X2_2420 ( .A(_abc_15724_n5652), .B(d_reg_25_), .Y(_abc_15724_n5654) );
  AND2X2 AND2X2_2421 ( .A(_abc_15724_n5655), .B(_abc_15724_n5653), .Y(_abc_15724_n5656) );
  AND2X2 AND2X2_2422 ( .A(_abc_15724_n3726_bF_buf4), .B(_abc_15724_n5656), .Y(_abc_15724_n5657) );
  AND2X2 AND2X2_2423 ( .A(_abc_15724_n5645), .B(_abc_15724_n5646), .Y(_abc_15724_n5658) );
  AND2X2 AND2X2_2424 ( .A(_abc_15724_n3737_bF_buf2), .B(_abc_15724_n5661), .Y(_abc_15724_n5662) );
  AND2X2 AND2X2_2425 ( .A(_abc_15724_n5664), .B(_abc_15724_n5650), .Y(_abc_15724_n5665) );
  AND2X2 AND2X2_2426 ( .A(_abc_15724_n5608), .B(_abc_15724_n5605), .Y(_abc_15724_n5666) );
  AND2X2 AND2X2_2427 ( .A(e_reg_25_), .B(a_reg_20_), .Y(_abc_15724_n5669) );
  AND2X2 AND2X2_2428 ( .A(_abc_15724_n5670), .B(_abc_15724_n5668), .Y(_abc_15724_n5671) );
  AND2X2 AND2X2_2429 ( .A(_abc_15724_n5671), .B(w_25_), .Y(_abc_15724_n5672) );
  AND2X2 AND2X2_243 ( .A(_auto_iopadmap_cc_313_execute_26059_45_), .B(d_reg_13_), .Y(_abc_15724_n1191_1) );
  AND2X2 AND2X2_2430 ( .A(_abc_15724_n5673), .B(_abc_15724_n5674), .Y(_abc_15724_n5675) );
  AND2X2 AND2X2_2431 ( .A(_abc_15724_n5667), .B(_abc_15724_n5675), .Y(_abc_15724_n5676) );
  AND2X2 AND2X2_2432 ( .A(_abc_15724_n5677), .B(_abc_15724_n5678), .Y(_abc_15724_n5679) );
  AND2X2 AND2X2_2433 ( .A(_abc_15724_n5665), .B(_abc_15724_n5679), .Y(_abc_15724_n5680) );
  AND2X2 AND2X2_2434 ( .A(_abc_15724_n5681), .B(_abc_15724_n5682), .Y(_abc_15724_n5683) );
  AND2X2 AND2X2_2435 ( .A(_abc_15724_n5643), .B(_abc_15724_n5683), .Y(_abc_15724_n5684) );
  AND2X2 AND2X2_2436 ( .A(_abc_15724_n5641), .B(_abc_15724_n5687), .Y(_abc_15724_n5688) );
  AND2X2 AND2X2_2437 ( .A(_abc_15724_n5689), .B(_abc_15724_n5690), .Y(_abc_15724_n5691) );
  AND2X2 AND2X2_2438 ( .A(_abc_15724_n5631), .B(_abc_15724_n5691), .Y(_abc_15724_n5694) );
  AND2X2 AND2X2_2439 ( .A(_abc_15724_n5691), .B(_abc_15724_n5628), .Y(_abc_15724_n5697) );
  AND2X2 AND2X2_244 ( .A(_abc_15724_n1192), .B(_abc_15724_n1190_1), .Y(_abc_15724_n1193_1) );
  AND2X2 AND2X2_2440 ( .A(_abc_15724_n5698), .B(round_ctr_inc_bF_buf1), .Y(_abc_15724_n5699) );
  AND2X2 AND2X2_2441 ( .A(_abc_15724_n5696), .B(_abc_15724_n5699), .Y(_abc_15724_n5700) );
  AND2X2 AND2X2_2442 ( .A(_abc_15724_n5693), .B(_abc_15724_n5700), .Y(_abc_15724_n5701) );
  AND2X2 AND2X2_2443 ( .A(_abc_15724_n2992_bF_buf2), .B(a_reg_25_), .Y(_abc_15724_n5702) );
  AND2X2 AND2X2_2444 ( .A(_abc_15724_n2994_bF_buf2), .B(_abc_15724_n2885), .Y(_abc_15724_n5703) );
  AND2X2 AND2X2_2445 ( .A(_abc_15724_n5698), .B(_abc_15724_n5689), .Y(_abc_15724_n5706) );
  AND2X2 AND2X2_2446 ( .A(_abc_15724_n5696), .B(_abc_15724_n5706), .Y(_abc_15724_n5707) );
  AND2X2 AND2X2_2447 ( .A(_abc_15724_n5681), .B(_abc_15724_n5677), .Y(_abc_15724_n5709) );
  AND2X2 AND2X2_2448 ( .A(c_reg_26_), .B(b_reg_26_), .Y(_abc_15724_n5711) );
  AND2X2 AND2X2_2449 ( .A(_abc_15724_n5714), .B(_abc_15724_n5712), .Y(_abc_15724_n5715) );
  AND2X2 AND2X2_245 ( .A(_abc_15724_n1180), .B(_abc_15724_n1193_1), .Y(_abc_15724_n1196) );
  AND2X2 AND2X2_2450 ( .A(_abc_15724_n3805_bF_buf2), .B(_abc_15724_n5715), .Y(_abc_15724_n5716) );
  AND2X2 AND2X2_2451 ( .A(_abc_15724_n5712), .B(_abc_15724_n5718), .Y(_abc_15724_n5719) );
  AND2X2 AND2X2_2452 ( .A(_abc_15724_n5719), .B(d_reg_26_), .Y(_abc_15724_n5721) );
  AND2X2 AND2X2_2453 ( .A(_abc_15724_n5722), .B(_abc_15724_n5720), .Y(_abc_15724_n5723) );
  AND2X2 AND2X2_2454 ( .A(_abc_15724_n3726_bF_buf3), .B(_abc_15724_n5723), .Y(_abc_15724_n5724) );
  AND2X2 AND2X2_2455 ( .A(_abc_15724_n5712), .B(_abc_15724_n5713), .Y(_abc_15724_n5725) );
  AND2X2 AND2X2_2456 ( .A(_abc_15724_n3737_bF_buf1), .B(_abc_15724_n5728), .Y(_abc_15724_n5729) );
  AND2X2 AND2X2_2457 ( .A(_abc_15724_n5731), .B(_abc_15724_n5717), .Y(_abc_15724_n5732) );
  AND2X2 AND2X2_2458 ( .A(_abc_15724_n5673), .B(_abc_15724_n5670), .Y(_abc_15724_n5733) );
  AND2X2 AND2X2_2459 ( .A(e_reg_26_), .B(a_reg_21_), .Y(_abc_15724_n5736) );
  AND2X2 AND2X2_246 ( .A(_abc_15724_n1176), .B(_abc_15724_n1196), .Y(_abc_15724_n1197_1) );
  AND2X2 AND2X2_2460 ( .A(_abc_15724_n5737), .B(_abc_15724_n5735), .Y(_abc_15724_n5738) );
  AND2X2 AND2X2_2461 ( .A(_abc_15724_n5738), .B(w_26_), .Y(_abc_15724_n5739) );
  AND2X2 AND2X2_2462 ( .A(_abc_15724_n5740), .B(_abc_15724_n5741), .Y(_abc_15724_n5742) );
  AND2X2 AND2X2_2463 ( .A(_abc_15724_n5734), .B(_abc_15724_n5742), .Y(_abc_15724_n5743) );
  AND2X2 AND2X2_2464 ( .A(_abc_15724_n5744), .B(_abc_15724_n5745), .Y(_abc_15724_n5746) );
  AND2X2 AND2X2_2465 ( .A(_abc_15724_n5732), .B(_abc_15724_n5746), .Y(_abc_15724_n5747) );
  AND2X2 AND2X2_2466 ( .A(_abc_15724_n5748), .B(_abc_15724_n5749), .Y(_abc_15724_n5750) );
  AND2X2 AND2X2_2467 ( .A(_abc_15724_n5710), .B(_abc_15724_n5750), .Y(_abc_15724_n5751) );
  AND2X2 AND2X2_2468 ( .A(_abc_15724_n5752), .B(_abc_15724_n5753), .Y(_abc_15724_n5754) );
  AND2X2 AND2X2_2469 ( .A(_abc_15724_n5755), .B(_abc_15724_n5006), .Y(_abc_15724_n5756) );
  AND2X2 AND2X2_247 ( .A(_abc_15724_n1193_1), .B(_abc_15724_n1178_1), .Y(_abc_15724_n1198_1) );
  AND2X2 AND2X2_2470 ( .A(_abc_15724_n5754), .B(_abc_15724_n5056), .Y(_abc_15724_n5757) );
  AND2X2 AND2X2_2471 ( .A(_abc_15724_n5759), .B(_abc_15724_n5685), .Y(_abc_15724_n5760) );
  AND2X2 AND2X2_2472 ( .A(_abc_15724_n5758), .B(_abc_15724_n5686), .Y(_abc_15724_n5761) );
  AND2X2 AND2X2_2473 ( .A(_abc_15724_n5765), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n5766) );
  AND2X2 AND2X2_2474 ( .A(_abc_15724_n5766), .B(_abc_15724_n5764), .Y(_abc_15724_n5767) );
  AND2X2 AND2X2_2475 ( .A(_abc_15724_n2992_bF_buf1), .B(a_reg_26_), .Y(_abc_15724_n5768) );
  AND2X2 AND2X2_2476 ( .A(_abc_15724_n2994_bF_buf1), .B(_abc_15724_n2902), .Y(_abc_15724_n5769) );
  AND2X2 AND2X2_2477 ( .A(_abc_15724_n5765), .B(_abc_15724_n5772), .Y(_abc_15724_n5773) );
  AND2X2 AND2X2_2478 ( .A(_abc_15724_n5748), .B(_abc_15724_n5744), .Y(_abc_15724_n5776) );
  AND2X2 AND2X2_2479 ( .A(c_reg_27_), .B(b_reg_27_), .Y(_abc_15724_n5778) );
  AND2X2 AND2X2_248 ( .A(_abc_15724_n1200_1), .B(digest_update_bF_buf11), .Y(_abc_15724_n1201) );
  AND2X2 AND2X2_2480 ( .A(_abc_15724_n5781), .B(_abc_15724_n5779), .Y(_abc_15724_n5782) );
  AND2X2 AND2X2_2481 ( .A(_abc_15724_n3805_bF_buf0), .B(_abc_15724_n5782), .Y(_abc_15724_n5783) );
  AND2X2 AND2X2_2482 ( .A(_abc_15724_n5779), .B(_abc_15724_n5785), .Y(_abc_15724_n5786) );
  AND2X2 AND2X2_2483 ( .A(_abc_15724_n5786), .B(d_reg_27_), .Y(_abc_15724_n5788) );
  AND2X2 AND2X2_2484 ( .A(_abc_15724_n5789), .B(_abc_15724_n5787), .Y(_abc_15724_n5790) );
  AND2X2 AND2X2_2485 ( .A(_abc_15724_n3726_bF_buf2), .B(_abc_15724_n5790), .Y(_abc_15724_n5791) );
  AND2X2 AND2X2_2486 ( .A(_abc_15724_n5779), .B(_abc_15724_n5780), .Y(_abc_15724_n5792) );
  AND2X2 AND2X2_2487 ( .A(_abc_15724_n3737_bF_buf0), .B(_abc_15724_n5795), .Y(_abc_15724_n5796) );
  AND2X2 AND2X2_2488 ( .A(_abc_15724_n5798), .B(_abc_15724_n5784), .Y(_abc_15724_n5799) );
  AND2X2 AND2X2_2489 ( .A(_abc_15724_n5740), .B(_abc_15724_n5737), .Y(_abc_15724_n5800) );
  AND2X2 AND2X2_249 ( .A(_abc_15724_n1201), .B(_abc_15724_n1195), .Y(_abc_15724_n1202) );
  AND2X2 AND2X2_2490 ( .A(e_reg_27_), .B(a_reg_22_), .Y(_abc_15724_n5803) );
  AND2X2 AND2X2_2491 ( .A(_abc_15724_n5804), .B(_abc_15724_n5802), .Y(_abc_15724_n5805) );
  AND2X2 AND2X2_2492 ( .A(_abc_15724_n5805), .B(w_27_), .Y(_abc_15724_n5806) );
  AND2X2 AND2X2_2493 ( .A(_abc_15724_n5807), .B(_abc_15724_n5808), .Y(_abc_15724_n5809) );
  AND2X2 AND2X2_2494 ( .A(_abc_15724_n5801), .B(_abc_15724_n5809), .Y(_abc_15724_n5810) );
  AND2X2 AND2X2_2495 ( .A(_abc_15724_n5811), .B(_abc_15724_n5812), .Y(_abc_15724_n5813) );
  AND2X2 AND2X2_2496 ( .A(_abc_15724_n5799), .B(_abc_15724_n5813), .Y(_abc_15724_n5814) );
  AND2X2 AND2X2_2497 ( .A(_abc_15724_n5815), .B(_abc_15724_n5816), .Y(_abc_15724_n5817) );
  AND2X2 AND2X2_2498 ( .A(_abc_15724_n5777), .B(_abc_15724_n5817), .Y(_abc_15724_n5818) );
  AND2X2 AND2X2_2499 ( .A(_abc_15724_n5775), .B(_abc_15724_n5821), .Y(_abc_15724_n5822) );
  AND2X2 AND2X2_25 ( .A(_abc_15724_n745), .B(_abc_15724_n737), .Y(_abc_15724_n746) );
  AND2X2 AND2X2_250 ( .A(_abc_15724_n1200_1), .B(_abc_15724_n1192), .Y(_abc_15724_n1204) );
  AND2X2 AND2X2_2500 ( .A(_abc_15724_n5823), .B(_abc_15724_n5824), .Y(_abc_15724_n5825) );
  AND2X2 AND2X2_2501 ( .A(_abc_15724_n5828), .B(round_ctr_inc_bF_buf12), .Y(_abc_15724_n5829) );
  AND2X2 AND2X2_2502 ( .A(_abc_15724_n5829), .B(_abc_15724_n5826), .Y(_abc_15724_n5830) );
  AND2X2 AND2X2_2503 ( .A(_abc_15724_n2992_bF_buf0), .B(a_reg_27_), .Y(_abc_15724_n5831) );
  AND2X2 AND2X2_2504 ( .A(_abc_15724_n906_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_155_), .Y(_abc_15724_n5832) );
  AND2X2 AND2X2_2505 ( .A(_abc_15724_n2994_bF_buf0), .B(_abc_15724_n5832), .Y(_abc_15724_n5833) );
  AND2X2 AND2X2_2506 ( .A(_abc_15724_n5763), .B(_abc_15724_n5825), .Y(_abc_15724_n5836) );
  AND2X2 AND2X2_2507 ( .A(_abc_15724_n5694), .B(_abc_15724_n5836), .Y(_abc_15724_n5837) );
  AND2X2 AND2X2_2508 ( .A(_abc_15724_n5840), .B(_abc_15724_n5836), .Y(_abc_15724_n5841) );
  AND2X2 AND2X2_2509 ( .A(_abc_15724_n5843), .B(_abc_15724_n5823), .Y(_abc_15724_n5844) );
  AND2X2 AND2X2_251 ( .A(_auto_iopadmap_cc_313_execute_26059_46_), .B(d_reg_14_), .Y(_abc_15724_n1207_1) );
  AND2X2 AND2X2_2510 ( .A(_abc_15724_n5842), .B(_abc_15724_n5844), .Y(_abc_15724_n5845) );
  AND2X2 AND2X2_2511 ( .A(_abc_15724_n5839), .B(_abc_15724_n5845), .Y(_abc_15724_n5846) );
  AND2X2 AND2X2_2512 ( .A(_abc_15724_n5815), .B(_abc_15724_n5811), .Y(_abc_15724_n5848) );
  AND2X2 AND2X2_2513 ( .A(c_reg_28_), .B(b_reg_28_), .Y(_abc_15724_n5850) );
  AND2X2 AND2X2_2514 ( .A(_abc_15724_n5853), .B(_abc_15724_n5851), .Y(_abc_15724_n5854) );
  AND2X2 AND2X2_2515 ( .A(_abc_15724_n3805_bF_buf3), .B(_abc_15724_n5854), .Y(_abc_15724_n5855) );
  AND2X2 AND2X2_2516 ( .A(_abc_15724_n5851), .B(_abc_15724_n5857), .Y(_abc_15724_n5858) );
  AND2X2 AND2X2_2517 ( .A(_abc_15724_n5858), .B(d_reg_28_), .Y(_abc_15724_n5860) );
  AND2X2 AND2X2_2518 ( .A(_abc_15724_n5861), .B(_abc_15724_n5859), .Y(_abc_15724_n5862) );
  AND2X2 AND2X2_2519 ( .A(_abc_15724_n3726_bF_buf1), .B(_abc_15724_n5862), .Y(_abc_15724_n5863) );
  AND2X2 AND2X2_252 ( .A(_abc_15724_n1208), .B(_abc_15724_n1206_1), .Y(_abc_15724_n1209_1) );
  AND2X2 AND2X2_2520 ( .A(_abc_15724_n5851), .B(_abc_15724_n5852), .Y(_abc_15724_n5864) );
  AND2X2 AND2X2_2521 ( .A(_abc_15724_n3737_bF_buf4), .B(_abc_15724_n5867), .Y(_abc_15724_n5868) );
  AND2X2 AND2X2_2522 ( .A(_abc_15724_n5870), .B(_abc_15724_n5856), .Y(_abc_15724_n5871) );
  AND2X2 AND2X2_2523 ( .A(_abc_15724_n5807), .B(_abc_15724_n5804), .Y(_abc_15724_n5872) );
  AND2X2 AND2X2_2524 ( .A(e_reg_28_), .B(a_reg_23_), .Y(_abc_15724_n5875) );
  AND2X2 AND2X2_2525 ( .A(_abc_15724_n5876), .B(_abc_15724_n5874), .Y(_abc_15724_n5877) );
  AND2X2 AND2X2_2526 ( .A(_abc_15724_n5877), .B(w_28_), .Y(_abc_15724_n5878) );
  AND2X2 AND2X2_2527 ( .A(_abc_15724_n5879), .B(_abc_15724_n5880), .Y(_abc_15724_n5881) );
  AND2X2 AND2X2_2528 ( .A(_abc_15724_n5873), .B(_abc_15724_n5881), .Y(_abc_15724_n5882) );
  AND2X2 AND2X2_2529 ( .A(_abc_15724_n5883), .B(_abc_15724_n5884), .Y(_abc_15724_n5885) );
  AND2X2 AND2X2_253 ( .A(_abc_15724_n1205), .B(_abc_15724_n1209_1), .Y(_abc_15724_n1211) );
  AND2X2 AND2X2_2530 ( .A(_abc_15724_n5871), .B(_abc_15724_n5885), .Y(_abc_15724_n5886) );
  AND2X2 AND2X2_2531 ( .A(_abc_15724_n5887), .B(_abc_15724_n5888), .Y(_abc_15724_n5889) );
  AND2X2 AND2X2_2532 ( .A(_abc_15724_n5849), .B(_abc_15724_n5889), .Y(_abc_15724_n5890) );
  AND2X2 AND2X2_2533 ( .A(_abc_15724_n5891), .B(_abc_15724_n5892), .Y(_abc_15724_n5893) );
  AND2X2 AND2X2_2534 ( .A(_abc_15724_n5893), .B(_abc_15724_n3805_bF_buf1), .Y(_abc_15724_n5894) );
  AND2X2 AND2X2_2535 ( .A(_abc_15724_n5895), .B(_abc_15724_n5896), .Y(_abc_15724_n5897) );
  AND2X2 AND2X2_2536 ( .A(_abc_15724_n5897), .B(_abc_15724_n5819), .Y(_abc_15724_n5898) );
  AND2X2 AND2X2_2537 ( .A(_abc_15724_n5899), .B(_abc_15724_n5900), .Y(_abc_15724_n5901) );
  AND2X2 AND2X2_2538 ( .A(_abc_15724_n5847), .B(_abc_15724_n5901), .Y(_abc_15724_n5903) );
  AND2X2 AND2X2_2539 ( .A(_abc_15724_n5904), .B(round_ctr_inc_bF_buf11), .Y(_abc_15724_n5905) );
  AND2X2 AND2X2_254 ( .A(_abc_15724_n1212), .B(_abc_15724_n1210), .Y(_abc_15724_n1213) );
  AND2X2 AND2X2_2540 ( .A(_abc_15724_n5905), .B(_abc_15724_n5902), .Y(_abc_15724_n5906) );
  AND2X2 AND2X2_2541 ( .A(_abc_15724_n2992_bF_buf11), .B(a_reg_28_), .Y(_abc_15724_n5907) );
  AND2X2 AND2X2_2542 ( .A(_abc_15724_n906_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_156_), .Y(_abc_15724_n5908) );
  AND2X2 AND2X2_2543 ( .A(_abc_15724_n2994_bF_buf11), .B(_abc_15724_n5908), .Y(_abc_15724_n5909) );
  AND2X2 AND2X2_2544 ( .A(_abc_15724_n5895), .B(_abc_15724_n5891), .Y(_abc_15724_n5912) );
  AND2X2 AND2X2_2545 ( .A(_abc_15724_n5887), .B(_abc_15724_n5883), .Y(_abc_15724_n5914) );
  AND2X2 AND2X2_2546 ( .A(c_reg_29_), .B(b_reg_29_), .Y(_abc_15724_n5916) );
  AND2X2 AND2X2_2547 ( .A(_abc_15724_n5919), .B(_abc_15724_n5917), .Y(_abc_15724_n5920) );
  AND2X2 AND2X2_2548 ( .A(_abc_15724_n3805_bF_buf4), .B(_abc_15724_n5920), .Y(_abc_15724_n5921) );
  AND2X2 AND2X2_2549 ( .A(_abc_15724_n5917), .B(_abc_15724_n5923), .Y(_abc_15724_n5924) );
  AND2X2 AND2X2_255 ( .A(_abc_15724_n1213), .B(digest_update_bF_buf10), .Y(_abc_15724_n1214) );
  AND2X2 AND2X2_2550 ( .A(_abc_15724_n5924), .B(d_reg_29_), .Y(_abc_15724_n5926) );
  AND2X2 AND2X2_2551 ( .A(_abc_15724_n5927), .B(_abc_15724_n5925), .Y(_abc_15724_n5928) );
  AND2X2 AND2X2_2552 ( .A(_abc_15724_n3726_bF_buf0), .B(_abc_15724_n5928), .Y(_abc_15724_n5929) );
  AND2X2 AND2X2_2553 ( .A(_abc_15724_n5917), .B(_abc_15724_n5918), .Y(_abc_15724_n5930) );
  AND2X2 AND2X2_2554 ( .A(_abc_15724_n3737_bF_buf3), .B(_abc_15724_n5933), .Y(_abc_15724_n5934) );
  AND2X2 AND2X2_2555 ( .A(_abc_15724_n5936), .B(_abc_15724_n5922), .Y(_abc_15724_n5937) );
  AND2X2 AND2X2_2556 ( .A(_abc_15724_n5879), .B(_abc_15724_n5876), .Y(_abc_15724_n5938) );
  AND2X2 AND2X2_2557 ( .A(e_reg_29_), .B(a_reg_24_), .Y(_abc_15724_n5941) );
  AND2X2 AND2X2_2558 ( .A(_abc_15724_n5942), .B(_abc_15724_n5940), .Y(_abc_15724_n5943) );
  AND2X2 AND2X2_2559 ( .A(_abc_15724_n5943), .B(w_29_), .Y(_abc_15724_n5944) );
  AND2X2 AND2X2_256 ( .A(_abc_15724_n1215_1), .B(_abc_15724_n850_bF_buf1), .Y(_abc_15724_n1216_1) );
  AND2X2 AND2X2_2560 ( .A(_abc_15724_n5945), .B(_abc_15724_n5946), .Y(_abc_15724_n5947) );
  AND2X2 AND2X2_2561 ( .A(_abc_15724_n5939), .B(_abc_15724_n5947), .Y(_abc_15724_n5948) );
  AND2X2 AND2X2_2562 ( .A(_abc_15724_n5949), .B(_abc_15724_n5950), .Y(_abc_15724_n5951) );
  AND2X2 AND2X2_2563 ( .A(_abc_15724_n5937), .B(_abc_15724_n5951), .Y(_abc_15724_n5952) );
  AND2X2 AND2X2_2564 ( .A(_abc_15724_n5953), .B(_abc_15724_n5954), .Y(_abc_15724_n5955) );
  AND2X2 AND2X2_2565 ( .A(_abc_15724_n5915), .B(_abc_15724_n5955), .Y(_abc_15724_n5956) );
  AND2X2 AND2X2_2566 ( .A(_abc_15724_n5957), .B(_abc_15724_n5958), .Y(_abc_15724_n5959) );
  AND2X2 AND2X2_2567 ( .A(_abc_15724_n5959), .B(_abc_15724_n4021), .Y(_abc_15724_n5960) );
  AND2X2 AND2X2_2568 ( .A(_abc_15724_n5961), .B(_abc_15724_n5962), .Y(_abc_15724_n5963) );
  AND2X2 AND2X2_2569 ( .A(_abc_15724_n5913), .B(_abc_15724_n5963), .Y(_abc_15724_n5964) );
  AND2X2 AND2X2_257 ( .A(_abc_15724_n1212), .B(_abc_15724_n1208), .Y(_abc_15724_n1218_1) );
  AND2X2 AND2X2_2570 ( .A(_abc_15724_n5965), .B(_abc_15724_n5966), .Y(_abc_15724_n5967) );
  AND2X2 AND2X2_2571 ( .A(_abc_15724_n5967), .B(_abc_15724_n5901), .Y(_abc_15724_n5970) );
  AND2X2 AND2X2_2572 ( .A(_abc_15724_n5967), .B(_abc_15724_n5898), .Y(_abc_15724_n5973) );
  AND2X2 AND2X2_2573 ( .A(_abc_15724_n5974), .B(round_ctr_inc_bF_buf10), .Y(_abc_15724_n5975) );
  AND2X2 AND2X2_2574 ( .A(_abc_15724_n5972), .B(_abc_15724_n5975), .Y(_abc_15724_n5976) );
  AND2X2 AND2X2_2575 ( .A(_abc_15724_n5969), .B(_abc_15724_n5976), .Y(_abc_15724_n5977) );
  AND2X2 AND2X2_2576 ( .A(_abc_15724_n2992_bF_buf10), .B(a_reg_29_), .Y(_abc_15724_n5978) );
  AND2X2 AND2X2_2577 ( .A(_abc_15724_n2994_bF_buf10), .B(_abc_15724_n2952), .Y(_abc_15724_n5979) );
  AND2X2 AND2X2_2578 ( .A(_abc_15724_n5974), .B(_abc_15724_n5965), .Y(_abc_15724_n5982) );
  AND2X2 AND2X2_2579 ( .A(_abc_15724_n5972), .B(_abc_15724_n5982), .Y(_abc_15724_n5983) );
  AND2X2 AND2X2_258 ( .A(_auto_iopadmap_cc_313_execute_26059_47_), .B(d_reg_15_), .Y(_abc_15724_n1220) );
  AND2X2 AND2X2_2580 ( .A(_abc_15724_n5961), .B(_abc_15724_n5957), .Y(_abc_15724_n5985) );
  AND2X2 AND2X2_2581 ( .A(_abc_15724_n5953), .B(_abc_15724_n5949), .Y(_abc_15724_n5987) );
  AND2X2 AND2X2_2582 ( .A(c_reg_30_), .B(b_reg_30_), .Y(_abc_15724_n5989) );
  AND2X2 AND2X2_2583 ( .A(_abc_15724_n5992), .B(_abc_15724_n5990), .Y(_abc_15724_n5993) );
  AND2X2 AND2X2_2584 ( .A(_abc_15724_n3805_bF_buf2), .B(_abc_15724_n5993), .Y(_abc_15724_n5994) );
  AND2X2 AND2X2_2585 ( .A(_abc_15724_n5990), .B(_abc_15724_n5996), .Y(_abc_15724_n5997) );
  AND2X2 AND2X2_2586 ( .A(_abc_15724_n5997), .B(d_reg_30_), .Y(_abc_15724_n5999) );
  AND2X2 AND2X2_2587 ( .A(_abc_15724_n6000), .B(_abc_15724_n5998), .Y(_abc_15724_n6001) );
  AND2X2 AND2X2_2588 ( .A(_abc_15724_n3726_bF_buf4), .B(_abc_15724_n6001), .Y(_abc_15724_n6002) );
  AND2X2 AND2X2_2589 ( .A(_abc_15724_n5990), .B(_abc_15724_n5991), .Y(_abc_15724_n6003) );
  AND2X2 AND2X2_259 ( .A(_abc_15724_n1221), .B(_abc_15724_n1219), .Y(_abc_15724_n1222) );
  AND2X2 AND2X2_2590 ( .A(_abc_15724_n3737_bF_buf2), .B(_abc_15724_n6006), .Y(_abc_15724_n6007) );
  AND2X2 AND2X2_2591 ( .A(_abc_15724_n6009), .B(_abc_15724_n5995), .Y(_abc_15724_n6010) );
  AND2X2 AND2X2_2592 ( .A(_abc_15724_n5945), .B(_abc_15724_n5942), .Y(_abc_15724_n6011) );
  AND2X2 AND2X2_2593 ( .A(e_reg_30_), .B(a_reg_25_), .Y(_abc_15724_n6014) );
  AND2X2 AND2X2_2594 ( .A(_abc_15724_n6015), .B(_abc_15724_n6013), .Y(_abc_15724_n6016) );
  AND2X2 AND2X2_2595 ( .A(_abc_15724_n6016), .B(w_30_), .Y(_abc_15724_n6017) );
  AND2X2 AND2X2_2596 ( .A(_abc_15724_n6018), .B(_abc_15724_n6019), .Y(_abc_15724_n6020) );
  AND2X2 AND2X2_2597 ( .A(_abc_15724_n6012), .B(_abc_15724_n6020), .Y(_abc_15724_n6021) );
  AND2X2 AND2X2_2598 ( .A(_abc_15724_n6022), .B(_abc_15724_n6023), .Y(_abc_15724_n6024) );
  AND2X2 AND2X2_2599 ( .A(_abc_15724_n6010), .B(_abc_15724_n6024), .Y(_abc_15724_n6025) );
  AND2X2 AND2X2_26 ( .A(_abc_15724_n731_1), .B(_abc_15724_n733), .Y(_abc_15724_n747) );
  AND2X2 AND2X2_260 ( .A(_abc_15724_n1218_1), .B(_abc_15724_n1222), .Y(_abc_15724_n1223) );
  AND2X2 AND2X2_2600 ( .A(_abc_15724_n6026), .B(_abc_15724_n6027), .Y(_abc_15724_n6028) );
  AND2X2 AND2X2_2601 ( .A(_abc_15724_n5988), .B(_abc_15724_n6028), .Y(_abc_15724_n6029) );
  AND2X2 AND2X2_2602 ( .A(_abc_15724_n6030), .B(_abc_15724_n6031), .Y(_abc_15724_n6032) );
  AND2X2 AND2X2_2603 ( .A(_abc_15724_n6032), .B(_abc_15724_n3725_bF_buf1), .Y(_abc_15724_n6033) );
  AND2X2 AND2X2_2604 ( .A(_abc_15724_n6034), .B(_abc_15724_n6035), .Y(_abc_15724_n6036) );
  AND2X2 AND2X2_2605 ( .A(_abc_15724_n5986), .B(_abc_15724_n6036), .Y(_abc_15724_n6037) );
  AND2X2 AND2X2_2606 ( .A(_abc_15724_n6038), .B(_abc_15724_n6039), .Y(_abc_15724_n6040) );
  AND2X2 AND2X2_2607 ( .A(_abc_15724_n6043), .B(round_ctr_inc_bF_buf9), .Y(_abc_15724_n6044) );
  AND2X2 AND2X2_2608 ( .A(_abc_15724_n6044), .B(_abc_15724_n6041), .Y(_abc_15724_n6045) );
  AND2X2 AND2X2_2609 ( .A(_abc_15724_n2992_bF_buf9), .B(a_reg_30_), .Y(_abc_15724_n6046) );
  AND2X2 AND2X2_261 ( .A(_abc_15724_n1224), .B(_abc_15724_n1225), .Y(_abc_15724_n1226) );
  AND2X2 AND2X2_2610 ( .A(_abc_15724_n2994_bF_buf9), .B(_abc_15724_n2972), .Y(_abc_15724_n6047) );
  AND2X2 AND2X2_2611 ( .A(_abc_15724_n6043), .B(_abc_15724_n6038), .Y(_abc_15724_n6050) );
  AND2X2 AND2X2_2612 ( .A(_abc_15724_n6034), .B(_abc_15724_n6030), .Y(_abc_15724_n6052) );
  AND2X2 AND2X2_2613 ( .A(_abc_15724_n6026), .B(_abc_15724_n6022), .Y(_abc_15724_n6053) );
  AND2X2 AND2X2_2614 ( .A(c_reg_31_), .B(b_reg_31_), .Y(_abc_15724_n6055) );
  AND2X2 AND2X2_2615 ( .A(_abc_15724_n6058), .B(_abc_15724_n6056), .Y(_abc_15724_n6059) );
  AND2X2 AND2X2_2616 ( .A(_abc_15724_n3805_bF_buf0), .B(_abc_15724_n6059), .Y(_abc_15724_n6060) );
  AND2X2 AND2X2_2617 ( .A(_abc_15724_n2003), .B(_abc_15724_n2480), .Y(_abc_15724_n6061) );
  AND2X2 AND2X2_2618 ( .A(_abc_15724_n6062), .B(_abc_15724_n6057), .Y(_abc_15724_n6063) );
  AND2X2 AND2X2_2619 ( .A(_abc_15724_n6056), .B(_abc_15724_n6057), .Y(_abc_15724_n6064) );
  AND2X2 AND2X2_262 ( .A(_abc_15724_n1227), .B(digest_update_bF_buf9), .Y(_abc_15724_n1228_1) );
  AND2X2 AND2X2_2620 ( .A(_abc_15724_n6066), .B(_abc_15724_n6056), .Y(_abc_15724_n6067) );
  AND2X2 AND2X2_2621 ( .A(_abc_15724_n3737_bF_buf1), .B(_abc_15724_n6066), .Y(_abc_15724_n6070) );
  AND2X2 AND2X2_2622 ( .A(_abc_15724_n6069), .B(_abc_15724_n6072), .Y(_abc_15724_n6073) );
  AND2X2 AND2X2_2623 ( .A(_abc_15724_n6018), .B(_abc_15724_n6015), .Y(_abc_15724_n6075) );
  AND2X2 AND2X2_2624 ( .A(e_reg_31_), .B(w_31_), .Y(_abc_15724_n6077) );
  AND2X2 AND2X2_2625 ( .A(_abc_15724_n6078), .B(_abc_15724_n6076), .Y(_abc_15724_n6079) );
  AND2X2 AND2X2_2626 ( .A(_abc_15724_n6079), .B(a_reg_26_), .Y(_abc_15724_n6080) );
  AND2X2 AND2X2_2627 ( .A(_abc_15724_n6081), .B(_abc_15724_n6082), .Y(_abc_15724_n6083) );
  AND2X2 AND2X2_2628 ( .A(_abc_15724_n6084), .B(_abc_15724_n6075), .Y(_abc_15724_n6085) );
  AND2X2 AND2X2_2629 ( .A(_abc_15724_n6086), .B(_abc_15724_n6087), .Y(_abc_15724_n6088) );
  AND2X2 AND2X2_263 ( .A(_abc_15724_n907_1_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_47_), .Y(_abc_15724_n1229_1) );
  AND2X2 AND2X2_2630 ( .A(_abc_15724_n6092), .B(_abc_15724_n6089), .Y(_abc_15724_n6093) );
  AND2X2 AND2X2_2631 ( .A(_abc_15724_n6094), .B(_abc_15724_n6054), .Y(_abc_15724_n6095) );
  AND2X2 AND2X2_2632 ( .A(_abc_15724_n6093), .B(_abc_15724_n6053), .Y(_abc_15724_n6096) );
  AND2X2 AND2X2_2633 ( .A(_abc_15724_n6099), .B(_abc_15724_n6100), .Y(_abc_15724_n6101) );
  AND2X2 AND2X2_2634 ( .A(_abc_15724_n6101), .B(_abc_15724_n6052), .Y(_abc_15724_n6102) );
  AND2X2 AND2X2_2635 ( .A(_abc_15724_n6103), .B(_abc_15724_n6104), .Y(_abc_15724_n6105) );
  AND2X2 AND2X2_2636 ( .A(_abc_15724_n6108), .B(round_ctr_inc_bF_buf8), .Y(_abc_15724_n6109) );
  AND2X2 AND2X2_2637 ( .A(_abc_15724_n6109), .B(_abc_15724_n6107), .Y(_abc_15724_n6110) );
  AND2X2 AND2X2_2638 ( .A(_abc_15724_n2992_bF_buf8), .B(a_reg_31_), .Y(_abc_15724_n6111) );
  AND2X2 AND2X2_2639 ( .A(_abc_15724_n906_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_159_), .Y(_abc_15724_n6112) );
  AND2X2 AND2X2_264 ( .A(_abc_15724_n907_1_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_48_), .Y(_abc_15724_n1231_1) );
  AND2X2 AND2X2_2640 ( .A(_abc_15724_n2994_bF_buf8), .B(_abc_15724_n6112), .Y(_abc_15724_n6113) );
  AND2X2 AND2X2_2641 ( .A(round_ctr_reg_1_), .B(round_ctr_reg_0_), .Y(_abc_15724_n6119) );
  AND2X2 AND2X2_2642 ( .A(_abc_15724_n3722), .B(_abc_15724_n6119), .Y(_abc_15724_n6120) );
  AND2X2 AND2X2_2643 ( .A(_abc_15724_n6120), .B(round_ctr_inc_bF_buf7), .Y(_abc_15724_n6121) );
  AND2X2 AND2X2_2644 ( .A(_abc_15724_n6121), .B(_abc_15724_n6118), .Y(_abc_15724_n3465) );
  AND2X2 AND2X2_2645 ( .A(_abc_15724_n6124), .B(round_ctr_inc_bF_buf6), .Y(_abc_15724_n6125) );
  AND2X2 AND2X2_2646 ( .A(_abc_15724_n6125), .B(_abc_15724_n907_1_bF_buf7), .Y(_abc_15724_n6126) );
  AND2X2 AND2X2_2647 ( .A(_abc_15724_n6129), .B(_auto_iopadmap_cc_313_execute_26222), .Y(_abc_15724_n6130) );
  AND2X2 AND2X2_2648 ( .A(_abc_15724_n2991), .B(_auto_iopadmap_cc_313_execute_26220), .Y(_abc_15724_n6132) );
  AND2X2 AND2X2_2649 ( .A(_abc_15724_n6135), .B(_abc_15724_n6136), .Y(round_ctr_reg_0__FF_INPUT) );
  AND2X2 AND2X2_265 ( .A(_abc_15724_n1209_1), .B(_abc_15724_n1222), .Y(_abc_15724_n1232) );
  AND2X2 AND2X2_2650 ( .A(_abc_15724_n2992_bF_buf6), .B(round_ctr_reg_1_), .Y(_abc_15724_n6138) );
  AND2X2 AND2X2_2651 ( .A(_abc_15724_n6139), .B(_abc_15724_n6140), .Y(_abc_15724_n6141) );
  AND2X2 AND2X2_2652 ( .A(_abc_15724_n6141), .B(round_ctr_inc_bF_buf4), .Y(_abc_15724_n6142) );
  AND2X2 AND2X2_2653 ( .A(_abc_15724_n2992_bF_buf5), .B(round_ctr_reg_2_), .Y(_abc_15724_n6144) );
  AND2X2 AND2X2_2654 ( .A(_abc_15724_n6119), .B(round_ctr_reg_2_), .Y(_abc_15724_n6145) );
  AND2X2 AND2X2_2655 ( .A(_abc_15724_n6146), .B(_abc_15724_n6147), .Y(_abc_15724_n6148) );
  AND2X2 AND2X2_2656 ( .A(_abc_15724_n6148), .B(round_ctr_inc_bF_buf3), .Y(_abc_15724_n6149) );
  AND2X2 AND2X2_2657 ( .A(_abc_15724_n2992_bF_buf4), .B(round_ctr_reg_3_), .Y(_abc_15724_n6151) );
  AND2X2 AND2X2_2658 ( .A(_abc_15724_n6152), .B(_abc_15724_n6123), .Y(_abc_15724_n6153) );
  AND2X2 AND2X2_2659 ( .A(_abc_15724_n6153), .B(round_ctr_inc_bF_buf2), .Y(_abc_15724_n6154) );
  AND2X2 AND2X2_266 ( .A(_abc_15724_n1196), .B(_abc_15724_n1232), .Y(_abc_15724_n1233) );
  AND2X2 AND2X2_2660 ( .A(_abc_15724_n6121), .B(round_ctr_reg_4_), .Y(_abc_15724_n6156) );
  AND2X2 AND2X2_2661 ( .A(_abc_15724_n6158), .B(round_ctr_reg_4_), .Y(_abc_15724_n6159) );
  AND2X2 AND2X2_2662 ( .A(_abc_15724_n6160), .B(_abc_15724_n6157), .Y(round_ctr_reg_4__FF_INPUT) );
  AND2X2 AND2X2_2663 ( .A(_abc_15724_n6120), .B(_abc_15724_n3700), .Y(_abc_15724_n6162) );
  AND2X2 AND2X2_2664 ( .A(round_ctr_inc_bF_buf1), .B(round_ctr_reg_5_), .Y(_abc_15724_n6164) );
  AND2X2 AND2X2_2665 ( .A(_abc_15724_n6165), .B(_abc_15724_n6163), .Y(_abc_15724_n6166) );
  AND2X2 AND2X2_2666 ( .A(_abc_15724_n2992_bF_buf3), .B(round_ctr_reg_5_), .Y(_abc_15724_n6167) );
  AND2X2 AND2X2_2667 ( .A(_abc_15724_n6158), .B(round_ctr_reg_6_), .Y(_abc_15724_n6169) );
  AND2X2 AND2X2_2668 ( .A(_abc_15724_n6162), .B(round_ctr_inc_bF_buf0), .Y(_abc_15724_n6170) );
  AND2X2 AND2X2_2669 ( .A(_abc_15724_n6170), .B(round_ctr_reg_6_), .Y(_abc_15724_n6172) );
  AND2X2 AND2X2_267 ( .A(_abc_15724_n1172), .B(_abc_15724_n1233), .Y(_abc_15724_n1234) );
  AND2X2 AND2X2_2670 ( .A(_abc_15724_n6171), .B(_abc_15724_n6173), .Y(round_ctr_reg_6__FF_INPUT) );
  AND2X2 AND2X2_2671 ( .A(_abc_15724_n6175), .B(_abc_15724_n6176), .Y(_abc_15724_n6177) );
  AND2X2 AND2X2_2672 ( .A(_abc_15724_n6178), .B(_abc_15724_n6179), .Y(H4_reg_0__FF_INPUT) );
  AND2X2 AND2X2_2673 ( .A(_abc_15724_n796), .B(_abc_15724_n6181), .Y(_abc_15724_n6182) );
  AND2X2 AND2X2_2674 ( .A(_abc_15724_n6182), .B(digest_update_bF_buf1), .Y(_abc_15724_n6183) );
  AND2X2 AND2X2_2675 ( .A(_abc_15724_n907_1_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_1_), .Y(_abc_15724_n6184) );
  AND2X2 AND2X2_2676 ( .A(_abc_15724_n6186), .B(_abc_15724_n6187), .Y(_abc_15724_n6188) );
  AND2X2 AND2X2_2677 ( .A(_abc_15724_n6188), .B(digest_update_bF_buf0), .Y(_abc_15724_n6189) );
  AND2X2 AND2X2_2678 ( .A(_abc_15724_n907_1_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_2_), .Y(_abc_15724_n6190) );
  AND2X2 AND2X2_2679 ( .A(_abc_15724_n6192), .B(_abc_15724_n788), .Y(_abc_15724_n6193) );
  AND2X2 AND2X2_268 ( .A(_abc_15724_n1235), .B(_abc_15724_n1232), .Y(_abc_15724_n1236) );
  AND2X2 AND2X2_2680 ( .A(_abc_15724_n6197), .B(_abc_15724_n6194), .Y(_abc_15724_n6198) );
  AND2X2 AND2X2_2681 ( .A(_abc_15724_n6198), .B(digest_update_bF_buf11), .Y(_abc_15724_n6199) );
  AND2X2 AND2X2_2682 ( .A(_abc_15724_n907_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_3_), .Y(_abc_15724_n6200) );
  AND2X2 AND2X2_2683 ( .A(_abc_15724_n6202), .B(_abc_15724_n6203), .Y(_abc_15724_n6204) );
  AND2X2 AND2X2_2684 ( .A(_abc_15724_n6205), .B(_abc_15724_n6206), .Y(H4_reg_4__FF_INPUT) );
  AND2X2 AND2X2_2685 ( .A(_abc_15724_n6210), .B(_abc_15724_n785), .Y(_abc_15724_n6211) );
  AND2X2 AND2X2_2686 ( .A(_abc_15724_n6209), .B(_abc_15724_n6211), .Y(_abc_15724_n6212) );
  AND2X2 AND2X2_2687 ( .A(_abc_15724_n810), .B(_abc_15724_n6213), .Y(_abc_15724_n6214) );
  AND2X2 AND2X2_2688 ( .A(_abc_15724_n6216), .B(_abc_15724_n6208), .Y(H4_reg_5__FF_INPUT) );
  AND2X2 AND2X2_2689 ( .A(_abc_15724_n812_1), .B(_abc_15724_n782), .Y(_abc_15724_n6219) );
  AND2X2 AND2X2_269 ( .A(_abc_15724_n1219), .B(_abc_15724_n1207_1), .Y(_abc_15724_n1237_1) );
  AND2X2 AND2X2_2690 ( .A(_abc_15724_n6220), .B(_abc_15724_n6218), .Y(_abc_15724_n6221) );
  AND2X2 AND2X2_2691 ( .A(_abc_15724_n6221), .B(digest_update_bF_buf8), .Y(_abc_15724_n6222) );
  AND2X2 AND2X2_2692 ( .A(_abc_15724_n3031), .B(_abc_15724_n850_bF_buf2), .Y(_abc_15724_n6223) );
  AND2X2 AND2X2_2693 ( .A(_abc_15724_n6220), .B(_abc_15724_n780_1), .Y(_abc_15724_n6225) );
  AND2X2 AND2X2_2694 ( .A(_abc_15724_n6227), .B(_abc_15724_n6229), .Y(_abc_15724_n6230) );
  AND2X2 AND2X2_2695 ( .A(_abc_15724_n6230), .B(digest_update_bF_buf7), .Y(_abc_15724_n6231) );
  AND2X2 AND2X2_2696 ( .A(_abc_15724_n3037), .B(_abc_15724_n850_bF_buf1), .Y(_abc_15724_n6232) );
  AND2X2 AND2X2_2697 ( .A(_abc_15724_n814), .B(_abc_15724_n819), .Y(_abc_15724_n6235) );
  AND2X2 AND2X2_2698 ( .A(_abc_15724_n6236), .B(_abc_15724_n6234), .Y(_abc_15724_n6237) );
  AND2X2 AND2X2_2699 ( .A(_abc_15724_n6237), .B(digest_update_bF_buf6), .Y(_abc_15724_n6238) );
  AND2X2 AND2X2_27 ( .A(_abc_15724_n740), .B(_abc_15724_n738_1), .Y(_abc_15724_n750) );
  AND2X2 AND2X2_270 ( .A(_abc_15724_n1174), .B(_abc_15724_n1233), .Y(_abc_15724_n1241) );
  AND2X2 AND2X2_2700 ( .A(_abc_15724_n3043), .B(_abc_15724_n850_bF_buf0), .Y(_abc_15724_n6239) );
  AND2X2 AND2X2_2701 ( .A(_abc_15724_n6236), .B(_abc_15724_n817), .Y(_abc_15724_n6241) );
  AND2X2 AND2X2_2702 ( .A(_abc_15724_n6241), .B(_abc_15724_n816), .Y(_abc_15724_n6242) );
  AND2X2 AND2X2_2703 ( .A(_abc_15724_n6244), .B(_abc_15724_n6243), .Y(_abc_15724_n6245) );
  AND2X2 AND2X2_2704 ( .A(_abc_15724_n6246), .B(digest_update_bF_buf5), .Y(_abc_15724_n6247) );
  AND2X2 AND2X2_2705 ( .A(_abc_15724_n907_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_9_), .Y(_abc_15724_n6248) );
  AND2X2 AND2X2_2706 ( .A(_abc_15724_n907_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_10_), .Y(_abc_15724_n6250) );
  AND2X2 AND2X2_2707 ( .A(_abc_15724_n814), .B(_abc_15724_n820), .Y(_abc_15724_n6251) );
  AND2X2 AND2X2_2708 ( .A(_abc_15724_n6252), .B(_abc_15724_n764), .Y(_abc_15724_n6254) );
  AND2X2 AND2X2_2709 ( .A(_abc_15724_n6255), .B(_abc_15724_n6253), .Y(_abc_15724_n6256) );
  AND2X2 AND2X2_271 ( .A(_abc_15724_n1115), .B(_abc_15724_n1241), .Y(_abc_15724_n1242) );
  AND2X2 AND2X2_2710 ( .A(_abc_15724_n6256), .B(digest_update_bF_buf4), .Y(_abc_15724_n6257) );
  AND2X2 AND2X2_2711 ( .A(_abc_15724_n6255), .B(_abc_15724_n762), .Y(_abc_15724_n6259) );
  AND2X2 AND2X2_2712 ( .A(_abc_15724_n6259), .B(_abc_15724_n761), .Y(_abc_15724_n6260) );
  AND2X2 AND2X2_2713 ( .A(_abc_15724_n6262), .B(_abc_15724_n6261), .Y(_abc_15724_n6263) );
  AND2X2 AND2X2_2714 ( .A(_abc_15724_n6264), .B(digest_update_bF_buf3), .Y(_abc_15724_n6265) );
  AND2X2 AND2X2_2715 ( .A(_abc_15724_n907_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_11_), .Y(_abc_15724_n6266) );
  AND2X2 AND2X2_2716 ( .A(_abc_15724_n907_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_12_), .Y(_abc_15724_n6268) );
  AND2X2 AND2X2_2717 ( .A(_abc_15724_n823), .B(_abc_15724_n752), .Y(_abc_15724_n6270) );
  AND2X2 AND2X2_2718 ( .A(_abc_15724_n6271), .B(_abc_15724_n6269), .Y(_abc_15724_n6272) );
  AND2X2 AND2X2_2719 ( .A(_abc_15724_n6272), .B(digest_update_bF_buf2), .Y(_abc_15724_n6273) );
  AND2X2 AND2X2_272 ( .A(_auto_iopadmap_cc_313_execute_26059_48_), .B(d_reg_16_), .Y(_abc_15724_n1245) );
  AND2X2 AND2X2_2720 ( .A(_abc_15724_n6271), .B(_abc_15724_n742), .Y(_abc_15724_n6275) );
  AND2X2 AND2X2_2721 ( .A(_abc_15724_n6277), .B(_abc_15724_n6279), .Y(_abc_15724_n6280) );
  AND2X2 AND2X2_2722 ( .A(_abc_15724_n6280), .B(digest_update_bF_buf1), .Y(_abc_15724_n6281) );
  AND2X2 AND2X2_2723 ( .A(_abc_15724_n3073), .B(_abc_15724_n850_bF_buf8), .Y(_abc_15724_n6282) );
  AND2X2 AND2X2_2724 ( .A(_abc_15724_n823), .B(_abc_15724_n753), .Y(_abc_15724_n6284) );
  AND2X2 AND2X2_2725 ( .A(_abc_15724_n6285), .B(_abc_15724_n736), .Y(_abc_15724_n6287) );
  AND2X2 AND2X2_2726 ( .A(_abc_15724_n6288), .B(_abc_15724_n6286), .Y(_abc_15724_n6289) );
  AND2X2 AND2X2_2727 ( .A(_abc_15724_n6289), .B(digest_update_bF_buf0), .Y(_abc_15724_n6290) );
  AND2X2 AND2X2_2728 ( .A(_abc_15724_n3079_1), .B(_abc_15724_n850_bF_buf7), .Y(_abc_15724_n6291) );
  AND2X2 AND2X2_2729 ( .A(_abc_15724_n6288), .B(_abc_15724_n734), .Y(_abc_15724_n6293) );
  AND2X2 AND2X2_273 ( .A(_abc_15724_n1246), .B(_abc_15724_n1244), .Y(_abc_15724_n1247) );
  AND2X2 AND2X2_2730 ( .A(_abc_15724_n6293), .B(_abc_15724_n732), .Y(_abc_15724_n6294) );
  AND2X2 AND2X2_2731 ( .A(_abc_15724_n6296), .B(_abc_15724_n6295), .Y(_abc_15724_n6297) );
  AND2X2 AND2X2_2732 ( .A(_abc_15724_n6298), .B(digest_update_bF_buf11), .Y(_abc_15724_n6299) );
  AND2X2 AND2X2_2733 ( .A(_abc_15724_n3085), .B(_abc_15724_n850_bF_buf6), .Y(_abc_15724_n6300) );
  AND2X2 AND2X2_2734 ( .A(_abc_15724_n907_1_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_16_), .Y(_abc_15724_n6302) );
  AND2X2 AND2X2_2735 ( .A(_abc_15724_n825_1), .B(_abc_15724_n828), .Y(_abc_15724_n6304) );
  AND2X2 AND2X2_2736 ( .A(_abc_15724_n6305), .B(_abc_15724_n6303), .Y(_abc_15724_n6306) );
  AND2X2 AND2X2_2737 ( .A(_abc_15724_n6306), .B(digest_update_bF_buf10), .Y(_abc_15724_n6307) );
  AND2X2 AND2X2_2738 ( .A(_abc_15724_n6305), .B(_abc_15724_n717), .Y(_abc_15724_n6309) );
  AND2X2 AND2X2_2739 ( .A(_abc_15724_n6311), .B(_abc_15724_n6312), .Y(_abc_15724_n6313) );
  AND2X2 AND2X2_274 ( .A(_abc_15724_n1243), .B(_abc_15724_n1247), .Y(_abc_15724_n1249) );
  AND2X2 AND2X2_2740 ( .A(_abc_15724_n6313), .B(digest_update_bF_buf9), .Y(_abc_15724_n6314) );
  AND2X2 AND2X2_2741 ( .A(_abc_15724_n3097), .B(_abc_15724_n850_bF_buf5), .Y(_abc_15724_n6315) );
  AND2X2 AND2X2_2742 ( .A(_abc_15724_n907_1_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_18_), .Y(_abc_15724_n6317) );
  AND2X2 AND2X2_2743 ( .A(_abc_15724_n825_1), .B(_abc_15724_n829), .Y(_abc_15724_n6318) );
  AND2X2 AND2X2_2744 ( .A(_abc_15724_n6319), .B(_abc_15724_n712), .Y(_abc_15724_n6321) );
  AND2X2 AND2X2_2745 ( .A(_abc_15724_n6322), .B(_abc_15724_n6320), .Y(_abc_15724_n6323) );
  AND2X2 AND2X2_2746 ( .A(_abc_15724_n6323), .B(digest_update_bF_buf8), .Y(_abc_15724_n6324) );
  AND2X2 AND2X2_2747 ( .A(_abc_15724_n6322), .B(_abc_15724_n710_1), .Y(_abc_15724_n6327) );
  AND2X2 AND2X2_2748 ( .A(_abc_15724_n6328), .B(_abc_15724_n6326), .Y(_abc_15724_n6329) );
  AND2X2 AND2X2_2749 ( .A(_abc_15724_n6327), .B(_abc_15724_n708_1), .Y(_abc_15724_n6330) );
  AND2X2 AND2X2_275 ( .A(_abc_15724_n1250_1), .B(_abc_15724_n1248), .Y(_abc_15724_n1251_1) );
  AND2X2 AND2X2_2750 ( .A(_abc_15724_n6331), .B(digest_update_bF_buf7), .Y(_abc_15724_n6332) );
  AND2X2 AND2X2_2751 ( .A(_abc_15724_n907_1_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_19_), .Y(_abc_15724_n6333) );
  AND2X2 AND2X2_2752 ( .A(_abc_15724_n834_1), .B(_abc_15724_n837_1), .Y(_abc_15724_n6335) );
  AND2X2 AND2X2_2753 ( .A(_abc_15724_n6336), .B(_abc_15724_n6337), .Y(_abc_15724_n6338) );
  AND2X2 AND2X2_2754 ( .A(_abc_15724_n6338), .B(digest_update_bF_buf6), .Y(_abc_15724_n6339) );
  AND2X2 AND2X2_2755 ( .A(_abc_15724_n3115), .B(_abc_15724_n850_bF_buf4), .Y(_abc_15724_n6340) );
  AND2X2 AND2X2_2756 ( .A(_abc_15724_n6336), .B(_abc_15724_n835), .Y(_abc_15724_n6343) );
  AND2X2 AND2X2_2757 ( .A(_abc_15724_n6345), .B(_abc_15724_n6347), .Y(_abc_15724_n6348) );
  AND2X2 AND2X2_2758 ( .A(_abc_15724_n6349), .B(_abc_15724_n6342), .Y(H4_reg_21__FF_INPUT) );
  AND2X2 AND2X2_2759 ( .A(w_mem_inst__abc_21378_n1589), .B(w_mem_inst__abc_21378_n1591), .Y(w_mem_inst__abc_21378_n1592) );
  AND2X2 AND2X2_276 ( .A(_abc_15724_n1251_1), .B(digest_update_bF_buf8), .Y(_abc_15724_n1252) );
  AND2X2 AND2X2_2760 ( .A(w_mem_inst_w_mem_2__31_), .B(w_mem_inst_w_mem_0__31_), .Y(w_mem_inst__abc_21378_n1595) );
  AND2X2 AND2X2_2761 ( .A(w_mem_inst__abc_21378_n1596), .B(w_mem_inst__abc_21378_n1594_1), .Y(w_mem_inst__abc_21378_n1597) );
  AND2X2 AND2X2_2762 ( .A(w_mem_inst__abc_21378_n1598), .B(w_mem_inst__abc_21378_n1600), .Y(w_mem_inst__abc_21378_n1601_1) );
  AND2X2 AND2X2_2763 ( .A(w_mem_inst_w_ctr_reg_1_), .B(w_mem_inst_w_ctr_reg_0_), .Y(w_mem_inst__abc_21378_n1603_1) );
  AND2X2 AND2X2_2764 ( .A(w_mem_inst_w_ctr_reg_3_), .B(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_21378_n1604) );
  AND2X2 AND2X2_2765 ( .A(w_mem_inst__abc_21378_n1603_1), .B(w_mem_inst__abc_21378_n1604), .Y(w_mem_inst__abc_21378_n1605) );
  AND2X2 AND2X2_2766 ( .A(w_mem_inst__abc_21378_n1605_bF_buf4), .B(w_mem_inst_w_mem_15__0_), .Y(w_mem_inst__abc_21378_n1606_1) );
  AND2X2 AND2X2_2767 ( .A(w_mem_inst__abc_21378_n1607_1), .B(w_mem_inst__abc_21378_n1608), .Y(w_mem_inst__abc_21378_n1609) );
  AND2X2 AND2X2_2768 ( .A(w_mem_inst__abc_21378_n1609), .B(w_mem_inst__abc_21378_n1603_1), .Y(w_mem_inst__abc_21378_n1610_1) );
  AND2X2 AND2X2_2769 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf4), .B(w_mem_inst_w_mem_3__0_), .Y(w_mem_inst__abc_21378_n1611_1) );
  AND2X2 AND2X2_277 ( .A(_abc_15724_n1250_1), .B(_abc_15724_n1246), .Y(_abc_15724_n1254) );
  AND2X2 AND2X2_2770 ( .A(w_mem_inst__abc_21378_n1607_1), .B(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_21378_n1613) );
  AND2X2 AND2X2_2771 ( .A(w_mem_inst__abc_21378_n1614_1), .B(w_mem_inst_w_ctr_reg_0_), .Y(w_mem_inst__abc_21378_n1615_1) );
  AND2X2 AND2X2_2772 ( .A(w_mem_inst__abc_21378_n1613), .B(w_mem_inst__abc_21378_n1615_1), .Y(w_mem_inst__abc_21378_n1616) );
  AND2X2 AND2X2_2773 ( .A(w_mem_inst__abc_21378_n1616_bF_buf4), .B(w_mem_inst_w_mem_5__0_), .Y(w_mem_inst__abc_21378_n1617) );
  AND2X2 AND2X2_2774 ( .A(w_mem_inst__abc_21378_n1609), .B(w_mem_inst__abc_21378_n1615_1), .Y(w_mem_inst__abc_21378_n1618_1) );
  AND2X2 AND2X2_2775 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf4), .B(w_mem_inst_w_mem_1__0_), .Y(w_mem_inst__abc_21378_n1619_1) );
  AND2X2 AND2X2_2776 ( .A(w_mem_inst__abc_21378_n1623_1), .B(w_mem_inst_w_ctr_reg_1_), .Y(w_mem_inst__abc_21378_n1624) );
  AND2X2 AND2X2_2777 ( .A(w_mem_inst__abc_21378_n1609), .B(w_mem_inst__abc_21378_n1624), .Y(w_mem_inst__abc_21378_n1625) );
  AND2X2 AND2X2_2778 ( .A(w_mem_inst__abc_21378_n1625_bF_buf4), .B(w_mem_inst_w_mem_2__0_), .Y(w_mem_inst__abc_21378_n1626_1) );
  AND2X2 AND2X2_2779 ( .A(w_mem_inst__abc_21378_n1615_1), .B(w_mem_inst__abc_21378_n1604), .Y(w_mem_inst__abc_21378_n1627_1) );
  AND2X2 AND2X2_278 ( .A(_auto_iopadmap_cc_313_execute_26059_49_), .B(d_reg_17_), .Y(_abc_15724_n1257) );
  AND2X2 AND2X2_2780 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf4), .B(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_21378_n1628) );
  AND2X2 AND2X2_2781 ( .A(w_mem_inst__abc_21378_n1624), .B(w_mem_inst__abc_21378_n1604), .Y(w_mem_inst__abc_21378_n1630_1) );
  AND2X2 AND2X2_2782 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf4), .B(w_mem_inst_w_mem_14__0_), .Y(w_mem_inst__abc_21378_n1631_1) );
  AND2X2 AND2X2_2783 ( .A(w_mem_inst__abc_21378_n1614_1), .B(w_mem_inst__abc_21378_n1623_1), .Y(w_mem_inst__abc_21378_n1632) );
  AND2X2 AND2X2_2784 ( .A(w_mem_inst__abc_21378_n1608), .B(w_mem_inst_w_ctr_reg_3_), .Y(w_mem_inst__abc_21378_n1633) );
  AND2X2 AND2X2_2785 ( .A(w_mem_inst__abc_21378_n1632), .B(w_mem_inst__abc_21378_n1633), .Y(w_mem_inst__abc_21378_n1634_1) );
  AND2X2 AND2X2_2786 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf4), .B(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_21378_n1635_1) );
  AND2X2 AND2X2_2787 ( .A(w_mem_inst__abc_21378_n1613), .B(w_mem_inst__abc_21378_n1624), .Y(w_mem_inst__abc_21378_n1638_1) );
  AND2X2 AND2X2_2788 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf4), .B(w_mem_inst_w_mem_6__0_), .Y(w_mem_inst__abc_21378_n1639_1) );
  AND2X2 AND2X2_2789 ( .A(w_mem_inst__abc_21378_n1613), .B(w_mem_inst__abc_21378_n1603_1), .Y(w_mem_inst__abc_21378_n1640) );
  AND2X2 AND2X2_279 ( .A(_abc_15724_n1258), .B(_abc_15724_n1256), .Y(_abc_15724_n1259_1) );
  AND2X2 AND2X2_2790 ( .A(w_mem_inst__abc_21378_n1640_bF_buf4), .B(w_mem_inst_w_mem_7__0_), .Y(w_mem_inst__abc_21378_n1641) );
  AND2X2 AND2X2_2791 ( .A(w_mem_inst__abc_21378_n1609), .B(w_mem_inst__abc_21378_n1632), .Y(w_mem_inst__abc_21378_n1643_1) );
  AND2X2 AND2X2_2792 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf4), .B(w_mem_inst_w_mem_0__0_), .Y(w_mem_inst__abc_21378_n1644) );
  AND2X2 AND2X2_2793 ( .A(w_mem_inst__abc_21378_n1633), .B(w_mem_inst__abc_21378_n1603_1), .Y(w_mem_inst__abc_21378_n1645) );
  AND2X2 AND2X2_2794 ( .A(w_mem_inst__abc_21378_n1645_bF_buf4), .B(w_mem_inst_w_mem_11__0_), .Y(w_mem_inst__abc_21378_n1646_1) );
  AND2X2 AND2X2_2795 ( .A(w_mem_inst__abc_21378_n1615_1), .B(w_mem_inst__abc_21378_n1633), .Y(w_mem_inst__abc_21378_n1649) );
  AND2X2 AND2X2_2796 ( .A(w_mem_inst__abc_21378_n1649_bF_buf4), .B(w_mem_inst_w_mem_9__0_), .Y(w_mem_inst__abc_21378_n1650_1) );
  AND2X2 AND2X2_2797 ( .A(w_mem_inst__abc_21378_n1624), .B(w_mem_inst__abc_21378_n1633), .Y(w_mem_inst__abc_21378_n1651_1) );
  AND2X2 AND2X2_2798 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf4), .B(w_mem_inst_w_mem_10__0_), .Y(w_mem_inst__abc_21378_n1652) );
  AND2X2 AND2X2_2799 ( .A(w_mem_inst__abc_21378_n1632), .B(w_mem_inst__abc_21378_n1613), .Y(w_mem_inst__abc_21378_n1654_1) );
  AND2X2 AND2X2_28 ( .A(_abc_15724_n742), .B(_abc_15724_n751), .Y(_abc_15724_n752) );
  AND2X2 AND2X2_280 ( .A(_abc_15724_n1260_1), .B(_abc_15724_n1262), .Y(_abc_15724_n1263) );
  AND2X2 AND2X2_2800 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf4), .B(w_mem_inst_w_mem_4__0_), .Y(w_mem_inst__abc_21378_n1655_1) );
  AND2X2 AND2X2_2801 ( .A(w_mem_inst__abc_21378_n1632), .B(w_mem_inst__abc_21378_n1604), .Y(w_mem_inst__abc_21378_n1656) );
  AND2X2 AND2X2_2802 ( .A(w_mem_inst__abc_21378_n1656_bF_buf4), .B(w_mem_inst_w_mem_12__0_), .Y(w_mem_inst__abc_21378_n1657) );
  AND2X2 AND2X2_2803 ( .A(w_mem_inst__abc_21378_n1662_1), .B(w_mem_inst__abc_21378_n1602), .Y(w_0_) );
  AND2X2 AND2X2_2804 ( .A(w_mem_inst__abc_21378_n1665), .B(w_mem_inst__abc_21378_n1667_1), .Y(w_mem_inst__abc_21378_n1668) );
  AND2X2 AND2X2_2805 ( .A(w_mem_inst_w_mem_2__0_), .B(w_mem_inst_w_mem_0__0_), .Y(w_mem_inst__abc_21378_n1671_1) );
  AND2X2 AND2X2_2806 ( .A(w_mem_inst__abc_21378_n1672), .B(w_mem_inst__abc_21378_n1670_1), .Y(w_mem_inst__abc_21378_n1673) );
  AND2X2 AND2X2_2807 ( .A(w_mem_inst__abc_21378_n1674_1), .B(w_mem_inst__abc_21378_n1676), .Y(w_mem_inst__abc_21378_n1677) );
  AND2X2 AND2X2_2808 ( .A(w_mem_inst__abc_21378_n1605_bF_buf3), .B(w_mem_inst_w_mem_15__1_), .Y(w_mem_inst__abc_21378_n1679_1) );
  AND2X2 AND2X2_2809 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf3), .B(w_mem_inst_w_mem_3__1_), .Y(w_mem_inst__abc_21378_n1680) );
  AND2X2 AND2X2_281 ( .A(_abc_15724_n1263), .B(digest_update_bF_buf7), .Y(_abc_15724_n1264) );
  AND2X2 AND2X2_2810 ( .A(w_mem_inst__abc_21378_n1616_bF_buf3), .B(w_mem_inst_w_mem_5__1_), .Y(w_mem_inst__abc_21378_n1682_1) );
  AND2X2 AND2X2_2811 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf3), .B(w_mem_inst_w_mem_1__1_), .Y(w_mem_inst__abc_21378_n1683_1) );
  AND2X2 AND2X2_2812 ( .A(w_mem_inst__abc_21378_n1625_bF_buf3), .B(w_mem_inst_w_mem_2__1_), .Y(w_mem_inst__abc_21378_n1687_1) );
  AND2X2 AND2X2_2813 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf3), .B(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_21378_n1688) );
  AND2X2 AND2X2_2814 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf3), .B(w_mem_inst_w_mem_14__1_), .Y(w_mem_inst__abc_21378_n1690_1) );
  AND2X2 AND2X2_2815 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf3), .B(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_21378_n1691_1) );
  AND2X2 AND2X2_2816 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf3), .B(w_mem_inst_w_mem_6__1_), .Y(w_mem_inst__abc_21378_n1694_1) );
  AND2X2 AND2X2_2817 ( .A(w_mem_inst__abc_21378_n1640_bF_buf3), .B(w_mem_inst_w_mem_7__1_), .Y(w_mem_inst__abc_21378_n1695_1) );
  AND2X2 AND2X2_2818 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf3), .B(w_mem_inst_w_mem_0__1_), .Y(w_mem_inst__abc_21378_n1697) );
  AND2X2 AND2X2_2819 ( .A(w_mem_inst__abc_21378_n1645_bF_buf3), .B(w_mem_inst_w_mem_11__1_), .Y(w_mem_inst__abc_21378_n1698_1) );
  AND2X2 AND2X2_282 ( .A(_abc_15724_n1265), .B(_abc_15724_n850_bF_buf0), .Y(_abc_15724_n1266) );
  AND2X2 AND2X2_2820 ( .A(w_mem_inst__abc_21378_n1649_bF_buf3), .B(w_mem_inst_w_mem_9__1_), .Y(w_mem_inst__abc_21378_n1701) );
  AND2X2 AND2X2_2821 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf3), .B(w_mem_inst_w_mem_10__1_), .Y(w_mem_inst__abc_21378_n1702_1) );
  AND2X2 AND2X2_2822 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf3), .B(w_mem_inst_w_mem_4__1_), .Y(w_mem_inst__abc_21378_n1704) );
  AND2X2 AND2X2_2823 ( .A(w_mem_inst__abc_21378_n1656_bF_buf3), .B(w_mem_inst_w_mem_12__1_), .Y(w_mem_inst__abc_21378_n1705) );
  AND2X2 AND2X2_2824 ( .A(w_mem_inst__abc_21378_n1710_1), .B(w_mem_inst__abc_21378_n1678_1), .Y(w_1_) );
  AND2X2 AND2X2_2825 ( .A(w_mem_inst__abc_21378_n1713), .B(w_mem_inst__abc_21378_n1715_1), .Y(w_mem_inst__abc_21378_n1716) );
  AND2X2 AND2X2_2826 ( .A(w_mem_inst_w_mem_2__1_), .B(w_mem_inst_w_mem_0__1_), .Y(w_mem_inst__abc_21378_n1719_1) );
  AND2X2 AND2X2_2827 ( .A(w_mem_inst__abc_21378_n1720), .B(w_mem_inst__abc_21378_n1718_1), .Y(w_mem_inst__abc_21378_n1721) );
  AND2X2 AND2X2_2828 ( .A(w_mem_inst__abc_21378_n1722_1), .B(w_mem_inst__abc_21378_n1724), .Y(w_mem_inst__abc_21378_n1725) );
  AND2X2 AND2X2_2829 ( .A(w_mem_inst__abc_21378_n1605_bF_buf2), .B(w_mem_inst_w_mem_15__2_), .Y(w_mem_inst__abc_21378_n1727_1) );
  AND2X2 AND2X2_283 ( .A(_abc_15724_n907_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_50_), .Y(_abc_15724_n1268) );
  AND2X2 AND2X2_2830 ( .A(w_mem_inst__abc_21378_n1649_bF_buf2), .B(w_mem_inst_w_mem_9__2_), .Y(w_mem_inst__abc_21378_n1728) );
  AND2X2 AND2X2_2831 ( .A(w_mem_inst__abc_21378_n1616_bF_buf2), .B(w_mem_inst_w_mem_5__2_), .Y(w_mem_inst__abc_21378_n1730_1) );
  AND2X2 AND2X2_2832 ( .A(w_mem_inst__abc_21378_n1656_bF_buf2), .B(w_mem_inst_w_mem_12__2_), .Y(w_mem_inst__abc_21378_n1731_1) );
  AND2X2 AND2X2_2833 ( .A(w_mem_inst__abc_21378_n1625_bF_buf2), .B(w_mem_inst_w_mem_2__2_), .Y(w_mem_inst__abc_21378_n1735_1) );
  AND2X2 AND2X2_2834 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf2), .B(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_21378_n1736) );
  AND2X2 AND2X2_2835 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf2), .B(w_mem_inst_w_mem_14__2_), .Y(w_mem_inst__abc_21378_n1738_1) );
  AND2X2 AND2X2_2836 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf2), .B(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_21378_n1739_1) );
  AND2X2 AND2X2_2837 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf2), .B(w_mem_inst_w_mem_6__2_), .Y(w_mem_inst__abc_21378_n1742_1) );
  AND2X2 AND2X2_2838 ( .A(w_mem_inst__abc_21378_n1645_bF_buf2), .B(w_mem_inst_w_mem_11__2_), .Y(w_mem_inst__abc_21378_n1743_1) );
  AND2X2 AND2X2_2839 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf2), .B(w_mem_inst_w_mem_0__2_), .Y(w_mem_inst__abc_21378_n1745) );
  AND2X2 AND2X2_284 ( .A(_auto_iopadmap_cc_313_execute_26059_50_), .B(d_reg_18_), .Y(_abc_15724_n1270) );
  AND2X2 AND2X2_2840 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf2), .B(w_mem_inst_w_mem_4__2_), .Y(w_mem_inst__abc_21378_n1746_1) );
  AND2X2 AND2X2_2841 ( .A(w_mem_inst__abc_21378_n1640_bF_buf2), .B(w_mem_inst_w_mem_7__2_), .Y(w_mem_inst__abc_21378_n1749) );
  AND2X2 AND2X2_2842 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf2), .B(w_mem_inst_w_mem_3__2_), .Y(w_mem_inst__abc_21378_n1750_1) );
  AND2X2 AND2X2_2843 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf2), .B(w_mem_inst_w_mem_1__2_), .Y(w_mem_inst__abc_21378_n1752) );
  AND2X2 AND2X2_2844 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf2), .B(w_mem_inst_w_mem_10__2_), .Y(w_mem_inst__abc_21378_n1753) );
  AND2X2 AND2X2_2845 ( .A(w_mem_inst__abc_21378_n1758_1), .B(w_mem_inst__abc_21378_n1726_1), .Y(w_2_) );
  AND2X2 AND2X2_2846 ( .A(w_mem_inst__abc_21378_n1761), .B(w_mem_inst__abc_21378_n1763_1), .Y(w_mem_inst__abc_21378_n1764) );
  AND2X2 AND2X2_2847 ( .A(w_mem_inst_w_mem_2__2_), .B(w_mem_inst_w_mem_0__2_), .Y(w_mem_inst__abc_21378_n1767_1) );
  AND2X2 AND2X2_2848 ( .A(w_mem_inst__abc_21378_n1768), .B(w_mem_inst__abc_21378_n1766_1), .Y(w_mem_inst__abc_21378_n1769) );
  AND2X2 AND2X2_2849 ( .A(w_mem_inst__abc_21378_n1770_1), .B(w_mem_inst__abc_21378_n1772), .Y(w_mem_inst__abc_21378_n1773) );
  AND2X2 AND2X2_285 ( .A(_abc_15724_n1271), .B(_abc_15724_n1269), .Y(_abc_15724_n1272) );
  AND2X2 AND2X2_2850 ( .A(w_mem_inst__abc_21378_n1605_bF_buf1), .B(w_mem_inst_w_mem_15__3_), .Y(w_mem_inst__abc_21378_n1775_1) );
  AND2X2 AND2X2_2851 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf1), .B(w_mem_inst_w_mem_3__3_), .Y(w_mem_inst__abc_21378_n1776) );
  AND2X2 AND2X2_2852 ( .A(w_mem_inst__abc_21378_n1616_bF_buf1), .B(w_mem_inst_w_mem_5__3_), .Y(w_mem_inst__abc_21378_n1778_1) );
  AND2X2 AND2X2_2853 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf1), .B(w_mem_inst_w_mem_1__3_), .Y(w_mem_inst__abc_21378_n1779_1) );
  AND2X2 AND2X2_2854 ( .A(w_mem_inst__abc_21378_n1625_bF_buf1), .B(w_mem_inst_w_mem_2__3_), .Y(w_mem_inst__abc_21378_n1783_1) );
  AND2X2 AND2X2_2855 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf1), .B(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_21378_n1784) );
  AND2X2 AND2X2_2856 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf1), .B(w_mem_inst_w_mem_14__3_), .Y(w_mem_inst__abc_21378_n1786_1) );
  AND2X2 AND2X2_2857 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf1), .B(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_21378_n1787_1) );
  AND2X2 AND2X2_2858 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf1), .B(w_mem_inst_w_mem_6__3_), .Y(w_mem_inst__abc_21378_n1790_1) );
  AND2X2 AND2X2_2859 ( .A(w_mem_inst__abc_21378_n1640_bF_buf1), .B(w_mem_inst_w_mem_7__3_), .Y(w_mem_inst__abc_21378_n1791_1) );
  AND2X2 AND2X2_286 ( .A(_abc_15724_n1246), .B(_abc_15724_n1258), .Y(_abc_15724_n1274_1) );
  AND2X2 AND2X2_2860 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf1), .B(w_mem_inst_w_mem_0__3_), .Y(w_mem_inst__abc_21378_n1793) );
  AND2X2 AND2X2_2861 ( .A(w_mem_inst__abc_21378_n1645_bF_buf1), .B(w_mem_inst_w_mem_11__3_), .Y(w_mem_inst__abc_21378_n1794_1) );
  AND2X2 AND2X2_2862 ( .A(w_mem_inst__abc_21378_n1649_bF_buf1), .B(w_mem_inst_w_mem_9__3_), .Y(w_mem_inst__abc_21378_n1797) );
  AND2X2 AND2X2_2863 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf1), .B(w_mem_inst_w_mem_10__3_), .Y(w_mem_inst__abc_21378_n1798_1) );
  AND2X2 AND2X2_2864 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf1), .B(w_mem_inst_w_mem_4__3_), .Y(w_mem_inst__abc_21378_n1800) );
  AND2X2 AND2X2_2865 ( .A(w_mem_inst__abc_21378_n1656_bF_buf1), .B(w_mem_inst_w_mem_12__3_), .Y(w_mem_inst__abc_21378_n1801) );
  AND2X2 AND2X2_2866 ( .A(w_mem_inst__abc_21378_n1806_1), .B(w_mem_inst__abc_21378_n1774_1), .Y(w_3_) );
  AND2X2 AND2X2_2867 ( .A(w_mem_inst__abc_21378_n1809), .B(w_mem_inst__abc_21378_n1811_1), .Y(w_mem_inst__abc_21378_n1812) );
  AND2X2 AND2X2_2868 ( .A(w_mem_inst_w_mem_2__3_), .B(w_mem_inst_w_mem_0__3_), .Y(w_mem_inst__abc_21378_n1815_1) );
  AND2X2 AND2X2_2869 ( .A(w_mem_inst__abc_21378_n1816), .B(w_mem_inst__abc_21378_n1814_1), .Y(w_mem_inst__abc_21378_n1817) );
  AND2X2 AND2X2_287 ( .A(_abc_15724_n1250_1), .B(_abc_15724_n1274_1), .Y(_abc_15724_n1275_1) );
  AND2X2 AND2X2_2870 ( .A(w_mem_inst__abc_21378_n1818_1), .B(w_mem_inst__abc_21378_n1820), .Y(w_mem_inst__abc_21378_n1821) );
  AND2X2 AND2X2_2871 ( .A(w_mem_inst__abc_21378_n1605_bF_buf0), .B(w_mem_inst_w_mem_15__4_), .Y(w_mem_inst__abc_21378_n1823_1) );
  AND2X2 AND2X2_2872 ( .A(w_mem_inst__abc_21378_n1649_bF_buf0), .B(w_mem_inst_w_mem_9__4_), .Y(w_mem_inst__abc_21378_n1824) );
  AND2X2 AND2X2_2873 ( .A(w_mem_inst__abc_21378_n1616_bF_buf0), .B(w_mem_inst_w_mem_5__4_), .Y(w_mem_inst__abc_21378_n1826_1) );
  AND2X2 AND2X2_2874 ( .A(w_mem_inst__abc_21378_n1656_bF_buf0), .B(w_mem_inst_w_mem_12__4_), .Y(w_mem_inst__abc_21378_n1827_1) );
  AND2X2 AND2X2_2875 ( .A(w_mem_inst__abc_21378_n1625_bF_buf0), .B(w_mem_inst_w_mem_2__4_), .Y(w_mem_inst__abc_21378_n1831_1) );
  AND2X2 AND2X2_2876 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf0), .B(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_21378_n1832) );
  AND2X2 AND2X2_2877 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf0), .B(w_mem_inst_w_mem_14__4_), .Y(w_mem_inst__abc_21378_n1834_1) );
  AND2X2 AND2X2_2878 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf0), .B(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_21378_n1835_1) );
  AND2X2 AND2X2_2879 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf0), .B(w_mem_inst_w_mem_6__4_), .Y(w_mem_inst__abc_21378_n1838_1) );
  AND2X2 AND2X2_288 ( .A(_abc_15724_n1277), .B(_abc_15724_n1272), .Y(_abc_15724_n1279) );
  AND2X2 AND2X2_2880 ( .A(w_mem_inst__abc_21378_n1645_bF_buf0), .B(w_mem_inst_w_mem_11__4_), .Y(w_mem_inst__abc_21378_n1839_1) );
  AND2X2 AND2X2_2881 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf0), .B(w_mem_inst_w_mem_0__4_), .Y(w_mem_inst__abc_21378_n1841) );
  AND2X2 AND2X2_2882 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf0), .B(w_mem_inst_w_mem_4__4_), .Y(w_mem_inst__abc_21378_n1842_1) );
  AND2X2 AND2X2_2883 ( .A(w_mem_inst__abc_21378_n1640_bF_buf0), .B(w_mem_inst_w_mem_7__4_), .Y(w_mem_inst__abc_21378_n1845) );
  AND2X2 AND2X2_2884 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf0), .B(w_mem_inst_w_mem_3__4_), .Y(w_mem_inst__abc_21378_n1846_1) );
  AND2X2 AND2X2_2885 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf0), .B(w_mem_inst_w_mem_1__4_), .Y(w_mem_inst__abc_21378_n1848) );
  AND2X2 AND2X2_2886 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf0), .B(w_mem_inst_w_mem_10__4_), .Y(w_mem_inst__abc_21378_n1849) );
  AND2X2 AND2X2_2887 ( .A(w_mem_inst__abc_21378_n1854_1), .B(w_mem_inst__abc_21378_n1822_1), .Y(w_4_) );
  AND2X2 AND2X2_2888 ( .A(w_mem_inst__abc_21378_n1857), .B(w_mem_inst__abc_21378_n1859_1), .Y(w_mem_inst__abc_21378_n1860) );
  AND2X2 AND2X2_2889 ( .A(w_mem_inst_w_mem_2__4_), .B(w_mem_inst_w_mem_0__4_), .Y(w_mem_inst__abc_21378_n1863_1) );
  AND2X2 AND2X2_289 ( .A(_abc_15724_n1280), .B(_abc_15724_n1278), .Y(_abc_15724_n1281) );
  AND2X2 AND2X2_2890 ( .A(w_mem_inst__abc_21378_n1864), .B(w_mem_inst__abc_21378_n1862_1), .Y(w_mem_inst__abc_21378_n1865) );
  AND2X2 AND2X2_2891 ( .A(w_mem_inst__abc_21378_n1866_1), .B(w_mem_inst__abc_21378_n1868), .Y(w_mem_inst__abc_21378_n1869) );
  AND2X2 AND2X2_2892 ( .A(w_mem_inst__abc_21378_n1605_bF_buf4), .B(w_mem_inst_w_mem_15__5_), .Y(w_mem_inst__abc_21378_n1871_1) );
  AND2X2 AND2X2_2893 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf4), .B(w_mem_inst_w_mem_3__5_), .Y(w_mem_inst__abc_21378_n1872) );
  AND2X2 AND2X2_2894 ( .A(w_mem_inst__abc_21378_n1616_bF_buf4), .B(w_mem_inst_w_mem_5__5_), .Y(w_mem_inst__abc_21378_n1874_1) );
  AND2X2 AND2X2_2895 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf4), .B(w_mem_inst_w_mem_1__5_), .Y(w_mem_inst__abc_21378_n1875_1) );
  AND2X2 AND2X2_2896 ( .A(w_mem_inst__abc_21378_n1625_bF_buf4), .B(w_mem_inst_w_mem_2__5_), .Y(w_mem_inst__abc_21378_n1879_1) );
  AND2X2 AND2X2_2897 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf4), .B(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_21378_n1880) );
  AND2X2 AND2X2_2898 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf4), .B(w_mem_inst_w_mem_14__5_), .Y(w_mem_inst__abc_21378_n1882_1) );
  AND2X2 AND2X2_2899 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf4), .B(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_21378_n1883_1) );
  AND2X2 AND2X2_29 ( .A(_abc_15724_n750), .B(_abc_15724_n752), .Y(_abc_15724_n753) );
  AND2X2 AND2X2_290 ( .A(_abc_15724_n1281), .B(digest_update_bF_buf6), .Y(_abc_15724_n1282) );
  AND2X2 AND2X2_2900 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf4), .B(w_mem_inst_w_mem_6__5_), .Y(w_mem_inst__abc_21378_n1886_1) );
  AND2X2 AND2X2_2901 ( .A(w_mem_inst__abc_21378_n1640_bF_buf4), .B(w_mem_inst_w_mem_7__5_), .Y(w_mem_inst__abc_21378_n1887_1) );
  AND2X2 AND2X2_2902 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf4), .B(w_mem_inst_w_mem_0__5_), .Y(w_mem_inst__abc_21378_n1889) );
  AND2X2 AND2X2_2903 ( .A(w_mem_inst__abc_21378_n1645_bF_buf4), .B(w_mem_inst_w_mem_11__5_), .Y(w_mem_inst__abc_21378_n1890_1) );
  AND2X2 AND2X2_2904 ( .A(w_mem_inst__abc_21378_n1649_bF_buf4), .B(w_mem_inst_w_mem_9__5_), .Y(w_mem_inst__abc_21378_n1893) );
  AND2X2 AND2X2_2905 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf4), .B(w_mem_inst_w_mem_10__5_), .Y(w_mem_inst__abc_21378_n1894_1) );
  AND2X2 AND2X2_2906 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf4), .B(w_mem_inst_w_mem_4__5_), .Y(w_mem_inst__abc_21378_n1896) );
  AND2X2 AND2X2_2907 ( .A(w_mem_inst__abc_21378_n1656_bF_buf4), .B(w_mem_inst_w_mem_12__5_), .Y(w_mem_inst__abc_21378_n1897) );
  AND2X2 AND2X2_2908 ( .A(w_mem_inst__abc_21378_n1902_1), .B(w_mem_inst__abc_21378_n1870_1), .Y(w_5_) );
  AND2X2 AND2X2_2909 ( .A(w_mem_inst__abc_21378_n1905), .B(w_mem_inst__abc_21378_n1907_1), .Y(w_mem_inst__abc_21378_n1908) );
  AND2X2 AND2X2_291 ( .A(_abc_15724_n1280), .B(_abc_15724_n1271), .Y(_abc_15724_n1284_1) );
  AND2X2 AND2X2_2910 ( .A(w_mem_inst_w_mem_2__5_), .B(w_mem_inst_w_mem_0__5_), .Y(w_mem_inst__abc_21378_n1911_1) );
  AND2X2 AND2X2_2911 ( .A(w_mem_inst__abc_21378_n1912), .B(w_mem_inst__abc_21378_n1910_1), .Y(w_mem_inst__abc_21378_n1913) );
  AND2X2 AND2X2_2912 ( .A(w_mem_inst__abc_21378_n1914_1), .B(w_mem_inst__abc_21378_n1916), .Y(w_mem_inst__abc_21378_n1917) );
  AND2X2 AND2X2_2913 ( .A(w_mem_inst__abc_21378_n1605_bF_buf3), .B(w_mem_inst_w_mem_15__6_), .Y(w_mem_inst__abc_21378_n1919_1) );
  AND2X2 AND2X2_2914 ( .A(w_mem_inst__abc_21378_n1649_bF_buf3), .B(w_mem_inst_w_mem_9__6_), .Y(w_mem_inst__abc_21378_n1920) );
  AND2X2 AND2X2_2915 ( .A(w_mem_inst__abc_21378_n1616_bF_buf3), .B(w_mem_inst_w_mem_5__6_), .Y(w_mem_inst__abc_21378_n1922_1) );
  AND2X2 AND2X2_2916 ( .A(w_mem_inst__abc_21378_n1656_bF_buf3), .B(w_mem_inst_w_mem_12__6_), .Y(w_mem_inst__abc_21378_n1923_1) );
  AND2X2 AND2X2_2917 ( .A(w_mem_inst__abc_21378_n1625_bF_buf3), .B(w_mem_inst_w_mem_2__6_), .Y(w_mem_inst__abc_21378_n1927_1) );
  AND2X2 AND2X2_2918 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf3), .B(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_21378_n1928) );
  AND2X2 AND2X2_2919 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf3), .B(w_mem_inst_w_mem_14__6_), .Y(w_mem_inst__abc_21378_n1930_1) );
  AND2X2 AND2X2_292 ( .A(_auto_iopadmap_cc_313_execute_26059_51_), .B(d_reg_19_), .Y(_abc_15724_n1286) );
  AND2X2 AND2X2_2920 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf3), .B(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_21378_n1931_1) );
  AND2X2 AND2X2_2921 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf3), .B(w_mem_inst_w_mem_6__6_), .Y(w_mem_inst__abc_21378_n1934_1) );
  AND2X2 AND2X2_2922 ( .A(w_mem_inst__abc_21378_n1645_bF_buf3), .B(w_mem_inst_w_mem_11__6_), .Y(w_mem_inst__abc_21378_n1935_1) );
  AND2X2 AND2X2_2923 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf3), .B(w_mem_inst_w_mem_0__6_), .Y(w_mem_inst__abc_21378_n1937) );
  AND2X2 AND2X2_2924 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf3), .B(w_mem_inst_w_mem_4__6_), .Y(w_mem_inst__abc_21378_n1938_1) );
  AND2X2 AND2X2_2925 ( .A(w_mem_inst__abc_21378_n1640_bF_buf3), .B(w_mem_inst_w_mem_7__6_), .Y(w_mem_inst__abc_21378_n1941) );
  AND2X2 AND2X2_2926 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf3), .B(w_mem_inst_w_mem_3__6_), .Y(w_mem_inst__abc_21378_n1942_1) );
  AND2X2 AND2X2_2927 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf3), .B(w_mem_inst_w_mem_1__6_), .Y(w_mem_inst__abc_21378_n1944) );
  AND2X2 AND2X2_2928 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf3), .B(w_mem_inst_w_mem_10__6_), .Y(w_mem_inst__abc_21378_n1945) );
  AND2X2 AND2X2_2929 ( .A(w_mem_inst__abc_21378_n1950_1), .B(w_mem_inst__abc_21378_n1918_1), .Y(w_6_) );
  AND2X2 AND2X2_293 ( .A(_abc_15724_n1287_1), .B(_abc_15724_n1285_1), .Y(_abc_15724_n1288) );
  AND2X2 AND2X2_2930 ( .A(w_mem_inst__abc_21378_n1953), .B(w_mem_inst__abc_21378_n1955_1), .Y(w_mem_inst__abc_21378_n1956) );
  AND2X2 AND2X2_2931 ( .A(w_mem_inst_w_mem_2__6_), .B(w_mem_inst_w_mem_0__6_), .Y(w_mem_inst__abc_21378_n1959_1) );
  AND2X2 AND2X2_2932 ( .A(w_mem_inst__abc_21378_n1960), .B(w_mem_inst__abc_21378_n1958_1), .Y(w_mem_inst__abc_21378_n1961) );
  AND2X2 AND2X2_2933 ( .A(w_mem_inst__abc_21378_n1962_1), .B(w_mem_inst__abc_21378_n1964), .Y(w_mem_inst__abc_21378_n1965) );
  AND2X2 AND2X2_2934 ( .A(w_mem_inst__abc_21378_n1605_bF_buf2), .B(w_mem_inst_w_mem_15__7_), .Y(w_mem_inst__abc_21378_n1967_1) );
  AND2X2 AND2X2_2935 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf2), .B(w_mem_inst_w_mem_3__7_), .Y(w_mem_inst__abc_21378_n1968) );
  AND2X2 AND2X2_2936 ( .A(w_mem_inst__abc_21378_n1616_bF_buf2), .B(w_mem_inst_w_mem_5__7_), .Y(w_mem_inst__abc_21378_n1970_1) );
  AND2X2 AND2X2_2937 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf2), .B(w_mem_inst_w_mem_1__7_), .Y(w_mem_inst__abc_21378_n1971_1) );
  AND2X2 AND2X2_2938 ( .A(w_mem_inst__abc_21378_n1625_bF_buf2), .B(w_mem_inst_w_mem_2__7_), .Y(w_mem_inst__abc_21378_n1975_1) );
  AND2X2 AND2X2_2939 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf2), .B(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_21378_n1976) );
  AND2X2 AND2X2_294 ( .A(_abc_15724_n1284_1), .B(_abc_15724_n1288), .Y(_abc_15724_n1289) );
  AND2X2 AND2X2_2940 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf2), .B(w_mem_inst_w_mem_14__7_), .Y(w_mem_inst__abc_21378_n1978_1) );
  AND2X2 AND2X2_2941 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf2), .B(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_21378_n1979_1) );
  AND2X2 AND2X2_2942 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf2), .B(w_mem_inst_w_mem_6__7_), .Y(w_mem_inst__abc_21378_n1982_1) );
  AND2X2 AND2X2_2943 ( .A(w_mem_inst__abc_21378_n1640_bF_buf2), .B(w_mem_inst_w_mem_7__7_), .Y(w_mem_inst__abc_21378_n1983_1) );
  AND2X2 AND2X2_2944 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf2), .B(w_mem_inst_w_mem_0__7_), .Y(w_mem_inst__abc_21378_n1985) );
  AND2X2 AND2X2_2945 ( .A(w_mem_inst__abc_21378_n1645_bF_buf2), .B(w_mem_inst_w_mem_11__7_), .Y(w_mem_inst__abc_21378_n1986_1) );
  AND2X2 AND2X2_2946 ( .A(w_mem_inst__abc_21378_n1649_bF_buf2), .B(w_mem_inst_w_mem_9__7_), .Y(w_mem_inst__abc_21378_n1989) );
  AND2X2 AND2X2_2947 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf2), .B(w_mem_inst_w_mem_10__7_), .Y(w_mem_inst__abc_21378_n1990_1) );
  AND2X2 AND2X2_2948 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf2), .B(w_mem_inst_w_mem_4__7_), .Y(w_mem_inst__abc_21378_n1992) );
  AND2X2 AND2X2_2949 ( .A(w_mem_inst__abc_21378_n1656_bF_buf2), .B(w_mem_inst_w_mem_12__7_), .Y(w_mem_inst__abc_21378_n1993) );
  AND2X2 AND2X2_295 ( .A(_abc_15724_n1290), .B(_abc_15724_n1291), .Y(_abc_15724_n1292) );
  AND2X2 AND2X2_2950 ( .A(w_mem_inst__abc_21378_n1998_1), .B(w_mem_inst__abc_21378_n1966_1), .Y(w_7_) );
  AND2X2 AND2X2_2951 ( .A(w_mem_inst__abc_21378_n2001), .B(w_mem_inst__abc_21378_n2003_1), .Y(w_mem_inst__abc_21378_n2004) );
  AND2X2 AND2X2_2952 ( .A(w_mem_inst_w_mem_2__7_), .B(w_mem_inst_w_mem_0__7_), .Y(w_mem_inst__abc_21378_n2007_1) );
  AND2X2 AND2X2_2953 ( .A(w_mem_inst__abc_21378_n2008), .B(w_mem_inst__abc_21378_n2006_1), .Y(w_mem_inst__abc_21378_n2009) );
  AND2X2 AND2X2_2954 ( .A(w_mem_inst__abc_21378_n2010_1), .B(w_mem_inst__abc_21378_n2012), .Y(w_mem_inst__abc_21378_n2013) );
  AND2X2 AND2X2_2955 ( .A(w_mem_inst__abc_21378_n1605_bF_buf1), .B(w_mem_inst_w_mem_15__8_), .Y(w_mem_inst__abc_21378_n2015_1) );
  AND2X2 AND2X2_2956 ( .A(w_mem_inst__abc_21378_n1649_bF_buf1), .B(w_mem_inst_w_mem_9__8_), .Y(w_mem_inst__abc_21378_n2016) );
  AND2X2 AND2X2_2957 ( .A(w_mem_inst__abc_21378_n1616_bF_buf1), .B(w_mem_inst_w_mem_5__8_), .Y(w_mem_inst__abc_21378_n2018_1) );
  AND2X2 AND2X2_2958 ( .A(w_mem_inst__abc_21378_n1656_bF_buf1), .B(w_mem_inst_w_mem_12__8_), .Y(w_mem_inst__abc_21378_n2019_1) );
  AND2X2 AND2X2_2959 ( .A(w_mem_inst__abc_21378_n1625_bF_buf1), .B(w_mem_inst_w_mem_2__8_), .Y(w_mem_inst__abc_21378_n2023_1) );
  AND2X2 AND2X2_296 ( .A(_abc_15724_n1293), .B(digest_update_bF_buf5), .Y(_abc_15724_n1294) );
  AND2X2 AND2X2_2960 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf1), .B(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_21378_n2024) );
  AND2X2 AND2X2_2961 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf1), .B(w_mem_inst_w_mem_14__8_), .Y(w_mem_inst__abc_21378_n2026_1) );
  AND2X2 AND2X2_2962 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf1), .B(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_21378_n2027_1) );
  AND2X2 AND2X2_2963 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf1), .B(w_mem_inst_w_mem_6__8_), .Y(w_mem_inst__abc_21378_n2030_1) );
  AND2X2 AND2X2_2964 ( .A(w_mem_inst__abc_21378_n1645_bF_buf1), .B(w_mem_inst_w_mem_11__8_), .Y(w_mem_inst__abc_21378_n2031_1) );
  AND2X2 AND2X2_2965 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf1), .B(w_mem_inst_w_mem_0__8_), .Y(w_mem_inst__abc_21378_n2033) );
  AND2X2 AND2X2_2966 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf1), .B(w_mem_inst_w_mem_4__8_), .Y(w_mem_inst__abc_21378_n2034_1) );
  AND2X2 AND2X2_2967 ( .A(w_mem_inst__abc_21378_n1640_bF_buf1), .B(w_mem_inst_w_mem_7__8_), .Y(w_mem_inst__abc_21378_n2037) );
  AND2X2 AND2X2_2968 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf1), .B(w_mem_inst_w_mem_3__8_), .Y(w_mem_inst__abc_21378_n2038_1) );
  AND2X2 AND2X2_2969 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf1), .B(w_mem_inst_w_mem_1__8_), .Y(w_mem_inst__abc_21378_n2040) );
  AND2X2 AND2X2_297 ( .A(_abc_15724_n907_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_51_), .Y(_abc_15724_n1295) );
  AND2X2 AND2X2_2970 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf1), .B(w_mem_inst_w_mem_10__8_), .Y(w_mem_inst__abc_21378_n2041) );
  AND2X2 AND2X2_2971 ( .A(w_mem_inst__abc_21378_n2046_1), .B(w_mem_inst__abc_21378_n2014_1), .Y(w_8_) );
  AND2X2 AND2X2_2972 ( .A(w_mem_inst__abc_21378_n2049), .B(w_mem_inst__abc_21378_n2051_1), .Y(w_mem_inst__abc_21378_n2052) );
  AND2X2 AND2X2_2973 ( .A(w_mem_inst_w_mem_2__8_), .B(w_mem_inst_w_mem_0__8_), .Y(w_mem_inst__abc_21378_n2055_1) );
  AND2X2 AND2X2_2974 ( .A(w_mem_inst__abc_21378_n2056), .B(w_mem_inst__abc_21378_n2054_1), .Y(w_mem_inst__abc_21378_n2057) );
  AND2X2 AND2X2_2975 ( .A(w_mem_inst__abc_21378_n2058_1), .B(w_mem_inst__abc_21378_n2060), .Y(w_mem_inst__abc_21378_n2061) );
  AND2X2 AND2X2_2976 ( .A(w_mem_inst__abc_21378_n1605_bF_buf0), .B(w_mem_inst_w_mem_15__9_), .Y(w_mem_inst__abc_21378_n2063_1) );
  AND2X2 AND2X2_2977 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf0), .B(w_mem_inst_w_mem_3__9_), .Y(w_mem_inst__abc_21378_n2064) );
  AND2X2 AND2X2_2978 ( .A(w_mem_inst__abc_21378_n1616_bF_buf0), .B(w_mem_inst_w_mem_5__9_), .Y(w_mem_inst__abc_21378_n2066_1) );
  AND2X2 AND2X2_2979 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf0), .B(w_mem_inst_w_mem_1__9_), .Y(w_mem_inst__abc_21378_n2067_1) );
  AND2X2 AND2X2_298 ( .A(_abc_15724_n1272), .B(_abc_15724_n1288), .Y(_abc_15724_n1298) );
  AND2X2 AND2X2_2980 ( .A(w_mem_inst__abc_21378_n1625_bF_buf0), .B(w_mem_inst_w_mem_2__9_), .Y(w_mem_inst__abc_21378_n2071_1) );
  AND2X2 AND2X2_2981 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf0), .B(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_21378_n2072) );
  AND2X2 AND2X2_2982 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf0), .B(w_mem_inst_w_mem_14__9_), .Y(w_mem_inst__abc_21378_n2074_1) );
  AND2X2 AND2X2_2983 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf0), .B(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_21378_n2075_1) );
  AND2X2 AND2X2_2984 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf0), .B(w_mem_inst_w_mem_6__9_), .Y(w_mem_inst__abc_21378_n2078_1) );
  AND2X2 AND2X2_2985 ( .A(w_mem_inst__abc_21378_n1640_bF_buf0), .B(w_mem_inst_w_mem_7__9_), .Y(w_mem_inst__abc_21378_n2079_1) );
  AND2X2 AND2X2_2986 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf0), .B(w_mem_inst_w_mem_0__9_), .Y(w_mem_inst__abc_21378_n2081) );
  AND2X2 AND2X2_2987 ( .A(w_mem_inst__abc_21378_n1645_bF_buf0), .B(w_mem_inst_w_mem_11__9_), .Y(w_mem_inst__abc_21378_n2082_1) );
  AND2X2 AND2X2_2988 ( .A(w_mem_inst__abc_21378_n1649_bF_buf0), .B(w_mem_inst_w_mem_9__9_), .Y(w_mem_inst__abc_21378_n2085) );
  AND2X2 AND2X2_2989 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf0), .B(w_mem_inst_w_mem_10__9_), .Y(w_mem_inst__abc_21378_n2086_1) );
  AND2X2 AND2X2_299 ( .A(_abc_15724_n1285_1), .B(_abc_15724_n1270), .Y(_abc_15724_n1301) );
  AND2X2 AND2X2_2990 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf0), .B(w_mem_inst_w_mem_4__9_), .Y(w_mem_inst__abc_21378_n2088) );
  AND2X2 AND2X2_2991 ( .A(w_mem_inst__abc_21378_n1656_bF_buf0), .B(w_mem_inst_w_mem_12__9_), .Y(w_mem_inst__abc_21378_n2089) );
  AND2X2 AND2X2_2992 ( .A(w_mem_inst__abc_21378_n2094_1), .B(w_mem_inst__abc_21378_n2062_1), .Y(w_9_) );
  AND2X2 AND2X2_2993 ( .A(w_mem_inst__abc_21378_n2097), .B(w_mem_inst__abc_21378_n2099_1), .Y(w_mem_inst__abc_21378_n2100) );
  AND2X2 AND2X2_2994 ( .A(w_mem_inst_w_mem_2__9_), .B(w_mem_inst_w_mem_0__9_), .Y(w_mem_inst__abc_21378_n2103_1) );
  AND2X2 AND2X2_2995 ( .A(w_mem_inst__abc_21378_n2104), .B(w_mem_inst__abc_21378_n2102_1), .Y(w_mem_inst__abc_21378_n2105) );
  AND2X2 AND2X2_2996 ( .A(w_mem_inst__abc_21378_n2106_1), .B(w_mem_inst__abc_21378_n2108), .Y(w_mem_inst__abc_21378_n2109) );
  AND2X2 AND2X2_2997 ( .A(w_mem_inst__abc_21378_n1605_bF_buf4), .B(w_mem_inst_w_mem_15__10_), .Y(w_mem_inst__abc_21378_n2111_1) );
  AND2X2 AND2X2_2998 ( .A(w_mem_inst__abc_21378_n1649_bF_buf4), .B(w_mem_inst_w_mem_9__10_), .Y(w_mem_inst__abc_21378_n2112) );
  AND2X2 AND2X2_2999 ( .A(w_mem_inst__abc_21378_n1616_bF_buf4), .B(w_mem_inst_w_mem_5__10_), .Y(w_mem_inst__abc_21378_n2114_1) );
  AND2X2 AND2X2_3 ( .A(_abc_15724_n700), .B(_abc_15724_n701), .Y(_abc_15724_n702) );
  AND2X2 AND2X2_30 ( .A(_abc_15724_n737), .B(_abc_15724_n753), .Y(_abc_15724_n754) );
  AND2X2 AND2X2_300 ( .A(_abc_15724_n1300), .B(_abc_15724_n1303), .Y(_abc_15724_n1304) );
  AND2X2 AND2X2_3000 ( .A(w_mem_inst__abc_21378_n1656_bF_buf4), .B(w_mem_inst_w_mem_12__10_), .Y(w_mem_inst__abc_21378_n2115_1) );
  AND2X2 AND2X2_3001 ( .A(w_mem_inst__abc_21378_n1625_bF_buf4), .B(w_mem_inst_w_mem_2__10_), .Y(w_mem_inst__abc_21378_n2119_1) );
  AND2X2 AND2X2_3002 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf4), .B(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_21378_n2120) );
  AND2X2 AND2X2_3003 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf4), .B(w_mem_inst_w_mem_14__10_), .Y(w_mem_inst__abc_21378_n2122_1) );
  AND2X2 AND2X2_3004 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf4), .B(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_21378_n2123_1) );
  AND2X2 AND2X2_3005 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf4), .B(w_mem_inst_w_mem_6__10_), .Y(w_mem_inst__abc_21378_n2126_1) );
  AND2X2 AND2X2_3006 ( .A(w_mem_inst__abc_21378_n1645_bF_buf4), .B(w_mem_inst_w_mem_11__10_), .Y(w_mem_inst__abc_21378_n2127_1) );
  AND2X2 AND2X2_3007 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf4), .B(w_mem_inst_w_mem_0__10_), .Y(w_mem_inst__abc_21378_n2129) );
  AND2X2 AND2X2_3008 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf4), .B(w_mem_inst_w_mem_4__10_), .Y(w_mem_inst__abc_21378_n2130_1) );
  AND2X2 AND2X2_3009 ( .A(w_mem_inst__abc_21378_n1640_bF_buf4), .B(w_mem_inst_w_mem_7__10_), .Y(w_mem_inst__abc_21378_n2133) );
  AND2X2 AND2X2_301 ( .A(_abc_15724_n1247), .B(_abc_15724_n1259_1), .Y(_abc_15724_n1306_1) );
  AND2X2 AND2X2_3010 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf4), .B(w_mem_inst_w_mem_3__10_), .Y(w_mem_inst__abc_21378_n2134_1) );
  AND2X2 AND2X2_3011 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf4), .B(w_mem_inst_w_mem_1__10_), .Y(w_mem_inst__abc_21378_n2136) );
  AND2X2 AND2X2_3012 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf4), .B(w_mem_inst_w_mem_10__10_), .Y(w_mem_inst__abc_21378_n2137) );
  AND2X2 AND2X2_3013 ( .A(w_mem_inst__abc_21378_n2142_1), .B(w_mem_inst__abc_21378_n2110_1), .Y(w_10_) );
  AND2X2 AND2X2_3014 ( .A(w_mem_inst__abc_21378_n2145), .B(w_mem_inst__abc_21378_n2147_1), .Y(w_mem_inst__abc_21378_n2148) );
  AND2X2 AND2X2_3015 ( .A(w_mem_inst_w_mem_2__10_), .B(w_mem_inst_w_mem_0__10_), .Y(w_mem_inst__abc_21378_n2151_1) );
  AND2X2 AND2X2_3016 ( .A(w_mem_inst__abc_21378_n2152), .B(w_mem_inst__abc_21378_n2150_1), .Y(w_mem_inst__abc_21378_n2153) );
  AND2X2 AND2X2_3017 ( .A(w_mem_inst__abc_21378_n2154_1), .B(w_mem_inst__abc_21378_n2156), .Y(w_mem_inst__abc_21378_n2157) );
  AND2X2 AND2X2_3018 ( .A(w_mem_inst__abc_21378_n1605_bF_buf3), .B(w_mem_inst_w_mem_15__11_), .Y(w_mem_inst__abc_21378_n2159_1) );
  AND2X2 AND2X2_3019 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf3), .B(w_mem_inst_w_mem_3__11_), .Y(w_mem_inst__abc_21378_n2160) );
  AND2X2 AND2X2_302 ( .A(_abc_15724_n1306_1), .B(_abc_15724_n1298), .Y(_abc_15724_n1307) );
  AND2X2 AND2X2_3020 ( .A(w_mem_inst__abc_21378_n1616_bF_buf3), .B(w_mem_inst_w_mem_5__11_), .Y(w_mem_inst__abc_21378_n2162_1) );
  AND2X2 AND2X2_3021 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf3), .B(w_mem_inst_w_mem_1__11_), .Y(w_mem_inst__abc_21378_n2163_1) );
  AND2X2 AND2X2_3022 ( .A(w_mem_inst__abc_21378_n1625_bF_buf3), .B(w_mem_inst_w_mem_2__11_), .Y(w_mem_inst__abc_21378_n2167_1) );
  AND2X2 AND2X2_3023 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf3), .B(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_21378_n2168) );
  AND2X2 AND2X2_3024 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf3), .B(w_mem_inst_w_mem_14__11_), .Y(w_mem_inst__abc_21378_n2170_1) );
  AND2X2 AND2X2_3025 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf3), .B(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_21378_n2171_1) );
  AND2X2 AND2X2_3026 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf3), .B(w_mem_inst_w_mem_6__11_), .Y(w_mem_inst__abc_21378_n2174_1) );
  AND2X2 AND2X2_3027 ( .A(w_mem_inst__abc_21378_n1640_bF_buf3), .B(w_mem_inst_w_mem_7__11_), .Y(w_mem_inst__abc_21378_n2175_1) );
  AND2X2 AND2X2_3028 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf3), .B(w_mem_inst_w_mem_0__11_), .Y(w_mem_inst__abc_21378_n2177) );
  AND2X2 AND2X2_3029 ( .A(w_mem_inst__abc_21378_n1645_bF_buf3), .B(w_mem_inst_w_mem_11__11_), .Y(w_mem_inst__abc_21378_n2178_1) );
  AND2X2 AND2X2_303 ( .A(_abc_15724_n1243), .B(_abc_15724_n1307), .Y(_abc_15724_n1308_1) );
  AND2X2 AND2X2_3030 ( .A(w_mem_inst__abc_21378_n1649_bF_buf3), .B(w_mem_inst_w_mem_9__11_), .Y(w_mem_inst__abc_21378_n2181) );
  AND2X2 AND2X2_3031 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf3), .B(w_mem_inst_w_mem_10__11_), .Y(w_mem_inst__abc_21378_n2182_1) );
  AND2X2 AND2X2_3032 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf3), .B(w_mem_inst_w_mem_4__11_), .Y(w_mem_inst__abc_21378_n2184) );
  AND2X2 AND2X2_3033 ( .A(w_mem_inst__abc_21378_n1656_bF_buf3), .B(w_mem_inst_w_mem_12__11_), .Y(w_mem_inst__abc_21378_n2185) );
  AND2X2 AND2X2_3034 ( .A(w_mem_inst__abc_21378_n2190_1), .B(w_mem_inst__abc_21378_n2158_1), .Y(w_11_) );
  AND2X2 AND2X2_3035 ( .A(w_mem_inst__abc_21378_n2193), .B(w_mem_inst__abc_21378_n2195_1), .Y(w_mem_inst__abc_21378_n2196) );
  AND2X2 AND2X2_3036 ( .A(w_mem_inst_w_mem_2__11_), .B(w_mem_inst_w_mem_0__11_), .Y(w_mem_inst__abc_21378_n2199_1) );
  AND2X2 AND2X2_3037 ( .A(w_mem_inst__abc_21378_n2200), .B(w_mem_inst__abc_21378_n2198_1), .Y(w_mem_inst__abc_21378_n2201) );
  AND2X2 AND2X2_3038 ( .A(w_mem_inst__abc_21378_n2202_1), .B(w_mem_inst__abc_21378_n2204), .Y(w_mem_inst__abc_21378_n2205) );
  AND2X2 AND2X2_3039 ( .A(w_mem_inst__abc_21378_n1605_bF_buf2), .B(w_mem_inst_w_mem_15__12_), .Y(w_mem_inst__abc_21378_n2207_1) );
  AND2X2 AND2X2_304 ( .A(_auto_iopadmap_cc_313_execute_26059_52_), .B(d_reg_20_), .Y(_abc_15724_n1311) );
  AND2X2 AND2X2_3040 ( .A(w_mem_inst__abc_21378_n1649_bF_buf2), .B(w_mem_inst_w_mem_9__12_), .Y(w_mem_inst__abc_21378_n2208) );
  AND2X2 AND2X2_3041 ( .A(w_mem_inst__abc_21378_n1616_bF_buf2), .B(w_mem_inst_w_mem_5__12_), .Y(w_mem_inst__abc_21378_n2210_1) );
  AND2X2 AND2X2_3042 ( .A(w_mem_inst__abc_21378_n1656_bF_buf2), .B(w_mem_inst_w_mem_12__12_), .Y(w_mem_inst__abc_21378_n2211_1) );
  AND2X2 AND2X2_3043 ( .A(w_mem_inst__abc_21378_n1625_bF_buf2), .B(w_mem_inst_w_mem_2__12_), .Y(w_mem_inst__abc_21378_n2215_1) );
  AND2X2 AND2X2_3044 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf2), .B(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_21378_n2216) );
  AND2X2 AND2X2_3045 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf2), .B(w_mem_inst_w_mem_14__12_), .Y(w_mem_inst__abc_21378_n2218_1) );
  AND2X2 AND2X2_3046 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf2), .B(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_21378_n2219_1) );
  AND2X2 AND2X2_3047 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf2), .B(w_mem_inst_w_mem_6__12_), .Y(w_mem_inst__abc_21378_n2222_1) );
  AND2X2 AND2X2_3048 ( .A(w_mem_inst__abc_21378_n1645_bF_buf2), .B(w_mem_inst_w_mem_11__12_), .Y(w_mem_inst__abc_21378_n2223_1) );
  AND2X2 AND2X2_3049 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf2), .B(w_mem_inst_w_mem_0__12_), .Y(w_mem_inst__abc_21378_n2225) );
  AND2X2 AND2X2_305 ( .A(_abc_15724_n1312), .B(_abc_15724_n1310), .Y(_abc_15724_n1313) );
  AND2X2 AND2X2_3050 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf2), .B(w_mem_inst_w_mem_4__12_), .Y(w_mem_inst__abc_21378_n2226_1) );
  AND2X2 AND2X2_3051 ( .A(w_mem_inst__abc_21378_n1640_bF_buf2), .B(w_mem_inst_w_mem_7__12_), .Y(w_mem_inst__abc_21378_n2229) );
  AND2X2 AND2X2_3052 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf2), .B(w_mem_inst_w_mem_3__12_), .Y(w_mem_inst__abc_21378_n2230_1) );
  AND2X2 AND2X2_3053 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf2), .B(w_mem_inst_w_mem_1__12_), .Y(w_mem_inst__abc_21378_n2232) );
  AND2X2 AND2X2_3054 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf2), .B(w_mem_inst_w_mem_10__12_), .Y(w_mem_inst__abc_21378_n2233) );
  AND2X2 AND2X2_3055 ( .A(w_mem_inst__abc_21378_n2238_1), .B(w_mem_inst__abc_21378_n2206_1), .Y(w_12_) );
  AND2X2 AND2X2_3056 ( .A(w_mem_inst__abc_21378_n2241), .B(w_mem_inst__abc_21378_n2243_1), .Y(w_mem_inst__abc_21378_n2244) );
  AND2X2 AND2X2_3057 ( .A(w_mem_inst_w_mem_2__12_), .B(w_mem_inst_w_mem_0__12_), .Y(w_mem_inst__abc_21378_n2247_1) );
  AND2X2 AND2X2_3058 ( .A(w_mem_inst__abc_21378_n2248), .B(w_mem_inst__abc_21378_n2246_1), .Y(w_mem_inst__abc_21378_n2249) );
  AND2X2 AND2X2_3059 ( .A(w_mem_inst__abc_21378_n2250_1), .B(w_mem_inst__abc_21378_n2252), .Y(w_mem_inst__abc_21378_n2253) );
  AND2X2 AND2X2_306 ( .A(_abc_15724_n1309), .B(_abc_15724_n1313), .Y(_abc_15724_n1315) );
  AND2X2 AND2X2_3060 ( .A(w_mem_inst__abc_21378_n1605_bF_buf1), .B(w_mem_inst_w_mem_15__13_), .Y(w_mem_inst__abc_21378_n2255_1) );
  AND2X2 AND2X2_3061 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf1), .B(w_mem_inst_w_mem_3__13_), .Y(w_mem_inst__abc_21378_n2256) );
  AND2X2 AND2X2_3062 ( .A(w_mem_inst__abc_21378_n1616_bF_buf1), .B(w_mem_inst_w_mem_5__13_), .Y(w_mem_inst__abc_21378_n2258_1) );
  AND2X2 AND2X2_3063 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf1), .B(w_mem_inst_w_mem_1__13_), .Y(w_mem_inst__abc_21378_n2259_1) );
  AND2X2 AND2X2_3064 ( .A(w_mem_inst__abc_21378_n1625_bF_buf1), .B(w_mem_inst_w_mem_2__13_), .Y(w_mem_inst__abc_21378_n2263_1) );
  AND2X2 AND2X2_3065 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf1), .B(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_21378_n2264) );
  AND2X2 AND2X2_3066 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf1), .B(w_mem_inst_w_mem_14__13_), .Y(w_mem_inst__abc_21378_n2266_1) );
  AND2X2 AND2X2_3067 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf1), .B(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_21378_n2267_1) );
  AND2X2 AND2X2_3068 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf1), .B(w_mem_inst_w_mem_6__13_), .Y(w_mem_inst__abc_21378_n2270_1) );
  AND2X2 AND2X2_3069 ( .A(w_mem_inst__abc_21378_n1640_bF_buf1), .B(w_mem_inst_w_mem_7__13_), .Y(w_mem_inst__abc_21378_n2271_1) );
  AND2X2 AND2X2_307 ( .A(_abc_15724_n1316), .B(_abc_15724_n1314), .Y(_abc_15724_n1317) );
  AND2X2 AND2X2_3070 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf1), .B(w_mem_inst_w_mem_0__13_), .Y(w_mem_inst__abc_21378_n2273) );
  AND2X2 AND2X2_3071 ( .A(w_mem_inst__abc_21378_n1645_bF_buf1), .B(w_mem_inst_w_mem_11__13_), .Y(w_mem_inst__abc_21378_n2274_1) );
  AND2X2 AND2X2_3072 ( .A(w_mem_inst__abc_21378_n1649_bF_buf1), .B(w_mem_inst_w_mem_9__13_), .Y(w_mem_inst__abc_21378_n2277) );
  AND2X2 AND2X2_3073 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf1), .B(w_mem_inst_w_mem_10__13_), .Y(w_mem_inst__abc_21378_n2278_1) );
  AND2X2 AND2X2_3074 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf1), .B(w_mem_inst_w_mem_4__13_), .Y(w_mem_inst__abc_21378_n2280) );
  AND2X2 AND2X2_3075 ( .A(w_mem_inst__abc_21378_n1656_bF_buf1), .B(w_mem_inst_w_mem_12__13_), .Y(w_mem_inst__abc_21378_n2281) );
  AND2X2 AND2X2_3076 ( .A(w_mem_inst__abc_21378_n2286_1), .B(w_mem_inst__abc_21378_n2254_1), .Y(w_13_) );
  AND2X2 AND2X2_3077 ( .A(w_mem_inst__abc_21378_n2289), .B(w_mem_inst__abc_21378_n2291_1), .Y(w_mem_inst__abc_21378_n2292) );
  AND2X2 AND2X2_3078 ( .A(w_mem_inst_w_mem_2__13_), .B(w_mem_inst_w_mem_0__13_), .Y(w_mem_inst__abc_21378_n2295_1) );
  AND2X2 AND2X2_3079 ( .A(w_mem_inst__abc_21378_n2296), .B(w_mem_inst__abc_21378_n2294_1), .Y(w_mem_inst__abc_21378_n2297) );
  AND2X2 AND2X2_308 ( .A(_abc_15724_n1317), .B(digest_update_bF_buf4), .Y(_abc_15724_n1318) );
  AND2X2 AND2X2_3080 ( .A(w_mem_inst__abc_21378_n2298_1), .B(w_mem_inst__abc_21378_n2300), .Y(w_mem_inst__abc_21378_n2301) );
  AND2X2 AND2X2_3081 ( .A(w_mem_inst__abc_21378_n1605_bF_buf0), .B(w_mem_inst_w_mem_15__14_), .Y(w_mem_inst__abc_21378_n2303_1) );
  AND2X2 AND2X2_3082 ( .A(w_mem_inst__abc_21378_n1649_bF_buf0), .B(w_mem_inst_w_mem_9__14_), .Y(w_mem_inst__abc_21378_n2304) );
  AND2X2 AND2X2_3083 ( .A(w_mem_inst__abc_21378_n1616_bF_buf0), .B(w_mem_inst_w_mem_5__14_), .Y(w_mem_inst__abc_21378_n2306_1) );
  AND2X2 AND2X2_3084 ( .A(w_mem_inst__abc_21378_n1656_bF_buf0), .B(w_mem_inst_w_mem_12__14_), .Y(w_mem_inst__abc_21378_n2307_1) );
  AND2X2 AND2X2_3085 ( .A(w_mem_inst__abc_21378_n1625_bF_buf0), .B(w_mem_inst_w_mem_2__14_), .Y(w_mem_inst__abc_21378_n2311_1) );
  AND2X2 AND2X2_3086 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf0), .B(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_21378_n2312) );
  AND2X2 AND2X2_3087 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf0), .B(w_mem_inst_w_mem_14__14_), .Y(w_mem_inst__abc_21378_n2314_1) );
  AND2X2 AND2X2_3088 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf0), .B(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_21378_n2315_1) );
  AND2X2 AND2X2_3089 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf0), .B(w_mem_inst_w_mem_6__14_), .Y(w_mem_inst__abc_21378_n2318_1) );
  AND2X2 AND2X2_309 ( .A(_abc_15724_n1319_1), .B(_abc_15724_n850_bF_buf8), .Y(_abc_15724_n1320_1) );
  AND2X2 AND2X2_3090 ( .A(w_mem_inst__abc_21378_n1645_bF_buf0), .B(w_mem_inst_w_mem_11__14_), .Y(w_mem_inst__abc_21378_n2319_1) );
  AND2X2 AND2X2_3091 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf0), .B(w_mem_inst_w_mem_0__14_), .Y(w_mem_inst__abc_21378_n2321) );
  AND2X2 AND2X2_3092 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf0), .B(w_mem_inst_w_mem_4__14_), .Y(w_mem_inst__abc_21378_n2322_1) );
  AND2X2 AND2X2_3093 ( .A(w_mem_inst__abc_21378_n1640_bF_buf0), .B(w_mem_inst_w_mem_7__14_), .Y(w_mem_inst__abc_21378_n2325) );
  AND2X2 AND2X2_3094 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf0), .B(w_mem_inst_w_mem_3__14_), .Y(w_mem_inst__abc_21378_n2326_1) );
  AND2X2 AND2X2_3095 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf0), .B(w_mem_inst_w_mem_1__14_), .Y(w_mem_inst__abc_21378_n2328) );
  AND2X2 AND2X2_3096 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf0), .B(w_mem_inst_w_mem_10__14_), .Y(w_mem_inst__abc_21378_n2329) );
  AND2X2 AND2X2_3097 ( .A(w_mem_inst__abc_21378_n2334_1), .B(w_mem_inst__abc_21378_n2302_1), .Y(w_14_) );
  AND2X2 AND2X2_3098 ( .A(w_mem_inst__abc_21378_n2337), .B(w_mem_inst__abc_21378_n2339_1), .Y(w_mem_inst__abc_21378_n2340) );
  AND2X2 AND2X2_3099 ( .A(w_mem_inst_w_mem_2__14_), .B(w_mem_inst_w_mem_0__14_), .Y(w_mem_inst__abc_21378_n2343_1) );
  AND2X2 AND2X2_31 ( .A(e_reg_11_), .B(_auto_iopadmap_cc_313_execute_26059_11_), .Y(_abc_15724_n755) );
  AND2X2 AND2X2_310 ( .A(_abc_15724_n1316), .B(_abc_15724_n1312), .Y(_abc_15724_n1322) );
  AND2X2 AND2X2_3100 ( .A(w_mem_inst__abc_21378_n2344), .B(w_mem_inst__abc_21378_n2342_1), .Y(w_mem_inst__abc_21378_n2345) );
  AND2X2 AND2X2_3101 ( .A(w_mem_inst__abc_21378_n2346_1), .B(w_mem_inst__abc_21378_n2348), .Y(w_mem_inst__abc_21378_n2349) );
  AND2X2 AND2X2_3102 ( .A(w_mem_inst__abc_21378_n1605_bF_buf4), .B(w_mem_inst_w_mem_15__15_), .Y(w_mem_inst__abc_21378_n2351_1) );
  AND2X2 AND2X2_3103 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf4), .B(w_mem_inst_w_mem_3__15_), .Y(w_mem_inst__abc_21378_n2352) );
  AND2X2 AND2X2_3104 ( .A(w_mem_inst__abc_21378_n1616_bF_buf4), .B(w_mem_inst_w_mem_5__15_), .Y(w_mem_inst__abc_21378_n2354_1) );
  AND2X2 AND2X2_3105 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf4), .B(w_mem_inst_w_mem_1__15_), .Y(w_mem_inst__abc_21378_n2355_1) );
  AND2X2 AND2X2_3106 ( .A(w_mem_inst__abc_21378_n1625_bF_buf4), .B(w_mem_inst_w_mem_2__15_), .Y(w_mem_inst__abc_21378_n2359_1) );
  AND2X2 AND2X2_3107 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf4), .B(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_21378_n2360) );
  AND2X2 AND2X2_3108 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf4), .B(w_mem_inst_w_mem_14__15_), .Y(w_mem_inst__abc_21378_n2362_1) );
  AND2X2 AND2X2_3109 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf4), .B(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_21378_n2363_1) );
  AND2X2 AND2X2_311 ( .A(_auto_iopadmap_cc_313_execute_26059_53_), .B(d_reg_21_), .Y(_abc_15724_n1324) );
  AND2X2 AND2X2_3110 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf4), .B(w_mem_inst_w_mem_6__15_), .Y(w_mem_inst__abc_21378_n2366_1) );
  AND2X2 AND2X2_3111 ( .A(w_mem_inst__abc_21378_n1640_bF_buf4), .B(w_mem_inst_w_mem_7__15_), .Y(w_mem_inst__abc_21378_n2367_1) );
  AND2X2 AND2X2_3112 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf4), .B(w_mem_inst_w_mem_0__15_), .Y(w_mem_inst__abc_21378_n2369) );
  AND2X2 AND2X2_3113 ( .A(w_mem_inst__abc_21378_n1645_bF_buf4), .B(w_mem_inst_w_mem_11__15_), .Y(w_mem_inst__abc_21378_n2370_1) );
  AND2X2 AND2X2_3114 ( .A(w_mem_inst__abc_21378_n1649_bF_buf4), .B(w_mem_inst_w_mem_9__15_), .Y(w_mem_inst__abc_21378_n2373) );
  AND2X2 AND2X2_3115 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf4), .B(w_mem_inst_w_mem_10__15_), .Y(w_mem_inst__abc_21378_n2374_1) );
  AND2X2 AND2X2_3116 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf4), .B(w_mem_inst_w_mem_4__15_), .Y(w_mem_inst__abc_21378_n2376) );
  AND2X2 AND2X2_3117 ( .A(w_mem_inst__abc_21378_n1656_bF_buf4), .B(w_mem_inst_w_mem_12__15_), .Y(w_mem_inst__abc_21378_n2377) );
  AND2X2 AND2X2_3118 ( .A(w_mem_inst__abc_21378_n2382_1), .B(w_mem_inst__abc_21378_n2350_1), .Y(w_15_) );
  AND2X2 AND2X2_3119 ( .A(w_mem_inst__abc_21378_n2385), .B(w_mem_inst__abc_21378_n2387_1), .Y(w_mem_inst__abc_21378_n2388) );
  AND2X2 AND2X2_312 ( .A(_abc_15724_n1325), .B(_abc_15724_n1323), .Y(_abc_15724_n1326) );
  AND2X2 AND2X2_3120 ( .A(w_mem_inst_w_mem_2__15_), .B(w_mem_inst_w_mem_0__15_), .Y(w_mem_inst__abc_21378_n2391_1) );
  AND2X2 AND2X2_3121 ( .A(w_mem_inst__abc_21378_n2392), .B(w_mem_inst__abc_21378_n2390_1), .Y(w_mem_inst__abc_21378_n2393) );
  AND2X2 AND2X2_3122 ( .A(w_mem_inst__abc_21378_n2394_1), .B(w_mem_inst__abc_21378_n2396), .Y(w_mem_inst__abc_21378_n2397) );
  AND2X2 AND2X2_3123 ( .A(w_mem_inst__abc_21378_n1605_bF_buf3), .B(w_mem_inst_w_mem_15__16_), .Y(w_mem_inst__abc_21378_n2399_1) );
  AND2X2 AND2X2_3124 ( .A(w_mem_inst__abc_21378_n1649_bF_buf3), .B(w_mem_inst_w_mem_9__16_), .Y(w_mem_inst__abc_21378_n2400) );
  AND2X2 AND2X2_3125 ( .A(w_mem_inst__abc_21378_n1616_bF_buf3), .B(w_mem_inst_w_mem_5__16_), .Y(w_mem_inst__abc_21378_n2402_1) );
  AND2X2 AND2X2_3126 ( .A(w_mem_inst__abc_21378_n1656_bF_buf3), .B(w_mem_inst_w_mem_12__16_), .Y(w_mem_inst__abc_21378_n2403_1) );
  AND2X2 AND2X2_3127 ( .A(w_mem_inst__abc_21378_n1625_bF_buf3), .B(w_mem_inst_w_mem_2__16_), .Y(w_mem_inst__abc_21378_n2407_1) );
  AND2X2 AND2X2_3128 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf3), .B(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_21378_n2408) );
  AND2X2 AND2X2_3129 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf3), .B(w_mem_inst_w_mem_14__16_), .Y(w_mem_inst__abc_21378_n2410_1) );
  AND2X2 AND2X2_313 ( .A(_abc_15724_n1322), .B(_abc_15724_n1326), .Y(_abc_15724_n1327) );
  AND2X2 AND2X2_3130 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf3), .B(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_21378_n2411_1) );
  AND2X2 AND2X2_3131 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf3), .B(w_mem_inst_w_mem_6__16_), .Y(w_mem_inst__abc_21378_n2414_1) );
  AND2X2 AND2X2_3132 ( .A(w_mem_inst__abc_21378_n1645_bF_buf3), .B(w_mem_inst_w_mem_11__16_), .Y(w_mem_inst__abc_21378_n2415_1) );
  AND2X2 AND2X2_3133 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf3), .B(w_mem_inst_w_mem_0__16_), .Y(w_mem_inst__abc_21378_n2417) );
  AND2X2 AND2X2_3134 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf3), .B(w_mem_inst_w_mem_4__16_), .Y(w_mem_inst__abc_21378_n2418_1) );
  AND2X2 AND2X2_3135 ( .A(w_mem_inst__abc_21378_n1640_bF_buf3), .B(w_mem_inst_w_mem_7__16_), .Y(w_mem_inst__abc_21378_n2421) );
  AND2X2 AND2X2_3136 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf3), .B(w_mem_inst_w_mem_3__16_), .Y(w_mem_inst__abc_21378_n2422_1) );
  AND2X2 AND2X2_3137 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf3), .B(w_mem_inst_w_mem_1__16_), .Y(w_mem_inst__abc_21378_n2424) );
  AND2X2 AND2X2_3138 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf3), .B(w_mem_inst_w_mem_10__16_), .Y(w_mem_inst__abc_21378_n2425) );
  AND2X2 AND2X2_3139 ( .A(w_mem_inst__abc_21378_n2430_1), .B(w_mem_inst__abc_21378_n2398_1), .Y(w_16_) );
  AND2X2 AND2X2_314 ( .A(_abc_15724_n1328), .B(_abc_15724_n1329_1), .Y(_abc_15724_n1330_1) );
  AND2X2 AND2X2_3140 ( .A(w_mem_inst__abc_21378_n2433), .B(w_mem_inst__abc_21378_n2435_1), .Y(w_mem_inst__abc_21378_n2436) );
  AND2X2 AND2X2_3141 ( .A(w_mem_inst_w_mem_2__16_), .B(w_mem_inst_w_mem_0__16_), .Y(w_mem_inst__abc_21378_n2439_1) );
  AND2X2 AND2X2_3142 ( .A(w_mem_inst__abc_21378_n2440), .B(w_mem_inst__abc_21378_n2438_1), .Y(w_mem_inst__abc_21378_n2441) );
  AND2X2 AND2X2_3143 ( .A(w_mem_inst__abc_21378_n2442_1), .B(w_mem_inst__abc_21378_n2444), .Y(w_mem_inst__abc_21378_n2445) );
  AND2X2 AND2X2_3144 ( .A(w_mem_inst__abc_21378_n1605_bF_buf2), .B(w_mem_inst_w_mem_15__17_), .Y(w_mem_inst__abc_21378_n2447_1) );
  AND2X2 AND2X2_3145 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf2), .B(w_mem_inst_w_mem_3__17_), .Y(w_mem_inst__abc_21378_n2448) );
  AND2X2 AND2X2_3146 ( .A(w_mem_inst__abc_21378_n1616_bF_buf2), .B(w_mem_inst_w_mem_5__17_), .Y(w_mem_inst__abc_21378_n2450_1) );
  AND2X2 AND2X2_3147 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf2), .B(w_mem_inst_w_mem_1__17_), .Y(w_mem_inst__abc_21378_n2451_1) );
  AND2X2 AND2X2_3148 ( .A(w_mem_inst__abc_21378_n1625_bF_buf2), .B(w_mem_inst_w_mem_2__17_), .Y(w_mem_inst__abc_21378_n2455_1) );
  AND2X2 AND2X2_3149 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf2), .B(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_21378_n2456) );
  AND2X2 AND2X2_315 ( .A(_abc_15724_n1331), .B(digest_update_bF_buf3), .Y(_abc_15724_n1332_1) );
  AND2X2 AND2X2_3150 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf2), .B(w_mem_inst_w_mem_14__17_), .Y(w_mem_inst__abc_21378_n2458_1) );
  AND2X2 AND2X2_3151 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf2), .B(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_21378_n2459_1) );
  AND2X2 AND2X2_3152 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf2), .B(w_mem_inst_w_mem_6__17_), .Y(w_mem_inst__abc_21378_n2462_1) );
  AND2X2 AND2X2_3153 ( .A(w_mem_inst__abc_21378_n1640_bF_buf2), .B(w_mem_inst_w_mem_7__17_), .Y(w_mem_inst__abc_21378_n2463_1) );
  AND2X2 AND2X2_3154 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf2), .B(w_mem_inst_w_mem_0__17_), .Y(w_mem_inst__abc_21378_n2465) );
  AND2X2 AND2X2_3155 ( .A(w_mem_inst__abc_21378_n1645_bF_buf2), .B(w_mem_inst_w_mem_11__17_), .Y(w_mem_inst__abc_21378_n2466_1) );
  AND2X2 AND2X2_3156 ( .A(w_mem_inst__abc_21378_n1649_bF_buf2), .B(w_mem_inst_w_mem_9__17_), .Y(w_mem_inst__abc_21378_n2469) );
  AND2X2 AND2X2_3157 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf2), .B(w_mem_inst_w_mem_10__17_), .Y(w_mem_inst__abc_21378_n2470_1) );
  AND2X2 AND2X2_3158 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf2), .B(w_mem_inst_w_mem_4__17_), .Y(w_mem_inst__abc_21378_n2472) );
  AND2X2 AND2X2_3159 ( .A(w_mem_inst__abc_21378_n1656_bF_buf2), .B(w_mem_inst_w_mem_12__17_), .Y(w_mem_inst__abc_21378_n2473) );
  AND2X2 AND2X2_316 ( .A(_abc_15724_n1333), .B(_abc_15724_n850_bF_buf7), .Y(_abc_15724_n1334) );
  AND2X2 AND2X2_3160 ( .A(w_mem_inst__abc_21378_n2478_1), .B(w_mem_inst__abc_21378_n2446_1), .Y(w_17_) );
  AND2X2 AND2X2_3161 ( .A(w_mem_inst__abc_21378_n2481), .B(w_mem_inst__abc_21378_n2483_1), .Y(w_mem_inst__abc_21378_n2484) );
  AND2X2 AND2X2_3162 ( .A(w_mem_inst_w_mem_2__17_), .B(w_mem_inst_w_mem_0__17_), .Y(w_mem_inst__abc_21378_n2487_1) );
  AND2X2 AND2X2_3163 ( .A(w_mem_inst__abc_21378_n2488), .B(w_mem_inst__abc_21378_n2486_1), .Y(w_mem_inst__abc_21378_n2489) );
  AND2X2 AND2X2_3164 ( .A(w_mem_inst__abc_21378_n2490_1), .B(w_mem_inst__abc_21378_n2492), .Y(w_mem_inst__abc_21378_n2493) );
  AND2X2 AND2X2_3165 ( .A(w_mem_inst__abc_21378_n1605_bF_buf1), .B(w_mem_inst_w_mem_15__18_), .Y(w_mem_inst__abc_21378_n2495_1) );
  AND2X2 AND2X2_3166 ( .A(w_mem_inst__abc_21378_n1649_bF_buf1), .B(w_mem_inst_w_mem_9__18_), .Y(w_mem_inst__abc_21378_n2496) );
  AND2X2 AND2X2_3167 ( .A(w_mem_inst__abc_21378_n1616_bF_buf1), .B(w_mem_inst_w_mem_5__18_), .Y(w_mem_inst__abc_21378_n2498_1) );
  AND2X2 AND2X2_3168 ( .A(w_mem_inst__abc_21378_n1656_bF_buf1), .B(w_mem_inst_w_mem_12__18_), .Y(w_mem_inst__abc_21378_n2499_1) );
  AND2X2 AND2X2_3169 ( .A(w_mem_inst__abc_21378_n1625_bF_buf1), .B(w_mem_inst_w_mem_2__18_), .Y(w_mem_inst__abc_21378_n2503_1) );
  AND2X2 AND2X2_317 ( .A(_abc_15724_n907_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_54_), .Y(_abc_15724_n1336) );
  AND2X2 AND2X2_3170 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf1), .B(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_21378_n2504) );
  AND2X2 AND2X2_3171 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf1), .B(w_mem_inst_w_mem_14__18_), .Y(w_mem_inst__abc_21378_n2506_1) );
  AND2X2 AND2X2_3172 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf1), .B(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_21378_n2507_1) );
  AND2X2 AND2X2_3173 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf1), .B(w_mem_inst_w_mem_6__18_), .Y(w_mem_inst__abc_21378_n2510_1) );
  AND2X2 AND2X2_3174 ( .A(w_mem_inst__abc_21378_n1645_bF_buf1), .B(w_mem_inst_w_mem_11__18_), .Y(w_mem_inst__abc_21378_n2511_1) );
  AND2X2 AND2X2_3175 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf1), .B(w_mem_inst_w_mem_0__18_), .Y(w_mem_inst__abc_21378_n2513) );
  AND2X2 AND2X2_3176 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf1), .B(w_mem_inst_w_mem_4__18_), .Y(w_mem_inst__abc_21378_n2514_1) );
  AND2X2 AND2X2_3177 ( .A(w_mem_inst__abc_21378_n1640_bF_buf1), .B(w_mem_inst_w_mem_7__18_), .Y(w_mem_inst__abc_21378_n2517) );
  AND2X2 AND2X2_3178 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf1), .B(w_mem_inst_w_mem_3__18_), .Y(w_mem_inst__abc_21378_n2518_1) );
  AND2X2 AND2X2_3179 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf1), .B(w_mem_inst_w_mem_1__18_), .Y(w_mem_inst__abc_21378_n2520) );
  AND2X2 AND2X2_318 ( .A(_auto_iopadmap_cc_313_execute_26059_54_), .B(d_reg_22_), .Y(_abc_15724_n1338) );
  AND2X2 AND2X2_3180 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf1), .B(w_mem_inst_w_mem_10__18_), .Y(w_mem_inst__abc_21378_n2521) );
  AND2X2 AND2X2_3181 ( .A(w_mem_inst__abc_21378_n2526_1), .B(w_mem_inst__abc_21378_n2494_1), .Y(w_18_) );
  AND2X2 AND2X2_3182 ( .A(w_mem_inst__abc_21378_n2529), .B(w_mem_inst__abc_21378_n2531_1), .Y(w_mem_inst__abc_21378_n2532) );
  AND2X2 AND2X2_3183 ( .A(w_mem_inst_w_mem_2__18_), .B(w_mem_inst_w_mem_0__18_), .Y(w_mem_inst__abc_21378_n2535_1) );
  AND2X2 AND2X2_3184 ( .A(w_mem_inst__abc_21378_n2536), .B(w_mem_inst__abc_21378_n2534_1), .Y(w_mem_inst__abc_21378_n2537) );
  AND2X2 AND2X2_3185 ( .A(w_mem_inst__abc_21378_n2538_1), .B(w_mem_inst__abc_21378_n2540), .Y(w_mem_inst__abc_21378_n2541) );
  AND2X2 AND2X2_3186 ( .A(w_mem_inst__abc_21378_n1605_bF_buf0), .B(w_mem_inst_w_mem_15__19_), .Y(w_mem_inst__abc_21378_n2543_1) );
  AND2X2 AND2X2_3187 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf0), .B(w_mem_inst_w_mem_3__19_), .Y(w_mem_inst__abc_21378_n2544) );
  AND2X2 AND2X2_3188 ( .A(w_mem_inst__abc_21378_n1616_bF_buf0), .B(w_mem_inst_w_mem_5__19_), .Y(w_mem_inst__abc_21378_n2546_1) );
  AND2X2 AND2X2_3189 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf0), .B(w_mem_inst_w_mem_1__19_), .Y(w_mem_inst__abc_21378_n2547_1) );
  AND2X2 AND2X2_319 ( .A(_abc_15724_n1339), .B(_abc_15724_n1337), .Y(_abc_15724_n1340_1) );
  AND2X2 AND2X2_3190 ( .A(w_mem_inst__abc_21378_n1625_bF_buf0), .B(w_mem_inst_w_mem_2__19_), .Y(w_mem_inst__abc_21378_n2551_1) );
  AND2X2 AND2X2_3191 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf0), .B(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_21378_n2552) );
  AND2X2 AND2X2_3192 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf0), .B(w_mem_inst_w_mem_14__19_), .Y(w_mem_inst__abc_21378_n2554_1) );
  AND2X2 AND2X2_3193 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf0), .B(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_21378_n2555_1) );
  AND2X2 AND2X2_3194 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf0), .B(w_mem_inst_w_mem_6__19_), .Y(w_mem_inst__abc_21378_n2558_1) );
  AND2X2 AND2X2_3195 ( .A(w_mem_inst__abc_21378_n1640_bF_buf0), .B(w_mem_inst_w_mem_7__19_), .Y(w_mem_inst__abc_21378_n2559_1) );
  AND2X2 AND2X2_3196 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf0), .B(w_mem_inst_w_mem_0__19_), .Y(w_mem_inst__abc_21378_n2561) );
  AND2X2 AND2X2_3197 ( .A(w_mem_inst__abc_21378_n1645_bF_buf0), .B(w_mem_inst_w_mem_11__19_), .Y(w_mem_inst__abc_21378_n2562_1) );
  AND2X2 AND2X2_3198 ( .A(w_mem_inst__abc_21378_n1649_bF_buf0), .B(w_mem_inst_w_mem_9__19_), .Y(w_mem_inst__abc_21378_n2565) );
  AND2X2 AND2X2_3199 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf0), .B(w_mem_inst_w_mem_10__19_), .Y(w_mem_inst__abc_21378_n2566_1) );
  AND2X2 AND2X2_32 ( .A(e_reg_10_), .B(_auto_iopadmap_cc_313_execute_26059_10_), .Y(_abc_15724_n757_1) );
  AND2X2 AND2X2_320 ( .A(_abc_15724_n1312), .B(_abc_15724_n1325), .Y(_abc_15724_n1342) );
  AND2X2 AND2X2_3200 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf0), .B(w_mem_inst_w_mem_4__19_), .Y(w_mem_inst__abc_21378_n2568) );
  AND2X2 AND2X2_3201 ( .A(w_mem_inst__abc_21378_n1656_bF_buf0), .B(w_mem_inst_w_mem_12__19_), .Y(w_mem_inst__abc_21378_n2569) );
  AND2X2 AND2X2_3202 ( .A(w_mem_inst__abc_21378_n2574_1), .B(w_mem_inst__abc_21378_n2542_1), .Y(w_19_) );
  AND2X2 AND2X2_3203 ( .A(w_mem_inst__abc_21378_n2577), .B(w_mem_inst__abc_21378_n2579_1), .Y(w_mem_inst__abc_21378_n2580) );
  AND2X2 AND2X2_3204 ( .A(w_mem_inst_w_mem_2__19_), .B(w_mem_inst_w_mem_0__19_), .Y(w_mem_inst__abc_21378_n2583_1) );
  AND2X2 AND2X2_3205 ( .A(w_mem_inst__abc_21378_n2584), .B(w_mem_inst__abc_21378_n2582_1), .Y(w_mem_inst__abc_21378_n2585) );
  AND2X2 AND2X2_3206 ( .A(w_mem_inst__abc_21378_n2586_1), .B(w_mem_inst__abc_21378_n2588), .Y(w_mem_inst__abc_21378_n2589) );
  AND2X2 AND2X2_3207 ( .A(w_mem_inst__abc_21378_n1605_bF_buf4), .B(w_mem_inst_w_mem_15__20_), .Y(w_mem_inst__abc_21378_n2591_1) );
  AND2X2 AND2X2_3208 ( .A(w_mem_inst__abc_21378_n1649_bF_buf4), .B(w_mem_inst_w_mem_9__20_), .Y(w_mem_inst__abc_21378_n2592) );
  AND2X2 AND2X2_3209 ( .A(w_mem_inst__abc_21378_n1616_bF_buf4), .B(w_mem_inst_w_mem_5__20_), .Y(w_mem_inst__abc_21378_n2594_1) );
  AND2X2 AND2X2_321 ( .A(_abc_15724_n1316), .B(_abc_15724_n1342), .Y(_abc_15724_n1343_1) );
  AND2X2 AND2X2_3210 ( .A(w_mem_inst__abc_21378_n1656_bF_buf4), .B(w_mem_inst_w_mem_12__20_), .Y(w_mem_inst__abc_21378_n2595_1) );
  AND2X2 AND2X2_3211 ( .A(w_mem_inst__abc_21378_n1625_bF_buf4), .B(w_mem_inst_w_mem_2__20_), .Y(w_mem_inst__abc_21378_n2599_1) );
  AND2X2 AND2X2_3212 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf4), .B(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_21378_n2600) );
  AND2X2 AND2X2_3213 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf4), .B(w_mem_inst_w_mem_14__20_), .Y(w_mem_inst__abc_21378_n2602_1) );
  AND2X2 AND2X2_3214 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf4), .B(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_21378_n2603_1) );
  AND2X2 AND2X2_3215 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf4), .B(w_mem_inst_w_mem_6__20_), .Y(w_mem_inst__abc_21378_n2606_1) );
  AND2X2 AND2X2_3216 ( .A(w_mem_inst__abc_21378_n1645_bF_buf4), .B(w_mem_inst_w_mem_11__20_), .Y(w_mem_inst__abc_21378_n2607_1) );
  AND2X2 AND2X2_3217 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf4), .B(w_mem_inst_w_mem_0__20_), .Y(w_mem_inst__abc_21378_n2609) );
  AND2X2 AND2X2_3218 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf4), .B(w_mem_inst_w_mem_4__20_), .Y(w_mem_inst__abc_21378_n2610_1) );
  AND2X2 AND2X2_3219 ( .A(w_mem_inst__abc_21378_n1640_bF_buf4), .B(w_mem_inst_w_mem_7__20_), .Y(w_mem_inst__abc_21378_n2613) );
  AND2X2 AND2X2_322 ( .A(_abc_15724_n1345), .B(_abc_15724_n1340_1), .Y(_abc_15724_n1346) );
  AND2X2 AND2X2_3220 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf4), .B(w_mem_inst_w_mem_3__20_), .Y(w_mem_inst__abc_21378_n2614_1) );
  AND2X2 AND2X2_3221 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf4), .B(w_mem_inst_w_mem_1__20_), .Y(w_mem_inst__abc_21378_n2616) );
  AND2X2 AND2X2_3222 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf4), .B(w_mem_inst_w_mem_10__20_), .Y(w_mem_inst__abc_21378_n2617) );
  AND2X2 AND2X2_3223 ( .A(w_mem_inst__abc_21378_n2622_1), .B(w_mem_inst__abc_21378_n2590_1), .Y(w_20_) );
  AND2X2 AND2X2_3224 ( .A(w_mem_inst__abc_21378_n2625), .B(w_mem_inst__abc_21378_n2627_1), .Y(w_mem_inst__abc_21378_n2628) );
  AND2X2 AND2X2_3225 ( .A(w_mem_inst_w_mem_2__20_), .B(w_mem_inst_w_mem_0__20_), .Y(w_mem_inst__abc_21378_n2631_1) );
  AND2X2 AND2X2_3226 ( .A(w_mem_inst__abc_21378_n2632), .B(w_mem_inst__abc_21378_n2630_1), .Y(w_mem_inst__abc_21378_n2633) );
  AND2X2 AND2X2_3227 ( .A(w_mem_inst__abc_21378_n2634_1), .B(w_mem_inst__abc_21378_n2636), .Y(w_mem_inst__abc_21378_n2637) );
  AND2X2 AND2X2_3228 ( .A(w_mem_inst__abc_21378_n1605_bF_buf3), .B(w_mem_inst_w_mem_15__21_), .Y(w_mem_inst__abc_21378_n2639_1) );
  AND2X2 AND2X2_3229 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf3), .B(w_mem_inst_w_mem_3__21_), .Y(w_mem_inst__abc_21378_n2640) );
  AND2X2 AND2X2_323 ( .A(_abc_15724_n1348), .B(digest_update_bF_buf2), .Y(_abc_15724_n1349) );
  AND2X2 AND2X2_3230 ( .A(w_mem_inst__abc_21378_n1616_bF_buf3), .B(w_mem_inst_w_mem_5__21_), .Y(w_mem_inst__abc_21378_n2642_1) );
  AND2X2 AND2X2_3231 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf3), .B(w_mem_inst_w_mem_1__21_), .Y(w_mem_inst__abc_21378_n2643_1) );
  AND2X2 AND2X2_3232 ( .A(w_mem_inst__abc_21378_n1625_bF_buf3), .B(w_mem_inst_w_mem_2__21_), .Y(w_mem_inst__abc_21378_n2647_1) );
  AND2X2 AND2X2_3233 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf3), .B(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_21378_n2648) );
  AND2X2 AND2X2_3234 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf3), .B(w_mem_inst_w_mem_14__21_), .Y(w_mem_inst__abc_21378_n2650_1) );
  AND2X2 AND2X2_3235 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf3), .B(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_21378_n2651_1) );
  AND2X2 AND2X2_3236 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf3), .B(w_mem_inst_w_mem_6__21_), .Y(w_mem_inst__abc_21378_n2654_1) );
  AND2X2 AND2X2_3237 ( .A(w_mem_inst__abc_21378_n1640_bF_buf3), .B(w_mem_inst_w_mem_7__21_), .Y(w_mem_inst__abc_21378_n2655_1) );
  AND2X2 AND2X2_3238 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf3), .B(w_mem_inst_w_mem_0__21_), .Y(w_mem_inst__abc_21378_n2657) );
  AND2X2 AND2X2_3239 ( .A(w_mem_inst__abc_21378_n1645_bF_buf3), .B(w_mem_inst_w_mem_11__21_), .Y(w_mem_inst__abc_21378_n2658_1) );
  AND2X2 AND2X2_324 ( .A(_abc_15724_n1349), .B(_abc_15724_n1347), .Y(_abc_15724_n1350_1) );
  AND2X2 AND2X2_3240 ( .A(w_mem_inst__abc_21378_n1649_bF_buf3), .B(w_mem_inst_w_mem_9__21_), .Y(w_mem_inst__abc_21378_n2661) );
  AND2X2 AND2X2_3241 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf3), .B(w_mem_inst_w_mem_10__21_), .Y(w_mem_inst__abc_21378_n2662_1) );
  AND2X2 AND2X2_3242 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf3), .B(w_mem_inst_w_mem_4__21_), .Y(w_mem_inst__abc_21378_n2664) );
  AND2X2 AND2X2_3243 ( .A(w_mem_inst__abc_21378_n1656_bF_buf3), .B(w_mem_inst_w_mem_12__21_), .Y(w_mem_inst__abc_21378_n2665) );
  AND2X2 AND2X2_3244 ( .A(w_mem_inst__abc_21378_n2670_1), .B(w_mem_inst__abc_21378_n2638_1), .Y(w_21_) );
  AND2X2 AND2X2_3245 ( .A(w_mem_inst__abc_21378_n2673), .B(w_mem_inst__abc_21378_n2675_1), .Y(w_mem_inst__abc_21378_n2676) );
  AND2X2 AND2X2_3246 ( .A(w_mem_inst_w_mem_2__21_), .B(w_mem_inst_w_mem_0__21_), .Y(w_mem_inst__abc_21378_n2679_1) );
  AND2X2 AND2X2_3247 ( .A(w_mem_inst__abc_21378_n2680), .B(w_mem_inst__abc_21378_n2678_1), .Y(w_mem_inst__abc_21378_n2681) );
  AND2X2 AND2X2_3248 ( .A(w_mem_inst__abc_21378_n2682_1), .B(w_mem_inst__abc_21378_n2684), .Y(w_mem_inst__abc_21378_n2685) );
  AND2X2 AND2X2_3249 ( .A(w_mem_inst__abc_21378_n1605_bF_buf2), .B(w_mem_inst_w_mem_15__22_), .Y(w_mem_inst__abc_21378_n2687_1) );
  AND2X2 AND2X2_325 ( .A(_abc_15724_n1347), .B(_abc_15724_n1339), .Y(_abc_15724_n1352_1) );
  AND2X2 AND2X2_3250 ( .A(w_mem_inst__abc_21378_n1649_bF_buf2), .B(w_mem_inst_w_mem_9__22_), .Y(w_mem_inst__abc_21378_n2688) );
  AND2X2 AND2X2_3251 ( .A(w_mem_inst__abc_21378_n1616_bF_buf2), .B(w_mem_inst_w_mem_5__22_), .Y(w_mem_inst__abc_21378_n2690_1) );
  AND2X2 AND2X2_3252 ( .A(w_mem_inst__abc_21378_n1656_bF_buf2), .B(w_mem_inst_w_mem_12__22_), .Y(w_mem_inst__abc_21378_n2691_1) );
  AND2X2 AND2X2_3253 ( .A(w_mem_inst__abc_21378_n1625_bF_buf2), .B(w_mem_inst_w_mem_2__22_), .Y(w_mem_inst__abc_21378_n2695_1) );
  AND2X2 AND2X2_3254 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf2), .B(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_21378_n2696) );
  AND2X2 AND2X2_3255 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf2), .B(w_mem_inst_w_mem_14__22_), .Y(w_mem_inst__abc_21378_n2698_1) );
  AND2X2 AND2X2_3256 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf2), .B(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_21378_n2699_1) );
  AND2X2 AND2X2_3257 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf2), .B(w_mem_inst_w_mem_6__22_), .Y(w_mem_inst__abc_21378_n2702_1) );
  AND2X2 AND2X2_3258 ( .A(w_mem_inst__abc_21378_n1645_bF_buf2), .B(w_mem_inst_w_mem_11__22_), .Y(w_mem_inst__abc_21378_n2703_1) );
  AND2X2 AND2X2_3259 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf2), .B(w_mem_inst_w_mem_0__22_), .Y(w_mem_inst__abc_21378_n2705) );
  AND2X2 AND2X2_326 ( .A(_auto_iopadmap_cc_313_execute_26059_55_), .B(d_reg_23_), .Y(_abc_15724_n1354) );
  AND2X2 AND2X2_3260 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf2), .B(w_mem_inst_w_mem_4__22_), .Y(w_mem_inst__abc_21378_n2706_1) );
  AND2X2 AND2X2_3261 ( .A(w_mem_inst__abc_21378_n1640_bF_buf2), .B(w_mem_inst_w_mem_7__22_), .Y(w_mem_inst__abc_21378_n2709) );
  AND2X2 AND2X2_3262 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf2), .B(w_mem_inst_w_mem_3__22_), .Y(w_mem_inst__abc_21378_n2710_1) );
  AND2X2 AND2X2_3263 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf2), .B(w_mem_inst_w_mem_1__22_), .Y(w_mem_inst__abc_21378_n2712) );
  AND2X2 AND2X2_3264 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf2), .B(w_mem_inst_w_mem_10__22_), .Y(w_mem_inst__abc_21378_n2713) );
  AND2X2 AND2X2_3265 ( .A(w_mem_inst__abc_21378_n2718_1), .B(w_mem_inst__abc_21378_n2686_1), .Y(w_22_) );
  AND2X2 AND2X2_3266 ( .A(w_mem_inst__abc_21378_n2721), .B(w_mem_inst__abc_21378_n2723_1), .Y(w_mem_inst__abc_21378_n2724) );
  AND2X2 AND2X2_3267 ( .A(w_mem_inst_w_mem_2__22_), .B(w_mem_inst_w_mem_0__22_), .Y(w_mem_inst__abc_21378_n2727_1) );
  AND2X2 AND2X2_3268 ( .A(w_mem_inst__abc_21378_n2728), .B(w_mem_inst__abc_21378_n2726_1), .Y(w_mem_inst__abc_21378_n2729) );
  AND2X2 AND2X2_3269 ( .A(w_mem_inst__abc_21378_n2730_1), .B(w_mem_inst__abc_21378_n2732), .Y(w_mem_inst__abc_21378_n2733) );
  AND2X2 AND2X2_327 ( .A(_abc_15724_n1355), .B(_abc_15724_n1353), .Y(_abc_15724_n1356) );
  AND2X2 AND2X2_3270 ( .A(w_mem_inst__abc_21378_n1605_bF_buf1), .B(w_mem_inst_w_mem_15__23_), .Y(w_mem_inst__abc_21378_n2735_1) );
  AND2X2 AND2X2_3271 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf1), .B(w_mem_inst_w_mem_3__23_), .Y(w_mem_inst__abc_21378_n2736) );
  AND2X2 AND2X2_3272 ( .A(w_mem_inst__abc_21378_n1616_bF_buf1), .B(w_mem_inst_w_mem_5__23_), .Y(w_mem_inst__abc_21378_n2738_1) );
  AND2X2 AND2X2_3273 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf1), .B(w_mem_inst_w_mem_1__23_), .Y(w_mem_inst__abc_21378_n2739_1) );
  AND2X2 AND2X2_3274 ( .A(w_mem_inst__abc_21378_n1625_bF_buf1), .B(w_mem_inst_w_mem_2__23_), .Y(w_mem_inst__abc_21378_n2743_1) );
  AND2X2 AND2X2_3275 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf1), .B(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_21378_n2744) );
  AND2X2 AND2X2_3276 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf1), .B(w_mem_inst_w_mem_14__23_), .Y(w_mem_inst__abc_21378_n2746_1) );
  AND2X2 AND2X2_3277 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf1), .B(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_21378_n2747_1) );
  AND2X2 AND2X2_3278 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf1), .B(w_mem_inst_w_mem_6__23_), .Y(w_mem_inst__abc_21378_n2750_1) );
  AND2X2 AND2X2_3279 ( .A(w_mem_inst__abc_21378_n1640_bF_buf1), .B(w_mem_inst_w_mem_7__23_), .Y(w_mem_inst__abc_21378_n2751_1) );
  AND2X2 AND2X2_328 ( .A(_abc_15724_n1360), .B(_abc_15724_n1358), .Y(_abc_15724_n1361) );
  AND2X2 AND2X2_3280 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf1), .B(w_mem_inst_w_mem_0__23_), .Y(w_mem_inst__abc_21378_n2753) );
  AND2X2 AND2X2_3281 ( .A(w_mem_inst__abc_21378_n1645_bF_buf1), .B(w_mem_inst_w_mem_11__23_), .Y(w_mem_inst__abc_21378_n2754_1) );
  AND2X2 AND2X2_3282 ( .A(w_mem_inst__abc_21378_n1649_bF_buf1), .B(w_mem_inst_w_mem_9__23_), .Y(w_mem_inst__abc_21378_n2757) );
  AND2X2 AND2X2_3283 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf1), .B(w_mem_inst_w_mem_10__23_), .Y(w_mem_inst__abc_21378_n2758_1) );
  AND2X2 AND2X2_3284 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf1), .B(w_mem_inst_w_mem_4__23_), .Y(w_mem_inst__abc_21378_n2760) );
  AND2X2 AND2X2_3285 ( .A(w_mem_inst__abc_21378_n1656_bF_buf1), .B(w_mem_inst_w_mem_12__23_), .Y(w_mem_inst__abc_21378_n2761) );
  AND2X2 AND2X2_3286 ( .A(w_mem_inst__abc_21378_n2766_1), .B(w_mem_inst__abc_21378_n2734_1), .Y(w_23_) );
  AND2X2 AND2X2_3287 ( .A(w_mem_inst__abc_21378_n2769), .B(w_mem_inst__abc_21378_n2771_1), .Y(w_mem_inst__abc_21378_n2772) );
  AND2X2 AND2X2_3288 ( .A(w_mem_inst_w_mem_2__23_), .B(w_mem_inst_w_mem_0__23_), .Y(w_mem_inst__abc_21378_n2775_1) );
  AND2X2 AND2X2_3289 ( .A(w_mem_inst__abc_21378_n2776), .B(w_mem_inst__abc_21378_n2774_1), .Y(w_mem_inst__abc_21378_n2777) );
  AND2X2 AND2X2_329 ( .A(_abc_15724_n1361), .B(digest_update_bF_buf1), .Y(_abc_15724_n1362) );
  AND2X2 AND2X2_3290 ( .A(w_mem_inst__abc_21378_n2778_1), .B(w_mem_inst__abc_21378_n2780), .Y(w_mem_inst__abc_21378_n2781) );
  AND2X2 AND2X2_3291 ( .A(w_mem_inst__abc_21378_n1605_bF_buf0), .B(w_mem_inst_w_mem_15__24_), .Y(w_mem_inst__abc_21378_n2783_1) );
  AND2X2 AND2X2_3292 ( .A(w_mem_inst__abc_21378_n1649_bF_buf0), .B(w_mem_inst_w_mem_9__24_), .Y(w_mem_inst__abc_21378_n2784) );
  AND2X2 AND2X2_3293 ( .A(w_mem_inst__abc_21378_n1616_bF_buf0), .B(w_mem_inst_w_mem_5__24_), .Y(w_mem_inst__abc_21378_n2786_1) );
  AND2X2 AND2X2_3294 ( .A(w_mem_inst__abc_21378_n1656_bF_buf0), .B(w_mem_inst_w_mem_12__24_), .Y(w_mem_inst__abc_21378_n2787_1) );
  AND2X2 AND2X2_3295 ( .A(w_mem_inst__abc_21378_n1625_bF_buf0), .B(w_mem_inst_w_mem_2__24_), .Y(w_mem_inst__abc_21378_n2791_1) );
  AND2X2 AND2X2_3296 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf0), .B(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_21378_n2792) );
  AND2X2 AND2X2_3297 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf0), .B(w_mem_inst_w_mem_14__24_), .Y(w_mem_inst__abc_21378_n2794_1) );
  AND2X2 AND2X2_3298 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf0), .B(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_21378_n2795_1) );
  AND2X2 AND2X2_3299 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf0), .B(w_mem_inst_w_mem_6__24_), .Y(w_mem_inst__abc_21378_n2798_1) );
  AND2X2 AND2X2_33 ( .A(_abc_15724_n756), .B(_abc_15724_n757_1), .Y(_abc_15724_n758_1) );
  AND2X2 AND2X2_330 ( .A(_abc_15724_n907_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_55_), .Y(_abc_15724_n1363) );
  AND2X2 AND2X2_3300 ( .A(w_mem_inst__abc_21378_n1645_bF_buf0), .B(w_mem_inst_w_mem_11__24_), .Y(w_mem_inst__abc_21378_n2799_1) );
  AND2X2 AND2X2_3301 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf0), .B(w_mem_inst_w_mem_0__24_), .Y(w_mem_inst__abc_21378_n2801) );
  AND2X2 AND2X2_3302 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf0), .B(w_mem_inst_w_mem_4__24_), .Y(w_mem_inst__abc_21378_n2802_1) );
  AND2X2 AND2X2_3303 ( .A(w_mem_inst__abc_21378_n1640_bF_buf0), .B(w_mem_inst_w_mem_7__24_), .Y(w_mem_inst__abc_21378_n2805) );
  AND2X2 AND2X2_3304 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf0), .B(w_mem_inst_w_mem_3__24_), .Y(w_mem_inst__abc_21378_n2806_1) );
  AND2X2 AND2X2_3305 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf0), .B(w_mem_inst_w_mem_1__24_), .Y(w_mem_inst__abc_21378_n2808) );
  AND2X2 AND2X2_3306 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf0), .B(w_mem_inst_w_mem_10__24_), .Y(w_mem_inst__abc_21378_n2809) );
  AND2X2 AND2X2_3307 ( .A(w_mem_inst__abc_21378_n2814_1), .B(w_mem_inst__abc_21378_n2782_1), .Y(w_24_) );
  AND2X2 AND2X2_3308 ( .A(w_mem_inst__abc_21378_n2817), .B(w_mem_inst__abc_21378_n2819_1), .Y(w_mem_inst__abc_21378_n2820) );
  AND2X2 AND2X2_3309 ( .A(w_mem_inst_w_mem_2__24_), .B(w_mem_inst_w_mem_0__24_), .Y(w_mem_inst__abc_21378_n2823_1) );
  AND2X2 AND2X2_331 ( .A(_abc_15724_n907_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_56_), .Y(_abc_15724_n1365) );
  AND2X2 AND2X2_3310 ( .A(w_mem_inst__abc_21378_n2824), .B(w_mem_inst__abc_21378_n2822_1), .Y(w_mem_inst__abc_21378_n2825) );
  AND2X2 AND2X2_3311 ( .A(w_mem_inst__abc_21378_n2826_1), .B(w_mem_inst__abc_21378_n2828), .Y(w_mem_inst__abc_21378_n2829) );
  AND2X2 AND2X2_3312 ( .A(w_mem_inst__abc_21378_n1605_bF_buf4), .B(w_mem_inst_w_mem_15__25_), .Y(w_mem_inst__abc_21378_n2831_1) );
  AND2X2 AND2X2_3313 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf4), .B(w_mem_inst_w_mem_3__25_), .Y(w_mem_inst__abc_21378_n2832) );
  AND2X2 AND2X2_3314 ( .A(w_mem_inst__abc_21378_n1616_bF_buf4), .B(w_mem_inst_w_mem_5__25_), .Y(w_mem_inst__abc_21378_n2834_1) );
  AND2X2 AND2X2_3315 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf4), .B(w_mem_inst_w_mem_1__25_), .Y(w_mem_inst__abc_21378_n2835_1) );
  AND2X2 AND2X2_3316 ( .A(w_mem_inst__abc_21378_n1625_bF_buf4), .B(w_mem_inst_w_mem_2__25_), .Y(w_mem_inst__abc_21378_n2839_1) );
  AND2X2 AND2X2_3317 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf4), .B(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_21378_n2840) );
  AND2X2 AND2X2_3318 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf4), .B(w_mem_inst_w_mem_14__25_), .Y(w_mem_inst__abc_21378_n2842_1) );
  AND2X2 AND2X2_3319 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf4), .B(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_21378_n2843_1) );
  AND2X2 AND2X2_332 ( .A(_abc_15724_n1313), .B(_abc_15724_n1326), .Y(_abc_15724_n1366) );
  AND2X2 AND2X2_3320 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf4), .B(w_mem_inst_w_mem_6__25_), .Y(w_mem_inst__abc_21378_n2846_1) );
  AND2X2 AND2X2_3321 ( .A(w_mem_inst__abc_21378_n1640_bF_buf4), .B(w_mem_inst_w_mem_7__25_), .Y(w_mem_inst__abc_21378_n2847_1) );
  AND2X2 AND2X2_3322 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf4), .B(w_mem_inst_w_mem_0__25_), .Y(w_mem_inst__abc_21378_n2849) );
  AND2X2 AND2X2_3323 ( .A(w_mem_inst__abc_21378_n1645_bF_buf4), .B(w_mem_inst_w_mem_11__25_), .Y(w_mem_inst__abc_21378_n2850_1) );
  AND2X2 AND2X2_3324 ( .A(w_mem_inst__abc_21378_n1649_bF_buf4), .B(w_mem_inst_w_mem_9__25_), .Y(w_mem_inst__abc_21378_n2853) );
  AND2X2 AND2X2_3325 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf4), .B(w_mem_inst_w_mem_10__25_), .Y(w_mem_inst__abc_21378_n2854_1) );
  AND2X2 AND2X2_3326 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf4), .B(w_mem_inst_w_mem_4__25_), .Y(w_mem_inst__abc_21378_n2856) );
  AND2X2 AND2X2_3327 ( .A(w_mem_inst__abc_21378_n1656_bF_buf4), .B(w_mem_inst_w_mem_12__25_), .Y(w_mem_inst__abc_21378_n2857) );
  AND2X2 AND2X2_3328 ( .A(w_mem_inst__abc_21378_n2862_1), .B(w_mem_inst__abc_21378_n2830_1), .Y(w_25_) );
  AND2X2 AND2X2_3329 ( .A(w_mem_inst__abc_21378_n2865), .B(w_mem_inst__abc_21378_n2867_1), .Y(w_mem_inst__abc_21378_n2868) );
  AND2X2 AND2X2_333 ( .A(_abc_15724_n1340_1), .B(_abc_15724_n1356), .Y(_abc_15724_n1367) );
  AND2X2 AND2X2_3330 ( .A(w_mem_inst_w_mem_2__25_), .B(w_mem_inst_w_mem_0__25_), .Y(w_mem_inst__abc_21378_n2871_1) );
  AND2X2 AND2X2_3331 ( .A(w_mem_inst__abc_21378_n2872), .B(w_mem_inst__abc_21378_n2870_1), .Y(w_mem_inst__abc_21378_n2873) );
  AND2X2 AND2X2_3332 ( .A(w_mem_inst__abc_21378_n2874_1), .B(w_mem_inst__abc_21378_n2876), .Y(w_mem_inst__abc_21378_n2877) );
  AND2X2 AND2X2_3333 ( .A(w_mem_inst__abc_21378_n1605_bF_buf3), .B(w_mem_inst_w_mem_15__26_), .Y(w_mem_inst__abc_21378_n2879_1) );
  AND2X2 AND2X2_3334 ( .A(w_mem_inst__abc_21378_n1649_bF_buf3), .B(w_mem_inst_w_mem_9__26_), .Y(w_mem_inst__abc_21378_n2880) );
  AND2X2 AND2X2_3335 ( .A(w_mem_inst__abc_21378_n1616_bF_buf3), .B(w_mem_inst_w_mem_5__26_), .Y(w_mem_inst__abc_21378_n2882_1) );
  AND2X2 AND2X2_3336 ( .A(w_mem_inst__abc_21378_n1656_bF_buf3), .B(w_mem_inst_w_mem_12__26_), .Y(w_mem_inst__abc_21378_n2883_1) );
  AND2X2 AND2X2_3337 ( .A(w_mem_inst__abc_21378_n1625_bF_buf3), .B(w_mem_inst_w_mem_2__26_), .Y(w_mem_inst__abc_21378_n2887_1) );
  AND2X2 AND2X2_3338 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf3), .B(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_21378_n2888) );
  AND2X2 AND2X2_3339 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf3), .B(w_mem_inst_w_mem_14__26_), .Y(w_mem_inst__abc_21378_n2890_1) );
  AND2X2 AND2X2_334 ( .A(_abc_15724_n1366), .B(_abc_15724_n1367), .Y(_abc_15724_n1368_1) );
  AND2X2 AND2X2_3340 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf3), .B(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_21378_n2891_1) );
  AND2X2 AND2X2_3341 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf3), .B(w_mem_inst_w_mem_6__26_), .Y(w_mem_inst__abc_21378_n2894_1) );
  AND2X2 AND2X2_3342 ( .A(w_mem_inst__abc_21378_n1645_bF_buf3), .B(w_mem_inst_w_mem_11__26_), .Y(w_mem_inst__abc_21378_n2895_1) );
  AND2X2 AND2X2_3343 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf3), .B(w_mem_inst_w_mem_0__26_), .Y(w_mem_inst__abc_21378_n2897) );
  AND2X2 AND2X2_3344 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf3), .B(w_mem_inst_w_mem_4__26_), .Y(w_mem_inst__abc_21378_n2898_1) );
  AND2X2 AND2X2_3345 ( .A(w_mem_inst__abc_21378_n1640_bF_buf3), .B(w_mem_inst_w_mem_7__26_), .Y(w_mem_inst__abc_21378_n2901) );
  AND2X2 AND2X2_3346 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf3), .B(w_mem_inst_w_mem_3__26_), .Y(w_mem_inst__abc_21378_n2902_1) );
  AND2X2 AND2X2_3347 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf3), .B(w_mem_inst_w_mem_1__26_), .Y(w_mem_inst__abc_21378_n2904) );
  AND2X2 AND2X2_3348 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf3), .B(w_mem_inst_w_mem_10__26_), .Y(w_mem_inst__abc_21378_n2905) );
  AND2X2 AND2X2_3349 ( .A(w_mem_inst__abc_21378_n2910_1), .B(w_mem_inst__abc_21378_n2878_1), .Y(w_26_) );
  AND2X2 AND2X2_335 ( .A(_abc_15724_n1305_1), .B(_abc_15724_n1368_1), .Y(_abc_15724_n1369_1) );
  AND2X2 AND2X2_3350 ( .A(w_mem_inst__abc_21378_n2913), .B(w_mem_inst__abc_21378_n2915_1), .Y(w_mem_inst__abc_21378_n2916) );
  AND2X2 AND2X2_3351 ( .A(w_mem_inst_w_mem_2__26_), .B(w_mem_inst_w_mem_0__26_), .Y(w_mem_inst__abc_21378_n2919_1) );
  AND2X2 AND2X2_3352 ( .A(w_mem_inst__abc_21378_n2920), .B(w_mem_inst__abc_21378_n2918_1), .Y(w_mem_inst__abc_21378_n2921) );
  AND2X2 AND2X2_3353 ( .A(w_mem_inst__abc_21378_n2922_1), .B(w_mem_inst__abc_21378_n2924), .Y(w_mem_inst__abc_21378_n2925) );
  AND2X2 AND2X2_3354 ( .A(w_mem_inst__abc_21378_n1605_bF_buf2), .B(w_mem_inst_w_mem_15__27_), .Y(w_mem_inst__abc_21378_n2927_1) );
  AND2X2 AND2X2_3355 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf2), .B(w_mem_inst_w_mem_3__27_), .Y(w_mem_inst__abc_21378_n2928) );
  AND2X2 AND2X2_3356 ( .A(w_mem_inst__abc_21378_n1616_bF_buf2), .B(w_mem_inst_w_mem_5__27_), .Y(w_mem_inst__abc_21378_n2930_1) );
  AND2X2 AND2X2_3357 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf2), .B(w_mem_inst_w_mem_1__27_), .Y(w_mem_inst__abc_21378_n2931_1) );
  AND2X2 AND2X2_3358 ( .A(w_mem_inst__abc_21378_n1625_bF_buf2), .B(w_mem_inst_w_mem_2__27_), .Y(w_mem_inst__abc_21378_n2935_1) );
  AND2X2 AND2X2_3359 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf2), .B(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_21378_n2936) );
  AND2X2 AND2X2_336 ( .A(_abc_15724_n1371_1), .B(_abc_15724_n1367), .Y(_abc_15724_n1372) );
  AND2X2 AND2X2_3360 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf2), .B(w_mem_inst_w_mem_14__27_), .Y(w_mem_inst__abc_21378_n2938_1) );
  AND2X2 AND2X2_3361 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf2), .B(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_21378_n2939_1) );
  AND2X2 AND2X2_3362 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf2), .B(w_mem_inst_w_mem_6__27_), .Y(w_mem_inst__abc_21378_n2942_1) );
  AND2X2 AND2X2_3363 ( .A(w_mem_inst__abc_21378_n1640_bF_buf2), .B(w_mem_inst_w_mem_7__27_), .Y(w_mem_inst__abc_21378_n2943_1) );
  AND2X2 AND2X2_3364 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf2), .B(w_mem_inst_w_mem_0__27_), .Y(w_mem_inst__abc_21378_n2945) );
  AND2X2 AND2X2_3365 ( .A(w_mem_inst__abc_21378_n1645_bF_buf2), .B(w_mem_inst_w_mem_11__27_), .Y(w_mem_inst__abc_21378_n2946_1) );
  AND2X2 AND2X2_3366 ( .A(w_mem_inst__abc_21378_n1649_bF_buf2), .B(w_mem_inst_w_mem_9__27_), .Y(w_mem_inst__abc_21378_n2949) );
  AND2X2 AND2X2_3367 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf2), .B(w_mem_inst_w_mem_10__27_), .Y(w_mem_inst__abc_21378_n2950_1) );
  AND2X2 AND2X2_3368 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf2), .B(w_mem_inst_w_mem_4__27_), .Y(w_mem_inst__abc_21378_n2952) );
  AND2X2 AND2X2_3369 ( .A(w_mem_inst__abc_21378_n1656_bF_buf2), .B(w_mem_inst_w_mem_12__27_), .Y(w_mem_inst__abc_21378_n2953) );
  AND2X2 AND2X2_337 ( .A(_abc_15724_n1353), .B(_abc_15724_n1338), .Y(_abc_15724_n1373) );
  AND2X2 AND2X2_3370 ( .A(w_mem_inst__abc_21378_n2958_1), .B(w_mem_inst__abc_21378_n2926_1), .Y(w_27_) );
  AND2X2 AND2X2_3371 ( .A(w_mem_inst__abc_21378_n2961), .B(w_mem_inst__abc_21378_n2963_1), .Y(w_mem_inst__abc_21378_n2964) );
  AND2X2 AND2X2_3372 ( .A(w_mem_inst_w_mem_2__27_), .B(w_mem_inst_w_mem_0__27_), .Y(w_mem_inst__abc_21378_n2967_1) );
  AND2X2 AND2X2_3373 ( .A(w_mem_inst__abc_21378_n2968), .B(w_mem_inst__abc_21378_n2966_1), .Y(w_mem_inst__abc_21378_n2969) );
  AND2X2 AND2X2_3374 ( .A(w_mem_inst__abc_21378_n2970_1), .B(w_mem_inst__abc_21378_n2972), .Y(w_mem_inst__abc_21378_n2973) );
  AND2X2 AND2X2_3375 ( .A(w_mem_inst__abc_21378_n1605_bF_buf1), .B(w_mem_inst_w_mem_15__28_), .Y(w_mem_inst__abc_21378_n2975_1) );
  AND2X2 AND2X2_3376 ( .A(w_mem_inst__abc_21378_n1649_bF_buf1), .B(w_mem_inst_w_mem_9__28_), .Y(w_mem_inst__abc_21378_n2976) );
  AND2X2 AND2X2_3377 ( .A(w_mem_inst__abc_21378_n1616_bF_buf1), .B(w_mem_inst_w_mem_5__28_), .Y(w_mem_inst__abc_21378_n2978_1) );
  AND2X2 AND2X2_3378 ( .A(w_mem_inst__abc_21378_n1656_bF_buf1), .B(w_mem_inst_w_mem_12__28_), .Y(w_mem_inst__abc_21378_n2979_1) );
  AND2X2 AND2X2_3379 ( .A(w_mem_inst__abc_21378_n1625_bF_buf1), .B(w_mem_inst_w_mem_2__28_), .Y(w_mem_inst__abc_21378_n2983_1) );
  AND2X2 AND2X2_338 ( .A(_abc_15724_n1307), .B(_abc_15724_n1368_1), .Y(_abc_15724_n1377_1) );
  AND2X2 AND2X2_3380 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf1), .B(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_21378_n2984) );
  AND2X2 AND2X2_3381 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf1), .B(w_mem_inst_w_mem_14__28_), .Y(w_mem_inst__abc_21378_n2986_1) );
  AND2X2 AND2X2_3382 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf1), .B(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_21378_n2987_1) );
  AND2X2 AND2X2_3383 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf1), .B(w_mem_inst_w_mem_6__28_), .Y(w_mem_inst__abc_21378_n2990_1) );
  AND2X2 AND2X2_3384 ( .A(w_mem_inst__abc_21378_n1645_bF_buf1), .B(w_mem_inst_w_mem_11__28_), .Y(w_mem_inst__abc_21378_n2991_1) );
  AND2X2 AND2X2_3385 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf1), .B(w_mem_inst_w_mem_0__28_), .Y(w_mem_inst__abc_21378_n2993) );
  AND2X2 AND2X2_3386 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf1), .B(w_mem_inst_w_mem_4__28_), .Y(w_mem_inst__abc_21378_n2994_1) );
  AND2X2 AND2X2_3387 ( .A(w_mem_inst__abc_21378_n1640_bF_buf1), .B(w_mem_inst_w_mem_7__28_), .Y(w_mem_inst__abc_21378_n2997) );
  AND2X2 AND2X2_3388 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf1), .B(w_mem_inst_w_mem_3__28_), .Y(w_mem_inst__abc_21378_n2998_1) );
  AND2X2 AND2X2_3389 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf1), .B(w_mem_inst_w_mem_1__28_), .Y(w_mem_inst__abc_21378_n3000) );
  AND2X2 AND2X2_339 ( .A(_abc_15724_n1243), .B(_abc_15724_n1377_1), .Y(_abc_15724_n1378_1) );
  AND2X2 AND2X2_3390 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf1), .B(w_mem_inst_w_mem_10__28_), .Y(w_mem_inst__abc_21378_n3001) );
  AND2X2 AND2X2_3391 ( .A(w_mem_inst__abc_21378_n3006_1), .B(w_mem_inst__abc_21378_n2974_1), .Y(w_28_) );
  AND2X2 AND2X2_3392 ( .A(w_mem_inst__abc_21378_n3009), .B(w_mem_inst__abc_21378_n3011_1), .Y(w_mem_inst__abc_21378_n3012) );
  AND2X2 AND2X2_3393 ( .A(w_mem_inst_w_mem_2__28_), .B(w_mem_inst_w_mem_0__28_), .Y(w_mem_inst__abc_21378_n3015_1) );
  AND2X2 AND2X2_3394 ( .A(w_mem_inst__abc_21378_n3016), .B(w_mem_inst__abc_21378_n3014_1), .Y(w_mem_inst__abc_21378_n3017) );
  AND2X2 AND2X2_3395 ( .A(w_mem_inst__abc_21378_n3018_1), .B(w_mem_inst__abc_21378_n3020), .Y(w_mem_inst__abc_21378_n3021) );
  AND2X2 AND2X2_3396 ( .A(w_mem_inst__abc_21378_n1605_bF_buf0), .B(w_mem_inst_w_mem_15__29_), .Y(w_mem_inst__abc_21378_n3023_1) );
  AND2X2 AND2X2_3397 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf0), .B(w_mem_inst_w_mem_3__29_), .Y(w_mem_inst__abc_21378_n3024) );
  AND2X2 AND2X2_3398 ( .A(w_mem_inst__abc_21378_n1616_bF_buf0), .B(w_mem_inst_w_mem_5__29_), .Y(w_mem_inst__abc_21378_n3026_1) );
  AND2X2 AND2X2_3399 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf0), .B(w_mem_inst_w_mem_1__29_), .Y(w_mem_inst__abc_21378_n3027_1) );
  AND2X2 AND2X2_34 ( .A(_abc_15724_n760_1), .B(_abc_15724_n756), .Y(_abc_15724_n761) );
  AND2X2 AND2X2_340 ( .A(_auto_iopadmap_cc_313_execute_26059_56_), .B(d_reg_24_), .Y(_abc_15724_n1381) );
  AND2X2 AND2X2_3400 ( .A(w_mem_inst__abc_21378_n1625_bF_buf0), .B(w_mem_inst_w_mem_2__29_), .Y(w_mem_inst__abc_21378_n3031_1) );
  AND2X2 AND2X2_3401 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf0), .B(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_21378_n3032) );
  AND2X2 AND2X2_3402 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf0), .B(w_mem_inst_w_mem_14__29_), .Y(w_mem_inst__abc_21378_n3034_1) );
  AND2X2 AND2X2_3403 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf0), .B(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_21378_n3035_1) );
  AND2X2 AND2X2_3404 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf0), .B(w_mem_inst_w_mem_6__29_), .Y(w_mem_inst__abc_21378_n3038_1) );
  AND2X2 AND2X2_3405 ( .A(w_mem_inst__abc_21378_n1640_bF_buf0), .B(w_mem_inst_w_mem_7__29_), .Y(w_mem_inst__abc_21378_n3039_1) );
  AND2X2 AND2X2_3406 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf0), .B(w_mem_inst_w_mem_0__29_), .Y(w_mem_inst__abc_21378_n3041) );
  AND2X2 AND2X2_3407 ( .A(w_mem_inst__abc_21378_n1645_bF_buf0), .B(w_mem_inst_w_mem_11__29_), .Y(w_mem_inst__abc_21378_n3042_1) );
  AND2X2 AND2X2_3408 ( .A(w_mem_inst__abc_21378_n1649_bF_buf0), .B(w_mem_inst_w_mem_9__29_), .Y(w_mem_inst__abc_21378_n3045) );
  AND2X2 AND2X2_3409 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf0), .B(w_mem_inst_w_mem_10__29_), .Y(w_mem_inst__abc_21378_n3046_1) );
  AND2X2 AND2X2_341 ( .A(_abc_15724_n1382), .B(_abc_15724_n1380), .Y(_abc_15724_n1383) );
  AND2X2 AND2X2_3410 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf0), .B(w_mem_inst_w_mem_4__29_), .Y(w_mem_inst__abc_21378_n3048) );
  AND2X2 AND2X2_3411 ( .A(w_mem_inst__abc_21378_n1656_bF_buf0), .B(w_mem_inst_w_mem_12__29_), .Y(w_mem_inst__abc_21378_n3049) );
  AND2X2 AND2X2_3412 ( .A(w_mem_inst__abc_21378_n3054_1), .B(w_mem_inst__abc_21378_n3022_1), .Y(w_29_) );
  AND2X2 AND2X2_3413 ( .A(w_mem_inst__abc_21378_n3057), .B(w_mem_inst__abc_21378_n3059_1), .Y(w_mem_inst__abc_21378_n3060) );
  AND2X2 AND2X2_3414 ( .A(w_mem_inst_w_mem_2__29_), .B(w_mem_inst_w_mem_0__29_), .Y(w_mem_inst__abc_21378_n3063_1) );
  AND2X2 AND2X2_3415 ( .A(w_mem_inst__abc_21378_n3064), .B(w_mem_inst__abc_21378_n3062_1), .Y(w_mem_inst__abc_21378_n3065) );
  AND2X2 AND2X2_3416 ( .A(w_mem_inst__abc_21378_n3066_1), .B(w_mem_inst__abc_21378_n3068), .Y(w_mem_inst__abc_21378_n3069) );
  AND2X2 AND2X2_3417 ( .A(w_mem_inst__abc_21378_n1605_bF_buf4), .B(w_mem_inst_w_mem_15__30_), .Y(w_mem_inst__abc_21378_n3071_1) );
  AND2X2 AND2X2_3418 ( .A(w_mem_inst__abc_21378_n1649_bF_buf4), .B(w_mem_inst_w_mem_9__30_), .Y(w_mem_inst__abc_21378_n3072) );
  AND2X2 AND2X2_3419 ( .A(w_mem_inst__abc_21378_n1616_bF_buf4), .B(w_mem_inst_w_mem_5__30_), .Y(w_mem_inst__abc_21378_n3074_1) );
  AND2X2 AND2X2_342 ( .A(_abc_15724_n1379_1), .B(_abc_15724_n1383), .Y(_abc_15724_n1385) );
  AND2X2 AND2X2_3420 ( .A(w_mem_inst__abc_21378_n1656_bF_buf4), .B(w_mem_inst_w_mem_12__30_), .Y(w_mem_inst__abc_21378_n3075_1) );
  AND2X2 AND2X2_3421 ( .A(w_mem_inst__abc_21378_n1625_bF_buf4), .B(w_mem_inst_w_mem_2__30_), .Y(w_mem_inst__abc_21378_n3079_1) );
  AND2X2 AND2X2_3422 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf4), .B(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_21378_n3080) );
  AND2X2 AND2X2_3423 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf4), .B(w_mem_inst_w_mem_14__30_), .Y(w_mem_inst__abc_21378_n3082_1) );
  AND2X2 AND2X2_3424 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf4), .B(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_21378_n3083_1) );
  AND2X2 AND2X2_3425 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf4), .B(w_mem_inst_w_mem_6__30_), .Y(w_mem_inst__abc_21378_n3086_1) );
  AND2X2 AND2X2_3426 ( .A(w_mem_inst__abc_21378_n1645_bF_buf4), .B(w_mem_inst_w_mem_11__30_), .Y(w_mem_inst__abc_21378_n3087_1) );
  AND2X2 AND2X2_3427 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf4), .B(w_mem_inst_w_mem_0__30_), .Y(w_mem_inst__abc_21378_n3089) );
  AND2X2 AND2X2_3428 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf4), .B(w_mem_inst_w_mem_4__30_), .Y(w_mem_inst__abc_21378_n3090_1) );
  AND2X2 AND2X2_3429 ( .A(w_mem_inst__abc_21378_n1640_bF_buf4), .B(w_mem_inst_w_mem_7__30_), .Y(w_mem_inst__abc_21378_n3093) );
  AND2X2 AND2X2_343 ( .A(_abc_15724_n1386), .B(_abc_15724_n1384), .Y(_abc_15724_n1387) );
  AND2X2 AND2X2_3430 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf4), .B(w_mem_inst_w_mem_3__30_), .Y(w_mem_inst__abc_21378_n3094_1) );
  AND2X2 AND2X2_3431 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf4), .B(w_mem_inst_w_mem_1__30_), .Y(w_mem_inst__abc_21378_n3096) );
  AND2X2 AND2X2_3432 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf4), .B(w_mem_inst_w_mem_10__30_), .Y(w_mem_inst__abc_21378_n3097) );
  AND2X2 AND2X2_3433 ( .A(w_mem_inst__abc_21378_n3102_1), .B(w_mem_inst__abc_21378_n3070_1), .Y(w_30_) );
  AND2X2 AND2X2_3434 ( .A(w_mem_inst__abc_21378_n3105), .B(w_mem_inst__abc_21378_n3107_1), .Y(w_mem_inst__abc_21378_n3108) );
  AND2X2 AND2X2_3435 ( .A(w_mem_inst_w_mem_2__30_), .B(w_mem_inst_w_mem_0__30_), .Y(w_mem_inst__abc_21378_n3111_1) );
  AND2X2 AND2X2_3436 ( .A(w_mem_inst__abc_21378_n3112), .B(w_mem_inst__abc_21378_n3110_1), .Y(w_mem_inst__abc_21378_n3113) );
  AND2X2 AND2X2_3437 ( .A(w_mem_inst__abc_21378_n3114_1), .B(w_mem_inst__abc_21378_n3116), .Y(w_mem_inst__abc_21378_n3117) );
  AND2X2 AND2X2_3438 ( .A(w_mem_inst__abc_21378_n1605_bF_buf3), .B(w_mem_inst_w_mem_15__31_), .Y(w_mem_inst__abc_21378_n3119_1) );
  AND2X2 AND2X2_3439 ( .A(w_mem_inst__abc_21378_n1610_1_bF_buf3), .B(w_mem_inst_w_mem_3__31_), .Y(w_mem_inst__abc_21378_n3120) );
  AND2X2 AND2X2_344 ( .A(_abc_15724_n1387), .B(digest_update_bF_buf0), .Y(_abc_15724_n1388) );
  AND2X2 AND2X2_3440 ( .A(w_mem_inst__abc_21378_n1616_bF_buf3), .B(w_mem_inst_w_mem_5__31_), .Y(w_mem_inst__abc_21378_n3122_1) );
  AND2X2 AND2X2_3441 ( .A(w_mem_inst__abc_21378_n1618_1_bF_buf3), .B(w_mem_inst_w_mem_1__31_), .Y(w_mem_inst__abc_21378_n3123_1) );
  AND2X2 AND2X2_3442 ( .A(w_mem_inst__abc_21378_n1625_bF_buf3), .B(w_mem_inst_w_mem_2__31_), .Y(w_mem_inst__abc_21378_n3127_1) );
  AND2X2 AND2X2_3443 ( .A(w_mem_inst__abc_21378_n1627_1_bF_buf3), .B(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_21378_n3128) );
  AND2X2 AND2X2_3444 ( .A(w_mem_inst__abc_21378_n1630_1_bF_buf3), .B(w_mem_inst_w_mem_14__31_), .Y(w_mem_inst__abc_21378_n3130_1) );
  AND2X2 AND2X2_3445 ( .A(w_mem_inst__abc_21378_n1634_1_bF_buf3), .B(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_21378_n3131_1) );
  AND2X2 AND2X2_3446 ( .A(w_mem_inst__abc_21378_n1638_1_bF_buf3), .B(w_mem_inst_w_mem_6__31_), .Y(w_mem_inst__abc_21378_n3134_1) );
  AND2X2 AND2X2_3447 ( .A(w_mem_inst__abc_21378_n1640_bF_buf3), .B(w_mem_inst_w_mem_7__31_), .Y(w_mem_inst__abc_21378_n3135_1) );
  AND2X2 AND2X2_3448 ( .A(w_mem_inst__abc_21378_n1643_1_bF_buf3), .B(w_mem_inst_w_mem_0__31_), .Y(w_mem_inst__abc_21378_n3137) );
  AND2X2 AND2X2_3449 ( .A(w_mem_inst__abc_21378_n1645_bF_buf3), .B(w_mem_inst_w_mem_11__31_), .Y(w_mem_inst__abc_21378_n3138_1) );
  AND2X2 AND2X2_345 ( .A(_abc_15724_n907_1_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_57_), .Y(_abc_15724_n1390_1) );
  AND2X2 AND2X2_3450 ( .A(w_mem_inst__abc_21378_n1649_bF_buf3), .B(w_mem_inst_w_mem_9__31_), .Y(w_mem_inst__abc_21378_n3141) );
  AND2X2 AND2X2_3451 ( .A(w_mem_inst__abc_21378_n1651_1_bF_buf3), .B(w_mem_inst_w_mem_10__31_), .Y(w_mem_inst__abc_21378_n3142_1) );
  AND2X2 AND2X2_3452 ( .A(w_mem_inst__abc_21378_n1654_1_bF_buf3), .B(w_mem_inst_w_mem_4__31_), .Y(w_mem_inst__abc_21378_n3144) );
  AND2X2 AND2X2_3453 ( .A(w_mem_inst__abc_21378_n1656_bF_buf3), .B(w_mem_inst_w_mem_12__31_), .Y(w_mem_inst__abc_21378_n3145) );
  AND2X2 AND2X2_3454 ( .A(w_mem_inst__abc_21378_n3150_1), .B(w_mem_inst__abc_21378_n3118_1), .Y(w_31_) );
  AND2X2 AND2X2_3455 ( .A(w_mem_inst__abc_21378_n1586_bF_buf1), .B(round_ctr_inc_bF_buf12), .Y(w_mem_inst__abc_21378_n3152) );
  AND2X2 AND2X2_3456 ( .A(w_mem_inst__abc_21378_n1601_1), .B(w_mem_inst__abc_21378_n3152_bF_buf63), .Y(w_mem_inst__abc_21378_n3153) );
  AND2X2 AND2X2_3457 ( .A(round_ctr_rst_bF_buf60), .B(\block[0] ), .Y(w_mem_inst__abc_21378_n3155_1) );
  AND2X2 AND2X2_3458 ( .A(w_mem_inst__abc_21378_n3156_bF_buf4), .B(w_mem_inst_w_mem_15__0_), .Y(w_mem_inst__abc_21378_n3157) );
  AND2X2 AND2X2_3459 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf63), .B(w_mem_inst__abc_21378_n3158_1), .Y(w_mem_inst__abc_21378_n3159_1) );
  AND2X2 AND2X2_346 ( .A(_auto_iopadmap_cc_313_execute_26059_57_), .B(d_reg_25_), .Y(_abc_15724_n1392) );
  AND2X2 AND2X2_3460 ( .A(w_mem_inst__abc_21378_n1677), .B(w_mem_inst__abc_21378_n3152_bF_buf61), .Y(w_mem_inst__abc_21378_n3161) );
  AND2X2 AND2X2_3461 ( .A(round_ctr_rst_bF_buf58), .B(\block[1] ), .Y(w_mem_inst__abc_21378_n3162_1) );
  AND2X2 AND2X2_3462 ( .A(w_mem_inst__abc_21378_n3156_bF_buf3), .B(w_mem_inst_w_mem_15__1_), .Y(w_mem_inst__abc_21378_n3163_1) );
  AND2X2 AND2X2_3463 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf62), .B(w_mem_inst__abc_21378_n3164), .Y(w_mem_inst__abc_21378_n3165) );
  AND2X2 AND2X2_3464 ( .A(round_ctr_rst_bF_buf57), .B(\block[2] ), .Y(w_mem_inst__abc_21378_n3167_1) );
  AND2X2 AND2X2_3465 ( .A(w_mem_inst__abc_21378_n3156_bF_buf2), .B(w_mem_inst_w_mem_15__2_), .Y(w_mem_inst__abc_21378_n3168) );
  AND2X2 AND2X2_3466 ( .A(w_mem_inst__abc_21378_n3171_1), .B(w_mem_inst__abc_21378_n3170_1), .Y(w_mem_inst__0w_mem_15__31_0__2_) );
  AND2X2 AND2X2_3467 ( .A(w_mem_inst__abc_21378_n1773), .B(w_mem_inst__abc_21378_n3152_bF_buf59), .Y(w_mem_inst__abc_21378_n3173) );
  AND2X2 AND2X2_3468 ( .A(round_ctr_rst_bF_buf56), .B(\block[3] ), .Y(w_mem_inst__abc_21378_n3174_1) );
  AND2X2 AND2X2_3469 ( .A(w_mem_inst__abc_21378_n3156_bF_buf1), .B(w_mem_inst_w_mem_15__3_), .Y(w_mem_inst__abc_21378_n3175_1) );
  AND2X2 AND2X2_347 ( .A(_abc_15724_n1393_1), .B(_abc_15724_n1391_1), .Y(_abc_15724_n1394) );
  AND2X2 AND2X2_3470 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf60), .B(w_mem_inst__abc_21378_n3176), .Y(w_mem_inst__abc_21378_n3177) );
  AND2X2 AND2X2_3471 ( .A(round_ctr_rst_bF_buf55), .B(\block[4] ), .Y(w_mem_inst__abc_21378_n3179_1) );
  AND2X2 AND2X2_3472 ( .A(w_mem_inst__abc_21378_n3156_bF_buf0), .B(w_mem_inst_w_mem_15__4_), .Y(w_mem_inst__abc_21378_n3180) );
  AND2X2 AND2X2_3473 ( .A(w_mem_inst__abc_21378_n3183_1), .B(w_mem_inst__abc_21378_n3182_1), .Y(w_mem_inst__0w_mem_15__31_0__4_) );
  AND2X2 AND2X2_3474 ( .A(w_mem_inst__abc_21378_n1869), .B(w_mem_inst__abc_21378_n3152_bF_buf57), .Y(w_mem_inst__abc_21378_n3185) );
  AND2X2 AND2X2_3475 ( .A(round_ctr_rst_bF_buf54), .B(\block[5] ), .Y(w_mem_inst__abc_21378_n3186_1) );
  AND2X2 AND2X2_3476 ( .A(w_mem_inst__abc_21378_n3156_bF_buf4), .B(w_mem_inst_w_mem_15__5_), .Y(w_mem_inst__abc_21378_n3187_1) );
  AND2X2 AND2X2_3477 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf58), .B(w_mem_inst__abc_21378_n3188), .Y(w_mem_inst__abc_21378_n3189) );
  AND2X2 AND2X2_3478 ( .A(w_mem_inst__abc_21378_n1917), .B(w_mem_inst__abc_21378_n3152_bF_buf56), .Y(w_mem_inst__abc_21378_n3191_1) );
  AND2X2 AND2X2_3479 ( .A(round_ctr_rst_bF_buf53), .B(\block[6] ), .Y(w_mem_inst__abc_21378_n3192) );
  AND2X2 AND2X2_348 ( .A(_abc_15724_n1109_1), .B(_abc_15724_n1102), .Y(_abc_15724_n1399_1) );
  AND2X2 AND2X2_3480 ( .A(w_mem_inst__abc_21378_n3156_bF_buf3), .B(w_mem_inst_w_mem_15__6_), .Y(w_mem_inst__abc_21378_n3193) );
  AND2X2 AND2X2_3481 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf57), .B(w_mem_inst__abc_21378_n3194_1), .Y(w_mem_inst__abc_21378_n3195_1) );
  AND2X2 AND2X2_3482 ( .A(w_mem_inst__abc_21378_n1965), .B(w_mem_inst__abc_21378_n3152_bF_buf55), .Y(w_mem_inst__abc_21378_n3197) );
  AND2X2 AND2X2_3483 ( .A(round_ctr_rst_bF_buf52), .B(\block[7] ), .Y(w_mem_inst__abc_21378_n3198_1) );
  AND2X2 AND2X2_3484 ( .A(w_mem_inst__abc_21378_n3156_bF_buf2), .B(w_mem_inst_w_mem_15__7_), .Y(w_mem_inst__abc_21378_n3199_1) );
  AND2X2 AND2X2_3485 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf56), .B(w_mem_inst__abc_21378_n3200), .Y(w_mem_inst__abc_21378_n3201) );
  AND2X2 AND2X2_3486 ( .A(w_mem_inst__abc_21378_n2013), .B(w_mem_inst__abc_21378_n3152_bF_buf54), .Y(w_mem_inst__abc_21378_n3203_1) );
  AND2X2 AND2X2_3487 ( .A(round_ctr_rst_bF_buf51), .B(\block[8] ), .Y(w_mem_inst__abc_21378_n3204) );
  AND2X2 AND2X2_3488 ( .A(w_mem_inst__abc_21378_n3156_bF_buf1), .B(w_mem_inst_w_mem_15__8_), .Y(w_mem_inst__abc_21378_n3205) );
  AND2X2 AND2X2_3489 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf55), .B(w_mem_inst__abc_21378_n3206_1), .Y(w_mem_inst__abc_21378_n3207_1) );
  AND2X2 AND2X2_349 ( .A(_abc_15724_n1401), .B(_abc_15724_n1398), .Y(_abc_15724_n1402_1) );
  AND2X2 AND2X2_3490 ( .A(w_mem_inst__abc_21378_n2061), .B(w_mem_inst__abc_21378_n3152_bF_buf53), .Y(w_mem_inst__abc_21378_n3209) );
  AND2X2 AND2X2_3491 ( .A(round_ctr_rst_bF_buf50), .B(\block[9] ), .Y(w_mem_inst__abc_21378_n3210_1) );
  AND2X2 AND2X2_3492 ( .A(w_mem_inst__abc_21378_n3156_bF_buf0), .B(w_mem_inst_w_mem_15__9_), .Y(w_mem_inst__abc_21378_n3211_1) );
  AND2X2 AND2X2_3493 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf54), .B(w_mem_inst__abc_21378_n3212), .Y(w_mem_inst__abc_21378_n3213) );
  AND2X2 AND2X2_3494 ( .A(round_ctr_rst_bF_buf49), .B(\block[10] ), .Y(w_mem_inst__abc_21378_n3215_1) );
  AND2X2 AND2X2_3495 ( .A(w_mem_inst__abc_21378_n3156_bF_buf4), .B(w_mem_inst_w_mem_15__10_), .Y(w_mem_inst__abc_21378_n3216) );
  AND2X2 AND2X2_3496 ( .A(w_mem_inst__abc_21378_n3219_1), .B(w_mem_inst__abc_21378_n3218_1), .Y(w_mem_inst__0w_mem_15__31_0__10_) );
  AND2X2 AND2X2_3497 ( .A(round_ctr_rst_bF_buf48), .B(\block[11] ), .Y(w_mem_inst__abc_21378_n3221) );
  AND2X2 AND2X2_3498 ( .A(w_mem_inst__abc_21378_n3156_bF_buf3), .B(w_mem_inst_w_mem_15__11_), .Y(w_mem_inst__abc_21378_n3222_1) );
  AND2X2 AND2X2_3499 ( .A(w_mem_inst__abc_21378_n3225), .B(w_mem_inst__abc_21378_n3224), .Y(w_mem_inst__0w_mem_15__31_0__11_) );
  AND2X2 AND2X2_35 ( .A(_abc_15724_n762), .B(_abc_15724_n763), .Y(_abc_15724_n764) );
  AND2X2 AND2X2_350 ( .A(_abc_15724_n1404), .B(_abc_15724_n1397), .Y(_abc_15724_n1405) );
  AND2X2 AND2X2_3500 ( .A(round_ctr_rst_bF_buf47), .B(\block[12] ), .Y(w_mem_inst__abc_21378_n3227_1) );
  AND2X2 AND2X2_3501 ( .A(w_mem_inst__abc_21378_n3156_bF_buf2), .B(w_mem_inst_w_mem_15__12_), .Y(w_mem_inst__abc_21378_n3228) );
  AND2X2 AND2X2_3502 ( .A(w_mem_inst__abc_21378_n3231_1), .B(w_mem_inst__abc_21378_n3230_1), .Y(w_mem_inst__0w_mem_15__31_0__12_) );
  AND2X2 AND2X2_3503 ( .A(w_mem_inst__abc_21378_n2253), .B(w_mem_inst__abc_21378_n3152_bF_buf49), .Y(w_mem_inst__abc_21378_n3233) );
  AND2X2 AND2X2_3504 ( .A(round_ctr_rst_bF_buf46), .B(\block[13] ), .Y(w_mem_inst__abc_21378_n3234_1) );
  AND2X2 AND2X2_3505 ( .A(w_mem_inst__abc_21378_n3156_bF_buf1), .B(w_mem_inst_w_mem_15__13_), .Y(w_mem_inst__abc_21378_n3235_1) );
  AND2X2 AND2X2_3506 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf50), .B(w_mem_inst__abc_21378_n3236), .Y(w_mem_inst__abc_21378_n3237) );
  AND2X2 AND2X2_3507 ( .A(w_mem_inst__abc_21378_n2301), .B(w_mem_inst__abc_21378_n3152_bF_buf48), .Y(w_mem_inst__abc_21378_n3239_1) );
  AND2X2 AND2X2_3508 ( .A(round_ctr_rst_bF_buf45), .B(\block[14] ), .Y(w_mem_inst__abc_21378_n3240) );
  AND2X2 AND2X2_3509 ( .A(w_mem_inst__abc_21378_n3156_bF_buf0), .B(w_mem_inst_w_mem_15__14_), .Y(w_mem_inst__abc_21378_n3241) );
  AND2X2 AND2X2_351 ( .A(_abc_15724_n1383), .B(_abc_15724_n1394), .Y(_abc_15724_n1406) );
  AND2X2 AND2X2_3510 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf49), .B(w_mem_inst__abc_21378_n3242_1), .Y(w_mem_inst__abc_21378_n3243_1) );
  AND2X2 AND2X2_3511 ( .A(w_mem_inst__abc_21378_n2349), .B(w_mem_inst__abc_21378_n3152_bF_buf47), .Y(w_mem_inst__abc_21378_n3245) );
  AND2X2 AND2X2_3512 ( .A(round_ctr_rst_bF_buf44), .B(\block[15] ), .Y(w_mem_inst__abc_21378_n3246_1) );
  AND2X2 AND2X2_3513 ( .A(w_mem_inst__abc_21378_n3156_bF_buf4), .B(w_mem_inst_w_mem_15__15_), .Y(w_mem_inst__abc_21378_n3247_1) );
  AND2X2 AND2X2_3514 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf48), .B(w_mem_inst__abc_21378_n3248), .Y(w_mem_inst__abc_21378_n3249) );
  AND2X2 AND2X2_3515 ( .A(w_mem_inst__abc_21378_n2397), .B(w_mem_inst__abc_21378_n3152_bF_buf46), .Y(w_mem_inst__abc_21378_n3251_1) );
  AND2X2 AND2X2_3516 ( .A(round_ctr_rst_bF_buf43), .B(\block[16] ), .Y(w_mem_inst__abc_21378_n3252) );
  AND2X2 AND2X2_3517 ( .A(w_mem_inst__abc_21378_n3156_bF_buf3), .B(w_mem_inst_w_mem_15__16_), .Y(w_mem_inst__abc_21378_n3253) );
  AND2X2 AND2X2_3518 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf47), .B(w_mem_inst__abc_21378_n3254_1), .Y(w_mem_inst__abc_21378_n3255_1) );
  AND2X2 AND2X2_3519 ( .A(w_mem_inst__abc_21378_n2445), .B(w_mem_inst__abc_21378_n3152_bF_buf45), .Y(w_mem_inst__abc_21378_n3257) );
  AND2X2 AND2X2_352 ( .A(_abc_15724_n1394), .B(_abc_15724_n1381), .Y(_abc_15724_n1409) );
  AND2X2 AND2X2_3520 ( .A(round_ctr_rst_bF_buf42), .B(\block[17] ), .Y(w_mem_inst__abc_21378_n3258_1) );
  AND2X2 AND2X2_3521 ( .A(w_mem_inst__abc_21378_n3156_bF_buf2), .B(w_mem_inst_w_mem_15__17_), .Y(w_mem_inst__abc_21378_n3259_1) );
  AND2X2 AND2X2_3522 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf46), .B(w_mem_inst__abc_21378_n3260), .Y(w_mem_inst__abc_21378_n3261) );
  AND2X2 AND2X2_3523 ( .A(round_ctr_rst_bF_buf41), .B(\block[18] ), .Y(w_mem_inst__abc_21378_n3263_1) );
  AND2X2 AND2X2_3524 ( .A(w_mem_inst__abc_21378_n3156_bF_buf1), .B(w_mem_inst_w_mem_15__18_), .Y(w_mem_inst__abc_21378_n3264) );
  AND2X2 AND2X2_3525 ( .A(w_mem_inst__abc_21378_n3267_1), .B(w_mem_inst__abc_21378_n3266_1), .Y(w_mem_inst__0w_mem_15__31_0__18_) );
  AND2X2 AND2X2_3526 ( .A(w_mem_inst__abc_21378_n2541), .B(w_mem_inst__abc_21378_n3152_bF_buf43), .Y(w_mem_inst__abc_21378_n3269) );
  AND2X2 AND2X2_3527 ( .A(round_ctr_rst_bF_buf40), .B(\block[19] ), .Y(w_mem_inst__abc_21378_n3270_1) );
  AND2X2 AND2X2_3528 ( .A(w_mem_inst__abc_21378_n3156_bF_buf0), .B(w_mem_inst_w_mem_15__19_), .Y(w_mem_inst__abc_21378_n3271_1) );
  AND2X2 AND2X2_3529 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf44), .B(w_mem_inst__abc_21378_n3272), .Y(w_mem_inst__abc_21378_n3273) );
  AND2X2 AND2X2_353 ( .A(_abc_15724_n1410), .B(digest_update_bF_buf11), .Y(_abc_15724_n1411) );
  AND2X2 AND2X2_3530 ( .A(w_mem_inst__abc_21378_n2589), .B(w_mem_inst__abc_21378_n3152_bF_buf42), .Y(w_mem_inst__abc_21378_n3275_1) );
  AND2X2 AND2X2_3531 ( .A(round_ctr_rst_bF_buf39), .B(\block[20] ), .Y(w_mem_inst__abc_21378_n3276) );
  AND2X2 AND2X2_3532 ( .A(w_mem_inst__abc_21378_n3156_bF_buf4), .B(w_mem_inst_w_mem_15__20_), .Y(w_mem_inst__abc_21378_n3277) );
  AND2X2 AND2X2_3533 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf43), .B(w_mem_inst__abc_21378_n3278_1), .Y(w_mem_inst__abc_21378_n3279_1) );
  AND2X2 AND2X2_3534 ( .A(w_mem_inst__abc_21378_n2637), .B(w_mem_inst__abc_21378_n3152_bF_buf41), .Y(w_mem_inst__abc_21378_n3281) );
  AND2X2 AND2X2_3535 ( .A(round_ctr_rst_bF_buf38), .B(\block[21] ), .Y(w_mem_inst__abc_21378_n3282_1) );
  AND2X2 AND2X2_3536 ( .A(w_mem_inst__abc_21378_n3156_bF_buf3), .B(w_mem_inst_w_mem_15__21_), .Y(w_mem_inst__abc_21378_n3283_1) );
  AND2X2 AND2X2_3537 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf42), .B(w_mem_inst__abc_21378_n3284), .Y(w_mem_inst__abc_21378_n3285) );
  AND2X2 AND2X2_3538 ( .A(w_mem_inst__abc_21378_n2685), .B(w_mem_inst__abc_21378_n3152_bF_buf40), .Y(w_mem_inst__abc_21378_n3287_1) );
  AND2X2 AND2X2_3539 ( .A(round_ctr_rst_bF_buf37), .B(\block[22] ), .Y(w_mem_inst__abc_21378_n3288) );
  AND2X2 AND2X2_354 ( .A(_abc_15724_n1408), .B(_abc_15724_n1411), .Y(_abc_15724_n1412) );
  AND2X2 AND2X2_3540 ( .A(w_mem_inst__abc_21378_n3156_bF_buf2), .B(w_mem_inst_w_mem_15__22_), .Y(w_mem_inst__abc_21378_n3289) );
  AND2X2 AND2X2_3541 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf41), .B(w_mem_inst__abc_21378_n3290_1), .Y(w_mem_inst__abc_21378_n3291_1) );
  AND2X2 AND2X2_3542 ( .A(w_mem_inst__abc_21378_n2733), .B(w_mem_inst__abc_21378_n3152_bF_buf39), .Y(w_mem_inst__abc_21378_n3293) );
  AND2X2 AND2X2_3543 ( .A(round_ctr_rst_bF_buf36), .B(\block[23] ), .Y(w_mem_inst__abc_21378_n3294_1) );
  AND2X2 AND2X2_3544 ( .A(w_mem_inst__abc_21378_n3156_bF_buf1), .B(w_mem_inst_w_mem_15__23_), .Y(w_mem_inst__abc_21378_n3295_1) );
  AND2X2 AND2X2_3545 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf40), .B(w_mem_inst__abc_21378_n3296), .Y(w_mem_inst__abc_21378_n3297) );
  AND2X2 AND2X2_3546 ( .A(w_mem_inst__abc_21378_n2781), .B(w_mem_inst__abc_21378_n3152_bF_buf38), .Y(w_mem_inst__abc_21378_n3299_1) );
  AND2X2 AND2X2_3547 ( .A(round_ctr_rst_bF_buf35), .B(\block[24] ), .Y(w_mem_inst__abc_21378_n3300) );
  AND2X2 AND2X2_3548 ( .A(w_mem_inst__abc_21378_n3156_bF_buf0), .B(w_mem_inst_w_mem_15__24_), .Y(w_mem_inst__abc_21378_n3301) );
  AND2X2 AND2X2_3549 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf39), .B(w_mem_inst__abc_21378_n3302_1), .Y(w_mem_inst__abc_21378_n3303_1) );
  AND2X2 AND2X2_355 ( .A(_abc_15724_n1412), .B(_abc_15724_n1396), .Y(_abc_15724_n1413_1) );
  AND2X2 AND2X2_3550 ( .A(round_ctr_rst_bF_buf34), .B(\block[25] ), .Y(w_mem_inst__abc_21378_n3305) );
  AND2X2 AND2X2_3551 ( .A(w_mem_inst__abc_21378_n3156_bF_buf4), .B(w_mem_inst_w_mem_15__25_), .Y(w_mem_inst__abc_21378_n3306_1) );
  AND2X2 AND2X2_3552 ( .A(w_mem_inst__abc_21378_n3309), .B(w_mem_inst__abc_21378_n3308), .Y(w_mem_inst__0w_mem_15__31_0__25_) );
  AND2X2 AND2X2_3553 ( .A(round_ctr_rst_bF_buf33), .B(\block[26] ), .Y(w_mem_inst__abc_21378_n3311_1) );
  AND2X2 AND2X2_3554 ( .A(w_mem_inst__abc_21378_n3156_bF_buf3), .B(w_mem_inst_w_mem_15__26_), .Y(w_mem_inst__abc_21378_n3312) );
  AND2X2 AND2X2_3555 ( .A(w_mem_inst__abc_21378_n3315_1), .B(w_mem_inst__abc_21378_n3314_1), .Y(w_mem_inst__0w_mem_15__31_0__26_) );
  AND2X2 AND2X2_3556 ( .A(round_ctr_rst_bF_buf32), .B(\block[27] ), .Y(w_mem_inst__abc_21378_n3317) );
  AND2X2 AND2X2_3557 ( .A(w_mem_inst__abc_21378_n3156_bF_buf2), .B(w_mem_inst_w_mem_15__27_), .Y(w_mem_inst__abc_21378_n3318_1) );
  AND2X2 AND2X2_3558 ( .A(w_mem_inst__abc_21378_n3321), .B(w_mem_inst__abc_21378_n3320), .Y(w_mem_inst__0w_mem_15__31_0__27_) );
  AND2X2 AND2X2_3559 ( .A(round_ctr_rst_bF_buf31), .B(\block[28] ), .Y(w_mem_inst__abc_21378_n3323_1) );
  AND2X2 AND2X2_356 ( .A(_abc_15724_n907_1_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_58_), .Y(_abc_15724_n1415) );
  AND2X2 AND2X2_3560 ( .A(w_mem_inst__abc_21378_n3156_bF_buf1), .B(w_mem_inst_w_mem_15__28_), .Y(w_mem_inst__abc_21378_n3324) );
  AND2X2 AND2X2_3561 ( .A(w_mem_inst__abc_21378_n3327_1), .B(w_mem_inst__abc_21378_n3326_1), .Y(w_mem_inst__0w_mem_15__31_0__28_) );
  AND2X2 AND2X2_3562 ( .A(w_mem_inst__abc_21378_n3021), .B(w_mem_inst__abc_21378_n3152_bF_buf33), .Y(w_mem_inst__abc_21378_n3329) );
  AND2X2 AND2X2_3563 ( .A(round_ctr_rst_bF_buf30), .B(\block[29] ), .Y(w_mem_inst__abc_21378_n3330_1) );
  AND2X2 AND2X2_3564 ( .A(w_mem_inst__abc_21378_n3156_bF_buf0), .B(w_mem_inst_w_mem_15__29_), .Y(w_mem_inst__abc_21378_n3331_1) );
  AND2X2 AND2X2_3565 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf34), .B(w_mem_inst__abc_21378_n3332), .Y(w_mem_inst__abc_21378_n3333) );
  AND2X2 AND2X2_3566 ( .A(w_mem_inst__abc_21378_n3069), .B(w_mem_inst__abc_21378_n3152_bF_buf32), .Y(w_mem_inst__abc_21378_n3335_1) );
  AND2X2 AND2X2_3567 ( .A(round_ctr_rst_bF_buf29), .B(\block[30] ), .Y(w_mem_inst__abc_21378_n3336) );
  AND2X2 AND2X2_3568 ( .A(w_mem_inst__abc_21378_n3156_bF_buf4), .B(w_mem_inst_w_mem_15__30_), .Y(w_mem_inst__abc_21378_n3337) );
  AND2X2 AND2X2_3569 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf33), .B(w_mem_inst__abc_21378_n3338_1), .Y(w_mem_inst__abc_21378_n3339_1) );
  AND2X2 AND2X2_357 ( .A(_abc_15724_n1379_1), .B(_abc_15724_n1406), .Y(_abc_15724_n1416_1) );
  AND2X2 AND2X2_3570 ( .A(w_mem_inst__abc_21378_n3117), .B(w_mem_inst__abc_21378_n3152_bF_buf31), .Y(w_mem_inst__abc_21378_n3341) );
  AND2X2 AND2X2_3571 ( .A(round_ctr_rst_bF_buf28), .B(\block[31] ), .Y(w_mem_inst__abc_21378_n3342_1) );
  AND2X2 AND2X2_3572 ( .A(w_mem_inst__abc_21378_n3156_bF_buf3), .B(w_mem_inst_w_mem_15__31_), .Y(w_mem_inst__abc_21378_n3343_1) );
  AND2X2 AND2X2_3573 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf32), .B(w_mem_inst__abc_21378_n3344), .Y(w_mem_inst__abc_21378_n3345) );
  AND2X2 AND2X2_3574 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf31), .B(w_mem_inst__abc_21378_n3156_bF_buf2), .Y(w_mem_inst__abc_21378_n3347_1) );
  AND2X2 AND2X2_3575 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf60), .B(w_mem_inst_w_mem_14__0_), .Y(w_mem_inst__abc_21378_n3348) );
  AND2X2 AND2X2_3576 ( .A(w_mem_inst__abc_21378_n3152_bF_buf30), .B(w_mem_inst_w_mem_15__0_), .Y(w_mem_inst__abc_21378_n3349) );
  AND2X2 AND2X2_3577 ( .A(round_ctr_rst_bF_buf27), .B(\block[32] ), .Y(w_mem_inst__abc_21378_n3350_1) );
  AND2X2 AND2X2_3578 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf30), .B(w_mem_inst__abc_21378_n3350_1), .Y(w_mem_inst__abc_21378_n3351_1) );
  AND2X2 AND2X2_3579 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf59), .B(w_mem_inst_w_mem_14__1_), .Y(w_mem_inst__abc_21378_n3354_1) );
  AND2X2 AND2X2_358 ( .A(_abc_15724_n1410), .B(_abc_15724_n1393_1), .Y(_abc_15724_n1417) );
  AND2X2 AND2X2_3580 ( .A(w_mem_inst__abc_21378_n3152_bF_buf29), .B(w_mem_inst_w_mem_15__1_), .Y(w_mem_inst__abc_21378_n3355_1) );
  AND2X2 AND2X2_3581 ( .A(round_ctr_rst_bF_buf26), .B(\block[33] ), .Y(w_mem_inst__abc_21378_n3356) );
  AND2X2 AND2X2_3582 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf29), .B(w_mem_inst__abc_21378_n3356), .Y(w_mem_inst__abc_21378_n3357) );
  AND2X2 AND2X2_3583 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf58), .B(w_mem_inst_w_mem_14__2_), .Y(w_mem_inst__abc_21378_n3360) );
  AND2X2 AND2X2_3584 ( .A(w_mem_inst__abc_21378_n3152_bF_buf28), .B(w_mem_inst_w_mem_15__2_), .Y(w_mem_inst__abc_21378_n3361) );
  AND2X2 AND2X2_3585 ( .A(round_ctr_rst_bF_buf25), .B(\block[34] ), .Y(w_mem_inst__abc_21378_n3362_1) );
  AND2X2 AND2X2_3586 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf28), .B(w_mem_inst__abc_21378_n3362_1), .Y(w_mem_inst__abc_21378_n3363_1) );
  AND2X2 AND2X2_3587 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf57), .B(w_mem_inst_w_mem_14__3_), .Y(w_mem_inst__abc_21378_n3366_1) );
  AND2X2 AND2X2_3588 ( .A(w_mem_inst__abc_21378_n3152_bF_buf27), .B(w_mem_inst_w_mem_15__3_), .Y(w_mem_inst__abc_21378_n3367_1) );
  AND2X2 AND2X2_3589 ( .A(round_ctr_rst_bF_buf24), .B(\block[35] ), .Y(w_mem_inst__abc_21378_n3368) );
  AND2X2 AND2X2_359 ( .A(_auto_iopadmap_cc_313_execute_26059_58_), .B(d_reg_26_), .Y(_abc_15724_n1421) );
  AND2X2 AND2X2_3590 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf27), .B(w_mem_inst__abc_21378_n3368), .Y(w_mem_inst__abc_21378_n3369) );
  AND2X2 AND2X2_3591 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf56), .B(w_mem_inst_w_mem_14__4_), .Y(w_mem_inst__abc_21378_n3372) );
  AND2X2 AND2X2_3592 ( .A(w_mem_inst__abc_21378_n3152_bF_buf26), .B(w_mem_inst_w_mem_15__4_), .Y(w_mem_inst__abc_21378_n3373) );
  AND2X2 AND2X2_3593 ( .A(round_ctr_rst_bF_buf23), .B(\block[36] ), .Y(w_mem_inst__abc_21378_n3374_1) );
  AND2X2 AND2X2_3594 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf26), .B(w_mem_inst__abc_21378_n3374_1), .Y(w_mem_inst__abc_21378_n3375_1) );
  AND2X2 AND2X2_3595 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf55), .B(w_mem_inst_w_mem_14__5_), .Y(w_mem_inst__abc_21378_n3378_1) );
  AND2X2 AND2X2_3596 ( .A(w_mem_inst__abc_21378_n3152_bF_buf25), .B(w_mem_inst_w_mem_15__5_), .Y(w_mem_inst__abc_21378_n3379_1) );
  AND2X2 AND2X2_3597 ( .A(round_ctr_rst_bF_buf22), .B(\block[37] ), .Y(w_mem_inst__abc_21378_n3380) );
  AND2X2 AND2X2_3598 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf25), .B(w_mem_inst__abc_21378_n3380), .Y(w_mem_inst__abc_21378_n3381) );
  AND2X2 AND2X2_3599 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf54), .B(w_mem_inst_w_mem_14__6_), .Y(w_mem_inst__abc_21378_n3384) );
  AND2X2 AND2X2_36 ( .A(_abc_15724_n761), .B(_abc_15724_n764), .Y(_abc_15724_n765) );
  AND2X2 AND2X2_360 ( .A(_abc_15724_n1422_1), .B(_abc_15724_n1420), .Y(_abc_15724_n1423_1) );
  AND2X2 AND2X2_3600 ( .A(w_mem_inst__abc_21378_n3152_bF_buf24), .B(w_mem_inst_w_mem_15__6_), .Y(w_mem_inst__abc_21378_n3385) );
  AND2X2 AND2X2_3601 ( .A(round_ctr_rst_bF_buf21), .B(\block[38] ), .Y(w_mem_inst__abc_21378_n3386_1) );
  AND2X2 AND2X2_3602 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf24), .B(w_mem_inst__abc_21378_n3386_1), .Y(w_mem_inst__abc_21378_n3387_1) );
  AND2X2 AND2X2_3603 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf53), .B(w_mem_inst_w_mem_14__7_), .Y(w_mem_inst__abc_21378_n3390_1) );
  AND2X2 AND2X2_3604 ( .A(w_mem_inst__abc_21378_n3152_bF_buf23), .B(w_mem_inst_w_mem_15__7_), .Y(w_mem_inst__abc_21378_n3391_1) );
  AND2X2 AND2X2_3605 ( .A(round_ctr_rst_bF_buf20), .B(\block[39] ), .Y(w_mem_inst__abc_21378_n3392) );
  AND2X2 AND2X2_3606 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf23), .B(w_mem_inst__abc_21378_n3392), .Y(w_mem_inst__abc_21378_n3393) );
  AND2X2 AND2X2_3607 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf52), .B(w_mem_inst_w_mem_14__8_), .Y(w_mem_inst__abc_21378_n3396) );
  AND2X2 AND2X2_3608 ( .A(w_mem_inst__abc_21378_n3152_bF_buf22), .B(w_mem_inst_w_mem_15__8_), .Y(w_mem_inst__abc_21378_n3397) );
  AND2X2 AND2X2_3609 ( .A(round_ctr_rst_bF_buf19), .B(\block[40] ), .Y(w_mem_inst__abc_21378_n3398_1) );
  AND2X2 AND2X2_361 ( .A(_abc_15724_n1419), .B(_abc_15724_n1423_1), .Y(_abc_15724_n1425) );
  AND2X2 AND2X2_3610 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf22), .B(w_mem_inst__abc_21378_n3398_1), .Y(w_mem_inst__abc_21378_n3399_1) );
  AND2X2 AND2X2_3611 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf51), .B(w_mem_inst_w_mem_14__9_), .Y(w_mem_inst__abc_21378_n3402_1) );
  AND2X2 AND2X2_3612 ( .A(w_mem_inst__abc_21378_n3152_bF_buf21), .B(w_mem_inst_w_mem_15__9_), .Y(w_mem_inst__abc_21378_n3403_1) );
  AND2X2 AND2X2_3613 ( .A(round_ctr_rst_bF_buf18), .B(\block[41] ), .Y(w_mem_inst__abc_21378_n3404) );
  AND2X2 AND2X2_3614 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf21), .B(w_mem_inst__abc_21378_n3404), .Y(w_mem_inst__abc_21378_n3405) );
  AND2X2 AND2X2_3615 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf50), .B(w_mem_inst_w_mem_14__10_), .Y(w_mem_inst__abc_21378_n3408) );
  AND2X2 AND2X2_3616 ( .A(w_mem_inst__abc_21378_n3152_bF_buf20), .B(w_mem_inst_w_mem_15__10_), .Y(w_mem_inst__abc_21378_n3409) );
  AND2X2 AND2X2_3617 ( .A(round_ctr_rst_bF_buf17), .B(\block[42] ), .Y(w_mem_inst__abc_21378_n3410_1) );
  AND2X2 AND2X2_3618 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf20), .B(w_mem_inst__abc_21378_n3410_1), .Y(w_mem_inst__abc_21378_n3411_1) );
  AND2X2 AND2X2_3619 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf49), .B(w_mem_inst_w_mem_14__11_), .Y(w_mem_inst__abc_21378_n3414_1) );
  AND2X2 AND2X2_362 ( .A(_abc_15724_n1426), .B(_abc_15724_n1424_1), .Y(_abc_15724_n1427) );
  AND2X2 AND2X2_3620 ( .A(w_mem_inst__abc_21378_n3152_bF_buf19), .B(w_mem_inst_w_mem_15__11_), .Y(w_mem_inst__abc_21378_n3415_1) );
  AND2X2 AND2X2_3621 ( .A(round_ctr_rst_bF_buf16), .B(\block[43] ), .Y(w_mem_inst__abc_21378_n3416) );
  AND2X2 AND2X2_3622 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf19), .B(w_mem_inst__abc_21378_n3416), .Y(w_mem_inst__abc_21378_n3417) );
  AND2X2 AND2X2_3623 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf48), .B(w_mem_inst_w_mem_14__12_), .Y(w_mem_inst__abc_21378_n3420) );
  AND2X2 AND2X2_3624 ( .A(w_mem_inst__abc_21378_n3152_bF_buf18), .B(w_mem_inst_w_mem_15__12_), .Y(w_mem_inst__abc_21378_n3421) );
  AND2X2 AND2X2_3625 ( .A(round_ctr_rst_bF_buf15), .B(\block[44] ), .Y(w_mem_inst__abc_21378_n3422_1) );
  AND2X2 AND2X2_3626 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf18), .B(w_mem_inst__abc_21378_n3422_1), .Y(w_mem_inst__abc_21378_n3423_1) );
  AND2X2 AND2X2_3627 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf47), .B(w_mem_inst_w_mem_14__13_), .Y(w_mem_inst__abc_21378_n3426_1) );
  AND2X2 AND2X2_3628 ( .A(w_mem_inst__abc_21378_n3152_bF_buf17), .B(w_mem_inst_w_mem_15__13_), .Y(w_mem_inst__abc_21378_n3427_1) );
  AND2X2 AND2X2_3629 ( .A(round_ctr_rst_bF_buf14), .B(\block[45] ), .Y(w_mem_inst__abc_21378_n3428) );
  AND2X2 AND2X2_363 ( .A(_abc_15724_n1427), .B(digest_update_bF_buf10), .Y(_abc_15724_n1428) );
  AND2X2 AND2X2_3630 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf17), .B(w_mem_inst__abc_21378_n3428), .Y(w_mem_inst__abc_21378_n3429) );
  AND2X2 AND2X2_3631 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf46), .B(w_mem_inst_w_mem_14__14_), .Y(w_mem_inst__abc_21378_n3432) );
  AND2X2 AND2X2_3632 ( .A(w_mem_inst__abc_21378_n3152_bF_buf16), .B(w_mem_inst_w_mem_15__14_), .Y(w_mem_inst__abc_21378_n3433) );
  AND2X2 AND2X2_3633 ( .A(round_ctr_rst_bF_buf13), .B(\block[46] ), .Y(w_mem_inst__abc_21378_n3434_1) );
  AND2X2 AND2X2_3634 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf16), .B(w_mem_inst__abc_21378_n3434_1), .Y(w_mem_inst__abc_21378_n3435_1) );
  AND2X2 AND2X2_3635 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf45), .B(w_mem_inst_w_mem_14__15_), .Y(w_mem_inst__abc_21378_n3438_1) );
  AND2X2 AND2X2_3636 ( .A(w_mem_inst__abc_21378_n3152_bF_buf15), .B(w_mem_inst_w_mem_15__15_), .Y(w_mem_inst__abc_21378_n3439_1) );
  AND2X2 AND2X2_3637 ( .A(round_ctr_rst_bF_buf12), .B(\block[47] ), .Y(w_mem_inst__abc_21378_n3440) );
  AND2X2 AND2X2_3638 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf15), .B(w_mem_inst__abc_21378_n3440), .Y(w_mem_inst__abc_21378_n3441) );
  AND2X2 AND2X2_3639 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf44), .B(w_mem_inst_w_mem_14__16_), .Y(w_mem_inst__abc_21378_n3444) );
  AND2X2 AND2X2_364 ( .A(_abc_15724_n907_1_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_59_), .Y(_abc_15724_n1430) );
  AND2X2 AND2X2_3640 ( .A(w_mem_inst__abc_21378_n3152_bF_buf14), .B(w_mem_inst_w_mem_15__16_), .Y(w_mem_inst__abc_21378_n3445) );
  AND2X2 AND2X2_3641 ( .A(round_ctr_rst_bF_buf11), .B(\block[48] ), .Y(w_mem_inst__abc_21378_n3446_1) );
  AND2X2 AND2X2_3642 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf14), .B(w_mem_inst__abc_21378_n3446_1), .Y(w_mem_inst__abc_21378_n3447_1) );
  AND2X2 AND2X2_3643 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf43), .B(w_mem_inst_w_mem_14__17_), .Y(w_mem_inst__abc_21378_n3450_1) );
  AND2X2 AND2X2_3644 ( .A(w_mem_inst__abc_21378_n3152_bF_buf13), .B(w_mem_inst_w_mem_15__17_), .Y(w_mem_inst__abc_21378_n3451_1) );
  AND2X2 AND2X2_3645 ( .A(round_ctr_rst_bF_buf10), .B(\block[49] ), .Y(w_mem_inst__abc_21378_n3452) );
  AND2X2 AND2X2_3646 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf13), .B(w_mem_inst__abc_21378_n3452), .Y(w_mem_inst__abc_21378_n3453) );
  AND2X2 AND2X2_3647 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf42), .B(w_mem_inst_w_mem_14__18_), .Y(w_mem_inst__abc_21378_n3456) );
  AND2X2 AND2X2_3648 ( .A(w_mem_inst__abc_21378_n3152_bF_buf12), .B(w_mem_inst_w_mem_15__18_), .Y(w_mem_inst__abc_21378_n3457) );
  AND2X2 AND2X2_3649 ( .A(round_ctr_rst_bF_buf9), .B(\block[50] ), .Y(w_mem_inst__abc_21378_n3458_1) );
  AND2X2 AND2X2_365 ( .A(_auto_iopadmap_cc_313_execute_26059_59_), .B(d_reg_27_), .Y(_abc_15724_n1432) );
  AND2X2 AND2X2_3650 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf12), .B(w_mem_inst__abc_21378_n3458_1), .Y(w_mem_inst__abc_21378_n3459_1) );
  AND2X2 AND2X2_3651 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf41), .B(w_mem_inst_w_mem_14__19_), .Y(w_mem_inst__abc_21378_n3462_1) );
  AND2X2 AND2X2_3652 ( .A(w_mem_inst__abc_21378_n3152_bF_buf11), .B(w_mem_inst_w_mem_15__19_), .Y(w_mem_inst__abc_21378_n3463_1) );
  AND2X2 AND2X2_3653 ( .A(round_ctr_rst_bF_buf8), .B(\block[51] ), .Y(w_mem_inst__abc_21378_n3464) );
  AND2X2 AND2X2_3654 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf11), .B(w_mem_inst__abc_21378_n3464), .Y(w_mem_inst__abc_21378_n3465) );
  AND2X2 AND2X2_3655 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf40), .B(w_mem_inst_w_mem_14__20_), .Y(w_mem_inst__abc_21378_n3468) );
  AND2X2 AND2X2_3656 ( .A(w_mem_inst__abc_21378_n3152_bF_buf10), .B(w_mem_inst_w_mem_15__20_), .Y(w_mem_inst__abc_21378_n3469) );
  AND2X2 AND2X2_3657 ( .A(round_ctr_rst_bF_buf7), .B(\block[52] ), .Y(w_mem_inst__abc_21378_n3470_1) );
  AND2X2 AND2X2_3658 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf10), .B(w_mem_inst__abc_21378_n3470_1), .Y(w_mem_inst__abc_21378_n3471_1) );
  AND2X2 AND2X2_3659 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf39), .B(w_mem_inst_w_mem_14__21_), .Y(w_mem_inst__abc_21378_n3474_1) );
  AND2X2 AND2X2_366 ( .A(_abc_15724_n1433), .B(_abc_15724_n1431), .Y(_abc_15724_n1434) );
  AND2X2 AND2X2_3660 ( .A(w_mem_inst__abc_21378_n3152_bF_buf9), .B(w_mem_inst_w_mem_15__21_), .Y(w_mem_inst__abc_21378_n3475_1) );
  AND2X2 AND2X2_3661 ( .A(round_ctr_rst_bF_buf6), .B(\block[53] ), .Y(w_mem_inst__abc_21378_n3476) );
  AND2X2 AND2X2_3662 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf9), .B(w_mem_inst__abc_21378_n3476), .Y(w_mem_inst__abc_21378_n3477) );
  AND2X2 AND2X2_3663 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf38), .B(w_mem_inst_w_mem_14__22_), .Y(w_mem_inst__abc_21378_n3480) );
  AND2X2 AND2X2_3664 ( .A(w_mem_inst__abc_21378_n3152_bF_buf8), .B(w_mem_inst_w_mem_15__22_), .Y(w_mem_inst__abc_21378_n3481) );
  AND2X2 AND2X2_3665 ( .A(round_ctr_rst_bF_buf5), .B(\block[54] ), .Y(w_mem_inst__abc_21378_n3482_1) );
  AND2X2 AND2X2_3666 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf8), .B(w_mem_inst__abc_21378_n3482_1), .Y(w_mem_inst__abc_21378_n3483_1) );
  AND2X2 AND2X2_3667 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf37), .B(w_mem_inst_w_mem_14__23_), .Y(w_mem_inst__abc_21378_n3486_1) );
  AND2X2 AND2X2_3668 ( .A(w_mem_inst__abc_21378_n3152_bF_buf7), .B(w_mem_inst_w_mem_15__23_), .Y(w_mem_inst__abc_21378_n3487_1) );
  AND2X2 AND2X2_3669 ( .A(round_ctr_rst_bF_buf4), .B(\block[55] ), .Y(w_mem_inst__abc_21378_n3488) );
  AND2X2 AND2X2_367 ( .A(_abc_15724_n1408), .B(_abc_15724_n1417), .Y(_abc_15724_n1437) );
  AND2X2 AND2X2_3670 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf7), .B(w_mem_inst__abc_21378_n3488), .Y(w_mem_inst__abc_21378_n3489) );
  AND2X2 AND2X2_3671 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf36), .B(w_mem_inst_w_mem_14__24_), .Y(w_mem_inst__abc_21378_n3492) );
  AND2X2 AND2X2_3672 ( .A(w_mem_inst__abc_21378_n3152_bF_buf6), .B(w_mem_inst_w_mem_15__24_), .Y(w_mem_inst__abc_21378_n3493) );
  AND2X2 AND2X2_3673 ( .A(round_ctr_rst_bF_buf3), .B(\block[56] ), .Y(w_mem_inst__abc_21378_n3494_1) );
  AND2X2 AND2X2_3674 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf6), .B(w_mem_inst__abc_21378_n3494_1), .Y(w_mem_inst__abc_21378_n3495_1) );
  AND2X2 AND2X2_3675 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf35), .B(w_mem_inst_w_mem_14__25_), .Y(w_mem_inst__abc_21378_n3498_1) );
  AND2X2 AND2X2_3676 ( .A(w_mem_inst__abc_21378_n3152_bF_buf5), .B(w_mem_inst_w_mem_15__25_), .Y(w_mem_inst__abc_21378_n3499_1) );
  AND2X2 AND2X2_3677 ( .A(round_ctr_rst_bF_buf2), .B(\block[57] ), .Y(w_mem_inst__abc_21378_n3500) );
  AND2X2 AND2X2_3678 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf5), .B(w_mem_inst__abc_21378_n3500), .Y(w_mem_inst__abc_21378_n3501) );
  AND2X2 AND2X2_3679 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf34), .B(w_mem_inst_w_mem_14__26_), .Y(w_mem_inst__abc_21378_n3504) );
  AND2X2 AND2X2_368 ( .A(_abc_15724_n1423_1), .B(_abc_15724_n1434), .Y(_abc_15724_n1438_1) );
  AND2X2 AND2X2_3680 ( .A(w_mem_inst__abc_21378_n3152_bF_buf4), .B(w_mem_inst_w_mem_15__26_), .Y(w_mem_inst__abc_21378_n3505) );
  AND2X2 AND2X2_3681 ( .A(round_ctr_rst_bF_buf1), .B(\block[58] ), .Y(w_mem_inst__abc_21378_n3506_1) );
  AND2X2 AND2X2_3682 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf4), .B(w_mem_inst__abc_21378_n3506_1), .Y(w_mem_inst__abc_21378_n3507_1) );
  AND2X2 AND2X2_3683 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf33), .B(w_mem_inst_w_mem_14__27_), .Y(w_mem_inst__abc_21378_n3510_1) );
  AND2X2 AND2X2_3684 ( .A(w_mem_inst__abc_21378_n3152_bF_buf3), .B(w_mem_inst_w_mem_15__27_), .Y(w_mem_inst__abc_21378_n3511_1) );
  AND2X2 AND2X2_3685 ( .A(round_ctr_rst_bF_buf0), .B(\block[59] ), .Y(w_mem_inst__abc_21378_n3512) );
  AND2X2 AND2X2_3686 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf3), .B(w_mem_inst__abc_21378_n3512), .Y(w_mem_inst__abc_21378_n3513) );
  AND2X2 AND2X2_3687 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf32), .B(w_mem_inst_w_mem_14__28_), .Y(w_mem_inst__abc_21378_n3516) );
  AND2X2 AND2X2_3688 ( .A(w_mem_inst__abc_21378_n3152_bF_buf2), .B(w_mem_inst_w_mem_15__28_), .Y(w_mem_inst__abc_21378_n3517) );
  AND2X2 AND2X2_3689 ( .A(round_ctr_rst_bF_buf63), .B(\block[60] ), .Y(w_mem_inst__abc_21378_n3518_1) );
  AND2X2 AND2X2_369 ( .A(_abc_15724_n1434), .B(_abc_15724_n1421), .Y(_abc_15724_n1441) );
  AND2X2 AND2X2_3690 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf2), .B(w_mem_inst__abc_21378_n3518_1), .Y(w_mem_inst__abc_21378_n3519_1) );
  AND2X2 AND2X2_3691 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf31), .B(w_mem_inst_w_mem_14__29_), .Y(w_mem_inst__abc_21378_n3522_1) );
  AND2X2 AND2X2_3692 ( .A(w_mem_inst__abc_21378_n3152_bF_buf1), .B(w_mem_inst_w_mem_15__29_), .Y(w_mem_inst__abc_21378_n3523_1) );
  AND2X2 AND2X2_3693 ( .A(round_ctr_rst_bF_buf62), .B(\block[61] ), .Y(w_mem_inst__abc_21378_n3524) );
  AND2X2 AND2X2_3694 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf1), .B(w_mem_inst__abc_21378_n3524), .Y(w_mem_inst__abc_21378_n3525) );
  AND2X2 AND2X2_3695 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf30), .B(w_mem_inst_w_mem_14__30_), .Y(w_mem_inst__abc_21378_n3528) );
  AND2X2 AND2X2_3696 ( .A(w_mem_inst__abc_21378_n3152_bF_buf0), .B(w_mem_inst_w_mem_15__30_), .Y(w_mem_inst__abc_21378_n3529) );
  AND2X2 AND2X2_3697 ( .A(round_ctr_rst_bF_buf61), .B(\block[62] ), .Y(w_mem_inst__abc_21378_n3530_1) );
  AND2X2 AND2X2_3698 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf0), .B(w_mem_inst__abc_21378_n3530_1), .Y(w_mem_inst__abc_21378_n3531_1) );
  AND2X2 AND2X2_3699 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf29), .B(w_mem_inst_w_mem_14__31_), .Y(w_mem_inst__abc_21378_n3534_1) );
  AND2X2 AND2X2_37 ( .A(e_reg_9_), .B(_auto_iopadmap_cc_313_execute_26059_9_), .Y(_abc_15724_n766_1) );
  AND2X2 AND2X2_370 ( .A(_abc_15724_n1442), .B(digest_update_bF_buf9), .Y(_abc_15724_n1443) );
  AND2X2 AND2X2_3700 ( .A(w_mem_inst__abc_21378_n3152_bF_buf63), .B(w_mem_inst_w_mem_15__31_), .Y(w_mem_inst__abc_21378_n3535_1) );
  AND2X2 AND2X2_3701 ( .A(round_ctr_rst_bF_buf60), .B(\block[63] ), .Y(w_mem_inst__abc_21378_n3536) );
  AND2X2 AND2X2_3702 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf63), .B(w_mem_inst__abc_21378_n3536), .Y(w_mem_inst__abc_21378_n3537) );
  AND2X2 AND2X2_3703 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf28), .B(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_21378_n3540) );
  AND2X2 AND2X2_3704 ( .A(w_mem_inst__abc_21378_n3152_bF_buf62), .B(w_mem_inst_w_mem_14__0_), .Y(w_mem_inst__abc_21378_n3541) );
  AND2X2 AND2X2_3705 ( .A(round_ctr_rst_bF_buf59), .B(\block[64] ), .Y(w_mem_inst__abc_21378_n3542_1) );
  AND2X2 AND2X2_3706 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf62), .B(w_mem_inst__abc_21378_n3542_1), .Y(w_mem_inst__abc_21378_n3543_1) );
  AND2X2 AND2X2_3707 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf27), .B(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_21378_n3546_1) );
  AND2X2 AND2X2_3708 ( .A(w_mem_inst__abc_21378_n3152_bF_buf61), .B(w_mem_inst_w_mem_14__1_), .Y(w_mem_inst__abc_21378_n3547_1) );
  AND2X2 AND2X2_3709 ( .A(round_ctr_rst_bF_buf58), .B(\block[65] ), .Y(w_mem_inst__abc_21378_n3548) );
  AND2X2 AND2X2_371 ( .A(_abc_15724_n1440), .B(_abc_15724_n1443), .Y(_abc_15724_n1444_1) );
  AND2X2 AND2X2_3710 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf61), .B(w_mem_inst__abc_21378_n3548), .Y(w_mem_inst__abc_21378_n3549) );
  AND2X2 AND2X2_3711 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf26), .B(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_21378_n3552) );
  AND2X2 AND2X2_3712 ( .A(w_mem_inst__abc_21378_n3152_bF_buf60), .B(w_mem_inst_w_mem_14__2_), .Y(w_mem_inst__abc_21378_n3553) );
  AND2X2 AND2X2_3713 ( .A(round_ctr_rst_bF_buf57), .B(\block[66] ), .Y(w_mem_inst__abc_21378_n3554_1) );
  AND2X2 AND2X2_3714 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf60), .B(w_mem_inst__abc_21378_n3554_1), .Y(w_mem_inst__abc_21378_n3555_1) );
  AND2X2 AND2X2_3715 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf25), .B(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_21378_n3558_1) );
  AND2X2 AND2X2_3716 ( .A(w_mem_inst__abc_21378_n3152_bF_buf59), .B(w_mem_inst_w_mem_14__3_), .Y(w_mem_inst__abc_21378_n3559_1) );
  AND2X2 AND2X2_3717 ( .A(round_ctr_rst_bF_buf56), .B(\block[67] ), .Y(w_mem_inst__abc_21378_n3560) );
  AND2X2 AND2X2_3718 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf59), .B(w_mem_inst__abc_21378_n3560), .Y(w_mem_inst__abc_21378_n3561) );
  AND2X2 AND2X2_3719 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf24), .B(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_21378_n3564) );
  AND2X2 AND2X2_372 ( .A(_abc_15724_n1444_1), .B(_abc_15724_n1436_1), .Y(_abc_15724_n1445_1) );
  AND2X2 AND2X2_3720 ( .A(w_mem_inst__abc_21378_n3152_bF_buf58), .B(w_mem_inst_w_mem_14__4_), .Y(w_mem_inst__abc_21378_n3565) );
  AND2X2 AND2X2_3721 ( .A(round_ctr_rst_bF_buf55), .B(\block[68] ), .Y(w_mem_inst__abc_21378_n3566_1) );
  AND2X2 AND2X2_3722 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf58), .B(w_mem_inst__abc_21378_n3566_1), .Y(w_mem_inst__abc_21378_n3567_1) );
  AND2X2 AND2X2_3723 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf23), .B(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_21378_n3570_1) );
  AND2X2 AND2X2_3724 ( .A(w_mem_inst__abc_21378_n3152_bF_buf57), .B(w_mem_inst_w_mem_14__5_), .Y(w_mem_inst__abc_21378_n3571_1) );
  AND2X2 AND2X2_3725 ( .A(round_ctr_rst_bF_buf54), .B(\block[69] ), .Y(w_mem_inst__abc_21378_n3572) );
  AND2X2 AND2X2_3726 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf57), .B(w_mem_inst__abc_21378_n3572), .Y(w_mem_inst__abc_21378_n3573) );
  AND2X2 AND2X2_3727 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf22), .B(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_21378_n3576) );
  AND2X2 AND2X2_3728 ( .A(w_mem_inst__abc_21378_n3152_bF_buf56), .B(w_mem_inst_w_mem_14__6_), .Y(w_mem_inst__abc_21378_n3577) );
  AND2X2 AND2X2_3729 ( .A(round_ctr_rst_bF_buf53), .B(\block[70] ), .Y(w_mem_inst__abc_21378_n3578_1) );
  AND2X2 AND2X2_373 ( .A(_abc_15724_n1419), .B(_abc_15724_n1438_1), .Y(_abc_15724_n1447) );
  AND2X2 AND2X2_3730 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf56), .B(w_mem_inst__abc_21378_n3578_1), .Y(w_mem_inst__abc_21378_n3579_1) );
  AND2X2 AND2X2_3731 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf21), .B(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_21378_n3582_1) );
  AND2X2 AND2X2_3732 ( .A(w_mem_inst__abc_21378_n3152_bF_buf55), .B(w_mem_inst_w_mem_14__7_), .Y(w_mem_inst__abc_21378_n3583_1) );
  AND2X2 AND2X2_3733 ( .A(round_ctr_rst_bF_buf52), .B(\block[71] ), .Y(w_mem_inst__abc_21378_n3584) );
  AND2X2 AND2X2_3734 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf55), .B(w_mem_inst__abc_21378_n3584), .Y(w_mem_inst__abc_21378_n3585) );
  AND2X2 AND2X2_3735 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf20), .B(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_21378_n3588) );
  AND2X2 AND2X2_3736 ( .A(w_mem_inst__abc_21378_n3152_bF_buf54), .B(w_mem_inst_w_mem_14__8_), .Y(w_mem_inst__abc_21378_n3589) );
  AND2X2 AND2X2_3737 ( .A(round_ctr_rst_bF_buf51), .B(\block[72] ), .Y(w_mem_inst__abc_21378_n3590_1) );
  AND2X2 AND2X2_3738 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf54), .B(w_mem_inst__abc_21378_n3590_1), .Y(w_mem_inst__abc_21378_n3591_1) );
  AND2X2 AND2X2_3739 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf19), .B(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_21378_n3594_1) );
  AND2X2 AND2X2_374 ( .A(_abc_15724_n1442), .B(_abc_15724_n1433), .Y(_abc_15724_n1448) );
  AND2X2 AND2X2_3740 ( .A(w_mem_inst__abc_21378_n3152_bF_buf53), .B(w_mem_inst_w_mem_14__9_), .Y(w_mem_inst__abc_21378_n3595_1) );
  AND2X2 AND2X2_3741 ( .A(round_ctr_rst_bF_buf50), .B(\block[73] ), .Y(w_mem_inst__abc_21378_n3596) );
  AND2X2 AND2X2_3742 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf53), .B(w_mem_inst__abc_21378_n3596), .Y(w_mem_inst__abc_21378_n3597) );
  AND2X2 AND2X2_3743 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf18), .B(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_21378_n3600) );
  AND2X2 AND2X2_3744 ( .A(w_mem_inst__abc_21378_n3152_bF_buf52), .B(w_mem_inst_w_mem_14__10_), .Y(w_mem_inst__abc_21378_n3601) );
  AND2X2 AND2X2_3745 ( .A(round_ctr_rst_bF_buf49), .B(\block[74] ), .Y(w_mem_inst__abc_21378_n3602_1) );
  AND2X2 AND2X2_3746 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf52), .B(w_mem_inst__abc_21378_n3602_1), .Y(w_mem_inst__abc_21378_n3603_1) );
  AND2X2 AND2X2_3747 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf17), .B(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_21378_n3606_1) );
  AND2X2 AND2X2_3748 ( .A(w_mem_inst__abc_21378_n3152_bF_buf51), .B(w_mem_inst_w_mem_14__11_), .Y(w_mem_inst__abc_21378_n3607_1) );
  AND2X2 AND2X2_3749 ( .A(round_ctr_rst_bF_buf48), .B(\block[75] ), .Y(w_mem_inst__abc_21378_n3608) );
  AND2X2 AND2X2_375 ( .A(_auto_iopadmap_cc_313_execute_26059_60_), .B(d_reg_28_), .Y(_abc_15724_n1452) );
  AND2X2 AND2X2_3750 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf51), .B(w_mem_inst__abc_21378_n3608), .Y(w_mem_inst__abc_21378_n3609) );
  AND2X2 AND2X2_3751 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf16), .B(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_21378_n3612) );
  AND2X2 AND2X2_3752 ( .A(w_mem_inst__abc_21378_n3152_bF_buf50), .B(w_mem_inst_w_mem_14__12_), .Y(w_mem_inst__abc_21378_n3613) );
  AND2X2 AND2X2_3753 ( .A(round_ctr_rst_bF_buf47), .B(\block[76] ), .Y(w_mem_inst__abc_21378_n3614_1) );
  AND2X2 AND2X2_3754 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf50), .B(w_mem_inst__abc_21378_n3614_1), .Y(w_mem_inst__abc_21378_n3615_1) );
  AND2X2 AND2X2_3755 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf15), .B(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_21378_n3618_1) );
  AND2X2 AND2X2_3756 ( .A(w_mem_inst__abc_21378_n3152_bF_buf49), .B(w_mem_inst_w_mem_14__13_), .Y(w_mem_inst__abc_21378_n3619_1) );
  AND2X2 AND2X2_3757 ( .A(round_ctr_rst_bF_buf46), .B(\block[77] ), .Y(w_mem_inst__abc_21378_n3620) );
  AND2X2 AND2X2_3758 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf49), .B(w_mem_inst__abc_21378_n3620), .Y(w_mem_inst__abc_21378_n3621) );
  AND2X2 AND2X2_3759 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf14), .B(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_21378_n3624) );
  AND2X2 AND2X2_376 ( .A(_abc_15724_n1453), .B(_abc_15724_n1451), .Y(_abc_15724_n1454) );
  AND2X2 AND2X2_3760 ( .A(w_mem_inst__abc_21378_n3152_bF_buf48), .B(w_mem_inst_w_mem_14__14_), .Y(w_mem_inst__abc_21378_n3625) );
  AND2X2 AND2X2_3761 ( .A(round_ctr_rst_bF_buf45), .B(\block[78] ), .Y(w_mem_inst__abc_21378_n3626_1) );
  AND2X2 AND2X2_3762 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf48), .B(w_mem_inst__abc_21378_n3626_1), .Y(w_mem_inst__abc_21378_n3627_1) );
  AND2X2 AND2X2_3763 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf13), .B(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_21378_n3630_1) );
  AND2X2 AND2X2_3764 ( .A(w_mem_inst__abc_21378_n3152_bF_buf47), .B(w_mem_inst_w_mem_14__15_), .Y(w_mem_inst__abc_21378_n3631_1) );
  AND2X2 AND2X2_3765 ( .A(round_ctr_rst_bF_buf44), .B(\block[79] ), .Y(w_mem_inst__abc_21378_n3632) );
  AND2X2 AND2X2_3766 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf47), .B(w_mem_inst__abc_21378_n3632), .Y(w_mem_inst__abc_21378_n3633) );
  AND2X2 AND2X2_3767 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf12), .B(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_21378_n3636) );
  AND2X2 AND2X2_3768 ( .A(w_mem_inst__abc_21378_n3152_bF_buf46), .B(w_mem_inst_w_mem_14__16_), .Y(w_mem_inst__abc_21378_n3637) );
  AND2X2 AND2X2_3769 ( .A(round_ctr_rst_bF_buf43), .B(\block[80] ), .Y(w_mem_inst__abc_21378_n3638_1) );
  AND2X2 AND2X2_377 ( .A(_abc_15724_n1440), .B(_abc_15724_n1448), .Y(_abc_15724_n1456) );
  AND2X2 AND2X2_3770 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf46), .B(w_mem_inst__abc_21378_n3638_1), .Y(w_mem_inst__abc_21378_n3639_1) );
  AND2X2 AND2X2_3771 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf11), .B(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_21378_n3642_1) );
  AND2X2 AND2X2_3772 ( .A(w_mem_inst__abc_21378_n3152_bF_buf45), .B(w_mem_inst_w_mem_14__17_), .Y(w_mem_inst__abc_21378_n3643_1) );
  AND2X2 AND2X2_3773 ( .A(round_ctr_rst_bF_buf42), .B(\block[81] ), .Y(w_mem_inst__abc_21378_n3644) );
  AND2X2 AND2X2_3774 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf45), .B(w_mem_inst__abc_21378_n3644), .Y(w_mem_inst__abc_21378_n3645) );
  AND2X2 AND2X2_3775 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf10), .B(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_21378_n3648) );
  AND2X2 AND2X2_3776 ( .A(w_mem_inst__abc_21378_n3152_bF_buf44), .B(w_mem_inst_w_mem_14__18_), .Y(w_mem_inst__abc_21378_n3649) );
  AND2X2 AND2X2_3777 ( .A(round_ctr_rst_bF_buf41), .B(\block[82] ), .Y(w_mem_inst__abc_21378_n3650_1) );
  AND2X2 AND2X2_3778 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf44), .B(w_mem_inst__abc_21378_n3650_1), .Y(w_mem_inst__abc_21378_n3651) );
  AND2X2 AND2X2_3779 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf9), .B(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_21378_n3654) );
  AND2X2 AND2X2_378 ( .A(_abc_15724_n1458), .B(_abc_15724_n1455), .Y(_abc_15724_n1459) );
  AND2X2 AND2X2_3780 ( .A(w_mem_inst__abc_21378_n3152_bF_buf43), .B(w_mem_inst_w_mem_14__19_), .Y(w_mem_inst__abc_21378_n3655) );
  AND2X2 AND2X2_3781 ( .A(round_ctr_rst_bF_buf40), .B(\block[83] ), .Y(w_mem_inst__abc_21378_n3656) );
  AND2X2 AND2X2_3782 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf43), .B(w_mem_inst__abc_21378_n3656), .Y(w_mem_inst__abc_21378_n3657_1) );
  AND2X2 AND2X2_3783 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf8), .B(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_21378_n3660) );
  AND2X2 AND2X2_3784 ( .A(w_mem_inst__abc_21378_n3152_bF_buf42), .B(w_mem_inst_w_mem_14__20_), .Y(w_mem_inst__abc_21378_n3661) );
  AND2X2 AND2X2_3785 ( .A(round_ctr_rst_bF_buf39), .B(\block[84] ), .Y(w_mem_inst__abc_21378_n3662_1) );
  AND2X2 AND2X2_3786 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf42), .B(w_mem_inst__abc_21378_n3662_1), .Y(w_mem_inst__abc_21378_n3663) );
  AND2X2 AND2X2_3787 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf7), .B(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_21378_n3666) );
  AND2X2 AND2X2_3788 ( .A(w_mem_inst__abc_21378_n3152_bF_buf41), .B(w_mem_inst_w_mem_14__21_), .Y(w_mem_inst__abc_21378_n3667) );
  AND2X2 AND2X2_3789 ( .A(round_ctr_rst_bF_buf38), .B(\block[85] ), .Y(w_mem_inst__abc_21378_n3668) );
  AND2X2 AND2X2_379 ( .A(_abc_15724_n1459), .B(digest_update_bF_buf8), .Y(_abc_15724_n1460) );
  AND2X2 AND2X2_3790 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf41), .B(w_mem_inst__abc_21378_n3668), .Y(w_mem_inst__abc_21378_n3669_1) );
  AND2X2 AND2X2_3791 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf6), .B(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_21378_n3672) );
  AND2X2 AND2X2_3792 ( .A(w_mem_inst__abc_21378_n3152_bF_buf40), .B(w_mem_inst_w_mem_14__22_), .Y(w_mem_inst__abc_21378_n3673_1) );
  AND2X2 AND2X2_3793 ( .A(round_ctr_rst_bF_buf37), .B(\block[86] ), .Y(w_mem_inst__abc_21378_n3674) );
  AND2X2 AND2X2_3794 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf40), .B(w_mem_inst__abc_21378_n3674), .Y(w_mem_inst__abc_21378_n3675) );
  AND2X2 AND2X2_3795 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf5), .B(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_21378_n3678) );
  AND2X2 AND2X2_3796 ( .A(w_mem_inst__abc_21378_n3152_bF_buf39), .B(w_mem_inst_w_mem_14__23_), .Y(w_mem_inst__abc_21378_n3679) );
  AND2X2 AND2X2_3797 ( .A(round_ctr_rst_bF_buf36), .B(\block[87] ), .Y(w_mem_inst__abc_21378_n3680) );
  AND2X2 AND2X2_3798 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf39), .B(w_mem_inst__abc_21378_n3680), .Y(w_mem_inst__abc_21378_n3681) );
  AND2X2 AND2X2_3799 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf4), .B(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_21378_n3684) );
  AND2X2 AND2X2_38 ( .A(_auto_iopadmap_cc_313_execute_26059_8_), .B(e_reg_8_), .Y(_abc_15724_n768) );
  AND2X2 AND2X2_380 ( .A(_abc_15724_n1461), .B(_abc_15724_n850_bF_buf6), .Y(_abc_15724_n1462_1) );
  AND2X2 AND2X2_3800 ( .A(w_mem_inst__abc_21378_n3152_bF_buf38), .B(w_mem_inst_w_mem_14__24_), .Y(w_mem_inst__abc_21378_n3685) );
  AND2X2 AND2X2_3801 ( .A(round_ctr_rst_bF_buf35), .B(\block[88] ), .Y(w_mem_inst__abc_21378_n3686) );
  AND2X2 AND2X2_3802 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf38), .B(w_mem_inst__abc_21378_n3686), .Y(w_mem_inst__abc_21378_n3687) );
  AND2X2 AND2X2_3803 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf3), .B(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_21378_n3690) );
  AND2X2 AND2X2_3804 ( .A(w_mem_inst__abc_21378_n3152_bF_buf37), .B(w_mem_inst_w_mem_14__25_), .Y(w_mem_inst__abc_21378_n3691) );
  AND2X2 AND2X2_3805 ( .A(round_ctr_rst_bF_buf34), .B(\block[89] ), .Y(w_mem_inst__abc_21378_n3692) );
  AND2X2 AND2X2_3806 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf37), .B(w_mem_inst__abc_21378_n3692), .Y(w_mem_inst__abc_21378_n3693) );
  AND2X2 AND2X2_3807 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf2), .B(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_21378_n3696) );
  AND2X2 AND2X2_3808 ( .A(w_mem_inst__abc_21378_n3152_bF_buf36), .B(w_mem_inst_w_mem_14__26_), .Y(w_mem_inst__abc_21378_n3697) );
  AND2X2 AND2X2_3809 ( .A(round_ctr_rst_bF_buf33), .B(\block[90] ), .Y(w_mem_inst__abc_21378_n3698) );
  AND2X2 AND2X2_381 ( .A(_abc_15724_n906_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_61_), .Y(_abc_15724_n1464_1) );
  AND2X2 AND2X2_3810 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf36), .B(w_mem_inst__abc_21378_n3698), .Y(w_mem_inst__abc_21378_n3699) );
  AND2X2 AND2X2_3811 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf1), .B(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_21378_n3702) );
  AND2X2 AND2X2_3812 ( .A(w_mem_inst__abc_21378_n3152_bF_buf35), .B(w_mem_inst_w_mem_14__27_), .Y(w_mem_inst__abc_21378_n3703) );
  AND2X2 AND2X2_3813 ( .A(round_ctr_rst_bF_buf32), .B(\block[91] ), .Y(w_mem_inst__abc_21378_n3704) );
  AND2X2 AND2X2_3814 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf35), .B(w_mem_inst__abc_21378_n3704), .Y(w_mem_inst__abc_21378_n3705) );
  AND2X2 AND2X2_3815 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf0), .B(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_21378_n3708) );
  AND2X2 AND2X2_3816 ( .A(w_mem_inst__abc_21378_n3152_bF_buf34), .B(w_mem_inst_w_mem_14__28_), .Y(w_mem_inst__abc_21378_n3709) );
  AND2X2 AND2X2_3817 ( .A(round_ctr_rst_bF_buf31), .B(\block[92] ), .Y(w_mem_inst__abc_21378_n3710) );
  AND2X2 AND2X2_3818 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf34), .B(w_mem_inst__abc_21378_n3710), .Y(w_mem_inst__abc_21378_n3711) );
  AND2X2 AND2X2_3819 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf60), .B(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_21378_n3714) );
  AND2X2 AND2X2_382 ( .A(_abc_15724_n1458), .B(_abc_15724_n1453), .Y(_abc_15724_n1466) );
  AND2X2 AND2X2_3820 ( .A(w_mem_inst__abc_21378_n3152_bF_buf33), .B(w_mem_inst_w_mem_14__29_), .Y(w_mem_inst__abc_21378_n3715) );
  AND2X2 AND2X2_3821 ( .A(round_ctr_rst_bF_buf30), .B(\block[93] ), .Y(w_mem_inst__abc_21378_n3716) );
  AND2X2 AND2X2_3822 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf33), .B(w_mem_inst__abc_21378_n3716), .Y(w_mem_inst__abc_21378_n3717) );
  AND2X2 AND2X2_3823 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf59), .B(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_21378_n3720) );
  AND2X2 AND2X2_3824 ( .A(w_mem_inst__abc_21378_n3152_bF_buf32), .B(w_mem_inst_w_mem_14__30_), .Y(w_mem_inst__abc_21378_n3721) );
  AND2X2 AND2X2_3825 ( .A(round_ctr_rst_bF_buf29), .B(\block[94] ), .Y(w_mem_inst__abc_21378_n3722) );
  AND2X2 AND2X2_3826 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf32), .B(w_mem_inst__abc_21378_n3722), .Y(w_mem_inst__abc_21378_n3723) );
  AND2X2 AND2X2_3827 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf58), .B(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_21378_n3726) );
  AND2X2 AND2X2_3828 ( .A(w_mem_inst__abc_21378_n3152_bF_buf31), .B(w_mem_inst_w_mem_14__31_), .Y(w_mem_inst__abc_21378_n3727) );
  AND2X2 AND2X2_3829 ( .A(round_ctr_rst_bF_buf28), .B(\block[95] ), .Y(w_mem_inst__abc_21378_n3728) );
  AND2X2 AND2X2_383 ( .A(_auto_iopadmap_cc_313_execute_26059_61_), .B(d_reg_29_), .Y(_abc_15724_n1468) );
  AND2X2 AND2X2_3830 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf31), .B(w_mem_inst__abc_21378_n3728), .Y(w_mem_inst__abc_21378_n3729) );
  AND2X2 AND2X2_3831 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf57), .B(w_mem_inst_w_mem_12__0_), .Y(w_mem_inst__abc_21378_n3732) );
  AND2X2 AND2X2_3832 ( .A(w_mem_inst__abc_21378_n3152_bF_buf30), .B(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_21378_n3733) );
  AND2X2 AND2X2_3833 ( .A(round_ctr_rst_bF_buf27), .B(\block[96] ), .Y(w_mem_inst__abc_21378_n3734) );
  AND2X2 AND2X2_3834 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf30), .B(w_mem_inst__abc_21378_n3734), .Y(w_mem_inst__abc_21378_n3735) );
  AND2X2 AND2X2_3835 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf56), .B(w_mem_inst_w_mem_12__1_), .Y(w_mem_inst__abc_21378_n3738) );
  AND2X2 AND2X2_3836 ( .A(w_mem_inst__abc_21378_n3152_bF_buf29), .B(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_21378_n3739) );
  AND2X2 AND2X2_3837 ( .A(round_ctr_rst_bF_buf26), .B(\block[97] ), .Y(w_mem_inst__abc_21378_n3740) );
  AND2X2 AND2X2_3838 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf29), .B(w_mem_inst__abc_21378_n3740), .Y(w_mem_inst__abc_21378_n3741) );
  AND2X2 AND2X2_3839 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf55), .B(w_mem_inst_w_mem_12__2_), .Y(w_mem_inst__abc_21378_n3744) );
  AND2X2 AND2X2_384 ( .A(_abc_15724_n1469), .B(_abc_15724_n1467), .Y(_abc_15724_n1470) );
  AND2X2 AND2X2_3840 ( .A(w_mem_inst__abc_21378_n3152_bF_buf28), .B(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_21378_n3745) );
  AND2X2 AND2X2_3841 ( .A(round_ctr_rst_bF_buf25), .B(\block[98] ), .Y(w_mem_inst__abc_21378_n3746) );
  AND2X2 AND2X2_3842 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf28), .B(w_mem_inst__abc_21378_n3746), .Y(w_mem_inst__abc_21378_n3747) );
  AND2X2 AND2X2_3843 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf54), .B(w_mem_inst_w_mem_12__3_), .Y(w_mem_inst__abc_21378_n3750) );
  AND2X2 AND2X2_3844 ( .A(w_mem_inst__abc_21378_n3152_bF_buf27), .B(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_21378_n3751) );
  AND2X2 AND2X2_3845 ( .A(round_ctr_rst_bF_buf24), .B(\block[99] ), .Y(w_mem_inst__abc_21378_n3752) );
  AND2X2 AND2X2_3846 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf27), .B(w_mem_inst__abc_21378_n3752), .Y(w_mem_inst__abc_21378_n3753) );
  AND2X2 AND2X2_3847 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf53), .B(w_mem_inst_w_mem_12__4_), .Y(w_mem_inst__abc_21378_n3756) );
  AND2X2 AND2X2_3848 ( .A(w_mem_inst__abc_21378_n3152_bF_buf26), .B(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_21378_n3757) );
  AND2X2 AND2X2_3849 ( .A(round_ctr_rst_bF_buf23), .B(\block[100] ), .Y(w_mem_inst__abc_21378_n3758) );
  AND2X2 AND2X2_385 ( .A(_abc_15724_n1466), .B(_abc_15724_n1470), .Y(_abc_15724_n1471) );
  AND2X2 AND2X2_3850 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf26), .B(w_mem_inst__abc_21378_n3758), .Y(w_mem_inst__abc_21378_n3759) );
  AND2X2 AND2X2_3851 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf52), .B(w_mem_inst_w_mem_12__5_), .Y(w_mem_inst__abc_21378_n3762) );
  AND2X2 AND2X2_3852 ( .A(w_mem_inst__abc_21378_n3152_bF_buf25), .B(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_21378_n3763) );
  AND2X2 AND2X2_3853 ( .A(round_ctr_rst_bF_buf22), .B(\block[101] ), .Y(w_mem_inst__abc_21378_n3764) );
  AND2X2 AND2X2_3854 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf25), .B(w_mem_inst__abc_21378_n3764), .Y(w_mem_inst__abc_21378_n3765) );
  AND2X2 AND2X2_3855 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf51), .B(w_mem_inst_w_mem_12__6_), .Y(w_mem_inst__abc_21378_n3768) );
  AND2X2 AND2X2_3856 ( .A(w_mem_inst__abc_21378_n3152_bF_buf24), .B(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_21378_n3769) );
  AND2X2 AND2X2_3857 ( .A(round_ctr_rst_bF_buf21), .B(\block[102] ), .Y(w_mem_inst__abc_21378_n3770) );
  AND2X2 AND2X2_3858 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf24), .B(w_mem_inst__abc_21378_n3770), .Y(w_mem_inst__abc_21378_n3771) );
  AND2X2 AND2X2_3859 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf50), .B(w_mem_inst_w_mem_12__7_), .Y(w_mem_inst__abc_21378_n3774) );
  AND2X2 AND2X2_386 ( .A(_abc_15724_n1450), .B(_abc_15724_n1454), .Y(_abc_15724_n1472_1) );
  AND2X2 AND2X2_3860 ( .A(w_mem_inst__abc_21378_n3152_bF_buf23), .B(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_21378_n3775) );
  AND2X2 AND2X2_3861 ( .A(round_ctr_rst_bF_buf20), .B(\block[103] ), .Y(w_mem_inst__abc_21378_n3776) );
  AND2X2 AND2X2_3862 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf23), .B(w_mem_inst__abc_21378_n3776), .Y(w_mem_inst__abc_21378_n3777) );
  AND2X2 AND2X2_3863 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf49), .B(w_mem_inst_w_mem_12__8_), .Y(w_mem_inst__abc_21378_n3780) );
  AND2X2 AND2X2_3864 ( .A(w_mem_inst__abc_21378_n3152_bF_buf22), .B(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_21378_n3781) );
  AND2X2 AND2X2_3865 ( .A(round_ctr_rst_bF_buf19), .B(\block[104] ), .Y(w_mem_inst__abc_21378_n3782) );
  AND2X2 AND2X2_3866 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf22), .B(w_mem_inst__abc_21378_n3782), .Y(w_mem_inst__abc_21378_n3783) );
  AND2X2 AND2X2_3867 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf48), .B(w_mem_inst_w_mem_12__9_), .Y(w_mem_inst__abc_21378_n3786) );
  AND2X2 AND2X2_3868 ( .A(w_mem_inst__abc_21378_n3152_bF_buf21), .B(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_21378_n3787) );
  AND2X2 AND2X2_3869 ( .A(round_ctr_rst_bF_buf18), .B(\block[105] ), .Y(w_mem_inst__abc_21378_n3788) );
  AND2X2 AND2X2_387 ( .A(_abc_15724_n1473_1), .B(_abc_15724_n1474_1), .Y(_abc_15724_n1475) );
  AND2X2 AND2X2_3870 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf21), .B(w_mem_inst__abc_21378_n3788), .Y(w_mem_inst__abc_21378_n3789) );
  AND2X2 AND2X2_3871 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf47), .B(w_mem_inst_w_mem_12__10_), .Y(w_mem_inst__abc_21378_n3792) );
  AND2X2 AND2X2_3872 ( .A(w_mem_inst__abc_21378_n3152_bF_buf20), .B(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_21378_n3793) );
  AND2X2 AND2X2_3873 ( .A(round_ctr_rst_bF_buf17), .B(\block[106] ), .Y(w_mem_inst__abc_21378_n3794) );
  AND2X2 AND2X2_3874 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf20), .B(w_mem_inst__abc_21378_n3794), .Y(w_mem_inst__abc_21378_n3795) );
  AND2X2 AND2X2_3875 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf46), .B(w_mem_inst_w_mem_12__11_), .Y(w_mem_inst__abc_21378_n3798) );
  AND2X2 AND2X2_3876 ( .A(w_mem_inst__abc_21378_n3152_bF_buf19), .B(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_21378_n3799) );
  AND2X2 AND2X2_3877 ( .A(round_ctr_rst_bF_buf16), .B(\block[107] ), .Y(w_mem_inst__abc_21378_n3800) );
  AND2X2 AND2X2_3878 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf19), .B(w_mem_inst__abc_21378_n3800), .Y(w_mem_inst__abc_21378_n3801) );
  AND2X2 AND2X2_3879 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf45), .B(w_mem_inst_w_mem_12__12_), .Y(w_mem_inst__abc_21378_n3804) );
  AND2X2 AND2X2_388 ( .A(_abc_15724_n1477), .B(_abc_15724_n1465), .Y(H3_reg_29__FF_INPUT) );
  AND2X2 AND2X2_3880 ( .A(w_mem_inst__abc_21378_n3152_bF_buf18), .B(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_21378_n3805) );
  AND2X2 AND2X2_3881 ( .A(round_ctr_rst_bF_buf15), .B(\block[108] ), .Y(w_mem_inst__abc_21378_n3806) );
  AND2X2 AND2X2_3882 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf18), .B(w_mem_inst__abc_21378_n3806), .Y(w_mem_inst__abc_21378_n3807) );
  AND2X2 AND2X2_3883 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf44), .B(w_mem_inst_w_mem_12__13_), .Y(w_mem_inst__abc_21378_n3810) );
  AND2X2 AND2X2_3884 ( .A(w_mem_inst__abc_21378_n3152_bF_buf17), .B(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_21378_n3811) );
  AND2X2 AND2X2_3885 ( .A(round_ctr_rst_bF_buf14), .B(\block[109] ), .Y(w_mem_inst__abc_21378_n3812) );
  AND2X2 AND2X2_3886 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf17), .B(w_mem_inst__abc_21378_n3812), .Y(w_mem_inst__abc_21378_n3813) );
  AND2X2 AND2X2_3887 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf43), .B(w_mem_inst_w_mem_12__14_), .Y(w_mem_inst__abc_21378_n3816) );
  AND2X2 AND2X2_3888 ( .A(w_mem_inst__abc_21378_n3152_bF_buf16), .B(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_21378_n3817) );
  AND2X2 AND2X2_3889 ( .A(round_ctr_rst_bF_buf13), .B(\block[110] ), .Y(w_mem_inst__abc_21378_n3818) );
  AND2X2 AND2X2_389 ( .A(_abc_15724_n907_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_62_), .Y(_abc_15724_n1479) );
  AND2X2 AND2X2_3890 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf16), .B(w_mem_inst__abc_21378_n3818), .Y(w_mem_inst__abc_21378_n3819) );
  AND2X2 AND2X2_3891 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf42), .B(w_mem_inst_w_mem_12__15_), .Y(w_mem_inst__abc_21378_n3822) );
  AND2X2 AND2X2_3892 ( .A(w_mem_inst__abc_21378_n3152_bF_buf15), .B(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_21378_n3823) );
  AND2X2 AND2X2_3893 ( .A(round_ctr_rst_bF_buf12), .B(\block[111] ), .Y(w_mem_inst__abc_21378_n3824) );
  AND2X2 AND2X2_3894 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf15), .B(w_mem_inst__abc_21378_n3824), .Y(w_mem_inst__abc_21378_n3825) );
  AND2X2 AND2X2_3895 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf41), .B(w_mem_inst_w_mem_12__16_), .Y(w_mem_inst__abc_21378_n3828) );
  AND2X2 AND2X2_3896 ( .A(w_mem_inst__abc_21378_n3152_bF_buf14), .B(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_21378_n3829) );
  AND2X2 AND2X2_3897 ( .A(round_ctr_rst_bF_buf11), .B(\block[112] ), .Y(w_mem_inst__abc_21378_n3830) );
  AND2X2 AND2X2_3898 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf14), .B(w_mem_inst__abc_21378_n3830), .Y(w_mem_inst__abc_21378_n3831) );
  AND2X2 AND2X2_3899 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf40), .B(w_mem_inst_w_mem_12__17_), .Y(w_mem_inst__abc_21378_n3834) );
  AND2X2 AND2X2_39 ( .A(_abc_15724_n767_1), .B(_abc_15724_n768), .Y(_abc_15724_n769_1) );
  AND2X2 AND2X2_390 ( .A(_auto_iopadmap_cc_313_execute_26059_62_), .B(d_reg_30_), .Y(_abc_15724_n1480) );
  AND2X2 AND2X2_3900 ( .A(w_mem_inst__abc_21378_n3152_bF_buf13), .B(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_21378_n3835) );
  AND2X2 AND2X2_3901 ( .A(round_ctr_rst_bF_buf10), .B(\block[113] ), .Y(w_mem_inst__abc_21378_n3836) );
  AND2X2 AND2X2_3902 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf13), .B(w_mem_inst__abc_21378_n3836), .Y(w_mem_inst__abc_21378_n3837) );
  AND2X2 AND2X2_3903 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf39), .B(w_mem_inst_w_mem_12__18_), .Y(w_mem_inst__abc_21378_n3840) );
  AND2X2 AND2X2_3904 ( .A(w_mem_inst__abc_21378_n3152_bF_buf12), .B(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_21378_n3841) );
  AND2X2 AND2X2_3905 ( .A(round_ctr_rst_bF_buf9), .B(\block[114] ), .Y(w_mem_inst__abc_21378_n3842) );
  AND2X2 AND2X2_3906 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf12), .B(w_mem_inst__abc_21378_n3842), .Y(w_mem_inst__abc_21378_n3843) );
  AND2X2 AND2X2_3907 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf38), .B(w_mem_inst_w_mem_12__19_), .Y(w_mem_inst__abc_21378_n3846) );
  AND2X2 AND2X2_3908 ( .A(w_mem_inst__abc_21378_n3152_bF_buf11), .B(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_21378_n3847) );
  AND2X2 AND2X2_3909 ( .A(round_ctr_rst_bF_buf8), .B(\block[115] ), .Y(w_mem_inst__abc_21378_n3848) );
  AND2X2 AND2X2_391 ( .A(_abc_15724_n1481), .B(_abc_15724_n1482), .Y(_abc_15724_n1483) );
  AND2X2 AND2X2_3910 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf11), .B(w_mem_inst__abc_21378_n3848), .Y(w_mem_inst__abc_21378_n3849) );
  AND2X2 AND2X2_3911 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf37), .B(w_mem_inst_w_mem_12__20_), .Y(w_mem_inst__abc_21378_n3852) );
  AND2X2 AND2X2_3912 ( .A(w_mem_inst__abc_21378_n3152_bF_buf10), .B(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_21378_n3853) );
  AND2X2 AND2X2_3913 ( .A(round_ctr_rst_bF_buf7), .B(\block[116] ), .Y(w_mem_inst__abc_21378_n3854) );
  AND2X2 AND2X2_3914 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf10), .B(w_mem_inst__abc_21378_n3854), .Y(w_mem_inst__abc_21378_n3855) );
  AND2X2 AND2X2_3915 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf36), .B(w_mem_inst_w_mem_12__21_), .Y(w_mem_inst__abc_21378_n3858) );
  AND2X2 AND2X2_3916 ( .A(w_mem_inst__abc_21378_n3152_bF_buf9), .B(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_21378_n3859) );
  AND2X2 AND2X2_3917 ( .A(round_ctr_rst_bF_buf6), .B(\block[117] ), .Y(w_mem_inst__abc_21378_n3860) );
  AND2X2 AND2X2_3918 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf9), .B(w_mem_inst__abc_21378_n3860), .Y(w_mem_inst__abc_21378_n3861) );
  AND2X2 AND2X2_3919 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf35), .B(w_mem_inst_w_mem_12__22_), .Y(w_mem_inst__abc_21378_n3864) );
  AND2X2 AND2X2_392 ( .A(_abc_15724_n1486), .B(_abc_15724_n1469), .Y(_abc_15724_n1487_1) );
  AND2X2 AND2X2_3920 ( .A(w_mem_inst__abc_21378_n3152_bF_buf8), .B(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_21378_n3865) );
  AND2X2 AND2X2_3921 ( .A(round_ctr_rst_bF_buf5), .B(\block[118] ), .Y(w_mem_inst__abc_21378_n3866) );
  AND2X2 AND2X2_3922 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf8), .B(w_mem_inst__abc_21378_n3866), .Y(w_mem_inst__abc_21378_n3867) );
  AND2X2 AND2X2_3923 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf34), .B(w_mem_inst_w_mem_12__23_), .Y(w_mem_inst__abc_21378_n3870) );
  AND2X2 AND2X2_3924 ( .A(w_mem_inst__abc_21378_n3152_bF_buf7), .B(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_21378_n3871) );
  AND2X2 AND2X2_3925 ( .A(round_ctr_rst_bF_buf4), .B(\block[119] ), .Y(w_mem_inst__abc_21378_n3872) );
  AND2X2 AND2X2_3926 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf7), .B(w_mem_inst__abc_21378_n3872), .Y(w_mem_inst__abc_21378_n3873) );
  AND2X2 AND2X2_3927 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf33), .B(w_mem_inst_w_mem_12__24_), .Y(w_mem_inst__abc_21378_n3876) );
  AND2X2 AND2X2_3928 ( .A(w_mem_inst__abc_21378_n3152_bF_buf6), .B(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_21378_n3877) );
  AND2X2 AND2X2_3929 ( .A(round_ctr_rst_bF_buf3), .B(\block[120] ), .Y(w_mem_inst__abc_21378_n3878) );
  AND2X2 AND2X2_393 ( .A(_abc_15724_n1473_1), .B(_abc_15724_n1467), .Y(_abc_15724_n1489) );
  AND2X2 AND2X2_3930 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf6), .B(w_mem_inst__abc_21378_n3878), .Y(w_mem_inst__abc_21378_n3879) );
  AND2X2 AND2X2_3931 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf32), .B(w_mem_inst_w_mem_12__25_), .Y(w_mem_inst__abc_21378_n3882) );
  AND2X2 AND2X2_3932 ( .A(w_mem_inst__abc_21378_n3152_bF_buf5), .B(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_21378_n3883) );
  AND2X2 AND2X2_3933 ( .A(round_ctr_rst_bF_buf2), .B(\block[121] ), .Y(w_mem_inst__abc_21378_n3884) );
  AND2X2 AND2X2_3934 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf5), .B(w_mem_inst__abc_21378_n3884), .Y(w_mem_inst__abc_21378_n3885) );
  AND2X2 AND2X2_3935 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf31), .B(w_mem_inst_w_mem_12__26_), .Y(w_mem_inst__abc_21378_n3888) );
  AND2X2 AND2X2_3936 ( .A(w_mem_inst__abc_21378_n3152_bF_buf4), .B(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_21378_n3889) );
  AND2X2 AND2X2_3937 ( .A(round_ctr_rst_bF_buf1), .B(\block[122] ), .Y(w_mem_inst__abc_21378_n3890) );
  AND2X2 AND2X2_3938 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf4), .B(w_mem_inst__abc_21378_n3890), .Y(w_mem_inst__abc_21378_n3891) );
  AND2X2 AND2X2_3939 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf30), .B(w_mem_inst_w_mem_12__27_), .Y(w_mem_inst__abc_21378_n3894) );
  AND2X2 AND2X2_394 ( .A(_abc_15724_n1491), .B(digest_update_bF_buf6), .Y(_abc_15724_n1492) );
  AND2X2 AND2X2_3940 ( .A(w_mem_inst__abc_21378_n3152_bF_buf3), .B(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_21378_n3895) );
  AND2X2 AND2X2_3941 ( .A(round_ctr_rst_bF_buf0), .B(\block[123] ), .Y(w_mem_inst__abc_21378_n3896) );
  AND2X2 AND2X2_3942 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf3), .B(w_mem_inst__abc_21378_n3896), .Y(w_mem_inst__abc_21378_n3897) );
  AND2X2 AND2X2_3943 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf29), .B(w_mem_inst_w_mem_12__28_), .Y(w_mem_inst__abc_21378_n3900) );
  AND2X2 AND2X2_3944 ( .A(w_mem_inst__abc_21378_n3152_bF_buf2), .B(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_21378_n3901) );
  AND2X2 AND2X2_3945 ( .A(round_ctr_rst_bF_buf63), .B(\block[124] ), .Y(w_mem_inst__abc_21378_n3902) );
  AND2X2 AND2X2_3946 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf2), .B(w_mem_inst__abc_21378_n3902), .Y(w_mem_inst__abc_21378_n3903) );
  AND2X2 AND2X2_3947 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf28), .B(w_mem_inst_w_mem_12__29_), .Y(w_mem_inst__abc_21378_n3906) );
  AND2X2 AND2X2_3948 ( .A(w_mem_inst__abc_21378_n3152_bF_buf1), .B(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_21378_n3907) );
  AND2X2 AND2X2_3949 ( .A(round_ctr_rst_bF_buf62), .B(\block[125] ), .Y(w_mem_inst__abc_21378_n3908) );
  AND2X2 AND2X2_395 ( .A(_abc_15724_n1492), .B(_abc_15724_n1488), .Y(_abc_15724_n1493_1) );
  AND2X2 AND2X2_3950 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf1), .B(w_mem_inst__abc_21378_n3908), .Y(w_mem_inst__abc_21378_n3909) );
  AND2X2 AND2X2_3951 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf27), .B(w_mem_inst_w_mem_12__30_), .Y(w_mem_inst__abc_21378_n3912) );
  AND2X2 AND2X2_3952 ( .A(w_mem_inst__abc_21378_n3152_bF_buf0), .B(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_21378_n3913) );
  AND2X2 AND2X2_3953 ( .A(round_ctr_rst_bF_buf61), .B(\block[126] ), .Y(w_mem_inst__abc_21378_n3914) );
  AND2X2 AND2X2_3954 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf0), .B(w_mem_inst__abc_21378_n3914), .Y(w_mem_inst__abc_21378_n3915) );
  AND2X2 AND2X2_3955 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf26), .B(w_mem_inst_w_mem_12__31_), .Y(w_mem_inst__abc_21378_n3918) );
  AND2X2 AND2X2_3956 ( .A(w_mem_inst__abc_21378_n3152_bF_buf63), .B(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_21378_n3919) );
  AND2X2 AND2X2_3957 ( .A(round_ctr_rst_bF_buf60), .B(\block[127] ), .Y(w_mem_inst__abc_21378_n3920) );
  AND2X2 AND2X2_3958 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf63), .B(w_mem_inst__abc_21378_n3920), .Y(w_mem_inst__abc_21378_n3921) );
  AND2X2 AND2X2_3959 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf25), .B(w_mem_inst_w_mem_11__0_), .Y(w_mem_inst__abc_21378_n3924) );
  AND2X2 AND2X2_396 ( .A(_abc_15724_n1488), .B(_abc_15724_n1481), .Y(_abc_15724_n1495) );
  AND2X2 AND2X2_3960 ( .A(w_mem_inst__abc_21378_n3152_bF_buf62), .B(w_mem_inst_w_mem_12__0_), .Y(w_mem_inst__abc_21378_n3925) );
  AND2X2 AND2X2_3961 ( .A(round_ctr_rst_bF_buf59), .B(\block[128] ), .Y(w_mem_inst__abc_21378_n3926) );
  AND2X2 AND2X2_3962 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf62), .B(w_mem_inst__abc_21378_n3926), .Y(w_mem_inst__abc_21378_n3927) );
  AND2X2 AND2X2_3963 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf24), .B(w_mem_inst_w_mem_11__1_), .Y(w_mem_inst__abc_21378_n3930) );
  AND2X2 AND2X2_3964 ( .A(w_mem_inst__abc_21378_n3152_bF_buf61), .B(w_mem_inst_w_mem_12__1_), .Y(w_mem_inst__abc_21378_n3931) );
  AND2X2 AND2X2_3965 ( .A(round_ctr_rst_bF_buf58), .B(\block[129] ), .Y(w_mem_inst__abc_21378_n3932) );
  AND2X2 AND2X2_3966 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf61), .B(w_mem_inst__abc_21378_n3932), .Y(w_mem_inst__abc_21378_n3933) );
  AND2X2 AND2X2_3967 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf23), .B(w_mem_inst_w_mem_11__2_), .Y(w_mem_inst__abc_21378_n3936) );
  AND2X2 AND2X2_3968 ( .A(w_mem_inst__abc_21378_n3152_bF_buf60), .B(w_mem_inst_w_mem_12__2_), .Y(w_mem_inst__abc_21378_n3937) );
  AND2X2 AND2X2_3969 ( .A(round_ctr_rst_bF_buf57), .B(\block[130] ), .Y(w_mem_inst__abc_21378_n3938) );
  AND2X2 AND2X2_397 ( .A(_auto_iopadmap_cc_313_execute_26059_63_), .B(d_reg_31_), .Y(_abc_15724_n1497) );
  AND2X2 AND2X2_3970 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf60), .B(w_mem_inst__abc_21378_n3938), .Y(w_mem_inst__abc_21378_n3939) );
  AND2X2 AND2X2_3971 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf22), .B(w_mem_inst_w_mem_11__3_), .Y(w_mem_inst__abc_21378_n3942) );
  AND2X2 AND2X2_3972 ( .A(w_mem_inst__abc_21378_n3152_bF_buf59), .B(w_mem_inst_w_mem_12__3_), .Y(w_mem_inst__abc_21378_n3943) );
  AND2X2 AND2X2_3973 ( .A(round_ctr_rst_bF_buf56), .B(\block[131] ), .Y(w_mem_inst__abc_21378_n3944) );
  AND2X2 AND2X2_3974 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf59), .B(w_mem_inst__abc_21378_n3944), .Y(w_mem_inst__abc_21378_n3945) );
  AND2X2 AND2X2_3975 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf21), .B(w_mem_inst_w_mem_11__4_), .Y(w_mem_inst__abc_21378_n3948) );
  AND2X2 AND2X2_3976 ( .A(w_mem_inst__abc_21378_n3152_bF_buf58), .B(w_mem_inst_w_mem_12__4_), .Y(w_mem_inst__abc_21378_n3949) );
  AND2X2 AND2X2_3977 ( .A(round_ctr_rst_bF_buf55), .B(\block[132] ), .Y(w_mem_inst__abc_21378_n3950) );
  AND2X2 AND2X2_3978 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf58), .B(w_mem_inst__abc_21378_n3950), .Y(w_mem_inst__abc_21378_n3951) );
  AND2X2 AND2X2_3979 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf20), .B(w_mem_inst_w_mem_11__5_), .Y(w_mem_inst__abc_21378_n3954) );
  AND2X2 AND2X2_398 ( .A(_abc_15724_n1498), .B(_abc_15724_n1496_1), .Y(_abc_15724_n1499) );
  AND2X2 AND2X2_3980 ( .A(w_mem_inst__abc_21378_n3152_bF_buf57), .B(w_mem_inst_w_mem_12__5_), .Y(w_mem_inst__abc_21378_n3955) );
  AND2X2 AND2X2_3981 ( .A(round_ctr_rst_bF_buf54), .B(\block[133] ), .Y(w_mem_inst__abc_21378_n3956) );
  AND2X2 AND2X2_3982 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf57), .B(w_mem_inst__abc_21378_n3956), .Y(w_mem_inst__abc_21378_n3957) );
  AND2X2 AND2X2_3983 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf19), .B(w_mem_inst_w_mem_11__6_), .Y(w_mem_inst__abc_21378_n3960) );
  AND2X2 AND2X2_3984 ( .A(w_mem_inst__abc_21378_n3152_bF_buf56), .B(w_mem_inst_w_mem_12__6_), .Y(w_mem_inst__abc_21378_n3961) );
  AND2X2 AND2X2_3985 ( .A(round_ctr_rst_bF_buf53), .B(\block[134] ), .Y(w_mem_inst__abc_21378_n3962) );
  AND2X2 AND2X2_3986 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf56), .B(w_mem_inst__abc_21378_n3962), .Y(w_mem_inst__abc_21378_n3963) );
  AND2X2 AND2X2_3987 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf18), .B(w_mem_inst_w_mem_11__7_), .Y(w_mem_inst__abc_21378_n3966) );
  AND2X2 AND2X2_3988 ( .A(w_mem_inst__abc_21378_n3152_bF_buf55), .B(w_mem_inst_w_mem_12__7_), .Y(w_mem_inst__abc_21378_n3967) );
  AND2X2 AND2X2_3989 ( .A(round_ctr_rst_bF_buf52), .B(\block[135] ), .Y(w_mem_inst__abc_21378_n3968) );
  AND2X2 AND2X2_399 ( .A(_abc_15724_n1495), .B(_abc_15724_n1499), .Y(_abc_15724_n1500) );
  AND2X2 AND2X2_3990 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf55), .B(w_mem_inst__abc_21378_n3968), .Y(w_mem_inst__abc_21378_n3969) );
  AND2X2 AND2X2_3991 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf17), .B(w_mem_inst_w_mem_11__8_), .Y(w_mem_inst__abc_21378_n3972) );
  AND2X2 AND2X2_3992 ( .A(w_mem_inst__abc_21378_n3152_bF_buf54), .B(w_mem_inst_w_mem_12__8_), .Y(w_mem_inst__abc_21378_n3973) );
  AND2X2 AND2X2_3993 ( .A(round_ctr_rst_bF_buf51), .B(\block[136] ), .Y(w_mem_inst__abc_21378_n3974) );
  AND2X2 AND2X2_3994 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf54), .B(w_mem_inst__abc_21378_n3974), .Y(w_mem_inst__abc_21378_n3975) );
  AND2X2 AND2X2_3995 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf16), .B(w_mem_inst_w_mem_11__9_), .Y(w_mem_inst__abc_21378_n3978) );
  AND2X2 AND2X2_3996 ( .A(w_mem_inst__abc_21378_n3152_bF_buf53), .B(w_mem_inst_w_mem_12__9_), .Y(w_mem_inst__abc_21378_n3979) );
  AND2X2 AND2X2_3997 ( .A(round_ctr_rst_bF_buf50), .B(\block[137] ), .Y(w_mem_inst__abc_21378_n3980) );
  AND2X2 AND2X2_3998 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf53), .B(w_mem_inst__abc_21378_n3980), .Y(w_mem_inst__abc_21378_n3981) );
  AND2X2 AND2X2_3999 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf15), .B(w_mem_inst_w_mem_11__10_), .Y(w_mem_inst__abc_21378_n3984) );
  AND2X2 AND2X2_4 ( .A(_abc_15724_n702), .B(_abc_15724_n699), .Y(_abc_15724_n703) );
  AND2X2 AND2X2_40 ( .A(_abc_15724_n765), .B(_abc_15724_n770), .Y(_abc_15724_n771) );
  AND2X2 AND2X2_400 ( .A(_abc_15724_n1490), .B(_abc_15724_n1483), .Y(_abc_15724_n1501) );
  AND2X2 AND2X2_4000 ( .A(w_mem_inst__abc_21378_n3152_bF_buf52), .B(w_mem_inst_w_mem_12__10_), .Y(w_mem_inst__abc_21378_n3985) );
  AND2X2 AND2X2_4001 ( .A(round_ctr_rst_bF_buf49), .B(\block[138] ), .Y(w_mem_inst__abc_21378_n3986) );
  AND2X2 AND2X2_4002 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf52), .B(w_mem_inst__abc_21378_n3986), .Y(w_mem_inst__abc_21378_n3987) );
  AND2X2 AND2X2_4003 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf14), .B(w_mem_inst_w_mem_11__11_), .Y(w_mem_inst__abc_21378_n3990) );
  AND2X2 AND2X2_4004 ( .A(w_mem_inst__abc_21378_n3152_bF_buf51), .B(w_mem_inst_w_mem_12__11_), .Y(w_mem_inst__abc_21378_n3991) );
  AND2X2 AND2X2_4005 ( .A(round_ctr_rst_bF_buf48), .B(\block[139] ), .Y(w_mem_inst__abc_21378_n3992) );
  AND2X2 AND2X2_4006 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf51), .B(w_mem_inst__abc_21378_n3992), .Y(w_mem_inst__abc_21378_n3993) );
  AND2X2 AND2X2_4007 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf13), .B(w_mem_inst_w_mem_11__12_), .Y(w_mem_inst__abc_21378_n3996) );
  AND2X2 AND2X2_4008 ( .A(w_mem_inst__abc_21378_n3152_bF_buf50), .B(w_mem_inst_w_mem_12__12_), .Y(w_mem_inst__abc_21378_n3997) );
  AND2X2 AND2X2_4009 ( .A(round_ctr_rst_bF_buf47), .B(\block[140] ), .Y(w_mem_inst__abc_21378_n3998) );
  AND2X2 AND2X2_401 ( .A(_abc_15724_n1502), .B(_abc_15724_n1503), .Y(_abc_15724_n1504) );
  AND2X2 AND2X2_4010 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf50), .B(w_mem_inst__abc_21378_n3998), .Y(w_mem_inst__abc_21378_n3999) );
  AND2X2 AND2X2_4011 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf12), .B(w_mem_inst_w_mem_11__13_), .Y(w_mem_inst__abc_21378_n4002) );
  AND2X2 AND2X2_4012 ( .A(w_mem_inst__abc_21378_n3152_bF_buf49), .B(w_mem_inst_w_mem_12__13_), .Y(w_mem_inst__abc_21378_n4003) );
  AND2X2 AND2X2_4013 ( .A(round_ctr_rst_bF_buf46), .B(\block[141] ), .Y(w_mem_inst__abc_21378_n4004) );
  AND2X2 AND2X2_4014 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf49), .B(w_mem_inst__abc_21378_n4004), .Y(w_mem_inst__abc_21378_n4005) );
  AND2X2 AND2X2_4015 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf11), .B(w_mem_inst_w_mem_11__14_), .Y(w_mem_inst__abc_21378_n4008) );
  AND2X2 AND2X2_4016 ( .A(w_mem_inst__abc_21378_n3152_bF_buf48), .B(w_mem_inst_w_mem_12__14_), .Y(w_mem_inst__abc_21378_n4009) );
  AND2X2 AND2X2_4017 ( .A(round_ctr_rst_bF_buf45), .B(\block[142] ), .Y(w_mem_inst__abc_21378_n4010) );
  AND2X2 AND2X2_4018 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf48), .B(w_mem_inst__abc_21378_n4010), .Y(w_mem_inst__abc_21378_n4011) );
  AND2X2 AND2X2_4019 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf10), .B(w_mem_inst_w_mem_11__15_), .Y(w_mem_inst__abc_21378_n4014) );
  AND2X2 AND2X2_402 ( .A(_abc_15724_n1505), .B(digest_update_bF_buf5), .Y(_abc_15724_n1506) );
  AND2X2 AND2X2_4020 ( .A(w_mem_inst__abc_21378_n3152_bF_buf47), .B(w_mem_inst_w_mem_12__15_), .Y(w_mem_inst__abc_21378_n4015) );
  AND2X2 AND2X2_4021 ( .A(round_ctr_rst_bF_buf44), .B(\block[143] ), .Y(w_mem_inst__abc_21378_n4016) );
  AND2X2 AND2X2_4022 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf47), .B(w_mem_inst__abc_21378_n4016), .Y(w_mem_inst__abc_21378_n4017) );
  AND2X2 AND2X2_4023 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf9), .B(w_mem_inst_w_mem_11__16_), .Y(w_mem_inst__abc_21378_n4020) );
  AND2X2 AND2X2_4024 ( .A(w_mem_inst__abc_21378_n3152_bF_buf46), .B(w_mem_inst_w_mem_12__16_), .Y(w_mem_inst__abc_21378_n4021) );
  AND2X2 AND2X2_4025 ( .A(round_ctr_rst_bF_buf43), .B(\block[144] ), .Y(w_mem_inst__abc_21378_n4022) );
  AND2X2 AND2X2_4026 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf46), .B(w_mem_inst__abc_21378_n4022), .Y(w_mem_inst__abc_21378_n4023) );
  AND2X2 AND2X2_4027 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf8), .B(w_mem_inst_w_mem_11__17_), .Y(w_mem_inst__abc_21378_n4026) );
  AND2X2 AND2X2_4028 ( .A(w_mem_inst__abc_21378_n3152_bF_buf45), .B(w_mem_inst_w_mem_12__17_), .Y(w_mem_inst__abc_21378_n4027) );
  AND2X2 AND2X2_4029 ( .A(round_ctr_rst_bF_buf42), .B(\block[145] ), .Y(w_mem_inst__abc_21378_n4028) );
  AND2X2 AND2X2_403 ( .A(_abc_15724_n907_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_63_), .Y(_abc_15724_n1507) );
  AND2X2 AND2X2_4030 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf45), .B(w_mem_inst__abc_21378_n4028), .Y(w_mem_inst__abc_21378_n4029) );
  AND2X2 AND2X2_4031 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf7), .B(w_mem_inst_w_mem_11__18_), .Y(w_mem_inst__abc_21378_n4032) );
  AND2X2 AND2X2_4032 ( .A(w_mem_inst__abc_21378_n3152_bF_buf44), .B(w_mem_inst_w_mem_12__18_), .Y(w_mem_inst__abc_21378_n4033) );
  AND2X2 AND2X2_4033 ( .A(round_ctr_rst_bF_buf41), .B(\block[146] ), .Y(w_mem_inst__abc_21378_n4034) );
  AND2X2 AND2X2_4034 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf44), .B(w_mem_inst__abc_21378_n4034), .Y(w_mem_inst__abc_21378_n4035) );
  AND2X2 AND2X2_4035 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf6), .B(w_mem_inst_w_mem_11__19_), .Y(w_mem_inst__abc_21378_n4038) );
  AND2X2 AND2X2_4036 ( .A(w_mem_inst__abc_21378_n3152_bF_buf43), .B(w_mem_inst_w_mem_12__19_), .Y(w_mem_inst__abc_21378_n4039) );
  AND2X2 AND2X2_4037 ( .A(round_ctr_rst_bF_buf40), .B(\block[147] ), .Y(w_mem_inst__abc_21378_n4040) );
  AND2X2 AND2X2_4038 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf43), .B(w_mem_inst__abc_21378_n4040), .Y(w_mem_inst__abc_21378_n4041) );
  AND2X2 AND2X2_4039 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf5), .B(w_mem_inst_w_mem_11__20_), .Y(w_mem_inst__abc_21378_n4044) );
  AND2X2 AND2X2_404 ( .A(_auto_iopadmap_cc_313_execute_26059_64_), .B(c_reg_0_), .Y(_abc_15724_n1510_1) );
  AND2X2 AND2X2_4040 ( .A(w_mem_inst__abc_21378_n3152_bF_buf42), .B(w_mem_inst_w_mem_12__20_), .Y(w_mem_inst__abc_21378_n4045) );
  AND2X2 AND2X2_4041 ( .A(round_ctr_rst_bF_buf39), .B(\block[148] ), .Y(w_mem_inst__abc_21378_n4046) );
  AND2X2 AND2X2_4042 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf42), .B(w_mem_inst__abc_21378_n4046), .Y(w_mem_inst__abc_21378_n4047) );
  AND2X2 AND2X2_4043 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf4), .B(w_mem_inst_w_mem_11__21_), .Y(w_mem_inst__abc_21378_n4050) );
  AND2X2 AND2X2_4044 ( .A(w_mem_inst__abc_21378_n3152_bF_buf41), .B(w_mem_inst_w_mem_12__21_), .Y(w_mem_inst__abc_21378_n4051) );
  AND2X2 AND2X2_4045 ( .A(round_ctr_rst_bF_buf38), .B(\block[149] ), .Y(w_mem_inst__abc_21378_n4052) );
  AND2X2 AND2X2_4046 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf41), .B(w_mem_inst__abc_21378_n4052), .Y(w_mem_inst__abc_21378_n4053) );
  AND2X2 AND2X2_4047 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf3), .B(w_mem_inst_w_mem_11__22_), .Y(w_mem_inst__abc_21378_n4056) );
  AND2X2 AND2X2_4048 ( .A(w_mem_inst__abc_21378_n3152_bF_buf40), .B(w_mem_inst_w_mem_12__22_), .Y(w_mem_inst__abc_21378_n4057) );
  AND2X2 AND2X2_4049 ( .A(round_ctr_rst_bF_buf37), .B(\block[150] ), .Y(w_mem_inst__abc_21378_n4058) );
  AND2X2 AND2X2_405 ( .A(_abc_15724_n1511), .B(_abc_15724_n1509_1), .Y(_abc_15724_n1512) );
  AND2X2 AND2X2_4050 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf40), .B(w_mem_inst__abc_21378_n4058), .Y(w_mem_inst__abc_21378_n4059) );
  AND2X2 AND2X2_4051 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf2), .B(w_mem_inst_w_mem_11__23_), .Y(w_mem_inst__abc_21378_n4062) );
  AND2X2 AND2X2_4052 ( .A(w_mem_inst__abc_21378_n3152_bF_buf39), .B(w_mem_inst_w_mem_12__23_), .Y(w_mem_inst__abc_21378_n4063) );
  AND2X2 AND2X2_4053 ( .A(round_ctr_rst_bF_buf36), .B(\block[151] ), .Y(w_mem_inst__abc_21378_n4064) );
  AND2X2 AND2X2_4054 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf39), .B(w_mem_inst__abc_21378_n4064), .Y(w_mem_inst__abc_21378_n4065) );
  AND2X2 AND2X2_4055 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf1), .B(w_mem_inst_w_mem_11__24_), .Y(w_mem_inst__abc_21378_n4068) );
  AND2X2 AND2X2_4056 ( .A(w_mem_inst__abc_21378_n3152_bF_buf38), .B(w_mem_inst_w_mem_12__24_), .Y(w_mem_inst__abc_21378_n4069) );
  AND2X2 AND2X2_4057 ( .A(round_ctr_rst_bF_buf35), .B(\block[152] ), .Y(w_mem_inst__abc_21378_n4070) );
  AND2X2 AND2X2_4058 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf38), .B(w_mem_inst__abc_21378_n4070), .Y(w_mem_inst__abc_21378_n4071) );
  AND2X2 AND2X2_4059 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf0), .B(w_mem_inst_w_mem_11__25_), .Y(w_mem_inst__abc_21378_n4074) );
  AND2X2 AND2X2_406 ( .A(_abc_15724_n906_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_64_), .Y(_abc_15724_n1514) );
  AND2X2 AND2X2_4060 ( .A(w_mem_inst__abc_21378_n3152_bF_buf37), .B(w_mem_inst_w_mem_12__25_), .Y(w_mem_inst__abc_21378_n4075) );
  AND2X2 AND2X2_4061 ( .A(round_ctr_rst_bF_buf34), .B(\block[153] ), .Y(w_mem_inst__abc_21378_n4076) );
  AND2X2 AND2X2_4062 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf37), .B(w_mem_inst__abc_21378_n4076), .Y(w_mem_inst__abc_21378_n4077) );
  AND2X2 AND2X2_4063 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf60), .B(w_mem_inst_w_mem_11__26_), .Y(w_mem_inst__abc_21378_n4080) );
  AND2X2 AND2X2_4064 ( .A(w_mem_inst__abc_21378_n3152_bF_buf36), .B(w_mem_inst_w_mem_12__26_), .Y(w_mem_inst__abc_21378_n4081) );
  AND2X2 AND2X2_4065 ( .A(round_ctr_rst_bF_buf33), .B(\block[154] ), .Y(w_mem_inst__abc_21378_n4082) );
  AND2X2 AND2X2_4066 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf36), .B(w_mem_inst__abc_21378_n4082), .Y(w_mem_inst__abc_21378_n4083) );
  AND2X2 AND2X2_4067 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf59), .B(w_mem_inst_w_mem_11__27_), .Y(w_mem_inst__abc_21378_n4086) );
  AND2X2 AND2X2_4068 ( .A(w_mem_inst__abc_21378_n3152_bF_buf35), .B(w_mem_inst_w_mem_12__27_), .Y(w_mem_inst__abc_21378_n4087) );
  AND2X2 AND2X2_4069 ( .A(round_ctr_rst_bF_buf32), .B(\block[155] ), .Y(w_mem_inst__abc_21378_n4088) );
  AND2X2 AND2X2_407 ( .A(_abc_15724_n1513), .B(_abc_15724_n1515), .Y(H2_reg_0__FF_INPUT) );
  AND2X2 AND2X2_4070 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf35), .B(w_mem_inst__abc_21378_n4088), .Y(w_mem_inst__abc_21378_n4089) );
  AND2X2 AND2X2_4071 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf58), .B(w_mem_inst_w_mem_11__28_), .Y(w_mem_inst__abc_21378_n4092) );
  AND2X2 AND2X2_4072 ( .A(w_mem_inst__abc_21378_n3152_bF_buf34), .B(w_mem_inst_w_mem_12__28_), .Y(w_mem_inst__abc_21378_n4093) );
  AND2X2 AND2X2_4073 ( .A(round_ctr_rst_bF_buf31), .B(\block[156] ), .Y(w_mem_inst__abc_21378_n4094) );
  AND2X2 AND2X2_4074 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf34), .B(w_mem_inst__abc_21378_n4094), .Y(w_mem_inst__abc_21378_n4095) );
  AND2X2 AND2X2_4075 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf57), .B(w_mem_inst_w_mem_11__29_), .Y(w_mem_inst__abc_21378_n4098) );
  AND2X2 AND2X2_4076 ( .A(w_mem_inst__abc_21378_n3152_bF_buf33), .B(w_mem_inst_w_mem_12__29_), .Y(w_mem_inst__abc_21378_n4099) );
  AND2X2 AND2X2_4077 ( .A(round_ctr_rst_bF_buf30), .B(\block[157] ), .Y(w_mem_inst__abc_21378_n4100) );
  AND2X2 AND2X2_4078 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf33), .B(w_mem_inst__abc_21378_n4100), .Y(w_mem_inst__abc_21378_n4101) );
  AND2X2 AND2X2_4079 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf56), .B(w_mem_inst_w_mem_11__30_), .Y(w_mem_inst__abc_21378_n4104) );
  AND2X2 AND2X2_408 ( .A(_auto_iopadmap_cc_313_execute_26059_65_), .B(c_reg_1_), .Y(_abc_15724_n1518_1) );
  AND2X2 AND2X2_4080 ( .A(w_mem_inst__abc_21378_n3152_bF_buf32), .B(w_mem_inst_w_mem_12__30_), .Y(w_mem_inst__abc_21378_n4105) );
  AND2X2 AND2X2_4081 ( .A(round_ctr_rst_bF_buf29), .B(\block[158] ), .Y(w_mem_inst__abc_21378_n4106) );
  AND2X2 AND2X2_4082 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf32), .B(w_mem_inst__abc_21378_n4106), .Y(w_mem_inst__abc_21378_n4107) );
  AND2X2 AND2X2_4083 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf55), .B(w_mem_inst_w_mem_11__31_), .Y(w_mem_inst__abc_21378_n4110) );
  AND2X2 AND2X2_4084 ( .A(w_mem_inst__abc_21378_n3152_bF_buf31), .B(w_mem_inst_w_mem_12__31_), .Y(w_mem_inst__abc_21378_n4111) );
  AND2X2 AND2X2_4085 ( .A(round_ctr_rst_bF_buf28), .B(\block[159] ), .Y(w_mem_inst__abc_21378_n4112) );
  AND2X2 AND2X2_4086 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf31), .B(w_mem_inst__abc_21378_n4112), .Y(w_mem_inst__abc_21378_n4113) );
  AND2X2 AND2X2_4087 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf54), .B(w_mem_inst_w_mem_10__0_), .Y(w_mem_inst__abc_21378_n4116) );
  AND2X2 AND2X2_4088 ( .A(w_mem_inst__abc_21378_n3152_bF_buf30), .B(w_mem_inst_w_mem_11__0_), .Y(w_mem_inst__abc_21378_n4117) );
  AND2X2 AND2X2_4089 ( .A(round_ctr_rst_bF_buf27), .B(\block[160] ), .Y(w_mem_inst__abc_21378_n4118) );
  AND2X2 AND2X2_409 ( .A(_abc_15724_n1519_1), .B(_abc_15724_n1517), .Y(_abc_15724_n1520_1) );
  AND2X2 AND2X2_4090 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf30), .B(w_mem_inst__abc_21378_n4118), .Y(w_mem_inst__abc_21378_n4119) );
  AND2X2 AND2X2_4091 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf53), .B(w_mem_inst_w_mem_10__1_), .Y(w_mem_inst__abc_21378_n4122) );
  AND2X2 AND2X2_4092 ( .A(w_mem_inst__abc_21378_n3152_bF_buf29), .B(w_mem_inst_w_mem_11__1_), .Y(w_mem_inst__abc_21378_n4123) );
  AND2X2 AND2X2_4093 ( .A(round_ctr_rst_bF_buf26), .B(\block[161] ), .Y(w_mem_inst__abc_21378_n4124) );
  AND2X2 AND2X2_4094 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf29), .B(w_mem_inst__abc_21378_n4124), .Y(w_mem_inst__abc_21378_n4125) );
  AND2X2 AND2X2_4095 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf52), .B(w_mem_inst_w_mem_10__2_), .Y(w_mem_inst__abc_21378_n4128) );
  AND2X2 AND2X2_4096 ( .A(w_mem_inst__abc_21378_n3152_bF_buf28), .B(w_mem_inst_w_mem_11__2_), .Y(w_mem_inst__abc_21378_n4129) );
  AND2X2 AND2X2_4097 ( .A(round_ctr_rst_bF_buf25), .B(\block[162] ), .Y(w_mem_inst__abc_21378_n4130) );
  AND2X2 AND2X2_4098 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf28), .B(w_mem_inst__abc_21378_n4130), .Y(w_mem_inst__abc_21378_n4131) );
  AND2X2 AND2X2_4099 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf51), .B(w_mem_inst_w_mem_10__3_), .Y(w_mem_inst__abc_21378_n4134) );
  AND2X2 AND2X2_41 ( .A(_auto_iopadmap_cc_313_execute_26059_7_), .B(e_reg_7_), .Y(_abc_15724_n773) );
  AND2X2 AND2X2_410 ( .A(_abc_15724_n1520_1), .B(_abc_15724_n1510_1), .Y(_abc_15724_n1521) );
  AND2X2 AND2X2_4100 ( .A(w_mem_inst__abc_21378_n3152_bF_buf27), .B(w_mem_inst_w_mem_11__3_), .Y(w_mem_inst__abc_21378_n4135) );
  AND2X2 AND2X2_4101 ( .A(round_ctr_rst_bF_buf24), .B(\block[163] ), .Y(w_mem_inst__abc_21378_n4136) );
  AND2X2 AND2X2_4102 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf27), .B(w_mem_inst__abc_21378_n4136), .Y(w_mem_inst__abc_21378_n4137) );
  AND2X2 AND2X2_4103 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf50), .B(w_mem_inst_w_mem_10__4_), .Y(w_mem_inst__abc_21378_n4140) );
  AND2X2 AND2X2_4104 ( .A(w_mem_inst__abc_21378_n3152_bF_buf26), .B(w_mem_inst_w_mem_11__4_), .Y(w_mem_inst__abc_21378_n4141) );
  AND2X2 AND2X2_4105 ( .A(round_ctr_rst_bF_buf23), .B(\block[164] ), .Y(w_mem_inst__abc_21378_n4142) );
  AND2X2 AND2X2_4106 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf26), .B(w_mem_inst__abc_21378_n4142), .Y(w_mem_inst__abc_21378_n4143) );
  AND2X2 AND2X2_4107 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf49), .B(w_mem_inst_w_mem_10__5_), .Y(w_mem_inst__abc_21378_n4146) );
  AND2X2 AND2X2_4108 ( .A(w_mem_inst__abc_21378_n3152_bF_buf25), .B(w_mem_inst_w_mem_11__5_), .Y(w_mem_inst__abc_21378_n4147) );
  AND2X2 AND2X2_4109 ( .A(round_ctr_rst_bF_buf22), .B(\block[165] ), .Y(w_mem_inst__abc_21378_n4148) );
  AND2X2 AND2X2_411 ( .A(_abc_15724_n1522), .B(_abc_15724_n1523), .Y(_abc_15724_n1524) );
  AND2X2 AND2X2_4110 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf25), .B(w_mem_inst__abc_21378_n4148), .Y(w_mem_inst__abc_21378_n4149) );
  AND2X2 AND2X2_4111 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf48), .B(w_mem_inst_w_mem_10__6_), .Y(w_mem_inst__abc_21378_n4152) );
  AND2X2 AND2X2_4112 ( .A(w_mem_inst__abc_21378_n3152_bF_buf24), .B(w_mem_inst_w_mem_11__6_), .Y(w_mem_inst__abc_21378_n4153) );
  AND2X2 AND2X2_4113 ( .A(round_ctr_rst_bF_buf21), .B(\block[166] ), .Y(w_mem_inst__abc_21378_n4154) );
  AND2X2 AND2X2_4114 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf24), .B(w_mem_inst__abc_21378_n4154), .Y(w_mem_inst__abc_21378_n4155) );
  AND2X2 AND2X2_4115 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf47), .B(w_mem_inst_w_mem_10__7_), .Y(w_mem_inst__abc_21378_n4158) );
  AND2X2 AND2X2_4116 ( .A(w_mem_inst__abc_21378_n3152_bF_buf23), .B(w_mem_inst_w_mem_11__7_), .Y(w_mem_inst__abc_21378_n4159) );
  AND2X2 AND2X2_4117 ( .A(round_ctr_rst_bF_buf20), .B(\block[167] ), .Y(w_mem_inst__abc_21378_n4160) );
  AND2X2 AND2X2_4118 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf23), .B(w_mem_inst__abc_21378_n4160), .Y(w_mem_inst__abc_21378_n4161) );
  AND2X2 AND2X2_4119 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf46), .B(w_mem_inst_w_mem_10__8_), .Y(w_mem_inst__abc_21378_n4164) );
  AND2X2 AND2X2_412 ( .A(_abc_15724_n1525), .B(_abc_15724_n1527), .Y(H2_reg_1__FF_INPUT) );
  AND2X2 AND2X2_4120 ( .A(w_mem_inst__abc_21378_n3152_bF_buf22), .B(w_mem_inst_w_mem_11__8_), .Y(w_mem_inst__abc_21378_n4165) );
  AND2X2 AND2X2_4121 ( .A(round_ctr_rst_bF_buf19), .B(\block[168] ), .Y(w_mem_inst__abc_21378_n4166) );
  AND2X2 AND2X2_4122 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf22), .B(w_mem_inst__abc_21378_n4166), .Y(w_mem_inst__abc_21378_n4167) );
  AND2X2 AND2X2_4123 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf45), .B(w_mem_inst_w_mem_10__9_), .Y(w_mem_inst__abc_21378_n4170) );
  AND2X2 AND2X2_4124 ( .A(w_mem_inst__abc_21378_n3152_bF_buf21), .B(w_mem_inst_w_mem_11__9_), .Y(w_mem_inst__abc_21378_n4171) );
  AND2X2 AND2X2_4125 ( .A(round_ctr_rst_bF_buf18), .B(\block[169] ), .Y(w_mem_inst__abc_21378_n4172) );
  AND2X2 AND2X2_4126 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf21), .B(w_mem_inst__abc_21378_n4172), .Y(w_mem_inst__abc_21378_n4173) );
  AND2X2 AND2X2_4127 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf44), .B(w_mem_inst_w_mem_10__10_), .Y(w_mem_inst__abc_21378_n4176) );
  AND2X2 AND2X2_4128 ( .A(w_mem_inst__abc_21378_n3152_bF_buf20), .B(w_mem_inst_w_mem_11__10_), .Y(w_mem_inst__abc_21378_n4177) );
  AND2X2 AND2X2_4129 ( .A(round_ctr_rst_bF_buf17), .B(\block[170] ), .Y(w_mem_inst__abc_21378_n4178) );
  AND2X2 AND2X2_413 ( .A(_abc_15724_n1522), .B(_abc_15724_n1519_1), .Y(_abc_15724_n1529) );
  AND2X2 AND2X2_4130 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf20), .B(w_mem_inst__abc_21378_n4178), .Y(w_mem_inst__abc_21378_n4179) );
  AND2X2 AND2X2_4131 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf43), .B(w_mem_inst_w_mem_10__11_), .Y(w_mem_inst__abc_21378_n4182) );
  AND2X2 AND2X2_4132 ( .A(w_mem_inst__abc_21378_n3152_bF_buf19), .B(w_mem_inst_w_mem_11__11_), .Y(w_mem_inst__abc_21378_n4183) );
  AND2X2 AND2X2_4133 ( .A(round_ctr_rst_bF_buf16), .B(\block[171] ), .Y(w_mem_inst__abc_21378_n4184) );
  AND2X2 AND2X2_4134 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf19), .B(w_mem_inst__abc_21378_n4184), .Y(w_mem_inst__abc_21378_n4185) );
  AND2X2 AND2X2_4135 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf42), .B(w_mem_inst_w_mem_10__12_), .Y(w_mem_inst__abc_21378_n4188) );
  AND2X2 AND2X2_4136 ( .A(w_mem_inst__abc_21378_n3152_bF_buf18), .B(w_mem_inst_w_mem_11__12_), .Y(w_mem_inst__abc_21378_n4189) );
  AND2X2 AND2X2_4137 ( .A(round_ctr_rst_bF_buf15), .B(\block[172] ), .Y(w_mem_inst__abc_21378_n4190) );
  AND2X2 AND2X2_4138 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf18), .B(w_mem_inst__abc_21378_n4190), .Y(w_mem_inst__abc_21378_n4191) );
  AND2X2 AND2X2_4139 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf41), .B(w_mem_inst_w_mem_10__13_), .Y(w_mem_inst__abc_21378_n4194) );
  AND2X2 AND2X2_414 ( .A(_auto_iopadmap_cc_313_execute_26059_66_), .B(c_reg_2_), .Y(_abc_15724_n1531_1) );
  AND2X2 AND2X2_4140 ( .A(w_mem_inst__abc_21378_n3152_bF_buf17), .B(w_mem_inst_w_mem_11__13_), .Y(w_mem_inst__abc_21378_n4195) );
  AND2X2 AND2X2_4141 ( .A(round_ctr_rst_bF_buf14), .B(\block[173] ), .Y(w_mem_inst__abc_21378_n4196) );
  AND2X2 AND2X2_4142 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf17), .B(w_mem_inst__abc_21378_n4196), .Y(w_mem_inst__abc_21378_n4197) );
  AND2X2 AND2X2_4143 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf40), .B(w_mem_inst_w_mem_10__14_), .Y(w_mem_inst__abc_21378_n4200) );
  AND2X2 AND2X2_4144 ( .A(w_mem_inst__abc_21378_n3152_bF_buf16), .B(w_mem_inst_w_mem_11__14_), .Y(w_mem_inst__abc_21378_n4201) );
  AND2X2 AND2X2_4145 ( .A(round_ctr_rst_bF_buf13), .B(\block[174] ), .Y(w_mem_inst__abc_21378_n4202) );
  AND2X2 AND2X2_4146 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf16), .B(w_mem_inst__abc_21378_n4202), .Y(w_mem_inst__abc_21378_n4203) );
  AND2X2 AND2X2_4147 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf39), .B(w_mem_inst_w_mem_10__15_), .Y(w_mem_inst__abc_21378_n4206) );
  AND2X2 AND2X2_4148 ( .A(w_mem_inst__abc_21378_n3152_bF_buf15), .B(w_mem_inst_w_mem_11__15_), .Y(w_mem_inst__abc_21378_n4207) );
  AND2X2 AND2X2_4149 ( .A(round_ctr_rst_bF_buf12), .B(\block[175] ), .Y(w_mem_inst__abc_21378_n4208) );
  AND2X2 AND2X2_415 ( .A(_abc_15724_n1532), .B(_abc_15724_n1530_1), .Y(_abc_15724_n1533_1) );
  AND2X2 AND2X2_4150 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf15), .B(w_mem_inst__abc_21378_n4208), .Y(w_mem_inst__abc_21378_n4209) );
  AND2X2 AND2X2_4151 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf38), .B(w_mem_inst_w_mem_10__16_), .Y(w_mem_inst__abc_21378_n4212) );
  AND2X2 AND2X2_4152 ( .A(w_mem_inst__abc_21378_n3152_bF_buf14), .B(w_mem_inst_w_mem_11__16_), .Y(w_mem_inst__abc_21378_n4213) );
  AND2X2 AND2X2_4153 ( .A(round_ctr_rst_bF_buf11), .B(\block[176] ), .Y(w_mem_inst__abc_21378_n4214) );
  AND2X2 AND2X2_4154 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf14), .B(w_mem_inst__abc_21378_n4214), .Y(w_mem_inst__abc_21378_n4215) );
  AND2X2 AND2X2_4155 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf37), .B(w_mem_inst_w_mem_10__17_), .Y(w_mem_inst__abc_21378_n4218) );
  AND2X2 AND2X2_4156 ( .A(w_mem_inst__abc_21378_n3152_bF_buf13), .B(w_mem_inst_w_mem_11__17_), .Y(w_mem_inst__abc_21378_n4219) );
  AND2X2 AND2X2_4157 ( .A(round_ctr_rst_bF_buf10), .B(\block[177] ), .Y(w_mem_inst__abc_21378_n4220) );
  AND2X2 AND2X2_4158 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf13), .B(w_mem_inst__abc_21378_n4220), .Y(w_mem_inst__abc_21378_n4221) );
  AND2X2 AND2X2_4159 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf36), .B(w_mem_inst_w_mem_10__18_), .Y(w_mem_inst__abc_21378_n4224) );
  AND2X2 AND2X2_416 ( .A(_abc_15724_n1537), .B(_abc_15724_n1535), .Y(_abc_15724_n1538_1) );
  AND2X2 AND2X2_4160 ( .A(w_mem_inst__abc_21378_n3152_bF_buf12), .B(w_mem_inst_w_mem_11__18_), .Y(w_mem_inst__abc_21378_n4225) );
  AND2X2 AND2X2_4161 ( .A(round_ctr_rst_bF_buf9), .B(\block[178] ), .Y(w_mem_inst__abc_21378_n4226) );
  AND2X2 AND2X2_4162 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf12), .B(w_mem_inst__abc_21378_n4226), .Y(w_mem_inst__abc_21378_n4227) );
  AND2X2 AND2X2_4163 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf35), .B(w_mem_inst_w_mem_10__19_), .Y(w_mem_inst__abc_21378_n4230) );
  AND2X2 AND2X2_4164 ( .A(w_mem_inst__abc_21378_n3152_bF_buf11), .B(w_mem_inst_w_mem_11__19_), .Y(w_mem_inst__abc_21378_n4231) );
  AND2X2 AND2X2_4165 ( .A(round_ctr_rst_bF_buf8), .B(\block[179] ), .Y(w_mem_inst__abc_21378_n4232) );
  AND2X2 AND2X2_4166 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf11), .B(w_mem_inst__abc_21378_n4232), .Y(w_mem_inst__abc_21378_n4233) );
  AND2X2 AND2X2_4167 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf34), .B(w_mem_inst_w_mem_10__20_), .Y(w_mem_inst__abc_21378_n4236) );
  AND2X2 AND2X2_4168 ( .A(w_mem_inst__abc_21378_n3152_bF_buf10), .B(w_mem_inst_w_mem_11__20_), .Y(w_mem_inst__abc_21378_n4237) );
  AND2X2 AND2X2_4169 ( .A(round_ctr_rst_bF_buf7), .B(\block[180] ), .Y(w_mem_inst__abc_21378_n4238) );
  AND2X2 AND2X2_417 ( .A(_abc_15724_n1539), .B(_abc_15724_n1541), .Y(H2_reg_2__FF_INPUT) );
  AND2X2 AND2X2_4170 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf10), .B(w_mem_inst__abc_21378_n4238), .Y(w_mem_inst__abc_21378_n4239) );
  AND2X2 AND2X2_4171 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf33), .B(w_mem_inst_w_mem_10__21_), .Y(w_mem_inst__abc_21378_n4242) );
  AND2X2 AND2X2_4172 ( .A(w_mem_inst__abc_21378_n3152_bF_buf9), .B(w_mem_inst_w_mem_11__21_), .Y(w_mem_inst__abc_21378_n4243) );
  AND2X2 AND2X2_4173 ( .A(round_ctr_rst_bF_buf6), .B(\block[181] ), .Y(w_mem_inst__abc_21378_n4244) );
  AND2X2 AND2X2_4174 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf9), .B(w_mem_inst__abc_21378_n4244), .Y(w_mem_inst__abc_21378_n4245) );
  AND2X2 AND2X2_4175 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf32), .B(w_mem_inst_w_mem_10__22_), .Y(w_mem_inst__abc_21378_n4248) );
  AND2X2 AND2X2_4176 ( .A(w_mem_inst__abc_21378_n3152_bF_buf8), .B(w_mem_inst_w_mem_11__22_), .Y(w_mem_inst__abc_21378_n4249) );
  AND2X2 AND2X2_4177 ( .A(round_ctr_rst_bF_buf5), .B(\block[182] ), .Y(w_mem_inst__abc_21378_n4250) );
  AND2X2 AND2X2_4178 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf8), .B(w_mem_inst__abc_21378_n4250), .Y(w_mem_inst__abc_21378_n4251) );
  AND2X2 AND2X2_4179 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf31), .B(w_mem_inst_w_mem_10__23_), .Y(w_mem_inst__abc_21378_n4254) );
  AND2X2 AND2X2_418 ( .A(_abc_15724_n1535), .B(_abc_15724_n1532), .Y(_abc_15724_n1543_1) );
  AND2X2 AND2X2_4180 ( .A(w_mem_inst__abc_21378_n3152_bF_buf7), .B(w_mem_inst_w_mem_11__23_), .Y(w_mem_inst__abc_21378_n4255) );
  AND2X2 AND2X2_4181 ( .A(round_ctr_rst_bF_buf4), .B(\block[183] ), .Y(w_mem_inst__abc_21378_n4256) );
  AND2X2 AND2X2_4182 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf7), .B(w_mem_inst__abc_21378_n4256), .Y(w_mem_inst__abc_21378_n4257) );
  AND2X2 AND2X2_4183 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf30), .B(w_mem_inst_w_mem_10__24_), .Y(w_mem_inst__abc_21378_n4260) );
  AND2X2 AND2X2_4184 ( .A(w_mem_inst__abc_21378_n3152_bF_buf6), .B(w_mem_inst_w_mem_11__24_), .Y(w_mem_inst__abc_21378_n4261) );
  AND2X2 AND2X2_4185 ( .A(round_ctr_rst_bF_buf3), .B(\block[184] ), .Y(w_mem_inst__abc_21378_n4262) );
  AND2X2 AND2X2_4186 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf6), .B(w_mem_inst__abc_21378_n4262), .Y(w_mem_inst__abc_21378_n4263) );
  AND2X2 AND2X2_4187 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf29), .B(w_mem_inst_w_mem_10__25_), .Y(w_mem_inst__abc_21378_n4266) );
  AND2X2 AND2X2_4188 ( .A(w_mem_inst__abc_21378_n3152_bF_buf5), .B(w_mem_inst_w_mem_11__25_), .Y(w_mem_inst__abc_21378_n4267) );
  AND2X2 AND2X2_4189 ( .A(round_ctr_rst_bF_buf2), .B(\block[185] ), .Y(w_mem_inst__abc_21378_n4268) );
  AND2X2 AND2X2_419 ( .A(_auto_iopadmap_cc_313_execute_26059_67_), .B(c_reg_3_), .Y(_abc_15724_n1545) );
  AND2X2 AND2X2_4190 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf5), .B(w_mem_inst__abc_21378_n4268), .Y(w_mem_inst__abc_21378_n4269) );
  AND2X2 AND2X2_4191 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf28), .B(w_mem_inst_w_mem_10__26_), .Y(w_mem_inst__abc_21378_n4272) );
  AND2X2 AND2X2_4192 ( .A(w_mem_inst__abc_21378_n3152_bF_buf4), .B(w_mem_inst_w_mem_11__26_), .Y(w_mem_inst__abc_21378_n4273) );
  AND2X2 AND2X2_4193 ( .A(round_ctr_rst_bF_buf1), .B(\block[186] ), .Y(w_mem_inst__abc_21378_n4274) );
  AND2X2 AND2X2_4194 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf4), .B(w_mem_inst__abc_21378_n4274), .Y(w_mem_inst__abc_21378_n4275) );
  AND2X2 AND2X2_4195 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf27), .B(w_mem_inst_w_mem_10__27_), .Y(w_mem_inst__abc_21378_n4278) );
  AND2X2 AND2X2_4196 ( .A(w_mem_inst__abc_21378_n3152_bF_buf3), .B(w_mem_inst_w_mem_11__27_), .Y(w_mem_inst__abc_21378_n4279) );
  AND2X2 AND2X2_4197 ( .A(round_ctr_rst_bF_buf0), .B(\block[187] ), .Y(w_mem_inst__abc_21378_n4280) );
  AND2X2 AND2X2_4198 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf3), .B(w_mem_inst__abc_21378_n4280), .Y(w_mem_inst__abc_21378_n4281) );
  AND2X2 AND2X2_4199 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf26), .B(w_mem_inst_w_mem_10__28_), .Y(w_mem_inst__abc_21378_n4284) );
  AND2X2 AND2X2_42 ( .A(_auto_iopadmap_cc_313_execute_26059_6_), .B(e_reg_6_), .Y(_abc_15724_n775) );
  AND2X2 AND2X2_420 ( .A(_abc_15724_n1546), .B(_abc_15724_n1544), .Y(_abc_15724_n1547) );
  AND2X2 AND2X2_4200 ( .A(w_mem_inst__abc_21378_n3152_bF_buf2), .B(w_mem_inst_w_mem_11__28_), .Y(w_mem_inst__abc_21378_n4285) );
  AND2X2 AND2X2_4201 ( .A(round_ctr_rst_bF_buf63), .B(\block[188] ), .Y(w_mem_inst__abc_21378_n4286) );
  AND2X2 AND2X2_4202 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf2), .B(w_mem_inst__abc_21378_n4286), .Y(w_mem_inst__abc_21378_n4287) );
  AND2X2 AND2X2_4203 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf25), .B(w_mem_inst_w_mem_10__29_), .Y(w_mem_inst__abc_21378_n4290) );
  AND2X2 AND2X2_4204 ( .A(w_mem_inst__abc_21378_n3152_bF_buf1), .B(w_mem_inst_w_mem_11__29_), .Y(w_mem_inst__abc_21378_n4291) );
  AND2X2 AND2X2_4205 ( .A(round_ctr_rst_bF_buf62), .B(\block[189] ), .Y(w_mem_inst__abc_21378_n4292) );
  AND2X2 AND2X2_4206 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf1), .B(w_mem_inst__abc_21378_n4292), .Y(w_mem_inst__abc_21378_n4293) );
  AND2X2 AND2X2_4207 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf24), .B(w_mem_inst_w_mem_10__30_), .Y(w_mem_inst__abc_21378_n4296) );
  AND2X2 AND2X2_4208 ( .A(w_mem_inst__abc_21378_n3152_bF_buf0), .B(w_mem_inst_w_mem_11__30_), .Y(w_mem_inst__abc_21378_n4297) );
  AND2X2 AND2X2_4209 ( .A(round_ctr_rst_bF_buf61), .B(\block[190] ), .Y(w_mem_inst__abc_21378_n4298) );
  AND2X2 AND2X2_421 ( .A(_abc_15724_n1543_1), .B(_abc_15724_n1547), .Y(_abc_15724_n1548_1) );
  AND2X2 AND2X2_4210 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf0), .B(w_mem_inst__abc_21378_n4298), .Y(w_mem_inst__abc_21378_n4299) );
  AND2X2 AND2X2_4211 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf23), .B(w_mem_inst_w_mem_10__31_), .Y(w_mem_inst__abc_21378_n4302) );
  AND2X2 AND2X2_4212 ( .A(w_mem_inst__abc_21378_n3152_bF_buf63), .B(w_mem_inst_w_mem_11__31_), .Y(w_mem_inst__abc_21378_n4303) );
  AND2X2 AND2X2_4213 ( .A(round_ctr_rst_bF_buf60), .B(\block[191] ), .Y(w_mem_inst__abc_21378_n4304) );
  AND2X2 AND2X2_4214 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf63), .B(w_mem_inst__abc_21378_n4304), .Y(w_mem_inst__abc_21378_n4305) );
  AND2X2 AND2X2_4215 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf22), .B(w_mem_inst_w_mem_9__0_), .Y(w_mem_inst__abc_21378_n4308) );
  AND2X2 AND2X2_4216 ( .A(w_mem_inst__abc_21378_n3152_bF_buf62), .B(w_mem_inst_w_mem_10__0_), .Y(w_mem_inst__abc_21378_n4309) );
  AND2X2 AND2X2_4217 ( .A(round_ctr_rst_bF_buf59), .B(\block[192] ), .Y(w_mem_inst__abc_21378_n4310) );
  AND2X2 AND2X2_4218 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf62), .B(w_mem_inst__abc_21378_n4310), .Y(w_mem_inst__abc_21378_n4311) );
  AND2X2 AND2X2_4219 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf21), .B(w_mem_inst_w_mem_9__1_), .Y(w_mem_inst__abc_21378_n4314) );
  AND2X2 AND2X2_422 ( .A(_abc_15724_n1549), .B(_abc_15724_n1550_1), .Y(_abc_15724_n1551) );
  AND2X2 AND2X2_4220 ( .A(w_mem_inst__abc_21378_n3152_bF_buf61), .B(w_mem_inst_w_mem_10__1_), .Y(w_mem_inst__abc_21378_n4315) );
  AND2X2 AND2X2_4221 ( .A(round_ctr_rst_bF_buf58), .B(\block[193] ), .Y(w_mem_inst__abc_21378_n4316) );
  AND2X2 AND2X2_4222 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf61), .B(w_mem_inst__abc_21378_n4316), .Y(w_mem_inst__abc_21378_n4317) );
  AND2X2 AND2X2_4223 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf20), .B(w_mem_inst_w_mem_9__2_), .Y(w_mem_inst__abc_21378_n4320) );
  AND2X2 AND2X2_4224 ( .A(w_mem_inst__abc_21378_n3152_bF_buf60), .B(w_mem_inst_w_mem_10__2_), .Y(w_mem_inst__abc_21378_n4321) );
  AND2X2 AND2X2_4225 ( .A(round_ctr_rst_bF_buf57), .B(\block[194] ), .Y(w_mem_inst__abc_21378_n4322) );
  AND2X2 AND2X2_4226 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf60), .B(w_mem_inst__abc_21378_n4322), .Y(w_mem_inst__abc_21378_n4323) );
  AND2X2 AND2X2_4227 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf19), .B(w_mem_inst_w_mem_9__3_), .Y(w_mem_inst__abc_21378_n4326) );
  AND2X2 AND2X2_4228 ( .A(w_mem_inst__abc_21378_n3152_bF_buf59), .B(w_mem_inst_w_mem_10__3_), .Y(w_mem_inst__abc_21378_n4327) );
  AND2X2 AND2X2_4229 ( .A(round_ctr_rst_bF_buf56), .B(\block[195] ), .Y(w_mem_inst__abc_21378_n4328) );
  AND2X2 AND2X2_423 ( .A(_abc_15724_n1552), .B(digest_update_bF_buf1), .Y(_abc_15724_n1553) );
  AND2X2 AND2X2_4230 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf59), .B(w_mem_inst__abc_21378_n4328), .Y(w_mem_inst__abc_21378_n4329) );
  AND2X2 AND2X2_4231 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf18), .B(w_mem_inst_w_mem_9__4_), .Y(w_mem_inst__abc_21378_n4332) );
  AND2X2 AND2X2_4232 ( .A(w_mem_inst__abc_21378_n3152_bF_buf58), .B(w_mem_inst_w_mem_10__4_), .Y(w_mem_inst__abc_21378_n4333) );
  AND2X2 AND2X2_4233 ( .A(round_ctr_rst_bF_buf55), .B(\block[196] ), .Y(w_mem_inst__abc_21378_n4334) );
  AND2X2 AND2X2_4234 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf58), .B(w_mem_inst__abc_21378_n4334), .Y(w_mem_inst__abc_21378_n4335) );
  AND2X2 AND2X2_4235 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf17), .B(w_mem_inst_w_mem_9__5_), .Y(w_mem_inst__abc_21378_n4338) );
  AND2X2 AND2X2_4236 ( .A(w_mem_inst__abc_21378_n3152_bF_buf57), .B(w_mem_inst_w_mem_10__5_), .Y(w_mem_inst__abc_21378_n4339) );
  AND2X2 AND2X2_4237 ( .A(round_ctr_rst_bF_buf54), .B(\block[197] ), .Y(w_mem_inst__abc_21378_n4340) );
  AND2X2 AND2X2_4238 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf57), .B(w_mem_inst__abc_21378_n4340), .Y(w_mem_inst__abc_21378_n4341) );
  AND2X2 AND2X2_4239 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf16), .B(w_mem_inst_w_mem_9__6_), .Y(w_mem_inst__abc_21378_n4344) );
  AND2X2 AND2X2_424 ( .A(_abc_15724_n1554), .B(_abc_15724_n850_bF_buf1), .Y(_abc_15724_n1555) );
  AND2X2 AND2X2_4240 ( .A(w_mem_inst__abc_21378_n3152_bF_buf56), .B(w_mem_inst_w_mem_10__6_), .Y(w_mem_inst__abc_21378_n4345) );
  AND2X2 AND2X2_4241 ( .A(round_ctr_rst_bF_buf53), .B(\block[198] ), .Y(w_mem_inst__abc_21378_n4346) );
  AND2X2 AND2X2_4242 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf56), .B(w_mem_inst__abc_21378_n4346), .Y(w_mem_inst__abc_21378_n4347) );
  AND2X2 AND2X2_4243 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf15), .B(w_mem_inst_w_mem_9__7_), .Y(w_mem_inst__abc_21378_n4350) );
  AND2X2 AND2X2_4244 ( .A(w_mem_inst__abc_21378_n3152_bF_buf55), .B(w_mem_inst_w_mem_10__7_), .Y(w_mem_inst__abc_21378_n4351) );
  AND2X2 AND2X2_4245 ( .A(round_ctr_rst_bF_buf52), .B(\block[199] ), .Y(w_mem_inst__abc_21378_n4352) );
  AND2X2 AND2X2_4246 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf55), .B(w_mem_inst__abc_21378_n4352), .Y(w_mem_inst__abc_21378_n4353) );
  AND2X2 AND2X2_4247 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf14), .B(w_mem_inst_w_mem_9__8_), .Y(w_mem_inst__abc_21378_n4356) );
  AND2X2 AND2X2_4248 ( .A(w_mem_inst__abc_21378_n3152_bF_buf54), .B(w_mem_inst_w_mem_10__8_), .Y(w_mem_inst__abc_21378_n4357) );
  AND2X2 AND2X2_4249 ( .A(round_ctr_rst_bF_buf51), .B(\block[200] ), .Y(w_mem_inst__abc_21378_n4358) );
  AND2X2 AND2X2_425 ( .A(_auto_iopadmap_cc_313_execute_26059_68_), .B(c_reg_4_), .Y(_abc_15724_n1558) );
  AND2X2 AND2X2_4250 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf54), .B(w_mem_inst__abc_21378_n4358), .Y(w_mem_inst__abc_21378_n4359) );
  AND2X2 AND2X2_4251 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf13), .B(w_mem_inst_w_mem_9__9_), .Y(w_mem_inst__abc_21378_n4362) );
  AND2X2 AND2X2_4252 ( .A(w_mem_inst__abc_21378_n3152_bF_buf53), .B(w_mem_inst_w_mem_10__9_), .Y(w_mem_inst__abc_21378_n4363) );
  AND2X2 AND2X2_4253 ( .A(round_ctr_rst_bF_buf50), .B(\block[201] ), .Y(w_mem_inst__abc_21378_n4364) );
  AND2X2 AND2X2_4254 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf53), .B(w_mem_inst__abc_21378_n4364), .Y(w_mem_inst__abc_21378_n4365) );
  AND2X2 AND2X2_4255 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf12), .B(w_mem_inst_w_mem_9__10_), .Y(w_mem_inst__abc_21378_n4368) );
  AND2X2 AND2X2_4256 ( .A(w_mem_inst__abc_21378_n3152_bF_buf52), .B(w_mem_inst_w_mem_10__10_), .Y(w_mem_inst__abc_21378_n4369) );
  AND2X2 AND2X2_4257 ( .A(round_ctr_rst_bF_buf49), .B(\block[202] ), .Y(w_mem_inst__abc_21378_n4370) );
  AND2X2 AND2X2_4258 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf52), .B(w_mem_inst__abc_21378_n4370), .Y(w_mem_inst__abc_21378_n4371) );
  AND2X2 AND2X2_4259 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf11), .B(w_mem_inst_w_mem_9__11_), .Y(w_mem_inst__abc_21378_n4374) );
  AND2X2 AND2X2_426 ( .A(_abc_15724_n1559), .B(_abc_15724_n1557_1), .Y(_abc_15724_n1560) );
  AND2X2 AND2X2_4260 ( .A(w_mem_inst__abc_21378_n3152_bF_buf51), .B(w_mem_inst_w_mem_10__11_), .Y(w_mem_inst__abc_21378_n4375) );
  AND2X2 AND2X2_4261 ( .A(round_ctr_rst_bF_buf48), .B(\block[203] ), .Y(w_mem_inst__abc_21378_n4376) );
  AND2X2 AND2X2_4262 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf51), .B(w_mem_inst__abc_21378_n4376), .Y(w_mem_inst__abc_21378_n4377) );
  AND2X2 AND2X2_4263 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf10), .B(w_mem_inst_w_mem_9__12_), .Y(w_mem_inst__abc_21378_n4380) );
  AND2X2 AND2X2_4264 ( .A(w_mem_inst__abc_21378_n3152_bF_buf50), .B(w_mem_inst_w_mem_10__12_), .Y(w_mem_inst__abc_21378_n4381) );
  AND2X2 AND2X2_4265 ( .A(round_ctr_rst_bF_buf47), .B(\block[204] ), .Y(w_mem_inst__abc_21378_n4382) );
  AND2X2 AND2X2_4266 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf50), .B(w_mem_inst__abc_21378_n4382), .Y(w_mem_inst__abc_21378_n4383) );
  AND2X2 AND2X2_4267 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf9), .B(w_mem_inst_w_mem_9__13_), .Y(w_mem_inst__abc_21378_n4386) );
  AND2X2 AND2X2_4268 ( .A(w_mem_inst__abc_21378_n3152_bF_buf49), .B(w_mem_inst_w_mem_10__13_), .Y(w_mem_inst__abc_21378_n4387) );
  AND2X2 AND2X2_4269 ( .A(round_ctr_rst_bF_buf46), .B(\block[205] ), .Y(w_mem_inst__abc_21378_n4388) );
  AND2X2 AND2X2_427 ( .A(_abc_15724_n1563_1), .B(_abc_15724_n1546), .Y(_abc_15724_n1564_1) );
  AND2X2 AND2X2_4270 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf49), .B(w_mem_inst__abc_21378_n4388), .Y(w_mem_inst__abc_21378_n4389) );
  AND2X2 AND2X2_4271 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf8), .B(w_mem_inst_w_mem_9__14_), .Y(w_mem_inst__abc_21378_n4392) );
  AND2X2 AND2X2_4272 ( .A(w_mem_inst__abc_21378_n3152_bF_buf48), .B(w_mem_inst_w_mem_10__14_), .Y(w_mem_inst__abc_21378_n4393) );
  AND2X2 AND2X2_4273 ( .A(round_ctr_rst_bF_buf45), .B(\block[206] ), .Y(w_mem_inst__abc_21378_n4394) );
  AND2X2 AND2X2_4274 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf48), .B(w_mem_inst__abc_21378_n4394), .Y(w_mem_inst__abc_21378_n4395) );
  AND2X2 AND2X2_4275 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf7), .B(w_mem_inst_w_mem_9__15_), .Y(w_mem_inst__abc_21378_n4398) );
  AND2X2 AND2X2_4276 ( .A(w_mem_inst__abc_21378_n3152_bF_buf47), .B(w_mem_inst_w_mem_10__15_), .Y(w_mem_inst__abc_21378_n4399) );
  AND2X2 AND2X2_4277 ( .A(round_ctr_rst_bF_buf44), .B(\block[207] ), .Y(w_mem_inst__abc_21378_n4400) );
  AND2X2 AND2X2_4278 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf47), .B(w_mem_inst__abc_21378_n4400), .Y(w_mem_inst__abc_21378_n4401) );
  AND2X2 AND2X2_4279 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf6), .B(w_mem_inst_w_mem_9__16_), .Y(w_mem_inst__abc_21378_n4404) );
  AND2X2 AND2X2_428 ( .A(_abc_15724_n1567), .B(_abc_15724_n1565), .Y(_abc_15724_n1568) );
  AND2X2 AND2X2_4280 ( .A(w_mem_inst__abc_21378_n3152_bF_buf46), .B(w_mem_inst_w_mem_10__16_), .Y(w_mem_inst__abc_21378_n4405) );
  AND2X2 AND2X2_4281 ( .A(round_ctr_rst_bF_buf43), .B(\block[208] ), .Y(w_mem_inst__abc_21378_n4406) );
  AND2X2 AND2X2_4282 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf46), .B(w_mem_inst__abc_21378_n4406), .Y(w_mem_inst__abc_21378_n4407) );
  AND2X2 AND2X2_4283 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf5), .B(w_mem_inst_w_mem_9__17_), .Y(w_mem_inst__abc_21378_n4410) );
  AND2X2 AND2X2_4284 ( .A(w_mem_inst__abc_21378_n3152_bF_buf45), .B(w_mem_inst_w_mem_10__17_), .Y(w_mem_inst__abc_21378_n4411) );
  AND2X2 AND2X2_4285 ( .A(round_ctr_rst_bF_buf42), .B(\block[209] ), .Y(w_mem_inst__abc_21378_n4412) );
  AND2X2 AND2X2_4286 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf45), .B(w_mem_inst__abc_21378_n4412), .Y(w_mem_inst__abc_21378_n4413) );
  AND2X2 AND2X2_4287 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf4), .B(w_mem_inst_w_mem_9__18_), .Y(w_mem_inst__abc_21378_n4416) );
  AND2X2 AND2X2_4288 ( .A(w_mem_inst__abc_21378_n3152_bF_buf44), .B(w_mem_inst_w_mem_10__18_), .Y(w_mem_inst__abc_21378_n4417) );
  AND2X2 AND2X2_4289 ( .A(round_ctr_rst_bF_buf41), .B(\block[210] ), .Y(w_mem_inst__abc_21378_n4418) );
  AND2X2 AND2X2_429 ( .A(_abc_15724_n1569), .B(_abc_15724_n1571_1), .Y(H2_reg_4__FF_INPUT) );
  AND2X2 AND2X2_4290 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf44), .B(w_mem_inst__abc_21378_n4418), .Y(w_mem_inst__abc_21378_n4419) );
  AND2X2 AND2X2_4291 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf3), .B(w_mem_inst_w_mem_9__19_), .Y(w_mem_inst__abc_21378_n4422) );
  AND2X2 AND2X2_4292 ( .A(w_mem_inst__abc_21378_n3152_bF_buf43), .B(w_mem_inst_w_mem_10__19_), .Y(w_mem_inst__abc_21378_n4423) );
  AND2X2 AND2X2_4293 ( .A(round_ctr_rst_bF_buf40), .B(\block[211] ), .Y(w_mem_inst__abc_21378_n4424) );
  AND2X2 AND2X2_4294 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf43), .B(w_mem_inst__abc_21378_n4424), .Y(w_mem_inst__abc_21378_n4425) );
  AND2X2 AND2X2_4295 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf2), .B(w_mem_inst_w_mem_9__20_), .Y(w_mem_inst__abc_21378_n4428) );
  AND2X2 AND2X2_4296 ( .A(w_mem_inst__abc_21378_n3152_bF_buf42), .B(w_mem_inst_w_mem_10__20_), .Y(w_mem_inst__abc_21378_n4429) );
  AND2X2 AND2X2_4297 ( .A(round_ctr_rst_bF_buf39), .B(\block[212] ), .Y(w_mem_inst__abc_21378_n4430) );
  AND2X2 AND2X2_4298 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf42), .B(w_mem_inst__abc_21378_n4430), .Y(w_mem_inst__abc_21378_n4431) );
  AND2X2 AND2X2_4299 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf1), .B(w_mem_inst_w_mem_9__21_), .Y(w_mem_inst__abc_21378_n4434) );
  AND2X2 AND2X2_43 ( .A(_abc_15724_n774), .B(_abc_15724_n775), .Y(_abc_15724_n776) );
  AND2X2 AND2X2_430 ( .A(_abc_15724_n1565), .B(_abc_15724_n1559), .Y(_abc_15724_n1573_1) );
  AND2X2 AND2X2_4300 ( .A(w_mem_inst__abc_21378_n3152_bF_buf41), .B(w_mem_inst_w_mem_10__21_), .Y(w_mem_inst__abc_21378_n4435) );
  AND2X2 AND2X2_4301 ( .A(round_ctr_rst_bF_buf38), .B(\block[213] ), .Y(w_mem_inst__abc_21378_n4436) );
  AND2X2 AND2X2_4302 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf41), .B(w_mem_inst__abc_21378_n4436), .Y(w_mem_inst__abc_21378_n4437) );
  AND2X2 AND2X2_4303 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf0), .B(w_mem_inst_w_mem_9__22_), .Y(w_mem_inst__abc_21378_n4440) );
  AND2X2 AND2X2_4304 ( .A(w_mem_inst__abc_21378_n3152_bF_buf40), .B(w_mem_inst_w_mem_10__22_), .Y(w_mem_inst__abc_21378_n4441) );
  AND2X2 AND2X2_4305 ( .A(round_ctr_rst_bF_buf37), .B(\block[214] ), .Y(w_mem_inst__abc_21378_n4442) );
  AND2X2 AND2X2_4306 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf40), .B(w_mem_inst__abc_21378_n4442), .Y(w_mem_inst__abc_21378_n4443) );
  AND2X2 AND2X2_4307 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf60), .B(w_mem_inst_w_mem_9__23_), .Y(w_mem_inst__abc_21378_n4446) );
  AND2X2 AND2X2_4308 ( .A(w_mem_inst__abc_21378_n3152_bF_buf39), .B(w_mem_inst_w_mem_10__23_), .Y(w_mem_inst__abc_21378_n4447) );
  AND2X2 AND2X2_4309 ( .A(round_ctr_rst_bF_buf36), .B(\block[215] ), .Y(w_mem_inst__abc_21378_n4448) );
  AND2X2 AND2X2_431 ( .A(_auto_iopadmap_cc_313_execute_26059_69_), .B(c_reg_5_), .Y(_abc_15724_n1576) );
  AND2X2 AND2X2_4310 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf39), .B(w_mem_inst__abc_21378_n4448), .Y(w_mem_inst__abc_21378_n4449) );
  AND2X2 AND2X2_4311 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf59), .B(w_mem_inst_w_mem_9__24_), .Y(w_mem_inst__abc_21378_n4452) );
  AND2X2 AND2X2_4312 ( .A(w_mem_inst__abc_21378_n3152_bF_buf38), .B(w_mem_inst_w_mem_10__24_), .Y(w_mem_inst__abc_21378_n4453) );
  AND2X2 AND2X2_4313 ( .A(round_ctr_rst_bF_buf35), .B(\block[216] ), .Y(w_mem_inst__abc_21378_n4454) );
  AND2X2 AND2X2_4314 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf38), .B(w_mem_inst__abc_21378_n4454), .Y(w_mem_inst__abc_21378_n4455) );
  AND2X2 AND2X2_4315 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf58), .B(w_mem_inst_w_mem_9__25_), .Y(w_mem_inst__abc_21378_n4458) );
  AND2X2 AND2X2_4316 ( .A(w_mem_inst__abc_21378_n3152_bF_buf37), .B(w_mem_inst_w_mem_10__25_), .Y(w_mem_inst__abc_21378_n4459) );
  AND2X2 AND2X2_4317 ( .A(round_ctr_rst_bF_buf34), .B(\block[217] ), .Y(w_mem_inst__abc_21378_n4460) );
  AND2X2 AND2X2_4318 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf37), .B(w_mem_inst__abc_21378_n4460), .Y(w_mem_inst__abc_21378_n4461) );
  AND2X2 AND2X2_4319 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf57), .B(w_mem_inst_w_mem_9__26_), .Y(w_mem_inst__abc_21378_n4464) );
  AND2X2 AND2X2_432 ( .A(_abc_15724_n1577), .B(_abc_15724_n1575), .Y(_abc_15724_n1578_1) );
  AND2X2 AND2X2_4320 ( .A(w_mem_inst__abc_21378_n3152_bF_buf36), .B(w_mem_inst_w_mem_10__26_), .Y(w_mem_inst__abc_21378_n4465) );
  AND2X2 AND2X2_4321 ( .A(round_ctr_rst_bF_buf33), .B(\block[218] ), .Y(w_mem_inst__abc_21378_n4466) );
  AND2X2 AND2X2_4322 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf36), .B(w_mem_inst__abc_21378_n4466), .Y(w_mem_inst__abc_21378_n4467) );
  AND2X2 AND2X2_4323 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf56), .B(w_mem_inst_w_mem_9__27_), .Y(w_mem_inst__abc_21378_n4470) );
  AND2X2 AND2X2_4324 ( .A(w_mem_inst__abc_21378_n3152_bF_buf35), .B(w_mem_inst_w_mem_10__27_), .Y(w_mem_inst__abc_21378_n4471) );
  AND2X2 AND2X2_4325 ( .A(round_ctr_rst_bF_buf32), .B(\block[219] ), .Y(w_mem_inst__abc_21378_n4472) );
  AND2X2 AND2X2_4326 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf35), .B(w_mem_inst__abc_21378_n4472), .Y(w_mem_inst__abc_21378_n4473) );
  AND2X2 AND2X2_4327 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf55), .B(w_mem_inst_w_mem_9__28_), .Y(w_mem_inst__abc_21378_n4476) );
  AND2X2 AND2X2_4328 ( .A(w_mem_inst__abc_21378_n3152_bF_buf34), .B(w_mem_inst_w_mem_10__28_), .Y(w_mem_inst__abc_21378_n4477) );
  AND2X2 AND2X2_4329 ( .A(round_ctr_rst_bF_buf31), .B(\block[220] ), .Y(w_mem_inst__abc_21378_n4478) );
  AND2X2 AND2X2_433 ( .A(_abc_15724_n1581_1), .B(digest_update_bF_buf11), .Y(_abc_15724_n1582) );
  AND2X2 AND2X2_4330 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf34), .B(w_mem_inst__abc_21378_n4478), .Y(w_mem_inst__abc_21378_n4479) );
  AND2X2 AND2X2_4331 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf54), .B(w_mem_inst_w_mem_9__29_), .Y(w_mem_inst__abc_21378_n4482) );
  AND2X2 AND2X2_4332 ( .A(w_mem_inst__abc_21378_n3152_bF_buf33), .B(w_mem_inst_w_mem_10__29_), .Y(w_mem_inst__abc_21378_n4483) );
  AND2X2 AND2X2_4333 ( .A(round_ctr_rst_bF_buf30), .B(\block[221] ), .Y(w_mem_inst__abc_21378_n4484) );
  AND2X2 AND2X2_4334 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf33), .B(w_mem_inst__abc_21378_n4484), .Y(w_mem_inst__abc_21378_n4485) );
  AND2X2 AND2X2_4335 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf53), .B(w_mem_inst_w_mem_9__30_), .Y(w_mem_inst__abc_21378_n4488) );
  AND2X2 AND2X2_4336 ( .A(w_mem_inst__abc_21378_n3152_bF_buf32), .B(w_mem_inst_w_mem_10__30_), .Y(w_mem_inst__abc_21378_n4489) );
  AND2X2 AND2X2_4337 ( .A(round_ctr_rst_bF_buf29), .B(\block[222] ), .Y(w_mem_inst__abc_21378_n4490) );
  AND2X2 AND2X2_4338 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf32), .B(w_mem_inst__abc_21378_n4490), .Y(w_mem_inst__abc_21378_n4491) );
  AND2X2 AND2X2_4339 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf52), .B(w_mem_inst_w_mem_9__31_), .Y(w_mem_inst__abc_21378_n4494) );
  AND2X2 AND2X2_434 ( .A(_abc_15724_n1582), .B(_abc_15724_n1579_1), .Y(_abc_15724_n1583) );
  AND2X2 AND2X2_4340 ( .A(w_mem_inst__abc_21378_n3152_bF_buf31), .B(w_mem_inst_w_mem_10__31_), .Y(w_mem_inst__abc_21378_n4495) );
  AND2X2 AND2X2_4341 ( .A(round_ctr_rst_bF_buf28), .B(\block[223] ), .Y(w_mem_inst__abc_21378_n4496) );
  AND2X2 AND2X2_4342 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf31), .B(w_mem_inst__abc_21378_n4496), .Y(w_mem_inst__abc_21378_n4497) );
  AND2X2 AND2X2_4343 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf51), .B(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_21378_n4500) );
  AND2X2 AND2X2_4344 ( .A(w_mem_inst__abc_21378_n3152_bF_buf30), .B(w_mem_inst_w_mem_9__0_), .Y(w_mem_inst__abc_21378_n4501) );
  AND2X2 AND2X2_4345 ( .A(round_ctr_rst_bF_buf27), .B(\block[224] ), .Y(w_mem_inst__abc_21378_n4502) );
  AND2X2 AND2X2_4346 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf30), .B(w_mem_inst__abc_21378_n4502), .Y(w_mem_inst__abc_21378_n4503) );
  AND2X2 AND2X2_4347 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf50), .B(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_21378_n4506) );
  AND2X2 AND2X2_4348 ( .A(w_mem_inst__abc_21378_n3152_bF_buf29), .B(w_mem_inst_w_mem_9__1_), .Y(w_mem_inst__abc_21378_n4507) );
  AND2X2 AND2X2_4349 ( .A(round_ctr_rst_bF_buf26), .B(\block[225] ), .Y(w_mem_inst__abc_21378_n4508) );
  AND2X2 AND2X2_435 ( .A(_abc_15724_n1584_1), .B(_abc_15724_n850_bF_buf8), .Y(_abc_15724_n1585_1) );
  AND2X2 AND2X2_4350 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf29), .B(w_mem_inst__abc_21378_n4508), .Y(w_mem_inst__abc_21378_n4509) );
  AND2X2 AND2X2_4351 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf49), .B(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_21378_n4512) );
  AND2X2 AND2X2_4352 ( .A(w_mem_inst__abc_21378_n3152_bF_buf28), .B(w_mem_inst_w_mem_9__2_), .Y(w_mem_inst__abc_21378_n4513) );
  AND2X2 AND2X2_4353 ( .A(round_ctr_rst_bF_buf25), .B(\block[226] ), .Y(w_mem_inst__abc_21378_n4514) );
  AND2X2 AND2X2_4354 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf28), .B(w_mem_inst__abc_21378_n4514), .Y(w_mem_inst__abc_21378_n4515) );
  AND2X2 AND2X2_4355 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf48), .B(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_21378_n4518) );
  AND2X2 AND2X2_4356 ( .A(w_mem_inst__abc_21378_n3152_bF_buf27), .B(w_mem_inst_w_mem_9__3_), .Y(w_mem_inst__abc_21378_n4519) );
  AND2X2 AND2X2_4357 ( .A(round_ctr_rst_bF_buf24), .B(\block[227] ), .Y(w_mem_inst__abc_21378_n4520) );
  AND2X2 AND2X2_4358 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf27), .B(w_mem_inst__abc_21378_n4520), .Y(w_mem_inst__abc_21378_n4521) );
  AND2X2 AND2X2_4359 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf47), .B(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_21378_n4524) );
  AND2X2 AND2X2_436 ( .A(_abc_15724_n1581_1), .B(_abc_15724_n1577), .Y(_abc_15724_n1587_1) );
  AND2X2 AND2X2_4360 ( .A(w_mem_inst__abc_21378_n3152_bF_buf26), .B(w_mem_inst_w_mem_9__4_), .Y(w_mem_inst__abc_21378_n4525) );
  AND2X2 AND2X2_4361 ( .A(round_ctr_rst_bF_buf23), .B(\block[228] ), .Y(w_mem_inst__abc_21378_n4526) );
  AND2X2 AND2X2_4362 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf26), .B(w_mem_inst__abc_21378_n4526), .Y(w_mem_inst__abc_21378_n4527) );
  AND2X2 AND2X2_4363 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf46), .B(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_21378_n4530) );
  AND2X2 AND2X2_4364 ( .A(w_mem_inst__abc_21378_n3152_bF_buf25), .B(w_mem_inst_w_mem_9__5_), .Y(w_mem_inst__abc_21378_n4531) );
  AND2X2 AND2X2_4365 ( .A(round_ctr_rst_bF_buf22), .B(\block[229] ), .Y(w_mem_inst__abc_21378_n4532) );
  AND2X2 AND2X2_4366 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf25), .B(w_mem_inst__abc_21378_n4532), .Y(w_mem_inst__abc_21378_n4533) );
  AND2X2 AND2X2_4367 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf45), .B(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_21378_n4536) );
  AND2X2 AND2X2_4368 ( .A(w_mem_inst__abc_21378_n3152_bF_buf24), .B(w_mem_inst_w_mem_9__6_), .Y(w_mem_inst__abc_21378_n4537) );
  AND2X2 AND2X2_4369 ( .A(round_ctr_rst_bF_buf21), .B(\block[230] ), .Y(w_mem_inst__abc_21378_n4538) );
  AND2X2 AND2X2_437 ( .A(_auto_iopadmap_cc_313_execute_26059_70_), .B(c_reg_6_), .Y(_abc_15724_n1590_1) );
  AND2X2 AND2X2_4370 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf24), .B(w_mem_inst__abc_21378_n4538), .Y(w_mem_inst__abc_21378_n4539) );
  AND2X2 AND2X2_4371 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf44), .B(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_21378_n4542) );
  AND2X2 AND2X2_4372 ( .A(w_mem_inst__abc_21378_n3152_bF_buf23), .B(w_mem_inst_w_mem_9__7_), .Y(w_mem_inst__abc_21378_n4543) );
  AND2X2 AND2X2_4373 ( .A(round_ctr_rst_bF_buf20), .B(\block[231] ), .Y(w_mem_inst__abc_21378_n4544) );
  AND2X2 AND2X2_4374 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf23), .B(w_mem_inst__abc_21378_n4544), .Y(w_mem_inst__abc_21378_n4545) );
  AND2X2 AND2X2_4375 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf43), .B(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_21378_n4548) );
  AND2X2 AND2X2_4376 ( .A(w_mem_inst__abc_21378_n3152_bF_buf22), .B(w_mem_inst_w_mem_9__8_), .Y(w_mem_inst__abc_21378_n4549) );
  AND2X2 AND2X2_4377 ( .A(round_ctr_rst_bF_buf19), .B(\block[232] ), .Y(w_mem_inst__abc_21378_n4550) );
  AND2X2 AND2X2_4378 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf22), .B(w_mem_inst__abc_21378_n4550), .Y(w_mem_inst__abc_21378_n4551) );
  AND2X2 AND2X2_4379 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf42), .B(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_21378_n4554) );
  AND2X2 AND2X2_438 ( .A(_abc_15724_n1591_1), .B(_abc_15724_n1589), .Y(_abc_15724_n1592) );
  AND2X2 AND2X2_4380 ( .A(w_mem_inst__abc_21378_n3152_bF_buf21), .B(w_mem_inst_w_mem_9__9_), .Y(w_mem_inst__abc_21378_n4555) );
  AND2X2 AND2X2_4381 ( .A(round_ctr_rst_bF_buf18), .B(\block[233] ), .Y(w_mem_inst__abc_21378_n4556) );
  AND2X2 AND2X2_4382 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf21), .B(w_mem_inst__abc_21378_n4556), .Y(w_mem_inst__abc_21378_n4557) );
  AND2X2 AND2X2_4383 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf41), .B(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_21378_n4560) );
  AND2X2 AND2X2_4384 ( .A(w_mem_inst__abc_21378_n3152_bF_buf20), .B(w_mem_inst_w_mem_9__10_), .Y(w_mem_inst__abc_21378_n4561) );
  AND2X2 AND2X2_4385 ( .A(round_ctr_rst_bF_buf17), .B(\block[234] ), .Y(w_mem_inst__abc_21378_n4562) );
  AND2X2 AND2X2_4386 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf20), .B(w_mem_inst__abc_21378_n4562), .Y(w_mem_inst__abc_21378_n4563) );
  AND2X2 AND2X2_4387 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf40), .B(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_21378_n4566) );
  AND2X2 AND2X2_4388 ( .A(w_mem_inst__abc_21378_n3152_bF_buf19), .B(w_mem_inst_w_mem_9__11_), .Y(w_mem_inst__abc_21378_n4567) );
  AND2X2 AND2X2_4389 ( .A(round_ctr_rst_bF_buf16), .B(\block[235] ), .Y(w_mem_inst__abc_21378_n4568) );
  AND2X2 AND2X2_439 ( .A(_abc_15724_n1595), .B(digest_update_bF_buf10), .Y(_abc_15724_n1596_1) );
  AND2X2 AND2X2_4390 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf19), .B(w_mem_inst__abc_21378_n4568), .Y(w_mem_inst__abc_21378_n4569) );
  AND2X2 AND2X2_4391 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf39), .B(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_21378_n4572) );
  AND2X2 AND2X2_4392 ( .A(w_mem_inst__abc_21378_n3152_bF_buf18), .B(w_mem_inst_w_mem_9__12_), .Y(w_mem_inst__abc_21378_n4573) );
  AND2X2 AND2X2_4393 ( .A(round_ctr_rst_bF_buf15), .B(\block[236] ), .Y(w_mem_inst__abc_21378_n4574) );
  AND2X2 AND2X2_4394 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf18), .B(w_mem_inst__abc_21378_n4574), .Y(w_mem_inst__abc_21378_n4575) );
  AND2X2 AND2X2_4395 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf38), .B(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_21378_n4578) );
  AND2X2 AND2X2_4396 ( .A(w_mem_inst__abc_21378_n3152_bF_buf17), .B(w_mem_inst_w_mem_9__13_), .Y(w_mem_inst__abc_21378_n4579) );
  AND2X2 AND2X2_4397 ( .A(round_ctr_rst_bF_buf14), .B(\block[237] ), .Y(w_mem_inst__abc_21378_n4580) );
  AND2X2 AND2X2_4398 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf17), .B(w_mem_inst__abc_21378_n4580), .Y(w_mem_inst__abc_21378_n4581) );
  AND2X2 AND2X2_4399 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf37), .B(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_21378_n4584) );
  AND2X2 AND2X2_44 ( .A(_abc_15724_n778), .B(_abc_15724_n774), .Y(_abc_15724_n779_1) );
  AND2X2 AND2X2_440 ( .A(_abc_15724_n1596_1), .B(_abc_15724_n1593_1), .Y(_abc_15724_n1597_1) );
  AND2X2 AND2X2_4400 ( .A(w_mem_inst__abc_21378_n3152_bF_buf16), .B(w_mem_inst_w_mem_9__14_), .Y(w_mem_inst__abc_21378_n4585) );
  AND2X2 AND2X2_4401 ( .A(round_ctr_rst_bF_buf13), .B(\block[238] ), .Y(w_mem_inst__abc_21378_n4586) );
  AND2X2 AND2X2_4402 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf16), .B(w_mem_inst__abc_21378_n4586), .Y(w_mem_inst__abc_21378_n4587) );
  AND2X2 AND2X2_4403 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf36), .B(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_21378_n4590) );
  AND2X2 AND2X2_4404 ( .A(w_mem_inst__abc_21378_n3152_bF_buf15), .B(w_mem_inst_w_mem_9__15_), .Y(w_mem_inst__abc_21378_n4591) );
  AND2X2 AND2X2_4405 ( .A(round_ctr_rst_bF_buf12), .B(\block[239] ), .Y(w_mem_inst__abc_21378_n4592) );
  AND2X2 AND2X2_4406 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf15), .B(w_mem_inst__abc_21378_n4592), .Y(w_mem_inst__abc_21378_n4593) );
  AND2X2 AND2X2_4407 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf35), .B(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_21378_n4596) );
  AND2X2 AND2X2_4408 ( .A(w_mem_inst__abc_21378_n3152_bF_buf14), .B(w_mem_inst_w_mem_9__16_), .Y(w_mem_inst__abc_21378_n4597) );
  AND2X2 AND2X2_4409 ( .A(round_ctr_rst_bF_buf11), .B(\block[240] ), .Y(w_mem_inst__abc_21378_n4598) );
  AND2X2 AND2X2_441 ( .A(_abc_15724_n1598), .B(_abc_15724_n850_bF_buf7), .Y(_abc_15724_n1599_1) );
  AND2X2 AND2X2_4410 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf14), .B(w_mem_inst__abc_21378_n4598), .Y(w_mem_inst__abc_21378_n4599) );
  AND2X2 AND2X2_4411 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf34), .B(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_21378_n4602) );
  AND2X2 AND2X2_4412 ( .A(w_mem_inst__abc_21378_n3152_bF_buf13), .B(w_mem_inst_w_mem_9__17_), .Y(w_mem_inst__abc_21378_n4603) );
  AND2X2 AND2X2_4413 ( .A(round_ctr_rst_bF_buf10), .B(\block[241] ), .Y(w_mem_inst__abc_21378_n4604) );
  AND2X2 AND2X2_4414 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf13), .B(w_mem_inst__abc_21378_n4604), .Y(w_mem_inst__abc_21378_n4605) );
  AND2X2 AND2X2_4415 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf33), .B(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_21378_n4608) );
  AND2X2 AND2X2_4416 ( .A(w_mem_inst__abc_21378_n3152_bF_buf12), .B(w_mem_inst_w_mem_9__18_), .Y(w_mem_inst__abc_21378_n4609) );
  AND2X2 AND2X2_4417 ( .A(round_ctr_rst_bF_buf9), .B(\block[242] ), .Y(w_mem_inst__abc_21378_n4610) );
  AND2X2 AND2X2_4418 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf12), .B(w_mem_inst__abc_21378_n4610), .Y(w_mem_inst__abc_21378_n4611) );
  AND2X2 AND2X2_4419 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf32), .B(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_21378_n4614) );
  AND2X2 AND2X2_442 ( .A(_abc_15724_n1595), .B(_abc_15724_n1591_1), .Y(_abc_15724_n1601) );
  AND2X2 AND2X2_4420 ( .A(w_mem_inst__abc_21378_n3152_bF_buf11), .B(w_mem_inst_w_mem_9__19_), .Y(w_mem_inst__abc_21378_n4615) );
  AND2X2 AND2X2_4421 ( .A(round_ctr_rst_bF_buf8), .B(\block[243] ), .Y(w_mem_inst__abc_21378_n4616) );
  AND2X2 AND2X2_4422 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf11), .B(w_mem_inst__abc_21378_n4616), .Y(w_mem_inst__abc_21378_n4617) );
  AND2X2 AND2X2_4423 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf31), .B(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_21378_n4620) );
  AND2X2 AND2X2_4424 ( .A(w_mem_inst__abc_21378_n3152_bF_buf10), .B(w_mem_inst_w_mem_9__20_), .Y(w_mem_inst__abc_21378_n4621) );
  AND2X2 AND2X2_4425 ( .A(round_ctr_rst_bF_buf7), .B(\block[244] ), .Y(w_mem_inst__abc_21378_n4622) );
  AND2X2 AND2X2_4426 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf10), .B(w_mem_inst__abc_21378_n4622), .Y(w_mem_inst__abc_21378_n4623) );
  AND2X2 AND2X2_4427 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf30), .B(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_21378_n4626) );
  AND2X2 AND2X2_4428 ( .A(w_mem_inst__abc_21378_n3152_bF_buf9), .B(w_mem_inst_w_mem_9__21_), .Y(w_mem_inst__abc_21378_n4627) );
  AND2X2 AND2X2_4429 ( .A(round_ctr_rst_bF_buf6), .B(\block[245] ), .Y(w_mem_inst__abc_21378_n4628) );
  AND2X2 AND2X2_443 ( .A(_auto_iopadmap_cc_313_execute_26059_71_), .B(c_reg_7_), .Y(_abc_15724_n1604) );
  AND2X2 AND2X2_4430 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf9), .B(w_mem_inst__abc_21378_n4628), .Y(w_mem_inst__abc_21378_n4629) );
  AND2X2 AND2X2_4431 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf29), .B(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_21378_n4632) );
  AND2X2 AND2X2_4432 ( .A(w_mem_inst__abc_21378_n3152_bF_buf8), .B(w_mem_inst_w_mem_9__22_), .Y(w_mem_inst__abc_21378_n4633) );
  AND2X2 AND2X2_4433 ( .A(round_ctr_rst_bF_buf5), .B(\block[246] ), .Y(w_mem_inst__abc_21378_n4634) );
  AND2X2 AND2X2_4434 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf8), .B(w_mem_inst__abc_21378_n4634), .Y(w_mem_inst__abc_21378_n4635) );
  AND2X2 AND2X2_4435 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf28), .B(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_21378_n4638) );
  AND2X2 AND2X2_4436 ( .A(w_mem_inst__abc_21378_n3152_bF_buf7), .B(w_mem_inst_w_mem_9__23_), .Y(w_mem_inst__abc_21378_n4639) );
  AND2X2 AND2X2_4437 ( .A(round_ctr_rst_bF_buf4), .B(\block[247] ), .Y(w_mem_inst__abc_21378_n4640) );
  AND2X2 AND2X2_4438 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf7), .B(w_mem_inst__abc_21378_n4640), .Y(w_mem_inst__abc_21378_n4641) );
  AND2X2 AND2X2_4439 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf27), .B(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_21378_n4644) );
  AND2X2 AND2X2_444 ( .A(_abc_15724_n1605), .B(_abc_15724_n1603_1), .Y(_abc_15724_n1606) );
  AND2X2 AND2X2_4440 ( .A(w_mem_inst__abc_21378_n3152_bF_buf6), .B(w_mem_inst_w_mem_9__24_), .Y(w_mem_inst__abc_21378_n4645) );
  AND2X2 AND2X2_4441 ( .A(round_ctr_rst_bF_buf3), .B(\block[248] ), .Y(w_mem_inst__abc_21378_n4646) );
  AND2X2 AND2X2_4442 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf6), .B(w_mem_inst__abc_21378_n4646), .Y(w_mem_inst__abc_21378_n4647) );
  AND2X2 AND2X2_4443 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf26), .B(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_21378_n4650) );
  AND2X2 AND2X2_4444 ( .A(w_mem_inst__abc_21378_n3152_bF_buf5), .B(w_mem_inst_w_mem_9__25_), .Y(w_mem_inst__abc_21378_n4651) );
  AND2X2 AND2X2_4445 ( .A(round_ctr_rst_bF_buf2), .B(\block[249] ), .Y(w_mem_inst__abc_21378_n4652) );
  AND2X2 AND2X2_4446 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf5), .B(w_mem_inst__abc_21378_n4652), .Y(w_mem_inst__abc_21378_n4653) );
  AND2X2 AND2X2_4447 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf25), .B(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_21378_n4656) );
  AND2X2 AND2X2_4448 ( .A(w_mem_inst__abc_21378_n3152_bF_buf4), .B(w_mem_inst_w_mem_9__26_), .Y(w_mem_inst__abc_21378_n4657) );
  AND2X2 AND2X2_4449 ( .A(round_ctr_rst_bF_buf1), .B(\block[250] ), .Y(w_mem_inst__abc_21378_n4658) );
  AND2X2 AND2X2_445 ( .A(_abc_15724_n1607), .B(_abc_15724_n1609_1), .Y(_abc_15724_n1610_1) );
  AND2X2 AND2X2_4450 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf4), .B(w_mem_inst__abc_21378_n4658), .Y(w_mem_inst__abc_21378_n4659) );
  AND2X2 AND2X2_4451 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf24), .B(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_21378_n4662) );
  AND2X2 AND2X2_4452 ( .A(w_mem_inst__abc_21378_n3152_bF_buf3), .B(w_mem_inst_w_mem_9__27_), .Y(w_mem_inst__abc_21378_n4663) );
  AND2X2 AND2X2_4453 ( .A(round_ctr_rst_bF_buf0), .B(\block[251] ), .Y(w_mem_inst__abc_21378_n4664) );
  AND2X2 AND2X2_4454 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf3), .B(w_mem_inst__abc_21378_n4664), .Y(w_mem_inst__abc_21378_n4665) );
  AND2X2 AND2X2_4455 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf23), .B(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_21378_n4668) );
  AND2X2 AND2X2_4456 ( .A(w_mem_inst__abc_21378_n3152_bF_buf2), .B(w_mem_inst_w_mem_9__28_), .Y(w_mem_inst__abc_21378_n4669) );
  AND2X2 AND2X2_4457 ( .A(round_ctr_rst_bF_buf63), .B(\block[252] ), .Y(w_mem_inst__abc_21378_n4670) );
  AND2X2 AND2X2_4458 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf2), .B(w_mem_inst__abc_21378_n4670), .Y(w_mem_inst__abc_21378_n4671) );
  AND2X2 AND2X2_4459 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf22), .B(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_21378_n4674) );
  AND2X2 AND2X2_446 ( .A(_abc_15724_n1610_1), .B(digest_update_bF_buf9), .Y(_abc_15724_n1611) );
  AND2X2 AND2X2_4460 ( .A(w_mem_inst__abc_21378_n3152_bF_buf1), .B(w_mem_inst_w_mem_9__29_), .Y(w_mem_inst__abc_21378_n4675) );
  AND2X2 AND2X2_4461 ( .A(round_ctr_rst_bF_buf62), .B(\block[253] ), .Y(w_mem_inst__abc_21378_n4676) );
  AND2X2 AND2X2_4462 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf1), .B(w_mem_inst__abc_21378_n4676), .Y(w_mem_inst__abc_21378_n4677) );
  AND2X2 AND2X2_4463 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf21), .B(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_21378_n4680) );
  AND2X2 AND2X2_4464 ( .A(w_mem_inst__abc_21378_n3152_bF_buf0), .B(w_mem_inst_w_mem_9__30_), .Y(w_mem_inst__abc_21378_n4681) );
  AND2X2 AND2X2_4465 ( .A(round_ctr_rst_bF_buf61), .B(\block[254] ), .Y(w_mem_inst__abc_21378_n4682) );
  AND2X2 AND2X2_4466 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf0), .B(w_mem_inst__abc_21378_n4682), .Y(w_mem_inst__abc_21378_n4683) );
  AND2X2 AND2X2_4467 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf20), .B(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_21378_n4686) );
  AND2X2 AND2X2_4468 ( .A(w_mem_inst__abc_21378_n3152_bF_buf63), .B(w_mem_inst_w_mem_9__31_), .Y(w_mem_inst__abc_21378_n4687) );
  AND2X2 AND2X2_4469 ( .A(round_ctr_rst_bF_buf60), .B(\block[255] ), .Y(w_mem_inst__abc_21378_n4688) );
  AND2X2 AND2X2_447 ( .A(_abc_15724_n1612), .B(_abc_15724_n850_bF_buf6), .Y(_abc_15724_n1613) );
  AND2X2 AND2X2_4470 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf63), .B(w_mem_inst__abc_21378_n4688), .Y(w_mem_inst__abc_21378_n4689) );
  AND2X2 AND2X2_4471 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf19), .B(w_mem_inst_w_mem_7__0_), .Y(w_mem_inst__abc_21378_n4692) );
  AND2X2 AND2X2_4472 ( .A(w_mem_inst__abc_21378_n3152_bF_buf62), .B(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_21378_n4693) );
  AND2X2 AND2X2_4473 ( .A(round_ctr_rst_bF_buf59), .B(\block[256] ), .Y(w_mem_inst__abc_21378_n4694) );
  AND2X2 AND2X2_4474 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf62), .B(w_mem_inst__abc_21378_n4694), .Y(w_mem_inst__abc_21378_n4695) );
  AND2X2 AND2X2_4475 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf18), .B(w_mem_inst_w_mem_7__1_), .Y(w_mem_inst__abc_21378_n4698) );
  AND2X2 AND2X2_4476 ( .A(w_mem_inst__abc_21378_n3152_bF_buf61), .B(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_21378_n4699) );
  AND2X2 AND2X2_4477 ( .A(round_ctr_rst_bF_buf58), .B(\block[257] ), .Y(w_mem_inst__abc_21378_n4700) );
  AND2X2 AND2X2_4478 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf61), .B(w_mem_inst__abc_21378_n4700), .Y(w_mem_inst__abc_21378_n4701) );
  AND2X2 AND2X2_4479 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf17), .B(w_mem_inst_w_mem_7__2_), .Y(w_mem_inst__abc_21378_n4704) );
  AND2X2 AND2X2_448 ( .A(_abc_15724_n907_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_72_), .Y(_abc_15724_n1615) );
  AND2X2 AND2X2_4480 ( .A(w_mem_inst__abc_21378_n3152_bF_buf60), .B(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_21378_n4705) );
  AND2X2 AND2X2_4481 ( .A(round_ctr_rst_bF_buf57), .B(\block[258] ), .Y(w_mem_inst__abc_21378_n4706) );
  AND2X2 AND2X2_4482 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf60), .B(w_mem_inst__abc_21378_n4706), .Y(w_mem_inst__abc_21378_n4707) );
  AND2X2 AND2X2_4483 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf16), .B(w_mem_inst_w_mem_7__3_), .Y(w_mem_inst__abc_21378_n4710) );
  AND2X2 AND2X2_4484 ( .A(w_mem_inst__abc_21378_n3152_bF_buf59), .B(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_21378_n4711) );
  AND2X2 AND2X2_4485 ( .A(round_ctr_rst_bF_buf56), .B(\block[259] ), .Y(w_mem_inst__abc_21378_n4712) );
  AND2X2 AND2X2_4486 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf59), .B(w_mem_inst__abc_21378_n4712), .Y(w_mem_inst__abc_21378_n4713) );
  AND2X2 AND2X2_4487 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf15), .B(w_mem_inst_w_mem_7__4_), .Y(w_mem_inst__abc_21378_n4716) );
  AND2X2 AND2X2_4488 ( .A(w_mem_inst__abc_21378_n3152_bF_buf58), .B(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_21378_n4717) );
  AND2X2 AND2X2_4489 ( .A(round_ctr_rst_bF_buf55), .B(\block[260] ), .Y(w_mem_inst__abc_21378_n4718) );
  AND2X2 AND2X2_449 ( .A(_auto_iopadmap_cc_313_execute_26059_72_), .B(c_reg_8_), .Y(_abc_15724_n1617_1) );
  AND2X2 AND2X2_4490 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf58), .B(w_mem_inst__abc_21378_n4718), .Y(w_mem_inst__abc_21378_n4719) );
  AND2X2 AND2X2_4491 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf14), .B(w_mem_inst_w_mem_7__5_), .Y(w_mem_inst__abc_21378_n4722) );
  AND2X2 AND2X2_4492 ( .A(w_mem_inst__abc_21378_n3152_bF_buf57), .B(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_21378_n4723) );
  AND2X2 AND2X2_4493 ( .A(round_ctr_rst_bF_buf54), .B(\block[261] ), .Y(w_mem_inst__abc_21378_n4724) );
  AND2X2 AND2X2_4494 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf57), .B(w_mem_inst__abc_21378_n4724), .Y(w_mem_inst__abc_21378_n4725) );
  AND2X2 AND2X2_4495 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf13), .B(w_mem_inst_w_mem_7__6_), .Y(w_mem_inst__abc_21378_n4728) );
  AND2X2 AND2X2_4496 ( .A(w_mem_inst__abc_21378_n3152_bF_buf56), .B(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_21378_n4729) );
  AND2X2 AND2X2_4497 ( .A(round_ctr_rst_bF_buf53), .B(\block[262] ), .Y(w_mem_inst__abc_21378_n4730) );
  AND2X2 AND2X2_4498 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf56), .B(w_mem_inst__abc_21378_n4730), .Y(w_mem_inst__abc_21378_n4731) );
  AND2X2 AND2X2_4499 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf12), .B(w_mem_inst_w_mem_7__7_), .Y(w_mem_inst__abc_21378_n4734) );
  AND2X2 AND2X2_45 ( .A(_abc_15724_n780_1), .B(_abc_15724_n781_1), .Y(_abc_15724_n782) );
  AND2X2 AND2X2_450 ( .A(_abc_15724_n1618), .B(_abc_15724_n1616_1), .Y(_abc_15724_n1619) );
  AND2X2 AND2X2_4500 ( .A(w_mem_inst__abc_21378_n3152_bF_buf55), .B(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_21378_n4735) );
  AND2X2 AND2X2_4501 ( .A(round_ctr_rst_bF_buf52), .B(\block[263] ), .Y(w_mem_inst__abc_21378_n4736) );
  AND2X2 AND2X2_4502 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf55), .B(w_mem_inst__abc_21378_n4736), .Y(w_mem_inst__abc_21378_n4737) );
  AND2X2 AND2X2_4503 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf11), .B(w_mem_inst_w_mem_7__8_), .Y(w_mem_inst__abc_21378_n4740) );
  AND2X2 AND2X2_4504 ( .A(w_mem_inst__abc_21378_n3152_bF_buf54), .B(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_21378_n4741) );
  AND2X2 AND2X2_4505 ( .A(round_ctr_rst_bF_buf51), .B(\block[264] ), .Y(w_mem_inst__abc_21378_n4742) );
  AND2X2 AND2X2_4506 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf54), .B(w_mem_inst__abc_21378_n4742), .Y(w_mem_inst__abc_21378_n4743) );
  AND2X2 AND2X2_4507 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf10), .B(w_mem_inst_w_mem_7__9_), .Y(w_mem_inst__abc_21378_n4746) );
  AND2X2 AND2X2_4508 ( .A(w_mem_inst__abc_21378_n3152_bF_buf53), .B(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_21378_n4747) );
  AND2X2 AND2X2_4509 ( .A(round_ctr_rst_bF_buf50), .B(\block[265] ), .Y(w_mem_inst__abc_21378_n4748) );
  AND2X2 AND2X2_451 ( .A(_abc_15724_n1591_1), .B(_abc_15724_n1605), .Y(_abc_15724_n1621) );
  AND2X2 AND2X2_4510 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf53), .B(w_mem_inst__abc_21378_n4748), .Y(w_mem_inst__abc_21378_n4749) );
  AND2X2 AND2X2_4511 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf9), .B(w_mem_inst_w_mem_7__10_), .Y(w_mem_inst__abc_21378_n4752) );
  AND2X2 AND2X2_4512 ( .A(w_mem_inst__abc_21378_n3152_bF_buf52), .B(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_21378_n4753) );
  AND2X2 AND2X2_4513 ( .A(round_ctr_rst_bF_buf49), .B(\block[266] ), .Y(w_mem_inst__abc_21378_n4754) );
  AND2X2 AND2X2_4514 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf52), .B(w_mem_inst__abc_21378_n4754), .Y(w_mem_inst__abc_21378_n4755) );
  AND2X2 AND2X2_4515 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf8), .B(w_mem_inst_w_mem_7__11_), .Y(w_mem_inst__abc_21378_n4758) );
  AND2X2 AND2X2_4516 ( .A(w_mem_inst__abc_21378_n3152_bF_buf51), .B(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_21378_n4759) );
  AND2X2 AND2X2_4517 ( .A(round_ctr_rst_bF_buf48), .B(\block[267] ), .Y(w_mem_inst__abc_21378_n4760) );
  AND2X2 AND2X2_4518 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf51), .B(w_mem_inst__abc_21378_n4760), .Y(w_mem_inst__abc_21378_n4761) );
  AND2X2 AND2X2_4519 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf7), .B(w_mem_inst_w_mem_7__12_), .Y(w_mem_inst__abc_21378_n4764) );
  AND2X2 AND2X2_452 ( .A(_abc_15724_n1595), .B(_abc_15724_n1621), .Y(_abc_15724_n1622) );
  AND2X2 AND2X2_4520 ( .A(w_mem_inst__abc_21378_n3152_bF_buf50), .B(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_21378_n4765) );
  AND2X2 AND2X2_4521 ( .A(round_ctr_rst_bF_buf47), .B(\block[268] ), .Y(w_mem_inst__abc_21378_n4766) );
  AND2X2 AND2X2_4522 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf50), .B(w_mem_inst__abc_21378_n4766), .Y(w_mem_inst__abc_21378_n4767) );
  AND2X2 AND2X2_4523 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf6), .B(w_mem_inst_w_mem_7__13_), .Y(w_mem_inst__abc_21378_n4770) );
  AND2X2 AND2X2_4524 ( .A(w_mem_inst__abc_21378_n3152_bF_buf49), .B(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_21378_n4771) );
  AND2X2 AND2X2_4525 ( .A(round_ctr_rst_bF_buf46), .B(\block[269] ), .Y(w_mem_inst__abc_21378_n4772) );
  AND2X2 AND2X2_4526 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf49), .B(w_mem_inst__abc_21378_n4772), .Y(w_mem_inst__abc_21378_n4773) );
  AND2X2 AND2X2_4527 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf5), .B(w_mem_inst_w_mem_7__14_), .Y(w_mem_inst__abc_21378_n4776) );
  AND2X2 AND2X2_4528 ( .A(w_mem_inst__abc_21378_n3152_bF_buf48), .B(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_21378_n4777) );
  AND2X2 AND2X2_4529 ( .A(round_ctr_rst_bF_buf45), .B(\block[270] ), .Y(w_mem_inst__abc_21378_n4778) );
  AND2X2 AND2X2_453 ( .A(_abc_15724_n1624_1), .B(_abc_15724_n1619), .Y(_abc_15724_n1626) );
  AND2X2 AND2X2_4530 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf48), .B(w_mem_inst__abc_21378_n4778), .Y(w_mem_inst__abc_21378_n4779) );
  AND2X2 AND2X2_4531 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf4), .B(w_mem_inst_w_mem_7__15_), .Y(w_mem_inst__abc_21378_n4782) );
  AND2X2 AND2X2_4532 ( .A(w_mem_inst__abc_21378_n3152_bF_buf47), .B(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_21378_n4783) );
  AND2X2 AND2X2_4533 ( .A(round_ctr_rst_bF_buf44), .B(\block[271] ), .Y(w_mem_inst__abc_21378_n4784) );
  AND2X2 AND2X2_4534 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf47), .B(w_mem_inst__abc_21378_n4784), .Y(w_mem_inst__abc_21378_n4785) );
  AND2X2 AND2X2_4535 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf3), .B(w_mem_inst_w_mem_7__16_), .Y(w_mem_inst__abc_21378_n4788) );
  AND2X2 AND2X2_4536 ( .A(w_mem_inst__abc_21378_n3152_bF_buf46), .B(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_21378_n4789) );
  AND2X2 AND2X2_4537 ( .A(round_ctr_rst_bF_buf43), .B(\block[272] ), .Y(w_mem_inst__abc_21378_n4790) );
  AND2X2 AND2X2_4538 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf46), .B(w_mem_inst__abc_21378_n4790), .Y(w_mem_inst__abc_21378_n4791) );
  AND2X2 AND2X2_4539 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf2), .B(w_mem_inst_w_mem_7__17_), .Y(w_mem_inst__abc_21378_n4794) );
  AND2X2 AND2X2_454 ( .A(_abc_15724_n1627), .B(_abc_15724_n1625), .Y(_abc_15724_n1628) );
  AND2X2 AND2X2_4540 ( .A(w_mem_inst__abc_21378_n3152_bF_buf45), .B(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_21378_n4795) );
  AND2X2 AND2X2_4541 ( .A(round_ctr_rst_bF_buf42), .B(\block[273] ), .Y(w_mem_inst__abc_21378_n4796) );
  AND2X2 AND2X2_4542 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf45), .B(w_mem_inst__abc_21378_n4796), .Y(w_mem_inst__abc_21378_n4797) );
  AND2X2 AND2X2_4543 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf1), .B(w_mem_inst_w_mem_7__18_), .Y(w_mem_inst__abc_21378_n4800) );
  AND2X2 AND2X2_4544 ( .A(w_mem_inst__abc_21378_n3152_bF_buf44), .B(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_21378_n4801) );
  AND2X2 AND2X2_4545 ( .A(round_ctr_rst_bF_buf41), .B(\block[274] ), .Y(w_mem_inst__abc_21378_n4802) );
  AND2X2 AND2X2_4546 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf44), .B(w_mem_inst__abc_21378_n4802), .Y(w_mem_inst__abc_21378_n4803) );
  AND2X2 AND2X2_4547 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf0), .B(w_mem_inst_w_mem_7__19_), .Y(w_mem_inst__abc_21378_n4806) );
  AND2X2 AND2X2_4548 ( .A(w_mem_inst__abc_21378_n3152_bF_buf43), .B(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_21378_n4807) );
  AND2X2 AND2X2_4549 ( .A(round_ctr_rst_bF_buf40), .B(\block[275] ), .Y(w_mem_inst__abc_21378_n4808) );
  AND2X2 AND2X2_455 ( .A(_abc_15724_n1628), .B(digest_update_bF_buf8), .Y(_abc_15724_n1629) );
  AND2X2 AND2X2_4550 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf43), .B(w_mem_inst__abc_21378_n4808), .Y(w_mem_inst__abc_21378_n4809) );
  AND2X2 AND2X2_4551 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf60), .B(w_mem_inst_w_mem_7__20_), .Y(w_mem_inst__abc_21378_n4812) );
  AND2X2 AND2X2_4552 ( .A(w_mem_inst__abc_21378_n3152_bF_buf42), .B(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_21378_n4813) );
  AND2X2 AND2X2_4553 ( .A(round_ctr_rst_bF_buf39), .B(\block[276] ), .Y(w_mem_inst__abc_21378_n4814) );
  AND2X2 AND2X2_4554 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf42), .B(w_mem_inst__abc_21378_n4814), .Y(w_mem_inst__abc_21378_n4815) );
  AND2X2 AND2X2_4555 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf59), .B(w_mem_inst_w_mem_7__21_), .Y(w_mem_inst__abc_21378_n4818) );
  AND2X2 AND2X2_4556 ( .A(w_mem_inst__abc_21378_n3152_bF_buf41), .B(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_21378_n4819) );
  AND2X2 AND2X2_4557 ( .A(round_ctr_rst_bF_buf38), .B(\block[277] ), .Y(w_mem_inst__abc_21378_n4820) );
  AND2X2 AND2X2_4558 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf41), .B(w_mem_inst__abc_21378_n4820), .Y(w_mem_inst__abc_21378_n4821) );
  AND2X2 AND2X2_4559 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf58), .B(w_mem_inst_w_mem_7__22_), .Y(w_mem_inst__abc_21378_n4824) );
  AND2X2 AND2X2_456 ( .A(_auto_iopadmap_cc_313_execute_26059_73_), .B(c_reg_9_), .Y(_abc_15724_n1632) );
  AND2X2 AND2X2_4560 ( .A(w_mem_inst__abc_21378_n3152_bF_buf40), .B(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_21378_n4825) );
  AND2X2 AND2X2_4561 ( .A(round_ctr_rst_bF_buf37), .B(\block[278] ), .Y(w_mem_inst__abc_21378_n4826) );
  AND2X2 AND2X2_4562 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf40), .B(w_mem_inst__abc_21378_n4826), .Y(w_mem_inst__abc_21378_n4827) );
  AND2X2 AND2X2_4563 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf57), .B(w_mem_inst_w_mem_7__23_), .Y(w_mem_inst__abc_21378_n4830) );
  AND2X2 AND2X2_4564 ( .A(w_mem_inst__abc_21378_n3152_bF_buf39), .B(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_21378_n4831) );
  AND2X2 AND2X2_4565 ( .A(round_ctr_rst_bF_buf36), .B(\block[279] ), .Y(w_mem_inst__abc_21378_n4832) );
  AND2X2 AND2X2_4566 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf39), .B(w_mem_inst__abc_21378_n4832), .Y(w_mem_inst__abc_21378_n4833) );
  AND2X2 AND2X2_4567 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf56), .B(w_mem_inst_w_mem_7__24_), .Y(w_mem_inst__abc_21378_n4836) );
  AND2X2 AND2X2_4568 ( .A(w_mem_inst__abc_21378_n3152_bF_buf38), .B(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_21378_n4837) );
  AND2X2 AND2X2_4569 ( .A(round_ctr_rst_bF_buf35), .B(\block[280] ), .Y(w_mem_inst__abc_21378_n4838) );
  AND2X2 AND2X2_457 ( .A(_abc_15724_n1633_1), .B(_abc_15724_n1631_1), .Y(_abc_15724_n1634) );
  AND2X2 AND2X2_4570 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf38), .B(w_mem_inst__abc_21378_n4838), .Y(w_mem_inst__abc_21378_n4839) );
  AND2X2 AND2X2_4571 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf55), .B(w_mem_inst_w_mem_7__25_), .Y(w_mem_inst__abc_21378_n4842) );
  AND2X2 AND2X2_4572 ( .A(w_mem_inst__abc_21378_n3152_bF_buf37), .B(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_21378_n4843) );
  AND2X2 AND2X2_4573 ( .A(round_ctr_rst_bF_buf34), .B(\block[281] ), .Y(w_mem_inst__abc_21378_n4844) );
  AND2X2 AND2X2_4574 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf37), .B(w_mem_inst__abc_21378_n4844), .Y(w_mem_inst__abc_21378_n4845) );
  AND2X2 AND2X2_4575 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf54), .B(w_mem_inst_w_mem_7__26_), .Y(w_mem_inst__abc_21378_n4848) );
  AND2X2 AND2X2_4576 ( .A(w_mem_inst__abc_21378_n3152_bF_buf36), .B(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_21378_n4849) );
  AND2X2 AND2X2_4577 ( .A(round_ctr_rst_bF_buf33), .B(\block[282] ), .Y(w_mem_inst__abc_21378_n4850) );
  AND2X2 AND2X2_4578 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf36), .B(w_mem_inst__abc_21378_n4850), .Y(w_mem_inst__abc_21378_n4851) );
  AND2X2 AND2X2_4579 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf53), .B(w_mem_inst_w_mem_7__27_), .Y(w_mem_inst__abc_21378_n4854) );
  AND2X2 AND2X2_458 ( .A(_abc_15724_n1627), .B(_abc_15724_n1618), .Y(_abc_15724_n1635) );
  AND2X2 AND2X2_4580 ( .A(w_mem_inst__abc_21378_n3152_bF_buf35), .B(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_21378_n4855) );
  AND2X2 AND2X2_4581 ( .A(round_ctr_rst_bF_buf32), .B(\block[283] ), .Y(w_mem_inst__abc_21378_n4856) );
  AND2X2 AND2X2_4582 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf35), .B(w_mem_inst__abc_21378_n4856), .Y(w_mem_inst__abc_21378_n4857) );
  AND2X2 AND2X2_4583 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf52), .B(w_mem_inst_w_mem_7__28_), .Y(w_mem_inst__abc_21378_n4860) );
  AND2X2 AND2X2_4584 ( .A(w_mem_inst__abc_21378_n3152_bF_buf34), .B(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_21378_n4861) );
  AND2X2 AND2X2_4585 ( .A(round_ctr_rst_bF_buf31), .B(\block[284] ), .Y(w_mem_inst__abc_21378_n4862) );
  AND2X2 AND2X2_4586 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf34), .B(w_mem_inst__abc_21378_n4862), .Y(w_mem_inst__abc_21378_n4863) );
  AND2X2 AND2X2_4587 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf51), .B(w_mem_inst_w_mem_7__29_), .Y(w_mem_inst__abc_21378_n4866) );
  AND2X2 AND2X2_4588 ( .A(w_mem_inst__abc_21378_n3152_bF_buf33), .B(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_21378_n4867) );
  AND2X2 AND2X2_4589 ( .A(round_ctr_rst_bF_buf30), .B(\block[285] ), .Y(w_mem_inst__abc_21378_n4868) );
  AND2X2 AND2X2_459 ( .A(_abc_15724_n1636_1), .B(_abc_15724_n1634), .Y(_abc_15724_n1638) );
  AND2X2 AND2X2_4590 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf33), .B(w_mem_inst__abc_21378_n4868), .Y(w_mem_inst__abc_21378_n4869) );
  AND2X2 AND2X2_4591 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf50), .B(w_mem_inst_w_mem_7__30_), .Y(w_mem_inst__abc_21378_n4872) );
  AND2X2 AND2X2_4592 ( .A(w_mem_inst__abc_21378_n3152_bF_buf32), .B(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_21378_n4873) );
  AND2X2 AND2X2_4593 ( .A(round_ctr_rst_bF_buf29), .B(\block[286] ), .Y(w_mem_inst__abc_21378_n4874) );
  AND2X2 AND2X2_4594 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf32), .B(w_mem_inst__abc_21378_n4874), .Y(w_mem_inst__abc_21378_n4875) );
  AND2X2 AND2X2_4595 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf49), .B(w_mem_inst_w_mem_7__31_), .Y(w_mem_inst__abc_21378_n4878) );
  AND2X2 AND2X2_4596 ( .A(w_mem_inst__abc_21378_n3152_bF_buf31), .B(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_21378_n4879) );
  AND2X2 AND2X2_4597 ( .A(round_ctr_rst_bF_buf28), .B(\block[287] ), .Y(w_mem_inst__abc_21378_n4880) );
  AND2X2 AND2X2_4598 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf31), .B(w_mem_inst__abc_21378_n4880), .Y(w_mem_inst__abc_21378_n4881) );
  AND2X2 AND2X2_4599 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf48), .B(w_mem_inst_w_mem_6__0_), .Y(w_mem_inst__abc_21378_n4884) );
  AND2X2 AND2X2_46 ( .A(_abc_15724_n779_1), .B(_abc_15724_n782), .Y(_abc_15724_n783) );
  AND2X2 AND2X2_460 ( .A(_abc_15724_n1639_1), .B(_abc_15724_n1637_1), .Y(_abc_15724_n1640) );
  AND2X2 AND2X2_4600 ( .A(w_mem_inst__abc_21378_n3152_bF_buf30), .B(w_mem_inst_w_mem_7__0_), .Y(w_mem_inst__abc_21378_n4885) );
  AND2X2 AND2X2_4601 ( .A(round_ctr_rst_bF_buf27), .B(\block[288] ), .Y(w_mem_inst__abc_21378_n4886) );
  AND2X2 AND2X2_4602 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf30), .B(w_mem_inst__abc_21378_n4886), .Y(w_mem_inst__abc_21378_n4887) );
  AND2X2 AND2X2_4603 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf47), .B(w_mem_inst_w_mem_6__1_), .Y(w_mem_inst__abc_21378_n4890) );
  AND2X2 AND2X2_4604 ( .A(w_mem_inst__abc_21378_n3152_bF_buf29), .B(w_mem_inst_w_mem_7__1_), .Y(w_mem_inst__abc_21378_n4891) );
  AND2X2 AND2X2_4605 ( .A(round_ctr_rst_bF_buf26), .B(\block[289] ), .Y(w_mem_inst__abc_21378_n4892) );
  AND2X2 AND2X2_4606 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf29), .B(w_mem_inst__abc_21378_n4892), .Y(w_mem_inst__abc_21378_n4893) );
  AND2X2 AND2X2_4607 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf46), .B(w_mem_inst_w_mem_6__2_), .Y(w_mem_inst__abc_21378_n4896) );
  AND2X2 AND2X2_4608 ( .A(w_mem_inst__abc_21378_n3152_bF_buf28), .B(w_mem_inst_w_mem_7__2_), .Y(w_mem_inst__abc_21378_n4897) );
  AND2X2 AND2X2_4609 ( .A(round_ctr_rst_bF_buf25), .B(\block[290] ), .Y(w_mem_inst__abc_21378_n4898) );
  AND2X2 AND2X2_461 ( .A(_abc_15724_n1640), .B(digest_update_bF_buf7), .Y(_abc_15724_n1641) );
  AND2X2 AND2X2_4610 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf28), .B(w_mem_inst__abc_21378_n4898), .Y(w_mem_inst__abc_21378_n4899) );
  AND2X2 AND2X2_4611 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf45), .B(w_mem_inst_w_mem_6__3_), .Y(w_mem_inst__abc_21378_n4902) );
  AND2X2 AND2X2_4612 ( .A(w_mem_inst__abc_21378_n3152_bF_buf27), .B(w_mem_inst_w_mem_7__3_), .Y(w_mem_inst__abc_21378_n4903) );
  AND2X2 AND2X2_4613 ( .A(round_ctr_rst_bF_buf24), .B(\block[291] ), .Y(w_mem_inst__abc_21378_n4904) );
  AND2X2 AND2X2_4614 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf27), .B(w_mem_inst__abc_21378_n4904), .Y(w_mem_inst__abc_21378_n4905) );
  AND2X2 AND2X2_4615 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf44), .B(w_mem_inst_w_mem_6__4_), .Y(w_mem_inst__abc_21378_n4908) );
  AND2X2 AND2X2_4616 ( .A(w_mem_inst__abc_21378_n3152_bF_buf26), .B(w_mem_inst_w_mem_7__4_), .Y(w_mem_inst__abc_21378_n4909) );
  AND2X2 AND2X2_4617 ( .A(round_ctr_rst_bF_buf23), .B(\block[292] ), .Y(w_mem_inst__abc_21378_n4910) );
  AND2X2 AND2X2_4618 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf26), .B(w_mem_inst__abc_21378_n4910), .Y(w_mem_inst__abc_21378_n4911) );
  AND2X2 AND2X2_4619 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf43), .B(w_mem_inst_w_mem_6__5_), .Y(w_mem_inst__abc_21378_n4914) );
  AND2X2 AND2X2_462 ( .A(_abc_15724_n907_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_73_), .Y(_abc_15724_n1642_1) );
  AND2X2 AND2X2_4620 ( .A(w_mem_inst__abc_21378_n3152_bF_buf25), .B(w_mem_inst_w_mem_7__5_), .Y(w_mem_inst__abc_21378_n4915) );
  AND2X2 AND2X2_4621 ( .A(round_ctr_rst_bF_buf22), .B(\block[293] ), .Y(w_mem_inst__abc_21378_n4916) );
  AND2X2 AND2X2_4622 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf25), .B(w_mem_inst__abc_21378_n4916), .Y(w_mem_inst__abc_21378_n4917) );
  AND2X2 AND2X2_4623 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf42), .B(w_mem_inst_w_mem_6__6_), .Y(w_mem_inst__abc_21378_n4920) );
  AND2X2 AND2X2_4624 ( .A(w_mem_inst__abc_21378_n3152_bF_buf24), .B(w_mem_inst_w_mem_7__6_), .Y(w_mem_inst__abc_21378_n4921) );
  AND2X2 AND2X2_4625 ( .A(round_ctr_rst_bF_buf21), .B(\block[294] ), .Y(w_mem_inst__abc_21378_n4922) );
  AND2X2 AND2X2_4626 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf24), .B(w_mem_inst__abc_21378_n4922), .Y(w_mem_inst__abc_21378_n4923) );
  AND2X2 AND2X2_4627 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf41), .B(w_mem_inst_w_mem_6__7_), .Y(w_mem_inst__abc_21378_n4926) );
  AND2X2 AND2X2_4628 ( .A(w_mem_inst__abc_21378_n3152_bF_buf23), .B(w_mem_inst_w_mem_7__7_), .Y(w_mem_inst__abc_21378_n4927) );
  AND2X2 AND2X2_4629 ( .A(round_ctr_rst_bF_buf20), .B(\block[295] ), .Y(w_mem_inst__abc_21378_n4928) );
  AND2X2 AND2X2_463 ( .A(_abc_15724_n1639_1), .B(_abc_15724_n1633_1), .Y(_abc_15724_n1644) );
  AND2X2 AND2X2_4630 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf23), .B(w_mem_inst__abc_21378_n4928), .Y(w_mem_inst__abc_21378_n4929) );
  AND2X2 AND2X2_4631 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf40), .B(w_mem_inst_w_mem_6__8_), .Y(w_mem_inst__abc_21378_n4932) );
  AND2X2 AND2X2_4632 ( .A(w_mem_inst__abc_21378_n3152_bF_buf22), .B(w_mem_inst_w_mem_7__8_), .Y(w_mem_inst__abc_21378_n4933) );
  AND2X2 AND2X2_4633 ( .A(round_ctr_rst_bF_buf19), .B(\block[296] ), .Y(w_mem_inst__abc_21378_n4934) );
  AND2X2 AND2X2_4634 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf22), .B(w_mem_inst__abc_21378_n4934), .Y(w_mem_inst__abc_21378_n4935) );
  AND2X2 AND2X2_4635 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf39), .B(w_mem_inst_w_mem_6__9_), .Y(w_mem_inst__abc_21378_n4938) );
  AND2X2 AND2X2_4636 ( .A(w_mem_inst__abc_21378_n3152_bF_buf21), .B(w_mem_inst_w_mem_7__9_), .Y(w_mem_inst__abc_21378_n4939) );
  AND2X2 AND2X2_4637 ( .A(round_ctr_rst_bF_buf18), .B(\block[297] ), .Y(w_mem_inst__abc_21378_n4940) );
  AND2X2 AND2X2_4638 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf21), .B(w_mem_inst__abc_21378_n4940), .Y(w_mem_inst__abc_21378_n4941) );
  AND2X2 AND2X2_4639 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf38), .B(w_mem_inst_w_mem_6__10_), .Y(w_mem_inst__abc_21378_n4944) );
  AND2X2 AND2X2_464 ( .A(_auto_iopadmap_cc_313_execute_26059_74_), .B(c_reg_10_), .Y(_abc_15724_n1647) );
  AND2X2 AND2X2_4640 ( .A(w_mem_inst__abc_21378_n3152_bF_buf20), .B(w_mem_inst_w_mem_7__10_), .Y(w_mem_inst__abc_21378_n4945) );
  AND2X2 AND2X2_4641 ( .A(round_ctr_rst_bF_buf17), .B(\block[298] ), .Y(w_mem_inst__abc_21378_n4946) );
  AND2X2 AND2X2_4642 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf20), .B(w_mem_inst__abc_21378_n4946), .Y(w_mem_inst__abc_21378_n4947) );
  AND2X2 AND2X2_4643 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf37), .B(w_mem_inst_w_mem_6__11_), .Y(w_mem_inst__abc_21378_n4950) );
  AND2X2 AND2X2_4644 ( .A(w_mem_inst__abc_21378_n3152_bF_buf19), .B(w_mem_inst_w_mem_7__11_), .Y(w_mem_inst__abc_21378_n4951) );
  AND2X2 AND2X2_4645 ( .A(round_ctr_rst_bF_buf16), .B(\block[299] ), .Y(w_mem_inst__abc_21378_n4952) );
  AND2X2 AND2X2_4646 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf19), .B(w_mem_inst__abc_21378_n4952), .Y(w_mem_inst__abc_21378_n4953) );
  AND2X2 AND2X2_4647 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf36), .B(w_mem_inst_w_mem_6__12_), .Y(w_mem_inst__abc_21378_n4956) );
  AND2X2 AND2X2_4648 ( .A(w_mem_inst__abc_21378_n3152_bF_buf18), .B(w_mem_inst_w_mem_7__12_), .Y(w_mem_inst__abc_21378_n4957) );
  AND2X2 AND2X2_4649 ( .A(round_ctr_rst_bF_buf15), .B(\block[300] ), .Y(w_mem_inst__abc_21378_n4958) );
  AND2X2 AND2X2_465 ( .A(_abc_15724_n1648_1), .B(_abc_15724_n1646), .Y(_abc_15724_n1649_1) );
  AND2X2 AND2X2_4650 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf18), .B(w_mem_inst__abc_21378_n4958), .Y(w_mem_inst__abc_21378_n4959) );
  AND2X2 AND2X2_4651 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf35), .B(w_mem_inst_w_mem_6__13_), .Y(w_mem_inst__abc_21378_n4962) );
  AND2X2 AND2X2_4652 ( .A(w_mem_inst__abc_21378_n3152_bF_buf17), .B(w_mem_inst_w_mem_7__13_), .Y(w_mem_inst__abc_21378_n4963) );
  AND2X2 AND2X2_4653 ( .A(round_ctr_rst_bF_buf14), .B(\block[301] ), .Y(w_mem_inst__abc_21378_n4964) );
  AND2X2 AND2X2_4654 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf17), .B(w_mem_inst__abc_21378_n4964), .Y(w_mem_inst__abc_21378_n4965) );
  AND2X2 AND2X2_4655 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf34), .B(w_mem_inst_w_mem_6__14_), .Y(w_mem_inst__abc_21378_n4968) );
  AND2X2 AND2X2_4656 ( .A(w_mem_inst__abc_21378_n3152_bF_buf16), .B(w_mem_inst_w_mem_7__14_), .Y(w_mem_inst__abc_21378_n4969) );
  AND2X2 AND2X2_4657 ( .A(round_ctr_rst_bF_buf13), .B(\block[302] ), .Y(w_mem_inst__abc_21378_n4970) );
  AND2X2 AND2X2_4658 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf16), .B(w_mem_inst__abc_21378_n4970), .Y(w_mem_inst__abc_21378_n4971) );
  AND2X2 AND2X2_4659 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf33), .B(w_mem_inst_w_mem_6__15_), .Y(w_mem_inst__abc_21378_n4974) );
  AND2X2 AND2X2_466 ( .A(_abc_15724_n1645_1), .B(_abc_15724_n1649_1), .Y(_abc_15724_n1651) );
  AND2X2 AND2X2_4660 ( .A(w_mem_inst__abc_21378_n3152_bF_buf15), .B(w_mem_inst_w_mem_7__15_), .Y(w_mem_inst__abc_21378_n4975) );
  AND2X2 AND2X2_4661 ( .A(round_ctr_rst_bF_buf12), .B(\block[303] ), .Y(w_mem_inst__abc_21378_n4976) );
  AND2X2 AND2X2_4662 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf15), .B(w_mem_inst__abc_21378_n4976), .Y(w_mem_inst__abc_21378_n4977) );
  AND2X2 AND2X2_4663 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf32), .B(w_mem_inst_w_mem_6__16_), .Y(w_mem_inst__abc_21378_n4980) );
  AND2X2 AND2X2_4664 ( .A(w_mem_inst__abc_21378_n3152_bF_buf14), .B(w_mem_inst_w_mem_7__16_), .Y(w_mem_inst__abc_21378_n4981) );
  AND2X2 AND2X2_4665 ( .A(round_ctr_rst_bF_buf11), .B(\block[304] ), .Y(w_mem_inst__abc_21378_n4982) );
  AND2X2 AND2X2_4666 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf14), .B(w_mem_inst__abc_21378_n4982), .Y(w_mem_inst__abc_21378_n4983) );
  AND2X2 AND2X2_4667 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf31), .B(w_mem_inst_w_mem_6__17_), .Y(w_mem_inst__abc_21378_n4986) );
  AND2X2 AND2X2_4668 ( .A(w_mem_inst__abc_21378_n3152_bF_buf13), .B(w_mem_inst_w_mem_7__17_), .Y(w_mem_inst__abc_21378_n4987) );
  AND2X2 AND2X2_4669 ( .A(round_ctr_rst_bF_buf10), .B(\block[305] ), .Y(w_mem_inst__abc_21378_n4988) );
  AND2X2 AND2X2_467 ( .A(_abc_15724_n1652), .B(_abc_15724_n1650), .Y(_abc_15724_n1653) );
  AND2X2 AND2X2_4670 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf13), .B(w_mem_inst__abc_21378_n4988), .Y(w_mem_inst__abc_21378_n4989) );
  AND2X2 AND2X2_4671 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf30), .B(w_mem_inst_w_mem_6__18_), .Y(w_mem_inst__abc_21378_n4992) );
  AND2X2 AND2X2_4672 ( .A(w_mem_inst__abc_21378_n3152_bF_buf12), .B(w_mem_inst_w_mem_7__18_), .Y(w_mem_inst__abc_21378_n4993) );
  AND2X2 AND2X2_4673 ( .A(round_ctr_rst_bF_buf9), .B(\block[306] ), .Y(w_mem_inst__abc_21378_n4994) );
  AND2X2 AND2X2_4674 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf12), .B(w_mem_inst__abc_21378_n4994), .Y(w_mem_inst__abc_21378_n4995) );
  AND2X2 AND2X2_4675 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf29), .B(w_mem_inst_w_mem_6__19_), .Y(w_mem_inst__abc_21378_n4998) );
  AND2X2 AND2X2_4676 ( .A(w_mem_inst__abc_21378_n3152_bF_buf11), .B(w_mem_inst_w_mem_7__19_), .Y(w_mem_inst__abc_21378_n4999) );
  AND2X2 AND2X2_4677 ( .A(round_ctr_rst_bF_buf8), .B(\block[307] ), .Y(w_mem_inst__abc_21378_n5000) );
  AND2X2 AND2X2_4678 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf11), .B(w_mem_inst__abc_21378_n5000), .Y(w_mem_inst__abc_21378_n5001) );
  AND2X2 AND2X2_4679 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf28), .B(w_mem_inst_w_mem_6__20_), .Y(w_mem_inst__abc_21378_n5004) );
  AND2X2 AND2X2_468 ( .A(_abc_15724_n1653), .B(digest_update_bF_buf6), .Y(_abc_15724_n1654) );
  AND2X2 AND2X2_4680 ( .A(w_mem_inst__abc_21378_n3152_bF_buf10), .B(w_mem_inst_w_mem_7__20_), .Y(w_mem_inst__abc_21378_n5005) );
  AND2X2 AND2X2_4681 ( .A(round_ctr_rst_bF_buf7), .B(\block[308] ), .Y(w_mem_inst__abc_21378_n5006) );
  AND2X2 AND2X2_4682 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf10), .B(w_mem_inst__abc_21378_n5006), .Y(w_mem_inst__abc_21378_n5007) );
  AND2X2 AND2X2_4683 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf27), .B(w_mem_inst_w_mem_6__21_), .Y(w_mem_inst__abc_21378_n5010) );
  AND2X2 AND2X2_4684 ( .A(w_mem_inst__abc_21378_n3152_bF_buf9), .B(w_mem_inst_w_mem_7__21_), .Y(w_mem_inst__abc_21378_n5011) );
  AND2X2 AND2X2_4685 ( .A(round_ctr_rst_bF_buf6), .B(\block[309] ), .Y(w_mem_inst__abc_21378_n5012) );
  AND2X2 AND2X2_4686 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf9), .B(w_mem_inst__abc_21378_n5012), .Y(w_mem_inst__abc_21378_n5013) );
  AND2X2 AND2X2_4687 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf26), .B(w_mem_inst_w_mem_6__22_), .Y(w_mem_inst__abc_21378_n5016) );
  AND2X2 AND2X2_4688 ( .A(w_mem_inst__abc_21378_n3152_bF_buf8), .B(w_mem_inst_w_mem_7__22_), .Y(w_mem_inst__abc_21378_n5017) );
  AND2X2 AND2X2_4689 ( .A(round_ctr_rst_bF_buf5), .B(\block[310] ), .Y(w_mem_inst__abc_21378_n5018) );
  AND2X2 AND2X2_469 ( .A(_abc_15724_n1655_1), .B(_abc_15724_n850_bF_buf5), .Y(_abc_15724_n1656_1) );
  AND2X2 AND2X2_4690 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf8), .B(w_mem_inst__abc_21378_n5018), .Y(w_mem_inst__abc_21378_n5019) );
  AND2X2 AND2X2_4691 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf25), .B(w_mem_inst_w_mem_6__23_), .Y(w_mem_inst__abc_21378_n5022) );
  AND2X2 AND2X2_4692 ( .A(w_mem_inst__abc_21378_n3152_bF_buf7), .B(w_mem_inst_w_mem_7__23_), .Y(w_mem_inst__abc_21378_n5023) );
  AND2X2 AND2X2_4693 ( .A(round_ctr_rst_bF_buf4), .B(\block[311] ), .Y(w_mem_inst__abc_21378_n5024) );
  AND2X2 AND2X2_4694 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf7), .B(w_mem_inst__abc_21378_n5024), .Y(w_mem_inst__abc_21378_n5025) );
  AND2X2 AND2X2_4695 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf24), .B(w_mem_inst_w_mem_6__24_), .Y(w_mem_inst__abc_21378_n5028) );
  AND2X2 AND2X2_4696 ( .A(w_mem_inst__abc_21378_n3152_bF_buf6), .B(w_mem_inst_w_mem_7__24_), .Y(w_mem_inst__abc_21378_n5029) );
  AND2X2 AND2X2_4697 ( .A(round_ctr_rst_bF_buf3), .B(\block[312] ), .Y(w_mem_inst__abc_21378_n5030) );
  AND2X2 AND2X2_4698 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf6), .B(w_mem_inst__abc_21378_n5030), .Y(w_mem_inst__abc_21378_n5031) );
  AND2X2 AND2X2_4699 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf23), .B(w_mem_inst_w_mem_6__25_), .Y(w_mem_inst__abc_21378_n5034) );
  AND2X2 AND2X2_47 ( .A(_auto_iopadmap_cc_313_execute_26059_5_), .B(e_reg_5_), .Y(_abc_15724_n784) );
  AND2X2 AND2X2_470 ( .A(_abc_15724_n1652), .B(_abc_15724_n1648_1), .Y(_abc_15724_n1658_1) );
  AND2X2 AND2X2_4700 ( .A(w_mem_inst__abc_21378_n3152_bF_buf5), .B(w_mem_inst_w_mem_7__25_), .Y(w_mem_inst__abc_21378_n5035) );
  AND2X2 AND2X2_4701 ( .A(round_ctr_rst_bF_buf2), .B(\block[313] ), .Y(w_mem_inst__abc_21378_n5036) );
  AND2X2 AND2X2_4702 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf5), .B(w_mem_inst__abc_21378_n5036), .Y(w_mem_inst__abc_21378_n5037) );
  AND2X2 AND2X2_4703 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf22), .B(w_mem_inst_w_mem_6__26_), .Y(w_mem_inst__abc_21378_n5040) );
  AND2X2 AND2X2_4704 ( .A(w_mem_inst__abc_21378_n3152_bF_buf4), .B(w_mem_inst_w_mem_7__26_), .Y(w_mem_inst__abc_21378_n5041) );
  AND2X2 AND2X2_4705 ( .A(round_ctr_rst_bF_buf1), .B(\block[314] ), .Y(w_mem_inst__abc_21378_n5042) );
  AND2X2 AND2X2_4706 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf4), .B(w_mem_inst__abc_21378_n5042), .Y(w_mem_inst__abc_21378_n5043) );
  AND2X2 AND2X2_4707 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf21), .B(w_mem_inst_w_mem_6__27_), .Y(w_mem_inst__abc_21378_n5046) );
  AND2X2 AND2X2_4708 ( .A(w_mem_inst__abc_21378_n3152_bF_buf3), .B(w_mem_inst_w_mem_7__27_), .Y(w_mem_inst__abc_21378_n5047) );
  AND2X2 AND2X2_4709 ( .A(round_ctr_rst_bF_buf0), .B(\block[315] ), .Y(w_mem_inst__abc_21378_n5048) );
  AND2X2 AND2X2_471 ( .A(_auto_iopadmap_cc_313_execute_26059_75_), .B(c_reg_11_), .Y(_abc_15724_n1660) );
  AND2X2 AND2X2_4710 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf3), .B(w_mem_inst__abc_21378_n5048), .Y(w_mem_inst__abc_21378_n5049) );
  AND2X2 AND2X2_4711 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf20), .B(w_mem_inst_w_mem_6__28_), .Y(w_mem_inst__abc_21378_n5052) );
  AND2X2 AND2X2_4712 ( .A(w_mem_inst__abc_21378_n3152_bF_buf2), .B(w_mem_inst_w_mem_7__28_), .Y(w_mem_inst__abc_21378_n5053) );
  AND2X2 AND2X2_4713 ( .A(round_ctr_rst_bF_buf63), .B(\block[316] ), .Y(w_mem_inst__abc_21378_n5054) );
  AND2X2 AND2X2_4714 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf2), .B(w_mem_inst__abc_21378_n5054), .Y(w_mem_inst__abc_21378_n5055) );
  AND2X2 AND2X2_4715 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf19), .B(w_mem_inst_w_mem_6__29_), .Y(w_mem_inst__abc_21378_n5058) );
  AND2X2 AND2X2_4716 ( .A(w_mem_inst__abc_21378_n3152_bF_buf1), .B(w_mem_inst_w_mem_7__29_), .Y(w_mem_inst__abc_21378_n5059) );
  AND2X2 AND2X2_4717 ( .A(round_ctr_rst_bF_buf62), .B(\block[317] ), .Y(w_mem_inst__abc_21378_n5060) );
  AND2X2 AND2X2_4718 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf1), .B(w_mem_inst__abc_21378_n5060), .Y(w_mem_inst__abc_21378_n5061) );
  AND2X2 AND2X2_4719 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf18), .B(w_mem_inst_w_mem_6__30_), .Y(w_mem_inst__abc_21378_n5064) );
  AND2X2 AND2X2_472 ( .A(_abc_15724_n1661_1), .B(_abc_15724_n1659), .Y(_abc_15724_n1662_1) );
  AND2X2 AND2X2_4720 ( .A(w_mem_inst__abc_21378_n3152_bF_buf0), .B(w_mem_inst_w_mem_7__30_), .Y(w_mem_inst__abc_21378_n5065) );
  AND2X2 AND2X2_4721 ( .A(round_ctr_rst_bF_buf61), .B(\block[318] ), .Y(w_mem_inst__abc_21378_n5066) );
  AND2X2 AND2X2_4722 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf0), .B(w_mem_inst__abc_21378_n5066), .Y(w_mem_inst__abc_21378_n5067) );
  AND2X2 AND2X2_4723 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf17), .B(w_mem_inst_w_mem_6__31_), .Y(w_mem_inst__abc_21378_n5070) );
  AND2X2 AND2X2_4724 ( .A(w_mem_inst__abc_21378_n3152_bF_buf63), .B(w_mem_inst_w_mem_7__31_), .Y(w_mem_inst__abc_21378_n5071) );
  AND2X2 AND2X2_4725 ( .A(round_ctr_rst_bF_buf60), .B(\block[319] ), .Y(w_mem_inst__abc_21378_n5072) );
  AND2X2 AND2X2_4726 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf63), .B(w_mem_inst__abc_21378_n5072), .Y(w_mem_inst__abc_21378_n5073) );
  AND2X2 AND2X2_4727 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf16), .B(w_mem_inst_w_mem_5__0_), .Y(w_mem_inst__abc_21378_n5076) );
  AND2X2 AND2X2_4728 ( .A(w_mem_inst__abc_21378_n3152_bF_buf62), .B(w_mem_inst_w_mem_6__0_), .Y(w_mem_inst__abc_21378_n5077) );
  AND2X2 AND2X2_4729 ( .A(round_ctr_rst_bF_buf59), .B(\block[320] ), .Y(w_mem_inst__abc_21378_n5078) );
  AND2X2 AND2X2_473 ( .A(_abc_15724_n1658_1), .B(_abc_15724_n1662_1), .Y(_abc_15724_n1663) );
  AND2X2 AND2X2_4730 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf62), .B(w_mem_inst__abc_21378_n5078), .Y(w_mem_inst__abc_21378_n5079) );
  AND2X2 AND2X2_4731 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf15), .B(w_mem_inst_w_mem_5__1_), .Y(w_mem_inst__abc_21378_n5082) );
  AND2X2 AND2X2_4732 ( .A(w_mem_inst__abc_21378_n3152_bF_buf61), .B(w_mem_inst_w_mem_6__1_), .Y(w_mem_inst__abc_21378_n5083) );
  AND2X2 AND2X2_4733 ( .A(round_ctr_rst_bF_buf58), .B(\block[321] ), .Y(w_mem_inst__abc_21378_n5084) );
  AND2X2 AND2X2_4734 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf61), .B(w_mem_inst__abc_21378_n5084), .Y(w_mem_inst__abc_21378_n5085) );
  AND2X2 AND2X2_4735 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf14), .B(w_mem_inst_w_mem_5__2_), .Y(w_mem_inst__abc_21378_n5088) );
  AND2X2 AND2X2_4736 ( .A(w_mem_inst__abc_21378_n3152_bF_buf60), .B(w_mem_inst_w_mem_6__2_), .Y(w_mem_inst__abc_21378_n5089) );
  AND2X2 AND2X2_4737 ( .A(round_ctr_rst_bF_buf57), .B(\block[322] ), .Y(w_mem_inst__abc_21378_n5090) );
  AND2X2 AND2X2_4738 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf60), .B(w_mem_inst__abc_21378_n5090), .Y(w_mem_inst__abc_21378_n5091) );
  AND2X2 AND2X2_4739 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf13), .B(w_mem_inst_w_mem_5__3_), .Y(w_mem_inst__abc_21378_n5094) );
  AND2X2 AND2X2_474 ( .A(_abc_15724_n1664), .B(_abc_15724_n1665), .Y(_abc_15724_n1666) );
  AND2X2 AND2X2_4740 ( .A(w_mem_inst__abc_21378_n3152_bF_buf59), .B(w_mem_inst_w_mem_6__3_), .Y(w_mem_inst__abc_21378_n5095) );
  AND2X2 AND2X2_4741 ( .A(round_ctr_rst_bF_buf56), .B(\block[323] ), .Y(w_mem_inst__abc_21378_n5096) );
  AND2X2 AND2X2_4742 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf59), .B(w_mem_inst__abc_21378_n5096), .Y(w_mem_inst__abc_21378_n5097) );
  AND2X2 AND2X2_4743 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf12), .B(w_mem_inst_w_mem_5__4_), .Y(w_mem_inst__abc_21378_n5100) );
  AND2X2 AND2X2_4744 ( .A(w_mem_inst__abc_21378_n3152_bF_buf58), .B(w_mem_inst_w_mem_6__4_), .Y(w_mem_inst__abc_21378_n5101) );
  AND2X2 AND2X2_4745 ( .A(round_ctr_rst_bF_buf55), .B(\block[324] ), .Y(w_mem_inst__abc_21378_n5102) );
  AND2X2 AND2X2_4746 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf58), .B(w_mem_inst__abc_21378_n5102), .Y(w_mem_inst__abc_21378_n5103) );
  AND2X2 AND2X2_4747 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf11), .B(w_mem_inst_w_mem_5__5_), .Y(w_mem_inst__abc_21378_n5106) );
  AND2X2 AND2X2_4748 ( .A(w_mem_inst__abc_21378_n3152_bF_buf57), .B(w_mem_inst_w_mem_6__5_), .Y(w_mem_inst__abc_21378_n5107) );
  AND2X2 AND2X2_4749 ( .A(round_ctr_rst_bF_buf54), .B(\block[325] ), .Y(w_mem_inst__abc_21378_n5108) );
  AND2X2 AND2X2_475 ( .A(_abc_15724_n1667), .B(digest_update_bF_buf5), .Y(_abc_15724_n1668_1) );
  AND2X2 AND2X2_4750 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf57), .B(w_mem_inst__abc_21378_n5108), .Y(w_mem_inst__abc_21378_n5109) );
  AND2X2 AND2X2_4751 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf10), .B(w_mem_inst_w_mem_5__6_), .Y(w_mem_inst__abc_21378_n5112) );
  AND2X2 AND2X2_4752 ( .A(w_mem_inst__abc_21378_n3152_bF_buf56), .B(w_mem_inst_w_mem_6__6_), .Y(w_mem_inst__abc_21378_n5113) );
  AND2X2 AND2X2_4753 ( .A(round_ctr_rst_bF_buf53), .B(\block[326] ), .Y(w_mem_inst__abc_21378_n5114) );
  AND2X2 AND2X2_4754 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf56), .B(w_mem_inst__abc_21378_n5114), .Y(w_mem_inst__abc_21378_n5115) );
  AND2X2 AND2X2_4755 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf9), .B(w_mem_inst_w_mem_5__7_), .Y(w_mem_inst__abc_21378_n5118) );
  AND2X2 AND2X2_4756 ( .A(w_mem_inst__abc_21378_n3152_bF_buf55), .B(w_mem_inst_w_mem_6__7_), .Y(w_mem_inst__abc_21378_n5119) );
  AND2X2 AND2X2_4757 ( .A(round_ctr_rst_bF_buf52), .B(\block[327] ), .Y(w_mem_inst__abc_21378_n5120) );
  AND2X2 AND2X2_4758 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf55), .B(w_mem_inst__abc_21378_n5120), .Y(w_mem_inst__abc_21378_n5121) );
  AND2X2 AND2X2_4759 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf8), .B(w_mem_inst_w_mem_5__8_), .Y(w_mem_inst__abc_21378_n5124) );
  AND2X2 AND2X2_476 ( .A(_abc_15724_n1669_1), .B(_abc_15724_n850_bF_buf4), .Y(_abc_15724_n1670) );
  AND2X2 AND2X2_4760 ( .A(w_mem_inst__abc_21378_n3152_bF_buf54), .B(w_mem_inst_w_mem_6__8_), .Y(w_mem_inst__abc_21378_n5125) );
  AND2X2 AND2X2_4761 ( .A(round_ctr_rst_bF_buf51), .B(\block[328] ), .Y(w_mem_inst__abc_21378_n5126) );
  AND2X2 AND2X2_4762 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf54), .B(w_mem_inst__abc_21378_n5126), .Y(w_mem_inst__abc_21378_n5127) );
  AND2X2 AND2X2_4763 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf7), .B(w_mem_inst_w_mem_5__9_), .Y(w_mem_inst__abc_21378_n5130) );
  AND2X2 AND2X2_4764 ( .A(w_mem_inst__abc_21378_n3152_bF_buf53), .B(w_mem_inst_w_mem_6__9_), .Y(w_mem_inst__abc_21378_n5131) );
  AND2X2 AND2X2_4765 ( .A(round_ctr_rst_bF_buf50), .B(\block[329] ), .Y(w_mem_inst__abc_21378_n5132) );
  AND2X2 AND2X2_4766 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf53), .B(w_mem_inst__abc_21378_n5132), .Y(w_mem_inst__abc_21378_n5133) );
  AND2X2 AND2X2_4767 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf6), .B(w_mem_inst_w_mem_5__10_), .Y(w_mem_inst__abc_21378_n5136) );
  AND2X2 AND2X2_4768 ( .A(w_mem_inst__abc_21378_n3152_bF_buf52), .B(w_mem_inst_w_mem_6__10_), .Y(w_mem_inst__abc_21378_n5137) );
  AND2X2 AND2X2_4769 ( .A(round_ctr_rst_bF_buf49), .B(\block[330] ), .Y(w_mem_inst__abc_21378_n5138) );
  AND2X2 AND2X2_477 ( .A(_abc_15724_n1619), .B(_abc_15724_n1634), .Y(_abc_15724_n1672) );
  AND2X2 AND2X2_4770 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf52), .B(w_mem_inst__abc_21378_n5138), .Y(w_mem_inst__abc_21378_n5139) );
  AND2X2 AND2X2_4771 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf5), .B(w_mem_inst_w_mem_5__11_), .Y(w_mem_inst__abc_21378_n5142) );
  AND2X2 AND2X2_4772 ( .A(w_mem_inst__abc_21378_n3152_bF_buf51), .B(w_mem_inst_w_mem_6__11_), .Y(w_mem_inst__abc_21378_n5143) );
  AND2X2 AND2X2_4773 ( .A(round_ctr_rst_bF_buf48), .B(\block[331] ), .Y(w_mem_inst__abc_21378_n5144) );
  AND2X2 AND2X2_4774 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf51), .B(w_mem_inst__abc_21378_n5144), .Y(w_mem_inst__abc_21378_n5145) );
  AND2X2 AND2X2_4775 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf4), .B(w_mem_inst_w_mem_5__12_), .Y(w_mem_inst__abc_21378_n5148) );
  AND2X2 AND2X2_4776 ( .A(w_mem_inst__abc_21378_n3152_bF_buf50), .B(w_mem_inst_w_mem_6__12_), .Y(w_mem_inst__abc_21378_n5149) );
  AND2X2 AND2X2_4777 ( .A(round_ctr_rst_bF_buf47), .B(\block[332] ), .Y(w_mem_inst__abc_21378_n5150) );
  AND2X2 AND2X2_4778 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf50), .B(w_mem_inst__abc_21378_n5150), .Y(w_mem_inst__abc_21378_n5151) );
  AND2X2 AND2X2_4779 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf3), .B(w_mem_inst_w_mem_5__13_), .Y(w_mem_inst__abc_21378_n5154) );
  AND2X2 AND2X2_478 ( .A(_abc_15724_n1649_1), .B(_abc_15724_n1662_1), .Y(_abc_15724_n1673) );
  AND2X2 AND2X2_4780 ( .A(w_mem_inst__abc_21378_n3152_bF_buf49), .B(w_mem_inst_w_mem_6__13_), .Y(w_mem_inst__abc_21378_n5155) );
  AND2X2 AND2X2_4781 ( .A(round_ctr_rst_bF_buf46), .B(\block[333] ), .Y(w_mem_inst__abc_21378_n5156) );
  AND2X2 AND2X2_4782 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf49), .B(w_mem_inst__abc_21378_n5156), .Y(w_mem_inst__abc_21378_n5157) );
  AND2X2 AND2X2_4783 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf2), .B(w_mem_inst_w_mem_5__14_), .Y(w_mem_inst__abc_21378_n5160) );
  AND2X2 AND2X2_4784 ( .A(w_mem_inst__abc_21378_n3152_bF_buf48), .B(w_mem_inst_w_mem_6__14_), .Y(w_mem_inst__abc_21378_n5161) );
  AND2X2 AND2X2_4785 ( .A(round_ctr_rst_bF_buf45), .B(\block[334] ), .Y(w_mem_inst__abc_21378_n5162) );
  AND2X2 AND2X2_4786 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf48), .B(w_mem_inst__abc_21378_n5162), .Y(w_mem_inst__abc_21378_n5163) );
  AND2X2 AND2X2_4787 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf1), .B(w_mem_inst_w_mem_5__15_), .Y(w_mem_inst__abc_21378_n5166) );
  AND2X2 AND2X2_4788 ( .A(w_mem_inst__abc_21378_n3152_bF_buf47), .B(w_mem_inst_w_mem_6__15_), .Y(w_mem_inst__abc_21378_n5167) );
  AND2X2 AND2X2_4789 ( .A(round_ctr_rst_bF_buf44), .B(\block[335] ), .Y(w_mem_inst__abc_21378_n5168) );
  AND2X2 AND2X2_479 ( .A(_abc_15724_n1672), .B(_abc_15724_n1673), .Y(_abc_15724_n1674) );
  AND2X2 AND2X2_4790 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf47), .B(w_mem_inst__abc_21378_n5168), .Y(w_mem_inst__abc_21378_n5169) );
  AND2X2 AND2X2_4791 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf0), .B(w_mem_inst_w_mem_5__16_), .Y(w_mem_inst__abc_21378_n5172) );
  AND2X2 AND2X2_4792 ( .A(w_mem_inst__abc_21378_n3152_bF_buf46), .B(w_mem_inst_w_mem_6__16_), .Y(w_mem_inst__abc_21378_n5173) );
  AND2X2 AND2X2_4793 ( .A(round_ctr_rst_bF_buf43), .B(\block[336] ), .Y(w_mem_inst__abc_21378_n5174) );
  AND2X2 AND2X2_4794 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf46), .B(w_mem_inst__abc_21378_n5174), .Y(w_mem_inst__abc_21378_n5175) );
  AND2X2 AND2X2_4795 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf60), .B(w_mem_inst_w_mem_5__17_), .Y(w_mem_inst__abc_21378_n5178) );
  AND2X2 AND2X2_4796 ( .A(w_mem_inst__abc_21378_n3152_bF_buf45), .B(w_mem_inst_w_mem_6__17_), .Y(w_mem_inst__abc_21378_n5179) );
  AND2X2 AND2X2_4797 ( .A(round_ctr_rst_bF_buf42), .B(\block[337] ), .Y(w_mem_inst__abc_21378_n5180) );
  AND2X2 AND2X2_4798 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf45), .B(w_mem_inst__abc_21378_n5180), .Y(w_mem_inst__abc_21378_n5181) );
  AND2X2 AND2X2_4799 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf59), .B(w_mem_inst_w_mem_5__18_), .Y(w_mem_inst__abc_21378_n5184) );
  AND2X2 AND2X2_48 ( .A(_auto_iopadmap_cc_313_execute_26059_4_), .B(e_reg_4_), .Y(_abc_15724_n786) );
  AND2X2 AND2X2_480 ( .A(_abc_15724_n1631_1), .B(_abc_15724_n1617_1), .Y(_abc_15724_n1677) );
  AND2X2 AND2X2_4800 ( .A(w_mem_inst__abc_21378_n3152_bF_buf44), .B(w_mem_inst_w_mem_6__18_), .Y(w_mem_inst__abc_21378_n5185) );
  AND2X2 AND2X2_4801 ( .A(round_ctr_rst_bF_buf41), .B(\block[338] ), .Y(w_mem_inst__abc_21378_n5186) );
  AND2X2 AND2X2_4802 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf44), .B(w_mem_inst__abc_21378_n5186), .Y(w_mem_inst__abc_21378_n5187) );
  AND2X2 AND2X2_4803 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf58), .B(w_mem_inst_w_mem_5__19_), .Y(w_mem_inst__abc_21378_n5190) );
  AND2X2 AND2X2_4804 ( .A(w_mem_inst__abc_21378_n3152_bF_buf43), .B(w_mem_inst_w_mem_6__19_), .Y(w_mem_inst__abc_21378_n5191) );
  AND2X2 AND2X2_4805 ( .A(round_ctr_rst_bF_buf40), .B(\block[339] ), .Y(w_mem_inst__abc_21378_n5192) );
  AND2X2 AND2X2_4806 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf43), .B(w_mem_inst__abc_21378_n5192), .Y(w_mem_inst__abc_21378_n5193) );
  AND2X2 AND2X2_4807 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf57), .B(w_mem_inst_w_mem_5__20_), .Y(w_mem_inst__abc_21378_n5196) );
  AND2X2 AND2X2_4808 ( .A(w_mem_inst__abc_21378_n3152_bF_buf42), .B(w_mem_inst_w_mem_6__20_), .Y(w_mem_inst__abc_21378_n5197) );
  AND2X2 AND2X2_4809 ( .A(round_ctr_rst_bF_buf39), .B(\block[340] ), .Y(w_mem_inst__abc_21378_n5198) );
  AND2X2 AND2X2_481 ( .A(_abc_15724_n1673), .B(_abc_15724_n1678_1), .Y(_abc_15724_n1679) );
  AND2X2 AND2X2_4810 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf42), .B(w_mem_inst__abc_21378_n5198), .Y(w_mem_inst__abc_21378_n5199) );
  AND2X2 AND2X2_4811 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf56), .B(w_mem_inst_w_mem_5__21_), .Y(w_mem_inst__abc_21378_n5202) );
  AND2X2 AND2X2_4812 ( .A(w_mem_inst__abc_21378_n3152_bF_buf41), .B(w_mem_inst_w_mem_6__21_), .Y(w_mem_inst__abc_21378_n5203) );
  AND2X2 AND2X2_4813 ( .A(round_ctr_rst_bF_buf38), .B(\block[341] ), .Y(w_mem_inst__abc_21378_n5204) );
  AND2X2 AND2X2_4814 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf41), .B(w_mem_inst__abc_21378_n5204), .Y(w_mem_inst__abc_21378_n5205) );
  AND2X2 AND2X2_4815 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf55), .B(w_mem_inst_w_mem_5__22_), .Y(w_mem_inst__abc_21378_n5208) );
  AND2X2 AND2X2_4816 ( .A(w_mem_inst__abc_21378_n3152_bF_buf40), .B(w_mem_inst_w_mem_6__22_), .Y(w_mem_inst__abc_21378_n5209) );
  AND2X2 AND2X2_4817 ( .A(round_ctr_rst_bF_buf37), .B(\block[342] ), .Y(w_mem_inst__abc_21378_n5210) );
  AND2X2 AND2X2_4818 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf40), .B(w_mem_inst__abc_21378_n5210), .Y(w_mem_inst__abc_21378_n5211) );
  AND2X2 AND2X2_4819 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf54), .B(w_mem_inst_w_mem_5__23_), .Y(w_mem_inst__abc_21378_n5214) );
  AND2X2 AND2X2_482 ( .A(_abc_15724_n1659), .B(_abc_15724_n1647), .Y(_abc_15724_n1680) );
  AND2X2 AND2X2_4820 ( .A(w_mem_inst__abc_21378_n3152_bF_buf39), .B(w_mem_inst_w_mem_6__23_), .Y(w_mem_inst__abc_21378_n5215) );
  AND2X2 AND2X2_4821 ( .A(round_ctr_rst_bF_buf36), .B(\block[343] ), .Y(w_mem_inst__abc_21378_n5216) );
  AND2X2 AND2X2_4822 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf39), .B(w_mem_inst__abc_21378_n5216), .Y(w_mem_inst__abc_21378_n5217) );
  AND2X2 AND2X2_4823 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf53), .B(w_mem_inst_w_mem_5__24_), .Y(w_mem_inst__abc_21378_n5220) );
  AND2X2 AND2X2_4824 ( .A(w_mem_inst__abc_21378_n3152_bF_buf38), .B(w_mem_inst_w_mem_6__24_), .Y(w_mem_inst__abc_21378_n5221) );
  AND2X2 AND2X2_4825 ( .A(round_ctr_rst_bF_buf35), .B(\block[344] ), .Y(w_mem_inst__abc_21378_n5222) );
  AND2X2 AND2X2_4826 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf38), .B(w_mem_inst__abc_21378_n5222), .Y(w_mem_inst__abc_21378_n5223) );
  AND2X2 AND2X2_4827 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf52), .B(w_mem_inst_w_mem_5__25_), .Y(w_mem_inst__abc_21378_n5226) );
  AND2X2 AND2X2_4828 ( .A(w_mem_inst__abc_21378_n3152_bF_buf37), .B(w_mem_inst_w_mem_6__25_), .Y(w_mem_inst__abc_21378_n5227) );
  AND2X2 AND2X2_4829 ( .A(round_ctr_rst_bF_buf34), .B(\block[345] ), .Y(w_mem_inst__abc_21378_n5228) );
  AND2X2 AND2X2_483 ( .A(_abc_15724_n1676_1), .B(_abc_15724_n1683), .Y(_abc_15724_n1684) );
  AND2X2 AND2X2_4830 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf37), .B(w_mem_inst__abc_21378_n5228), .Y(w_mem_inst__abc_21378_n5229) );
  AND2X2 AND2X2_4831 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf51), .B(w_mem_inst_w_mem_5__26_), .Y(w_mem_inst__abc_21378_n5232) );
  AND2X2 AND2X2_4832 ( .A(w_mem_inst__abc_21378_n3152_bF_buf36), .B(w_mem_inst_w_mem_6__26_), .Y(w_mem_inst__abc_21378_n5233) );
  AND2X2 AND2X2_4833 ( .A(round_ctr_rst_bF_buf33), .B(\block[346] ), .Y(w_mem_inst__abc_21378_n5234) );
  AND2X2 AND2X2_4834 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf36), .B(w_mem_inst__abc_21378_n5234), .Y(w_mem_inst__abc_21378_n5235) );
  AND2X2 AND2X2_4835 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf50), .B(w_mem_inst_w_mem_5__27_), .Y(w_mem_inst__abc_21378_n5238) );
  AND2X2 AND2X2_4836 ( .A(w_mem_inst__abc_21378_n3152_bF_buf35), .B(w_mem_inst_w_mem_6__27_), .Y(w_mem_inst__abc_21378_n5239) );
  AND2X2 AND2X2_4837 ( .A(round_ctr_rst_bF_buf32), .B(\block[347] ), .Y(w_mem_inst__abc_21378_n5240) );
  AND2X2 AND2X2_4838 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf35), .B(w_mem_inst__abc_21378_n5240), .Y(w_mem_inst__abc_21378_n5241) );
  AND2X2 AND2X2_4839 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf49), .B(w_mem_inst_w_mem_5__28_), .Y(w_mem_inst__abc_21378_n5244) );
  AND2X2 AND2X2_484 ( .A(_auto_iopadmap_cc_313_execute_26059_76_), .B(c_reg_12_), .Y(_abc_15724_n1687) );
  AND2X2 AND2X2_4840 ( .A(w_mem_inst__abc_21378_n3152_bF_buf34), .B(w_mem_inst_w_mem_6__28_), .Y(w_mem_inst__abc_21378_n5245) );
  AND2X2 AND2X2_4841 ( .A(round_ctr_rst_bF_buf31), .B(\block[348] ), .Y(w_mem_inst__abc_21378_n5246) );
  AND2X2 AND2X2_4842 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf34), .B(w_mem_inst__abc_21378_n5246), .Y(w_mem_inst__abc_21378_n5247) );
  AND2X2 AND2X2_4843 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf48), .B(w_mem_inst_w_mem_5__29_), .Y(w_mem_inst__abc_21378_n5250) );
  AND2X2 AND2X2_4844 ( .A(w_mem_inst__abc_21378_n3152_bF_buf33), .B(w_mem_inst_w_mem_6__29_), .Y(w_mem_inst__abc_21378_n5251) );
  AND2X2 AND2X2_4845 ( .A(round_ctr_rst_bF_buf30), .B(\block[349] ), .Y(w_mem_inst__abc_21378_n5252) );
  AND2X2 AND2X2_4846 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf33), .B(w_mem_inst__abc_21378_n5252), .Y(w_mem_inst__abc_21378_n5253) );
  AND2X2 AND2X2_4847 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf47), .B(w_mem_inst_w_mem_5__30_), .Y(w_mem_inst__abc_21378_n5256) );
  AND2X2 AND2X2_4848 ( .A(w_mem_inst__abc_21378_n3152_bF_buf32), .B(w_mem_inst_w_mem_6__30_), .Y(w_mem_inst__abc_21378_n5257) );
  AND2X2 AND2X2_4849 ( .A(round_ctr_rst_bF_buf29), .B(\block[350] ), .Y(w_mem_inst__abc_21378_n5258) );
  AND2X2 AND2X2_485 ( .A(_abc_15724_n1688_1), .B(_abc_15724_n1686), .Y(_abc_15724_n1689) );
  AND2X2 AND2X2_4850 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf32), .B(w_mem_inst__abc_21378_n5258), .Y(w_mem_inst__abc_21378_n5259) );
  AND2X2 AND2X2_4851 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf46), .B(w_mem_inst_w_mem_5__31_), .Y(w_mem_inst__abc_21378_n5262) );
  AND2X2 AND2X2_4852 ( .A(w_mem_inst__abc_21378_n3152_bF_buf31), .B(w_mem_inst_w_mem_6__31_), .Y(w_mem_inst__abc_21378_n5263) );
  AND2X2 AND2X2_4853 ( .A(round_ctr_rst_bF_buf28), .B(\block[351] ), .Y(w_mem_inst__abc_21378_n5264) );
  AND2X2 AND2X2_4854 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf31), .B(w_mem_inst__abc_21378_n5264), .Y(w_mem_inst__abc_21378_n5265) );
  AND2X2 AND2X2_4855 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf45), .B(w_mem_inst_w_mem_4__0_), .Y(w_mem_inst__abc_21378_n5268) );
  AND2X2 AND2X2_4856 ( .A(w_mem_inst__abc_21378_n3152_bF_buf30), .B(w_mem_inst_w_mem_5__0_), .Y(w_mem_inst__abc_21378_n5269) );
  AND2X2 AND2X2_4857 ( .A(round_ctr_rst_bF_buf27), .B(\block[352] ), .Y(w_mem_inst__abc_21378_n5270) );
  AND2X2 AND2X2_4858 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf30), .B(w_mem_inst__abc_21378_n5270), .Y(w_mem_inst__abc_21378_n5271) );
  AND2X2 AND2X2_4859 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf44), .B(w_mem_inst_w_mem_4__1_), .Y(w_mem_inst__abc_21378_n5274) );
  AND2X2 AND2X2_486 ( .A(_abc_15724_n1685), .B(_abc_15724_n1689), .Y(_abc_15724_n1691) );
  AND2X2 AND2X2_4860 ( .A(w_mem_inst__abc_21378_n3152_bF_buf29), .B(w_mem_inst_w_mem_5__1_), .Y(w_mem_inst__abc_21378_n5275) );
  AND2X2 AND2X2_4861 ( .A(round_ctr_rst_bF_buf26), .B(\block[353] ), .Y(w_mem_inst__abc_21378_n5276) );
  AND2X2 AND2X2_4862 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf29), .B(w_mem_inst__abc_21378_n5276), .Y(w_mem_inst__abc_21378_n5277) );
  AND2X2 AND2X2_4863 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf43), .B(w_mem_inst_w_mem_4__2_), .Y(w_mem_inst__abc_21378_n5280) );
  AND2X2 AND2X2_4864 ( .A(w_mem_inst__abc_21378_n3152_bF_buf28), .B(w_mem_inst_w_mem_5__2_), .Y(w_mem_inst__abc_21378_n5281) );
  AND2X2 AND2X2_4865 ( .A(round_ctr_rst_bF_buf25), .B(\block[354] ), .Y(w_mem_inst__abc_21378_n5282) );
  AND2X2 AND2X2_4866 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf28), .B(w_mem_inst__abc_21378_n5282), .Y(w_mem_inst__abc_21378_n5283) );
  AND2X2 AND2X2_4867 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf42), .B(w_mem_inst_w_mem_4__3_), .Y(w_mem_inst__abc_21378_n5286) );
  AND2X2 AND2X2_4868 ( .A(w_mem_inst__abc_21378_n3152_bF_buf27), .B(w_mem_inst_w_mem_5__3_), .Y(w_mem_inst__abc_21378_n5287) );
  AND2X2 AND2X2_4869 ( .A(round_ctr_rst_bF_buf24), .B(\block[355] ), .Y(w_mem_inst__abc_21378_n5288) );
  AND2X2 AND2X2_487 ( .A(_abc_15724_n1692_1), .B(_abc_15724_n1690), .Y(_abc_15724_n1693) );
  AND2X2 AND2X2_4870 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf27), .B(w_mem_inst__abc_21378_n5288), .Y(w_mem_inst__abc_21378_n5289) );
  AND2X2 AND2X2_4871 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf41), .B(w_mem_inst_w_mem_4__4_), .Y(w_mem_inst__abc_21378_n5292) );
  AND2X2 AND2X2_4872 ( .A(w_mem_inst__abc_21378_n3152_bF_buf26), .B(w_mem_inst_w_mem_5__4_), .Y(w_mem_inst__abc_21378_n5293) );
  AND2X2 AND2X2_4873 ( .A(round_ctr_rst_bF_buf23), .B(\block[356] ), .Y(w_mem_inst__abc_21378_n5294) );
  AND2X2 AND2X2_4874 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf26), .B(w_mem_inst__abc_21378_n5294), .Y(w_mem_inst__abc_21378_n5295) );
  AND2X2 AND2X2_4875 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf40), .B(w_mem_inst_w_mem_4__5_), .Y(w_mem_inst__abc_21378_n5298) );
  AND2X2 AND2X2_4876 ( .A(w_mem_inst__abc_21378_n3152_bF_buf25), .B(w_mem_inst_w_mem_5__5_), .Y(w_mem_inst__abc_21378_n5299) );
  AND2X2 AND2X2_4877 ( .A(round_ctr_rst_bF_buf22), .B(\block[357] ), .Y(w_mem_inst__abc_21378_n5300) );
  AND2X2 AND2X2_4878 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf25), .B(w_mem_inst__abc_21378_n5300), .Y(w_mem_inst__abc_21378_n5301) );
  AND2X2 AND2X2_4879 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf39), .B(w_mem_inst_w_mem_4__6_), .Y(w_mem_inst__abc_21378_n5304) );
  AND2X2 AND2X2_488 ( .A(_abc_15724_n1693), .B(digest_update_bF_buf4), .Y(_abc_15724_n1694) );
  AND2X2 AND2X2_4880 ( .A(w_mem_inst__abc_21378_n3152_bF_buf24), .B(w_mem_inst_w_mem_5__6_), .Y(w_mem_inst__abc_21378_n5305) );
  AND2X2 AND2X2_4881 ( .A(round_ctr_rst_bF_buf21), .B(\block[358] ), .Y(w_mem_inst__abc_21378_n5306) );
  AND2X2 AND2X2_4882 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf24), .B(w_mem_inst__abc_21378_n5306), .Y(w_mem_inst__abc_21378_n5307) );
  AND2X2 AND2X2_4883 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf38), .B(w_mem_inst_w_mem_4__7_), .Y(w_mem_inst__abc_21378_n5310) );
  AND2X2 AND2X2_4884 ( .A(w_mem_inst__abc_21378_n3152_bF_buf23), .B(w_mem_inst_w_mem_5__7_), .Y(w_mem_inst__abc_21378_n5311) );
  AND2X2 AND2X2_4885 ( .A(round_ctr_rst_bF_buf20), .B(\block[359] ), .Y(w_mem_inst__abc_21378_n5312) );
  AND2X2 AND2X2_4886 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf23), .B(w_mem_inst__abc_21378_n5312), .Y(w_mem_inst__abc_21378_n5313) );
  AND2X2 AND2X2_4887 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf37), .B(w_mem_inst_w_mem_4__8_), .Y(w_mem_inst__abc_21378_n5316) );
  AND2X2 AND2X2_4888 ( .A(w_mem_inst__abc_21378_n3152_bF_buf22), .B(w_mem_inst_w_mem_5__8_), .Y(w_mem_inst__abc_21378_n5317) );
  AND2X2 AND2X2_4889 ( .A(round_ctr_rst_bF_buf19), .B(\block[360] ), .Y(w_mem_inst__abc_21378_n5318) );
  AND2X2 AND2X2_489 ( .A(_abc_15724_n1695), .B(_abc_15724_n850_bF_buf3), .Y(_abc_15724_n1696_1) );
  AND2X2 AND2X2_4890 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf22), .B(w_mem_inst__abc_21378_n5318), .Y(w_mem_inst__abc_21378_n5319) );
  AND2X2 AND2X2_4891 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf36), .B(w_mem_inst_w_mem_4__9_), .Y(w_mem_inst__abc_21378_n5322) );
  AND2X2 AND2X2_4892 ( .A(w_mem_inst__abc_21378_n3152_bF_buf21), .B(w_mem_inst_w_mem_5__9_), .Y(w_mem_inst__abc_21378_n5323) );
  AND2X2 AND2X2_4893 ( .A(round_ctr_rst_bF_buf18), .B(\block[361] ), .Y(w_mem_inst__abc_21378_n5324) );
  AND2X2 AND2X2_4894 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf21), .B(w_mem_inst__abc_21378_n5324), .Y(w_mem_inst__abc_21378_n5325) );
  AND2X2 AND2X2_4895 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf35), .B(w_mem_inst_w_mem_4__10_), .Y(w_mem_inst__abc_21378_n5328) );
  AND2X2 AND2X2_4896 ( .A(w_mem_inst__abc_21378_n3152_bF_buf20), .B(w_mem_inst_w_mem_5__10_), .Y(w_mem_inst__abc_21378_n5329) );
  AND2X2 AND2X2_4897 ( .A(round_ctr_rst_bF_buf17), .B(\block[362] ), .Y(w_mem_inst__abc_21378_n5330) );
  AND2X2 AND2X2_4898 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf20), .B(w_mem_inst__abc_21378_n5330), .Y(w_mem_inst__abc_21378_n5331) );
  AND2X2 AND2X2_4899 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf34), .B(w_mem_inst_w_mem_4__11_), .Y(w_mem_inst__abc_21378_n5334) );
  AND2X2 AND2X2_49 ( .A(e_reg_3_), .B(_auto_iopadmap_cc_313_execute_26059_3_), .Y(_abc_15724_n787) );
  AND2X2 AND2X2_490 ( .A(_auto_iopadmap_cc_313_execute_26059_77_), .B(c_reg_13_), .Y(_abc_15724_n1699) );
  AND2X2 AND2X2_4900 ( .A(w_mem_inst__abc_21378_n3152_bF_buf19), .B(w_mem_inst_w_mem_5__11_), .Y(w_mem_inst__abc_21378_n5335) );
  AND2X2 AND2X2_4901 ( .A(round_ctr_rst_bF_buf16), .B(\block[363] ), .Y(w_mem_inst__abc_21378_n5336) );
  AND2X2 AND2X2_4902 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf19), .B(w_mem_inst__abc_21378_n5336), .Y(w_mem_inst__abc_21378_n5337) );
  AND2X2 AND2X2_4903 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf33), .B(w_mem_inst_w_mem_4__12_), .Y(w_mem_inst__abc_21378_n5340) );
  AND2X2 AND2X2_4904 ( .A(w_mem_inst__abc_21378_n3152_bF_buf18), .B(w_mem_inst_w_mem_5__12_), .Y(w_mem_inst__abc_21378_n5341) );
  AND2X2 AND2X2_4905 ( .A(round_ctr_rst_bF_buf15), .B(\block[364] ), .Y(w_mem_inst__abc_21378_n5342) );
  AND2X2 AND2X2_4906 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf18), .B(w_mem_inst__abc_21378_n5342), .Y(w_mem_inst__abc_21378_n5343) );
  AND2X2 AND2X2_4907 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf32), .B(w_mem_inst_w_mem_4__13_), .Y(w_mem_inst__abc_21378_n5346) );
  AND2X2 AND2X2_4908 ( .A(w_mem_inst__abc_21378_n3152_bF_buf17), .B(w_mem_inst_w_mem_5__13_), .Y(w_mem_inst__abc_21378_n5347) );
  AND2X2 AND2X2_4909 ( .A(round_ctr_rst_bF_buf14), .B(\block[365] ), .Y(w_mem_inst__abc_21378_n5348) );
  AND2X2 AND2X2_491 ( .A(_abc_15724_n1700_1), .B(_abc_15724_n1698), .Y(_abc_15724_n1701) );
  AND2X2 AND2X2_4910 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf17), .B(w_mem_inst__abc_21378_n5348), .Y(w_mem_inst__abc_21378_n5349) );
  AND2X2 AND2X2_4911 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf31), .B(w_mem_inst_w_mem_4__14_), .Y(w_mem_inst__abc_21378_n5352) );
  AND2X2 AND2X2_4912 ( .A(w_mem_inst__abc_21378_n3152_bF_buf16), .B(w_mem_inst_w_mem_5__14_), .Y(w_mem_inst__abc_21378_n5353) );
  AND2X2 AND2X2_4913 ( .A(round_ctr_rst_bF_buf13), .B(\block[366] ), .Y(w_mem_inst__abc_21378_n5354) );
  AND2X2 AND2X2_4914 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf16), .B(w_mem_inst__abc_21378_n5354), .Y(w_mem_inst__abc_21378_n5355) );
  AND2X2 AND2X2_4915 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf30), .B(w_mem_inst_w_mem_4__15_), .Y(w_mem_inst__abc_21378_n5358) );
  AND2X2 AND2X2_4916 ( .A(w_mem_inst__abc_21378_n3152_bF_buf15), .B(w_mem_inst_w_mem_5__15_), .Y(w_mem_inst__abc_21378_n5359) );
  AND2X2 AND2X2_4917 ( .A(round_ctr_rst_bF_buf12), .B(\block[367] ), .Y(w_mem_inst__abc_21378_n5360) );
  AND2X2 AND2X2_4918 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf15), .B(w_mem_inst__abc_21378_n5360), .Y(w_mem_inst__abc_21378_n5361) );
  AND2X2 AND2X2_4919 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf29), .B(w_mem_inst_w_mem_4__16_), .Y(w_mem_inst__abc_21378_n5364) );
  AND2X2 AND2X2_492 ( .A(_abc_15724_n1692_1), .B(_abc_15724_n1688_1), .Y(_abc_15724_n1702) );
  AND2X2 AND2X2_4920 ( .A(w_mem_inst__abc_21378_n3152_bF_buf14), .B(w_mem_inst_w_mem_5__16_), .Y(w_mem_inst__abc_21378_n5365) );
  AND2X2 AND2X2_4921 ( .A(round_ctr_rst_bF_buf11), .B(\block[368] ), .Y(w_mem_inst__abc_21378_n5366) );
  AND2X2 AND2X2_4922 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf14), .B(w_mem_inst__abc_21378_n5366), .Y(w_mem_inst__abc_21378_n5367) );
  AND2X2 AND2X2_4923 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf28), .B(w_mem_inst_w_mem_4__17_), .Y(w_mem_inst__abc_21378_n5370) );
  AND2X2 AND2X2_4924 ( .A(w_mem_inst__abc_21378_n3152_bF_buf13), .B(w_mem_inst_w_mem_5__17_), .Y(w_mem_inst__abc_21378_n5371) );
  AND2X2 AND2X2_4925 ( .A(round_ctr_rst_bF_buf10), .B(\block[369] ), .Y(w_mem_inst__abc_21378_n5372) );
  AND2X2 AND2X2_4926 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf13), .B(w_mem_inst__abc_21378_n5372), .Y(w_mem_inst__abc_21378_n5373) );
  AND2X2 AND2X2_4927 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf27), .B(w_mem_inst_w_mem_4__18_), .Y(w_mem_inst__abc_21378_n5376) );
  AND2X2 AND2X2_4928 ( .A(w_mem_inst__abc_21378_n3152_bF_buf12), .B(w_mem_inst_w_mem_5__18_), .Y(w_mem_inst__abc_21378_n5377) );
  AND2X2 AND2X2_4929 ( .A(round_ctr_rst_bF_buf9), .B(\block[370] ), .Y(w_mem_inst__abc_21378_n5378) );
  AND2X2 AND2X2_493 ( .A(_abc_15724_n1703), .B(_abc_15724_n1701), .Y(_abc_15724_n1705) );
  AND2X2 AND2X2_4930 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf12), .B(w_mem_inst__abc_21378_n5378), .Y(w_mem_inst__abc_21378_n5379) );
  AND2X2 AND2X2_4931 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf26), .B(w_mem_inst_w_mem_4__19_), .Y(w_mem_inst__abc_21378_n5382) );
  AND2X2 AND2X2_4932 ( .A(w_mem_inst__abc_21378_n3152_bF_buf11), .B(w_mem_inst_w_mem_5__19_), .Y(w_mem_inst__abc_21378_n5383) );
  AND2X2 AND2X2_4933 ( .A(round_ctr_rst_bF_buf8), .B(\block[371] ), .Y(w_mem_inst__abc_21378_n5384) );
  AND2X2 AND2X2_4934 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf11), .B(w_mem_inst__abc_21378_n5384), .Y(w_mem_inst__abc_21378_n5385) );
  AND2X2 AND2X2_4935 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf25), .B(w_mem_inst_w_mem_4__20_), .Y(w_mem_inst__abc_21378_n5388) );
  AND2X2 AND2X2_4936 ( .A(w_mem_inst__abc_21378_n3152_bF_buf10), .B(w_mem_inst_w_mem_5__20_), .Y(w_mem_inst__abc_21378_n5389) );
  AND2X2 AND2X2_4937 ( .A(round_ctr_rst_bF_buf7), .B(\block[372] ), .Y(w_mem_inst__abc_21378_n5390) );
  AND2X2 AND2X2_4938 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf10), .B(w_mem_inst__abc_21378_n5390), .Y(w_mem_inst__abc_21378_n5391) );
  AND2X2 AND2X2_4939 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf24), .B(w_mem_inst_w_mem_4__21_), .Y(w_mem_inst__abc_21378_n5394) );
  AND2X2 AND2X2_494 ( .A(_abc_15724_n1706), .B(_abc_15724_n1704_1), .Y(_abc_15724_n1707) );
  AND2X2 AND2X2_4940 ( .A(w_mem_inst__abc_21378_n3152_bF_buf9), .B(w_mem_inst_w_mem_5__21_), .Y(w_mem_inst__abc_21378_n5395) );
  AND2X2 AND2X2_4941 ( .A(round_ctr_rst_bF_buf6), .B(\block[373] ), .Y(w_mem_inst__abc_21378_n5396) );
  AND2X2 AND2X2_4942 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf9), .B(w_mem_inst__abc_21378_n5396), .Y(w_mem_inst__abc_21378_n5397) );
  AND2X2 AND2X2_4943 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf23), .B(w_mem_inst_w_mem_4__22_), .Y(w_mem_inst__abc_21378_n5400) );
  AND2X2 AND2X2_4944 ( .A(w_mem_inst__abc_21378_n3152_bF_buf8), .B(w_mem_inst_w_mem_5__22_), .Y(w_mem_inst__abc_21378_n5401) );
  AND2X2 AND2X2_4945 ( .A(round_ctr_rst_bF_buf5), .B(\block[374] ), .Y(w_mem_inst__abc_21378_n5402) );
  AND2X2 AND2X2_4946 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf8), .B(w_mem_inst__abc_21378_n5402), .Y(w_mem_inst__abc_21378_n5403) );
  AND2X2 AND2X2_4947 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf22), .B(w_mem_inst_w_mem_4__23_), .Y(w_mem_inst__abc_21378_n5406) );
  AND2X2 AND2X2_4948 ( .A(w_mem_inst__abc_21378_n3152_bF_buf7), .B(w_mem_inst_w_mem_5__23_), .Y(w_mem_inst__abc_21378_n5407) );
  AND2X2 AND2X2_4949 ( .A(round_ctr_rst_bF_buf4), .B(\block[375] ), .Y(w_mem_inst__abc_21378_n5408) );
  AND2X2 AND2X2_495 ( .A(_abc_15724_n1707), .B(digest_update_bF_buf3), .Y(_abc_15724_n1708) );
  AND2X2 AND2X2_4950 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf7), .B(w_mem_inst__abc_21378_n5408), .Y(w_mem_inst__abc_21378_n5409) );
  AND2X2 AND2X2_4951 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf21), .B(w_mem_inst_w_mem_4__24_), .Y(w_mem_inst__abc_21378_n5412) );
  AND2X2 AND2X2_4952 ( .A(w_mem_inst__abc_21378_n3152_bF_buf6), .B(w_mem_inst_w_mem_5__24_), .Y(w_mem_inst__abc_21378_n5413) );
  AND2X2 AND2X2_4953 ( .A(round_ctr_rst_bF_buf3), .B(\block[376] ), .Y(w_mem_inst__abc_21378_n5414) );
  AND2X2 AND2X2_4954 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf6), .B(w_mem_inst__abc_21378_n5414), .Y(w_mem_inst__abc_21378_n5415) );
  AND2X2 AND2X2_4955 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf20), .B(w_mem_inst_w_mem_4__25_), .Y(w_mem_inst__abc_21378_n5418) );
  AND2X2 AND2X2_4956 ( .A(w_mem_inst__abc_21378_n3152_bF_buf5), .B(w_mem_inst_w_mem_5__25_), .Y(w_mem_inst__abc_21378_n5419) );
  AND2X2 AND2X2_4957 ( .A(round_ctr_rst_bF_buf2), .B(\block[377] ), .Y(w_mem_inst__abc_21378_n5420) );
  AND2X2 AND2X2_4958 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf5), .B(w_mem_inst__abc_21378_n5420), .Y(w_mem_inst__abc_21378_n5421) );
  AND2X2 AND2X2_4959 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf19), .B(w_mem_inst_w_mem_4__26_), .Y(w_mem_inst__abc_21378_n5424) );
  AND2X2 AND2X2_496 ( .A(_abc_15724_n907_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_77_), .Y(_abc_15724_n1709_1) );
  AND2X2 AND2X2_4960 ( .A(w_mem_inst__abc_21378_n3152_bF_buf4), .B(w_mem_inst_w_mem_5__26_), .Y(w_mem_inst__abc_21378_n5425) );
  AND2X2 AND2X2_4961 ( .A(round_ctr_rst_bF_buf1), .B(\block[378] ), .Y(w_mem_inst__abc_21378_n5426) );
  AND2X2 AND2X2_4962 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf4), .B(w_mem_inst__abc_21378_n5426), .Y(w_mem_inst__abc_21378_n5427) );
  AND2X2 AND2X2_4963 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf18), .B(w_mem_inst_w_mem_4__27_), .Y(w_mem_inst__abc_21378_n5430) );
  AND2X2 AND2X2_4964 ( .A(w_mem_inst__abc_21378_n3152_bF_buf3), .B(w_mem_inst_w_mem_5__27_), .Y(w_mem_inst__abc_21378_n5431) );
  AND2X2 AND2X2_4965 ( .A(round_ctr_rst_bF_buf0), .B(\block[379] ), .Y(w_mem_inst__abc_21378_n5432) );
  AND2X2 AND2X2_4966 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf3), .B(w_mem_inst__abc_21378_n5432), .Y(w_mem_inst__abc_21378_n5433) );
  AND2X2 AND2X2_4967 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf17), .B(w_mem_inst_w_mem_4__28_), .Y(w_mem_inst__abc_21378_n5436) );
  AND2X2 AND2X2_4968 ( .A(w_mem_inst__abc_21378_n3152_bF_buf2), .B(w_mem_inst_w_mem_5__28_), .Y(w_mem_inst__abc_21378_n5437) );
  AND2X2 AND2X2_4969 ( .A(round_ctr_rst_bF_buf63), .B(\block[380] ), .Y(w_mem_inst__abc_21378_n5438) );
  AND2X2 AND2X2_497 ( .A(_abc_15724_n1706), .B(_abc_15724_n1700_1), .Y(_abc_15724_n1711) );
  AND2X2 AND2X2_4970 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf2), .B(w_mem_inst__abc_21378_n5438), .Y(w_mem_inst__abc_21378_n5439) );
  AND2X2 AND2X2_4971 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf16), .B(w_mem_inst_w_mem_4__29_), .Y(w_mem_inst__abc_21378_n5442) );
  AND2X2 AND2X2_4972 ( .A(w_mem_inst__abc_21378_n3152_bF_buf1), .B(w_mem_inst_w_mem_5__29_), .Y(w_mem_inst__abc_21378_n5443) );
  AND2X2 AND2X2_4973 ( .A(round_ctr_rst_bF_buf62), .B(\block[381] ), .Y(w_mem_inst__abc_21378_n5444) );
  AND2X2 AND2X2_4974 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf1), .B(w_mem_inst__abc_21378_n5444), .Y(w_mem_inst__abc_21378_n5445) );
  AND2X2 AND2X2_4975 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf15), .B(w_mem_inst_w_mem_4__30_), .Y(w_mem_inst__abc_21378_n5448) );
  AND2X2 AND2X2_4976 ( .A(w_mem_inst__abc_21378_n3152_bF_buf0), .B(w_mem_inst_w_mem_5__30_), .Y(w_mem_inst__abc_21378_n5449) );
  AND2X2 AND2X2_4977 ( .A(round_ctr_rst_bF_buf61), .B(\block[382] ), .Y(w_mem_inst__abc_21378_n5450) );
  AND2X2 AND2X2_4978 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf0), .B(w_mem_inst__abc_21378_n5450), .Y(w_mem_inst__abc_21378_n5451) );
  AND2X2 AND2X2_4979 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf14), .B(w_mem_inst_w_mem_4__31_), .Y(w_mem_inst__abc_21378_n5454) );
  AND2X2 AND2X2_498 ( .A(_auto_iopadmap_cc_313_execute_26059_78_), .B(c_reg_14_), .Y(_abc_15724_n1714_1) );
  AND2X2 AND2X2_4980 ( .A(w_mem_inst__abc_21378_n3152_bF_buf63), .B(w_mem_inst_w_mem_5__31_), .Y(w_mem_inst__abc_21378_n5455) );
  AND2X2 AND2X2_4981 ( .A(round_ctr_rst_bF_buf60), .B(\block[383] ), .Y(w_mem_inst__abc_21378_n5456) );
  AND2X2 AND2X2_4982 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf63), .B(w_mem_inst__abc_21378_n5456), .Y(w_mem_inst__abc_21378_n5457) );
  AND2X2 AND2X2_4983 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf13), .B(w_mem_inst_w_mem_3__0_), .Y(w_mem_inst__abc_21378_n5460) );
  AND2X2 AND2X2_4984 ( .A(w_mem_inst__abc_21378_n3152_bF_buf62), .B(w_mem_inst_w_mem_4__0_), .Y(w_mem_inst__abc_21378_n5461) );
  AND2X2 AND2X2_4985 ( .A(round_ctr_rst_bF_buf59), .B(\block[384] ), .Y(w_mem_inst__abc_21378_n5462) );
  AND2X2 AND2X2_4986 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf62), .B(w_mem_inst__abc_21378_n5462), .Y(w_mem_inst__abc_21378_n5463) );
  AND2X2 AND2X2_4987 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf12), .B(w_mem_inst_w_mem_3__1_), .Y(w_mem_inst__abc_21378_n5466) );
  AND2X2 AND2X2_4988 ( .A(w_mem_inst__abc_21378_n3152_bF_buf61), .B(w_mem_inst_w_mem_4__1_), .Y(w_mem_inst__abc_21378_n5467) );
  AND2X2 AND2X2_4989 ( .A(round_ctr_rst_bF_buf58), .B(\block[385] ), .Y(w_mem_inst__abc_21378_n5468) );
  AND2X2 AND2X2_499 ( .A(_abc_15724_n1715), .B(_abc_15724_n1713), .Y(_abc_15724_n1716) );
  AND2X2 AND2X2_4990 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf61), .B(w_mem_inst__abc_21378_n5468), .Y(w_mem_inst__abc_21378_n5469) );
  AND2X2 AND2X2_4991 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf11), .B(w_mem_inst_w_mem_3__2_), .Y(w_mem_inst__abc_21378_n5472) );
  AND2X2 AND2X2_4992 ( .A(w_mem_inst__abc_21378_n3152_bF_buf60), .B(w_mem_inst_w_mem_4__2_), .Y(w_mem_inst__abc_21378_n5473) );
  AND2X2 AND2X2_4993 ( .A(round_ctr_rst_bF_buf57), .B(\block[386] ), .Y(w_mem_inst__abc_21378_n5474) );
  AND2X2 AND2X2_4994 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf60), .B(w_mem_inst__abc_21378_n5474), .Y(w_mem_inst__abc_21378_n5475) );
  AND2X2 AND2X2_4995 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf10), .B(w_mem_inst_w_mem_3__3_), .Y(w_mem_inst__abc_21378_n5478) );
  AND2X2 AND2X2_4996 ( .A(w_mem_inst__abc_21378_n3152_bF_buf59), .B(w_mem_inst_w_mem_4__3_), .Y(w_mem_inst__abc_21378_n5479) );
  AND2X2 AND2X2_4997 ( .A(round_ctr_rst_bF_buf56), .B(\block[387] ), .Y(w_mem_inst__abc_21378_n5480) );
  AND2X2 AND2X2_4998 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf59), .B(w_mem_inst__abc_21378_n5480), .Y(w_mem_inst__abc_21378_n5481) );
  AND2X2 AND2X2_4999 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf9), .B(w_mem_inst_w_mem_3__4_), .Y(w_mem_inst__abc_21378_n5484) );
  AND2X2 AND2X2_5 ( .A(e_reg_19_), .B(_auto_iopadmap_cc_313_execute_26059_19_), .Y(_abc_15724_n705) );
  AND2X2 AND2X2_50 ( .A(e_reg_2_), .B(_auto_iopadmap_cc_313_execute_26059_2_), .Y(_abc_15724_n789_1) );
  AND2X2 AND2X2_500 ( .A(_abc_15724_n1712), .B(_abc_15724_n1716), .Y(_abc_15724_n1718) );
  AND2X2 AND2X2_5000 ( .A(w_mem_inst__abc_21378_n3152_bF_buf58), .B(w_mem_inst_w_mem_4__4_), .Y(w_mem_inst__abc_21378_n5485) );
  AND2X2 AND2X2_5001 ( .A(round_ctr_rst_bF_buf55), .B(\block[388] ), .Y(w_mem_inst__abc_21378_n5486) );
  AND2X2 AND2X2_5002 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf58), .B(w_mem_inst__abc_21378_n5486), .Y(w_mem_inst__abc_21378_n5487) );
  AND2X2 AND2X2_5003 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf8), .B(w_mem_inst_w_mem_3__5_), .Y(w_mem_inst__abc_21378_n5490) );
  AND2X2 AND2X2_5004 ( .A(w_mem_inst__abc_21378_n3152_bF_buf57), .B(w_mem_inst_w_mem_4__5_), .Y(w_mem_inst__abc_21378_n5491) );
  AND2X2 AND2X2_5005 ( .A(round_ctr_rst_bF_buf54), .B(\block[389] ), .Y(w_mem_inst__abc_21378_n5492) );
  AND2X2 AND2X2_5006 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf57), .B(w_mem_inst__abc_21378_n5492), .Y(w_mem_inst__abc_21378_n5493) );
  AND2X2 AND2X2_5007 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf7), .B(w_mem_inst_w_mem_3__6_), .Y(w_mem_inst__abc_21378_n5496) );
  AND2X2 AND2X2_5008 ( .A(w_mem_inst__abc_21378_n3152_bF_buf56), .B(w_mem_inst_w_mem_4__6_), .Y(w_mem_inst__abc_21378_n5497) );
  AND2X2 AND2X2_5009 ( .A(round_ctr_rst_bF_buf53), .B(\block[390] ), .Y(w_mem_inst__abc_21378_n5498) );
  AND2X2 AND2X2_501 ( .A(_abc_15724_n1719_1), .B(_abc_15724_n1717), .Y(_abc_15724_n1720) );
  AND2X2 AND2X2_5010 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf56), .B(w_mem_inst__abc_21378_n5498), .Y(w_mem_inst__abc_21378_n5499) );
  AND2X2 AND2X2_5011 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf6), .B(w_mem_inst_w_mem_3__7_), .Y(w_mem_inst__abc_21378_n5502) );
  AND2X2 AND2X2_5012 ( .A(w_mem_inst__abc_21378_n3152_bF_buf55), .B(w_mem_inst_w_mem_4__7_), .Y(w_mem_inst__abc_21378_n5503) );
  AND2X2 AND2X2_5013 ( .A(round_ctr_rst_bF_buf52), .B(\block[391] ), .Y(w_mem_inst__abc_21378_n5504) );
  AND2X2 AND2X2_5014 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf55), .B(w_mem_inst__abc_21378_n5504), .Y(w_mem_inst__abc_21378_n5505) );
  AND2X2 AND2X2_5015 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf5), .B(w_mem_inst_w_mem_3__8_), .Y(w_mem_inst__abc_21378_n5508) );
  AND2X2 AND2X2_5016 ( .A(w_mem_inst__abc_21378_n3152_bF_buf54), .B(w_mem_inst_w_mem_4__8_), .Y(w_mem_inst__abc_21378_n5509) );
  AND2X2 AND2X2_5017 ( .A(round_ctr_rst_bF_buf51), .B(\block[392] ), .Y(w_mem_inst__abc_21378_n5510) );
  AND2X2 AND2X2_5018 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf54), .B(w_mem_inst__abc_21378_n5510), .Y(w_mem_inst__abc_21378_n5511) );
  AND2X2 AND2X2_5019 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf4), .B(w_mem_inst_w_mem_3__9_), .Y(w_mem_inst__abc_21378_n5514) );
  AND2X2 AND2X2_502 ( .A(_abc_15724_n1720), .B(digest_update_bF_buf2), .Y(_abc_15724_n1721) );
  AND2X2 AND2X2_5020 ( .A(w_mem_inst__abc_21378_n3152_bF_buf53), .B(w_mem_inst_w_mem_4__9_), .Y(w_mem_inst__abc_21378_n5515) );
  AND2X2 AND2X2_5021 ( .A(round_ctr_rst_bF_buf50), .B(\block[393] ), .Y(w_mem_inst__abc_21378_n5516) );
  AND2X2 AND2X2_5022 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf53), .B(w_mem_inst__abc_21378_n5516), .Y(w_mem_inst__abc_21378_n5517) );
  AND2X2 AND2X2_5023 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf3), .B(w_mem_inst_w_mem_3__10_), .Y(w_mem_inst__abc_21378_n5520) );
  AND2X2 AND2X2_5024 ( .A(w_mem_inst__abc_21378_n3152_bF_buf52), .B(w_mem_inst_w_mem_4__10_), .Y(w_mem_inst__abc_21378_n5521) );
  AND2X2 AND2X2_5025 ( .A(round_ctr_rst_bF_buf49), .B(\block[394] ), .Y(w_mem_inst__abc_21378_n5522) );
  AND2X2 AND2X2_5026 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf52), .B(w_mem_inst__abc_21378_n5522), .Y(w_mem_inst__abc_21378_n5523) );
  AND2X2 AND2X2_5027 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf2), .B(w_mem_inst_w_mem_3__11_), .Y(w_mem_inst__abc_21378_n5526) );
  AND2X2 AND2X2_5028 ( .A(w_mem_inst__abc_21378_n3152_bF_buf51), .B(w_mem_inst_w_mem_4__11_), .Y(w_mem_inst__abc_21378_n5527) );
  AND2X2 AND2X2_5029 ( .A(round_ctr_rst_bF_buf48), .B(\block[395] ), .Y(w_mem_inst__abc_21378_n5528) );
  AND2X2 AND2X2_503 ( .A(_abc_15724_n1722), .B(_abc_15724_n850_bF_buf2), .Y(_abc_15724_n1723) );
  AND2X2 AND2X2_5030 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf51), .B(w_mem_inst__abc_21378_n5528), .Y(w_mem_inst__abc_21378_n5529) );
  AND2X2 AND2X2_5031 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf1), .B(w_mem_inst_w_mem_3__12_), .Y(w_mem_inst__abc_21378_n5532) );
  AND2X2 AND2X2_5032 ( .A(w_mem_inst__abc_21378_n3152_bF_buf50), .B(w_mem_inst_w_mem_4__12_), .Y(w_mem_inst__abc_21378_n5533) );
  AND2X2 AND2X2_5033 ( .A(round_ctr_rst_bF_buf47), .B(\block[396] ), .Y(w_mem_inst__abc_21378_n5534) );
  AND2X2 AND2X2_5034 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf50), .B(w_mem_inst__abc_21378_n5534), .Y(w_mem_inst__abc_21378_n5535) );
  AND2X2 AND2X2_5035 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf0), .B(w_mem_inst_w_mem_3__13_), .Y(w_mem_inst__abc_21378_n5538) );
  AND2X2 AND2X2_5036 ( .A(w_mem_inst__abc_21378_n3152_bF_buf49), .B(w_mem_inst_w_mem_4__13_), .Y(w_mem_inst__abc_21378_n5539) );
  AND2X2 AND2X2_5037 ( .A(round_ctr_rst_bF_buf46), .B(\block[397] ), .Y(w_mem_inst__abc_21378_n5540) );
  AND2X2 AND2X2_5038 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf49), .B(w_mem_inst__abc_21378_n5540), .Y(w_mem_inst__abc_21378_n5541) );
  AND2X2 AND2X2_5039 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf60), .B(w_mem_inst_w_mem_3__14_), .Y(w_mem_inst__abc_21378_n5544) );
  AND2X2 AND2X2_504 ( .A(_abc_15724_n1719_1), .B(_abc_15724_n1715), .Y(_abc_15724_n1725) );
  AND2X2 AND2X2_5040 ( .A(w_mem_inst__abc_21378_n3152_bF_buf48), .B(w_mem_inst_w_mem_4__14_), .Y(w_mem_inst__abc_21378_n5545) );
  AND2X2 AND2X2_5041 ( .A(round_ctr_rst_bF_buf45), .B(\block[398] ), .Y(w_mem_inst__abc_21378_n5546) );
  AND2X2 AND2X2_5042 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf48), .B(w_mem_inst__abc_21378_n5546), .Y(w_mem_inst__abc_21378_n5547) );
  AND2X2 AND2X2_5043 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf59), .B(w_mem_inst_w_mem_3__15_), .Y(w_mem_inst__abc_21378_n5550) );
  AND2X2 AND2X2_5044 ( .A(w_mem_inst__abc_21378_n3152_bF_buf47), .B(w_mem_inst_w_mem_4__15_), .Y(w_mem_inst__abc_21378_n5551) );
  AND2X2 AND2X2_5045 ( .A(round_ctr_rst_bF_buf44), .B(\block[399] ), .Y(w_mem_inst__abc_21378_n5552) );
  AND2X2 AND2X2_5046 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf47), .B(w_mem_inst__abc_21378_n5552), .Y(w_mem_inst__abc_21378_n5553) );
  AND2X2 AND2X2_5047 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf58), .B(w_mem_inst_w_mem_3__16_), .Y(w_mem_inst__abc_21378_n5556) );
  AND2X2 AND2X2_5048 ( .A(w_mem_inst__abc_21378_n3152_bF_buf46), .B(w_mem_inst_w_mem_4__16_), .Y(w_mem_inst__abc_21378_n5557) );
  AND2X2 AND2X2_5049 ( .A(round_ctr_rst_bF_buf43), .B(\block[400] ), .Y(w_mem_inst__abc_21378_n5558) );
  AND2X2 AND2X2_505 ( .A(_auto_iopadmap_cc_313_execute_26059_79_), .B(c_reg_15_), .Y(_abc_15724_n1728_1) );
  AND2X2 AND2X2_5050 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf46), .B(w_mem_inst__abc_21378_n5558), .Y(w_mem_inst__abc_21378_n5559) );
  AND2X2 AND2X2_5051 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf57), .B(w_mem_inst_w_mem_3__17_), .Y(w_mem_inst__abc_21378_n5562) );
  AND2X2 AND2X2_5052 ( .A(w_mem_inst__abc_21378_n3152_bF_buf45), .B(w_mem_inst_w_mem_4__17_), .Y(w_mem_inst__abc_21378_n5563) );
  AND2X2 AND2X2_5053 ( .A(round_ctr_rst_bF_buf42), .B(\block[401] ), .Y(w_mem_inst__abc_21378_n5564) );
  AND2X2 AND2X2_5054 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf45), .B(w_mem_inst__abc_21378_n5564), .Y(w_mem_inst__abc_21378_n5565) );
  AND2X2 AND2X2_5055 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf56), .B(w_mem_inst_w_mem_3__18_), .Y(w_mem_inst__abc_21378_n5568) );
  AND2X2 AND2X2_5056 ( .A(w_mem_inst__abc_21378_n3152_bF_buf44), .B(w_mem_inst_w_mem_4__18_), .Y(w_mem_inst__abc_21378_n5569) );
  AND2X2 AND2X2_5057 ( .A(round_ctr_rst_bF_buf41), .B(\block[402] ), .Y(w_mem_inst__abc_21378_n5570) );
  AND2X2 AND2X2_5058 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf44), .B(w_mem_inst__abc_21378_n5570), .Y(w_mem_inst__abc_21378_n5571) );
  AND2X2 AND2X2_5059 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf55), .B(w_mem_inst_w_mem_3__19_), .Y(w_mem_inst__abc_21378_n5574) );
  AND2X2 AND2X2_506 ( .A(_abc_15724_n1729), .B(_abc_15724_n1727), .Y(_abc_15724_n1730) );
  AND2X2 AND2X2_5060 ( .A(w_mem_inst__abc_21378_n3152_bF_buf43), .B(w_mem_inst_w_mem_4__19_), .Y(w_mem_inst__abc_21378_n5575) );
  AND2X2 AND2X2_5061 ( .A(round_ctr_rst_bF_buf40), .B(\block[403] ), .Y(w_mem_inst__abc_21378_n5576) );
  AND2X2 AND2X2_5062 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf43), .B(w_mem_inst__abc_21378_n5576), .Y(w_mem_inst__abc_21378_n5577) );
  AND2X2 AND2X2_5063 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf54), .B(w_mem_inst_w_mem_3__20_), .Y(w_mem_inst__abc_21378_n5580) );
  AND2X2 AND2X2_5064 ( .A(w_mem_inst__abc_21378_n3152_bF_buf42), .B(w_mem_inst_w_mem_4__20_), .Y(w_mem_inst__abc_21378_n5581) );
  AND2X2 AND2X2_5065 ( .A(round_ctr_rst_bF_buf39), .B(\block[404] ), .Y(w_mem_inst__abc_21378_n5582) );
  AND2X2 AND2X2_5066 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf42), .B(w_mem_inst__abc_21378_n5582), .Y(w_mem_inst__abc_21378_n5583) );
  AND2X2 AND2X2_5067 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf53), .B(w_mem_inst_w_mem_3__21_), .Y(w_mem_inst__abc_21378_n5586) );
  AND2X2 AND2X2_5068 ( .A(w_mem_inst__abc_21378_n3152_bF_buf41), .B(w_mem_inst_w_mem_4__21_), .Y(w_mem_inst__abc_21378_n5587) );
  AND2X2 AND2X2_5069 ( .A(round_ctr_rst_bF_buf38), .B(\block[405] ), .Y(w_mem_inst__abc_21378_n5588) );
  AND2X2 AND2X2_507 ( .A(_abc_15724_n1731), .B(_abc_15724_n1733), .Y(_abc_15724_n1734) );
  AND2X2 AND2X2_5070 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf41), .B(w_mem_inst__abc_21378_n5588), .Y(w_mem_inst__abc_21378_n5589) );
  AND2X2 AND2X2_5071 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf52), .B(w_mem_inst_w_mem_3__22_), .Y(w_mem_inst__abc_21378_n5592) );
  AND2X2 AND2X2_5072 ( .A(w_mem_inst__abc_21378_n3152_bF_buf40), .B(w_mem_inst_w_mem_4__22_), .Y(w_mem_inst__abc_21378_n5593) );
  AND2X2 AND2X2_5073 ( .A(round_ctr_rst_bF_buf37), .B(\block[406] ), .Y(w_mem_inst__abc_21378_n5594) );
  AND2X2 AND2X2_5074 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf40), .B(w_mem_inst__abc_21378_n5594), .Y(w_mem_inst__abc_21378_n5595) );
  AND2X2 AND2X2_5075 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf51), .B(w_mem_inst_w_mem_3__23_), .Y(w_mem_inst__abc_21378_n5598) );
  AND2X2 AND2X2_5076 ( .A(w_mem_inst__abc_21378_n3152_bF_buf39), .B(w_mem_inst_w_mem_4__23_), .Y(w_mem_inst__abc_21378_n5599) );
  AND2X2 AND2X2_5077 ( .A(round_ctr_rst_bF_buf36), .B(\block[407] ), .Y(w_mem_inst__abc_21378_n5600) );
  AND2X2 AND2X2_5078 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf39), .B(w_mem_inst__abc_21378_n5600), .Y(w_mem_inst__abc_21378_n5601) );
  AND2X2 AND2X2_5079 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf50), .B(w_mem_inst_w_mem_3__24_), .Y(w_mem_inst__abc_21378_n5604) );
  AND2X2 AND2X2_508 ( .A(_abc_15724_n1734), .B(digest_update_bF_buf1), .Y(_abc_15724_n1735) );
  AND2X2 AND2X2_5080 ( .A(w_mem_inst__abc_21378_n3152_bF_buf38), .B(w_mem_inst_w_mem_4__24_), .Y(w_mem_inst__abc_21378_n5605) );
  AND2X2 AND2X2_5081 ( .A(round_ctr_rst_bF_buf35), .B(\block[408] ), .Y(w_mem_inst__abc_21378_n5606) );
  AND2X2 AND2X2_5082 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf38), .B(w_mem_inst__abc_21378_n5606), .Y(w_mem_inst__abc_21378_n5607) );
  AND2X2 AND2X2_5083 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf49), .B(w_mem_inst_w_mem_3__25_), .Y(w_mem_inst__abc_21378_n5610) );
  AND2X2 AND2X2_5084 ( .A(w_mem_inst__abc_21378_n3152_bF_buf37), .B(w_mem_inst_w_mem_4__25_), .Y(w_mem_inst__abc_21378_n5611) );
  AND2X2 AND2X2_5085 ( .A(round_ctr_rst_bF_buf34), .B(\block[409] ), .Y(w_mem_inst__abc_21378_n5612) );
  AND2X2 AND2X2_5086 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf37), .B(w_mem_inst__abc_21378_n5612), .Y(w_mem_inst__abc_21378_n5613) );
  AND2X2 AND2X2_5087 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf48), .B(w_mem_inst_w_mem_3__26_), .Y(w_mem_inst__abc_21378_n5616) );
  AND2X2 AND2X2_5088 ( .A(w_mem_inst__abc_21378_n3152_bF_buf36), .B(w_mem_inst_w_mem_4__26_), .Y(w_mem_inst__abc_21378_n5617) );
  AND2X2 AND2X2_5089 ( .A(round_ctr_rst_bF_buf33), .B(\block[410] ), .Y(w_mem_inst__abc_21378_n5618) );
  AND2X2 AND2X2_509 ( .A(_abc_15724_n1736), .B(_abc_15724_n850_bF_buf1), .Y(_abc_15724_n1737_1) );
  AND2X2 AND2X2_5090 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf36), .B(w_mem_inst__abc_21378_n5618), .Y(w_mem_inst__abc_21378_n5619) );
  AND2X2 AND2X2_5091 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf47), .B(w_mem_inst_w_mem_3__27_), .Y(w_mem_inst__abc_21378_n5622) );
  AND2X2 AND2X2_5092 ( .A(w_mem_inst__abc_21378_n3152_bF_buf35), .B(w_mem_inst_w_mem_4__27_), .Y(w_mem_inst__abc_21378_n5623) );
  AND2X2 AND2X2_5093 ( .A(round_ctr_rst_bF_buf32), .B(\block[411] ), .Y(w_mem_inst__abc_21378_n5624) );
  AND2X2 AND2X2_5094 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf35), .B(w_mem_inst__abc_21378_n5624), .Y(w_mem_inst__abc_21378_n5625) );
  AND2X2 AND2X2_5095 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf46), .B(w_mem_inst_w_mem_3__28_), .Y(w_mem_inst__abc_21378_n5628) );
  AND2X2 AND2X2_5096 ( .A(w_mem_inst__abc_21378_n3152_bF_buf34), .B(w_mem_inst_w_mem_4__28_), .Y(w_mem_inst__abc_21378_n5629) );
  AND2X2 AND2X2_5097 ( .A(round_ctr_rst_bF_buf31), .B(\block[412] ), .Y(w_mem_inst__abc_21378_n5630) );
  AND2X2 AND2X2_5098 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf34), .B(w_mem_inst__abc_21378_n5630), .Y(w_mem_inst__abc_21378_n5631) );
  AND2X2 AND2X2_5099 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf45), .B(w_mem_inst_w_mem_3__29_), .Y(w_mem_inst__abc_21378_n5634) );
  AND2X2 AND2X2_51 ( .A(e_reg_1_), .B(_auto_iopadmap_cc_313_execute_26059_1_), .Y(_abc_15724_n790_1) );
  AND2X2 AND2X2_510 ( .A(_abc_15724_n907_1_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_80_), .Y(_abc_15724_n1739) );
  AND2X2 AND2X2_5100 ( .A(w_mem_inst__abc_21378_n3152_bF_buf33), .B(w_mem_inst_w_mem_4__29_), .Y(w_mem_inst__abc_21378_n5635) );
  AND2X2 AND2X2_5101 ( .A(round_ctr_rst_bF_buf30), .B(\block[413] ), .Y(w_mem_inst__abc_21378_n5636) );
  AND2X2 AND2X2_5102 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf33), .B(w_mem_inst__abc_21378_n5636), .Y(w_mem_inst__abc_21378_n5637) );
  AND2X2 AND2X2_5103 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf44), .B(w_mem_inst_w_mem_3__30_), .Y(w_mem_inst__abc_21378_n5640) );
  AND2X2 AND2X2_5104 ( .A(w_mem_inst__abc_21378_n3152_bF_buf32), .B(w_mem_inst_w_mem_4__30_), .Y(w_mem_inst__abc_21378_n5641) );
  AND2X2 AND2X2_5105 ( .A(round_ctr_rst_bF_buf29), .B(\block[414] ), .Y(w_mem_inst__abc_21378_n5642) );
  AND2X2 AND2X2_5106 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf32), .B(w_mem_inst__abc_21378_n5642), .Y(w_mem_inst__abc_21378_n5643) );
  AND2X2 AND2X2_5107 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf43), .B(w_mem_inst_w_mem_3__31_), .Y(w_mem_inst__abc_21378_n5646) );
  AND2X2 AND2X2_5108 ( .A(w_mem_inst__abc_21378_n3152_bF_buf31), .B(w_mem_inst_w_mem_4__31_), .Y(w_mem_inst__abc_21378_n5647) );
  AND2X2 AND2X2_5109 ( .A(round_ctr_rst_bF_buf28), .B(\block[415] ), .Y(w_mem_inst__abc_21378_n5648) );
  AND2X2 AND2X2_511 ( .A(_abc_15724_n1698), .B(_abc_15724_n1687), .Y(_abc_15724_n1740) );
  AND2X2 AND2X2_5110 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf31), .B(w_mem_inst__abc_21378_n5648), .Y(w_mem_inst__abc_21378_n5649) );
  AND2X2 AND2X2_5111 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf42), .B(w_mem_inst_w_mem_2__0_), .Y(w_mem_inst__abc_21378_n5652) );
  AND2X2 AND2X2_5112 ( .A(w_mem_inst__abc_21378_n3152_bF_buf30), .B(w_mem_inst_w_mem_3__0_), .Y(w_mem_inst__abc_21378_n5653) );
  AND2X2 AND2X2_5113 ( .A(round_ctr_rst_bF_buf27), .B(\block[416] ), .Y(w_mem_inst__abc_21378_n5654) );
  AND2X2 AND2X2_5114 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf30), .B(w_mem_inst__abc_21378_n5654), .Y(w_mem_inst__abc_21378_n5655) );
  AND2X2 AND2X2_5115 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf41), .B(w_mem_inst_w_mem_2__1_), .Y(w_mem_inst__abc_21378_n5658) );
  AND2X2 AND2X2_5116 ( .A(w_mem_inst__abc_21378_n3152_bF_buf29), .B(w_mem_inst_w_mem_3__1_), .Y(w_mem_inst__abc_21378_n5659) );
  AND2X2 AND2X2_5117 ( .A(round_ctr_rst_bF_buf26), .B(\block[417] ), .Y(w_mem_inst__abc_21378_n5660) );
  AND2X2 AND2X2_5118 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf29), .B(w_mem_inst__abc_21378_n5660), .Y(w_mem_inst__abc_21378_n5661) );
  AND2X2 AND2X2_5119 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf40), .B(w_mem_inst_w_mem_2__2_), .Y(w_mem_inst__abc_21378_n5664) );
  AND2X2 AND2X2_512 ( .A(_abc_15724_n1716), .B(_abc_15724_n1730), .Y(_abc_15724_n1742) );
  AND2X2 AND2X2_5120 ( .A(w_mem_inst__abc_21378_n3152_bF_buf28), .B(w_mem_inst_w_mem_3__2_), .Y(w_mem_inst__abc_21378_n5665) );
  AND2X2 AND2X2_5121 ( .A(round_ctr_rst_bF_buf25), .B(\block[418] ), .Y(w_mem_inst__abc_21378_n5666) );
  AND2X2 AND2X2_5122 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf28), .B(w_mem_inst__abc_21378_n5666), .Y(w_mem_inst__abc_21378_n5667) );
  AND2X2 AND2X2_5123 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf39), .B(w_mem_inst_w_mem_2__3_), .Y(w_mem_inst__abc_21378_n5670) );
  AND2X2 AND2X2_5124 ( .A(w_mem_inst__abc_21378_n3152_bF_buf27), .B(w_mem_inst_w_mem_3__3_), .Y(w_mem_inst__abc_21378_n5671) );
  AND2X2 AND2X2_5125 ( .A(round_ctr_rst_bF_buf24), .B(\block[419] ), .Y(w_mem_inst__abc_21378_n5672) );
  AND2X2 AND2X2_5126 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf27), .B(w_mem_inst__abc_21378_n5672), .Y(w_mem_inst__abc_21378_n5673) );
  AND2X2 AND2X2_5127 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf38), .B(w_mem_inst_w_mem_2__4_), .Y(w_mem_inst__abc_21378_n5676) );
  AND2X2 AND2X2_5128 ( .A(w_mem_inst__abc_21378_n3152_bF_buf26), .B(w_mem_inst_w_mem_3__4_), .Y(w_mem_inst__abc_21378_n5677) );
  AND2X2 AND2X2_5129 ( .A(round_ctr_rst_bF_buf23), .B(\block[420] ), .Y(w_mem_inst__abc_21378_n5678) );
  AND2X2 AND2X2_513 ( .A(_abc_15724_n1742), .B(_abc_15724_n1741_1), .Y(_abc_15724_n1743) );
  AND2X2 AND2X2_5130 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf26), .B(w_mem_inst__abc_21378_n5678), .Y(w_mem_inst__abc_21378_n5679) );
  AND2X2 AND2X2_5131 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf37), .B(w_mem_inst_w_mem_2__5_), .Y(w_mem_inst__abc_21378_n5682) );
  AND2X2 AND2X2_5132 ( .A(w_mem_inst__abc_21378_n3152_bF_buf25), .B(w_mem_inst_w_mem_3__5_), .Y(w_mem_inst__abc_21378_n5683) );
  AND2X2 AND2X2_5133 ( .A(round_ctr_rst_bF_buf22), .B(\block[421] ), .Y(w_mem_inst__abc_21378_n5684) );
  AND2X2 AND2X2_5134 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf25), .B(w_mem_inst__abc_21378_n5684), .Y(w_mem_inst__abc_21378_n5685) );
  AND2X2 AND2X2_5135 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf36), .B(w_mem_inst_w_mem_2__6_), .Y(w_mem_inst__abc_21378_n5688) );
  AND2X2 AND2X2_5136 ( .A(w_mem_inst__abc_21378_n3152_bF_buf24), .B(w_mem_inst_w_mem_3__6_), .Y(w_mem_inst__abc_21378_n5689) );
  AND2X2 AND2X2_5137 ( .A(round_ctr_rst_bF_buf21), .B(\block[422] ), .Y(w_mem_inst__abc_21378_n5690) );
  AND2X2 AND2X2_5138 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf24), .B(w_mem_inst__abc_21378_n5690), .Y(w_mem_inst__abc_21378_n5691) );
  AND2X2 AND2X2_5139 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf35), .B(w_mem_inst_w_mem_2__7_), .Y(w_mem_inst__abc_21378_n5694) );
  AND2X2 AND2X2_514 ( .A(_abc_15724_n1727), .B(_abc_15724_n1714_1), .Y(_abc_15724_n1744) );
  AND2X2 AND2X2_5140 ( .A(w_mem_inst__abc_21378_n3152_bF_buf23), .B(w_mem_inst_w_mem_3__7_), .Y(w_mem_inst__abc_21378_n5695) );
  AND2X2 AND2X2_5141 ( .A(round_ctr_rst_bF_buf20), .B(\block[423] ), .Y(w_mem_inst__abc_21378_n5696) );
  AND2X2 AND2X2_5142 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf23), .B(w_mem_inst__abc_21378_n5696), .Y(w_mem_inst__abc_21378_n5697) );
  AND2X2 AND2X2_5143 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf34), .B(w_mem_inst_w_mem_2__8_), .Y(w_mem_inst__abc_21378_n5700) );
  AND2X2 AND2X2_5144 ( .A(w_mem_inst__abc_21378_n3152_bF_buf22), .B(w_mem_inst_w_mem_3__8_), .Y(w_mem_inst__abc_21378_n5701) );
  AND2X2 AND2X2_5145 ( .A(round_ctr_rst_bF_buf19), .B(\block[424] ), .Y(w_mem_inst__abc_21378_n5702) );
  AND2X2 AND2X2_5146 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf22), .B(w_mem_inst__abc_21378_n5702), .Y(w_mem_inst__abc_21378_n5703) );
  AND2X2 AND2X2_5147 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf33), .B(w_mem_inst_w_mem_2__9_), .Y(w_mem_inst__abc_21378_n5706) );
  AND2X2 AND2X2_5148 ( .A(w_mem_inst__abc_21378_n3152_bF_buf21), .B(w_mem_inst_w_mem_3__9_), .Y(w_mem_inst__abc_21378_n5707) );
  AND2X2 AND2X2_5149 ( .A(round_ctr_rst_bF_buf18), .B(\block[425] ), .Y(w_mem_inst__abc_21378_n5708) );
  AND2X2 AND2X2_515 ( .A(_abc_15724_n1689), .B(_abc_15724_n1701), .Y(_abc_15724_n1748) );
  AND2X2 AND2X2_5150 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf21), .B(w_mem_inst__abc_21378_n5708), .Y(w_mem_inst__abc_21378_n5709) );
  AND2X2 AND2X2_5151 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf32), .B(w_mem_inst_w_mem_2__10_), .Y(w_mem_inst__abc_21378_n5712) );
  AND2X2 AND2X2_5152 ( .A(w_mem_inst__abc_21378_n3152_bF_buf20), .B(w_mem_inst_w_mem_3__10_), .Y(w_mem_inst__abc_21378_n5713) );
  AND2X2 AND2X2_5153 ( .A(round_ctr_rst_bF_buf17), .B(\block[426] ), .Y(w_mem_inst__abc_21378_n5714) );
  AND2X2 AND2X2_5154 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf20), .B(w_mem_inst__abc_21378_n5714), .Y(w_mem_inst__abc_21378_n5715) );
  AND2X2 AND2X2_5155 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf31), .B(w_mem_inst_w_mem_2__11_), .Y(w_mem_inst__abc_21378_n5718) );
  AND2X2 AND2X2_5156 ( .A(w_mem_inst__abc_21378_n3152_bF_buf19), .B(w_mem_inst_w_mem_3__11_), .Y(w_mem_inst__abc_21378_n5719) );
  AND2X2 AND2X2_5157 ( .A(round_ctr_rst_bF_buf16), .B(\block[427] ), .Y(w_mem_inst__abc_21378_n5720) );
  AND2X2 AND2X2_5158 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf19), .B(w_mem_inst__abc_21378_n5720), .Y(w_mem_inst__abc_21378_n5721) );
  AND2X2 AND2X2_5159 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf30), .B(w_mem_inst_w_mem_2__12_), .Y(w_mem_inst__abc_21378_n5724) );
  AND2X2 AND2X2_516 ( .A(_abc_15724_n1748), .B(_abc_15724_n1742), .Y(_abc_15724_n1749) );
  AND2X2 AND2X2_5160 ( .A(w_mem_inst__abc_21378_n3152_bF_buf18), .B(w_mem_inst_w_mem_3__12_), .Y(w_mem_inst__abc_21378_n5725) );
  AND2X2 AND2X2_5161 ( .A(round_ctr_rst_bF_buf15), .B(\block[428] ), .Y(w_mem_inst__abc_21378_n5726) );
  AND2X2 AND2X2_5162 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf18), .B(w_mem_inst__abc_21378_n5726), .Y(w_mem_inst__abc_21378_n5727) );
  AND2X2 AND2X2_5163 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf29), .B(w_mem_inst_w_mem_2__13_), .Y(w_mem_inst__abc_21378_n5730) );
  AND2X2 AND2X2_5164 ( .A(w_mem_inst__abc_21378_n3152_bF_buf17), .B(w_mem_inst_w_mem_3__13_), .Y(w_mem_inst__abc_21378_n5731) );
  AND2X2 AND2X2_5165 ( .A(round_ctr_rst_bF_buf14), .B(\block[429] ), .Y(w_mem_inst__abc_21378_n5732) );
  AND2X2 AND2X2_5166 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf17), .B(w_mem_inst__abc_21378_n5732), .Y(w_mem_inst__abc_21378_n5733) );
  AND2X2 AND2X2_5167 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf28), .B(w_mem_inst_w_mem_2__14_), .Y(w_mem_inst__abc_21378_n5736) );
  AND2X2 AND2X2_5168 ( .A(w_mem_inst__abc_21378_n3152_bF_buf16), .B(w_mem_inst_w_mem_3__14_), .Y(w_mem_inst__abc_21378_n5737) );
  AND2X2 AND2X2_5169 ( .A(round_ctr_rst_bF_buf13), .B(\block[430] ), .Y(w_mem_inst__abc_21378_n5738) );
  AND2X2 AND2X2_517 ( .A(_abc_15724_n1751), .B(_abc_15724_n1747), .Y(_abc_15724_n1752) );
  AND2X2 AND2X2_5170 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf16), .B(w_mem_inst__abc_21378_n5738), .Y(w_mem_inst__abc_21378_n5739) );
  AND2X2 AND2X2_5171 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf27), .B(w_mem_inst_w_mem_2__15_), .Y(w_mem_inst__abc_21378_n5742) );
  AND2X2 AND2X2_5172 ( .A(w_mem_inst__abc_21378_n3152_bF_buf15), .B(w_mem_inst_w_mem_3__15_), .Y(w_mem_inst__abc_21378_n5743) );
  AND2X2 AND2X2_5173 ( .A(round_ctr_rst_bF_buf12), .B(\block[431] ), .Y(w_mem_inst__abc_21378_n5744) );
  AND2X2 AND2X2_5174 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf15), .B(w_mem_inst__abc_21378_n5744), .Y(w_mem_inst__abc_21378_n5745) );
  AND2X2 AND2X2_5175 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf26), .B(w_mem_inst_w_mem_2__16_), .Y(w_mem_inst__abc_21378_n5748) );
  AND2X2 AND2X2_5176 ( .A(w_mem_inst__abc_21378_n3152_bF_buf14), .B(w_mem_inst_w_mem_3__16_), .Y(w_mem_inst__abc_21378_n5749) );
  AND2X2 AND2X2_5177 ( .A(round_ctr_rst_bF_buf11), .B(\block[432] ), .Y(w_mem_inst__abc_21378_n5750) );
  AND2X2 AND2X2_5178 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf14), .B(w_mem_inst__abc_21378_n5750), .Y(w_mem_inst__abc_21378_n5751) );
  AND2X2 AND2X2_5179 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf25), .B(w_mem_inst_w_mem_2__17_), .Y(w_mem_inst__abc_21378_n5754) );
  AND2X2 AND2X2_518 ( .A(_auto_iopadmap_cc_313_execute_26059_80_), .B(c_reg_16_), .Y(_abc_15724_n1755) );
  AND2X2 AND2X2_5180 ( .A(w_mem_inst__abc_21378_n3152_bF_buf13), .B(w_mem_inst_w_mem_3__17_), .Y(w_mem_inst__abc_21378_n5755) );
  AND2X2 AND2X2_5181 ( .A(round_ctr_rst_bF_buf10), .B(\block[433] ), .Y(w_mem_inst__abc_21378_n5756) );
  AND2X2 AND2X2_5182 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf13), .B(w_mem_inst__abc_21378_n5756), .Y(w_mem_inst__abc_21378_n5757) );
  AND2X2 AND2X2_5183 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf24), .B(w_mem_inst_w_mem_2__18_), .Y(w_mem_inst__abc_21378_n5760) );
  AND2X2 AND2X2_5184 ( .A(w_mem_inst__abc_21378_n3152_bF_buf12), .B(w_mem_inst_w_mem_3__18_), .Y(w_mem_inst__abc_21378_n5761) );
  AND2X2 AND2X2_5185 ( .A(round_ctr_rst_bF_buf9), .B(\block[434] ), .Y(w_mem_inst__abc_21378_n5762) );
  AND2X2 AND2X2_5186 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf12), .B(w_mem_inst__abc_21378_n5762), .Y(w_mem_inst__abc_21378_n5763) );
  AND2X2 AND2X2_5187 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf23), .B(w_mem_inst_w_mem_2__19_), .Y(w_mem_inst__abc_21378_n5766) );
  AND2X2 AND2X2_5188 ( .A(w_mem_inst__abc_21378_n3152_bF_buf11), .B(w_mem_inst_w_mem_3__19_), .Y(w_mem_inst__abc_21378_n5767) );
  AND2X2 AND2X2_5189 ( .A(round_ctr_rst_bF_buf8), .B(\block[435] ), .Y(w_mem_inst__abc_21378_n5768) );
  AND2X2 AND2X2_519 ( .A(_abc_15724_n1756), .B(_abc_15724_n1754_1), .Y(_abc_15724_n1757) );
  AND2X2 AND2X2_5190 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf11), .B(w_mem_inst__abc_21378_n5768), .Y(w_mem_inst__abc_21378_n5769) );
  AND2X2 AND2X2_5191 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf22), .B(w_mem_inst_w_mem_2__20_), .Y(w_mem_inst__abc_21378_n5772) );
  AND2X2 AND2X2_5192 ( .A(w_mem_inst__abc_21378_n3152_bF_buf10), .B(w_mem_inst_w_mem_3__20_), .Y(w_mem_inst__abc_21378_n5773) );
  AND2X2 AND2X2_5193 ( .A(round_ctr_rst_bF_buf7), .B(\block[436] ), .Y(w_mem_inst__abc_21378_n5774) );
  AND2X2 AND2X2_5194 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf10), .B(w_mem_inst__abc_21378_n5774), .Y(w_mem_inst__abc_21378_n5775) );
  AND2X2 AND2X2_5195 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf21), .B(w_mem_inst_w_mem_2__21_), .Y(w_mem_inst__abc_21378_n5778) );
  AND2X2 AND2X2_5196 ( .A(w_mem_inst__abc_21378_n3152_bF_buf9), .B(w_mem_inst_w_mem_3__21_), .Y(w_mem_inst__abc_21378_n5779) );
  AND2X2 AND2X2_5197 ( .A(round_ctr_rst_bF_buf6), .B(\block[437] ), .Y(w_mem_inst__abc_21378_n5780) );
  AND2X2 AND2X2_5198 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf9), .B(w_mem_inst__abc_21378_n5780), .Y(w_mem_inst__abc_21378_n5781) );
  AND2X2 AND2X2_5199 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf20), .B(w_mem_inst_w_mem_2__22_), .Y(w_mem_inst__abc_21378_n5784) );
  AND2X2 AND2X2_52 ( .A(e_reg_0_), .B(_auto_iopadmap_cc_313_execute_26059_0_), .Y(_abc_15724_n792) );
  AND2X2 AND2X2_520 ( .A(_abc_15724_n1753), .B(_abc_15724_n1757), .Y(_abc_15724_n1759) );
  AND2X2 AND2X2_5200 ( .A(w_mem_inst__abc_21378_n3152_bF_buf8), .B(w_mem_inst_w_mem_3__22_), .Y(w_mem_inst__abc_21378_n5785) );
  AND2X2 AND2X2_5201 ( .A(round_ctr_rst_bF_buf5), .B(\block[438] ), .Y(w_mem_inst__abc_21378_n5786) );
  AND2X2 AND2X2_5202 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf8), .B(w_mem_inst__abc_21378_n5786), .Y(w_mem_inst__abc_21378_n5787) );
  AND2X2 AND2X2_5203 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf19), .B(w_mem_inst_w_mem_2__23_), .Y(w_mem_inst__abc_21378_n5790) );
  AND2X2 AND2X2_5204 ( .A(w_mem_inst__abc_21378_n3152_bF_buf7), .B(w_mem_inst_w_mem_3__23_), .Y(w_mem_inst__abc_21378_n5791) );
  AND2X2 AND2X2_5205 ( .A(round_ctr_rst_bF_buf4), .B(\block[439] ), .Y(w_mem_inst__abc_21378_n5792) );
  AND2X2 AND2X2_5206 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf7), .B(w_mem_inst__abc_21378_n5792), .Y(w_mem_inst__abc_21378_n5793) );
  AND2X2 AND2X2_5207 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf18), .B(w_mem_inst_w_mem_2__24_), .Y(w_mem_inst__abc_21378_n5796) );
  AND2X2 AND2X2_5208 ( .A(w_mem_inst__abc_21378_n3152_bF_buf6), .B(w_mem_inst_w_mem_3__24_), .Y(w_mem_inst__abc_21378_n5797) );
  AND2X2 AND2X2_5209 ( .A(round_ctr_rst_bF_buf3), .B(\block[440] ), .Y(w_mem_inst__abc_21378_n5798) );
  AND2X2 AND2X2_521 ( .A(_abc_15724_n1760), .B(_abc_15724_n1758_1), .Y(_abc_15724_n1761) );
  AND2X2 AND2X2_5210 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf6), .B(w_mem_inst__abc_21378_n5798), .Y(w_mem_inst__abc_21378_n5799) );
  AND2X2 AND2X2_5211 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf17), .B(w_mem_inst_w_mem_2__25_), .Y(w_mem_inst__abc_21378_n5802) );
  AND2X2 AND2X2_5212 ( .A(w_mem_inst__abc_21378_n3152_bF_buf5), .B(w_mem_inst_w_mem_3__25_), .Y(w_mem_inst__abc_21378_n5803) );
  AND2X2 AND2X2_5213 ( .A(round_ctr_rst_bF_buf2), .B(\block[441] ), .Y(w_mem_inst__abc_21378_n5804) );
  AND2X2 AND2X2_5214 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf5), .B(w_mem_inst__abc_21378_n5804), .Y(w_mem_inst__abc_21378_n5805) );
  AND2X2 AND2X2_5215 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf16), .B(w_mem_inst_w_mem_2__26_), .Y(w_mem_inst__abc_21378_n5808) );
  AND2X2 AND2X2_5216 ( .A(w_mem_inst__abc_21378_n3152_bF_buf4), .B(w_mem_inst_w_mem_3__26_), .Y(w_mem_inst__abc_21378_n5809) );
  AND2X2 AND2X2_5217 ( .A(round_ctr_rst_bF_buf1), .B(\block[442] ), .Y(w_mem_inst__abc_21378_n5810) );
  AND2X2 AND2X2_5218 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf4), .B(w_mem_inst__abc_21378_n5810), .Y(w_mem_inst__abc_21378_n5811) );
  AND2X2 AND2X2_5219 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf15), .B(w_mem_inst_w_mem_2__27_), .Y(w_mem_inst__abc_21378_n5814) );
  AND2X2 AND2X2_522 ( .A(_abc_15724_n1761), .B(digest_update_bF_buf0), .Y(_abc_15724_n1762_1) );
  AND2X2 AND2X2_5220 ( .A(w_mem_inst__abc_21378_n3152_bF_buf3), .B(w_mem_inst_w_mem_3__27_), .Y(w_mem_inst__abc_21378_n5815) );
  AND2X2 AND2X2_5221 ( .A(round_ctr_rst_bF_buf0), .B(\block[443] ), .Y(w_mem_inst__abc_21378_n5816) );
  AND2X2 AND2X2_5222 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf3), .B(w_mem_inst__abc_21378_n5816), .Y(w_mem_inst__abc_21378_n5817) );
  AND2X2 AND2X2_5223 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf14), .B(w_mem_inst_w_mem_2__28_), .Y(w_mem_inst__abc_21378_n5820) );
  AND2X2 AND2X2_5224 ( .A(w_mem_inst__abc_21378_n3152_bF_buf2), .B(w_mem_inst_w_mem_3__28_), .Y(w_mem_inst__abc_21378_n5821) );
  AND2X2 AND2X2_5225 ( .A(round_ctr_rst_bF_buf63), .B(\block[444] ), .Y(w_mem_inst__abc_21378_n5822) );
  AND2X2 AND2X2_5226 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf2), .B(w_mem_inst__abc_21378_n5822), .Y(w_mem_inst__abc_21378_n5823) );
  AND2X2 AND2X2_5227 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf13), .B(w_mem_inst_w_mem_2__29_), .Y(w_mem_inst__abc_21378_n5826) );
  AND2X2 AND2X2_5228 ( .A(w_mem_inst__abc_21378_n3152_bF_buf1), .B(w_mem_inst_w_mem_3__29_), .Y(w_mem_inst__abc_21378_n5827) );
  AND2X2 AND2X2_5229 ( .A(round_ctr_rst_bF_buf62), .B(\block[445] ), .Y(w_mem_inst__abc_21378_n5828) );
  AND2X2 AND2X2_523 ( .A(_abc_15724_n1760), .B(_abc_15724_n1756), .Y(_abc_15724_n1764) );
  AND2X2 AND2X2_5230 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf1), .B(w_mem_inst__abc_21378_n5828), .Y(w_mem_inst__abc_21378_n5829) );
  AND2X2 AND2X2_5231 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf12), .B(w_mem_inst_w_mem_2__30_), .Y(w_mem_inst__abc_21378_n5832) );
  AND2X2 AND2X2_5232 ( .A(w_mem_inst__abc_21378_n3152_bF_buf0), .B(w_mem_inst_w_mem_3__30_), .Y(w_mem_inst__abc_21378_n5833) );
  AND2X2 AND2X2_5233 ( .A(round_ctr_rst_bF_buf61), .B(\block[446] ), .Y(w_mem_inst__abc_21378_n5834) );
  AND2X2 AND2X2_5234 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf0), .B(w_mem_inst__abc_21378_n5834), .Y(w_mem_inst__abc_21378_n5835) );
  AND2X2 AND2X2_5235 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf11), .B(w_mem_inst_w_mem_2__31_), .Y(w_mem_inst__abc_21378_n5838) );
  AND2X2 AND2X2_5236 ( .A(w_mem_inst__abc_21378_n3152_bF_buf63), .B(w_mem_inst_w_mem_3__31_), .Y(w_mem_inst__abc_21378_n5839) );
  AND2X2 AND2X2_5237 ( .A(round_ctr_rst_bF_buf60), .B(\block[447] ), .Y(w_mem_inst__abc_21378_n5840) );
  AND2X2 AND2X2_5238 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf63), .B(w_mem_inst__abc_21378_n5840), .Y(w_mem_inst__abc_21378_n5841) );
  AND2X2 AND2X2_5239 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf10), .B(w_mem_inst_w_mem_1__0_), .Y(w_mem_inst__abc_21378_n5844) );
  AND2X2 AND2X2_524 ( .A(_auto_iopadmap_cc_313_execute_26059_81_), .B(c_reg_17_), .Y(_abc_15724_n1767_1) );
  AND2X2 AND2X2_5240 ( .A(w_mem_inst__abc_21378_n3152_bF_buf62), .B(w_mem_inst_w_mem_2__0_), .Y(w_mem_inst__abc_21378_n5845) );
  AND2X2 AND2X2_5241 ( .A(round_ctr_rst_bF_buf59), .B(\block[448] ), .Y(w_mem_inst__abc_21378_n5846) );
  AND2X2 AND2X2_5242 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf62), .B(w_mem_inst__abc_21378_n5846), .Y(w_mem_inst__abc_21378_n5847) );
  AND2X2 AND2X2_5243 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf9), .B(w_mem_inst_w_mem_1__1_), .Y(w_mem_inst__abc_21378_n5850) );
  AND2X2 AND2X2_5244 ( .A(w_mem_inst__abc_21378_n3152_bF_buf61), .B(w_mem_inst_w_mem_2__1_), .Y(w_mem_inst__abc_21378_n5851) );
  AND2X2 AND2X2_5245 ( .A(round_ctr_rst_bF_buf58), .B(\block[449] ), .Y(w_mem_inst__abc_21378_n5852) );
  AND2X2 AND2X2_5246 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf61), .B(w_mem_inst__abc_21378_n5852), .Y(w_mem_inst__abc_21378_n5853) );
  AND2X2 AND2X2_5247 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf8), .B(w_mem_inst_w_mem_1__2_), .Y(w_mem_inst__abc_21378_n5856) );
  AND2X2 AND2X2_5248 ( .A(w_mem_inst__abc_21378_n3152_bF_buf60), .B(w_mem_inst_w_mem_2__2_), .Y(w_mem_inst__abc_21378_n5857) );
  AND2X2 AND2X2_5249 ( .A(round_ctr_rst_bF_buf57), .B(\block[450] ), .Y(w_mem_inst__abc_21378_n5858) );
  AND2X2 AND2X2_525 ( .A(_abc_15724_n1768), .B(_abc_15724_n1766), .Y(_abc_15724_n1769) );
  AND2X2 AND2X2_5250 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf60), .B(w_mem_inst__abc_21378_n5858), .Y(w_mem_inst__abc_21378_n5859) );
  AND2X2 AND2X2_5251 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf7), .B(w_mem_inst_w_mem_1__3_), .Y(w_mem_inst__abc_21378_n5862) );
  AND2X2 AND2X2_5252 ( .A(w_mem_inst__abc_21378_n3152_bF_buf59), .B(w_mem_inst_w_mem_2__3_), .Y(w_mem_inst__abc_21378_n5863) );
  AND2X2 AND2X2_5253 ( .A(round_ctr_rst_bF_buf56), .B(\block[451] ), .Y(w_mem_inst__abc_21378_n5864) );
  AND2X2 AND2X2_5254 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf59), .B(w_mem_inst__abc_21378_n5864), .Y(w_mem_inst__abc_21378_n5865) );
  AND2X2 AND2X2_5255 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf6), .B(w_mem_inst_w_mem_1__4_), .Y(w_mem_inst__abc_21378_n5868) );
  AND2X2 AND2X2_5256 ( .A(w_mem_inst__abc_21378_n3152_bF_buf58), .B(w_mem_inst_w_mem_2__4_), .Y(w_mem_inst__abc_21378_n5869) );
  AND2X2 AND2X2_5257 ( .A(round_ctr_rst_bF_buf55), .B(\block[452] ), .Y(w_mem_inst__abc_21378_n5870) );
  AND2X2 AND2X2_5258 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf58), .B(w_mem_inst__abc_21378_n5870), .Y(w_mem_inst__abc_21378_n5871) );
  AND2X2 AND2X2_5259 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf5), .B(w_mem_inst_w_mem_1__5_), .Y(w_mem_inst__abc_21378_n5874) );
  AND2X2 AND2X2_526 ( .A(_abc_15724_n1770), .B(_abc_15724_n1772_1), .Y(_abc_15724_n1773) );
  AND2X2 AND2X2_5260 ( .A(w_mem_inst__abc_21378_n3152_bF_buf57), .B(w_mem_inst_w_mem_2__5_), .Y(w_mem_inst__abc_21378_n5875) );
  AND2X2 AND2X2_5261 ( .A(round_ctr_rst_bF_buf54), .B(\block[453] ), .Y(w_mem_inst__abc_21378_n5876) );
  AND2X2 AND2X2_5262 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf57), .B(w_mem_inst__abc_21378_n5876), .Y(w_mem_inst__abc_21378_n5877) );
  AND2X2 AND2X2_5263 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf4), .B(w_mem_inst_w_mem_1__6_), .Y(w_mem_inst__abc_21378_n5880) );
  AND2X2 AND2X2_5264 ( .A(w_mem_inst__abc_21378_n3152_bF_buf56), .B(w_mem_inst_w_mem_2__6_), .Y(w_mem_inst__abc_21378_n5881) );
  AND2X2 AND2X2_5265 ( .A(round_ctr_rst_bF_buf53), .B(\block[454] ), .Y(w_mem_inst__abc_21378_n5882) );
  AND2X2 AND2X2_5266 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf56), .B(w_mem_inst__abc_21378_n5882), .Y(w_mem_inst__abc_21378_n5883) );
  AND2X2 AND2X2_5267 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf3), .B(w_mem_inst_w_mem_1__7_), .Y(w_mem_inst__abc_21378_n5886) );
  AND2X2 AND2X2_5268 ( .A(w_mem_inst__abc_21378_n3152_bF_buf55), .B(w_mem_inst_w_mem_2__7_), .Y(w_mem_inst__abc_21378_n5887) );
  AND2X2 AND2X2_5269 ( .A(round_ctr_rst_bF_buf52), .B(\block[455] ), .Y(w_mem_inst__abc_21378_n5888) );
  AND2X2 AND2X2_527 ( .A(_abc_15724_n1773), .B(digest_update_bF_buf11), .Y(_abc_15724_n1774) );
  AND2X2 AND2X2_5270 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf55), .B(w_mem_inst__abc_21378_n5888), .Y(w_mem_inst__abc_21378_n5889) );
  AND2X2 AND2X2_5271 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf2), .B(w_mem_inst_w_mem_1__8_), .Y(w_mem_inst__abc_21378_n5892) );
  AND2X2 AND2X2_5272 ( .A(w_mem_inst__abc_21378_n3152_bF_buf54), .B(w_mem_inst_w_mem_2__8_), .Y(w_mem_inst__abc_21378_n5893) );
  AND2X2 AND2X2_5273 ( .A(round_ctr_rst_bF_buf51), .B(\block[456] ), .Y(w_mem_inst__abc_21378_n5894) );
  AND2X2 AND2X2_5274 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf54), .B(w_mem_inst__abc_21378_n5894), .Y(w_mem_inst__abc_21378_n5895) );
  AND2X2 AND2X2_5275 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf1), .B(w_mem_inst_w_mem_1__9_), .Y(w_mem_inst__abc_21378_n5898) );
  AND2X2 AND2X2_5276 ( .A(w_mem_inst__abc_21378_n3152_bF_buf53), .B(w_mem_inst_w_mem_2__9_), .Y(w_mem_inst__abc_21378_n5899) );
  AND2X2 AND2X2_5277 ( .A(round_ctr_rst_bF_buf50), .B(\block[457] ), .Y(w_mem_inst__abc_21378_n5900) );
  AND2X2 AND2X2_5278 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf53), .B(w_mem_inst__abc_21378_n5900), .Y(w_mem_inst__abc_21378_n5901) );
  AND2X2 AND2X2_5279 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf0), .B(w_mem_inst_w_mem_1__10_), .Y(w_mem_inst__abc_21378_n5904) );
  AND2X2 AND2X2_528 ( .A(_abc_15724_n1775), .B(_abc_15724_n850_bF_buf0), .Y(_abc_15724_n1776) );
  AND2X2 AND2X2_5280 ( .A(w_mem_inst__abc_21378_n3152_bF_buf52), .B(w_mem_inst_w_mem_2__10_), .Y(w_mem_inst__abc_21378_n5905) );
  AND2X2 AND2X2_5281 ( .A(round_ctr_rst_bF_buf49), .B(\block[458] ), .Y(w_mem_inst__abc_21378_n5906) );
  AND2X2 AND2X2_5282 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf52), .B(w_mem_inst__abc_21378_n5906), .Y(w_mem_inst__abc_21378_n5907) );
  AND2X2 AND2X2_5283 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf60), .B(w_mem_inst_w_mem_1__11_), .Y(w_mem_inst__abc_21378_n5910) );
  AND2X2 AND2X2_5284 ( .A(w_mem_inst__abc_21378_n3152_bF_buf51), .B(w_mem_inst_w_mem_2__11_), .Y(w_mem_inst__abc_21378_n5911) );
  AND2X2 AND2X2_5285 ( .A(round_ctr_rst_bF_buf48), .B(\block[459] ), .Y(w_mem_inst__abc_21378_n5912) );
  AND2X2 AND2X2_5286 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf51), .B(w_mem_inst__abc_21378_n5912), .Y(w_mem_inst__abc_21378_n5913) );
  AND2X2 AND2X2_5287 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf59), .B(w_mem_inst_w_mem_1__12_), .Y(w_mem_inst__abc_21378_n5916) );
  AND2X2 AND2X2_5288 ( .A(w_mem_inst__abc_21378_n3152_bF_buf50), .B(w_mem_inst_w_mem_2__12_), .Y(w_mem_inst__abc_21378_n5917) );
  AND2X2 AND2X2_5289 ( .A(round_ctr_rst_bF_buf47), .B(\block[460] ), .Y(w_mem_inst__abc_21378_n5918) );
  AND2X2 AND2X2_529 ( .A(_abc_15724_n907_1_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_82_), .Y(_abc_15724_n1778) );
  AND2X2 AND2X2_5290 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf50), .B(w_mem_inst__abc_21378_n5918), .Y(w_mem_inst__abc_21378_n5919) );
  AND2X2 AND2X2_5291 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf58), .B(w_mem_inst_w_mem_1__13_), .Y(w_mem_inst__abc_21378_n5922) );
  AND2X2 AND2X2_5292 ( .A(w_mem_inst__abc_21378_n3152_bF_buf49), .B(w_mem_inst_w_mem_2__13_), .Y(w_mem_inst__abc_21378_n5923) );
  AND2X2 AND2X2_5293 ( .A(round_ctr_rst_bF_buf46), .B(\block[461] ), .Y(w_mem_inst__abc_21378_n5924) );
  AND2X2 AND2X2_5294 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf49), .B(w_mem_inst__abc_21378_n5924), .Y(w_mem_inst__abc_21378_n5925) );
  AND2X2 AND2X2_5295 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf57), .B(w_mem_inst_w_mem_1__14_), .Y(w_mem_inst__abc_21378_n5928) );
  AND2X2 AND2X2_5296 ( .A(w_mem_inst__abc_21378_n3152_bF_buf48), .B(w_mem_inst_w_mem_2__14_), .Y(w_mem_inst__abc_21378_n5929) );
  AND2X2 AND2X2_5297 ( .A(round_ctr_rst_bF_buf45), .B(\block[462] ), .Y(w_mem_inst__abc_21378_n5930) );
  AND2X2 AND2X2_5298 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf48), .B(w_mem_inst__abc_21378_n5930), .Y(w_mem_inst__abc_21378_n5931) );
  AND2X2 AND2X2_5299 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf56), .B(w_mem_inst_w_mem_1__15_), .Y(w_mem_inst__abc_21378_n5934) );
  AND2X2 AND2X2_53 ( .A(_abc_15724_n791_1), .B(_abc_15724_n793), .Y(_abc_15724_n794) );
  AND2X2 AND2X2_530 ( .A(_abc_15724_n1779), .B(_abc_15724_n1768), .Y(_abc_15724_n1780) );
  AND2X2 AND2X2_5300 ( .A(w_mem_inst__abc_21378_n3152_bF_buf47), .B(w_mem_inst_w_mem_2__15_), .Y(w_mem_inst__abc_21378_n5935) );
  AND2X2 AND2X2_5301 ( .A(round_ctr_rst_bF_buf44), .B(\block[463] ), .Y(w_mem_inst__abc_21378_n5936) );
  AND2X2 AND2X2_5302 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf47), .B(w_mem_inst__abc_21378_n5936), .Y(w_mem_inst__abc_21378_n5937) );
  AND2X2 AND2X2_5303 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf55), .B(w_mem_inst_w_mem_1__16_), .Y(w_mem_inst__abc_21378_n5940) );
  AND2X2 AND2X2_5304 ( .A(w_mem_inst__abc_21378_n3152_bF_buf46), .B(w_mem_inst_w_mem_2__16_), .Y(w_mem_inst__abc_21378_n5941) );
  AND2X2 AND2X2_5305 ( .A(round_ctr_rst_bF_buf43), .B(\block[464] ), .Y(w_mem_inst__abc_21378_n5942) );
  AND2X2 AND2X2_5306 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf46), .B(w_mem_inst__abc_21378_n5942), .Y(w_mem_inst__abc_21378_n5943) );
  AND2X2 AND2X2_5307 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf54), .B(w_mem_inst_w_mem_1__17_), .Y(w_mem_inst__abc_21378_n5946) );
  AND2X2 AND2X2_5308 ( .A(w_mem_inst__abc_21378_n3152_bF_buf45), .B(w_mem_inst_w_mem_2__17_), .Y(w_mem_inst__abc_21378_n5947) );
  AND2X2 AND2X2_5309 ( .A(round_ctr_rst_bF_buf42), .B(\block[465] ), .Y(w_mem_inst__abc_21378_n5948) );
  AND2X2 AND2X2_531 ( .A(_abc_15724_n1757), .B(_abc_15724_n1769), .Y(_abc_15724_n1782) );
  AND2X2 AND2X2_5310 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf45), .B(w_mem_inst__abc_21378_n5948), .Y(w_mem_inst__abc_21378_n5949) );
  AND2X2 AND2X2_5311 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf53), .B(w_mem_inst_w_mem_1__18_), .Y(w_mem_inst__abc_21378_n5952) );
  AND2X2 AND2X2_5312 ( .A(w_mem_inst__abc_21378_n3152_bF_buf44), .B(w_mem_inst_w_mem_2__18_), .Y(w_mem_inst__abc_21378_n5953) );
  AND2X2 AND2X2_5313 ( .A(round_ctr_rst_bF_buf41), .B(\block[466] ), .Y(w_mem_inst__abc_21378_n5954) );
  AND2X2 AND2X2_5314 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf44), .B(w_mem_inst__abc_21378_n5954), .Y(w_mem_inst__abc_21378_n5955) );
  AND2X2 AND2X2_5315 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf52), .B(w_mem_inst_w_mem_1__19_), .Y(w_mem_inst__abc_21378_n5958) );
  AND2X2 AND2X2_5316 ( .A(w_mem_inst__abc_21378_n3152_bF_buf43), .B(w_mem_inst_w_mem_2__19_), .Y(w_mem_inst__abc_21378_n5959) );
  AND2X2 AND2X2_5317 ( .A(round_ctr_rst_bF_buf40), .B(\block[467] ), .Y(w_mem_inst__abc_21378_n5960) );
  AND2X2 AND2X2_5318 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf43), .B(w_mem_inst__abc_21378_n5960), .Y(w_mem_inst__abc_21378_n5961) );
  AND2X2 AND2X2_5319 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf51), .B(w_mem_inst_w_mem_1__20_), .Y(w_mem_inst__abc_21378_n5964) );
  AND2X2 AND2X2_532 ( .A(_abc_15724_n1753), .B(_abc_15724_n1782), .Y(_abc_15724_n1783) );
  AND2X2 AND2X2_5320 ( .A(w_mem_inst__abc_21378_n3152_bF_buf42), .B(w_mem_inst_w_mem_2__20_), .Y(w_mem_inst__abc_21378_n5965) );
  AND2X2 AND2X2_5321 ( .A(round_ctr_rst_bF_buf39), .B(\block[468] ), .Y(w_mem_inst__abc_21378_n5966) );
  AND2X2 AND2X2_5322 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf42), .B(w_mem_inst__abc_21378_n5966), .Y(w_mem_inst__abc_21378_n5967) );
  AND2X2 AND2X2_5323 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf50), .B(w_mem_inst_w_mem_1__21_), .Y(w_mem_inst__abc_21378_n5970) );
  AND2X2 AND2X2_5324 ( .A(w_mem_inst__abc_21378_n3152_bF_buf41), .B(w_mem_inst_w_mem_2__21_), .Y(w_mem_inst__abc_21378_n5971) );
  AND2X2 AND2X2_5325 ( .A(round_ctr_rst_bF_buf38), .B(\block[469] ), .Y(w_mem_inst__abc_21378_n5972) );
  AND2X2 AND2X2_5326 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf41), .B(w_mem_inst__abc_21378_n5972), .Y(w_mem_inst__abc_21378_n5973) );
  AND2X2 AND2X2_5327 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf49), .B(w_mem_inst_w_mem_1__22_), .Y(w_mem_inst__abc_21378_n5976) );
  AND2X2 AND2X2_5328 ( .A(w_mem_inst__abc_21378_n3152_bF_buf40), .B(w_mem_inst_w_mem_2__22_), .Y(w_mem_inst__abc_21378_n5977) );
  AND2X2 AND2X2_5329 ( .A(round_ctr_rst_bF_buf37), .B(\block[470] ), .Y(w_mem_inst__abc_21378_n5978) );
  AND2X2 AND2X2_533 ( .A(_auto_iopadmap_cc_313_execute_26059_82_), .B(c_reg_18_), .Y(_abc_15724_n1786_1) );
  AND2X2 AND2X2_5330 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf40), .B(w_mem_inst__abc_21378_n5978), .Y(w_mem_inst__abc_21378_n5979) );
  AND2X2 AND2X2_5331 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf48), .B(w_mem_inst_w_mem_1__23_), .Y(w_mem_inst__abc_21378_n5982) );
  AND2X2 AND2X2_5332 ( .A(w_mem_inst__abc_21378_n3152_bF_buf39), .B(w_mem_inst_w_mem_2__23_), .Y(w_mem_inst__abc_21378_n5983) );
  AND2X2 AND2X2_5333 ( .A(round_ctr_rst_bF_buf36), .B(\block[471] ), .Y(w_mem_inst__abc_21378_n5984) );
  AND2X2 AND2X2_5334 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf39), .B(w_mem_inst__abc_21378_n5984), .Y(w_mem_inst__abc_21378_n5985) );
  AND2X2 AND2X2_5335 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf47), .B(w_mem_inst_w_mem_1__24_), .Y(w_mem_inst__abc_21378_n5988) );
  AND2X2 AND2X2_5336 ( .A(w_mem_inst__abc_21378_n3152_bF_buf38), .B(w_mem_inst_w_mem_2__24_), .Y(w_mem_inst__abc_21378_n5989) );
  AND2X2 AND2X2_5337 ( .A(round_ctr_rst_bF_buf35), .B(\block[472] ), .Y(w_mem_inst__abc_21378_n5990) );
  AND2X2 AND2X2_5338 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf38), .B(w_mem_inst__abc_21378_n5990), .Y(w_mem_inst__abc_21378_n5991) );
  AND2X2 AND2X2_5339 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf46), .B(w_mem_inst_w_mem_1__25_), .Y(w_mem_inst__abc_21378_n5994) );
  AND2X2 AND2X2_534 ( .A(_abc_15724_n1787), .B(_abc_15724_n1785), .Y(_abc_15724_n1788) );
  AND2X2 AND2X2_5340 ( .A(w_mem_inst__abc_21378_n3152_bF_buf37), .B(w_mem_inst_w_mem_2__25_), .Y(w_mem_inst__abc_21378_n5995) );
  AND2X2 AND2X2_5341 ( .A(round_ctr_rst_bF_buf34), .B(\block[473] ), .Y(w_mem_inst__abc_21378_n5996) );
  AND2X2 AND2X2_5342 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf37), .B(w_mem_inst__abc_21378_n5996), .Y(w_mem_inst__abc_21378_n5997) );
  AND2X2 AND2X2_5343 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf45), .B(w_mem_inst_w_mem_1__26_), .Y(w_mem_inst__abc_21378_n6000) );
  AND2X2 AND2X2_5344 ( .A(w_mem_inst__abc_21378_n3152_bF_buf36), .B(w_mem_inst_w_mem_2__26_), .Y(w_mem_inst__abc_21378_n6001) );
  AND2X2 AND2X2_5345 ( .A(round_ctr_rst_bF_buf33), .B(\block[474] ), .Y(w_mem_inst__abc_21378_n6002) );
  AND2X2 AND2X2_5346 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf36), .B(w_mem_inst__abc_21378_n6002), .Y(w_mem_inst__abc_21378_n6003) );
  AND2X2 AND2X2_5347 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf44), .B(w_mem_inst_w_mem_1__27_), .Y(w_mem_inst__abc_21378_n6006) );
  AND2X2 AND2X2_5348 ( .A(w_mem_inst__abc_21378_n3152_bF_buf35), .B(w_mem_inst_w_mem_2__27_), .Y(w_mem_inst__abc_21378_n6007) );
  AND2X2 AND2X2_5349 ( .A(round_ctr_rst_bF_buf32), .B(\block[475] ), .Y(w_mem_inst__abc_21378_n6008) );
  AND2X2 AND2X2_535 ( .A(_abc_15724_n1784), .B(_abc_15724_n1788), .Y(_abc_15724_n1790_1) );
  AND2X2 AND2X2_5350 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf35), .B(w_mem_inst__abc_21378_n6008), .Y(w_mem_inst__abc_21378_n6009) );
  AND2X2 AND2X2_5351 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf43), .B(w_mem_inst_w_mem_1__28_), .Y(w_mem_inst__abc_21378_n6012) );
  AND2X2 AND2X2_5352 ( .A(w_mem_inst__abc_21378_n3152_bF_buf34), .B(w_mem_inst_w_mem_2__28_), .Y(w_mem_inst__abc_21378_n6013) );
  AND2X2 AND2X2_5353 ( .A(round_ctr_rst_bF_buf31), .B(\block[476] ), .Y(w_mem_inst__abc_21378_n6014) );
  AND2X2 AND2X2_5354 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf34), .B(w_mem_inst__abc_21378_n6014), .Y(w_mem_inst__abc_21378_n6015) );
  AND2X2 AND2X2_5355 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf42), .B(w_mem_inst_w_mem_1__29_), .Y(w_mem_inst__abc_21378_n6018) );
  AND2X2 AND2X2_5356 ( .A(w_mem_inst__abc_21378_n3152_bF_buf33), .B(w_mem_inst_w_mem_2__29_), .Y(w_mem_inst__abc_21378_n6019) );
  AND2X2 AND2X2_5357 ( .A(round_ctr_rst_bF_buf30), .B(\block[477] ), .Y(w_mem_inst__abc_21378_n6020) );
  AND2X2 AND2X2_5358 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf33), .B(w_mem_inst__abc_21378_n6020), .Y(w_mem_inst__abc_21378_n6021) );
  AND2X2 AND2X2_5359 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf41), .B(w_mem_inst_w_mem_1__30_), .Y(w_mem_inst__abc_21378_n6024) );
  AND2X2 AND2X2_536 ( .A(_abc_15724_n1791), .B(_abc_15724_n1789), .Y(_abc_15724_n1792) );
  AND2X2 AND2X2_5360 ( .A(w_mem_inst__abc_21378_n3152_bF_buf32), .B(w_mem_inst_w_mem_2__30_), .Y(w_mem_inst__abc_21378_n6025) );
  AND2X2 AND2X2_5361 ( .A(round_ctr_rst_bF_buf29), .B(\block[478] ), .Y(w_mem_inst__abc_21378_n6026) );
  AND2X2 AND2X2_5362 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf32), .B(w_mem_inst__abc_21378_n6026), .Y(w_mem_inst__abc_21378_n6027) );
  AND2X2 AND2X2_5363 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf40), .B(w_mem_inst_w_mem_1__31_), .Y(w_mem_inst__abc_21378_n6030) );
  AND2X2 AND2X2_5364 ( .A(w_mem_inst__abc_21378_n3152_bF_buf31), .B(w_mem_inst_w_mem_2__31_), .Y(w_mem_inst__abc_21378_n6031) );
  AND2X2 AND2X2_5365 ( .A(round_ctr_rst_bF_buf28), .B(\block[479] ), .Y(w_mem_inst__abc_21378_n6032) );
  AND2X2 AND2X2_5366 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf31), .B(w_mem_inst__abc_21378_n6032), .Y(w_mem_inst__abc_21378_n6033) );
  AND2X2 AND2X2_5367 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf39), .B(w_mem_inst_w_mem_0__0_), .Y(w_mem_inst__abc_21378_n6036) );
  AND2X2 AND2X2_5368 ( .A(w_mem_inst__abc_21378_n3152_bF_buf30), .B(w_mem_inst_w_mem_1__0_), .Y(w_mem_inst__abc_21378_n6037) );
  AND2X2 AND2X2_5369 ( .A(round_ctr_rst_bF_buf27), .B(\block[480] ), .Y(w_mem_inst__abc_21378_n6038) );
  AND2X2 AND2X2_537 ( .A(_abc_15724_n1792), .B(digest_update_bF_buf10), .Y(_abc_15724_n1793) );
  AND2X2 AND2X2_5370 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf30), .B(w_mem_inst__abc_21378_n6038), .Y(w_mem_inst__abc_21378_n6039) );
  AND2X2 AND2X2_5371 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf38), .B(w_mem_inst_w_mem_0__1_), .Y(w_mem_inst__abc_21378_n6042) );
  AND2X2 AND2X2_5372 ( .A(w_mem_inst__abc_21378_n3152_bF_buf29), .B(w_mem_inst_w_mem_1__1_), .Y(w_mem_inst__abc_21378_n6043) );
  AND2X2 AND2X2_5373 ( .A(round_ctr_rst_bF_buf26), .B(\block[481] ), .Y(w_mem_inst__abc_21378_n6044) );
  AND2X2 AND2X2_5374 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf29), .B(w_mem_inst__abc_21378_n6044), .Y(w_mem_inst__abc_21378_n6045) );
  AND2X2 AND2X2_5375 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf37), .B(w_mem_inst_w_mem_0__2_), .Y(w_mem_inst__abc_21378_n6048) );
  AND2X2 AND2X2_5376 ( .A(w_mem_inst__abc_21378_n3152_bF_buf28), .B(w_mem_inst_w_mem_1__2_), .Y(w_mem_inst__abc_21378_n6049) );
  AND2X2 AND2X2_5377 ( .A(round_ctr_rst_bF_buf25), .B(\block[482] ), .Y(w_mem_inst__abc_21378_n6050) );
  AND2X2 AND2X2_5378 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf28), .B(w_mem_inst__abc_21378_n6050), .Y(w_mem_inst__abc_21378_n6051) );
  AND2X2 AND2X2_5379 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf36), .B(w_mem_inst_w_mem_0__3_), .Y(w_mem_inst__abc_21378_n6054) );
  AND2X2 AND2X2_538 ( .A(_abc_15724_n1791), .B(_abc_15724_n1787), .Y(_abc_15724_n1795_1) );
  AND2X2 AND2X2_5380 ( .A(w_mem_inst__abc_21378_n3152_bF_buf27), .B(w_mem_inst_w_mem_1__3_), .Y(w_mem_inst__abc_21378_n6055) );
  AND2X2 AND2X2_5381 ( .A(round_ctr_rst_bF_buf24), .B(\block[483] ), .Y(w_mem_inst__abc_21378_n6056) );
  AND2X2 AND2X2_5382 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf27), .B(w_mem_inst__abc_21378_n6056), .Y(w_mem_inst__abc_21378_n6057) );
  AND2X2 AND2X2_5383 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf35), .B(w_mem_inst_w_mem_0__4_), .Y(w_mem_inst__abc_21378_n6060) );
  AND2X2 AND2X2_5384 ( .A(w_mem_inst__abc_21378_n3152_bF_buf26), .B(w_mem_inst_w_mem_1__4_), .Y(w_mem_inst__abc_21378_n6061) );
  AND2X2 AND2X2_5385 ( .A(round_ctr_rst_bF_buf23), .B(\block[484] ), .Y(w_mem_inst__abc_21378_n6062) );
  AND2X2 AND2X2_5386 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf26), .B(w_mem_inst__abc_21378_n6062), .Y(w_mem_inst__abc_21378_n6063) );
  AND2X2 AND2X2_5387 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf34), .B(w_mem_inst_w_mem_0__5_), .Y(w_mem_inst__abc_21378_n6066) );
  AND2X2 AND2X2_5388 ( .A(w_mem_inst__abc_21378_n3152_bF_buf25), .B(w_mem_inst_w_mem_1__5_), .Y(w_mem_inst__abc_21378_n6067) );
  AND2X2 AND2X2_5389 ( .A(round_ctr_rst_bF_buf22), .B(\block[485] ), .Y(w_mem_inst__abc_21378_n6068) );
  AND2X2 AND2X2_539 ( .A(_auto_iopadmap_cc_313_execute_26059_83_), .B(c_reg_19_), .Y(_abc_15724_n1798) );
  AND2X2 AND2X2_5390 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf25), .B(w_mem_inst__abc_21378_n6068), .Y(w_mem_inst__abc_21378_n6069) );
  AND2X2 AND2X2_5391 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf33), .B(w_mem_inst_w_mem_0__6_), .Y(w_mem_inst__abc_21378_n6072) );
  AND2X2 AND2X2_5392 ( .A(w_mem_inst__abc_21378_n3152_bF_buf24), .B(w_mem_inst_w_mem_1__6_), .Y(w_mem_inst__abc_21378_n6073) );
  AND2X2 AND2X2_5393 ( .A(round_ctr_rst_bF_buf21), .B(\block[486] ), .Y(w_mem_inst__abc_21378_n6074) );
  AND2X2 AND2X2_5394 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf24), .B(w_mem_inst__abc_21378_n6074), .Y(w_mem_inst__abc_21378_n6075) );
  AND2X2 AND2X2_5395 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf32), .B(w_mem_inst_w_mem_0__7_), .Y(w_mem_inst__abc_21378_n6078) );
  AND2X2 AND2X2_5396 ( .A(w_mem_inst__abc_21378_n3152_bF_buf23), .B(w_mem_inst_w_mem_1__7_), .Y(w_mem_inst__abc_21378_n6079) );
  AND2X2 AND2X2_5397 ( .A(round_ctr_rst_bF_buf20), .B(\block[487] ), .Y(w_mem_inst__abc_21378_n6080) );
  AND2X2 AND2X2_5398 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf23), .B(w_mem_inst__abc_21378_n6080), .Y(w_mem_inst__abc_21378_n6081) );
  AND2X2 AND2X2_5399 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf31), .B(w_mem_inst_w_mem_0__8_), .Y(w_mem_inst__abc_21378_n6084) );
  AND2X2 AND2X2_54 ( .A(_abc_15724_n794), .B(_abc_15724_n792), .Y(_abc_15724_n795) );
  AND2X2 AND2X2_540 ( .A(_abc_15724_n1799_1), .B(_abc_15724_n1797), .Y(_abc_15724_n1800) );
  AND2X2 AND2X2_5400 ( .A(w_mem_inst__abc_21378_n3152_bF_buf22), .B(w_mem_inst_w_mem_1__8_), .Y(w_mem_inst__abc_21378_n6085) );
  AND2X2 AND2X2_5401 ( .A(round_ctr_rst_bF_buf19), .B(\block[488] ), .Y(w_mem_inst__abc_21378_n6086) );
  AND2X2 AND2X2_5402 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf22), .B(w_mem_inst__abc_21378_n6086), .Y(w_mem_inst__abc_21378_n6087) );
  AND2X2 AND2X2_5403 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf30), .B(w_mem_inst_w_mem_0__9_), .Y(w_mem_inst__abc_21378_n6090) );
  AND2X2 AND2X2_5404 ( .A(w_mem_inst__abc_21378_n3152_bF_buf21), .B(w_mem_inst_w_mem_1__9_), .Y(w_mem_inst__abc_21378_n6091) );
  AND2X2 AND2X2_5405 ( .A(round_ctr_rst_bF_buf18), .B(\block[489] ), .Y(w_mem_inst__abc_21378_n6092) );
  AND2X2 AND2X2_5406 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf21), .B(w_mem_inst__abc_21378_n6092), .Y(w_mem_inst__abc_21378_n6093) );
  AND2X2 AND2X2_5407 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf29), .B(w_mem_inst_w_mem_0__10_), .Y(w_mem_inst__abc_21378_n6096) );
  AND2X2 AND2X2_5408 ( .A(w_mem_inst__abc_21378_n3152_bF_buf20), .B(w_mem_inst_w_mem_1__10_), .Y(w_mem_inst__abc_21378_n6097) );
  AND2X2 AND2X2_5409 ( .A(round_ctr_rst_bF_buf17), .B(\block[490] ), .Y(w_mem_inst__abc_21378_n6098) );
  AND2X2 AND2X2_541 ( .A(_abc_15724_n1801), .B(_abc_15724_n1803), .Y(_abc_15724_n1804_1) );
  AND2X2 AND2X2_5410 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf20), .B(w_mem_inst__abc_21378_n6098), .Y(w_mem_inst__abc_21378_n6099) );
  AND2X2 AND2X2_5411 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf28), .B(w_mem_inst_w_mem_0__11_), .Y(w_mem_inst__abc_21378_n6102) );
  AND2X2 AND2X2_5412 ( .A(w_mem_inst__abc_21378_n3152_bF_buf19), .B(w_mem_inst_w_mem_1__11_), .Y(w_mem_inst__abc_21378_n6103) );
  AND2X2 AND2X2_5413 ( .A(round_ctr_rst_bF_buf16), .B(\block[491] ), .Y(w_mem_inst__abc_21378_n6104) );
  AND2X2 AND2X2_5414 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf19), .B(w_mem_inst__abc_21378_n6104), .Y(w_mem_inst__abc_21378_n6105) );
  AND2X2 AND2X2_5415 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf27), .B(w_mem_inst_w_mem_0__12_), .Y(w_mem_inst__abc_21378_n6108) );
  AND2X2 AND2X2_5416 ( .A(w_mem_inst__abc_21378_n3152_bF_buf18), .B(w_mem_inst_w_mem_1__12_), .Y(w_mem_inst__abc_21378_n6109) );
  AND2X2 AND2X2_5417 ( .A(round_ctr_rst_bF_buf15), .B(\block[492] ), .Y(w_mem_inst__abc_21378_n6110) );
  AND2X2 AND2X2_5418 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf18), .B(w_mem_inst__abc_21378_n6110), .Y(w_mem_inst__abc_21378_n6111) );
  AND2X2 AND2X2_5419 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf26), .B(w_mem_inst_w_mem_0__13_), .Y(w_mem_inst__abc_21378_n6114) );
  AND2X2 AND2X2_542 ( .A(_abc_15724_n1804_1), .B(digest_update_bF_buf9), .Y(_abc_15724_n1805) );
  AND2X2 AND2X2_5420 ( .A(w_mem_inst__abc_21378_n3152_bF_buf17), .B(w_mem_inst_w_mem_1__13_), .Y(w_mem_inst__abc_21378_n6115) );
  AND2X2 AND2X2_5421 ( .A(round_ctr_rst_bF_buf14), .B(\block[493] ), .Y(w_mem_inst__abc_21378_n6116) );
  AND2X2 AND2X2_5422 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf17), .B(w_mem_inst__abc_21378_n6116), .Y(w_mem_inst__abc_21378_n6117) );
  AND2X2 AND2X2_5423 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf25), .B(w_mem_inst_w_mem_0__14_), .Y(w_mem_inst__abc_21378_n6120) );
  AND2X2 AND2X2_5424 ( .A(w_mem_inst__abc_21378_n3152_bF_buf16), .B(w_mem_inst_w_mem_1__14_), .Y(w_mem_inst__abc_21378_n6121) );
  AND2X2 AND2X2_5425 ( .A(round_ctr_rst_bF_buf13), .B(\block[494] ), .Y(w_mem_inst__abc_21378_n6122) );
  AND2X2 AND2X2_5426 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf16), .B(w_mem_inst__abc_21378_n6122), .Y(w_mem_inst__abc_21378_n6123) );
  AND2X2 AND2X2_5427 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf24), .B(w_mem_inst_w_mem_0__15_), .Y(w_mem_inst__abc_21378_n6126) );
  AND2X2 AND2X2_5428 ( .A(w_mem_inst__abc_21378_n3152_bF_buf15), .B(w_mem_inst_w_mem_1__15_), .Y(w_mem_inst__abc_21378_n6127) );
  AND2X2 AND2X2_5429 ( .A(round_ctr_rst_bF_buf12), .B(\block[495] ), .Y(w_mem_inst__abc_21378_n6128) );
  AND2X2 AND2X2_543 ( .A(_abc_15724_n1806), .B(_abc_15724_n850_bF_buf8), .Y(_abc_15724_n1807) );
  AND2X2 AND2X2_5430 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf15), .B(w_mem_inst__abc_21378_n6128), .Y(w_mem_inst__abc_21378_n6129) );
  AND2X2 AND2X2_5431 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf23), .B(w_mem_inst_w_mem_0__16_), .Y(w_mem_inst__abc_21378_n6132) );
  AND2X2 AND2X2_5432 ( .A(w_mem_inst__abc_21378_n3152_bF_buf14), .B(w_mem_inst_w_mem_1__16_), .Y(w_mem_inst__abc_21378_n6133) );
  AND2X2 AND2X2_5433 ( .A(round_ctr_rst_bF_buf11), .B(\block[496] ), .Y(w_mem_inst__abc_21378_n6134) );
  AND2X2 AND2X2_5434 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf14), .B(w_mem_inst__abc_21378_n6134), .Y(w_mem_inst__abc_21378_n6135) );
  AND2X2 AND2X2_5435 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf22), .B(w_mem_inst_w_mem_0__17_), .Y(w_mem_inst__abc_21378_n6138) );
  AND2X2 AND2X2_5436 ( .A(w_mem_inst__abc_21378_n3152_bF_buf13), .B(w_mem_inst_w_mem_1__17_), .Y(w_mem_inst__abc_21378_n6139) );
  AND2X2 AND2X2_5437 ( .A(round_ctr_rst_bF_buf10), .B(\block[497] ), .Y(w_mem_inst__abc_21378_n6140) );
  AND2X2 AND2X2_5438 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf13), .B(w_mem_inst__abc_21378_n6140), .Y(w_mem_inst__abc_21378_n6141) );
  AND2X2 AND2X2_5439 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf21), .B(w_mem_inst_w_mem_0__18_), .Y(w_mem_inst__abc_21378_n6144) );
  AND2X2 AND2X2_544 ( .A(_abc_15724_n1788), .B(_abc_15724_n1800), .Y(_abc_15724_n1809_1) );
  AND2X2 AND2X2_5440 ( .A(w_mem_inst__abc_21378_n3152_bF_buf12), .B(w_mem_inst_w_mem_1__18_), .Y(w_mem_inst__abc_21378_n6145) );
  AND2X2 AND2X2_5441 ( .A(round_ctr_rst_bF_buf9), .B(\block[498] ), .Y(w_mem_inst__abc_21378_n6146) );
  AND2X2 AND2X2_5442 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf12), .B(w_mem_inst__abc_21378_n6146), .Y(w_mem_inst__abc_21378_n6147) );
  AND2X2 AND2X2_5443 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf20), .B(w_mem_inst_w_mem_0__19_), .Y(w_mem_inst__abc_21378_n6150) );
  AND2X2 AND2X2_5444 ( .A(w_mem_inst__abc_21378_n3152_bF_buf11), .B(w_mem_inst_w_mem_1__19_), .Y(w_mem_inst__abc_21378_n6151) );
  AND2X2 AND2X2_5445 ( .A(round_ctr_rst_bF_buf8), .B(\block[499] ), .Y(w_mem_inst__abc_21378_n6152) );
  AND2X2 AND2X2_5446 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf11), .B(w_mem_inst__abc_21378_n6152), .Y(w_mem_inst__abc_21378_n6153) );
  AND2X2 AND2X2_5447 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf19), .B(w_mem_inst_w_mem_0__20_), .Y(w_mem_inst__abc_21378_n6156) );
  AND2X2 AND2X2_5448 ( .A(w_mem_inst__abc_21378_n3152_bF_buf10), .B(w_mem_inst_w_mem_1__20_), .Y(w_mem_inst__abc_21378_n6157) );
  AND2X2 AND2X2_5449 ( .A(round_ctr_rst_bF_buf7), .B(\block[500] ), .Y(w_mem_inst__abc_21378_n6158) );
  AND2X2 AND2X2_545 ( .A(_abc_15724_n1782), .B(_abc_15724_n1809_1), .Y(_abc_15724_n1810) );
  AND2X2 AND2X2_5450 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf10), .B(w_mem_inst__abc_21378_n6158), .Y(w_mem_inst__abc_21378_n6159) );
  AND2X2 AND2X2_5451 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf18), .B(w_mem_inst_w_mem_0__21_), .Y(w_mem_inst__abc_21378_n6162) );
  AND2X2 AND2X2_5452 ( .A(w_mem_inst__abc_21378_n3152_bF_buf9), .B(w_mem_inst_w_mem_1__21_), .Y(w_mem_inst__abc_21378_n6163) );
  AND2X2 AND2X2_5453 ( .A(round_ctr_rst_bF_buf6), .B(\block[501] ), .Y(w_mem_inst__abc_21378_n6164) );
  AND2X2 AND2X2_5454 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf9), .B(w_mem_inst__abc_21378_n6164), .Y(w_mem_inst__abc_21378_n6165) );
  AND2X2 AND2X2_5455 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf17), .B(w_mem_inst_w_mem_0__22_), .Y(w_mem_inst__abc_21378_n6168) );
  AND2X2 AND2X2_5456 ( .A(w_mem_inst__abc_21378_n3152_bF_buf8), .B(w_mem_inst_w_mem_1__22_), .Y(w_mem_inst__abc_21378_n6169) );
  AND2X2 AND2X2_5457 ( .A(round_ctr_rst_bF_buf5), .B(\block[502] ), .Y(w_mem_inst__abc_21378_n6170) );
  AND2X2 AND2X2_5458 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf8), .B(w_mem_inst__abc_21378_n6170), .Y(w_mem_inst__abc_21378_n6171) );
  AND2X2 AND2X2_5459 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf16), .B(w_mem_inst_w_mem_0__23_), .Y(w_mem_inst__abc_21378_n6174) );
  AND2X2 AND2X2_546 ( .A(_abc_15724_n1781_1), .B(_abc_15724_n1809_1), .Y(_abc_15724_n1813_1) );
  AND2X2 AND2X2_5460 ( .A(w_mem_inst__abc_21378_n3152_bF_buf7), .B(w_mem_inst_w_mem_1__23_), .Y(w_mem_inst__abc_21378_n6175) );
  AND2X2 AND2X2_5461 ( .A(round_ctr_rst_bF_buf4), .B(\block[503] ), .Y(w_mem_inst__abc_21378_n6176) );
  AND2X2 AND2X2_5462 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf7), .B(w_mem_inst__abc_21378_n6176), .Y(w_mem_inst__abc_21378_n6177) );
  AND2X2 AND2X2_5463 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf15), .B(w_mem_inst_w_mem_0__24_), .Y(w_mem_inst__abc_21378_n6180) );
  AND2X2 AND2X2_5464 ( .A(w_mem_inst__abc_21378_n3152_bF_buf6), .B(w_mem_inst_w_mem_1__24_), .Y(w_mem_inst__abc_21378_n6181) );
  AND2X2 AND2X2_5465 ( .A(round_ctr_rst_bF_buf3), .B(\block[504] ), .Y(w_mem_inst__abc_21378_n6182) );
  AND2X2 AND2X2_5466 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf6), .B(w_mem_inst__abc_21378_n6182), .Y(w_mem_inst__abc_21378_n6183) );
  AND2X2 AND2X2_5467 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf14), .B(w_mem_inst_w_mem_0__25_), .Y(w_mem_inst__abc_21378_n6186) );
  AND2X2 AND2X2_5468 ( .A(w_mem_inst__abc_21378_n3152_bF_buf5), .B(w_mem_inst_w_mem_1__25_), .Y(w_mem_inst__abc_21378_n6187) );
  AND2X2 AND2X2_5469 ( .A(round_ctr_rst_bF_buf2), .B(\block[505] ), .Y(w_mem_inst__abc_21378_n6188) );
  AND2X2 AND2X2_547 ( .A(_abc_15724_n1797), .B(_abc_15724_n1786_1), .Y(_abc_15724_n1814) );
  AND2X2 AND2X2_5470 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf5), .B(w_mem_inst__abc_21378_n6188), .Y(w_mem_inst__abc_21378_n6189) );
  AND2X2 AND2X2_5471 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf13), .B(w_mem_inst_w_mem_0__26_), .Y(w_mem_inst__abc_21378_n6192) );
  AND2X2 AND2X2_5472 ( .A(w_mem_inst__abc_21378_n3152_bF_buf4), .B(w_mem_inst_w_mem_1__26_), .Y(w_mem_inst__abc_21378_n6193) );
  AND2X2 AND2X2_5473 ( .A(round_ctr_rst_bF_buf1), .B(\block[506] ), .Y(w_mem_inst__abc_21378_n6194) );
  AND2X2 AND2X2_5474 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf4), .B(w_mem_inst__abc_21378_n6194), .Y(w_mem_inst__abc_21378_n6195) );
  AND2X2 AND2X2_5475 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf12), .B(w_mem_inst_w_mem_0__27_), .Y(w_mem_inst__abc_21378_n6198) );
  AND2X2 AND2X2_5476 ( .A(w_mem_inst__abc_21378_n3152_bF_buf3), .B(w_mem_inst_w_mem_1__27_), .Y(w_mem_inst__abc_21378_n6199) );
  AND2X2 AND2X2_5477 ( .A(round_ctr_rst_bF_buf0), .B(\block[507] ), .Y(w_mem_inst__abc_21378_n6200) );
  AND2X2 AND2X2_5478 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf3), .B(w_mem_inst__abc_21378_n6200), .Y(w_mem_inst__abc_21378_n6201) );
  AND2X2 AND2X2_5479 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf11), .B(w_mem_inst_w_mem_0__28_), .Y(w_mem_inst__abc_21378_n6204) );
  AND2X2 AND2X2_548 ( .A(_abc_15724_n1812), .B(_abc_15724_n1817), .Y(_abc_15724_n1818_1) );
  AND2X2 AND2X2_5480 ( .A(w_mem_inst__abc_21378_n3152_bF_buf2), .B(w_mem_inst_w_mem_1__28_), .Y(w_mem_inst__abc_21378_n6205) );
  AND2X2 AND2X2_5481 ( .A(round_ctr_rst_bF_buf63), .B(\block[508] ), .Y(w_mem_inst__abc_21378_n6206) );
  AND2X2 AND2X2_5482 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf2), .B(w_mem_inst__abc_21378_n6206), .Y(w_mem_inst__abc_21378_n6207) );
  AND2X2 AND2X2_5483 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf10), .B(w_mem_inst_w_mem_0__29_), .Y(w_mem_inst__abc_21378_n6210) );
  AND2X2 AND2X2_5484 ( .A(w_mem_inst__abc_21378_n3152_bF_buf1), .B(w_mem_inst_w_mem_1__29_), .Y(w_mem_inst__abc_21378_n6211) );
  AND2X2 AND2X2_5485 ( .A(round_ctr_rst_bF_buf62), .B(\block[509] ), .Y(w_mem_inst__abc_21378_n6212) );
  AND2X2 AND2X2_5486 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf1), .B(w_mem_inst__abc_21378_n6212), .Y(w_mem_inst__abc_21378_n6213) );
  AND2X2 AND2X2_5487 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf9), .B(w_mem_inst_w_mem_0__30_), .Y(w_mem_inst__abc_21378_n6216) );
  AND2X2 AND2X2_5488 ( .A(w_mem_inst__abc_21378_n3152_bF_buf0), .B(w_mem_inst_w_mem_1__30_), .Y(w_mem_inst__abc_21378_n6217) );
  AND2X2 AND2X2_5489 ( .A(round_ctr_rst_bF_buf61), .B(\block[510] ), .Y(w_mem_inst__abc_21378_n6218) );
  AND2X2 AND2X2_549 ( .A(_auto_iopadmap_cc_313_execute_26059_84_), .B(c_reg_20_), .Y(_abc_15724_n1821) );
  AND2X2 AND2X2_5490 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf0), .B(w_mem_inst__abc_21378_n6218), .Y(w_mem_inst__abc_21378_n6219) );
  AND2X2 AND2X2_5491 ( .A(w_mem_inst__abc_21378_n3347_1_bF_buf8), .B(w_mem_inst_w_mem_0__31_), .Y(w_mem_inst__abc_21378_n6222) );
  AND2X2 AND2X2_5492 ( .A(w_mem_inst__abc_21378_n3152_bF_buf63), .B(w_mem_inst_w_mem_1__31_), .Y(w_mem_inst__abc_21378_n6223) );
  AND2X2 AND2X2_5493 ( .A(round_ctr_rst_bF_buf60), .B(\block[511] ), .Y(w_mem_inst__abc_21378_n6224) );
  AND2X2 AND2X2_5494 ( .A(w_mem_inst__abc_21378_n3154_1_bF_buf63), .B(w_mem_inst__abc_21378_n6224), .Y(w_mem_inst__abc_21378_n6225) );
  AND2X2 AND2X2_5495 ( .A(w_mem_inst__abc_21378_n6229), .B(w_mem_inst__abc_21378_n3156_bF_buf1), .Y(w_mem_inst__abc_21378_n6230) );
  AND2X2 AND2X2_5496 ( .A(w_mem_inst__abc_21378_n6231), .B(w_mem_inst__abc_21378_n6228), .Y(w_mem_inst_w_ctr_reg_0__FF_INPUT) );
  AND2X2 AND2X2_5497 ( .A(w_mem_inst__abc_21378_n6230), .B(w_mem_inst_w_ctr_reg_1_), .Y(w_mem_inst__abc_21378_n6233) );
  AND2X2 AND2X2_5498 ( .A(w_mem_inst__abc_21378_n6234), .B(round_ctr_inc_bF_buf9), .Y(w_mem_inst__abc_21378_n6235) );
  AND2X2 AND2X2_5499 ( .A(w_mem_inst__abc_21378_n6237), .B(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_21378_n6238) );
  AND2X2 AND2X2_55 ( .A(_abc_15724_n796), .B(_abc_15724_n791_1), .Y(_abc_15724_n797) );
  AND2X2 AND2X2_550 ( .A(_abc_15724_n1822), .B(_abc_15724_n1820), .Y(_abc_15724_n1823_1) );
  AND2X2 AND2X2_5500 ( .A(w_mem_inst__abc_21378_n1603_1), .B(round_ctr_inc_bF_buf7), .Y(w_mem_inst__abc_21378_n6239) );
  AND2X2 AND2X2_5501 ( .A(w_mem_inst__abc_21378_n1603_1), .B(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_21378_n6241) );
  AND2X2 AND2X2_5502 ( .A(w_mem_inst__abc_21378_n6241), .B(round_ctr_inc_bF_buf6), .Y(w_mem_inst__abc_21378_n6242) );
  AND2X2 AND2X2_5503 ( .A(w_mem_inst__abc_21378_n6240), .B(w_mem_inst__abc_21378_n6243), .Y(w_mem_inst_w_ctr_reg_2__FF_INPUT) );
  AND2X2 AND2X2_5504 ( .A(w_mem_inst__abc_21378_n6237), .B(w_mem_inst_w_ctr_reg_3_), .Y(w_mem_inst__abc_21378_n6245) );
  AND2X2 AND2X2_5505 ( .A(w_mem_inst__abc_21378_n1605_bF_buf2), .B(round_ctr_inc_bF_buf5), .Y(w_mem_inst__abc_21378_n6247) );
  AND2X2 AND2X2_5506 ( .A(w_mem_inst__abc_21378_n6246), .B(w_mem_inst__abc_21378_n6248), .Y(w_mem_inst_w_ctr_reg_3__FF_INPUT) );
  AND2X2 AND2X2_5507 ( .A(w_mem_inst__abc_21378_n6237), .B(w_mem_inst_w_ctr_reg_4_), .Y(w_mem_inst__abc_21378_n6250) );
  AND2X2 AND2X2_5508 ( .A(w_mem_inst__abc_21378_n6247), .B(w_mem_inst_w_ctr_reg_4_), .Y(w_mem_inst__abc_21378_n6252) );
  AND2X2 AND2X2_5509 ( .A(w_mem_inst__abc_21378_n6253), .B(w_mem_inst__abc_21378_n6251), .Y(w_mem_inst_w_ctr_reg_4__FF_INPUT) );
  AND2X2 AND2X2_551 ( .A(_abc_15724_n1819), .B(_abc_15724_n1823_1), .Y(_abc_15724_n1825) );
  AND2X2 AND2X2_5510 ( .A(w_mem_inst__abc_21378_n6237), .B(w_mem_inst_w_ctr_reg_5_), .Y(w_mem_inst__abc_21378_n6255) );
  AND2X2 AND2X2_5511 ( .A(w_mem_inst__abc_21378_n6252), .B(w_mem_inst_w_ctr_reg_5_), .Y(w_mem_inst__abc_21378_n6257) );
  AND2X2 AND2X2_5512 ( .A(w_mem_inst__abc_21378_n6258), .B(w_mem_inst__abc_21378_n6256), .Y(w_mem_inst_w_ctr_reg_5__FF_INPUT) );
  AND2X2 AND2X2_5513 ( .A(w_mem_inst__abc_21378_n6237), .B(w_mem_inst_w_ctr_reg_6_), .Y(w_mem_inst__abc_21378_n6260) );
  AND2X2 AND2X2_5514 ( .A(w_mem_inst__abc_21378_n6257), .B(w_mem_inst_w_ctr_reg_6_), .Y(w_mem_inst__abc_21378_n6262) );
  AND2X2 AND2X2_5515 ( .A(w_mem_inst__abc_21378_n6263), .B(w_mem_inst__abc_21378_n6261), .Y(w_mem_inst_w_ctr_reg_6__FF_INPUT) );
  AND2X2 AND2X2_552 ( .A(_abc_15724_n1826), .B(_abc_15724_n1824), .Y(_abc_15724_n1827_1) );
  AND2X2 AND2X2_553 ( .A(_abc_15724_n1827_1), .B(digest_update_bF_buf8), .Y(_abc_15724_n1828) );
  AND2X2 AND2X2_554 ( .A(_abc_15724_n1829), .B(_abc_15724_n850_bF_buf7), .Y(_abc_15724_n1830) );
  AND2X2 AND2X2_555 ( .A(_abc_15724_n1826), .B(_abc_15724_n1822), .Y(_abc_15724_n1832) );
  AND2X2 AND2X2_556 ( .A(_auto_iopadmap_cc_313_execute_26059_85_), .B(c_reg_21_), .Y(_abc_15724_n1835) );
  AND2X2 AND2X2_557 ( .A(_abc_15724_n1836_1), .B(_abc_15724_n1834), .Y(_abc_15724_n1837) );
  AND2X2 AND2X2_558 ( .A(_abc_15724_n1838), .B(_abc_15724_n1840), .Y(_abc_15724_n1841_1) );
  AND2X2 AND2X2_559 ( .A(_abc_15724_n1841_1), .B(digest_update_bF_buf7), .Y(_abc_15724_n1842) );
  AND2X2 AND2X2_56 ( .A(_abc_15724_n799), .B(_abc_15724_n800), .Y(_abc_15724_n801) );
  AND2X2 AND2X2_560 ( .A(_abc_15724_n1843), .B(_abc_15724_n850_bF_buf6), .Y(_abc_15724_n1844) );
  AND2X2 AND2X2_561 ( .A(_abc_15724_n907_1_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_86_), .Y(_abc_15724_n1846_1) );
  AND2X2 AND2X2_562 ( .A(_abc_15724_n1847), .B(_abc_15724_n1836_1), .Y(_abc_15724_n1848) );
  AND2X2 AND2X2_563 ( .A(_abc_15724_n1823_1), .B(_abc_15724_n1837), .Y(_abc_15724_n1850) );
  AND2X2 AND2X2_564 ( .A(_abc_15724_n1819), .B(_abc_15724_n1850), .Y(_abc_15724_n1851_1) );
  AND2X2 AND2X2_565 ( .A(_auto_iopadmap_cc_313_execute_26059_86_), .B(c_reg_22_), .Y(_abc_15724_n1854) );
  AND2X2 AND2X2_566 ( .A(_abc_15724_n1855), .B(_abc_15724_n1853), .Y(_abc_15724_n1856_1) );
  AND2X2 AND2X2_567 ( .A(_abc_15724_n1852), .B(_abc_15724_n1856_1), .Y(_abc_15724_n1857) );
  AND2X2 AND2X2_568 ( .A(_abc_15724_n1859), .B(digest_update_bF_buf6), .Y(_abc_15724_n1860) );
  AND2X2 AND2X2_569 ( .A(_abc_15724_n1860), .B(_abc_15724_n1858), .Y(_abc_15724_n1861_1) );
  AND2X2 AND2X2_57 ( .A(_abc_15724_n798), .B(_abc_15724_n801), .Y(_abc_15724_n802) );
  AND2X2 AND2X2_570 ( .A(_abc_15724_n1858), .B(_abc_15724_n1855), .Y(_abc_15724_n1863) );
  AND2X2 AND2X2_571 ( .A(_auto_iopadmap_cc_313_execute_26059_87_), .B(c_reg_23_), .Y(_abc_15724_n1866) );
  AND2X2 AND2X2_572 ( .A(_abc_15724_n1867), .B(_abc_15724_n1865_1), .Y(_abc_15724_n1868) );
  AND2X2 AND2X2_573 ( .A(_abc_15724_n1869), .B(_abc_15724_n1871), .Y(_abc_15724_n1872) );
  AND2X2 AND2X2_574 ( .A(_abc_15724_n1872), .B(digest_update_bF_buf5), .Y(_abc_15724_n1873) );
  AND2X2 AND2X2_575 ( .A(_abc_15724_n1874), .B(_abc_15724_n850_bF_buf5), .Y(_abc_15724_n1875_1) );
  AND2X2 AND2X2_576 ( .A(_abc_15724_n907_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_88_), .Y(_abc_15724_n1877) );
  AND2X2 AND2X2_577 ( .A(_abc_15724_n1856_1), .B(_abc_15724_n1868), .Y(_abc_15724_n1878) );
  AND2X2 AND2X2_578 ( .A(_abc_15724_n1849), .B(_abc_15724_n1878), .Y(_abc_15724_n1879) );
  AND2X2 AND2X2_579 ( .A(_abc_15724_n1865_1), .B(_abc_15724_n1854), .Y(_abc_15724_n1880_1) );
  AND2X2 AND2X2_58 ( .A(_abc_15724_n803_1), .B(_abc_15724_n788), .Y(_abc_15724_n804_1) );
  AND2X2 AND2X2_580 ( .A(_abc_15724_n1850), .B(_abc_15724_n1878), .Y(_abc_15724_n1884) );
  AND2X2 AND2X2_581 ( .A(_abc_15724_n1886), .B(_abc_15724_n1883), .Y(_abc_15724_n1887) );
  AND2X2 AND2X2_582 ( .A(_auto_iopadmap_cc_313_execute_26059_88_), .B(c_reg_24_), .Y(_abc_15724_n1890) );
  AND2X2 AND2X2_583 ( .A(_abc_15724_n1891), .B(_abc_15724_n1889_1), .Y(_abc_15724_n1892) );
  AND2X2 AND2X2_584 ( .A(_abc_15724_n1888), .B(_abc_15724_n1892), .Y(_abc_15724_n1894) );
  AND2X2 AND2X2_585 ( .A(_abc_15724_n1895), .B(_abc_15724_n1893_1), .Y(_abc_15724_n1896) );
  AND2X2 AND2X2_586 ( .A(_abc_15724_n1896), .B(digest_update_bF_buf4), .Y(_abc_15724_n1897_1) );
  AND2X2 AND2X2_587 ( .A(_abc_15724_n907_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_89_), .Y(_abc_15724_n1899) );
  AND2X2 AND2X2_588 ( .A(_auto_iopadmap_cc_313_execute_26059_89_), .B(c_reg_25_), .Y(_abc_15724_n1901_1) );
  AND2X2 AND2X2_589 ( .A(_abc_15724_n1902), .B(_abc_15724_n1900), .Y(_abc_15724_n1903) );
  AND2X2 AND2X2_59 ( .A(_abc_15724_n806_1), .B(_abc_15724_n807), .Y(_abc_15724_n808) );
  AND2X2 AND2X2_590 ( .A(_abc_15724_n1892), .B(_abc_15724_n1903), .Y(_abc_15724_n1906) );
  AND2X2 AND2X2_591 ( .A(_abc_15724_n1888), .B(_abc_15724_n1906), .Y(_abc_15724_n1907) );
  AND2X2 AND2X2_592 ( .A(_abc_15724_n1903), .B(_abc_15724_n1890), .Y(_abc_15724_n1909_1) );
  AND2X2 AND2X2_593 ( .A(_abc_15724_n1910), .B(digest_update_bF_buf3), .Y(_abc_15724_n1911) );
  AND2X2 AND2X2_594 ( .A(_abc_15724_n1908), .B(_abc_15724_n1911), .Y(_abc_15724_n1912) );
  AND2X2 AND2X2_595 ( .A(_abc_15724_n1912), .B(_abc_15724_n1905_1), .Y(_abc_15724_n1913_1) );
  AND2X2 AND2X2_596 ( .A(_abc_15724_n907_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_90_), .Y(_abc_15724_n1915) );
  AND2X2 AND2X2_597 ( .A(_abc_15724_n1910), .B(_abc_15724_n1902), .Y(_abc_15724_n1916) );
  AND2X2 AND2X2_598 ( .A(_abc_15724_n1908), .B(_abc_15724_n1916), .Y(_abc_15724_n1917) );
  AND2X2 AND2X2_599 ( .A(_auto_iopadmap_cc_313_execute_26059_90_), .B(c_reg_26_), .Y(_abc_15724_n1920) );
  AND2X2 AND2X2_6 ( .A(_abc_15724_n706), .B(_abc_15724_n707), .Y(_abc_15724_n708_1) );
  AND2X2 AND2X2_60 ( .A(_abc_15724_n805), .B(_abc_15724_n808), .Y(_abc_15724_n809) );
  AND2X2 AND2X2_600 ( .A(_abc_15724_n1921), .B(_abc_15724_n1919), .Y(_abc_15724_n1922) );
  AND2X2 AND2X2_601 ( .A(_abc_15724_n1918_1), .B(_abc_15724_n1922), .Y(_abc_15724_n1924) );
  AND2X2 AND2X2_602 ( .A(_abc_15724_n1925), .B(_abc_15724_n1923_1), .Y(_abc_15724_n1926) );
  AND2X2 AND2X2_603 ( .A(_abc_15724_n1926), .B(digest_update_bF_buf2), .Y(_abc_15724_n1927_1) );
  AND2X2 AND2X2_604 ( .A(_auto_iopadmap_cc_313_execute_26059_91_), .B(c_reg_27_), .Y(_abc_15724_n1931_1) );
  AND2X2 AND2X2_605 ( .A(_abc_15724_n1932), .B(_abc_15724_n1930), .Y(_abc_15724_n1933) );
  AND2X2 AND2X2_606 ( .A(_abc_15724_n1937), .B(_abc_15724_n1934), .Y(_abc_15724_n1938) );
  AND2X2 AND2X2_607 ( .A(_abc_15724_n1938), .B(digest_update_bF_buf1), .Y(_abc_15724_n1939) );
  AND2X2 AND2X2_608 ( .A(_abc_15724_n1940_1), .B(_abc_15724_n850_bF_buf4), .Y(_abc_15724_n1941) );
  AND2X2 AND2X2_609 ( .A(_abc_15724_n1930), .B(_abc_15724_n1920), .Y(_abc_15724_n1943) );
  AND2X2 AND2X2_61 ( .A(_abc_15724_n810), .B(_abc_15724_n785), .Y(_abc_15724_n811) );
  AND2X2 AND2X2_610 ( .A(_abc_15724_n1922), .B(_abc_15724_n1933), .Y(_abc_15724_n1946) );
  AND2X2 AND2X2_611 ( .A(_abc_15724_n1948_1), .B(_abc_15724_n1945), .Y(_abc_15724_n1949) );
  AND2X2 AND2X2_612 ( .A(_abc_15724_n1906), .B(_abc_15724_n1946), .Y(_abc_15724_n1950) );
  AND2X2 AND2X2_613 ( .A(_abc_15724_n1952), .B(_abc_15724_n1949), .Y(_abc_15724_n1953_1) );
  AND2X2 AND2X2_614 ( .A(_auto_iopadmap_cc_313_execute_26059_92_), .B(c_reg_28_), .Y(_abc_15724_n1956) );
  AND2X2 AND2X2_615 ( .A(_abc_15724_n1957_1), .B(_abc_15724_n1955), .Y(_abc_15724_n1958) );
  AND2X2 AND2X2_616 ( .A(_abc_15724_n1954), .B(_abc_15724_n1958), .Y(_abc_15724_n1960) );
  AND2X2 AND2X2_617 ( .A(_abc_15724_n1961), .B(_abc_15724_n1959), .Y(_abc_15724_n1962_1) );
  AND2X2 AND2X2_618 ( .A(_abc_15724_n1962_1), .B(digest_update_bF_buf0), .Y(_abc_15724_n1963) );
  AND2X2 AND2X2_619 ( .A(_abc_15724_n1964), .B(_abc_15724_n850_bF_buf3), .Y(_abc_15724_n1965) );
  AND2X2 AND2X2_62 ( .A(_abc_15724_n812_1), .B(_abc_15724_n783), .Y(_abc_15724_n813_1) );
  AND2X2 AND2X2_620 ( .A(_abc_15724_n907_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_93_), .Y(_abc_15724_n1967) );
  AND2X2 AND2X2_621 ( .A(_abc_15724_n1961), .B(_abc_15724_n1957_1), .Y(_abc_15724_n1968) );
  AND2X2 AND2X2_622 ( .A(_auto_iopadmap_cc_313_execute_26059_93_), .B(c_reg_29_), .Y(_abc_15724_n1970_1) );
  AND2X2 AND2X2_623 ( .A(_abc_15724_n1971), .B(_abc_15724_n1969), .Y(_abc_15724_n1972) );
  AND2X2 AND2X2_624 ( .A(_abc_15724_n1976), .B(_abc_15724_n1974_1), .Y(_abc_15724_n1977) );
  AND2X2 AND2X2_625 ( .A(_abc_15724_n1977), .B(digest_update_bF_buf11), .Y(_abc_15724_n1978) );
  AND2X2 AND2X2_626 ( .A(_abc_15724_n907_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_94_), .Y(_abc_15724_n1980) );
  AND2X2 AND2X2_627 ( .A(_auto_iopadmap_cc_313_execute_26059_94_), .B(c_reg_30_), .Y(_abc_15724_n1981) );
  AND2X2 AND2X2_628 ( .A(_abc_15724_n1982), .B(_abc_15724_n1983_1), .Y(_abc_15724_n1984) );
  AND2X2 AND2X2_629 ( .A(_abc_15724_n1972), .B(_abc_15724_n1956), .Y(_abc_15724_n1986) );
  AND2X2 AND2X2_63 ( .A(_abc_15724_n815_1), .B(_abc_15724_n767_1), .Y(_abc_15724_n816) );
  AND2X2 AND2X2_630 ( .A(_abc_15724_n1958), .B(_abc_15724_n1972), .Y(_abc_15724_n1989) );
  AND2X2 AND2X2_631 ( .A(_abc_15724_n1991), .B(_abc_15724_n1988_1), .Y(_abc_15724_n1992) );
  AND2X2 AND2X2_632 ( .A(_abc_15724_n1995), .B(digest_update_bF_buf10), .Y(_abc_15724_n1996) );
  AND2X2 AND2X2_633 ( .A(_abc_15724_n1996), .B(_abc_15724_n1993_1), .Y(_abc_15724_n1997) );
  AND2X2 AND2X2_634 ( .A(_abc_15724_n1993_1), .B(_abc_15724_n1982), .Y(_abc_15724_n1999) );
  AND2X2 AND2X2_635 ( .A(_abc_15724_n2002_1), .B(_abc_15724_n2004), .Y(_abc_15724_n2005) );
  AND2X2 AND2X2_636 ( .A(_abc_15724_n2007), .B(_abc_15724_n2008), .Y(_abc_15724_n2009) );
  AND2X2 AND2X2_637 ( .A(_abc_15724_n2009), .B(digest_update_bF_buf9), .Y(_abc_15724_n2010) );
  AND2X2 AND2X2_638 ( .A(_abc_15724_n2011_1), .B(_abc_15724_n850_bF_buf2), .Y(_abc_15724_n2012) );
  AND2X2 AND2X2_639 ( .A(_auto_iopadmap_cc_313_execute_26059_96_), .B(b_reg_0_), .Y(_abc_15724_n2015) );
  AND2X2 AND2X2_64 ( .A(_abc_15724_n817), .B(_abc_15724_n818), .Y(_abc_15724_n819) );
  AND2X2 AND2X2_640 ( .A(_abc_15724_n2016_1), .B(digest_update_bF_buf8), .Y(_abc_15724_n2017) );
  AND2X2 AND2X2_641 ( .A(_abc_15724_n2017), .B(_abc_15724_n2014), .Y(_abc_15724_n2018) );
  AND2X2 AND2X2_642 ( .A(_abc_15724_n2019), .B(_abc_15724_n850_bF_buf1), .Y(_abc_15724_n2020_1) );
  AND2X2 AND2X2_643 ( .A(_auto_iopadmap_cc_313_execute_26059_97_), .B(b_reg_1_), .Y(_abc_15724_n2023) );
  AND2X2 AND2X2_644 ( .A(_abc_15724_n2024_1), .B(_abc_15724_n2022), .Y(_abc_15724_n2025) );
  AND2X2 AND2X2_645 ( .A(_abc_15724_n2025), .B(_abc_15724_n2015), .Y(_abc_15724_n2027) );
  AND2X2 AND2X2_646 ( .A(_abc_15724_n2028), .B(_abc_15724_n2026), .Y(_abc_15724_n2029_1) );
  AND2X2 AND2X2_647 ( .A(_abc_15724_n2029_1), .B(digest_update_bF_buf7), .Y(_abc_15724_n2030) );
  AND2X2 AND2X2_648 ( .A(_abc_15724_n907_1_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_97_), .Y(_abc_15724_n2031) );
  AND2X2 AND2X2_649 ( .A(_abc_15724_n2028), .B(_abc_15724_n2024_1), .Y(_abc_15724_n2033) );
  AND2X2 AND2X2_65 ( .A(_abc_15724_n816), .B(_abc_15724_n819), .Y(_abc_15724_n820) );
  AND2X2 AND2X2_650 ( .A(_auto_iopadmap_cc_313_execute_26059_98_), .B(b_reg_2_), .Y(_abc_15724_n2036) );
  AND2X2 AND2X2_651 ( .A(_abc_15724_n2037), .B(_abc_15724_n2035), .Y(_abc_15724_n2038_1) );
  AND2X2 AND2X2_652 ( .A(_abc_15724_n2034_1), .B(_abc_15724_n2038_1), .Y(_abc_15724_n2039) );
  AND2X2 AND2X2_653 ( .A(_abc_15724_n2040), .B(_abc_15724_n2041), .Y(_abc_15724_n2042) );
  AND2X2 AND2X2_654 ( .A(_abc_15724_n2042), .B(digest_update_bF_buf6), .Y(_abc_15724_n2043_1) );
  AND2X2 AND2X2_655 ( .A(_abc_15724_n907_1_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_98_), .Y(_abc_15724_n2044) );
  AND2X2 AND2X2_656 ( .A(_auto_iopadmap_cc_313_execute_26059_99_), .B(b_reg_3_), .Y(_abc_15724_n2048_1) );
  AND2X2 AND2X2_657 ( .A(_abc_15724_n2049), .B(_abc_15724_n2047), .Y(_abc_15724_n2050) );
  AND2X2 AND2X2_658 ( .A(_abc_15724_n2054), .B(_abc_15724_n2051), .Y(_abc_15724_n2055) );
  AND2X2 AND2X2_659 ( .A(_abc_15724_n2055), .B(digest_update_bF_buf5), .Y(_abc_15724_n2056) );
  AND2X2 AND2X2_66 ( .A(_abc_15724_n765), .B(_abc_15724_n820), .Y(_abc_15724_n821) );
  AND2X2 AND2X2_660 ( .A(_abc_15724_n2057_1), .B(_abc_15724_n850_bF_buf0), .Y(_abc_15724_n2058) );
  AND2X2 AND2X2_661 ( .A(_auto_iopadmap_cc_313_execute_26059_100_), .B(b_reg_4_), .Y(_abc_15724_n2061_1) );
  AND2X2 AND2X2_662 ( .A(_abc_15724_n2062), .B(_abc_15724_n2060), .Y(_abc_15724_n2063) );
  AND2X2 AND2X2_663 ( .A(_abc_15724_n2046), .B(_abc_15724_n2047), .Y(_abc_15724_n2064) );
  AND2X2 AND2X2_664 ( .A(_abc_15724_n2065_1), .B(_abc_15724_n2063), .Y(_abc_15724_n2066) );
  AND2X2 AND2X2_665 ( .A(_abc_15724_n2067), .B(_abc_15724_n2068), .Y(_abc_15724_n2069) );
  AND2X2 AND2X2_666 ( .A(_abc_15724_n2069), .B(digest_update_bF_buf4), .Y(_abc_15724_n2070_1) );
  AND2X2 AND2X2_667 ( .A(_abc_15724_n907_1_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_100_), .Y(_abc_15724_n2071) );
  AND2X2 AND2X2_668 ( .A(_abc_15724_n907_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_101_), .Y(_abc_15724_n2073) );
  AND2X2 AND2X2_669 ( .A(_auto_iopadmap_cc_313_execute_26059_101_), .B(b_reg_5_), .Y(_abc_15724_n2076) );
  AND2X2 AND2X2_67 ( .A(_abc_15724_n814), .B(_abc_15724_n821), .Y(_abc_15724_n822) );
  AND2X2 AND2X2_670 ( .A(_abc_15724_n2077), .B(_abc_15724_n2075), .Y(_abc_15724_n2078) );
  AND2X2 AND2X2_671 ( .A(_abc_15724_n2074_1), .B(_abc_15724_n2078), .Y(_abc_15724_n2079_1) );
  AND2X2 AND2X2_672 ( .A(_abc_15724_n2081), .B(digest_update_bF_buf3), .Y(_abc_15724_n2082) );
  AND2X2 AND2X2_673 ( .A(_abc_15724_n2082), .B(_abc_15724_n2080), .Y(_abc_15724_n2083_1) );
  AND2X2 AND2X2_674 ( .A(_abc_15724_n907_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_102_), .Y(_abc_15724_n2085) );
  AND2X2 AND2X2_675 ( .A(_auto_iopadmap_cc_313_execute_26059_102_), .B(b_reg_6_), .Y(_abc_15724_n2088_1) );
  AND2X2 AND2X2_676 ( .A(_abc_15724_n2089), .B(_abc_15724_n2087), .Y(_abc_15724_n2090) );
  AND2X2 AND2X2_677 ( .A(_abc_15724_n2086), .B(_abc_15724_n2090), .Y(_abc_15724_n2092_1) );
  AND2X2 AND2X2_678 ( .A(_abc_15724_n2093), .B(_abc_15724_n2091), .Y(_abc_15724_n2094) );
  AND2X2 AND2X2_679 ( .A(_abc_15724_n2094), .B(digest_update_bF_buf2), .Y(_abc_15724_n2095) );
  AND2X2 AND2X2_68 ( .A(_abc_15724_n823), .B(_abc_15724_n754), .Y(_abc_15724_n824_1) );
  AND2X2 AND2X2_680 ( .A(_auto_iopadmap_cc_313_execute_26059_103_), .B(b_reg_7_), .Y(_abc_15724_n2102) );
  AND2X2 AND2X2_681 ( .A(_abc_15724_n2103), .B(_abc_15724_n2101_1), .Y(_abc_15724_n2104) );
  AND2X2 AND2X2_682 ( .A(_abc_15724_n2100), .B(_abc_15724_n2104), .Y(_abc_15724_n2105_1) );
  AND2X2 AND2X2_683 ( .A(_abc_15724_n2099), .B(_abc_15724_n2106), .Y(_abc_15724_n2107) );
  AND2X2 AND2X2_684 ( .A(_abc_15724_n2109_1), .B(_abc_15724_n2098), .Y(H1_reg_7__FF_INPUT) );
  AND2X2 AND2X2_685 ( .A(_auto_iopadmap_cc_313_execute_26059_104_), .B(b_reg_8_), .Y(_abc_15724_n2112) );
  AND2X2 AND2X2_686 ( .A(_abc_15724_n2113), .B(_abc_15724_n2111), .Y(_abc_15724_n2114_1) );
  AND2X2 AND2X2_687 ( .A(_abc_15724_n2099), .B(_abc_15724_n2101_1), .Y(_abc_15724_n2115) );
  AND2X2 AND2X2_688 ( .A(_abc_15724_n2116), .B(_abc_15724_n2114_1), .Y(_abc_15724_n2118) );
  AND2X2 AND2X2_689 ( .A(_abc_15724_n2119_1), .B(_abc_15724_n2117), .Y(_abc_15724_n2120) );
  AND2X2 AND2X2_69 ( .A(_abc_15724_n717), .B(_abc_15724_n827), .Y(_abc_15724_n828) );
  AND2X2 AND2X2_690 ( .A(_abc_15724_n2120), .B(digest_update_bF_buf0), .Y(_abc_15724_n2121) );
  AND2X2 AND2X2_691 ( .A(_abc_15724_n2122), .B(_abc_15724_n850_bF_buf7), .Y(_abc_15724_n2123_1) );
  AND2X2 AND2X2_692 ( .A(_abc_15724_n2119_1), .B(_abc_15724_n2113), .Y(_abc_15724_n2125) );
  AND2X2 AND2X2_693 ( .A(_auto_iopadmap_cc_313_execute_26059_105_), .B(b_reg_9_), .Y(_abc_15724_n2128) );
  AND2X2 AND2X2_694 ( .A(_abc_15724_n2129), .B(_abc_15724_n2127_1), .Y(_abc_15724_n2130) );
  AND2X2 AND2X2_695 ( .A(_abc_15724_n2131_1), .B(_abc_15724_n2133), .Y(_abc_15724_n2134) );
  AND2X2 AND2X2_696 ( .A(_abc_15724_n2134), .B(digest_update_bF_buf11), .Y(_abc_15724_n2135_1) );
  AND2X2 AND2X2_697 ( .A(_abc_15724_n2136), .B(_abc_15724_n850_bF_buf6), .Y(_abc_15724_n2137) );
  AND2X2 AND2X2_698 ( .A(_abc_15724_n907_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_106_), .Y(_abc_15724_n2139_1) );
  AND2X2 AND2X2_699 ( .A(_abc_15724_n2140), .B(_abc_15724_n2129), .Y(_abc_15724_n2141) );
  AND2X2 AND2X2_7 ( .A(e_reg_18_), .B(_auto_iopadmap_cc_313_execute_26059_18_), .Y(_abc_15724_n709_1) );
  AND2X2 AND2X2_70 ( .A(_abc_15724_n719_1), .B(_abc_15724_n828), .Y(_abc_15724_n829) );
  AND2X2 AND2X2_700 ( .A(_abc_15724_n2114_1), .B(_abc_15724_n2130), .Y(_abc_15724_n2143_1) );
  AND2X2 AND2X2_701 ( .A(_abc_15724_n2116), .B(_abc_15724_n2143_1), .Y(_abc_15724_n2144) );
  AND2X2 AND2X2_702 ( .A(_auto_iopadmap_cc_313_execute_26059_106_), .B(b_reg_10_), .Y(_abc_15724_n2147) );
  AND2X2 AND2X2_703 ( .A(_abc_15724_n2148_1), .B(_abc_15724_n2146), .Y(_abc_15724_n2149) );
  AND2X2 AND2X2_704 ( .A(_abc_15724_n2145), .B(_abc_15724_n2149), .Y(_abc_15724_n2151) );
  AND2X2 AND2X2_705 ( .A(_abc_15724_n2152_1), .B(_abc_15724_n2150), .Y(_abc_15724_n2153) );
  AND2X2 AND2X2_706 ( .A(_abc_15724_n2153), .B(digest_update_bF_buf10), .Y(_abc_15724_n2154) );
  AND2X2 AND2X2_707 ( .A(_abc_15724_n2152_1), .B(_abc_15724_n2148_1), .Y(_abc_15724_n2156_1) );
  AND2X2 AND2X2_708 ( .A(_auto_iopadmap_cc_313_execute_26059_107_), .B(b_reg_11_), .Y(_abc_15724_n2159) );
  AND2X2 AND2X2_709 ( .A(_abc_15724_n2160_1), .B(_abc_15724_n2158), .Y(_abc_15724_n2161) );
  AND2X2 AND2X2_71 ( .A(_abc_15724_n713), .B(_abc_15724_n829), .Y(_abc_15724_n830) );
  AND2X2 AND2X2_710 ( .A(_abc_15724_n2162), .B(_abc_15724_n2164), .Y(_abc_15724_n2165) );
  AND2X2 AND2X2_711 ( .A(_abc_15724_n2165), .B(digest_update_bF_buf9), .Y(_abc_15724_n2166) );
  AND2X2 AND2X2_712 ( .A(_abc_15724_n2167), .B(_abc_15724_n850_bF_buf5), .Y(_abc_15724_n2168_1) );
  AND2X2 AND2X2_713 ( .A(_abc_15724_n907_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_108_), .Y(_abc_15724_n2170) );
  AND2X2 AND2X2_714 ( .A(_abc_15724_n2149), .B(_abc_15724_n2161), .Y(_abc_15724_n2171_1) );
  AND2X2 AND2X2_715 ( .A(_abc_15724_n2143_1), .B(_abc_15724_n2171_1), .Y(_abc_15724_n2172_1) );
  AND2X2 AND2X2_716 ( .A(_abc_15724_n2116), .B(_abc_15724_n2172_1), .Y(_abc_15724_n2173) );
  AND2X2 AND2X2_717 ( .A(_abc_15724_n2142), .B(_abc_15724_n2171_1), .Y(_abc_15724_n2174) );
  AND2X2 AND2X2_718 ( .A(_abc_15724_n2158), .B(_abc_15724_n2147), .Y(_abc_15724_n2175) );
  AND2X2 AND2X2_719 ( .A(_auto_iopadmap_cc_313_execute_26059_108_), .B(b_reg_12_), .Y(_abc_15724_n2180_1) );
  AND2X2 AND2X2_72 ( .A(_abc_15724_n832_1), .B(_abc_15724_n728), .Y(_abc_15724_n833_1) );
  AND2X2 AND2X2_720 ( .A(_abc_15724_n2181), .B(_abc_15724_n2179), .Y(_abc_15724_n2182_1) );
  AND2X2 AND2X2_721 ( .A(_abc_15724_n2178), .B(_abc_15724_n2182_1), .Y(_abc_15724_n2184) );
  AND2X2 AND2X2_722 ( .A(_abc_15724_n2185), .B(_abc_15724_n2183), .Y(_abc_15724_n2186) );
  AND2X2 AND2X2_723 ( .A(_abc_15724_n2186), .B(digest_update_bF_buf8), .Y(_abc_15724_n2187) );
  AND2X2 AND2X2_724 ( .A(_abc_15724_n2185), .B(_abc_15724_n2181), .Y(_abc_15724_n2189) );
  AND2X2 AND2X2_725 ( .A(_auto_iopadmap_cc_313_execute_26059_109_), .B(b_reg_13_), .Y(_abc_15724_n2192) );
  AND2X2 AND2X2_726 ( .A(_abc_15724_n2193), .B(_abc_15724_n2191), .Y(_abc_15724_n2194) );
  AND2X2 AND2X2_727 ( .A(_abc_15724_n2195_1), .B(_abc_15724_n2197), .Y(_abc_15724_n2198) );
  AND2X2 AND2X2_728 ( .A(_abc_15724_n2198), .B(digest_update_bF_buf7), .Y(_abc_15724_n2199) );
  AND2X2 AND2X2_729 ( .A(_abc_15724_n2200), .B(_abc_15724_n850_bF_buf4), .Y(_abc_15724_n2201) );
  AND2X2 AND2X2_73 ( .A(_abc_15724_n835), .B(_abc_15724_n836), .Y(_abc_15724_n837_1) );
  AND2X2 AND2X2_730 ( .A(_abc_15724_n907_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_110_), .Y(_abc_15724_n2203) );
  AND2X2 AND2X2_731 ( .A(_abc_15724_n2204), .B(_abc_15724_n2193), .Y(_abc_15724_n2205) );
  AND2X2 AND2X2_732 ( .A(_abc_15724_n2182_1), .B(_abc_15724_n2194), .Y(_abc_15724_n2207) );
  AND2X2 AND2X2_733 ( .A(_abc_15724_n2178), .B(_abc_15724_n2207), .Y(_abc_15724_n2208) );
  AND2X2 AND2X2_734 ( .A(_auto_iopadmap_cc_313_execute_26059_110_), .B(b_reg_14_), .Y(_abc_15724_n2211) );
  AND2X2 AND2X2_735 ( .A(_abc_15724_n2212), .B(_abc_15724_n2210), .Y(_abc_15724_n2213) );
  AND2X2 AND2X2_736 ( .A(_abc_15724_n2209), .B(_abc_15724_n2213), .Y(_abc_15724_n2214) );
  AND2X2 AND2X2_737 ( .A(_abc_15724_n2216), .B(digest_update_bF_buf6), .Y(_abc_15724_n2217) );
  AND2X2 AND2X2_738 ( .A(_abc_15724_n2217), .B(_abc_15724_n2215), .Y(_abc_15724_n2218) );
  AND2X2 AND2X2_739 ( .A(_abc_15724_n2215), .B(_abc_15724_n2212), .Y(_abc_15724_n2220) );
  AND2X2 AND2X2_74 ( .A(_abc_15724_n837_1), .B(_abc_15724_n702), .Y(_abc_15724_n838_1) );
  AND2X2 AND2X2_740 ( .A(_auto_iopadmap_cc_313_execute_26059_111_), .B(b_reg_15_), .Y(_abc_15724_n2223) );
  AND2X2 AND2X2_741 ( .A(_abc_15724_n2224), .B(_abc_15724_n2222), .Y(_abc_15724_n2225) );
  AND2X2 AND2X2_742 ( .A(_abc_15724_n2226), .B(_abc_15724_n2228), .Y(_abc_15724_n2229) );
  AND2X2 AND2X2_743 ( .A(_abc_15724_n2229), .B(digest_update_bF_buf5), .Y(_abc_15724_n2230) );
  AND2X2 AND2X2_744 ( .A(_abc_15724_n2231), .B(_abc_15724_n850_bF_buf3), .Y(_abc_15724_n2232) );
  AND2X2 AND2X2_745 ( .A(_abc_15724_n2213), .B(_abc_15724_n2225), .Y(_abc_15724_n2234) );
  AND2X2 AND2X2_746 ( .A(_abc_15724_n2206), .B(_abc_15724_n2234), .Y(_abc_15724_n2235) );
  AND2X2 AND2X2_747 ( .A(_abc_15724_n2222), .B(_abc_15724_n2211), .Y(_abc_15724_n2236) );
  AND2X2 AND2X2_748 ( .A(_abc_15724_n2207), .B(_abc_15724_n2234), .Y(_abc_15724_n2239) );
  AND2X2 AND2X2_749 ( .A(_abc_15724_n2178), .B(_abc_15724_n2239), .Y(_abc_15724_n2240) );
  AND2X2 AND2X2_75 ( .A(_abc_15724_n834_1), .B(_abc_15724_n838_1), .Y(_abc_15724_n839) );
  AND2X2 AND2X2_750 ( .A(_auto_iopadmap_cc_313_execute_26059_112_), .B(b_reg_16_), .Y(_abc_15724_n2243) );
  AND2X2 AND2X2_751 ( .A(_abc_15724_n2244), .B(_abc_15724_n2242), .Y(_abc_15724_n2245) );
  AND2X2 AND2X2_752 ( .A(_abc_15724_n2241), .B(_abc_15724_n2245), .Y(_abc_15724_n2247) );
  AND2X2 AND2X2_753 ( .A(_abc_15724_n2248), .B(_abc_15724_n2246_1), .Y(_abc_15724_n2249) );
  AND2X2 AND2X2_754 ( .A(_abc_15724_n2249), .B(digest_update_bF_buf4), .Y(_abc_15724_n2250_1) );
  AND2X2 AND2X2_755 ( .A(_abc_15724_n2251), .B(_abc_15724_n850_bF_buf2), .Y(_abc_15724_n2252) );
  AND2X2 AND2X2_756 ( .A(_auto_iopadmap_cc_313_execute_26059_113_), .B(b_reg_17_), .Y(_abc_15724_n2255) );
  AND2X2 AND2X2_757 ( .A(_abc_15724_n2256), .B(_abc_15724_n2254), .Y(_abc_15724_n2257) );
  AND2X2 AND2X2_758 ( .A(_abc_15724_n2248), .B(_abc_15724_n2244), .Y(_abc_15724_n2258) );
  AND2X2 AND2X2_759 ( .A(_abc_15724_n2259), .B(_abc_15724_n2257), .Y(_abc_15724_n2261) );
  AND2X2 AND2X2_76 ( .A(e_reg_22_), .B(_auto_iopadmap_cc_313_execute_26059_22_), .Y(_abc_15724_n842) );
  AND2X2 AND2X2_760 ( .A(_abc_15724_n2262), .B(_abc_15724_n2260), .Y(_abc_15724_n2263) );
  AND2X2 AND2X2_761 ( .A(_abc_15724_n2263), .B(digest_update_bF_buf3), .Y(_abc_15724_n2264) );
  AND2X2 AND2X2_762 ( .A(_abc_15724_n907_1_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_113_), .Y(_abc_15724_n2265) );
  AND2X2 AND2X2_763 ( .A(_abc_15724_n2262), .B(_abc_15724_n2256), .Y(_abc_15724_n2267) );
  AND2X2 AND2X2_764 ( .A(_auto_iopadmap_cc_313_execute_26059_114_), .B(b_reg_18_), .Y(_abc_15724_n2270) );
  AND2X2 AND2X2_765 ( .A(_abc_15724_n2271), .B(_abc_15724_n2269), .Y(_abc_15724_n2272) );
  AND2X2 AND2X2_766 ( .A(_abc_15724_n2268), .B(_abc_15724_n2272), .Y(_abc_15724_n2274) );
  AND2X2 AND2X2_767 ( .A(_abc_15724_n2275), .B(_abc_15724_n2273), .Y(_abc_15724_n2276) );
  AND2X2 AND2X2_768 ( .A(_abc_15724_n2276), .B(digest_update_bF_buf2), .Y(_abc_15724_n2277) );
  AND2X2 AND2X2_769 ( .A(_abc_15724_n2278), .B(_abc_15724_n850_bF_buf1), .Y(_abc_15724_n2279) );
  AND2X2 AND2X2_77 ( .A(_abc_15724_n843), .B(_abc_15724_n841), .Y(_abc_15724_n844_1) );
  AND2X2 AND2X2_770 ( .A(_auto_iopadmap_cc_313_execute_26059_115_), .B(b_reg_19_), .Y(_abc_15724_n2283) );
  AND2X2 AND2X2_771 ( .A(_abc_15724_n2284), .B(_abc_15724_n2282), .Y(_abc_15724_n2285) );
  AND2X2 AND2X2_772 ( .A(_abc_15724_n2289), .B(_abc_15724_n2286), .Y(_abc_15724_n2290) );
  AND2X2 AND2X2_773 ( .A(_abc_15724_n2290), .B(digest_update_bF_buf1), .Y(_abc_15724_n2291_1) );
  AND2X2 AND2X2_774 ( .A(_abc_15724_n2292), .B(_abc_15724_n850_bF_buf0), .Y(_abc_15724_n2293) );
  AND2X2 AND2X2_775 ( .A(_abc_15724_n907_1_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_116_), .Y(_abc_15724_n2295) );
  AND2X2 AND2X2_776 ( .A(_abc_15724_n2254), .B(_abc_15724_n2243), .Y(_abc_15724_n2296) );
  AND2X2 AND2X2_777 ( .A(_abc_15724_n2272), .B(_abc_15724_n2285), .Y(_abc_15724_n2298) );
  AND2X2 AND2X2_778 ( .A(_abc_15724_n2298), .B(_abc_15724_n2297), .Y(_abc_15724_n2299) );
  AND2X2 AND2X2_779 ( .A(_abc_15724_n2282), .B(_abc_15724_n2270), .Y(_abc_15724_n2300) );
  AND2X2 AND2X2_78 ( .A(_abc_15724_n840_1), .B(_abc_15724_n844_1), .Y(_abc_15724_n846) );
  AND2X2 AND2X2_780 ( .A(_abc_15724_n2245), .B(_abc_15724_n2257), .Y(_abc_15724_n2303) );
  AND2X2 AND2X2_781 ( .A(_abc_15724_n2303), .B(_abc_15724_n2298), .Y(_abc_15724_n2304) );
  AND2X2 AND2X2_782 ( .A(_abc_15724_n2241), .B(_abc_15724_n2304), .Y(_abc_15724_n2305) );
  AND2X2 AND2X2_783 ( .A(_auto_iopadmap_cc_313_execute_26059_116_), .B(b_reg_20_), .Y(_abc_15724_n2308) );
  AND2X2 AND2X2_784 ( .A(_abc_15724_n2309), .B(_abc_15724_n2307), .Y(_abc_15724_n2310) );
  AND2X2 AND2X2_785 ( .A(_abc_15724_n2306), .B(_abc_15724_n2310), .Y(_abc_15724_n2312) );
  AND2X2 AND2X2_786 ( .A(_abc_15724_n2313), .B(_abc_15724_n2311), .Y(_abc_15724_n2314) );
  AND2X2 AND2X2_787 ( .A(_abc_15724_n2314), .B(digest_update_bF_buf0), .Y(_abc_15724_n2315) );
  AND2X2 AND2X2_788 ( .A(_abc_15724_n907_1_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_117_), .Y(_abc_15724_n2317) );
  AND2X2 AND2X2_789 ( .A(_auto_iopadmap_cc_313_execute_26059_117_), .B(b_reg_21_), .Y(_abc_15724_n2319) );
  AND2X2 AND2X2_79 ( .A(_abc_15724_n847_1), .B(_abc_15724_n845_1), .Y(_abc_15724_n848) );
  AND2X2 AND2X2_790 ( .A(_abc_15724_n2320), .B(_abc_15724_n2318), .Y(_abc_15724_n2321) );
  AND2X2 AND2X2_791 ( .A(_abc_15724_n2322), .B(_abc_15724_n2321), .Y(_abc_15724_n2324) );
  AND2X2 AND2X2_792 ( .A(_abc_15724_n2325), .B(digest_update_bF_buf11), .Y(_abc_15724_n2326_1) );
  AND2X2 AND2X2_793 ( .A(_abc_15724_n2326_1), .B(_abc_15724_n2323), .Y(_abc_15724_n2327) );
  AND2X2 AND2X2_794 ( .A(_auto_iopadmap_cc_313_execute_26059_118_), .B(b_reg_22_), .Y(_abc_15724_n2331) );
  AND2X2 AND2X2_795 ( .A(_abc_15724_n2332), .B(_abc_15724_n2330_1), .Y(_abc_15724_n2333) );
  AND2X2 AND2X2_796 ( .A(_abc_15724_n2329), .B(_abc_15724_n2333), .Y(_abc_15724_n2335) );
  AND2X2 AND2X2_797 ( .A(_abc_15724_n2336), .B(_abc_15724_n2334), .Y(_abc_15724_n2337) );
  AND2X2 AND2X2_798 ( .A(_abc_15724_n2337), .B(digest_update_bF_buf10), .Y(_abc_15724_n2338) );
  AND2X2 AND2X2_799 ( .A(_abc_15724_n2339), .B(_abc_15724_n850_bF_buf8), .Y(_abc_15724_n2340) );
  AND2X2 AND2X2_8 ( .A(_abc_15724_n710_1), .B(_abc_15724_n711), .Y(_abc_15724_n712) );
  AND2X2 AND2X2_80 ( .A(_abc_15724_n848), .B(digest_update_bF_buf11), .Y(_abc_15724_n849) );
  AND2X2 AND2X2_800 ( .A(_auto_iopadmap_cc_313_execute_26059_119_), .B(b_reg_23_), .Y(_abc_15724_n2345) );
  AND2X2 AND2X2_801 ( .A(_abc_15724_n2346), .B(_abc_15724_n2344), .Y(_abc_15724_n2347) );
  AND2X2 AND2X2_802 ( .A(_abc_15724_n2343), .B(_abc_15724_n2347), .Y(_abc_15724_n2348) );
  AND2X2 AND2X2_803 ( .A(_abc_15724_n2342), .B(_abc_15724_n2349), .Y(_abc_15724_n2350) );
  AND2X2 AND2X2_804 ( .A(_abc_15724_n2351), .B(digest_update_bF_buf9), .Y(_abc_15724_n2352) );
  AND2X2 AND2X2_805 ( .A(_abc_15724_n2353), .B(_abc_15724_n850_bF_buf7), .Y(_abc_15724_n2354) );
  AND2X2 AND2X2_806 ( .A(_abc_15724_n2310), .B(_abc_15724_n2321), .Y(_abc_15724_n2356) );
  AND2X2 AND2X2_807 ( .A(_abc_15724_n2333), .B(_abc_15724_n2347), .Y(_abc_15724_n2357) );
  AND2X2 AND2X2_808 ( .A(_abc_15724_n2356), .B(_abc_15724_n2357), .Y(_abc_15724_n2358) );
  AND2X2 AND2X2_809 ( .A(_abc_15724_n2304), .B(_abc_15724_n2358), .Y(_abc_15724_n2359) );
  AND2X2 AND2X2_81 ( .A(init), .B(_auto_iopadmap_cc_313_execute_26222), .Y(_abc_15724_n851) );
  AND2X2 AND2X2_810 ( .A(_abc_15724_n2241), .B(_abc_15724_n2359), .Y(_abc_15724_n2360) );
  AND2X2 AND2X2_811 ( .A(_abc_15724_n2302), .B(_abc_15724_n2358), .Y(_abc_15724_n2361) );
  AND2X2 AND2X2_812 ( .A(_abc_15724_n2344), .B(_abc_15724_n2331), .Y(_abc_15724_n2362) );
  AND2X2 AND2X2_813 ( .A(_abc_15724_n2318), .B(_abc_15724_n2308), .Y(_abc_15724_n2364) );
  AND2X2 AND2X2_814 ( .A(_abc_15724_n2357), .B(_abc_15724_n2365), .Y(_abc_15724_n2366_1) );
  AND2X2 AND2X2_815 ( .A(_auto_iopadmap_cc_313_execute_26059_120_), .B(b_reg_24_), .Y(_abc_15724_n2371) );
  AND2X2 AND2X2_816 ( .A(_abc_15724_n2372), .B(_abc_15724_n2370_1), .Y(_abc_15724_n2373) );
  AND2X2 AND2X2_817 ( .A(_abc_15724_n2369), .B(_abc_15724_n2373), .Y(_abc_15724_n2375) );
  AND2X2 AND2X2_818 ( .A(_abc_15724_n2376), .B(_abc_15724_n2374), .Y(_abc_15724_n2377) );
  AND2X2 AND2X2_819 ( .A(_abc_15724_n2377), .B(digest_update_bF_buf8), .Y(_abc_15724_n2378) );
  AND2X2 AND2X2_82 ( .A(_abc_15724_n852), .B(_abc_15724_n850_bF_buf8), .Y(_abc_15724_n853_1) );
  AND2X2 AND2X2_820 ( .A(_abc_15724_n2379), .B(_abc_15724_n850_bF_buf6), .Y(_abc_15724_n2380) );
  AND2X2 AND2X2_821 ( .A(_abc_15724_n2376), .B(_abc_15724_n2372), .Y(_abc_15724_n2382) );
  AND2X2 AND2X2_822 ( .A(_auto_iopadmap_cc_313_execute_26059_121_), .B(b_reg_25_), .Y(_abc_15724_n2385) );
  AND2X2 AND2X2_823 ( .A(_abc_15724_n2386), .B(_abc_15724_n2384), .Y(_abc_15724_n2387) );
  AND2X2 AND2X2_824 ( .A(_abc_15724_n2388), .B(_abc_15724_n2390), .Y(_abc_15724_n2391) );
  AND2X2 AND2X2_825 ( .A(_abc_15724_n2391), .B(digest_update_bF_buf7), .Y(_abc_15724_n2392) );
  AND2X2 AND2X2_826 ( .A(_abc_15724_n2393), .B(_abc_15724_n850_bF_buf5), .Y(_abc_15724_n2394) );
  AND2X2 AND2X2_827 ( .A(_abc_15724_n2373), .B(_abc_15724_n2387), .Y(_abc_15724_n2396) );
  AND2X2 AND2X2_828 ( .A(_abc_15724_n2369), .B(_abc_15724_n2396), .Y(_abc_15724_n2397) );
  AND2X2 AND2X2_829 ( .A(_abc_15724_n2384), .B(_abc_15724_n2371), .Y(_abc_15724_n2398) );
  AND2X2 AND2X2_83 ( .A(e_reg_23_), .B(_auto_iopadmap_cc_313_execute_26059_23_), .Y(_abc_15724_n857) );
  AND2X2 AND2X2_830 ( .A(_auto_iopadmap_cc_313_execute_26059_122_), .B(b_reg_26_), .Y(_abc_15724_n2402) );
  AND2X2 AND2X2_831 ( .A(_abc_15724_n2403), .B(_abc_15724_n2401), .Y(_abc_15724_n2404) );
  AND2X2 AND2X2_832 ( .A(_abc_15724_n2400), .B(_abc_15724_n2404), .Y(_abc_15724_n2406_1) );
  AND2X2 AND2X2_833 ( .A(_abc_15724_n2407), .B(_abc_15724_n2405), .Y(_abc_15724_n2408) );
  AND2X2 AND2X2_834 ( .A(_abc_15724_n2408), .B(digest_update_bF_buf6), .Y(_abc_15724_n2409) );
  AND2X2 AND2X2_835 ( .A(_abc_15724_n2410), .B(_abc_15724_n850_bF_buf4), .Y(_abc_15724_n2411) );
  AND2X2 AND2X2_836 ( .A(_abc_15724_n2407), .B(_abc_15724_n2403), .Y(_abc_15724_n2413) );
  AND2X2 AND2X2_837 ( .A(_auto_iopadmap_cc_313_execute_26059_123_), .B(b_reg_27_), .Y(_abc_15724_n2416) );
  AND2X2 AND2X2_838 ( .A(_abc_15724_n2417), .B(_abc_15724_n2415), .Y(_abc_15724_n2418) );
  AND2X2 AND2X2_839 ( .A(_abc_15724_n2419), .B(_abc_15724_n2421), .Y(_abc_15724_n2422) );
  AND2X2 AND2X2_84 ( .A(_abc_15724_n858), .B(_abc_15724_n856), .Y(_abc_15724_n859) );
  AND2X2 AND2X2_840 ( .A(_abc_15724_n2422), .B(digest_update_bF_buf5), .Y(_abc_15724_n2423) );
  AND2X2 AND2X2_841 ( .A(_abc_15724_n2424), .B(_abc_15724_n850_bF_buf3), .Y(_abc_15724_n2425) );
  AND2X2 AND2X2_842 ( .A(_abc_15724_n907_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_124_), .Y(_abc_15724_n2427) );
  AND2X2 AND2X2_843 ( .A(_abc_15724_n2415), .B(_abc_15724_n2402), .Y(_abc_15724_n2428) );
  AND2X2 AND2X2_844 ( .A(_abc_15724_n2404), .B(_abc_15724_n2418), .Y(_abc_15724_n2430) );
  AND2X2 AND2X2_845 ( .A(_abc_15724_n2430), .B(_abc_15724_n2399), .Y(_abc_15724_n2431) );
  AND2X2 AND2X2_846 ( .A(_abc_15724_n2396), .B(_abc_15724_n2430), .Y(_abc_15724_n2433) );
  AND2X2 AND2X2_847 ( .A(_abc_15724_n2369), .B(_abc_15724_n2433), .Y(_abc_15724_n2434) );
  AND2X2 AND2X2_848 ( .A(_auto_iopadmap_cc_313_execute_26059_124_), .B(b_reg_28_), .Y(_abc_15724_n2437) );
  AND2X2 AND2X2_849 ( .A(_abc_15724_n2438), .B(_abc_15724_n2436), .Y(_abc_15724_n2439) );
  AND2X2 AND2X2_85 ( .A(_abc_15724_n863_1), .B(_abc_15724_n860), .Y(_abc_15724_n864_1) );
  AND2X2 AND2X2_850 ( .A(_abc_15724_n2435), .B(_abc_15724_n2439), .Y(_abc_15724_n2441) );
  AND2X2 AND2X2_851 ( .A(_abc_15724_n2442), .B(_abc_15724_n2440), .Y(_abc_15724_n2443) );
  AND2X2 AND2X2_852 ( .A(_abc_15724_n2443), .B(digest_update_bF_buf4), .Y(_abc_15724_n2444) );
  AND2X2 AND2X2_853 ( .A(_abc_15724_n2442), .B(_abc_15724_n2438), .Y(_abc_15724_n2446) );
  AND2X2 AND2X2_854 ( .A(_auto_iopadmap_cc_313_execute_26059_125_), .B(b_reg_29_), .Y(_abc_15724_n2448) );
  AND2X2 AND2X2_855 ( .A(_abc_15724_n2449_1), .B(_abc_15724_n2447), .Y(_abc_15724_n2450) );
  AND2X2 AND2X2_856 ( .A(_abc_15724_n2446), .B(_abc_15724_n2450), .Y(_abc_15724_n2451) );
  AND2X2 AND2X2_857 ( .A(_abc_15724_n2452), .B(_abc_15724_n2453), .Y(_abc_15724_n2454) );
  AND2X2 AND2X2_858 ( .A(_abc_15724_n2455), .B(digest_update_bF_buf3), .Y(_abc_15724_n2456) );
  AND2X2 AND2X2_859 ( .A(_abc_15724_n2457), .B(_abc_15724_n850_bF_buf2), .Y(_abc_15724_n2458) );
  AND2X2 AND2X2_86 ( .A(_abc_15724_n864_1), .B(digest_update_bF_buf9), .Y(_abc_15724_n865) );
  AND2X2 AND2X2_860 ( .A(_auto_iopadmap_cc_313_execute_26059_126_), .B(b_reg_30_), .Y(_abc_15724_n2461) );
  AND2X2 AND2X2_861 ( .A(_abc_15724_n2462), .B(_abc_15724_n2460), .Y(_abc_15724_n2463) );
  AND2X2 AND2X2_862 ( .A(_abc_15724_n2450), .B(_abc_15724_n2437), .Y(_abc_15724_n2464) );
  AND2X2 AND2X2_863 ( .A(_abc_15724_n2439), .B(_abc_15724_n2450), .Y(_abc_15724_n2466) );
  AND2X2 AND2X2_864 ( .A(_abc_15724_n2435), .B(_abc_15724_n2466), .Y(_abc_15724_n2467) );
  AND2X2 AND2X2_865 ( .A(_abc_15724_n2468), .B(_abc_15724_n2463), .Y(_abc_15724_n2470) );
  AND2X2 AND2X2_866 ( .A(_abc_15724_n2471), .B(_abc_15724_n2469), .Y(_abc_15724_n2472) );
  AND2X2 AND2X2_867 ( .A(_abc_15724_n2472), .B(digest_update_bF_buf2), .Y(_abc_15724_n2473) );
  AND2X2 AND2X2_868 ( .A(_abc_15724_n2474), .B(_abc_15724_n850_bF_buf1), .Y(_abc_15724_n2475) );
  AND2X2 AND2X2_869 ( .A(_abc_15724_n2479), .B(_abc_15724_n2481), .Y(_abc_15724_n2482) );
  AND2X2 AND2X2_87 ( .A(_abc_15724_n866_1), .B(_abc_15724_n850_bF_buf7), .Y(_abc_15724_n867) );
  AND2X2 AND2X2_870 ( .A(_abc_15724_n2486), .B(_abc_15724_n2484_1), .Y(_abc_15724_n2487) );
  AND2X2 AND2X2_871 ( .A(_abc_15724_n2487), .B(digest_update_bF_buf1), .Y(_abc_15724_n2488_1) );
  AND2X2 AND2X2_872 ( .A(_abc_15724_n2489), .B(_abc_15724_n850_bF_buf0), .Y(_abc_15724_n2490) );
  AND2X2 AND2X2_873 ( .A(_auto_iopadmap_cc_313_execute_26059_128_), .B(a_reg_0_), .Y(_abc_15724_n2493) );
  AND2X2 AND2X2_874 ( .A(_abc_15724_n2494), .B(digest_update_bF_buf0), .Y(_abc_15724_n2495) );
  AND2X2 AND2X2_875 ( .A(_abc_15724_n2495), .B(_abc_15724_n2492), .Y(_abc_15724_n2496) );
  AND2X2 AND2X2_876 ( .A(_abc_15724_n2497), .B(_abc_15724_n850_bF_buf8), .Y(_abc_15724_n2498) );
  AND2X2 AND2X2_877 ( .A(_auto_iopadmap_cc_313_execute_26059_129_), .B(a_reg_1_), .Y(_abc_15724_n2501) );
  AND2X2 AND2X2_878 ( .A(_abc_15724_n2502), .B(_abc_15724_n2500), .Y(_abc_15724_n2503) );
  AND2X2 AND2X2_879 ( .A(_abc_15724_n2503), .B(_abc_15724_n2493), .Y(_abc_15724_n2505) );
  AND2X2 AND2X2_88 ( .A(_abc_15724_n844_1), .B(_abc_15724_n859), .Y(_abc_15724_n869) );
  AND2X2 AND2X2_880 ( .A(_abc_15724_n2506), .B(_abc_15724_n2504), .Y(_abc_15724_n2507) );
  AND2X2 AND2X2_881 ( .A(_abc_15724_n2507), .B(digest_update_bF_buf11), .Y(_abc_15724_n2508) );
  AND2X2 AND2X2_882 ( .A(_abc_15724_n907_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_129_), .Y(_abc_15724_n2509) );
  AND2X2 AND2X2_883 ( .A(_abc_15724_n2506), .B(_abc_15724_n2502), .Y(_abc_15724_n2511) );
  AND2X2 AND2X2_884 ( .A(_auto_iopadmap_cc_313_execute_26059_130_), .B(a_reg_2_), .Y(_abc_15724_n2513) );
  AND2X2 AND2X2_885 ( .A(_abc_15724_n2514), .B(_abc_15724_n2512), .Y(_abc_15724_n2515) );
  AND2X2 AND2X2_886 ( .A(_abc_15724_n2519), .B(_abc_15724_n2517), .Y(_abc_15724_n2520) );
  AND2X2 AND2X2_887 ( .A(_abc_15724_n2520), .B(digest_update_bF_buf10), .Y(_abc_15724_n2521) );
  AND2X2 AND2X2_888 ( .A(_abc_15724_n907_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_130_), .Y(_abc_15724_n2522) );
  AND2X2 AND2X2_889 ( .A(_abc_15724_n2517), .B(_abc_15724_n2514), .Y(_abc_15724_n2524_1) );
  AND2X2 AND2X2_89 ( .A(_abc_15724_n838_1), .B(_abc_15724_n869), .Y(_abc_15724_n870) );
  AND2X2 AND2X2_890 ( .A(_auto_iopadmap_cc_313_execute_26059_131_), .B(a_reg_3_), .Y(_abc_15724_n2527_1) );
  AND2X2 AND2X2_891 ( .A(_abc_15724_n2528), .B(_abc_15724_n2526), .Y(_abc_15724_n2529) );
  AND2X2 AND2X2_892 ( .A(_abc_15724_n2530), .B(_abc_15724_n2532), .Y(_abc_15724_n2533) );
  AND2X2 AND2X2_893 ( .A(_abc_15724_n2533), .B(digest_update_bF_buf9), .Y(_abc_15724_n2534) );
  AND2X2 AND2X2_894 ( .A(_abc_15724_n907_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_131_), .Y(_abc_15724_n2535) );
  AND2X2 AND2X2_895 ( .A(_auto_iopadmap_cc_313_execute_26059_132_), .B(a_reg_4_), .Y(_abc_15724_n2538) );
  AND2X2 AND2X2_896 ( .A(_abc_15724_n2539), .B(_abc_15724_n2537), .Y(_abc_15724_n2540) );
  AND2X2 AND2X2_897 ( .A(_abc_15724_n2543), .B(_abc_15724_n2528), .Y(_abc_15724_n2544) );
  AND2X2 AND2X2_898 ( .A(_abc_15724_n2547), .B(_abc_15724_n2545), .Y(_abc_15724_n2548) );
  AND2X2 AND2X2_899 ( .A(_abc_15724_n2548), .B(digest_update_bF_buf8), .Y(_abc_15724_n2549) );
  AND2X2 AND2X2_9 ( .A(_abc_15724_n708_1), .B(_abc_15724_n712), .Y(_abc_15724_n713) );
  AND2X2 AND2X2_90 ( .A(_abc_15724_n830), .B(_abc_15724_n870), .Y(_abc_15724_n871) );
  AND2X2 AND2X2_900 ( .A(_abc_15724_n907_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_132_), .Y(_abc_15724_n2550) );
  AND2X2 AND2X2_901 ( .A(_abc_15724_n907_1_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_133_), .Y(_abc_15724_n2552) );
  AND2X2 AND2X2_902 ( .A(_abc_15724_n2545), .B(_abc_15724_n2539), .Y(_abc_15724_n2553) );
  AND2X2 AND2X2_903 ( .A(_auto_iopadmap_cc_313_execute_26059_133_), .B(a_reg_5_), .Y(_abc_15724_n2555) );
  AND2X2 AND2X2_904 ( .A(_abc_15724_n2556), .B(_abc_15724_n2554), .Y(_abc_15724_n2557) );
  AND2X2 AND2X2_905 ( .A(_abc_15724_n2561), .B(digest_update_bF_buf7), .Y(_abc_15724_n2562) );
  AND2X2 AND2X2_906 ( .A(_abc_15724_n2562), .B(_abc_15724_n2559), .Y(_abc_15724_n2563) );
  AND2X2 AND2X2_907 ( .A(_abc_15724_n907_1_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_134_), .Y(_abc_15724_n2565) );
  AND2X2 AND2X2_908 ( .A(_abc_15724_n2559), .B(_abc_15724_n2556), .Y(_abc_15724_n2566) );
  AND2X2 AND2X2_909 ( .A(_auto_iopadmap_cc_313_execute_26059_134_), .B(a_reg_6_), .Y(_abc_15724_n2569) );
  AND2X2 AND2X2_91 ( .A(_abc_15724_n825_1), .B(_abc_15724_n871), .Y(_abc_15724_n872) );
  AND2X2 AND2X2_910 ( .A(_abc_15724_n2570_1), .B(_abc_15724_n2568), .Y(_abc_15724_n2571) );
  AND2X2 AND2X2_911 ( .A(_abc_15724_n2574), .B(digest_update_bF_buf6), .Y(_abc_15724_n2575) );
  AND2X2 AND2X2_912 ( .A(_abc_15724_n2575), .B(_abc_15724_n2572), .Y(_abc_15724_n2576) );
  AND2X2 AND2X2_913 ( .A(_abc_15724_n907_1_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_135_), .Y(_abc_15724_n2578) );
  AND2X2 AND2X2_914 ( .A(_auto_iopadmap_cc_313_execute_26059_135_), .B(a_reg_7_), .Y(_abc_15724_n2581) );
  AND2X2 AND2X2_915 ( .A(_abc_15724_n2582), .B(_abc_15724_n2580), .Y(_abc_15724_n2583) );
  AND2X2 AND2X2_916 ( .A(_abc_15724_n2583), .B(_abc_15724_n2569), .Y(_abc_15724_n2588) );
  AND2X2 AND2X2_917 ( .A(_abc_15724_n2589), .B(digest_update_bF_buf5), .Y(_abc_15724_n2590) );
  AND2X2 AND2X2_918 ( .A(_abc_15724_n2587), .B(_abc_15724_n2590), .Y(_abc_15724_n2591) );
  AND2X2 AND2X2_919 ( .A(_abc_15724_n2591), .B(_abc_15724_n2585), .Y(_abc_15724_n2592) );
  AND2X2 AND2X2_92 ( .A(_abc_15724_n727), .B(_abc_15724_n870), .Y(_abc_15724_n873) );
  AND2X2 AND2X2_920 ( .A(_abc_15724_n2589), .B(_abc_15724_n2582), .Y(_abc_15724_n2594) );
  AND2X2 AND2X2_921 ( .A(_abc_15724_n2587), .B(_abc_15724_n2594), .Y(_abc_15724_n2595) );
  AND2X2 AND2X2_922 ( .A(_auto_iopadmap_cc_313_execute_26059_136_), .B(a_reg_8_), .Y(_abc_15724_n2598) );
  AND2X2 AND2X2_923 ( .A(_abc_15724_n2599), .B(_abc_15724_n2597), .Y(_abc_15724_n2600) );
  AND2X2 AND2X2_924 ( .A(_abc_15724_n2596), .B(_abc_15724_n2600), .Y(_abc_15724_n2602) );
  AND2X2 AND2X2_925 ( .A(_abc_15724_n2603), .B(_abc_15724_n2601), .Y(_abc_15724_n2604) );
  AND2X2 AND2X2_926 ( .A(_abc_15724_n2604), .B(digest_update_bF_buf4), .Y(_abc_15724_n2605) );
  AND2X2 AND2X2_927 ( .A(_abc_15724_n2606), .B(_abc_15724_n850_bF_buf7), .Y(_abc_15724_n2607_1) );
  AND2X2 AND2X2_928 ( .A(_abc_15724_n2603), .B(_abc_15724_n2599), .Y(_abc_15724_n2609) );
  AND2X2 AND2X2_929 ( .A(_auto_iopadmap_cc_313_execute_26059_137_), .B(a_reg_9_), .Y(_abc_15724_n2612_1) );
  AND2X2 AND2X2_93 ( .A(_abc_15724_n704), .B(_abc_15724_n869), .Y(_abc_15724_n874) );
  AND2X2 AND2X2_930 ( .A(_abc_15724_n2613), .B(_abc_15724_n2611), .Y(_abc_15724_n2614) );
  AND2X2 AND2X2_931 ( .A(_abc_15724_n2615), .B(_abc_15724_n2617), .Y(_abc_15724_n2618) );
  AND2X2 AND2X2_932 ( .A(_abc_15724_n2618), .B(digest_update_bF_buf3), .Y(_abc_15724_n2619) );
  AND2X2 AND2X2_933 ( .A(_abc_15724_n2620), .B(_abc_15724_n850_bF_buf6), .Y(_abc_15724_n2621) );
  AND2X2 AND2X2_934 ( .A(_abc_15724_n907_1_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_138_), .Y(_abc_15724_n2623) );
  AND2X2 AND2X2_935 ( .A(_auto_iopadmap_cc_313_execute_26059_138_), .B(a_reg_10_), .Y(_abc_15724_n2625) );
  AND2X2 AND2X2_936 ( .A(_abc_15724_n2626), .B(_abc_15724_n2624), .Y(_abc_15724_n2627) );
  AND2X2 AND2X2_937 ( .A(_abc_15724_n2628), .B(_abc_15724_n2613), .Y(_abc_15724_n2629) );
  AND2X2 AND2X2_938 ( .A(_abc_15724_n2600), .B(_abc_15724_n2614), .Y(_abc_15724_n2631) );
  AND2X2 AND2X2_939 ( .A(_abc_15724_n2596), .B(_abc_15724_n2631), .Y(_abc_15724_n2632) );
  AND2X2 AND2X2_94 ( .A(_abc_15724_n856), .B(_abc_15724_n842), .Y(_abc_15724_n875_1) );
  AND2X2 AND2X2_940 ( .A(_abc_15724_n2633), .B(_abc_15724_n2627), .Y(_abc_15724_n2635) );
  AND2X2 AND2X2_941 ( .A(_abc_15724_n2636), .B(_abc_15724_n2634), .Y(_abc_15724_n2637) );
  AND2X2 AND2X2_942 ( .A(_abc_15724_n2637), .B(digest_update_bF_buf2), .Y(_abc_15724_n2638) );
  AND2X2 AND2X2_943 ( .A(_abc_15724_n2636), .B(_abc_15724_n2626), .Y(_abc_15724_n2640) );
  AND2X2 AND2X2_944 ( .A(_auto_iopadmap_cc_313_execute_26059_139_), .B(a_reg_11_), .Y(_abc_15724_n2642) );
  AND2X2 AND2X2_945 ( .A(_abc_15724_n2643), .B(_abc_15724_n2641), .Y(_abc_15724_n2644) );
  AND2X2 AND2X2_946 ( .A(_abc_15724_n2640), .B(_abc_15724_n2644), .Y(_abc_15724_n2645) );
  AND2X2 AND2X2_947 ( .A(_abc_15724_n2646), .B(_abc_15724_n2647), .Y(_abc_15724_n2648_1) );
  AND2X2 AND2X2_948 ( .A(_abc_15724_n2649), .B(digest_update_bF_buf1), .Y(_abc_15724_n2650) );
  AND2X2 AND2X2_949 ( .A(_abc_15724_n907_1_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_139_), .Y(_abc_15724_n2651) );
  AND2X2 AND2X2_95 ( .A(e_reg_24_), .B(_auto_iopadmap_cc_313_execute_26059_24_), .Y(_abc_15724_n881) );
  AND2X2 AND2X2_950 ( .A(_abc_15724_n907_1_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_140_), .Y(_abc_15724_n2653) );
  AND2X2 AND2X2_951 ( .A(_abc_15724_n2627), .B(_abc_15724_n2644), .Y(_abc_15724_n2654) );
  AND2X2 AND2X2_952 ( .A(_abc_15724_n2631), .B(_abc_15724_n2654), .Y(_abc_15724_n2655) );
  AND2X2 AND2X2_953 ( .A(_abc_15724_n2630), .B(_abc_15724_n2654), .Y(_abc_15724_n2658) );
  AND2X2 AND2X2_954 ( .A(_abc_15724_n2641), .B(_abc_15724_n2625), .Y(_abc_15724_n2659) );
  AND2X2 AND2X2_955 ( .A(_abc_15724_n2657), .B(_abc_15724_n2662), .Y(_abc_15724_n2663) );
  AND2X2 AND2X2_956 ( .A(_auto_iopadmap_cc_313_execute_26059_140_), .B(a_reg_12_), .Y(_abc_15724_n2666) );
  AND2X2 AND2X2_957 ( .A(_abc_15724_n2667), .B(_abc_15724_n2665), .Y(_abc_15724_n2668) );
  AND2X2 AND2X2_958 ( .A(_abc_15724_n2664), .B(_abc_15724_n2668), .Y(_abc_15724_n2670) );
  AND2X2 AND2X2_959 ( .A(_abc_15724_n2671), .B(_abc_15724_n2669), .Y(_abc_15724_n2672) );
  AND2X2 AND2X2_96 ( .A(_abc_15724_n882), .B(_abc_15724_n880), .Y(_abc_15724_n883) );
  AND2X2 AND2X2_960 ( .A(_abc_15724_n2672), .B(digest_update_bF_buf0), .Y(_abc_15724_n2673) );
  AND2X2 AND2X2_961 ( .A(_abc_15724_n2671), .B(_abc_15724_n2667), .Y(_abc_15724_n2675) );
  AND2X2 AND2X2_962 ( .A(_auto_iopadmap_cc_313_execute_26059_141_), .B(a_reg_13_), .Y(_abc_15724_n2678) );
  AND2X2 AND2X2_963 ( .A(_abc_15724_n2679), .B(_abc_15724_n2677), .Y(_abc_15724_n2680) );
  AND2X2 AND2X2_964 ( .A(_abc_15724_n2681), .B(_abc_15724_n2683), .Y(_abc_15724_n2684) );
  AND2X2 AND2X2_965 ( .A(_abc_15724_n2684), .B(digest_update_bF_buf11), .Y(_abc_15724_n2685) );
  AND2X2 AND2X2_966 ( .A(_abc_15724_n2686), .B(_abc_15724_n850_bF_buf5), .Y(_abc_15724_n2687_1) );
  AND2X2 AND2X2_967 ( .A(_abc_15724_n907_1_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_142_), .Y(_abc_15724_n2689) );
  AND2X2 AND2X2_968 ( .A(_auto_iopadmap_cc_313_execute_26059_142_), .B(a_reg_14_), .Y(_abc_15724_n2691_1) );
  AND2X2 AND2X2_969 ( .A(_abc_15724_n2692), .B(_abc_15724_n2690), .Y(_abc_15724_n2693) );
  AND2X2 AND2X2_97 ( .A(_abc_15724_n879), .B(_abc_15724_n883), .Y(_abc_15724_n885_1) );
  AND2X2 AND2X2_970 ( .A(_abc_15724_n2667), .B(_abc_15724_n2679), .Y(_abc_15724_n2695) );
  AND2X2 AND2X2_971 ( .A(_abc_15724_n2671), .B(_abc_15724_n2695), .Y(_abc_15724_n2696) );
  AND2X2 AND2X2_972 ( .A(_abc_15724_n2698), .B(_abc_15724_n2693), .Y(_abc_15724_n2699) );
  AND2X2 AND2X2_973 ( .A(_abc_15724_n2701), .B(digest_update_bF_buf10), .Y(_abc_15724_n2702) );
  AND2X2 AND2X2_974 ( .A(_abc_15724_n2702), .B(_abc_15724_n2700), .Y(_abc_15724_n2703) );
  AND2X2 AND2X2_975 ( .A(_abc_15724_n2700), .B(_abc_15724_n2692), .Y(_abc_15724_n2705) );
  AND2X2 AND2X2_976 ( .A(_auto_iopadmap_cc_313_execute_26059_143_), .B(a_reg_15_), .Y(_abc_15724_n2707) );
  AND2X2 AND2X2_977 ( .A(_abc_15724_n2708), .B(_abc_15724_n2706), .Y(_abc_15724_n2709) );
  AND2X2 AND2X2_978 ( .A(_abc_15724_n2713), .B(_abc_15724_n2711), .Y(_abc_15724_n2714) );
  AND2X2 AND2X2_979 ( .A(_abc_15724_n2714), .B(digest_update_bF_buf9), .Y(_abc_15724_n2715) );
  AND2X2 AND2X2_98 ( .A(_abc_15724_n886), .B(_abc_15724_n884_1), .Y(_abc_15724_n887_1) );
  AND2X2 AND2X2_980 ( .A(_abc_15724_n907_1_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_143_), .Y(_abc_15724_n2716) );
  AND2X2 AND2X2_981 ( .A(_abc_15724_n2706), .B(_abc_15724_n2691_1), .Y(_abc_15724_n2718) );
  AND2X2 AND2X2_982 ( .A(_abc_15724_n2693), .B(_abc_15724_n2709), .Y(_abc_15724_n2722) );
  AND2X2 AND2X2_983 ( .A(_abc_15724_n2724), .B(_abc_15724_n2720), .Y(_abc_15724_n2725) );
  AND2X2 AND2X2_984 ( .A(_abc_15724_n2668), .B(_abc_15724_n2680), .Y(_abc_15724_n2726) );
  AND2X2 AND2X2_985 ( .A(_abc_15724_n2726), .B(_abc_15724_n2722), .Y(_abc_15724_n2727) );
  AND2X2 AND2X2_986 ( .A(_abc_15724_n2729), .B(_abc_15724_n2725), .Y(_abc_15724_n2730) );
  AND2X2 AND2X2_987 ( .A(_auto_iopadmap_cc_313_execute_26059_144_), .B(a_reg_16_), .Y(_abc_15724_n2733) );
  AND2X2 AND2X2_988 ( .A(_abc_15724_n2734_1), .B(_abc_15724_n2732), .Y(_abc_15724_n2735) );
  AND2X2 AND2X2_989 ( .A(_abc_15724_n2731_1), .B(_abc_15724_n2735), .Y(_abc_15724_n2737) );
  AND2X2 AND2X2_99 ( .A(_abc_15724_n887_1), .B(digest_update_bF_buf8), .Y(_abc_15724_n888) );
  AND2X2 AND2X2_990 ( .A(_abc_15724_n2738), .B(_abc_15724_n2736), .Y(_abc_15724_n2739) );
  AND2X2 AND2X2_991 ( .A(_abc_15724_n2739), .B(digest_update_bF_buf8), .Y(_abc_15724_n2740) );
  AND2X2 AND2X2_992 ( .A(_abc_15724_n2741), .B(_abc_15724_n850_bF_buf4), .Y(_abc_15724_n2742) );
  AND2X2 AND2X2_993 ( .A(_auto_iopadmap_cc_313_execute_26059_145_), .B(a_reg_17_), .Y(_abc_15724_n2745) );
  AND2X2 AND2X2_994 ( .A(_abc_15724_n2746), .B(_abc_15724_n2744), .Y(_abc_15724_n2747) );
  AND2X2 AND2X2_995 ( .A(_abc_15724_n2738), .B(_abc_15724_n2734_1), .Y(_abc_15724_n2748) );
  AND2X2 AND2X2_996 ( .A(_abc_15724_n2749), .B(_abc_15724_n2747), .Y(_abc_15724_n2751) );
  AND2X2 AND2X2_997 ( .A(_abc_15724_n2752), .B(_abc_15724_n2750), .Y(_abc_15724_n2753) );
  AND2X2 AND2X2_998 ( .A(_abc_15724_n2753), .B(digest_update_bF_buf7), .Y(_abc_15724_n2754) );
  AND2X2 AND2X2_999 ( .A(_abc_15724_n907_1_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_145_), .Y(_abc_15724_n2755) );
  BUFX2 BUFX2_1 ( .A(w_mem_inst__abc_21378_n3347_1), .Y(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6) );
  BUFX2 BUFX2_10 ( .A(clk), .Y(clk_hier0_bF_buf6) );
  BUFX2 BUFX2_100 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf60) );
  BUFX2 BUFX2_101 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf59) );
  BUFX2 BUFX2_102 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf58) );
  BUFX2 BUFX2_103 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf57) );
  BUFX2 BUFX2_104 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf56) );
  BUFX2 BUFX2_105 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf55) );
  BUFX2 BUFX2_106 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf54) );
  BUFX2 BUFX2_107 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf53) );
  BUFX2 BUFX2_108 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf52) );
  BUFX2 BUFX2_109 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf51) );
  BUFX2 BUFX2_11 ( .A(clk), .Y(clk_hier0_bF_buf5) );
  BUFX2 BUFX2_110 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf50) );
  BUFX2 BUFX2_111 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf49) );
  BUFX2 BUFX2_112 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf48) );
  BUFX2 BUFX2_113 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf47) );
  BUFX2 BUFX2_114 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf46) );
  BUFX2 BUFX2_115 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf45) );
  BUFX2 BUFX2_116 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf44) );
  BUFX2 BUFX2_117 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf43) );
  BUFX2 BUFX2_118 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf42) );
  BUFX2 BUFX2_119 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf41) );
  BUFX2 BUFX2_12 ( .A(clk), .Y(clk_hier0_bF_buf4) );
  BUFX2 BUFX2_120 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf40) );
  BUFX2 BUFX2_121 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf39) );
  BUFX2 BUFX2_122 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf38) );
  BUFX2 BUFX2_123 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf37) );
  BUFX2 BUFX2_124 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf36) );
  BUFX2 BUFX2_125 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf35) );
  BUFX2 BUFX2_126 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf34) );
  BUFX2 BUFX2_127 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf33) );
  BUFX2 BUFX2_128 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf32) );
  BUFX2 BUFX2_129 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf31) );
  BUFX2 BUFX2_13 ( .A(clk), .Y(clk_hier0_bF_buf3) );
  BUFX2 BUFX2_130 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf30) );
  BUFX2 BUFX2_131 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf29) );
  BUFX2 BUFX2_132 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf28) );
  BUFX2 BUFX2_133 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf27) );
  BUFX2 BUFX2_134 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf26) );
  BUFX2 BUFX2_135 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf25) );
  BUFX2 BUFX2_136 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf24) );
  BUFX2 BUFX2_137 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf23) );
  BUFX2 BUFX2_138 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf22) );
  BUFX2 BUFX2_139 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf21) );
  BUFX2 BUFX2_14 ( .A(clk), .Y(clk_hier0_bF_buf2) );
  BUFX2 BUFX2_140 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf20) );
  BUFX2 BUFX2_141 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf19) );
  BUFX2 BUFX2_142 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf18) );
  BUFX2 BUFX2_143 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf17) );
  BUFX2 BUFX2_144 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf16) );
  BUFX2 BUFX2_145 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf15) );
  BUFX2 BUFX2_146 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf14) );
  BUFX2 BUFX2_147 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf13) );
  BUFX2 BUFX2_148 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf12) );
  BUFX2 BUFX2_149 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf11) );
  BUFX2 BUFX2_15 ( .A(clk), .Y(clk_hier0_bF_buf1) );
  BUFX2 BUFX2_150 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf10) );
  BUFX2 BUFX2_151 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf9) );
  BUFX2 BUFX2_152 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf8) );
  BUFX2 BUFX2_153 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf7) );
  BUFX2 BUFX2_154 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf6) );
  BUFX2 BUFX2_155 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf5) );
  BUFX2 BUFX2_156 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf4) );
  BUFX2 BUFX2_157 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf3) );
  BUFX2 BUFX2_158 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf2) );
  BUFX2 BUFX2_159 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf1) );
  BUFX2 BUFX2_16 ( .A(clk), .Y(clk_hier0_bF_buf0) );
  BUFX2 BUFX2_160 ( .A(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3347_1_bF_buf0) );
  BUFX2 BUFX2_161 ( .A(w_mem_inst__abc_21378_n1638_1), .Y(w_mem_inst__abc_21378_n1638_1_bF_buf4) );
  BUFX2 BUFX2_162 ( .A(w_mem_inst__abc_21378_n1638_1), .Y(w_mem_inst__abc_21378_n1638_1_bF_buf3) );
  BUFX2 BUFX2_163 ( .A(w_mem_inst__abc_21378_n1638_1), .Y(w_mem_inst__abc_21378_n1638_1_bF_buf2) );
  BUFX2 BUFX2_164 ( .A(w_mem_inst__abc_21378_n1638_1), .Y(w_mem_inst__abc_21378_n1638_1_bF_buf1) );
  BUFX2 BUFX2_165 ( .A(w_mem_inst__abc_21378_n1638_1), .Y(w_mem_inst__abc_21378_n1638_1_bF_buf0) );
  BUFX2 BUFX2_166 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf88) );
  BUFX2 BUFX2_167 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf87) );
  BUFX2 BUFX2_168 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf86) );
  BUFX2 BUFX2_169 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf85) );
  BUFX2 BUFX2_17 ( .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf7) );
  BUFX2 BUFX2_170 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf84) );
  BUFX2 BUFX2_171 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf83) );
  BUFX2 BUFX2_172 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf82) );
  BUFX2 BUFX2_173 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf81) );
  BUFX2 BUFX2_174 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf80) );
  BUFX2 BUFX2_175 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf79) );
  BUFX2 BUFX2_176 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf78) );
  BUFX2 BUFX2_177 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf77) );
  BUFX2 BUFX2_178 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf76) );
  BUFX2 BUFX2_179 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf75) );
  BUFX2 BUFX2_18 ( .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf6) );
  BUFX2 BUFX2_180 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf74) );
  BUFX2 BUFX2_181 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf73) );
  BUFX2 BUFX2_182 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf72) );
  BUFX2 BUFX2_183 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf71) );
  BUFX2 BUFX2_184 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf70) );
  BUFX2 BUFX2_185 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf69) );
  BUFX2 BUFX2_186 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf68) );
  BUFX2 BUFX2_187 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf67) );
  BUFX2 BUFX2_188 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf66) );
  BUFX2 BUFX2_189 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf65) );
  BUFX2 BUFX2_19 ( .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf5) );
  BUFX2 BUFX2_190 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf64) );
  BUFX2 BUFX2_191 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf63) );
  BUFX2 BUFX2_192 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf62) );
  BUFX2 BUFX2_193 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf61) );
  BUFX2 BUFX2_194 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf60) );
  BUFX2 BUFX2_195 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf59) );
  BUFX2 BUFX2_196 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf58) );
  BUFX2 BUFX2_197 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf57) );
  BUFX2 BUFX2_198 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf56) );
  BUFX2 BUFX2_199 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf55) );
  BUFX2 BUFX2_2 ( .A(w_mem_inst__abc_21378_n3347_1), .Y(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf5) );
  BUFX2 BUFX2_20 ( .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf4) );
  BUFX2 BUFX2_200 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf54) );
  BUFX2 BUFX2_201 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf53) );
  BUFX2 BUFX2_202 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf52) );
  BUFX2 BUFX2_203 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf51) );
  BUFX2 BUFX2_204 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf50) );
  BUFX2 BUFX2_205 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf49) );
  BUFX2 BUFX2_206 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf48) );
  BUFX2 BUFX2_207 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf47) );
  BUFX2 BUFX2_208 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf46) );
  BUFX2 BUFX2_209 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf45) );
  BUFX2 BUFX2_21 ( .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf3) );
  BUFX2 BUFX2_210 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf44) );
  BUFX2 BUFX2_211 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf43) );
  BUFX2 BUFX2_212 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf42) );
  BUFX2 BUFX2_213 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf41) );
  BUFX2 BUFX2_214 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf40) );
  BUFX2 BUFX2_215 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf39) );
  BUFX2 BUFX2_216 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf38) );
  BUFX2 BUFX2_217 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf37) );
  BUFX2 BUFX2_218 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf36) );
  BUFX2 BUFX2_219 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf35) );
  BUFX2 BUFX2_22 ( .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf2) );
  BUFX2 BUFX2_220 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf34) );
  BUFX2 BUFX2_221 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf33) );
  BUFX2 BUFX2_222 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf32) );
  BUFX2 BUFX2_223 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf31) );
  BUFX2 BUFX2_224 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf30) );
  BUFX2 BUFX2_225 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf29) );
  BUFX2 BUFX2_226 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf28) );
  BUFX2 BUFX2_227 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf27) );
  BUFX2 BUFX2_228 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf26) );
  BUFX2 BUFX2_229 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf25) );
  BUFX2 BUFX2_23 ( .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf1) );
  BUFX2 BUFX2_230 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf24) );
  BUFX2 BUFX2_231 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf23) );
  BUFX2 BUFX2_232 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf22) );
  BUFX2 BUFX2_233 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf21) );
  BUFX2 BUFX2_234 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf20) );
  BUFX2 BUFX2_235 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf19) );
  BUFX2 BUFX2_236 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf18) );
  BUFX2 BUFX2_237 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf17) );
  BUFX2 BUFX2_238 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf16) );
  BUFX2 BUFX2_239 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf15) );
  BUFX2 BUFX2_24 ( .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf0) );
  BUFX2 BUFX2_240 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf14) );
  BUFX2 BUFX2_241 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf13) );
  BUFX2 BUFX2_242 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf12) );
  BUFX2 BUFX2_243 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf11) );
  BUFX2 BUFX2_244 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf10) );
  BUFX2 BUFX2_245 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf9) );
  BUFX2 BUFX2_246 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf8) );
  BUFX2 BUFX2_247 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf7) );
  BUFX2 BUFX2_248 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf6) );
  BUFX2 BUFX2_249 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf5) );
  BUFX2 BUFX2_25 ( .A(reset_n), .Y(reset_n_hier0_bF_buf8) );
  BUFX2 BUFX2_250 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf4) );
  BUFX2 BUFX2_251 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf3) );
  BUFX2 BUFX2_252 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf2) );
  BUFX2 BUFX2_253 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf1) );
  BUFX2 BUFX2_254 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf0) );
  BUFX2 BUFX2_255 ( .A(w_mem_inst__abc_21378_n1616), .Y(w_mem_inst__abc_21378_n1616_bF_buf4) );
  BUFX2 BUFX2_256 ( .A(w_mem_inst__abc_21378_n1616), .Y(w_mem_inst__abc_21378_n1616_bF_buf3) );
  BUFX2 BUFX2_257 ( .A(w_mem_inst__abc_21378_n1616), .Y(w_mem_inst__abc_21378_n1616_bF_buf2) );
  BUFX2 BUFX2_258 ( .A(w_mem_inst__abc_21378_n1616), .Y(w_mem_inst__abc_21378_n1616_bF_buf1) );
  BUFX2 BUFX2_259 ( .A(w_mem_inst__abc_21378_n1616), .Y(w_mem_inst__abc_21378_n1616_bF_buf0) );
  BUFX2 BUFX2_26 ( .A(reset_n), .Y(reset_n_hier0_bF_buf7) );
  BUFX2 BUFX2_260 ( .A(w_mem_inst__abc_21378_n1586), .Y(w_mem_inst__abc_21378_n1586_bF_buf4) );
  BUFX2 BUFX2_261 ( .A(w_mem_inst__abc_21378_n1586), .Y(w_mem_inst__abc_21378_n1586_bF_buf3) );
  BUFX2 BUFX2_262 ( .A(w_mem_inst__abc_21378_n1586), .Y(w_mem_inst__abc_21378_n1586_bF_buf2) );
  BUFX2 BUFX2_263 ( .A(w_mem_inst__abc_21378_n1586), .Y(w_mem_inst__abc_21378_n1586_bF_buf1) );
  BUFX2 BUFX2_264 ( .A(w_mem_inst__abc_21378_n1586), .Y(w_mem_inst__abc_21378_n1586_bF_buf0) );
  BUFX2 BUFX2_265 ( .A(w_mem_inst__abc_21378_n1587), .Y(w_mem_inst__abc_21378_n1587_bF_buf4) );
  BUFX2 BUFX2_266 ( .A(w_mem_inst__abc_21378_n1587), .Y(w_mem_inst__abc_21378_n1587_bF_buf3) );
  BUFX2 BUFX2_267 ( .A(w_mem_inst__abc_21378_n1587), .Y(w_mem_inst__abc_21378_n1587_bF_buf2) );
  BUFX2 BUFX2_268 ( .A(w_mem_inst__abc_21378_n1587), .Y(w_mem_inst__abc_21378_n1587_bF_buf1) );
  BUFX2 BUFX2_269 ( .A(w_mem_inst__abc_21378_n1587), .Y(w_mem_inst__abc_21378_n1587_bF_buf0) );
  BUFX2 BUFX2_27 ( .A(reset_n), .Y(reset_n_hier0_bF_buf6) );
  BUFX2 BUFX2_270 ( .A(w_mem_inst__abc_21378_n1643_1), .Y(w_mem_inst__abc_21378_n1643_1_bF_buf4) );
  BUFX2 BUFX2_271 ( .A(w_mem_inst__abc_21378_n1643_1), .Y(w_mem_inst__abc_21378_n1643_1_bF_buf3) );
  BUFX2 BUFX2_272 ( .A(w_mem_inst__abc_21378_n1643_1), .Y(w_mem_inst__abc_21378_n1643_1_bF_buf2) );
  BUFX2 BUFX2_273 ( .A(w_mem_inst__abc_21378_n1643_1), .Y(w_mem_inst__abc_21378_n1643_1_bF_buf1) );
  BUFX2 BUFX2_274 ( .A(w_mem_inst__abc_21378_n1643_1), .Y(w_mem_inst__abc_21378_n1643_1_bF_buf0) );
  BUFX2 BUFX2_275 ( .A(w_mem_inst__abc_21378_n1618_1), .Y(w_mem_inst__abc_21378_n1618_1_bF_buf4) );
  BUFX2 BUFX2_276 ( .A(w_mem_inst__abc_21378_n1618_1), .Y(w_mem_inst__abc_21378_n1618_1_bF_buf3) );
  BUFX2 BUFX2_277 ( .A(w_mem_inst__abc_21378_n1618_1), .Y(w_mem_inst__abc_21378_n1618_1_bF_buf2) );
  BUFX2 BUFX2_278 ( .A(w_mem_inst__abc_21378_n1618_1), .Y(w_mem_inst__abc_21378_n1618_1_bF_buf1) );
  BUFX2 BUFX2_279 ( .A(w_mem_inst__abc_21378_n1618_1), .Y(w_mem_inst__abc_21378_n1618_1_bF_buf0) );
  BUFX2 BUFX2_28 ( .A(reset_n), .Y(reset_n_hier0_bF_buf5) );
  BUFX2 BUFX2_280 ( .A(_abc_15724_n3737), .Y(_abc_15724_n3737_bF_buf4) );
  BUFX2 BUFX2_281 ( .A(_abc_15724_n3737), .Y(_abc_15724_n3737_bF_buf3) );
  BUFX2 BUFX2_282 ( .A(_abc_15724_n3737), .Y(_abc_15724_n3737_bF_buf2) );
  BUFX2 BUFX2_283 ( .A(_abc_15724_n3737), .Y(_abc_15724_n3737_bF_buf1) );
  BUFX2 BUFX2_284 ( .A(_abc_15724_n3737), .Y(_abc_15724_n3737_bF_buf0) );
  BUFX2 BUFX2_285 ( .A(w_mem_inst__abc_21378_n1605), .Y(w_mem_inst__abc_21378_n1605_bF_buf4) );
  BUFX2 BUFX2_286 ( .A(w_mem_inst__abc_21378_n1605), .Y(w_mem_inst__abc_21378_n1605_bF_buf3) );
  BUFX2 BUFX2_287 ( .A(w_mem_inst__abc_21378_n1605), .Y(w_mem_inst__abc_21378_n1605_bF_buf2) );
  BUFX2 BUFX2_288 ( .A(w_mem_inst__abc_21378_n1605), .Y(w_mem_inst__abc_21378_n1605_bF_buf1) );
  BUFX2 BUFX2_289 ( .A(w_mem_inst__abc_21378_n1605), .Y(w_mem_inst__abc_21378_n1605_bF_buf0) );
  BUFX2 BUFX2_29 ( .A(reset_n), .Y(reset_n_hier0_bF_buf4) );
  BUFX2 BUFX2_290 ( .A(w_mem_inst__abc_21378_n1630_1), .Y(w_mem_inst__abc_21378_n1630_1_bF_buf4) );
  BUFX2 BUFX2_291 ( .A(w_mem_inst__abc_21378_n1630_1), .Y(w_mem_inst__abc_21378_n1630_1_bF_buf3) );
  BUFX2 BUFX2_292 ( .A(w_mem_inst__abc_21378_n1630_1), .Y(w_mem_inst__abc_21378_n1630_1_bF_buf2) );
  BUFX2 BUFX2_293 ( .A(w_mem_inst__abc_21378_n1630_1), .Y(w_mem_inst__abc_21378_n1630_1_bF_buf1) );
  BUFX2 BUFX2_294 ( .A(w_mem_inst__abc_21378_n1630_1), .Y(w_mem_inst__abc_21378_n1630_1_bF_buf0) );
  BUFX2 BUFX2_295 ( .A(w_mem_inst__abc_21378_n1610_1), .Y(w_mem_inst__abc_21378_n1610_1_bF_buf4) );
  BUFX2 BUFX2_296 ( .A(w_mem_inst__abc_21378_n1610_1), .Y(w_mem_inst__abc_21378_n1610_1_bF_buf3) );
  BUFX2 BUFX2_297 ( .A(w_mem_inst__abc_21378_n1610_1), .Y(w_mem_inst__abc_21378_n1610_1_bF_buf2) );
  BUFX2 BUFX2_298 ( .A(w_mem_inst__abc_21378_n1610_1), .Y(w_mem_inst__abc_21378_n1610_1_bF_buf1) );
  BUFX2 BUFX2_299 ( .A(w_mem_inst__abc_21378_n1610_1), .Y(w_mem_inst__abc_21378_n1610_1_bF_buf0) );
  BUFX2 BUFX2_3 ( .A(w_mem_inst__abc_21378_n3347_1), .Y(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf4) );
  BUFX2 BUFX2_30 ( .A(reset_n), .Y(reset_n_hier0_bF_buf3) );
  BUFX2 BUFX2_300 ( .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf63) );
  BUFX2 BUFX2_301 ( .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf62) );
  BUFX2 BUFX2_302 ( .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf61) );
  BUFX2 BUFX2_303 ( .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf60) );
  BUFX2 BUFX2_304 ( .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf59) );
  BUFX2 BUFX2_305 ( .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf58) );
  BUFX2 BUFX2_306 ( .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf57) );
  BUFX2 BUFX2_307 ( .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf56) );
  BUFX2 BUFX2_308 ( .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf55) );
  BUFX2 BUFX2_309 ( .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf54) );
  BUFX2 BUFX2_31 ( .A(reset_n), .Y(reset_n_hier0_bF_buf2) );
  BUFX2 BUFX2_310 ( .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf53) );
  BUFX2 BUFX2_311 ( .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf52) );
  BUFX2 BUFX2_312 ( .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf51) );
  BUFX2 BUFX2_313 ( .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf50) );
  BUFX2 BUFX2_314 ( .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf49) );
  BUFX2 BUFX2_315 ( .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf48) );
  BUFX2 BUFX2_316 ( .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf47) );
  BUFX2 BUFX2_317 ( .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf46) );
  BUFX2 BUFX2_318 ( .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf45) );
  BUFX2 BUFX2_319 ( .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf44) );
  BUFX2 BUFX2_32 ( .A(reset_n), .Y(reset_n_hier0_bF_buf1) );
  BUFX2 BUFX2_320 ( .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf43) );
  BUFX2 BUFX2_321 ( .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf42) );
  BUFX2 BUFX2_322 ( .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf41) );
  BUFX2 BUFX2_323 ( .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf40) );
  BUFX2 BUFX2_324 ( .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf39) );
  BUFX2 BUFX2_325 ( .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf38) );
  BUFX2 BUFX2_326 ( .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf37) );
  BUFX2 BUFX2_327 ( .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf36) );
  BUFX2 BUFX2_328 ( .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf35) );
  BUFX2 BUFX2_329 ( .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf34) );
  BUFX2 BUFX2_33 ( .A(reset_n), .Y(reset_n_hier0_bF_buf0) );
  BUFX2 BUFX2_330 ( .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf33) );
  BUFX2 BUFX2_331 ( .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf32) );
  BUFX2 BUFX2_332 ( .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf31) );
  BUFX2 BUFX2_333 ( .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf30) );
  BUFX2 BUFX2_334 ( .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf29) );
  BUFX2 BUFX2_335 ( .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf28) );
  BUFX2 BUFX2_336 ( .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf27) );
  BUFX2 BUFX2_337 ( .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf26) );
  BUFX2 BUFX2_338 ( .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf25) );
  BUFX2 BUFX2_339 ( .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf24) );
  BUFX2 BUFX2_34 ( .A(w_mem_inst__abc_21378_n3154_1), .Y(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf7) );
  BUFX2 BUFX2_340 ( .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf23) );
  BUFX2 BUFX2_341 ( .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf22) );
  BUFX2 BUFX2_342 ( .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf21) );
  BUFX2 BUFX2_343 ( .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf20) );
  BUFX2 BUFX2_344 ( .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf19) );
  BUFX2 BUFX2_345 ( .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf18) );
  BUFX2 BUFX2_346 ( .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf17) );
  BUFX2 BUFX2_347 ( .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf16) );
  BUFX2 BUFX2_348 ( .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf15) );
  BUFX2 BUFX2_349 ( .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf14) );
  BUFX2 BUFX2_35 ( .A(w_mem_inst__abc_21378_n3154_1), .Y(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf6) );
  BUFX2 BUFX2_350 ( .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf13) );
  BUFX2 BUFX2_351 ( .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf12) );
  BUFX2 BUFX2_352 ( .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf11) );
  BUFX2 BUFX2_353 ( .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf10) );
  BUFX2 BUFX2_354 ( .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf9) );
  BUFX2 BUFX2_355 ( .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf8) );
  BUFX2 BUFX2_356 ( .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf7) );
  BUFX2 BUFX2_357 ( .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf6) );
  BUFX2 BUFX2_358 ( .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf5) );
  BUFX2 BUFX2_359 ( .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf4) );
  BUFX2 BUFX2_36 ( .A(w_mem_inst__abc_21378_n3154_1), .Y(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf5) );
  BUFX2 BUFX2_360 ( .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf3) );
  BUFX2 BUFX2_361 ( .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf2) );
  BUFX2 BUFX2_362 ( .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf1) );
  BUFX2 BUFX2_363 ( .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf0) );
  BUFX2 BUFX2_364 ( .A(w_mem_inst__abc_21378_n1627_1), .Y(w_mem_inst__abc_21378_n1627_1_bF_buf4) );
  BUFX2 BUFX2_365 ( .A(w_mem_inst__abc_21378_n1627_1), .Y(w_mem_inst__abc_21378_n1627_1_bF_buf3) );
  BUFX2 BUFX2_366 ( .A(w_mem_inst__abc_21378_n1627_1), .Y(w_mem_inst__abc_21378_n1627_1_bF_buf2) );
  BUFX2 BUFX2_367 ( .A(w_mem_inst__abc_21378_n1627_1), .Y(w_mem_inst__abc_21378_n1627_1_bF_buf1) );
  BUFX2 BUFX2_368 ( .A(w_mem_inst__abc_21378_n1627_1), .Y(w_mem_inst__abc_21378_n1627_1_bF_buf0) );
  BUFX2 BUFX2_369 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf11) );
  BUFX2 BUFX2_37 ( .A(w_mem_inst__abc_21378_n3154_1), .Y(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf4) );
  BUFX2 BUFX2_370 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf10) );
  BUFX2 BUFX2_371 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf9) );
  BUFX2 BUFX2_372 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf8) );
  BUFX2 BUFX2_373 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf7) );
  BUFX2 BUFX2_374 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf6) );
  BUFX2 BUFX2_375 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf5) );
  BUFX2 BUFX2_376 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf4) );
  BUFX2 BUFX2_377 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf3) );
  BUFX2 BUFX2_378 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf2) );
  BUFX2 BUFX2_379 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf1) );
  BUFX2 BUFX2_38 ( .A(w_mem_inst__abc_21378_n3154_1), .Y(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf3) );
  BUFX2 BUFX2_380 ( .A(_abc_15724_n2992), .Y(_abc_15724_n2992_bF_buf0) );
  BUFX2 BUFX2_381 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf11) );
  BUFX2 BUFX2_382 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf10) );
  BUFX2 BUFX2_383 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf9) );
  BUFX2 BUFX2_384 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf8) );
  BUFX2 BUFX2_385 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf7) );
  BUFX2 BUFX2_386 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf6) );
  BUFX2 BUFX2_387 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf5) );
  BUFX2 BUFX2_388 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf4) );
  BUFX2 BUFX2_389 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf3) );
  BUFX2 BUFX2_39 ( .A(w_mem_inst__abc_21378_n3154_1), .Y(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf2) );
  BUFX2 BUFX2_390 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf2) );
  BUFX2 BUFX2_391 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf1) );
  BUFX2 BUFX2_392 ( .A(_abc_15724_n2994), .Y(_abc_15724_n2994_bF_buf0) );
  BUFX2 BUFX2_393 ( .A(_abc_15724_n850), .Y(_abc_15724_n850_bF_buf8) );
  BUFX2 BUFX2_394 ( .A(_abc_15724_n850), .Y(_abc_15724_n850_bF_buf7) );
  BUFX2 BUFX2_395 ( .A(_abc_15724_n850), .Y(_abc_15724_n850_bF_buf6) );
  BUFX2 BUFX2_396 ( .A(_abc_15724_n850), .Y(_abc_15724_n850_bF_buf5) );
  BUFX2 BUFX2_397 ( .A(_abc_15724_n850), .Y(_abc_15724_n850_bF_buf4) );
  BUFX2 BUFX2_398 ( .A(_abc_15724_n850), .Y(_abc_15724_n850_bF_buf3) );
  BUFX2 BUFX2_399 ( .A(_abc_15724_n850), .Y(_abc_15724_n850_bF_buf2) );
  BUFX2 BUFX2_4 ( .A(w_mem_inst__abc_21378_n3347_1), .Y(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf3) );
  BUFX2 BUFX2_40 ( .A(w_mem_inst__abc_21378_n3154_1), .Y(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf1) );
  BUFX2 BUFX2_400 ( .A(_abc_15724_n850), .Y(_abc_15724_n850_bF_buf1) );
  BUFX2 BUFX2_401 ( .A(_abc_15724_n850), .Y(_abc_15724_n850_bF_buf0) );
  BUFX2 BUFX2_402 ( .A(_abc_15724_n851), .Y(_abc_15724_n851_bF_buf8) );
  BUFX2 BUFX2_403 ( .A(_abc_15724_n851), .Y(_abc_15724_n851_bF_buf7) );
  BUFX2 BUFX2_404 ( .A(_abc_15724_n851), .Y(_abc_15724_n851_bF_buf6) );
  BUFX2 BUFX2_405 ( .A(_abc_15724_n851), .Y(_abc_15724_n851_bF_buf5) );
  BUFX2 BUFX2_406 ( .A(_abc_15724_n851), .Y(_abc_15724_n851_bF_buf4) );
  BUFX2 BUFX2_407 ( .A(_abc_15724_n851), .Y(_abc_15724_n851_bF_buf3) );
  BUFX2 BUFX2_408 ( .A(_abc_15724_n851), .Y(_abc_15724_n851_bF_buf2) );
  BUFX2 BUFX2_409 ( .A(_abc_15724_n851), .Y(_abc_15724_n851_bF_buf1) );
  BUFX2 BUFX2_41 ( .A(w_mem_inst__abc_21378_n3154_1), .Y(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf0) );
  BUFX2 BUFX2_410 ( .A(_abc_15724_n851), .Y(_abc_15724_n851_bF_buf0) );
  BUFX2 BUFX2_411 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf88) );
  BUFX2 BUFX2_412 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf87) );
  BUFX2 BUFX2_413 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf86) );
  BUFX2 BUFX2_414 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf85) );
  BUFX2 BUFX2_415 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf84) );
  BUFX2 BUFX2_416 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf83) );
  BUFX2 BUFX2_417 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf82) );
  BUFX2 BUFX2_418 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf81) );
  BUFX2 BUFX2_419 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf80) );
  BUFX2 BUFX2_42 ( .A(w_mem_inst__abc_21378_n3152), .Y(w_mem_inst__abc_21378_n3152_hier0_bF_buf7) );
  BUFX2 BUFX2_420 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf79) );
  BUFX2 BUFX2_421 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf78) );
  BUFX2 BUFX2_422 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf77) );
  BUFX2 BUFX2_423 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf76) );
  BUFX2 BUFX2_424 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf75) );
  BUFX2 BUFX2_425 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf74) );
  BUFX2 BUFX2_426 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf73) );
  BUFX2 BUFX2_427 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf72) );
  BUFX2 BUFX2_428 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf71) );
  BUFX2 BUFX2_429 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf70) );
  BUFX2 BUFX2_43 ( .A(w_mem_inst__abc_21378_n3152), .Y(w_mem_inst__abc_21378_n3152_hier0_bF_buf6) );
  BUFX2 BUFX2_430 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf69) );
  BUFX2 BUFX2_431 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf68) );
  BUFX2 BUFX2_432 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf67) );
  BUFX2 BUFX2_433 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf66) );
  BUFX2 BUFX2_434 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf65) );
  BUFX2 BUFX2_435 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf64) );
  BUFX2 BUFX2_436 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf63) );
  BUFX2 BUFX2_437 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf62) );
  BUFX2 BUFX2_438 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf61) );
  BUFX2 BUFX2_439 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf60) );
  BUFX2 BUFX2_44 ( .A(w_mem_inst__abc_21378_n3152), .Y(w_mem_inst__abc_21378_n3152_hier0_bF_buf5) );
  BUFX2 BUFX2_440 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf59) );
  BUFX2 BUFX2_441 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf58) );
  BUFX2 BUFX2_442 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf57) );
  BUFX2 BUFX2_443 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf56) );
  BUFX2 BUFX2_444 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf55) );
  BUFX2 BUFX2_445 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf54) );
  BUFX2 BUFX2_446 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf53) );
  BUFX2 BUFX2_447 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf52) );
  BUFX2 BUFX2_448 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf51) );
  BUFX2 BUFX2_449 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf50) );
  BUFX2 BUFX2_45 ( .A(w_mem_inst__abc_21378_n3152), .Y(w_mem_inst__abc_21378_n3152_hier0_bF_buf4) );
  BUFX2 BUFX2_450 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf49) );
  BUFX2 BUFX2_451 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf48) );
  BUFX2 BUFX2_452 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf47) );
  BUFX2 BUFX2_453 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf46) );
  BUFX2 BUFX2_454 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf45) );
  BUFX2 BUFX2_455 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf44) );
  BUFX2 BUFX2_456 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf43) );
  BUFX2 BUFX2_457 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf42) );
  BUFX2 BUFX2_458 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf41) );
  BUFX2 BUFX2_459 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf40) );
  BUFX2 BUFX2_46 ( .A(w_mem_inst__abc_21378_n3152), .Y(w_mem_inst__abc_21378_n3152_hier0_bF_buf3) );
  BUFX2 BUFX2_460 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf39) );
  BUFX2 BUFX2_461 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf38) );
  BUFX2 BUFX2_462 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf37) );
  BUFX2 BUFX2_463 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf36) );
  BUFX2 BUFX2_464 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf35) );
  BUFX2 BUFX2_465 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf34) );
  BUFX2 BUFX2_466 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf33) );
  BUFX2 BUFX2_467 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf32) );
  BUFX2 BUFX2_468 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf31) );
  BUFX2 BUFX2_469 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf30) );
  BUFX2 BUFX2_47 ( .A(w_mem_inst__abc_21378_n3152), .Y(w_mem_inst__abc_21378_n3152_hier0_bF_buf2) );
  BUFX2 BUFX2_470 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf29) );
  BUFX2 BUFX2_471 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf28) );
  BUFX2 BUFX2_472 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf27) );
  BUFX2 BUFX2_473 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf26) );
  BUFX2 BUFX2_474 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf25) );
  BUFX2 BUFX2_475 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf24) );
  BUFX2 BUFX2_476 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf23) );
  BUFX2 BUFX2_477 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf22) );
  BUFX2 BUFX2_478 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf21) );
  BUFX2 BUFX2_479 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf20) );
  BUFX2 BUFX2_48 ( .A(w_mem_inst__abc_21378_n3152), .Y(w_mem_inst__abc_21378_n3152_hier0_bF_buf1) );
  BUFX2 BUFX2_480 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf19) );
  BUFX2 BUFX2_481 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf18) );
  BUFX2 BUFX2_482 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf17) );
  BUFX2 BUFX2_483 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf16) );
  BUFX2 BUFX2_484 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf15) );
  BUFX2 BUFX2_485 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf14) );
  BUFX2 BUFX2_486 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf13) );
  BUFX2 BUFX2_487 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf12) );
  BUFX2 BUFX2_488 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf11) );
  BUFX2 BUFX2_489 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf10) );
  BUFX2 BUFX2_49 ( .A(w_mem_inst__abc_21378_n3152), .Y(w_mem_inst__abc_21378_n3152_hier0_bF_buf0) );
  BUFX2 BUFX2_490 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf9) );
  BUFX2 BUFX2_491 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf8) );
  BUFX2 BUFX2_492 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf7) );
  BUFX2 BUFX2_493 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf6) );
  BUFX2 BUFX2_494 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf5) );
  BUFX2 BUFX2_495 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf4) );
  BUFX2 BUFX2_496 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf3) );
  BUFX2 BUFX2_497 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf2) );
  BUFX2 BUFX2_498 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf1) );
  BUFX2 BUFX2_499 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf0) );
  BUFX2 BUFX2_5 ( .A(w_mem_inst__abc_21378_n3347_1), .Y(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf2) );
  BUFX2 BUFX2_50 ( .A(w_mem_inst__abc_21378_n1651_1), .Y(w_mem_inst__abc_21378_n1651_1_bF_buf4) );
  BUFX2 BUFX2_500 ( .A(w_mem_inst__abc_21378_n1654_1), .Y(w_mem_inst__abc_21378_n1654_1_bF_buf4) );
  BUFX2 BUFX2_501 ( .A(w_mem_inst__abc_21378_n1654_1), .Y(w_mem_inst__abc_21378_n1654_1_bF_buf3) );
  BUFX2 BUFX2_502 ( .A(w_mem_inst__abc_21378_n1654_1), .Y(w_mem_inst__abc_21378_n1654_1_bF_buf2) );
  BUFX2 BUFX2_503 ( .A(w_mem_inst__abc_21378_n1654_1), .Y(w_mem_inst__abc_21378_n1654_1_bF_buf1) );
  BUFX2 BUFX2_504 ( .A(w_mem_inst__abc_21378_n1654_1), .Y(w_mem_inst__abc_21378_n1654_1_bF_buf0) );
  BUFX2 BUFX2_505 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf63) );
  BUFX2 BUFX2_506 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf62) );
  BUFX2 BUFX2_507 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf61) );
  BUFX2 BUFX2_508 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf60) );
  BUFX2 BUFX2_509 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf59) );
  BUFX2 BUFX2_51 ( .A(w_mem_inst__abc_21378_n1651_1), .Y(w_mem_inst__abc_21378_n1651_1_bF_buf3) );
  BUFX2 BUFX2_510 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf58) );
  BUFX2 BUFX2_511 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf57) );
  BUFX2 BUFX2_512 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf56) );
  BUFX2 BUFX2_513 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf55) );
  BUFX2 BUFX2_514 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf54) );
  BUFX2 BUFX2_515 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf53) );
  BUFX2 BUFX2_516 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf52) );
  BUFX2 BUFX2_517 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf51) );
  BUFX2 BUFX2_518 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf50) );
  BUFX2 BUFX2_519 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf49) );
  BUFX2 BUFX2_52 ( .A(w_mem_inst__abc_21378_n1651_1), .Y(w_mem_inst__abc_21378_n1651_1_bF_buf2) );
  BUFX2 BUFX2_520 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf48) );
  BUFX2 BUFX2_521 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf47) );
  BUFX2 BUFX2_522 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf46) );
  BUFX2 BUFX2_523 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf45) );
  BUFX2 BUFX2_524 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf44) );
  BUFX2 BUFX2_525 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf43) );
  BUFX2 BUFX2_526 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf42) );
  BUFX2 BUFX2_527 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf41) );
  BUFX2 BUFX2_528 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf40) );
  BUFX2 BUFX2_529 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf39) );
  BUFX2 BUFX2_53 ( .A(w_mem_inst__abc_21378_n1651_1), .Y(w_mem_inst__abc_21378_n1651_1_bF_buf1) );
  BUFX2 BUFX2_530 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf38) );
  BUFX2 BUFX2_531 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf37) );
  BUFX2 BUFX2_532 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf36) );
  BUFX2 BUFX2_533 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf35) );
  BUFX2 BUFX2_534 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf34) );
  BUFX2 BUFX2_535 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf33) );
  BUFX2 BUFX2_536 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf32) );
  BUFX2 BUFX2_537 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf31) );
  BUFX2 BUFX2_538 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf30) );
  BUFX2 BUFX2_539 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf29) );
  BUFX2 BUFX2_54 ( .A(w_mem_inst__abc_21378_n1651_1), .Y(w_mem_inst__abc_21378_n1651_1_bF_buf0) );
  BUFX2 BUFX2_540 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf28) );
  BUFX2 BUFX2_541 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf27) );
  BUFX2 BUFX2_542 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf26) );
  BUFX2 BUFX2_543 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf25) );
  BUFX2 BUFX2_544 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf24) );
  BUFX2 BUFX2_545 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf23) );
  BUFX2 BUFX2_546 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf22) );
  BUFX2 BUFX2_547 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf21) );
  BUFX2 BUFX2_548 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf20) );
  BUFX2 BUFX2_549 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf19) );
  BUFX2 BUFX2_55 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf12) );
  BUFX2 BUFX2_550 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf18) );
  BUFX2 BUFX2_551 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf17) );
  BUFX2 BUFX2_552 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf16) );
  BUFX2 BUFX2_553 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf15) );
  BUFX2 BUFX2_554 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf14) );
  BUFX2 BUFX2_555 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf13) );
  BUFX2 BUFX2_556 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf12) );
  BUFX2 BUFX2_557 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf11) );
  BUFX2 BUFX2_558 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf10) );
  BUFX2 BUFX2_559 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf9) );
  BUFX2 BUFX2_56 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf11) );
  BUFX2 BUFX2_560 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf8) );
  BUFX2 BUFX2_561 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf7) );
  BUFX2 BUFX2_562 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf6) );
  BUFX2 BUFX2_563 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf5) );
  BUFX2 BUFX2_564 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf4) );
  BUFX2 BUFX2_565 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf3) );
  BUFX2 BUFX2_566 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf2) );
  BUFX2 BUFX2_567 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf1) );
  BUFX2 BUFX2_568 ( .A(w_mem_inst__abc_21378_n3154_1_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3154_1_bF_buf0) );
  BUFX2 BUFX2_569 ( .A(w_mem_inst__abc_21378_n1656), .Y(w_mem_inst__abc_21378_n1656_bF_buf4) );
  BUFX2 BUFX2_57 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf10) );
  BUFX2 BUFX2_570 ( .A(w_mem_inst__abc_21378_n1656), .Y(w_mem_inst__abc_21378_n1656_bF_buf3) );
  BUFX2 BUFX2_571 ( .A(w_mem_inst__abc_21378_n1656), .Y(w_mem_inst__abc_21378_n1656_bF_buf2) );
  BUFX2 BUFX2_572 ( .A(w_mem_inst__abc_21378_n1656), .Y(w_mem_inst__abc_21378_n1656_bF_buf1) );
  BUFX2 BUFX2_573 ( .A(w_mem_inst__abc_21378_n1656), .Y(w_mem_inst__abc_21378_n1656_bF_buf0) );
  BUFX2 BUFX2_574 ( .A(digest_update), .Y(digest_update_bF_buf11) );
  BUFX2 BUFX2_575 ( .A(digest_update), .Y(digest_update_bF_buf10) );
  BUFX2 BUFX2_576 ( .A(digest_update), .Y(digest_update_bF_buf9) );
  BUFX2 BUFX2_577 ( .A(digest_update), .Y(digest_update_bF_buf8) );
  BUFX2 BUFX2_578 ( .A(digest_update), .Y(digest_update_bF_buf7) );
  BUFX2 BUFX2_579 ( .A(digest_update), .Y(digest_update_bF_buf6) );
  BUFX2 BUFX2_58 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf9) );
  BUFX2 BUFX2_580 ( .A(digest_update), .Y(digest_update_bF_buf5) );
  BUFX2 BUFX2_581 ( .A(digest_update), .Y(digest_update_bF_buf4) );
  BUFX2 BUFX2_582 ( .A(digest_update), .Y(digest_update_bF_buf3) );
  BUFX2 BUFX2_583 ( .A(digest_update), .Y(digest_update_bF_buf2) );
  BUFX2 BUFX2_584 ( .A(digest_update), .Y(digest_update_bF_buf1) );
  BUFX2 BUFX2_585 ( .A(digest_update), .Y(digest_update_bF_buf0) );
  BUFX2 BUFX2_586 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3152_bF_buf63) );
  BUFX2 BUFX2_587 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3152_bF_buf62) );
  BUFX2 BUFX2_588 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3152_bF_buf61) );
  BUFX2 BUFX2_589 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3152_bF_buf60) );
  BUFX2 BUFX2_59 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf8) );
  BUFX2 BUFX2_590 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3152_bF_buf59) );
  BUFX2 BUFX2_591 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3152_bF_buf58) );
  BUFX2 BUFX2_592 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3152_bF_buf57) );
  BUFX2 BUFX2_593 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3152_bF_buf56) );
  BUFX2 BUFX2_594 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3152_bF_buf55) );
  BUFX2 BUFX2_595 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3152_bF_buf54) );
  BUFX2 BUFX2_596 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3152_bF_buf53) );
  BUFX2 BUFX2_597 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3152_bF_buf52) );
  BUFX2 BUFX2_598 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3152_bF_buf51) );
  BUFX2 BUFX2_599 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3152_bF_buf50) );
  BUFX2 BUFX2_6 ( .A(w_mem_inst__abc_21378_n3347_1), .Y(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf1) );
  BUFX2 BUFX2_60 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf7) );
  BUFX2 BUFX2_600 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3152_bF_buf49) );
  BUFX2 BUFX2_601 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3152_bF_buf48) );
  BUFX2 BUFX2_602 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3152_bF_buf47) );
  BUFX2 BUFX2_603 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3152_bF_buf46) );
  BUFX2 BUFX2_604 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3152_bF_buf45) );
  BUFX2 BUFX2_605 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3152_bF_buf44) );
  BUFX2 BUFX2_606 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3152_bF_buf43) );
  BUFX2 BUFX2_607 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3152_bF_buf42) );
  BUFX2 BUFX2_608 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3152_bF_buf41) );
  BUFX2 BUFX2_609 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3152_bF_buf40) );
  BUFX2 BUFX2_61 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf6) );
  BUFX2 BUFX2_610 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3152_bF_buf39) );
  BUFX2 BUFX2_611 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3152_bF_buf38) );
  BUFX2 BUFX2_612 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3152_bF_buf37) );
  BUFX2 BUFX2_613 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3152_bF_buf36) );
  BUFX2 BUFX2_614 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3152_bF_buf35) );
  BUFX2 BUFX2_615 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3152_bF_buf34) );
  BUFX2 BUFX2_616 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3152_bF_buf33) );
  BUFX2 BUFX2_617 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3152_bF_buf32) );
  BUFX2 BUFX2_618 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3152_bF_buf31) );
  BUFX2 BUFX2_619 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3152_bF_buf30) );
  BUFX2 BUFX2_62 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf5) );
  BUFX2 BUFX2_620 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3152_bF_buf29) );
  BUFX2 BUFX2_621 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3152_bF_buf28) );
  BUFX2 BUFX2_622 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3152_bF_buf27) );
  BUFX2 BUFX2_623 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3152_bF_buf26) );
  BUFX2 BUFX2_624 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3152_bF_buf25) );
  BUFX2 BUFX2_625 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3152_bF_buf24) );
  BUFX2 BUFX2_626 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3152_bF_buf23) );
  BUFX2 BUFX2_627 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3152_bF_buf22) );
  BUFX2 BUFX2_628 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3152_bF_buf21) );
  BUFX2 BUFX2_629 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3152_bF_buf20) );
  BUFX2 BUFX2_63 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf4) );
  BUFX2 BUFX2_630 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3152_bF_buf19) );
  BUFX2 BUFX2_631 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3152_bF_buf18) );
  BUFX2 BUFX2_632 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3152_bF_buf17) );
  BUFX2 BUFX2_633 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3152_bF_buf16) );
  BUFX2 BUFX2_634 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3152_bF_buf15) );
  BUFX2 BUFX2_635 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3152_bF_buf14) );
  BUFX2 BUFX2_636 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3152_bF_buf13) );
  BUFX2 BUFX2_637 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3152_bF_buf12) );
  BUFX2 BUFX2_638 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3152_bF_buf11) );
  BUFX2 BUFX2_639 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3152_bF_buf10) );
  BUFX2 BUFX2_64 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf3) );
  BUFX2 BUFX2_640 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3152_bF_buf9) );
  BUFX2 BUFX2_641 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3152_bF_buf8) );
  BUFX2 BUFX2_642 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf7), .Y(w_mem_inst__abc_21378_n3152_bF_buf7) );
  BUFX2 BUFX2_643 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf6), .Y(w_mem_inst__abc_21378_n3152_bF_buf6) );
  BUFX2 BUFX2_644 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf5), .Y(w_mem_inst__abc_21378_n3152_bF_buf5) );
  BUFX2 BUFX2_645 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf4), .Y(w_mem_inst__abc_21378_n3152_bF_buf4) );
  BUFX2 BUFX2_646 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf3), .Y(w_mem_inst__abc_21378_n3152_bF_buf3) );
  BUFX2 BUFX2_647 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf2), .Y(w_mem_inst__abc_21378_n3152_bF_buf2) );
  BUFX2 BUFX2_648 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf1), .Y(w_mem_inst__abc_21378_n3152_bF_buf1) );
  BUFX2 BUFX2_649 ( .A(w_mem_inst__abc_21378_n3152_hier0_bF_buf0), .Y(w_mem_inst__abc_21378_n3152_bF_buf0) );
  BUFX2 BUFX2_65 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf2) );
  BUFX2 BUFX2_650 ( .A(w_mem_inst__abc_21378_n3156), .Y(w_mem_inst__abc_21378_n3156_bF_buf4) );
  BUFX2 BUFX2_651 ( .A(w_mem_inst__abc_21378_n3156), .Y(w_mem_inst__abc_21378_n3156_bF_buf3) );
  BUFX2 BUFX2_652 ( .A(w_mem_inst__abc_21378_n3156), .Y(w_mem_inst__abc_21378_n3156_bF_buf2) );
  BUFX2 BUFX2_653 ( .A(w_mem_inst__abc_21378_n3156), .Y(w_mem_inst__abc_21378_n3156_bF_buf1) );
  BUFX2 BUFX2_654 ( .A(w_mem_inst__abc_21378_n3156), .Y(w_mem_inst__abc_21378_n3156_bF_buf0) );
  BUFX2 BUFX2_655 ( .A(w_mem_inst__abc_21378_n1625), .Y(w_mem_inst__abc_21378_n1625_bF_buf4) );
  BUFX2 BUFX2_656 ( .A(w_mem_inst__abc_21378_n1625), .Y(w_mem_inst__abc_21378_n1625_bF_buf3) );
  BUFX2 BUFX2_657 ( .A(w_mem_inst__abc_21378_n1625), .Y(w_mem_inst__abc_21378_n1625_bF_buf2) );
  BUFX2 BUFX2_658 ( .A(w_mem_inst__abc_21378_n1625), .Y(w_mem_inst__abc_21378_n1625_bF_buf1) );
  BUFX2 BUFX2_659 ( .A(w_mem_inst__abc_21378_n1625), .Y(w_mem_inst__abc_21378_n1625_bF_buf0) );
  BUFX2 BUFX2_66 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf1) );
  BUFX2 BUFX2_660 ( .A(w_mem_inst__abc_21378_n1634_1), .Y(w_mem_inst__abc_21378_n1634_1_bF_buf4) );
  BUFX2 BUFX2_661 ( .A(w_mem_inst__abc_21378_n1634_1), .Y(w_mem_inst__abc_21378_n1634_1_bF_buf3) );
  BUFX2 BUFX2_662 ( .A(w_mem_inst__abc_21378_n1634_1), .Y(w_mem_inst__abc_21378_n1634_1_bF_buf2) );
  BUFX2 BUFX2_663 ( .A(w_mem_inst__abc_21378_n1634_1), .Y(w_mem_inst__abc_21378_n1634_1_bF_buf1) );
  BUFX2 BUFX2_664 ( .A(w_mem_inst__abc_21378_n1634_1), .Y(w_mem_inst__abc_21378_n1634_1_bF_buf0) );
  BUFX2 BUFX2_665 ( .A(_abc_15724_n3721), .Y(_abc_15724_n3721_bF_buf4) );
  BUFX2 BUFX2_666 ( .A(_abc_15724_n3721), .Y(_abc_15724_n3721_bF_buf3) );
  BUFX2 BUFX2_667 ( .A(_abc_15724_n3721), .Y(_abc_15724_n3721_bF_buf2) );
  BUFX2 BUFX2_668 ( .A(_abc_15724_n3721), .Y(_abc_15724_n3721_bF_buf1) );
  BUFX2 BUFX2_669 ( .A(_abc_15724_n3721), .Y(_abc_15724_n3721_bF_buf0) );
  BUFX2 BUFX2_67 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf0) );
  BUFX2 BUFX2_670 ( .A(_abc_15724_n3725), .Y(_abc_15724_n3725_bF_buf3) );
  BUFX2 BUFX2_671 ( .A(_abc_15724_n3725), .Y(_abc_15724_n3725_bF_buf2) );
  BUFX2 BUFX2_672 ( .A(_abc_15724_n3725), .Y(_abc_15724_n3725_bF_buf1) );
  BUFX2 BUFX2_673 ( .A(_abc_15724_n3725), .Y(_abc_15724_n3725_bF_buf0) );
  BUFX2 BUFX2_674 ( .A(_abc_15724_n3726), .Y(_abc_15724_n3726_bF_buf4) );
  BUFX2 BUFX2_675 ( .A(_abc_15724_n3726), .Y(_abc_15724_n3726_bF_buf3) );
  BUFX2 BUFX2_676 ( .A(_abc_15724_n3726), .Y(_abc_15724_n3726_bF_buf2) );
  BUFX2 BUFX2_677 ( .A(_abc_15724_n3726), .Y(_abc_15724_n3726_bF_buf1) );
  BUFX2 BUFX2_678 ( .A(_abc_15724_n3726), .Y(_abc_15724_n3726_bF_buf0) );
  BUFX2 BUFX2_679 ( .A(_abc_15724_n906), .Y(_abc_15724_n906_bF_buf8) );
  BUFX2 BUFX2_68 ( .A(_abc_15724_n907_1), .Y(_abc_15724_n907_1_bF_buf7) );
  BUFX2 BUFX2_680 ( .A(_abc_15724_n906), .Y(_abc_15724_n906_bF_buf7) );
  BUFX2 BUFX2_681 ( .A(_abc_15724_n906), .Y(_abc_15724_n906_bF_buf6) );
  BUFX2 BUFX2_682 ( .A(_abc_15724_n906), .Y(_abc_15724_n906_bF_buf5) );
  BUFX2 BUFX2_683 ( .A(_abc_15724_n906), .Y(_abc_15724_n906_bF_buf4) );
  BUFX2 BUFX2_684 ( .A(_abc_15724_n906), .Y(_abc_15724_n906_bF_buf3) );
  BUFX2 BUFX2_685 ( .A(_abc_15724_n906), .Y(_abc_15724_n906_bF_buf2) );
  BUFX2 BUFX2_686 ( .A(_abc_15724_n906), .Y(_abc_15724_n906_bF_buf1) );
  BUFX2 BUFX2_687 ( .A(_abc_15724_n906), .Y(_abc_15724_n906_bF_buf0) );
  BUFX2 BUFX2_688 ( .A(_auto_iopadmap_cc_313_execute_26059_0_), .Y(\digest[0] ) );
  BUFX2 BUFX2_689 ( .A(_auto_iopadmap_cc_313_execute_26059_1_), .Y(\digest[1] ) );
  BUFX2 BUFX2_69 ( .A(_abc_15724_n907_1), .Y(_abc_15724_n907_1_bF_buf6) );
  BUFX2 BUFX2_690 ( .A(_auto_iopadmap_cc_313_execute_26059_2_), .Y(\digest[2] ) );
  BUFX2 BUFX2_691 ( .A(_auto_iopadmap_cc_313_execute_26059_3_), .Y(\digest[3] ) );
  BUFX2 BUFX2_692 ( .A(_auto_iopadmap_cc_313_execute_26059_4_), .Y(\digest[4] ) );
  BUFX2 BUFX2_693 ( .A(_auto_iopadmap_cc_313_execute_26059_5_), .Y(\digest[5] ) );
  BUFX2 BUFX2_694 ( .A(_auto_iopadmap_cc_313_execute_26059_6_), .Y(\digest[6] ) );
  BUFX2 BUFX2_695 ( .A(_auto_iopadmap_cc_313_execute_26059_7_), .Y(\digest[7] ) );
  BUFX2 BUFX2_696 ( .A(_auto_iopadmap_cc_313_execute_26059_8_), .Y(\digest[8] ) );
  BUFX2 BUFX2_697 ( .A(_auto_iopadmap_cc_313_execute_26059_9_), .Y(\digest[9] ) );
  BUFX2 BUFX2_698 ( .A(_auto_iopadmap_cc_313_execute_26059_10_), .Y(\digest[10] ) );
  BUFX2 BUFX2_699 ( .A(_auto_iopadmap_cc_313_execute_26059_11_), .Y(\digest[11] ) );
  BUFX2 BUFX2_7 ( .A(w_mem_inst__abc_21378_n3347_1), .Y(w_mem_inst__abc_21378_n3347_1_hier0_bF_buf0) );
  BUFX2 BUFX2_70 ( .A(_abc_15724_n907_1), .Y(_abc_15724_n907_1_bF_buf5) );
  BUFX2 BUFX2_700 ( .A(_auto_iopadmap_cc_313_execute_26059_12_), .Y(\digest[12] ) );
  BUFX2 BUFX2_701 ( .A(_auto_iopadmap_cc_313_execute_26059_13_), .Y(\digest[13] ) );
  BUFX2 BUFX2_702 ( .A(_auto_iopadmap_cc_313_execute_26059_14_), .Y(\digest[14] ) );
  BUFX2 BUFX2_703 ( .A(_auto_iopadmap_cc_313_execute_26059_15_), .Y(\digest[15] ) );
  BUFX2 BUFX2_704 ( .A(_auto_iopadmap_cc_313_execute_26059_16_), .Y(\digest[16] ) );
  BUFX2 BUFX2_705 ( .A(_auto_iopadmap_cc_313_execute_26059_17_), .Y(\digest[17] ) );
  BUFX2 BUFX2_706 ( .A(_auto_iopadmap_cc_313_execute_26059_18_), .Y(\digest[18] ) );
  BUFX2 BUFX2_707 ( .A(_auto_iopadmap_cc_313_execute_26059_19_), .Y(\digest[19] ) );
  BUFX2 BUFX2_708 ( .A(_auto_iopadmap_cc_313_execute_26059_20_), .Y(\digest[20] ) );
  BUFX2 BUFX2_709 ( .A(_auto_iopadmap_cc_313_execute_26059_21_), .Y(\digest[21] ) );
  BUFX2 BUFX2_71 ( .A(_abc_15724_n907_1), .Y(_abc_15724_n907_1_bF_buf4) );
  BUFX2 BUFX2_710 ( .A(_auto_iopadmap_cc_313_execute_26059_22_), .Y(\digest[22] ) );
  BUFX2 BUFX2_711 ( .A(_auto_iopadmap_cc_313_execute_26059_23_), .Y(\digest[23] ) );
  BUFX2 BUFX2_712 ( .A(_auto_iopadmap_cc_313_execute_26059_24_), .Y(\digest[24] ) );
  BUFX2 BUFX2_713 ( .A(_auto_iopadmap_cc_313_execute_26059_25_), .Y(\digest[25] ) );
  BUFX2 BUFX2_714 ( .A(_auto_iopadmap_cc_313_execute_26059_26_), .Y(\digest[26] ) );
  BUFX2 BUFX2_715 ( .A(_auto_iopadmap_cc_313_execute_26059_27_), .Y(\digest[27] ) );
  BUFX2 BUFX2_716 ( .A(_auto_iopadmap_cc_313_execute_26059_28_), .Y(\digest[28] ) );
  BUFX2 BUFX2_717 ( .A(_auto_iopadmap_cc_313_execute_26059_29_), .Y(\digest[29] ) );
  BUFX2 BUFX2_718 ( .A(_auto_iopadmap_cc_313_execute_26059_30_), .Y(\digest[30] ) );
  BUFX2 BUFX2_719 ( .A(_auto_iopadmap_cc_313_execute_26059_31_), .Y(\digest[31] ) );
  BUFX2 BUFX2_72 ( .A(_abc_15724_n907_1), .Y(_abc_15724_n907_1_bF_buf3) );
  BUFX2 BUFX2_720 ( .A(_auto_iopadmap_cc_313_execute_26059_32_), .Y(\digest[32] ) );
  BUFX2 BUFX2_721 ( .A(_auto_iopadmap_cc_313_execute_26059_33_), .Y(\digest[33] ) );
  BUFX2 BUFX2_722 ( .A(_auto_iopadmap_cc_313_execute_26059_34_), .Y(\digest[34] ) );
  BUFX2 BUFX2_723 ( .A(_auto_iopadmap_cc_313_execute_26059_35_), .Y(\digest[35] ) );
  BUFX2 BUFX2_724 ( .A(_auto_iopadmap_cc_313_execute_26059_36_), .Y(\digest[36] ) );
  BUFX2 BUFX2_725 ( .A(_auto_iopadmap_cc_313_execute_26059_37_), .Y(\digest[37] ) );
  BUFX2 BUFX2_726 ( .A(_auto_iopadmap_cc_313_execute_26059_38_), .Y(\digest[38] ) );
  BUFX2 BUFX2_727 ( .A(_auto_iopadmap_cc_313_execute_26059_39_), .Y(\digest[39] ) );
  BUFX2 BUFX2_728 ( .A(_auto_iopadmap_cc_313_execute_26059_40_), .Y(\digest[40] ) );
  BUFX2 BUFX2_729 ( .A(_auto_iopadmap_cc_313_execute_26059_41_), .Y(\digest[41] ) );
  BUFX2 BUFX2_73 ( .A(_abc_15724_n907_1), .Y(_abc_15724_n907_1_bF_buf2) );
  BUFX2 BUFX2_730 ( .A(_auto_iopadmap_cc_313_execute_26059_42_), .Y(\digest[42] ) );
  BUFX2 BUFX2_731 ( .A(_auto_iopadmap_cc_313_execute_26059_43_), .Y(\digest[43] ) );
  BUFX2 BUFX2_732 ( .A(_auto_iopadmap_cc_313_execute_26059_44_), .Y(\digest[44] ) );
  BUFX2 BUFX2_733 ( .A(_auto_iopadmap_cc_313_execute_26059_45_), .Y(\digest[45] ) );
  BUFX2 BUFX2_734 ( .A(_auto_iopadmap_cc_313_execute_26059_46_), .Y(\digest[46] ) );
  BUFX2 BUFX2_735 ( .A(_auto_iopadmap_cc_313_execute_26059_47_), .Y(\digest[47] ) );
  BUFX2 BUFX2_736 ( .A(_auto_iopadmap_cc_313_execute_26059_48_), .Y(\digest[48] ) );
  BUFX2 BUFX2_737 ( .A(_auto_iopadmap_cc_313_execute_26059_49_), .Y(\digest[49] ) );
  BUFX2 BUFX2_738 ( .A(_auto_iopadmap_cc_313_execute_26059_50_), .Y(\digest[50] ) );
  BUFX2 BUFX2_739 ( .A(_auto_iopadmap_cc_313_execute_26059_51_), .Y(\digest[51] ) );
  BUFX2 BUFX2_74 ( .A(_abc_15724_n907_1), .Y(_abc_15724_n907_1_bF_buf1) );
  BUFX2 BUFX2_740 ( .A(_auto_iopadmap_cc_313_execute_26059_52_), .Y(\digest[52] ) );
  BUFX2 BUFX2_741 ( .A(_auto_iopadmap_cc_313_execute_26059_53_), .Y(\digest[53] ) );
  BUFX2 BUFX2_742 ( .A(_auto_iopadmap_cc_313_execute_26059_54_), .Y(\digest[54] ) );
  BUFX2 BUFX2_743 ( .A(_auto_iopadmap_cc_313_execute_26059_55_), .Y(\digest[55] ) );
  BUFX2 BUFX2_744 ( .A(_auto_iopadmap_cc_313_execute_26059_56_), .Y(\digest[56] ) );
  BUFX2 BUFX2_745 ( .A(_auto_iopadmap_cc_313_execute_26059_57_), .Y(\digest[57] ) );
  BUFX2 BUFX2_746 ( .A(_auto_iopadmap_cc_313_execute_26059_58_), .Y(\digest[58] ) );
  BUFX2 BUFX2_747 ( .A(_auto_iopadmap_cc_313_execute_26059_59_), .Y(\digest[59] ) );
  BUFX2 BUFX2_748 ( .A(_auto_iopadmap_cc_313_execute_26059_60_), .Y(\digest[60] ) );
  BUFX2 BUFX2_749 ( .A(_auto_iopadmap_cc_313_execute_26059_61_), .Y(\digest[61] ) );
  BUFX2 BUFX2_75 ( .A(_abc_15724_n907_1), .Y(_abc_15724_n907_1_bF_buf0) );
  BUFX2 BUFX2_750 ( .A(_auto_iopadmap_cc_313_execute_26059_62_), .Y(\digest[62] ) );
  BUFX2 BUFX2_751 ( .A(_auto_iopadmap_cc_313_execute_26059_63_), .Y(\digest[63] ) );
  BUFX2 BUFX2_752 ( .A(_auto_iopadmap_cc_313_execute_26059_64_), .Y(\digest[64] ) );
  BUFX2 BUFX2_753 ( .A(_auto_iopadmap_cc_313_execute_26059_65_), .Y(\digest[65] ) );
  BUFX2 BUFX2_754 ( .A(_auto_iopadmap_cc_313_execute_26059_66_), .Y(\digest[66] ) );
  BUFX2 BUFX2_755 ( .A(_auto_iopadmap_cc_313_execute_26059_67_), .Y(\digest[67] ) );
  BUFX2 BUFX2_756 ( .A(_auto_iopadmap_cc_313_execute_26059_68_), .Y(\digest[68] ) );
  BUFX2 BUFX2_757 ( .A(_auto_iopadmap_cc_313_execute_26059_69_), .Y(\digest[69] ) );
  BUFX2 BUFX2_758 ( .A(_auto_iopadmap_cc_313_execute_26059_70_), .Y(\digest[70] ) );
  BUFX2 BUFX2_759 ( .A(_auto_iopadmap_cc_313_execute_26059_71_), .Y(\digest[71] ) );
  BUFX2 BUFX2_76 ( .A(_abc_15724_n3805), .Y(_abc_15724_n3805_bF_buf4) );
  BUFX2 BUFX2_760 ( .A(_auto_iopadmap_cc_313_execute_26059_72_), .Y(\digest[72] ) );
  BUFX2 BUFX2_761 ( .A(_auto_iopadmap_cc_313_execute_26059_73_), .Y(\digest[73] ) );
  BUFX2 BUFX2_762 ( .A(_auto_iopadmap_cc_313_execute_26059_74_), .Y(\digest[74] ) );
  BUFX2 BUFX2_763 ( .A(_auto_iopadmap_cc_313_execute_26059_75_), .Y(\digest[75] ) );
  BUFX2 BUFX2_764 ( .A(_auto_iopadmap_cc_313_execute_26059_76_), .Y(\digest[76] ) );
  BUFX2 BUFX2_765 ( .A(_auto_iopadmap_cc_313_execute_26059_77_), .Y(\digest[77] ) );
  BUFX2 BUFX2_766 ( .A(_auto_iopadmap_cc_313_execute_26059_78_), .Y(\digest[78] ) );
  BUFX2 BUFX2_767 ( .A(_auto_iopadmap_cc_313_execute_26059_79_), .Y(\digest[79] ) );
  BUFX2 BUFX2_768 ( .A(_auto_iopadmap_cc_313_execute_26059_80_), .Y(\digest[80] ) );
  BUFX2 BUFX2_769 ( .A(_auto_iopadmap_cc_313_execute_26059_81_), .Y(\digest[81] ) );
  BUFX2 BUFX2_77 ( .A(_abc_15724_n3805), .Y(_abc_15724_n3805_bF_buf3) );
  BUFX2 BUFX2_770 ( .A(_auto_iopadmap_cc_313_execute_26059_82_), .Y(\digest[82] ) );
  BUFX2 BUFX2_771 ( .A(_auto_iopadmap_cc_313_execute_26059_83_), .Y(\digest[83] ) );
  BUFX2 BUFX2_772 ( .A(_auto_iopadmap_cc_313_execute_26059_84_), .Y(\digest[84] ) );
  BUFX2 BUFX2_773 ( .A(_auto_iopadmap_cc_313_execute_26059_85_), .Y(\digest[85] ) );
  BUFX2 BUFX2_774 ( .A(_auto_iopadmap_cc_313_execute_26059_86_), .Y(\digest[86] ) );
  BUFX2 BUFX2_775 ( .A(_auto_iopadmap_cc_313_execute_26059_87_), .Y(\digest[87] ) );
  BUFX2 BUFX2_776 ( .A(_auto_iopadmap_cc_313_execute_26059_88_), .Y(\digest[88] ) );
  BUFX2 BUFX2_777 ( .A(_auto_iopadmap_cc_313_execute_26059_89_), .Y(\digest[89] ) );
  BUFX2 BUFX2_778 ( .A(_auto_iopadmap_cc_313_execute_26059_90_), .Y(\digest[90] ) );
  BUFX2 BUFX2_779 ( .A(_auto_iopadmap_cc_313_execute_26059_91_), .Y(\digest[91] ) );
  BUFX2 BUFX2_78 ( .A(_abc_15724_n3805), .Y(_abc_15724_n3805_bF_buf2) );
  BUFX2 BUFX2_780 ( .A(_auto_iopadmap_cc_313_execute_26059_92_), .Y(\digest[92] ) );
  BUFX2 BUFX2_781 ( .A(_auto_iopadmap_cc_313_execute_26059_93_), .Y(\digest[93] ) );
  BUFX2 BUFX2_782 ( .A(_auto_iopadmap_cc_313_execute_26059_94_), .Y(\digest[94] ) );
  BUFX2 BUFX2_783 ( .A(_auto_iopadmap_cc_313_execute_26059_95_), .Y(\digest[95] ) );
  BUFX2 BUFX2_784 ( .A(_auto_iopadmap_cc_313_execute_26059_96_), .Y(\digest[96] ) );
  BUFX2 BUFX2_785 ( .A(_auto_iopadmap_cc_313_execute_26059_97_), .Y(\digest[97] ) );
  BUFX2 BUFX2_786 ( .A(_auto_iopadmap_cc_313_execute_26059_98_), .Y(\digest[98] ) );
  BUFX2 BUFX2_787 ( .A(_auto_iopadmap_cc_313_execute_26059_99_), .Y(\digest[99] ) );
  BUFX2 BUFX2_788 ( .A(_auto_iopadmap_cc_313_execute_26059_100_), .Y(\digest[100] ) );
  BUFX2 BUFX2_789 ( .A(_auto_iopadmap_cc_313_execute_26059_101_), .Y(\digest[101] ) );
  BUFX2 BUFX2_79 ( .A(_abc_15724_n3805), .Y(_abc_15724_n3805_bF_buf1) );
  BUFX2 BUFX2_790 ( .A(_auto_iopadmap_cc_313_execute_26059_102_), .Y(\digest[102] ) );
  BUFX2 BUFX2_791 ( .A(_auto_iopadmap_cc_313_execute_26059_103_), .Y(\digest[103] ) );
  BUFX2 BUFX2_792 ( .A(_auto_iopadmap_cc_313_execute_26059_104_), .Y(\digest[104] ) );
  BUFX2 BUFX2_793 ( .A(_auto_iopadmap_cc_313_execute_26059_105_), .Y(\digest[105] ) );
  BUFX2 BUFX2_794 ( .A(_auto_iopadmap_cc_313_execute_26059_106_), .Y(\digest[106] ) );
  BUFX2 BUFX2_795 ( .A(_auto_iopadmap_cc_313_execute_26059_107_), .Y(\digest[107] ) );
  BUFX2 BUFX2_796 ( .A(_auto_iopadmap_cc_313_execute_26059_108_), .Y(\digest[108] ) );
  BUFX2 BUFX2_797 ( .A(_auto_iopadmap_cc_313_execute_26059_109_), .Y(\digest[109] ) );
  BUFX2 BUFX2_798 ( .A(_auto_iopadmap_cc_313_execute_26059_110_), .Y(\digest[110] ) );
  BUFX2 BUFX2_799 ( .A(_auto_iopadmap_cc_313_execute_26059_111_), .Y(\digest[111] ) );
  BUFX2 BUFX2_8 ( .A(clk), .Y(clk_hier0_bF_buf8) );
  BUFX2 BUFX2_80 ( .A(_abc_15724_n3805), .Y(_abc_15724_n3805_bF_buf0) );
  BUFX2 BUFX2_800 ( .A(_auto_iopadmap_cc_313_execute_26059_112_), .Y(\digest[112] ) );
  BUFX2 BUFX2_801 ( .A(_auto_iopadmap_cc_313_execute_26059_113_), .Y(\digest[113] ) );
  BUFX2 BUFX2_802 ( .A(_auto_iopadmap_cc_313_execute_26059_114_), .Y(\digest[114] ) );
  BUFX2 BUFX2_803 ( .A(_auto_iopadmap_cc_313_execute_26059_115_), .Y(\digest[115] ) );
  BUFX2 BUFX2_804 ( .A(_auto_iopadmap_cc_313_execute_26059_116_), .Y(\digest[116] ) );
  BUFX2 BUFX2_805 ( .A(_auto_iopadmap_cc_313_execute_26059_117_), .Y(\digest[117] ) );
  BUFX2 BUFX2_806 ( .A(_auto_iopadmap_cc_313_execute_26059_118_), .Y(\digest[118] ) );
  BUFX2 BUFX2_807 ( .A(_auto_iopadmap_cc_313_execute_26059_119_), .Y(\digest[119] ) );
  BUFX2 BUFX2_808 ( .A(_auto_iopadmap_cc_313_execute_26059_120_), .Y(\digest[120] ) );
  BUFX2 BUFX2_809 ( .A(_auto_iopadmap_cc_313_execute_26059_121_), .Y(\digest[121] ) );
  BUFX2 BUFX2_81 ( .A(_abc_15724_n3806), .Y(_abc_15724_n3806_bF_buf3) );
  BUFX2 BUFX2_810 ( .A(_auto_iopadmap_cc_313_execute_26059_122_), .Y(\digest[122] ) );
  BUFX2 BUFX2_811 ( .A(_auto_iopadmap_cc_313_execute_26059_123_), .Y(\digest[123] ) );
  BUFX2 BUFX2_812 ( .A(_auto_iopadmap_cc_313_execute_26059_124_), .Y(\digest[124] ) );
  BUFX2 BUFX2_813 ( .A(_auto_iopadmap_cc_313_execute_26059_125_), .Y(\digest[125] ) );
  BUFX2 BUFX2_814 ( .A(_auto_iopadmap_cc_313_execute_26059_126_), .Y(\digest[126] ) );
  BUFX2 BUFX2_815 ( .A(_auto_iopadmap_cc_313_execute_26059_127_), .Y(\digest[127] ) );
  BUFX2 BUFX2_816 ( .A(_auto_iopadmap_cc_313_execute_26059_128_), .Y(\digest[128] ) );
  BUFX2 BUFX2_817 ( .A(_auto_iopadmap_cc_313_execute_26059_129_), .Y(\digest[129] ) );
  BUFX2 BUFX2_818 ( .A(_auto_iopadmap_cc_313_execute_26059_130_), .Y(\digest[130] ) );
  BUFX2 BUFX2_819 ( .A(_auto_iopadmap_cc_313_execute_26059_131_), .Y(\digest[131] ) );
  BUFX2 BUFX2_82 ( .A(_abc_15724_n3806), .Y(_abc_15724_n3806_bF_buf2) );
  BUFX2 BUFX2_820 ( .A(_auto_iopadmap_cc_313_execute_26059_132_), .Y(\digest[132] ) );
  BUFX2 BUFX2_821 ( .A(_auto_iopadmap_cc_313_execute_26059_133_), .Y(\digest[133] ) );
  BUFX2 BUFX2_822 ( .A(_auto_iopadmap_cc_313_execute_26059_134_), .Y(\digest[134] ) );
  BUFX2 BUFX2_823 ( .A(_auto_iopadmap_cc_313_execute_26059_135_), .Y(\digest[135] ) );
  BUFX2 BUFX2_824 ( .A(_auto_iopadmap_cc_313_execute_26059_136_), .Y(\digest[136] ) );
  BUFX2 BUFX2_825 ( .A(_auto_iopadmap_cc_313_execute_26059_137_), .Y(\digest[137] ) );
  BUFX2 BUFX2_826 ( .A(_auto_iopadmap_cc_313_execute_26059_138_), .Y(\digest[138] ) );
  BUFX2 BUFX2_827 ( .A(_auto_iopadmap_cc_313_execute_26059_139_), .Y(\digest[139] ) );
  BUFX2 BUFX2_828 ( .A(_auto_iopadmap_cc_313_execute_26059_140_), .Y(\digest[140] ) );
  BUFX2 BUFX2_829 ( .A(_auto_iopadmap_cc_313_execute_26059_141_), .Y(\digest[141] ) );
  BUFX2 BUFX2_83 ( .A(_abc_15724_n3806), .Y(_abc_15724_n3806_bF_buf1) );
  BUFX2 BUFX2_830 ( .A(_auto_iopadmap_cc_313_execute_26059_142_), .Y(\digest[142] ) );
  BUFX2 BUFX2_831 ( .A(_auto_iopadmap_cc_313_execute_26059_143_), .Y(\digest[143] ) );
  BUFX2 BUFX2_832 ( .A(_auto_iopadmap_cc_313_execute_26059_144_), .Y(\digest[144] ) );
  BUFX2 BUFX2_833 ( .A(_auto_iopadmap_cc_313_execute_26059_145_), .Y(\digest[145] ) );
  BUFX2 BUFX2_834 ( .A(_auto_iopadmap_cc_313_execute_26059_146_), .Y(\digest[146] ) );
  BUFX2 BUFX2_835 ( .A(_auto_iopadmap_cc_313_execute_26059_147_), .Y(\digest[147] ) );
  BUFX2 BUFX2_836 ( .A(_auto_iopadmap_cc_313_execute_26059_148_), .Y(\digest[148] ) );
  BUFX2 BUFX2_837 ( .A(_auto_iopadmap_cc_313_execute_26059_149_), .Y(\digest[149] ) );
  BUFX2 BUFX2_838 ( .A(_auto_iopadmap_cc_313_execute_26059_150_), .Y(\digest[150] ) );
  BUFX2 BUFX2_839 ( .A(_auto_iopadmap_cc_313_execute_26059_151_), .Y(\digest[151] ) );
  BUFX2 BUFX2_84 ( .A(_abc_15724_n3806), .Y(_abc_15724_n3806_bF_buf0) );
  BUFX2 BUFX2_840 ( .A(_auto_iopadmap_cc_313_execute_26059_152_), .Y(\digest[152] ) );
  BUFX2 BUFX2_841 ( .A(_auto_iopadmap_cc_313_execute_26059_153_), .Y(\digest[153] ) );
  BUFX2 BUFX2_842 ( .A(_auto_iopadmap_cc_313_execute_26059_154_), .Y(\digest[154] ) );
  BUFX2 BUFX2_843 ( .A(_auto_iopadmap_cc_313_execute_26059_155_), .Y(\digest[155] ) );
  BUFX2 BUFX2_844 ( .A(_auto_iopadmap_cc_313_execute_26059_156_), .Y(\digest[156] ) );
  BUFX2 BUFX2_845 ( .A(_auto_iopadmap_cc_313_execute_26059_157_), .Y(\digest[157] ) );
  BUFX2 BUFX2_846 ( .A(_auto_iopadmap_cc_313_execute_26059_158_), .Y(\digest[158] ) );
  BUFX2 BUFX2_847 ( .A(_auto_iopadmap_cc_313_execute_26059_159_), .Y(\digest[159] ) );
  BUFX2 BUFX2_848 ( .A(_auto_iopadmap_cc_313_execute_26220), .Y(digest_valid) );
  BUFX2 BUFX2_849 ( .A(_auto_iopadmap_cc_313_execute_26222), .Y(ready) );
  BUFX2 BUFX2_85 ( .A(w_mem_inst__abc_21378_n1640), .Y(w_mem_inst__abc_21378_n1640_bF_buf4) );
  BUFX2 BUFX2_86 ( .A(w_mem_inst__abc_21378_n1640), .Y(w_mem_inst__abc_21378_n1640_bF_buf3) );
  BUFX2 BUFX2_87 ( .A(w_mem_inst__abc_21378_n1640), .Y(w_mem_inst__abc_21378_n1640_bF_buf2) );
  BUFX2 BUFX2_88 ( .A(w_mem_inst__abc_21378_n1640), .Y(w_mem_inst__abc_21378_n1640_bF_buf1) );
  BUFX2 BUFX2_89 ( .A(w_mem_inst__abc_21378_n1640), .Y(w_mem_inst__abc_21378_n1640_bF_buf0) );
  BUFX2 BUFX2_9 ( .A(clk), .Y(clk_hier0_bF_buf7) );
  BUFX2 BUFX2_90 ( .A(w_mem_inst__abc_21378_n1645), .Y(w_mem_inst__abc_21378_n1645_bF_buf4) );
  BUFX2 BUFX2_91 ( .A(w_mem_inst__abc_21378_n1645), .Y(w_mem_inst__abc_21378_n1645_bF_buf3) );
  BUFX2 BUFX2_92 ( .A(w_mem_inst__abc_21378_n1645), .Y(w_mem_inst__abc_21378_n1645_bF_buf2) );
  BUFX2 BUFX2_93 ( .A(w_mem_inst__abc_21378_n1645), .Y(w_mem_inst__abc_21378_n1645_bF_buf1) );
  BUFX2 BUFX2_94 ( .A(w_mem_inst__abc_21378_n1645), .Y(w_mem_inst__abc_21378_n1645_bF_buf0) );
  BUFX2 BUFX2_95 ( .A(w_mem_inst__abc_21378_n1649), .Y(w_mem_inst__abc_21378_n1649_bF_buf4) );
  BUFX2 BUFX2_96 ( .A(w_mem_inst__abc_21378_n1649), .Y(w_mem_inst__abc_21378_n1649_bF_buf3) );
  BUFX2 BUFX2_97 ( .A(w_mem_inst__abc_21378_n1649), .Y(w_mem_inst__abc_21378_n1649_bF_buf2) );
  BUFX2 BUFX2_98 ( .A(w_mem_inst__abc_21378_n1649), .Y(w_mem_inst__abc_21378_n1649_bF_buf1) );
  BUFX2 BUFX2_99 ( .A(w_mem_inst__abc_21378_n1649), .Y(w_mem_inst__abc_21378_n1649_bF_buf0) );
  DFFSR DFFSR_1 ( .CLK(clk_bF_buf88), .D(a_reg_0__FF_INPUT), .Q(a_reg_0_), .R(reset_n_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_10 ( .CLK(clk_bF_buf79), .D(a_reg_9__FF_INPUT), .Q(a_reg_9_), .R(reset_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_100 ( .CLK(clk_bF_buf78), .D(d_reg_3__FF_INPUT), .Q(d_reg_3_), .R(reset_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_101 ( .CLK(clk_bF_buf77), .D(d_reg_4__FF_INPUT), .Q(d_reg_4_), .R(reset_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_102 ( .CLK(clk_bF_buf76), .D(d_reg_5__FF_INPUT), .Q(d_reg_5_), .R(reset_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_103 ( .CLK(clk_bF_buf75), .D(d_reg_6__FF_INPUT), .Q(d_reg_6_), .R(reset_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_104 ( .CLK(clk_bF_buf74), .D(d_reg_7__FF_INPUT), .Q(d_reg_7_), .R(reset_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_105 ( .CLK(clk_bF_buf73), .D(d_reg_8__FF_INPUT), .Q(d_reg_8_), .R(reset_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_106 ( .CLK(clk_bF_buf72), .D(d_reg_9__FF_INPUT), .Q(d_reg_9_), .R(reset_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_107 ( .CLK(clk_bF_buf71), .D(d_reg_10__FF_INPUT), .Q(d_reg_10_), .R(reset_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_108 ( .CLK(clk_bF_buf70), .D(d_reg_11__FF_INPUT), .Q(d_reg_11_), .R(reset_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_109 ( .CLK(clk_bF_buf69), .D(d_reg_12__FF_INPUT), .Q(d_reg_12_), .R(reset_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_11 ( .CLK(clk_bF_buf78), .D(a_reg_10__FF_INPUT), .Q(a_reg_10_), .R(reset_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_110 ( .CLK(clk_bF_buf68), .D(d_reg_13__FF_INPUT), .Q(d_reg_13_), .R(reset_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_111 ( .CLK(clk_bF_buf67), .D(d_reg_14__FF_INPUT), .Q(d_reg_14_), .R(reset_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_112 ( .CLK(clk_bF_buf66), .D(d_reg_15__FF_INPUT), .Q(d_reg_15_), .R(reset_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_113 ( .CLK(clk_bF_buf65), .D(d_reg_16__FF_INPUT), .Q(d_reg_16_), .R(reset_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_114 ( .CLK(clk_bF_buf64), .D(d_reg_17__FF_INPUT), .Q(d_reg_17_), .R(reset_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_115 ( .CLK(clk_bF_buf63), .D(d_reg_18__FF_INPUT), .Q(d_reg_18_), .R(reset_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_116 ( .CLK(clk_bF_buf62), .D(d_reg_19__FF_INPUT), .Q(d_reg_19_), .R(reset_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_117 ( .CLK(clk_bF_buf61), .D(d_reg_20__FF_INPUT), .Q(d_reg_20_), .R(reset_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_118 ( .CLK(clk_bF_buf60), .D(d_reg_21__FF_INPUT), .Q(d_reg_21_), .R(reset_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_119 ( .CLK(clk_bF_buf59), .D(d_reg_22__FF_INPUT), .Q(d_reg_22_), .R(reset_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_12 ( .CLK(clk_bF_buf77), .D(a_reg_11__FF_INPUT), .Q(a_reg_11_), .R(reset_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_120 ( .CLK(clk_bF_buf58), .D(d_reg_23__FF_INPUT), .Q(d_reg_23_), .R(reset_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_121 ( .CLK(clk_bF_buf57), .D(d_reg_24__FF_INPUT), .Q(d_reg_24_), .R(reset_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_122 ( .CLK(clk_bF_buf56), .D(d_reg_25__FF_INPUT), .Q(d_reg_25_), .R(reset_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_123 ( .CLK(clk_bF_buf55), .D(d_reg_26__FF_INPUT), .Q(d_reg_26_), .R(reset_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_124 ( .CLK(clk_bF_buf54), .D(d_reg_27__FF_INPUT), .Q(d_reg_27_), .R(reset_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_125 ( .CLK(clk_bF_buf53), .D(d_reg_28__FF_INPUT), .Q(d_reg_28_), .R(reset_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_126 ( .CLK(clk_bF_buf52), .D(d_reg_29__FF_INPUT), .Q(d_reg_29_), .R(reset_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_127 ( .CLK(clk_bF_buf51), .D(d_reg_30__FF_INPUT), .Q(d_reg_30_), .R(reset_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_128 ( .CLK(clk_bF_buf50), .D(d_reg_31__FF_INPUT), .Q(d_reg_31_), .R(reset_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_129 ( .CLK(clk_bF_buf49), .D(e_reg_0__FF_INPUT), .Q(e_reg_0_), .R(reset_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_13 ( .CLK(clk_bF_buf76), .D(a_reg_12__FF_INPUT), .Q(a_reg_12_), .R(reset_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_130 ( .CLK(clk_bF_buf48), .D(e_reg_1__FF_INPUT), .Q(e_reg_1_), .R(reset_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_131 ( .CLK(clk_bF_buf47), .D(e_reg_2__FF_INPUT), .Q(e_reg_2_), .R(reset_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_132 ( .CLK(clk_bF_buf46), .D(e_reg_3__FF_INPUT), .Q(e_reg_3_), .R(reset_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_133 ( .CLK(clk_bF_buf45), .D(e_reg_4__FF_INPUT), .Q(e_reg_4_), .R(reset_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_134 ( .CLK(clk_bF_buf44), .D(e_reg_5__FF_INPUT), .Q(e_reg_5_), .R(reset_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_135 ( .CLK(clk_bF_buf43), .D(e_reg_6__FF_INPUT), .Q(e_reg_6_), .R(reset_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_136 ( .CLK(clk_bF_buf42), .D(e_reg_7__FF_INPUT), .Q(e_reg_7_), .R(reset_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_137 ( .CLK(clk_bF_buf41), .D(e_reg_8__FF_INPUT), .Q(e_reg_8_), .R(reset_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_138 ( .CLK(clk_bF_buf40), .D(e_reg_9__FF_INPUT), .Q(e_reg_9_), .R(reset_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_139 ( .CLK(clk_bF_buf39), .D(e_reg_10__FF_INPUT), .Q(e_reg_10_), .R(reset_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_14 ( .CLK(clk_bF_buf75), .D(a_reg_13__FF_INPUT), .Q(a_reg_13_), .R(reset_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_140 ( .CLK(clk_bF_buf38), .D(e_reg_11__FF_INPUT), .Q(e_reg_11_), .R(reset_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_141 ( .CLK(clk_bF_buf37), .D(e_reg_12__FF_INPUT), .Q(e_reg_12_), .R(reset_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_142 ( .CLK(clk_bF_buf36), .D(e_reg_13__FF_INPUT), .Q(e_reg_13_), .R(reset_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_143 ( .CLK(clk_bF_buf35), .D(e_reg_14__FF_INPUT), .Q(e_reg_14_), .R(reset_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_144 ( .CLK(clk_bF_buf34), .D(e_reg_15__FF_INPUT), .Q(e_reg_15_), .R(reset_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_145 ( .CLK(clk_bF_buf33), .D(e_reg_16__FF_INPUT), .Q(e_reg_16_), .R(reset_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_146 ( .CLK(clk_bF_buf32), .D(e_reg_17__FF_INPUT), .Q(e_reg_17_), .R(reset_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_147 ( .CLK(clk_bF_buf31), .D(e_reg_18__FF_INPUT), .Q(e_reg_18_), .R(reset_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_148 ( .CLK(clk_bF_buf30), .D(e_reg_19__FF_INPUT), .Q(e_reg_19_), .R(reset_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_149 ( .CLK(clk_bF_buf29), .D(e_reg_20__FF_INPUT), .Q(e_reg_20_), .R(reset_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_15 ( .CLK(clk_bF_buf74), .D(a_reg_14__FF_INPUT), .Q(a_reg_14_), .R(reset_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_150 ( .CLK(clk_bF_buf28), .D(e_reg_21__FF_INPUT), .Q(e_reg_21_), .R(reset_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_151 ( .CLK(clk_bF_buf27), .D(e_reg_22__FF_INPUT), .Q(e_reg_22_), .R(reset_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_152 ( .CLK(clk_bF_buf26), .D(e_reg_23__FF_INPUT), .Q(e_reg_23_), .R(reset_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_153 ( .CLK(clk_bF_buf25), .D(e_reg_24__FF_INPUT), .Q(e_reg_24_), .R(reset_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_154 ( .CLK(clk_bF_buf24), .D(e_reg_25__FF_INPUT), .Q(e_reg_25_), .R(reset_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_155 ( .CLK(clk_bF_buf23), .D(e_reg_26__FF_INPUT), .Q(e_reg_26_), .R(reset_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_156 ( .CLK(clk_bF_buf22), .D(e_reg_27__FF_INPUT), .Q(e_reg_27_), .R(reset_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_157 ( .CLK(clk_bF_buf21), .D(e_reg_28__FF_INPUT), .Q(e_reg_28_), .R(reset_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_158 ( .CLK(clk_bF_buf20), .D(e_reg_29__FF_INPUT), .Q(e_reg_29_), .R(reset_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_159 ( .CLK(clk_bF_buf19), .D(e_reg_30__FF_INPUT), .Q(e_reg_30_), .R(reset_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_16 ( .CLK(clk_bF_buf73), .D(a_reg_15__FF_INPUT), .Q(a_reg_15_), .R(reset_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_160 ( .CLK(clk_bF_buf18), .D(e_reg_31__FF_INPUT), .Q(e_reg_31_), .R(reset_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_161 ( .CLK(clk_bF_buf17), .D(H0_reg_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_128_), .R(reset_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_162 ( .CLK(clk_bF_buf16), .D(H0_reg_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_129_), .R(reset_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_163 ( .CLK(clk_bF_buf15), .D(H0_reg_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_130_), .R(reset_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_164 ( .CLK(clk_bF_buf14), .D(H0_reg_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_131_), .R(reset_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_165 ( .CLK(clk_bF_buf13), .D(H0_reg_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_132_), .R(reset_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_166 ( .CLK(clk_bF_buf12), .D(H0_reg_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_133_), .R(reset_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_167 ( .CLK(clk_bF_buf11), .D(H0_reg_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_134_), .R(reset_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_168 ( .CLK(clk_bF_buf10), .D(H0_reg_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_135_), .R(reset_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_169 ( .CLK(clk_bF_buf9), .D(H0_reg_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_136_), .R(reset_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_17 ( .CLK(clk_bF_buf72), .D(a_reg_16__FF_INPUT), .Q(a_reg_16_), .R(reset_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_170 ( .CLK(clk_bF_buf8), .D(H0_reg_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_137_), .R(reset_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_171 ( .CLK(clk_bF_buf7), .D(H0_reg_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_138_), .R(reset_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_172 ( .CLK(clk_bF_buf6), .D(H0_reg_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_139_), .R(reset_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_173 ( .CLK(clk_bF_buf5), .D(H0_reg_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_140_), .R(reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_174 ( .CLK(clk_bF_buf4), .D(H0_reg_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_141_), .R(reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_175 ( .CLK(clk_bF_buf3), .D(H0_reg_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_142_), .R(reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_176 ( .CLK(clk_bF_buf2), .D(H0_reg_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_143_), .R(reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_177 ( .CLK(clk_bF_buf1), .D(H0_reg_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_144_), .R(reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_178 ( .CLK(clk_bF_buf0), .D(H0_reg_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_145_), .R(reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_179 ( .CLK(clk_bF_buf88), .D(H0_reg_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_146_), .R(reset_n_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_18 ( .CLK(clk_bF_buf71), .D(a_reg_17__FF_INPUT), .Q(a_reg_17_), .R(reset_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_180 ( .CLK(clk_bF_buf87), .D(H0_reg_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_147_), .R(reset_n_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_181 ( .CLK(clk_bF_buf86), .D(H0_reg_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_148_), .R(reset_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_182 ( .CLK(clk_bF_buf85), .D(H0_reg_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_149_), .R(reset_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_183 ( .CLK(clk_bF_buf84), .D(H0_reg_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_150_), .R(reset_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_184 ( .CLK(clk_bF_buf83), .D(H0_reg_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_151_), .R(reset_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_185 ( .CLK(clk_bF_buf82), .D(H0_reg_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_152_), .R(reset_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_186 ( .CLK(clk_bF_buf81), .D(H0_reg_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_153_), .R(reset_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_187 ( .CLK(clk_bF_buf80), .D(H0_reg_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_154_), .R(reset_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_188 ( .CLK(clk_bF_buf79), .D(H0_reg_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_155_), .R(reset_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_189 ( .CLK(clk_bF_buf78), .D(H0_reg_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_156_), .R(reset_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_19 ( .CLK(clk_bF_buf70), .D(a_reg_18__FF_INPUT), .Q(a_reg_18_), .R(reset_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_190 ( .CLK(clk_bF_buf77), .D(H0_reg_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_157_), .R(reset_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_191 ( .CLK(clk_bF_buf76), .D(H0_reg_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_158_), .R(reset_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_192 ( .CLK(clk_bF_buf75), .D(H0_reg_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_159_), .R(reset_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_193 ( .CLK(clk_bF_buf74), .D(H1_reg_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_96_), .R(reset_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_194 ( .CLK(clk_bF_buf73), .D(H1_reg_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_97_), .R(reset_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_195 ( .CLK(clk_bF_buf72), .D(H1_reg_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_98_), .R(reset_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_196 ( .CLK(clk_bF_buf71), .D(H1_reg_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_99_), .R(reset_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_197 ( .CLK(clk_bF_buf70), .D(H1_reg_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_100_), .R(reset_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_198 ( .CLK(clk_bF_buf69), .D(H1_reg_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_101_), .R(reset_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_199 ( .CLK(clk_bF_buf68), .D(H1_reg_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_102_), .R(reset_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_2 ( .CLK(clk_bF_buf87), .D(a_reg_1__FF_INPUT), .Q(a_reg_1_), .R(reset_n_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_20 ( .CLK(clk_bF_buf69), .D(a_reg_19__FF_INPUT), .Q(a_reg_19_), .R(reset_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_200 ( .CLK(clk_bF_buf67), .D(H1_reg_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_103_), .R(reset_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_201 ( .CLK(clk_bF_buf66), .D(H1_reg_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_104_), .R(reset_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_202 ( .CLK(clk_bF_buf65), .D(H1_reg_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_105_), .R(reset_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_203 ( .CLK(clk_bF_buf64), .D(H1_reg_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_106_), .R(reset_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_204 ( .CLK(clk_bF_buf63), .D(H1_reg_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_107_), .R(reset_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_205 ( .CLK(clk_bF_buf62), .D(H1_reg_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_108_), .R(reset_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_206 ( .CLK(clk_bF_buf61), .D(H1_reg_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_109_), .R(reset_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_207 ( .CLK(clk_bF_buf60), .D(H1_reg_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_110_), .R(reset_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_208 ( .CLK(clk_bF_buf59), .D(H1_reg_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_111_), .R(reset_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_209 ( .CLK(clk_bF_buf58), .D(H1_reg_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_112_), .R(reset_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_21 ( .CLK(clk_bF_buf68), .D(a_reg_20__FF_INPUT), .Q(a_reg_20_), .R(reset_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_210 ( .CLK(clk_bF_buf57), .D(H1_reg_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_113_), .R(reset_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_211 ( .CLK(clk_bF_buf56), .D(H1_reg_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_114_), .R(reset_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_212 ( .CLK(clk_bF_buf55), .D(H1_reg_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_115_), .R(reset_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_213 ( .CLK(clk_bF_buf54), .D(H1_reg_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_116_), .R(reset_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_214 ( .CLK(clk_bF_buf53), .D(H1_reg_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_117_), .R(reset_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_215 ( .CLK(clk_bF_buf52), .D(H1_reg_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_118_), .R(reset_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_216 ( .CLK(clk_bF_buf51), .D(H1_reg_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_119_), .R(reset_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_217 ( .CLK(clk_bF_buf50), .D(H1_reg_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_120_), .R(reset_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_218 ( .CLK(clk_bF_buf49), .D(H1_reg_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_121_), .R(reset_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_219 ( .CLK(clk_bF_buf48), .D(H1_reg_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_122_), .R(reset_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_22 ( .CLK(clk_bF_buf67), .D(a_reg_21__FF_INPUT), .Q(a_reg_21_), .R(reset_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_220 ( .CLK(clk_bF_buf47), .D(H1_reg_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_123_), .R(reset_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_221 ( .CLK(clk_bF_buf46), .D(H1_reg_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_124_), .R(reset_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_222 ( .CLK(clk_bF_buf45), .D(H1_reg_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_125_), .R(reset_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_223 ( .CLK(clk_bF_buf44), .D(H1_reg_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_126_), .R(reset_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_224 ( .CLK(clk_bF_buf43), .D(H1_reg_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_127_), .R(reset_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_225 ( .CLK(clk_bF_buf42), .D(H2_reg_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_64_), .R(reset_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_226 ( .CLK(clk_bF_buf41), .D(H2_reg_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_65_), .R(reset_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_227 ( .CLK(clk_bF_buf40), .D(H2_reg_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_66_), .R(reset_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_228 ( .CLK(clk_bF_buf39), .D(H2_reg_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_67_), .R(reset_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_229 ( .CLK(clk_bF_buf38), .D(H2_reg_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_68_), .R(reset_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_23 ( .CLK(clk_bF_buf66), .D(a_reg_22__FF_INPUT), .Q(a_reg_22_), .R(reset_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_230 ( .CLK(clk_bF_buf37), .D(H2_reg_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_69_), .R(reset_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_231 ( .CLK(clk_bF_buf36), .D(H2_reg_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_70_), .R(reset_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_232 ( .CLK(clk_bF_buf35), .D(H2_reg_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_71_), .R(reset_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_233 ( .CLK(clk_bF_buf34), .D(H2_reg_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_72_), .R(reset_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_234 ( .CLK(clk_bF_buf33), .D(H2_reg_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_73_), .R(reset_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_235 ( .CLK(clk_bF_buf32), .D(H2_reg_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_74_), .R(reset_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_236 ( .CLK(clk_bF_buf31), .D(H2_reg_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_75_), .R(reset_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_237 ( .CLK(clk_bF_buf30), .D(H2_reg_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_76_), .R(reset_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_238 ( .CLK(clk_bF_buf29), .D(H2_reg_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_77_), .R(reset_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_239 ( .CLK(clk_bF_buf28), .D(H2_reg_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_78_), .R(reset_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_24 ( .CLK(clk_bF_buf65), .D(a_reg_23__FF_INPUT), .Q(a_reg_23_), .R(reset_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_240 ( .CLK(clk_bF_buf27), .D(H2_reg_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_79_), .R(reset_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_241 ( .CLK(clk_bF_buf26), .D(H2_reg_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_80_), .R(reset_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_242 ( .CLK(clk_bF_buf25), .D(H2_reg_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_81_), .R(reset_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_243 ( .CLK(clk_bF_buf24), .D(H2_reg_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_82_), .R(reset_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_244 ( .CLK(clk_bF_buf23), .D(H2_reg_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_83_), .R(reset_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_245 ( .CLK(clk_bF_buf22), .D(H2_reg_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_84_), .R(reset_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_246 ( .CLK(clk_bF_buf21), .D(H2_reg_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_85_), .R(reset_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_247 ( .CLK(clk_bF_buf20), .D(H2_reg_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_86_), .R(reset_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_248 ( .CLK(clk_bF_buf19), .D(H2_reg_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_87_), .R(reset_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_249 ( .CLK(clk_bF_buf18), .D(H2_reg_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_88_), .R(reset_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_25 ( .CLK(clk_bF_buf64), .D(a_reg_24__FF_INPUT), .Q(a_reg_24_), .R(reset_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_250 ( .CLK(clk_bF_buf17), .D(H2_reg_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_89_), .R(reset_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_251 ( .CLK(clk_bF_buf16), .D(H2_reg_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_90_), .R(reset_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_252 ( .CLK(clk_bF_buf15), .D(H2_reg_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_91_), .R(reset_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_253 ( .CLK(clk_bF_buf14), .D(H2_reg_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_92_), .R(reset_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_254 ( .CLK(clk_bF_buf13), .D(H2_reg_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_93_), .R(reset_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_255 ( .CLK(clk_bF_buf12), .D(H2_reg_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_94_), .R(reset_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_256 ( .CLK(clk_bF_buf11), .D(H2_reg_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_95_), .R(reset_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_257 ( .CLK(clk_bF_buf10), .D(H3_reg_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_32_), .R(reset_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_258 ( .CLK(clk_bF_buf9), .D(H3_reg_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_33_), .R(reset_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_259 ( .CLK(clk_bF_buf8), .D(H3_reg_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_34_), .R(reset_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_26 ( .CLK(clk_bF_buf63), .D(a_reg_25__FF_INPUT), .Q(a_reg_25_), .R(reset_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_260 ( .CLK(clk_bF_buf7), .D(H3_reg_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_35_), .R(reset_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_261 ( .CLK(clk_bF_buf6), .D(H3_reg_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_36_), .R(reset_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_262 ( .CLK(clk_bF_buf5), .D(H3_reg_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_37_), .R(reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_263 ( .CLK(clk_bF_buf4), .D(H3_reg_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_38_), .R(reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_264 ( .CLK(clk_bF_buf3), .D(H3_reg_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_39_), .R(reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_265 ( .CLK(clk_bF_buf2), .D(H3_reg_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_40_), .R(reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_266 ( .CLK(clk_bF_buf1), .D(H3_reg_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_41_), .R(reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_267 ( .CLK(clk_bF_buf0), .D(H3_reg_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_42_), .R(reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_268 ( .CLK(clk_bF_buf88), .D(H3_reg_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_43_), .R(reset_n_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_269 ( .CLK(clk_bF_buf87), .D(H3_reg_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_44_), .R(reset_n_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_27 ( .CLK(clk_bF_buf62), .D(a_reg_26__FF_INPUT), .Q(a_reg_26_), .R(reset_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_270 ( .CLK(clk_bF_buf86), .D(H3_reg_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_45_), .R(reset_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_271 ( .CLK(clk_bF_buf85), .D(H3_reg_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_46_), .R(reset_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_272 ( .CLK(clk_bF_buf84), .D(H3_reg_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_47_), .R(reset_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_273 ( .CLK(clk_bF_buf83), .D(H3_reg_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_48_), .R(reset_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_274 ( .CLK(clk_bF_buf82), .D(H3_reg_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_49_), .R(reset_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_275 ( .CLK(clk_bF_buf81), .D(H3_reg_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_50_), .R(reset_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_276 ( .CLK(clk_bF_buf80), .D(H3_reg_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_51_), .R(reset_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_277 ( .CLK(clk_bF_buf79), .D(H3_reg_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_52_), .R(reset_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_278 ( .CLK(clk_bF_buf78), .D(H3_reg_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_53_), .R(reset_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_279 ( .CLK(clk_bF_buf77), .D(H3_reg_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_54_), .R(reset_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_28 ( .CLK(clk_bF_buf61), .D(a_reg_27__FF_INPUT), .Q(a_reg_27_), .R(reset_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_280 ( .CLK(clk_bF_buf76), .D(H3_reg_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_55_), .R(reset_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_281 ( .CLK(clk_bF_buf75), .D(H3_reg_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_56_), .R(reset_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_282 ( .CLK(clk_bF_buf74), .D(H3_reg_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_57_), .R(reset_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_283 ( .CLK(clk_bF_buf73), .D(H3_reg_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_58_), .R(reset_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_284 ( .CLK(clk_bF_buf72), .D(H3_reg_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_59_), .R(reset_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_285 ( .CLK(clk_bF_buf71), .D(H3_reg_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_60_), .R(reset_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_286 ( .CLK(clk_bF_buf70), .D(H3_reg_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_61_), .R(reset_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_287 ( .CLK(clk_bF_buf69), .D(H3_reg_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_62_), .R(reset_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_288 ( .CLK(clk_bF_buf68), .D(H3_reg_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_63_), .R(reset_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_289 ( .CLK(clk_bF_buf67), .D(H4_reg_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_0_), .R(reset_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_29 ( .CLK(clk_bF_buf60), .D(a_reg_28__FF_INPUT), .Q(a_reg_28_), .R(reset_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_290 ( .CLK(clk_bF_buf66), .D(H4_reg_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_1_), .R(reset_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_291 ( .CLK(clk_bF_buf65), .D(H4_reg_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_2_), .R(reset_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_292 ( .CLK(clk_bF_buf64), .D(H4_reg_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_3_), .R(reset_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_293 ( .CLK(clk_bF_buf63), .D(H4_reg_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_4_), .R(reset_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_294 ( .CLK(clk_bF_buf62), .D(H4_reg_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_5_), .R(reset_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_295 ( .CLK(clk_bF_buf61), .D(H4_reg_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_6_), .R(reset_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_296 ( .CLK(clk_bF_buf60), .D(H4_reg_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_7_), .R(reset_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_297 ( .CLK(clk_bF_buf59), .D(H4_reg_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_8_), .R(reset_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_298 ( .CLK(clk_bF_buf58), .D(H4_reg_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_9_), .R(reset_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_299 ( .CLK(clk_bF_buf57), .D(H4_reg_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_10_), .R(reset_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_3 ( .CLK(clk_bF_buf86), .D(a_reg_2__FF_INPUT), .Q(a_reg_2_), .R(reset_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_30 ( .CLK(clk_bF_buf59), .D(a_reg_29__FF_INPUT), .Q(a_reg_29_), .R(reset_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_300 ( .CLK(clk_bF_buf56), .D(H4_reg_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_11_), .R(reset_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_301 ( .CLK(clk_bF_buf55), .D(H4_reg_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_12_), .R(reset_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_302 ( .CLK(clk_bF_buf54), .D(H4_reg_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_13_), .R(reset_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_303 ( .CLK(clk_bF_buf53), .D(H4_reg_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_14_), .R(reset_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_304 ( .CLK(clk_bF_buf52), .D(H4_reg_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_15_), .R(reset_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_305 ( .CLK(clk_bF_buf51), .D(H4_reg_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_16_), .R(reset_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_306 ( .CLK(clk_bF_buf50), .D(H4_reg_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_17_), .R(reset_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_307 ( .CLK(clk_bF_buf49), .D(H4_reg_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_18_), .R(reset_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_308 ( .CLK(clk_bF_buf48), .D(H4_reg_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_19_), .R(reset_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_309 ( .CLK(clk_bF_buf47), .D(H4_reg_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_20_), .R(reset_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_31 ( .CLK(clk_bF_buf58), .D(a_reg_30__FF_INPUT), .Q(a_reg_30_), .R(reset_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_310 ( .CLK(clk_bF_buf46), .D(H4_reg_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_21_), .R(reset_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_311 ( .CLK(clk_bF_buf45), .D(H4_reg_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_22_), .R(reset_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_312 ( .CLK(clk_bF_buf44), .D(H4_reg_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_23_), .R(reset_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_313 ( .CLK(clk_bF_buf43), .D(H4_reg_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_24_), .R(reset_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_314 ( .CLK(clk_bF_buf42), .D(H4_reg_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_25_), .R(reset_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_315 ( .CLK(clk_bF_buf41), .D(H4_reg_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_26_), .R(reset_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_316 ( .CLK(clk_bF_buf40), .D(H4_reg_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_27_), .R(reset_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_317 ( .CLK(clk_bF_buf39), .D(H4_reg_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_28_), .R(reset_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_318 ( .CLK(clk_bF_buf38), .D(H4_reg_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_29_), .R(reset_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_319 ( .CLK(clk_bF_buf37), .D(H4_reg_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_30_), .R(reset_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_32 ( .CLK(clk_bF_buf57), .D(a_reg_31__FF_INPUT), .Q(a_reg_31_), .R(reset_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_320 ( .CLK(clk_bF_buf36), .D(H4_reg_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26059_31_), .R(reset_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_321 ( .CLK(clk_bF_buf35), .D(round_ctr_reg_0__FF_INPUT), .Q(round_ctr_reg_0_), .R(reset_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_322 ( .CLK(clk_bF_buf34), .D(round_ctr_reg_1__FF_INPUT), .Q(round_ctr_reg_1_), .R(reset_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_323 ( .CLK(clk_bF_buf33), .D(round_ctr_reg_2__FF_INPUT), .Q(round_ctr_reg_2_), .R(reset_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_324 ( .CLK(clk_bF_buf32), .D(round_ctr_reg_3__FF_INPUT), .Q(round_ctr_reg_3_), .R(reset_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_325 ( .CLK(clk_bF_buf31), .D(round_ctr_reg_4__FF_INPUT), .Q(round_ctr_reg_4_), .R(reset_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_326 ( .CLK(clk_bF_buf30), .D(round_ctr_reg_5__FF_INPUT), .Q(round_ctr_reg_5_), .R(reset_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_327 ( .CLK(clk_bF_buf29), .D(round_ctr_reg_6__FF_INPUT), .Q(round_ctr_reg_6_), .R(reset_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_328 ( .CLK(clk_bF_buf28), .D(digest_valid_reg_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_26220), .R(reset_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_329 ( .CLK(clk_bF_buf27), .D(_abc_15724_n3489), .Q(_auto_iopadmap_cc_313_execute_26222), .R(1'b1), .S(reset_n_bF_buf27) );
  DFFSR DFFSR_33 ( .CLK(clk_bF_buf56), .D(b_reg_0__FF_INPUT), .Q(b_reg_0_), .R(reset_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_330 ( .CLK(clk_bF_buf26), .D(_abc_15724_n3465), .Q(digest_update), .R(reset_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_331 ( .CLK(clk_bF_buf25), .D(_abc_15724_n3483), .Q(round_ctr_inc), .R(reset_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_332 ( .CLK(clk_bF_buf24), .D(w_mem_inst_w_ctr_reg_0__FF_INPUT), .Q(w_mem_inst_w_ctr_reg_0_), .R(reset_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_333 ( .CLK(clk_bF_buf23), .D(w_mem_inst_w_ctr_reg_1__FF_INPUT), .Q(w_mem_inst_w_ctr_reg_1_), .R(reset_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_334 ( .CLK(clk_bF_buf22), .D(w_mem_inst_w_ctr_reg_2__FF_INPUT), .Q(w_mem_inst_w_ctr_reg_2_), .R(reset_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_335 ( .CLK(clk_bF_buf21), .D(w_mem_inst_w_ctr_reg_3__FF_INPUT), .Q(w_mem_inst_w_ctr_reg_3_), .R(reset_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_336 ( .CLK(clk_bF_buf20), .D(w_mem_inst_w_ctr_reg_4__FF_INPUT), .Q(w_mem_inst_w_ctr_reg_4_), .R(reset_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_337 ( .CLK(clk_bF_buf19), .D(w_mem_inst_w_ctr_reg_5__FF_INPUT), .Q(w_mem_inst_w_ctr_reg_5_), .R(reset_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_338 ( .CLK(clk_bF_buf18), .D(w_mem_inst_w_ctr_reg_6__FF_INPUT), .Q(w_mem_inst_w_ctr_reg_6_), .R(reset_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_339 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_0__31_0__0_), .Q(w_mem_inst_w_mem_0__0_), .R(reset_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_34 ( .CLK(clk_bF_buf55), .D(b_reg_1__FF_INPUT), .Q(b_reg_1_), .R(reset_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_340 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_0__31_0__1_), .Q(w_mem_inst_w_mem_0__1_), .R(reset_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_341 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_0__31_0__2_), .Q(w_mem_inst_w_mem_0__2_), .R(reset_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_342 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_0__31_0__3_), .Q(w_mem_inst_w_mem_0__3_), .R(reset_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_343 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_0__31_0__4_), .Q(w_mem_inst_w_mem_0__4_), .R(reset_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_344 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_0__31_0__5_), .Q(w_mem_inst_w_mem_0__5_), .R(reset_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_345 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_0__31_0__6_), .Q(w_mem_inst_w_mem_0__6_), .R(reset_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_346 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_0__31_0__7_), .Q(w_mem_inst_w_mem_0__7_), .R(reset_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_347 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_0__31_0__8_), .Q(w_mem_inst_w_mem_0__8_), .R(reset_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_348 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_0__31_0__9_), .Q(w_mem_inst_w_mem_0__9_), .R(reset_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_349 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_0__31_0__10_), .Q(w_mem_inst_w_mem_0__10_), .R(reset_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_35 ( .CLK(clk_bF_buf54), .D(b_reg_2__FF_INPUT), .Q(b_reg_2_), .R(reset_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_350 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_0__31_0__11_), .Q(w_mem_inst_w_mem_0__11_), .R(reset_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_351 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_0__31_0__12_), .Q(w_mem_inst_w_mem_0__12_), .R(reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_352 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_0__31_0__13_), .Q(w_mem_inst_w_mem_0__13_), .R(reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_353 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_0__31_0__14_), .Q(w_mem_inst_w_mem_0__14_), .R(reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_354 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_0__31_0__15_), .Q(w_mem_inst_w_mem_0__15_), .R(reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_355 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_0__31_0__16_), .Q(w_mem_inst_w_mem_0__16_), .R(reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_356 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_0__31_0__17_), .Q(w_mem_inst_w_mem_0__17_), .R(reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_357 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_0__31_0__18_), .Q(w_mem_inst_w_mem_0__18_), .R(reset_n_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_358 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_0__31_0__19_), .Q(w_mem_inst_w_mem_0__19_), .R(reset_n_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_359 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_0__31_0__20_), .Q(w_mem_inst_w_mem_0__20_), .R(reset_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_36 ( .CLK(clk_bF_buf53), .D(b_reg_3__FF_INPUT), .Q(b_reg_3_), .R(reset_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_360 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_0__31_0__21_), .Q(w_mem_inst_w_mem_0__21_), .R(reset_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_361 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_0__31_0__22_), .Q(w_mem_inst_w_mem_0__22_), .R(reset_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_362 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_0__31_0__23_), .Q(w_mem_inst_w_mem_0__23_), .R(reset_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_363 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_0__31_0__24_), .Q(w_mem_inst_w_mem_0__24_), .R(reset_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_364 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_0__31_0__25_), .Q(w_mem_inst_w_mem_0__25_), .R(reset_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_365 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_0__31_0__26_), .Q(w_mem_inst_w_mem_0__26_), .R(reset_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_366 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_0__31_0__27_), .Q(w_mem_inst_w_mem_0__27_), .R(reset_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_367 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_0__31_0__28_), .Q(w_mem_inst_w_mem_0__28_), .R(reset_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_368 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_0__31_0__29_), .Q(w_mem_inst_w_mem_0__29_), .R(reset_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_369 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_0__31_0__30_), .Q(w_mem_inst_w_mem_0__30_), .R(reset_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_37 ( .CLK(clk_bF_buf52), .D(b_reg_4__FF_INPUT), .Q(b_reg_4_), .R(reset_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_370 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_0__31_0__31_), .Q(w_mem_inst_w_mem_0__31_), .R(reset_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_371 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_1__31_0__0_), .Q(w_mem_inst_w_mem_1__0_), .R(reset_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_372 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_1__31_0__1_), .Q(w_mem_inst_w_mem_1__1_), .R(reset_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_373 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_1__31_0__2_), .Q(w_mem_inst_w_mem_1__2_), .R(reset_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_374 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_1__31_0__3_), .Q(w_mem_inst_w_mem_1__3_), .R(reset_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_375 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_1__31_0__4_), .Q(w_mem_inst_w_mem_1__4_), .R(reset_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_376 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_1__31_0__5_), .Q(w_mem_inst_w_mem_1__5_), .R(reset_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_377 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_1__31_0__6_), .Q(w_mem_inst_w_mem_1__6_), .R(reset_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_378 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_1__31_0__7_), .Q(w_mem_inst_w_mem_1__7_), .R(reset_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_379 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_1__31_0__8_), .Q(w_mem_inst_w_mem_1__8_), .R(reset_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_38 ( .CLK(clk_bF_buf51), .D(b_reg_5__FF_INPUT), .Q(b_reg_5_), .R(reset_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_380 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_1__31_0__9_), .Q(w_mem_inst_w_mem_1__9_), .R(reset_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_381 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_1__31_0__10_), .Q(w_mem_inst_w_mem_1__10_), .R(reset_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_382 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_1__31_0__11_), .Q(w_mem_inst_w_mem_1__11_), .R(reset_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_383 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_1__31_0__12_), .Q(w_mem_inst_w_mem_1__12_), .R(reset_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_384 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_1__31_0__13_), .Q(w_mem_inst_w_mem_1__13_), .R(reset_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_385 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_1__31_0__14_), .Q(w_mem_inst_w_mem_1__14_), .R(reset_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_386 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_1__31_0__15_), .Q(w_mem_inst_w_mem_1__15_), .R(reset_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_387 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_1__31_0__16_), .Q(w_mem_inst_w_mem_1__16_), .R(reset_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_388 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_1__31_0__17_), .Q(w_mem_inst_w_mem_1__17_), .R(reset_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_389 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_1__31_0__18_), .Q(w_mem_inst_w_mem_1__18_), .R(reset_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_39 ( .CLK(clk_bF_buf50), .D(b_reg_6__FF_INPUT), .Q(b_reg_6_), .R(reset_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_390 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_1__31_0__19_), .Q(w_mem_inst_w_mem_1__19_), .R(reset_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_391 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_1__31_0__20_), .Q(w_mem_inst_w_mem_1__20_), .R(reset_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_392 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_1__31_0__21_), .Q(w_mem_inst_w_mem_1__21_), .R(reset_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_393 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_1__31_0__22_), .Q(w_mem_inst_w_mem_1__22_), .R(reset_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_394 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_1__31_0__23_), .Q(w_mem_inst_w_mem_1__23_), .R(reset_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_395 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_1__31_0__24_), .Q(w_mem_inst_w_mem_1__24_), .R(reset_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_396 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_1__31_0__25_), .Q(w_mem_inst_w_mem_1__25_), .R(reset_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_397 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_1__31_0__26_), .Q(w_mem_inst_w_mem_1__26_), .R(reset_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_398 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_1__31_0__27_), .Q(w_mem_inst_w_mem_1__27_), .R(reset_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_399 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_1__31_0__28_), .Q(w_mem_inst_w_mem_1__28_), .R(reset_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_4 ( .CLK(clk_bF_buf85), .D(a_reg_3__FF_INPUT), .Q(a_reg_3_), .R(reset_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_40 ( .CLK(clk_bF_buf49), .D(b_reg_7__FF_INPUT), .Q(b_reg_7_), .R(reset_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_400 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_1__31_0__29_), .Q(w_mem_inst_w_mem_1__29_), .R(reset_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_401 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_1__31_0__30_), .Q(w_mem_inst_w_mem_1__30_), .R(reset_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_402 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_1__31_0__31_), .Q(w_mem_inst_w_mem_1__31_), .R(reset_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_403 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_2__31_0__0_), .Q(w_mem_inst_w_mem_2__0_), .R(reset_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_404 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_2__31_0__1_), .Q(w_mem_inst_w_mem_2__1_), .R(reset_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_405 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_2__31_0__2_), .Q(w_mem_inst_w_mem_2__2_), .R(reset_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_406 ( .CLK(clk_bF_buf39), .D(w_mem_inst__0w_mem_2__31_0__3_), .Q(w_mem_inst_w_mem_2__3_), .R(reset_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_407 ( .CLK(clk_bF_buf38), .D(w_mem_inst__0w_mem_2__31_0__4_), .Q(w_mem_inst_w_mem_2__4_), .R(reset_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_408 ( .CLK(clk_bF_buf37), .D(w_mem_inst__0w_mem_2__31_0__5_), .Q(w_mem_inst_w_mem_2__5_), .R(reset_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_409 ( .CLK(clk_bF_buf36), .D(w_mem_inst__0w_mem_2__31_0__6_), .Q(w_mem_inst_w_mem_2__6_), .R(reset_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_41 ( .CLK(clk_bF_buf48), .D(b_reg_8__FF_INPUT), .Q(b_reg_8_), .R(reset_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_410 ( .CLK(clk_bF_buf35), .D(w_mem_inst__0w_mem_2__31_0__7_), .Q(w_mem_inst_w_mem_2__7_), .R(reset_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_411 ( .CLK(clk_bF_buf34), .D(w_mem_inst__0w_mem_2__31_0__8_), .Q(w_mem_inst_w_mem_2__8_), .R(reset_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_412 ( .CLK(clk_bF_buf33), .D(w_mem_inst__0w_mem_2__31_0__9_), .Q(w_mem_inst_w_mem_2__9_), .R(reset_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_413 ( .CLK(clk_bF_buf32), .D(w_mem_inst__0w_mem_2__31_0__10_), .Q(w_mem_inst_w_mem_2__10_), .R(reset_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_414 ( .CLK(clk_bF_buf31), .D(w_mem_inst__0w_mem_2__31_0__11_), .Q(w_mem_inst_w_mem_2__11_), .R(reset_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_415 ( .CLK(clk_bF_buf30), .D(w_mem_inst__0w_mem_2__31_0__12_), .Q(w_mem_inst_w_mem_2__12_), .R(reset_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_416 ( .CLK(clk_bF_buf29), .D(w_mem_inst__0w_mem_2__31_0__13_), .Q(w_mem_inst_w_mem_2__13_), .R(reset_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_417 ( .CLK(clk_bF_buf28), .D(w_mem_inst__0w_mem_2__31_0__14_), .Q(w_mem_inst_w_mem_2__14_), .R(reset_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_418 ( .CLK(clk_bF_buf27), .D(w_mem_inst__0w_mem_2__31_0__15_), .Q(w_mem_inst_w_mem_2__15_), .R(reset_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_419 ( .CLK(clk_bF_buf26), .D(w_mem_inst__0w_mem_2__31_0__16_), .Q(w_mem_inst_w_mem_2__16_), .R(reset_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_42 ( .CLK(clk_bF_buf47), .D(b_reg_9__FF_INPUT), .Q(b_reg_9_), .R(reset_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_420 ( .CLK(clk_bF_buf25), .D(w_mem_inst__0w_mem_2__31_0__17_), .Q(w_mem_inst_w_mem_2__17_), .R(reset_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_421 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_mem_2__31_0__18_), .Q(w_mem_inst_w_mem_2__18_), .R(reset_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_422 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_mem_2__31_0__19_), .Q(w_mem_inst_w_mem_2__19_), .R(reset_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_423 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_mem_2__31_0__20_), .Q(w_mem_inst_w_mem_2__20_), .R(reset_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_424 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_mem_2__31_0__21_), .Q(w_mem_inst_w_mem_2__21_), .R(reset_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_425 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_mem_2__31_0__22_), .Q(w_mem_inst_w_mem_2__22_), .R(reset_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_426 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_mem_2__31_0__23_), .Q(w_mem_inst_w_mem_2__23_), .R(reset_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_427 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_mem_2__31_0__24_), .Q(w_mem_inst_w_mem_2__24_), .R(reset_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_428 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_2__31_0__25_), .Q(w_mem_inst_w_mem_2__25_), .R(reset_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_429 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_2__31_0__26_), .Q(w_mem_inst_w_mem_2__26_), .R(reset_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_43 ( .CLK(clk_bF_buf46), .D(b_reg_10__FF_INPUT), .Q(b_reg_10_), .R(reset_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_430 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_2__31_0__27_), .Q(w_mem_inst_w_mem_2__27_), .R(reset_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_431 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_2__31_0__28_), .Q(w_mem_inst_w_mem_2__28_), .R(reset_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_432 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_2__31_0__29_), .Q(w_mem_inst_w_mem_2__29_), .R(reset_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_433 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_2__31_0__30_), .Q(w_mem_inst_w_mem_2__30_), .R(reset_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_434 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_2__31_0__31_), .Q(w_mem_inst_w_mem_2__31_), .R(reset_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_435 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_3__31_0__0_), .Q(w_mem_inst_w_mem_3__0_), .R(reset_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_436 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_3__31_0__1_), .Q(w_mem_inst_w_mem_3__1_), .R(reset_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_437 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_3__31_0__2_), .Q(w_mem_inst_w_mem_3__2_), .R(reset_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_438 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_3__31_0__3_), .Q(w_mem_inst_w_mem_3__3_), .R(reset_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_439 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_3__31_0__4_), .Q(w_mem_inst_w_mem_3__4_), .R(reset_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_44 ( .CLK(clk_bF_buf45), .D(b_reg_11__FF_INPUT), .Q(b_reg_11_), .R(reset_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_440 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_3__31_0__5_), .Q(w_mem_inst_w_mem_3__5_), .R(reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_441 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_3__31_0__6_), .Q(w_mem_inst_w_mem_3__6_), .R(reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_442 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_3__31_0__7_), .Q(w_mem_inst_w_mem_3__7_), .R(reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_443 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_3__31_0__8_), .Q(w_mem_inst_w_mem_3__8_), .R(reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_444 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_3__31_0__9_), .Q(w_mem_inst_w_mem_3__9_), .R(reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_445 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_3__31_0__10_), .Q(w_mem_inst_w_mem_3__10_), .R(reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_446 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_3__31_0__11_), .Q(w_mem_inst_w_mem_3__11_), .R(reset_n_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_447 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_3__31_0__12_), .Q(w_mem_inst_w_mem_3__12_), .R(reset_n_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_448 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_3__31_0__13_), .Q(w_mem_inst_w_mem_3__13_), .R(reset_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_449 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_3__31_0__14_), .Q(w_mem_inst_w_mem_3__14_), .R(reset_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_45 ( .CLK(clk_bF_buf44), .D(b_reg_12__FF_INPUT), .Q(b_reg_12_), .R(reset_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_450 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_3__31_0__15_), .Q(w_mem_inst_w_mem_3__15_), .R(reset_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_451 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_3__31_0__16_), .Q(w_mem_inst_w_mem_3__16_), .R(reset_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_452 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_3__31_0__17_), .Q(w_mem_inst_w_mem_3__17_), .R(reset_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_453 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_3__31_0__18_), .Q(w_mem_inst_w_mem_3__18_), .R(reset_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_454 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_3__31_0__19_), .Q(w_mem_inst_w_mem_3__19_), .R(reset_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_455 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_3__31_0__20_), .Q(w_mem_inst_w_mem_3__20_), .R(reset_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_456 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_3__31_0__21_), .Q(w_mem_inst_w_mem_3__21_), .R(reset_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_457 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_3__31_0__22_), .Q(w_mem_inst_w_mem_3__22_), .R(reset_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_458 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_3__31_0__23_), .Q(w_mem_inst_w_mem_3__23_), .R(reset_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_459 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_3__31_0__24_), .Q(w_mem_inst_w_mem_3__24_), .R(reset_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_46 ( .CLK(clk_bF_buf43), .D(b_reg_13__FF_INPUT), .Q(b_reg_13_), .R(reset_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_460 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_3__31_0__25_), .Q(w_mem_inst_w_mem_3__25_), .R(reset_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_461 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_3__31_0__26_), .Q(w_mem_inst_w_mem_3__26_), .R(reset_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_462 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_3__31_0__27_), .Q(w_mem_inst_w_mem_3__27_), .R(reset_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_463 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_3__31_0__28_), .Q(w_mem_inst_w_mem_3__28_), .R(reset_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_464 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_3__31_0__29_), .Q(w_mem_inst_w_mem_3__29_), .R(reset_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_465 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_3__31_0__30_), .Q(w_mem_inst_w_mem_3__30_), .R(reset_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_466 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_3__31_0__31_), .Q(w_mem_inst_w_mem_3__31_), .R(reset_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_467 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_4__31_0__0_), .Q(w_mem_inst_w_mem_4__0_), .R(reset_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_468 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_4__31_0__1_), .Q(w_mem_inst_w_mem_4__1_), .R(reset_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_469 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_4__31_0__2_), .Q(w_mem_inst_w_mem_4__2_), .R(reset_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_47 ( .CLK(clk_bF_buf42), .D(b_reg_14__FF_INPUT), .Q(b_reg_14_), .R(reset_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_470 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_4__31_0__3_), .Q(w_mem_inst_w_mem_4__3_), .R(reset_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_471 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_4__31_0__4_), .Q(w_mem_inst_w_mem_4__4_), .R(reset_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_472 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_4__31_0__5_), .Q(w_mem_inst_w_mem_4__5_), .R(reset_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_473 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_4__31_0__6_), .Q(w_mem_inst_w_mem_4__6_), .R(reset_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_474 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_4__31_0__7_), .Q(w_mem_inst_w_mem_4__7_), .R(reset_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_475 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_4__31_0__8_), .Q(w_mem_inst_w_mem_4__8_), .R(reset_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_476 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_4__31_0__9_), .Q(w_mem_inst_w_mem_4__9_), .R(reset_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_477 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_4__31_0__10_), .Q(w_mem_inst_w_mem_4__10_), .R(reset_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_478 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_4__31_0__11_), .Q(w_mem_inst_w_mem_4__11_), .R(reset_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_479 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_4__31_0__12_), .Q(w_mem_inst_w_mem_4__12_), .R(reset_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_48 ( .CLK(clk_bF_buf41), .D(b_reg_15__FF_INPUT), .Q(b_reg_15_), .R(reset_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_480 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_4__31_0__13_), .Q(w_mem_inst_w_mem_4__13_), .R(reset_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_481 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_4__31_0__14_), .Q(w_mem_inst_w_mem_4__14_), .R(reset_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_482 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_4__31_0__15_), .Q(w_mem_inst_w_mem_4__15_), .R(reset_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_483 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_4__31_0__16_), .Q(w_mem_inst_w_mem_4__16_), .R(reset_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_484 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_4__31_0__17_), .Q(w_mem_inst_w_mem_4__17_), .R(reset_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_485 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_4__31_0__18_), .Q(w_mem_inst_w_mem_4__18_), .R(reset_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_486 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_4__31_0__19_), .Q(w_mem_inst_w_mem_4__19_), .R(reset_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_487 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_4__31_0__20_), .Q(w_mem_inst_w_mem_4__20_), .R(reset_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_488 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_4__31_0__21_), .Q(w_mem_inst_w_mem_4__21_), .R(reset_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_489 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_4__31_0__22_), .Q(w_mem_inst_w_mem_4__22_), .R(reset_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_49 ( .CLK(clk_bF_buf40), .D(b_reg_16__FF_INPUT), .Q(b_reg_16_), .R(reset_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_490 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_4__31_0__23_), .Q(w_mem_inst_w_mem_4__23_), .R(reset_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_491 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_4__31_0__24_), .Q(w_mem_inst_w_mem_4__24_), .R(reset_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_492 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_4__31_0__25_), .Q(w_mem_inst_w_mem_4__25_), .R(reset_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_493 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_4__31_0__26_), .Q(w_mem_inst_w_mem_4__26_), .R(reset_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_494 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_4__31_0__27_), .Q(w_mem_inst_w_mem_4__27_), .R(reset_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_495 ( .CLK(clk_bF_buf39), .D(w_mem_inst__0w_mem_4__31_0__28_), .Q(w_mem_inst_w_mem_4__28_), .R(reset_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_496 ( .CLK(clk_bF_buf38), .D(w_mem_inst__0w_mem_4__31_0__29_), .Q(w_mem_inst_w_mem_4__29_), .R(reset_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_497 ( .CLK(clk_bF_buf37), .D(w_mem_inst__0w_mem_4__31_0__30_), .Q(w_mem_inst_w_mem_4__30_), .R(reset_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_498 ( .CLK(clk_bF_buf36), .D(w_mem_inst__0w_mem_4__31_0__31_), .Q(w_mem_inst_w_mem_4__31_), .R(reset_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_499 ( .CLK(clk_bF_buf35), .D(w_mem_inst__0w_mem_5__31_0__0_), .Q(w_mem_inst_w_mem_5__0_), .R(reset_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_5 ( .CLK(clk_bF_buf84), .D(a_reg_4__FF_INPUT), .Q(a_reg_4_), .R(reset_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_50 ( .CLK(clk_bF_buf39), .D(b_reg_17__FF_INPUT), .Q(b_reg_17_), .R(reset_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_500 ( .CLK(clk_bF_buf34), .D(w_mem_inst__0w_mem_5__31_0__1_), .Q(w_mem_inst_w_mem_5__1_), .R(reset_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_501 ( .CLK(clk_bF_buf33), .D(w_mem_inst__0w_mem_5__31_0__2_), .Q(w_mem_inst_w_mem_5__2_), .R(reset_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_502 ( .CLK(clk_bF_buf32), .D(w_mem_inst__0w_mem_5__31_0__3_), .Q(w_mem_inst_w_mem_5__3_), .R(reset_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_503 ( .CLK(clk_bF_buf31), .D(w_mem_inst__0w_mem_5__31_0__4_), .Q(w_mem_inst_w_mem_5__4_), .R(reset_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_504 ( .CLK(clk_bF_buf30), .D(w_mem_inst__0w_mem_5__31_0__5_), .Q(w_mem_inst_w_mem_5__5_), .R(reset_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_505 ( .CLK(clk_bF_buf29), .D(w_mem_inst__0w_mem_5__31_0__6_), .Q(w_mem_inst_w_mem_5__6_), .R(reset_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_506 ( .CLK(clk_bF_buf28), .D(w_mem_inst__0w_mem_5__31_0__7_), .Q(w_mem_inst_w_mem_5__7_), .R(reset_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_507 ( .CLK(clk_bF_buf27), .D(w_mem_inst__0w_mem_5__31_0__8_), .Q(w_mem_inst_w_mem_5__8_), .R(reset_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_508 ( .CLK(clk_bF_buf26), .D(w_mem_inst__0w_mem_5__31_0__9_), .Q(w_mem_inst_w_mem_5__9_), .R(reset_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_509 ( .CLK(clk_bF_buf25), .D(w_mem_inst__0w_mem_5__31_0__10_), .Q(w_mem_inst_w_mem_5__10_), .R(reset_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_51 ( .CLK(clk_bF_buf38), .D(b_reg_18__FF_INPUT), .Q(b_reg_18_), .R(reset_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_510 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_mem_5__31_0__11_), .Q(w_mem_inst_w_mem_5__11_), .R(reset_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_511 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_mem_5__31_0__12_), .Q(w_mem_inst_w_mem_5__12_), .R(reset_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_512 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_mem_5__31_0__13_), .Q(w_mem_inst_w_mem_5__13_), .R(reset_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_513 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_mem_5__31_0__14_), .Q(w_mem_inst_w_mem_5__14_), .R(reset_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_514 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_mem_5__31_0__15_), .Q(w_mem_inst_w_mem_5__15_), .R(reset_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_515 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_mem_5__31_0__16_), .Q(w_mem_inst_w_mem_5__16_), .R(reset_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_516 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_mem_5__31_0__17_), .Q(w_mem_inst_w_mem_5__17_), .R(reset_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_517 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_5__31_0__18_), .Q(w_mem_inst_w_mem_5__18_), .R(reset_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_518 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_5__31_0__19_), .Q(w_mem_inst_w_mem_5__19_), .R(reset_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_519 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_5__31_0__20_), .Q(w_mem_inst_w_mem_5__20_), .R(reset_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_52 ( .CLK(clk_bF_buf37), .D(b_reg_19__FF_INPUT), .Q(b_reg_19_), .R(reset_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_520 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_5__31_0__21_), .Q(w_mem_inst_w_mem_5__21_), .R(reset_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_521 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_5__31_0__22_), .Q(w_mem_inst_w_mem_5__22_), .R(reset_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_522 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_5__31_0__23_), .Q(w_mem_inst_w_mem_5__23_), .R(reset_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_523 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_5__31_0__24_), .Q(w_mem_inst_w_mem_5__24_), .R(reset_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_524 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_5__31_0__25_), .Q(w_mem_inst_w_mem_5__25_), .R(reset_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_525 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_5__31_0__26_), .Q(w_mem_inst_w_mem_5__26_), .R(reset_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_526 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_5__31_0__27_), .Q(w_mem_inst_w_mem_5__27_), .R(reset_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_527 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_5__31_0__28_), .Q(w_mem_inst_w_mem_5__28_), .R(reset_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_528 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_5__31_0__29_), .Q(w_mem_inst_w_mem_5__29_), .R(reset_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_529 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_5__31_0__30_), .Q(w_mem_inst_w_mem_5__30_), .R(reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_53 ( .CLK(clk_bF_buf36), .D(b_reg_20__FF_INPUT), .Q(b_reg_20_), .R(reset_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_530 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_5__31_0__31_), .Q(w_mem_inst_w_mem_5__31_), .R(reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_531 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_6__31_0__0_), .Q(w_mem_inst_w_mem_6__0_), .R(reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_532 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_6__31_0__1_), .Q(w_mem_inst_w_mem_6__1_), .R(reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_533 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_6__31_0__2_), .Q(w_mem_inst_w_mem_6__2_), .R(reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_534 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_6__31_0__3_), .Q(w_mem_inst_w_mem_6__3_), .R(reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_535 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_6__31_0__4_), .Q(w_mem_inst_w_mem_6__4_), .R(reset_n_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_536 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_6__31_0__5_), .Q(w_mem_inst_w_mem_6__5_), .R(reset_n_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_537 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_6__31_0__6_), .Q(w_mem_inst_w_mem_6__6_), .R(reset_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_538 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_6__31_0__7_), .Q(w_mem_inst_w_mem_6__7_), .R(reset_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_539 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_6__31_0__8_), .Q(w_mem_inst_w_mem_6__8_), .R(reset_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_54 ( .CLK(clk_bF_buf35), .D(b_reg_21__FF_INPUT), .Q(b_reg_21_), .R(reset_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_540 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_6__31_0__9_), .Q(w_mem_inst_w_mem_6__9_), .R(reset_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_541 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_6__31_0__10_), .Q(w_mem_inst_w_mem_6__10_), .R(reset_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_542 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_6__31_0__11_), .Q(w_mem_inst_w_mem_6__11_), .R(reset_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_543 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_6__31_0__12_), .Q(w_mem_inst_w_mem_6__12_), .R(reset_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_544 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_6__31_0__13_), .Q(w_mem_inst_w_mem_6__13_), .R(reset_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_545 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_6__31_0__14_), .Q(w_mem_inst_w_mem_6__14_), .R(reset_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_546 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_6__31_0__15_), .Q(w_mem_inst_w_mem_6__15_), .R(reset_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_547 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_6__31_0__16_), .Q(w_mem_inst_w_mem_6__16_), .R(reset_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_548 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_6__31_0__17_), .Q(w_mem_inst_w_mem_6__17_), .R(reset_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_549 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_6__31_0__18_), .Q(w_mem_inst_w_mem_6__18_), .R(reset_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_55 ( .CLK(clk_bF_buf34), .D(b_reg_22__FF_INPUT), .Q(b_reg_22_), .R(reset_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_550 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_6__31_0__19_), .Q(w_mem_inst_w_mem_6__19_), .R(reset_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_551 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_6__31_0__20_), .Q(w_mem_inst_w_mem_6__20_), .R(reset_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_552 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_6__31_0__21_), .Q(w_mem_inst_w_mem_6__21_), .R(reset_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_553 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_6__31_0__22_), .Q(w_mem_inst_w_mem_6__22_), .R(reset_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_554 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_6__31_0__23_), .Q(w_mem_inst_w_mem_6__23_), .R(reset_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_555 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_6__31_0__24_), .Q(w_mem_inst_w_mem_6__24_), .R(reset_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_556 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_6__31_0__25_), .Q(w_mem_inst_w_mem_6__25_), .R(reset_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_557 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_6__31_0__26_), .Q(w_mem_inst_w_mem_6__26_), .R(reset_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_558 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_6__31_0__27_), .Q(w_mem_inst_w_mem_6__27_), .R(reset_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_559 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_6__31_0__28_), .Q(w_mem_inst_w_mem_6__28_), .R(reset_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_56 ( .CLK(clk_bF_buf33), .D(b_reg_23__FF_INPUT), .Q(b_reg_23_), .R(reset_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_560 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_6__31_0__29_), .Q(w_mem_inst_w_mem_6__29_), .R(reset_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_561 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_6__31_0__30_), .Q(w_mem_inst_w_mem_6__30_), .R(reset_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_562 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_6__31_0__31_), .Q(w_mem_inst_w_mem_6__31_), .R(reset_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_563 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_7__31_0__0_), .Q(w_mem_inst_w_mem_7__0_), .R(reset_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_564 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_7__31_0__1_), .Q(w_mem_inst_w_mem_7__1_), .R(reset_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_565 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_7__31_0__2_), .Q(w_mem_inst_w_mem_7__2_), .R(reset_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_566 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_7__31_0__3_), .Q(w_mem_inst_w_mem_7__3_), .R(reset_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_567 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_7__31_0__4_), .Q(w_mem_inst_w_mem_7__4_), .R(reset_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_568 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_7__31_0__5_), .Q(w_mem_inst_w_mem_7__5_), .R(reset_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_569 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_7__31_0__6_), .Q(w_mem_inst_w_mem_7__6_), .R(reset_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_57 ( .CLK(clk_bF_buf32), .D(b_reg_24__FF_INPUT), .Q(b_reg_24_), .R(reset_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_570 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_7__31_0__7_), .Q(w_mem_inst_w_mem_7__7_), .R(reset_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_571 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_7__31_0__8_), .Q(w_mem_inst_w_mem_7__8_), .R(reset_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_572 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_7__31_0__9_), .Q(w_mem_inst_w_mem_7__9_), .R(reset_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_573 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_7__31_0__10_), .Q(w_mem_inst_w_mem_7__10_), .R(reset_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_574 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_7__31_0__11_), .Q(w_mem_inst_w_mem_7__11_), .R(reset_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_575 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_7__31_0__12_), .Q(w_mem_inst_w_mem_7__12_), .R(reset_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_576 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_7__31_0__13_), .Q(w_mem_inst_w_mem_7__13_), .R(reset_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_577 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_7__31_0__14_), .Q(w_mem_inst_w_mem_7__14_), .R(reset_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_578 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_7__31_0__15_), .Q(w_mem_inst_w_mem_7__15_), .R(reset_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_579 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_7__31_0__16_), .Q(w_mem_inst_w_mem_7__16_), .R(reset_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_58 ( .CLK(clk_bF_buf31), .D(b_reg_25__FF_INPUT), .Q(b_reg_25_), .R(reset_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_580 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_7__31_0__17_), .Q(w_mem_inst_w_mem_7__17_), .R(reset_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_581 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_7__31_0__18_), .Q(w_mem_inst_w_mem_7__18_), .R(reset_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_582 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_7__31_0__19_), .Q(w_mem_inst_w_mem_7__19_), .R(reset_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_583 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_7__31_0__20_), .Q(w_mem_inst_w_mem_7__20_), .R(reset_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_584 ( .CLK(clk_bF_buf39), .D(w_mem_inst__0w_mem_7__31_0__21_), .Q(w_mem_inst_w_mem_7__21_), .R(reset_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_585 ( .CLK(clk_bF_buf38), .D(w_mem_inst__0w_mem_7__31_0__22_), .Q(w_mem_inst_w_mem_7__22_), .R(reset_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_586 ( .CLK(clk_bF_buf37), .D(w_mem_inst__0w_mem_7__31_0__23_), .Q(w_mem_inst_w_mem_7__23_), .R(reset_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_587 ( .CLK(clk_bF_buf36), .D(w_mem_inst__0w_mem_7__31_0__24_), .Q(w_mem_inst_w_mem_7__24_), .R(reset_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_588 ( .CLK(clk_bF_buf35), .D(w_mem_inst__0w_mem_7__31_0__25_), .Q(w_mem_inst_w_mem_7__25_), .R(reset_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_589 ( .CLK(clk_bF_buf34), .D(w_mem_inst__0w_mem_7__31_0__26_), .Q(w_mem_inst_w_mem_7__26_), .R(reset_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_59 ( .CLK(clk_bF_buf30), .D(b_reg_26__FF_INPUT), .Q(b_reg_26_), .R(reset_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_590 ( .CLK(clk_bF_buf33), .D(w_mem_inst__0w_mem_7__31_0__27_), .Q(w_mem_inst_w_mem_7__27_), .R(reset_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_591 ( .CLK(clk_bF_buf32), .D(w_mem_inst__0w_mem_7__31_0__28_), .Q(w_mem_inst_w_mem_7__28_), .R(reset_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_592 ( .CLK(clk_bF_buf31), .D(w_mem_inst__0w_mem_7__31_0__29_), .Q(w_mem_inst_w_mem_7__29_), .R(reset_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_593 ( .CLK(clk_bF_buf30), .D(w_mem_inst__0w_mem_7__31_0__30_), .Q(w_mem_inst_w_mem_7__30_), .R(reset_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_594 ( .CLK(clk_bF_buf29), .D(w_mem_inst__0w_mem_7__31_0__31_), .Q(w_mem_inst_w_mem_7__31_), .R(reset_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_595 ( .CLK(clk_bF_buf28), .D(w_mem_inst__0w_mem_8__31_0__0_), .Q(w_mem_inst_w_mem_8__0_), .R(reset_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_596 ( .CLK(clk_bF_buf27), .D(w_mem_inst__0w_mem_8__31_0__1_), .Q(w_mem_inst_w_mem_8__1_), .R(reset_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_597 ( .CLK(clk_bF_buf26), .D(w_mem_inst__0w_mem_8__31_0__2_), .Q(w_mem_inst_w_mem_8__2_), .R(reset_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_598 ( .CLK(clk_bF_buf25), .D(w_mem_inst__0w_mem_8__31_0__3_), .Q(w_mem_inst_w_mem_8__3_), .R(reset_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_599 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_mem_8__31_0__4_), .Q(w_mem_inst_w_mem_8__4_), .R(reset_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_6 ( .CLK(clk_bF_buf83), .D(a_reg_5__FF_INPUT), .Q(a_reg_5_), .R(reset_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_60 ( .CLK(clk_bF_buf29), .D(b_reg_27__FF_INPUT), .Q(b_reg_27_), .R(reset_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_600 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_mem_8__31_0__5_), .Q(w_mem_inst_w_mem_8__5_), .R(reset_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_601 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_mem_8__31_0__6_), .Q(w_mem_inst_w_mem_8__6_), .R(reset_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_602 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_mem_8__31_0__7_), .Q(w_mem_inst_w_mem_8__7_), .R(reset_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_603 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_mem_8__31_0__8_), .Q(w_mem_inst_w_mem_8__8_), .R(reset_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_604 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_mem_8__31_0__9_), .Q(w_mem_inst_w_mem_8__9_), .R(reset_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_605 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_mem_8__31_0__10_), .Q(w_mem_inst_w_mem_8__10_), .R(reset_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_606 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_8__31_0__11_), .Q(w_mem_inst_w_mem_8__11_), .R(reset_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_607 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_8__31_0__12_), .Q(w_mem_inst_w_mem_8__12_), .R(reset_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_608 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_8__31_0__13_), .Q(w_mem_inst_w_mem_8__13_), .R(reset_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_609 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_8__31_0__14_), .Q(w_mem_inst_w_mem_8__14_), .R(reset_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_61 ( .CLK(clk_bF_buf28), .D(b_reg_28__FF_INPUT), .Q(b_reg_28_), .R(reset_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_610 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_8__31_0__15_), .Q(w_mem_inst_w_mem_8__15_), .R(reset_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_611 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_8__31_0__16_), .Q(w_mem_inst_w_mem_8__16_), .R(reset_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_612 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_8__31_0__17_), .Q(w_mem_inst_w_mem_8__17_), .R(reset_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_613 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_8__31_0__18_), .Q(w_mem_inst_w_mem_8__18_), .R(reset_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_614 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_8__31_0__19_), .Q(w_mem_inst_w_mem_8__19_), .R(reset_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_615 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_8__31_0__20_), .Q(w_mem_inst_w_mem_8__20_), .R(reset_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_616 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_8__31_0__21_), .Q(w_mem_inst_w_mem_8__21_), .R(reset_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_617 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_8__31_0__22_), .Q(w_mem_inst_w_mem_8__22_), .R(reset_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_618 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_8__31_0__23_), .Q(w_mem_inst_w_mem_8__23_), .R(reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_619 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_8__31_0__24_), .Q(w_mem_inst_w_mem_8__24_), .R(reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_62 ( .CLK(clk_bF_buf27), .D(b_reg_29__FF_INPUT), .Q(b_reg_29_), .R(reset_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_620 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_8__31_0__25_), .Q(w_mem_inst_w_mem_8__25_), .R(reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_621 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_8__31_0__26_), .Q(w_mem_inst_w_mem_8__26_), .R(reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_622 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_8__31_0__27_), .Q(w_mem_inst_w_mem_8__27_), .R(reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_623 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_8__31_0__28_), .Q(w_mem_inst_w_mem_8__28_), .R(reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_624 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_8__31_0__29_), .Q(w_mem_inst_w_mem_8__29_), .R(reset_n_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_625 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_8__31_0__30_), .Q(w_mem_inst_w_mem_8__30_), .R(reset_n_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_626 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_8__31_0__31_), .Q(w_mem_inst_w_mem_8__31_), .R(reset_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_627 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_9__31_0__0_), .Q(w_mem_inst_w_mem_9__0_), .R(reset_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_628 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_9__31_0__1_), .Q(w_mem_inst_w_mem_9__1_), .R(reset_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_629 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_9__31_0__2_), .Q(w_mem_inst_w_mem_9__2_), .R(reset_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_63 ( .CLK(clk_bF_buf26), .D(b_reg_30__FF_INPUT), .Q(b_reg_30_), .R(reset_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_630 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_9__31_0__3_), .Q(w_mem_inst_w_mem_9__3_), .R(reset_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_631 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_9__31_0__4_), .Q(w_mem_inst_w_mem_9__4_), .R(reset_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_632 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_9__31_0__5_), .Q(w_mem_inst_w_mem_9__5_), .R(reset_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_633 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_9__31_0__6_), .Q(w_mem_inst_w_mem_9__6_), .R(reset_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_634 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_9__31_0__7_), .Q(w_mem_inst_w_mem_9__7_), .R(reset_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_635 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_9__31_0__8_), .Q(w_mem_inst_w_mem_9__8_), .R(reset_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_636 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_9__31_0__9_), .Q(w_mem_inst_w_mem_9__9_), .R(reset_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_637 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_9__31_0__10_), .Q(w_mem_inst_w_mem_9__10_), .R(reset_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_638 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_9__31_0__11_), .Q(w_mem_inst_w_mem_9__11_), .R(reset_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_639 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_9__31_0__12_), .Q(w_mem_inst_w_mem_9__12_), .R(reset_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_64 ( .CLK(clk_bF_buf25), .D(b_reg_31__FF_INPUT), .Q(b_reg_31_), .R(reset_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_640 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_9__31_0__13_), .Q(w_mem_inst_w_mem_9__13_), .R(reset_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_641 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_9__31_0__14_), .Q(w_mem_inst_w_mem_9__14_), .R(reset_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_642 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_9__31_0__15_), .Q(w_mem_inst_w_mem_9__15_), .R(reset_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_643 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_9__31_0__16_), .Q(w_mem_inst_w_mem_9__16_), .R(reset_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_644 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_9__31_0__17_), .Q(w_mem_inst_w_mem_9__17_), .R(reset_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_645 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_9__31_0__18_), .Q(w_mem_inst_w_mem_9__18_), .R(reset_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_646 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_9__31_0__19_), .Q(w_mem_inst_w_mem_9__19_), .R(reset_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_647 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_9__31_0__20_), .Q(w_mem_inst_w_mem_9__20_), .R(reset_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_648 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_9__31_0__21_), .Q(w_mem_inst_w_mem_9__21_), .R(reset_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_649 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_9__31_0__22_), .Q(w_mem_inst_w_mem_9__22_), .R(reset_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_65 ( .CLK(clk_bF_buf24), .D(c_reg_0__FF_INPUT), .Q(c_reg_0_), .R(reset_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_650 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_9__31_0__23_), .Q(w_mem_inst_w_mem_9__23_), .R(reset_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_651 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_9__31_0__24_), .Q(w_mem_inst_w_mem_9__24_), .R(reset_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_652 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_9__31_0__25_), .Q(w_mem_inst_w_mem_9__25_), .R(reset_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_653 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_9__31_0__26_), .Q(w_mem_inst_w_mem_9__26_), .R(reset_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_654 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_9__31_0__27_), .Q(w_mem_inst_w_mem_9__27_), .R(reset_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_655 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_9__31_0__28_), .Q(w_mem_inst_w_mem_9__28_), .R(reset_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_656 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_9__31_0__29_), .Q(w_mem_inst_w_mem_9__29_), .R(reset_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_657 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_9__31_0__30_), .Q(w_mem_inst_w_mem_9__30_), .R(reset_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_658 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_9__31_0__31_), .Q(w_mem_inst_w_mem_9__31_), .R(reset_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_659 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_10__31_0__0_), .Q(w_mem_inst_w_mem_10__0_), .R(reset_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_66 ( .CLK(clk_bF_buf23), .D(c_reg_1__FF_INPUT), .Q(c_reg_1_), .R(reset_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_660 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_10__31_0__1_), .Q(w_mem_inst_w_mem_10__1_), .R(reset_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_661 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_10__31_0__2_), .Q(w_mem_inst_w_mem_10__2_), .R(reset_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_662 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_10__31_0__3_), .Q(w_mem_inst_w_mem_10__3_), .R(reset_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_663 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_10__31_0__4_), .Q(w_mem_inst_w_mem_10__4_), .R(reset_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_664 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_10__31_0__5_), .Q(w_mem_inst_w_mem_10__5_), .R(reset_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_665 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_10__31_0__6_), .Q(w_mem_inst_w_mem_10__6_), .R(reset_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_666 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_10__31_0__7_), .Q(w_mem_inst_w_mem_10__7_), .R(reset_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_667 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_10__31_0__8_), .Q(w_mem_inst_w_mem_10__8_), .R(reset_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_668 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_10__31_0__9_), .Q(w_mem_inst_w_mem_10__9_), .R(reset_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_669 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_10__31_0__10_), .Q(w_mem_inst_w_mem_10__10_), .R(reset_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_67 ( .CLK(clk_bF_buf22), .D(c_reg_2__FF_INPUT), .Q(c_reg_2_), .R(reset_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_670 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_10__31_0__11_), .Q(w_mem_inst_w_mem_10__11_), .R(reset_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_671 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_10__31_0__12_), .Q(w_mem_inst_w_mem_10__12_), .R(reset_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_672 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_10__31_0__13_), .Q(w_mem_inst_w_mem_10__13_), .R(reset_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_673 ( .CLK(clk_bF_buf39), .D(w_mem_inst__0w_mem_10__31_0__14_), .Q(w_mem_inst_w_mem_10__14_), .R(reset_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_674 ( .CLK(clk_bF_buf38), .D(w_mem_inst__0w_mem_10__31_0__15_), .Q(w_mem_inst_w_mem_10__15_), .R(reset_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_675 ( .CLK(clk_bF_buf37), .D(w_mem_inst__0w_mem_10__31_0__16_), .Q(w_mem_inst_w_mem_10__16_), .R(reset_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_676 ( .CLK(clk_bF_buf36), .D(w_mem_inst__0w_mem_10__31_0__17_), .Q(w_mem_inst_w_mem_10__17_), .R(reset_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_677 ( .CLK(clk_bF_buf35), .D(w_mem_inst__0w_mem_10__31_0__18_), .Q(w_mem_inst_w_mem_10__18_), .R(reset_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_678 ( .CLK(clk_bF_buf34), .D(w_mem_inst__0w_mem_10__31_0__19_), .Q(w_mem_inst_w_mem_10__19_), .R(reset_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_679 ( .CLK(clk_bF_buf33), .D(w_mem_inst__0w_mem_10__31_0__20_), .Q(w_mem_inst_w_mem_10__20_), .R(reset_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_68 ( .CLK(clk_bF_buf21), .D(c_reg_3__FF_INPUT), .Q(c_reg_3_), .R(reset_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_680 ( .CLK(clk_bF_buf32), .D(w_mem_inst__0w_mem_10__31_0__21_), .Q(w_mem_inst_w_mem_10__21_), .R(reset_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_681 ( .CLK(clk_bF_buf31), .D(w_mem_inst__0w_mem_10__31_0__22_), .Q(w_mem_inst_w_mem_10__22_), .R(reset_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_682 ( .CLK(clk_bF_buf30), .D(w_mem_inst__0w_mem_10__31_0__23_), .Q(w_mem_inst_w_mem_10__23_), .R(reset_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_683 ( .CLK(clk_bF_buf29), .D(w_mem_inst__0w_mem_10__31_0__24_), .Q(w_mem_inst_w_mem_10__24_), .R(reset_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_684 ( .CLK(clk_bF_buf28), .D(w_mem_inst__0w_mem_10__31_0__25_), .Q(w_mem_inst_w_mem_10__25_), .R(reset_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_685 ( .CLK(clk_bF_buf27), .D(w_mem_inst__0w_mem_10__31_0__26_), .Q(w_mem_inst_w_mem_10__26_), .R(reset_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_686 ( .CLK(clk_bF_buf26), .D(w_mem_inst__0w_mem_10__31_0__27_), .Q(w_mem_inst_w_mem_10__27_), .R(reset_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_687 ( .CLK(clk_bF_buf25), .D(w_mem_inst__0w_mem_10__31_0__28_), .Q(w_mem_inst_w_mem_10__28_), .R(reset_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_688 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_mem_10__31_0__29_), .Q(w_mem_inst_w_mem_10__29_), .R(reset_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_689 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_mem_10__31_0__30_), .Q(w_mem_inst_w_mem_10__30_), .R(reset_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_69 ( .CLK(clk_bF_buf20), .D(c_reg_4__FF_INPUT), .Q(c_reg_4_), .R(reset_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_690 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_mem_10__31_0__31_), .Q(w_mem_inst_w_mem_10__31_), .R(reset_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_691 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_mem_11__31_0__0_), .Q(w_mem_inst_w_mem_11__0_), .R(reset_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_692 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_mem_11__31_0__1_), .Q(w_mem_inst_w_mem_11__1_), .R(reset_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_693 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_mem_11__31_0__2_), .Q(w_mem_inst_w_mem_11__2_), .R(reset_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_694 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_mem_11__31_0__3_), .Q(w_mem_inst_w_mem_11__3_), .R(reset_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_695 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_11__31_0__4_), .Q(w_mem_inst_w_mem_11__4_), .R(reset_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_696 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_11__31_0__5_), .Q(w_mem_inst_w_mem_11__5_), .R(reset_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_697 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_11__31_0__6_), .Q(w_mem_inst_w_mem_11__6_), .R(reset_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_698 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_11__31_0__7_), .Q(w_mem_inst_w_mem_11__7_), .R(reset_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_699 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_11__31_0__8_), .Q(w_mem_inst_w_mem_11__8_), .R(reset_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_7 ( .CLK(clk_bF_buf82), .D(a_reg_6__FF_INPUT), .Q(a_reg_6_), .R(reset_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_70 ( .CLK(clk_bF_buf19), .D(c_reg_5__FF_INPUT), .Q(c_reg_5_), .R(reset_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_700 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_11__31_0__9_), .Q(w_mem_inst_w_mem_11__9_), .R(reset_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_701 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_11__31_0__10_), .Q(w_mem_inst_w_mem_11__10_), .R(reset_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_702 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_11__31_0__11_), .Q(w_mem_inst_w_mem_11__11_), .R(reset_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_703 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_11__31_0__12_), .Q(w_mem_inst_w_mem_11__12_), .R(reset_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_704 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_11__31_0__13_), .Q(w_mem_inst_w_mem_11__13_), .R(reset_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_705 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_11__31_0__14_), .Q(w_mem_inst_w_mem_11__14_), .R(reset_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_706 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_11__31_0__15_), .Q(w_mem_inst_w_mem_11__15_), .R(reset_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_707 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_11__31_0__16_), .Q(w_mem_inst_w_mem_11__16_), .R(reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_708 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_11__31_0__17_), .Q(w_mem_inst_w_mem_11__17_), .R(reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_709 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_11__31_0__18_), .Q(w_mem_inst_w_mem_11__18_), .R(reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_71 ( .CLK(clk_bF_buf18), .D(c_reg_6__FF_INPUT), .Q(c_reg_6_), .R(reset_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_710 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_11__31_0__19_), .Q(w_mem_inst_w_mem_11__19_), .R(reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_711 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_11__31_0__20_), .Q(w_mem_inst_w_mem_11__20_), .R(reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_712 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_11__31_0__21_), .Q(w_mem_inst_w_mem_11__21_), .R(reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_713 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_11__31_0__22_), .Q(w_mem_inst_w_mem_11__22_), .R(reset_n_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_714 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_11__31_0__23_), .Q(w_mem_inst_w_mem_11__23_), .R(reset_n_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_715 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_11__31_0__24_), .Q(w_mem_inst_w_mem_11__24_), .R(reset_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_716 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_11__31_0__25_), .Q(w_mem_inst_w_mem_11__25_), .R(reset_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_717 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_11__31_0__26_), .Q(w_mem_inst_w_mem_11__26_), .R(reset_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_718 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_11__31_0__27_), .Q(w_mem_inst_w_mem_11__27_), .R(reset_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_719 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_11__31_0__28_), .Q(w_mem_inst_w_mem_11__28_), .R(reset_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_72 ( .CLK(clk_bF_buf17), .D(c_reg_7__FF_INPUT), .Q(c_reg_7_), .R(reset_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_720 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_11__31_0__29_), .Q(w_mem_inst_w_mem_11__29_), .R(reset_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_721 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_11__31_0__30_), .Q(w_mem_inst_w_mem_11__30_), .R(reset_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_722 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_11__31_0__31_), .Q(w_mem_inst_w_mem_11__31_), .R(reset_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_723 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_12__31_0__0_), .Q(w_mem_inst_w_mem_12__0_), .R(reset_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_724 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_12__31_0__1_), .Q(w_mem_inst_w_mem_12__1_), .R(reset_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_725 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_12__31_0__2_), .Q(w_mem_inst_w_mem_12__2_), .R(reset_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_726 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_12__31_0__3_), .Q(w_mem_inst_w_mem_12__3_), .R(reset_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_727 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_12__31_0__4_), .Q(w_mem_inst_w_mem_12__4_), .R(reset_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_728 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_12__31_0__5_), .Q(w_mem_inst_w_mem_12__5_), .R(reset_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_729 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_12__31_0__6_), .Q(w_mem_inst_w_mem_12__6_), .R(reset_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_73 ( .CLK(clk_bF_buf16), .D(c_reg_8__FF_INPUT), .Q(c_reg_8_), .R(reset_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_730 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_12__31_0__7_), .Q(w_mem_inst_w_mem_12__7_), .R(reset_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_731 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_12__31_0__8_), .Q(w_mem_inst_w_mem_12__8_), .R(reset_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_732 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_12__31_0__9_), .Q(w_mem_inst_w_mem_12__9_), .R(reset_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_733 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_12__31_0__10_), .Q(w_mem_inst_w_mem_12__10_), .R(reset_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_734 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_12__31_0__11_), .Q(w_mem_inst_w_mem_12__11_), .R(reset_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_735 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_12__31_0__12_), .Q(w_mem_inst_w_mem_12__12_), .R(reset_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_736 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_12__31_0__13_), .Q(w_mem_inst_w_mem_12__13_), .R(reset_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_737 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_12__31_0__14_), .Q(w_mem_inst_w_mem_12__14_), .R(reset_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_738 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_12__31_0__15_), .Q(w_mem_inst_w_mem_12__15_), .R(reset_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_739 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_12__31_0__16_), .Q(w_mem_inst_w_mem_12__16_), .R(reset_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_74 ( .CLK(clk_bF_buf15), .D(c_reg_9__FF_INPUT), .Q(c_reg_9_), .R(reset_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_740 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_12__31_0__17_), .Q(w_mem_inst_w_mem_12__17_), .R(reset_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_741 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_12__31_0__18_), .Q(w_mem_inst_w_mem_12__18_), .R(reset_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_742 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_12__31_0__19_), .Q(w_mem_inst_w_mem_12__19_), .R(reset_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_743 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_12__31_0__20_), .Q(w_mem_inst_w_mem_12__20_), .R(reset_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_744 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_12__31_0__21_), .Q(w_mem_inst_w_mem_12__21_), .R(reset_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_745 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_12__31_0__22_), .Q(w_mem_inst_w_mem_12__22_), .R(reset_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_746 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_12__31_0__23_), .Q(w_mem_inst_w_mem_12__23_), .R(reset_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_747 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_12__31_0__24_), .Q(w_mem_inst_w_mem_12__24_), .R(reset_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_748 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_12__31_0__25_), .Q(w_mem_inst_w_mem_12__25_), .R(reset_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_749 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_12__31_0__26_), .Q(w_mem_inst_w_mem_12__26_), .R(reset_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_75 ( .CLK(clk_bF_buf14), .D(c_reg_10__FF_INPUT), .Q(c_reg_10_), .R(reset_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_750 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_12__31_0__27_), .Q(w_mem_inst_w_mem_12__27_), .R(reset_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_751 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_12__31_0__28_), .Q(w_mem_inst_w_mem_12__28_), .R(reset_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_752 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_12__31_0__29_), .Q(w_mem_inst_w_mem_12__29_), .R(reset_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_753 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_12__31_0__30_), .Q(w_mem_inst_w_mem_12__30_), .R(reset_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_754 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_12__31_0__31_), .Q(w_mem_inst_w_mem_12__31_), .R(reset_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_755 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_13__31_0__0_), .Q(w_mem_inst_w_mem_13__0_), .R(reset_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_756 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_13__31_0__1_), .Q(w_mem_inst_w_mem_13__1_), .R(reset_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_757 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_13__31_0__2_), .Q(w_mem_inst_w_mem_13__2_), .R(reset_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_758 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_13__31_0__3_), .Q(w_mem_inst_w_mem_13__3_), .R(reset_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_759 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_13__31_0__4_), .Q(w_mem_inst_w_mem_13__4_), .R(reset_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_76 ( .CLK(clk_bF_buf13), .D(c_reg_11__FF_INPUT), .Q(c_reg_11_), .R(reset_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_760 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_13__31_0__5_), .Q(w_mem_inst_w_mem_13__5_), .R(reset_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_761 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_13__31_0__6_), .Q(w_mem_inst_w_mem_13__6_), .R(reset_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_762 ( .CLK(clk_bF_buf39), .D(w_mem_inst__0w_mem_13__31_0__7_), .Q(w_mem_inst_w_mem_13__7_), .R(reset_n_bF_buf39), .S(1'b1) );
  DFFSR DFFSR_763 ( .CLK(clk_bF_buf38), .D(w_mem_inst__0w_mem_13__31_0__8_), .Q(w_mem_inst_w_mem_13__8_), .R(reset_n_bF_buf38), .S(1'b1) );
  DFFSR DFFSR_764 ( .CLK(clk_bF_buf37), .D(w_mem_inst__0w_mem_13__31_0__9_), .Q(w_mem_inst_w_mem_13__9_), .R(reset_n_bF_buf37), .S(1'b1) );
  DFFSR DFFSR_765 ( .CLK(clk_bF_buf36), .D(w_mem_inst__0w_mem_13__31_0__10_), .Q(w_mem_inst_w_mem_13__10_), .R(reset_n_bF_buf36), .S(1'b1) );
  DFFSR DFFSR_766 ( .CLK(clk_bF_buf35), .D(w_mem_inst__0w_mem_13__31_0__11_), .Q(w_mem_inst_w_mem_13__11_), .R(reset_n_bF_buf35), .S(1'b1) );
  DFFSR DFFSR_767 ( .CLK(clk_bF_buf34), .D(w_mem_inst__0w_mem_13__31_0__12_), .Q(w_mem_inst_w_mem_13__12_), .R(reset_n_bF_buf34), .S(1'b1) );
  DFFSR DFFSR_768 ( .CLK(clk_bF_buf33), .D(w_mem_inst__0w_mem_13__31_0__13_), .Q(w_mem_inst_w_mem_13__13_), .R(reset_n_bF_buf33), .S(1'b1) );
  DFFSR DFFSR_769 ( .CLK(clk_bF_buf32), .D(w_mem_inst__0w_mem_13__31_0__14_), .Q(w_mem_inst_w_mem_13__14_), .R(reset_n_bF_buf32), .S(1'b1) );
  DFFSR DFFSR_77 ( .CLK(clk_bF_buf12), .D(c_reg_12__FF_INPUT), .Q(c_reg_12_), .R(reset_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_770 ( .CLK(clk_bF_buf31), .D(w_mem_inst__0w_mem_13__31_0__15_), .Q(w_mem_inst_w_mem_13__15_), .R(reset_n_bF_buf31), .S(1'b1) );
  DFFSR DFFSR_771 ( .CLK(clk_bF_buf30), .D(w_mem_inst__0w_mem_13__31_0__16_), .Q(w_mem_inst_w_mem_13__16_), .R(reset_n_bF_buf30), .S(1'b1) );
  DFFSR DFFSR_772 ( .CLK(clk_bF_buf29), .D(w_mem_inst__0w_mem_13__31_0__17_), .Q(w_mem_inst_w_mem_13__17_), .R(reset_n_bF_buf29), .S(1'b1) );
  DFFSR DFFSR_773 ( .CLK(clk_bF_buf28), .D(w_mem_inst__0w_mem_13__31_0__18_), .Q(w_mem_inst_w_mem_13__18_), .R(reset_n_bF_buf28), .S(1'b1) );
  DFFSR DFFSR_774 ( .CLK(clk_bF_buf27), .D(w_mem_inst__0w_mem_13__31_0__19_), .Q(w_mem_inst_w_mem_13__19_), .R(reset_n_bF_buf27), .S(1'b1) );
  DFFSR DFFSR_775 ( .CLK(clk_bF_buf26), .D(w_mem_inst__0w_mem_13__31_0__20_), .Q(w_mem_inst_w_mem_13__20_), .R(reset_n_bF_buf26), .S(1'b1) );
  DFFSR DFFSR_776 ( .CLK(clk_bF_buf25), .D(w_mem_inst__0w_mem_13__31_0__21_), .Q(w_mem_inst_w_mem_13__21_), .R(reset_n_bF_buf25), .S(1'b1) );
  DFFSR DFFSR_777 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_mem_13__31_0__22_), .Q(w_mem_inst_w_mem_13__22_), .R(reset_n_bF_buf24), .S(1'b1) );
  DFFSR DFFSR_778 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_mem_13__31_0__23_), .Q(w_mem_inst_w_mem_13__23_), .R(reset_n_bF_buf23), .S(1'b1) );
  DFFSR DFFSR_779 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_mem_13__31_0__24_), .Q(w_mem_inst_w_mem_13__24_), .R(reset_n_bF_buf22), .S(1'b1) );
  DFFSR DFFSR_78 ( .CLK(clk_bF_buf11), .D(c_reg_13__FF_INPUT), .Q(c_reg_13_), .R(reset_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_780 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_mem_13__31_0__25_), .Q(w_mem_inst_w_mem_13__25_), .R(reset_n_bF_buf21), .S(1'b1) );
  DFFSR DFFSR_781 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_mem_13__31_0__26_), .Q(w_mem_inst_w_mem_13__26_), .R(reset_n_bF_buf20), .S(1'b1) );
  DFFSR DFFSR_782 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_mem_13__31_0__27_), .Q(w_mem_inst_w_mem_13__27_), .R(reset_n_bF_buf19), .S(1'b1) );
  DFFSR DFFSR_783 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_mem_13__31_0__28_), .Q(w_mem_inst_w_mem_13__28_), .R(reset_n_bF_buf18), .S(1'b1) );
  DFFSR DFFSR_784 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_13__31_0__29_), .Q(w_mem_inst_w_mem_13__29_), .R(reset_n_bF_buf17), .S(1'b1) );
  DFFSR DFFSR_785 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_13__31_0__30_), .Q(w_mem_inst_w_mem_13__30_), .R(reset_n_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_786 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_13__31_0__31_), .Q(w_mem_inst_w_mem_13__31_), .R(reset_n_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_787 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_14__31_0__0_), .Q(w_mem_inst_w_mem_14__0_), .R(reset_n_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_788 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_14__31_0__1_), .Q(w_mem_inst_w_mem_14__1_), .R(reset_n_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_789 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_14__31_0__2_), .Q(w_mem_inst_w_mem_14__2_), .R(reset_n_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_79 ( .CLK(clk_bF_buf10), .D(c_reg_14__FF_INPUT), .Q(c_reg_14_), .R(reset_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_790 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_14__31_0__3_), .Q(w_mem_inst_w_mem_14__3_), .R(reset_n_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_791 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_14__31_0__4_), .Q(w_mem_inst_w_mem_14__4_), .R(reset_n_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_792 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_14__31_0__5_), .Q(w_mem_inst_w_mem_14__5_), .R(reset_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_793 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_14__31_0__6_), .Q(w_mem_inst_w_mem_14__6_), .R(reset_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_794 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_14__31_0__7_), .Q(w_mem_inst_w_mem_14__7_), .R(reset_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_795 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_14__31_0__8_), .Q(w_mem_inst_w_mem_14__8_), .R(reset_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_796 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_14__31_0__9_), .Q(w_mem_inst_w_mem_14__9_), .R(reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_797 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_14__31_0__10_), .Q(w_mem_inst_w_mem_14__10_), .R(reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_798 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_14__31_0__11_), .Q(w_mem_inst_w_mem_14__11_), .R(reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_799 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_14__31_0__12_), .Q(w_mem_inst_w_mem_14__12_), .R(reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_8 ( .CLK(clk_bF_buf81), .D(a_reg_7__FF_INPUT), .Q(a_reg_7_), .R(reset_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_80 ( .CLK(clk_bF_buf9), .D(c_reg_15__FF_INPUT), .Q(c_reg_15_), .R(reset_n_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_800 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_14__31_0__13_), .Q(w_mem_inst_w_mem_14__13_), .R(reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_801 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_14__31_0__14_), .Q(w_mem_inst_w_mem_14__14_), .R(reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_802 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_14__31_0__15_), .Q(w_mem_inst_w_mem_14__15_), .R(reset_n_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_803 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_14__31_0__16_), .Q(w_mem_inst_w_mem_14__16_), .R(reset_n_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_804 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_14__31_0__17_), .Q(w_mem_inst_w_mem_14__17_), .R(reset_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_805 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_14__31_0__18_), .Q(w_mem_inst_w_mem_14__18_), .R(reset_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_806 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_14__31_0__19_), .Q(w_mem_inst_w_mem_14__19_), .R(reset_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_807 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_14__31_0__20_), .Q(w_mem_inst_w_mem_14__20_), .R(reset_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_808 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_14__31_0__21_), .Q(w_mem_inst_w_mem_14__21_), .R(reset_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_809 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_14__31_0__22_), .Q(w_mem_inst_w_mem_14__22_), .R(reset_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_81 ( .CLK(clk_bF_buf8), .D(c_reg_16__FF_INPUT), .Q(c_reg_16_), .R(reset_n_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_810 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_14__31_0__23_), .Q(w_mem_inst_w_mem_14__23_), .R(reset_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_811 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_14__31_0__24_), .Q(w_mem_inst_w_mem_14__24_), .R(reset_n_bF_buf79), .S(1'b1) );
  DFFSR DFFSR_812 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_14__31_0__25_), .Q(w_mem_inst_w_mem_14__25_), .R(reset_n_bF_buf78), .S(1'b1) );
  DFFSR DFFSR_813 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_14__31_0__26_), .Q(w_mem_inst_w_mem_14__26_), .R(reset_n_bF_buf77), .S(1'b1) );
  DFFSR DFFSR_814 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_14__31_0__27_), .Q(w_mem_inst_w_mem_14__27_), .R(reset_n_bF_buf76), .S(1'b1) );
  DFFSR DFFSR_815 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_14__31_0__28_), .Q(w_mem_inst_w_mem_14__28_), .R(reset_n_bF_buf75), .S(1'b1) );
  DFFSR DFFSR_816 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_14__31_0__29_), .Q(w_mem_inst_w_mem_14__29_), .R(reset_n_bF_buf74), .S(1'b1) );
  DFFSR DFFSR_817 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_14__31_0__30_), .Q(w_mem_inst_w_mem_14__30_), .R(reset_n_bF_buf73), .S(1'b1) );
  DFFSR DFFSR_818 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_14__31_0__31_), .Q(w_mem_inst_w_mem_14__31_), .R(reset_n_bF_buf72), .S(1'b1) );
  DFFSR DFFSR_819 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_15__31_0__0_), .Q(w_mem_inst_w_mem_15__0_), .R(reset_n_bF_buf71), .S(1'b1) );
  DFFSR DFFSR_82 ( .CLK(clk_bF_buf7), .D(c_reg_17__FF_INPUT), .Q(c_reg_17_), .R(reset_n_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_820 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_15__31_0__1_), .Q(w_mem_inst_w_mem_15__1_), .R(reset_n_bF_buf70), .S(1'b1) );
  DFFSR DFFSR_821 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_15__31_0__2_), .Q(w_mem_inst_w_mem_15__2_), .R(reset_n_bF_buf69), .S(1'b1) );
  DFFSR DFFSR_822 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_15__31_0__3_), .Q(w_mem_inst_w_mem_15__3_), .R(reset_n_bF_buf68), .S(1'b1) );
  DFFSR DFFSR_823 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_15__31_0__4_), .Q(w_mem_inst_w_mem_15__4_), .R(reset_n_bF_buf67), .S(1'b1) );
  DFFSR DFFSR_824 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_15__31_0__5_), .Q(w_mem_inst_w_mem_15__5_), .R(reset_n_bF_buf66), .S(1'b1) );
  DFFSR DFFSR_825 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_15__31_0__6_), .Q(w_mem_inst_w_mem_15__6_), .R(reset_n_bF_buf65), .S(1'b1) );
  DFFSR DFFSR_826 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_15__31_0__7_), .Q(w_mem_inst_w_mem_15__7_), .R(reset_n_bF_buf64), .S(1'b1) );
  DFFSR DFFSR_827 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_15__31_0__8_), .Q(w_mem_inst_w_mem_15__8_), .R(reset_n_bF_buf63), .S(1'b1) );
  DFFSR DFFSR_828 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_15__31_0__9_), .Q(w_mem_inst_w_mem_15__9_), .R(reset_n_bF_buf62), .S(1'b1) );
  DFFSR DFFSR_829 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_15__31_0__10_), .Q(w_mem_inst_w_mem_15__10_), .R(reset_n_bF_buf61), .S(1'b1) );
  DFFSR DFFSR_83 ( .CLK(clk_bF_buf6), .D(c_reg_18__FF_INPUT), .Q(c_reg_18_), .R(reset_n_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_830 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_15__31_0__11_), .Q(w_mem_inst_w_mem_15__11_), .R(reset_n_bF_buf60), .S(1'b1) );
  DFFSR DFFSR_831 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_15__31_0__12_), .Q(w_mem_inst_w_mem_15__12_), .R(reset_n_bF_buf59), .S(1'b1) );
  DFFSR DFFSR_832 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_15__31_0__13_), .Q(w_mem_inst_w_mem_15__13_), .R(reset_n_bF_buf58), .S(1'b1) );
  DFFSR DFFSR_833 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_15__31_0__14_), .Q(w_mem_inst_w_mem_15__14_), .R(reset_n_bF_buf57), .S(1'b1) );
  DFFSR DFFSR_834 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_15__31_0__15_), .Q(w_mem_inst_w_mem_15__15_), .R(reset_n_bF_buf56), .S(1'b1) );
  DFFSR DFFSR_835 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_15__31_0__16_), .Q(w_mem_inst_w_mem_15__16_), .R(reset_n_bF_buf55), .S(1'b1) );
  DFFSR DFFSR_836 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_15__31_0__17_), .Q(w_mem_inst_w_mem_15__17_), .R(reset_n_bF_buf54), .S(1'b1) );
  DFFSR DFFSR_837 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_15__31_0__18_), .Q(w_mem_inst_w_mem_15__18_), .R(reset_n_bF_buf53), .S(1'b1) );
  DFFSR DFFSR_838 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_15__31_0__19_), .Q(w_mem_inst_w_mem_15__19_), .R(reset_n_bF_buf52), .S(1'b1) );
  DFFSR DFFSR_839 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_15__31_0__20_), .Q(w_mem_inst_w_mem_15__20_), .R(reset_n_bF_buf51), .S(1'b1) );
  DFFSR DFFSR_84 ( .CLK(clk_bF_buf5), .D(c_reg_19__FF_INPUT), .Q(c_reg_19_), .R(reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_840 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_15__31_0__21_), .Q(w_mem_inst_w_mem_15__21_), .R(reset_n_bF_buf50), .S(1'b1) );
  DFFSR DFFSR_841 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_15__31_0__22_), .Q(w_mem_inst_w_mem_15__22_), .R(reset_n_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_842 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_15__31_0__23_), .Q(w_mem_inst_w_mem_15__23_), .R(reset_n_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_843 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_15__31_0__24_), .Q(w_mem_inst_w_mem_15__24_), .R(reset_n_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_844 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_15__31_0__25_), .Q(w_mem_inst_w_mem_15__25_), .R(reset_n_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_845 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_15__31_0__26_), .Q(w_mem_inst_w_mem_15__26_), .R(reset_n_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_846 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_15__31_0__27_), .Q(w_mem_inst_w_mem_15__27_), .R(reset_n_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_847 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_15__31_0__28_), .Q(w_mem_inst_w_mem_15__28_), .R(reset_n_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_848 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_15__31_0__29_), .Q(w_mem_inst_w_mem_15__29_), .R(reset_n_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_849 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_15__31_0__30_), .Q(w_mem_inst_w_mem_15__30_), .R(reset_n_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_85 ( .CLK(clk_bF_buf4), .D(c_reg_20__FF_INPUT), .Q(c_reg_20_), .R(reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_850 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_15__31_0__31_), .Q(w_mem_inst_w_mem_15__31_), .R(reset_n_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_86 ( .CLK(clk_bF_buf3), .D(c_reg_21__FF_INPUT), .Q(c_reg_21_), .R(reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_87 ( .CLK(clk_bF_buf2), .D(c_reg_22__FF_INPUT), .Q(c_reg_22_), .R(reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_88 ( .CLK(clk_bF_buf1), .D(c_reg_23__FF_INPUT), .Q(c_reg_23_), .R(reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_89 ( .CLK(clk_bF_buf0), .D(c_reg_24__FF_INPUT), .Q(c_reg_24_), .R(reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_9 ( .CLK(clk_bF_buf80), .D(a_reg_8__FF_INPUT), .Q(a_reg_8_), .R(reset_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_90 ( .CLK(clk_bF_buf88), .D(c_reg_25__FF_INPUT), .Q(c_reg_25_), .R(reset_n_bF_buf88), .S(1'b1) );
  DFFSR DFFSR_91 ( .CLK(clk_bF_buf87), .D(c_reg_26__FF_INPUT), .Q(c_reg_26_), .R(reset_n_bF_buf87), .S(1'b1) );
  DFFSR DFFSR_92 ( .CLK(clk_bF_buf86), .D(c_reg_27__FF_INPUT), .Q(c_reg_27_), .R(reset_n_bF_buf86), .S(1'b1) );
  DFFSR DFFSR_93 ( .CLK(clk_bF_buf85), .D(c_reg_28__FF_INPUT), .Q(c_reg_28_), .R(reset_n_bF_buf85), .S(1'b1) );
  DFFSR DFFSR_94 ( .CLK(clk_bF_buf84), .D(c_reg_29__FF_INPUT), .Q(c_reg_29_), .R(reset_n_bF_buf84), .S(1'b1) );
  DFFSR DFFSR_95 ( .CLK(clk_bF_buf83), .D(c_reg_30__FF_INPUT), .Q(c_reg_30_), .R(reset_n_bF_buf83), .S(1'b1) );
  DFFSR DFFSR_96 ( .CLK(clk_bF_buf82), .D(c_reg_31__FF_INPUT), .Q(c_reg_31_), .R(reset_n_bF_buf82), .S(1'b1) );
  DFFSR DFFSR_97 ( .CLK(clk_bF_buf81), .D(d_reg_0__FF_INPUT), .Q(d_reg_0_), .R(reset_n_bF_buf81), .S(1'b1) );
  DFFSR DFFSR_98 ( .CLK(clk_bF_buf80), .D(d_reg_1__FF_INPUT), .Q(d_reg_1_), .R(reset_n_bF_buf80), .S(1'b1) );
  DFFSR DFFSR_99 ( .CLK(clk_bF_buf79), .D(d_reg_2__FF_INPUT), .Q(d_reg_2_), .R(reset_n_bF_buf79), .S(1'b1) );
  INVX1 INVX1_1 ( .A(_abc_15724_n698), .Y(_abc_15724_n700) );
  INVX1 INVX1_10 ( .A(_abc_15724_n733), .Y(_abc_15724_n734) );
  INVX1 INVX1_100 ( .A(_abc_15724_n1256), .Y(_abc_15724_n1273) );
  INVX1 INVX1_1000 ( .A(_abc_15724_n6053), .Y(_abc_15724_n6054) );
  INVX1 INVX1_1001 ( .A(_abc_15724_n6055), .Y(_abc_15724_n6056) );
  INVX1 INVX1_1002 ( .A(d_reg_31_), .Y(_abc_15724_n6057) );
  INVX1 INVX1_1003 ( .A(_abc_15724_n6065), .Y(_abc_15724_n6066) );
  INVX1 INVX1_1004 ( .A(_abc_15724_n6071), .Y(_abc_15724_n6072) );
  INVX1 INVX1_1005 ( .A(_abc_15724_n6077), .Y(_abc_15724_n6078) );
  INVX1 INVX1_1006 ( .A(_abc_15724_n6080), .Y(_abc_15724_n6081) );
  INVX1 INVX1_1007 ( .A(_abc_15724_n6083), .Y(_abc_15724_n6084) );
  INVX1 INVX1_1008 ( .A(_abc_15724_n6085), .Y(_abc_15724_n6086) );
  INVX1 INVX1_1009 ( .A(_abc_15724_n6074), .Y(_abc_15724_n6090) );
  INVX1 INVX1_101 ( .A(_abc_15724_n1276_1), .Y(_abc_15724_n1277) );
  INVX1 INVX1_1010 ( .A(_abc_15724_n6088), .Y(_abc_15724_n6091) );
  INVX1 INVX1_1011 ( .A(_abc_15724_n6093), .Y(_abc_15724_n6094) );
  INVX1 INVX1_1012 ( .A(_abc_15724_n6097), .Y(_abc_15724_n6098) );
  INVX1 INVX1_1013 ( .A(_abc_15724_n6102), .Y(_abc_15724_n6103) );
  INVX1 INVX1_1014 ( .A(_abc_15724_n6105), .Y(_abc_15724_n6106) );
  INVX1 INVX1_1015 ( .A(_abc_15724_n6117), .Y(_abc_15724_n6118) );
  INVX1 INVX1_1016 ( .A(_abc_15724_n6120), .Y(_abc_15724_n6123) );
  INVX1 INVX1_1017 ( .A(_abc_15724_n2988), .Y(_abc_15724_n6128) );
  INVX1 INVX1_1018 ( .A(round_ctr_reg_0_), .Y(_abc_15724_n6134) );
  INVX1 INVX1_1019 ( .A(_abc_15724_n6119), .Y(_abc_15724_n6139) );
  INVX1 INVX1_102 ( .A(_abc_15724_n1279), .Y(_abc_15724_n1280) );
  INVX1 INVX1_1020 ( .A(_abc_15724_n6145), .Y(_abc_15724_n6146) );
  INVX1 INVX1_1021 ( .A(_abc_15724_n6156), .Y(_abc_15724_n6157) );
  INVX1 INVX1_1022 ( .A(_abc_15724_n2994_bF_buf7), .Y(_abc_15724_n6158) );
  INVX1 INVX1_1023 ( .A(_abc_15724_n6162), .Y(_abc_15724_n6163) );
  INVX1 INVX1_1024 ( .A(_abc_15724_n6172), .Y(_abc_15724_n6173) );
  INVX1 INVX1_1025 ( .A(_abc_15724_n792), .Y(_abc_15724_n6175) );
  INVX1 INVX1_1026 ( .A(_abc_15724_n802), .Y(_abc_15724_n6186) );
  INVX1 INVX1_1027 ( .A(_abc_15724_n787), .Y(_abc_15724_n6192) );
  INVX1 INVX1_1028 ( .A(_abc_15724_n803_1), .Y(_abc_15724_n6195) );
  INVX1 INVX1_1029 ( .A(_abc_15724_n6193), .Y(_abc_15724_n6196) );
  INVX1 INVX1_103 ( .A(_abc_15724_n1286), .Y(_abc_15724_n1287_1) );
  INVX1 INVX1_1030 ( .A(_abc_15724_n809), .Y(_abc_15724_n6202) );
  INVX1 INVX1_1031 ( .A(_abc_15724_n810), .Y(_abc_15724_n6209) );
  INVX1 INVX1_1032 ( .A(_abc_15724_n784), .Y(_abc_15724_n6210) );
  INVX1 INVX1_1033 ( .A(_abc_15724_n6211), .Y(_abc_15724_n6213) );
  INVX1 INVX1_1034 ( .A(_abc_15724_n6219), .Y(_abc_15724_n6220) );
  INVX1 INVX1_1035 ( .A(_abc_15724_n6225), .Y(_abc_15724_n6226) );
  INVX1 INVX1_1036 ( .A(_abc_15724_n779_1), .Y(_abc_15724_n6228) );
  INVX1 INVX1_1037 ( .A(_abc_15724_n6235), .Y(_abc_15724_n6236) );
  INVX1 INVX1_1038 ( .A(_abc_15724_n816), .Y(_abc_15724_n6243) );
  INVX1 INVX1_1039 ( .A(_abc_15724_n6241), .Y(_abc_15724_n6244) );
  INVX1 INVX1_104 ( .A(_abc_15724_n1284_1), .Y(_abc_15724_n1290) );
  INVX1 INVX1_1040 ( .A(_abc_15724_n6254), .Y(_abc_15724_n6255) );
  INVX1 INVX1_1041 ( .A(_abc_15724_n761), .Y(_abc_15724_n6261) );
  INVX1 INVX1_1042 ( .A(_abc_15724_n6259), .Y(_abc_15724_n6262) );
  INVX1 INVX1_1043 ( .A(_abc_15724_n6270), .Y(_abc_15724_n6271) );
  INVX1 INVX1_1044 ( .A(_abc_15724_n6275), .Y(_abc_15724_n6276) );
  INVX1 INVX1_1045 ( .A(_abc_15724_n750), .Y(_abc_15724_n6278) );
  INVX1 INVX1_1046 ( .A(_abc_15724_n6287), .Y(_abc_15724_n6288) );
  INVX1 INVX1_1047 ( .A(_abc_15724_n732), .Y(_abc_15724_n6295) );
  INVX1 INVX1_1048 ( .A(_abc_15724_n6293), .Y(_abc_15724_n6296) );
  INVX1 INVX1_1049 ( .A(_abc_15724_n6304), .Y(_abc_15724_n6305) );
  INVX1 INVX1_105 ( .A(_abc_15724_n1288), .Y(_abc_15724_n1291) );
  INVX1 INVX1_1050 ( .A(_abc_15724_n6309), .Y(_abc_15724_n6310) );
  INVX1 INVX1_1051 ( .A(_abc_15724_n6321), .Y(_abc_15724_n6322) );
  INVX1 INVX1_1052 ( .A(_abc_15724_n708_1), .Y(_abc_15724_n6326) );
  INVX1 INVX1_1053 ( .A(_abc_15724_n6327), .Y(_abc_15724_n6328) );
  INVX1 INVX1_1054 ( .A(_abc_15724_n6335), .Y(_abc_15724_n6336) );
  INVX1 INVX1_1055 ( .A(_abc_15724_n6343), .Y(_abc_15724_n6344) );
  INVX1 INVX1_1056 ( .A(_abc_15724_n702), .Y(_abc_15724_n6346) );
  INVX1 INVX1_1057 ( .A(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_21378_n1588) );
  INVX1 INVX1_1058 ( .A(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_21378_n1590) );
  INVX1 INVX1_1059 ( .A(w_mem_inst__abc_21378_n1592), .Y(w_mem_inst__abc_21378_n1593) );
  INVX1 INVX1_106 ( .A(_abc_15724_n1298), .Y(_abc_15724_n1299_1) );
  INVX1 INVX1_1060 ( .A(w_mem_inst__abc_21378_n1595), .Y(w_mem_inst__abc_21378_n1596) );
  INVX1 INVX1_1061 ( .A(w_mem_inst__abc_21378_n1597), .Y(w_mem_inst__abc_21378_n1599_1) );
  INVX1 INVX1_1062 ( .A(w_mem_inst_w_ctr_reg_3_), .Y(w_mem_inst__abc_21378_n1607_1) );
  INVX1 INVX1_1063 ( .A(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_21378_n1608) );
  INVX1 INVX1_1064 ( .A(w_mem_inst_w_ctr_reg_1_), .Y(w_mem_inst__abc_21378_n1614_1) );
  INVX1 INVX1_1065 ( .A(w_mem_inst_w_ctr_reg_0_), .Y(w_mem_inst__abc_21378_n1623_1) );
  INVX1 INVX1_1066 ( .A(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_21378_n1664) );
  INVX1 INVX1_1067 ( .A(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_21378_n1666_1) );
  INVX1 INVX1_1068 ( .A(w_mem_inst__abc_21378_n1668), .Y(w_mem_inst__abc_21378_n1669) );
  INVX1 INVX1_1069 ( .A(w_mem_inst__abc_21378_n1671_1), .Y(w_mem_inst__abc_21378_n1672) );
  INVX1 INVX1_107 ( .A(_abc_15724_n1302), .Y(_abc_15724_n1303) );
  INVX1 INVX1_1070 ( .A(w_mem_inst__abc_21378_n1673), .Y(w_mem_inst__abc_21378_n1675_1) );
  INVX1 INVX1_1071 ( .A(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_21378_n1712) );
  INVX1 INVX1_1072 ( .A(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_21378_n1714_1) );
  INVX1 INVX1_1073 ( .A(w_mem_inst__abc_21378_n1716), .Y(w_mem_inst__abc_21378_n1717) );
  INVX1 INVX1_1074 ( .A(w_mem_inst__abc_21378_n1719_1), .Y(w_mem_inst__abc_21378_n1720) );
  INVX1 INVX1_1075 ( .A(w_mem_inst__abc_21378_n1721), .Y(w_mem_inst__abc_21378_n1723_1) );
  INVX1 INVX1_1076 ( .A(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_21378_n1760) );
  INVX1 INVX1_1077 ( .A(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_21378_n1762_1) );
  INVX1 INVX1_1078 ( .A(w_mem_inst__abc_21378_n1764), .Y(w_mem_inst__abc_21378_n1765) );
  INVX1 INVX1_1079 ( .A(w_mem_inst__abc_21378_n1767_1), .Y(w_mem_inst__abc_21378_n1768) );
  INVX1 INVX1_108 ( .A(_abc_15724_n1304), .Y(_abc_15724_n1305_1) );
  INVX1 INVX1_1080 ( .A(w_mem_inst__abc_21378_n1769), .Y(w_mem_inst__abc_21378_n1771_1) );
  INVX1 INVX1_1081 ( .A(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_21378_n1808) );
  INVX1 INVX1_1082 ( .A(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_21378_n1810_1) );
  INVX1 INVX1_1083 ( .A(w_mem_inst__abc_21378_n1812), .Y(w_mem_inst__abc_21378_n1813) );
  INVX1 INVX1_1084 ( .A(w_mem_inst__abc_21378_n1815_1), .Y(w_mem_inst__abc_21378_n1816) );
  INVX1 INVX1_1085 ( .A(w_mem_inst__abc_21378_n1817), .Y(w_mem_inst__abc_21378_n1819_1) );
  INVX1 INVX1_1086 ( .A(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_21378_n1856) );
  INVX1 INVX1_1087 ( .A(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_21378_n1858_1) );
  INVX1 INVX1_1088 ( .A(w_mem_inst__abc_21378_n1860), .Y(w_mem_inst__abc_21378_n1861) );
  INVX1 INVX1_1089 ( .A(w_mem_inst__abc_21378_n1863_1), .Y(w_mem_inst__abc_21378_n1864) );
  INVX1 INVX1_109 ( .A(_abc_15724_n1311), .Y(_abc_15724_n1312) );
  INVX1 INVX1_1090 ( .A(w_mem_inst__abc_21378_n1865), .Y(w_mem_inst__abc_21378_n1867_1) );
  INVX1 INVX1_1091 ( .A(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_21378_n1904) );
  INVX1 INVX1_1092 ( .A(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_21378_n1906_1) );
  INVX1 INVX1_1093 ( .A(w_mem_inst__abc_21378_n1908), .Y(w_mem_inst__abc_21378_n1909) );
  INVX1 INVX1_1094 ( .A(w_mem_inst__abc_21378_n1911_1), .Y(w_mem_inst__abc_21378_n1912) );
  INVX1 INVX1_1095 ( .A(w_mem_inst__abc_21378_n1913), .Y(w_mem_inst__abc_21378_n1915_1) );
  INVX1 INVX1_1096 ( .A(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_21378_n1952) );
  INVX1 INVX1_1097 ( .A(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_21378_n1954_1) );
  INVX1 INVX1_1098 ( .A(w_mem_inst__abc_21378_n1956), .Y(w_mem_inst__abc_21378_n1957) );
  INVX1 INVX1_1099 ( .A(w_mem_inst__abc_21378_n1959_1), .Y(w_mem_inst__abc_21378_n1960) );
  INVX1 INVX1_11 ( .A(_abc_15724_n739_1), .Y(_abc_15724_n740) );
  INVX1 INVX1_110 ( .A(_abc_15724_n1315), .Y(_abc_15724_n1316) );
  INVX1 INVX1_1100 ( .A(w_mem_inst__abc_21378_n1961), .Y(w_mem_inst__abc_21378_n1963_1) );
  INVX1 INVX1_1101 ( .A(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_21378_n2000) );
  INVX1 INVX1_1102 ( .A(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_21378_n2002_1) );
  INVX1 INVX1_1103 ( .A(w_mem_inst__abc_21378_n2004), .Y(w_mem_inst__abc_21378_n2005) );
  INVX1 INVX1_1104 ( .A(w_mem_inst__abc_21378_n2007_1), .Y(w_mem_inst__abc_21378_n2008) );
  INVX1 INVX1_1105 ( .A(w_mem_inst__abc_21378_n2009), .Y(w_mem_inst__abc_21378_n2011_1) );
  INVX1 INVX1_1106 ( .A(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_21378_n2048) );
  INVX1 INVX1_1107 ( .A(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_21378_n2050_1) );
  INVX1 INVX1_1108 ( .A(w_mem_inst__abc_21378_n2052), .Y(w_mem_inst__abc_21378_n2053) );
  INVX1 INVX1_1109 ( .A(w_mem_inst__abc_21378_n2055_1), .Y(w_mem_inst__abc_21378_n2056) );
  INVX1 INVX1_111 ( .A(_abc_15724_n1324), .Y(_abc_15724_n1325) );
  INVX1 INVX1_1110 ( .A(w_mem_inst__abc_21378_n2057), .Y(w_mem_inst__abc_21378_n2059_1) );
  INVX1 INVX1_1111 ( .A(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_21378_n2096) );
  INVX1 INVX1_1112 ( .A(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_21378_n2098_1) );
  INVX1 INVX1_1113 ( .A(w_mem_inst__abc_21378_n2100), .Y(w_mem_inst__abc_21378_n2101) );
  INVX1 INVX1_1114 ( .A(w_mem_inst__abc_21378_n2103_1), .Y(w_mem_inst__abc_21378_n2104) );
  INVX1 INVX1_1115 ( .A(w_mem_inst__abc_21378_n2105), .Y(w_mem_inst__abc_21378_n2107_1) );
  INVX1 INVX1_1116 ( .A(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_21378_n2144) );
  INVX1 INVX1_1117 ( .A(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_21378_n2146_1) );
  INVX1 INVX1_1118 ( .A(w_mem_inst__abc_21378_n2148), .Y(w_mem_inst__abc_21378_n2149) );
  INVX1 INVX1_1119 ( .A(w_mem_inst__abc_21378_n2151_1), .Y(w_mem_inst__abc_21378_n2152) );
  INVX1 INVX1_112 ( .A(_abc_15724_n1322), .Y(_abc_15724_n1328) );
  INVX1 INVX1_1120 ( .A(w_mem_inst__abc_21378_n2153), .Y(w_mem_inst__abc_21378_n2155_1) );
  INVX1 INVX1_1121 ( .A(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_21378_n2192) );
  INVX1 INVX1_1122 ( .A(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_21378_n2194_1) );
  INVX1 INVX1_1123 ( .A(w_mem_inst__abc_21378_n2196), .Y(w_mem_inst__abc_21378_n2197) );
  INVX1 INVX1_1124 ( .A(w_mem_inst__abc_21378_n2199_1), .Y(w_mem_inst__abc_21378_n2200) );
  INVX1 INVX1_1125 ( .A(w_mem_inst__abc_21378_n2201), .Y(w_mem_inst__abc_21378_n2203_1) );
  INVX1 INVX1_1126 ( .A(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_21378_n2240) );
  INVX1 INVX1_1127 ( .A(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_21378_n2242_1) );
  INVX1 INVX1_1128 ( .A(w_mem_inst__abc_21378_n2244), .Y(w_mem_inst__abc_21378_n2245) );
  INVX1 INVX1_1129 ( .A(w_mem_inst__abc_21378_n2247_1), .Y(w_mem_inst__abc_21378_n2248) );
  INVX1 INVX1_113 ( .A(_abc_15724_n1326), .Y(_abc_15724_n1329_1) );
  INVX1 INVX1_1130 ( .A(w_mem_inst__abc_21378_n2249), .Y(w_mem_inst__abc_21378_n2251_1) );
  INVX1 INVX1_1131 ( .A(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_21378_n2288) );
  INVX1 INVX1_1132 ( .A(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_21378_n2290_1) );
  INVX1 INVX1_1133 ( .A(w_mem_inst__abc_21378_n2292), .Y(w_mem_inst__abc_21378_n2293) );
  INVX1 INVX1_1134 ( .A(w_mem_inst__abc_21378_n2295_1), .Y(w_mem_inst__abc_21378_n2296) );
  INVX1 INVX1_1135 ( .A(w_mem_inst__abc_21378_n2297), .Y(w_mem_inst__abc_21378_n2299_1) );
  INVX1 INVX1_1136 ( .A(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_21378_n2336) );
  INVX1 INVX1_1137 ( .A(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_21378_n2338_1) );
  INVX1 INVX1_1138 ( .A(w_mem_inst__abc_21378_n2340), .Y(w_mem_inst__abc_21378_n2341) );
  INVX1 INVX1_1139 ( .A(w_mem_inst__abc_21378_n2343_1), .Y(w_mem_inst__abc_21378_n2344) );
  INVX1 INVX1_114 ( .A(_abc_15724_n1338), .Y(_abc_15724_n1339) );
  INVX1 INVX1_1140 ( .A(w_mem_inst__abc_21378_n2345), .Y(w_mem_inst__abc_21378_n2347_1) );
  INVX1 INVX1_1141 ( .A(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_21378_n2384) );
  INVX1 INVX1_1142 ( .A(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_21378_n2386_1) );
  INVX1 INVX1_1143 ( .A(w_mem_inst__abc_21378_n2388), .Y(w_mem_inst__abc_21378_n2389) );
  INVX1 INVX1_1144 ( .A(w_mem_inst__abc_21378_n2391_1), .Y(w_mem_inst__abc_21378_n2392) );
  INVX1 INVX1_1145 ( .A(w_mem_inst__abc_21378_n2393), .Y(w_mem_inst__abc_21378_n2395_1) );
  INVX1 INVX1_1146 ( .A(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_21378_n2432) );
  INVX1 INVX1_1147 ( .A(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_21378_n2434_1) );
  INVX1 INVX1_1148 ( .A(w_mem_inst__abc_21378_n2436), .Y(w_mem_inst__abc_21378_n2437) );
  INVX1 INVX1_1149 ( .A(w_mem_inst__abc_21378_n2439_1), .Y(w_mem_inst__abc_21378_n2440) );
  INVX1 INVX1_115 ( .A(_abc_15724_n1323), .Y(_abc_15724_n1341_1) );
  INVX1 INVX1_1150 ( .A(w_mem_inst__abc_21378_n2441), .Y(w_mem_inst__abc_21378_n2443_1) );
  INVX1 INVX1_1151 ( .A(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_21378_n2480) );
  INVX1 INVX1_1152 ( .A(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_21378_n2482_1) );
  INVX1 INVX1_1153 ( .A(w_mem_inst__abc_21378_n2484), .Y(w_mem_inst__abc_21378_n2485) );
  INVX1 INVX1_1154 ( .A(w_mem_inst__abc_21378_n2487_1), .Y(w_mem_inst__abc_21378_n2488) );
  INVX1 INVX1_1155 ( .A(w_mem_inst__abc_21378_n2489), .Y(w_mem_inst__abc_21378_n2491_1) );
  INVX1 INVX1_1156 ( .A(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_21378_n2528) );
  INVX1 INVX1_1157 ( .A(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_21378_n2530_1) );
  INVX1 INVX1_1158 ( .A(w_mem_inst__abc_21378_n2532), .Y(w_mem_inst__abc_21378_n2533) );
  INVX1 INVX1_1159 ( .A(w_mem_inst__abc_21378_n2535_1), .Y(w_mem_inst__abc_21378_n2536) );
  INVX1 INVX1_116 ( .A(_abc_15724_n1344), .Y(_abc_15724_n1345) );
  INVX1 INVX1_1160 ( .A(w_mem_inst__abc_21378_n2537), .Y(w_mem_inst__abc_21378_n2539_1) );
  INVX1 INVX1_1161 ( .A(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_21378_n2576) );
  INVX1 INVX1_1162 ( .A(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_21378_n2578_1) );
  INVX1 INVX1_1163 ( .A(w_mem_inst__abc_21378_n2580), .Y(w_mem_inst__abc_21378_n2581) );
  INVX1 INVX1_1164 ( .A(w_mem_inst__abc_21378_n2583_1), .Y(w_mem_inst__abc_21378_n2584) );
  INVX1 INVX1_1165 ( .A(w_mem_inst__abc_21378_n2585), .Y(w_mem_inst__abc_21378_n2587_1) );
  INVX1 INVX1_1166 ( .A(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_21378_n2624) );
  INVX1 INVX1_1167 ( .A(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_21378_n2626_1) );
  INVX1 INVX1_1168 ( .A(w_mem_inst__abc_21378_n2628), .Y(w_mem_inst__abc_21378_n2629) );
  INVX1 INVX1_1169 ( .A(w_mem_inst__abc_21378_n2631_1), .Y(w_mem_inst__abc_21378_n2632) );
  INVX1 INVX1_117 ( .A(_abc_15724_n1346), .Y(_abc_15724_n1347) );
  INVX1 INVX1_1170 ( .A(w_mem_inst__abc_21378_n2633), .Y(w_mem_inst__abc_21378_n2635_1) );
  INVX1 INVX1_1171 ( .A(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_21378_n2672) );
  INVX1 INVX1_1172 ( .A(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_21378_n2674_1) );
  INVX1 INVX1_1173 ( .A(w_mem_inst__abc_21378_n2676), .Y(w_mem_inst__abc_21378_n2677) );
  INVX1 INVX1_1174 ( .A(w_mem_inst__abc_21378_n2679_1), .Y(w_mem_inst__abc_21378_n2680) );
  INVX1 INVX1_1175 ( .A(w_mem_inst__abc_21378_n2681), .Y(w_mem_inst__abc_21378_n2683_1) );
  INVX1 INVX1_1176 ( .A(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_21378_n2720) );
  INVX1 INVX1_1177 ( .A(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_21378_n2722_1) );
  INVX1 INVX1_1178 ( .A(w_mem_inst__abc_21378_n2724), .Y(w_mem_inst__abc_21378_n2725) );
  INVX1 INVX1_1179 ( .A(w_mem_inst__abc_21378_n2727_1), .Y(w_mem_inst__abc_21378_n2728) );
  INVX1 INVX1_118 ( .A(_abc_15724_n1354), .Y(_abc_15724_n1355) );
  INVX1 INVX1_1180 ( .A(w_mem_inst__abc_21378_n2729), .Y(w_mem_inst__abc_21378_n2731_1) );
  INVX1 INVX1_1181 ( .A(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_21378_n2768) );
  INVX1 INVX1_1182 ( .A(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_21378_n2770_1) );
  INVX1 INVX1_1183 ( .A(w_mem_inst__abc_21378_n2772), .Y(w_mem_inst__abc_21378_n2773) );
  INVX1 INVX1_1184 ( .A(w_mem_inst__abc_21378_n2775_1), .Y(w_mem_inst__abc_21378_n2776) );
  INVX1 INVX1_1185 ( .A(w_mem_inst__abc_21378_n2777), .Y(w_mem_inst__abc_21378_n2779_1) );
  INVX1 INVX1_1186 ( .A(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_21378_n2816) );
  INVX1 INVX1_1187 ( .A(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_21378_n2818_1) );
  INVX1 INVX1_1188 ( .A(w_mem_inst__abc_21378_n2820), .Y(w_mem_inst__abc_21378_n2821) );
  INVX1 INVX1_1189 ( .A(w_mem_inst__abc_21378_n2823_1), .Y(w_mem_inst__abc_21378_n2824) );
  INVX1 INVX1_119 ( .A(_abc_15724_n1356), .Y(_abc_15724_n1357) );
  INVX1 INVX1_1190 ( .A(w_mem_inst__abc_21378_n2825), .Y(w_mem_inst__abc_21378_n2827_1) );
  INVX1 INVX1_1191 ( .A(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_21378_n2864) );
  INVX1 INVX1_1192 ( .A(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_21378_n2866_1) );
  INVX1 INVX1_1193 ( .A(w_mem_inst__abc_21378_n2868), .Y(w_mem_inst__abc_21378_n2869) );
  INVX1 INVX1_1194 ( .A(w_mem_inst__abc_21378_n2871_1), .Y(w_mem_inst__abc_21378_n2872) );
  INVX1 INVX1_1195 ( .A(w_mem_inst__abc_21378_n2873), .Y(w_mem_inst__abc_21378_n2875_1) );
  INVX1 INVX1_1196 ( .A(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_21378_n2912) );
  INVX1 INVX1_1197 ( .A(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_21378_n2914_1) );
  INVX1 INVX1_1198 ( .A(w_mem_inst__abc_21378_n2916), .Y(w_mem_inst__abc_21378_n2917) );
  INVX1 INVX1_1199 ( .A(w_mem_inst__abc_21378_n2919_1), .Y(w_mem_inst__abc_21378_n2920) );
  INVX1 INVX1_12 ( .A(_abc_15724_n741_1), .Y(_abc_15724_n742) );
  INVX1 INVX1_120 ( .A(_abc_15724_n1352_1), .Y(_abc_15724_n1359) );
  INVX1 INVX1_1200 ( .A(w_mem_inst__abc_21378_n2921), .Y(w_mem_inst__abc_21378_n2923_1) );
  INVX1 INVX1_1201 ( .A(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_21378_n2960) );
  INVX1 INVX1_1202 ( .A(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_21378_n2962_1) );
  INVX1 INVX1_1203 ( .A(w_mem_inst__abc_21378_n2964), .Y(w_mem_inst__abc_21378_n2965) );
  INVX1 INVX1_1204 ( .A(w_mem_inst__abc_21378_n2967_1), .Y(w_mem_inst__abc_21378_n2968) );
  INVX1 INVX1_1205 ( .A(w_mem_inst__abc_21378_n2969), .Y(w_mem_inst__abc_21378_n2971_1) );
  INVX1 INVX1_1206 ( .A(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_21378_n3008) );
  INVX1 INVX1_1207 ( .A(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_21378_n3010_1) );
  INVX1 INVX1_1208 ( .A(w_mem_inst__abc_21378_n3012), .Y(w_mem_inst__abc_21378_n3013) );
  INVX1 INVX1_1209 ( .A(w_mem_inst__abc_21378_n3015_1), .Y(w_mem_inst__abc_21378_n3016) );
  INVX1 INVX1_121 ( .A(_abc_15724_n1370), .Y(_abc_15724_n1371_1) );
  INVX1 INVX1_1210 ( .A(w_mem_inst__abc_21378_n3017), .Y(w_mem_inst__abc_21378_n3019_1) );
  INVX1 INVX1_1211 ( .A(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_21378_n3056) );
  INVX1 INVX1_1212 ( .A(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_21378_n3058_1) );
  INVX1 INVX1_1213 ( .A(w_mem_inst__abc_21378_n3060), .Y(w_mem_inst__abc_21378_n3061) );
  INVX1 INVX1_1214 ( .A(w_mem_inst__abc_21378_n3063_1), .Y(w_mem_inst__abc_21378_n3064) );
  INVX1 INVX1_1215 ( .A(w_mem_inst__abc_21378_n3065), .Y(w_mem_inst__abc_21378_n3067_1) );
  INVX1 INVX1_1216 ( .A(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_21378_n3104) );
  INVX1 INVX1_1217 ( .A(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_21378_n3106_1) );
  INVX1 INVX1_1218 ( .A(w_mem_inst__abc_21378_n3108), .Y(w_mem_inst__abc_21378_n3109) );
  INVX1 INVX1_1219 ( .A(w_mem_inst__abc_21378_n3111_1), .Y(w_mem_inst__abc_21378_n3112) );
  INVX1 INVX1_122 ( .A(_abc_15724_n1381), .Y(_abc_15724_n1382) );
  INVX1 INVX1_1220 ( .A(w_mem_inst__abc_21378_n3113), .Y(w_mem_inst__abc_21378_n3115_1) );
  INVX1 INVX1_1221 ( .A(round_ctr_inc_bF_buf10), .Y(w_mem_inst__abc_21378_n6229) );
  INVX1 INVX1_1222 ( .A(w_mem_inst__abc_21378_n6242), .Y(w_mem_inst__abc_21378_n6243) );
  INVX1 INVX1_1223 ( .A(w_mem_inst__abc_21378_n6247), .Y(w_mem_inst__abc_21378_n6248) );
  INVX1 INVX1_1224 ( .A(w_mem_inst__abc_21378_n6252), .Y(w_mem_inst__abc_21378_n6253) );
  INVX1 INVX1_1225 ( .A(w_mem_inst__abc_21378_n6257), .Y(w_mem_inst__abc_21378_n6258) );
  INVX1 INVX1_1226 ( .A(w_mem_inst__abc_21378_n6262), .Y(w_mem_inst__abc_21378_n6263) );
  INVX1 INVX1_123 ( .A(_abc_15724_n1385), .Y(_abc_15724_n1386) );
  INVX1 INVX1_124 ( .A(_abc_15724_n1392), .Y(_abc_15724_n1393_1) );
  INVX1 INVX1_125 ( .A(_abc_15724_n1376), .Y(_abc_15724_n1397) );
  INVX1 INVX1_126 ( .A(_abc_15724_n1240_1), .Y(_abc_15724_n1398) );
  INVX1 INVX1_127 ( .A(_abc_15724_n1241), .Y(_abc_15724_n1400_1) );
  INVX1 INVX1_128 ( .A(_abc_15724_n1377_1), .Y(_abc_15724_n1403) );
  INVX1 INVX1_129 ( .A(_abc_15724_n1406), .Y(_abc_15724_n1407) );
  INVX1 INVX1_13 ( .A(_abc_15724_n743), .Y(_abc_15724_n744) );
  INVX1 INVX1_130 ( .A(_abc_15724_n1409), .Y(_abc_15724_n1410) );
  INVX1 INVX1_131 ( .A(_abc_15724_n1417), .Y(_abc_15724_n1418) );
  INVX1 INVX1_132 ( .A(_abc_15724_n1421), .Y(_abc_15724_n1422_1) );
  INVX1 INVX1_133 ( .A(_abc_15724_n1425), .Y(_abc_15724_n1426) );
  INVX1 INVX1_134 ( .A(_abc_15724_n1432), .Y(_abc_15724_n1433) );
  INVX1 INVX1_135 ( .A(_abc_15724_n1438_1), .Y(_abc_15724_n1439) );
  INVX1 INVX1_136 ( .A(_abc_15724_n1441), .Y(_abc_15724_n1442) );
  INVX1 INVX1_137 ( .A(_abc_15724_n1448), .Y(_abc_15724_n1449) );
  INVX1 INVX1_138 ( .A(_abc_15724_n1452), .Y(_abc_15724_n1453) );
  INVX1 INVX1_139 ( .A(_abc_15724_n1454), .Y(_abc_15724_n1457) );
  INVX1 INVX1_14 ( .A(_abc_15724_n755), .Y(_abc_15724_n760_1) );
  INVX1 INVX1_140 ( .A(_abc_15724_n1468), .Y(_abc_15724_n1469) );
  INVX1 INVX1_141 ( .A(_abc_15724_n1470), .Y(_abc_15724_n1474_1) );
  INVX1 INVX1_142 ( .A(_abc_15724_n1480), .Y(_abc_15724_n1481) );
  INVX1 INVX1_143 ( .A(_abc_15724_n1483), .Y(_abc_15724_n1484_1) );
  INVX1 INVX1_144 ( .A(_abc_15724_n1467), .Y(_abc_15724_n1485_1) );
  INVX1 INVX1_145 ( .A(_abc_15724_n1497), .Y(_abc_15724_n1498) );
  INVX1 INVX1_146 ( .A(_abc_15724_n1499), .Y(_abc_15724_n1503) );
  INVX1 INVX1_147 ( .A(_abc_15724_n1510_1), .Y(_abc_15724_n1511) );
  INVX1 INVX1_148 ( .A(_abc_15724_n1518_1), .Y(_abc_15724_n1519_1) );
  INVX1 INVX1_149 ( .A(_abc_15724_n1521), .Y(_abc_15724_n1522) );
  INVX1 INVX1_15 ( .A(_abc_15724_n757_1), .Y(_abc_15724_n762) );
  INVX1 INVX1_150 ( .A(_abc_15724_n1531_1), .Y(_abc_15724_n1532) );
  INVX1 INVX1_151 ( .A(_abc_15724_n1533_1), .Y(_abc_15724_n1534) );
  INVX1 INVX1_152 ( .A(_abc_15724_n1529), .Y(_abc_15724_n1536) );
  INVX1 INVX1_153 ( .A(_abc_15724_n1545), .Y(_abc_15724_n1546) );
  INVX1 INVX1_154 ( .A(_abc_15724_n1543_1), .Y(_abc_15724_n1549) );
  INVX1 INVX1_155 ( .A(_abc_15724_n1547), .Y(_abc_15724_n1550_1) );
  INVX1 INVX1_156 ( .A(_abc_15724_n1558), .Y(_abc_15724_n1559) );
  INVX1 INVX1_157 ( .A(_abc_15724_n1560), .Y(_abc_15724_n1561) );
  INVX1 INVX1_158 ( .A(_abc_15724_n1544), .Y(_abc_15724_n1562) );
  INVX1 INVX1_159 ( .A(_abc_15724_n1564_1), .Y(_abc_15724_n1566) );
  INVX1 INVX1_16 ( .A(_abc_15724_n773), .Y(_abc_15724_n778) );
  INVX1 INVX1_160 ( .A(_abc_15724_n1573_1), .Y(_abc_15724_n1574) );
  INVX1 INVX1_161 ( .A(_abc_15724_n1576), .Y(_abc_15724_n1577) );
  INVX1 INVX1_162 ( .A(_abc_15724_n1578_1), .Y(_abc_15724_n1580) );
  INVX1 INVX1_163 ( .A(_abc_15724_n1587_1), .Y(_abc_15724_n1588) );
  INVX1 INVX1_164 ( .A(_abc_15724_n1590_1), .Y(_abc_15724_n1591_1) );
  INVX1 INVX1_165 ( .A(_abc_15724_n1592), .Y(_abc_15724_n1594) );
  INVX1 INVX1_166 ( .A(_abc_15724_n1601), .Y(_abc_15724_n1602_1) );
  INVX1 INVX1_167 ( .A(_abc_15724_n1604), .Y(_abc_15724_n1605) );
  INVX1 INVX1_168 ( .A(_abc_15724_n1606), .Y(_abc_15724_n1608) );
  INVX1 INVX1_169 ( .A(_abc_15724_n1617_1), .Y(_abc_15724_n1618) );
  INVX1 INVX1_17 ( .A(_abc_15724_n775), .Y(_abc_15724_n780_1) );
  INVX1 INVX1_170 ( .A(_abc_15724_n1603_1), .Y(_abc_15724_n1620) );
  INVX1 INVX1_171 ( .A(_abc_15724_n1623_1), .Y(_abc_15724_n1624_1) );
  INVX1 INVX1_172 ( .A(_abc_15724_n1626), .Y(_abc_15724_n1627) );
  INVX1 INVX1_173 ( .A(_abc_15724_n1632), .Y(_abc_15724_n1633_1) );
  INVX1 INVX1_174 ( .A(_abc_15724_n1635), .Y(_abc_15724_n1636_1) );
  INVX1 INVX1_175 ( .A(_abc_15724_n1638), .Y(_abc_15724_n1639_1) );
  INVX1 INVX1_176 ( .A(_abc_15724_n1644), .Y(_abc_15724_n1645_1) );
  INVX1 INVX1_177 ( .A(_abc_15724_n1647), .Y(_abc_15724_n1648_1) );
  INVX1 INVX1_178 ( .A(_abc_15724_n1651), .Y(_abc_15724_n1652) );
  INVX1 INVX1_179 ( .A(_abc_15724_n1660), .Y(_abc_15724_n1661_1) );
  INVX1 INVX1_18 ( .A(_abc_15724_n790_1), .Y(_abc_15724_n791_1) );
  INVX1 INVX1_180 ( .A(_abc_15724_n1658_1), .Y(_abc_15724_n1664) );
  INVX1 INVX1_181 ( .A(_abc_15724_n1662_1), .Y(_abc_15724_n1665) );
  INVX1 INVX1_182 ( .A(_abc_15724_n1674), .Y(_abc_15724_n1675_1) );
  INVX1 INVX1_183 ( .A(_abc_15724_n1682_1), .Y(_abc_15724_n1683) );
  INVX1 INVX1_184 ( .A(_abc_15724_n1684), .Y(_abc_15724_n1685) );
  INVX1 INVX1_185 ( .A(_abc_15724_n1687), .Y(_abc_15724_n1688_1) );
  INVX1 INVX1_186 ( .A(_abc_15724_n1691), .Y(_abc_15724_n1692_1) );
  INVX1 INVX1_187 ( .A(_abc_15724_n1699), .Y(_abc_15724_n1700_1) );
  INVX1 INVX1_188 ( .A(_abc_15724_n1702), .Y(_abc_15724_n1703) );
  INVX1 INVX1_189 ( .A(_abc_15724_n1705), .Y(_abc_15724_n1706) );
  INVX1 INVX1_19 ( .A(_abc_15724_n795), .Y(_abc_15724_n796) );
  INVX1 INVX1_190 ( .A(_abc_15724_n1711), .Y(_abc_15724_n1712) );
  INVX1 INVX1_191 ( .A(_abc_15724_n1714_1), .Y(_abc_15724_n1715) );
  INVX1 INVX1_192 ( .A(_abc_15724_n1718), .Y(_abc_15724_n1719_1) );
  INVX1 INVX1_193 ( .A(_abc_15724_n1725), .Y(_abc_15724_n1726) );
  INVX1 INVX1_194 ( .A(_abc_15724_n1728_1), .Y(_abc_15724_n1729) );
  INVX1 INVX1_195 ( .A(_abc_15724_n1730), .Y(_abc_15724_n1732_1) );
  INVX1 INVX1_196 ( .A(_abc_15724_n1746), .Y(_abc_15724_n1747) );
  INVX1 INVX1_197 ( .A(_abc_15724_n1749), .Y(_abc_15724_n1750_1) );
  INVX1 INVX1_198 ( .A(_abc_15724_n1752), .Y(_abc_15724_n1753) );
  INVX1 INVX1_199 ( .A(_abc_15724_n1755), .Y(_abc_15724_n1756) );
  INVX1 INVX1_2 ( .A(_abc_15724_n705), .Y(_abc_15724_n706) );
  INVX1 INVX1_20 ( .A(_abc_15724_n797), .Y(_abc_15724_n798) );
  INVX1 INVX1_200 ( .A(_abc_15724_n1759), .Y(_abc_15724_n1760) );
  INVX1 INVX1_201 ( .A(_abc_15724_n1764), .Y(_abc_15724_n1765) );
  INVX1 INVX1_202 ( .A(_abc_15724_n1767_1), .Y(_abc_15724_n1768) );
  INVX1 INVX1_203 ( .A(_abc_15724_n1769), .Y(_abc_15724_n1771) );
  INVX1 INVX1_204 ( .A(_abc_15724_n1780), .Y(_abc_15724_n1781_1) );
  INVX1 INVX1_205 ( .A(_abc_15724_n1786_1), .Y(_abc_15724_n1787) );
  INVX1 INVX1_206 ( .A(_abc_15724_n1790_1), .Y(_abc_15724_n1791) );
  INVX1 INVX1_207 ( .A(_abc_15724_n1795_1), .Y(_abc_15724_n1796) );
  INVX1 INVX1_208 ( .A(_abc_15724_n1798), .Y(_abc_15724_n1799_1) );
  INVX1 INVX1_209 ( .A(_abc_15724_n1800), .Y(_abc_15724_n1802) );
  INVX1 INVX1_21 ( .A(_abc_15724_n789_1), .Y(_abc_15724_n799) );
  INVX1 INVX1_210 ( .A(_abc_15724_n1810), .Y(_abc_15724_n1811) );
  INVX1 INVX1_211 ( .A(_abc_15724_n1816), .Y(_abc_15724_n1817) );
  INVX1 INVX1_212 ( .A(_abc_15724_n1818_1), .Y(_abc_15724_n1819) );
  INVX1 INVX1_213 ( .A(_abc_15724_n1821), .Y(_abc_15724_n1822) );
  INVX1 INVX1_214 ( .A(_abc_15724_n1825), .Y(_abc_15724_n1826) );
  INVX1 INVX1_215 ( .A(_abc_15724_n1832), .Y(_abc_15724_n1833) );
  INVX1 INVX1_216 ( .A(_abc_15724_n1835), .Y(_abc_15724_n1836_1) );
  INVX1 INVX1_217 ( .A(_abc_15724_n1837), .Y(_abc_15724_n1839) );
  INVX1 INVX1_218 ( .A(_abc_15724_n1848), .Y(_abc_15724_n1849) );
  INVX1 INVX1_219 ( .A(_abc_15724_n1854), .Y(_abc_15724_n1855) );
  INVX1 INVX1_22 ( .A(_abc_15724_n786), .Y(_abc_15724_n806_1) );
  INVX1 INVX1_220 ( .A(_abc_15724_n1857), .Y(_abc_15724_n1858) );
  INVX1 INVX1_221 ( .A(_abc_15724_n1863), .Y(_abc_15724_n1864) );
  INVX1 INVX1_222 ( .A(_abc_15724_n1866), .Y(_abc_15724_n1867) );
  INVX1 INVX1_223 ( .A(_abc_15724_n1868), .Y(_abc_15724_n1870_1) );
  INVX1 INVX1_224 ( .A(_abc_15724_n1882), .Y(_abc_15724_n1883) );
  INVX1 INVX1_225 ( .A(_abc_15724_n1884), .Y(_abc_15724_n1885_1) );
  INVX1 INVX1_226 ( .A(_abc_15724_n1887), .Y(_abc_15724_n1888) );
  INVX1 INVX1_227 ( .A(_abc_15724_n1890), .Y(_abc_15724_n1891) );
  INVX1 INVX1_228 ( .A(_abc_15724_n1894), .Y(_abc_15724_n1895) );
  INVX1 INVX1_229 ( .A(_abc_15724_n1901_1), .Y(_abc_15724_n1902) );
  INVX1 INVX1_23 ( .A(_abc_15724_n766_1), .Y(_abc_15724_n815_1) );
  INVX1 INVX1_230 ( .A(_abc_15724_n1907), .Y(_abc_15724_n1908) );
  INVX1 INVX1_231 ( .A(_abc_15724_n1909_1), .Y(_abc_15724_n1910) );
  INVX1 INVX1_232 ( .A(_abc_15724_n1917), .Y(_abc_15724_n1918_1) );
  INVX1 INVX1_233 ( .A(_abc_15724_n1920), .Y(_abc_15724_n1921) );
  INVX1 INVX1_234 ( .A(_abc_15724_n1924), .Y(_abc_15724_n1925) );
  INVX1 INVX1_235 ( .A(_abc_15724_n1931_1), .Y(_abc_15724_n1932) );
  INVX1 INVX1_236 ( .A(_abc_15724_n1929), .Y(_abc_15724_n1935_1) );
  INVX1 INVX1_237 ( .A(_abc_15724_n1933), .Y(_abc_15724_n1936) );
  INVX1 INVX1_238 ( .A(_abc_15724_n1944_1), .Y(_abc_15724_n1945) );
  INVX1 INVX1_239 ( .A(_abc_15724_n1946), .Y(_abc_15724_n1947) );
  INVX1 INVX1_24 ( .A(_abc_15724_n768), .Y(_abc_15724_n817) );
  INVX1 INVX1_240 ( .A(_abc_15724_n1950), .Y(_abc_15724_n1951) );
  INVX1 INVX1_241 ( .A(_abc_15724_n1953_1), .Y(_abc_15724_n1954) );
  INVX1 INVX1_242 ( .A(_abc_15724_n1956), .Y(_abc_15724_n1957_1) );
  INVX1 INVX1_243 ( .A(_abc_15724_n1960), .Y(_abc_15724_n1961) );
  INVX1 INVX1_244 ( .A(_abc_15724_n1970_1), .Y(_abc_15724_n1971) );
  INVX1 INVX1_245 ( .A(_abc_15724_n1972), .Y(_abc_15724_n1973) );
  INVX1 INVX1_246 ( .A(_abc_15724_n1968), .Y(_abc_15724_n1975) );
  INVX1 INVX1_247 ( .A(_abc_15724_n1981), .Y(_abc_15724_n1982) );
  INVX1 INVX1_248 ( .A(_abc_15724_n1984), .Y(_abc_15724_n1985) );
  INVX1 INVX1_249 ( .A(_abc_15724_n1987), .Y(_abc_15724_n1988_1) );
  INVX1 INVX1_25 ( .A(_abc_15724_n825_1), .Y(_abc_15724_n826_1) );
  INVX1 INVX1_250 ( .A(_abc_15724_n1989), .Y(_abc_15724_n1990) );
  INVX1 INVX1_251 ( .A(_abc_15724_n1992), .Y(_abc_15724_n1994) );
  INVX1 INVX1_252 ( .A(_abc_15724_n1999), .Y(_abc_15724_n2000) );
  INVX1 INVX1_253 ( .A(_auto_iopadmap_cc_313_execute_26059_95_), .Y(_abc_15724_n2001) );
  INVX1 INVX1_254 ( .A(c_reg_31_), .Y(_abc_15724_n2003) );
  INVX1 INVX1_255 ( .A(_abc_15724_n2005), .Y(_abc_15724_n2006_1) );
  INVX1 INVX1_256 ( .A(_abc_15724_n2015), .Y(_abc_15724_n2016_1) );
  INVX1 INVX1_257 ( .A(_abc_15724_n2023), .Y(_abc_15724_n2024_1) );
  INVX1 INVX1_258 ( .A(_abc_15724_n2027), .Y(_abc_15724_n2028) );
  INVX1 INVX1_259 ( .A(_abc_15724_n2033), .Y(_abc_15724_n2034_1) );
  INVX1 INVX1_26 ( .A(_abc_15724_n830), .Y(_abc_15724_n831) );
  INVX1 INVX1_260 ( .A(_abc_15724_n2036), .Y(_abc_15724_n2037) );
  INVX1 INVX1_261 ( .A(_abc_15724_n2039), .Y(_abc_15724_n2040) );
  INVX1 INVX1_262 ( .A(_abc_15724_n2048_1), .Y(_abc_15724_n2049) );
  INVX1 INVX1_263 ( .A(_abc_15724_n2046), .Y(_abc_15724_n2052) );
  INVX1 INVX1_264 ( .A(_abc_15724_n2050), .Y(_abc_15724_n2053_1) );
  INVX1 INVX1_265 ( .A(_abc_15724_n2061_1), .Y(_abc_15724_n2062) );
  INVX1 INVX1_266 ( .A(_abc_15724_n2066), .Y(_abc_15724_n2067) );
  INVX1 INVX1_267 ( .A(_abc_15724_n2076), .Y(_abc_15724_n2077) );
  INVX1 INVX1_268 ( .A(_abc_15724_n2079_1), .Y(_abc_15724_n2080) );
  INVX1 INVX1_269 ( .A(_abc_15724_n2088_1), .Y(_abc_15724_n2089) );
  INVX1 INVX1_27 ( .A(_abc_15724_n833_1), .Y(_abc_15724_n834_1) );
  INVX1 INVX1_270 ( .A(_abc_15724_n2092_1), .Y(_abc_15724_n2093) );
  INVX1 INVX1_271 ( .A(_abc_15724_n2099), .Y(_abc_15724_n2100) );
  INVX1 INVX1_272 ( .A(_abc_15724_n2102), .Y(_abc_15724_n2103) );
  INVX1 INVX1_273 ( .A(_abc_15724_n2104), .Y(_abc_15724_n2106) );
  INVX1 INVX1_274 ( .A(_abc_15724_n2112), .Y(_abc_15724_n2113) );
  INVX1 INVX1_275 ( .A(_abc_15724_n2118), .Y(_abc_15724_n2119_1) );
  INVX1 INVX1_276 ( .A(_abc_15724_n2125), .Y(_abc_15724_n2126) );
  INVX1 INVX1_277 ( .A(_abc_15724_n2128), .Y(_abc_15724_n2129) );
  INVX1 INVX1_278 ( .A(_abc_15724_n2130), .Y(_abc_15724_n2132) );
  INVX1 INVX1_279 ( .A(_abc_15724_n2141), .Y(_abc_15724_n2142) );
  INVX1 INVX1_28 ( .A(_abc_15724_n699), .Y(_abc_15724_n835) );
  INVX1 INVX1_280 ( .A(_abc_15724_n2147), .Y(_abc_15724_n2148_1) );
  INVX1 INVX1_281 ( .A(_abc_15724_n2151), .Y(_abc_15724_n2152_1) );
  INVX1 INVX1_282 ( .A(_abc_15724_n2156_1), .Y(_abc_15724_n2157) );
  INVX1 INVX1_283 ( .A(_abc_15724_n2159), .Y(_abc_15724_n2160_1) );
  INVX1 INVX1_284 ( .A(_abc_15724_n2161), .Y(_abc_15724_n2163_1) );
  INVX1 INVX1_285 ( .A(_abc_15724_n2180_1), .Y(_abc_15724_n2181) );
  INVX1 INVX1_286 ( .A(_abc_15724_n2184), .Y(_abc_15724_n2185) );
  INVX1 INVX1_287 ( .A(_abc_15724_n2189), .Y(_abc_15724_n2190) );
  INVX1 INVX1_288 ( .A(_abc_15724_n2192), .Y(_abc_15724_n2193) );
  INVX1 INVX1_289 ( .A(_abc_15724_n2194), .Y(_abc_15724_n2196) );
  INVX1 INVX1_29 ( .A(_abc_15724_n842), .Y(_abc_15724_n843) );
  INVX1 INVX1_290 ( .A(_abc_15724_n2205), .Y(_abc_15724_n2206) );
  INVX1 INVX1_291 ( .A(_abc_15724_n2211), .Y(_abc_15724_n2212) );
  INVX1 INVX1_292 ( .A(_abc_15724_n2214), .Y(_abc_15724_n2215) );
  INVX1 INVX1_293 ( .A(_abc_15724_n2220), .Y(_abc_15724_n2221) );
  INVX1 INVX1_294 ( .A(_abc_15724_n2223), .Y(_abc_15724_n2224) );
  INVX1 INVX1_295 ( .A(_abc_15724_n2225), .Y(_abc_15724_n2227) );
  INVX1 INVX1_296 ( .A(_abc_15724_n2243), .Y(_abc_15724_n2244) );
  INVX1 INVX1_297 ( .A(_abc_15724_n2247), .Y(_abc_15724_n2248) );
  INVX1 INVX1_298 ( .A(_abc_15724_n2255), .Y(_abc_15724_n2256) );
  INVX1 INVX1_299 ( .A(_abc_15724_n2258), .Y(_abc_15724_n2259) );
  INVX1 INVX1_3 ( .A(_abc_15724_n709_1), .Y(_abc_15724_n710_1) );
  INVX1 INVX1_30 ( .A(_abc_15724_n846), .Y(_abc_15724_n847_1) );
  INVX1 INVX1_300 ( .A(_abc_15724_n2261), .Y(_abc_15724_n2262) );
  INVX1 INVX1_301 ( .A(_abc_15724_n2267), .Y(_abc_15724_n2268) );
  INVX1 INVX1_302 ( .A(_abc_15724_n2270), .Y(_abc_15724_n2271) );
  INVX1 INVX1_303 ( .A(_abc_15724_n2274), .Y(_abc_15724_n2275) );
  INVX1 INVX1_304 ( .A(_abc_15724_n2283), .Y(_abc_15724_n2284) );
  INVX1 INVX1_305 ( .A(_abc_15724_n2281), .Y(_abc_15724_n2287_1) );
  INVX1 INVX1_306 ( .A(_abc_15724_n2285), .Y(_abc_15724_n2288) );
  INVX1 INVX1_307 ( .A(_abc_15724_n2308), .Y(_abc_15724_n2309) );
  INVX1 INVX1_308 ( .A(_abc_15724_n2312), .Y(_abc_15724_n2313) );
  INVX1 INVX1_309 ( .A(_abc_15724_n2319), .Y(_abc_15724_n2320) );
  INVX1 INVX1_31 ( .A(_abc_15724_n857), .Y(_abc_15724_n858) );
  INVX1 INVX1_310 ( .A(_abc_15724_n2324), .Y(_abc_15724_n2325) );
  INVX1 INVX1_311 ( .A(_abc_15724_n2331), .Y(_abc_15724_n2332) );
  INVX1 INVX1_312 ( .A(_abc_15724_n2335), .Y(_abc_15724_n2336) );
  INVX1 INVX1_313 ( .A(_abc_15724_n2342), .Y(_abc_15724_n2343) );
  INVX1 INVX1_314 ( .A(_abc_15724_n2345), .Y(_abc_15724_n2346) );
  INVX1 INVX1_315 ( .A(_abc_15724_n2347), .Y(_abc_15724_n2349) );
  INVX1 INVX1_316 ( .A(_abc_15724_n2371), .Y(_abc_15724_n2372) );
  INVX1 INVX1_317 ( .A(_abc_15724_n2375), .Y(_abc_15724_n2376) );
  INVX1 INVX1_318 ( .A(_abc_15724_n2382), .Y(_abc_15724_n2383) );
  INVX1 INVX1_319 ( .A(_abc_15724_n2385), .Y(_abc_15724_n2386) );
  INVX1 INVX1_32 ( .A(_abc_15724_n855_1), .Y(_abc_15724_n861) );
  INVX1 INVX1_320 ( .A(_abc_15724_n2387), .Y(_abc_15724_n2389) );
  INVX1 INVX1_321 ( .A(_abc_15724_n2402), .Y(_abc_15724_n2403) );
  INVX1 INVX1_322 ( .A(_abc_15724_n2406_1), .Y(_abc_15724_n2407) );
  INVX1 INVX1_323 ( .A(_abc_15724_n2413), .Y(_abc_15724_n2414) );
  INVX1 INVX1_324 ( .A(_abc_15724_n2416), .Y(_abc_15724_n2417) );
  INVX1 INVX1_325 ( .A(_abc_15724_n2418), .Y(_abc_15724_n2420) );
  INVX1 INVX1_326 ( .A(_abc_15724_n2437), .Y(_abc_15724_n2438) );
  INVX1 INVX1_327 ( .A(_abc_15724_n2441), .Y(_abc_15724_n2442) );
  INVX1 INVX1_328 ( .A(_abc_15724_n2448), .Y(_abc_15724_n2449_1) );
  INVX1 INVX1_329 ( .A(_abc_15724_n2446), .Y(_abc_15724_n2452) );
  INVX1 INVX1_33 ( .A(_abc_15724_n859), .Y(_abc_15724_n862) );
  INVX1 INVX1_330 ( .A(_abc_15724_n2450), .Y(_abc_15724_n2453) );
  INVX1 INVX1_331 ( .A(_abc_15724_n2461), .Y(_abc_15724_n2462) );
  INVX1 INVX1_332 ( .A(_abc_15724_n2470), .Y(_abc_15724_n2471) );
  INVX1 INVX1_333 ( .A(_auto_iopadmap_cc_313_execute_26059_127_), .Y(_abc_15724_n2478) );
  INVX1 INVX1_334 ( .A(b_reg_31_), .Y(_abc_15724_n2480) );
  INVX1 INVX1_335 ( .A(_abc_15724_n2482), .Y(_abc_15724_n2483) );
  INVX1 INVX1_336 ( .A(_abc_15724_n2477), .Y(_abc_15724_n2485) );
  INVX1 INVX1_337 ( .A(_abc_15724_n2493), .Y(_abc_15724_n2494) );
  INVX1 INVX1_338 ( .A(_abc_15724_n2501), .Y(_abc_15724_n2502) );
  INVX1 INVX1_339 ( .A(_abc_15724_n2505), .Y(_abc_15724_n2506) );
  INVX1 INVX1_34 ( .A(_abc_15724_n881), .Y(_abc_15724_n882) );
  INVX1 INVX1_340 ( .A(_abc_15724_n2513), .Y(_abc_15724_n2514) );
  INVX1 INVX1_341 ( .A(_abc_15724_n2515), .Y(_abc_15724_n2516) );
  INVX1 INVX1_342 ( .A(_abc_15724_n2511), .Y(_abc_15724_n2518) );
  INVX1 INVX1_343 ( .A(_abc_15724_n2524_1), .Y(_abc_15724_n2525) );
  INVX1 INVX1_344 ( .A(_abc_15724_n2527_1), .Y(_abc_15724_n2528) );
  INVX1 INVX1_345 ( .A(_abc_15724_n2529), .Y(_abc_15724_n2531) );
  INVX1 INVX1_346 ( .A(_abc_15724_n2538), .Y(_abc_15724_n2539) );
  INVX1 INVX1_347 ( .A(_abc_15724_n2540), .Y(_abc_15724_n2541) );
  INVX1 INVX1_348 ( .A(_abc_15724_n2526), .Y(_abc_15724_n2542) );
  INVX1 INVX1_349 ( .A(_abc_15724_n2544), .Y(_abc_15724_n2546) );
  INVX1 INVX1_35 ( .A(_abc_15724_n885_1), .Y(_abc_15724_n886) );
  INVX1 INVX1_350 ( .A(_abc_15724_n2555), .Y(_abc_15724_n2556) );
  INVX1 INVX1_351 ( .A(_abc_15724_n2557), .Y(_abc_15724_n2558) );
  INVX1 INVX1_352 ( .A(_abc_15724_n2553), .Y(_abc_15724_n2560) );
  INVX1 INVX1_353 ( .A(_abc_15724_n2566), .Y(_abc_15724_n2567) );
  INVX1 INVX1_354 ( .A(_abc_15724_n2569), .Y(_abc_15724_n2570_1) );
  INVX1 INVX1_355 ( .A(_abc_15724_n2571), .Y(_abc_15724_n2573_1) );
  INVX1 INVX1_356 ( .A(_abc_15724_n2574), .Y(_abc_15724_n2579) );
  INVX1 INVX1_357 ( .A(_abc_15724_n2581), .Y(_abc_15724_n2582) );
  INVX1 INVX1_358 ( .A(_abc_15724_n2583), .Y(_abc_15724_n2586) );
  INVX1 INVX1_359 ( .A(_abc_15724_n2588), .Y(_abc_15724_n2589) );
  INVX1 INVX1_36 ( .A(_abc_15724_n892), .Y(_abc_15724_n893) );
  INVX1 INVX1_360 ( .A(_abc_15724_n2595), .Y(_abc_15724_n2596) );
  INVX1 INVX1_361 ( .A(_abc_15724_n2598), .Y(_abc_15724_n2599) );
  INVX1 INVX1_362 ( .A(_abc_15724_n2602), .Y(_abc_15724_n2603) );
  INVX1 INVX1_363 ( .A(_abc_15724_n2609), .Y(_abc_15724_n2610) );
  INVX1 INVX1_364 ( .A(_abc_15724_n2612_1), .Y(_abc_15724_n2613) );
  INVX1 INVX1_365 ( .A(_abc_15724_n2614), .Y(_abc_15724_n2616) );
  INVX1 INVX1_366 ( .A(_abc_15724_n2625), .Y(_abc_15724_n2626) );
  INVX1 INVX1_367 ( .A(_abc_15724_n2629), .Y(_abc_15724_n2630) );
  INVX1 INVX1_368 ( .A(_abc_15724_n2635), .Y(_abc_15724_n2636) );
  INVX1 INVX1_369 ( .A(_abc_15724_n2642), .Y(_abc_15724_n2643) );
  INVX1 INVX1_37 ( .A(_abc_15724_n895), .Y(_abc_15724_n896) );
  INVX1 INVX1_370 ( .A(_abc_15724_n2640), .Y(_abc_15724_n2646) );
  INVX1 INVX1_371 ( .A(_abc_15724_n2644), .Y(_abc_15724_n2647) );
  INVX1 INVX1_372 ( .A(_abc_15724_n2655), .Y(_abc_15724_n2656) );
  INVX1 INVX1_373 ( .A(_abc_15724_n2661), .Y(_abc_15724_n2662) );
  INVX1 INVX1_374 ( .A(_abc_15724_n2663), .Y(_abc_15724_n2664) );
  INVX1 INVX1_375 ( .A(_abc_15724_n2666), .Y(_abc_15724_n2667) );
  INVX1 INVX1_376 ( .A(_abc_15724_n2670), .Y(_abc_15724_n2671) );
  INVX1 INVX1_377 ( .A(_abc_15724_n2675), .Y(_abc_15724_n2676) );
  INVX1 INVX1_378 ( .A(_abc_15724_n2678), .Y(_abc_15724_n2679) );
  INVX1 INVX1_379 ( .A(_abc_15724_n2680), .Y(_abc_15724_n2682) );
  INVX1 INVX1_38 ( .A(_abc_15724_n897_1), .Y(_abc_15724_n899_1) );
  INVX1 INVX1_380 ( .A(_abc_15724_n2691_1), .Y(_abc_15724_n2692) );
  INVX1 INVX1_381 ( .A(_abc_15724_n2677), .Y(_abc_15724_n2694) );
  INVX1 INVX1_382 ( .A(_abc_15724_n2697), .Y(_abc_15724_n2698) );
  INVX1 INVX1_383 ( .A(_abc_15724_n2699), .Y(_abc_15724_n2700) );
  INVX1 INVX1_384 ( .A(_abc_15724_n2707), .Y(_abc_15724_n2708) );
  INVX1 INVX1_385 ( .A(_abc_15724_n2709), .Y(_abc_15724_n2710) );
  INVX1 INVX1_386 ( .A(_abc_15724_n2705), .Y(_abc_15724_n2712) );
  INVX1 INVX1_387 ( .A(_abc_15724_n2719), .Y(_abc_15724_n2720) );
  INVX1 INVX1_388 ( .A(_abc_15724_n2722), .Y(_abc_15724_n2723) );
  INVX1 INVX1_389 ( .A(_abc_15724_n2727), .Y(_abc_15724_n2728) );
  INVX1 INVX1_39 ( .A(_abc_15724_n915), .Y(_abc_15724_n916) );
  INVX1 INVX1_390 ( .A(_abc_15724_n2730), .Y(_abc_15724_n2731_1) );
  INVX1 INVX1_391 ( .A(_abc_15724_n2733), .Y(_abc_15724_n2734_1) );
  INVX1 INVX1_392 ( .A(_abc_15724_n2737), .Y(_abc_15724_n2738) );
  INVX1 INVX1_393 ( .A(_abc_15724_n2745), .Y(_abc_15724_n2746) );
  INVX1 INVX1_394 ( .A(_abc_15724_n2748), .Y(_abc_15724_n2749) );
  INVX1 INVX1_395 ( .A(_abc_15724_n2751), .Y(_abc_15724_n2752) );
  INVX1 INVX1_396 ( .A(_abc_15724_n2757), .Y(_abc_15724_n2758) );
  INVX1 INVX1_397 ( .A(_abc_15724_n2760), .Y(_abc_15724_n2761) );
  INVX1 INVX1_398 ( .A(_abc_15724_n2764), .Y(_abc_15724_n2765) );
  INVX1 INVX1_399 ( .A(_abc_15724_n2773), .Y(_abc_15724_n2774) );
  INVX1 INVX1_4 ( .A(_abc_15724_n714), .Y(_abc_15724_n715) );
  INVX1 INVX1_40 ( .A(_abc_15724_n919), .Y(_abc_15724_n920) );
  INVX1 INVX1_400 ( .A(_abc_15724_n2771), .Y(_abc_15724_n2777) );
  INVX1 INVX1_401 ( .A(_abc_15724_n2775), .Y(_abc_15724_n2778) );
  INVX1 INVX1_402 ( .A(_abc_15724_n2787), .Y(_abc_15724_n2788) );
  INVX1 INVX1_403 ( .A(_abc_15724_n2795), .Y(_abc_15724_n2796) );
  INVX1 INVX1_404 ( .A(_abc_15724_n2797), .Y(_abc_15724_n2798) );
  INVX1 INVX1_405 ( .A(_abc_15724_n2800), .Y(_abc_15724_n2801) );
  INVX1 INVX1_406 ( .A(_abc_15724_n2804), .Y(_abc_15724_n2805) );
  INVX1 INVX1_407 ( .A(_abc_15724_n2810), .Y(_abc_15724_n2811) );
  INVX1 INVX1_408 ( .A(_abc_15724_n2813), .Y(_abc_15724_n2814) );
  INVX1 INVX1_409 ( .A(_abc_15724_n2816), .Y(_abc_15724_n2817) );
  INVX1 INVX1_41 ( .A(_abc_15724_n926), .Y(_abc_15724_n927) );
  INVX1 INVX1_410 ( .A(_abc_15724_n2824), .Y(_abc_15724_n2825) );
  INVX1 INVX1_411 ( .A(_abc_15724_n2828), .Y(_abc_15724_n2829) );
  INVX1 INVX1_412 ( .A(_abc_15724_n2835), .Y(_abc_15724_n2836) );
  INVX1 INVX1_413 ( .A(_abc_15724_n2838), .Y(_abc_15724_n2839) );
  INVX1 INVX1_414 ( .A(_abc_15724_n2840), .Y(_abc_15724_n2842) );
  INVX1 INVX1_415 ( .A(_abc_15724_n2854), .Y(_abc_15724_n2855) );
  INVX1 INVX1_416 ( .A(_abc_15724_n2857), .Y(_abc_15724_n2858) );
  INVX1 INVX1_417 ( .A(_abc_15724_n2860), .Y(_abc_15724_n2861) );
  INVX1 INVX1_418 ( .A(_abc_15724_n2863), .Y(_abc_15724_n2864) );
  INVX1 INVX1_419 ( .A(_abc_15724_n2867), .Y(_abc_15724_n2868) );
  INVX1 INVX1_42 ( .A(_abc_15724_n932_1), .Y(_abc_15724_n933) );
  INVX1 INVX1_420 ( .A(_abc_15724_n2874), .Y(_abc_15724_n2875) );
  INVX1 INVX1_421 ( .A(_abc_15724_n2877), .Y(_abc_15724_n2878) );
  INVX1 INVX1_422 ( .A(_abc_15724_n2879), .Y(_abc_15724_n2881) );
  INVX1 INVX1_423 ( .A(_abc_15724_n2894_1), .Y(_abc_15724_n2895) );
  INVX1 INVX1_424 ( .A(_abc_15724_n2898), .Y(_abc_15724_n2899) );
  INVX1 INVX1_425 ( .A(_abc_15724_n2907), .Y(_abc_15724_n2908) );
  INVX1 INVX1_426 ( .A(_abc_15724_n2909), .Y(_abc_15724_n2912) );
  INVX1 INVX1_427 ( .A(_abc_15724_n2919), .Y(_abc_15724_n2920) );
  INVX1 INVX1_428 ( .A(_abc_15724_n2923), .Y(_abc_15724_n2924) );
  INVX1 INVX1_429 ( .A(_abc_15724_n2926), .Y(_abc_15724_n2927_1) );
  INVX1 INVX1_43 ( .A(_abc_15724_n934_1), .Y(_abc_15724_n935) );
  INVX1 INVX1_430 ( .A(_abc_15724_n2929), .Y(_abc_15724_n2930_1) );
  INVX1 INVX1_431 ( .A(_abc_15724_n2932), .Y(_abc_15724_n2933) );
  INVX1 INVX1_432 ( .A(_abc_15724_n2936), .Y(_abc_15724_n2937) );
  INVX1 INVX1_433 ( .A(_abc_15724_n2943), .Y(_abc_15724_n2944) );
  INVX1 INVX1_434 ( .A(_abc_15724_n2945), .Y(_abc_15724_n2946) );
  INVX1 INVX1_435 ( .A(_abc_15724_n2941), .Y(_abc_15724_n2948) );
  INVX1 INVX1_436 ( .A(_abc_15724_n2956), .Y(_abc_15724_n2957) );
  INVX1 INVX1_437 ( .A(_abc_15724_n2960), .Y(_abc_15724_n2961) );
  INVX1 INVX1_438 ( .A(_abc_15724_n2962), .Y(_abc_15724_n2963) );
  INVX1 INVX1_439 ( .A(_abc_15724_n2965), .Y(_abc_15724_n2966) );
  INVX1 INVX1_44 ( .A(_abc_15724_n941), .Y(_abc_15724_n942) );
  INVX1 INVX1_440 ( .A(_abc_15724_n2958), .Y(_abc_15724_n2968_1) );
  INVX1 INVX1_441 ( .A(_abc_15724_n2977), .Y(_abc_15724_n2978) );
  INVX1 INVX1_442 ( .A(_abc_15724_n2975), .Y(_abc_15724_n2981) );
  INVX1 INVX1_443 ( .A(_abc_15724_n2979), .Y(_abc_15724_n2982) );
  INVX1 INVX1_444 ( .A(round_ctr_inc_bF_buf12), .Y(_abc_15724_n2990) );
  INVX1 INVX1_445 ( .A(round_ctr_rst_bF_buf63), .Y(_abc_15724_n2991) );
  INVX1 INVX1_446 ( .A(_abc_15724_n3700), .Y(_abc_15724_n3701) );
  INVX1 INVX1_447 ( .A(round_ctr_reg_6_), .Y(_abc_15724_n3702) );
  INVX1 INVX1_448 ( .A(_abc_15724_n3703), .Y(_abc_15724_n3704) );
  INVX1 INVX1_449 ( .A(d_reg_0_), .Y(_abc_15724_n3707) );
  INVX1 INVX1_45 ( .A(_abc_15724_n945_1), .Y(_abc_15724_n946) );
  INVX1 INVX1_450 ( .A(c_reg_0_), .Y(_abc_15724_n3709) );
  INVX1 INVX1_451 ( .A(b_reg_0_), .Y(_abc_15724_n3710) );
  INVX1 INVX1_452 ( .A(_abc_15724_n3712), .Y(_abc_15724_n3713) );
  INVX1 INVX1_453 ( .A(_abc_15724_n3727), .Y(_abc_15724_n3728) );
  INVX1 INVX1_454 ( .A(_abc_15724_n3723), .Y(_abc_15724_n3735) );
  INVX1 INVX1_455 ( .A(_abc_15724_n3711), .Y(_abc_15724_n3738) );
  INVX1 INVX1_456 ( .A(_abc_15724_n3741), .Y(_abc_15724_n3742) );
  INVX1 INVX1_457 ( .A(_abc_15724_n3744), .Y(_abc_15724_n3745) );
  INVX1 INVX1_458 ( .A(_abc_15724_n3747), .Y(_abc_15724_n3748) );
  INVX1 INVX1_459 ( .A(w_0_), .Y(_abc_15724_n3751) );
  INVX1 INVX1_46 ( .A(_abc_15724_n949), .Y(_abc_15724_n950) );
  INVX1 INVX1_460 ( .A(_abc_15724_n3749), .Y(_abc_15724_n3752) );
  INVX1 INVX1_461 ( .A(_abc_15724_n3754), .Y(_abc_15724_n3755) );
  INVX1 INVX1_462 ( .A(_abc_15724_n3758), .Y(_abc_15724_n3759) );
  INVX1 INVX1_463 ( .A(_abc_15724_n3761), .Y(_abc_15724_n3762) );
  INVX1 INVX1_464 ( .A(c_reg_1_), .Y(_abc_15724_n3770) );
  INVX1 INVX1_465 ( .A(b_reg_1_), .Y(_abc_15724_n3771) );
  INVX1 INVX1_466 ( .A(_abc_15724_n3776), .Y(_abc_15724_n3777) );
  INVX1 INVX1_467 ( .A(_abc_15724_n3773), .Y(_abc_15724_n3780) );
  INVX1 INVX1_468 ( .A(_abc_15724_n3784), .Y(_abc_15724_n3785) );
  INVX1 INVX1_469 ( .A(_abc_15724_n3786), .Y(_abc_15724_n3787) );
  INVX1 INVX1_47 ( .A(_abc_15724_n956_1), .Y(_abc_15724_n957) );
  INVX1 INVX1_470 ( .A(_abc_15724_n3793), .Y(_abc_15724_n3794) );
  INVX1 INVX1_471 ( .A(_abc_15724_n3796), .Y(_abc_15724_n3797) );
  INVX1 INVX1_472 ( .A(_abc_15724_n3800), .Y(_abc_15724_n3801) );
  INVX1 INVX1_473 ( .A(_abc_15724_n3774), .Y(_abc_15724_n3807) );
  INVX1 INVX1_474 ( .A(_abc_15724_n3791), .Y(_abc_15724_n3814) );
  INVX1 INVX1_475 ( .A(_abc_15724_n3798), .Y(_abc_15724_n3815) );
  INVX1 INVX1_476 ( .A(_abc_15724_n3832), .Y(_abc_15724_n3834) );
  INVX1 INVX1_477 ( .A(_abc_15724_n3833), .Y(_abc_15724_n3843) );
  INVX1 INVX1_478 ( .A(c_reg_2_), .Y(_abc_15724_n3847) );
  INVX1 INVX1_479 ( .A(b_reg_2_), .Y(_abc_15724_n3848) );
  INVX1 INVX1_48 ( .A(_abc_15724_n959), .Y(_abc_15724_n960) );
  INVX1 INVX1_480 ( .A(_abc_15724_n3851), .Y(_abc_15724_n3852) );
  INVX1 INVX1_481 ( .A(d_reg_2_), .Y(_abc_15724_n3854) );
  INVX1 INVX1_482 ( .A(_abc_15724_n3850), .Y(_abc_15724_n3858) );
  INVX1 INVX1_483 ( .A(_abc_15724_n3869), .Y(_abc_15724_n3870) );
  INVX1 INVX1_484 ( .A(_abc_15724_n3872), .Y(_abc_15724_n3873) );
  INVX1 INVX1_485 ( .A(_abc_15724_n3867), .Y(_abc_15724_n3877) );
  INVX1 INVX1_486 ( .A(_abc_15724_n3874), .Y(_abc_15724_n3878) );
  INVX1 INVX1_487 ( .A(_abc_15724_n3855), .Y(_abc_15724_n3884) );
  INVX1 INVX1_488 ( .A(_abc_15724_n3862), .Y(_abc_15724_n3887) );
  INVX1 INVX1_489 ( .A(_abc_15724_n3863), .Y(_abc_15724_n3888) );
  INVX1 INVX1_49 ( .A(_abc_15724_n961), .Y(_abc_15724_n963) );
  INVX1 INVX1_490 ( .A(_abc_15724_n3876), .Y(_abc_15724_n3892) );
  INVX1 INVX1_491 ( .A(_abc_15724_n3821), .Y(_abc_15724_n3911) );
  INVX1 INVX1_492 ( .A(_abc_15724_n3917), .Y(_abc_15724_n3918) );
  INVX1 INVX1_493 ( .A(_abc_15724_n3920), .Y(_abc_15724_n3928) );
  INVX1 INVX1_494 ( .A(_abc_15724_n3897), .Y(_abc_15724_n3930) );
  INVX1 INVX1_495 ( .A(d_reg_3_), .Y(_abc_15724_n3933) );
  INVX1 INVX1_496 ( .A(c_reg_3_), .Y(_abc_15724_n3934) );
  INVX1 INVX1_497 ( .A(b_reg_3_), .Y(_abc_15724_n3935) );
  INVX1 INVX1_498 ( .A(_abc_15724_n3939), .Y(_abc_15724_n3940) );
  INVX1 INVX1_499 ( .A(_abc_15724_n3937), .Y(_abc_15724_n3944) );
  INVX1 INVX1_5 ( .A(_abc_15724_n716), .Y(_abc_15724_n717) );
  INVX1 INVX1_50 ( .A(_abc_15724_n969), .Y(_abc_15724_n970) );
  INVX1 INVX1_500 ( .A(_abc_15724_n3948), .Y(_abc_15724_n3949) );
  INVX1 INVX1_501 ( .A(_abc_15724_n3950), .Y(_abc_15724_n3951) );
  INVX1 INVX1_502 ( .A(_abc_15724_n3957), .Y(_abc_15724_n3958) );
  INVX1 INVX1_503 ( .A(_abc_15724_n3960), .Y(_abc_15724_n3961) );
  INVX1 INVX1_504 ( .A(_abc_15724_n3964), .Y(_abc_15724_n3965) );
  INVX1 INVX1_505 ( .A(_abc_15724_n3941), .Y(_abc_15724_n3969) );
  INVX1 INVX1_506 ( .A(_abc_15724_n3955), .Y(_abc_15724_n3975) );
  INVX1 INVX1_507 ( .A(_abc_15724_n3962), .Y(_abc_15724_n3976) );
  INVX1 INVX1_508 ( .A(_abc_15724_n4001), .Y(_abc_15724_n4002) );
  INVX1 INVX1_509 ( .A(_abc_15724_n3929), .Y(_abc_15724_n4006) );
  INVX1 INVX1_51 ( .A(_abc_15724_n978), .Y(_abc_15724_n979_1) );
  INVX1 INVX1_510 ( .A(_abc_15724_n3995), .Y(_abc_15724_n4016) );
  INVX1 INVX1_511 ( .A(_abc_15724_n4018), .Y(_abc_15724_n4019) );
  INVX1 INVX1_512 ( .A(d_reg_4_), .Y(_abc_15724_n4024) );
  INVX1 INVX1_513 ( .A(c_reg_4_), .Y(_abc_15724_n4025) );
  INVX1 INVX1_514 ( .A(b_reg_4_), .Y(_abc_15724_n4026) );
  INVX1 INVX1_515 ( .A(_abc_15724_n4031), .Y(_abc_15724_n4032) );
  INVX1 INVX1_516 ( .A(_abc_15724_n4028), .Y(_abc_15724_n4035) );
  INVX1 INVX1_517 ( .A(_abc_15724_n4046), .Y(_abc_15724_n4047) );
  INVX1 INVX1_518 ( .A(_abc_15724_n4049), .Y(_abc_15724_n4050) );
  INVX1 INVX1_519 ( .A(_abc_15724_n4044), .Y(_abc_15724_n4054) );
  INVX1 INVX1_52 ( .A(e_reg_31_), .Y(_abc_15724_n986) );
  INVX1 INVX1_520 ( .A(_abc_15724_n4051), .Y(_abc_15724_n4055) );
  INVX1 INVX1_521 ( .A(_abc_15724_n4030), .Y(_abc_15724_n4060) );
  INVX1 INVX1_522 ( .A(_abc_15724_n4039), .Y(_abc_15724_n4063) );
  INVX1 INVX1_523 ( .A(_abc_15724_n4040), .Y(_abc_15724_n4064) );
  INVX1 INVX1_524 ( .A(_abc_15724_n4053), .Y(_abc_15724_n4068) );
  INVX1 INVX1_525 ( .A(_abc_15724_n4086), .Y(_abc_15724_n4087) );
  INVX1 INVX1_526 ( .A(_abc_15724_n4089), .Y(_abc_15724_n4090) );
  INVX1 INVX1_527 ( .A(_abc_15724_n4092), .Y(_abc_15724_n4093) );
  INVX1 INVX1_528 ( .A(d_reg_5_), .Y(_abc_15724_n4103) );
  INVX1 INVX1_529 ( .A(c_reg_5_), .Y(_abc_15724_n4104) );
  INVX1 INVX1_53 ( .A(_auto_iopadmap_cc_313_execute_26059_31_), .Y(_abc_15724_n988_1) );
  INVX1 INVX1_530 ( .A(b_reg_5_), .Y(_abc_15724_n4105) );
  INVX1 INVX1_531 ( .A(_abc_15724_n4110), .Y(_abc_15724_n4111) );
  INVX1 INVX1_532 ( .A(_abc_15724_n4107), .Y(_abc_15724_n4114) );
  INVX1 INVX1_533 ( .A(_abc_15724_n4125), .Y(_abc_15724_n4126) );
  INVX1 INVX1_534 ( .A(_abc_15724_n4128), .Y(_abc_15724_n4129) );
  INVX1 INVX1_535 ( .A(_abc_15724_n4123), .Y(_abc_15724_n4133) );
  INVX1 INVX1_536 ( .A(_abc_15724_n4130), .Y(_abc_15724_n4134) );
  INVX1 INVX1_537 ( .A(_abc_15724_n4109), .Y(_abc_15724_n4139) );
  INVX1 INVX1_538 ( .A(_abc_15724_n4118), .Y(_abc_15724_n4142) );
  INVX1 INVX1_539 ( .A(_abc_15724_n4119), .Y(_abc_15724_n4143) );
  INVX1 INVX1_54 ( .A(_abc_15724_n990), .Y(_abc_15724_n991) );
  INVX1 INVX1_540 ( .A(_abc_15724_n4132), .Y(_abc_15724_n4147) );
  INVX1 INVX1_541 ( .A(_abc_15724_n4172), .Y(_abc_15724_n4173) );
  INVX1 INVX1_542 ( .A(_abc_15724_n4176), .Y(_abc_15724_n4177) );
  INVX1 INVX1_543 ( .A(_abc_15724_n4178), .Y(_abc_15724_n4179) );
  INVX1 INVX1_544 ( .A(_abc_15724_n4165), .Y(_abc_15724_n4189) );
  INVX1 INVX1_545 ( .A(_abc_15724_n4191), .Y(_abc_15724_n4192) );
  INVX1 INVX1_546 ( .A(_abc_15724_n4193), .Y(_abc_15724_n4194) );
  INVX1 INVX1_547 ( .A(d_reg_6_), .Y(_abc_15724_n4196) );
  INVX1 INVX1_548 ( .A(c_reg_6_), .Y(_abc_15724_n4197) );
  INVX1 INVX1_549 ( .A(b_reg_6_), .Y(_abc_15724_n4198) );
  INVX1 INVX1_55 ( .A(_abc_15724_n985), .Y(_abc_15724_n993) );
  INVX1 INVX1_550 ( .A(_abc_15724_n4202), .Y(_abc_15724_n4203) );
  INVX1 INVX1_551 ( .A(_abc_15724_n4210), .Y(_abc_15724_n4211) );
  INVX1 INVX1_552 ( .A(_abc_15724_n4200), .Y(_abc_15724_n4212) );
  INVX1 INVX1_553 ( .A(_abc_15724_n4214), .Y(_abc_15724_n4215) );
  INVX1 INVX1_554 ( .A(_abc_15724_n4218), .Y(_abc_15724_n4219) );
  INVX1 INVX1_555 ( .A(_abc_15724_n4220), .Y(_abc_15724_n4221) );
  INVX1 INVX1_556 ( .A(_abc_15724_n4223), .Y(_abc_15724_n4224) );
  INVX1 INVX1_557 ( .A(_abc_15724_n4226), .Y(_abc_15724_n4227) );
  INVX1 INVX1_558 ( .A(_abc_15724_n4229), .Y(_abc_15724_n4231) );
  INVX1 INVX1_559 ( .A(_abc_15724_n4230), .Y(_abc_15724_n4235) );
  INVX1 INVX1_56 ( .A(_abc_15724_n1001), .Y(_abc_15724_n1002) );
  INVX1 INVX1_560 ( .A(_abc_15724_n4232), .Y(_abc_15724_n4236) );
  INVX1 INVX1_561 ( .A(_abc_15724_n4195), .Y(_abc_15724_n4241) );
  INVX1 INVX1_562 ( .A(_abc_15724_n4258), .Y(_abc_15724_n4259) );
  INVX1 INVX1_563 ( .A(_abc_15724_n4260), .Y(_abc_15724_n4261) );
  INVX1 INVX1_564 ( .A(_abc_15724_n4253), .Y(_abc_15724_n4270) );
  INVX1 INVX1_565 ( .A(_abc_15724_n4271), .Y(_abc_15724_n4272) );
  INVX1 INVX1_566 ( .A(_abc_15724_n4274), .Y(_abc_15724_n4275) );
  INVX1 INVX1_567 ( .A(d_reg_7_), .Y(_abc_15724_n4276) );
  INVX1 INVX1_568 ( .A(c_reg_7_), .Y(_abc_15724_n4277) );
  INVX1 INVX1_569 ( .A(b_reg_7_), .Y(_abc_15724_n4278) );
  INVX1 INVX1_57 ( .A(_auto_iopadmap_cc_313_execute_26059_33_), .Y(_abc_15724_n1008) );
  INVX1 INVX1_570 ( .A(_abc_15724_n4283), .Y(_abc_15724_n4284) );
  INVX1 INVX1_571 ( .A(_abc_15724_n4280), .Y(_abc_15724_n4287) );
  INVX1 INVX1_572 ( .A(_abc_15724_n4298), .Y(_abc_15724_n4299) );
  INVX1 INVX1_573 ( .A(_abc_15724_n4301), .Y(_abc_15724_n4302) );
  INVX1 INVX1_574 ( .A(_abc_15724_n4296), .Y(_abc_15724_n4306) );
  INVX1 INVX1_575 ( .A(_abc_15724_n4303), .Y(_abc_15724_n4307) );
  INVX1 INVX1_576 ( .A(_abc_15724_n4282), .Y(_abc_15724_n4312) );
  INVX1 INVX1_577 ( .A(_abc_15724_n4291), .Y(_abc_15724_n4315) );
  INVX1 INVX1_578 ( .A(_abc_15724_n4292), .Y(_abc_15724_n4316) );
  INVX1 INVX1_579 ( .A(_abc_15724_n4305), .Y(_abc_15724_n4320) );
  INVX1 INVX1_58 ( .A(d_reg_1_), .Y(_abc_15724_n1009) );
  INVX1 INVX1_580 ( .A(_abc_15724_n4324), .Y(_abc_15724_n4325) );
  INVX1 INVX1_581 ( .A(_abc_15724_n4328), .Y(_abc_15724_n4331) );
  INVX1 INVX1_582 ( .A(_abc_15724_n4333), .Y(_abc_15724_n4334) );
  INVX1 INVX1_583 ( .A(_abc_15724_n4329), .Y(_abc_15724_n4348) );
  INVX1 INVX1_584 ( .A(_abc_15724_n4352), .Y(_abc_15724_n4353) );
  INVX1 INVX1_585 ( .A(d_reg_8_), .Y(_abc_15724_n4356) );
  INVX1 INVX1_586 ( .A(c_reg_8_), .Y(_abc_15724_n4357) );
  INVX1 INVX1_587 ( .A(b_reg_8_), .Y(_abc_15724_n4358) );
  INVX1 INVX1_588 ( .A(_abc_15724_n4363), .Y(_abc_15724_n4364) );
  INVX1 INVX1_589 ( .A(_abc_15724_n4360), .Y(_abc_15724_n4367) );
  INVX1 INVX1_59 ( .A(_abc_15724_n1011), .Y(_abc_15724_n1015_1) );
  INVX1 INVX1_590 ( .A(_abc_15724_n4378), .Y(_abc_15724_n4379) );
  INVX1 INVX1_591 ( .A(_abc_15724_n4381), .Y(_abc_15724_n4382) );
  INVX1 INVX1_592 ( .A(_abc_15724_n4376), .Y(_abc_15724_n4386) );
  INVX1 INVX1_593 ( .A(_abc_15724_n4383), .Y(_abc_15724_n4387) );
  INVX1 INVX1_594 ( .A(_abc_15724_n4362), .Y(_abc_15724_n4392) );
  INVX1 INVX1_595 ( .A(_abc_15724_n4371), .Y(_abc_15724_n4395) );
  INVX1 INVX1_596 ( .A(_abc_15724_n4372), .Y(_abc_15724_n4396) );
  INVX1 INVX1_597 ( .A(_abc_15724_n4385), .Y(_abc_15724_n4400) );
  INVX1 INVX1_598 ( .A(_abc_15724_n4418), .Y(_abc_15724_n4419) );
  INVX1 INVX1_599 ( .A(_abc_15724_n4421), .Y(_abc_15724_n4422) );
  INVX1 INVX1_6 ( .A(_abc_15724_n719_1), .Y(_abc_15724_n720) );
  INVX1 INVX1_60 ( .A(_abc_15724_n1025_1), .Y(_abc_15724_n1026_1) );
  INVX1 INVX1_600 ( .A(_abc_15724_n4423), .Y(_abc_15724_n4424) );
  INVX1 INVX1_601 ( .A(d_reg_9_), .Y(_abc_15724_n4434) );
  INVX1 INVX1_602 ( .A(c_reg_9_), .Y(_abc_15724_n4435) );
  INVX1 INVX1_603 ( .A(b_reg_9_), .Y(_abc_15724_n4436) );
  INVX1 INVX1_604 ( .A(_abc_15724_n4441), .Y(_abc_15724_n4442) );
  INVX1 INVX1_605 ( .A(_abc_15724_n4438), .Y(_abc_15724_n4445) );
  INVX1 INVX1_606 ( .A(_abc_15724_n4456), .Y(_abc_15724_n4457) );
  INVX1 INVX1_607 ( .A(_abc_15724_n4459), .Y(_abc_15724_n4460) );
  INVX1 INVX1_608 ( .A(_abc_15724_n4454), .Y(_abc_15724_n4464) );
  INVX1 INVX1_609 ( .A(_abc_15724_n4461), .Y(_abc_15724_n4465) );
  INVX1 INVX1_61 ( .A(_abc_15724_n1027), .Y(_abc_15724_n1028) );
  INVX1 INVX1_610 ( .A(_abc_15724_n4440), .Y(_abc_15724_n4470) );
  INVX1 INVX1_611 ( .A(_abc_15724_n4449), .Y(_abc_15724_n4473) );
  INVX1 INVX1_612 ( .A(_abc_15724_n4450), .Y(_abc_15724_n4474) );
  INVX1 INVX1_613 ( .A(_abc_15724_n4463), .Y(_abc_15724_n4478) );
  INVX1 INVX1_614 ( .A(_abc_15724_n4503), .Y(_abc_15724_n4504) );
  INVX1 INVX1_615 ( .A(_abc_15724_n4505), .Y(_abc_15724_n4506) );
  INVX1 INVX1_616 ( .A(_abc_15724_n4496), .Y(_abc_15724_n4517) );
  INVX1 INVX1_617 ( .A(_abc_15724_n4518), .Y(_abc_15724_n4519) );
  INVX1 INVX1_618 ( .A(_abc_15724_n4521), .Y(_abc_15724_n4522) );
  INVX1 INVX1_619 ( .A(d_reg_10_), .Y(_abc_15724_n4524) );
  INVX1 INVX1_62 ( .A(_abc_15724_n1040), .Y(_abc_15724_n1041) );
  INVX1 INVX1_620 ( .A(c_reg_10_), .Y(_abc_15724_n4525) );
  INVX1 INVX1_621 ( .A(b_reg_10_), .Y(_abc_15724_n4526) );
  INVX1 INVX1_622 ( .A(_abc_15724_n4530), .Y(_abc_15724_n4531) );
  INVX1 INVX1_623 ( .A(_abc_15724_n4534), .Y(_abc_15724_n4535) );
  INVX1 INVX1_624 ( .A(_abc_15724_n4528), .Y(_abc_15724_n4540) );
  INVX1 INVX1_625 ( .A(_abc_15724_n4546), .Y(_abc_15724_n4547) );
  INVX1 INVX1_626 ( .A(_abc_15724_n4549), .Y(_abc_15724_n4550) );
  INVX1 INVX1_627 ( .A(_abc_15724_n4552), .Y(_abc_15724_n4553) );
  INVX1 INVX1_628 ( .A(_abc_15724_n4557), .Y(_abc_15724_n4558) );
  INVX1 INVX1_629 ( .A(_abc_15724_n4544), .Y(_abc_15724_n4561) );
  INVX1 INVX1_63 ( .A(_abc_15724_n1042), .Y(_abc_15724_n1043) );
  INVX1 INVX1_630 ( .A(_abc_15724_n4556), .Y(_abc_15724_n4563) );
  INVX1 INVX1_631 ( .A(_abc_15724_n4523), .Y(_abc_15724_n4568) );
  INVX1 INVX1_632 ( .A(_abc_15724_n4585), .Y(_abc_15724_n4586) );
  INVX1 INVX1_633 ( .A(_abc_15724_n4587), .Y(_abc_15724_n4588) );
  INVX1 INVX1_634 ( .A(_abc_15724_n4580), .Y(_abc_15724_n4597) );
  INVX1 INVX1_635 ( .A(d_reg_11_), .Y(_abc_15724_n4601) );
  INVX1 INVX1_636 ( .A(c_reg_11_), .Y(_abc_15724_n4602) );
  INVX1 INVX1_637 ( .A(b_reg_11_), .Y(_abc_15724_n4603) );
  INVX1 INVX1_638 ( .A(_abc_15724_n4607), .Y(_abc_15724_n4608) );
  INVX1 INVX1_639 ( .A(_abc_15724_n4605), .Y(_abc_15724_n4616) );
  INVX1 INVX1_64 ( .A(_abc_15724_n1053), .Y(_abc_15724_n1054) );
  INVX1 INVX1_640 ( .A(_abc_15724_n4620), .Y(_abc_15724_n4621) );
  INVX1 INVX1_641 ( .A(_abc_15724_n4623), .Y(_abc_15724_n4624) );
  INVX1 INVX1_642 ( .A(_abc_15724_n4626), .Y(_abc_15724_n4627) );
  INVX1 INVX1_643 ( .A(_abc_15724_n4629), .Y(_abc_15724_n4630) );
  INVX1 INVX1_644 ( .A(_abc_15724_n4633), .Y(_abc_15724_n4634) );
  INVX1 INVX1_645 ( .A(_abc_15724_n4611), .Y(_abc_15724_n4638) );
  INVX1 INVX1_646 ( .A(_abc_15724_n4635), .Y(_abc_15724_n4640) );
  INVX1 INVX1_647 ( .A(_abc_15724_n4598), .Y(_abc_15724_n4665) );
  INVX1 INVX1_648 ( .A(_abc_15724_n4663), .Y(_abc_15724_n4666) );
  INVX1 INVX1_649 ( .A(_abc_15724_n4657), .Y(_abc_15724_n4679) );
  INVX1 INVX1_65 ( .A(_abc_15724_n1055), .Y(_abc_15724_n1056) );
  INVX1 INVX1_650 ( .A(_abc_15724_n4684), .Y(_abc_15724_n4685) );
  INVX1 INVX1_651 ( .A(d_reg_12_), .Y(_abc_15724_n4688) );
  INVX1 INVX1_652 ( .A(c_reg_12_), .Y(_abc_15724_n4689) );
  INVX1 INVX1_653 ( .A(b_reg_12_), .Y(_abc_15724_n4690) );
  INVX1 INVX1_654 ( .A(_abc_15724_n4694), .Y(_abc_15724_n4695) );
  INVX1 INVX1_655 ( .A(_abc_15724_n4698), .Y(_abc_15724_n4699) );
  INVX1 INVX1_656 ( .A(_abc_15724_n4692), .Y(_abc_15724_n4704) );
  INVX1 INVX1_657 ( .A(_abc_15724_n4709), .Y(_abc_15724_n4710) );
  INVX1 INVX1_658 ( .A(_abc_15724_n4711), .Y(_abc_15724_n4712) );
  INVX1 INVX1_659 ( .A(_abc_15724_n4714), .Y(_abc_15724_n4715) );
  INVX1 INVX1_66 ( .A(_abc_15724_n1039_1), .Y(_abc_15724_n1057) );
  INVX1 INVX1_660 ( .A(_abc_15724_n4717), .Y(_abc_15724_n4718) );
  INVX1 INVX1_661 ( .A(_abc_15724_n4721), .Y(_abc_15724_n4722) );
  INVX1 INVX1_662 ( .A(_abc_15724_n4723), .Y(_abc_15724_n4726) );
  INVX1 INVX1_663 ( .A(_abc_15724_n4743), .Y(_abc_15724_n4744) );
  INVX1 INVX1_664 ( .A(_abc_15724_n4746), .Y(_abc_15724_n4747) );
  INVX1 INVX1_665 ( .A(_abc_15724_n4749), .Y(_abc_15724_n4750) );
  INVX1 INVX1_666 ( .A(d_reg_13_), .Y(_abc_15724_n4760) );
  INVX1 INVX1_667 ( .A(c_reg_13_), .Y(_abc_15724_n4761) );
  INVX1 INVX1_668 ( .A(b_reg_13_), .Y(_abc_15724_n4762) );
  INVX1 INVX1_669 ( .A(_abc_15724_n4766), .Y(_abc_15724_n4767) );
  INVX1 INVX1_67 ( .A(_abc_15724_n1072), .Y(_abc_15724_n1073) );
  INVX1 INVX1_670 ( .A(_abc_15724_n4770), .Y(_abc_15724_n4771) );
  INVX1 INVX1_671 ( .A(_abc_15724_n4764), .Y(_abc_15724_n4776) );
  INVX1 INVX1_672 ( .A(_abc_15724_n4782), .Y(_abc_15724_n4783) );
  INVX1 INVX1_673 ( .A(_abc_15724_n4785), .Y(_abc_15724_n4786) );
  INVX1 INVX1_674 ( .A(_abc_15724_n4788), .Y(_abc_15724_n4789) );
  INVX1 INVX1_675 ( .A(_abc_15724_n4793), .Y(_abc_15724_n4794) );
  INVX1 INVX1_676 ( .A(_abc_15724_n4781), .Y(_abc_15724_n4797) );
  INVX1 INVX1_677 ( .A(_abc_15724_n4792), .Y(_abc_15724_n4798) );
  INVX1 INVX1_678 ( .A(_abc_15724_n4822), .Y(_abc_15724_n4823) );
  INVX1 INVX1_679 ( .A(_abc_15724_n4826), .Y(_abc_15724_n4827) );
  INVX1 INVX1_68 ( .A(_abc_15724_n1074), .Y(_abc_15724_n1077) );
  INVX1 INVX1_680 ( .A(_abc_15724_n4828), .Y(_abc_15724_n4829) );
  INVX1 INVX1_681 ( .A(_abc_15724_n4815), .Y(_abc_15724_n4838) );
  INVX1 INVX1_682 ( .A(_abc_15724_n4840), .Y(_abc_15724_n4841) );
  INVX1 INVX1_683 ( .A(_abc_15724_n4842), .Y(_abc_15724_n4843) );
  INVX1 INVX1_684 ( .A(d_reg_14_), .Y(_abc_15724_n4845) );
  INVX1 INVX1_685 ( .A(c_reg_14_), .Y(_abc_15724_n4846) );
  INVX1 INVX1_686 ( .A(b_reg_14_), .Y(_abc_15724_n4847) );
  INVX1 INVX1_687 ( .A(_abc_15724_n4849), .Y(_abc_15724_n4852) );
  INVX1 INVX1_688 ( .A(_abc_15724_n4854), .Y(_abc_15724_n4855) );
  INVX1 INVX1_689 ( .A(_abc_15724_n4862), .Y(_abc_15724_n4863) );
  INVX1 INVX1_69 ( .A(_abc_15724_n1087), .Y(_abc_15724_n1088) );
  INVX1 INVX1_690 ( .A(_abc_15724_n4866), .Y(_abc_15724_n4867) );
  INVX1 INVX1_691 ( .A(_abc_15724_n4869), .Y(_abc_15724_n4870) );
  INVX1 INVX1_692 ( .A(_abc_15724_n4872), .Y(_abc_15724_n4873) );
  INVX1 INVX1_693 ( .A(_abc_15724_n4876), .Y(_abc_15724_n4877) );
  INVX1 INVX1_694 ( .A(_abc_15724_n4879), .Y(_abc_15724_n4880) );
  INVX1 INVX1_695 ( .A(_abc_15724_n4882), .Y(_abc_15724_n4883) );
  INVX1 INVX1_696 ( .A(_abc_15724_n4844), .Y(_abc_15724_n4886) );
  INVX1 INVX1_697 ( .A(_abc_15724_n4881), .Y(_abc_15724_n4887) );
  INVX1 INVX1_698 ( .A(_abc_15724_n4902), .Y(_abc_15724_n4903) );
  INVX1 INVX1_699 ( .A(_abc_15724_n4904), .Y(_abc_15724_n4905) );
  INVX1 INVX1_7 ( .A(_abc_15724_n722), .Y(_abc_15724_n723) );
  INVX1 INVX1_70 ( .A(_abc_15724_n1089), .Y(_abc_15724_n1092_1) );
  INVX1 INVX1_700 ( .A(_abc_15724_n4897), .Y(_abc_15724_n4914) );
  INVX1 INVX1_701 ( .A(_abc_15724_n4915), .Y(_abc_15724_n4916) );
  INVX1 INVX1_702 ( .A(_abc_15724_n4918), .Y(_abc_15724_n4919) );
  INVX1 INVX1_703 ( .A(_abc_15724_n4920), .Y(_abc_15724_n4921) );
  INVX1 INVX1_704 ( .A(d_reg_15_), .Y(_abc_15724_n4922) );
  INVX1 INVX1_705 ( .A(_abc_15724_n4929), .Y(_abc_15724_n4930) );
  INVX1 INVX1_706 ( .A(_abc_15724_n4932), .Y(_abc_15724_n4933) );
  INVX1 INVX1_707 ( .A(_abc_15724_n4926), .Y(_abc_15724_n4935) );
  INVX1 INVX1_708 ( .A(_abc_15724_n4943), .Y(_abc_15724_n4944) );
  INVX1 INVX1_709 ( .A(_abc_15724_n4946), .Y(_abc_15724_n4947) );
  INVX1 INVX1_71 ( .A(_abc_15724_n1101), .Y(_abc_15724_n1102) );
  INVX1 INVX1_710 ( .A(_abc_15724_n4950), .Y(_abc_15724_n4951) );
  INVX1 INVX1_711 ( .A(_abc_15724_n4953), .Y(_abc_15724_n4954) );
  INVX1 INVX1_712 ( .A(_abc_15724_n4925), .Y(_abc_15724_n4956) );
  INVX1 INVX1_713 ( .A(_abc_15724_n4938), .Y(_abc_15724_n4957) );
  INVX1 INVX1_714 ( .A(_abc_15724_n4980), .Y(_abc_15724_n4981) );
  INVX1 INVX1_715 ( .A(_abc_15724_n4979), .Y(_abc_15724_n4996) );
  INVX1 INVX1_716 ( .A(_abc_15724_n4998), .Y(_abc_15724_n4999) );
  INVX1 INVX1_717 ( .A(_abc_15724_n5003), .Y(_abc_15724_n5004) );
  INVX1 INVX1_718 ( .A(_abc_15724_n5007), .Y(_abc_15724_n5008) );
  INVX1 INVX1_719 ( .A(c_reg_16_), .Y(_abc_15724_n5009) );
  INVX1 INVX1_72 ( .A(_abc_15724_n1103), .Y(_abc_15724_n1107) );
  INVX1 INVX1_720 ( .A(b_reg_16_), .Y(_abc_15724_n5010) );
  INVX1 INVX1_721 ( .A(_abc_15724_n5011), .Y(_abc_15724_n5012) );
  INVX1 INVX1_722 ( .A(_abc_15724_n5013), .Y(_abc_15724_n5014) );
  INVX1 INVX1_723 ( .A(_abc_15724_n5019), .Y(_abc_15724_n5020) );
  INVX1 INVX1_724 ( .A(_abc_15724_n5022), .Y(_abc_15724_n5023) );
  INVX1 INVX1_725 ( .A(_abc_15724_n5017), .Y(_abc_15724_n5024) );
  INVX1 INVX1_726 ( .A(_abc_15724_n5028), .Y(_abc_15724_n5029) );
  INVX1 INVX1_727 ( .A(_abc_15724_n5032), .Y(_abc_15724_n5033) );
  INVX1 INVX1_728 ( .A(_abc_15724_n5035), .Y(_abc_15724_n5036) );
  INVX1 INVX1_729 ( .A(_abc_15724_n5038), .Y(_abc_15724_n5039) );
  INVX1 INVX1_73 ( .A(_abc_15724_n1117), .Y(_abc_15724_n1118) );
  INVX1 INVX1_730 ( .A(_abc_15724_n5042), .Y(_abc_15724_n5043) );
  INVX1 INVX1_731 ( .A(_abc_15724_n5045), .Y(_abc_15724_n5046) );
  INVX1 INVX1_732 ( .A(_abc_15724_n5048), .Y(_abc_15724_n5049) );
  INVX1 INVX1_733 ( .A(_abc_15724_n5050), .Y(_abc_15724_n5051) );
  INVX1 INVX1_734 ( .A(_abc_15724_n5006), .Y(_abc_15724_n5056) );
  INVX1 INVX1_735 ( .A(_abc_15724_n5054), .Y(_abc_15724_n5057) );
  INVX1 INVX1_736 ( .A(_abc_15724_n5060), .Y(_abc_15724_n5061) );
  INVX1 INVX1_737 ( .A(_abc_15724_n5063), .Y(_abc_15724_n5064) );
  INVX1 INVX1_738 ( .A(_abc_15724_n5066), .Y(_abc_15724_n5067) );
  INVX1 INVX1_739 ( .A(_abc_15724_n5052), .Y(_abc_15724_n5074) );
  INVX1 INVX1_74 ( .A(_abc_15724_n1121_1), .Y(_abc_15724_n1122) );
  INVX1 INVX1_740 ( .A(_abc_15724_n5077), .Y(_abc_15724_n5078) );
  INVX1 INVX1_741 ( .A(_abc_15724_n5079), .Y(_abc_15724_n5080) );
  INVX1 INVX1_742 ( .A(d_reg_17_), .Y(_abc_15724_n5081) );
  INVX1 INVX1_743 ( .A(_abc_15724_n5084), .Y(_abc_15724_n5085) );
  INVX1 INVX1_744 ( .A(_abc_15724_n5089), .Y(_abc_15724_n5090) );
  INVX1 INVX1_745 ( .A(_abc_15724_n5099), .Y(_abc_15724_n5100) );
  INVX1 INVX1_746 ( .A(_abc_15724_n5102), .Y(_abc_15724_n5103) );
  INVX1 INVX1_747 ( .A(_abc_15724_n5105), .Y(_abc_15724_n5106) );
  INVX1 INVX1_748 ( .A(_abc_15724_n5109), .Y(_abc_15724_n5110) );
  INVX1 INVX1_749 ( .A(_abc_15724_n5113), .Y(_abc_15724_n5114) );
  INVX1 INVX1_75 ( .A(_abc_15724_n1127), .Y(_abc_15724_n1128) );
  INVX1 INVX1_750 ( .A(_abc_15724_n5117), .Y(_abc_15724_n5118) );
  INVX1 INVX1_751 ( .A(_abc_15724_n5120), .Y(_abc_15724_n5121) );
  INVX1 INVX1_752 ( .A(_abc_15724_n5126), .Y(_abc_15724_n5127) );
  INVX1 INVX1_753 ( .A(_abc_15724_n5130), .Y(_abc_15724_n5131) );
  INVX1 INVX1_754 ( .A(_abc_15724_n5140), .Y(_abc_15724_n5141) );
  INVX1 INVX1_755 ( .A(_abc_15724_n5143), .Y(_abc_15724_n5144) );
  INVX1 INVX1_756 ( .A(d_reg_18_), .Y(_abc_15724_n5145) );
  INVX1 INVX1_757 ( .A(c_reg_18_), .Y(_abc_15724_n5146) );
  INVX1 INVX1_758 ( .A(b_reg_18_), .Y(_abc_15724_n5147) );
  INVX1 INVX1_759 ( .A(_abc_15724_n5149), .Y(_abc_15724_n5152) );
  INVX1 INVX1_76 ( .A(_abc_15724_n1130), .Y(_abc_15724_n1131_1) );
  INVX1 INVX1_760 ( .A(_abc_15724_n5154), .Y(_abc_15724_n5155) );
  INVX1 INVX1_761 ( .A(_abc_15724_n5162), .Y(_abc_15724_n5163) );
  INVX1 INVX1_762 ( .A(_abc_15724_n5166), .Y(_abc_15724_n5167) );
  INVX1 INVX1_763 ( .A(_abc_15724_n5169), .Y(_abc_15724_n5170) );
  INVX1 INVX1_764 ( .A(_abc_15724_n5172), .Y(_abc_15724_n5173) );
  INVX1 INVX1_765 ( .A(_abc_15724_n5176), .Y(_abc_15724_n5177) );
  INVX1 INVX1_766 ( .A(_abc_15724_n5179), .Y(_abc_15724_n5180) );
  INVX1 INVX1_767 ( .A(_abc_15724_n5182), .Y(_abc_15724_n5183) );
  INVX1 INVX1_768 ( .A(_abc_15724_n5184), .Y(_abc_15724_n5185) );
  INVX1 INVX1_769 ( .A(_abc_15724_n5188), .Y(_abc_15724_n5189) );
  INVX1 INVX1_77 ( .A(_abc_15724_n1133_1), .Y(_abc_15724_n1134) );
  INVX1 INVX1_770 ( .A(_abc_15724_n5142), .Y(_abc_15724_n5191) );
  INVX1 INVX1_771 ( .A(_abc_15724_n5193), .Y(_abc_15724_n5194) );
  INVX1 INVX1_772 ( .A(_abc_15724_n5190), .Y(_abc_15724_n5203) );
  INVX1 INVX1_773 ( .A(_abc_15724_n5204), .Y(_abc_15724_n5205) );
  INVX1 INVX1_774 ( .A(_abc_15724_n5206), .Y(_abc_15724_n5207) );
  INVX1 INVX1_775 ( .A(d_reg_19_), .Y(_abc_15724_n5208) );
  INVX1 INVX1_776 ( .A(c_reg_19_), .Y(_abc_15724_n5209) );
  INVX1 INVX1_777 ( .A(b_reg_19_), .Y(_abc_15724_n5210) );
  INVX1 INVX1_778 ( .A(_abc_15724_n5214), .Y(_abc_15724_n5215) );
  INVX1 INVX1_779 ( .A(_abc_15724_n5218), .Y(_abc_15724_n5219) );
  INVX1 INVX1_78 ( .A(_abc_15724_n1139), .Y(_abc_15724_n1140) );
  INVX1 INVX1_780 ( .A(_abc_15724_n5212), .Y(_abc_15724_n5220) );
  INVX1 INVX1_781 ( .A(_abc_15724_n5229), .Y(_abc_15724_n5230) );
  INVX1 INVX1_782 ( .A(_abc_15724_n5232), .Y(_abc_15724_n5233) );
  INVX1 INVX1_783 ( .A(_abc_15724_n5235), .Y(_abc_15724_n5236) );
  INVX1 INVX1_784 ( .A(_abc_15724_n5239), .Y(_abc_15724_n5240) );
  INVX1 INVX1_785 ( .A(_abc_15724_n5242), .Y(_abc_15724_n5243) );
  INVX1 INVX1_786 ( .A(_abc_15724_n5244), .Y(_abc_15724_n5245) );
  INVX1 INVX1_787 ( .A(_abc_15724_n5248), .Y(_abc_15724_n5249) );
  INVX1 INVX1_788 ( .A(_abc_15724_n5252), .Y(_abc_15724_n5253) );
  INVX1 INVX1_789 ( .A(_abc_15724_n5186), .Y(_abc_15724_n5257) );
  INVX1 INVX1_79 ( .A(_abc_15724_n1142_1), .Y(_abc_15724_n1143) );
  INVX1 INVX1_790 ( .A(_abc_15724_n5255), .Y(_abc_15724_n5258) );
  INVX1 INVX1_791 ( .A(_abc_15724_n5260), .Y(_abc_15724_n5261) );
  INVX1 INVX1_792 ( .A(_abc_15724_n5259), .Y(_abc_15724_n5271) );
  INVX1 INVX1_793 ( .A(_abc_15724_n5273), .Y(_abc_15724_n5274) );
  INVX1 INVX1_794 ( .A(_abc_15724_n5128), .Y(_abc_15724_n5280) );
  INVX1 INVX1_795 ( .A(_abc_15724_n5284), .Y(_abc_15724_n5285) );
  INVX1 INVX1_796 ( .A(_abc_15724_n5286), .Y(_abc_15724_n5287) );
  INVX1 INVX1_797 ( .A(_abc_15724_n5288), .Y(_abc_15724_n5289) );
  INVX1 INVX1_798 ( .A(d_reg_20_), .Y(_abc_15724_n5290) );
  INVX1 INVX1_799 ( .A(c_reg_20_), .Y(_abc_15724_n5291) );
  INVX1 INVX1_8 ( .A(_abc_15724_n727), .Y(_abc_15724_n728) );
  INVX1 INVX1_80 ( .A(_abc_15724_n1146), .Y(_abc_15724_n1147) );
  INVX1 INVX1_800 ( .A(b_reg_20_), .Y(_abc_15724_n5292) );
  INVX1 INVX1_801 ( .A(_abc_15724_n5294), .Y(_abc_15724_n5297) );
  INVX1 INVX1_802 ( .A(_abc_15724_n5299), .Y(_abc_15724_n5300) );
  INVX1 INVX1_803 ( .A(_abc_15724_n5307), .Y(_abc_15724_n5308) );
  INVX1 INVX1_804 ( .A(_abc_15724_n5311), .Y(_abc_15724_n5312) );
  INVX1 INVX1_805 ( .A(_abc_15724_n5314), .Y(_abc_15724_n5315) );
  INVX1 INVX1_806 ( .A(_abc_15724_n5317), .Y(_abc_15724_n5318) );
  INVX1 INVX1_807 ( .A(_abc_15724_n5321), .Y(_abc_15724_n5322) );
  INVX1 INVX1_808 ( .A(_abc_15724_n5324), .Y(_abc_15724_n5325) );
  INVX1 INVX1_809 ( .A(_abc_15724_n5327), .Y(_abc_15724_n5328) );
  INVX1 INVX1_81 ( .A(_abc_15724_n1155_1), .Y(_abc_15724_n1156_1) );
  INVX1 INVX1_810 ( .A(_abc_15724_n5329), .Y(_abc_15724_n5330) );
  INVX1 INVX1_811 ( .A(_abc_15724_n5335), .Y(_abc_15724_n5336) );
  INVX1 INVX1_812 ( .A(_abc_15724_n5337), .Y(_abc_15724_n5338) );
  INVX1 INVX1_813 ( .A(_abc_15724_n5341), .Y(_abc_15724_n5342) );
  INVX1 INVX1_814 ( .A(_abc_15724_n5344), .Y(_abc_15724_n5352) );
  INVX1 INVX1_815 ( .A(_abc_15724_n5331), .Y(_abc_15724_n5353) );
  INVX1 INVX1_816 ( .A(_abc_15724_n5354), .Y(_abc_15724_n5355) );
  INVX1 INVX1_817 ( .A(_abc_15724_n5356), .Y(_abc_15724_n5357) );
  INVX1 INVX1_818 ( .A(d_reg_21_), .Y(_abc_15724_n5358) );
  INVX1 INVX1_819 ( .A(c_reg_21_), .Y(_abc_15724_n5359) );
  INVX1 INVX1_82 ( .A(_abc_15724_n1153), .Y(_abc_15724_n1159) );
  INVX1 INVX1_820 ( .A(b_reg_21_), .Y(_abc_15724_n5360) );
  INVX1 INVX1_821 ( .A(_abc_15724_n5362), .Y(_abc_15724_n5365) );
  INVX1 INVX1_822 ( .A(_abc_15724_n5367), .Y(_abc_15724_n5368) );
  INVX1 INVX1_823 ( .A(_abc_15724_n5375), .Y(_abc_15724_n5376) );
  INVX1 INVX1_824 ( .A(_abc_15724_n5379), .Y(_abc_15724_n5380) );
  INVX1 INVX1_825 ( .A(_abc_15724_n5382), .Y(_abc_15724_n5383) );
  INVX1 INVX1_826 ( .A(_abc_15724_n5385), .Y(_abc_15724_n5386) );
  INVX1 INVX1_827 ( .A(_abc_15724_n5389), .Y(_abc_15724_n5390) );
  INVX1 INVX1_828 ( .A(_abc_15724_n5392), .Y(_abc_15724_n5393) );
  INVX1 INVX1_829 ( .A(_abc_15724_n5394), .Y(_abc_15724_n5395) );
  INVX1 INVX1_83 ( .A(_abc_15724_n1157_1), .Y(_abc_15724_n1160) );
  INVX1 INVX1_830 ( .A(_abc_15724_n5398), .Y(_abc_15724_n5399) );
  INVX1 INVX1_831 ( .A(_abc_15724_n5401), .Y(_abc_15724_n5402) );
  INVX1 INVX1_832 ( .A(_abc_15724_n5405), .Y(_abc_15724_n5406) );
  INVX1 INVX1_833 ( .A(_abc_15724_n5409), .Y(_abc_15724_n5410) );
  INVX1 INVX1_834 ( .A(_abc_15724_n5339), .Y(_abc_15724_n5415) );
  INVX1 INVX1_835 ( .A(_abc_15724_n5407), .Y(_abc_15724_n5425) );
  INVX1 INVX1_836 ( .A(_abc_15724_n5427), .Y(_abc_15724_n5428) );
  INVX1 INVX1_837 ( .A(_abc_15724_n5404), .Y(_abc_15724_n5429) );
  INVX1 INVX1_838 ( .A(_abc_15724_n5430), .Y(_abc_15724_n5431) );
  INVX1 INVX1_839 ( .A(_abc_15724_n5432), .Y(_abc_15724_n5433) );
  INVX1 INVX1_84 ( .A(_abc_15724_n1178_1), .Y(_abc_15724_n1179_1) );
  INVX1 INVX1_840 ( .A(d_reg_22_), .Y(_abc_15724_n5434) );
  INVX1 INVX1_841 ( .A(c_reg_22_), .Y(_abc_15724_n5435) );
  INVX1 INVX1_842 ( .A(b_reg_22_), .Y(_abc_15724_n5436) );
  INVX1 INVX1_843 ( .A(_abc_15724_n5438), .Y(_abc_15724_n5441) );
  INVX1 INVX1_844 ( .A(_abc_15724_n5443), .Y(_abc_15724_n5444) );
  INVX1 INVX1_845 ( .A(_abc_15724_n5451), .Y(_abc_15724_n5452) );
  INVX1 INVX1_846 ( .A(_abc_15724_n5455), .Y(_abc_15724_n5456) );
  INVX1 INVX1_847 ( .A(_abc_15724_n5458), .Y(_abc_15724_n5459) );
  INVX1 INVX1_848 ( .A(_abc_15724_n5461), .Y(_abc_15724_n5462) );
  INVX1 INVX1_849 ( .A(_abc_15724_n5465), .Y(_abc_15724_n5466) );
  INVX1 INVX1_85 ( .A(_abc_15724_n1182), .Y(_abc_15724_n1183) );
  INVX1 INVX1_850 ( .A(_abc_15724_n5468), .Y(_abc_15724_n5469) );
  INVX1 INVX1_851 ( .A(_abc_15724_n5470), .Y(_abc_15724_n5471) );
  INVX1 INVX1_852 ( .A(_abc_15724_n5474), .Y(_abc_15724_n5475) );
  INVX1 INVX1_853 ( .A(_abc_15724_n5477), .Y(_abc_15724_n5478) );
  INVX1 INVX1_854 ( .A(_abc_15724_n5481), .Y(_abc_15724_n5482) );
  INVX1 INVX1_855 ( .A(_abc_15724_n5485), .Y(_abc_15724_n5486) );
  INVX1 INVX1_856 ( .A(_abc_15724_n5483), .Y(_abc_15724_n5495) );
  INVX1 INVX1_857 ( .A(_abc_15724_n5496), .Y(_abc_15724_n5497) );
  INVX1 INVX1_858 ( .A(_abc_15724_n5499), .Y(_abc_15724_n5500) );
  INVX1 INVX1_859 ( .A(_abc_15724_n5501), .Y(_abc_15724_n5502) );
  INVX1 INVX1_86 ( .A(_abc_15724_n1191_1), .Y(_abc_15724_n1192) );
  INVX1 INVX1_860 ( .A(d_reg_23_), .Y(_abc_15724_n5503) );
  INVX1 INVX1_861 ( .A(_abc_15724_n5506), .Y(_abc_15724_n5507) );
  INVX1 INVX1_862 ( .A(_abc_15724_n5511), .Y(_abc_15724_n5512) );
  INVX1 INVX1_863 ( .A(_abc_15724_n5521), .Y(_abc_15724_n5522) );
  INVX1 INVX1_864 ( .A(_abc_15724_n5524), .Y(_abc_15724_n5525) );
  INVX1 INVX1_865 ( .A(_abc_15724_n5527), .Y(_abc_15724_n5528) );
  INVX1 INVX1_866 ( .A(_abc_15724_n5531), .Y(_abc_15724_n5532) );
  INVX1 INVX1_867 ( .A(_abc_15724_n5535), .Y(_abc_15724_n5536) );
  INVX1 INVX1_868 ( .A(_abc_15724_n5539), .Y(_abc_15724_n5540) );
  INVX1 INVX1_869 ( .A(_abc_15724_n5543), .Y(_abc_15724_n5544) );
  INVX1 INVX1_87 ( .A(_abc_15724_n1199), .Y(_abc_15724_n1200_1) );
  INVX1 INVX1_870 ( .A(_abc_15724_n5498), .Y(_abc_15724_n5548) );
  INVX1 INVX1_871 ( .A(_abc_15724_n5546), .Y(_abc_15724_n5549) );
  INVX1 INVX1_872 ( .A(_abc_15724_n5551), .Y(_abc_15724_n5552) );
  INVX1 INVX1_873 ( .A(_abc_15724_n5547), .Y(_abc_15724_n5566) );
  INVX1 INVX1_874 ( .A(_abc_15724_n5573), .Y(_abc_15724_n5574) );
  INVX1 INVX1_875 ( .A(_abc_15724_n5575), .Y(_abc_15724_n5576) );
  INVX1 INVX1_876 ( .A(_abc_15724_n5577), .Y(_abc_15724_n5578) );
  INVX1 INVX1_877 ( .A(_abc_15724_n5579), .Y(_abc_15724_n5580) );
  INVX1 INVX1_878 ( .A(d_reg_24_), .Y(_abc_15724_n5581) );
  INVX1 INVX1_879 ( .A(_abc_15724_n5584), .Y(_abc_15724_n5585) );
  INVX1 INVX1_88 ( .A(_abc_15724_n1204), .Y(_abc_15724_n1205) );
  INVX1 INVX1_880 ( .A(_abc_15724_n5589), .Y(_abc_15724_n5590) );
  INVX1 INVX1_881 ( .A(_abc_15724_n5586), .Y(_abc_15724_n5594) );
  INVX1 INVX1_882 ( .A(_abc_15724_n5595), .Y(_abc_15724_n5596) );
  INVX1 INVX1_883 ( .A(_abc_15724_n5601), .Y(_abc_15724_n5602) );
  INVX1 INVX1_884 ( .A(_abc_15724_n5604), .Y(_abc_15724_n5605) );
  INVX1 INVX1_885 ( .A(_abc_15724_n5607), .Y(_abc_15724_n5608) );
  INVX1 INVX1_886 ( .A(_abc_15724_n5611), .Y(_abc_15724_n5612) );
  INVX1 INVX1_887 ( .A(_abc_15724_n5615), .Y(_abc_15724_n5616) );
  INVX1 INVX1_888 ( .A(_abc_15724_n5619), .Y(_abc_15724_n5620) );
  INVX1 INVX1_889 ( .A(_abc_15724_n5622), .Y(_abc_15724_n5623) );
  INVX1 INVX1_89 ( .A(_abc_15724_n1207_1), .Y(_abc_15724_n1208) );
  INVX1 INVX1_890 ( .A(_abc_15724_n5626), .Y(_abc_15724_n5627) );
  INVX1 INVX1_891 ( .A(_abc_15724_n5630), .Y(_abc_15724_n5631) );
  INVX1 INVX1_892 ( .A(_abc_15724_n5632), .Y(_abc_15724_n5633) );
  INVX1 INVX1_893 ( .A(_abc_15724_n5642), .Y(_abc_15724_n5643) );
  INVX1 INVX1_894 ( .A(_abc_15724_n5644), .Y(_abc_15724_n5645) );
  INVX1 INVX1_895 ( .A(d_reg_25_), .Y(_abc_15724_n5646) );
  INVX1 INVX1_896 ( .A(_abc_15724_n5649), .Y(_abc_15724_n5650) );
  INVX1 INVX1_897 ( .A(_abc_15724_n5654), .Y(_abc_15724_n5655) );
  INVX1 INVX1_898 ( .A(_abc_15724_n5651), .Y(_abc_15724_n5659) );
  INVX1 INVX1_899 ( .A(_abc_15724_n5660), .Y(_abc_15724_n5661) );
  INVX1 INVX1_9 ( .A(_abc_15724_n729_1), .Y(_abc_15724_n730_1) );
  INVX1 INVX1_90 ( .A(_abc_15724_n1211), .Y(_abc_15724_n1212) );
  INVX1 INVX1_900 ( .A(_abc_15724_n5666), .Y(_abc_15724_n5667) );
  INVX1 INVX1_901 ( .A(_abc_15724_n5669), .Y(_abc_15724_n5670) );
  INVX1 INVX1_902 ( .A(_abc_15724_n5672), .Y(_abc_15724_n5673) );
  INVX1 INVX1_903 ( .A(_abc_15724_n5676), .Y(_abc_15724_n5677) );
  INVX1 INVX1_904 ( .A(_abc_15724_n5680), .Y(_abc_15724_n5681) );
  INVX1 INVX1_905 ( .A(_abc_15724_n5685), .Y(_abc_15724_n5686) );
  INVX1 INVX1_906 ( .A(_abc_15724_n5688), .Y(_abc_15724_n5689) );
  INVX1 INVX1_907 ( .A(_abc_15724_n5694), .Y(_abc_15724_n5695) );
  INVX1 INVX1_908 ( .A(_abc_15724_n5697), .Y(_abc_15724_n5698) );
  INVX1 INVX1_909 ( .A(_abc_15724_n5707), .Y(_abc_15724_n5708) );
  INVX1 INVX1_91 ( .A(_abc_15724_n1220), .Y(_abc_15724_n1221) );
  INVX1 INVX1_910 ( .A(_abc_15724_n5709), .Y(_abc_15724_n5710) );
  INVX1 INVX1_911 ( .A(_abc_15724_n5711), .Y(_abc_15724_n5712) );
  INVX1 INVX1_912 ( .A(d_reg_26_), .Y(_abc_15724_n5713) );
  INVX1 INVX1_913 ( .A(_abc_15724_n5716), .Y(_abc_15724_n5717) );
  INVX1 INVX1_914 ( .A(_abc_15724_n5721), .Y(_abc_15724_n5722) );
  INVX1 INVX1_915 ( .A(_abc_15724_n5718), .Y(_abc_15724_n5726) );
  INVX1 INVX1_916 ( .A(_abc_15724_n5727), .Y(_abc_15724_n5728) );
  INVX1 INVX1_917 ( .A(_abc_15724_n5733), .Y(_abc_15724_n5734) );
  INVX1 INVX1_918 ( .A(_abc_15724_n5736), .Y(_abc_15724_n5737) );
  INVX1 INVX1_919 ( .A(_abc_15724_n5739), .Y(_abc_15724_n5740) );
  INVX1 INVX1_92 ( .A(_abc_15724_n1218_1), .Y(_abc_15724_n1224) );
  INVX1 INVX1_920 ( .A(_abc_15724_n5743), .Y(_abc_15724_n5744) );
  INVX1 INVX1_921 ( .A(_abc_15724_n5747), .Y(_abc_15724_n5748) );
  INVX1 INVX1_922 ( .A(_abc_15724_n5751), .Y(_abc_15724_n5752) );
  INVX1 INVX1_923 ( .A(_abc_15724_n5754), .Y(_abc_15724_n5755) );
  INVX1 INVX1_924 ( .A(_abc_15724_n5758), .Y(_abc_15724_n5759) );
  INVX1 INVX1_925 ( .A(_abc_15724_n5762), .Y(_abc_15724_n5763) );
  INVX1 INVX1_926 ( .A(_abc_15724_n5760), .Y(_abc_15724_n5772) );
  INVX1 INVX1_927 ( .A(_abc_15724_n5773), .Y(_abc_15724_n5774) );
  INVX1 INVX1_928 ( .A(_abc_15724_n5776), .Y(_abc_15724_n5777) );
  INVX1 INVX1_929 ( .A(_abc_15724_n5778), .Y(_abc_15724_n5779) );
  INVX1 INVX1_93 ( .A(_abc_15724_n1222), .Y(_abc_15724_n1225) );
  INVX1 INVX1_930 ( .A(d_reg_27_), .Y(_abc_15724_n5780) );
  INVX1 INVX1_931 ( .A(_abc_15724_n5783), .Y(_abc_15724_n5784) );
  INVX1 INVX1_932 ( .A(_abc_15724_n5788), .Y(_abc_15724_n5789) );
  INVX1 INVX1_933 ( .A(_abc_15724_n5785), .Y(_abc_15724_n5793) );
  INVX1 INVX1_934 ( .A(_abc_15724_n5794), .Y(_abc_15724_n5795) );
  INVX1 INVX1_935 ( .A(_abc_15724_n5800), .Y(_abc_15724_n5801) );
  INVX1 INVX1_936 ( .A(_abc_15724_n5803), .Y(_abc_15724_n5804) );
  INVX1 INVX1_937 ( .A(_abc_15724_n5806), .Y(_abc_15724_n5807) );
  INVX1 INVX1_938 ( .A(_abc_15724_n5810), .Y(_abc_15724_n5811) );
  INVX1 INVX1_939 ( .A(_abc_15724_n5814), .Y(_abc_15724_n5815) );
  INVX1 INVX1_94 ( .A(_abc_15724_n1245), .Y(_abc_15724_n1246) );
  INVX1 INVX1_940 ( .A(_abc_15724_n5819), .Y(_abc_15724_n5820) );
  INVX1 INVX1_941 ( .A(_abc_15724_n5822), .Y(_abc_15724_n5823) );
  INVX1 INVX1_942 ( .A(_abc_15724_n5825), .Y(_abc_15724_n5827) );
  INVX1 INVX1_943 ( .A(_abc_15724_n5837), .Y(_abc_15724_n5838) );
  INVX1 INVX1_944 ( .A(_abc_15724_n5706), .Y(_abc_15724_n5840) );
  INVX1 INVX1_945 ( .A(_abc_15724_n5841), .Y(_abc_15724_n5842) );
  INVX1 INVX1_946 ( .A(_abc_15724_n5846), .Y(_abc_15724_n5847) );
  INVX1 INVX1_947 ( .A(_abc_15724_n5848), .Y(_abc_15724_n5849) );
  INVX1 INVX1_948 ( .A(_abc_15724_n5850), .Y(_abc_15724_n5851) );
  INVX1 INVX1_949 ( .A(d_reg_28_), .Y(_abc_15724_n5852) );
  INVX1 INVX1_95 ( .A(_abc_15724_n1249), .Y(_abc_15724_n1250_1) );
  INVX1 INVX1_950 ( .A(_abc_15724_n5855), .Y(_abc_15724_n5856) );
  INVX1 INVX1_951 ( .A(_abc_15724_n5860), .Y(_abc_15724_n5861) );
  INVX1 INVX1_952 ( .A(_abc_15724_n5857), .Y(_abc_15724_n5865) );
  INVX1 INVX1_953 ( .A(_abc_15724_n5866), .Y(_abc_15724_n5867) );
  INVX1 INVX1_954 ( .A(_abc_15724_n5872), .Y(_abc_15724_n5873) );
  INVX1 INVX1_955 ( .A(_abc_15724_n5875), .Y(_abc_15724_n5876) );
  INVX1 INVX1_956 ( .A(_abc_15724_n5878), .Y(_abc_15724_n5879) );
  INVX1 INVX1_957 ( .A(_abc_15724_n5882), .Y(_abc_15724_n5883) );
  INVX1 INVX1_958 ( .A(_abc_15724_n5886), .Y(_abc_15724_n5887) );
  INVX1 INVX1_959 ( .A(_abc_15724_n5890), .Y(_abc_15724_n5891) );
  INVX1 INVX1_96 ( .A(_abc_15724_n1254), .Y(_abc_15724_n1255) );
  INVX1 INVX1_960 ( .A(_abc_15724_n5894), .Y(_abc_15724_n5895) );
  INVX1 INVX1_961 ( .A(_abc_15724_n5898), .Y(_abc_15724_n5899) );
  INVX1 INVX1_962 ( .A(_abc_15724_n5903), .Y(_abc_15724_n5904) );
  INVX1 INVX1_963 ( .A(_abc_15724_n5912), .Y(_abc_15724_n5913) );
  INVX1 INVX1_964 ( .A(_abc_15724_n5914), .Y(_abc_15724_n5915) );
  INVX1 INVX1_965 ( .A(_abc_15724_n5916), .Y(_abc_15724_n5917) );
  INVX1 INVX1_966 ( .A(d_reg_29_), .Y(_abc_15724_n5918) );
  INVX1 INVX1_967 ( .A(_abc_15724_n5921), .Y(_abc_15724_n5922) );
  INVX1 INVX1_968 ( .A(_abc_15724_n5926), .Y(_abc_15724_n5927) );
  INVX1 INVX1_969 ( .A(_abc_15724_n5923), .Y(_abc_15724_n5931) );
  INVX1 INVX1_97 ( .A(_abc_15724_n1257), .Y(_abc_15724_n1258) );
  INVX1 INVX1_970 ( .A(_abc_15724_n5932), .Y(_abc_15724_n5933) );
  INVX1 INVX1_971 ( .A(_abc_15724_n5938), .Y(_abc_15724_n5939) );
  INVX1 INVX1_972 ( .A(_abc_15724_n5941), .Y(_abc_15724_n5942) );
  INVX1 INVX1_973 ( .A(_abc_15724_n5944), .Y(_abc_15724_n5945) );
  INVX1 INVX1_974 ( .A(_abc_15724_n5948), .Y(_abc_15724_n5949) );
  INVX1 INVX1_975 ( .A(_abc_15724_n5952), .Y(_abc_15724_n5953) );
  INVX1 INVX1_976 ( .A(_abc_15724_n5956), .Y(_abc_15724_n5957) );
  INVX1 INVX1_977 ( .A(_abc_15724_n5960), .Y(_abc_15724_n5961) );
  INVX1 INVX1_978 ( .A(_abc_15724_n5964), .Y(_abc_15724_n5965) );
  INVX1 INVX1_979 ( .A(_abc_15724_n5970), .Y(_abc_15724_n5971) );
  INVX1 INVX1_98 ( .A(_abc_15724_n1259_1), .Y(_abc_15724_n1261_1) );
  INVX1 INVX1_980 ( .A(_abc_15724_n5973), .Y(_abc_15724_n5974) );
  INVX1 INVX1_981 ( .A(_abc_15724_n5983), .Y(_abc_15724_n5984) );
  INVX1 INVX1_982 ( .A(_abc_15724_n5985), .Y(_abc_15724_n5986) );
  INVX1 INVX1_983 ( .A(_abc_15724_n5987), .Y(_abc_15724_n5988) );
  INVX1 INVX1_984 ( .A(_abc_15724_n5989), .Y(_abc_15724_n5990) );
  INVX1 INVX1_985 ( .A(d_reg_30_), .Y(_abc_15724_n5991) );
  INVX1 INVX1_986 ( .A(_abc_15724_n5994), .Y(_abc_15724_n5995) );
  INVX1 INVX1_987 ( .A(_abc_15724_n5999), .Y(_abc_15724_n6000) );
  INVX1 INVX1_988 ( .A(_abc_15724_n5996), .Y(_abc_15724_n6004) );
  INVX1 INVX1_989 ( .A(_abc_15724_n6005), .Y(_abc_15724_n6006) );
  INVX1 INVX1_99 ( .A(_abc_15724_n1270), .Y(_abc_15724_n1271) );
  INVX1 INVX1_990 ( .A(_abc_15724_n6011), .Y(_abc_15724_n6012) );
  INVX1 INVX1_991 ( .A(_abc_15724_n6014), .Y(_abc_15724_n6015) );
  INVX1 INVX1_992 ( .A(_abc_15724_n6017), .Y(_abc_15724_n6018) );
  INVX1 INVX1_993 ( .A(_abc_15724_n6021), .Y(_abc_15724_n6022) );
  INVX1 INVX1_994 ( .A(_abc_15724_n6025), .Y(_abc_15724_n6026) );
  INVX1 INVX1_995 ( .A(_abc_15724_n6029), .Y(_abc_15724_n6030) );
  INVX1 INVX1_996 ( .A(_abc_15724_n6033), .Y(_abc_15724_n6034) );
  INVX1 INVX1_997 ( .A(_abc_15724_n6037), .Y(_abc_15724_n6038) );
  INVX1 INVX1_998 ( .A(_abc_15724_n6040), .Y(_abc_15724_n6042) );
  INVX1 INVX1_999 ( .A(_abc_15724_n6050), .Y(_abc_15724_n6051) );
  INVX2 INVX2_1 ( .A(_abc_15724_n4021), .Y(_abc_15724_n4022) );
  INVX8 INVX8_1 ( .A(digest_update_bF_buf10), .Y(_abc_15724_n850) );
  INVX8 INVX8_2 ( .A(_abc_15724_n851_bF_buf4), .Y(_abc_15724_n906) );
  INVX8 INVX8_3 ( .A(_abc_15724_n3721_bF_buf1), .Y(_abc_15724_n3805) );
  INVX8 INVX8_4 ( .A(w_mem_inst__abc_21378_n1586_bF_buf4), .Y(w_mem_inst__abc_21378_n1587) );
  INVX8 INVX8_5 ( .A(w_mem_inst__abc_21378_n3152_bF_buf62), .Y(w_mem_inst__abc_21378_n3154_1) );
  INVX8 INVX8_6 ( .A(round_ctr_rst_bF_buf59), .Y(w_mem_inst__abc_21378_n3156) );
  OR2X2 OR2X2_1 ( .A(e_reg_21_), .B(_auto_iopadmap_cc_313_execute_26059_21_), .Y(_abc_15724_n701) );
  OR2X2 OR2X2_10 ( .A(_auto_iopadmap_cc_313_execute_26059_14_), .B(e_reg_14_), .Y(_abc_15724_n735) );
  OR2X2 OR2X2_100 ( .A(_auto_iopadmap_cc_313_execute_26059_33_), .B(d_reg_1_), .Y(_abc_15724_n1014) );
  OR2X2 OR2X2_1000 ( .A(_abc_15724_n3711), .B(_abc_15724_n3708), .Y(_abc_15724_n3712) );
  OR2X2 OR2X2_1001 ( .A(_abc_15724_n3714), .B(_abc_15724_n3715), .Y(_abc_15724_n3716) );
  OR2X2 OR2X2_1002 ( .A(_abc_15724_n3717), .B(round_ctr_reg_6_), .Y(_abc_15724_n3718) );
  OR2X2 OR2X2_1003 ( .A(_abc_15724_n3719), .B(round_ctr_reg_5_), .Y(_abc_15724_n3720) );
  OR2X2 OR2X2_1004 ( .A(_abc_15724_n3718), .B(_abc_15724_n3720), .Y(_abc_15724_n3721) );
  OR2X2 OR2X2_1005 ( .A(_abc_15724_n3723), .B(round_ctr_reg_6_), .Y(_abc_15724_n3724) );
  OR2X2 OR2X2_1006 ( .A(_abc_15724_n3706), .B(_abc_15724_n3724), .Y(_abc_15724_n3725) );
  OR2X2 OR2X2_1007 ( .A(_abc_15724_n3730), .B(_abc_15724_n3729), .Y(_abc_15724_n3731) );
  OR2X2 OR2X2_1008 ( .A(_abc_15724_n3721_bF_buf3), .B(_abc_15724_n3731), .Y(_abc_15724_n3732) );
  OR2X2 OR2X2_1009 ( .A(_abc_15724_n3703), .B(round_ctr_reg_6_), .Y(_abc_15724_n3733) );
  OR2X2 OR2X2_101 ( .A(_abc_15724_n1016_1), .B(_abc_15724_n1001), .Y(_abc_15724_n1017) );
  OR2X2 OR2X2_1010 ( .A(_abc_15724_n3733), .B(_abc_15724_n3700), .Y(_abc_15724_n3734) );
  OR2X2 OR2X2_1011 ( .A(_abc_15724_n3708), .B(d_reg_0_), .Y(_abc_15724_n3739) );
  OR2X2 OR2X2_1012 ( .A(a_reg_27_), .B(e_reg_0_), .Y(_abc_15724_n3746) );
  OR2X2 OR2X2_1013 ( .A(_abc_15724_n3753), .B(_abc_15724_n3750), .Y(_abc_15724_n3754) );
  OR2X2 OR2X2_1014 ( .A(_abc_15724_n3756), .B(_abc_15724_n3757), .Y(_abc_15724_n3758) );
  OR2X2 OR2X2_1015 ( .A(_abc_15724_n3759), .B(_abc_15724_n3706), .Y(_abc_15724_n3760) );
  OR2X2 OR2X2_1016 ( .A(_abc_15724_n3765), .B(_abc_15724_n3766), .Y(_abc_15724_n3767) );
  OR2X2 OR2X2_1017 ( .A(_abc_15724_n3764), .B(_abc_15724_n3767), .Y(a_reg_0__FF_INPUT) );
  OR2X2 OR2X2_1018 ( .A(_abc_15724_n3744), .B(_abc_15724_n3754), .Y(_abc_15724_n3769) );
  OR2X2 OR2X2_1019 ( .A(_abc_15724_n3772), .B(_abc_15724_n3773), .Y(_abc_15724_n3774) );
  OR2X2 OR2X2_102 ( .A(_abc_15724_n1018_1), .B(_abc_15724_n850_bF_buf8), .Y(_abc_15724_n1019) );
  OR2X2 OR2X2_1020 ( .A(_abc_15724_n3774), .B(_abc_15724_n1009), .Y(_abc_15724_n3775) );
  OR2X2 OR2X2_1021 ( .A(_abc_15724_n3781), .B(_abc_15724_n3782), .Y(_abc_15724_n3783) );
  OR2X2 OR2X2_1022 ( .A(_abc_15724_n3783), .B(_abc_15724_n3721_bF_buf2), .Y(_abc_15724_n3784) );
  OR2X2 OR2X2_1023 ( .A(_abc_15724_n3781), .B(_abc_15724_n3772), .Y(_abc_15724_n3786) );
  OR2X2 OR2X2_1024 ( .A(_abc_15724_n3788), .B(_abc_15724_n3785), .Y(_abc_15724_n3789) );
  OR2X2 OR2X2_1025 ( .A(_abc_15724_n3789), .B(_abc_15724_n3779), .Y(_abc_15724_n3790) );
  OR2X2 OR2X2_1026 ( .A(_abc_15724_n3750), .B(_abc_15724_n3747), .Y(_abc_15724_n3791) );
  OR2X2 OR2X2_1027 ( .A(a_reg_28_), .B(e_reg_1_), .Y(_abc_15724_n3792) );
  OR2X2 OR2X2_1028 ( .A(_abc_15724_n3795), .B(w_1_), .Y(_abc_15724_n3798) );
  OR2X2 OR2X2_1029 ( .A(_abc_15724_n3799), .B(_abc_15724_n3791), .Y(_abc_15724_n3802) );
  OR2X2 OR2X2_103 ( .A(_abc_15724_n851_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_33_), .Y(_abc_15724_n1020) );
  OR2X2 OR2X2_1030 ( .A(_abc_15724_n3737_bF_buf2), .B(_abc_15724_n3805_bF_buf4), .Y(_abc_15724_n3806) );
  OR2X2 OR2X2_1031 ( .A(_abc_15724_n3808), .B(_abc_15724_n3776), .Y(_abc_15724_n3809) );
  OR2X2 OR2X2_1032 ( .A(_abc_15724_n3806_bF_buf3), .B(_abc_15724_n3809), .Y(_abc_15724_n3810) );
  OR2X2 OR2X2_1033 ( .A(_abc_15724_n3725_bF_buf2), .B(_abc_15724_n3786), .Y(_abc_15724_n3811) );
  OR2X2 OR2X2_1034 ( .A(_abc_15724_n3815), .B(_abc_15724_n3796), .Y(_abc_15724_n3816) );
  OR2X2 OR2X2_1035 ( .A(_abc_15724_n3817), .B(_abc_15724_n3800), .Y(_abc_15724_n3818) );
  OR2X2 OR2X2_1036 ( .A(_abc_15724_n3804), .B(_abc_15724_n3819), .Y(_abc_15724_n3820) );
  OR2X2 OR2X2_1037 ( .A(_abc_15724_n3820), .B(_abc_15724_n3769), .Y(_abc_15724_n3821) );
  OR2X2 OR2X2_1038 ( .A(_abc_15724_n3813), .B(_abc_15724_n3818), .Y(_abc_15724_n3822) );
  OR2X2 OR2X2_1039 ( .A(_abc_15724_n3790), .B(_abc_15724_n3803), .Y(_abc_15724_n3823) );
  OR2X2 OR2X2_104 ( .A(_abc_15724_n1020), .B(digest_update_bF_buf11), .Y(_abc_15724_n1021) );
  OR2X2 OR2X2_1040 ( .A(_abc_15724_n3824), .B(_abc_15724_n3756), .Y(_abc_15724_n3825) );
  OR2X2 OR2X2_1041 ( .A(_abc_15724_n3820), .B(_abc_15724_n3756), .Y(_abc_15724_n3828) );
  OR2X2 OR2X2_1042 ( .A(_abc_15724_n3824), .B(_abc_15724_n3769), .Y(_abc_15724_n3829) );
  OR2X2 OR2X2_1043 ( .A(_abc_15724_n3827), .B(_abc_15724_n3831), .Y(_abc_15724_n3832) );
  OR2X2 OR2X2_1044 ( .A(_abc_15724_n3832), .B(_abc_15724_n3762), .Y(_abc_15724_n3833) );
  OR2X2 OR2X2_1045 ( .A(_abc_15724_n3834), .B(_abc_15724_n3761), .Y(_abc_15724_n3835) );
  OR2X2 OR2X2_1046 ( .A(_abc_15724_n3838), .B(_abc_15724_n3840), .Y(_abc_15724_n3841) );
  OR2X2 OR2X2_1047 ( .A(_abc_15724_n3837), .B(_abc_15724_n3841), .Y(a_reg_1__FF_INPUT) );
  OR2X2 OR2X2_1048 ( .A(_abc_15724_n3830), .B(_abc_15724_n3736), .Y(_abc_15724_n3844) );
  OR2X2 OR2X2_1049 ( .A(_abc_15724_n3849), .B(_abc_15724_n3850), .Y(_abc_15724_n3851) );
  OR2X2 OR2X2_105 ( .A(_auto_iopadmap_cc_313_execute_26059_34_), .B(d_reg_2_), .Y(_abc_15724_n1024_1) );
  OR2X2 OR2X2_1050 ( .A(_abc_15724_n3853), .B(_abc_15724_n3855), .Y(_abc_15724_n3856) );
  OR2X2 OR2X2_1051 ( .A(_abc_15724_n3806_bF_buf2), .B(_abc_15724_n3856), .Y(_abc_15724_n3857) );
  OR2X2 OR2X2_1052 ( .A(_abc_15724_n3859), .B(_abc_15724_n3860), .Y(_abc_15724_n3861) );
  OR2X2 OR2X2_1053 ( .A(_abc_15724_n3861), .B(_abc_15724_n3721_bF_buf0), .Y(_abc_15724_n3862) );
  OR2X2 OR2X2_1054 ( .A(_abc_15724_n3859), .B(_abc_15724_n3849), .Y(_abc_15724_n3863) );
  OR2X2 OR2X2_1055 ( .A(_abc_15724_n3725_bF_buf1), .B(_abc_15724_n3863), .Y(_abc_15724_n3864) );
  OR2X2 OR2X2_1056 ( .A(_abc_15724_n3796), .B(_abc_15724_n3793), .Y(_abc_15724_n3867) );
  OR2X2 OR2X2_1057 ( .A(a_reg_29_), .B(e_reg_2_), .Y(_abc_15724_n3868) );
  OR2X2 OR2X2_1058 ( .A(_abc_15724_n3871), .B(w_2_), .Y(_abc_15724_n3874) );
  OR2X2 OR2X2_1059 ( .A(_abc_15724_n3878), .B(_abc_15724_n3872), .Y(_abc_15724_n3879) );
  OR2X2 OR2X2_106 ( .A(_abc_15724_n1023), .B(_abc_15724_n1028), .Y(_abc_15724_n1029) );
  OR2X2 OR2X2_1060 ( .A(_abc_15724_n3880), .B(_abc_15724_n3876), .Y(_abc_15724_n3881) );
  OR2X2 OR2X2_1061 ( .A(_abc_15724_n3851), .B(_abc_15724_n3854), .Y(_abc_15724_n3883) );
  OR2X2 OR2X2_1062 ( .A(_abc_15724_n3889), .B(_abc_15724_n3887), .Y(_abc_15724_n3890) );
  OR2X2 OR2X2_1063 ( .A(_abc_15724_n3890), .B(_abc_15724_n3886), .Y(_abc_15724_n3891) );
  OR2X2 OR2X2_1064 ( .A(_abc_15724_n3875), .B(_abc_15724_n3867), .Y(_abc_15724_n3893) );
  OR2X2 OR2X2_1065 ( .A(_abc_15724_n3895), .B(_abc_15724_n3882), .Y(_abc_15724_n3896) );
  OR2X2 OR2X2_1066 ( .A(_abc_15724_n3896), .B(_abc_15724_n3846), .Y(_abc_15724_n3897) );
  OR2X2 OR2X2_1067 ( .A(_abc_15724_n3804), .B(_abc_15724_n3800), .Y(_abc_15724_n3898) );
  OR2X2 OR2X2_1068 ( .A(_abc_15724_n3891), .B(_abc_15724_n3894), .Y(_abc_15724_n3899) );
  OR2X2 OR2X2_1069 ( .A(_abc_15724_n3866), .B(_abc_15724_n3881), .Y(_abc_15724_n3900) );
  OR2X2 OR2X2_107 ( .A(_abc_15724_n1030), .B(_abc_15724_n1011), .Y(_abc_15724_n1031) );
  OR2X2 OR2X2_1070 ( .A(_abc_15724_n3898), .B(_abc_15724_n3901), .Y(_abc_15724_n3902) );
  OR2X2 OR2X2_1071 ( .A(_abc_15724_n3903), .B(_abc_15724_n3734), .Y(_abc_15724_n3904) );
  OR2X2 OR2X2_1072 ( .A(_abc_15724_n3901), .B(_abc_15724_n3846), .Y(_abc_15724_n3905) );
  OR2X2 OR2X2_1073 ( .A(_abc_15724_n3896), .B(_abc_15724_n3898), .Y(_abc_15724_n3906) );
  OR2X2 OR2X2_1074 ( .A(_abc_15724_n3907), .B(_abc_15724_n3706), .Y(_abc_15724_n3908) );
  OR2X2 OR2X2_1075 ( .A(_abc_15724_n3909), .B(_abc_15724_n3845), .Y(_abc_15724_n3910) );
  OR2X2 OR2X2_1076 ( .A(_abc_15724_n3827), .B(_abc_15724_n3911), .Y(_abc_15724_n3912) );
  OR2X2 OR2X2_1077 ( .A(_abc_15724_n3913), .B(_abc_15724_n3914), .Y(_abc_15724_n3915) );
  OR2X2 OR2X2_1078 ( .A(_abc_15724_n3915), .B(_abc_15724_n3912), .Y(_abc_15724_n3916) );
  OR2X2 OR2X2_1079 ( .A(_abc_15724_n3918), .B(_abc_15724_n3843), .Y(_abc_15724_n3919) );
  OR2X2 OR2X2_108 ( .A(_abc_15724_n1031), .B(_abc_15724_n1027), .Y(_abc_15724_n1032) );
  OR2X2 OR2X2_1080 ( .A(_abc_15724_n3917), .B(_abc_15724_n3833), .Y(_abc_15724_n3920) );
  OR2X2 OR2X2_1081 ( .A(_abc_15724_n3923), .B(_abc_15724_n3925), .Y(_abc_15724_n3926) );
  OR2X2 OR2X2_1082 ( .A(_abc_15724_n3922), .B(_abc_15724_n3926), .Y(a_reg_2__FF_INPUT) );
  OR2X2 OR2X2_1083 ( .A(_abc_15724_n3914), .B(_abc_15724_n3930), .Y(_abc_15724_n3931) );
  OR2X2 OR2X2_1084 ( .A(_abc_15724_n3895), .B(_abc_15724_n3876), .Y(_abc_15724_n3932) );
  OR2X2 OR2X2_1085 ( .A(_abc_15724_n3936), .B(_abc_15724_n3937), .Y(_abc_15724_n3938) );
  OR2X2 OR2X2_1086 ( .A(_abc_15724_n3938), .B(_abc_15724_n3933), .Y(_abc_15724_n3941) );
  OR2X2 OR2X2_1087 ( .A(_abc_15724_n3945), .B(_abc_15724_n3946), .Y(_abc_15724_n3947) );
  OR2X2 OR2X2_1088 ( .A(_abc_15724_n3947), .B(_abc_15724_n3721_bF_buf4), .Y(_abc_15724_n3948) );
  OR2X2 OR2X2_1089 ( .A(_abc_15724_n3945), .B(_abc_15724_n3936), .Y(_abc_15724_n3950) );
  OR2X2 OR2X2_109 ( .A(_abc_15724_n1033), .B(_abc_15724_n850_bF_buf7), .Y(_abc_15724_n1034) );
  OR2X2 OR2X2_1090 ( .A(_abc_15724_n3952), .B(_abc_15724_n3949), .Y(_abc_15724_n3953) );
  OR2X2 OR2X2_1091 ( .A(_abc_15724_n3953), .B(_abc_15724_n3943), .Y(_abc_15724_n3954) );
  OR2X2 OR2X2_1092 ( .A(_abc_15724_n3872), .B(_abc_15724_n3869), .Y(_abc_15724_n3955) );
  OR2X2 OR2X2_1093 ( .A(a_reg_30_), .B(e_reg_3_), .Y(_abc_15724_n3956) );
  OR2X2 OR2X2_1094 ( .A(_abc_15724_n3959), .B(w_3_), .Y(_abc_15724_n3962) );
  OR2X2 OR2X2_1095 ( .A(_abc_15724_n3963), .B(_abc_15724_n3955), .Y(_abc_15724_n3966) );
  OR2X2 OR2X2_1096 ( .A(_abc_15724_n3954), .B(_abc_15724_n3967), .Y(_abc_15724_n3968) );
  OR2X2 OR2X2_1097 ( .A(_abc_15724_n3969), .B(_abc_15724_n3939), .Y(_abc_15724_n3970) );
  OR2X2 OR2X2_1098 ( .A(_abc_15724_n3806_bF_buf1), .B(_abc_15724_n3970), .Y(_abc_15724_n3971) );
  OR2X2 OR2X2_1099 ( .A(_abc_15724_n3725_bF_buf0), .B(_abc_15724_n3950), .Y(_abc_15724_n3972) );
  OR2X2 OR2X2_11 ( .A(_auto_iopadmap_cc_313_execute_26059_13_), .B(e_reg_13_), .Y(_abc_15724_n738_1) );
  OR2X2 OR2X2_110 ( .A(_abc_15724_n851_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_34_), .Y(_abc_15724_n1035) );
  OR2X2 OR2X2_1100 ( .A(_abc_15724_n3976), .B(_abc_15724_n3960), .Y(_abc_15724_n3977) );
  OR2X2 OR2X2_1101 ( .A(_abc_15724_n3978), .B(_abc_15724_n3964), .Y(_abc_15724_n3979) );
  OR2X2 OR2X2_1102 ( .A(_abc_15724_n3974), .B(_abc_15724_n3979), .Y(_abc_15724_n3980) );
  OR2X2 OR2X2_1103 ( .A(_abc_15724_n3985), .B(_abc_15724_n3984), .Y(_abc_15724_n3986) );
  OR2X2 OR2X2_1104 ( .A(_abc_15724_n3982), .B(_abc_15724_n3987), .Y(_abc_15724_n3988) );
  OR2X2 OR2X2_1105 ( .A(_abc_15724_n3988), .B(_abc_15724_n3726_bF_buf0), .Y(_abc_15724_n3989) );
  OR2X2 OR2X2_1106 ( .A(_abc_15724_n3986), .B(_abc_15724_n3983), .Y(_abc_15724_n3990) );
  OR2X2 OR2X2_1107 ( .A(_abc_15724_n3932), .B(_abc_15724_n3981), .Y(_abc_15724_n3991) );
  OR2X2 OR2X2_1108 ( .A(_abc_15724_n3992), .B(_abc_15724_n3806_bF_buf0), .Y(_abc_15724_n3993) );
  OR2X2 OR2X2_1109 ( .A(_abc_15724_n3998), .B(_abc_15724_n3997), .Y(_abc_15724_n3999) );
  OR2X2 OR2X2_111 ( .A(_abc_15724_n1035), .B(digest_update_bF_buf10), .Y(_abc_15724_n1036) );
  OR2X2 OR2X2_1110 ( .A(_abc_15724_n4000), .B(_abc_15724_n3995), .Y(_abc_15724_n4001) );
  OR2X2 OR2X2_1111 ( .A(_abc_15724_n4002), .B(_abc_15724_n3929), .Y(_abc_15724_n4003) );
  OR2X2 OR2X2_1112 ( .A(_abc_15724_n4003), .B(_abc_15724_n3928), .Y(_abc_15724_n4004) );
  OR2X2 OR2X2_1113 ( .A(_abc_15724_n3920), .B(_abc_15724_n4001), .Y(_abc_15724_n4005) );
  OR2X2 OR2X2_1114 ( .A(_abc_15724_n4001), .B(_abc_15724_n4006), .Y(_abc_15724_n4007) );
  OR2X2 OR2X2_1115 ( .A(_abc_15724_n4011), .B(_abc_15724_n4013), .Y(_abc_15724_n4014) );
  OR2X2 OR2X2_1116 ( .A(_abc_15724_n4010), .B(_abc_15724_n4014), .Y(a_reg_3__FF_INPUT) );
  OR2X2 OR2X2_1117 ( .A(_abc_15724_n4027), .B(_abc_15724_n4028), .Y(_abc_15724_n4029) );
  OR2X2 OR2X2_1118 ( .A(_abc_15724_n4029), .B(_abc_15724_n4024), .Y(_abc_15724_n4031) );
  OR2X2 OR2X2_1119 ( .A(_abc_15724_n4032), .B(_abc_15724_n4030), .Y(_abc_15724_n4033) );
  OR2X2 OR2X2_112 ( .A(_auto_iopadmap_cc_313_execute_26059_35_), .B(d_reg_3_), .Y(_abc_15724_n1039_1) );
  OR2X2 OR2X2_1120 ( .A(_abc_15724_n3806_bF_buf2), .B(_abc_15724_n4033), .Y(_abc_15724_n4034) );
  OR2X2 OR2X2_1121 ( .A(_abc_15724_n4036), .B(_abc_15724_n4037), .Y(_abc_15724_n4038) );
  OR2X2 OR2X2_1122 ( .A(_abc_15724_n4038), .B(_abc_15724_n3721_bF_buf2), .Y(_abc_15724_n4039) );
  OR2X2 OR2X2_1123 ( .A(_abc_15724_n4036), .B(_abc_15724_n4027), .Y(_abc_15724_n4040) );
  OR2X2 OR2X2_1124 ( .A(_abc_15724_n3725_bF_buf3), .B(_abc_15724_n4040), .Y(_abc_15724_n4041) );
  OR2X2 OR2X2_1125 ( .A(_abc_15724_n3960), .B(_abc_15724_n3957), .Y(_abc_15724_n4044) );
  OR2X2 OR2X2_1126 ( .A(a_reg_31_), .B(e_reg_4_), .Y(_abc_15724_n4045) );
  OR2X2 OR2X2_1127 ( .A(_abc_15724_n4048), .B(w_4_), .Y(_abc_15724_n4051) );
  OR2X2 OR2X2_1128 ( .A(_abc_15724_n4055), .B(_abc_15724_n4049), .Y(_abc_15724_n4056) );
  OR2X2 OR2X2_1129 ( .A(_abc_15724_n4057), .B(_abc_15724_n4053), .Y(_abc_15724_n4058) );
  OR2X2 OR2X2_113 ( .A(_abc_15724_n1038_1), .B(_abc_15724_n1043), .Y(_abc_15724_n1044) );
  OR2X2 OR2X2_1130 ( .A(_abc_15724_n4065), .B(_abc_15724_n4063), .Y(_abc_15724_n4066) );
  OR2X2 OR2X2_1131 ( .A(_abc_15724_n4066), .B(_abc_15724_n4062), .Y(_abc_15724_n4067) );
  OR2X2 OR2X2_1132 ( .A(_abc_15724_n4052), .B(_abc_15724_n4044), .Y(_abc_15724_n4069) );
  OR2X2 OR2X2_1133 ( .A(_abc_15724_n4071), .B(_abc_15724_n4059), .Y(_abc_15724_n4072) );
  OR2X2 OR2X2_1134 ( .A(_abc_15724_n4072), .B(_abc_15724_n4023), .Y(_abc_15724_n4073) );
  OR2X2 OR2X2_1135 ( .A(_abc_15724_n3985), .B(_abc_15724_n3964), .Y(_abc_15724_n4074) );
  OR2X2 OR2X2_1136 ( .A(_abc_15724_n4067), .B(_abc_15724_n4070), .Y(_abc_15724_n4075) );
  OR2X2 OR2X2_1137 ( .A(_abc_15724_n4043), .B(_abc_15724_n4058), .Y(_abc_15724_n4076) );
  OR2X2 OR2X2_1138 ( .A(_abc_15724_n4074), .B(_abc_15724_n4077), .Y(_abc_15724_n4078) );
  OR2X2 OR2X2_1139 ( .A(_abc_15724_n4081), .B(_abc_15724_n4082), .Y(_abc_15724_n4083) );
  OR2X2 OR2X2_114 ( .A(_abc_15724_n1045), .B(_abc_15724_n1025_1), .Y(_abc_15724_n1046) );
  OR2X2 OR2X2_1140 ( .A(_abc_15724_n4084), .B(_abc_15724_n4080), .Y(_abc_15724_n4085) );
  OR2X2 OR2X2_1141 ( .A(_abc_15724_n4085), .B(_abc_15724_n4020), .Y(_abc_15724_n4086) );
  OR2X2 OR2X2_1142 ( .A(_abc_15724_n4087), .B(_abc_15724_n4088), .Y(_abc_15724_n4089) );
  OR2X2 OR2X2_1143 ( .A(_abc_15724_n4019), .B(_abc_15724_n4090), .Y(_abc_15724_n4091) );
  OR2X2 OR2X2_1144 ( .A(_abc_15724_n4096), .B(_abc_15724_n4098), .Y(_abc_15724_n4099) );
  OR2X2 OR2X2_1145 ( .A(_abc_15724_n4095), .B(_abc_15724_n4099), .Y(a_reg_4__FF_INPUT) );
  OR2X2 OR2X2_1146 ( .A(_abc_15724_n4080), .B(_abc_15724_n4081), .Y(_abc_15724_n4101) );
  OR2X2 OR2X2_1147 ( .A(_abc_15724_n4106), .B(_abc_15724_n4107), .Y(_abc_15724_n4108) );
  OR2X2 OR2X2_1148 ( .A(_abc_15724_n4108), .B(_abc_15724_n4103), .Y(_abc_15724_n4110) );
  OR2X2 OR2X2_1149 ( .A(_abc_15724_n4111), .B(_abc_15724_n4109), .Y(_abc_15724_n4112) );
  OR2X2 OR2X2_115 ( .A(_abc_15724_n1046), .B(_abc_15724_n1042), .Y(_abc_15724_n1047_1) );
  OR2X2 OR2X2_1150 ( .A(_abc_15724_n3806_bF_buf1), .B(_abc_15724_n4112), .Y(_abc_15724_n4113) );
  OR2X2 OR2X2_1151 ( .A(_abc_15724_n4115), .B(_abc_15724_n4116), .Y(_abc_15724_n4117) );
  OR2X2 OR2X2_1152 ( .A(_abc_15724_n4117), .B(_abc_15724_n3721_bF_buf1), .Y(_abc_15724_n4118) );
  OR2X2 OR2X2_1153 ( .A(_abc_15724_n4115), .B(_abc_15724_n4106), .Y(_abc_15724_n4119) );
  OR2X2 OR2X2_1154 ( .A(_abc_15724_n3725_bF_buf2), .B(_abc_15724_n4119), .Y(_abc_15724_n4120) );
  OR2X2 OR2X2_1155 ( .A(_abc_15724_n4049), .B(_abc_15724_n4046), .Y(_abc_15724_n4123) );
  OR2X2 OR2X2_1156 ( .A(a_reg_0_), .B(e_reg_5_), .Y(_abc_15724_n4124) );
  OR2X2 OR2X2_1157 ( .A(_abc_15724_n4127), .B(w_5_), .Y(_abc_15724_n4130) );
  OR2X2 OR2X2_1158 ( .A(_abc_15724_n4134), .B(_abc_15724_n4128), .Y(_abc_15724_n4135) );
  OR2X2 OR2X2_1159 ( .A(_abc_15724_n4136), .B(_abc_15724_n4132), .Y(_abc_15724_n4137) );
  OR2X2 OR2X2_116 ( .A(_abc_15724_n1049), .B(_abc_15724_n1050_1), .Y(H3_reg_3__FF_INPUT) );
  OR2X2 OR2X2_1160 ( .A(_abc_15724_n4144), .B(_abc_15724_n4142), .Y(_abc_15724_n4145) );
  OR2X2 OR2X2_1161 ( .A(_abc_15724_n4145), .B(_abc_15724_n4141), .Y(_abc_15724_n4146) );
  OR2X2 OR2X2_1162 ( .A(_abc_15724_n4131), .B(_abc_15724_n4123), .Y(_abc_15724_n4148) );
  OR2X2 OR2X2_1163 ( .A(_abc_15724_n4150), .B(_abc_15724_n4138), .Y(_abc_15724_n4151) );
  OR2X2 OR2X2_1164 ( .A(_abc_15724_n4151), .B(_abc_15724_n4102), .Y(_abc_15724_n4152) );
  OR2X2 OR2X2_1165 ( .A(_abc_15724_n4071), .B(_abc_15724_n4053), .Y(_abc_15724_n4153) );
  OR2X2 OR2X2_1166 ( .A(_abc_15724_n4146), .B(_abc_15724_n4149), .Y(_abc_15724_n4154) );
  OR2X2 OR2X2_1167 ( .A(_abc_15724_n4122), .B(_abc_15724_n4137), .Y(_abc_15724_n4155) );
  OR2X2 OR2X2_1168 ( .A(_abc_15724_n4153), .B(_abc_15724_n4156), .Y(_abc_15724_n4157) );
  OR2X2 OR2X2_1169 ( .A(_abc_15724_n4158), .B(_abc_15724_n4021), .Y(_abc_15724_n4159) );
  OR2X2 OR2X2_117 ( .A(_auto_iopadmap_cc_313_execute_26059_36_), .B(d_reg_4_), .Y(_abc_15724_n1052) );
  OR2X2 OR2X2_1170 ( .A(_abc_15724_n4160), .B(_abc_15724_n4161), .Y(_abc_15724_n4162) );
  OR2X2 OR2X2_1171 ( .A(_abc_15724_n4162), .B(_abc_15724_n4022), .Y(_abc_15724_n4163) );
  OR2X2 OR2X2_1172 ( .A(_abc_15724_n4083), .B(_abc_15724_n4021), .Y(_abc_15724_n4166) );
  OR2X2 OR2X2_1173 ( .A(_abc_15724_n4168), .B(_abc_15724_n4169), .Y(_abc_15724_n4170) );
  OR2X2 OR2X2_1174 ( .A(_abc_15724_n4171), .B(_abc_15724_n4165), .Y(_abc_15724_n4172) );
  OR2X2 OR2X2_1175 ( .A(_abc_15724_n4173), .B(_abc_15724_n4087), .Y(_abc_15724_n4174) );
  OR2X2 OR2X2_1176 ( .A(_abc_15724_n4092), .B(_abc_15724_n4174), .Y(_abc_15724_n4175) );
  OR2X2 OR2X2_1177 ( .A(_abc_15724_n4089), .B(_abc_15724_n4172), .Y(_abc_15724_n4176) );
  OR2X2 OR2X2_1178 ( .A(_abc_15724_n4172), .B(_abc_15724_n4086), .Y(_abc_15724_n4180) );
  OR2X2 OR2X2_1179 ( .A(_abc_15724_n4184), .B(_abc_15724_n4186), .Y(_abc_15724_n4187) );
  OR2X2 OR2X2_118 ( .A(_abc_15724_n1038_1), .B(_abc_15724_n1057), .Y(_abc_15724_n1058) );
  OR2X2 OR2X2_1180 ( .A(_abc_15724_n4183), .B(_abc_15724_n4187), .Y(a_reg_5__FF_INPUT) );
  OR2X2 OR2X2_1181 ( .A(_abc_15724_n4199), .B(_abc_15724_n4200), .Y(_abc_15724_n4201) );
  OR2X2 OR2X2_1182 ( .A(_abc_15724_n4201), .B(_abc_15724_n4196), .Y(_abc_15724_n4204) );
  OR2X2 OR2X2_1183 ( .A(_abc_15724_n4207), .B(_abc_15724_n4208), .Y(_abc_15724_n4209) );
  OR2X2 OR2X2_1184 ( .A(_abc_15724_n3721_bF_buf0), .B(_abc_15724_n4209), .Y(_abc_15724_n4210) );
  OR2X2 OR2X2_1185 ( .A(_abc_15724_n4213), .B(_abc_15724_n4199), .Y(_abc_15724_n4214) );
  OR2X2 OR2X2_1186 ( .A(_abc_15724_n4216), .B(_abc_15724_n4211), .Y(_abc_15724_n4217) );
  OR2X2 OR2X2_1187 ( .A(_abc_15724_n4217), .B(_abc_15724_n4206), .Y(_abc_15724_n4218) );
  OR2X2 OR2X2_1188 ( .A(a_reg_1_), .B(e_reg_6_), .Y(_abc_15724_n4222) );
  OR2X2 OR2X2_1189 ( .A(_abc_15724_n4225), .B(w_6_), .Y(_abc_15724_n4228) );
  OR2X2 OR2X2_119 ( .A(_abc_15724_n1059), .B(_abc_15724_n1056), .Y(_abc_15724_n1060_1) );
  OR2X2 OR2X2_1190 ( .A(_abc_15724_n4232), .B(_abc_15724_n4230), .Y(_abc_15724_n4233) );
  OR2X2 OR2X2_1191 ( .A(_abc_15724_n4234), .B(_abc_15724_n4238), .Y(_abc_15724_n4239) );
  OR2X2 OR2X2_1192 ( .A(_abc_15724_n4239), .B(_abc_15724_n4195), .Y(_abc_15724_n4240) );
  OR2X2 OR2X2_1193 ( .A(_abc_15724_n4237), .B(_abc_15724_n4218), .Y(_abc_15724_n4242) );
  OR2X2 OR2X2_1194 ( .A(_abc_15724_n4219), .B(_abc_15724_n4233), .Y(_abc_15724_n4243) );
  OR2X2 OR2X2_1195 ( .A(_abc_15724_n4244), .B(_abc_15724_n4241), .Y(_abc_15724_n4245) );
  OR2X2 OR2X2_1196 ( .A(_abc_15724_n4246), .B(_abc_15724_n3734), .Y(_abc_15724_n4247) );
  OR2X2 OR2X2_1197 ( .A(_abc_15724_n4248), .B(_abc_15724_n4249), .Y(_abc_15724_n4250) );
  OR2X2 OR2X2_1198 ( .A(_abc_15724_n4250), .B(_abc_15724_n3706), .Y(_abc_15724_n4251) );
  OR2X2 OR2X2_1199 ( .A(_abc_15724_n4254), .B(_abc_15724_n4255), .Y(_abc_15724_n4256) );
  OR2X2 OR2X2_12 ( .A(_abc_15724_n747), .B(_abc_15724_n729_1), .Y(_abc_15724_n748) );
  OR2X2 OR2X2_120 ( .A(_abc_15724_n1061_1), .B(_abc_15724_n1040), .Y(_abc_15724_n1062) );
  OR2X2 OR2X2_1200 ( .A(_abc_15724_n4257), .B(_abc_15724_n4253), .Y(_abc_15724_n4258) );
  OR2X2 OR2X2_1201 ( .A(_abc_15724_n4192), .B(_abc_15724_n4259), .Y(_abc_15724_n4262) );
  OR2X2 OR2X2_1202 ( .A(_abc_15724_n4265), .B(_abc_15724_n4267), .Y(_abc_15724_n4268) );
  OR2X2 OR2X2_1203 ( .A(_abc_15724_n4264), .B(_abc_15724_n4268), .Y(a_reg_6__FF_INPUT) );
  OR2X2 OR2X2_1204 ( .A(_abc_15724_n4255), .B(_abc_15724_n4248), .Y(_abc_15724_n4273) );
  OR2X2 OR2X2_1205 ( .A(_abc_15724_n4279), .B(_abc_15724_n4280), .Y(_abc_15724_n4281) );
  OR2X2 OR2X2_1206 ( .A(_abc_15724_n4281), .B(_abc_15724_n4276), .Y(_abc_15724_n4283) );
  OR2X2 OR2X2_1207 ( .A(_abc_15724_n4284), .B(_abc_15724_n4282), .Y(_abc_15724_n4285) );
  OR2X2 OR2X2_1208 ( .A(_abc_15724_n3806_bF_buf0), .B(_abc_15724_n4285), .Y(_abc_15724_n4286) );
  OR2X2 OR2X2_1209 ( .A(_abc_15724_n4288), .B(_abc_15724_n4289), .Y(_abc_15724_n4290) );
  OR2X2 OR2X2_121 ( .A(_abc_15724_n1062), .B(_abc_15724_n1055), .Y(_abc_15724_n1063_1) );
  OR2X2 OR2X2_1210 ( .A(_abc_15724_n4290), .B(_abc_15724_n3721_bF_buf4), .Y(_abc_15724_n4291) );
  OR2X2 OR2X2_1211 ( .A(_abc_15724_n4288), .B(_abc_15724_n4279), .Y(_abc_15724_n4292) );
  OR2X2 OR2X2_1212 ( .A(_abc_15724_n3725_bF_buf1), .B(_abc_15724_n4292), .Y(_abc_15724_n4293) );
  OR2X2 OR2X2_1213 ( .A(_abc_15724_n4226), .B(_abc_15724_n4223), .Y(_abc_15724_n4296) );
  OR2X2 OR2X2_1214 ( .A(a_reg_2_), .B(e_reg_7_), .Y(_abc_15724_n4297) );
  OR2X2 OR2X2_1215 ( .A(_abc_15724_n4300), .B(w_7_), .Y(_abc_15724_n4303) );
  OR2X2 OR2X2_1216 ( .A(_abc_15724_n4307), .B(_abc_15724_n4301), .Y(_abc_15724_n4308) );
  OR2X2 OR2X2_1217 ( .A(_abc_15724_n4309), .B(_abc_15724_n4305), .Y(_abc_15724_n4310) );
  OR2X2 OR2X2_1218 ( .A(_abc_15724_n4317), .B(_abc_15724_n4315), .Y(_abc_15724_n4318) );
  OR2X2 OR2X2_1219 ( .A(_abc_15724_n4318), .B(_abc_15724_n4314), .Y(_abc_15724_n4319) );
  OR2X2 OR2X2_122 ( .A(_abc_15724_n1064), .B(_abc_15724_n850_bF_buf6), .Y(_abc_15724_n1065) );
  OR2X2 OR2X2_1220 ( .A(_abc_15724_n4304), .B(_abc_15724_n4296), .Y(_abc_15724_n4321) );
  OR2X2 OR2X2_1221 ( .A(_abc_15724_n4323), .B(_abc_15724_n4311), .Y(_abc_15724_n4324) );
  OR2X2 OR2X2_1222 ( .A(_abc_15724_n4326), .B(_abc_15724_n4327), .Y(_abc_15724_n4328) );
  OR2X2 OR2X2_1223 ( .A(_abc_15724_n4332), .B(_abc_15724_n4329), .Y(_abc_15724_n4333) );
  OR2X2 OR2X2_1224 ( .A(_abc_15724_n4272), .B(_abc_15724_n4334), .Y(_abc_15724_n4335) );
  OR2X2 OR2X2_1225 ( .A(_abc_15724_n4271), .B(_abc_15724_n4333), .Y(_abc_15724_n4336) );
  OR2X2 OR2X2_1226 ( .A(_abc_15724_n4339), .B(_abc_15724_n4341), .Y(_abc_15724_n4342) );
  OR2X2 OR2X2_1227 ( .A(_abc_15724_n4338), .B(_abc_15724_n4342), .Y(a_reg_7__FF_INPUT) );
  OR2X2 OR2X2_1228 ( .A(_abc_15724_n4258), .B(_abc_15724_n4333), .Y(_abc_15724_n4344) );
  OR2X2 OR2X2_1229 ( .A(_abc_15724_n4176), .B(_abc_15724_n4344), .Y(_abc_15724_n4345) );
  OR2X2 OR2X2_123 ( .A(_abc_15724_n851_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_36_), .Y(_abc_15724_n1066) );
  OR2X2 OR2X2_1230 ( .A(_abc_15724_n4018), .B(_abc_15724_n4345), .Y(_abc_15724_n4346) );
  OR2X2 OR2X2_1231 ( .A(_abc_15724_n4190), .B(_abc_15724_n4344), .Y(_abc_15724_n4347) );
  OR2X2 OR2X2_1232 ( .A(_abc_15724_n4349), .B(_abc_15724_n4332), .Y(_abc_15724_n4350) );
  OR2X2 OR2X2_1233 ( .A(_abc_15724_n4295), .B(_abc_15724_n4310), .Y(_abc_15724_n4354) );
  OR2X2 OR2X2_1234 ( .A(_abc_15724_n4359), .B(_abc_15724_n4360), .Y(_abc_15724_n4361) );
  OR2X2 OR2X2_1235 ( .A(_abc_15724_n4361), .B(_abc_15724_n4356), .Y(_abc_15724_n4363) );
  OR2X2 OR2X2_1236 ( .A(_abc_15724_n4364), .B(_abc_15724_n4362), .Y(_abc_15724_n4365) );
  OR2X2 OR2X2_1237 ( .A(_abc_15724_n3806_bF_buf3), .B(_abc_15724_n4365), .Y(_abc_15724_n4366) );
  OR2X2 OR2X2_1238 ( .A(_abc_15724_n4368), .B(_abc_15724_n4369), .Y(_abc_15724_n4370) );
  OR2X2 OR2X2_1239 ( .A(_abc_15724_n4370), .B(_abc_15724_n3721_bF_buf3), .Y(_abc_15724_n4371) );
  OR2X2 OR2X2_124 ( .A(_abc_15724_n1066), .B(digest_update_bF_buf8), .Y(_abc_15724_n1067) );
  OR2X2 OR2X2_1240 ( .A(_abc_15724_n4368), .B(_abc_15724_n4359), .Y(_abc_15724_n4372) );
  OR2X2 OR2X2_1241 ( .A(_abc_15724_n3725_bF_buf0), .B(_abc_15724_n4372), .Y(_abc_15724_n4373) );
  OR2X2 OR2X2_1242 ( .A(_abc_15724_n4301), .B(_abc_15724_n4298), .Y(_abc_15724_n4376) );
  OR2X2 OR2X2_1243 ( .A(a_reg_3_), .B(e_reg_8_), .Y(_abc_15724_n4377) );
  OR2X2 OR2X2_1244 ( .A(_abc_15724_n4380), .B(w_8_), .Y(_abc_15724_n4383) );
  OR2X2 OR2X2_1245 ( .A(_abc_15724_n4387), .B(_abc_15724_n4381), .Y(_abc_15724_n4388) );
  OR2X2 OR2X2_1246 ( .A(_abc_15724_n4389), .B(_abc_15724_n4385), .Y(_abc_15724_n4390) );
  OR2X2 OR2X2_1247 ( .A(_abc_15724_n4397), .B(_abc_15724_n4395), .Y(_abc_15724_n4398) );
  OR2X2 OR2X2_1248 ( .A(_abc_15724_n4398), .B(_abc_15724_n4394), .Y(_abc_15724_n4399) );
  OR2X2 OR2X2_1249 ( .A(_abc_15724_n4384), .B(_abc_15724_n4376), .Y(_abc_15724_n4401) );
  OR2X2 OR2X2_125 ( .A(_abc_15724_n1069_1), .B(_abc_15724_n1053), .Y(_abc_15724_n1070_1) );
  OR2X2 OR2X2_1250 ( .A(_abc_15724_n4403), .B(_abc_15724_n4391), .Y(_abc_15724_n4404) );
  OR2X2 OR2X2_1251 ( .A(_abc_15724_n4404), .B(_abc_15724_n4355), .Y(_abc_15724_n4405) );
  OR2X2 OR2X2_1252 ( .A(_abc_15724_n4323), .B(_abc_15724_n4305), .Y(_abc_15724_n4406) );
  OR2X2 OR2X2_1253 ( .A(_abc_15724_n4399), .B(_abc_15724_n4402), .Y(_abc_15724_n4407) );
  OR2X2 OR2X2_1254 ( .A(_abc_15724_n4375), .B(_abc_15724_n4390), .Y(_abc_15724_n4408) );
  OR2X2 OR2X2_1255 ( .A(_abc_15724_n4406), .B(_abc_15724_n4409), .Y(_abc_15724_n4410) );
  OR2X2 OR2X2_1256 ( .A(_abc_15724_n4413), .B(_abc_15724_n4414), .Y(_abc_15724_n4415) );
  OR2X2 OR2X2_1257 ( .A(_abc_15724_n4416), .B(_abc_15724_n4412), .Y(_abc_15724_n4417) );
  OR2X2 OR2X2_1258 ( .A(_abc_15724_n4417), .B(_abc_15724_n4327), .Y(_abc_15724_n4418) );
  OR2X2 OR2X2_1259 ( .A(_abc_15724_n4419), .B(_abc_15724_n4420), .Y(_abc_15724_n4421) );
  OR2X2 OR2X2_126 ( .A(_auto_iopadmap_cc_313_execute_26059_37_), .B(d_reg_5_), .Y(_abc_15724_n1071_1) );
  OR2X2 OR2X2_1260 ( .A(_abc_15724_n4353), .B(_abc_15724_n4422), .Y(_abc_15724_n4425) );
  OR2X2 OR2X2_1261 ( .A(_abc_15724_n4428), .B(_abc_15724_n4429), .Y(_abc_15724_n4430) );
  OR2X2 OR2X2_1262 ( .A(_abc_15724_n4427), .B(_abc_15724_n4430), .Y(a_reg_8__FF_INPUT) );
  OR2X2 OR2X2_1263 ( .A(_abc_15724_n4412), .B(_abc_15724_n4413), .Y(_abc_15724_n4432) );
  OR2X2 OR2X2_1264 ( .A(_abc_15724_n4437), .B(_abc_15724_n4438), .Y(_abc_15724_n4439) );
  OR2X2 OR2X2_1265 ( .A(_abc_15724_n4439), .B(_abc_15724_n4434), .Y(_abc_15724_n4441) );
  OR2X2 OR2X2_1266 ( .A(_abc_15724_n4442), .B(_abc_15724_n4440), .Y(_abc_15724_n4443) );
  OR2X2 OR2X2_1267 ( .A(_abc_15724_n3806_bF_buf2), .B(_abc_15724_n4443), .Y(_abc_15724_n4444) );
  OR2X2 OR2X2_1268 ( .A(_abc_15724_n4446), .B(_abc_15724_n4447), .Y(_abc_15724_n4448) );
  OR2X2 OR2X2_1269 ( .A(_abc_15724_n4448), .B(_abc_15724_n3721_bF_buf2), .Y(_abc_15724_n4449) );
  OR2X2 OR2X2_127 ( .A(_abc_15724_n1070_1), .B(_abc_15724_n1074), .Y(_abc_15724_n1075) );
  OR2X2 OR2X2_1270 ( .A(_abc_15724_n4446), .B(_abc_15724_n4437), .Y(_abc_15724_n4450) );
  OR2X2 OR2X2_1271 ( .A(_abc_15724_n3725_bF_buf2), .B(_abc_15724_n4450), .Y(_abc_15724_n4451) );
  OR2X2 OR2X2_1272 ( .A(_abc_15724_n4381), .B(_abc_15724_n4378), .Y(_abc_15724_n4454) );
  OR2X2 OR2X2_1273 ( .A(a_reg_4_), .B(e_reg_9_), .Y(_abc_15724_n4455) );
  OR2X2 OR2X2_1274 ( .A(_abc_15724_n4458), .B(w_9_), .Y(_abc_15724_n4461) );
  OR2X2 OR2X2_1275 ( .A(_abc_15724_n4465), .B(_abc_15724_n4459), .Y(_abc_15724_n4466) );
  OR2X2 OR2X2_1276 ( .A(_abc_15724_n4467), .B(_abc_15724_n4463), .Y(_abc_15724_n4468) );
  OR2X2 OR2X2_1277 ( .A(_abc_15724_n4475), .B(_abc_15724_n4473), .Y(_abc_15724_n4476) );
  OR2X2 OR2X2_1278 ( .A(_abc_15724_n4476), .B(_abc_15724_n4472), .Y(_abc_15724_n4477) );
  OR2X2 OR2X2_1279 ( .A(_abc_15724_n4462), .B(_abc_15724_n4454), .Y(_abc_15724_n4479) );
  OR2X2 OR2X2_128 ( .A(_abc_15724_n1076), .B(_abc_15724_n1077), .Y(_abc_15724_n1078) );
  OR2X2 OR2X2_1280 ( .A(_abc_15724_n4481), .B(_abc_15724_n4469), .Y(_abc_15724_n4482) );
  OR2X2 OR2X2_1281 ( .A(_abc_15724_n4482), .B(_abc_15724_n4433), .Y(_abc_15724_n4483) );
  OR2X2 OR2X2_1282 ( .A(_abc_15724_n4403), .B(_abc_15724_n4385), .Y(_abc_15724_n4484) );
  OR2X2 OR2X2_1283 ( .A(_abc_15724_n4477), .B(_abc_15724_n4480), .Y(_abc_15724_n4485) );
  OR2X2 OR2X2_1284 ( .A(_abc_15724_n4453), .B(_abc_15724_n4468), .Y(_abc_15724_n4486) );
  OR2X2 OR2X2_1285 ( .A(_abc_15724_n4484), .B(_abc_15724_n4487), .Y(_abc_15724_n4488) );
  OR2X2 OR2X2_1286 ( .A(_abc_15724_n4489), .B(_abc_15724_n4021), .Y(_abc_15724_n4490) );
  OR2X2 OR2X2_1287 ( .A(_abc_15724_n4491), .B(_abc_15724_n4492), .Y(_abc_15724_n4493) );
  OR2X2 OR2X2_1288 ( .A(_abc_15724_n4493), .B(_abc_15724_n4022), .Y(_abc_15724_n4494) );
  OR2X2 OR2X2_1289 ( .A(_abc_15724_n4415), .B(_abc_15724_n3737_bF_buf2), .Y(_abc_15724_n4497) );
  OR2X2 OR2X2_129 ( .A(_abc_15724_n851_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_37_), .Y(_abc_15724_n1081) );
  OR2X2 OR2X2_1290 ( .A(_abc_15724_n4499), .B(_abc_15724_n4500), .Y(_abc_15724_n4501) );
  OR2X2 OR2X2_1291 ( .A(_abc_15724_n4502), .B(_abc_15724_n4496), .Y(_abc_15724_n4503) );
  OR2X2 OR2X2_1292 ( .A(_abc_15724_n4504), .B(_abc_15724_n4419), .Y(_abc_15724_n4507) );
  OR2X2 OR2X2_1293 ( .A(_abc_15724_n4423), .B(_abc_15724_n4507), .Y(_abc_15724_n4508) );
  OR2X2 OR2X2_1294 ( .A(_abc_15724_n4503), .B(_abc_15724_n4418), .Y(_abc_15724_n4509) );
  OR2X2 OR2X2_1295 ( .A(_abc_15724_n4513), .B(_abc_15724_n4514), .Y(_abc_15724_n4515) );
  OR2X2 OR2X2_1296 ( .A(_abc_15724_n4512), .B(_abc_15724_n4515), .Y(a_reg_9__FF_INPUT) );
  OR2X2 OR2X2_1297 ( .A(_abc_15724_n4505), .B(_abc_15724_n4519), .Y(_abc_15724_n4520) );
  OR2X2 OR2X2_1298 ( .A(_abc_15724_n4527), .B(_abc_15724_n4528), .Y(_abc_15724_n4529) );
  OR2X2 OR2X2_1299 ( .A(_abc_15724_n4529), .B(_abc_15724_n4524), .Y(_abc_15724_n4532) );
  OR2X2 OR2X2_13 ( .A(_abc_15724_n746), .B(_abc_15724_n748), .Y(_abc_15724_n749) );
  OR2X2 OR2X2_130 ( .A(_abc_15724_n1080), .B(_abc_15724_n1082_1), .Y(H3_reg_5__FF_INPUT) );
  OR2X2 OR2X2_1300 ( .A(_abc_15724_n4536), .B(_abc_15724_n4537), .Y(_abc_15724_n4538) );
  OR2X2 OR2X2_1301 ( .A(_abc_15724_n3721_bF_buf1), .B(_abc_15724_n4538), .Y(_abc_15724_n4539) );
  OR2X2 OR2X2_1302 ( .A(_abc_15724_n4541), .B(_abc_15724_n4527), .Y(_abc_15724_n4542) );
  OR2X2 OR2X2_1303 ( .A(_abc_15724_n3725_bF_buf1), .B(_abc_15724_n4542), .Y(_abc_15724_n4543) );
  OR2X2 OR2X2_1304 ( .A(a_reg_5_), .B(e_reg_10_), .Y(_abc_15724_n4548) );
  OR2X2 OR2X2_1305 ( .A(_abc_15724_n4551), .B(w_10_), .Y(_abc_15724_n4554) );
  OR2X2 OR2X2_1306 ( .A(_abc_15724_n4547), .B(_abc_15724_n4555), .Y(_abc_15724_n4557) );
  OR2X2 OR2X2_1307 ( .A(_abc_15724_n4558), .B(_abc_15724_n4556), .Y(_abc_15724_n4559) );
  OR2X2 OR2X2_1308 ( .A(_abc_15724_n4561), .B(_abc_15724_n4534), .Y(_abc_15724_n4562) );
  OR2X2 OR2X2_1309 ( .A(_abc_15724_n4560), .B(_abc_15724_n4565), .Y(_abc_15724_n4566) );
  OR2X2 OR2X2_131 ( .A(_abc_15724_n1084_1), .B(_abc_15724_n1072), .Y(_abc_15724_n1085) );
  OR2X2 OR2X2_1310 ( .A(_abc_15724_n4566), .B(_abc_15724_n4523), .Y(_abc_15724_n4567) );
  OR2X2 OR2X2_1311 ( .A(_abc_15724_n4562), .B(_abc_15724_n4564), .Y(_abc_15724_n4569) );
  OR2X2 OR2X2_1312 ( .A(_abc_15724_n4559), .B(_abc_15724_n4545), .Y(_abc_15724_n4570) );
  OR2X2 OR2X2_1313 ( .A(_abc_15724_n4571), .B(_abc_15724_n4568), .Y(_abc_15724_n4572) );
  OR2X2 OR2X2_1314 ( .A(_abc_15724_n4573), .B(_abc_15724_n3737_bF_buf1), .Y(_abc_15724_n4574) );
  OR2X2 OR2X2_1315 ( .A(_abc_15724_n4576), .B(_abc_15724_n4575), .Y(_abc_15724_n4577) );
  OR2X2 OR2X2_1316 ( .A(_abc_15724_n4577), .B(_abc_15724_n3725_bF_buf0), .Y(_abc_15724_n4578) );
  OR2X2 OR2X2_1317 ( .A(_abc_15724_n4581), .B(_abc_15724_n4582), .Y(_abc_15724_n4583) );
  OR2X2 OR2X2_1318 ( .A(_abc_15724_n4584), .B(_abc_15724_n4580), .Y(_abc_15724_n4585) );
  OR2X2 OR2X2_1319 ( .A(_abc_15724_n4520), .B(_abc_15724_n4586), .Y(_abc_15724_n4589) );
  OR2X2 OR2X2_132 ( .A(_auto_iopadmap_cc_313_execute_26059_38_), .B(d_reg_6_), .Y(_abc_15724_n1086) );
  OR2X2 OR2X2_1320 ( .A(_abc_15724_n4592), .B(_abc_15724_n4594), .Y(_abc_15724_n4595) );
  OR2X2 OR2X2_1321 ( .A(_abc_15724_n4591), .B(_abc_15724_n4595), .Y(a_reg_10__FF_INPUT) );
  OR2X2 OR2X2_1322 ( .A(_abc_15724_n4582), .B(_abc_15724_n4575), .Y(_abc_15724_n4599) );
  OR2X2 OR2X2_1323 ( .A(_abc_15724_n4565), .B(_abc_15724_n4556), .Y(_abc_15724_n4600) );
  OR2X2 OR2X2_1324 ( .A(_abc_15724_n4604), .B(_abc_15724_n4605), .Y(_abc_15724_n4606) );
  OR2X2 OR2X2_1325 ( .A(_abc_15724_n4606), .B(_abc_15724_n4601), .Y(_abc_15724_n4609) );
  OR2X2 OR2X2_1326 ( .A(_abc_15724_n4612), .B(_abc_15724_n4613), .Y(_abc_15724_n4614) );
  OR2X2 OR2X2_1327 ( .A(_abc_15724_n3721_bF_buf0), .B(_abc_15724_n4614), .Y(_abc_15724_n4615) );
  OR2X2 OR2X2_1328 ( .A(_abc_15724_n4617), .B(_abc_15724_n4604), .Y(_abc_15724_n4618) );
  OR2X2 OR2X2_1329 ( .A(_abc_15724_n3725_bF_buf2), .B(_abc_15724_n4618), .Y(_abc_15724_n4619) );
  OR2X2 OR2X2_133 ( .A(_abc_15724_n1085), .B(_abc_15724_n1089), .Y(_abc_15724_n1090_1) );
  OR2X2 OR2X2_1330 ( .A(_abc_15724_n4621), .B(_abc_15724_n4611), .Y(_abc_15724_n4622) );
  OR2X2 OR2X2_1331 ( .A(a_reg_6_), .B(e_reg_11_), .Y(_abc_15724_n4625) );
  OR2X2 OR2X2_1332 ( .A(_abc_15724_n4628), .B(w_11_), .Y(_abc_15724_n4631) );
  OR2X2 OR2X2_1333 ( .A(_abc_15724_n4624), .B(_abc_15724_n4632), .Y(_abc_15724_n4635) );
  OR2X2 OR2X2_1334 ( .A(_abc_15724_n4622), .B(_abc_15724_n4636), .Y(_abc_15724_n4637) );
  OR2X2 OR2X2_1335 ( .A(_abc_15724_n4640), .B(_abc_15724_n4633), .Y(_abc_15724_n4641) );
  OR2X2 OR2X2_1336 ( .A(_abc_15724_n4641), .B(_abc_15724_n4639), .Y(_abc_15724_n4642) );
  OR2X2 OR2X2_1337 ( .A(_abc_15724_n4646), .B(_abc_15724_n4647), .Y(_abc_15724_n4648) );
  OR2X2 OR2X2_1338 ( .A(_abc_15724_n4649), .B(_abc_15724_n4644), .Y(_abc_15724_n4650) );
  OR2X2 OR2X2_1339 ( .A(_abc_15724_n4650), .B(_abc_15724_n3724), .Y(_abc_15724_n4651) );
  OR2X2 OR2X2_134 ( .A(_abc_15724_n1091_1), .B(_abc_15724_n1092_1), .Y(_abc_15724_n1093) );
  OR2X2 OR2X2_1340 ( .A(_abc_15724_n4648), .B(_abc_15724_n4645), .Y(_abc_15724_n4652) );
  OR2X2 OR2X2_1341 ( .A(_abc_15724_n4643), .B(_abc_15724_n4600), .Y(_abc_15724_n4653) );
  OR2X2 OR2X2_1342 ( .A(_abc_15724_n4654), .B(_abc_15724_n3736), .Y(_abc_15724_n4655) );
  OR2X2 OR2X2_1343 ( .A(_abc_15724_n4660), .B(_abc_15724_n4659), .Y(_abc_15724_n4661) );
  OR2X2 OR2X2_1344 ( .A(_abc_15724_n4662), .B(_abc_15724_n4657), .Y(_abc_15724_n4663) );
  OR2X2 OR2X2_1345 ( .A(_abc_15724_n4598), .B(_abc_15724_n4663), .Y(_abc_15724_n4664) );
  OR2X2 OR2X2_1346 ( .A(_abc_15724_n4665), .B(_abc_15724_n4666), .Y(_abc_15724_n4667) );
  OR2X2 OR2X2_1347 ( .A(_abc_15724_n4670), .B(_abc_15724_n4672), .Y(_abc_15724_n4673) );
  OR2X2 OR2X2_1348 ( .A(_abc_15724_n4669), .B(_abc_15724_n4673), .Y(a_reg_11__FF_INPUT) );
  OR2X2 OR2X2_1349 ( .A(_abc_15724_n4421), .B(_abc_15724_n4503), .Y(_abc_15724_n4675) );
  OR2X2 OR2X2_135 ( .A(_abc_15724_n851_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_38_), .Y(_abc_15724_n1096) );
  OR2X2 OR2X2_1350 ( .A(_abc_15724_n4663), .B(_abc_15724_n4585), .Y(_abc_15724_n4676) );
  OR2X2 OR2X2_1351 ( .A(_abc_15724_n4676), .B(_abc_15724_n4675), .Y(_abc_15724_n4677) );
  OR2X2 OR2X2_1352 ( .A(_abc_15724_n4352), .B(_abc_15724_n4677), .Y(_abc_15724_n4678) );
  OR2X2 OR2X2_1353 ( .A(_abc_15724_n4597), .B(_abc_15724_n4662), .Y(_abc_15724_n4680) );
  OR2X2 OR2X2_1354 ( .A(_abc_15724_n4518), .B(_abc_15724_n4676), .Y(_abc_15724_n4682) );
  OR2X2 OR2X2_1355 ( .A(_abc_15724_n4647), .B(_abc_15724_n4633), .Y(_abc_15724_n4687) );
  OR2X2 OR2X2_1356 ( .A(_abc_15724_n4691), .B(_abc_15724_n4692), .Y(_abc_15724_n4693) );
  OR2X2 OR2X2_1357 ( .A(_abc_15724_n4693), .B(_abc_15724_n4688), .Y(_abc_15724_n4696) );
  OR2X2 OR2X2_1358 ( .A(_abc_15724_n4700), .B(_abc_15724_n4701), .Y(_abc_15724_n4702) );
  OR2X2 OR2X2_1359 ( .A(_abc_15724_n3721_bF_buf4), .B(_abc_15724_n4702), .Y(_abc_15724_n4703) );
  OR2X2 OR2X2_136 ( .A(_abc_15724_n1095), .B(_abc_15724_n1097), .Y(H3_reg_6__FF_INPUT) );
  OR2X2 OR2X2_1360 ( .A(_abc_15724_n4705), .B(_abc_15724_n4691), .Y(_abc_15724_n4706) );
  OR2X2 OR2X2_1361 ( .A(_abc_15724_n3725_bF_buf1), .B(_abc_15724_n4706), .Y(_abc_15724_n4707) );
  OR2X2 OR2X2_1362 ( .A(a_reg_7_), .B(e_reg_12_), .Y(_abc_15724_n4713) );
  OR2X2 OR2X2_1363 ( .A(_abc_15724_n4716), .B(w_12_), .Y(_abc_15724_n4719) );
  OR2X2 OR2X2_1364 ( .A(_abc_15724_n4712), .B(_abc_15724_n4720), .Y(_abc_15724_n4723) );
  OR2X2 OR2X2_1365 ( .A(_abc_15724_n4710), .B(_abc_15724_n4724), .Y(_abc_15724_n4725) );
  OR2X2 OR2X2_1366 ( .A(_abc_15724_n4726), .B(_abc_15724_n4721), .Y(_abc_15724_n4727) );
  OR2X2 OR2X2_1367 ( .A(_abc_15724_n4727), .B(_abc_15724_n4709), .Y(_abc_15724_n4728) );
  OR2X2 OR2X2_1368 ( .A(_abc_15724_n4733), .B(_abc_15724_n4732), .Y(_abc_15724_n4734) );
  OR2X2 OR2X2_1369 ( .A(_abc_15724_n4730), .B(_abc_15724_n4735), .Y(_abc_15724_n4736) );
  OR2X2 OR2X2_137 ( .A(_auto_iopadmap_cc_313_execute_26059_39_), .B(d_reg_7_), .Y(_abc_15724_n1100) );
  OR2X2 OR2X2_1370 ( .A(_abc_15724_n4734), .B(_abc_15724_n4731), .Y(_abc_15724_n4738) );
  OR2X2 OR2X2_1371 ( .A(_abc_15724_n4729), .B(_abc_15724_n4687), .Y(_abc_15724_n4739) );
  OR2X2 OR2X2_1372 ( .A(_abc_15724_n4737), .B(_abc_15724_n4741), .Y(_abc_15724_n4742) );
  OR2X2 OR2X2_1373 ( .A(_abc_15724_n4742), .B(_abc_15724_n4686), .Y(_abc_15724_n4743) );
  OR2X2 OR2X2_1374 ( .A(_abc_15724_n4744), .B(_abc_15724_n4745), .Y(_abc_15724_n4746) );
  OR2X2 OR2X2_1375 ( .A(_abc_15724_n4685), .B(_abc_15724_n4747), .Y(_abc_15724_n4748) );
  OR2X2 OR2X2_1376 ( .A(_abc_15724_n4753), .B(_abc_15724_n4755), .Y(_abc_15724_n4756) );
  OR2X2 OR2X2_1377 ( .A(_abc_15724_n4752), .B(_abc_15724_n4756), .Y(a_reg_12__FF_INPUT) );
  OR2X2 OR2X2_1378 ( .A(_abc_15724_n4741), .B(_abc_15724_n4730), .Y(_abc_15724_n4758) );
  OR2X2 OR2X2_1379 ( .A(_abc_15724_n4763), .B(_abc_15724_n4764), .Y(_abc_15724_n4765) );
  OR2X2 OR2X2_138 ( .A(_abc_15724_n1104), .B(_abc_15724_n1087), .Y(_abc_15724_n1105) );
  OR2X2 OR2X2_1380 ( .A(_abc_15724_n4765), .B(_abc_15724_n4760), .Y(_abc_15724_n4768) );
  OR2X2 OR2X2_1381 ( .A(_abc_15724_n4772), .B(_abc_15724_n4773), .Y(_abc_15724_n4774) );
  OR2X2 OR2X2_1382 ( .A(_abc_15724_n3721_bF_buf3), .B(_abc_15724_n4774), .Y(_abc_15724_n4775) );
  OR2X2 OR2X2_1383 ( .A(_abc_15724_n4777), .B(_abc_15724_n4763), .Y(_abc_15724_n4778) );
  OR2X2 OR2X2_1384 ( .A(_abc_15724_n3725_bF_buf0), .B(_abc_15724_n4778), .Y(_abc_15724_n4779) );
  OR2X2 OR2X2_1385 ( .A(a_reg_8_), .B(e_reg_13_), .Y(_abc_15724_n4784) );
  OR2X2 OR2X2_1386 ( .A(_abc_15724_n4787), .B(w_13_), .Y(_abc_15724_n4790) );
  OR2X2 OR2X2_1387 ( .A(_abc_15724_n4783), .B(_abc_15724_n4791), .Y(_abc_15724_n4793) );
  OR2X2 OR2X2_1388 ( .A(_abc_15724_n4794), .B(_abc_15724_n4792), .Y(_abc_15724_n4795) );
  OR2X2 OR2X2_1389 ( .A(_abc_15724_n4800), .B(_abc_15724_n4796), .Y(_abc_15724_n4801) );
  OR2X2 OR2X2_139 ( .A(_abc_15724_n1105), .B(_abc_15724_n1103), .Y(_abc_15724_n1106) );
  OR2X2 OR2X2_1390 ( .A(_abc_15724_n4801), .B(_abc_15724_n4759), .Y(_abc_15724_n4802) );
  OR2X2 OR2X2_1391 ( .A(_abc_15724_n4733), .B(_abc_15724_n4721), .Y(_abc_15724_n4803) );
  OR2X2 OR2X2_1392 ( .A(_abc_15724_n4797), .B(_abc_15724_n4799), .Y(_abc_15724_n4804) );
  OR2X2 OR2X2_1393 ( .A(_abc_15724_n4795), .B(_abc_15724_n4781), .Y(_abc_15724_n4805) );
  OR2X2 OR2X2_1394 ( .A(_abc_15724_n4803), .B(_abc_15724_n4806), .Y(_abc_15724_n4807) );
  OR2X2 OR2X2_1395 ( .A(_abc_15724_n4808), .B(_abc_15724_n3736), .Y(_abc_15724_n4809) );
  OR2X2 OR2X2_1396 ( .A(_abc_15724_n4810), .B(_abc_15724_n4811), .Y(_abc_15724_n4812) );
  OR2X2 OR2X2_1397 ( .A(_abc_15724_n4812), .B(_abc_15724_n3724), .Y(_abc_15724_n4813) );
  OR2X2 OR2X2_1398 ( .A(_abc_15724_n4736), .B(_abc_15724_n3726_bF_buf2), .Y(_abc_15724_n4816) );
  OR2X2 OR2X2_1399 ( .A(_abc_15724_n4818), .B(_abc_15724_n4819), .Y(_abc_15724_n4820) );
  OR2X2 OR2X2_14 ( .A(e_reg_12_), .B(_auto_iopadmap_cc_313_execute_26059_12_), .Y(_abc_15724_n751) );
  OR2X2 OR2X2_140 ( .A(_abc_15724_n1108), .B(_abc_15724_n1107), .Y(_abc_15724_n1109_1) );
  OR2X2 OR2X2_1400 ( .A(_abc_15724_n4821), .B(_abc_15724_n4815), .Y(_abc_15724_n4822) );
  OR2X2 OR2X2_1401 ( .A(_abc_15724_n4823), .B(_abc_15724_n4744), .Y(_abc_15724_n4824) );
  OR2X2 OR2X2_1402 ( .A(_abc_15724_n4749), .B(_abc_15724_n4824), .Y(_abc_15724_n4825) );
  OR2X2 OR2X2_1403 ( .A(_abc_15724_n4746), .B(_abc_15724_n4822), .Y(_abc_15724_n4826) );
  OR2X2 OR2X2_1404 ( .A(_abc_15724_n4822), .B(_abc_15724_n4743), .Y(_abc_15724_n4830) );
  OR2X2 OR2X2_1405 ( .A(_abc_15724_n4834), .B(_abc_15724_n4835), .Y(_abc_15724_n4836) );
  OR2X2 OR2X2_1406 ( .A(_abc_15724_n4833), .B(_abc_15724_n4836), .Y(a_reg_13__FF_INPUT) );
  OR2X2 OR2X2_1407 ( .A(_abc_15724_n4848), .B(_abc_15724_n4849), .Y(_abc_15724_n4850) );
  OR2X2 OR2X2_1408 ( .A(_abc_15724_n4853), .B(_abc_15724_n4848), .Y(_abc_15724_n4854) );
  OR2X2 OR2X2_1409 ( .A(_abc_15724_n4856), .B(_abc_15724_n4851), .Y(_abc_15724_n4857) );
  OR2X2 OR2X2_141 ( .A(_abc_15724_n1111_1), .B(_abc_15724_n1099), .Y(H3_reg_7__FF_INPUT) );
  OR2X2 OR2X2_1410 ( .A(_abc_15724_n4857), .B(_abc_15724_n3806_bF_buf0), .Y(_abc_15724_n4858) );
  OR2X2 OR2X2_1411 ( .A(_abc_15724_n4853), .B(_abc_15724_n4859), .Y(_abc_15724_n4860) );
  OR2X2 OR2X2_1412 ( .A(_abc_15724_n4860), .B(_abc_15724_n3721_bF_buf2), .Y(_abc_15724_n4861) );
  OR2X2 OR2X2_1413 ( .A(a_reg_9_), .B(e_reg_14_), .Y(_abc_15724_n4868) );
  OR2X2 OR2X2_1414 ( .A(_abc_15724_n4871), .B(w_14_), .Y(_abc_15724_n4874) );
  OR2X2 OR2X2_1415 ( .A(_abc_15724_n4867), .B(_abc_15724_n4875), .Y(_abc_15724_n4878) );
  OR2X2 OR2X2_1416 ( .A(_abc_15724_n4880), .B(_abc_15724_n4865), .Y(_abc_15724_n4882) );
  OR2X2 OR2X2_1417 ( .A(_abc_15724_n4883), .B(_abc_15724_n4881), .Y(_abc_15724_n4884) );
  OR2X2 OR2X2_1418 ( .A(_abc_15724_n4884), .B(_abc_15724_n4844), .Y(_abc_15724_n4885) );
  OR2X2 OR2X2_1419 ( .A(_abc_15724_n4888), .B(_abc_15724_n4886), .Y(_abc_15724_n4889) );
  OR2X2 OR2X2_142 ( .A(_abc_15724_n1114), .B(_abc_15724_n1101), .Y(_abc_15724_n1115) );
  OR2X2 OR2X2_1420 ( .A(_abc_15724_n4890), .B(_abc_15724_n3725_bF_buf3), .Y(_abc_15724_n4891) );
  OR2X2 OR2X2_1421 ( .A(_abc_15724_n4893), .B(_abc_15724_n4892), .Y(_abc_15724_n4894) );
  OR2X2 OR2X2_1422 ( .A(_abc_15724_n4894), .B(_abc_15724_n3737_bF_buf3), .Y(_abc_15724_n4895) );
  OR2X2 OR2X2_1423 ( .A(_abc_15724_n4898), .B(_abc_15724_n4899), .Y(_abc_15724_n4900) );
  OR2X2 OR2X2_1424 ( .A(_abc_15724_n4901), .B(_abc_15724_n4897), .Y(_abc_15724_n4902) );
  OR2X2 OR2X2_1425 ( .A(_abc_15724_n4841), .B(_abc_15724_n4903), .Y(_abc_15724_n4906) );
  OR2X2 OR2X2_1426 ( .A(_abc_15724_n4909), .B(_abc_15724_n4911), .Y(_abc_15724_n4912) );
  OR2X2 OR2X2_1427 ( .A(_abc_15724_n4908), .B(_abc_15724_n4912), .Y(a_reg_14__FF_INPUT) );
  OR2X2 OR2X2_1428 ( .A(_abc_15724_n4899), .B(_abc_15724_n4892), .Y(_abc_15724_n4917) );
  OR2X2 OR2X2_1429 ( .A(_abc_15724_n4922), .B(b_reg_15_), .Y(_abc_15724_n4923) );
  OR2X2 OR2X2_143 ( .A(_auto_iopadmap_cc_313_execute_26059_40_), .B(d_reg_8_), .Y(_abc_15724_n1116) );
  OR2X2 OR2X2_1430 ( .A(c_reg_15_), .B(b_reg_15_), .Y(_abc_15724_n4926) );
  OR2X2 OR2X2_1431 ( .A(_abc_15724_n4927), .B(d_reg_15_), .Y(_abc_15724_n4928) );
  OR2X2 OR2X2_1432 ( .A(_abc_15724_n4934), .B(_abc_15724_n4935), .Y(_abc_15724_n4936) );
  OR2X2 OR2X2_1433 ( .A(_abc_15724_n3725_bF_buf1), .B(_abc_15724_n4936), .Y(_abc_15724_n4937) );
  OR2X2 OR2X2_1434 ( .A(_abc_15724_n4939), .B(_abc_15724_n4925), .Y(_abc_15724_n4940) );
  OR2X2 OR2X2_1435 ( .A(_abc_15724_n4872), .B(_abc_15724_n4869), .Y(_abc_15724_n4941) );
  OR2X2 OR2X2_1436 ( .A(a_reg_10_), .B(e_reg_15_), .Y(_abc_15724_n4942) );
  OR2X2 OR2X2_1437 ( .A(_abc_15724_n4945), .B(w_15_), .Y(_abc_15724_n4948) );
  OR2X2 OR2X2_1438 ( .A(_abc_15724_n4949), .B(_abc_15724_n4941), .Y(_abc_15724_n4952) );
  OR2X2 OR2X2_1439 ( .A(_abc_15724_n4940), .B(_abc_15724_n4954), .Y(_abc_15724_n4955) );
  OR2X2 OR2X2_144 ( .A(_abc_15724_n1115), .B(_abc_15724_n1119_1), .Y(_abc_15724_n1120_1) );
  OR2X2 OR2X2_1440 ( .A(_abc_15724_n4957), .B(_abc_15724_n4932), .Y(_abc_15724_n4958) );
  OR2X2 OR2X2_1441 ( .A(_abc_15724_n4959), .B(_abc_15724_n4953), .Y(_abc_15724_n4960) );
  OR2X2 OR2X2_1442 ( .A(_abc_15724_n4963), .B(_abc_15724_n4964), .Y(_abc_15724_n4965) );
  OR2X2 OR2X2_1443 ( .A(_abc_15724_n4962), .B(_abc_15724_n4966), .Y(_abc_15724_n4967) );
  OR2X2 OR2X2_1444 ( .A(_abc_15724_n4967), .B(_abc_15724_n3805_bF_buf2), .Y(_abc_15724_n4968) );
  OR2X2 OR2X2_1445 ( .A(_abc_15724_n4965), .B(_abc_15724_n4918), .Y(_abc_15724_n4969) );
  OR2X2 OR2X2_1446 ( .A(_abc_15724_n4961), .B(_abc_15724_n4919), .Y(_abc_15724_n4970) );
  OR2X2 OR2X2_1447 ( .A(_abc_15724_n4971), .B(_abc_15724_n3721_bF_buf0), .Y(_abc_15724_n4972) );
  OR2X2 OR2X2_1448 ( .A(_abc_15724_n4977), .B(_abc_15724_n4976), .Y(_abc_15724_n4978) );
  OR2X2 OR2X2_1449 ( .A(_abc_15724_n4979), .B(_abc_15724_n4974), .Y(_abc_15724_n4980) );
  OR2X2 OR2X2_145 ( .A(_abc_15724_n1124), .B(_abc_15724_n1113), .Y(H3_reg_8__FF_INPUT) );
  OR2X2 OR2X2_1450 ( .A(_abc_15724_n4916), .B(_abc_15724_n4981), .Y(_abc_15724_n4982) );
  OR2X2 OR2X2_1451 ( .A(_abc_15724_n4915), .B(_abc_15724_n4980), .Y(_abc_15724_n4983) );
  OR2X2 OR2X2_1452 ( .A(_abc_15724_n4986), .B(_abc_15724_n4988), .Y(_abc_15724_n4989) );
  OR2X2 OR2X2_1453 ( .A(_abc_15724_n4985), .B(_abc_15724_n4989), .Y(a_reg_15__FF_INPUT) );
  OR2X2 OR2X2_1454 ( .A(_abc_15724_n4902), .B(_abc_15724_n4980), .Y(_abc_15724_n4991) );
  OR2X2 OR2X2_1455 ( .A(_abc_15724_n4991), .B(_abc_15724_n4826), .Y(_abc_15724_n4992) );
  OR2X2 OR2X2_1456 ( .A(_abc_15724_n4992), .B(_abc_15724_n4677), .Y(_abc_15724_n4993) );
  OR2X2 OR2X2_1457 ( .A(_abc_15724_n4352), .B(_abc_15724_n4993), .Y(_abc_15724_n4994) );
  OR2X2 OR2X2_1458 ( .A(_abc_15724_n4839), .B(_abc_15724_n4991), .Y(_abc_15724_n4995) );
  OR2X2 OR2X2_1459 ( .A(_abc_15724_n4997), .B(_abc_15724_n4974), .Y(_abc_15724_n4998) );
  OR2X2 OR2X2_146 ( .A(_auto_iopadmap_cc_313_execute_26059_41_), .B(d_reg_9_), .Y(_abc_15724_n1126) );
  OR2X2 OR2X2_1460 ( .A(_abc_15724_n4683), .B(_abc_15724_n4992), .Y(_abc_15724_n5001) );
  OR2X2 OR2X2_1461 ( .A(_abc_15724_n5015), .B(d_reg_16_), .Y(_abc_15724_n5016) );
  OR2X2 OR2X2_1462 ( .A(_abc_15724_n5013), .B(d_reg_16_), .Y(_abc_15724_n5017) );
  OR2X2 OR2X2_1463 ( .A(_abc_15724_n5024), .B(_abc_15724_n5025), .Y(_abc_15724_n5026) );
  OR2X2 OR2X2_1464 ( .A(_abc_15724_n5026), .B(_abc_15724_n3721_bF_buf3), .Y(_abc_15724_n5027) );
  OR2X2 OR2X2_1465 ( .A(a_reg_11_), .B(e_reg_16_), .Y(_abc_15724_n5034) );
  OR2X2 OR2X2_1466 ( .A(_abc_15724_n5037), .B(w_16_), .Y(_abc_15724_n5040) );
  OR2X2 OR2X2_1467 ( .A(_abc_15724_n5033), .B(_abc_15724_n5041), .Y(_abc_15724_n5044) );
  OR2X2 OR2X2_1468 ( .A(_abc_15724_n5046), .B(_abc_15724_n5031), .Y(_abc_15724_n5048) );
  OR2X2 OR2X2_1469 ( .A(_abc_15724_n5049), .B(_abc_15724_n5047), .Y(_abc_15724_n5050) );
  OR2X2 OR2X2_147 ( .A(_abc_15724_n1131_1), .B(_abc_15724_n1129), .Y(_abc_15724_n1132_1) );
  OR2X2 OR2X2_1470 ( .A(_abc_15724_n5052), .B(_abc_15724_n5053), .Y(_abc_15724_n5054) );
  OR2X2 OR2X2_1471 ( .A(_abc_15724_n5058), .B(_abc_15724_n5055), .Y(_abc_15724_n5059) );
  OR2X2 OR2X2_1472 ( .A(_abc_15724_n5059), .B(_abc_15724_n5005), .Y(_abc_15724_n5060) );
  OR2X2 OR2X2_1473 ( .A(_abc_15724_n5061), .B(_abc_15724_n5062), .Y(_abc_15724_n5063) );
  OR2X2 OR2X2_1474 ( .A(_abc_15724_n5004), .B(_abc_15724_n5064), .Y(_abc_15724_n5065) );
  OR2X2 OR2X2_1475 ( .A(_abc_15724_n5070), .B(_abc_15724_n5071), .Y(_abc_15724_n5072) );
  OR2X2 OR2X2_1476 ( .A(_abc_15724_n5069), .B(_abc_15724_n5072), .Y(a_reg_16__FF_INPUT) );
  OR2X2 OR2X2_1477 ( .A(_abc_15724_n5054), .B(_abc_15724_n5006), .Y(_abc_15724_n5075) );
  OR2X2 OR2X2_1478 ( .A(_abc_15724_n5081), .B(b_reg_17_), .Y(_abc_15724_n5082) );
  OR2X2 OR2X2_1479 ( .A(c_reg_17_), .B(b_reg_17_), .Y(_abc_15724_n5086) );
  OR2X2 OR2X2_148 ( .A(_abc_15724_n1136), .B(_abc_15724_n1137), .Y(H3_reg_9__FF_INPUT) );
  OR2X2 OR2X2_1480 ( .A(_abc_15724_n5087), .B(d_reg_17_), .Y(_abc_15724_n5088) );
  OR2X2 OR2X2_1481 ( .A(_abc_15724_n5079), .B(d_reg_17_), .Y(_abc_15724_n5093) );
  OR2X2 OR2X2_1482 ( .A(_abc_15724_n5095), .B(_abc_15724_n3805_bF_buf4), .Y(_abc_15724_n5096) );
  OR2X2 OR2X2_1483 ( .A(_abc_15724_n5096), .B(_abc_15724_n5092), .Y(_abc_15724_n5097) );
  OR2X2 OR2X2_1484 ( .A(a_reg_12_), .B(e_reg_17_), .Y(_abc_15724_n5101) );
  OR2X2 OR2X2_1485 ( .A(_abc_15724_n5104), .B(w_17_), .Y(_abc_15724_n5107) );
  OR2X2 OR2X2_1486 ( .A(_abc_15724_n5100), .B(_abc_15724_n5108), .Y(_abc_15724_n5111) );
  OR2X2 OR2X2_1487 ( .A(_abc_15724_n5098), .B(_abc_15724_n5112), .Y(_abc_15724_n5115) );
  OR2X2 OR2X2_1488 ( .A(_abc_15724_n5078), .B(_abc_15724_n5116), .Y(_abc_15724_n5119) );
  OR2X2 OR2X2_1489 ( .A(_abc_15724_n5122), .B(_abc_15724_n5123), .Y(_abc_15724_n5124) );
  OR2X2 OR2X2_149 ( .A(_auto_iopadmap_cc_313_execute_26059_42_), .B(d_reg_10_), .Y(_abc_15724_n1141_1) );
  OR2X2 OR2X2_1490 ( .A(_abc_15724_n5124), .B(_abc_15724_n5076), .Y(_abc_15724_n5125) );
  OR2X2 OR2X2_1491 ( .A(_abc_15724_n5066), .B(_abc_15724_n5061), .Y(_abc_15724_n5129) );
  OR2X2 OR2X2_1492 ( .A(_abc_15724_n5129), .B(_abc_15724_n5128), .Y(_abc_15724_n5132) );
  OR2X2 OR2X2_1493 ( .A(_abc_15724_n5135), .B(_abc_15724_n5137), .Y(_abc_15724_n5138) );
  OR2X2 OR2X2_1494 ( .A(_abc_15724_n5134), .B(_abc_15724_n5138), .Y(a_reg_17__FF_INPUT) );
  OR2X2 OR2X2_1495 ( .A(_abc_15724_n5123), .B(_abc_15724_n5117), .Y(_abc_15724_n5142) );
  OR2X2 OR2X2_1496 ( .A(_abc_15724_n5148), .B(_abc_15724_n5149), .Y(_abc_15724_n5150) );
  OR2X2 OR2X2_1497 ( .A(_abc_15724_n5153), .B(_abc_15724_n5148), .Y(_abc_15724_n5154) );
  OR2X2 OR2X2_1498 ( .A(_abc_15724_n5156), .B(_abc_15724_n5151), .Y(_abc_15724_n5157) );
  OR2X2 OR2X2_1499 ( .A(_abc_15724_n5157), .B(_abc_15724_n3806_bF_buf3), .Y(_abc_15724_n5158) );
  OR2X2 OR2X2_15 ( .A(e_reg_11_), .B(_auto_iopadmap_cc_313_execute_26059_11_), .Y(_abc_15724_n756) );
  OR2X2 OR2X2_150 ( .A(_abc_15724_n1140), .B(_abc_15724_n1144_1), .Y(_abc_15724_n1145) );
  OR2X2 OR2X2_1500 ( .A(_abc_15724_n5153), .B(_abc_15724_n5159), .Y(_abc_15724_n5160) );
  OR2X2 OR2X2_1501 ( .A(_abc_15724_n5160), .B(_abc_15724_n3721_bF_buf2), .Y(_abc_15724_n5161) );
  OR2X2 OR2X2_1502 ( .A(a_reg_13_), .B(e_reg_18_), .Y(_abc_15724_n5168) );
  OR2X2 OR2X2_1503 ( .A(_abc_15724_n5171), .B(w_18_), .Y(_abc_15724_n5174) );
  OR2X2 OR2X2_1504 ( .A(_abc_15724_n5167), .B(_abc_15724_n5175), .Y(_abc_15724_n5178) );
  OR2X2 OR2X2_1505 ( .A(_abc_15724_n5180), .B(_abc_15724_n5165), .Y(_abc_15724_n5182) );
  OR2X2 OR2X2_1506 ( .A(_abc_15724_n5183), .B(_abc_15724_n5181), .Y(_abc_15724_n5184) );
  OR2X2 OR2X2_1507 ( .A(_abc_15724_n5186), .B(_abc_15724_n5187), .Y(_abc_15724_n5188) );
  OR2X2 OR2X2_1508 ( .A(_abc_15724_n5192), .B(_abc_15724_n5190), .Y(_abc_15724_n5193) );
  OR2X2 OR2X2_1509 ( .A(_abc_15724_n5141), .B(_abc_15724_n5194), .Y(_abc_15724_n5195) );
  OR2X2 OR2X2_151 ( .A(_abc_15724_n851_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_42_), .Y(_abc_15724_n1150) );
  OR2X2 OR2X2_1510 ( .A(_abc_15724_n5140), .B(_abc_15724_n5193), .Y(_abc_15724_n5196) );
  OR2X2 OR2X2_1511 ( .A(_abc_15724_n5199), .B(_abc_15724_n5200), .Y(_abc_15724_n5201) );
  OR2X2 OR2X2_1512 ( .A(_abc_15724_n5198), .B(_abc_15724_n5201), .Y(a_reg_18__FF_INPUT) );
  OR2X2 OR2X2_1513 ( .A(_abc_15724_n5211), .B(_abc_15724_n5212), .Y(_abc_15724_n5213) );
  OR2X2 OR2X2_1514 ( .A(_abc_15724_n5213), .B(_abc_15724_n5208), .Y(_abc_15724_n5216) );
  OR2X2 OR2X2_1515 ( .A(_abc_15724_n5221), .B(_abc_15724_n5222), .Y(_abc_15724_n5223) );
  OR2X2 OR2X2_1516 ( .A(_abc_15724_n5223), .B(_abc_15724_n3721_bF_buf1), .Y(_abc_15724_n5224) );
  OR2X2 OR2X2_1517 ( .A(_abc_15724_n5221), .B(_abc_15724_n5211), .Y(_abc_15724_n5225) );
  OR2X2 OR2X2_1518 ( .A(_abc_15724_n3725_bF_buf3), .B(_abc_15724_n5225), .Y(_abc_15724_n5226) );
  OR2X2 OR2X2_1519 ( .A(a_reg_14_), .B(e_reg_19_), .Y(_abc_15724_n5231) );
  OR2X2 OR2X2_152 ( .A(_abc_15724_n1149), .B(_abc_15724_n1151), .Y(H3_reg_10__FF_INPUT) );
  OR2X2 OR2X2_1520 ( .A(_abc_15724_n5234), .B(w_19_), .Y(_abc_15724_n5237) );
  OR2X2 OR2X2_1521 ( .A(_abc_15724_n5230), .B(_abc_15724_n5238), .Y(_abc_15724_n5241) );
  OR2X2 OR2X2_1522 ( .A(_abc_15724_n5243), .B(_abc_15724_n5228), .Y(_abc_15724_n5246) );
  OR2X2 OR2X2_1523 ( .A(_abc_15724_n5207), .B(_abc_15724_n5247), .Y(_abc_15724_n5250) );
  OR2X2 OR2X2_1524 ( .A(_abc_15724_n5251), .B(_abc_15724_n5056), .Y(_abc_15724_n5254) );
  OR2X2 OR2X2_1525 ( .A(_abc_15724_n5259), .B(_abc_15724_n5256), .Y(_abc_15724_n5260) );
  OR2X2 OR2X2_1526 ( .A(_abc_15724_n5205), .B(_abc_15724_n5261), .Y(_abc_15724_n5262) );
  OR2X2 OR2X2_1527 ( .A(_abc_15724_n5204), .B(_abc_15724_n5260), .Y(_abc_15724_n5263) );
  OR2X2 OR2X2_1528 ( .A(_abc_15724_n5266), .B(_abc_15724_n5268), .Y(_abc_15724_n5269) );
  OR2X2 OR2X2_1529 ( .A(_abc_15724_n5265), .B(_abc_15724_n5269), .Y(a_reg_19__FF_INPUT) );
  OR2X2 OR2X2_153 ( .A(_auto_iopadmap_cc_313_execute_26059_43_), .B(d_reg_11_), .Y(_abc_15724_n1154) );
  OR2X2 OR2X2_1530 ( .A(_abc_15724_n5256), .B(_abc_15724_n5190), .Y(_abc_15724_n5272) );
  OR2X2 OR2X2_1531 ( .A(_abc_15724_n5275), .B(_abc_15724_n5126), .Y(_abc_15724_n5276) );
  OR2X2 OR2X2_1532 ( .A(_abc_15724_n5260), .B(_abc_15724_n5193), .Y(_abc_15724_n5277) );
  OR2X2 OR2X2_1533 ( .A(_abc_15724_n5277), .B(_abc_15724_n5276), .Y(_abc_15724_n5278) );
  OR2X2 OR2X2_1534 ( .A(_abc_15724_n5280), .B(_abc_15724_n5063), .Y(_abc_15724_n5281) );
  OR2X2 OR2X2_1535 ( .A(_abc_15724_n5281), .B(_abc_15724_n5277), .Y(_abc_15724_n5282) );
  OR2X2 OR2X2_1536 ( .A(_abc_15724_n5003), .B(_abc_15724_n5282), .Y(_abc_15724_n5283) );
  OR2X2 OR2X2_1537 ( .A(_abc_15724_n5293), .B(_abc_15724_n5294), .Y(_abc_15724_n5295) );
  OR2X2 OR2X2_1538 ( .A(_abc_15724_n5298), .B(_abc_15724_n5293), .Y(_abc_15724_n5299) );
  OR2X2 OR2X2_1539 ( .A(_abc_15724_n5301), .B(_abc_15724_n5296), .Y(_abc_15724_n5302) );
  OR2X2 OR2X2_154 ( .A(_abc_15724_n1161), .B(_abc_15724_n1158), .Y(_abc_15724_n1162) );
  OR2X2 OR2X2_1540 ( .A(_abc_15724_n5302), .B(_abc_15724_n3806_bF_buf2), .Y(_abc_15724_n5303) );
  OR2X2 OR2X2_1541 ( .A(_abc_15724_n5298), .B(_abc_15724_n5304), .Y(_abc_15724_n5305) );
  OR2X2 OR2X2_1542 ( .A(_abc_15724_n5305), .B(_abc_15724_n3721_bF_buf0), .Y(_abc_15724_n5306) );
  OR2X2 OR2X2_1543 ( .A(a_reg_15_), .B(e_reg_20_), .Y(_abc_15724_n5313) );
  OR2X2 OR2X2_1544 ( .A(_abc_15724_n5316), .B(w_20_), .Y(_abc_15724_n5319) );
  OR2X2 OR2X2_1545 ( .A(_abc_15724_n5312), .B(_abc_15724_n5320), .Y(_abc_15724_n5323) );
  OR2X2 OR2X2_1546 ( .A(_abc_15724_n5325), .B(_abc_15724_n5310), .Y(_abc_15724_n5327) );
  OR2X2 OR2X2_1547 ( .A(_abc_15724_n5328), .B(_abc_15724_n5326), .Y(_abc_15724_n5329) );
  OR2X2 OR2X2_1548 ( .A(_abc_15724_n5331), .B(_abc_15724_n5332), .Y(_abc_15724_n5333) );
  OR2X2 OR2X2_1549 ( .A(_abc_15724_n5333), .B(_abc_15724_n5006), .Y(_abc_15724_n5335) );
  OR2X2 OR2X2_155 ( .A(_abc_15724_n1163), .B(_abc_15724_n1164), .Y(H3_reg_11__FF_INPUT) );
  OR2X2 OR2X2_1550 ( .A(_abc_15724_n5336), .B(_abc_15724_n5334), .Y(_abc_15724_n5337) );
  OR2X2 OR2X2_1551 ( .A(_abc_15724_n5339), .B(_abc_15724_n5340), .Y(_abc_15724_n5341) );
  OR2X2 OR2X2_1552 ( .A(_abc_15724_n5285), .B(_abc_15724_n5342), .Y(_abc_15724_n5343) );
  OR2X2 OR2X2_1553 ( .A(_abc_15724_n5284), .B(_abc_15724_n5341), .Y(_abc_15724_n5344) );
  OR2X2 OR2X2_1554 ( .A(_abc_15724_n5347), .B(_abc_15724_n5349), .Y(_abc_15724_n5350) );
  OR2X2 OR2X2_1555 ( .A(_abc_15724_n5346), .B(_abc_15724_n5350), .Y(a_reg_20__FF_INPUT) );
  OR2X2 OR2X2_1556 ( .A(_abc_15724_n5361), .B(_abc_15724_n5362), .Y(_abc_15724_n5363) );
  OR2X2 OR2X2_1557 ( .A(_abc_15724_n5366), .B(_abc_15724_n5361), .Y(_abc_15724_n5367) );
  OR2X2 OR2X2_1558 ( .A(_abc_15724_n5369), .B(_abc_15724_n5364), .Y(_abc_15724_n5370) );
  OR2X2 OR2X2_1559 ( .A(_abc_15724_n5370), .B(_abc_15724_n3806_bF_buf1), .Y(_abc_15724_n5371) );
  OR2X2 OR2X2_156 ( .A(_abc_15724_n1166_1), .B(_abc_15724_n1127), .Y(_abc_15724_n1167_1) );
  OR2X2 OR2X2_1560 ( .A(_abc_15724_n5366), .B(_abc_15724_n5372), .Y(_abc_15724_n5373) );
  OR2X2 OR2X2_1561 ( .A(_abc_15724_n5373), .B(_abc_15724_n3721_bF_buf4), .Y(_abc_15724_n5374) );
  OR2X2 OR2X2_1562 ( .A(e_reg_21_), .B(a_reg_16_), .Y(_abc_15724_n5381) );
  OR2X2 OR2X2_1563 ( .A(_abc_15724_n5384), .B(w_21_), .Y(_abc_15724_n5387) );
  OR2X2 OR2X2_1564 ( .A(_abc_15724_n5380), .B(_abc_15724_n5388), .Y(_abc_15724_n5391) );
  OR2X2 OR2X2_1565 ( .A(_abc_15724_n5393), .B(_abc_15724_n5378), .Y(_abc_15724_n5396) );
  OR2X2 OR2X2_1566 ( .A(_abc_15724_n5357), .B(_abc_15724_n5397), .Y(_abc_15724_n5400) );
  OR2X2 OR2X2_1567 ( .A(_abc_15724_n5403), .B(_abc_15724_n5404), .Y(_abc_15724_n5405) );
  OR2X2 OR2X2_1568 ( .A(_abc_15724_n5407), .B(_abc_15724_n5408), .Y(_abc_15724_n5409) );
  OR2X2 OR2X2_1569 ( .A(_abc_15724_n5410), .B(_abc_15724_n5339), .Y(_abc_15724_n5411) );
  OR2X2 OR2X2_157 ( .A(_abc_15724_n1170), .B(_abc_15724_n1155_1), .Y(_abc_15724_n1171) );
  OR2X2 OR2X2_1570 ( .A(_abc_15724_n5352), .B(_abc_15724_n5411), .Y(_abc_15724_n5412) );
  OR2X2 OR2X2_1571 ( .A(_abc_15724_n5341), .B(_abc_15724_n5409), .Y(_abc_15724_n5413) );
  OR2X2 OR2X2_1572 ( .A(_abc_15724_n5284), .B(_abc_15724_n5413), .Y(_abc_15724_n5414) );
  OR2X2 OR2X2_1573 ( .A(_abc_15724_n5409), .B(_abc_15724_n5415), .Y(_abc_15724_n5416) );
  OR2X2 OR2X2_1574 ( .A(_abc_15724_n5420), .B(_abc_15724_n5422), .Y(_abc_15724_n5423) );
  OR2X2 OR2X2_1575 ( .A(_abc_15724_n5419), .B(_abc_15724_n5423), .Y(a_reg_21__FF_INPUT) );
  OR2X2 OR2X2_1576 ( .A(_abc_15724_n5437), .B(_abc_15724_n5438), .Y(_abc_15724_n5439) );
  OR2X2 OR2X2_1577 ( .A(_abc_15724_n5442), .B(_abc_15724_n5437), .Y(_abc_15724_n5443) );
  OR2X2 OR2X2_1578 ( .A(_abc_15724_n5445), .B(_abc_15724_n5440), .Y(_abc_15724_n5446) );
  OR2X2 OR2X2_1579 ( .A(_abc_15724_n5446), .B(_abc_15724_n3806_bF_buf0), .Y(_abc_15724_n5447) );
  OR2X2 OR2X2_158 ( .A(_abc_15724_n1169), .B(_abc_15724_n1171), .Y(_abc_15724_n1172) );
  OR2X2 OR2X2_1580 ( .A(_abc_15724_n5442), .B(_abc_15724_n5448), .Y(_abc_15724_n5449) );
  OR2X2 OR2X2_1581 ( .A(_abc_15724_n5449), .B(_abc_15724_n3721_bF_buf3), .Y(_abc_15724_n5450) );
  OR2X2 OR2X2_1582 ( .A(e_reg_22_), .B(a_reg_17_), .Y(_abc_15724_n5457) );
  OR2X2 OR2X2_1583 ( .A(_abc_15724_n5460), .B(w_22_), .Y(_abc_15724_n5463) );
  OR2X2 OR2X2_1584 ( .A(_abc_15724_n5456), .B(_abc_15724_n5464), .Y(_abc_15724_n5467) );
  OR2X2 OR2X2_1585 ( .A(_abc_15724_n5469), .B(_abc_15724_n5454), .Y(_abc_15724_n5472) );
  OR2X2 OR2X2_1586 ( .A(_abc_15724_n5433), .B(_abc_15724_n5473), .Y(_abc_15724_n5476) );
  OR2X2 OR2X2_1587 ( .A(_abc_15724_n5479), .B(_abc_15724_n5480), .Y(_abc_15724_n5481) );
  OR2X2 OR2X2_1588 ( .A(_abc_15724_n5483), .B(_abc_15724_n5484), .Y(_abc_15724_n5485) );
  OR2X2 OR2X2_1589 ( .A(_abc_15724_n5428), .B(_abc_15724_n5486), .Y(_abc_15724_n5487) );
  OR2X2 OR2X2_159 ( .A(_abc_15724_n1175), .B(_abc_15724_n1172), .Y(_abc_15724_n1176) );
  OR2X2 OR2X2_1590 ( .A(_abc_15724_n5427), .B(_abc_15724_n5485), .Y(_abc_15724_n5488) );
  OR2X2 OR2X2_1591 ( .A(_abc_15724_n5491), .B(_abc_15724_n5492), .Y(_abc_15724_n5493) );
  OR2X2 OR2X2_1592 ( .A(_abc_15724_n5490), .B(_abc_15724_n5493), .Y(a_reg_22__FF_INPUT) );
  OR2X2 OR2X2_1593 ( .A(_abc_15724_n5480), .B(_abc_15724_n5474), .Y(_abc_15724_n5498) );
  OR2X2 OR2X2_1594 ( .A(_abc_15724_n5503), .B(b_reg_23_), .Y(_abc_15724_n5504) );
  OR2X2 OR2X2_1595 ( .A(c_reg_23_), .B(b_reg_23_), .Y(_abc_15724_n5508) );
  OR2X2 OR2X2_1596 ( .A(_abc_15724_n5509), .B(d_reg_23_), .Y(_abc_15724_n5510) );
  OR2X2 OR2X2_1597 ( .A(_abc_15724_n5501), .B(d_reg_23_), .Y(_abc_15724_n5515) );
  OR2X2 OR2X2_1598 ( .A(_abc_15724_n5517), .B(_abc_15724_n3805_bF_buf2), .Y(_abc_15724_n5518) );
  OR2X2 OR2X2_1599 ( .A(_abc_15724_n5518), .B(_abc_15724_n5514), .Y(_abc_15724_n5519) );
  OR2X2 OR2X2_16 ( .A(_abc_15724_n758_1), .B(_abc_15724_n755), .Y(_abc_15724_n759) );
  OR2X2 OR2X2_160 ( .A(_auto_iopadmap_cc_313_execute_26059_44_), .B(d_reg_12_), .Y(_abc_15724_n1177_1) );
  OR2X2 OR2X2_1600 ( .A(e_reg_23_), .B(a_reg_18_), .Y(_abc_15724_n5523) );
  OR2X2 OR2X2_1601 ( .A(_abc_15724_n5526), .B(w_23_), .Y(_abc_15724_n5529) );
  OR2X2 OR2X2_1602 ( .A(_abc_15724_n5522), .B(_abc_15724_n5530), .Y(_abc_15724_n5533) );
  OR2X2 OR2X2_1603 ( .A(_abc_15724_n5520), .B(_abc_15724_n5534), .Y(_abc_15724_n5537) );
  OR2X2 OR2X2_1604 ( .A(_abc_15724_n5500), .B(_abc_15724_n5538), .Y(_abc_15724_n5541) );
  OR2X2 OR2X2_1605 ( .A(_abc_15724_n5542), .B(_abc_15724_n3706), .Y(_abc_15724_n5545) );
  OR2X2 OR2X2_1606 ( .A(_abc_15724_n5550), .B(_abc_15724_n5547), .Y(_abc_15724_n5551) );
  OR2X2 OR2X2_1607 ( .A(_abc_15724_n5497), .B(_abc_15724_n5552), .Y(_abc_15724_n5553) );
  OR2X2 OR2X2_1608 ( .A(_abc_15724_n5496), .B(_abc_15724_n5551), .Y(_abc_15724_n5554) );
  OR2X2 OR2X2_1609 ( .A(_abc_15724_n5557), .B(_abc_15724_n5559), .Y(_abc_15724_n5560) );
  OR2X2 OR2X2_161 ( .A(_abc_15724_n1176), .B(_abc_15724_n1180), .Y(_abc_15724_n1181) );
  OR2X2 OR2X2_1610 ( .A(_abc_15724_n5556), .B(_abc_15724_n5560), .Y(a_reg_23__FF_INPUT) );
  OR2X2 OR2X2_1611 ( .A(_abc_15724_n5485), .B(_abc_15724_n5551), .Y(_abc_15724_n5562) );
  OR2X2 OR2X2_1612 ( .A(_abc_15724_n5413), .B(_abc_15724_n5562), .Y(_abc_15724_n5563) );
  OR2X2 OR2X2_1613 ( .A(_abc_15724_n5279), .B(_abc_15724_n5563), .Y(_abc_15724_n5564) );
  OR2X2 OR2X2_1614 ( .A(_abc_15724_n5426), .B(_abc_15724_n5562), .Y(_abc_15724_n5565) );
  OR2X2 OR2X2_1615 ( .A(_abc_15724_n5495), .B(_abc_15724_n5550), .Y(_abc_15724_n5567) );
  OR2X2 OR2X2_1616 ( .A(_abc_15724_n5282), .B(_abc_15724_n5563), .Y(_abc_15724_n5571) );
  OR2X2 OR2X2_1617 ( .A(_abc_15724_n5003), .B(_abc_15724_n5571), .Y(_abc_15724_n5572) );
  OR2X2 OR2X2_1618 ( .A(_abc_15724_n5581), .B(b_reg_24_), .Y(_abc_15724_n5582) );
  OR2X2 OR2X2_1619 ( .A(c_reg_24_), .B(b_reg_24_), .Y(_abc_15724_n5586) );
  OR2X2 OR2X2_162 ( .A(_abc_15724_n851_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_44_), .Y(_abc_15724_n1186_1) );
  OR2X2 OR2X2_1620 ( .A(_abc_15724_n5587), .B(d_reg_24_), .Y(_abc_15724_n5588) );
  OR2X2 OR2X2_1621 ( .A(_abc_15724_n5593), .B(_abc_15724_n5594), .Y(_abc_15724_n5595) );
  OR2X2 OR2X2_1622 ( .A(_abc_15724_n5597), .B(_abc_15724_n3805_bF_buf0), .Y(_abc_15724_n5598) );
  OR2X2 OR2X2_1623 ( .A(_abc_15724_n5598), .B(_abc_15724_n5592), .Y(_abc_15724_n5599) );
  OR2X2 OR2X2_1624 ( .A(e_reg_24_), .B(a_reg_19_), .Y(_abc_15724_n5603) );
  OR2X2 OR2X2_1625 ( .A(_abc_15724_n5606), .B(w_24_), .Y(_abc_15724_n5609) );
  OR2X2 OR2X2_1626 ( .A(_abc_15724_n5602), .B(_abc_15724_n5610), .Y(_abc_15724_n5613) );
  OR2X2 OR2X2_1627 ( .A(_abc_15724_n5600), .B(_abc_15724_n5614), .Y(_abc_15724_n5617) );
  OR2X2 OR2X2_1628 ( .A(_abc_15724_n5578), .B(_abc_15724_n5618), .Y(_abc_15724_n5621) );
  OR2X2 OR2X2_1629 ( .A(_abc_15724_n5624), .B(_abc_15724_n5625), .Y(_abc_15724_n5626) );
  OR2X2 OR2X2_163 ( .A(_abc_15724_n1185_1), .B(_abc_15724_n1187_1), .Y(H3_reg_12__FF_INPUT) );
  OR2X2 OR2X2_1630 ( .A(_abc_15724_n5628), .B(_abc_15724_n5629), .Y(_abc_15724_n5630) );
  OR2X2 OR2X2_1631 ( .A(_abc_15724_n5574), .B(_abc_15724_n5631), .Y(_abc_15724_n5634) );
  OR2X2 OR2X2_1632 ( .A(_abc_15724_n5637), .B(_abc_15724_n5638), .Y(_abc_15724_n5639) );
  OR2X2 OR2X2_1633 ( .A(_abc_15724_n5636), .B(_abc_15724_n5639), .Y(a_reg_24__FF_INPUT) );
  OR2X2 OR2X2_1634 ( .A(_abc_15724_n5625), .B(_abc_15724_n5619), .Y(_abc_15724_n5641) );
  OR2X2 OR2X2_1635 ( .A(_abc_15724_n5646), .B(b_reg_25_), .Y(_abc_15724_n5647) );
  OR2X2 OR2X2_1636 ( .A(c_reg_25_), .B(b_reg_25_), .Y(_abc_15724_n5651) );
  OR2X2 OR2X2_1637 ( .A(_abc_15724_n5652), .B(d_reg_25_), .Y(_abc_15724_n5653) );
  OR2X2 OR2X2_1638 ( .A(_abc_15724_n5658), .B(_abc_15724_n5659), .Y(_abc_15724_n5660) );
  OR2X2 OR2X2_1639 ( .A(_abc_15724_n5662), .B(_abc_15724_n3805_bF_buf3), .Y(_abc_15724_n5663) );
  OR2X2 OR2X2_164 ( .A(_auto_iopadmap_cc_313_execute_26059_45_), .B(d_reg_13_), .Y(_abc_15724_n1190_1) );
  OR2X2 OR2X2_1640 ( .A(_abc_15724_n5663), .B(_abc_15724_n5657), .Y(_abc_15724_n5664) );
  OR2X2 OR2X2_1641 ( .A(e_reg_25_), .B(a_reg_20_), .Y(_abc_15724_n5668) );
  OR2X2 OR2X2_1642 ( .A(_abc_15724_n5671), .B(w_25_), .Y(_abc_15724_n5674) );
  OR2X2 OR2X2_1643 ( .A(_abc_15724_n5667), .B(_abc_15724_n5675), .Y(_abc_15724_n5678) );
  OR2X2 OR2X2_1644 ( .A(_abc_15724_n5665), .B(_abc_15724_n5679), .Y(_abc_15724_n5682) );
  OR2X2 OR2X2_1645 ( .A(_abc_15724_n5643), .B(_abc_15724_n5683), .Y(_abc_15724_n5685) );
  OR2X2 OR2X2_1646 ( .A(_abc_15724_n5686), .B(_abc_15724_n5684), .Y(_abc_15724_n5687) );
  OR2X2 OR2X2_1647 ( .A(_abc_15724_n5641), .B(_abc_15724_n5687), .Y(_abc_15724_n5690) );
  OR2X2 OR2X2_1648 ( .A(_abc_15724_n5691), .B(_abc_15724_n5628), .Y(_abc_15724_n5692) );
  OR2X2 OR2X2_1649 ( .A(_abc_15724_n5632), .B(_abc_15724_n5692), .Y(_abc_15724_n5693) );
  OR2X2 OR2X2_165 ( .A(_abc_15724_n1193_1), .B(_abc_15724_n1178_1), .Y(_abc_15724_n1194) );
  OR2X2 OR2X2_1650 ( .A(_abc_15724_n5573), .B(_abc_15724_n5695), .Y(_abc_15724_n5696) );
  OR2X2 OR2X2_1651 ( .A(_abc_15724_n5702), .B(_abc_15724_n5703), .Y(_abc_15724_n5704) );
  OR2X2 OR2X2_1652 ( .A(_abc_15724_n5701), .B(_abc_15724_n5704), .Y(a_reg_25__FF_INPUT) );
  OR2X2 OR2X2_1653 ( .A(_abc_15724_n5713), .B(b_reg_26_), .Y(_abc_15724_n5714) );
  OR2X2 OR2X2_1654 ( .A(c_reg_26_), .B(b_reg_26_), .Y(_abc_15724_n5718) );
  OR2X2 OR2X2_1655 ( .A(_abc_15724_n5719), .B(d_reg_26_), .Y(_abc_15724_n5720) );
  OR2X2 OR2X2_1656 ( .A(_abc_15724_n5725), .B(_abc_15724_n5726), .Y(_abc_15724_n5727) );
  OR2X2 OR2X2_1657 ( .A(_abc_15724_n5729), .B(_abc_15724_n3805_bF_buf1), .Y(_abc_15724_n5730) );
  OR2X2 OR2X2_1658 ( .A(_abc_15724_n5730), .B(_abc_15724_n5724), .Y(_abc_15724_n5731) );
  OR2X2 OR2X2_1659 ( .A(e_reg_26_), .B(a_reg_21_), .Y(_abc_15724_n5735) );
  OR2X2 OR2X2_166 ( .A(_abc_15724_n1182), .B(_abc_15724_n1194), .Y(_abc_15724_n1195) );
  OR2X2 OR2X2_1660 ( .A(_abc_15724_n5738), .B(w_26_), .Y(_abc_15724_n5741) );
  OR2X2 OR2X2_1661 ( .A(_abc_15724_n5734), .B(_abc_15724_n5742), .Y(_abc_15724_n5745) );
  OR2X2 OR2X2_1662 ( .A(_abc_15724_n5732), .B(_abc_15724_n5746), .Y(_abc_15724_n5749) );
  OR2X2 OR2X2_1663 ( .A(_abc_15724_n5710), .B(_abc_15724_n5750), .Y(_abc_15724_n5753) );
  OR2X2 OR2X2_1664 ( .A(_abc_15724_n5756), .B(_abc_15724_n5757), .Y(_abc_15724_n5758) );
  OR2X2 OR2X2_1665 ( .A(_abc_15724_n5760), .B(_abc_15724_n5761), .Y(_abc_15724_n5762) );
  OR2X2 OR2X2_1666 ( .A(_abc_15724_n5708), .B(_abc_15724_n5763), .Y(_abc_15724_n5764) );
  OR2X2 OR2X2_1667 ( .A(_abc_15724_n5707), .B(_abc_15724_n5762), .Y(_abc_15724_n5765) );
  OR2X2 OR2X2_1668 ( .A(_abc_15724_n5768), .B(_abc_15724_n5769), .Y(_abc_15724_n5770) );
  OR2X2 OR2X2_1669 ( .A(_abc_15724_n5767), .B(_abc_15724_n5770), .Y(a_reg_26__FF_INPUT) );
  OR2X2 OR2X2_167 ( .A(_abc_15724_n1197_1), .B(_abc_15724_n1198_1), .Y(_abc_15724_n1199) );
  OR2X2 OR2X2_1670 ( .A(_abc_15724_n5757), .B(_abc_15724_n5751), .Y(_abc_15724_n5775) );
  OR2X2 OR2X2_1671 ( .A(_abc_15724_n5780), .B(b_reg_27_), .Y(_abc_15724_n5781) );
  OR2X2 OR2X2_1672 ( .A(c_reg_27_), .B(b_reg_27_), .Y(_abc_15724_n5785) );
  OR2X2 OR2X2_1673 ( .A(_abc_15724_n5786), .B(d_reg_27_), .Y(_abc_15724_n5787) );
  OR2X2 OR2X2_1674 ( .A(_abc_15724_n5792), .B(_abc_15724_n5793), .Y(_abc_15724_n5794) );
  OR2X2 OR2X2_1675 ( .A(_abc_15724_n5796), .B(_abc_15724_n3805_bF_buf4), .Y(_abc_15724_n5797) );
  OR2X2 OR2X2_1676 ( .A(_abc_15724_n5797), .B(_abc_15724_n5791), .Y(_abc_15724_n5798) );
  OR2X2 OR2X2_1677 ( .A(e_reg_27_), .B(a_reg_22_), .Y(_abc_15724_n5802) );
  OR2X2 OR2X2_1678 ( .A(_abc_15724_n5805), .B(w_27_), .Y(_abc_15724_n5808) );
  OR2X2 OR2X2_1679 ( .A(_abc_15724_n5801), .B(_abc_15724_n5809), .Y(_abc_15724_n5812) );
  OR2X2 OR2X2_168 ( .A(_abc_15724_n1202), .B(_abc_15724_n1189), .Y(H3_reg_13__FF_INPUT) );
  OR2X2 OR2X2_1680 ( .A(_abc_15724_n5799), .B(_abc_15724_n5813), .Y(_abc_15724_n5816) );
  OR2X2 OR2X2_1681 ( .A(_abc_15724_n5777), .B(_abc_15724_n5817), .Y(_abc_15724_n5819) );
  OR2X2 OR2X2_1682 ( .A(_abc_15724_n5820), .B(_abc_15724_n5818), .Y(_abc_15724_n5821) );
  OR2X2 OR2X2_1683 ( .A(_abc_15724_n5775), .B(_abc_15724_n5821), .Y(_abc_15724_n5824) );
  OR2X2 OR2X2_1684 ( .A(_abc_15724_n5774), .B(_abc_15724_n5825), .Y(_abc_15724_n5826) );
  OR2X2 OR2X2_1685 ( .A(_abc_15724_n5773), .B(_abc_15724_n5827), .Y(_abc_15724_n5828) );
  OR2X2 OR2X2_1686 ( .A(_abc_15724_n5831), .B(_abc_15724_n5833), .Y(_abc_15724_n5834) );
  OR2X2 OR2X2_1687 ( .A(_abc_15724_n5830), .B(_abc_15724_n5834), .Y(a_reg_27__FF_INPUT) );
  OR2X2 OR2X2_1688 ( .A(_abc_15724_n5573), .B(_abc_15724_n5838), .Y(_abc_15724_n5839) );
  OR2X2 OR2X2_1689 ( .A(_abc_15724_n5827), .B(_abc_15724_n5772), .Y(_abc_15724_n5843) );
  OR2X2 OR2X2_169 ( .A(_auto_iopadmap_cc_313_execute_26059_46_), .B(d_reg_14_), .Y(_abc_15724_n1206_1) );
  OR2X2 OR2X2_1690 ( .A(_abc_15724_n5852), .B(b_reg_28_), .Y(_abc_15724_n5853) );
  OR2X2 OR2X2_1691 ( .A(c_reg_28_), .B(b_reg_28_), .Y(_abc_15724_n5857) );
  OR2X2 OR2X2_1692 ( .A(_abc_15724_n5858), .B(d_reg_28_), .Y(_abc_15724_n5859) );
  OR2X2 OR2X2_1693 ( .A(_abc_15724_n5864), .B(_abc_15724_n5865), .Y(_abc_15724_n5866) );
  OR2X2 OR2X2_1694 ( .A(_abc_15724_n5868), .B(_abc_15724_n3805_bF_buf2), .Y(_abc_15724_n5869) );
  OR2X2 OR2X2_1695 ( .A(_abc_15724_n5869), .B(_abc_15724_n5863), .Y(_abc_15724_n5870) );
  OR2X2 OR2X2_1696 ( .A(e_reg_28_), .B(a_reg_23_), .Y(_abc_15724_n5874) );
  OR2X2 OR2X2_1697 ( .A(_abc_15724_n5877), .B(w_28_), .Y(_abc_15724_n5880) );
  OR2X2 OR2X2_1698 ( .A(_abc_15724_n5873), .B(_abc_15724_n5881), .Y(_abc_15724_n5884) );
  OR2X2 OR2X2_1699 ( .A(_abc_15724_n5871), .B(_abc_15724_n5885), .Y(_abc_15724_n5888) );
  OR2X2 OR2X2_17 ( .A(e_reg_10_), .B(_auto_iopadmap_cc_313_execute_26059_10_), .Y(_abc_15724_n763) );
  OR2X2 OR2X2_170 ( .A(_abc_15724_n1205), .B(_abc_15724_n1209_1), .Y(_abc_15724_n1210) );
  OR2X2 OR2X2_1700 ( .A(_abc_15724_n5849), .B(_abc_15724_n5889), .Y(_abc_15724_n5892) );
  OR2X2 OR2X2_1701 ( .A(_abc_15724_n5893), .B(_abc_15724_n3805_bF_buf0), .Y(_abc_15724_n5896) );
  OR2X2 OR2X2_1702 ( .A(_abc_15724_n5897), .B(_abc_15724_n5819), .Y(_abc_15724_n5900) );
  OR2X2 OR2X2_1703 ( .A(_abc_15724_n5847), .B(_abc_15724_n5901), .Y(_abc_15724_n5902) );
  OR2X2 OR2X2_1704 ( .A(_abc_15724_n5907), .B(_abc_15724_n5909), .Y(_abc_15724_n5910) );
  OR2X2 OR2X2_1705 ( .A(_abc_15724_n5906), .B(_abc_15724_n5910), .Y(a_reg_28__FF_INPUT) );
  OR2X2 OR2X2_1706 ( .A(_abc_15724_n5918), .B(b_reg_29_), .Y(_abc_15724_n5919) );
  OR2X2 OR2X2_1707 ( .A(c_reg_29_), .B(b_reg_29_), .Y(_abc_15724_n5923) );
  OR2X2 OR2X2_1708 ( .A(_abc_15724_n5924), .B(d_reg_29_), .Y(_abc_15724_n5925) );
  OR2X2 OR2X2_1709 ( .A(_abc_15724_n5930), .B(_abc_15724_n5931), .Y(_abc_15724_n5932) );
  OR2X2 OR2X2_171 ( .A(_abc_15724_n851_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_46_), .Y(_abc_15724_n1215_1) );
  OR2X2 OR2X2_1710 ( .A(_abc_15724_n5934), .B(_abc_15724_n3805_bF_buf3), .Y(_abc_15724_n5935) );
  OR2X2 OR2X2_1711 ( .A(_abc_15724_n5935), .B(_abc_15724_n5929), .Y(_abc_15724_n5936) );
  OR2X2 OR2X2_1712 ( .A(e_reg_29_), .B(a_reg_24_), .Y(_abc_15724_n5940) );
  OR2X2 OR2X2_1713 ( .A(_abc_15724_n5943), .B(w_29_), .Y(_abc_15724_n5946) );
  OR2X2 OR2X2_1714 ( .A(_abc_15724_n5939), .B(_abc_15724_n5947), .Y(_abc_15724_n5950) );
  OR2X2 OR2X2_1715 ( .A(_abc_15724_n5937), .B(_abc_15724_n5951), .Y(_abc_15724_n5954) );
  OR2X2 OR2X2_1716 ( .A(_abc_15724_n5915), .B(_abc_15724_n5955), .Y(_abc_15724_n5958) );
  OR2X2 OR2X2_1717 ( .A(_abc_15724_n5959), .B(_abc_15724_n4021), .Y(_abc_15724_n5962) );
  OR2X2 OR2X2_1718 ( .A(_abc_15724_n5913), .B(_abc_15724_n5963), .Y(_abc_15724_n5966) );
  OR2X2 OR2X2_1719 ( .A(_abc_15724_n5967), .B(_abc_15724_n5898), .Y(_abc_15724_n5968) );
  OR2X2 OR2X2_172 ( .A(_abc_15724_n1214), .B(_abc_15724_n1216_1), .Y(H3_reg_14__FF_INPUT) );
  OR2X2 OR2X2_1720 ( .A(_abc_15724_n5903), .B(_abc_15724_n5968), .Y(_abc_15724_n5969) );
  OR2X2 OR2X2_1721 ( .A(_abc_15724_n5846), .B(_abc_15724_n5971), .Y(_abc_15724_n5972) );
  OR2X2 OR2X2_1722 ( .A(_abc_15724_n5978), .B(_abc_15724_n5979), .Y(_abc_15724_n5980) );
  OR2X2 OR2X2_1723 ( .A(_abc_15724_n5977), .B(_abc_15724_n5980), .Y(a_reg_29__FF_INPUT) );
  OR2X2 OR2X2_1724 ( .A(_abc_15724_n5991), .B(b_reg_30_), .Y(_abc_15724_n5992) );
  OR2X2 OR2X2_1725 ( .A(c_reg_30_), .B(b_reg_30_), .Y(_abc_15724_n5996) );
  OR2X2 OR2X2_1726 ( .A(_abc_15724_n5997), .B(d_reg_30_), .Y(_abc_15724_n5998) );
  OR2X2 OR2X2_1727 ( .A(_abc_15724_n6003), .B(_abc_15724_n6004), .Y(_abc_15724_n6005) );
  OR2X2 OR2X2_1728 ( .A(_abc_15724_n6007), .B(_abc_15724_n3805_bF_buf1), .Y(_abc_15724_n6008) );
  OR2X2 OR2X2_1729 ( .A(_abc_15724_n6008), .B(_abc_15724_n6002), .Y(_abc_15724_n6009) );
  OR2X2 OR2X2_173 ( .A(_auto_iopadmap_cc_313_execute_26059_47_), .B(d_reg_15_), .Y(_abc_15724_n1219) );
  OR2X2 OR2X2_1730 ( .A(e_reg_30_), .B(a_reg_25_), .Y(_abc_15724_n6013) );
  OR2X2 OR2X2_1731 ( .A(_abc_15724_n6016), .B(w_30_), .Y(_abc_15724_n6019) );
  OR2X2 OR2X2_1732 ( .A(_abc_15724_n6012), .B(_abc_15724_n6020), .Y(_abc_15724_n6023) );
  OR2X2 OR2X2_1733 ( .A(_abc_15724_n6010), .B(_abc_15724_n6024), .Y(_abc_15724_n6027) );
  OR2X2 OR2X2_1734 ( .A(_abc_15724_n5988), .B(_abc_15724_n6028), .Y(_abc_15724_n6031) );
  OR2X2 OR2X2_1735 ( .A(_abc_15724_n6032), .B(_abc_15724_n3725_bF_buf0), .Y(_abc_15724_n6035) );
  OR2X2 OR2X2_1736 ( .A(_abc_15724_n5986), .B(_abc_15724_n6036), .Y(_abc_15724_n6039) );
  OR2X2 OR2X2_1737 ( .A(_abc_15724_n5984), .B(_abc_15724_n6040), .Y(_abc_15724_n6041) );
  OR2X2 OR2X2_1738 ( .A(_abc_15724_n5983), .B(_abc_15724_n6042), .Y(_abc_15724_n6043) );
  OR2X2 OR2X2_1739 ( .A(_abc_15724_n6046), .B(_abc_15724_n6047), .Y(_abc_15724_n6048) );
  OR2X2 OR2X2_174 ( .A(_abc_15724_n1226), .B(_abc_15724_n1223), .Y(_abc_15724_n1227) );
  OR2X2 OR2X2_1740 ( .A(_abc_15724_n6045), .B(_abc_15724_n6048), .Y(a_reg_30__FF_INPUT) );
  OR2X2 OR2X2_1741 ( .A(_abc_15724_n6057), .B(b_reg_31_), .Y(_abc_15724_n6058) );
  OR2X2 OR2X2_1742 ( .A(_abc_15724_n6061), .B(_abc_15724_n6055), .Y(_abc_15724_n6062) );
  OR2X2 OR2X2_1743 ( .A(_abc_15724_n6064), .B(_abc_15724_n6061), .Y(_abc_15724_n6065) );
  OR2X2 OR2X2_1744 ( .A(_abc_15724_n6067), .B(_abc_15724_n6063), .Y(_abc_15724_n6068) );
  OR2X2 OR2X2_1745 ( .A(_abc_15724_n6068), .B(_abc_15724_n3806_bF_buf2), .Y(_abc_15724_n6069) );
  OR2X2 OR2X2_1746 ( .A(_abc_15724_n6070), .B(_abc_15724_n3805_bF_buf4), .Y(_abc_15724_n6071) );
  OR2X2 OR2X2_1747 ( .A(_abc_15724_n6073), .B(_abc_15724_n6060), .Y(_abc_15724_n6074) );
  OR2X2 OR2X2_1748 ( .A(e_reg_31_), .B(w_31_), .Y(_abc_15724_n6076) );
  OR2X2 OR2X2_1749 ( .A(_abc_15724_n6079), .B(a_reg_26_), .Y(_abc_15724_n6082) );
  OR2X2 OR2X2_175 ( .A(_abc_15724_n1228_1), .B(_abc_15724_n1229_1), .Y(H3_reg_15__FF_INPUT) );
  OR2X2 OR2X2_1750 ( .A(_abc_15724_n6084), .B(_abc_15724_n6075), .Y(_abc_15724_n6087) );
  OR2X2 OR2X2_1751 ( .A(_abc_15724_n6074), .B(_abc_15724_n6088), .Y(_abc_15724_n6089) );
  OR2X2 OR2X2_1752 ( .A(_abc_15724_n6090), .B(_abc_15724_n6091), .Y(_abc_15724_n6092) );
  OR2X2 OR2X2_1753 ( .A(_abc_15724_n6095), .B(_abc_15724_n6096), .Y(_abc_15724_n6097) );
  OR2X2 OR2X2_1754 ( .A(_abc_15724_n6098), .B(_abc_15724_n3734), .Y(_abc_15724_n6099) );
  OR2X2 OR2X2_1755 ( .A(_abc_15724_n6097), .B(_abc_15724_n3706), .Y(_abc_15724_n6100) );
  OR2X2 OR2X2_1756 ( .A(_abc_15724_n6101), .B(_abc_15724_n6052), .Y(_abc_15724_n6104) );
  OR2X2 OR2X2_1757 ( .A(_abc_15724_n6051), .B(_abc_15724_n6106), .Y(_abc_15724_n6107) );
  OR2X2 OR2X2_1758 ( .A(_abc_15724_n6050), .B(_abc_15724_n6105), .Y(_abc_15724_n6108) );
  OR2X2 OR2X2_1759 ( .A(_abc_15724_n6111), .B(_abc_15724_n6113), .Y(_abc_15724_n6114) );
  OR2X2 OR2X2_176 ( .A(_abc_15724_n1198_1), .B(_abc_15724_n1191_1), .Y(_abc_15724_n1235) );
  OR2X2 OR2X2_1760 ( .A(_abc_15724_n6110), .B(_abc_15724_n6114), .Y(a_reg_31__FF_INPUT) );
  OR2X2 OR2X2_1761 ( .A(round_ctr_reg_5_), .B(round_ctr_reg_4_), .Y(_abc_15724_n6116) );
  OR2X2 OR2X2_1762 ( .A(_abc_15724_n6116), .B(_abc_15724_n3702), .Y(_abc_15724_n6117) );
  OR2X2 OR2X2_1763 ( .A(_abc_15724_n6123), .B(_abc_15724_n6117), .Y(_abc_15724_n6124) );
  OR2X2 OR2X2_1764 ( .A(_abc_15724_n6126), .B(round_ctr_rst_bF_buf61), .Y(_abc_15724_n3483) );
  OR2X2 OR2X2_1765 ( .A(_abc_15724_n6125), .B(_abc_15724_n6128), .Y(_abc_15724_n6129) );
  OR2X2 OR2X2_1766 ( .A(_abc_15724_n6130), .B(digest_update_bF_buf4), .Y(_abc_15724_n3489) );
  OR2X2 OR2X2_1767 ( .A(_abc_15724_n6132), .B(digest_update_bF_buf3), .Y(digest_valid_reg_FF_INPUT) );
  OR2X2 OR2X2_1768 ( .A(_abc_15724_n2992_bF_buf7), .B(_abc_15724_n6134), .Y(_abc_15724_n6135) );
  OR2X2 OR2X2_1769 ( .A(round_ctr_inc_bF_buf5), .B(round_ctr_reg_0_), .Y(_abc_15724_n6136) );
  OR2X2 OR2X2_177 ( .A(_abc_15724_n1237_1), .B(_abc_15724_n1220), .Y(_abc_15724_n1238_1) );
  OR2X2 OR2X2_1770 ( .A(round_ctr_reg_1_), .B(round_ctr_reg_0_), .Y(_abc_15724_n6140) );
  OR2X2 OR2X2_1771 ( .A(_abc_15724_n6138), .B(_abc_15724_n6142), .Y(round_ctr_reg_1__FF_INPUT) );
  OR2X2 OR2X2_1772 ( .A(_abc_15724_n6119), .B(round_ctr_reg_2_), .Y(_abc_15724_n6147) );
  OR2X2 OR2X2_1773 ( .A(_abc_15724_n6144), .B(_abc_15724_n6149), .Y(round_ctr_reg_2__FF_INPUT) );
  OR2X2 OR2X2_1774 ( .A(_abc_15724_n6145), .B(round_ctr_reg_3_), .Y(_abc_15724_n6152) );
  OR2X2 OR2X2_1775 ( .A(_abc_15724_n6154), .B(_abc_15724_n6151), .Y(round_ctr_reg_3__FF_INPUT) );
  OR2X2 OR2X2_1776 ( .A(_abc_15724_n6159), .B(_abc_15724_n6121), .Y(_abc_15724_n6160) );
  OR2X2 OR2X2_1777 ( .A(_abc_15724_n6156), .B(_abc_15724_n6164), .Y(_abc_15724_n6165) );
  OR2X2 OR2X2_1778 ( .A(_abc_15724_n6166), .B(_abc_15724_n6167), .Y(round_ctr_reg_5__FF_INPUT) );
  OR2X2 OR2X2_1779 ( .A(_abc_15724_n6169), .B(_abc_15724_n6170), .Y(_abc_15724_n6171) );
  OR2X2 OR2X2_178 ( .A(_abc_15724_n1236), .B(_abc_15724_n1238_1), .Y(_abc_15724_n1239) );
  OR2X2 OR2X2_1780 ( .A(e_reg_0_), .B(_auto_iopadmap_cc_313_execute_26059_0_), .Y(_abc_15724_n6176) );
  OR2X2 OR2X2_1781 ( .A(_abc_15724_n6177), .B(_abc_15724_n850_bF_buf5), .Y(_abc_15724_n6178) );
  OR2X2 OR2X2_1782 ( .A(_abc_15724_n2995), .B(digest_update_bF_buf2), .Y(_abc_15724_n6179) );
  OR2X2 OR2X2_1783 ( .A(_abc_15724_n794), .B(_abc_15724_n792), .Y(_abc_15724_n6181) );
  OR2X2 OR2X2_1784 ( .A(_abc_15724_n6183), .B(_abc_15724_n6184), .Y(H4_reg_1__FF_INPUT) );
  OR2X2 OR2X2_1785 ( .A(_abc_15724_n798), .B(_abc_15724_n801), .Y(_abc_15724_n6187) );
  OR2X2 OR2X2_1786 ( .A(_abc_15724_n6189), .B(_abc_15724_n6190), .Y(H4_reg_2__FF_INPUT) );
  OR2X2 OR2X2_1787 ( .A(_abc_15724_n803_1), .B(_abc_15724_n6193), .Y(_abc_15724_n6194) );
  OR2X2 OR2X2_1788 ( .A(_abc_15724_n6195), .B(_abc_15724_n6196), .Y(_abc_15724_n6197) );
  OR2X2 OR2X2_1789 ( .A(_abc_15724_n6199), .B(_abc_15724_n6200), .Y(H4_reg_3__FF_INPUT) );
  OR2X2 OR2X2_179 ( .A(_abc_15724_n1239), .B(_abc_15724_n1234), .Y(_abc_15724_n1240_1) );
  OR2X2 OR2X2_1790 ( .A(_abc_15724_n805), .B(_abc_15724_n808), .Y(_abc_15724_n6203) );
  OR2X2 OR2X2_1791 ( .A(_abc_15724_n6204), .B(_abc_15724_n850_bF_buf4), .Y(_abc_15724_n6205) );
  OR2X2 OR2X2_1792 ( .A(_abc_15724_n3019), .B(digest_update_bF_buf10), .Y(_abc_15724_n6206) );
  OR2X2 OR2X2_1793 ( .A(_abc_15724_n3025), .B(digest_update_bF_buf9), .Y(_abc_15724_n6208) );
  OR2X2 OR2X2_1794 ( .A(_abc_15724_n6214), .B(_abc_15724_n850_bF_buf3), .Y(_abc_15724_n6215) );
  OR2X2 OR2X2_1795 ( .A(_abc_15724_n6215), .B(_abc_15724_n6212), .Y(_abc_15724_n6216) );
  OR2X2 OR2X2_1796 ( .A(_abc_15724_n812_1), .B(_abc_15724_n782), .Y(_abc_15724_n6218) );
  OR2X2 OR2X2_1797 ( .A(_abc_15724_n6222), .B(_abc_15724_n6223), .Y(H4_reg_6__FF_INPUT) );
  OR2X2 OR2X2_1798 ( .A(_abc_15724_n6226), .B(_abc_15724_n779_1), .Y(_abc_15724_n6227) );
  OR2X2 OR2X2_1799 ( .A(_abc_15724_n6225), .B(_abc_15724_n6228), .Y(_abc_15724_n6229) );
  OR2X2 OR2X2_18 ( .A(e_reg_9_), .B(_auto_iopadmap_cc_313_execute_26059_9_), .Y(_abc_15724_n767_1) );
  OR2X2 OR2X2_180 ( .A(_abc_15724_n1242), .B(_abc_15724_n1240_1), .Y(_abc_15724_n1243) );
  OR2X2 OR2X2_1800 ( .A(_abc_15724_n6231), .B(_abc_15724_n6232), .Y(H4_reg_7__FF_INPUT) );
  OR2X2 OR2X2_1801 ( .A(_abc_15724_n814), .B(_abc_15724_n819), .Y(_abc_15724_n6234) );
  OR2X2 OR2X2_1802 ( .A(_abc_15724_n6238), .B(_abc_15724_n6239), .Y(H4_reg_8__FF_INPUT) );
  OR2X2 OR2X2_1803 ( .A(_abc_15724_n6245), .B(_abc_15724_n6242), .Y(_abc_15724_n6246) );
  OR2X2 OR2X2_1804 ( .A(_abc_15724_n6247), .B(_abc_15724_n6248), .Y(H4_reg_9__FF_INPUT) );
  OR2X2 OR2X2_1805 ( .A(_abc_15724_n6251), .B(_abc_15724_n770), .Y(_abc_15724_n6252) );
  OR2X2 OR2X2_1806 ( .A(_abc_15724_n6252), .B(_abc_15724_n764), .Y(_abc_15724_n6253) );
  OR2X2 OR2X2_1807 ( .A(_abc_15724_n6257), .B(_abc_15724_n6250), .Y(H4_reg_10__FF_INPUT) );
  OR2X2 OR2X2_1808 ( .A(_abc_15724_n6263), .B(_abc_15724_n6260), .Y(_abc_15724_n6264) );
  OR2X2 OR2X2_1809 ( .A(_abc_15724_n6265), .B(_abc_15724_n6266), .Y(H4_reg_11__FF_INPUT) );
  OR2X2 OR2X2_181 ( .A(_auto_iopadmap_cc_313_execute_26059_48_), .B(d_reg_16_), .Y(_abc_15724_n1244) );
  OR2X2 OR2X2_1810 ( .A(_abc_15724_n823), .B(_abc_15724_n752), .Y(_abc_15724_n6269) );
  OR2X2 OR2X2_1811 ( .A(_abc_15724_n6273), .B(_abc_15724_n6268), .Y(H4_reg_12__FF_INPUT) );
  OR2X2 OR2X2_1812 ( .A(_abc_15724_n6276), .B(_abc_15724_n750), .Y(_abc_15724_n6277) );
  OR2X2 OR2X2_1813 ( .A(_abc_15724_n6275), .B(_abc_15724_n6278), .Y(_abc_15724_n6279) );
  OR2X2 OR2X2_1814 ( .A(_abc_15724_n6281), .B(_abc_15724_n6282), .Y(H4_reg_13__FF_INPUT) );
  OR2X2 OR2X2_1815 ( .A(_abc_15724_n6284), .B(_abc_15724_n745), .Y(_abc_15724_n6285) );
  OR2X2 OR2X2_1816 ( .A(_abc_15724_n6285), .B(_abc_15724_n736), .Y(_abc_15724_n6286) );
  OR2X2 OR2X2_1817 ( .A(_abc_15724_n6290), .B(_abc_15724_n6291), .Y(H4_reg_14__FF_INPUT) );
  OR2X2 OR2X2_1818 ( .A(_abc_15724_n6297), .B(_abc_15724_n6294), .Y(_abc_15724_n6298) );
  OR2X2 OR2X2_1819 ( .A(_abc_15724_n6299), .B(_abc_15724_n6300), .Y(H4_reg_15__FF_INPUT) );
  OR2X2 OR2X2_182 ( .A(_abc_15724_n1243), .B(_abc_15724_n1247), .Y(_abc_15724_n1248) );
  OR2X2 OR2X2_1820 ( .A(_abc_15724_n825_1), .B(_abc_15724_n828), .Y(_abc_15724_n6303) );
  OR2X2 OR2X2_1821 ( .A(_abc_15724_n6307), .B(_abc_15724_n6302), .Y(H4_reg_16__FF_INPUT) );
  OR2X2 OR2X2_1822 ( .A(_abc_15724_n6310), .B(_abc_15724_n719_1), .Y(_abc_15724_n6311) );
  OR2X2 OR2X2_1823 ( .A(_abc_15724_n6309), .B(_abc_15724_n720), .Y(_abc_15724_n6312) );
  OR2X2 OR2X2_1824 ( .A(_abc_15724_n6314), .B(_abc_15724_n6315), .Y(H4_reg_17__FF_INPUT) );
  OR2X2 OR2X2_1825 ( .A(_abc_15724_n6318), .B(_abc_15724_n723), .Y(_abc_15724_n6319) );
  OR2X2 OR2X2_1826 ( .A(_abc_15724_n6319), .B(_abc_15724_n712), .Y(_abc_15724_n6320) );
  OR2X2 OR2X2_1827 ( .A(_abc_15724_n6324), .B(_abc_15724_n6317), .Y(H4_reg_18__FF_INPUT) );
  OR2X2 OR2X2_1828 ( .A(_abc_15724_n6329), .B(_abc_15724_n6330), .Y(_abc_15724_n6331) );
  OR2X2 OR2X2_1829 ( .A(_abc_15724_n6332), .B(_abc_15724_n6333), .Y(H4_reg_19__FF_INPUT) );
  OR2X2 OR2X2_183 ( .A(_abc_15724_n1252), .B(_abc_15724_n1231_1), .Y(H3_reg_16__FF_INPUT) );
  OR2X2 OR2X2_1830 ( .A(_abc_15724_n834_1), .B(_abc_15724_n837_1), .Y(_abc_15724_n6337) );
  OR2X2 OR2X2_1831 ( .A(_abc_15724_n6339), .B(_abc_15724_n6340), .Y(H4_reg_20__FF_INPUT) );
  OR2X2 OR2X2_1832 ( .A(_abc_15724_n3121), .B(digest_update_bF_buf5), .Y(_abc_15724_n6342) );
  OR2X2 OR2X2_1833 ( .A(_abc_15724_n6344), .B(_abc_15724_n702), .Y(_abc_15724_n6345) );
  OR2X2 OR2X2_1834 ( .A(_abc_15724_n6343), .B(_abc_15724_n6346), .Y(_abc_15724_n6347) );
  OR2X2 OR2X2_1835 ( .A(_abc_15724_n6348), .B(_abc_15724_n850_bF_buf3), .Y(_abc_15724_n6349) );
  OR2X2 OR2X2_1836 ( .A(w_mem_inst_w_ctr_reg_5_), .B(w_mem_inst_w_ctr_reg_4_), .Y(w_mem_inst__abc_21378_n1585) );
  OR2X2 OR2X2_1837 ( .A(w_mem_inst__abc_21378_n1585), .B(w_mem_inst_w_ctr_reg_6_), .Y(w_mem_inst__abc_21378_n1586) );
  OR2X2 OR2X2_1838 ( .A(w_mem_inst__abc_21378_n1588), .B(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_21378_n1589) );
  OR2X2 OR2X2_1839 ( .A(w_mem_inst__abc_21378_n1590), .B(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_21378_n1591) );
  OR2X2 OR2X2_184 ( .A(_auto_iopadmap_cc_313_execute_26059_49_), .B(d_reg_17_), .Y(_abc_15724_n1256) );
  OR2X2 OR2X2_1840 ( .A(w_mem_inst_w_mem_2__31_), .B(w_mem_inst_w_mem_0__31_), .Y(w_mem_inst__abc_21378_n1594_1) );
  OR2X2 OR2X2_1841 ( .A(w_mem_inst__abc_21378_n1593), .B(w_mem_inst__abc_21378_n1597), .Y(w_mem_inst__abc_21378_n1598) );
  OR2X2 OR2X2_1842 ( .A(w_mem_inst__abc_21378_n1599_1), .B(w_mem_inst__abc_21378_n1592), .Y(w_mem_inst__abc_21378_n1600) );
  OR2X2 OR2X2_1843 ( .A(w_mem_inst__abc_21378_n1601_1), .B(w_mem_inst__abc_21378_n1587_bF_buf4), .Y(w_mem_inst__abc_21378_n1602) );
  OR2X2 OR2X2_1844 ( .A(w_mem_inst__abc_21378_n1611_1), .B(w_mem_inst__abc_21378_n1586_bF_buf3), .Y(w_mem_inst__abc_21378_n1612) );
  OR2X2 OR2X2_1845 ( .A(w_mem_inst__abc_21378_n1617), .B(w_mem_inst__abc_21378_n1619_1), .Y(w_mem_inst__abc_21378_n1620) );
  OR2X2 OR2X2_1846 ( .A(w_mem_inst__abc_21378_n1620), .B(w_mem_inst__abc_21378_n1612), .Y(w_mem_inst__abc_21378_n1621) );
  OR2X2 OR2X2_1847 ( .A(w_mem_inst__abc_21378_n1621), .B(w_mem_inst__abc_21378_n1606_1), .Y(w_mem_inst__abc_21378_n1622_1) );
  OR2X2 OR2X2_1848 ( .A(w_mem_inst__abc_21378_n1626_1), .B(w_mem_inst__abc_21378_n1628), .Y(w_mem_inst__abc_21378_n1629) );
  OR2X2 OR2X2_1849 ( .A(w_mem_inst__abc_21378_n1635_1), .B(w_mem_inst__abc_21378_n1631_1), .Y(w_mem_inst__abc_21378_n1636) );
  OR2X2 OR2X2_185 ( .A(_abc_15724_n1255), .B(_abc_15724_n1259_1), .Y(_abc_15724_n1260_1) );
  OR2X2 OR2X2_1850 ( .A(w_mem_inst__abc_21378_n1629), .B(w_mem_inst__abc_21378_n1636), .Y(w_mem_inst__abc_21378_n1637) );
  OR2X2 OR2X2_1851 ( .A(w_mem_inst__abc_21378_n1639_1), .B(w_mem_inst__abc_21378_n1641), .Y(w_mem_inst__abc_21378_n1642_1) );
  OR2X2 OR2X2_1852 ( .A(w_mem_inst__abc_21378_n1644), .B(w_mem_inst__abc_21378_n1646_1), .Y(w_mem_inst__abc_21378_n1647_1) );
  OR2X2 OR2X2_1853 ( .A(w_mem_inst__abc_21378_n1642_1), .B(w_mem_inst__abc_21378_n1647_1), .Y(w_mem_inst__abc_21378_n1648) );
  OR2X2 OR2X2_1854 ( .A(w_mem_inst__abc_21378_n1650_1), .B(w_mem_inst__abc_21378_n1652), .Y(w_mem_inst__abc_21378_n1653) );
  OR2X2 OR2X2_1855 ( .A(w_mem_inst__abc_21378_n1655_1), .B(w_mem_inst__abc_21378_n1657), .Y(w_mem_inst__abc_21378_n1658_1) );
  OR2X2 OR2X2_1856 ( .A(w_mem_inst__abc_21378_n1653), .B(w_mem_inst__abc_21378_n1658_1), .Y(w_mem_inst__abc_21378_n1659_1) );
  OR2X2 OR2X2_1857 ( .A(w_mem_inst__abc_21378_n1659_1), .B(w_mem_inst__abc_21378_n1648), .Y(w_mem_inst__abc_21378_n1660) );
  OR2X2 OR2X2_1858 ( .A(w_mem_inst__abc_21378_n1660), .B(w_mem_inst__abc_21378_n1637), .Y(w_mem_inst__abc_21378_n1661) );
  OR2X2 OR2X2_1859 ( .A(w_mem_inst__abc_21378_n1661), .B(w_mem_inst__abc_21378_n1622_1), .Y(w_mem_inst__abc_21378_n1662_1) );
  OR2X2 OR2X2_186 ( .A(_abc_15724_n1254), .B(_abc_15724_n1261_1), .Y(_abc_15724_n1262) );
  OR2X2 OR2X2_1860 ( .A(w_mem_inst__abc_21378_n1664), .B(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_21378_n1665) );
  OR2X2 OR2X2_1861 ( .A(w_mem_inst__abc_21378_n1666_1), .B(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_21378_n1667_1) );
  OR2X2 OR2X2_1862 ( .A(w_mem_inst_w_mem_2__0_), .B(w_mem_inst_w_mem_0__0_), .Y(w_mem_inst__abc_21378_n1670_1) );
  OR2X2 OR2X2_1863 ( .A(w_mem_inst__abc_21378_n1669), .B(w_mem_inst__abc_21378_n1673), .Y(w_mem_inst__abc_21378_n1674_1) );
  OR2X2 OR2X2_1864 ( .A(w_mem_inst__abc_21378_n1675_1), .B(w_mem_inst__abc_21378_n1668), .Y(w_mem_inst__abc_21378_n1676) );
  OR2X2 OR2X2_1865 ( .A(w_mem_inst__abc_21378_n1677), .B(w_mem_inst__abc_21378_n1587_bF_buf3), .Y(w_mem_inst__abc_21378_n1678_1) );
  OR2X2 OR2X2_1866 ( .A(w_mem_inst__abc_21378_n1680), .B(w_mem_inst__abc_21378_n1586_bF_buf2), .Y(w_mem_inst__abc_21378_n1681) );
  OR2X2 OR2X2_1867 ( .A(w_mem_inst__abc_21378_n1682_1), .B(w_mem_inst__abc_21378_n1683_1), .Y(w_mem_inst__abc_21378_n1684) );
  OR2X2 OR2X2_1868 ( .A(w_mem_inst__abc_21378_n1684), .B(w_mem_inst__abc_21378_n1681), .Y(w_mem_inst__abc_21378_n1685) );
  OR2X2 OR2X2_1869 ( .A(w_mem_inst__abc_21378_n1685), .B(w_mem_inst__abc_21378_n1679_1), .Y(w_mem_inst__abc_21378_n1686_1) );
  OR2X2 OR2X2_187 ( .A(_abc_15724_n851_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_49_), .Y(_abc_15724_n1265) );
  OR2X2 OR2X2_1870 ( .A(w_mem_inst__abc_21378_n1687_1), .B(w_mem_inst__abc_21378_n1688), .Y(w_mem_inst__abc_21378_n1689) );
  OR2X2 OR2X2_1871 ( .A(w_mem_inst__abc_21378_n1691_1), .B(w_mem_inst__abc_21378_n1690_1), .Y(w_mem_inst__abc_21378_n1692) );
  OR2X2 OR2X2_1872 ( .A(w_mem_inst__abc_21378_n1689), .B(w_mem_inst__abc_21378_n1692), .Y(w_mem_inst__abc_21378_n1693) );
  OR2X2 OR2X2_1873 ( .A(w_mem_inst__abc_21378_n1694_1), .B(w_mem_inst__abc_21378_n1695_1), .Y(w_mem_inst__abc_21378_n1696) );
  OR2X2 OR2X2_1874 ( .A(w_mem_inst__abc_21378_n1697), .B(w_mem_inst__abc_21378_n1698_1), .Y(w_mem_inst__abc_21378_n1699_1) );
  OR2X2 OR2X2_1875 ( .A(w_mem_inst__abc_21378_n1696), .B(w_mem_inst__abc_21378_n1699_1), .Y(w_mem_inst__abc_21378_n1700) );
  OR2X2 OR2X2_1876 ( .A(w_mem_inst__abc_21378_n1701), .B(w_mem_inst__abc_21378_n1702_1), .Y(w_mem_inst__abc_21378_n1703_1) );
  OR2X2 OR2X2_1877 ( .A(w_mem_inst__abc_21378_n1704), .B(w_mem_inst__abc_21378_n1705), .Y(w_mem_inst__abc_21378_n1706_1) );
  OR2X2 OR2X2_1878 ( .A(w_mem_inst__abc_21378_n1703_1), .B(w_mem_inst__abc_21378_n1706_1), .Y(w_mem_inst__abc_21378_n1707_1) );
  OR2X2 OR2X2_1879 ( .A(w_mem_inst__abc_21378_n1707_1), .B(w_mem_inst__abc_21378_n1700), .Y(w_mem_inst__abc_21378_n1708) );
  OR2X2 OR2X2_188 ( .A(_abc_15724_n1264), .B(_abc_15724_n1266), .Y(H3_reg_17__FF_INPUT) );
  OR2X2 OR2X2_1880 ( .A(w_mem_inst__abc_21378_n1708), .B(w_mem_inst__abc_21378_n1693), .Y(w_mem_inst__abc_21378_n1709) );
  OR2X2 OR2X2_1881 ( .A(w_mem_inst__abc_21378_n1709), .B(w_mem_inst__abc_21378_n1686_1), .Y(w_mem_inst__abc_21378_n1710_1) );
  OR2X2 OR2X2_1882 ( .A(w_mem_inst__abc_21378_n1712), .B(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_21378_n1713) );
  OR2X2 OR2X2_1883 ( .A(w_mem_inst__abc_21378_n1714_1), .B(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_21378_n1715_1) );
  OR2X2 OR2X2_1884 ( .A(w_mem_inst_w_mem_2__1_), .B(w_mem_inst_w_mem_0__1_), .Y(w_mem_inst__abc_21378_n1718_1) );
  OR2X2 OR2X2_1885 ( .A(w_mem_inst__abc_21378_n1717), .B(w_mem_inst__abc_21378_n1721), .Y(w_mem_inst__abc_21378_n1722_1) );
  OR2X2 OR2X2_1886 ( .A(w_mem_inst__abc_21378_n1723_1), .B(w_mem_inst__abc_21378_n1716), .Y(w_mem_inst__abc_21378_n1724) );
  OR2X2 OR2X2_1887 ( .A(w_mem_inst__abc_21378_n1725), .B(w_mem_inst__abc_21378_n1587_bF_buf2), .Y(w_mem_inst__abc_21378_n1726_1) );
  OR2X2 OR2X2_1888 ( .A(w_mem_inst__abc_21378_n1728), .B(w_mem_inst__abc_21378_n1586_bF_buf1), .Y(w_mem_inst__abc_21378_n1729) );
  OR2X2 OR2X2_1889 ( .A(w_mem_inst__abc_21378_n1730_1), .B(w_mem_inst__abc_21378_n1731_1), .Y(w_mem_inst__abc_21378_n1732) );
  OR2X2 OR2X2_189 ( .A(_auto_iopadmap_cc_313_execute_26059_50_), .B(d_reg_18_), .Y(_abc_15724_n1269) );
  OR2X2 OR2X2_1890 ( .A(w_mem_inst__abc_21378_n1732), .B(w_mem_inst__abc_21378_n1729), .Y(w_mem_inst__abc_21378_n1733) );
  OR2X2 OR2X2_1891 ( .A(w_mem_inst__abc_21378_n1733), .B(w_mem_inst__abc_21378_n1727_1), .Y(w_mem_inst__abc_21378_n1734_1) );
  OR2X2 OR2X2_1892 ( .A(w_mem_inst__abc_21378_n1735_1), .B(w_mem_inst__abc_21378_n1736), .Y(w_mem_inst__abc_21378_n1737) );
  OR2X2 OR2X2_1893 ( .A(w_mem_inst__abc_21378_n1739_1), .B(w_mem_inst__abc_21378_n1738_1), .Y(w_mem_inst__abc_21378_n1740) );
  OR2X2 OR2X2_1894 ( .A(w_mem_inst__abc_21378_n1737), .B(w_mem_inst__abc_21378_n1740), .Y(w_mem_inst__abc_21378_n1741) );
  OR2X2 OR2X2_1895 ( .A(w_mem_inst__abc_21378_n1742_1), .B(w_mem_inst__abc_21378_n1743_1), .Y(w_mem_inst__abc_21378_n1744) );
  OR2X2 OR2X2_1896 ( .A(w_mem_inst__abc_21378_n1745), .B(w_mem_inst__abc_21378_n1746_1), .Y(w_mem_inst__abc_21378_n1747_1) );
  OR2X2 OR2X2_1897 ( .A(w_mem_inst__abc_21378_n1747_1), .B(w_mem_inst__abc_21378_n1744), .Y(w_mem_inst__abc_21378_n1748) );
  OR2X2 OR2X2_1898 ( .A(w_mem_inst__abc_21378_n1750_1), .B(w_mem_inst__abc_21378_n1749), .Y(w_mem_inst__abc_21378_n1751_1) );
  OR2X2 OR2X2_1899 ( .A(w_mem_inst__abc_21378_n1752), .B(w_mem_inst__abc_21378_n1753), .Y(w_mem_inst__abc_21378_n1754_1) );
  OR2X2 OR2X2_19 ( .A(_abc_15724_n769_1), .B(_abc_15724_n766_1), .Y(_abc_15724_n770) );
  OR2X2 OR2X2_190 ( .A(_abc_15724_n1275_1), .B(_abc_15724_n1273), .Y(_abc_15724_n1276_1) );
  OR2X2 OR2X2_1900 ( .A(w_mem_inst__abc_21378_n1754_1), .B(w_mem_inst__abc_21378_n1751_1), .Y(w_mem_inst__abc_21378_n1755_1) );
  OR2X2 OR2X2_1901 ( .A(w_mem_inst__abc_21378_n1748), .B(w_mem_inst__abc_21378_n1755_1), .Y(w_mem_inst__abc_21378_n1756) );
  OR2X2 OR2X2_1902 ( .A(w_mem_inst__abc_21378_n1756), .B(w_mem_inst__abc_21378_n1741), .Y(w_mem_inst__abc_21378_n1757) );
  OR2X2 OR2X2_1903 ( .A(w_mem_inst__abc_21378_n1757), .B(w_mem_inst__abc_21378_n1734_1), .Y(w_mem_inst__abc_21378_n1758_1) );
  OR2X2 OR2X2_1904 ( .A(w_mem_inst__abc_21378_n1760), .B(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_21378_n1761) );
  OR2X2 OR2X2_1905 ( .A(w_mem_inst__abc_21378_n1762_1), .B(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_21378_n1763_1) );
  OR2X2 OR2X2_1906 ( .A(w_mem_inst_w_mem_2__2_), .B(w_mem_inst_w_mem_0__2_), .Y(w_mem_inst__abc_21378_n1766_1) );
  OR2X2 OR2X2_1907 ( .A(w_mem_inst__abc_21378_n1765), .B(w_mem_inst__abc_21378_n1769), .Y(w_mem_inst__abc_21378_n1770_1) );
  OR2X2 OR2X2_1908 ( .A(w_mem_inst__abc_21378_n1771_1), .B(w_mem_inst__abc_21378_n1764), .Y(w_mem_inst__abc_21378_n1772) );
  OR2X2 OR2X2_1909 ( .A(w_mem_inst__abc_21378_n1773), .B(w_mem_inst__abc_21378_n1587_bF_buf1), .Y(w_mem_inst__abc_21378_n1774_1) );
  OR2X2 OR2X2_191 ( .A(_abc_15724_n1277), .B(_abc_15724_n1272), .Y(_abc_15724_n1278) );
  OR2X2 OR2X2_1910 ( .A(w_mem_inst__abc_21378_n1776), .B(w_mem_inst__abc_21378_n1586_bF_buf0), .Y(w_mem_inst__abc_21378_n1777) );
  OR2X2 OR2X2_1911 ( .A(w_mem_inst__abc_21378_n1778_1), .B(w_mem_inst__abc_21378_n1779_1), .Y(w_mem_inst__abc_21378_n1780) );
  OR2X2 OR2X2_1912 ( .A(w_mem_inst__abc_21378_n1780), .B(w_mem_inst__abc_21378_n1777), .Y(w_mem_inst__abc_21378_n1781) );
  OR2X2 OR2X2_1913 ( .A(w_mem_inst__abc_21378_n1781), .B(w_mem_inst__abc_21378_n1775_1), .Y(w_mem_inst__abc_21378_n1782_1) );
  OR2X2 OR2X2_1914 ( .A(w_mem_inst__abc_21378_n1783_1), .B(w_mem_inst__abc_21378_n1784), .Y(w_mem_inst__abc_21378_n1785) );
  OR2X2 OR2X2_1915 ( .A(w_mem_inst__abc_21378_n1787_1), .B(w_mem_inst__abc_21378_n1786_1), .Y(w_mem_inst__abc_21378_n1788) );
  OR2X2 OR2X2_1916 ( .A(w_mem_inst__abc_21378_n1785), .B(w_mem_inst__abc_21378_n1788), .Y(w_mem_inst__abc_21378_n1789) );
  OR2X2 OR2X2_1917 ( .A(w_mem_inst__abc_21378_n1790_1), .B(w_mem_inst__abc_21378_n1791_1), .Y(w_mem_inst__abc_21378_n1792) );
  OR2X2 OR2X2_1918 ( .A(w_mem_inst__abc_21378_n1793), .B(w_mem_inst__abc_21378_n1794_1), .Y(w_mem_inst__abc_21378_n1795_1) );
  OR2X2 OR2X2_1919 ( .A(w_mem_inst__abc_21378_n1792), .B(w_mem_inst__abc_21378_n1795_1), .Y(w_mem_inst__abc_21378_n1796) );
  OR2X2 OR2X2_192 ( .A(_abc_15724_n1282), .B(_abc_15724_n1268), .Y(H3_reg_18__FF_INPUT) );
  OR2X2 OR2X2_1920 ( .A(w_mem_inst__abc_21378_n1797), .B(w_mem_inst__abc_21378_n1798_1), .Y(w_mem_inst__abc_21378_n1799_1) );
  OR2X2 OR2X2_1921 ( .A(w_mem_inst__abc_21378_n1800), .B(w_mem_inst__abc_21378_n1801), .Y(w_mem_inst__abc_21378_n1802_1) );
  OR2X2 OR2X2_1922 ( .A(w_mem_inst__abc_21378_n1799_1), .B(w_mem_inst__abc_21378_n1802_1), .Y(w_mem_inst__abc_21378_n1803_1) );
  OR2X2 OR2X2_1923 ( .A(w_mem_inst__abc_21378_n1803_1), .B(w_mem_inst__abc_21378_n1796), .Y(w_mem_inst__abc_21378_n1804) );
  OR2X2 OR2X2_1924 ( .A(w_mem_inst__abc_21378_n1804), .B(w_mem_inst__abc_21378_n1789), .Y(w_mem_inst__abc_21378_n1805) );
  OR2X2 OR2X2_1925 ( .A(w_mem_inst__abc_21378_n1805), .B(w_mem_inst__abc_21378_n1782_1), .Y(w_mem_inst__abc_21378_n1806_1) );
  OR2X2 OR2X2_1926 ( .A(w_mem_inst__abc_21378_n1808), .B(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_21378_n1809) );
  OR2X2 OR2X2_1927 ( .A(w_mem_inst__abc_21378_n1810_1), .B(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_21378_n1811_1) );
  OR2X2 OR2X2_1928 ( .A(w_mem_inst_w_mem_2__3_), .B(w_mem_inst_w_mem_0__3_), .Y(w_mem_inst__abc_21378_n1814_1) );
  OR2X2 OR2X2_1929 ( .A(w_mem_inst__abc_21378_n1813), .B(w_mem_inst__abc_21378_n1817), .Y(w_mem_inst__abc_21378_n1818_1) );
  OR2X2 OR2X2_193 ( .A(_auto_iopadmap_cc_313_execute_26059_51_), .B(d_reg_19_), .Y(_abc_15724_n1285_1) );
  OR2X2 OR2X2_1930 ( .A(w_mem_inst__abc_21378_n1819_1), .B(w_mem_inst__abc_21378_n1812), .Y(w_mem_inst__abc_21378_n1820) );
  OR2X2 OR2X2_1931 ( .A(w_mem_inst__abc_21378_n1821), .B(w_mem_inst__abc_21378_n1587_bF_buf0), .Y(w_mem_inst__abc_21378_n1822_1) );
  OR2X2 OR2X2_1932 ( .A(w_mem_inst__abc_21378_n1824), .B(w_mem_inst__abc_21378_n1586_bF_buf4), .Y(w_mem_inst__abc_21378_n1825) );
  OR2X2 OR2X2_1933 ( .A(w_mem_inst__abc_21378_n1826_1), .B(w_mem_inst__abc_21378_n1827_1), .Y(w_mem_inst__abc_21378_n1828) );
  OR2X2 OR2X2_1934 ( .A(w_mem_inst__abc_21378_n1828), .B(w_mem_inst__abc_21378_n1825), .Y(w_mem_inst__abc_21378_n1829) );
  OR2X2 OR2X2_1935 ( .A(w_mem_inst__abc_21378_n1829), .B(w_mem_inst__abc_21378_n1823_1), .Y(w_mem_inst__abc_21378_n1830_1) );
  OR2X2 OR2X2_1936 ( .A(w_mem_inst__abc_21378_n1831_1), .B(w_mem_inst__abc_21378_n1832), .Y(w_mem_inst__abc_21378_n1833) );
  OR2X2 OR2X2_1937 ( .A(w_mem_inst__abc_21378_n1835_1), .B(w_mem_inst__abc_21378_n1834_1), .Y(w_mem_inst__abc_21378_n1836) );
  OR2X2 OR2X2_1938 ( .A(w_mem_inst__abc_21378_n1833), .B(w_mem_inst__abc_21378_n1836), .Y(w_mem_inst__abc_21378_n1837) );
  OR2X2 OR2X2_1939 ( .A(w_mem_inst__abc_21378_n1838_1), .B(w_mem_inst__abc_21378_n1839_1), .Y(w_mem_inst__abc_21378_n1840) );
  OR2X2 OR2X2_194 ( .A(_abc_15724_n1292), .B(_abc_15724_n1289), .Y(_abc_15724_n1293) );
  OR2X2 OR2X2_1940 ( .A(w_mem_inst__abc_21378_n1841), .B(w_mem_inst__abc_21378_n1842_1), .Y(w_mem_inst__abc_21378_n1843_1) );
  OR2X2 OR2X2_1941 ( .A(w_mem_inst__abc_21378_n1843_1), .B(w_mem_inst__abc_21378_n1840), .Y(w_mem_inst__abc_21378_n1844) );
  OR2X2 OR2X2_1942 ( .A(w_mem_inst__abc_21378_n1846_1), .B(w_mem_inst__abc_21378_n1845), .Y(w_mem_inst__abc_21378_n1847_1) );
  OR2X2 OR2X2_1943 ( .A(w_mem_inst__abc_21378_n1848), .B(w_mem_inst__abc_21378_n1849), .Y(w_mem_inst__abc_21378_n1850_1) );
  OR2X2 OR2X2_1944 ( .A(w_mem_inst__abc_21378_n1850_1), .B(w_mem_inst__abc_21378_n1847_1), .Y(w_mem_inst__abc_21378_n1851_1) );
  OR2X2 OR2X2_1945 ( .A(w_mem_inst__abc_21378_n1844), .B(w_mem_inst__abc_21378_n1851_1), .Y(w_mem_inst__abc_21378_n1852) );
  OR2X2 OR2X2_1946 ( .A(w_mem_inst__abc_21378_n1852), .B(w_mem_inst__abc_21378_n1837), .Y(w_mem_inst__abc_21378_n1853) );
  OR2X2 OR2X2_1947 ( .A(w_mem_inst__abc_21378_n1853), .B(w_mem_inst__abc_21378_n1830_1), .Y(w_mem_inst__abc_21378_n1854_1) );
  OR2X2 OR2X2_1948 ( .A(w_mem_inst__abc_21378_n1856), .B(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_21378_n1857) );
  OR2X2 OR2X2_1949 ( .A(w_mem_inst__abc_21378_n1858_1), .B(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_21378_n1859_1) );
  OR2X2 OR2X2_195 ( .A(_abc_15724_n1294), .B(_abc_15724_n1295), .Y(H3_reg_19__FF_INPUT) );
  OR2X2 OR2X2_1950 ( .A(w_mem_inst_w_mem_2__4_), .B(w_mem_inst_w_mem_0__4_), .Y(w_mem_inst__abc_21378_n1862_1) );
  OR2X2 OR2X2_1951 ( .A(w_mem_inst__abc_21378_n1861), .B(w_mem_inst__abc_21378_n1865), .Y(w_mem_inst__abc_21378_n1866_1) );
  OR2X2 OR2X2_1952 ( .A(w_mem_inst__abc_21378_n1867_1), .B(w_mem_inst__abc_21378_n1860), .Y(w_mem_inst__abc_21378_n1868) );
  OR2X2 OR2X2_1953 ( .A(w_mem_inst__abc_21378_n1869), .B(w_mem_inst__abc_21378_n1587_bF_buf4), .Y(w_mem_inst__abc_21378_n1870_1) );
  OR2X2 OR2X2_1954 ( .A(w_mem_inst__abc_21378_n1872), .B(w_mem_inst__abc_21378_n1586_bF_buf3), .Y(w_mem_inst__abc_21378_n1873) );
  OR2X2 OR2X2_1955 ( .A(w_mem_inst__abc_21378_n1874_1), .B(w_mem_inst__abc_21378_n1875_1), .Y(w_mem_inst__abc_21378_n1876) );
  OR2X2 OR2X2_1956 ( .A(w_mem_inst__abc_21378_n1876), .B(w_mem_inst__abc_21378_n1873), .Y(w_mem_inst__abc_21378_n1877) );
  OR2X2 OR2X2_1957 ( .A(w_mem_inst__abc_21378_n1877), .B(w_mem_inst__abc_21378_n1871_1), .Y(w_mem_inst__abc_21378_n1878_1) );
  OR2X2 OR2X2_1958 ( .A(w_mem_inst__abc_21378_n1879_1), .B(w_mem_inst__abc_21378_n1880), .Y(w_mem_inst__abc_21378_n1881) );
  OR2X2 OR2X2_1959 ( .A(w_mem_inst__abc_21378_n1883_1), .B(w_mem_inst__abc_21378_n1882_1), .Y(w_mem_inst__abc_21378_n1884) );
  OR2X2 OR2X2_196 ( .A(_abc_15724_n1274_1), .B(_abc_15724_n1273), .Y(_abc_15724_n1297_1) );
  OR2X2 OR2X2_1960 ( .A(w_mem_inst__abc_21378_n1881), .B(w_mem_inst__abc_21378_n1884), .Y(w_mem_inst__abc_21378_n1885) );
  OR2X2 OR2X2_1961 ( .A(w_mem_inst__abc_21378_n1886_1), .B(w_mem_inst__abc_21378_n1887_1), .Y(w_mem_inst__abc_21378_n1888) );
  OR2X2 OR2X2_1962 ( .A(w_mem_inst__abc_21378_n1889), .B(w_mem_inst__abc_21378_n1890_1), .Y(w_mem_inst__abc_21378_n1891_1) );
  OR2X2 OR2X2_1963 ( .A(w_mem_inst__abc_21378_n1888), .B(w_mem_inst__abc_21378_n1891_1), .Y(w_mem_inst__abc_21378_n1892) );
  OR2X2 OR2X2_1964 ( .A(w_mem_inst__abc_21378_n1893), .B(w_mem_inst__abc_21378_n1894_1), .Y(w_mem_inst__abc_21378_n1895_1) );
  OR2X2 OR2X2_1965 ( .A(w_mem_inst__abc_21378_n1896), .B(w_mem_inst__abc_21378_n1897), .Y(w_mem_inst__abc_21378_n1898_1) );
  OR2X2 OR2X2_1966 ( .A(w_mem_inst__abc_21378_n1895_1), .B(w_mem_inst__abc_21378_n1898_1), .Y(w_mem_inst__abc_21378_n1899_1) );
  OR2X2 OR2X2_1967 ( .A(w_mem_inst__abc_21378_n1899_1), .B(w_mem_inst__abc_21378_n1892), .Y(w_mem_inst__abc_21378_n1900) );
  OR2X2 OR2X2_1968 ( .A(w_mem_inst__abc_21378_n1900), .B(w_mem_inst__abc_21378_n1885), .Y(w_mem_inst__abc_21378_n1901) );
  OR2X2 OR2X2_1969 ( .A(w_mem_inst__abc_21378_n1901), .B(w_mem_inst__abc_21378_n1878_1), .Y(w_mem_inst__abc_21378_n1902_1) );
  OR2X2 OR2X2_197 ( .A(_abc_15724_n1299_1), .B(_abc_15724_n1297_1), .Y(_abc_15724_n1300) );
  OR2X2 OR2X2_1970 ( .A(w_mem_inst__abc_21378_n1904), .B(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_21378_n1905) );
  OR2X2 OR2X2_1971 ( .A(w_mem_inst__abc_21378_n1906_1), .B(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_21378_n1907_1) );
  OR2X2 OR2X2_1972 ( .A(w_mem_inst_w_mem_2__5_), .B(w_mem_inst_w_mem_0__5_), .Y(w_mem_inst__abc_21378_n1910_1) );
  OR2X2 OR2X2_1973 ( .A(w_mem_inst__abc_21378_n1909), .B(w_mem_inst__abc_21378_n1913), .Y(w_mem_inst__abc_21378_n1914_1) );
  OR2X2 OR2X2_1974 ( .A(w_mem_inst__abc_21378_n1915_1), .B(w_mem_inst__abc_21378_n1908), .Y(w_mem_inst__abc_21378_n1916) );
  OR2X2 OR2X2_1975 ( .A(w_mem_inst__abc_21378_n1917), .B(w_mem_inst__abc_21378_n1587_bF_buf3), .Y(w_mem_inst__abc_21378_n1918_1) );
  OR2X2 OR2X2_1976 ( .A(w_mem_inst__abc_21378_n1920), .B(w_mem_inst__abc_21378_n1586_bF_buf2), .Y(w_mem_inst__abc_21378_n1921) );
  OR2X2 OR2X2_1977 ( .A(w_mem_inst__abc_21378_n1922_1), .B(w_mem_inst__abc_21378_n1923_1), .Y(w_mem_inst__abc_21378_n1924) );
  OR2X2 OR2X2_1978 ( .A(w_mem_inst__abc_21378_n1924), .B(w_mem_inst__abc_21378_n1921), .Y(w_mem_inst__abc_21378_n1925) );
  OR2X2 OR2X2_1979 ( .A(w_mem_inst__abc_21378_n1925), .B(w_mem_inst__abc_21378_n1919_1), .Y(w_mem_inst__abc_21378_n1926_1) );
  OR2X2 OR2X2_198 ( .A(_abc_15724_n1301), .B(_abc_15724_n1286), .Y(_abc_15724_n1302) );
  OR2X2 OR2X2_1980 ( .A(w_mem_inst__abc_21378_n1927_1), .B(w_mem_inst__abc_21378_n1928), .Y(w_mem_inst__abc_21378_n1929) );
  OR2X2 OR2X2_1981 ( .A(w_mem_inst__abc_21378_n1931_1), .B(w_mem_inst__abc_21378_n1930_1), .Y(w_mem_inst__abc_21378_n1932) );
  OR2X2 OR2X2_1982 ( .A(w_mem_inst__abc_21378_n1929), .B(w_mem_inst__abc_21378_n1932), .Y(w_mem_inst__abc_21378_n1933) );
  OR2X2 OR2X2_1983 ( .A(w_mem_inst__abc_21378_n1934_1), .B(w_mem_inst__abc_21378_n1935_1), .Y(w_mem_inst__abc_21378_n1936) );
  OR2X2 OR2X2_1984 ( .A(w_mem_inst__abc_21378_n1937), .B(w_mem_inst__abc_21378_n1938_1), .Y(w_mem_inst__abc_21378_n1939_1) );
  OR2X2 OR2X2_1985 ( .A(w_mem_inst__abc_21378_n1939_1), .B(w_mem_inst__abc_21378_n1936), .Y(w_mem_inst__abc_21378_n1940) );
  OR2X2 OR2X2_1986 ( .A(w_mem_inst__abc_21378_n1942_1), .B(w_mem_inst__abc_21378_n1941), .Y(w_mem_inst__abc_21378_n1943_1) );
  OR2X2 OR2X2_1987 ( .A(w_mem_inst__abc_21378_n1944), .B(w_mem_inst__abc_21378_n1945), .Y(w_mem_inst__abc_21378_n1946_1) );
  OR2X2 OR2X2_1988 ( .A(w_mem_inst__abc_21378_n1946_1), .B(w_mem_inst__abc_21378_n1943_1), .Y(w_mem_inst__abc_21378_n1947_1) );
  OR2X2 OR2X2_1989 ( .A(w_mem_inst__abc_21378_n1940), .B(w_mem_inst__abc_21378_n1947_1), .Y(w_mem_inst__abc_21378_n1948) );
  OR2X2 OR2X2_199 ( .A(_abc_15724_n1308_1), .B(_abc_15724_n1305_1), .Y(_abc_15724_n1309) );
  OR2X2 OR2X2_1990 ( .A(w_mem_inst__abc_21378_n1948), .B(w_mem_inst__abc_21378_n1933), .Y(w_mem_inst__abc_21378_n1949) );
  OR2X2 OR2X2_1991 ( .A(w_mem_inst__abc_21378_n1949), .B(w_mem_inst__abc_21378_n1926_1), .Y(w_mem_inst__abc_21378_n1950_1) );
  OR2X2 OR2X2_1992 ( .A(w_mem_inst__abc_21378_n1952), .B(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_21378_n1953) );
  OR2X2 OR2X2_1993 ( .A(w_mem_inst__abc_21378_n1954_1), .B(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_21378_n1955_1) );
  OR2X2 OR2X2_1994 ( .A(w_mem_inst_w_mem_2__6_), .B(w_mem_inst_w_mem_0__6_), .Y(w_mem_inst__abc_21378_n1958_1) );
  OR2X2 OR2X2_1995 ( .A(w_mem_inst__abc_21378_n1957), .B(w_mem_inst__abc_21378_n1961), .Y(w_mem_inst__abc_21378_n1962_1) );
  OR2X2 OR2X2_1996 ( .A(w_mem_inst__abc_21378_n1963_1), .B(w_mem_inst__abc_21378_n1956), .Y(w_mem_inst__abc_21378_n1964) );
  OR2X2 OR2X2_1997 ( .A(w_mem_inst__abc_21378_n1965), .B(w_mem_inst__abc_21378_n1587_bF_buf2), .Y(w_mem_inst__abc_21378_n1966_1) );
  OR2X2 OR2X2_1998 ( .A(w_mem_inst__abc_21378_n1968), .B(w_mem_inst__abc_21378_n1586_bF_buf1), .Y(w_mem_inst__abc_21378_n1969) );
  OR2X2 OR2X2_1999 ( .A(w_mem_inst__abc_21378_n1970_1), .B(w_mem_inst__abc_21378_n1971_1), .Y(w_mem_inst__abc_21378_n1972) );
  OR2X2 OR2X2_2 ( .A(_abc_15724_n703), .B(_abc_15724_n698), .Y(_abc_15724_n704) );
  OR2X2 OR2X2_20 ( .A(_abc_15724_n771), .B(_abc_15724_n759), .Y(_abc_15724_n772) );
  OR2X2 OR2X2_200 ( .A(_auto_iopadmap_cc_313_execute_26059_52_), .B(d_reg_20_), .Y(_abc_15724_n1310) );
  OR2X2 OR2X2_2000 ( .A(w_mem_inst__abc_21378_n1972), .B(w_mem_inst__abc_21378_n1969), .Y(w_mem_inst__abc_21378_n1973) );
  OR2X2 OR2X2_2001 ( .A(w_mem_inst__abc_21378_n1973), .B(w_mem_inst__abc_21378_n1967_1), .Y(w_mem_inst__abc_21378_n1974_1) );
  OR2X2 OR2X2_2002 ( .A(w_mem_inst__abc_21378_n1975_1), .B(w_mem_inst__abc_21378_n1976), .Y(w_mem_inst__abc_21378_n1977) );
  OR2X2 OR2X2_2003 ( .A(w_mem_inst__abc_21378_n1979_1), .B(w_mem_inst__abc_21378_n1978_1), .Y(w_mem_inst__abc_21378_n1980) );
  OR2X2 OR2X2_2004 ( .A(w_mem_inst__abc_21378_n1977), .B(w_mem_inst__abc_21378_n1980), .Y(w_mem_inst__abc_21378_n1981) );
  OR2X2 OR2X2_2005 ( .A(w_mem_inst__abc_21378_n1982_1), .B(w_mem_inst__abc_21378_n1983_1), .Y(w_mem_inst__abc_21378_n1984) );
  OR2X2 OR2X2_2006 ( .A(w_mem_inst__abc_21378_n1985), .B(w_mem_inst__abc_21378_n1986_1), .Y(w_mem_inst__abc_21378_n1987_1) );
  OR2X2 OR2X2_2007 ( .A(w_mem_inst__abc_21378_n1984), .B(w_mem_inst__abc_21378_n1987_1), .Y(w_mem_inst__abc_21378_n1988) );
  OR2X2 OR2X2_2008 ( .A(w_mem_inst__abc_21378_n1989), .B(w_mem_inst__abc_21378_n1990_1), .Y(w_mem_inst__abc_21378_n1991_1) );
  OR2X2 OR2X2_2009 ( .A(w_mem_inst__abc_21378_n1992), .B(w_mem_inst__abc_21378_n1993), .Y(w_mem_inst__abc_21378_n1994_1) );
  OR2X2 OR2X2_201 ( .A(_abc_15724_n1309), .B(_abc_15724_n1313), .Y(_abc_15724_n1314) );
  OR2X2 OR2X2_2010 ( .A(w_mem_inst__abc_21378_n1991_1), .B(w_mem_inst__abc_21378_n1994_1), .Y(w_mem_inst__abc_21378_n1995_1) );
  OR2X2 OR2X2_2011 ( .A(w_mem_inst__abc_21378_n1995_1), .B(w_mem_inst__abc_21378_n1988), .Y(w_mem_inst__abc_21378_n1996) );
  OR2X2 OR2X2_2012 ( .A(w_mem_inst__abc_21378_n1996), .B(w_mem_inst__abc_21378_n1981), .Y(w_mem_inst__abc_21378_n1997) );
  OR2X2 OR2X2_2013 ( .A(w_mem_inst__abc_21378_n1997), .B(w_mem_inst__abc_21378_n1974_1), .Y(w_mem_inst__abc_21378_n1998_1) );
  OR2X2 OR2X2_2014 ( .A(w_mem_inst__abc_21378_n2000), .B(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_21378_n2001) );
  OR2X2 OR2X2_2015 ( .A(w_mem_inst__abc_21378_n2002_1), .B(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_21378_n2003_1) );
  OR2X2 OR2X2_2016 ( .A(w_mem_inst_w_mem_2__7_), .B(w_mem_inst_w_mem_0__7_), .Y(w_mem_inst__abc_21378_n2006_1) );
  OR2X2 OR2X2_2017 ( .A(w_mem_inst__abc_21378_n2005), .B(w_mem_inst__abc_21378_n2009), .Y(w_mem_inst__abc_21378_n2010_1) );
  OR2X2 OR2X2_2018 ( .A(w_mem_inst__abc_21378_n2011_1), .B(w_mem_inst__abc_21378_n2004), .Y(w_mem_inst__abc_21378_n2012) );
  OR2X2 OR2X2_2019 ( .A(w_mem_inst__abc_21378_n2013), .B(w_mem_inst__abc_21378_n1587_bF_buf1), .Y(w_mem_inst__abc_21378_n2014_1) );
  OR2X2 OR2X2_202 ( .A(_abc_15724_n851_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_52_), .Y(_abc_15724_n1319_1) );
  OR2X2 OR2X2_2020 ( .A(w_mem_inst__abc_21378_n2016), .B(w_mem_inst__abc_21378_n1586_bF_buf0), .Y(w_mem_inst__abc_21378_n2017) );
  OR2X2 OR2X2_2021 ( .A(w_mem_inst__abc_21378_n2018_1), .B(w_mem_inst__abc_21378_n2019_1), .Y(w_mem_inst__abc_21378_n2020) );
  OR2X2 OR2X2_2022 ( .A(w_mem_inst__abc_21378_n2020), .B(w_mem_inst__abc_21378_n2017), .Y(w_mem_inst__abc_21378_n2021) );
  OR2X2 OR2X2_2023 ( .A(w_mem_inst__abc_21378_n2021), .B(w_mem_inst__abc_21378_n2015_1), .Y(w_mem_inst__abc_21378_n2022_1) );
  OR2X2 OR2X2_2024 ( .A(w_mem_inst__abc_21378_n2023_1), .B(w_mem_inst__abc_21378_n2024), .Y(w_mem_inst__abc_21378_n2025) );
  OR2X2 OR2X2_2025 ( .A(w_mem_inst__abc_21378_n2027_1), .B(w_mem_inst__abc_21378_n2026_1), .Y(w_mem_inst__abc_21378_n2028) );
  OR2X2 OR2X2_2026 ( .A(w_mem_inst__abc_21378_n2025), .B(w_mem_inst__abc_21378_n2028), .Y(w_mem_inst__abc_21378_n2029) );
  OR2X2 OR2X2_2027 ( .A(w_mem_inst__abc_21378_n2030_1), .B(w_mem_inst__abc_21378_n2031_1), .Y(w_mem_inst__abc_21378_n2032) );
  OR2X2 OR2X2_2028 ( .A(w_mem_inst__abc_21378_n2033), .B(w_mem_inst__abc_21378_n2034_1), .Y(w_mem_inst__abc_21378_n2035_1) );
  OR2X2 OR2X2_2029 ( .A(w_mem_inst__abc_21378_n2035_1), .B(w_mem_inst__abc_21378_n2032), .Y(w_mem_inst__abc_21378_n2036) );
  OR2X2 OR2X2_203 ( .A(_abc_15724_n1318), .B(_abc_15724_n1320_1), .Y(H3_reg_20__FF_INPUT) );
  OR2X2 OR2X2_2030 ( .A(w_mem_inst__abc_21378_n2038_1), .B(w_mem_inst__abc_21378_n2037), .Y(w_mem_inst__abc_21378_n2039_1) );
  OR2X2 OR2X2_2031 ( .A(w_mem_inst__abc_21378_n2040), .B(w_mem_inst__abc_21378_n2041), .Y(w_mem_inst__abc_21378_n2042_1) );
  OR2X2 OR2X2_2032 ( .A(w_mem_inst__abc_21378_n2042_1), .B(w_mem_inst__abc_21378_n2039_1), .Y(w_mem_inst__abc_21378_n2043_1) );
  OR2X2 OR2X2_2033 ( .A(w_mem_inst__abc_21378_n2036), .B(w_mem_inst__abc_21378_n2043_1), .Y(w_mem_inst__abc_21378_n2044) );
  OR2X2 OR2X2_2034 ( .A(w_mem_inst__abc_21378_n2044), .B(w_mem_inst__abc_21378_n2029), .Y(w_mem_inst__abc_21378_n2045) );
  OR2X2 OR2X2_2035 ( .A(w_mem_inst__abc_21378_n2045), .B(w_mem_inst__abc_21378_n2022_1), .Y(w_mem_inst__abc_21378_n2046_1) );
  OR2X2 OR2X2_2036 ( .A(w_mem_inst__abc_21378_n2048), .B(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_21378_n2049) );
  OR2X2 OR2X2_2037 ( .A(w_mem_inst__abc_21378_n2050_1), .B(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_21378_n2051_1) );
  OR2X2 OR2X2_2038 ( .A(w_mem_inst_w_mem_2__8_), .B(w_mem_inst_w_mem_0__8_), .Y(w_mem_inst__abc_21378_n2054_1) );
  OR2X2 OR2X2_2039 ( .A(w_mem_inst__abc_21378_n2053), .B(w_mem_inst__abc_21378_n2057), .Y(w_mem_inst__abc_21378_n2058_1) );
  OR2X2 OR2X2_204 ( .A(_auto_iopadmap_cc_313_execute_26059_53_), .B(d_reg_21_), .Y(_abc_15724_n1323) );
  OR2X2 OR2X2_2040 ( .A(w_mem_inst__abc_21378_n2059_1), .B(w_mem_inst__abc_21378_n2052), .Y(w_mem_inst__abc_21378_n2060) );
  OR2X2 OR2X2_2041 ( .A(w_mem_inst__abc_21378_n2061), .B(w_mem_inst__abc_21378_n1587_bF_buf0), .Y(w_mem_inst__abc_21378_n2062_1) );
  OR2X2 OR2X2_2042 ( .A(w_mem_inst__abc_21378_n2064), .B(w_mem_inst__abc_21378_n1586_bF_buf4), .Y(w_mem_inst__abc_21378_n2065) );
  OR2X2 OR2X2_2043 ( .A(w_mem_inst__abc_21378_n2066_1), .B(w_mem_inst__abc_21378_n2067_1), .Y(w_mem_inst__abc_21378_n2068) );
  OR2X2 OR2X2_2044 ( .A(w_mem_inst__abc_21378_n2068), .B(w_mem_inst__abc_21378_n2065), .Y(w_mem_inst__abc_21378_n2069) );
  OR2X2 OR2X2_2045 ( .A(w_mem_inst__abc_21378_n2069), .B(w_mem_inst__abc_21378_n2063_1), .Y(w_mem_inst__abc_21378_n2070_1) );
  OR2X2 OR2X2_2046 ( .A(w_mem_inst__abc_21378_n2071_1), .B(w_mem_inst__abc_21378_n2072), .Y(w_mem_inst__abc_21378_n2073) );
  OR2X2 OR2X2_2047 ( .A(w_mem_inst__abc_21378_n2075_1), .B(w_mem_inst__abc_21378_n2074_1), .Y(w_mem_inst__abc_21378_n2076) );
  OR2X2 OR2X2_2048 ( .A(w_mem_inst__abc_21378_n2073), .B(w_mem_inst__abc_21378_n2076), .Y(w_mem_inst__abc_21378_n2077) );
  OR2X2 OR2X2_2049 ( .A(w_mem_inst__abc_21378_n2078_1), .B(w_mem_inst__abc_21378_n2079_1), .Y(w_mem_inst__abc_21378_n2080) );
  OR2X2 OR2X2_205 ( .A(_abc_15724_n1330_1), .B(_abc_15724_n1327), .Y(_abc_15724_n1331) );
  OR2X2 OR2X2_2050 ( .A(w_mem_inst__abc_21378_n2081), .B(w_mem_inst__abc_21378_n2082_1), .Y(w_mem_inst__abc_21378_n2083_1) );
  OR2X2 OR2X2_2051 ( .A(w_mem_inst__abc_21378_n2080), .B(w_mem_inst__abc_21378_n2083_1), .Y(w_mem_inst__abc_21378_n2084) );
  OR2X2 OR2X2_2052 ( .A(w_mem_inst__abc_21378_n2085), .B(w_mem_inst__abc_21378_n2086_1), .Y(w_mem_inst__abc_21378_n2087_1) );
  OR2X2 OR2X2_2053 ( .A(w_mem_inst__abc_21378_n2088), .B(w_mem_inst__abc_21378_n2089), .Y(w_mem_inst__abc_21378_n2090_1) );
  OR2X2 OR2X2_2054 ( .A(w_mem_inst__abc_21378_n2087_1), .B(w_mem_inst__abc_21378_n2090_1), .Y(w_mem_inst__abc_21378_n2091_1) );
  OR2X2 OR2X2_2055 ( .A(w_mem_inst__abc_21378_n2091_1), .B(w_mem_inst__abc_21378_n2084), .Y(w_mem_inst__abc_21378_n2092) );
  OR2X2 OR2X2_2056 ( .A(w_mem_inst__abc_21378_n2092), .B(w_mem_inst__abc_21378_n2077), .Y(w_mem_inst__abc_21378_n2093) );
  OR2X2 OR2X2_2057 ( .A(w_mem_inst__abc_21378_n2093), .B(w_mem_inst__abc_21378_n2070_1), .Y(w_mem_inst__abc_21378_n2094_1) );
  OR2X2 OR2X2_2058 ( .A(w_mem_inst__abc_21378_n2096), .B(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_21378_n2097) );
  OR2X2 OR2X2_2059 ( .A(w_mem_inst__abc_21378_n2098_1), .B(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_21378_n2099_1) );
  OR2X2 OR2X2_206 ( .A(_abc_15724_n851_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_53_), .Y(_abc_15724_n1333) );
  OR2X2 OR2X2_2060 ( .A(w_mem_inst_w_mem_2__9_), .B(w_mem_inst_w_mem_0__9_), .Y(w_mem_inst__abc_21378_n2102_1) );
  OR2X2 OR2X2_2061 ( .A(w_mem_inst__abc_21378_n2101), .B(w_mem_inst__abc_21378_n2105), .Y(w_mem_inst__abc_21378_n2106_1) );
  OR2X2 OR2X2_2062 ( .A(w_mem_inst__abc_21378_n2107_1), .B(w_mem_inst__abc_21378_n2100), .Y(w_mem_inst__abc_21378_n2108) );
  OR2X2 OR2X2_2063 ( .A(w_mem_inst__abc_21378_n2109), .B(w_mem_inst__abc_21378_n1587_bF_buf4), .Y(w_mem_inst__abc_21378_n2110_1) );
  OR2X2 OR2X2_2064 ( .A(w_mem_inst__abc_21378_n2112), .B(w_mem_inst__abc_21378_n1586_bF_buf3), .Y(w_mem_inst__abc_21378_n2113) );
  OR2X2 OR2X2_2065 ( .A(w_mem_inst__abc_21378_n2114_1), .B(w_mem_inst__abc_21378_n2115_1), .Y(w_mem_inst__abc_21378_n2116) );
  OR2X2 OR2X2_2066 ( .A(w_mem_inst__abc_21378_n2116), .B(w_mem_inst__abc_21378_n2113), .Y(w_mem_inst__abc_21378_n2117) );
  OR2X2 OR2X2_2067 ( .A(w_mem_inst__abc_21378_n2117), .B(w_mem_inst__abc_21378_n2111_1), .Y(w_mem_inst__abc_21378_n2118_1) );
  OR2X2 OR2X2_2068 ( .A(w_mem_inst__abc_21378_n2119_1), .B(w_mem_inst__abc_21378_n2120), .Y(w_mem_inst__abc_21378_n2121) );
  OR2X2 OR2X2_2069 ( .A(w_mem_inst__abc_21378_n2123_1), .B(w_mem_inst__abc_21378_n2122_1), .Y(w_mem_inst__abc_21378_n2124) );
  OR2X2 OR2X2_207 ( .A(_abc_15724_n1332_1), .B(_abc_15724_n1334), .Y(H3_reg_21__FF_INPUT) );
  OR2X2 OR2X2_2070 ( .A(w_mem_inst__abc_21378_n2121), .B(w_mem_inst__abc_21378_n2124), .Y(w_mem_inst__abc_21378_n2125) );
  OR2X2 OR2X2_2071 ( .A(w_mem_inst__abc_21378_n2126_1), .B(w_mem_inst__abc_21378_n2127_1), .Y(w_mem_inst__abc_21378_n2128) );
  OR2X2 OR2X2_2072 ( .A(w_mem_inst__abc_21378_n2129), .B(w_mem_inst__abc_21378_n2130_1), .Y(w_mem_inst__abc_21378_n2131_1) );
  OR2X2 OR2X2_2073 ( .A(w_mem_inst__abc_21378_n2131_1), .B(w_mem_inst__abc_21378_n2128), .Y(w_mem_inst__abc_21378_n2132) );
  OR2X2 OR2X2_2074 ( .A(w_mem_inst__abc_21378_n2134_1), .B(w_mem_inst__abc_21378_n2133), .Y(w_mem_inst__abc_21378_n2135_1) );
  OR2X2 OR2X2_2075 ( .A(w_mem_inst__abc_21378_n2136), .B(w_mem_inst__abc_21378_n2137), .Y(w_mem_inst__abc_21378_n2138_1) );
  OR2X2 OR2X2_2076 ( .A(w_mem_inst__abc_21378_n2138_1), .B(w_mem_inst__abc_21378_n2135_1), .Y(w_mem_inst__abc_21378_n2139_1) );
  OR2X2 OR2X2_2077 ( .A(w_mem_inst__abc_21378_n2132), .B(w_mem_inst__abc_21378_n2139_1), .Y(w_mem_inst__abc_21378_n2140) );
  OR2X2 OR2X2_2078 ( .A(w_mem_inst__abc_21378_n2140), .B(w_mem_inst__abc_21378_n2125), .Y(w_mem_inst__abc_21378_n2141) );
  OR2X2 OR2X2_2079 ( .A(w_mem_inst__abc_21378_n2141), .B(w_mem_inst__abc_21378_n2118_1), .Y(w_mem_inst__abc_21378_n2142_1) );
  OR2X2 OR2X2_208 ( .A(_auto_iopadmap_cc_313_execute_26059_54_), .B(d_reg_22_), .Y(_abc_15724_n1337) );
  OR2X2 OR2X2_2080 ( .A(w_mem_inst__abc_21378_n2144), .B(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_21378_n2145) );
  OR2X2 OR2X2_2081 ( .A(w_mem_inst__abc_21378_n2146_1), .B(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_21378_n2147_1) );
  OR2X2 OR2X2_2082 ( .A(w_mem_inst_w_mem_2__10_), .B(w_mem_inst_w_mem_0__10_), .Y(w_mem_inst__abc_21378_n2150_1) );
  OR2X2 OR2X2_2083 ( .A(w_mem_inst__abc_21378_n2149), .B(w_mem_inst__abc_21378_n2153), .Y(w_mem_inst__abc_21378_n2154_1) );
  OR2X2 OR2X2_2084 ( .A(w_mem_inst__abc_21378_n2155_1), .B(w_mem_inst__abc_21378_n2148), .Y(w_mem_inst__abc_21378_n2156) );
  OR2X2 OR2X2_2085 ( .A(w_mem_inst__abc_21378_n2157), .B(w_mem_inst__abc_21378_n1587_bF_buf3), .Y(w_mem_inst__abc_21378_n2158_1) );
  OR2X2 OR2X2_2086 ( .A(w_mem_inst__abc_21378_n2160), .B(w_mem_inst__abc_21378_n1586_bF_buf2), .Y(w_mem_inst__abc_21378_n2161) );
  OR2X2 OR2X2_2087 ( .A(w_mem_inst__abc_21378_n2162_1), .B(w_mem_inst__abc_21378_n2163_1), .Y(w_mem_inst__abc_21378_n2164) );
  OR2X2 OR2X2_2088 ( .A(w_mem_inst__abc_21378_n2164), .B(w_mem_inst__abc_21378_n2161), .Y(w_mem_inst__abc_21378_n2165) );
  OR2X2 OR2X2_2089 ( .A(w_mem_inst__abc_21378_n2165), .B(w_mem_inst__abc_21378_n2159_1), .Y(w_mem_inst__abc_21378_n2166_1) );
  OR2X2 OR2X2_209 ( .A(_abc_15724_n1343_1), .B(_abc_15724_n1341_1), .Y(_abc_15724_n1344) );
  OR2X2 OR2X2_2090 ( .A(w_mem_inst__abc_21378_n2167_1), .B(w_mem_inst__abc_21378_n2168), .Y(w_mem_inst__abc_21378_n2169) );
  OR2X2 OR2X2_2091 ( .A(w_mem_inst__abc_21378_n2171_1), .B(w_mem_inst__abc_21378_n2170_1), .Y(w_mem_inst__abc_21378_n2172) );
  OR2X2 OR2X2_2092 ( .A(w_mem_inst__abc_21378_n2169), .B(w_mem_inst__abc_21378_n2172), .Y(w_mem_inst__abc_21378_n2173) );
  OR2X2 OR2X2_2093 ( .A(w_mem_inst__abc_21378_n2174_1), .B(w_mem_inst__abc_21378_n2175_1), .Y(w_mem_inst__abc_21378_n2176) );
  OR2X2 OR2X2_2094 ( .A(w_mem_inst__abc_21378_n2177), .B(w_mem_inst__abc_21378_n2178_1), .Y(w_mem_inst__abc_21378_n2179_1) );
  OR2X2 OR2X2_2095 ( .A(w_mem_inst__abc_21378_n2176), .B(w_mem_inst__abc_21378_n2179_1), .Y(w_mem_inst__abc_21378_n2180) );
  OR2X2 OR2X2_2096 ( .A(w_mem_inst__abc_21378_n2181), .B(w_mem_inst__abc_21378_n2182_1), .Y(w_mem_inst__abc_21378_n2183_1) );
  OR2X2 OR2X2_2097 ( .A(w_mem_inst__abc_21378_n2184), .B(w_mem_inst__abc_21378_n2185), .Y(w_mem_inst__abc_21378_n2186_1) );
  OR2X2 OR2X2_2098 ( .A(w_mem_inst__abc_21378_n2183_1), .B(w_mem_inst__abc_21378_n2186_1), .Y(w_mem_inst__abc_21378_n2187_1) );
  OR2X2 OR2X2_2099 ( .A(w_mem_inst__abc_21378_n2187_1), .B(w_mem_inst__abc_21378_n2180), .Y(w_mem_inst__abc_21378_n2188) );
  OR2X2 OR2X2_21 ( .A(_auto_iopadmap_cc_313_execute_26059_7_), .B(e_reg_7_), .Y(_abc_15724_n774) );
  OR2X2 OR2X2_210 ( .A(_abc_15724_n1345), .B(_abc_15724_n1340_1), .Y(_abc_15724_n1348) );
  OR2X2 OR2X2_2100 ( .A(w_mem_inst__abc_21378_n2188), .B(w_mem_inst__abc_21378_n2173), .Y(w_mem_inst__abc_21378_n2189) );
  OR2X2 OR2X2_2101 ( .A(w_mem_inst__abc_21378_n2189), .B(w_mem_inst__abc_21378_n2166_1), .Y(w_mem_inst__abc_21378_n2190_1) );
  OR2X2 OR2X2_2102 ( .A(w_mem_inst__abc_21378_n2192), .B(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_21378_n2193) );
  OR2X2 OR2X2_2103 ( .A(w_mem_inst__abc_21378_n2194_1), .B(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_21378_n2195_1) );
  OR2X2 OR2X2_2104 ( .A(w_mem_inst_w_mem_2__11_), .B(w_mem_inst_w_mem_0__11_), .Y(w_mem_inst__abc_21378_n2198_1) );
  OR2X2 OR2X2_2105 ( .A(w_mem_inst__abc_21378_n2197), .B(w_mem_inst__abc_21378_n2201), .Y(w_mem_inst__abc_21378_n2202_1) );
  OR2X2 OR2X2_2106 ( .A(w_mem_inst__abc_21378_n2203_1), .B(w_mem_inst__abc_21378_n2196), .Y(w_mem_inst__abc_21378_n2204) );
  OR2X2 OR2X2_2107 ( .A(w_mem_inst__abc_21378_n2205), .B(w_mem_inst__abc_21378_n1587_bF_buf2), .Y(w_mem_inst__abc_21378_n2206_1) );
  OR2X2 OR2X2_2108 ( .A(w_mem_inst__abc_21378_n2208), .B(w_mem_inst__abc_21378_n1586_bF_buf1), .Y(w_mem_inst__abc_21378_n2209) );
  OR2X2 OR2X2_2109 ( .A(w_mem_inst__abc_21378_n2210_1), .B(w_mem_inst__abc_21378_n2211_1), .Y(w_mem_inst__abc_21378_n2212) );
  OR2X2 OR2X2_211 ( .A(_abc_15724_n1350_1), .B(_abc_15724_n1336), .Y(H3_reg_22__FF_INPUT) );
  OR2X2 OR2X2_2110 ( .A(w_mem_inst__abc_21378_n2212), .B(w_mem_inst__abc_21378_n2209), .Y(w_mem_inst__abc_21378_n2213) );
  OR2X2 OR2X2_2111 ( .A(w_mem_inst__abc_21378_n2213), .B(w_mem_inst__abc_21378_n2207_1), .Y(w_mem_inst__abc_21378_n2214_1) );
  OR2X2 OR2X2_2112 ( .A(w_mem_inst__abc_21378_n2215_1), .B(w_mem_inst__abc_21378_n2216), .Y(w_mem_inst__abc_21378_n2217) );
  OR2X2 OR2X2_2113 ( .A(w_mem_inst__abc_21378_n2219_1), .B(w_mem_inst__abc_21378_n2218_1), .Y(w_mem_inst__abc_21378_n2220) );
  OR2X2 OR2X2_2114 ( .A(w_mem_inst__abc_21378_n2217), .B(w_mem_inst__abc_21378_n2220), .Y(w_mem_inst__abc_21378_n2221) );
  OR2X2 OR2X2_2115 ( .A(w_mem_inst__abc_21378_n2222_1), .B(w_mem_inst__abc_21378_n2223_1), .Y(w_mem_inst__abc_21378_n2224) );
  OR2X2 OR2X2_2116 ( .A(w_mem_inst__abc_21378_n2225), .B(w_mem_inst__abc_21378_n2226_1), .Y(w_mem_inst__abc_21378_n2227_1) );
  OR2X2 OR2X2_2117 ( .A(w_mem_inst__abc_21378_n2227_1), .B(w_mem_inst__abc_21378_n2224), .Y(w_mem_inst__abc_21378_n2228) );
  OR2X2 OR2X2_2118 ( .A(w_mem_inst__abc_21378_n2230_1), .B(w_mem_inst__abc_21378_n2229), .Y(w_mem_inst__abc_21378_n2231_1) );
  OR2X2 OR2X2_2119 ( .A(w_mem_inst__abc_21378_n2232), .B(w_mem_inst__abc_21378_n2233), .Y(w_mem_inst__abc_21378_n2234_1) );
  OR2X2 OR2X2_212 ( .A(_auto_iopadmap_cc_313_execute_26059_55_), .B(d_reg_23_), .Y(_abc_15724_n1353) );
  OR2X2 OR2X2_2120 ( .A(w_mem_inst__abc_21378_n2234_1), .B(w_mem_inst__abc_21378_n2231_1), .Y(w_mem_inst__abc_21378_n2235_1) );
  OR2X2 OR2X2_2121 ( .A(w_mem_inst__abc_21378_n2228), .B(w_mem_inst__abc_21378_n2235_1), .Y(w_mem_inst__abc_21378_n2236) );
  OR2X2 OR2X2_2122 ( .A(w_mem_inst__abc_21378_n2236), .B(w_mem_inst__abc_21378_n2221), .Y(w_mem_inst__abc_21378_n2237) );
  OR2X2 OR2X2_2123 ( .A(w_mem_inst__abc_21378_n2237), .B(w_mem_inst__abc_21378_n2214_1), .Y(w_mem_inst__abc_21378_n2238_1) );
  OR2X2 OR2X2_2124 ( .A(w_mem_inst__abc_21378_n2240), .B(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_21378_n2241) );
  OR2X2 OR2X2_2125 ( .A(w_mem_inst__abc_21378_n2242_1), .B(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_21378_n2243_1) );
  OR2X2 OR2X2_2126 ( .A(w_mem_inst_w_mem_2__12_), .B(w_mem_inst_w_mem_0__12_), .Y(w_mem_inst__abc_21378_n2246_1) );
  OR2X2 OR2X2_2127 ( .A(w_mem_inst__abc_21378_n2245), .B(w_mem_inst__abc_21378_n2249), .Y(w_mem_inst__abc_21378_n2250_1) );
  OR2X2 OR2X2_2128 ( .A(w_mem_inst__abc_21378_n2251_1), .B(w_mem_inst__abc_21378_n2244), .Y(w_mem_inst__abc_21378_n2252) );
  OR2X2 OR2X2_2129 ( .A(w_mem_inst__abc_21378_n2253), .B(w_mem_inst__abc_21378_n1587_bF_buf1), .Y(w_mem_inst__abc_21378_n2254_1) );
  OR2X2 OR2X2_213 ( .A(_abc_15724_n1352_1), .B(_abc_15724_n1357), .Y(_abc_15724_n1358) );
  OR2X2 OR2X2_2130 ( .A(w_mem_inst__abc_21378_n2256), .B(w_mem_inst__abc_21378_n1586_bF_buf0), .Y(w_mem_inst__abc_21378_n2257) );
  OR2X2 OR2X2_2131 ( .A(w_mem_inst__abc_21378_n2258_1), .B(w_mem_inst__abc_21378_n2259_1), .Y(w_mem_inst__abc_21378_n2260) );
  OR2X2 OR2X2_2132 ( .A(w_mem_inst__abc_21378_n2260), .B(w_mem_inst__abc_21378_n2257), .Y(w_mem_inst__abc_21378_n2261) );
  OR2X2 OR2X2_2133 ( .A(w_mem_inst__abc_21378_n2261), .B(w_mem_inst__abc_21378_n2255_1), .Y(w_mem_inst__abc_21378_n2262_1) );
  OR2X2 OR2X2_2134 ( .A(w_mem_inst__abc_21378_n2263_1), .B(w_mem_inst__abc_21378_n2264), .Y(w_mem_inst__abc_21378_n2265) );
  OR2X2 OR2X2_2135 ( .A(w_mem_inst__abc_21378_n2267_1), .B(w_mem_inst__abc_21378_n2266_1), .Y(w_mem_inst__abc_21378_n2268) );
  OR2X2 OR2X2_2136 ( .A(w_mem_inst__abc_21378_n2265), .B(w_mem_inst__abc_21378_n2268), .Y(w_mem_inst__abc_21378_n2269) );
  OR2X2 OR2X2_2137 ( .A(w_mem_inst__abc_21378_n2270_1), .B(w_mem_inst__abc_21378_n2271_1), .Y(w_mem_inst__abc_21378_n2272) );
  OR2X2 OR2X2_2138 ( .A(w_mem_inst__abc_21378_n2273), .B(w_mem_inst__abc_21378_n2274_1), .Y(w_mem_inst__abc_21378_n2275_1) );
  OR2X2 OR2X2_2139 ( .A(w_mem_inst__abc_21378_n2272), .B(w_mem_inst__abc_21378_n2275_1), .Y(w_mem_inst__abc_21378_n2276) );
  OR2X2 OR2X2_214 ( .A(_abc_15724_n1359), .B(_abc_15724_n1356), .Y(_abc_15724_n1360) );
  OR2X2 OR2X2_2140 ( .A(w_mem_inst__abc_21378_n2277), .B(w_mem_inst__abc_21378_n2278_1), .Y(w_mem_inst__abc_21378_n2279_1) );
  OR2X2 OR2X2_2141 ( .A(w_mem_inst__abc_21378_n2280), .B(w_mem_inst__abc_21378_n2281), .Y(w_mem_inst__abc_21378_n2282_1) );
  OR2X2 OR2X2_2142 ( .A(w_mem_inst__abc_21378_n2279_1), .B(w_mem_inst__abc_21378_n2282_1), .Y(w_mem_inst__abc_21378_n2283_1) );
  OR2X2 OR2X2_2143 ( .A(w_mem_inst__abc_21378_n2283_1), .B(w_mem_inst__abc_21378_n2276), .Y(w_mem_inst__abc_21378_n2284) );
  OR2X2 OR2X2_2144 ( .A(w_mem_inst__abc_21378_n2284), .B(w_mem_inst__abc_21378_n2269), .Y(w_mem_inst__abc_21378_n2285) );
  OR2X2 OR2X2_2145 ( .A(w_mem_inst__abc_21378_n2285), .B(w_mem_inst__abc_21378_n2262_1), .Y(w_mem_inst__abc_21378_n2286_1) );
  OR2X2 OR2X2_2146 ( .A(w_mem_inst__abc_21378_n2288), .B(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_21378_n2289) );
  OR2X2 OR2X2_2147 ( .A(w_mem_inst__abc_21378_n2290_1), .B(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_21378_n2291_1) );
  OR2X2 OR2X2_2148 ( .A(w_mem_inst_w_mem_2__13_), .B(w_mem_inst_w_mem_0__13_), .Y(w_mem_inst__abc_21378_n2294_1) );
  OR2X2 OR2X2_2149 ( .A(w_mem_inst__abc_21378_n2293), .B(w_mem_inst__abc_21378_n2297), .Y(w_mem_inst__abc_21378_n2298_1) );
  OR2X2 OR2X2_215 ( .A(_abc_15724_n1362), .B(_abc_15724_n1363), .Y(H3_reg_23__FF_INPUT) );
  OR2X2 OR2X2_2150 ( .A(w_mem_inst__abc_21378_n2299_1), .B(w_mem_inst__abc_21378_n2292), .Y(w_mem_inst__abc_21378_n2300) );
  OR2X2 OR2X2_2151 ( .A(w_mem_inst__abc_21378_n2301), .B(w_mem_inst__abc_21378_n1587_bF_buf0), .Y(w_mem_inst__abc_21378_n2302_1) );
  OR2X2 OR2X2_2152 ( .A(w_mem_inst__abc_21378_n2304), .B(w_mem_inst__abc_21378_n1586_bF_buf4), .Y(w_mem_inst__abc_21378_n2305) );
  OR2X2 OR2X2_2153 ( .A(w_mem_inst__abc_21378_n2306_1), .B(w_mem_inst__abc_21378_n2307_1), .Y(w_mem_inst__abc_21378_n2308) );
  OR2X2 OR2X2_2154 ( .A(w_mem_inst__abc_21378_n2308), .B(w_mem_inst__abc_21378_n2305), .Y(w_mem_inst__abc_21378_n2309) );
  OR2X2 OR2X2_2155 ( .A(w_mem_inst__abc_21378_n2309), .B(w_mem_inst__abc_21378_n2303_1), .Y(w_mem_inst__abc_21378_n2310_1) );
  OR2X2 OR2X2_2156 ( .A(w_mem_inst__abc_21378_n2311_1), .B(w_mem_inst__abc_21378_n2312), .Y(w_mem_inst__abc_21378_n2313) );
  OR2X2 OR2X2_2157 ( .A(w_mem_inst__abc_21378_n2315_1), .B(w_mem_inst__abc_21378_n2314_1), .Y(w_mem_inst__abc_21378_n2316) );
  OR2X2 OR2X2_2158 ( .A(w_mem_inst__abc_21378_n2313), .B(w_mem_inst__abc_21378_n2316), .Y(w_mem_inst__abc_21378_n2317) );
  OR2X2 OR2X2_2159 ( .A(w_mem_inst__abc_21378_n2318_1), .B(w_mem_inst__abc_21378_n2319_1), .Y(w_mem_inst__abc_21378_n2320) );
  OR2X2 OR2X2_216 ( .A(_abc_15724_n1342), .B(_abc_15724_n1341_1), .Y(_abc_15724_n1370) );
  OR2X2 OR2X2_2160 ( .A(w_mem_inst__abc_21378_n2321), .B(w_mem_inst__abc_21378_n2322_1), .Y(w_mem_inst__abc_21378_n2323_1) );
  OR2X2 OR2X2_2161 ( .A(w_mem_inst__abc_21378_n2323_1), .B(w_mem_inst__abc_21378_n2320), .Y(w_mem_inst__abc_21378_n2324) );
  OR2X2 OR2X2_2162 ( .A(w_mem_inst__abc_21378_n2326_1), .B(w_mem_inst__abc_21378_n2325), .Y(w_mem_inst__abc_21378_n2327_1) );
  OR2X2 OR2X2_2163 ( .A(w_mem_inst__abc_21378_n2328), .B(w_mem_inst__abc_21378_n2329), .Y(w_mem_inst__abc_21378_n2330_1) );
  OR2X2 OR2X2_2164 ( .A(w_mem_inst__abc_21378_n2330_1), .B(w_mem_inst__abc_21378_n2327_1), .Y(w_mem_inst__abc_21378_n2331_1) );
  OR2X2 OR2X2_2165 ( .A(w_mem_inst__abc_21378_n2324), .B(w_mem_inst__abc_21378_n2331_1), .Y(w_mem_inst__abc_21378_n2332) );
  OR2X2 OR2X2_2166 ( .A(w_mem_inst__abc_21378_n2332), .B(w_mem_inst__abc_21378_n2317), .Y(w_mem_inst__abc_21378_n2333) );
  OR2X2 OR2X2_2167 ( .A(w_mem_inst__abc_21378_n2333), .B(w_mem_inst__abc_21378_n2310_1), .Y(w_mem_inst__abc_21378_n2334_1) );
  OR2X2 OR2X2_2168 ( .A(w_mem_inst__abc_21378_n2336), .B(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_21378_n2337) );
  OR2X2 OR2X2_2169 ( .A(w_mem_inst__abc_21378_n2338_1), .B(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_21378_n2339_1) );
  OR2X2 OR2X2_217 ( .A(_abc_15724_n1373), .B(_abc_15724_n1354), .Y(_abc_15724_n1374) );
  OR2X2 OR2X2_2170 ( .A(w_mem_inst_w_mem_2__14_), .B(w_mem_inst_w_mem_0__14_), .Y(w_mem_inst__abc_21378_n2342_1) );
  OR2X2 OR2X2_2171 ( .A(w_mem_inst__abc_21378_n2341), .B(w_mem_inst__abc_21378_n2345), .Y(w_mem_inst__abc_21378_n2346_1) );
  OR2X2 OR2X2_2172 ( .A(w_mem_inst__abc_21378_n2347_1), .B(w_mem_inst__abc_21378_n2340), .Y(w_mem_inst__abc_21378_n2348) );
  OR2X2 OR2X2_2173 ( .A(w_mem_inst__abc_21378_n2349), .B(w_mem_inst__abc_21378_n1587_bF_buf4), .Y(w_mem_inst__abc_21378_n2350_1) );
  OR2X2 OR2X2_2174 ( .A(w_mem_inst__abc_21378_n2352), .B(w_mem_inst__abc_21378_n1586_bF_buf3), .Y(w_mem_inst__abc_21378_n2353) );
  OR2X2 OR2X2_2175 ( .A(w_mem_inst__abc_21378_n2354_1), .B(w_mem_inst__abc_21378_n2355_1), .Y(w_mem_inst__abc_21378_n2356) );
  OR2X2 OR2X2_2176 ( .A(w_mem_inst__abc_21378_n2356), .B(w_mem_inst__abc_21378_n2353), .Y(w_mem_inst__abc_21378_n2357) );
  OR2X2 OR2X2_2177 ( .A(w_mem_inst__abc_21378_n2357), .B(w_mem_inst__abc_21378_n2351_1), .Y(w_mem_inst__abc_21378_n2358_1) );
  OR2X2 OR2X2_2178 ( .A(w_mem_inst__abc_21378_n2359_1), .B(w_mem_inst__abc_21378_n2360), .Y(w_mem_inst__abc_21378_n2361) );
  OR2X2 OR2X2_2179 ( .A(w_mem_inst__abc_21378_n2363_1), .B(w_mem_inst__abc_21378_n2362_1), .Y(w_mem_inst__abc_21378_n2364) );
  OR2X2 OR2X2_218 ( .A(_abc_15724_n1372), .B(_abc_15724_n1374), .Y(_abc_15724_n1375) );
  OR2X2 OR2X2_2180 ( .A(w_mem_inst__abc_21378_n2361), .B(w_mem_inst__abc_21378_n2364), .Y(w_mem_inst__abc_21378_n2365) );
  OR2X2 OR2X2_2181 ( .A(w_mem_inst__abc_21378_n2366_1), .B(w_mem_inst__abc_21378_n2367_1), .Y(w_mem_inst__abc_21378_n2368) );
  OR2X2 OR2X2_2182 ( .A(w_mem_inst__abc_21378_n2369), .B(w_mem_inst__abc_21378_n2370_1), .Y(w_mem_inst__abc_21378_n2371_1) );
  OR2X2 OR2X2_2183 ( .A(w_mem_inst__abc_21378_n2368), .B(w_mem_inst__abc_21378_n2371_1), .Y(w_mem_inst__abc_21378_n2372) );
  OR2X2 OR2X2_2184 ( .A(w_mem_inst__abc_21378_n2373), .B(w_mem_inst__abc_21378_n2374_1), .Y(w_mem_inst__abc_21378_n2375_1) );
  OR2X2 OR2X2_2185 ( .A(w_mem_inst__abc_21378_n2376), .B(w_mem_inst__abc_21378_n2377), .Y(w_mem_inst__abc_21378_n2378_1) );
  OR2X2 OR2X2_2186 ( .A(w_mem_inst__abc_21378_n2375_1), .B(w_mem_inst__abc_21378_n2378_1), .Y(w_mem_inst__abc_21378_n2379_1) );
  OR2X2 OR2X2_2187 ( .A(w_mem_inst__abc_21378_n2379_1), .B(w_mem_inst__abc_21378_n2372), .Y(w_mem_inst__abc_21378_n2380) );
  OR2X2 OR2X2_2188 ( .A(w_mem_inst__abc_21378_n2380), .B(w_mem_inst__abc_21378_n2365), .Y(w_mem_inst__abc_21378_n2381) );
  OR2X2 OR2X2_2189 ( .A(w_mem_inst__abc_21378_n2381), .B(w_mem_inst__abc_21378_n2358_1), .Y(w_mem_inst__abc_21378_n2382_1) );
  OR2X2 OR2X2_219 ( .A(_abc_15724_n1369_1), .B(_abc_15724_n1375), .Y(_abc_15724_n1376) );
  OR2X2 OR2X2_2190 ( .A(w_mem_inst__abc_21378_n2384), .B(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_21378_n2385) );
  OR2X2 OR2X2_2191 ( .A(w_mem_inst__abc_21378_n2386_1), .B(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_21378_n2387_1) );
  OR2X2 OR2X2_2192 ( .A(w_mem_inst_w_mem_2__15_), .B(w_mem_inst_w_mem_0__15_), .Y(w_mem_inst__abc_21378_n2390_1) );
  OR2X2 OR2X2_2193 ( .A(w_mem_inst__abc_21378_n2389), .B(w_mem_inst__abc_21378_n2393), .Y(w_mem_inst__abc_21378_n2394_1) );
  OR2X2 OR2X2_2194 ( .A(w_mem_inst__abc_21378_n2395_1), .B(w_mem_inst__abc_21378_n2388), .Y(w_mem_inst__abc_21378_n2396) );
  OR2X2 OR2X2_2195 ( .A(w_mem_inst__abc_21378_n2397), .B(w_mem_inst__abc_21378_n1587_bF_buf3), .Y(w_mem_inst__abc_21378_n2398_1) );
  OR2X2 OR2X2_2196 ( .A(w_mem_inst__abc_21378_n2400), .B(w_mem_inst__abc_21378_n1586_bF_buf2), .Y(w_mem_inst__abc_21378_n2401) );
  OR2X2 OR2X2_2197 ( .A(w_mem_inst__abc_21378_n2402_1), .B(w_mem_inst__abc_21378_n2403_1), .Y(w_mem_inst__abc_21378_n2404) );
  OR2X2 OR2X2_2198 ( .A(w_mem_inst__abc_21378_n2404), .B(w_mem_inst__abc_21378_n2401), .Y(w_mem_inst__abc_21378_n2405) );
  OR2X2 OR2X2_2199 ( .A(w_mem_inst__abc_21378_n2405), .B(w_mem_inst__abc_21378_n2399_1), .Y(w_mem_inst__abc_21378_n2406_1) );
  OR2X2 OR2X2_22 ( .A(_abc_15724_n776), .B(_abc_15724_n773), .Y(_abc_15724_n777) );
  OR2X2 OR2X2_220 ( .A(_abc_15724_n1378_1), .B(_abc_15724_n1376), .Y(_abc_15724_n1379_1) );
  OR2X2 OR2X2_2200 ( .A(w_mem_inst__abc_21378_n2407_1), .B(w_mem_inst__abc_21378_n2408), .Y(w_mem_inst__abc_21378_n2409) );
  OR2X2 OR2X2_2201 ( .A(w_mem_inst__abc_21378_n2411_1), .B(w_mem_inst__abc_21378_n2410_1), .Y(w_mem_inst__abc_21378_n2412) );
  OR2X2 OR2X2_2202 ( .A(w_mem_inst__abc_21378_n2409), .B(w_mem_inst__abc_21378_n2412), .Y(w_mem_inst__abc_21378_n2413) );
  OR2X2 OR2X2_2203 ( .A(w_mem_inst__abc_21378_n2414_1), .B(w_mem_inst__abc_21378_n2415_1), .Y(w_mem_inst__abc_21378_n2416) );
  OR2X2 OR2X2_2204 ( .A(w_mem_inst__abc_21378_n2417), .B(w_mem_inst__abc_21378_n2418_1), .Y(w_mem_inst__abc_21378_n2419_1) );
  OR2X2 OR2X2_2205 ( .A(w_mem_inst__abc_21378_n2419_1), .B(w_mem_inst__abc_21378_n2416), .Y(w_mem_inst__abc_21378_n2420) );
  OR2X2 OR2X2_2206 ( .A(w_mem_inst__abc_21378_n2422_1), .B(w_mem_inst__abc_21378_n2421), .Y(w_mem_inst__abc_21378_n2423_1) );
  OR2X2 OR2X2_2207 ( .A(w_mem_inst__abc_21378_n2424), .B(w_mem_inst__abc_21378_n2425), .Y(w_mem_inst__abc_21378_n2426_1) );
  OR2X2 OR2X2_2208 ( .A(w_mem_inst__abc_21378_n2426_1), .B(w_mem_inst__abc_21378_n2423_1), .Y(w_mem_inst__abc_21378_n2427_1) );
  OR2X2 OR2X2_2209 ( .A(w_mem_inst__abc_21378_n2420), .B(w_mem_inst__abc_21378_n2427_1), .Y(w_mem_inst__abc_21378_n2428) );
  OR2X2 OR2X2_221 ( .A(_auto_iopadmap_cc_313_execute_26059_56_), .B(d_reg_24_), .Y(_abc_15724_n1380) );
  OR2X2 OR2X2_2210 ( .A(w_mem_inst__abc_21378_n2428), .B(w_mem_inst__abc_21378_n2413), .Y(w_mem_inst__abc_21378_n2429) );
  OR2X2 OR2X2_2211 ( .A(w_mem_inst__abc_21378_n2429), .B(w_mem_inst__abc_21378_n2406_1), .Y(w_mem_inst__abc_21378_n2430_1) );
  OR2X2 OR2X2_2212 ( .A(w_mem_inst__abc_21378_n2432), .B(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_21378_n2433) );
  OR2X2 OR2X2_2213 ( .A(w_mem_inst__abc_21378_n2434_1), .B(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_21378_n2435_1) );
  OR2X2 OR2X2_2214 ( .A(w_mem_inst_w_mem_2__16_), .B(w_mem_inst_w_mem_0__16_), .Y(w_mem_inst__abc_21378_n2438_1) );
  OR2X2 OR2X2_2215 ( .A(w_mem_inst__abc_21378_n2437), .B(w_mem_inst__abc_21378_n2441), .Y(w_mem_inst__abc_21378_n2442_1) );
  OR2X2 OR2X2_2216 ( .A(w_mem_inst__abc_21378_n2443_1), .B(w_mem_inst__abc_21378_n2436), .Y(w_mem_inst__abc_21378_n2444) );
  OR2X2 OR2X2_2217 ( .A(w_mem_inst__abc_21378_n2445), .B(w_mem_inst__abc_21378_n1587_bF_buf2), .Y(w_mem_inst__abc_21378_n2446_1) );
  OR2X2 OR2X2_2218 ( .A(w_mem_inst__abc_21378_n2448), .B(w_mem_inst__abc_21378_n1586_bF_buf1), .Y(w_mem_inst__abc_21378_n2449) );
  OR2X2 OR2X2_2219 ( .A(w_mem_inst__abc_21378_n2450_1), .B(w_mem_inst__abc_21378_n2451_1), .Y(w_mem_inst__abc_21378_n2452) );
  OR2X2 OR2X2_222 ( .A(_abc_15724_n1379_1), .B(_abc_15724_n1383), .Y(_abc_15724_n1384) );
  OR2X2 OR2X2_2220 ( .A(w_mem_inst__abc_21378_n2452), .B(w_mem_inst__abc_21378_n2449), .Y(w_mem_inst__abc_21378_n2453) );
  OR2X2 OR2X2_2221 ( .A(w_mem_inst__abc_21378_n2453), .B(w_mem_inst__abc_21378_n2447_1), .Y(w_mem_inst__abc_21378_n2454_1) );
  OR2X2 OR2X2_2222 ( .A(w_mem_inst__abc_21378_n2455_1), .B(w_mem_inst__abc_21378_n2456), .Y(w_mem_inst__abc_21378_n2457) );
  OR2X2 OR2X2_2223 ( .A(w_mem_inst__abc_21378_n2459_1), .B(w_mem_inst__abc_21378_n2458_1), .Y(w_mem_inst__abc_21378_n2460) );
  OR2X2 OR2X2_2224 ( .A(w_mem_inst__abc_21378_n2457), .B(w_mem_inst__abc_21378_n2460), .Y(w_mem_inst__abc_21378_n2461) );
  OR2X2 OR2X2_2225 ( .A(w_mem_inst__abc_21378_n2462_1), .B(w_mem_inst__abc_21378_n2463_1), .Y(w_mem_inst__abc_21378_n2464) );
  OR2X2 OR2X2_2226 ( .A(w_mem_inst__abc_21378_n2465), .B(w_mem_inst__abc_21378_n2466_1), .Y(w_mem_inst__abc_21378_n2467_1) );
  OR2X2 OR2X2_2227 ( .A(w_mem_inst__abc_21378_n2464), .B(w_mem_inst__abc_21378_n2467_1), .Y(w_mem_inst__abc_21378_n2468) );
  OR2X2 OR2X2_2228 ( .A(w_mem_inst__abc_21378_n2469), .B(w_mem_inst__abc_21378_n2470_1), .Y(w_mem_inst__abc_21378_n2471_1) );
  OR2X2 OR2X2_2229 ( .A(w_mem_inst__abc_21378_n2472), .B(w_mem_inst__abc_21378_n2473), .Y(w_mem_inst__abc_21378_n2474_1) );
  OR2X2 OR2X2_223 ( .A(_abc_15724_n1388), .B(_abc_15724_n1365), .Y(H3_reg_24__FF_INPUT) );
  OR2X2 OR2X2_2230 ( .A(w_mem_inst__abc_21378_n2471_1), .B(w_mem_inst__abc_21378_n2474_1), .Y(w_mem_inst__abc_21378_n2475_1) );
  OR2X2 OR2X2_2231 ( .A(w_mem_inst__abc_21378_n2475_1), .B(w_mem_inst__abc_21378_n2468), .Y(w_mem_inst__abc_21378_n2476) );
  OR2X2 OR2X2_2232 ( .A(w_mem_inst__abc_21378_n2476), .B(w_mem_inst__abc_21378_n2461), .Y(w_mem_inst__abc_21378_n2477) );
  OR2X2 OR2X2_2233 ( .A(w_mem_inst__abc_21378_n2477), .B(w_mem_inst__abc_21378_n2454_1), .Y(w_mem_inst__abc_21378_n2478_1) );
  OR2X2 OR2X2_2234 ( .A(w_mem_inst__abc_21378_n2480), .B(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_21378_n2481) );
  OR2X2 OR2X2_2235 ( .A(w_mem_inst__abc_21378_n2482_1), .B(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_21378_n2483_1) );
  OR2X2 OR2X2_2236 ( .A(w_mem_inst_w_mem_2__17_), .B(w_mem_inst_w_mem_0__17_), .Y(w_mem_inst__abc_21378_n2486_1) );
  OR2X2 OR2X2_2237 ( .A(w_mem_inst__abc_21378_n2485), .B(w_mem_inst__abc_21378_n2489), .Y(w_mem_inst__abc_21378_n2490_1) );
  OR2X2 OR2X2_2238 ( .A(w_mem_inst__abc_21378_n2491_1), .B(w_mem_inst__abc_21378_n2484), .Y(w_mem_inst__abc_21378_n2492) );
  OR2X2 OR2X2_2239 ( .A(w_mem_inst__abc_21378_n2493), .B(w_mem_inst__abc_21378_n1587_bF_buf1), .Y(w_mem_inst__abc_21378_n2494_1) );
  OR2X2 OR2X2_224 ( .A(_auto_iopadmap_cc_313_execute_26059_57_), .B(d_reg_25_), .Y(_abc_15724_n1391_1) );
  OR2X2 OR2X2_2240 ( .A(w_mem_inst__abc_21378_n2496), .B(w_mem_inst__abc_21378_n1586_bF_buf0), .Y(w_mem_inst__abc_21378_n2497) );
  OR2X2 OR2X2_2241 ( .A(w_mem_inst__abc_21378_n2498_1), .B(w_mem_inst__abc_21378_n2499_1), .Y(w_mem_inst__abc_21378_n2500) );
  OR2X2 OR2X2_2242 ( .A(w_mem_inst__abc_21378_n2500), .B(w_mem_inst__abc_21378_n2497), .Y(w_mem_inst__abc_21378_n2501) );
  OR2X2 OR2X2_2243 ( .A(w_mem_inst__abc_21378_n2501), .B(w_mem_inst__abc_21378_n2495_1), .Y(w_mem_inst__abc_21378_n2502_1) );
  OR2X2 OR2X2_2244 ( .A(w_mem_inst__abc_21378_n2503_1), .B(w_mem_inst__abc_21378_n2504), .Y(w_mem_inst__abc_21378_n2505) );
  OR2X2 OR2X2_2245 ( .A(w_mem_inst__abc_21378_n2507_1), .B(w_mem_inst__abc_21378_n2506_1), .Y(w_mem_inst__abc_21378_n2508) );
  OR2X2 OR2X2_2246 ( .A(w_mem_inst__abc_21378_n2505), .B(w_mem_inst__abc_21378_n2508), .Y(w_mem_inst__abc_21378_n2509) );
  OR2X2 OR2X2_2247 ( .A(w_mem_inst__abc_21378_n2510_1), .B(w_mem_inst__abc_21378_n2511_1), .Y(w_mem_inst__abc_21378_n2512) );
  OR2X2 OR2X2_2248 ( .A(w_mem_inst__abc_21378_n2513), .B(w_mem_inst__abc_21378_n2514_1), .Y(w_mem_inst__abc_21378_n2515_1) );
  OR2X2 OR2X2_2249 ( .A(w_mem_inst__abc_21378_n2515_1), .B(w_mem_inst__abc_21378_n2512), .Y(w_mem_inst__abc_21378_n2516) );
  OR2X2 OR2X2_225 ( .A(_abc_15724_n1394), .B(_abc_15724_n1381), .Y(_abc_15724_n1395) );
  OR2X2 OR2X2_2250 ( .A(w_mem_inst__abc_21378_n2518_1), .B(w_mem_inst__abc_21378_n2517), .Y(w_mem_inst__abc_21378_n2519_1) );
  OR2X2 OR2X2_2251 ( .A(w_mem_inst__abc_21378_n2520), .B(w_mem_inst__abc_21378_n2521), .Y(w_mem_inst__abc_21378_n2522_1) );
  OR2X2 OR2X2_2252 ( .A(w_mem_inst__abc_21378_n2522_1), .B(w_mem_inst__abc_21378_n2519_1), .Y(w_mem_inst__abc_21378_n2523_1) );
  OR2X2 OR2X2_2253 ( .A(w_mem_inst__abc_21378_n2516), .B(w_mem_inst__abc_21378_n2523_1), .Y(w_mem_inst__abc_21378_n2524) );
  OR2X2 OR2X2_2254 ( .A(w_mem_inst__abc_21378_n2524), .B(w_mem_inst__abc_21378_n2509), .Y(w_mem_inst__abc_21378_n2525) );
  OR2X2 OR2X2_2255 ( .A(w_mem_inst__abc_21378_n2525), .B(w_mem_inst__abc_21378_n2502_1), .Y(w_mem_inst__abc_21378_n2526_1) );
  OR2X2 OR2X2_2256 ( .A(w_mem_inst__abc_21378_n2528), .B(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_21378_n2529) );
  OR2X2 OR2X2_2257 ( .A(w_mem_inst__abc_21378_n2530_1), .B(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_21378_n2531_1) );
  OR2X2 OR2X2_2258 ( .A(w_mem_inst_w_mem_2__18_), .B(w_mem_inst_w_mem_0__18_), .Y(w_mem_inst__abc_21378_n2534_1) );
  OR2X2 OR2X2_2259 ( .A(w_mem_inst__abc_21378_n2533), .B(w_mem_inst__abc_21378_n2537), .Y(w_mem_inst__abc_21378_n2538_1) );
  OR2X2 OR2X2_226 ( .A(_abc_15724_n1385), .B(_abc_15724_n1395), .Y(_abc_15724_n1396) );
  OR2X2 OR2X2_2260 ( .A(w_mem_inst__abc_21378_n2539_1), .B(w_mem_inst__abc_21378_n2532), .Y(w_mem_inst__abc_21378_n2540) );
  OR2X2 OR2X2_2261 ( .A(w_mem_inst__abc_21378_n2541), .B(w_mem_inst__abc_21378_n1587_bF_buf0), .Y(w_mem_inst__abc_21378_n2542_1) );
  OR2X2 OR2X2_2262 ( .A(w_mem_inst__abc_21378_n2544), .B(w_mem_inst__abc_21378_n1586_bF_buf4), .Y(w_mem_inst__abc_21378_n2545) );
  OR2X2 OR2X2_2263 ( .A(w_mem_inst__abc_21378_n2546_1), .B(w_mem_inst__abc_21378_n2547_1), .Y(w_mem_inst__abc_21378_n2548) );
  OR2X2 OR2X2_2264 ( .A(w_mem_inst__abc_21378_n2548), .B(w_mem_inst__abc_21378_n2545), .Y(w_mem_inst__abc_21378_n2549) );
  OR2X2 OR2X2_2265 ( .A(w_mem_inst__abc_21378_n2549), .B(w_mem_inst__abc_21378_n2543_1), .Y(w_mem_inst__abc_21378_n2550_1) );
  OR2X2 OR2X2_2266 ( .A(w_mem_inst__abc_21378_n2551_1), .B(w_mem_inst__abc_21378_n2552), .Y(w_mem_inst__abc_21378_n2553) );
  OR2X2 OR2X2_2267 ( .A(w_mem_inst__abc_21378_n2555_1), .B(w_mem_inst__abc_21378_n2554_1), .Y(w_mem_inst__abc_21378_n2556) );
  OR2X2 OR2X2_2268 ( .A(w_mem_inst__abc_21378_n2553), .B(w_mem_inst__abc_21378_n2556), .Y(w_mem_inst__abc_21378_n2557) );
  OR2X2 OR2X2_2269 ( .A(w_mem_inst__abc_21378_n2558_1), .B(w_mem_inst__abc_21378_n2559_1), .Y(w_mem_inst__abc_21378_n2560) );
  OR2X2 OR2X2_227 ( .A(_abc_15724_n1399_1), .B(_abc_15724_n1400_1), .Y(_abc_15724_n1401) );
  OR2X2 OR2X2_2270 ( .A(w_mem_inst__abc_21378_n2561), .B(w_mem_inst__abc_21378_n2562_1), .Y(w_mem_inst__abc_21378_n2563_1) );
  OR2X2 OR2X2_2271 ( .A(w_mem_inst__abc_21378_n2560), .B(w_mem_inst__abc_21378_n2563_1), .Y(w_mem_inst__abc_21378_n2564) );
  OR2X2 OR2X2_2272 ( .A(w_mem_inst__abc_21378_n2565), .B(w_mem_inst__abc_21378_n2566_1), .Y(w_mem_inst__abc_21378_n2567_1) );
  OR2X2 OR2X2_2273 ( .A(w_mem_inst__abc_21378_n2568), .B(w_mem_inst__abc_21378_n2569), .Y(w_mem_inst__abc_21378_n2570_1) );
  OR2X2 OR2X2_2274 ( .A(w_mem_inst__abc_21378_n2567_1), .B(w_mem_inst__abc_21378_n2570_1), .Y(w_mem_inst__abc_21378_n2571_1) );
  OR2X2 OR2X2_2275 ( .A(w_mem_inst__abc_21378_n2571_1), .B(w_mem_inst__abc_21378_n2564), .Y(w_mem_inst__abc_21378_n2572) );
  OR2X2 OR2X2_2276 ( .A(w_mem_inst__abc_21378_n2572), .B(w_mem_inst__abc_21378_n2557), .Y(w_mem_inst__abc_21378_n2573) );
  OR2X2 OR2X2_2277 ( .A(w_mem_inst__abc_21378_n2573), .B(w_mem_inst__abc_21378_n2550_1), .Y(w_mem_inst__abc_21378_n2574_1) );
  OR2X2 OR2X2_2278 ( .A(w_mem_inst__abc_21378_n2576), .B(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_21378_n2577) );
  OR2X2 OR2X2_2279 ( .A(w_mem_inst__abc_21378_n2578_1), .B(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_21378_n2579_1) );
  OR2X2 OR2X2_228 ( .A(_abc_15724_n1402_1), .B(_abc_15724_n1403), .Y(_abc_15724_n1404) );
  OR2X2 OR2X2_2280 ( .A(w_mem_inst_w_mem_2__19_), .B(w_mem_inst_w_mem_0__19_), .Y(w_mem_inst__abc_21378_n2582_1) );
  OR2X2 OR2X2_2281 ( .A(w_mem_inst__abc_21378_n2581), .B(w_mem_inst__abc_21378_n2585), .Y(w_mem_inst__abc_21378_n2586_1) );
  OR2X2 OR2X2_2282 ( .A(w_mem_inst__abc_21378_n2587_1), .B(w_mem_inst__abc_21378_n2580), .Y(w_mem_inst__abc_21378_n2588) );
  OR2X2 OR2X2_2283 ( .A(w_mem_inst__abc_21378_n2589), .B(w_mem_inst__abc_21378_n1587_bF_buf4), .Y(w_mem_inst__abc_21378_n2590_1) );
  OR2X2 OR2X2_2284 ( .A(w_mem_inst__abc_21378_n2592), .B(w_mem_inst__abc_21378_n1586_bF_buf3), .Y(w_mem_inst__abc_21378_n2593) );
  OR2X2 OR2X2_2285 ( .A(w_mem_inst__abc_21378_n2594_1), .B(w_mem_inst__abc_21378_n2595_1), .Y(w_mem_inst__abc_21378_n2596) );
  OR2X2 OR2X2_2286 ( .A(w_mem_inst__abc_21378_n2596), .B(w_mem_inst__abc_21378_n2593), .Y(w_mem_inst__abc_21378_n2597) );
  OR2X2 OR2X2_2287 ( .A(w_mem_inst__abc_21378_n2597), .B(w_mem_inst__abc_21378_n2591_1), .Y(w_mem_inst__abc_21378_n2598_1) );
  OR2X2 OR2X2_2288 ( .A(w_mem_inst__abc_21378_n2599_1), .B(w_mem_inst__abc_21378_n2600), .Y(w_mem_inst__abc_21378_n2601) );
  OR2X2 OR2X2_2289 ( .A(w_mem_inst__abc_21378_n2603_1), .B(w_mem_inst__abc_21378_n2602_1), .Y(w_mem_inst__abc_21378_n2604) );
  OR2X2 OR2X2_229 ( .A(_abc_15724_n1405), .B(_abc_15724_n1407), .Y(_abc_15724_n1408) );
  OR2X2 OR2X2_2290 ( .A(w_mem_inst__abc_21378_n2601), .B(w_mem_inst__abc_21378_n2604), .Y(w_mem_inst__abc_21378_n2605) );
  OR2X2 OR2X2_2291 ( .A(w_mem_inst__abc_21378_n2606_1), .B(w_mem_inst__abc_21378_n2607_1), .Y(w_mem_inst__abc_21378_n2608) );
  OR2X2 OR2X2_2292 ( .A(w_mem_inst__abc_21378_n2609), .B(w_mem_inst__abc_21378_n2610_1), .Y(w_mem_inst__abc_21378_n2611_1) );
  OR2X2 OR2X2_2293 ( .A(w_mem_inst__abc_21378_n2611_1), .B(w_mem_inst__abc_21378_n2608), .Y(w_mem_inst__abc_21378_n2612) );
  OR2X2 OR2X2_2294 ( .A(w_mem_inst__abc_21378_n2614_1), .B(w_mem_inst__abc_21378_n2613), .Y(w_mem_inst__abc_21378_n2615_1) );
  OR2X2 OR2X2_2295 ( .A(w_mem_inst__abc_21378_n2616), .B(w_mem_inst__abc_21378_n2617), .Y(w_mem_inst__abc_21378_n2618_1) );
  OR2X2 OR2X2_2296 ( .A(w_mem_inst__abc_21378_n2618_1), .B(w_mem_inst__abc_21378_n2615_1), .Y(w_mem_inst__abc_21378_n2619_1) );
  OR2X2 OR2X2_2297 ( .A(w_mem_inst__abc_21378_n2612), .B(w_mem_inst__abc_21378_n2619_1), .Y(w_mem_inst__abc_21378_n2620) );
  OR2X2 OR2X2_2298 ( .A(w_mem_inst__abc_21378_n2620), .B(w_mem_inst__abc_21378_n2605), .Y(w_mem_inst__abc_21378_n2621) );
  OR2X2 OR2X2_2299 ( .A(w_mem_inst__abc_21378_n2621), .B(w_mem_inst__abc_21378_n2598_1), .Y(w_mem_inst__abc_21378_n2622_1) );
  OR2X2 OR2X2_23 ( .A(_auto_iopadmap_cc_313_execute_26059_6_), .B(e_reg_6_), .Y(_abc_15724_n781_1) );
  OR2X2 OR2X2_230 ( .A(_abc_15724_n1413_1), .B(_abc_15724_n1390_1), .Y(H3_reg_25__FF_INPUT) );
  OR2X2 OR2X2_2300 ( .A(w_mem_inst__abc_21378_n2624), .B(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_21378_n2625) );
  OR2X2 OR2X2_2301 ( .A(w_mem_inst__abc_21378_n2626_1), .B(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_21378_n2627_1) );
  OR2X2 OR2X2_2302 ( .A(w_mem_inst_w_mem_2__20_), .B(w_mem_inst_w_mem_0__20_), .Y(w_mem_inst__abc_21378_n2630_1) );
  OR2X2 OR2X2_2303 ( .A(w_mem_inst__abc_21378_n2629), .B(w_mem_inst__abc_21378_n2633), .Y(w_mem_inst__abc_21378_n2634_1) );
  OR2X2 OR2X2_2304 ( .A(w_mem_inst__abc_21378_n2635_1), .B(w_mem_inst__abc_21378_n2628), .Y(w_mem_inst__abc_21378_n2636) );
  OR2X2 OR2X2_2305 ( .A(w_mem_inst__abc_21378_n2637), .B(w_mem_inst__abc_21378_n1587_bF_buf3), .Y(w_mem_inst__abc_21378_n2638_1) );
  OR2X2 OR2X2_2306 ( .A(w_mem_inst__abc_21378_n2640), .B(w_mem_inst__abc_21378_n1586_bF_buf2), .Y(w_mem_inst__abc_21378_n2641) );
  OR2X2 OR2X2_2307 ( .A(w_mem_inst__abc_21378_n2642_1), .B(w_mem_inst__abc_21378_n2643_1), .Y(w_mem_inst__abc_21378_n2644) );
  OR2X2 OR2X2_2308 ( .A(w_mem_inst__abc_21378_n2644), .B(w_mem_inst__abc_21378_n2641), .Y(w_mem_inst__abc_21378_n2645) );
  OR2X2 OR2X2_2309 ( .A(w_mem_inst__abc_21378_n2645), .B(w_mem_inst__abc_21378_n2639_1), .Y(w_mem_inst__abc_21378_n2646_1) );
  OR2X2 OR2X2_231 ( .A(_abc_15724_n1416_1), .B(_abc_15724_n1418), .Y(_abc_15724_n1419) );
  OR2X2 OR2X2_2310 ( .A(w_mem_inst__abc_21378_n2647_1), .B(w_mem_inst__abc_21378_n2648), .Y(w_mem_inst__abc_21378_n2649) );
  OR2X2 OR2X2_2311 ( .A(w_mem_inst__abc_21378_n2651_1), .B(w_mem_inst__abc_21378_n2650_1), .Y(w_mem_inst__abc_21378_n2652) );
  OR2X2 OR2X2_2312 ( .A(w_mem_inst__abc_21378_n2649), .B(w_mem_inst__abc_21378_n2652), .Y(w_mem_inst__abc_21378_n2653) );
  OR2X2 OR2X2_2313 ( .A(w_mem_inst__abc_21378_n2654_1), .B(w_mem_inst__abc_21378_n2655_1), .Y(w_mem_inst__abc_21378_n2656) );
  OR2X2 OR2X2_2314 ( .A(w_mem_inst__abc_21378_n2657), .B(w_mem_inst__abc_21378_n2658_1), .Y(w_mem_inst__abc_21378_n2659_1) );
  OR2X2 OR2X2_2315 ( .A(w_mem_inst__abc_21378_n2656), .B(w_mem_inst__abc_21378_n2659_1), .Y(w_mem_inst__abc_21378_n2660) );
  OR2X2 OR2X2_2316 ( .A(w_mem_inst__abc_21378_n2661), .B(w_mem_inst__abc_21378_n2662_1), .Y(w_mem_inst__abc_21378_n2663_1) );
  OR2X2 OR2X2_2317 ( .A(w_mem_inst__abc_21378_n2664), .B(w_mem_inst__abc_21378_n2665), .Y(w_mem_inst__abc_21378_n2666_1) );
  OR2X2 OR2X2_2318 ( .A(w_mem_inst__abc_21378_n2663_1), .B(w_mem_inst__abc_21378_n2666_1), .Y(w_mem_inst__abc_21378_n2667_1) );
  OR2X2 OR2X2_2319 ( .A(w_mem_inst__abc_21378_n2667_1), .B(w_mem_inst__abc_21378_n2660), .Y(w_mem_inst__abc_21378_n2668) );
  OR2X2 OR2X2_232 ( .A(_auto_iopadmap_cc_313_execute_26059_58_), .B(d_reg_26_), .Y(_abc_15724_n1420) );
  OR2X2 OR2X2_2320 ( .A(w_mem_inst__abc_21378_n2668), .B(w_mem_inst__abc_21378_n2653), .Y(w_mem_inst__abc_21378_n2669) );
  OR2X2 OR2X2_2321 ( .A(w_mem_inst__abc_21378_n2669), .B(w_mem_inst__abc_21378_n2646_1), .Y(w_mem_inst__abc_21378_n2670_1) );
  OR2X2 OR2X2_2322 ( .A(w_mem_inst__abc_21378_n2672), .B(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_21378_n2673) );
  OR2X2 OR2X2_2323 ( .A(w_mem_inst__abc_21378_n2674_1), .B(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_21378_n2675_1) );
  OR2X2 OR2X2_2324 ( .A(w_mem_inst_w_mem_2__21_), .B(w_mem_inst_w_mem_0__21_), .Y(w_mem_inst__abc_21378_n2678_1) );
  OR2X2 OR2X2_2325 ( .A(w_mem_inst__abc_21378_n2677), .B(w_mem_inst__abc_21378_n2681), .Y(w_mem_inst__abc_21378_n2682_1) );
  OR2X2 OR2X2_2326 ( .A(w_mem_inst__abc_21378_n2683_1), .B(w_mem_inst__abc_21378_n2676), .Y(w_mem_inst__abc_21378_n2684) );
  OR2X2 OR2X2_2327 ( .A(w_mem_inst__abc_21378_n2685), .B(w_mem_inst__abc_21378_n1587_bF_buf2), .Y(w_mem_inst__abc_21378_n2686_1) );
  OR2X2 OR2X2_2328 ( .A(w_mem_inst__abc_21378_n2688), .B(w_mem_inst__abc_21378_n1586_bF_buf1), .Y(w_mem_inst__abc_21378_n2689) );
  OR2X2 OR2X2_2329 ( .A(w_mem_inst__abc_21378_n2690_1), .B(w_mem_inst__abc_21378_n2691_1), .Y(w_mem_inst__abc_21378_n2692) );
  OR2X2 OR2X2_233 ( .A(_abc_15724_n1419), .B(_abc_15724_n1423_1), .Y(_abc_15724_n1424_1) );
  OR2X2 OR2X2_2330 ( .A(w_mem_inst__abc_21378_n2692), .B(w_mem_inst__abc_21378_n2689), .Y(w_mem_inst__abc_21378_n2693) );
  OR2X2 OR2X2_2331 ( .A(w_mem_inst__abc_21378_n2693), .B(w_mem_inst__abc_21378_n2687_1), .Y(w_mem_inst__abc_21378_n2694_1) );
  OR2X2 OR2X2_2332 ( .A(w_mem_inst__abc_21378_n2695_1), .B(w_mem_inst__abc_21378_n2696), .Y(w_mem_inst__abc_21378_n2697) );
  OR2X2 OR2X2_2333 ( .A(w_mem_inst__abc_21378_n2699_1), .B(w_mem_inst__abc_21378_n2698_1), .Y(w_mem_inst__abc_21378_n2700) );
  OR2X2 OR2X2_2334 ( .A(w_mem_inst__abc_21378_n2697), .B(w_mem_inst__abc_21378_n2700), .Y(w_mem_inst__abc_21378_n2701) );
  OR2X2 OR2X2_2335 ( .A(w_mem_inst__abc_21378_n2702_1), .B(w_mem_inst__abc_21378_n2703_1), .Y(w_mem_inst__abc_21378_n2704) );
  OR2X2 OR2X2_2336 ( .A(w_mem_inst__abc_21378_n2705), .B(w_mem_inst__abc_21378_n2706_1), .Y(w_mem_inst__abc_21378_n2707_1) );
  OR2X2 OR2X2_2337 ( .A(w_mem_inst__abc_21378_n2707_1), .B(w_mem_inst__abc_21378_n2704), .Y(w_mem_inst__abc_21378_n2708) );
  OR2X2 OR2X2_2338 ( .A(w_mem_inst__abc_21378_n2710_1), .B(w_mem_inst__abc_21378_n2709), .Y(w_mem_inst__abc_21378_n2711_1) );
  OR2X2 OR2X2_2339 ( .A(w_mem_inst__abc_21378_n2712), .B(w_mem_inst__abc_21378_n2713), .Y(w_mem_inst__abc_21378_n2714_1) );
  OR2X2 OR2X2_234 ( .A(_abc_15724_n1428), .B(_abc_15724_n1415), .Y(H3_reg_26__FF_INPUT) );
  OR2X2 OR2X2_2340 ( .A(w_mem_inst__abc_21378_n2714_1), .B(w_mem_inst__abc_21378_n2711_1), .Y(w_mem_inst__abc_21378_n2715_1) );
  OR2X2 OR2X2_2341 ( .A(w_mem_inst__abc_21378_n2708), .B(w_mem_inst__abc_21378_n2715_1), .Y(w_mem_inst__abc_21378_n2716) );
  OR2X2 OR2X2_2342 ( .A(w_mem_inst__abc_21378_n2716), .B(w_mem_inst__abc_21378_n2701), .Y(w_mem_inst__abc_21378_n2717) );
  OR2X2 OR2X2_2343 ( .A(w_mem_inst__abc_21378_n2717), .B(w_mem_inst__abc_21378_n2694_1), .Y(w_mem_inst__abc_21378_n2718_1) );
  OR2X2 OR2X2_2344 ( .A(w_mem_inst__abc_21378_n2720), .B(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_21378_n2721) );
  OR2X2 OR2X2_2345 ( .A(w_mem_inst__abc_21378_n2722_1), .B(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_21378_n2723_1) );
  OR2X2 OR2X2_2346 ( .A(w_mem_inst_w_mem_2__22_), .B(w_mem_inst_w_mem_0__22_), .Y(w_mem_inst__abc_21378_n2726_1) );
  OR2X2 OR2X2_2347 ( .A(w_mem_inst__abc_21378_n2725), .B(w_mem_inst__abc_21378_n2729), .Y(w_mem_inst__abc_21378_n2730_1) );
  OR2X2 OR2X2_2348 ( .A(w_mem_inst__abc_21378_n2731_1), .B(w_mem_inst__abc_21378_n2724), .Y(w_mem_inst__abc_21378_n2732) );
  OR2X2 OR2X2_2349 ( .A(w_mem_inst__abc_21378_n2733), .B(w_mem_inst__abc_21378_n1587_bF_buf1), .Y(w_mem_inst__abc_21378_n2734_1) );
  OR2X2 OR2X2_235 ( .A(_auto_iopadmap_cc_313_execute_26059_59_), .B(d_reg_27_), .Y(_abc_15724_n1431) );
  OR2X2 OR2X2_2350 ( .A(w_mem_inst__abc_21378_n2736), .B(w_mem_inst__abc_21378_n1586_bF_buf0), .Y(w_mem_inst__abc_21378_n2737) );
  OR2X2 OR2X2_2351 ( .A(w_mem_inst__abc_21378_n2738_1), .B(w_mem_inst__abc_21378_n2739_1), .Y(w_mem_inst__abc_21378_n2740) );
  OR2X2 OR2X2_2352 ( .A(w_mem_inst__abc_21378_n2740), .B(w_mem_inst__abc_21378_n2737), .Y(w_mem_inst__abc_21378_n2741) );
  OR2X2 OR2X2_2353 ( .A(w_mem_inst__abc_21378_n2741), .B(w_mem_inst__abc_21378_n2735_1), .Y(w_mem_inst__abc_21378_n2742_1) );
  OR2X2 OR2X2_2354 ( .A(w_mem_inst__abc_21378_n2743_1), .B(w_mem_inst__abc_21378_n2744), .Y(w_mem_inst__abc_21378_n2745) );
  OR2X2 OR2X2_2355 ( .A(w_mem_inst__abc_21378_n2747_1), .B(w_mem_inst__abc_21378_n2746_1), .Y(w_mem_inst__abc_21378_n2748) );
  OR2X2 OR2X2_2356 ( .A(w_mem_inst__abc_21378_n2745), .B(w_mem_inst__abc_21378_n2748), .Y(w_mem_inst__abc_21378_n2749) );
  OR2X2 OR2X2_2357 ( .A(w_mem_inst__abc_21378_n2750_1), .B(w_mem_inst__abc_21378_n2751_1), .Y(w_mem_inst__abc_21378_n2752) );
  OR2X2 OR2X2_2358 ( .A(w_mem_inst__abc_21378_n2753), .B(w_mem_inst__abc_21378_n2754_1), .Y(w_mem_inst__abc_21378_n2755_1) );
  OR2X2 OR2X2_2359 ( .A(w_mem_inst__abc_21378_n2752), .B(w_mem_inst__abc_21378_n2755_1), .Y(w_mem_inst__abc_21378_n2756) );
  OR2X2 OR2X2_236 ( .A(_abc_15724_n1434), .B(_abc_15724_n1421), .Y(_abc_15724_n1435_1) );
  OR2X2 OR2X2_2360 ( .A(w_mem_inst__abc_21378_n2757), .B(w_mem_inst__abc_21378_n2758_1), .Y(w_mem_inst__abc_21378_n2759_1) );
  OR2X2 OR2X2_2361 ( .A(w_mem_inst__abc_21378_n2760), .B(w_mem_inst__abc_21378_n2761), .Y(w_mem_inst__abc_21378_n2762_1) );
  OR2X2 OR2X2_2362 ( .A(w_mem_inst__abc_21378_n2759_1), .B(w_mem_inst__abc_21378_n2762_1), .Y(w_mem_inst__abc_21378_n2763_1) );
  OR2X2 OR2X2_2363 ( .A(w_mem_inst__abc_21378_n2763_1), .B(w_mem_inst__abc_21378_n2756), .Y(w_mem_inst__abc_21378_n2764) );
  OR2X2 OR2X2_2364 ( .A(w_mem_inst__abc_21378_n2764), .B(w_mem_inst__abc_21378_n2749), .Y(w_mem_inst__abc_21378_n2765) );
  OR2X2 OR2X2_2365 ( .A(w_mem_inst__abc_21378_n2765), .B(w_mem_inst__abc_21378_n2742_1), .Y(w_mem_inst__abc_21378_n2766_1) );
  OR2X2 OR2X2_2366 ( .A(w_mem_inst__abc_21378_n2768), .B(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_21378_n2769) );
  OR2X2 OR2X2_2367 ( .A(w_mem_inst__abc_21378_n2770_1), .B(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_21378_n2771_1) );
  OR2X2 OR2X2_2368 ( .A(w_mem_inst_w_mem_2__23_), .B(w_mem_inst_w_mem_0__23_), .Y(w_mem_inst__abc_21378_n2774_1) );
  OR2X2 OR2X2_2369 ( .A(w_mem_inst__abc_21378_n2773), .B(w_mem_inst__abc_21378_n2777), .Y(w_mem_inst__abc_21378_n2778_1) );
  OR2X2 OR2X2_237 ( .A(_abc_15724_n1425), .B(_abc_15724_n1435_1), .Y(_abc_15724_n1436_1) );
  OR2X2 OR2X2_2370 ( .A(w_mem_inst__abc_21378_n2779_1), .B(w_mem_inst__abc_21378_n2772), .Y(w_mem_inst__abc_21378_n2780) );
  OR2X2 OR2X2_2371 ( .A(w_mem_inst__abc_21378_n2781), .B(w_mem_inst__abc_21378_n1587_bF_buf0), .Y(w_mem_inst__abc_21378_n2782_1) );
  OR2X2 OR2X2_2372 ( .A(w_mem_inst__abc_21378_n2784), .B(w_mem_inst__abc_21378_n1586_bF_buf4), .Y(w_mem_inst__abc_21378_n2785) );
  OR2X2 OR2X2_2373 ( .A(w_mem_inst__abc_21378_n2786_1), .B(w_mem_inst__abc_21378_n2787_1), .Y(w_mem_inst__abc_21378_n2788) );
  OR2X2 OR2X2_2374 ( .A(w_mem_inst__abc_21378_n2788), .B(w_mem_inst__abc_21378_n2785), .Y(w_mem_inst__abc_21378_n2789) );
  OR2X2 OR2X2_2375 ( .A(w_mem_inst__abc_21378_n2789), .B(w_mem_inst__abc_21378_n2783_1), .Y(w_mem_inst__abc_21378_n2790_1) );
  OR2X2 OR2X2_2376 ( .A(w_mem_inst__abc_21378_n2791_1), .B(w_mem_inst__abc_21378_n2792), .Y(w_mem_inst__abc_21378_n2793) );
  OR2X2 OR2X2_2377 ( .A(w_mem_inst__abc_21378_n2795_1), .B(w_mem_inst__abc_21378_n2794_1), .Y(w_mem_inst__abc_21378_n2796) );
  OR2X2 OR2X2_2378 ( .A(w_mem_inst__abc_21378_n2793), .B(w_mem_inst__abc_21378_n2796), .Y(w_mem_inst__abc_21378_n2797) );
  OR2X2 OR2X2_2379 ( .A(w_mem_inst__abc_21378_n2798_1), .B(w_mem_inst__abc_21378_n2799_1), .Y(w_mem_inst__abc_21378_n2800) );
  OR2X2 OR2X2_238 ( .A(_abc_15724_n1437), .B(_abc_15724_n1439), .Y(_abc_15724_n1440) );
  OR2X2 OR2X2_2380 ( .A(w_mem_inst__abc_21378_n2801), .B(w_mem_inst__abc_21378_n2802_1), .Y(w_mem_inst__abc_21378_n2803_1) );
  OR2X2 OR2X2_2381 ( .A(w_mem_inst__abc_21378_n2803_1), .B(w_mem_inst__abc_21378_n2800), .Y(w_mem_inst__abc_21378_n2804) );
  OR2X2 OR2X2_2382 ( .A(w_mem_inst__abc_21378_n2806_1), .B(w_mem_inst__abc_21378_n2805), .Y(w_mem_inst__abc_21378_n2807_1) );
  OR2X2 OR2X2_2383 ( .A(w_mem_inst__abc_21378_n2808), .B(w_mem_inst__abc_21378_n2809), .Y(w_mem_inst__abc_21378_n2810_1) );
  OR2X2 OR2X2_2384 ( .A(w_mem_inst__abc_21378_n2810_1), .B(w_mem_inst__abc_21378_n2807_1), .Y(w_mem_inst__abc_21378_n2811_1) );
  OR2X2 OR2X2_2385 ( .A(w_mem_inst__abc_21378_n2804), .B(w_mem_inst__abc_21378_n2811_1), .Y(w_mem_inst__abc_21378_n2812) );
  OR2X2 OR2X2_2386 ( .A(w_mem_inst__abc_21378_n2812), .B(w_mem_inst__abc_21378_n2797), .Y(w_mem_inst__abc_21378_n2813) );
  OR2X2 OR2X2_2387 ( .A(w_mem_inst__abc_21378_n2813), .B(w_mem_inst__abc_21378_n2790_1), .Y(w_mem_inst__abc_21378_n2814_1) );
  OR2X2 OR2X2_2388 ( .A(w_mem_inst__abc_21378_n2816), .B(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_21378_n2817) );
  OR2X2 OR2X2_2389 ( .A(w_mem_inst__abc_21378_n2818_1), .B(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_21378_n2819_1) );
  OR2X2 OR2X2_239 ( .A(_abc_15724_n1445_1), .B(_abc_15724_n1430), .Y(H3_reg_27__FF_INPUT) );
  OR2X2 OR2X2_2390 ( .A(w_mem_inst_w_mem_2__24_), .B(w_mem_inst_w_mem_0__24_), .Y(w_mem_inst__abc_21378_n2822_1) );
  OR2X2 OR2X2_2391 ( .A(w_mem_inst__abc_21378_n2821), .B(w_mem_inst__abc_21378_n2825), .Y(w_mem_inst__abc_21378_n2826_1) );
  OR2X2 OR2X2_2392 ( .A(w_mem_inst__abc_21378_n2827_1), .B(w_mem_inst__abc_21378_n2820), .Y(w_mem_inst__abc_21378_n2828) );
  OR2X2 OR2X2_2393 ( .A(w_mem_inst__abc_21378_n2829), .B(w_mem_inst__abc_21378_n1587_bF_buf4), .Y(w_mem_inst__abc_21378_n2830_1) );
  OR2X2 OR2X2_2394 ( .A(w_mem_inst__abc_21378_n2832), .B(w_mem_inst__abc_21378_n1586_bF_buf3), .Y(w_mem_inst__abc_21378_n2833) );
  OR2X2 OR2X2_2395 ( .A(w_mem_inst__abc_21378_n2834_1), .B(w_mem_inst__abc_21378_n2835_1), .Y(w_mem_inst__abc_21378_n2836) );
  OR2X2 OR2X2_2396 ( .A(w_mem_inst__abc_21378_n2836), .B(w_mem_inst__abc_21378_n2833), .Y(w_mem_inst__abc_21378_n2837) );
  OR2X2 OR2X2_2397 ( .A(w_mem_inst__abc_21378_n2837), .B(w_mem_inst__abc_21378_n2831_1), .Y(w_mem_inst__abc_21378_n2838_1) );
  OR2X2 OR2X2_2398 ( .A(w_mem_inst__abc_21378_n2839_1), .B(w_mem_inst__abc_21378_n2840), .Y(w_mem_inst__abc_21378_n2841) );
  OR2X2 OR2X2_2399 ( .A(w_mem_inst__abc_21378_n2843_1), .B(w_mem_inst__abc_21378_n2842_1), .Y(w_mem_inst__abc_21378_n2844) );
  OR2X2 OR2X2_24 ( .A(_auto_iopadmap_cc_313_execute_26059_5_), .B(e_reg_5_), .Y(_abc_15724_n785) );
  OR2X2 OR2X2_240 ( .A(_abc_15724_n1447), .B(_abc_15724_n1449), .Y(_abc_15724_n1450) );
  OR2X2 OR2X2_2400 ( .A(w_mem_inst__abc_21378_n2841), .B(w_mem_inst__abc_21378_n2844), .Y(w_mem_inst__abc_21378_n2845) );
  OR2X2 OR2X2_2401 ( .A(w_mem_inst__abc_21378_n2846_1), .B(w_mem_inst__abc_21378_n2847_1), .Y(w_mem_inst__abc_21378_n2848) );
  OR2X2 OR2X2_2402 ( .A(w_mem_inst__abc_21378_n2849), .B(w_mem_inst__abc_21378_n2850_1), .Y(w_mem_inst__abc_21378_n2851_1) );
  OR2X2 OR2X2_2403 ( .A(w_mem_inst__abc_21378_n2848), .B(w_mem_inst__abc_21378_n2851_1), .Y(w_mem_inst__abc_21378_n2852) );
  OR2X2 OR2X2_2404 ( .A(w_mem_inst__abc_21378_n2853), .B(w_mem_inst__abc_21378_n2854_1), .Y(w_mem_inst__abc_21378_n2855_1) );
  OR2X2 OR2X2_2405 ( .A(w_mem_inst__abc_21378_n2856), .B(w_mem_inst__abc_21378_n2857), .Y(w_mem_inst__abc_21378_n2858_1) );
  OR2X2 OR2X2_2406 ( .A(w_mem_inst__abc_21378_n2855_1), .B(w_mem_inst__abc_21378_n2858_1), .Y(w_mem_inst__abc_21378_n2859_1) );
  OR2X2 OR2X2_2407 ( .A(w_mem_inst__abc_21378_n2859_1), .B(w_mem_inst__abc_21378_n2852), .Y(w_mem_inst__abc_21378_n2860) );
  OR2X2 OR2X2_2408 ( .A(w_mem_inst__abc_21378_n2860), .B(w_mem_inst__abc_21378_n2845), .Y(w_mem_inst__abc_21378_n2861) );
  OR2X2 OR2X2_2409 ( .A(w_mem_inst__abc_21378_n2861), .B(w_mem_inst__abc_21378_n2838_1), .Y(w_mem_inst__abc_21378_n2862_1) );
  OR2X2 OR2X2_241 ( .A(_auto_iopadmap_cc_313_execute_26059_60_), .B(d_reg_28_), .Y(_abc_15724_n1451) );
  OR2X2 OR2X2_2410 ( .A(w_mem_inst__abc_21378_n2864), .B(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_21378_n2865) );
  OR2X2 OR2X2_2411 ( .A(w_mem_inst__abc_21378_n2866_1), .B(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_21378_n2867_1) );
  OR2X2 OR2X2_2412 ( .A(w_mem_inst_w_mem_2__25_), .B(w_mem_inst_w_mem_0__25_), .Y(w_mem_inst__abc_21378_n2870_1) );
  OR2X2 OR2X2_2413 ( .A(w_mem_inst__abc_21378_n2869), .B(w_mem_inst__abc_21378_n2873), .Y(w_mem_inst__abc_21378_n2874_1) );
  OR2X2 OR2X2_2414 ( .A(w_mem_inst__abc_21378_n2875_1), .B(w_mem_inst__abc_21378_n2868), .Y(w_mem_inst__abc_21378_n2876) );
  OR2X2 OR2X2_2415 ( .A(w_mem_inst__abc_21378_n2877), .B(w_mem_inst__abc_21378_n1587_bF_buf3), .Y(w_mem_inst__abc_21378_n2878_1) );
  OR2X2 OR2X2_2416 ( .A(w_mem_inst__abc_21378_n2880), .B(w_mem_inst__abc_21378_n1586_bF_buf2), .Y(w_mem_inst__abc_21378_n2881) );
  OR2X2 OR2X2_2417 ( .A(w_mem_inst__abc_21378_n2882_1), .B(w_mem_inst__abc_21378_n2883_1), .Y(w_mem_inst__abc_21378_n2884) );
  OR2X2 OR2X2_2418 ( .A(w_mem_inst__abc_21378_n2884), .B(w_mem_inst__abc_21378_n2881), .Y(w_mem_inst__abc_21378_n2885) );
  OR2X2 OR2X2_2419 ( .A(w_mem_inst__abc_21378_n2885), .B(w_mem_inst__abc_21378_n2879_1), .Y(w_mem_inst__abc_21378_n2886_1) );
  OR2X2 OR2X2_242 ( .A(_abc_15724_n1450), .B(_abc_15724_n1454), .Y(_abc_15724_n1455) );
  OR2X2 OR2X2_2420 ( .A(w_mem_inst__abc_21378_n2887_1), .B(w_mem_inst__abc_21378_n2888), .Y(w_mem_inst__abc_21378_n2889) );
  OR2X2 OR2X2_2421 ( .A(w_mem_inst__abc_21378_n2891_1), .B(w_mem_inst__abc_21378_n2890_1), .Y(w_mem_inst__abc_21378_n2892) );
  OR2X2 OR2X2_2422 ( .A(w_mem_inst__abc_21378_n2889), .B(w_mem_inst__abc_21378_n2892), .Y(w_mem_inst__abc_21378_n2893) );
  OR2X2 OR2X2_2423 ( .A(w_mem_inst__abc_21378_n2894_1), .B(w_mem_inst__abc_21378_n2895_1), .Y(w_mem_inst__abc_21378_n2896) );
  OR2X2 OR2X2_2424 ( .A(w_mem_inst__abc_21378_n2897), .B(w_mem_inst__abc_21378_n2898_1), .Y(w_mem_inst__abc_21378_n2899_1) );
  OR2X2 OR2X2_2425 ( .A(w_mem_inst__abc_21378_n2899_1), .B(w_mem_inst__abc_21378_n2896), .Y(w_mem_inst__abc_21378_n2900) );
  OR2X2 OR2X2_2426 ( .A(w_mem_inst__abc_21378_n2902_1), .B(w_mem_inst__abc_21378_n2901), .Y(w_mem_inst__abc_21378_n2903_1) );
  OR2X2 OR2X2_2427 ( .A(w_mem_inst__abc_21378_n2904), .B(w_mem_inst__abc_21378_n2905), .Y(w_mem_inst__abc_21378_n2906_1) );
  OR2X2 OR2X2_2428 ( .A(w_mem_inst__abc_21378_n2906_1), .B(w_mem_inst__abc_21378_n2903_1), .Y(w_mem_inst__abc_21378_n2907_1) );
  OR2X2 OR2X2_2429 ( .A(w_mem_inst__abc_21378_n2900), .B(w_mem_inst__abc_21378_n2907_1), .Y(w_mem_inst__abc_21378_n2908) );
  OR2X2 OR2X2_243 ( .A(_abc_15724_n1456), .B(_abc_15724_n1457), .Y(_abc_15724_n1458) );
  OR2X2 OR2X2_2430 ( .A(w_mem_inst__abc_21378_n2908), .B(w_mem_inst__abc_21378_n2893), .Y(w_mem_inst__abc_21378_n2909) );
  OR2X2 OR2X2_2431 ( .A(w_mem_inst__abc_21378_n2909), .B(w_mem_inst__abc_21378_n2886_1), .Y(w_mem_inst__abc_21378_n2910_1) );
  OR2X2 OR2X2_2432 ( .A(w_mem_inst__abc_21378_n2912), .B(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_21378_n2913) );
  OR2X2 OR2X2_2433 ( .A(w_mem_inst__abc_21378_n2914_1), .B(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_21378_n2915_1) );
  OR2X2 OR2X2_2434 ( .A(w_mem_inst_w_mem_2__26_), .B(w_mem_inst_w_mem_0__26_), .Y(w_mem_inst__abc_21378_n2918_1) );
  OR2X2 OR2X2_2435 ( .A(w_mem_inst__abc_21378_n2917), .B(w_mem_inst__abc_21378_n2921), .Y(w_mem_inst__abc_21378_n2922_1) );
  OR2X2 OR2X2_2436 ( .A(w_mem_inst__abc_21378_n2923_1), .B(w_mem_inst__abc_21378_n2916), .Y(w_mem_inst__abc_21378_n2924) );
  OR2X2 OR2X2_2437 ( .A(w_mem_inst__abc_21378_n2925), .B(w_mem_inst__abc_21378_n1587_bF_buf2), .Y(w_mem_inst__abc_21378_n2926_1) );
  OR2X2 OR2X2_2438 ( .A(w_mem_inst__abc_21378_n2928), .B(w_mem_inst__abc_21378_n1586_bF_buf1), .Y(w_mem_inst__abc_21378_n2929) );
  OR2X2 OR2X2_2439 ( .A(w_mem_inst__abc_21378_n2930_1), .B(w_mem_inst__abc_21378_n2931_1), .Y(w_mem_inst__abc_21378_n2932) );
  OR2X2 OR2X2_244 ( .A(_abc_15724_n851_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_60_), .Y(_abc_15724_n1461) );
  OR2X2 OR2X2_2440 ( .A(w_mem_inst__abc_21378_n2932), .B(w_mem_inst__abc_21378_n2929), .Y(w_mem_inst__abc_21378_n2933) );
  OR2X2 OR2X2_2441 ( .A(w_mem_inst__abc_21378_n2933), .B(w_mem_inst__abc_21378_n2927_1), .Y(w_mem_inst__abc_21378_n2934_1) );
  OR2X2 OR2X2_2442 ( .A(w_mem_inst__abc_21378_n2935_1), .B(w_mem_inst__abc_21378_n2936), .Y(w_mem_inst__abc_21378_n2937) );
  OR2X2 OR2X2_2443 ( .A(w_mem_inst__abc_21378_n2939_1), .B(w_mem_inst__abc_21378_n2938_1), .Y(w_mem_inst__abc_21378_n2940) );
  OR2X2 OR2X2_2444 ( .A(w_mem_inst__abc_21378_n2937), .B(w_mem_inst__abc_21378_n2940), .Y(w_mem_inst__abc_21378_n2941) );
  OR2X2 OR2X2_2445 ( .A(w_mem_inst__abc_21378_n2942_1), .B(w_mem_inst__abc_21378_n2943_1), .Y(w_mem_inst__abc_21378_n2944) );
  OR2X2 OR2X2_2446 ( .A(w_mem_inst__abc_21378_n2945), .B(w_mem_inst__abc_21378_n2946_1), .Y(w_mem_inst__abc_21378_n2947_1) );
  OR2X2 OR2X2_2447 ( .A(w_mem_inst__abc_21378_n2944), .B(w_mem_inst__abc_21378_n2947_1), .Y(w_mem_inst__abc_21378_n2948) );
  OR2X2 OR2X2_2448 ( .A(w_mem_inst__abc_21378_n2949), .B(w_mem_inst__abc_21378_n2950_1), .Y(w_mem_inst__abc_21378_n2951_1) );
  OR2X2 OR2X2_2449 ( .A(w_mem_inst__abc_21378_n2952), .B(w_mem_inst__abc_21378_n2953), .Y(w_mem_inst__abc_21378_n2954_1) );
  OR2X2 OR2X2_245 ( .A(_abc_15724_n1460), .B(_abc_15724_n1462_1), .Y(H3_reg_28__FF_INPUT) );
  OR2X2 OR2X2_2450 ( .A(w_mem_inst__abc_21378_n2951_1), .B(w_mem_inst__abc_21378_n2954_1), .Y(w_mem_inst__abc_21378_n2955_1) );
  OR2X2 OR2X2_2451 ( .A(w_mem_inst__abc_21378_n2955_1), .B(w_mem_inst__abc_21378_n2948), .Y(w_mem_inst__abc_21378_n2956) );
  OR2X2 OR2X2_2452 ( .A(w_mem_inst__abc_21378_n2956), .B(w_mem_inst__abc_21378_n2941), .Y(w_mem_inst__abc_21378_n2957) );
  OR2X2 OR2X2_2453 ( .A(w_mem_inst__abc_21378_n2957), .B(w_mem_inst__abc_21378_n2934_1), .Y(w_mem_inst__abc_21378_n2958_1) );
  OR2X2 OR2X2_2454 ( .A(w_mem_inst__abc_21378_n2960), .B(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_21378_n2961) );
  OR2X2 OR2X2_2455 ( .A(w_mem_inst__abc_21378_n2962_1), .B(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_21378_n2963_1) );
  OR2X2 OR2X2_2456 ( .A(w_mem_inst_w_mem_2__27_), .B(w_mem_inst_w_mem_0__27_), .Y(w_mem_inst__abc_21378_n2966_1) );
  OR2X2 OR2X2_2457 ( .A(w_mem_inst__abc_21378_n2965), .B(w_mem_inst__abc_21378_n2969), .Y(w_mem_inst__abc_21378_n2970_1) );
  OR2X2 OR2X2_2458 ( .A(w_mem_inst__abc_21378_n2971_1), .B(w_mem_inst__abc_21378_n2964), .Y(w_mem_inst__abc_21378_n2972) );
  OR2X2 OR2X2_2459 ( .A(w_mem_inst__abc_21378_n2973), .B(w_mem_inst__abc_21378_n1587_bF_buf1), .Y(w_mem_inst__abc_21378_n2974_1) );
  OR2X2 OR2X2_246 ( .A(_abc_15724_n1464_1), .B(digest_update_bF_buf7), .Y(_abc_15724_n1465) );
  OR2X2 OR2X2_2460 ( .A(w_mem_inst__abc_21378_n2976), .B(w_mem_inst__abc_21378_n1586_bF_buf0), .Y(w_mem_inst__abc_21378_n2977) );
  OR2X2 OR2X2_2461 ( .A(w_mem_inst__abc_21378_n2978_1), .B(w_mem_inst__abc_21378_n2979_1), .Y(w_mem_inst__abc_21378_n2980) );
  OR2X2 OR2X2_2462 ( .A(w_mem_inst__abc_21378_n2980), .B(w_mem_inst__abc_21378_n2977), .Y(w_mem_inst__abc_21378_n2981) );
  OR2X2 OR2X2_2463 ( .A(w_mem_inst__abc_21378_n2981), .B(w_mem_inst__abc_21378_n2975_1), .Y(w_mem_inst__abc_21378_n2982_1) );
  OR2X2 OR2X2_2464 ( .A(w_mem_inst__abc_21378_n2983_1), .B(w_mem_inst__abc_21378_n2984), .Y(w_mem_inst__abc_21378_n2985) );
  OR2X2 OR2X2_2465 ( .A(w_mem_inst__abc_21378_n2987_1), .B(w_mem_inst__abc_21378_n2986_1), .Y(w_mem_inst__abc_21378_n2988) );
  OR2X2 OR2X2_2466 ( .A(w_mem_inst__abc_21378_n2985), .B(w_mem_inst__abc_21378_n2988), .Y(w_mem_inst__abc_21378_n2989) );
  OR2X2 OR2X2_2467 ( .A(w_mem_inst__abc_21378_n2990_1), .B(w_mem_inst__abc_21378_n2991_1), .Y(w_mem_inst__abc_21378_n2992) );
  OR2X2 OR2X2_2468 ( .A(w_mem_inst__abc_21378_n2993), .B(w_mem_inst__abc_21378_n2994_1), .Y(w_mem_inst__abc_21378_n2995_1) );
  OR2X2 OR2X2_2469 ( .A(w_mem_inst__abc_21378_n2995_1), .B(w_mem_inst__abc_21378_n2992), .Y(w_mem_inst__abc_21378_n2996) );
  OR2X2 OR2X2_247 ( .A(_auto_iopadmap_cc_313_execute_26059_61_), .B(d_reg_29_), .Y(_abc_15724_n1467) );
  OR2X2 OR2X2_2470 ( .A(w_mem_inst__abc_21378_n2998_1), .B(w_mem_inst__abc_21378_n2997), .Y(w_mem_inst__abc_21378_n2999_1) );
  OR2X2 OR2X2_2471 ( .A(w_mem_inst__abc_21378_n3000), .B(w_mem_inst__abc_21378_n3001), .Y(w_mem_inst__abc_21378_n3002_1) );
  OR2X2 OR2X2_2472 ( .A(w_mem_inst__abc_21378_n3002_1), .B(w_mem_inst__abc_21378_n2999_1), .Y(w_mem_inst__abc_21378_n3003_1) );
  OR2X2 OR2X2_2473 ( .A(w_mem_inst__abc_21378_n2996), .B(w_mem_inst__abc_21378_n3003_1), .Y(w_mem_inst__abc_21378_n3004) );
  OR2X2 OR2X2_2474 ( .A(w_mem_inst__abc_21378_n3004), .B(w_mem_inst__abc_21378_n2989), .Y(w_mem_inst__abc_21378_n3005) );
  OR2X2 OR2X2_2475 ( .A(w_mem_inst__abc_21378_n3005), .B(w_mem_inst__abc_21378_n2982_1), .Y(w_mem_inst__abc_21378_n3006_1) );
  OR2X2 OR2X2_2476 ( .A(w_mem_inst__abc_21378_n3008), .B(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_21378_n3009) );
  OR2X2 OR2X2_2477 ( .A(w_mem_inst__abc_21378_n3010_1), .B(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_21378_n3011_1) );
  OR2X2 OR2X2_2478 ( .A(w_mem_inst_w_mem_2__28_), .B(w_mem_inst_w_mem_0__28_), .Y(w_mem_inst__abc_21378_n3014_1) );
  OR2X2 OR2X2_2479 ( .A(w_mem_inst__abc_21378_n3013), .B(w_mem_inst__abc_21378_n3017), .Y(w_mem_inst__abc_21378_n3018_1) );
  OR2X2 OR2X2_248 ( .A(_abc_15724_n1472_1), .B(_abc_15724_n1452), .Y(_abc_15724_n1473_1) );
  OR2X2 OR2X2_2480 ( .A(w_mem_inst__abc_21378_n3019_1), .B(w_mem_inst__abc_21378_n3012), .Y(w_mem_inst__abc_21378_n3020) );
  OR2X2 OR2X2_2481 ( .A(w_mem_inst__abc_21378_n3021), .B(w_mem_inst__abc_21378_n1587_bF_buf0), .Y(w_mem_inst__abc_21378_n3022_1) );
  OR2X2 OR2X2_2482 ( .A(w_mem_inst__abc_21378_n3024), .B(w_mem_inst__abc_21378_n1586_bF_buf4), .Y(w_mem_inst__abc_21378_n3025) );
  OR2X2 OR2X2_2483 ( .A(w_mem_inst__abc_21378_n3026_1), .B(w_mem_inst__abc_21378_n3027_1), .Y(w_mem_inst__abc_21378_n3028) );
  OR2X2 OR2X2_2484 ( .A(w_mem_inst__abc_21378_n3028), .B(w_mem_inst__abc_21378_n3025), .Y(w_mem_inst__abc_21378_n3029) );
  OR2X2 OR2X2_2485 ( .A(w_mem_inst__abc_21378_n3029), .B(w_mem_inst__abc_21378_n3023_1), .Y(w_mem_inst__abc_21378_n3030_1) );
  OR2X2 OR2X2_2486 ( .A(w_mem_inst__abc_21378_n3031_1), .B(w_mem_inst__abc_21378_n3032), .Y(w_mem_inst__abc_21378_n3033) );
  OR2X2 OR2X2_2487 ( .A(w_mem_inst__abc_21378_n3035_1), .B(w_mem_inst__abc_21378_n3034_1), .Y(w_mem_inst__abc_21378_n3036) );
  OR2X2 OR2X2_2488 ( .A(w_mem_inst__abc_21378_n3033), .B(w_mem_inst__abc_21378_n3036), .Y(w_mem_inst__abc_21378_n3037) );
  OR2X2 OR2X2_2489 ( .A(w_mem_inst__abc_21378_n3038_1), .B(w_mem_inst__abc_21378_n3039_1), .Y(w_mem_inst__abc_21378_n3040) );
  OR2X2 OR2X2_249 ( .A(_abc_15724_n1475), .B(_abc_15724_n850_bF_buf5), .Y(_abc_15724_n1476) );
  OR2X2 OR2X2_2490 ( .A(w_mem_inst__abc_21378_n3041), .B(w_mem_inst__abc_21378_n3042_1), .Y(w_mem_inst__abc_21378_n3043_1) );
  OR2X2 OR2X2_2491 ( .A(w_mem_inst__abc_21378_n3040), .B(w_mem_inst__abc_21378_n3043_1), .Y(w_mem_inst__abc_21378_n3044) );
  OR2X2 OR2X2_2492 ( .A(w_mem_inst__abc_21378_n3045), .B(w_mem_inst__abc_21378_n3046_1), .Y(w_mem_inst__abc_21378_n3047_1) );
  OR2X2 OR2X2_2493 ( .A(w_mem_inst__abc_21378_n3048), .B(w_mem_inst__abc_21378_n3049), .Y(w_mem_inst__abc_21378_n3050_1) );
  OR2X2 OR2X2_2494 ( .A(w_mem_inst__abc_21378_n3047_1), .B(w_mem_inst__abc_21378_n3050_1), .Y(w_mem_inst__abc_21378_n3051_1) );
  OR2X2 OR2X2_2495 ( .A(w_mem_inst__abc_21378_n3051_1), .B(w_mem_inst__abc_21378_n3044), .Y(w_mem_inst__abc_21378_n3052) );
  OR2X2 OR2X2_2496 ( .A(w_mem_inst__abc_21378_n3052), .B(w_mem_inst__abc_21378_n3037), .Y(w_mem_inst__abc_21378_n3053) );
  OR2X2 OR2X2_2497 ( .A(w_mem_inst__abc_21378_n3053), .B(w_mem_inst__abc_21378_n3030_1), .Y(w_mem_inst__abc_21378_n3054_1) );
  OR2X2 OR2X2_2498 ( .A(w_mem_inst__abc_21378_n3056), .B(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_21378_n3057) );
  OR2X2 OR2X2_2499 ( .A(w_mem_inst__abc_21378_n3058_1), .B(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_21378_n3059_1) );
  OR2X2 OR2X2_25 ( .A(e_reg_3_), .B(_auto_iopadmap_cc_313_execute_26059_3_), .Y(_abc_15724_n788) );
  OR2X2 OR2X2_250 ( .A(_abc_15724_n1476), .B(_abc_15724_n1471), .Y(_abc_15724_n1477) );
  OR2X2 OR2X2_2500 ( .A(w_mem_inst_w_mem_2__29_), .B(w_mem_inst_w_mem_0__29_), .Y(w_mem_inst__abc_21378_n3062_1) );
  OR2X2 OR2X2_2501 ( .A(w_mem_inst__abc_21378_n3061), .B(w_mem_inst__abc_21378_n3065), .Y(w_mem_inst__abc_21378_n3066_1) );
  OR2X2 OR2X2_2502 ( .A(w_mem_inst__abc_21378_n3067_1), .B(w_mem_inst__abc_21378_n3060), .Y(w_mem_inst__abc_21378_n3068) );
  OR2X2 OR2X2_2503 ( .A(w_mem_inst__abc_21378_n3069), .B(w_mem_inst__abc_21378_n1587_bF_buf4), .Y(w_mem_inst__abc_21378_n3070_1) );
  OR2X2 OR2X2_2504 ( .A(w_mem_inst__abc_21378_n3072), .B(w_mem_inst__abc_21378_n1586_bF_buf3), .Y(w_mem_inst__abc_21378_n3073) );
  OR2X2 OR2X2_2505 ( .A(w_mem_inst__abc_21378_n3074_1), .B(w_mem_inst__abc_21378_n3075_1), .Y(w_mem_inst__abc_21378_n3076) );
  OR2X2 OR2X2_2506 ( .A(w_mem_inst__abc_21378_n3076), .B(w_mem_inst__abc_21378_n3073), .Y(w_mem_inst__abc_21378_n3077) );
  OR2X2 OR2X2_2507 ( .A(w_mem_inst__abc_21378_n3077), .B(w_mem_inst__abc_21378_n3071_1), .Y(w_mem_inst__abc_21378_n3078_1) );
  OR2X2 OR2X2_2508 ( .A(w_mem_inst__abc_21378_n3079_1), .B(w_mem_inst__abc_21378_n3080), .Y(w_mem_inst__abc_21378_n3081) );
  OR2X2 OR2X2_2509 ( .A(w_mem_inst__abc_21378_n3083_1), .B(w_mem_inst__abc_21378_n3082_1), .Y(w_mem_inst__abc_21378_n3084) );
  OR2X2 OR2X2_251 ( .A(_auto_iopadmap_cc_313_execute_26059_62_), .B(d_reg_30_), .Y(_abc_15724_n1482) );
  OR2X2 OR2X2_2510 ( .A(w_mem_inst__abc_21378_n3081), .B(w_mem_inst__abc_21378_n3084), .Y(w_mem_inst__abc_21378_n3085) );
  OR2X2 OR2X2_2511 ( .A(w_mem_inst__abc_21378_n3086_1), .B(w_mem_inst__abc_21378_n3087_1), .Y(w_mem_inst__abc_21378_n3088) );
  OR2X2 OR2X2_2512 ( .A(w_mem_inst__abc_21378_n3089), .B(w_mem_inst__abc_21378_n3090_1), .Y(w_mem_inst__abc_21378_n3091_1) );
  OR2X2 OR2X2_2513 ( .A(w_mem_inst__abc_21378_n3091_1), .B(w_mem_inst__abc_21378_n3088), .Y(w_mem_inst__abc_21378_n3092) );
  OR2X2 OR2X2_2514 ( .A(w_mem_inst__abc_21378_n3094_1), .B(w_mem_inst__abc_21378_n3093), .Y(w_mem_inst__abc_21378_n3095_1) );
  OR2X2 OR2X2_2515 ( .A(w_mem_inst__abc_21378_n3096), .B(w_mem_inst__abc_21378_n3097), .Y(w_mem_inst__abc_21378_n3098_1) );
  OR2X2 OR2X2_2516 ( .A(w_mem_inst__abc_21378_n3098_1), .B(w_mem_inst__abc_21378_n3095_1), .Y(w_mem_inst__abc_21378_n3099_1) );
  OR2X2 OR2X2_2517 ( .A(w_mem_inst__abc_21378_n3092), .B(w_mem_inst__abc_21378_n3099_1), .Y(w_mem_inst__abc_21378_n3100) );
  OR2X2 OR2X2_2518 ( .A(w_mem_inst__abc_21378_n3100), .B(w_mem_inst__abc_21378_n3085), .Y(w_mem_inst__abc_21378_n3101) );
  OR2X2 OR2X2_2519 ( .A(w_mem_inst__abc_21378_n3101), .B(w_mem_inst__abc_21378_n3078_1), .Y(w_mem_inst__abc_21378_n3102_1) );
  OR2X2 OR2X2_252 ( .A(_abc_15724_n1466), .B(_abc_15724_n1485_1), .Y(_abc_15724_n1486) );
  OR2X2 OR2X2_2520 ( .A(w_mem_inst__abc_21378_n3104), .B(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_21378_n3105) );
  OR2X2 OR2X2_2521 ( .A(w_mem_inst__abc_21378_n3106_1), .B(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_21378_n3107_1) );
  OR2X2 OR2X2_2522 ( .A(w_mem_inst_w_mem_2__30_), .B(w_mem_inst_w_mem_0__30_), .Y(w_mem_inst__abc_21378_n3110_1) );
  OR2X2 OR2X2_2523 ( .A(w_mem_inst__abc_21378_n3109), .B(w_mem_inst__abc_21378_n3113), .Y(w_mem_inst__abc_21378_n3114_1) );
  OR2X2 OR2X2_2524 ( .A(w_mem_inst__abc_21378_n3115_1), .B(w_mem_inst__abc_21378_n3108), .Y(w_mem_inst__abc_21378_n3116) );
  OR2X2 OR2X2_2525 ( .A(w_mem_inst__abc_21378_n3117), .B(w_mem_inst__abc_21378_n1587_bF_buf3), .Y(w_mem_inst__abc_21378_n3118_1) );
  OR2X2 OR2X2_2526 ( .A(w_mem_inst__abc_21378_n3120), .B(w_mem_inst__abc_21378_n1586_bF_buf2), .Y(w_mem_inst__abc_21378_n3121) );
  OR2X2 OR2X2_2527 ( .A(w_mem_inst__abc_21378_n3122_1), .B(w_mem_inst__abc_21378_n3123_1), .Y(w_mem_inst__abc_21378_n3124) );
  OR2X2 OR2X2_2528 ( .A(w_mem_inst__abc_21378_n3124), .B(w_mem_inst__abc_21378_n3121), .Y(w_mem_inst__abc_21378_n3125) );
  OR2X2 OR2X2_2529 ( .A(w_mem_inst__abc_21378_n3125), .B(w_mem_inst__abc_21378_n3119_1), .Y(w_mem_inst__abc_21378_n3126_1) );
  OR2X2 OR2X2_253 ( .A(_abc_15724_n1487_1), .B(_abc_15724_n1484_1), .Y(_abc_15724_n1488) );
  OR2X2 OR2X2_2530 ( .A(w_mem_inst__abc_21378_n3127_1), .B(w_mem_inst__abc_21378_n3128), .Y(w_mem_inst__abc_21378_n3129) );
  OR2X2 OR2X2_2531 ( .A(w_mem_inst__abc_21378_n3131_1), .B(w_mem_inst__abc_21378_n3130_1), .Y(w_mem_inst__abc_21378_n3132) );
  OR2X2 OR2X2_2532 ( .A(w_mem_inst__abc_21378_n3129), .B(w_mem_inst__abc_21378_n3132), .Y(w_mem_inst__abc_21378_n3133) );
  OR2X2 OR2X2_2533 ( .A(w_mem_inst__abc_21378_n3134_1), .B(w_mem_inst__abc_21378_n3135_1), .Y(w_mem_inst__abc_21378_n3136) );
  OR2X2 OR2X2_2534 ( .A(w_mem_inst__abc_21378_n3137), .B(w_mem_inst__abc_21378_n3138_1), .Y(w_mem_inst__abc_21378_n3139_1) );
  OR2X2 OR2X2_2535 ( .A(w_mem_inst__abc_21378_n3136), .B(w_mem_inst__abc_21378_n3139_1), .Y(w_mem_inst__abc_21378_n3140) );
  OR2X2 OR2X2_2536 ( .A(w_mem_inst__abc_21378_n3141), .B(w_mem_inst__abc_21378_n3142_1), .Y(w_mem_inst__abc_21378_n3143_1) );
  OR2X2 OR2X2_2537 ( .A(w_mem_inst__abc_21378_n3144), .B(w_mem_inst__abc_21378_n3145), .Y(w_mem_inst__abc_21378_n3146_1) );
  OR2X2 OR2X2_2538 ( .A(w_mem_inst__abc_21378_n3143_1), .B(w_mem_inst__abc_21378_n3146_1), .Y(w_mem_inst__abc_21378_n3147_1) );
  OR2X2 OR2X2_2539 ( .A(w_mem_inst__abc_21378_n3147_1), .B(w_mem_inst__abc_21378_n3140), .Y(w_mem_inst__abc_21378_n3148) );
  OR2X2 OR2X2_254 ( .A(_abc_15724_n1489), .B(_abc_15724_n1468), .Y(_abc_15724_n1490) );
  OR2X2 OR2X2_2540 ( .A(w_mem_inst__abc_21378_n3148), .B(w_mem_inst__abc_21378_n3133), .Y(w_mem_inst__abc_21378_n3149) );
  OR2X2 OR2X2_2541 ( .A(w_mem_inst__abc_21378_n3149), .B(w_mem_inst__abc_21378_n3126_1), .Y(w_mem_inst__abc_21378_n3150_1) );
  OR2X2 OR2X2_2542 ( .A(w_mem_inst__abc_21378_n3157), .B(w_mem_inst__abc_21378_n3155_1), .Y(w_mem_inst__abc_21378_n3158_1) );
  OR2X2 OR2X2_2543 ( .A(w_mem_inst__abc_21378_n3153), .B(w_mem_inst__abc_21378_n3159_1), .Y(w_mem_inst__0w_mem_15__31_0__0_) );
  OR2X2 OR2X2_2544 ( .A(w_mem_inst__abc_21378_n3163_1), .B(w_mem_inst__abc_21378_n3162_1), .Y(w_mem_inst__abc_21378_n3164) );
  OR2X2 OR2X2_2545 ( .A(w_mem_inst__abc_21378_n3161), .B(w_mem_inst__abc_21378_n3165), .Y(w_mem_inst__0w_mem_15__31_0__1_) );
  OR2X2 OR2X2_2546 ( .A(w_mem_inst__abc_21378_n3168), .B(w_mem_inst__abc_21378_n3167_1), .Y(w_mem_inst__abc_21378_n3169) );
  OR2X2 OR2X2_2547 ( .A(w_mem_inst__abc_21378_n3152_bF_buf60), .B(w_mem_inst__abc_21378_n3169), .Y(w_mem_inst__abc_21378_n3170_1) );
  OR2X2 OR2X2_2548 ( .A(w_mem_inst__abc_21378_n1725), .B(w_mem_inst__abc_21378_n3154_1_bF_buf61), .Y(w_mem_inst__abc_21378_n3171_1) );
  OR2X2 OR2X2_2549 ( .A(w_mem_inst__abc_21378_n3175_1), .B(w_mem_inst__abc_21378_n3174_1), .Y(w_mem_inst__abc_21378_n3176) );
  OR2X2 OR2X2_255 ( .A(_abc_15724_n1490), .B(_abc_15724_n1483), .Y(_abc_15724_n1491) );
  OR2X2 OR2X2_2550 ( .A(w_mem_inst__abc_21378_n3173), .B(w_mem_inst__abc_21378_n3177), .Y(w_mem_inst__0w_mem_15__31_0__3_) );
  OR2X2 OR2X2_2551 ( .A(w_mem_inst__abc_21378_n3180), .B(w_mem_inst__abc_21378_n3179_1), .Y(w_mem_inst__abc_21378_n3181) );
  OR2X2 OR2X2_2552 ( .A(w_mem_inst__abc_21378_n3152_bF_buf58), .B(w_mem_inst__abc_21378_n3181), .Y(w_mem_inst__abc_21378_n3182_1) );
  OR2X2 OR2X2_2553 ( .A(w_mem_inst__abc_21378_n1821), .B(w_mem_inst__abc_21378_n3154_1_bF_buf59), .Y(w_mem_inst__abc_21378_n3183_1) );
  OR2X2 OR2X2_2554 ( .A(w_mem_inst__abc_21378_n3187_1), .B(w_mem_inst__abc_21378_n3186_1), .Y(w_mem_inst__abc_21378_n3188) );
  OR2X2 OR2X2_2555 ( .A(w_mem_inst__abc_21378_n3185), .B(w_mem_inst__abc_21378_n3189), .Y(w_mem_inst__0w_mem_15__31_0__5_) );
  OR2X2 OR2X2_2556 ( .A(w_mem_inst__abc_21378_n3193), .B(w_mem_inst__abc_21378_n3192), .Y(w_mem_inst__abc_21378_n3194_1) );
  OR2X2 OR2X2_2557 ( .A(w_mem_inst__abc_21378_n3191_1), .B(w_mem_inst__abc_21378_n3195_1), .Y(w_mem_inst__0w_mem_15__31_0__6_) );
  OR2X2 OR2X2_2558 ( .A(w_mem_inst__abc_21378_n3199_1), .B(w_mem_inst__abc_21378_n3198_1), .Y(w_mem_inst__abc_21378_n3200) );
  OR2X2 OR2X2_2559 ( .A(w_mem_inst__abc_21378_n3197), .B(w_mem_inst__abc_21378_n3201), .Y(w_mem_inst__0w_mem_15__31_0__7_) );
  OR2X2 OR2X2_256 ( .A(_abc_15724_n1493_1), .B(_abc_15724_n1479), .Y(H3_reg_30__FF_INPUT) );
  OR2X2 OR2X2_2560 ( .A(w_mem_inst__abc_21378_n3205), .B(w_mem_inst__abc_21378_n3204), .Y(w_mem_inst__abc_21378_n3206_1) );
  OR2X2 OR2X2_2561 ( .A(w_mem_inst__abc_21378_n3203_1), .B(w_mem_inst__abc_21378_n3207_1), .Y(w_mem_inst__0w_mem_15__31_0__8_) );
  OR2X2 OR2X2_2562 ( .A(w_mem_inst__abc_21378_n3211_1), .B(w_mem_inst__abc_21378_n3210_1), .Y(w_mem_inst__abc_21378_n3212) );
  OR2X2 OR2X2_2563 ( .A(w_mem_inst__abc_21378_n3209), .B(w_mem_inst__abc_21378_n3213), .Y(w_mem_inst__0w_mem_15__31_0__9_) );
  OR2X2 OR2X2_2564 ( .A(w_mem_inst__abc_21378_n3216), .B(w_mem_inst__abc_21378_n3215_1), .Y(w_mem_inst__abc_21378_n3217) );
  OR2X2 OR2X2_2565 ( .A(w_mem_inst__abc_21378_n3152_bF_buf52), .B(w_mem_inst__abc_21378_n3217), .Y(w_mem_inst__abc_21378_n3218_1) );
  OR2X2 OR2X2_2566 ( .A(w_mem_inst__abc_21378_n2109), .B(w_mem_inst__abc_21378_n3154_1_bF_buf53), .Y(w_mem_inst__abc_21378_n3219_1) );
  OR2X2 OR2X2_2567 ( .A(w_mem_inst__abc_21378_n3222_1), .B(w_mem_inst__abc_21378_n3221), .Y(w_mem_inst__abc_21378_n3223_1) );
  OR2X2 OR2X2_2568 ( .A(w_mem_inst__abc_21378_n3152_bF_buf51), .B(w_mem_inst__abc_21378_n3223_1), .Y(w_mem_inst__abc_21378_n3224) );
  OR2X2 OR2X2_2569 ( .A(w_mem_inst__abc_21378_n2157), .B(w_mem_inst__abc_21378_n3154_1_bF_buf52), .Y(w_mem_inst__abc_21378_n3225) );
  OR2X2 OR2X2_257 ( .A(_auto_iopadmap_cc_313_execute_26059_63_), .B(d_reg_31_), .Y(_abc_15724_n1496_1) );
  OR2X2 OR2X2_2570 ( .A(w_mem_inst__abc_21378_n3228), .B(w_mem_inst__abc_21378_n3227_1), .Y(w_mem_inst__abc_21378_n3229) );
  OR2X2 OR2X2_2571 ( .A(w_mem_inst__abc_21378_n3152_bF_buf50), .B(w_mem_inst__abc_21378_n3229), .Y(w_mem_inst__abc_21378_n3230_1) );
  OR2X2 OR2X2_2572 ( .A(w_mem_inst__abc_21378_n2205), .B(w_mem_inst__abc_21378_n3154_1_bF_buf51), .Y(w_mem_inst__abc_21378_n3231_1) );
  OR2X2 OR2X2_2573 ( .A(w_mem_inst__abc_21378_n3235_1), .B(w_mem_inst__abc_21378_n3234_1), .Y(w_mem_inst__abc_21378_n3236) );
  OR2X2 OR2X2_2574 ( .A(w_mem_inst__abc_21378_n3233), .B(w_mem_inst__abc_21378_n3237), .Y(w_mem_inst__0w_mem_15__31_0__13_) );
  OR2X2 OR2X2_2575 ( .A(w_mem_inst__abc_21378_n3241), .B(w_mem_inst__abc_21378_n3240), .Y(w_mem_inst__abc_21378_n3242_1) );
  OR2X2 OR2X2_2576 ( .A(w_mem_inst__abc_21378_n3239_1), .B(w_mem_inst__abc_21378_n3243_1), .Y(w_mem_inst__0w_mem_15__31_0__14_) );
  OR2X2 OR2X2_2577 ( .A(w_mem_inst__abc_21378_n3247_1), .B(w_mem_inst__abc_21378_n3246_1), .Y(w_mem_inst__abc_21378_n3248) );
  OR2X2 OR2X2_2578 ( .A(w_mem_inst__abc_21378_n3245), .B(w_mem_inst__abc_21378_n3249), .Y(w_mem_inst__0w_mem_15__31_0__15_) );
  OR2X2 OR2X2_2579 ( .A(w_mem_inst__abc_21378_n3253), .B(w_mem_inst__abc_21378_n3252), .Y(w_mem_inst__abc_21378_n3254_1) );
  OR2X2 OR2X2_258 ( .A(_abc_15724_n1501), .B(_abc_15724_n1480), .Y(_abc_15724_n1502) );
  OR2X2 OR2X2_2580 ( .A(w_mem_inst__abc_21378_n3251_1), .B(w_mem_inst__abc_21378_n3255_1), .Y(w_mem_inst__0w_mem_15__31_0__16_) );
  OR2X2 OR2X2_2581 ( .A(w_mem_inst__abc_21378_n3259_1), .B(w_mem_inst__abc_21378_n3258_1), .Y(w_mem_inst__abc_21378_n3260) );
  OR2X2 OR2X2_2582 ( .A(w_mem_inst__abc_21378_n3257), .B(w_mem_inst__abc_21378_n3261), .Y(w_mem_inst__0w_mem_15__31_0__17_) );
  OR2X2 OR2X2_2583 ( .A(w_mem_inst__abc_21378_n3264), .B(w_mem_inst__abc_21378_n3263_1), .Y(w_mem_inst__abc_21378_n3265) );
  OR2X2 OR2X2_2584 ( .A(w_mem_inst__abc_21378_n3152_bF_buf44), .B(w_mem_inst__abc_21378_n3265), .Y(w_mem_inst__abc_21378_n3266_1) );
  OR2X2 OR2X2_2585 ( .A(w_mem_inst__abc_21378_n2493), .B(w_mem_inst__abc_21378_n3154_1_bF_buf45), .Y(w_mem_inst__abc_21378_n3267_1) );
  OR2X2 OR2X2_2586 ( .A(w_mem_inst__abc_21378_n3271_1), .B(w_mem_inst__abc_21378_n3270_1), .Y(w_mem_inst__abc_21378_n3272) );
  OR2X2 OR2X2_2587 ( .A(w_mem_inst__abc_21378_n3269), .B(w_mem_inst__abc_21378_n3273), .Y(w_mem_inst__0w_mem_15__31_0__19_) );
  OR2X2 OR2X2_2588 ( .A(w_mem_inst__abc_21378_n3277), .B(w_mem_inst__abc_21378_n3276), .Y(w_mem_inst__abc_21378_n3278_1) );
  OR2X2 OR2X2_2589 ( .A(w_mem_inst__abc_21378_n3275_1), .B(w_mem_inst__abc_21378_n3279_1), .Y(w_mem_inst__0w_mem_15__31_0__20_) );
  OR2X2 OR2X2_259 ( .A(_abc_15724_n1500), .B(_abc_15724_n1504), .Y(_abc_15724_n1505) );
  OR2X2 OR2X2_2590 ( .A(w_mem_inst__abc_21378_n3283_1), .B(w_mem_inst__abc_21378_n3282_1), .Y(w_mem_inst__abc_21378_n3284) );
  OR2X2 OR2X2_2591 ( .A(w_mem_inst__abc_21378_n3281), .B(w_mem_inst__abc_21378_n3285), .Y(w_mem_inst__0w_mem_15__31_0__21_) );
  OR2X2 OR2X2_2592 ( .A(w_mem_inst__abc_21378_n3289), .B(w_mem_inst__abc_21378_n3288), .Y(w_mem_inst__abc_21378_n3290_1) );
  OR2X2 OR2X2_2593 ( .A(w_mem_inst__abc_21378_n3287_1), .B(w_mem_inst__abc_21378_n3291_1), .Y(w_mem_inst__0w_mem_15__31_0__22_) );
  OR2X2 OR2X2_2594 ( .A(w_mem_inst__abc_21378_n3295_1), .B(w_mem_inst__abc_21378_n3294_1), .Y(w_mem_inst__abc_21378_n3296) );
  OR2X2 OR2X2_2595 ( .A(w_mem_inst__abc_21378_n3293), .B(w_mem_inst__abc_21378_n3297), .Y(w_mem_inst__0w_mem_15__31_0__23_) );
  OR2X2 OR2X2_2596 ( .A(w_mem_inst__abc_21378_n3301), .B(w_mem_inst__abc_21378_n3300), .Y(w_mem_inst__abc_21378_n3302_1) );
  OR2X2 OR2X2_2597 ( .A(w_mem_inst__abc_21378_n3299_1), .B(w_mem_inst__abc_21378_n3303_1), .Y(w_mem_inst__0w_mem_15__31_0__24_) );
  OR2X2 OR2X2_2598 ( .A(w_mem_inst__abc_21378_n3306_1), .B(w_mem_inst__abc_21378_n3305), .Y(w_mem_inst__abc_21378_n3307_1) );
  OR2X2 OR2X2_2599 ( .A(w_mem_inst__abc_21378_n3152_bF_buf37), .B(w_mem_inst__abc_21378_n3307_1), .Y(w_mem_inst__abc_21378_n3308) );
  OR2X2 OR2X2_26 ( .A(e_reg_1_), .B(_auto_iopadmap_cc_313_execute_26059_1_), .Y(_abc_15724_n793) );
  OR2X2 OR2X2_260 ( .A(_abc_15724_n1506), .B(_abc_15724_n1507), .Y(H3_reg_31__FF_INPUT) );
  OR2X2 OR2X2_2600 ( .A(w_mem_inst__abc_21378_n2829), .B(w_mem_inst__abc_21378_n3154_1_bF_buf38), .Y(w_mem_inst__abc_21378_n3309) );
  OR2X2 OR2X2_2601 ( .A(w_mem_inst__abc_21378_n3312), .B(w_mem_inst__abc_21378_n3311_1), .Y(w_mem_inst__abc_21378_n3313) );
  OR2X2 OR2X2_2602 ( .A(w_mem_inst__abc_21378_n3152_bF_buf36), .B(w_mem_inst__abc_21378_n3313), .Y(w_mem_inst__abc_21378_n3314_1) );
  OR2X2 OR2X2_2603 ( .A(w_mem_inst__abc_21378_n2877), .B(w_mem_inst__abc_21378_n3154_1_bF_buf37), .Y(w_mem_inst__abc_21378_n3315_1) );
  OR2X2 OR2X2_2604 ( .A(w_mem_inst__abc_21378_n3318_1), .B(w_mem_inst__abc_21378_n3317), .Y(w_mem_inst__abc_21378_n3319_1) );
  OR2X2 OR2X2_2605 ( .A(w_mem_inst__abc_21378_n3152_bF_buf35), .B(w_mem_inst__abc_21378_n3319_1), .Y(w_mem_inst__abc_21378_n3320) );
  OR2X2 OR2X2_2606 ( .A(w_mem_inst__abc_21378_n2925), .B(w_mem_inst__abc_21378_n3154_1_bF_buf36), .Y(w_mem_inst__abc_21378_n3321) );
  OR2X2 OR2X2_2607 ( .A(w_mem_inst__abc_21378_n3324), .B(w_mem_inst__abc_21378_n3323_1), .Y(w_mem_inst__abc_21378_n3325) );
  OR2X2 OR2X2_2608 ( .A(w_mem_inst__abc_21378_n3152_bF_buf34), .B(w_mem_inst__abc_21378_n3325), .Y(w_mem_inst__abc_21378_n3326_1) );
  OR2X2 OR2X2_2609 ( .A(w_mem_inst__abc_21378_n2973), .B(w_mem_inst__abc_21378_n3154_1_bF_buf35), .Y(w_mem_inst__abc_21378_n3327_1) );
  OR2X2 OR2X2_261 ( .A(_auto_iopadmap_cc_313_execute_26059_64_), .B(c_reg_0_), .Y(_abc_15724_n1509_1) );
  OR2X2 OR2X2_2610 ( .A(w_mem_inst__abc_21378_n3331_1), .B(w_mem_inst__abc_21378_n3330_1), .Y(w_mem_inst__abc_21378_n3332) );
  OR2X2 OR2X2_2611 ( .A(w_mem_inst__abc_21378_n3329), .B(w_mem_inst__abc_21378_n3333), .Y(w_mem_inst__0w_mem_15__31_0__29_) );
  OR2X2 OR2X2_2612 ( .A(w_mem_inst__abc_21378_n3337), .B(w_mem_inst__abc_21378_n3336), .Y(w_mem_inst__abc_21378_n3338_1) );
  OR2X2 OR2X2_2613 ( .A(w_mem_inst__abc_21378_n3335_1), .B(w_mem_inst__abc_21378_n3339_1), .Y(w_mem_inst__0w_mem_15__31_0__30_) );
  OR2X2 OR2X2_2614 ( .A(w_mem_inst__abc_21378_n3343_1), .B(w_mem_inst__abc_21378_n3342_1), .Y(w_mem_inst__abc_21378_n3344) );
  OR2X2 OR2X2_2615 ( .A(w_mem_inst__abc_21378_n3341), .B(w_mem_inst__abc_21378_n3345), .Y(w_mem_inst__0w_mem_15__31_0__31_) );
  OR2X2 OR2X2_2616 ( .A(w_mem_inst__abc_21378_n3351_1), .B(w_mem_inst__abc_21378_n3349), .Y(w_mem_inst__abc_21378_n3352) );
  OR2X2 OR2X2_2617 ( .A(w_mem_inst__abc_21378_n3352), .B(w_mem_inst__abc_21378_n3348), .Y(w_mem_inst__0w_mem_14__31_0__0_) );
  OR2X2 OR2X2_2618 ( .A(w_mem_inst__abc_21378_n3357), .B(w_mem_inst__abc_21378_n3355_1), .Y(w_mem_inst__abc_21378_n3358_1) );
  OR2X2 OR2X2_2619 ( .A(w_mem_inst__abc_21378_n3358_1), .B(w_mem_inst__abc_21378_n3354_1), .Y(w_mem_inst__0w_mem_14__31_0__1_) );
  OR2X2 OR2X2_262 ( .A(_abc_15724_n1512), .B(_abc_15724_n850_bF_buf4), .Y(_abc_15724_n1513) );
  OR2X2 OR2X2_2620 ( .A(w_mem_inst__abc_21378_n3363_1), .B(w_mem_inst__abc_21378_n3361), .Y(w_mem_inst__abc_21378_n3364) );
  OR2X2 OR2X2_2621 ( .A(w_mem_inst__abc_21378_n3364), .B(w_mem_inst__abc_21378_n3360), .Y(w_mem_inst__0w_mem_14__31_0__2_) );
  OR2X2 OR2X2_2622 ( .A(w_mem_inst__abc_21378_n3369), .B(w_mem_inst__abc_21378_n3367_1), .Y(w_mem_inst__abc_21378_n3370_1) );
  OR2X2 OR2X2_2623 ( .A(w_mem_inst__abc_21378_n3370_1), .B(w_mem_inst__abc_21378_n3366_1), .Y(w_mem_inst__0w_mem_14__31_0__3_) );
  OR2X2 OR2X2_2624 ( .A(w_mem_inst__abc_21378_n3375_1), .B(w_mem_inst__abc_21378_n3373), .Y(w_mem_inst__abc_21378_n3376) );
  OR2X2 OR2X2_2625 ( .A(w_mem_inst__abc_21378_n3376), .B(w_mem_inst__abc_21378_n3372), .Y(w_mem_inst__0w_mem_14__31_0__4_) );
  OR2X2 OR2X2_2626 ( .A(w_mem_inst__abc_21378_n3381), .B(w_mem_inst__abc_21378_n3379_1), .Y(w_mem_inst__abc_21378_n3382_1) );
  OR2X2 OR2X2_2627 ( .A(w_mem_inst__abc_21378_n3382_1), .B(w_mem_inst__abc_21378_n3378_1), .Y(w_mem_inst__0w_mem_14__31_0__5_) );
  OR2X2 OR2X2_2628 ( .A(w_mem_inst__abc_21378_n3387_1), .B(w_mem_inst__abc_21378_n3385), .Y(w_mem_inst__abc_21378_n3388) );
  OR2X2 OR2X2_2629 ( .A(w_mem_inst__abc_21378_n3388), .B(w_mem_inst__abc_21378_n3384), .Y(w_mem_inst__0w_mem_14__31_0__6_) );
  OR2X2 OR2X2_263 ( .A(_abc_15724_n1514), .B(digest_update_bF_buf4), .Y(_abc_15724_n1515) );
  OR2X2 OR2X2_2630 ( .A(w_mem_inst__abc_21378_n3393), .B(w_mem_inst__abc_21378_n3391_1), .Y(w_mem_inst__abc_21378_n3394_1) );
  OR2X2 OR2X2_2631 ( .A(w_mem_inst__abc_21378_n3394_1), .B(w_mem_inst__abc_21378_n3390_1), .Y(w_mem_inst__0w_mem_14__31_0__7_) );
  OR2X2 OR2X2_2632 ( .A(w_mem_inst__abc_21378_n3399_1), .B(w_mem_inst__abc_21378_n3397), .Y(w_mem_inst__abc_21378_n3400) );
  OR2X2 OR2X2_2633 ( .A(w_mem_inst__abc_21378_n3400), .B(w_mem_inst__abc_21378_n3396), .Y(w_mem_inst__0w_mem_14__31_0__8_) );
  OR2X2 OR2X2_2634 ( .A(w_mem_inst__abc_21378_n3405), .B(w_mem_inst__abc_21378_n3403_1), .Y(w_mem_inst__abc_21378_n3406_1) );
  OR2X2 OR2X2_2635 ( .A(w_mem_inst__abc_21378_n3406_1), .B(w_mem_inst__abc_21378_n3402_1), .Y(w_mem_inst__0w_mem_14__31_0__9_) );
  OR2X2 OR2X2_2636 ( .A(w_mem_inst__abc_21378_n3411_1), .B(w_mem_inst__abc_21378_n3409), .Y(w_mem_inst__abc_21378_n3412) );
  OR2X2 OR2X2_2637 ( .A(w_mem_inst__abc_21378_n3412), .B(w_mem_inst__abc_21378_n3408), .Y(w_mem_inst__0w_mem_14__31_0__10_) );
  OR2X2 OR2X2_2638 ( .A(w_mem_inst__abc_21378_n3417), .B(w_mem_inst__abc_21378_n3415_1), .Y(w_mem_inst__abc_21378_n3418_1) );
  OR2X2 OR2X2_2639 ( .A(w_mem_inst__abc_21378_n3418_1), .B(w_mem_inst__abc_21378_n3414_1), .Y(w_mem_inst__0w_mem_14__31_0__11_) );
  OR2X2 OR2X2_264 ( .A(_auto_iopadmap_cc_313_execute_26059_65_), .B(c_reg_1_), .Y(_abc_15724_n1517) );
  OR2X2 OR2X2_2640 ( .A(w_mem_inst__abc_21378_n3423_1), .B(w_mem_inst__abc_21378_n3421), .Y(w_mem_inst__abc_21378_n3424) );
  OR2X2 OR2X2_2641 ( .A(w_mem_inst__abc_21378_n3424), .B(w_mem_inst__abc_21378_n3420), .Y(w_mem_inst__0w_mem_14__31_0__12_) );
  OR2X2 OR2X2_2642 ( .A(w_mem_inst__abc_21378_n3429), .B(w_mem_inst__abc_21378_n3427_1), .Y(w_mem_inst__abc_21378_n3430_1) );
  OR2X2 OR2X2_2643 ( .A(w_mem_inst__abc_21378_n3430_1), .B(w_mem_inst__abc_21378_n3426_1), .Y(w_mem_inst__0w_mem_14__31_0__13_) );
  OR2X2 OR2X2_2644 ( .A(w_mem_inst__abc_21378_n3435_1), .B(w_mem_inst__abc_21378_n3433), .Y(w_mem_inst__abc_21378_n3436) );
  OR2X2 OR2X2_2645 ( .A(w_mem_inst__abc_21378_n3436), .B(w_mem_inst__abc_21378_n3432), .Y(w_mem_inst__0w_mem_14__31_0__14_) );
  OR2X2 OR2X2_2646 ( .A(w_mem_inst__abc_21378_n3441), .B(w_mem_inst__abc_21378_n3439_1), .Y(w_mem_inst__abc_21378_n3442_1) );
  OR2X2 OR2X2_2647 ( .A(w_mem_inst__abc_21378_n3442_1), .B(w_mem_inst__abc_21378_n3438_1), .Y(w_mem_inst__0w_mem_14__31_0__15_) );
  OR2X2 OR2X2_2648 ( .A(w_mem_inst__abc_21378_n3447_1), .B(w_mem_inst__abc_21378_n3445), .Y(w_mem_inst__abc_21378_n3448) );
  OR2X2 OR2X2_2649 ( .A(w_mem_inst__abc_21378_n3448), .B(w_mem_inst__abc_21378_n3444), .Y(w_mem_inst__0w_mem_14__31_0__16_) );
  OR2X2 OR2X2_265 ( .A(_abc_15724_n1520_1), .B(_abc_15724_n1510_1), .Y(_abc_15724_n1523) );
  OR2X2 OR2X2_2650 ( .A(w_mem_inst__abc_21378_n3453), .B(w_mem_inst__abc_21378_n3451_1), .Y(w_mem_inst__abc_21378_n3454_1) );
  OR2X2 OR2X2_2651 ( .A(w_mem_inst__abc_21378_n3454_1), .B(w_mem_inst__abc_21378_n3450_1), .Y(w_mem_inst__0w_mem_14__31_0__17_) );
  OR2X2 OR2X2_2652 ( .A(w_mem_inst__abc_21378_n3459_1), .B(w_mem_inst__abc_21378_n3457), .Y(w_mem_inst__abc_21378_n3460) );
  OR2X2 OR2X2_2653 ( .A(w_mem_inst__abc_21378_n3460), .B(w_mem_inst__abc_21378_n3456), .Y(w_mem_inst__0w_mem_14__31_0__18_) );
  OR2X2 OR2X2_2654 ( .A(w_mem_inst__abc_21378_n3465), .B(w_mem_inst__abc_21378_n3463_1), .Y(w_mem_inst__abc_21378_n3466_1) );
  OR2X2 OR2X2_2655 ( .A(w_mem_inst__abc_21378_n3466_1), .B(w_mem_inst__abc_21378_n3462_1), .Y(w_mem_inst__0w_mem_14__31_0__19_) );
  OR2X2 OR2X2_2656 ( .A(w_mem_inst__abc_21378_n3471_1), .B(w_mem_inst__abc_21378_n3469), .Y(w_mem_inst__abc_21378_n3472) );
  OR2X2 OR2X2_2657 ( .A(w_mem_inst__abc_21378_n3472), .B(w_mem_inst__abc_21378_n3468), .Y(w_mem_inst__0w_mem_14__31_0__20_) );
  OR2X2 OR2X2_2658 ( .A(w_mem_inst__abc_21378_n3477), .B(w_mem_inst__abc_21378_n3475_1), .Y(w_mem_inst__abc_21378_n3478_1) );
  OR2X2 OR2X2_2659 ( .A(w_mem_inst__abc_21378_n3478_1), .B(w_mem_inst__abc_21378_n3474_1), .Y(w_mem_inst__0w_mem_14__31_0__21_) );
  OR2X2 OR2X2_266 ( .A(_abc_15724_n1524), .B(_abc_15724_n850_bF_buf3), .Y(_abc_15724_n1525) );
  OR2X2 OR2X2_2660 ( .A(w_mem_inst__abc_21378_n3483_1), .B(w_mem_inst__abc_21378_n3481), .Y(w_mem_inst__abc_21378_n3484) );
  OR2X2 OR2X2_2661 ( .A(w_mem_inst__abc_21378_n3484), .B(w_mem_inst__abc_21378_n3480), .Y(w_mem_inst__0w_mem_14__31_0__22_) );
  OR2X2 OR2X2_2662 ( .A(w_mem_inst__abc_21378_n3489), .B(w_mem_inst__abc_21378_n3487_1), .Y(w_mem_inst__abc_21378_n3490_1) );
  OR2X2 OR2X2_2663 ( .A(w_mem_inst__abc_21378_n3490_1), .B(w_mem_inst__abc_21378_n3486_1), .Y(w_mem_inst__0w_mem_14__31_0__23_) );
  OR2X2 OR2X2_2664 ( .A(w_mem_inst__abc_21378_n3495_1), .B(w_mem_inst__abc_21378_n3493), .Y(w_mem_inst__abc_21378_n3496) );
  OR2X2 OR2X2_2665 ( .A(w_mem_inst__abc_21378_n3496), .B(w_mem_inst__abc_21378_n3492), .Y(w_mem_inst__0w_mem_14__31_0__24_) );
  OR2X2 OR2X2_2666 ( .A(w_mem_inst__abc_21378_n3501), .B(w_mem_inst__abc_21378_n3499_1), .Y(w_mem_inst__abc_21378_n3502_1) );
  OR2X2 OR2X2_2667 ( .A(w_mem_inst__abc_21378_n3502_1), .B(w_mem_inst__abc_21378_n3498_1), .Y(w_mem_inst__0w_mem_14__31_0__25_) );
  OR2X2 OR2X2_2668 ( .A(w_mem_inst__abc_21378_n3507_1), .B(w_mem_inst__abc_21378_n3505), .Y(w_mem_inst__abc_21378_n3508) );
  OR2X2 OR2X2_2669 ( .A(w_mem_inst__abc_21378_n3508), .B(w_mem_inst__abc_21378_n3504), .Y(w_mem_inst__0w_mem_14__31_0__26_) );
  OR2X2 OR2X2_267 ( .A(_abc_15724_n851_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_65_), .Y(_abc_15724_n1526) );
  OR2X2 OR2X2_2670 ( .A(w_mem_inst__abc_21378_n3513), .B(w_mem_inst__abc_21378_n3511_1), .Y(w_mem_inst__abc_21378_n3514_1) );
  OR2X2 OR2X2_2671 ( .A(w_mem_inst__abc_21378_n3514_1), .B(w_mem_inst__abc_21378_n3510_1), .Y(w_mem_inst__0w_mem_14__31_0__27_) );
  OR2X2 OR2X2_2672 ( .A(w_mem_inst__abc_21378_n3519_1), .B(w_mem_inst__abc_21378_n3517), .Y(w_mem_inst__abc_21378_n3520) );
  OR2X2 OR2X2_2673 ( .A(w_mem_inst__abc_21378_n3520), .B(w_mem_inst__abc_21378_n3516), .Y(w_mem_inst__0w_mem_14__31_0__28_) );
  OR2X2 OR2X2_2674 ( .A(w_mem_inst__abc_21378_n3525), .B(w_mem_inst__abc_21378_n3523_1), .Y(w_mem_inst__abc_21378_n3526_1) );
  OR2X2 OR2X2_2675 ( .A(w_mem_inst__abc_21378_n3526_1), .B(w_mem_inst__abc_21378_n3522_1), .Y(w_mem_inst__0w_mem_14__31_0__29_) );
  OR2X2 OR2X2_2676 ( .A(w_mem_inst__abc_21378_n3531_1), .B(w_mem_inst__abc_21378_n3529), .Y(w_mem_inst__abc_21378_n3532) );
  OR2X2 OR2X2_2677 ( .A(w_mem_inst__abc_21378_n3532), .B(w_mem_inst__abc_21378_n3528), .Y(w_mem_inst__0w_mem_14__31_0__30_) );
  OR2X2 OR2X2_2678 ( .A(w_mem_inst__abc_21378_n3537), .B(w_mem_inst__abc_21378_n3535_1), .Y(w_mem_inst__abc_21378_n3538_1) );
  OR2X2 OR2X2_2679 ( .A(w_mem_inst__abc_21378_n3538_1), .B(w_mem_inst__abc_21378_n3534_1), .Y(w_mem_inst__0w_mem_14__31_0__31_) );
  OR2X2 OR2X2_268 ( .A(_abc_15724_n1526), .B(digest_update_bF_buf3), .Y(_abc_15724_n1527) );
  OR2X2 OR2X2_2680 ( .A(w_mem_inst__abc_21378_n3543_1), .B(w_mem_inst__abc_21378_n3541), .Y(w_mem_inst__abc_21378_n3544) );
  OR2X2 OR2X2_2681 ( .A(w_mem_inst__abc_21378_n3544), .B(w_mem_inst__abc_21378_n3540), .Y(w_mem_inst__0w_mem_13__31_0__0_) );
  OR2X2 OR2X2_2682 ( .A(w_mem_inst__abc_21378_n3549), .B(w_mem_inst__abc_21378_n3547_1), .Y(w_mem_inst__abc_21378_n3550_1) );
  OR2X2 OR2X2_2683 ( .A(w_mem_inst__abc_21378_n3550_1), .B(w_mem_inst__abc_21378_n3546_1), .Y(w_mem_inst__0w_mem_13__31_0__1_) );
  OR2X2 OR2X2_2684 ( .A(w_mem_inst__abc_21378_n3555_1), .B(w_mem_inst__abc_21378_n3553), .Y(w_mem_inst__abc_21378_n3556) );
  OR2X2 OR2X2_2685 ( .A(w_mem_inst__abc_21378_n3556), .B(w_mem_inst__abc_21378_n3552), .Y(w_mem_inst__0w_mem_13__31_0__2_) );
  OR2X2 OR2X2_2686 ( .A(w_mem_inst__abc_21378_n3561), .B(w_mem_inst__abc_21378_n3559_1), .Y(w_mem_inst__abc_21378_n3562_1) );
  OR2X2 OR2X2_2687 ( .A(w_mem_inst__abc_21378_n3562_1), .B(w_mem_inst__abc_21378_n3558_1), .Y(w_mem_inst__0w_mem_13__31_0__3_) );
  OR2X2 OR2X2_2688 ( .A(w_mem_inst__abc_21378_n3567_1), .B(w_mem_inst__abc_21378_n3565), .Y(w_mem_inst__abc_21378_n3568) );
  OR2X2 OR2X2_2689 ( .A(w_mem_inst__abc_21378_n3568), .B(w_mem_inst__abc_21378_n3564), .Y(w_mem_inst__0w_mem_13__31_0__4_) );
  OR2X2 OR2X2_269 ( .A(_auto_iopadmap_cc_313_execute_26059_66_), .B(c_reg_2_), .Y(_abc_15724_n1530_1) );
  OR2X2 OR2X2_2690 ( .A(w_mem_inst__abc_21378_n3573), .B(w_mem_inst__abc_21378_n3571_1), .Y(w_mem_inst__abc_21378_n3574_1) );
  OR2X2 OR2X2_2691 ( .A(w_mem_inst__abc_21378_n3574_1), .B(w_mem_inst__abc_21378_n3570_1), .Y(w_mem_inst__0w_mem_13__31_0__5_) );
  OR2X2 OR2X2_2692 ( .A(w_mem_inst__abc_21378_n3579_1), .B(w_mem_inst__abc_21378_n3577), .Y(w_mem_inst__abc_21378_n3580) );
  OR2X2 OR2X2_2693 ( .A(w_mem_inst__abc_21378_n3580), .B(w_mem_inst__abc_21378_n3576), .Y(w_mem_inst__0w_mem_13__31_0__6_) );
  OR2X2 OR2X2_2694 ( .A(w_mem_inst__abc_21378_n3585), .B(w_mem_inst__abc_21378_n3583_1), .Y(w_mem_inst__abc_21378_n3586_1) );
  OR2X2 OR2X2_2695 ( .A(w_mem_inst__abc_21378_n3586_1), .B(w_mem_inst__abc_21378_n3582_1), .Y(w_mem_inst__0w_mem_13__31_0__7_) );
  OR2X2 OR2X2_2696 ( .A(w_mem_inst__abc_21378_n3591_1), .B(w_mem_inst__abc_21378_n3589), .Y(w_mem_inst__abc_21378_n3592) );
  OR2X2 OR2X2_2697 ( .A(w_mem_inst__abc_21378_n3592), .B(w_mem_inst__abc_21378_n3588), .Y(w_mem_inst__0w_mem_13__31_0__8_) );
  OR2X2 OR2X2_2698 ( .A(w_mem_inst__abc_21378_n3597), .B(w_mem_inst__abc_21378_n3595_1), .Y(w_mem_inst__abc_21378_n3598_1) );
  OR2X2 OR2X2_2699 ( .A(w_mem_inst__abc_21378_n3598_1), .B(w_mem_inst__abc_21378_n3594_1), .Y(w_mem_inst__0w_mem_13__31_0__9_) );
  OR2X2 OR2X2_27 ( .A(e_reg_2_), .B(_auto_iopadmap_cc_313_execute_26059_2_), .Y(_abc_15724_n800) );
  OR2X2 OR2X2_270 ( .A(_abc_15724_n1529), .B(_abc_15724_n1534), .Y(_abc_15724_n1535) );
  OR2X2 OR2X2_2700 ( .A(w_mem_inst__abc_21378_n3603_1), .B(w_mem_inst__abc_21378_n3601), .Y(w_mem_inst__abc_21378_n3604) );
  OR2X2 OR2X2_2701 ( .A(w_mem_inst__abc_21378_n3604), .B(w_mem_inst__abc_21378_n3600), .Y(w_mem_inst__0w_mem_13__31_0__10_) );
  OR2X2 OR2X2_2702 ( .A(w_mem_inst__abc_21378_n3609), .B(w_mem_inst__abc_21378_n3607_1), .Y(w_mem_inst__abc_21378_n3610_1) );
  OR2X2 OR2X2_2703 ( .A(w_mem_inst__abc_21378_n3610_1), .B(w_mem_inst__abc_21378_n3606_1), .Y(w_mem_inst__0w_mem_13__31_0__11_) );
  OR2X2 OR2X2_2704 ( .A(w_mem_inst__abc_21378_n3615_1), .B(w_mem_inst__abc_21378_n3613), .Y(w_mem_inst__abc_21378_n3616) );
  OR2X2 OR2X2_2705 ( .A(w_mem_inst__abc_21378_n3616), .B(w_mem_inst__abc_21378_n3612), .Y(w_mem_inst__0w_mem_13__31_0__12_) );
  OR2X2 OR2X2_2706 ( .A(w_mem_inst__abc_21378_n3621), .B(w_mem_inst__abc_21378_n3619_1), .Y(w_mem_inst__abc_21378_n3622_1) );
  OR2X2 OR2X2_2707 ( .A(w_mem_inst__abc_21378_n3622_1), .B(w_mem_inst__abc_21378_n3618_1), .Y(w_mem_inst__0w_mem_13__31_0__13_) );
  OR2X2 OR2X2_2708 ( .A(w_mem_inst__abc_21378_n3627_1), .B(w_mem_inst__abc_21378_n3625), .Y(w_mem_inst__abc_21378_n3628) );
  OR2X2 OR2X2_2709 ( .A(w_mem_inst__abc_21378_n3628), .B(w_mem_inst__abc_21378_n3624), .Y(w_mem_inst__0w_mem_13__31_0__14_) );
  OR2X2 OR2X2_271 ( .A(_abc_15724_n1536), .B(_abc_15724_n1533_1), .Y(_abc_15724_n1537) );
  OR2X2 OR2X2_2710 ( .A(w_mem_inst__abc_21378_n3633), .B(w_mem_inst__abc_21378_n3631_1), .Y(w_mem_inst__abc_21378_n3634_1) );
  OR2X2 OR2X2_2711 ( .A(w_mem_inst__abc_21378_n3634_1), .B(w_mem_inst__abc_21378_n3630_1), .Y(w_mem_inst__0w_mem_13__31_0__15_) );
  OR2X2 OR2X2_2712 ( .A(w_mem_inst__abc_21378_n3639_1), .B(w_mem_inst__abc_21378_n3637), .Y(w_mem_inst__abc_21378_n3640) );
  OR2X2 OR2X2_2713 ( .A(w_mem_inst__abc_21378_n3640), .B(w_mem_inst__abc_21378_n3636), .Y(w_mem_inst__0w_mem_13__31_0__16_) );
  OR2X2 OR2X2_2714 ( .A(w_mem_inst__abc_21378_n3645), .B(w_mem_inst__abc_21378_n3643_1), .Y(w_mem_inst__abc_21378_n3646_1) );
  OR2X2 OR2X2_2715 ( .A(w_mem_inst__abc_21378_n3646_1), .B(w_mem_inst__abc_21378_n3642_1), .Y(w_mem_inst__0w_mem_13__31_0__17_) );
  OR2X2 OR2X2_2716 ( .A(w_mem_inst__abc_21378_n3651), .B(w_mem_inst__abc_21378_n3649), .Y(w_mem_inst__abc_21378_n3652) );
  OR2X2 OR2X2_2717 ( .A(w_mem_inst__abc_21378_n3652), .B(w_mem_inst__abc_21378_n3648), .Y(w_mem_inst__0w_mem_13__31_0__18_) );
  OR2X2 OR2X2_2718 ( .A(w_mem_inst__abc_21378_n3657_1), .B(w_mem_inst__abc_21378_n3655), .Y(w_mem_inst__abc_21378_n3658) );
  OR2X2 OR2X2_2719 ( .A(w_mem_inst__abc_21378_n3658), .B(w_mem_inst__abc_21378_n3654), .Y(w_mem_inst__0w_mem_13__31_0__19_) );
  OR2X2 OR2X2_272 ( .A(_abc_15724_n1538_1), .B(_abc_15724_n850_bF_buf2), .Y(_abc_15724_n1539) );
  OR2X2 OR2X2_2720 ( .A(w_mem_inst__abc_21378_n3663), .B(w_mem_inst__abc_21378_n3661), .Y(w_mem_inst__abc_21378_n3664) );
  OR2X2 OR2X2_2721 ( .A(w_mem_inst__abc_21378_n3664), .B(w_mem_inst__abc_21378_n3660), .Y(w_mem_inst__0w_mem_13__31_0__20_) );
  OR2X2 OR2X2_2722 ( .A(w_mem_inst__abc_21378_n3669_1), .B(w_mem_inst__abc_21378_n3667), .Y(w_mem_inst__abc_21378_n3670) );
  OR2X2 OR2X2_2723 ( .A(w_mem_inst__abc_21378_n3670), .B(w_mem_inst__abc_21378_n3666), .Y(w_mem_inst__0w_mem_13__31_0__21_) );
  OR2X2 OR2X2_2724 ( .A(w_mem_inst__abc_21378_n3675), .B(w_mem_inst__abc_21378_n3673_1), .Y(w_mem_inst__abc_21378_n3676) );
  OR2X2 OR2X2_2725 ( .A(w_mem_inst__abc_21378_n3676), .B(w_mem_inst__abc_21378_n3672), .Y(w_mem_inst__0w_mem_13__31_0__22_) );
  OR2X2 OR2X2_2726 ( .A(w_mem_inst__abc_21378_n3681), .B(w_mem_inst__abc_21378_n3679), .Y(w_mem_inst__abc_21378_n3682) );
  OR2X2 OR2X2_2727 ( .A(w_mem_inst__abc_21378_n3682), .B(w_mem_inst__abc_21378_n3678), .Y(w_mem_inst__0w_mem_13__31_0__23_) );
  OR2X2 OR2X2_2728 ( .A(w_mem_inst__abc_21378_n3687), .B(w_mem_inst__abc_21378_n3685), .Y(w_mem_inst__abc_21378_n3688) );
  OR2X2 OR2X2_2729 ( .A(w_mem_inst__abc_21378_n3688), .B(w_mem_inst__abc_21378_n3684), .Y(w_mem_inst__0w_mem_13__31_0__24_) );
  OR2X2 OR2X2_273 ( .A(_abc_15724_n851_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_66_), .Y(_abc_15724_n1540_1) );
  OR2X2 OR2X2_2730 ( .A(w_mem_inst__abc_21378_n3693), .B(w_mem_inst__abc_21378_n3691), .Y(w_mem_inst__abc_21378_n3694) );
  OR2X2 OR2X2_2731 ( .A(w_mem_inst__abc_21378_n3694), .B(w_mem_inst__abc_21378_n3690), .Y(w_mem_inst__0w_mem_13__31_0__25_) );
  OR2X2 OR2X2_2732 ( .A(w_mem_inst__abc_21378_n3699), .B(w_mem_inst__abc_21378_n3697), .Y(w_mem_inst__abc_21378_n3700) );
  OR2X2 OR2X2_2733 ( .A(w_mem_inst__abc_21378_n3700), .B(w_mem_inst__abc_21378_n3696), .Y(w_mem_inst__0w_mem_13__31_0__26_) );
  OR2X2 OR2X2_2734 ( .A(w_mem_inst__abc_21378_n3705), .B(w_mem_inst__abc_21378_n3703), .Y(w_mem_inst__abc_21378_n3706) );
  OR2X2 OR2X2_2735 ( .A(w_mem_inst__abc_21378_n3706), .B(w_mem_inst__abc_21378_n3702), .Y(w_mem_inst__0w_mem_13__31_0__27_) );
  OR2X2 OR2X2_2736 ( .A(w_mem_inst__abc_21378_n3711), .B(w_mem_inst__abc_21378_n3709), .Y(w_mem_inst__abc_21378_n3712) );
  OR2X2 OR2X2_2737 ( .A(w_mem_inst__abc_21378_n3712), .B(w_mem_inst__abc_21378_n3708), .Y(w_mem_inst__0w_mem_13__31_0__28_) );
  OR2X2 OR2X2_2738 ( .A(w_mem_inst__abc_21378_n3717), .B(w_mem_inst__abc_21378_n3715), .Y(w_mem_inst__abc_21378_n3718) );
  OR2X2 OR2X2_2739 ( .A(w_mem_inst__abc_21378_n3718), .B(w_mem_inst__abc_21378_n3714), .Y(w_mem_inst__0w_mem_13__31_0__29_) );
  OR2X2 OR2X2_274 ( .A(_abc_15724_n1540_1), .B(digest_update_bF_buf2), .Y(_abc_15724_n1541) );
  OR2X2 OR2X2_2740 ( .A(w_mem_inst__abc_21378_n3723), .B(w_mem_inst__abc_21378_n3721), .Y(w_mem_inst__abc_21378_n3724) );
  OR2X2 OR2X2_2741 ( .A(w_mem_inst__abc_21378_n3724), .B(w_mem_inst__abc_21378_n3720), .Y(w_mem_inst__0w_mem_13__31_0__30_) );
  OR2X2 OR2X2_2742 ( .A(w_mem_inst__abc_21378_n3729), .B(w_mem_inst__abc_21378_n3727), .Y(w_mem_inst__abc_21378_n3730) );
  OR2X2 OR2X2_2743 ( .A(w_mem_inst__abc_21378_n3730), .B(w_mem_inst__abc_21378_n3726), .Y(w_mem_inst__0w_mem_13__31_0__31_) );
  OR2X2 OR2X2_2744 ( .A(w_mem_inst__abc_21378_n3735), .B(w_mem_inst__abc_21378_n3733), .Y(w_mem_inst__abc_21378_n3736) );
  OR2X2 OR2X2_2745 ( .A(w_mem_inst__abc_21378_n3736), .B(w_mem_inst__abc_21378_n3732), .Y(w_mem_inst__0w_mem_12__31_0__0_) );
  OR2X2 OR2X2_2746 ( .A(w_mem_inst__abc_21378_n3741), .B(w_mem_inst__abc_21378_n3739), .Y(w_mem_inst__abc_21378_n3742) );
  OR2X2 OR2X2_2747 ( .A(w_mem_inst__abc_21378_n3742), .B(w_mem_inst__abc_21378_n3738), .Y(w_mem_inst__0w_mem_12__31_0__1_) );
  OR2X2 OR2X2_2748 ( .A(w_mem_inst__abc_21378_n3747), .B(w_mem_inst__abc_21378_n3745), .Y(w_mem_inst__abc_21378_n3748) );
  OR2X2 OR2X2_2749 ( .A(w_mem_inst__abc_21378_n3748), .B(w_mem_inst__abc_21378_n3744), .Y(w_mem_inst__0w_mem_12__31_0__2_) );
  OR2X2 OR2X2_275 ( .A(_auto_iopadmap_cc_313_execute_26059_67_), .B(c_reg_3_), .Y(_abc_15724_n1544) );
  OR2X2 OR2X2_2750 ( .A(w_mem_inst__abc_21378_n3753), .B(w_mem_inst__abc_21378_n3751), .Y(w_mem_inst__abc_21378_n3754) );
  OR2X2 OR2X2_2751 ( .A(w_mem_inst__abc_21378_n3754), .B(w_mem_inst__abc_21378_n3750), .Y(w_mem_inst__0w_mem_12__31_0__3_) );
  OR2X2 OR2X2_2752 ( .A(w_mem_inst__abc_21378_n3759), .B(w_mem_inst__abc_21378_n3757), .Y(w_mem_inst__abc_21378_n3760) );
  OR2X2 OR2X2_2753 ( .A(w_mem_inst__abc_21378_n3760), .B(w_mem_inst__abc_21378_n3756), .Y(w_mem_inst__0w_mem_12__31_0__4_) );
  OR2X2 OR2X2_2754 ( .A(w_mem_inst__abc_21378_n3765), .B(w_mem_inst__abc_21378_n3763), .Y(w_mem_inst__abc_21378_n3766) );
  OR2X2 OR2X2_2755 ( .A(w_mem_inst__abc_21378_n3766), .B(w_mem_inst__abc_21378_n3762), .Y(w_mem_inst__0w_mem_12__31_0__5_) );
  OR2X2 OR2X2_2756 ( .A(w_mem_inst__abc_21378_n3771), .B(w_mem_inst__abc_21378_n3769), .Y(w_mem_inst__abc_21378_n3772) );
  OR2X2 OR2X2_2757 ( .A(w_mem_inst__abc_21378_n3772), .B(w_mem_inst__abc_21378_n3768), .Y(w_mem_inst__0w_mem_12__31_0__6_) );
  OR2X2 OR2X2_2758 ( .A(w_mem_inst__abc_21378_n3777), .B(w_mem_inst__abc_21378_n3775), .Y(w_mem_inst__abc_21378_n3778) );
  OR2X2 OR2X2_2759 ( .A(w_mem_inst__abc_21378_n3778), .B(w_mem_inst__abc_21378_n3774), .Y(w_mem_inst__0w_mem_12__31_0__7_) );
  OR2X2 OR2X2_276 ( .A(_abc_15724_n1551), .B(_abc_15724_n1548_1), .Y(_abc_15724_n1552) );
  OR2X2 OR2X2_2760 ( .A(w_mem_inst__abc_21378_n3783), .B(w_mem_inst__abc_21378_n3781), .Y(w_mem_inst__abc_21378_n3784) );
  OR2X2 OR2X2_2761 ( .A(w_mem_inst__abc_21378_n3784), .B(w_mem_inst__abc_21378_n3780), .Y(w_mem_inst__0w_mem_12__31_0__8_) );
  OR2X2 OR2X2_2762 ( .A(w_mem_inst__abc_21378_n3789), .B(w_mem_inst__abc_21378_n3787), .Y(w_mem_inst__abc_21378_n3790) );
  OR2X2 OR2X2_2763 ( .A(w_mem_inst__abc_21378_n3790), .B(w_mem_inst__abc_21378_n3786), .Y(w_mem_inst__0w_mem_12__31_0__9_) );
  OR2X2 OR2X2_2764 ( .A(w_mem_inst__abc_21378_n3795), .B(w_mem_inst__abc_21378_n3793), .Y(w_mem_inst__abc_21378_n3796) );
  OR2X2 OR2X2_2765 ( .A(w_mem_inst__abc_21378_n3796), .B(w_mem_inst__abc_21378_n3792), .Y(w_mem_inst__0w_mem_12__31_0__10_) );
  OR2X2 OR2X2_2766 ( .A(w_mem_inst__abc_21378_n3801), .B(w_mem_inst__abc_21378_n3799), .Y(w_mem_inst__abc_21378_n3802) );
  OR2X2 OR2X2_2767 ( .A(w_mem_inst__abc_21378_n3802), .B(w_mem_inst__abc_21378_n3798), .Y(w_mem_inst__0w_mem_12__31_0__11_) );
  OR2X2 OR2X2_2768 ( .A(w_mem_inst__abc_21378_n3807), .B(w_mem_inst__abc_21378_n3805), .Y(w_mem_inst__abc_21378_n3808) );
  OR2X2 OR2X2_2769 ( .A(w_mem_inst__abc_21378_n3808), .B(w_mem_inst__abc_21378_n3804), .Y(w_mem_inst__0w_mem_12__31_0__12_) );
  OR2X2 OR2X2_277 ( .A(_abc_15724_n851_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_67_), .Y(_abc_15724_n1554) );
  OR2X2 OR2X2_2770 ( .A(w_mem_inst__abc_21378_n3813), .B(w_mem_inst__abc_21378_n3811), .Y(w_mem_inst__abc_21378_n3814) );
  OR2X2 OR2X2_2771 ( .A(w_mem_inst__abc_21378_n3814), .B(w_mem_inst__abc_21378_n3810), .Y(w_mem_inst__0w_mem_12__31_0__13_) );
  OR2X2 OR2X2_2772 ( .A(w_mem_inst__abc_21378_n3819), .B(w_mem_inst__abc_21378_n3817), .Y(w_mem_inst__abc_21378_n3820) );
  OR2X2 OR2X2_2773 ( .A(w_mem_inst__abc_21378_n3820), .B(w_mem_inst__abc_21378_n3816), .Y(w_mem_inst__0w_mem_12__31_0__14_) );
  OR2X2 OR2X2_2774 ( .A(w_mem_inst__abc_21378_n3825), .B(w_mem_inst__abc_21378_n3823), .Y(w_mem_inst__abc_21378_n3826) );
  OR2X2 OR2X2_2775 ( .A(w_mem_inst__abc_21378_n3826), .B(w_mem_inst__abc_21378_n3822), .Y(w_mem_inst__0w_mem_12__31_0__15_) );
  OR2X2 OR2X2_2776 ( .A(w_mem_inst__abc_21378_n3831), .B(w_mem_inst__abc_21378_n3829), .Y(w_mem_inst__abc_21378_n3832) );
  OR2X2 OR2X2_2777 ( .A(w_mem_inst__abc_21378_n3832), .B(w_mem_inst__abc_21378_n3828), .Y(w_mem_inst__0w_mem_12__31_0__16_) );
  OR2X2 OR2X2_2778 ( .A(w_mem_inst__abc_21378_n3837), .B(w_mem_inst__abc_21378_n3835), .Y(w_mem_inst__abc_21378_n3838) );
  OR2X2 OR2X2_2779 ( .A(w_mem_inst__abc_21378_n3838), .B(w_mem_inst__abc_21378_n3834), .Y(w_mem_inst__0w_mem_12__31_0__17_) );
  OR2X2 OR2X2_278 ( .A(_abc_15724_n1553), .B(_abc_15724_n1555), .Y(H2_reg_3__FF_INPUT) );
  OR2X2 OR2X2_2780 ( .A(w_mem_inst__abc_21378_n3843), .B(w_mem_inst__abc_21378_n3841), .Y(w_mem_inst__abc_21378_n3844) );
  OR2X2 OR2X2_2781 ( .A(w_mem_inst__abc_21378_n3844), .B(w_mem_inst__abc_21378_n3840), .Y(w_mem_inst__0w_mem_12__31_0__18_) );
  OR2X2 OR2X2_2782 ( .A(w_mem_inst__abc_21378_n3849), .B(w_mem_inst__abc_21378_n3847), .Y(w_mem_inst__abc_21378_n3850) );
  OR2X2 OR2X2_2783 ( .A(w_mem_inst__abc_21378_n3850), .B(w_mem_inst__abc_21378_n3846), .Y(w_mem_inst__0w_mem_12__31_0__19_) );
  OR2X2 OR2X2_2784 ( .A(w_mem_inst__abc_21378_n3855), .B(w_mem_inst__abc_21378_n3853), .Y(w_mem_inst__abc_21378_n3856) );
  OR2X2 OR2X2_2785 ( .A(w_mem_inst__abc_21378_n3856), .B(w_mem_inst__abc_21378_n3852), .Y(w_mem_inst__0w_mem_12__31_0__20_) );
  OR2X2 OR2X2_2786 ( .A(w_mem_inst__abc_21378_n3861), .B(w_mem_inst__abc_21378_n3859), .Y(w_mem_inst__abc_21378_n3862) );
  OR2X2 OR2X2_2787 ( .A(w_mem_inst__abc_21378_n3862), .B(w_mem_inst__abc_21378_n3858), .Y(w_mem_inst__0w_mem_12__31_0__21_) );
  OR2X2 OR2X2_2788 ( .A(w_mem_inst__abc_21378_n3867), .B(w_mem_inst__abc_21378_n3865), .Y(w_mem_inst__abc_21378_n3868) );
  OR2X2 OR2X2_2789 ( .A(w_mem_inst__abc_21378_n3868), .B(w_mem_inst__abc_21378_n3864), .Y(w_mem_inst__0w_mem_12__31_0__22_) );
  OR2X2 OR2X2_279 ( .A(_auto_iopadmap_cc_313_execute_26059_68_), .B(c_reg_4_), .Y(_abc_15724_n1557_1) );
  OR2X2 OR2X2_2790 ( .A(w_mem_inst__abc_21378_n3873), .B(w_mem_inst__abc_21378_n3871), .Y(w_mem_inst__abc_21378_n3874) );
  OR2X2 OR2X2_2791 ( .A(w_mem_inst__abc_21378_n3874), .B(w_mem_inst__abc_21378_n3870), .Y(w_mem_inst__0w_mem_12__31_0__23_) );
  OR2X2 OR2X2_2792 ( .A(w_mem_inst__abc_21378_n3879), .B(w_mem_inst__abc_21378_n3877), .Y(w_mem_inst__abc_21378_n3880) );
  OR2X2 OR2X2_2793 ( .A(w_mem_inst__abc_21378_n3880), .B(w_mem_inst__abc_21378_n3876), .Y(w_mem_inst__0w_mem_12__31_0__24_) );
  OR2X2 OR2X2_2794 ( .A(w_mem_inst__abc_21378_n3885), .B(w_mem_inst__abc_21378_n3883), .Y(w_mem_inst__abc_21378_n3886) );
  OR2X2 OR2X2_2795 ( .A(w_mem_inst__abc_21378_n3886), .B(w_mem_inst__abc_21378_n3882), .Y(w_mem_inst__0w_mem_12__31_0__25_) );
  OR2X2 OR2X2_2796 ( .A(w_mem_inst__abc_21378_n3891), .B(w_mem_inst__abc_21378_n3889), .Y(w_mem_inst__abc_21378_n3892) );
  OR2X2 OR2X2_2797 ( .A(w_mem_inst__abc_21378_n3892), .B(w_mem_inst__abc_21378_n3888), .Y(w_mem_inst__0w_mem_12__31_0__26_) );
  OR2X2 OR2X2_2798 ( .A(w_mem_inst__abc_21378_n3897), .B(w_mem_inst__abc_21378_n3895), .Y(w_mem_inst__abc_21378_n3898) );
  OR2X2 OR2X2_2799 ( .A(w_mem_inst__abc_21378_n3898), .B(w_mem_inst__abc_21378_n3894), .Y(w_mem_inst__0w_mem_12__31_0__27_) );
  OR2X2 OR2X2_28 ( .A(_abc_15724_n802), .B(_abc_15724_n789_1), .Y(_abc_15724_n803_1) );
  OR2X2 OR2X2_280 ( .A(_abc_15724_n1543_1), .B(_abc_15724_n1562), .Y(_abc_15724_n1563_1) );
  OR2X2 OR2X2_2800 ( .A(w_mem_inst__abc_21378_n3903), .B(w_mem_inst__abc_21378_n3901), .Y(w_mem_inst__abc_21378_n3904) );
  OR2X2 OR2X2_2801 ( .A(w_mem_inst__abc_21378_n3904), .B(w_mem_inst__abc_21378_n3900), .Y(w_mem_inst__0w_mem_12__31_0__28_) );
  OR2X2 OR2X2_2802 ( .A(w_mem_inst__abc_21378_n3909), .B(w_mem_inst__abc_21378_n3907), .Y(w_mem_inst__abc_21378_n3910) );
  OR2X2 OR2X2_2803 ( .A(w_mem_inst__abc_21378_n3910), .B(w_mem_inst__abc_21378_n3906), .Y(w_mem_inst__0w_mem_12__31_0__29_) );
  OR2X2 OR2X2_2804 ( .A(w_mem_inst__abc_21378_n3915), .B(w_mem_inst__abc_21378_n3913), .Y(w_mem_inst__abc_21378_n3916) );
  OR2X2 OR2X2_2805 ( .A(w_mem_inst__abc_21378_n3916), .B(w_mem_inst__abc_21378_n3912), .Y(w_mem_inst__0w_mem_12__31_0__30_) );
  OR2X2 OR2X2_2806 ( .A(w_mem_inst__abc_21378_n3921), .B(w_mem_inst__abc_21378_n3919), .Y(w_mem_inst__abc_21378_n3922) );
  OR2X2 OR2X2_2807 ( .A(w_mem_inst__abc_21378_n3922), .B(w_mem_inst__abc_21378_n3918), .Y(w_mem_inst__0w_mem_12__31_0__31_) );
  OR2X2 OR2X2_2808 ( .A(w_mem_inst__abc_21378_n3927), .B(w_mem_inst__abc_21378_n3925), .Y(w_mem_inst__abc_21378_n3928) );
  OR2X2 OR2X2_2809 ( .A(w_mem_inst__abc_21378_n3928), .B(w_mem_inst__abc_21378_n3924), .Y(w_mem_inst__0w_mem_11__31_0__0_) );
  OR2X2 OR2X2_281 ( .A(_abc_15724_n1564_1), .B(_abc_15724_n1561), .Y(_abc_15724_n1565) );
  OR2X2 OR2X2_2810 ( .A(w_mem_inst__abc_21378_n3933), .B(w_mem_inst__abc_21378_n3931), .Y(w_mem_inst__abc_21378_n3934) );
  OR2X2 OR2X2_2811 ( .A(w_mem_inst__abc_21378_n3934), .B(w_mem_inst__abc_21378_n3930), .Y(w_mem_inst__0w_mem_11__31_0__1_) );
  OR2X2 OR2X2_2812 ( .A(w_mem_inst__abc_21378_n3939), .B(w_mem_inst__abc_21378_n3937), .Y(w_mem_inst__abc_21378_n3940) );
  OR2X2 OR2X2_2813 ( .A(w_mem_inst__abc_21378_n3940), .B(w_mem_inst__abc_21378_n3936), .Y(w_mem_inst__0w_mem_11__31_0__2_) );
  OR2X2 OR2X2_2814 ( .A(w_mem_inst__abc_21378_n3945), .B(w_mem_inst__abc_21378_n3943), .Y(w_mem_inst__abc_21378_n3946) );
  OR2X2 OR2X2_2815 ( .A(w_mem_inst__abc_21378_n3946), .B(w_mem_inst__abc_21378_n3942), .Y(w_mem_inst__0w_mem_11__31_0__3_) );
  OR2X2 OR2X2_2816 ( .A(w_mem_inst__abc_21378_n3951), .B(w_mem_inst__abc_21378_n3949), .Y(w_mem_inst__abc_21378_n3952) );
  OR2X2 OR2X2_2817 ( .A(w_mem_inst__abc_21378_n3952), .B(w_mem_inst__abc_21378_n3948), .Y(w_mem_inst__0w_mem_11__31_0__4_) );
  OR2X2 OR2X2_2818 ( .A(w_mem_inst__abc_21378_n3957), .B(w_mem_inst__abc_21378_n3955), .Y(w_mem_inst__abc_21378_n3958) );
  OR2X2 OR2X2_2819 ( .A(w_mem_inst__abc_21378_n3958), .B(w_mem_inst__abc_21378_n3954), .Y(w_mem_inst__0w_mem_11__31_0__5_) );
  OR2X2 OR2X2_282 ( .A(_abc_15724_n1566), .B(_abc_15724_n1560), .Y(_abc_15724_n1567) );
  OR2X2 OR2X2_2820 ( .A(w_mem_inst__abc_21378_n3963), .B(w_mem_inst__abc_21378_n3961), .Y(w_mem_inst__abc_21378_n3964) );
  OR2X2 OR2X2_2821 ( .A(w_mem_inst__abc_21378_n3964), .B(w_mem_inst__abc_21378_n3960), .Y(w_mem_inst__0w_mem_11__31_0__6_) );
  OR2X2 OR2X2_2822 ( .A(w_mem_inst__abc_21378_n3969), .B(w_mem_inst__abc_21378_n3967), .Y(w_mem_inst__abc_21378_n3970) );
  OR2X2 OR2X2_2823 ( .A(w_mem_inst__abc_21378_n3970), .B(w_mem_inst__abc_21378_n3966), .Y(w_mem_inst__0w_mem_11__31_0__7_) );
  OR2X2 OR2X2_2824 ( .A(w_mem_inst__abc_21378_n3975), .B(w_mem_inst__abc_21378_n3973), .Y(w_mem_inst__abc_21378_n3976) );
  OR2X2 OR2X2_2825 ( .A(w_mem_inst__abc_21378_n3976), .B(w_mem_inst__abc_21378_n3972), .Y(w_mem_inst__0w_mem_11__31_0__8_) );
  OR2X2 OR2X2_2826 ( .A(w_mem_inst__abc_21378_n3981), .B(w_mem_inst__abc_21378_n3979), .Y(w_mem_inst__abc_21378_n3982) );
  OR2X2 OR2X2_2827 ( .A(w_mem_inst__abc_21378_n3982), .B(w_mem_inst__abc_21378_n3978), .Y(w_mem_inst__0w_mem_11__31_0__9_) );
  OR2X2 OR2X2_2828 ( .A(w_mem_inst__abc_21378_n3987), .B(w_mem_inst__abc_21378_n3985), .Y(w_mem_inst__abc_21378_n3988) );
  OR2X2 OR2X2_2829 ( .A(w_mem_inst__abc_21378_n3988), .B(w_mem_inst__abc_21378_n3984), .Y(w_mem_inst__0w_mem_11__31_0__10_) );
  OR2X2 OR2X2_283 ( .A(_abc_15724_n1568), .B(_abc_15724_n850_bF_buf0), .Y(_abc_15724_n1569) );
  OR2X2 OR2X2_2830 ( .A(w_mem_inst__abc_21378_n3993), .B(w_mem_inst__abc_21378_n3991), .Y(w_mem_inst__abc_21378_n3994) );
  OR2X2 OR2X2_2831 ( .A(w_mem_inst__abc_21378_n3994), .B(w_mem_inst__abc_21378_n3990), .Y(w_mem_inst__0w_mem_11__31_0__11_) );
  OR2X2 OR2X2_2832 ( .A(w_mem_inst__abc_21378_n3999), .B(w_mem_inst__abc_21378_n3997), .Y(w_mem_inst__abc_21378_n4000) );
  OR2X2 OR2X2_2833 ( .A(w_mem_inst__abc_21378_n4000), .B(w_mem_inst__abc_21378_n3996), .Y(w_mem_inst__0w_mem_11__31_0__12_) );
  OR2X2 OR2X2_2834 ( .A(w_mem_inst__abc_21378_n4005), .B(w_mem_inst__abc_21378_n4003), .Y(w_mem_inst__abc_21378_n4006) );
  OR2X2 OR2X2_2835 ( .A(w_mem_inst__abc_21378_n4006), .B(w_mem_inst__abc_21378_n4002), .Y(w_mem_inst__0w_mem_11__31_0__13_) );
  OR2X2 OR2X2_2836 ( .A(w_mem_inst__abc_21378_n4011), .B(w_mem_inst__abc_21378_n4009), .Y(w_mem_inst__abc_21378_n4012) );
  OR2X2 OR2X2_2837 ( .A(w_mem_inst__abc_21378_n4012), .B(w_mem_inst__abc_21378_n4008), .Y(w_mem_inst__0w_mem_11__31_0__14_) );
  OR2X2 OR2X2_2838 ( .A(w_mem_inst__abc_21378_n4017), .B(w_mem_inst__abc_21378_n4015), .Y(w_mem_inst__abc_21378_n4018) );
  OR2X2 OR2X2_2839 ( .A(w_mem_inst__abc_21378_n4018), .B(w_mem_inst__abc_21378_n4014), .Y(w_mem_inst__0w_mem_11__31_0__15_) );
  OR2X2 OR2X2_284 ( .A(_abc_15724_n851_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_68_), .Y(_abc_15724_n1570_1) );
  OR2X2 OR2X2_2840 ( .A(w_mem_inst__abc_21378_n4023), .B(w_mem_inst__abc_21378_n4021), .Y(w_mem_inst__abc_21378_n4024) );
  OR2X2 OR2X2_2841 ( .A(w_mem_inst__abc_21378_n4024), .B(w_mem_inst__abc_21378_n4020), .Y(w_mem_inst__0w_mem_11__31_0__16_) );
  OR2X2 OR2X2_2842 ( .A(w_mem_inst__abc_21378_n4029), .B(w_mem_inst__abc_21378_n4027), .Y(w_mem_inst__abc_21378_n4030) );
  OR2X2 OR2X2_2843 ( .A(w_mem_inst__abc_21378_n4030), .B(w_mem_inst__abc_21378_n4026), .Y(w_mem_inst__0w_mem_11__31_0__17_) );
  OR2X2 OR2X2_2844 ( .A(w_mem_inst__abc_21378_n4035), .B(w_mem_inst__abc_21378_n4033), .Y(w_mem_inst__abc_21378_n4036) );
  OR2X2 OR2X2_2845 ( .A(w_mem_inst__abc_21378_n4036), .B(w_mem_inst__abc_21378_n4032), .Y(w_mem_inst__0w_mem_11__31_0__18_) );
  OR2X2 OR2X2_2846 ( .A(w_mem_inst__abc_21378_n4041), .B(w_mem_inst__abc_21378_n4039), .Y(w_mem_inst__abc_21378_n4042) );
  OR2X2 OR2X2_2847 ( .A(w_mem_inst__abc_21378_n4042), .B(w_mem_inst__abc_21378_n4038), .Y(w_mem_inst__0w_mem_11__31_0__19_) );
  OR2X2 OR2X2_2848 ( .A(w_mem_inst__abc_21378_n4047), .B(w_mem_inst__abc_21378_n4045), .Y(w_mem_inst__abc_21378_n4048) );
  OR2X2 OR2X2_2849 ( .A(w_mem_inst__abc_21378_n4048), .B(w_mem_inst__abc_21378_n4044), .Y(w_mem_inst__0w_mem_11__31_0__20_) );
  OR2X2 OR2X2_285 ( .A(_abc_15724_n1570_1), .B(digest_update_bF_buf0), .Y(_abc_15724_n1571_1) );
  OR2X2 OR2X2_2850 ( .A(w_mem_inst__abc_21378_n4053), .B(w_mem_inst__abc_21378_n4051), .Y(w_mem_inst__abc_21378_n4054) );
  OR2X2 OR2X2_2851 ( .A(w_mem_inst__abc_21378_n4054), .B(w_mem_inst__abc_21378_n4050), .Y(w_mem_inst__0w_mem_11__31_0__21_) );
  OR2X2 OR2X2_2852 ( .A(w_mem_inst__abc_21378_n4059), .B(w_mem_inst__abc_21378_n4057), .Y(w_mem_inst__abc_21378_n4060) );
  OR2X2 OR2X2_2853 ( .A(w_mem_inst__abc_21378_n4060), .B(w_mem_inst__abc_21378_n4056), .Y(w_mem_inst__0w_mem_11__31_0__22_) );
  OR2X2 OR2X2_2854 ( .A(w_mem_inst__abc_21378_n4065), .B(w_mem_inst__abc_21378_n4063), .Y(w_mem_inst__abc_21378_n4066) );
  OR2X2 OR2X2_2855 ( .A(w_mem_inst__abc_21378_n4066), .B(w_mem_inst__abc_21378_n4062), .Y(w_mem_inst__0w_mem_11__31_0__23_) );
  OR2X2 OR2X2_2856 ( .A(w_mem_inst__abc_21378_n4071), .B(w_mem_inst__abc_21378_n4069), .Y(w_mem_inst__abc_21378_n4072) );
  OR2X2 OR2X2_2857 ( .A(w_mem_inst__abc_21378_n4072), .B(w_mem_inst__abc_21378_n4068), .Y(w_mem_inst__0w_mem_11__31_0__24_) );
  OR2X2 OR2X2_2858 ( .A(w_mem_inst__abc_21378_n4077), .B(w_mem_inst__abc_21378_n4075), .Y(w_mem_inst__abc_21378_n4078) );
  OR2X2 OR2X2_2859 ( .A(w_mem_inst__abc_21378_n4078), .B(w_mem_inst__abc_21378_n4074), .Y(w_mem_inst__0w_mem_11__31_0__25_) );
  OR2X2 OR2X2_286 ( .A(_auto_iopadmap_cc_313_execute_26059_69_), .B(c_reg_5_), .Y(_abc_15724_n1575) );
  OR2X2 OR2X2_2860 ( .A(w_mem_inst__abc_21378_n4083), .B(w_mem_inst__abc_21378_n4081), .Y(w_mem_inst__abc_21378_n4084) );
  OR2X2 OR2X2_2861 ( .A(w_mem_inst__abc_21378_n4084), .B(w_mem_inst__abc_21378_n4080), .Y(w_mem_inst__0w_mem_11__31_0__26_) );
  OR2X2 OR2X2_2862 ( .A(w_mem_inst__abc_21378_n4089), .B(w_mem_inst__abc_21378_n4087), .Y(w_mem_inst__abc_21378_n4090) );
  OR2X2 OR2X2_2863 ( .A(w_mem_inst__abc_21378_n4090), .B(w_mem_inst__abc_21378_n4086), .Y(w_mem_inst__0w_mem_11__31_0__27_) );
  OR2X2 OR2X2_2864 ( .A(w_mem_inst__abc_21378_n4095), .B(w_mem_inst__abc_21378_n4093), .Y(w_mem_inst__abc_21378_n4096) );
  OR2X2 OR2X2_2865 ( .A(w_mem_inst__abc_21378_n4096), .B(w_mem_inst__abc_21378_n4092), .Y(w_mem_inst__0w_mem_11__31_0__28_) );
  OR2X2 OR2X2_2866 ( .A(w_mem_inst__abc_21378_n4101), .B(w_mem_inst__abc_21378_n4099), .Y(w_mem_inst__abc_21378_n4102) );
  OR2X2 OR2X2_2867 ( .A(w_mem_inst__abc_21378_n4102), .B(w_mem_inst__abc_21378_n4098), .Y(w_mem_inst__0w_mem_11__31_0__29_) );
  OR2X2 OR2X2_2868 ( .A(w_mem_inst__abc_21378_n4107), .B(w_mem_inst__abc_21378_n4105), .Y(w_mem_inst__abc_21378_n4108) );
  OR2X2 OR2X2_2869 ( .A(w_mem_inst__abc_21378_n4108), .B(w_mem_inst__abc_21378_n4104), .Y(w_mem_inst__0w_mem_11__31_0__30_) );
  OR2X2 OR2X2_287 ( .A(_abc_15724_n1574), .B(_abc_15724_n1578_1), .Y(_abc_15724_n1579_1) );
  OR2X2 OR2X2_2870 ( .A(w_mem_inst__abc_21378_n4113), .B(w_mem_inst__abc_21378_n4111), .Y(w_mem_inst__abc_21378_n4114) );
  OR2X2 OR2X2_2871 ( .A(w_mem_inst__abc_21378_n4114), .B(w_mem_inst__abc_21378_n4110), .Y(w_mem_inst__0w_mem_11__31_0__31_) );
  OR2X2 OR2X2_2872 ( .A(w_mem_inst__abc_21378_n4119), .B(w_mem_inst__abc_21378_n4117), .Y(w_mem_inst__abc_21378_n4120) );
  OR2X2 OR2X2_2873 ( .A(w_mem_inst__abc_21378_n4120), .B(w_mem_inst__abc_21378_n4116), .Y(w_mem_inst__0w_mem_10__31_0__0_) );
  OR2X2 OR2X2_2874 ( .A(w_mem_inst__abc_21378_n4125), .B(w_mem_inst__abc_21378_n4123), .Y(w_mem_inst__abc_21378_n4126) );
  OR2X2 OR2X2_2875 ( .A(w_mem_inst__abc_21378_n4126), .B(w_mem_inst__abc_21378_n4122), .Y(w_mem_inst__0w_mem_10__31_0__1_) );
  OR2X2 OR2X2_2876 ( .A(w_mem_inst__abc_21378_n4131), .B(w_mem_inst__abc_21378_n4129), .Y(w_mem_inst__abc_21378_n4132) );
  OR2X2 OR2X2_2877 ( .A(w_mem_inst__abc_21378_n4132), .B(w_mem_inst__abc_21378_n4128), .Y(w_mem_inst__0w_mem_10__31_0__2_) );
  OR2X2 OR2X2_2878 ( .A(w_mem_inst__abc_21378_n4137), .B(w_mem_inst__abc_21378_n4135), .Y(w_mem_inst__abc_21378_n4138) );
  OR2X2 OR2X2_2879 ( .A(w_mem_inst__abc_21378_n4138), .B(w_mem_inst__abc_21378_n4134), .Y(w_mem_inst__0w_mem_10__31_0__3_) );
  OR2X2 OR2X2_288 ( .A(_abc_15724_n1573_1), .B(_abc_15724_n1580), .Y(_abc_15724_n1581_1) );
  OR2X2 OR2X2_2880 ( .A(w_mem_inst__abc_21378_n4143), .B(w_mem_inst__abc_21378_n4141), .Y(w_mem_inst__abc_21378_n4144) );
  OR2X2 OR2X2_2881 ( .A(w_mem_inst__abc_21378_n4144), .B(w_mem_inst__abc_21378_n4140), .Y(w_mem_inst__0w_mem_10__31_0__4_) );
  OR2X2 OR2X2_2882 ( .A(w_mem_inst__abc_21378_n4149), .B(w_mem_inst__abc_21378_n4147), .Y(w_mem_inst__abc_21378_n4150) );
  OR2X2 OR2X2_2883 ( .A(w_mem_inst__abc_21378_n4150), .B(w_mem_inst__abc_21378_n4146), .Y(w_mem_inst__0w_mem_10__31_0__5_) );
  OR2X2 OR2X2_2884 ( .A(w_mem_inst__abc_21378_n4155), .B(w_mem_inst__abc_21378_n4153), .Y(w_mem_inst__abc_21378_n4156) );
  OR2X2 OR2X2_2885 ( .A(w_mem_inst__abc_21378_n4156), .B(w_mem_inst__abc_21378_n4152), .Y(w_mem_inst__0w_mem_10__31_0__6_) );
  OR2X2 OR2X2_2886 ( .A(w_mem_inst__abc_21378_n4161), .B(w_mem_inst__abc_21378_n4159), .Y(w_mem_inst__abc_21378_n4162) );
  OR2X2 OR2X2_2887 ( .A(w_mem_inst__abc_21378_n4162), .B(w_mem_inst__abc_21378_n4158), .Y(w_mem_inst__0w_mem_10__31_0__7_) );
  OR2X2 OR2X2_2888 ( .A(w_mem_inst__abc_21378_n4167), .B(w_mem_inst__abc_21378_n4165), .Y(w_mem_inst__abc_21378_n4168) );
  OR2X2 OR2X2_2889 ( .A(w_mem_inst__abc_21378_n4168), .B(w_mem_inst__abc_21378_n4164), .Y(w_mem_inst__0w_mem_10__31_0__8_) );
  OR2X2 OR2X2_289 ( .A(_abc_15724_n851_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_69_), .Y(_abc_15724_n1584_1) );
  OR2X2 OR2X2_2890 ( .A(w_mem_inst__abc_21378_n4173), .B(w_mem_inst__abc_21378_n4171), .Y(w_mem_inst__abc_21378_n4174) );
  OR2X2 OR2X2_2891 ( .A(w_mem_inst__abc_21378_n4174), .B(w_mem_inst__abc_21378_n4170), .Y(w_mem_inst__0w_mem_10__31_0__9_) );
  OR2X2 OR2X2_2892 ( .A(w_mem_inst__abc_21378_n4179), .B(w_mem_inst__abc_21378_n4177), .Y(w_mem_inst__abc_21378_n4180) );
  OR2X2 OR2X2_2893 ( .A(w_mem_inst__abc_21378_n4180), .B(w_mem_inst__abc_21378_n4176), .Y(w_mem_inst__0w_mem_10__31_0__10_) );
  OR2X2 OR2X2_2894 ( .A(w_mem_inst__abc_21378_n4185), .B(w_mem_inst__abc_21378_n4183), .Y(w_mem_inst__abc_21378_n4186) );
  OR2X2 OR2X2_2895 ( .A(w_mem_inst__abc_21378_n4186), .B(w_mem_inst__abc_21378_n4182), .Y(w_mem_inst__0w_mem_10__31_0__11_) );
  OR2X2 OR2X2_2896 ( .A(w_mem_inst__abc_21378_n4191), .B(w_mem_inst__abc_21378_n4189), .Y(w_mem_inst__abc_21378_n4192) );
  OR2X2 OR2X2_2897 ( .A(w_mem_inst__abc_21378_n4192), .B(w_mem_inst__abc_21378_n4188), .Y(w_mem_inst__0w_mem_10__31_0__12_) );
  OR2X2 OR2X2_2898 ( .A(w_mem_inst__abc_21378_n4197), .B(w_mem_inst__abc_21378_n4195), .Y(w_mem_inst__abc_21378_n4198) );
  OR2X2 OR2X2_2899 ( .A(w_mem_inst__abc_21378_n4198), .B(w_mem_inst__abc_21378_n4194), .Y(w_mem_inst__0w_mem_10__31_0__13_) );
  OR2X2 OR2X2_29 ( .A(_abc_15724_n804_1), .B(_abc_15724_n787), .Y(_abc_15724_n805) );
  OR2X2 OR2X2_290 ( .A(_abc_15724_n1583), .B(_abc_15724_n1585_1), .Y(H2_reg_5__FF_INPUT) );
  OR2X2 OR2X2_2900 ( .A(w_mem_inst__abc_21378_n4203), .B(w_mem_inst__abc_21378_n4201), .Y(w_mem_inst__abc_21378_n4204) );
  OR2X2 OR2X2_2901 ( .A(w_mem_inst__abc_21378_n4204), .B(w_mem_inst__abc_21378_n4200), .Y(w_mem_inst__0w_mem_10__31_0__14_) );
  OR2X2 OR2X2_2902 ( .A(w_mem_inst__abc_21378_n4209), .B(w_mem_inst__abc_21378_n4207), .Y(w_mem_inst__abc_21378_n4210) );
  OR2X2 OR2X2_2903 ( .A(w_mem_inst__abc_21378_n4210), .B(w_mem_inst__abc_21378_n4206), .Y(w_mem_inst__0w_mem_10__31_0__15_) );
  OR2X2 OR2X2_2904 ( .A(w_mem_inst__abc_21378_n4215), .B(w_mem_inst__abc_21378_n4213), .Y(w_mem_inst__abc_21378_n4216) );
  OR2X2 OR2X2_2905 ( .A(w_mem_inst__abc_21378_n4216), .B(w_mem_inst__abc_21378_n4212), .Y(w_mem_inst__0w_mem_10__31_0__16_) );
  OR2X2 OR2X2_2906 ( .A(w_mem_inst__abc_21378_n4221), .B(w_mem_inst__abc_21378_n4219), .Y(w_mem_inst__abc_21378_n4222) );
  OR2X2 OR2X2_2907 ( .A(w_mem_inst__abc_21378_n4222), .B(w_mem_inst__abc_21378_n4218), .Y(w_mem_inst__0w_mem_10__31_0__17_) );
  OR2X2 OR2X2_2908 ( .A(w_mem_inst__abc_21378_n4227), .B(w_mem_inst__abc_21378_n4225), .Y(w_mem_inst__abc_21378_n4228) );
  OR2X2 OR2X2_2909 ( .A(w_mem_inst__abc_21378_n4228), .B(w_mem_inst__abc_21378_n4224), .Y(w_mem_inst__0w_mem_10__31_0__18_) );
  OR2X2 OR2X2_291 ( .A(_auto_iopadmap_cc_313_execute_26059_70_), .B(c_reg_6_), .Y(_abc_15724_n1589) );
  OR2X2 OR2X2_2910 ( .A(w_mem_inst__abc_21378_n4233), .B(w_mem_inst__abc_21378_n4231), .Y(w_mem_inst__abc_21378_n4234) );
  OR2X2 OR2X2_2911 ( .A(w_mem_inst__abc_21378_n4234), .B(w_mem_inst__abc_21378_n4230), .Y(w_mem_inst__0w_mem_10__31_0__19_) );
  OR2X2 OR2X2_2912 ( .A(w_mem_inst__abc_21378_n4239), .B(w_mem_inst__abc_21378_n4237), .Y(w_mem_inst__abc_21378_n4240) );
  OR2X2 OR2X2_2913 ( .A(w_mem_inst__abc_21378_n4240), .B(w_mem_inst__abc_21378_n4236), .Y(w_mem_inst__0w_mem_10__31_0__20_) );
  OR2X2 OR2X2_2914 ( .A(w_mem_inst__abc_21378_n4245), .B(w_mem_inst__abc_21378_n4243), .Y(w_mem_inst__abc_21378_n4246) );
  OR2X2 OR2X2_2915 ( .A(w_mem_inst__abc_21378_n4246), .B(w_mem_inst__abc_21378_n4242), .Y(w_mem_inst__0w_mem_10__31_0__21_) );
  OR2X2 OR2X2_2916 ( .A(w_mem_inst__abc_21378_n4251), .B(w_mem_inst__abc_21378_n4249), .Y(w_mem_inst__abc_21378_n4252) );
  OR2X2 OR2X2_2917 ( .A(w_mem_inst__abc_21378_n4252), .B(w_mem_inst__abc_21378_n4248), .Y(w_mem_inst__0w_mem_10__31_0__22_) );
  OR2X2 OR2X2_2918 ( .A(w_mem_inst__abc_21378_n4257), .B(w_mem_inst__abc_21378_n4255), .Y(w_mem_inst__abc_21378_n4258) );
  OR2X2 OR2X2_2919 ( .A(w_mem_inst__abc_21378_n4258), .B(w_mem_inst__abc_21378_n4254), .Y(w_mem_inst__0w_mem_10__31_0__23_) );
  OR2X2 OR2X2_292 ( .A(_abc_15724_n1588), .B(_abc_15724_n1592), .Y(_abc_15724_n1593_1) );
  OR2X2 OR2X2_2920 ( .A(w_mem_inst__abc_21378_n4263), .B(w_mem_inst__abc_21378_n4261), .Y(w_mem_inst__abc_21378_n4264) );
  OR2X2 OR2X2_2921 ( .A(w_mem_inst__abc_21378_n4264), .B(w_mem_inst__abc_21378_n4260), .Y(w_mem_inst__0w_mem_10__31_0__24_) );
  OR2X2 OR2X2_2922 ( .A(w_mem_inst__abc_21378_n4269), .B(w_mem_inst__abc_21378_n4267), .Y(w_mem_inst__abc_21378_n4270) );
  OR2X2 OR2X2_2923 ( .A(w_mem_inst__abc_21378_n4270), .B(w_mem_inst__abc_21378_n4266), .Y(w_mem_inst__0w_mem_10__31_0__25_) );
  OR2X2 OR2X2_2924 ( .A(w_mem_inst__abc_21378_n4275), .B(w_mem_inst__abc_21378_n4273), .Y(w_mem_inst__abc_21378_n4276) );
  OR2X2 OR2X2_2925 ( .A(w_mem_inst__abc_21378_n4276), .B(w_mem_inst__abc_21378_n4272), .Y(w_mem_inst__0w_mem_10__31_0__26_) );
  OR2X2 OR2X2_2926 ( .A(w_mem_inst__abc_21378_n4281), .B(w_mem_inst__abc_21378_n4279), .Y(w_mem_inst__abc_21378_n4282) );
  OR2X2 OR2X2_2927 ( .A(w_mem_inst__abc_21378_n4282), .B(w_mem_inst__abc_21378_n4278), .Y(w_mem_inst__0w_mem_10__31_0__27_) );
  OR2X2 OR2X2_2928 ( .A(w_mem_inst__abc_21378_n4287), .B(w_mem_inst__abc_21378_n4285), .Y(w_mem_inst__abc_21378_n4288) );
  OR2X2 OR2X2_2929 ( .A(w_mem_inst__abc_21378_n4288), .B(w_mem_inst__abc_21378_n4284), .Y(w_mem_inst__0w_mem_10__31_0__28_) );
  OR2X2 OR2X2_293 ( .A(_abc_15724_n1587_1), .B(_abc_15724_n1594), .Y(_abc_15724_n1595) );
  OR2X2 OR2X2_2930 ( .A(w_mem_inst__abc_21378_n4293), .B(w_mem_inst__abc_21378_n4291), .Y(w_mem_inst__abc_21378_n4294) );
  OR2X2 OR2X2_2931 ( .A(w_mem_inst__abc_21378_n4294), .B(w_mem_inst__abc_21378_n4290), .Y(w_mem_inst__0w_mem_10__31_0__29_) );
  OR2X2 OR2X2_2932 ( .A(w_mem_inst__abc_21378_n4299), .B(w_mem_inst__abc_21378_n4297), .Y(w_mem_inst__abc_21378_n4300) );
  OR2X2 OR2X2_2933 ( .A(w_mem_inst__abc_21378_n4300), .B(w_mem_inst__abc_21378_n4296), .Y(w_mem_inst__0w_mem_10__31_0__30_) );
  OR2X2 OR2X2_2934 ( .A(w_mem_inst__abc_21378_n4305), .B(w_mem_inst__abc_21378_n4303), .Y(w_mem_inst__abc_21378_n4306) );
  OR2X2 OR2X2_2935 ( .A(w_mem_inst__abc_21378_n4306), .B(w_mem_inst__abc_21378_n4302), .Y(w_mem_inst__0w_mem_10__31_0__31_) );
  OR2X2 OR2X2_2936 ( .A(w_mem_inst__abc_21378_n4311), .B(w_mem_inst__abc_21378_n4309), .Y(w_mem_inst__abc_21378_n4312) );
  OR2X2 OR2X2_2937 ( .A(w_mem_inst__abc_21378_n4312), .B(w_mem_inst__abc_21378_n4308), .Y(w_mem_inst__0w_mem_9__31_0__0_) );
  OR2X2 OR2X2_2938 ( .A(w_mem_inst__abc_21378_n4317), .B(w_mem_inst__abc_21378_n4315), .Y(w_mem_inst__abc_21378_n4318) );
  OR2X2 OR2X2_2939 ( .A(w_mem_inst__abc_21378_n4318), .B(w_mem_inst__abc_21378_n4314), .Y(w_mem_inst__0w_mem_9__31_0__1_) );
  OR2X2 OR2X2_294 ( .A(_abc_15724_n851_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_70_), .Y(_abc_15724_n1598) );
  OR2X2 OR2X2_2940 ( .A(w_mem_inst__abc_21378_n4323), .B(w_mem_inst__abc_21378_n4321), .Y(w_mem_inst__abc_21378_n4324) );
  OR2X2 OR2X2_2941 ( .A(w_mem_inst__abc_21378_n4324), .B(w_mem_inst__abc_21378_n4320), .Y(w_mem_inst__0w_mem_9__31_0__2_) );
  OR2X2 OR2X2_2942 ( .A(w_mem_inst__abc_21378_n4329), .B(w_mem_inst__abc_21378_n4327), .Y(w_mem_inst__abc_21378_n4330) );
  OR2X2 OR2X2_2943 ( .A(w_mem_inst__abc_21378_n4330), .B(w_mem_inst__abc_21378_n4326), .Y(w_mem_inst__0w_mem_9__31_0__3_) );
  OR2X2 OR2X2_2944 ( .A(w_mem_inst__abc_21378_n4335), .B(w_mem_inst__abc_21378_n4333), .Y(w_mem_inst__abc_21378_n4336) );
  OR2X2 OR2X2_2945 ( .A(w_mem_inst__abc_21378_n4336), .B(w_mem_inst__abc_21378_n4332), .Y(w_mem_inst__0w_mem_9__31_0__4_) );
  OR2X2 OR2X2_2946 ( .A(w_mem_inst__abc_21378_n4341), .B(w_mem_inst__abc_21378_n4339), .Y(w_mem_inst__abc_21378_n4342) );
  OR2X2 OR2X2_2947 ( .A(w_mem_inst__abc_21378_n4342), .B(w_mem_inst__abc_21378_n4338), .Y(w_mem_inst__0w_mem_9__31_0__5_) );
  OR2X2 OR2X2_2948 ( .A(w_mem_inst__abc_21378_n4347), .B(w_mem_inst__abc_21378_n4345), .Y(w_mem_inst__abc_21378_n4348) );
  OR2X2 OR2X2_2949 ( .A(w_mem_inst__abc_21378_n4348), .B(w_mem_inst__abc_21378_n4344), .Y(w_mem_inst__0w_mem_9__31_0__6_) );
  OR2X2 OR2X2_295 ( .A(_abc_15724_n1597_1), .B(_abc_15724_n1599_1), .Y(H2_reg_6__FF_INPUT) );
  OR2X2 OR2X2_2950 ( .A(w_mem_inst__abc_21378_n4353), .B(w_mem_inst__abc_21378_n4351), .Y(w_mem_inst__abc_21378_n4354) );
  OR2X2 OR2X2_2951 ( .A(w_mem_inst__abc_21378_n4354), .B(w_mem_inst__abc_21378_n4350), .Y(w_mem_inst__0w_mem_9__31_0__7_) );
  OR2X2 OR2X2_2952 ( .A(w_mem_inst__abc_21378_n4359), .B(w_mem_inst__abc_21378_n4357), .Y(w_mem_inst__abc_21378_n4360) );
  OR2X2 OR2X2_2953 ( .A(w_mem_inst__abc_21378_n4360), .B(w_mem_inst__abc_21378_n4356), .Y(w_mem_inst__0w_mem_9__31_0__8_) );
  OR2X2 OR2X2_2954 ( .A(w_mem_inst__abc_21378_n4365), .B(w_mem_inst__abc_21378_n4363), .Y(w_mem_inst__abc_21378_n4366) );
  OR2X2 OR2X2_2955 ( .A(w_mem_inst__abc_21378_n4366), .B(w_mem_inst__abc_21378_n4362), .Y(w_mem_inst__0w_mem_9__31_0__9_) );
  OR2X2 OR2X2_2956 ( .A(w_mem_inst__abc_21378_n4371), .B(w_mem_inst__abc_21378_n4369), .Y(w_mem_inst__abc_21378_n4372) );
  OR2X2 OR2X2_2957 ( .A(w_mem_inst__abc_21378_n4372), .B(w_mem_inst__abc_21378_n4368), .Y(w_mem_inst__0w_mem_9__31_0__10_) );
  OR2X2 OR2X2_2958 ( .A(w_mem_inst__abc_21378_n4377), .B(w_mem_inst__abc_21378_n4375), .Y(w_mem_inst__abc_21378_n4378) );
  OR2X2 OR2X2_2959 ( .A(w_mem_inst__abc_21378_n4378), .B(w_mem_inst__abc_21378_n4374), .Y(w_mem_inst__0w_mem_9__31_0__11_) );
  OR2X2 OR2X2_296 ( .A(_auto_iopadmap_cc_313_execute_26059_71_), .B(c_reg_7_), .Y(_abc_15724_n1603_1) );
  OR2X2 OR2X2_2960 ( .A(w_mem_inst__abc_21378_n4383), .B(w_mem_inst__abc_21378_n4381), .Y(w_mem_inst__abc_21378_n4384) );
  OR2X2 OR2X2_2961 ( .A(w_mem_inst__abc_21378_n4384), .B(w_mem_inst__abc_21378_n4380), .Y(w_mem_inst__0w_mem_9__31_0__12_) );
  OR2X2 OR2X2_2962 ( .A(w_mem_inst__abc_21378_n4389), .B(w_mem_inst__abc_21378_n4387), .Y(w_mem_inst__abc_21378_n4390) );
  OR2X2 OR2X2_2963 ( .A(w_mem_inst__abc_21378_n4390), .B(w_mem_inst__abc_21378_n4386), .Y(w_mem_inst__0w_mem_9__31_0__13_) );
  OR2X2 OR2X2_2964 ( .A(w_mem_inst__abc_21378_n4395), .B(w_mem_inst__abc_21378_n4393), .Y(w_mem_inst__abc_21378_n4396) );
  OR2X2 OR2X2_2965 ( .A(w_mem_inst__abc_21378_n4396), .B(w_mem_inst__abc_21378_n4392), .Y(w_mem_inst__0w_mem_9__31_0__14_) );
  OR2X2 OR2X2_2966 ( .A(w_mem_inst__abc_21378_n4401), .B(w_mem_inst__abc_21378_n4399), .Y(w_mem_inst__abc_21378_n4402) );
  OR2X2 OR2X2_2967 ( .A(w_mem_inst__abc_21378_n4402), .B(w_mem_inst__abc_21378_n4398), .Y(w_mem_inst__0w_mem_9__31_0__15_) );
  OR2X2 OR2X2_2968 ( .A(w_mem_inst__abc_21378_n4407), .B(w_mem_inst__abc_21378_n4405), .Y(w_mem_inst__abc_21378_n4408) );
  OR2X2 OR2X2_2969 ( .A(w_mem_inst__abc_21378_n4408), .B(w_mem_inst__abc_21378_n4404), .Y(w_mem_inst__0w_mem_9__31_0__16_) );
  OR2X2 OR2X2_297 ( .A(_abc_15724_n1602_1), .B(_abc_15724_n1606), .Y(_abc_15724_n1607) );
  OR2X2 OR2X2_2970 ( .A(w_mem_inst__abc_21378_n4413), .B(w_mem_inst__abc_21378_n4411), .Y(w_mem_inst__abc_21378_n4414) );
  OR2X2 OR2X2_2971 ( .A(w_mem_inst__abc_21378_n4414), .B(w_mem_inst__abc_21378_n4410), .Y(w_mem_inst__0w_mem_9__31_0__17_) );
  OR2X2 OR2X2_2972 ( .A(w_mem_inst__abc_21378_n4419), .B(w_mem_inst__abc_21378_n4417), .Y(w_mem_inst__abc_21378_n4420) );
  OR2X2 OR2X2_2973 ( .A(w_mem_inst__abc_21378_n4420), .B(w_mem_inst__abc_21378_n4416), .Y(w_mem_inst__0w_mem_9__31_0__18_) );
  OR2X2 OR2X2_2974 ( .A(w_mem_inst__abc_21378_n4425), .B(w_mem_inst__abc_21378_n4423), .Y(w_mem_inst__abc_21378_n4426) );
  OR2X2 OR2X2_2975 ( .A(w_mem_inst__abc_21378_n4426), .B(w_mem_inst__abc_21378_n4422), .Y(w_mem_inst__0w_mem_9__31_0__19_) );
  OR2X2 OR2X2_2976 ( .A(w_mem_inst__abc_21378_n4431), .B(w_mem_inst__abc_21378_n4429), .Y(w_mem_inst__abc_21378_n4432) );
  OR2X2 OR2X2_2977 ( .A(w_mem_inst__abc_21378_n4432), .B(w_mem_inst__abc_21378_n4428), .Y(w_mem_inst__0w_mem_9__31_0__20_) );
  OR2X2 OR2X2_2978 ( .A(w_mem_inst__abc_21378_n4437), .B(w_mem_inst__abc_21378_n4435), .Y(w_mem_inst__abc_21378_n4438) );
  OR2X2 OR2X2_2979 ( .A(w_mem_inst__abc_21378_n4438), .B(w_mem_inst__abc_21378_n4434), .Y(w_mem_inst__0w_mem_9__31_0__21_) );
  OR2X2 OR2X2_298 ( .A(_abc_15724_n1601), .B(_abc_15724_n1608), .Y(_abc_15724_n1609_1) );
  OR2X2 OR2X2_2980 ( .A(w_mem_inst__abc_21378_n4443), .B(w_mem_inst__abc_21378_n4441), .Y(w_mem_inst__abc_21378_n4444) );
  OR2X2 OR2X2_2981 ( .A(w_mem_inst__abc_21378_n4444), .B(w_mem_inst__abc_21378_n4440), .Y(w_mem_inst__0w_mem_9__31_0__22_) );
  OR2X2 OR2X2_2982 ( .A(w_mem_inst__abc_21378_n4449), .B(w_mem_inst__abc_21378_n4447), .Y(w_mem_inst__abc_21378_n4450) );
  OR2X2 OR2X2_2983 ( .A(w_mem_inst__abc_21378_n4450), .B(w_mem_inst__abc_21378_n4446), .Y(w_mem_inst__0w_mem_9__31_0__23_) );
  OR2X2 OR2X2_2984 ( .A(w_mem_inst__abc_21378_n4455), .B(w_mem_inst__abc_21378_n4453), .Y(w_mem_inst__abc_21378_n4456) );
  OR2X2 OR2X2_2985 ( .A(w_mem_inst__abc_21378_n4456), .B(w_mem_inst__abc_21378_n4452), .Y(w_mem_inst__0w_mem_9__31_0__24_) );
  OR2X2 OR2X2_2986 ( .A(w_mem_inst__abc_21378_n4461), .B(w_mem_inst__abc_21378_n4459), .Y(w_mem_inst__abc_21378_n4462) );
  OR2X2 OR2X2_2987 ( .A(w_mem_inst__abc_21378_n4462), .B(w_mem_inst__abc_21378_n4458), .Y(w_mem_inst__0w_mem_9__31_0__25_) );
  OR2X2 OR2X2_2988 ( .A(w_mem_inst__abc_21378_n4467), .B(w_mem_inst__abc_21378_n4465), .Y(w_mem_inst__abc_21378_n4468) );
  OR2X2 OR2X2_2989 ( .A(w_mem_inst__abc_21378_n4468), .B(w_mem_inst__abc_21378_n4464), .Y(w_mem_inst__0w_mem_9__31_0__26_) );
  OR2X2 OR2X2_299 ( .A(_abc_15724_n851_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_71_), .Y(_abc_15724_n1612) );
  OR2X2 OR2X2_2990 ( .A(w_mem_inst__abc_21378_n4473), .B(w_mem_inst__abc_21378_n4471), .Y(w_mem_inst__abc_21378_n4474) );
  OR2X2 OR2X2_2991 ( .A(w_mem_inst__abc_21378_n4474), .B(w_mem_inst__abc_21378_n4470), .Y(w_mem_inst__0w_mem_9__31_0__27_) );
  OR2X2 OR2X2_2992 ( .A(w_mem_inst__abc_21378_n4479), .B(w_mem_inst__abc_21378_n4477), .Y(w_mem_inst__abc_21378_n4480) );
  OR2X2 OR2X2_2993 ( .A(w_mem_inst__abc_21378_n4480), .B(w_mem_inst__abc_21378_n4476), .Y(w_mem_inst__0w_mem_9__31_0__28_) );
  OR2X2 OR2X2_2994 ( .A(w_mem_inst__abc_21378_n4485), .B(w_mem_inst__abc_21378_n4483), .Y(w_mem_inst__abc_21378_n4486) );
  OR2X2 OR2X2_2995 ( .A(w_mem_inst__abc_21378_n4486), .B(w_mem_inst__abc_21378_n4482), .Y(w_mem_inst__0w_mem_9__31_0__29_) );
  OR2X2 OR2X2_2996 ( .A(w_mem_inst__abc_21378_n4491), .B(w_mem_inst__abc_21378_n4489), .Y(w_mem_inst__abc_21378_n4492) );
  OR2X2 OR2X2_2997 ( .A(w_mem_inst__abc_21378_n4492), .B(w_mem_inst__abc_21378_n4488), .Y(w_mem_inst__0w_mem_9__31_0__30_) );
  OR2X2 OR2X2_2998 ( .A(w_mem_inst__abc_21378_n4497), .B(w_mem_inst__abc_21378_n4495), .Y(w_mem_inst__abc_21378_n4498) );
  OR2X2 OR2X2_2999 ( .A(w_mem_inst__abc_21378_n4498), .B(w_mem_inst__abc_21378_n4494), .Y(w_mem_inst__0w_mem_9__31_0__31_) );
  OR2X2 OR2X2_3 ( .A(e_reg_19_), .B(_auto_iopadmap_cc_313_execute_26059_19_), .Y(_abc_15724_n707) );
  OR2X2 OR2X2_30 ( .A(_auto_iopadmap_cc_313_execute_26059_4_), .B(e_reg_4_), .Y(_abc_15724_n807) );
  OR2X2 OR2X2_300 ( .A(_abc_15724_n1611), .B(_abc_15724_n1613), .Y(H2_reg_7__FF_INPUT) );
  OR2X2 OR2X2_3000 ( .A(w_mem_inst__abc_21378_n4503), .B(w_mem_inst__abc_21378_n4501), .Y(w_mem_inst__abc_21378_n4504) );
  OR2X2 OR2X2_3001 ( .A(w_mem_inst__abc_21378_n4504), .B(w_mem_inst__abc_21378_n4500), .Y(w_mem_inst__0w_mem_8__31_0__0_) );
  OR2X2 OR2X2_3002 ( .A(w_mem_inst__abc_21378_n4509), .B(w_mem_inst__abc_21378_n4507), .Y(w_mem_inst__abc_21378_n4510) );
  OR2X2 OR2X2_3003 ( .A(w_mem_inst__abc_21378_n4510), .B(w_mem_inst__abc_21378_n4506), .Y(w_mem_inst__0w_mem_8__31_0__1_) );
  OR2X2 OR2X2_3004 ( .A(w_mem_inst__abc_21378_n4515), .B(w_mem_inst__abc_21378_n4513), .Y(w_mem_inst__abc_21378_n4516) );
  OR2X2 OR2X2_3005 ( .A(w_mem_inst__abc_21378_n4516), .B(w_mem_inst__abc_21378_n4512), .Y(w_mem_inst__0w_mem_8__31_0__2_) );
  OR2X2 OR2X2_3006 ( .A(w_mem_inst__abc_21378_n4521), .B(w_mem_inst__abc_21378_n4519), .Y(w_mem_inst__abc_21378_n4522) );
  OR2X2 OR2X2_3007 ( .A(w_mem_inst__abc_21378_n4522), .B(w_mem_inst__abc_21378_n4518), .Y(w_mem_inst__0w_mem_8__31_0__3_) );
  OR2X2 OR2X2_3008 ( .A(w_mem_inst__abc_21378_n4527), .B(w_mem_inst__abc_21378_n4525), .Y(w_mem_inst__abc_21378_n4528) );
  OR2X2 OR2X2_3009 ( .A(w_mem_inst__abc_21378_n4528), .B(w_mem_inst__abc_21378_n4524), .Y(w_mem_inst__0w_mem_8__31_0__4_) );
  OR2X2 OR2X2_301 ( .A(_auto_iopadmap_cc_313_execute_26059_72_), .B(c_reg_8_), .Y(_abc_15724_n1616_1) );
  OR2X2 OR2X2_3010 ( .A(w_mem_inst__abc_21378_n4533), .B(w_mem_inst__abc_21378_n4531), .Y(w_mem_inst__abc_21378_n4534) );
  OR2X2 OR2X2_3011 ( .A(w_mem_inst__abc_21378_n4534), .B(w_mem_inst__abc_21378_n4530), .Y(w_mem_inst__0w_mem_8__31_0__5_) );
  OR2X2 OR2X2_3012 ( .A(w_mem_inst__abc_21378_n4539), .B(w_mem_inst__abc_21378_n4537), .Y(w_mem_inst__abc_21378_n4540) );
  OR2X2 OR2X2_3013 ( .A(w_mem_inst__abc_21378_n4540), .B(w_mem_inst__abc_21378_n4536), .Y(w_mem_inst__0w_mem_8__31_0__6_) );
  OR2X2 OR2X2_3014 ( .A(w_mem_inst__abc_21378_n4545), .B(w_mem_inst__abc_21378_n4543), .Y(w_mem_inst__abc_21378_n4546) );
  OR2X2 OR2X2_3015 ( .A(w_mem_inst__abc_21378_n4546), .B(w_mem_inst__abc_21378_n4542), .Y(w_mem_inst__0w_mem_8__31_0__7_) );
  OR2X2 OR2X2_3016 ( .A(w_mem_inst__abc_21378_n4551), .B(w_mem_inst__abc_21378_n4549), .Y(w_mem_inst__abc_21378_n4552) );
  OR2X2 OR2X2_3017 ( .A(w_mem_inst__abc_21378_n4552), .B(w_mem_inst__abc_21378_n4548), .Y(w_mem_inst__0w_mem_8__31_0__8_) );
  OR2X2 OR2X2_3018 ( .A(w_mem_inst__abc_21378_n4557), .B(w_mem_inst__abc_21378_n4555), .Y(w_mem_inst__abc_21378_n4558) );
  OR2X2 OR2X2_3019 ( .A(w_mem_inst__abc_21378_n4558), .B(w_mem_inst__abc_21378_n4554), .Y(w_mem_inst__0w_mem_8__31_0__9_) );
  OR2X2 OR2X2_302 ( .A(_abc_15724_n1622), .B(_abc_15724_n1620), .Y(_abc_15724_n1623_1) );
  OR2X2 OR2X2_3020 ( .A(w_mem_inst__abc_21378_n4563), .B(w_mem_inst__abc_21378_n4561), .Y(w_mem_inst__abc_21378_n4564) );
  OR2X2 OR2X2_3021 ( .A(w_mem_inst__abc_21378_n4564), .B(w_mem_inst__abc_21378_n4560), .Y(w_mem_inst__0w_mem_8__31_0__10_) );
  OR2X2 OR2X2_3022 ( .A(w_mem_inst__abc_21378_n4569), .B(w_mem_inst__abc_21378_n4567), .Y(w_mem_inst__abc_21378_n4570) );
  OR2X2 OR2X2_3023 ( .A(w_mem_inst__abc_21378_n4570), .B(w_mem_inst__abc_21378_n4566), .Y(w_mem_inst__0w_mem_8__31_0__11_) );
  OR2X2 OR2X2_3024 ( .A(w_mem_inst__abc_21378_n4575), .B(w_mem_inst__abc_21378_n4573), .Y(w_mem_inst__abc_21378_n4576) );
  OR2X2 OR2X2_3025 ( .A(w_mem_inst__abc_21378_n4576), .B(w_mem_inst__abc_21378_n4572), .Y(w_mem_inst__0w_mem_8__31_0__12_) );
  OR2X2 OR2X2_3026 ( .A(w_mem_inst__abc_21378_n4581), .B(w_mem_inst__abc_21378_n4579), .Y(w_mem_inst__abc_21378_n4582) );
  OR2X2 OR2X2_3027 ( .A(w_mem_inst__abc_21378_n4582), .B(w_mem_inst__abc_21378_n4578), .Y(w_mem_inst__0w_mem_8__31_0__13_) );
  OR2X2 OR2X2_3028 ( .A(w_mem_inst__abc_21378_n4587), .B(w_mem_inst__abc_21378_n4585), .Y(w_mem_inst__abc_21378_n4588) );
  OR2X2 OR2X2_3029 ( .A(w_mem_inst__abc_21378_n4588), .B(w_mem_inst__abc_21378_n4584), .Y(w_mem_inst__0w_mem_8__31_0__14_) );
  OR2X2 OR2X2_303 ( .A(_abc_15724_n1624_1), .B(_abc_15724_n1619), .Y(_abc_15724_n1625) );
  OR2X2 OR2X2_3030 ( .A(w_mem_inst__abc_21378_n4593), .B(w_mem_inst__abc_21378_n4591), .Y(w_mem_inst__abc_21378_n4594) );
  OR2X2 OR2X2_3031 ( .A(w_mem_inst__abc_21378_n4594), .B(w_mem_inst__abc_21378_n4590), .Y(w_mem_inst__0w_mem_8__31_0__15_) );
  OR2X2 OR2X2_3032 ( .A(w_mem_inst__abc_21378_n4599), .B(w_mem_inst__abc_21378_n4597), .Y(w_mem_inst__abc_21378_n4600) );
  OR2X2 OR2X2_3033 ( .A(w_mem_inst__abc_21378_n4600), .B(w_mem_inst__abc_21378_n4596), .Y(w_mem_inst__0w_mem_8__31_0__16_) );
  OR2X2 OR2X2_3034 ( .A(w_mem_inst__abc_21378_n4605), .B(w_mem_inst__abc_21378_n4603), .Y(w_mem_inst__abc_21378_n4606) );
  OR2X2 OR2X2_3035 ( .A(w_mem_inst__abc_21378_n4606), .B(w_mem_inst__abc_21378_n4602), .Y(w_mem_inst__0w_mem_8__31_0__17_) );
  OR2X2 OR2X2_3036 ( .A(w_mem_inst__abc_21378_n4611), .B(w_mem_inst__abc_21378_n4609), .Y(w_mem_inst__abc_21378_n4612) );
  OR2X2 OR2X2_3037 ( .A(w_mem_inst__abc_21378_n4612), .B(w_mem_inst__abc_21378_n4608), .Y(w_mem_inst__0w_mem_8__31_0__18_) );
  OR2X2 OR2X2_3038 ( .A(w_mem_inst__abc_21378_n4617), .B(w_mem_inst__abc_21378_n4615), .Y(w_mem_inst__abc_21378_n4618) );
  OR2X2 OR2X2_3039 ( .A(w_mem_inst__abc_21378_n4618), .B(w_mem_inst__abc_21378_n4614), .Y(w_mem_inst__0w_mem_8__31_0__19_) );
  OR2X2 OR2X2_304 ( .A(_abc_15724_n1629), .B(_abc_15724_n1615), .Y(H2_reg_8__FF_INPUT) );
  OR2X2 OR2X2_3040 ( .A(w_mem_inst__abc_21378_n4623), .B(w_mem_inst__abc_21378_n4621), .Y(w_mem_inst__abc_21378_n4624) );
  OR2X2 OR2X2_3041 ( .A(w_mem_inst__abc_21378_n4624), .B(w_mem_inst__abc_21378_n4620), .Y(w_mem_inst__0w_mem_8__31_0__20_) );
  OR2X2 OR2X2_3042 ( .A(w_mem_inst__abc_21378_n4629), .B(w_mem_inst__abc_21378_n4627), .Y(w_mem_inst__abc_21378_n4630) );
  OR2X2 OR2X2_3043 ( .A(w_mem_inst__abc_21378_n4630), .B(w_mem_inst__abc_21378_n4626), .Y(w_mem_inst__0w_mem_8__31_0__21_) );
  OR2X2 OR2X2_3044 ( .A(w_mem_inst__abc_21378_n4635), .B(w_mem_inst__abc_21378_n4633), .Y(w_mem_inst__abc_21378_n4636) );
  OR2X2 OR2X2_3045 ( .A(w_mem_inst__abc_21378_n4636), .B(w_mem_inst__abc_21378_n4632), .Y(w_mem_inst__0w_mem_8__31_0__22_) );
  OR2X2 OR2X2_3046 ( .A(w_mem_inst__abc_21378_n4641), .B(w_mem_inst__abc_21378_n4639), .Y(w_mem_inst__abc_21378_n4642) );
  OR2X2 OR2X2_3047 ( .A(w_mem_inst__abc_21378_n4642), .B(w_mem_inst__abc_21378_n4638), .Y(w_mem_inst__0w_mem_8__31_0__23_) );
  OR2X2 OR2X2_3048 ( .A(w_mem_inst__abc_21378_n4647), .B(w_mem_inst__abc_21378_n4645), .Y(w_mem_inst__abc_21378_n4648) );
  OR2X2 OR2X2_3049 ( .A(w_mem_inst__abc_21378_n4648), .B(w_mem_inst__abc_21378_n4644), .Y(w_mem_inst__0w_mem_8__31_0__24_) );
  OR2X2 OR2X2_305 ( .A(_auto_iopadmap_cc_313_execute_26059_73_), .B(c_reg_9_), .Y(_abc_15724_n1631_1) );
  OR2X2 OR2X2_3050 ( .A(w_mem_inst__abc_21378_n4653), .B(w_mem_inst__abc_21378_n4651), .Y(w_mem_inst__abc_21378_n4654) );
  OR2X2 OR2X2_3051 ( .A(w_mem_inst__abc_21378_n4654), .B(w_mem_inst__abc_21378_n4650), .Y(w_mem_inst__0w_mem_8__31_0__25_) );
  OR2X2 OR2X2_3052 ( .A(w_mem_inst__abc_21378_n4659), .B(w_mem_inst__abc_21378_n4657), .Y(w_mem_inst__abc_21378_n4660) );
  OR2X2 OR2X2_3053 ( .A(w_mem_inst__abc_21378_n4660), .B(w_mem_inst__abc_21378_n4656), .Y(w_mem_inst__0w_mem_8__31_0__26_) );
  OR2X2 OR2X2_3054 ( .A(w_mem_inst__abc_21378_n4665), .B(w_mem_inst__abc_21378_n4663), .Y(w_mem_inst__abc_21378_n4666) );
  OR2X2 OR2X2_3055 ( .A(w_mem_inst__abc_21378_n4666), .B(w_mem_inst__abc_21378_n4662), .Y(w_mem_inst__0w_mem_8__31_0__27_) );
  OR2X2 OR2X2_3056 ( .A(w_mem_inst__abc_21378_n4671), .B(w_mem_inst__abc_21378_n4669), .Y(w_mem_inst__abc_21378_n4672) );
  OR2X2 OR2X2_3057 ( .A(w_mem_inst__abc_21378_n4672), .B(w_mem_inst__abc_21378_n4668), .Y(w_mem_inst__0w_mem_8__31_0__28_) );
  OR2X2 OR2X2_3058 ( .A(w_mem_inst__abc_21378_n4677), .B(w_mem_inst__abc_21378_n4675), .Y(w_mem_inst__abc_21378_n4678) );
  OR2X2 OR2X2_3059 ( .A(w_mem_inst__abc_21378_n4678), .B(w_mem_inst__abc_21378_n4674), .Y(w_mem_inst__0w_mem_8__31_0__29_) );
  OR2X2 OR2X2_306 ( .A(_abc_15724_n1636_1), .B(_abc_15724_n1634), .Y(_abc_15724_n1637_1) );
  OR2X2 OR2X2_3060 ( .A(w_mem_inst__abc_21378_n4683), .B(w_mem_inst__abc_21378_n4681), .Y(w_mem_inst__abc_21378_n4684) );
  OR2X2 OR2X2_3061 ( .A(w_mem_inst__abc_21378_n4684), .B(w_mem_inst__abc_21378_n4680), .Y(w_mem_inst__0w_mem_8__31_0__30_) );
  OR2X2 OR2X2_3062 ( .A(w_mem_inst__abc_21378_n4689), .B(w_mem_inst__abc_21378_n4687), .Y(w_mem_inst__abc_21378_n4690) );
  OR2X2 OR2X2_3063 ( .A(w_mem_inst__abc_21378_n4690), .B(w_mem_inst__abc_21378_n4686), .Y(w_mem_inst__0w_mem_8__31_0__31_) );
  OR2X2 OR2X2_3064 ( .A(w_mem_inst__abc_21378_n4695), .B(w_mem_inst__abc_21378_n4693), .Y(w_mem_inst__abc_21378_n4696) );
  OR2X2 OR2X2_3065 ( .A(w_mem_inst__abc_21378_n4696), .B(w_mem_inst__abc_21378_n4692), .Y(w_mem_inst__0w_mem_7__31_0__0_) );
  OR2X2 OR2X2_3066 ( .A(w_mem_inst__abc_21378_n4701), .B(w_mem_inst__abc_21378_n4699), .Y(w_mem_inst__abc_21378_n4702) );
  OR2X2 OR2X2_3067 ( .A(w_mem_inst__abc_21378_n4702), .B(w_mem_inst__abc_21378_n4698), .Y(w_mem_inst__0w_mem_7__31_0__1_) );
  OR2X2 OR2X2_3068 ( .A(w_mem_inst__abc_21378_n4707), .B(w_mem_inst__abc_21378_n4705), .Y(w_mem_inst__abc_21378_n4708) );
  OR2X2 OR2X2_3069 ( .A(w_mem_inst__abc_21378_n4708), .B(w_mem_inst__abc_21378_n4704), .Y(w_mem_inst__0w_mem_7__31_0__2_) );
  OR2X2 OR2X2_307 ( .A(_abc_15724_n1641), .B(_abc_15724_n1642_1), .Y(H2_reg_9__FF_INPUT) );
  OR2X2 OR2X2_3070 ( .A(w_mem_inst__abc_21378_n4713), .B(w_mem_inst__abc_21378_n4711), .Y(w_mem_inst__abc_21378_n4714) );
  OR2X2 OR2X2_3071 ( .A(w_mem_inst__abc_21378_n4714), .B(w_mem_inst__abc_21378_n4710), .Y(w_mem_inst__0w_mem_7__31_0__3_) );
  OR2X2 OR2X2_3072 ( .A(w_mem_inst__abc_21378_n4719), .B(w_mem_inst__abc_21378_n4717), .Y(w_mem_inst__abc_21378_n4720) );
  OR2X2 OR2X2_3073 ( .A(w_mem_inst__abc_21378_n4720), .B(w_mem_inst__abc_21378_n4716), .Y(w_mem_inst__0w_mem_7__31_0__4_) );
  OR2X2 OR2X2_3074 ( .A(w_mem_inst__abc_21378_n4725), .B(w_mem_inst__abc_21378_n4723), .Y(w_mem_inst__abc_21378_n4726) );
  OR2X2 OR2X2_3075 ( .A(w_mem_inst__abc_21378_n4726), .B(w_mem_inst__abc_21378_n4722), .Y(w_mem_inst__0w_mem_7__31_0__5_) );
  OR2X2 OR2X2_3076 ( .A(w_mem_inst__abc_21378_n4731), .B(w_mem_inst__abc_21378_n4729), .Y(w_mem_inst__abc_21378_n4732) );
  OR2X2 OR2X2_3077 ( .A(w_mem_inst__abc_21378_n4732), .B(w_mem_inst__abc_21378_n4728), .Y(w_mem_inst__0w_mem_7__31_0__6_) );
  OR2X2 OR2X2_3078 ( .A(w_mem_inst__abc_21378_n4737), .B(w_mem_inst__abc_21378_n4735), .Y(w_mem_inst__abc_21378_n4738) );
  OR2X2 OR2X2_3079 ( .A(w_mem_inst__abc_21378_n4738), .B(w_mem_inst__abc_21378_n4734), .Y(w_mem_inst__0w_mem_7__31_0__7_) );
  OR2X2 OR2X2_308 ( .A(_auto_iopadmap_cc_313_execute_26059_74_), .B(c_reg_10_), .Y(_abc_15724_n1646) );
  OR2X2 OR2X2_3080 ( .A(w_mem_inst__abc_21378_n4743), .B(w_mem_inst__abc_21378_n4741), .Y(w_mem_inst__abc_21378_n4744) );
  OR2X2 OR2X2_3081 ( .A(w_mem_inst__abc_21378_n4744), .B(w_mem_inst__abc_21378_n4740), .Y(w_mem_inst__0w_mem_7__31_0__8_) );
  OR2X2 OR2X2_3082 ( .A(w_mem_inst__abc_21378_n4749), .B(w_mem_inst__abc_21378_n4747), .Y(w_mem_inst__abc_21378_n4750) );
  OR2X2 OR2X2_3083 ( .A(w_mem_inst__abc_21378_n4750), .B(w_mem_inst__abc_21378_n4746), .Y(w_mem_inst__0w_mem_7__31_0__9_) );
  OR2X2 OR2X2_3084 ( .A(w_mem_inst__abc_21378_n4755), .B(w_mem_inst__abc_21378_n4753), .Y(w_mem_inst__abc_21378_n4756) );
  OR2X2 OR2X2_3085 ( .A(w_mem_inst__abc_21378_n4756), .B(w_mem_inst__abc_21378_n4752), .Y(w_mem_inst__0w_mem_7__31_0__10_) );
  OR2X2 OR2X2_3086 ( .A(w_mem_inst__abc_21378_n4761), .B(w_mem_inst__abc_21378_n4759), .Y(w_mem_inst__abc_21378_n4762) );
  OR2X2 OR2X2_3087 ( .A(w_mem_inst__abc_21378_n4762), .B(w_mem_inst__abc_21378_n4758), .Y(w_mem_inst__0w_mem_7__31_0__11_) );
  OR2X2 OR2X2_3088 ( .A(w_mem_inst__abc_21378_n4767), .B(w_mem_inst__abc_21378_n4765), .Y(w_mem_inst__abc_21378_n4768) );
  OR2X2 OR2X2_3089 ( .A(w_mem_inst__abc_21378_n4768), .B(w_mem_inst__abc_21378_n4764), .Y(w_mem_inst__0w_mem_7__31_0__12_) );
  OR2X2 OR2X2_309 ( .A(_abc_15724_n1645_1), .B(_abc_15724_n1649_1), .Y(_abc_15724_n1650) );
  OR2X2 OR2X2_3090 ( .A(w_mem_inst__abc_21378_n4773), .B(w_mem_inst__abc_21378_n4771), .Y(w_mem_inst__abc_21378_n4774) );
  OR2X2 OR2X2_3091 ( .A(w_mem_inst__abc_21378_n4774), .B(w_mem_inst__abc_21378_n4770), .Y(w_mem_inst__0w_mem_7__31_0__13_) );
  OR2X2 OR2X2_3092 ( .A(w_mem_inst__abc_21378_n4779), .B(w_mem_inst__abc_21378_n4777), .Y(w_mem_inst__abc_21378_n4780) );
  OR2X2 OR2X2_3093 ( .A(w_mem_inst__abc_21378_n4780), .B(w_mem_inst__abc_21378_n4776), .Y(w_mem_inst__0w_mem_7__31_0__14_) );
  OR2X2 OR2X2_3094 ( .A(w_mem_inst__abc_21378_n4785), .B(w_mem_inst__abc_21378_n4783), .Y(w_mem_inst__abc_21378_n4786) );
  OR2X2 OR2X2_3095 ( .A(w_mem_inst__abc_21378_n4786), .B(w_mem_inst__abc_21378_n4782), .Y(w_mem_inst__0w_mem_7__31_0__15_) );
  OR2X2 OR2X2_3096 ( .A(w_mem_inst__abc_21378_n4791), .B(w_mem_inst__abc_21378_n4789), .Y(w_mem_inst__abc_21378_n4792) );
  OR2X2 OR2X2_3097 ( .A(w_mem_inst__abc_21378_n4792), .B(w_mem_inst__abc_21378_n4788), .Y(w_mem_inst__0w_mem_7__31_0__16_) );
  OR2X2 OR2X2_3098 ( .A(w_mem_inst__abc_21378_n4797), .B(w_mem_inst__abc_21378_n4795), .Y(w_mem_inst__abc_21378_n4798) );
  OR2X2 OR2X2_3099 ( .A(w_mem_inst__abc_21378_n4798), .B(w_mem_inst__abc_21378_n4794), .Y(w_mem_inst__0w_mem_7__31_0__17_) );
  OR2X2 OR2X2_31 ( .A(_abc_15724_n809), .B(_abc_15724_n786), .Y(_abc_15724_n810) );
  OR2X2 OR2X2_310 ( .A(_abc_15724_n851_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_74_), .Y(_abc_15724_n1655_1) );
  OR2X2 OR2X2_3100 ( .A(w_mem_inst__abc_21378_n4803), .B(w_mem_inst__abc_21378_n4801), .Y(w_mem_inst__abc_21378_n4804) );
  OR2X2 OR2X2_3101 ( .A(w_mem_inst__abc_21378_n4804), .B(w_mem_inst__abc_21378_n4800), .Y(w_mem_inst__0w_mem_7__31_0__18_) );
  OR2X2 OR2X2_3102 ( .A(w_mem_inst__abc_21378_n4809), .B(w_mem_inst__abc_21378_n4807), .Y(w_mem_inst__abc_21378_n4810) );
  OR2X2 OR2X2_3103 ( .A(w_mem_inst__abc_21378_n4810), .B(w_mem_inst__abc_21378_n4806), .Y(w_mem_inst__0w_mem_7__31_0__19_) );
  OR2X2 OR2X2_3104 ( .A(w_mem_inst__abc_21378_n4815), .B(w_mem_inst__abc_21378_n4813), .Y(w_mem_inst__abc_21378_n4816) );
  OR2X2 OR2X2_3105 ( .A(w_mem_inst__abc_21378_n4816), .B(w_mem_inst__abc_21378_n4812), .Y(w_mem_inst__0w_mem_7__31_0__20_) );
  OR2X2 OR2X2_3106 ( .A(w_mem_inst__abc_21378_n4821), .B(w_mem_inst__abc_21378_n4819), .Y(w_mem_inst__abc_21378_n4822) );
  OR2X2 OR2X2_3107 ( .A(w_mem_inst__abc_21378_n4822), .B(w_mem_inst__abc_21378_n4818), .Y(w_mem_inst__0w_mem_7__31_0__21_) );
  OR2X2 OR2X2_3108 ( .A(w_mem_inst__abc_21378_n4827), .B(w_mem_inst__abc_21378_n4825), .Y(w_mem_inst__abc_21378_n4828) );
  OR2X2 OR2X2_3109 ( .A(w_mem_inst__abc_21378_n4828), .B(w_mem_inst__abc_21378_n4824), .Y(w_mem_inst__0w_mem_7__31_0__22_) );
  OR2X2 OR2X2_311 ( .A(_abc_15724_n1654), .B(_abc_15724_n1656_1), .Y(H2_reg_10__FF_INPUT) );
  OR2X2 OR2X2_3110 ( .A(w_mem_inst__abc_21378_n4833), .B(w_mem_inst__abc_21378_n4831), .Y(w_mem_inst__abc_21378_n4834) );
  OR2X2 OR2X2_3111 ( .A(w_mem_inst__abc_21378_n4834), .B(w_mem_inst__abc_21378_n4830), .Y(w_mem_inst__0w_mem_7__31_0__23_) );
  OR2X2 OR2X2_3112 ( .A(w_mem_inst__abc_21378_n4839), .B(w_mem_inst__abc_21378_n4837), .Y(w_mem_inst__abc_21378_n4840) );
  OR2X2 OR2X2_3113 ( .A(w_mem_inst__abc_21378_n4840), .B(w_mem_inst__abc_21378_n4836), .Y(w_mem_inst__0w_mem_7__31_0__24_) );
  OR2X2 OR2X2_3114 ( .A(w_mem_inst__abc_21378_n4845), .B(w_mem_inst__abc_21378_n4843), .Y(w_mem_inst__abc_21378_n4846) );
  OR2X2 OR2X2_3115 ( .A(w_mem_inst__abc_21378_n4846), .B(w_mem_inst__abc_21378_n4842), .Y(w_mem_inst__0w_mem_7__31_0__25_) );
  OR2X2 OR2X2_3116 ( .A(w_mem_inst__abc_21378_n4851), .B(w_mem_inst__abc_21378_n4849), .Y(w_mem_inst__abc_21378_n4852) );
  OR2X2 OR2X2_3117 ( .A(w_mem_inst__abc_21378_n4852), .B(w_mem_inst__abc_21378_n4848), .Y(w_mem_inst__0w_mem_7__31_0__26_) );
  OR2X2 OR2X2_3118 ( .A(w_mem_inst__abc_21378_n4857), .B(w_mem_inst__abc_21378_n4855), .Y(w_mem_inst__abc_21378_n4858) );
  OR2X2 OR2X2_3119 ( .A(w_mem_inst__abc_21378_n4858), .B(w_mem_inst__abc_21378_n4854), .Y(w_mem_inst__0w_mem_7__31_0__27_) );
  OR2X2 OR2X2_312 ( .A(_auto_iopadmap_cc_313_execute_26059_75_), .B(c_reg_11_), .Y(_abc_15724_n1659) );
  OR2X2 OR2X2_3120 ( .A(w_mem_inst__abc_21378_n4863), .B(w_mem_inst__abc_21378_n4861), .Y(w_mem_inst__abc_21378_n4864) );
  OR2X2 OR2X2_3121 ( .A(w_mem_inst__abc_21378_n4864), .B(w_mem_inst__abc_21378_n4860), .Y(w_mem_inst__0w_mem_7__31_0__28_) );
  OR2X2 OR2X2_3122 ( .A(w_mem_inst__abc_21378_n4869), .B(w_mem_inst__abc_21378_n4867), .Y(w_mem_inst__abc_21378_n4870) );
  OR2X2 OR2X2_3123 ( .A(w_mem_inst__abc_21378_n4870), .B(w_mem_inst__abc_21378_n4866), .Y(w_mem_inst__0w_mem_7__31_0__29_) );
  OR2X2 OR2X2_3124 ( .A(w_mem_inst__abc_21378_n4875), .B(w_mem_inst__abc_21378_n4873), .Y(w_mem_inst__abc_21378_n4876) );
  OR2X2 OR2X2_3125 ( .A(w_mem_inst__abc_21378_n4876), .B(w_mem_inst__abc_21378_n4872), .Y(w_mem_inst__0w_mem_7__31_0__30_) );
  OR2X2 OR2X2_3126 ( .A(w_mem_inst__abc_21378_n4881), .B(w_mem_inst__abc_21378_n4879), .Y(w_mem_inst__abc_21378_n4882) );
  OR2X2 OR2X2_3127 ( .A(w_mem_inst__abc_21378_n4882), .B(w_mem_inst__abc_21378_n4878), .Y(w_mem_inst__0w_mem_7__31_0__31_) );
  OR2X2 OR2X2_3128 ( .A(w_mem_inst__abc_21378_n4887), .B(w_mem_inst__abc_21378_n4885), .Y(w_mem_inst__abc_21378_n4888) );
  OR2X2 OR2X2_3129 ( .A(w_mem_inst__abc_21378_n4888), .B(w_mem_inst__abc_21378_n4884), .Y(w_mem_inst__0w_mem_6__31_0__0_) );
  OR2X2 OR2X2_313 ( .A(_abc_15724_n1666), .B(_abc_15724_n1663), .Y(_abc_15724_n1667) );
  OR2X2 OR2X2_3130 ( .A(w_mem_inst__abc_21378_n4893), .B(w_mem_inst__abc_21378_n4891), .Y(w_mem_inst__abc_21378_n4894) );
  OR2X2 OR2X2_3131 ( .A(w_mem_inst__abc_21378_n4894), .B(w_mem_inst__abc_21378_n4890), .Y(w_mem_inst__0w_mem_6__31_0__1_) );
  OR2X2 OR2X2_3132 ( .A(w_mem_inst__abc_21378_n4899), .B(w_mem_inst__abc_21378_n4897), .Y(w_mem_inst__abc_21378_n4900) );
  OR2X2 OR2X2_3133 ( .A(w_mem_inst__abc_21378_n4900), .B(w_mem_inst__abc_21378_n4896), .Y(w_mem_inst__0w_mem_6__31_0__2_) );
  OR2X2 OR2X2_3134 ( .A(w_mem_inst__abc_21378_n4905), .B(w_mem_inst__abc_21378_n4903), .Y(w_mem_inst__abc_21378_n4906) );
  OR2X2 OR2X2_3135 ( .A(w_mem_inst__abc_21378_n4906), .B(w_mem_inst__abc_21378_n4902), .Y(w_mem_inst__0w_mem_6__31_0__3_) );
  OR2X2 OR2X2_3136 ( .A(w_mem_inst__abc_21378_n4911), .B(w_mem_inst__abc_21378_n4909), .Y(w_mem_inst__abc_21378_n4912) );
  OR2X2 OR2X2_3137 ( .A(w_mem_inst__abc_21378_n4912), .B(w_mem_inst__abc_21378_n4908), .Y(w_mem_inst__0w_mem_6__31_0__4_) );
  OR2X2 OR2X2_3138 ( .A(w_mem_inst__abc_21378_n4917), .B(w_mem_inst__abc_21378_n4915), .Y(w_mem_inst__abc_21378_n4918) );
  OR2X2 OR2X2_3139 ( .A(w_mem_inst__abc_21378_n4918), .B(w_mem_inst__abc_21378_n4914), .Y(w_mem_inst__0w_mem_6__31_0__5_) );
  OR2X2 OR2X2_314 ( .A(_abc_15724_n851_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_75_), .Y(_abc_15724_n1669_1) );
  OR2X2 OR2X2_3140 ( .A(w_mem_inst__abc_21378_n4923), .B(w_mem_inst__abc_21378_n4921), .Y(w_mem_inst__abc_21378_n4924) );
  OR2X2 OR2X2_3141 ( .A(w_mem_inst__abc_21378_n4924), .B(w_mem_inst__abc_21378_n4920), .Y(w_mem_inst__0w_mem_6__31_0__6_) );
  OR2X2 OR2X2_3142 ( .A(w_mem_inst__abc_21378_n4929), .B(w_mem_inst__abc_21378_n4927), .Y(w_mem_inst__abc_21378_n4930) );
  OR2X2 OR2X2_3143 ( .A(w_mem_inst__abc_21378_n4930), .B(w_mem_inst__abc_21378_n4926), .Y(w_mem_inst__0w_mem_6__31_0__7_) );
  OR2X2 OR2X2_3144 ( .A(w_mem_inst__abc_21378_n4935), .B(w_mem_inst__abc_21378_n4933), .Y(w_mem_inst__abc_21378_n4936) );
  OR2X2 OR2X2_3145 ( .A(w_mem_inst__abc_21378_n4936), .B(w_mem_inst__abc_21378_n4932), .Y(w_mem_inst__0w_mem_6__31_0__8_) );
  OR2X2 OR2X2_3146 ( .A(w_mem_inst__abc_21378_n4941), .B(w_mem_inst__abc_21378_n4939), .Y(w_mem_inst__abc_21378_n4942) );
  OR2X2 OR2X2_3147 ( .A(w_mem_inst__abc_21378_n4942), .B(w_mem_inst__abc_21378_n4938), .Y(w_mem_inst__0w_mem_6__31_0__9_) );
  OR2X2 OR2X2_3148 ( .A(w_mem_inst__abc_21378_n4947), .B(w_mem_inst__abc_21378_n4945), .Y(w_mem_inst__abc_21378_n4948) );
  OR2X2 OR2X2_3149 ( .A(w_mem_inst__abc_21378_n4948), .B(w_mem_inst__abc_21378_n4944), .Y(w_mem_inst__0w_mem_6__31_0__10_) );
  OR2X2 OR2X2_315 ( .A(_abc_15724_n1668_1), .B(_abc_15724_n1670), .Y(H2_reg_11__FF_INPUT) );
  OR2X2 OR2X2_3150 ( .A(w_mem_inst__abc_21378_n4953), .B(w_mem_inst__abc_21378_n4951), .Y(w_mem_inst__abc_21378_n4954) );
  OR2X2 OR2X2_3151 ( .A(w_mem_inst__abc_21378_n4954), .B(w_mem_inst__abc_21378_n4950), .Y(w_mem_inst__0w_mem_6__31_0__11_) );
  OR2X2 OR2X2_3152 ( .A(w_mem_inst__abc_21378_n4959), .B(w_mem_inst__abc_21378_n4957), .Y(w_mem_inst__abc_21378_n4960) );
  OR2X2 OR2X2_3153 ( .A(w_mem_inst__abc_21378_n4960), .B(w_mem_inst__abc_21378_n4956), .Y(w_mem_inst__0w_mem_6__31_0__12_) );
  OR2X2 OR2X2_3154 ( .A(w_mem_inst__abc_21378_n4965), .B(w_mem_inst__abc_21378_n4963), .Y(w_mem_inst__abc_21378_n4966) );
  OR2X2 OR2X2_3155 ( .A(w_mem_inst__abc_21378_n4966), .B(w_mem_inst__abc_21378_n4962), .Y(w_mem_inst__0w_mem_6__31_0__13_) );
  OR2X2 OR2X2_3156 ( .A(w_mem_inst__abc_21378_n4971), .B(w_mem_inst__abc_21378_n4969), .Y(w_mem_inst__abc_21378_n4972) );
  OR2X2 OR2X2_3157 ( .A(w_mem_inst__abc_21378_n4972), .B(w_mem_inst__abc_21378_n4968), .Y(w_mem_inst__0w_mem_6__31_0__14_) );
  OR2X2 OR2X2_3158 ( .A(w_mem_inst__abc_21378_n4977), .B(w_mem_inst__abc_21378_n4975), .Y(w_mem_inst__abc_21378_n4978) );
  OR2X2 OR2X2_3159 ( .A(w_mem_inst__abc_21378_n4978), .B(w_mem_inst__abc_21378_n4974), .Y(w_mem_inst__0w_mem_6__31_0__15_) );
  OR2X2 OR2X2_316 ( .A(_abc_15724_n1623_1), .B(_abc_15724_n1675_1), .Y(_abc_15724_n1676_1) );
  OR2X2 OR2X2_3160 ( .A(w_mem_inst__abc_21378_n4983), .B(w_mem_inst__abc_21378_n4981), .Y(w_mem_inst__abc_21378_n4984) );
  OR2X2 OR2X2_3161 ( .A(w_mem_inst__abc_21378_n4984), .B(w_mem_inst__abc_21378_n4980), .Y(w_mem_inst__0w_mem_6__31_0__16_) );
  OR2X2 OR2X2_3162 ( .A(w_mem_inst__abc_21378_n4989), .B(w_mem_inst__abc_21378_n4987), .Y(w_mem_inst__abc_21378_n4990) );
  OR2X2 OR2X2_3163 ( .A(w_mem_inst__abc_21378_n4990), .B(w_mem_inst__abc_21378_n4986), .Y(w_mem_inst__0w_mem_6__31_0__17_) );
  OR2X2 OR2X2_3164 ( .A(w_mem_inst__abc_21378_n4995), .B(w_mem_inst__abc_21378_n4993), .Y(w_mem_inst__abc_21378_n4996) );
  OR2X2 OR2X2_3165 ( .A(w_mem_inst__abc_21378_n4996), .B(w_mem_inst__abc_21378_n4992), .Y(w_mem_inst__0w_mem_6__31_0__18_) );
  OR2X2 OR2X2_3166 ( .A(w_mem_inst__abc_21378_n5001), .B(w_mem_inst__abc_21378_n4999), .Y(w_mem_inst__abc_21378_n5002) );
  OR2X2 OR2X2_3167 ( .A(w_mem_inst__abc_21378_n5002), .B(w_mem_inst__abc_21378_n4998), .Y(w_mem_inst__0w_mem_6__31_0__19_) );
  OR2X2 OR2X2_3168 ( .A(w_mem_inst__abc_21378_n5007), .B(w_mem_inst__abc_21378_n5005), .Y(w_mem_inst__abc_21378_n5008) );
  OR2X2 OR2X2_3169 ( .A(w_mem_inst__abc_21378_n5008), .B(w_mem_inst__abc_21378_n5004), .Y(w_mem_inst__0w_mem_6__31_0__20_) );
  OR2X2 OR2X2_317 ( .A(_abc_15724_n1677), .B(_abc_15724_n1632), .Y(_abc_15724_n1678_1) );
  OR2X2 OR2X2_3170 ( .A(w_mem_inst__abc_21378_n5013), .B(w_mem_inst__abc_21378_n5011), .Y(w_mem_inst__abc_21378_n5014) );
  OR2X2 OR2X2_3171 ( .A(w_mem_inst__abc_21378_n5014), .B(w_mem_inst__abc_21378_n5010), .Y(w_mem_inst__0w_mem_6__31_0__21_) );
  OR2X2 OR2X2_3172 ( .A(w_mem_inst__abc_21378_n5019), .B(w_mem_inst__abc_21378_n5017), .Y(w_mem_inst__abc_21378_n5020) );
  OR2X2 OR2X2_3173 ( .A(w_mem_inst__abc_21378_n5020), .B(w_mem_inst__abc_21378_n5016), .Y(w_mem_inst__0w_mem_6__31_0__22_) );
  OR2X2 OR2X2_3174 ( .A(w_mem_inst__abc_21378_n5025), .B(w_mem_inst__abc_21378_n5023), .Y(w_mem_inst__abc_21378_n5026) );
  OR2X2 OR2X2_3175 ( .A(w_mem_inst__abc_21378_n5026), .B(w_mem_inst__abc_21378_n5022), .Y(w_mem_inst__0w_mem_6__31_0__23_) );
  OR2X2 OR2X2_3176 ( .A(w_mem_inst__abc_21378_n5031), .B(w_mem_inst__abc_21378_n5029), .Y(w_mem_inst__abc_21378_n5032) );
  OR2X2 OR2X2_3177 ( .A(w_mem_inst__abc_21378_n5032), .B(w_mem_inst__abc_21378_n5028), .Y(w_mem_inst__0w_mem_6__31_0__24_) );
  OR2X2 OR2X2_3178 ( .A(w_mem_inst__abc_21378_n5037), .B(w_mem_inst__abc_21378_n5035), .Y(w_mem_inst__abc_21378_n5038) );
  OR2X2 OR2X2_3179 ( .A(w_mem_inst__abc_21378_n5038), .B(w_mem_inst__abc_21378_n5034), .Y(w_mem_inst__0w_mem_6__31_0__25_) );
  OR2X2 OR2X2_318 ( .A(_abc_15724_n1680), .B(_abc_15724_n1660), .Y(_abc_15724_n1681_1) );
  OR2X2 OR2X2_3180 ( .A(w_mem_inst__abc_21378_n5043), .B(w_mem_inst__abc_21378_n5041), .Y(w_mem_inst__abc_21378_n5044) );
  OR2X2 OR2X2_3181 ( .A(w_mem_inst__abc_21378_n5044), .B(w_mem_inst__abc_21378_n5040), .Y(w_mem_inst__0w_mem_6__31_0__26_) );
  OR2X2 OR2X2_3182 ( .A(w_mem_inst__abc_21378_n5049), .B(w_mem_inst__abc_21378_n5047), .Y(w_mem_inst__abc_21378_n5050) );
  OR2X2 OR2X2_3183 ( .A(w_mem_inst__abc_21378_n5050), .B(w_mem_inst__abc_21378_n5046), .Y(w_mem_inst__0w_mem_6__31_0__27_) );
  OR2X2 OR2X2_3184 ( .A(w_mem_inst__abc_21378_n5055), .B(w_mem_inst__abc_21378_n5053), .Y(w_mem_inst__abc_21378_n5056) );
  OR2X2 OR2X2_3185 ( .A(w_mem_inst__abc_21378_n5056), .B(w_mem_inst__abc_21378_n5052), .Y(w_mem_inst__0w_mem_6__31_0__28_) );
  OR2X2 OR2X2_3186 ( .A(w_mem_inst__abc_21378_n5061), .B(w_mem_inst__abc_21378_n5059), .Y(w_mem_inst__abc_21378_n5062) );
  OR2X2 OR2X2_3187 ( .A(w_mem_inst__abc_21378_n5062), .B(w_mem_inst__abc_21378_n5058), .Y(w_mem_inst__0w_mem_6__31_0__29_) );
  OR2X2 OR2X2_3188 ( .A(w_mem_inst__abc_21378_n5067), .B(w_mem_inst__abc_21378_n5065), .Y(w_mem_inst__abc_21378_n5068) );
  OR2X2 OR2X2_3189 ( .A(w_mem_inst__abc_21378_n5068), .B(w_mem_inst__abc_21378_n5064), .Y(w_mem_inst__0w_mem_6__31_0__30_) );
  OR2X2 OR2X2_319 ( .A(_abc_15724_n1679), .B(_abc_15724_n1681_1), .Y(_abc_15724_n1682_1) );
  OR2X2 OR2X2_3190 ( .A(w_mem_inst__abc_21378_n5073), .B(w_mem_inst__abc_21378_n5071), .Y(w_mem_inst__abc_21378_n5074) );
  OR2X2 OR2X2_3191 ( .A(w_mem_inst__abc_21378_n5074), .B(w_mem_inst__abc_21378_n5070), .Y(w_mem_inst__0w_mem_6__31_0__31_) );
  OR2X2 OR2X2_3192 ( .A(w_mem_inst__abc_21378_n5079), .B(w_mem_inst__abc_21378_n5077), .Y(w_mem_inst__abc_21378_n5080) );
  OR2X2 OR2X2_3193 ( .A(w_mem_inst__abc_21378_n5080), .B(w_mem_inst__abc_21378_n5076), .Y(w_mem_inst__0w_mem_5__31_0__0_) );
  OR2X2 OR2X2_3194 ( .A(w_mem_inst__abc_21378_n5085), .B(w_mem_inst__abc_21378_n5083), .Y(w_mem_inst__abc_21378_n5086) );
  OR2X2 OR2X2_3195 ( .A(w_mem_inst__abc_21378_n5086), .B(w_mem_inst__abc_21378_n5082), .Y(w_mem_inst__0w_mem_5__31_0__1_) );
  OR2X2 OR2X2_3196 ( .A(w_mem_inst__abc_21378_n5091), .B(w_mem_inst__abc_21378_n5089), .Y(w_mem_inst__abc_21378_n5092) );
  OR2X2 OR2X2_3197 ( .A(w_mem_inst__abc_21378_n5092), .B(w_mem_inst__abc_21378_n5088), .Y(w_mem_inst__0w_mem_5__31_0__2_) );
  OR2X2 OR2X2_3198 ( .A(w_mem_inst__abc_21378_n5097), .B(w_mem_inst__abc_21378_n5095), .Y(w_mem_inst__abc_21378_n5098) );
  OR2X2 OR2X2_3199 ( .A(w_mem_inst__abc_21378_n5098), .B(w_mem_inst__abc_21378_n5094), .Y(w_mem_inst__0w_mem_5__31_0__3_) );
  OR2X2 OR2X2_32 ( .A(_abc_15724_n811), .B(_abc_15724_n784), .Y(_abc_15724_n812_1) );
  OR2X2 OR2X2_320 ( .A(_auto_iopadmap_cc_313_execute_26059_76_), .B(c_reg_12_), .Y(_abc_15724_n1686) );
  OR2X2 OR2X2_3200 ( .A(w_mem_inst__abc_21378_n5103), .B(w_mem_inst__abc_21378_n5101), .Y(w_mem_inst__abc_21378_n5104) );
  OR2X2 OR2X2_3201 ( .A(w_mem_inst__abc_21378_n5104), .B(w_mem_inst__abc_21378_n5100), .Y(w_mem_inst__0w_mem_5__31_0__4_) );
  OR2X2 OR2X2_3202 ( .A(w_mem_inst__abc_21378_n5109), .B(w_mem_inst__abc_21378_n5107), .Y(w_mem_inst__abc_21378_n5110) );
  OR2X2 OR2X2_3203 ( .A(w_mem_inst__abc_21378_n5110), .B(w_mem_inst__abc_21378_n5106), .Y(w_mem_inst__0w_mem_5__31_0__5_) );
  OR2X2 OR2X2_3204 ( .A(w_mem_inst__abc_21378_n5115), .B(w_mem_inst__abc_21378_n5113), .Y(w_mem_inst__abc_21378_n5116) );
  OR2X2 OR2X2_3205 ( .A(w_mem_inst__abc_21378_n5116), .B(w_mem_inst__abc_21378_n5112), .Y(w_mem_inst__0w_mem_5__31_0__6_) );
  OR2X2 OR2X2_3206 ( .A(w_mem_inst__abc_21378_n5121), .B(w_mem_inst__abc_21378_n5119), .Y(w_mem_inst__abc_21378_n5122) );
  OR2X2 OR2X2_3207 ( .A(w_mem_inst__abc_21378_n5122), .B(w_mem_inst__abc_21378_n5118), .Y(w_mem_inst__0w_mem_5__31_0__7_) );
  OR2X2 OR2X2_3208 ( .A(w_mem_inst__abc_21378_n5127), .B(w_mem_inst__abc_21378_n5125), .Y(w_mem_inst__abc_21378_n5128) );
  OR2X2 OR2X2_3209 ( .A(w_mem_inst__abc_21378_n5128), .B(w_mem_inst__abc_21378_n5124), .Y(w_mem_inst__0w_mem_5__31_0__8_) );
  OR2X2 OR2X2_321 ( .A(_abc_15724_n1685), .B(_abc_15724_n1689), .Y(_abc_15724_n1690) );
  OR2X2 OR2X2_3210 ( .A(w_mem_inst__abc_21378_n5133), .B(w_mem_inst__abc_21378_n5131), .Y(w_mem_inst__abc_21378_n5134) );
  OR2X2 OR2X2_3211 ( .A(w_mem_inst__abc_21378_n5134), .B(w_mem_inst__abc_21378_n5130), .Y(w_mem_inst__0w_mem_5__31_0__9_) );
  OR2X2 OR2X2_3212 ( .A(w_mem_inst__abc_21378_n5139), .B(w_mem_inst__abc_21378_n5137), .Y(w_mem_inst__abc_21378_n5140) );
  OR2X2 OR2X2_3213 ( .A(w_mem_inst__abc_21378_n5140), .B(w_mem_inst__abc_21378_n5136), .Y(w_mem_inst__0w_mem_5__31_0__10_) );
  OR2X2 OR2X2_3214 ( .A(w_mem_inst__abc_21378_n5145), .B(w_mem_inst__abc_21378_n5143), .Y(w_mem_inst__abc_21378_n5146) );
  OR2X2 OR2X2_3215 ( .A(w_mem_inst__abc_21378_n5146), .B(w_mem_inst__abc_21378_n5142), .Y(w_mem_inst__0w_mem_5__31_0__11_) );
  OR2X2 OR2X2_3216 ( .A(w_mem_inst__abc_21378_n5151), .B(w_mem_inst__abc_21378_n5149), .Y(w_mem_inst__abc_21378_n5152) );
  OR2X2 OR2X2_3217 ( .A(w_mem_inst__abc_21378_n5152), .B(w_mem_inst__abc_21378_n5148), .Y(w_mem_inst__0w_mem_5__31_0__12_) );
  OR2X2 OR2X2_3218 ( .A(w_mem_inst__abc_21378_n5157), .B(w_mem_inst__abc_21378_n5155), .Y(w_mem_inst__abc_21378_n5158) );
  OR2X2 OR2X2_3219 ( .A(w_mem_inst__abc_21378_n5158), .B(w_mem_inst__abc_21378_n5154), .Y(w_mem_inst__0w_mem_5__31_0__13_) );
  OR2X2 OR2X2_322 ( .A(_abc_15724_n851_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_76_), .Y(_abc_15724_n1695) );
  OR2X2 OR2X2_3220 ( .A(w_mem_inst__abc_21378_n5163), .B(w_mem_inst__abc_21378_n5161), .Y(w_mem_inst__abc_21378_n5164) );
  OR2X2 OR2X2_3221 ( .A(w_mem_inst__abc_21378_n5164), .B(w_mem_inst__abc_21378_n5160), .Y(w_mem_inst__0w_mem_5__31_0__14_) );
  OR2X2 OR2X2_3222 ( .A(w_mem_inst__abc_21378_n5169), .B(w_mem_inst__abc_21378_n5167), .Y(w_mem_inst__abc_21378_n5170) );
  OR2X2 OR2X2_3223 ( .A(w_mem_inst__abc_21378_n5170), .B(w_mem_inst__abc_21378_n5166), .Y(w_mem_inst__0w_mem_5__31_0__15_) );
  OR2X2 OR2X2_3224 ( .A(w_mem_inst__abc_21378_n5175), .B(w_mem_inst__abc_21378_n5173), .Y(w_mem_inst__abc_21378_n5176) );
  OR2X2 OR2X2_3225 ( .A(w_mem_inst__abc_21378_n5176), .B(w_mem_inst__abc_21378_n5172), .Y(w_mem_inst__0w_mem_5__31_0__16_) );
  OR2X2 OR2X2_3226 ( .A(w_mem_inst__abc_21378_n5181), .B(w_mem_inst__abc_21378_n5179), .Y(w_mem_inst__abc_21378_n5182) );
  OR2X2 OR2X2_3227 ( .A(w_mem_inst__abc_21378_n5182), .B(w_mem_inst__abc_21378_n5178), .Y(w_mem_inst__0w_mem_5__31_0__17_) );
  OR2X2 OR2X2_3228 ( .A(w_mem_inst__abc_21378_n5187), .B(w_mem_inst__abc_21378_n5185), .Y(w_mem_inst__abc_21378_n5188) );
  OR2X2 OR2X2_3229 ( .A(w_mem_inst__abc_21378_n5188), .B(w_mem_inst__abc_21378_n5184), .Y(w_mem_inst__0w_mem_5__31_0__18_) );
  OR2X2 OR2X2_323 ( .A(_abc_15724_n1694), .B(_abc_15724_n1696_1), .Y(H2_reg_12__FF_INPUT) );
  OR2X2 OR2X2_3230 ( .A(w_mem_inst__abc_21378_n5193), .B(w_mem_inst__abc_21378_n5191), .Y(w_mem_inst__abc_21378_n5194) );
  OR2X2 OR2X2_3231 ( .A(w_mem_inst__abc_21378_n5194), .B(w_mem_inst__abc_21378_n5190), .Y(w_mem_inst__0w_mem_5__31_0__19_) );
  OR2X2 OR2X2_3232 ( .A(w_mem_inst__abc_21378_n5199), .B(w_mem_inst__abc_21378_n5197), .Y(w_mem_inst__abc_21378_n5200) );
  OR2X2 OR2X2_3233 ( .A(w_mem_inst__abc_21378_n5200), .B(w_mem_inst__abc_21378_n5196), .Y(w_mem_inst__0w_mem_5__31_0__20_) );
  OR2X2 OR2X2_3234 ( .A(w_mem_inst__abc_21378_n5205), .B(w_mem_inst__abc_21378_n5203), .Y(w_mem_inst__abc_21378_n5206) );
  OR2X2 OR2X2_3235 ( .A(w_mem_inst__abc_21378_n5206), .B(w_mem_inst__abc_21378_n5202), .Y(w_mem_inst__0w_mem_5__31_0__21_) );
  OR2X2 OR2X2_3236 ( .A(w_mem_inst__abc_21378_n5211), .B(w_mem_inst__abc_21378_n5209), .Y(w_mem_inst__abc_21378_n5212) );
  OR2X2 OR2X2_3237 ( .A(w_mem_inst__abc_21378_n5212), .B(w_mem_inst__abc_21378_n5208), .Y(w_mem_inst__0w_mem_5__31_0__22_) );
  OR2X2 OR2X2_3238 ( .A(w_mem_inst__abc_21378_n5217), .B(w_mem_inst__abc_21378_n5215), .Y(w_mem_inst__abc_21378_n5218) );
  OR2X2 OR2X2_3239 ( .A(w_mem_inst__abc_21378_n5218), .B(w_mem_inst__abc_21378_n5214), .Y(w_mem_inst__0w_mem_5__31_0__23_) );
  OR2X2 OR2X2_324 ( .A(_auto_iopadmap_cc_313_execute_26059_77_), .B(c_reg_13_), .Y(_abc_15724_n1698) );
  OR2X2 OR2X2_3240 ( .A(w_mem_inst__abc_21378_n5223), .B(w_mem_inst__abc_21378_n5221), .Y(w_mem_inst__abc_21378_n5224) );
  OR2X2 OR2X2_3241 ( .A(w_mem_inst__abc_21378_n5224), .B(w_mem_inst__abc_21378_n5220), .Y(w_mem_inst__0w_mem_5__31_0__24_) );
  OR2X2 OR2X2_3242 ( .A(w_mem_inst__abc_21378_n5229), .B(w_mem_inst__abc_21378_n5227), .Y(w_mem_inst__abc_21378_n5230) );
  OR2X2 OR2X2_3243 ( .A(w_mem_inst__abc_21378_n5230), .B(w_mem_inst__abc_21378_n5226), .Y(w_mem_inst__0w_mem_5__31_0__25_) );
  OR2X2 OR2X2_3244 ( .A(w_mem_inst__abc_21378_n5235), .B(w_mem_inst__abc_21378_n5233), .Y(w_mem_inst__abc_21378_n5236) );
  OR2X2 OR2X2_3245 ( .A(w_mem_inst__abc_21378_n5236), .B(w_mem_inst__abc_21378_n5232), .Y(w_mem_inst__0w_mem_5__31_0__26_) );
  OR2X2 OR2X2_3246 ( .A(w_mem_inst__abc_21378_n5241), .B(w_mem_inst__abc_21378_n5239), .Y(w_mem_inst__abc_21378_n5242) );
  OR2X2 OR2X2_3247 ( .A(w_mem_inst__abc_21378_n5242), .B(w_mem_inst__abc_21378_n5238), .Y(w_mem_inst__0w_mem_5__31_0__27_) );
  OR2X2 OR2X2_3248 ( .A(w_mem_inst__abc_21378_n5247), .B(w_mem_inst__abc_21378_n5245), .Y(w_mem_inst__abc_21378_n5248) );
  OR2X2 OR2X2_3249 ( .A(w_mem_inst__abc_21378_n5248), .B(w_mem_inst__abc_21378_n5244), .Y(w_mem_inst__0w_mem_5__31_0__28_) );
  OR2X2 OR2X2_325 ( .A(_abc_15724_n1703), .B(_abc_15724_n1701), .Y(_abc_15724_n1704_1) );
  OR2X2 OR2X2_3250 ( .A(w_mem_inst__abc_21378_n5253), .B(w_mem_inst__abc_21378_n5251), .Y(w_mem_inst__abc_21378_n5254) );
  OR2X2 OR2X2_3251 ( .A(w_mem_inst__abc_21378_n5254), .B(w_mem_inst__abc_21378_n5250), .Y(w_mem_inst__0w_mem_5__31_0__29_) );
  OR2X2 OR2X2_3252 ( .A(w_mem_inst__abc_21378_n5259), .B(w_mem_inst__abc_21378_n5257), .Y(w_mem_inst__abc_21378_n5260) );
  OR2X2 OR2X2_3253 ( .A(w_mem_inst__abc_21378_n5260), .B(w_mem_inst__abc_21378_n5256), .Y(w_mem_inst__0w_mem_5__31_0__30_) );
  OR2X2 OR2X2_3254 ( .A(w_mem_inst__abc_21378_n5265), .B(w_mem_inst__abc_21378_n5263), .Y(w_mem_inst__abc_21378_n5266) );
  OR2X2 OR2X2_3255 ( .A(w_mem_inst__abc_21378_n5266), .B(w_mem_inst__abc_21378_n5262), .Y(w_mem_inst__0w_mem_5__31_0__31_) );
  OR2X2 OR2X2_3256 ( .A(w_mem_inst__abc_21378_n5271), .B(w_mem_inst__abc_21378_n5269), .Y(w_mem_inst__abc_21378_n5272) );
  OR2X2 OR2X2_3257 ( .A(w_mem_inst__abc_21378_n5272), .B(w_mem_inst__abc_21378_n5268), .Y(w_mem_inst__0w_mem_4__31_0__0_) );
  OR2X2 OR2X2_3258 ( .A(w_mem_inst__abc_21378_n5277), .B(w_mem_inst__abc_21378_n5275), .Y(w_mem_inst__abc_21378_n5278) );
  OR2X2 OR2X2_3259 ( .A(w_mem_inst__abc_21378_n5278), .B(w_mem_inst__abc_21378_n5274), .Y(w_mem_inst__0w_mem_4__31_0__1_) );
  OR2X2 OR2X2_326 ( .A(_abc_15724_n1708), .B(_abc_15724_n1709_1), .Y(H2_reg_13__FF_INPUT) );
  OR2X2 OR2X2_3260 ( .A(w_mem_inst__abc_21378_n5283), .B(w_mem_inst__abc_21378_n5281), .Y(w_mem_inst__abc_21378_n5284) );
  OR2X2 OR2X2_3261 ( .A(w_mem_inst__abc_21378_n5284), .B(w_mem_inst__abc_21378_n5280), .Y(w_mem_inst__0w_mem_4__31_0__2_) );
  OR2X2 OR2X2_3262 ( .A(w_mem_inst__abc_21378_n5289), .B(w_mem_inst__abc_21378_n5287), .Y(w_mem_inst__abc_21378_n5290) );
  OR2X2 OR2X2_3263 ( .A(w_mem_inst__abc_21378_n5290), .B(w_mem_inst__abc_21378_n5286), .Y(w_mem_inst__0w_mem_4__31_0__3_) );
  OR2X2 OR2X2_3264 ( .A(w_mem_inst__abc_21378_n5295), .B(w_mem_inst__abc_21378_n5293), .Y(w_mem_inst__abc_21378_n5296) );
  OR2X2 OR2X2_3265 ( .A(w_mem_inst__abc_21378_n5296), .B(w_mem_inst__abc_21378_n5292), .Y(w_mem_inst__0w_mem_4__31_0__4_) );
  OR2X2 OR2X2_3266 ( .A(w_mem_inst__abc_21378_n5301), .B(w_mem_inst__abc_21378_n5299), .Y(w_mem_inst__abc_21378_n5302) );
  OR2X2 OR2X2_3267 ( .A(w_mem_inst__abc_21378_n5302), .B(w_mem_inst__abc_21378_n5298), .Y(w_mem_inst__0w_mem_4__31_0__5_) );
  OR2X2 OR2X2_3268 ( .A(w_mem_inst__abc_21378_n5307), .B(w_mem_inst__abc_21378_n5305), .Y(w_mem_inst__abc_21378_n5308) );
  OR2X2 OR2X2_3269 ( .A(w_mem_inst__abc_21378_n5308), .B(w_mem_inst__abc_21378_n5304), .Y(w_mem_inst__0w_mem_4__31_0__6_) );
  OR2X2 OR2X2_327 ( .A(_auto_iopadmap_cc_313_execute_26059_78_), .B(c_reg_14_), .Y(_abc_15724_n1713) );
  OR2X2 OR2X2_3270 ( .A(w_mem_inst__abc_21378_n5313), .B(w_mem_inst__abc_21378_n5311), .Y(w_mem_inst__abc_21378_n5314) );
  OR2X2 OR2X2_3271 ( .A(w_mem_inst__abc_21378_n5314), .B(w_mem_inst__abc_21378_n5310), .Y(w_mem_inst__0w_mem_4__31_0__7_) );
  OR2X2 OR2X2_3272 ( .A(w_mem_inst__abc_21378_n5319), .B(w_mem_inst__abc_21378_n5317), .Y(w_mem_inst__abc_21378_n5320) );
  OR2X2 OR2X2_3273 ( .A(w_mem_inst__abc_21378_n5320), .B(w_mem_inst__abc_21378_n5316), .Y(w_mem_inst__0w_mem_4__31_0__8_) );
  OR2X2 OR2X2_3274 ( .A(w_mem_inst__abc_21378_n5325), .B(w_mem_inst__abc_21378_n5323), .Y(w_mem_inst__abc_21378_n5326) );
  OR2X2 OR2X2_3275 ( .A(w_mem_inst__abc_21378_n5326), .B(w_mem_inst__abc_21378_n5322), .Y(w_mem_inst__0w_mem_4__31_0__9_) );
  OR2X2 OR2X2_3276 ( .A(w_mem_inst__abc_21378_n5331), .B(w_mem_inst__abc_21378_n5329), .Y(w_mem_inst__abc_21378_n5332) );
  OR2X2 OR2X2_3277 ( .A(w_mem_inst__abc_21378_n5332), .B(w_mem_inst__abc_21378_n5328), .Y(w_mem_inst__0w_mem_4__31_0__10_) );
  OR2X2 OR2X2_3278 ( .A(w_mem_inst__abc_21378_n5337), .B(w_mem_inst__abc_21378_n5335), .Y(w_mem_inst__abc_21378_n5338) );
  OR2X2 OR2X2_3279 ( .A(w_mem_inst__abc_21378_n5338), .B(w_mem_inst__abc_21378_n5334), .Y(w_mem_inst__0w_mem_4__31_0__11_) );
  OR2X2 OR2X2_328 ( .A(_abc_15724_n1712), .B(_abc_15724_n1716), .Y(_abc_15724_n1717) );
  OR2X2 OR2X2_3280 ( .A(w_mem_inst__abc_21378_n5343), .B(w_mem_inst__abc_21378_n5341), .Y(w_mem_inst__abc_21378_n5344) );
  OR2X2 OR2X2_3281 ( .A(w_mem_inst__abc_21378_n5344), .B(w_mem_inst__abc_21378_n5340), .Y(w_mem_inst__0w_mem_4__31_0__12_) );
  OR2X2 OR2X2_3282 ( .A(w_mem_inst__abc_21378_n5349), .B(w_mem_inst__abc_21378_n5347), .Y(w_mem_inst__abc_21378_n5350) );
  OR2X2 OR2X2_3283 ( .A(w_mem_inst__abc_21378_n5350), .B(w_mem_inst__abc_21378_n5346), .Y(w_mem_inst__0w_mem_4__31_0__13_) );
  OR2X2 OR2X2_3284 ( .A(w_mem_inst__abc_21378_n5355), .B(w_mem_inst__abc_21378_n5353), .Y(w_mem_inst__abc_21378_n5356) );
  OR2X2 OR2X2_3285 ( .A(w_mem_inst__abc_21378_n5356), .B(w_mem_inst__abc_21378_n5352), .Y(w_mem_inst__0w_mem_4__31_0__14_) );
  OR2X2 OR2X2_3286 ( .A(w_mem_inst__abc_21378_n5361), .B(w_mem_inst__abc_21378_n5359), .Y(w_mem_inst__abc_21378_n5362) );
  OR2X2 OR2X2_3287 ( .A(w_mem_inst__abc_21378_n5362), .B(w_mem_inst__abc_21378_n5358), .Y(w_mem_inst__0w_mem_4__31_0__15_) );
  OR2X2 OR2X2_3288 ( .A(w_mem_inst__abc_21378_n5367), .B(w_mem_inst__abc_21378_n5365), .Y(w_mem_inst__abc_21378_n5368) );
  OR2X2 OR2X2_3289 ( .A(w_mem_inst__abc_21378_n5368), .B(w_mem_inst__abc_21378_n5364), .Y(w_mem_inst__0w_mem_4__31_0__16_) );
  OR2X2 OR2X2_329 ( .A(_abc_15724_n851_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_78_), .Y(_abc_15724_n1722) );
  OR2X2 OR2X2_3290 ( .A(w_mem_inst__abc_21378_n5373), .B(w_mem_inst__abc_21378_n5371), .Y(w_mem_inst__abc_21378_n5374) );
  OR2X2 OR2X2_3291 ( .A(w_mem_inst__abc_21378_n5374), .B(w_mem_inst__abc_21378_n5370), .Y(w_mem_inst__0w_mem_4__31_0__17_) );
  OR2X2 OR2X2_3292 ( .A(w_mem_inst__abc_21378_n5379), .B(w_mem_inst__abc_21378_n5377), .Y(w_mem_inst__abc_21378_n5380) );
  OR2X2 OR2X2_3293 ( .A(w_mem_inst__abc_21378_n5380), .B(w_mem_inst__abc_21378_n5376), .Y(w_mem_inst__0w_mem_4__31_0__18_) );
  OR2X2 OR2X2_3294 ( .A(w_mem_inst__abc_21378_n5385), .B(w_mem_inst__abc_21378_n5383), .Y(w_mem_inst__abc_21378_n5386) );
  OR2X2 OR2X2_3295 ( .A(w_mem_inst__abc_21378_n5386), .B(w_mem_inst__abc_21378_n5382), .Y(w_mem_inst__0w_mem_4__31_0__19_) );
  OR2X2 OR2X2_3296 ( .A(w_mem_inst__abc_21378_n5391), .B(w_mem_inst__abc_21378_n5389), .Y(w_mem_inst__abc_21378_n5392) );
  OR2X2 OR2X2_3297 ( .A(w_mem_inst__abc_21378_n5392), .B(w_mem_inst__abc_21378_n5388), .Y(w_mem_inst__0w_mem_4__31_0__20_) );
  OR2X2 OR2X2_3298 ( .A(w_mem_inst__abc_21378_n5397), .B(w_mem_inst__abc_21378_n5395), .Y(w_mem_inst__abc_21378_n5398) );
  OR2X2 OR2X2_3299 ( .A(w_mem_inst__abc_21378_n5398), .B(w_mem_inst__abc_21378_n5394), .Y(w_mem_inst__0w_mem_4__31_0__21_) );
  OR2X2 OR2X2_33 ( .A(_abc_15724_n813_1), .B(_abc_15724_n777), .Y(_abc_15724_n814) );
  OR2X2 OR2X2_330 ( .A(_abc_15724_n1721), .B(_abc_15724_n1723), .Y(H2_reg_14__FF_INPUT) );
  OR2X2 OR2X2_3300 ( .A(w_mem_inst__abc_21378_n5403), .B(w_mem_inst__abc_21378_n5401), .Y(w_mem_inst__abc_21378_n5404) );
  OR2X2 OR2X2_3301 ( .A(w_mem_inst__abc_21378_n5404), .B(w_mem_inst__abc_21378_n5400), .Y(w_mem_inst__0w_mem_4__31_0__22_) );
  OR2X2 OR2X2_3302 ( .A(w_mem_inst__abc_21378_n5409), .B(w_mem_inst__abc_21378_n5407), .Y(w_mem_inst__abc_21378_n5410) );
  OR2X2 OR2X2_3303 ( .A(w_mem_inst__abc_21378_n5410), .B(w_mem_inst__abc_21378_n5406), .Y(w_mem_inst__0w_mem_4__31_0__23_) );
  OR2X2 OR2X2_3304 ( .A(w_mem_inst__abc_21378_n5415), .B(w_mem_inst__abc_21378_n5413), .Y(w_mem_inst__abc_21378_n5416) );
  OR2X2 OR2X2_3305 ( .A(w_mem_inst__abc_21378_n5416), .B(w_mem_inst__abc_21378_n5412), .Y(w_mem_inst__0w_mem_4__31_0__24_) );
  OR2X2 OR2X2_3306 ( .A(w_mem_inst__abc_21378_n5421), .B(w_mem_inst__abc_21378_n5419), .Y(w_mem_inst__abc_21378_n5422) );
  OR2X2 OR2X2_3307 ( .A(w_mem_inst__abc_21378_n5422), .B(w_mem_inst__abc_21378_n5418), .Y(w_mem_inst__0w_mem_4__31_0__25_) );
  OR2X2 OR2X2_3308 ( .A(w_mem_inst__abc_21378_n5427), .B(w_mem_inst__abc_21378_n5425), .Y(w_mem_inst__abc_21378_n5428) );
  OR2X2 OR2X2_3309 ( .A(w_mem_inst__abc_21378_n5428), .B(w_mem_inst__abc_21378_n5424), .Y(w_mem_inst__0w_mem_4__31_0__26_) );
  OR2X2 OR2X2_331 ( .A(_auto_iopadmap_cc_313_execute_26059_79_), .B(c_reg_15_), .Y(_abc_15724_n1727) );
  OR2X2 OR2X2_3310 ( .A(w_mem_inst__abc_21378_n5433), .B(w_mem_inst__abc_21378_n5431), .Y(w_mem_inst__abc_21378_n5434) );
  OR2X2 OR2X2_3311 ( .A(w_mem_inst__abc_21378_n5434), .B(w_mem_inst__abc_21378_n5430), .Y(w_mem_inst__0w_mem_4__31_0__27_) );
  OR2X2 OR2X2_3312 ( .A(w_mem_inst__abc_21378_n5439), .B(w_mem_inst__abc_21378_n5437), .Y(w_mem_inst__abc_21378_n5440) );
  OR2X2 OR2X2_3313 ( .A(w_mem_inst__abc_21378_n5440), .B(w_mem_inst__abc_21378_n5436), .Y(w_mem_inst__0w_mem_4__31_0__28_) );
  OR2X2 OR2X2_3314 ( .A(w_mem_inst__abc_21378_n5445), .B(w_mem_inst__abc_21378_n5443), .Y(w_mem_inst__abc_21378_n5446) );
  OR2X2 OR2X2_3315 ( .A(w_mem_inst__abc_21378_n5446), .B(w_mem_inst__abc_21378_n5442), .Y(w_mem_inst__0w_mem_4__31_0__29_) );
  OR2X2 OR2X2_3316 ( .A(w_mem_inst__abc_21378_n5451), .B(w_mem_inst__abc_21378_n5449), .Y(w_mem_inst__abc_21378_n5452) );
  OR2X2 OR2X2_3317 ( .A(w_mem_inst__abc_21378_n5452), .B(w_mem_inst__abc_21378_n5448), .Y(w_mem_inst__0w_mem_4__31_0__30_) );
  OR2X2 OR2X2_3318 ( .A(w_mem_inst__abc_21378_n5457), .B(w_mem_inst__abc_21378_n5455), .Y(w_mem_inst__abc_21378_n5458) );
  OR2X2 OR2X2_3319 ( .A(w_mem_inst__abc_21378_n5458), .B(w_mem_inst__abc_21378_n5454), .Y(w_mem_inst__0w_mem_4__31_0__31_) );
  OR2X2 OR2X2_332 ( .A(_abc_15724_n1726), .B(_abc_15724_n1730), .Y(_abc_15724_n1731) );
  OR2X2 OR2X2_3320 ( .A(w_mem_inst__abc_21378_n5463), .B(w_mem_inst__abc_21378_n5461), .Y(w_mem_inst__abc_21378_n5464) );
  OR2X2 OR2X2_3321 ( .A(w_mem_inst__abc_21378_n5464), .B(w_mem_inst__abc_21378_n5460), .Y(w_mem_inst__0w_mem_3__31_0__0_) );
  OR2X2 OR2X2_3322 ( .A(w_mem_inst__abc_21378_n5469), .B(w_mem_inst__abc_21378_n5467), .Y(w_mem_inst__abc_21378_n5470) );
  OR2X2 OR2X2_3323 ( .A(w_mem_inst__abc_21378_n5470), .B(w_mem_inst__abc_21378_n5466), .Y(w_mem_inst__0w_mem_3__31_0__1_) );
  OR2X2 OR2X2_3324 ( .A(w_mem_inst__abc_21378_n5475), .B(w_mem_inst__abc_21378_n5473), .Y(w_mem_inst__abc_21378_n5476) );
  OR2X2 OR2X2_3325 ( .A(w_mem_inst__abc_21378_n5476), .B(w_mem_inst__abc_21378_n5472), .Y(w_mem_inst__0w_mem_3__31_0__2_) );
  OR2X2 OR2X2_3326 ( .A(w_mem_inst__abc_21378_n5481), .B(w_mem_inst__abc_21378_n5479), .Y(w_mem_inst__abc_21378_n5482) );
  OR2X2 OR2X2_3327 ( .A(w_mem_inst__abc_21378_n5482), .B(w_mem_inst__abc_21378_n5478), .Y(w_mem_inst__0w_mem_3__31_0__3_) );
  OR2X2 OR2X2_3328 ( .A(w_mem_inst__abc_21378_n5487), .B(w_mem_inst__abc_21378_n5485), .Y(w_mem_inst__abc_21378_n5488) );
  OR2X2 OR2X2_3329 ( .A(w_mem_inst__abc_21378_n5488), .B(w_mem_inst__abc_21378_n5484), .Y(w_mem_inst__0w_mem_3__31_0__4_) );
  OR2X2 OR2X2_333 ( .A(_abc_15724_n1725), .B(_abc_15724_n1732_1), .Y(_abc_15724_n1733) );
  OR2X2 OR2X2_3330 ( .A(w_mem_inst__abc_21378_n5493), .B(w_mem_inst__abc_21378_n5491), .Y(w_mem_inst__abc_21378_n5494) );
  OR2X2 OR2X2_3331 ( .A(w_mem_inst__abc_21378_n5494), .B(w_mem_inst__abc_21378_n5490), .Y(w_mem_inst__0w_mem_3__31_0__5_) );
  OR2X2 OR2X2_3332 ( .A(w_mem_inst__abc_21378_n5499), .B(w_mem_inst__abc_21378_n5497), .Y(w_mem_inst__abc_21378_n5500) );
  OR2X2 OR2X2_3333 ( .A(w_mem_inst__abc_21378_n5500), .B(w_mem_inst__abc_21378_n5496), .Y(w_mem_inst__0w_mem_3__31_0__6_) );
  OR2X2 OR2X2_3334 ( .A(w_mem_inst__abc_21378_n5505), .B(w_mem_inst__abc_21378_n5503), .Y(w_mem_inst__abc_21378_n5506) );
  OR2X2 OR2X2_3335 ( .A(w_mem_inst__abc_21378_n5506), .B(w_mem_inst__abc_21378_n5502), .Y(w_mem_inst__0w_mem_3__31_0__7_) );
  OR2X2 OR2X2_3336 ( .A(w_mem_inst__abc_21378_n5511), .B(w_mem_inst__abc_21378_n5509), .Y(w_mem_inst__abc_21378_n5512) );
  OR2X2 OR2X2_3337 ( .A(w_mem_inst__abc_21378_n5512), .B(w_mem_inst__abc_21378_n5508), .Y(w_mem_inst__0w_mem_3__31_0__8_) );
  OR2X2 OR2X2_3338 ( .A(w_mem_inst__abc_21378_n5517), .B(w_mem_inst__abc_21378_n5515), .Y(w_mem_inst__abc_21378_n5518) );
  OR2X2 OR2X2_3339 ( .A(w_mem_inst__abc_21378_n5518), .B(w_mem_inst__abc_21378_n5514), .Y(w_mem_inst__0w_mem_3__31_0__9_) );
  OR2X2 OR2X2_334 ( .A(_abc_15724_n851_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_79_), .Y(_abc_15724_n1736) );
  OR2X2 OR2X2_3340 ( .A(w_mem_inst__abc_21378_n5523), .B(w_mem_inst__abc_21378_n5521), .Y(w_mem_inst__abc_21378_n5524) );
  OR2X2 OR2X2_3341 ( .A(w_mem_inst__abc_21378_n5524), .B(w_mem_inst__abc_21378_n5520), .Y(w_mem_inst__0w_mem_3__31_0__10_) );
  OR2X2 OR2X2_3342 ( .A(w_mem_inst__abc_21378_n5529), .B(w_mem_inst__abc_21378_n5527), .Y(w_mem_inst__abc_21378_n5530) );
  OR2X2 OR2X2_3343 ( .A(w_mem_inst__abc_21378_n5530), .B(w_mem_inst__abc_21378_n5526), .Y(w_mem_inst__0w_mem_3__31_0__11_) );
  OR2X2 OR2X2_3344 ( .A(w_mem_inst__abc_21378_n5535), .B(w_mem_inst__abc_21378_n5533), .Y(w_mem_inst__abc_21378_n5536) );
  OR2X2 OR2X2_3345 ( .A(w_mem_inst__abc_21378_n5536), .B(w_mem_inst__abc_21378_n5532), .Y(w_mem_inst__0w_mem_3__31_0__12_) );
  OR2X2 OR2X2_3346 ( .A(w_mem_inst__abc_21378_n5541), .B(w_mem_inst__abc_21378_n5539), .Y(w_mem_inst__abc_21378_n5542) );
  OR2X2 OR2X2_3347 ( .A(w_mem_inst__abc_21378_n5542), .B(w_mem_inst__abc_21378_n5538), .Y(w_mem_inst__0w_mem_3__31_0__13_) );
  OR2X2 OR2X2_3348 ( .A(w_mem_inst__abc_21378_n5547), .B(w_mem_inst__abc_21378_n5545), .Y(w_mem_inst__abc_21378_n5548) );
  OR2X2 OR2X2_3349 ( .A(w_mem_inst__abc_21378_n5548), .B(w_mem_inst__abc_21378_n5544), .Y(w_mem_inst__0w_mem_3__31_0__14_) );
  OR2X2 OR2X2_335 ( .A(_abc_15724_n1735), .B(_abc_15724_n1737_1), .Y(H2_reg_15__FF_INPUT) );
  OR2X2 OR2X2_3350 ( .A(w_mem_inst__abc_21378_n5553), .B(w_mem_inst__abc_21378_n5551), .Y(w_mem_inst__abc_21378_n5554) );
  OR2X2 OR2X2_3351 ( .A(w_mem_inst__abc_21378_n5554), .B(w_mem_inst__abc_21378_n5550), .Y(w_mem_inst__0w_mem_3__31_0__15_) );
  OR2X2 OR2X2_3352 ( .A(w_mem_inst__abc_21378_n5559), .B(w_mem_inst__abc_21378_n5557), .Y(w_mem_inst__abc_21378_n5560) );
  OR2X2 OR2X2_3353 ( .A(w_mem_inst__abc_21378_n5560), .B(w_mem_inst__abc_21378_n5556), .Y(w_mem_inst__0w_mem_3__31_0__16_) );
  OR2X2 OR2X2_3354 ( .A(w_mem_inst__abc_21378_n5565), .B(w_mem_inst__abc_21378_n5563), .Y(w_mem_inst__abc_21378_n5566) );
  OR2X2 OR2X2_3355 ( .A(w_mem_inst__abc_21378_n5566), .B(w_mem_inst__abc_21378_n5562), .Y(w_mem_inst__0w_mem_3__31_0__17_) );
  OR2X2 OR2X2_3356 ( .A(w_mem_inst__abc_21378_n5571), .B(w_mem_inst__abc_21378_n5569), .Y(w_mem_inst__abc_21378_n5572) );
  OR2X2 OR2X2_3357 ( .A(w_mem_inst__abc_21378_n5572), .B(w_mem_inst__abc_21378_n5568), .Y(w_mem_inst__0w_mem_3__31_0__18_) );
  OR2X2 OR2X2_3358 ( .A(w_mem_inst__abc_21378_n5577), .B(w_mem_inst__abc_21378_n5575), .Y(w_mem_inst__abc_21378_n5578) );
  OR2X2 OR2X2_3359 ( .A(w_mem_inst__abc_21378_n5578), .B(w_mem_inst__abc_21378_n5574), .Y(w_mem_inst__0w_mem_3__31_0__19_) );
  OR2X2 OR2X2_336 ( .A(_abc_15724_n1740), .B(_abc_15724_n1699), .Y(_abc_15724_n1741_1) );
  OR2X2 OR2X2_3360 ( .A(w_mem_inst__abc_21378_n5583), .B(w_mem_inst__abc_21378_n5581), .Y(w_mem_inst__abc_21378_n5584) );
  OR2X2 OR2X2_3361 ( .A(w_mem_inst__abc_21378_n5584), .B(w_mem_inst__abc_21378_n5580), .Y(w_mem_inst__0w_mem_3__31_0__20_) );
  OR2X2 OR2X2_3362 ( .A(w_mem_inst__abc_21378_n5589), .B(w_mem_inst__abc_21378_n5587), .Y(w_mem_inst__abc_21378_n5590) );
  OR2X2 OR2X2_3363 ( .A(w_mem_inst__abc_21378_n5590), .B(w_mem_inst__abc_21378_n5586), .Y(w_mem_inst__0w_mem_3__31_0__21_) );
  OR2X2 OR2X2_3364 ( .A(w_mem_inst__abc_21378_n5595), .B(w_mem_inst__abc_21378_n5593), .Y(w_mem_inst__abc_21378_n5596) );
  OR2X2 OR2X2_3365 ( .A(w_mem_inst__abc_21378_n5596), .B(w_mem_inst__abc_21378_n5592), .Y(w_mem_inst__0w_mem_3__31_0__22_) );
  OR2X2 OR2X2_3366 ( .A(w_mem_inst__abc_21378_n5601), .B(w_mem_inst__abc_21378_n5599), .Y(w_mem_inst__abc_21378_n5602) );
  OR2X2 OR2X2_3367 ( .A(w_mem_inst__abc_21378_n5602), .B(w_mem_inst__abc_21378_n5598), .Y(w_mem_inst__0w_mem_3__31_0__23_) );
  OR2X2 OR2X2_3368 ( .A(w_mem_inst__abc_21378_n5607), .B(w_mem_inst__abc_21378_n5605), .Y(w_mem_inst__abc_21378_n5608) );
  OR2X2 OR2X2_3369 ( .A(w_mem_inst__abc_21378_n5608), .B(w_mem_inst__abc_21378_n5604), .Y(w_mem_inst__0w_mem_3__31_0__24_) );
  OR2X2 OR2X2_337 ( .A(_abc_15724_n1744), .B(_abc_15724_n1728_1), .Y(_abc_15724_n1745_1) );
  OR2X2 OR2X2_3370 ( .A(w_mem_inst__abc_21378_n5613), .B(w_mem_inst__abc_21378_n5611), .Y(w_mem_inst__abc_21378_n5614) );
  OR2X2 OR2X2_3371 ( .A(w_mem_inst__abc_21378_n5614), .B(w_mem_inst__abc_21378_n5610), .Y(w_mem_inst__0w_mem_3__31_0__25_) );
  OR2X2 OR2X2_3372 ( .A(w_mem_inst__abc_21378_n5619), .B(w_mem_inst__abc_21378_n5617), .Y(w_mem_inst__abc_21378_n5620) );
  OR2X2 OR2X2_3373 ( .A(w_mem_inst__abc_21378_n5620), .B(w_mem_inst__abc_21378_n5616), .Y(w_mem_inst__0w_mem_3__31_0__26_) );
  OR2X2 OR2X2_3374 ( .A(w_mem_inst__abc_21378_n5625), .B(w_mem_inst__abc_21378_n5623), .Y(w_mem_inst__abc_21378_n5626) );
  OR2X2 OR2X2_3375 ( .A(w_mem_inst__abc_21378_n5626), .B(w_mem_inst__abc_21378_n5622), .Y(w_mem_inst__0w_mem_3__31_0__27_) );
  OR2X2 OR2X2_3376 ( .A(w_mem_inst__abc_21378_n5631), .B(w_mem_inst__abc_21378_n5629), .Y(w_mem_inst__abc_21378_n5632) );
  OR2X2 OR2X2_3377 ( .A(w_mem_inst__abc_21378_n5632), .B(w_mem_inst__abc_21378_n5628), .Y(w_mem_inst__0w_mem_3__31_0__28_) );
  OR2X2 OR2X2_3378 ( .A(w_mem_inst__abc_21378_n5637), .B(w_mem_inst__abc_21378_n5635), .Y(w_mem_inst__abc_21378_n5638) );
  OR2X2 OR2X2_3379 ( .A(w_mem_inst__abc_21378_n5638), .B(w_mem_inst__abc_21378_n5634), .Y(w_mem_inst__0w_mem_3__31_0__29_) );
  OR2X2 OR2X2_338 ( .A(_abc_15724_n1743), .B(_abc_15724_n1745_1), .Y(_abc_15724_n1746) );
  OR2X2 OR2X2_3380 ( .A(w_mem_inst__abc_21378_n5643), .B(w_mem_inst__abc_21378_n5641), .Y(w_mem_inst__abc_21378_n5644) );
  OR2X2 OR2X2_3381 ( .A(w_mem_inst__abc_21378_n5644), .B(w_mem_inst__abc_21378_n5640), .Y(w_mem_inst__0w_mem_3__31_0__30_) );
  OR2X2 OR2X2_3382 ( .A(w_mem_inst__abc_21378_n5649), .B(w_mem_inst__abc_21378_n5647), .Y(w_mem_inst__abc_21378_n5650) );
  OR2X2 OR2X2_3383 ( .A(w_mem_inst__abc_21378_n5650), .B(w_mem_inst__abc_21378_n5646), .Y(w_mem_inst__0w_mem_3__31_0__31_) );
  OR2X2 OR2X2_3384 ( .A(w_mem_inst__abc_21378_n5655), .B(w_mem_inst__abc_21378_n5653), .Y(w_mem_inst__abc_21378_n5656) );
  OR2X2 OR2X2_3385 ( .A(w_mem_inst__abc_21378_n5656), .B(w_mem_inst__abc_21378_n5652), .Y(w_mem_inst__0w_mem_2__31_0__0_) );
  OR2X2 OR2X2_3386 ( .A(w_mem_inst__abc_21378_n5661), .B(w_mem_inst__abc_21378_n5659), .Y(w_mem_inst__abc_21378_n5662) );
  OR2X2 OR2X2_3387 ( .A(w_mem_inst__abc_21378_n5662), .B(w_mem_inst__abc_21378_n5658), .Y(w_mem_inst__0w_mem_2__31_0__1_) );
  OR2X2 OR2X2_3388 ( .A(w_mem_inst__abc_21378_n5667), .B(w_mem_inst__abc_21378_n5665), .Y(w_mem_inst__abc_21378_n5668) );
  OR2X2 OR2X2_3389 ( .A(w_mem_inst__abc_21378_n5668), .B(w_mem_inst__abc_21378_n5664), .Y(w_mem_inst__0w_mem_2__31_0__2_) );
  OR2X2 OR2X2_339 ( .A(_abc_15724_n1684), .B(_abc_15724_n1750_1), .Y(_abc_15724_n1751) );
  OR2X2 OR2X2_3390 ( .A(w_mem_inst__abc_21378_n5673), .B(w_mem_inst__abc_21378_n5671), .Y(w_mem_inst__abc_21378_n5674) );
  OR2X2 OR2X2_3391 ( .A(w_mem_inst__abc_21378_n5674), .B(w_mem_inst__abc_21378_n5670), .Y(w_mem_inst__0w_mem_2__31_0__3_) );
  OR2X2 OR2X2_3392 ( .A(w_mem_inst__abc_21378_n5679), .B(w_mem_inst__abc_21378_n5677), .Y(w_mem_inst__abc_21378_n5680) );
  OR2X2 OR2X2_3393 ( .A(w_mem_inst__abc_21378_n5680), .B(w_mem_inst__abc_21378_n5676), .Y(w_mem_inst__0w_mem_2__31_0__4_) );
  OR2X2 OR2X2_3394 ( .A(w_mem_inst__abc_21378_n5685), .B(w_mem_inst__abc_21378_n5683), .Y(w_mem_inst__abc_21378_n5686) );
  OR2X2 OR2X2_3395 ( .A(w_mem_inst__abc_21378_n5686), .B(w_mem_inst__abc_21378_n5682), .Y(w_mem_inst__0w_mem_2__31_0__5_) );
  OR2X2 OR2X2_3396 ( .A(w_mem_inst__abc_21378_n5691), .B(w_mem_inst__abc_21378_n5689), .Y(w_mem_inst__abc_21378_n5692) );
  OR2X2 OR2X2_3397 ( .A(w_mem_inst__abc_21378_n5692), .B(w_mem_inst__abc_21378_n5688), .Y(w_mem_inst__0w_mem_2__31_0__6_) );
  OR2X2 OR2X2_3398 ( .A(w_mem_inst__abc_21378_n5697), .B(w_mem_inst__abc_21378_n5695), .Y(w_mem_inst__abc_21378_n5698) );
  OR2X2 OR2X2_3399 ( .A(w_mem_inst__abc_21378_n5698), .B(w_mem_inst__abc_21378_n5694), .Y(w_mem_inst__0w_mem_2__31_0__7_) );
  OR2X2 OR2X2_34 ( .A(_auto_iopadmap_cc_313_execute_26059_8_), .B(e_reg_8_), .Y(_abc_15724_n818) );
  OR2X2 OR2X2_340 ( .A(_auto_iopadmap_cc_313_execute_26059_80_), .B(c_reg_16_), .Y(_abc_15724_n1754_1) );
  OR2X2 OR2X2_3400 ( .A(w_mem_inst__abc_21378_n5703), .B(w_mem_inst__abc_21378_n5701), .Y(w_mem_inst__abc_21378_n5704) );
  OR2X2 OR2X2_3401 ( .A(w_mem_inst__abc_21378_n5704), .B(w_mem_inst__abc_21378_n5700), .Y(w_mem_inst__0w_mem_2__31_0__8_) );
  OR2X2 OR2X2_3402 ( .A(w_mem_inst__abc_21378_n5709), .B(w_mem_inst__abc_21378_n5707), .Y(w_mem_inst__abc_21378_n5710) );
  OR2X2 OR2X2_3403 ( .A(w_mem_inst__abc_21378_n5710), .B(w_mem_inst__abc_21378_n5706), .Y(w_mem_inst__0w_mem_2__31_0__9_) );
  OR2X2 OR2X2_3404 ( .A(w_mem_inst__abc_21378_n5715), .B(w_mem_inst__abc_21378_n5713), .Y(w_mem_inst__abc_21378_n5716) );
  OR2X2 OR2X2_3405 ( .A(w_mem_inst__abc_21378_n5716), .B(w_mem_inst__abc_21378_n5712), .Y(w_mem_inst__0w_mem_2__31_0__10_) );
  OR2X2 OR2X2_3406 ( .A(w_mem_inst__abc_21378_n5721), .B(w_mem_inst__abc_21378_n5719), .Y(w_mem_inst__abc_21378_n5722) );
  OR2X2 OR2X2_3407 ( .A(w_mem_inst__abc_21378_n5722), .B(w_mem_inst__abc_21378_n5718), .Y(w_mem_inst__0w_mem_2__31_0__11_) );
  OR2X2 OR2X2_3408 ( .A(w_mem_inst__abc_21378_n5727), .B(w_mem_inst__abc_21378_n5725), .Y(w_mem_inst__abc_21378_n5728) );
  OR2X2 OR2X2_3409 ( .A(w_mem_inst__abc_21378_n5728), .B(w_mem_inst__abc_21378_n5724), .Y(w_mem_inst__0w_mem_2__31_0__12_) );
  OR2X2 OR2X2_341 ( .A(_abc_15724_n1753), .B(_abc_15724_n1757), .Y(_abc_15724_n1758_1) );
  OR2X2 OR2X2_3410 ( .A(w_mem_inst__abc_21378_n5733), .B(w_mem_inst__abc_21378_n5731), .Y(w_mem_inst__abc_21378_n5734) );
  OR2X2 OR2X2_3411 ( .A(w_mem_inst__abc_21378_n5734), .B(w_mem_inst__abc_21378_n5730), .Y(w_mem_inst__0w_mem_2__31_0__13_) );
  OR2X2 OR2X2_3412 ( .A(w_mem_inst__abc_21378_n5739), .B(w_mem_inst__abc_21378_n5737), .Y(w_mem_inst__abc_21378_n5740) );
  OR2X2 OR2X2_3413 ( .A(w_mem_inst__abc_21378_n5740), .B(w_mem_inst__abc_21378_n5736), .Y(w_mem_inst__0w_mem_2__31_0__14_) );
  OR2X2 OR2X2_3414 ( .A(w_mem_inst__abc_21378_n5745), .B(w_mem_inst__abc_21378_n5743), .Y(w_mem_inst__abc_21378_n5746) );
  OR2X2 OR2X2_3415 ( .A(w_mem_inst__abc_21378_n5746), .B(w_mem_inst__abc_21378_n5742), .Y(w_mem_inst__0w_mem_2__31_0__15_) );
  OR2X2 OR2X2_3416 ( .A(w_mem_inst__abc_21378_n5751), .B(w_mem_inst__abc_21378_n5749), .Y(w_mem_inst__abc_21378_n5752) );
  OR2X2 OR2X2_3417 ( .A(w_mem_inst__abc_21378_n5752), .B(w_mem_inst__abc_21378_n5748), .Y(w_mem_inst__0w_mem_2__31_0__16_) );
  OR2X2 OR2X2_3418 ( .A(w_mem_inst__abc_21378_n5757), .B(w_mem_inst__abc_21378_n5755), .Y(w_mem_inst__abc_21378_n5758) );
  OR2X2 OR2X2_3419 ( .A(w_mem_inst__abc_21378_n5758), .B(w_mem_inst__abc_21378_n5754), .Y(w_mem_inst__0w_mem_2__31_0__17_) );
  OR2X2 OR2X2_342 ( .A(_abc_15724_n1762_1), .B(_abc_15724_n1739), .Y(H2_reg_16__FF_INPUT) );
  OR2X2 OR2X2_3420 ( .A(w_mem_inst__abc_21378_n5763), .B(w_mem_inst__abc_21378_n5761), .Y(w_mem_inst__abc_21378_n5764) );
  OR2X2 OR2X2_3421 ( .A(w_mem_inst__abc_21378_n5764), .B(w_mem_inst__abc_21378_n5760), .Y(w_mem_inst__0w_mem_2__31_0__18_) );
  OR2X2 OR2X2_3422 ( .A(w_mem_inst__abc_21378_n5769), .B(w_mem_inst__abc_21378_n5767), .Y(w_mem_inst__abc_21378_n5770) );
  OR2X2 OR2X2_3423 ( .A(w_mem_inst__abc_21378_n5770), .B(w_mem_inst__abc_21378_n5766), .Y(w_mem_inst__0w_mem_2__31_0__19_) );
  OR2X2 OR2X2_3424 ( .A(w_mem_inst__abc_21378_n5775), .B(w_mem_inst__abc_21378_n5773), .Y(w_mem_inst__abc_21378_n5776) );
  OR2X2 OR2X2_3425 ( .A(w_mem_inst__abc_21378_n5776), .B(w_mem_inst__abc_21378_n5772), .Y(w_mem_inst__0w_mem_2__31_0__20_) );
  OR2X2 OR2X2_3426 ( .A(w_mem_inst__abc_21378_n5781), .B(w_mem_inst__abc_21378_n5779), .Y(w_mem_inst__abc_21378_n5782) );
  OR2X2 OR2X2_3427 ( .A(w_mem_inst__abc_21378_n5782), .B(w_mem_inst__abc_21378_n5778), .Y(w_mem_inst__0w_mem_2__31_0__21_) );
  OR2X2 OR2X2_3428 ( .A(w_mem_inst__abc_21378_n5787), .B(w_mem_inst__abc_21378_n5785), .Y(w_mem_inst__abc_21378_n5788) );
  OR2X2 OR2X2_3429 ( .A(w_mem_inst__abc_21378_n5788), .B(w_mem_inst__abc_21378_n5784), .Y(w_mem_inst__0w_mem_2__31_0__22_) );
  OR2X2 OR2X2_343 ( .A(_auto_iopadmap_cc_313_execute_26059_81_), .B(c_reg_17_), .Y(_abc_15724_n1766) );
  OR2X2 OR2X2_3430 ( .A(w_mem_inst__abc_21378_n5793), .B(w_mem_inst__abc_21378_n5791), .Y(w_mem_inst__abc_21378_n5794) );
  OR2X2 OR2X2_3431 ( .A(w_mem_inst__abc_21378_n5794), .B(w_mem_inst__abc_21378_n5790), .Y(w_mem_inst__0w_mem_2__31_0__23_) );
  OR2X2 OR2X2_3432 ( .A(w_mem_inst__abc_21378_n5799), .B(w_mem_inst__abc_21378_n5797), .Y(w_mem_inst__abc_21378_n5800) );
  OR2X2 OR2X2_3433 ( .A(w_mem_inst__abc_21378_n5800), .B(w_mem_inst__abc_21378_n5796), .Y(w_mem_inst__0w_mem_2__31_0__24_) );
  OR2X2 OR2X2_3434 ( .A(w_mem_inst__abc_21378_n5805), .B(w_mem_inst__abc_21378_n5803), .Y(w_mem_inst__abc_21378_n5806) );
  OR2X2 OR2X2_3435 ( .A(w_mem_inst__abc_21378_n5806), .B(w_mem_inst__abc_21378_n5802), .Y(w_mem_inst__0w_mem_2__31_0__25_) );
  OR2X2 OR2X2_3436 ( .A(w_mem_inst__abc_21378_n5811), .B(w_mem_inst__abc_21378_n5809), .Y(w_mem_inst__abc_21378_n5812) );
  OR2X2 OR2X2_3437 ( .A(w_mem_inst__abc_21378_n5812), .B(w_mem_inst__abc_21378_n5808), .Y(w_mem_inst__0w_mem_2__31_0__26_) );
  OR2X2 OR2X2_3438 ( .A(w_mem_inst__abc_21378_n5817), .B(w_mem_inst__abc_21378_n5815), .Y(w_mem_inst__abc_21378_n5818) );
  OR2X2 OR2X2_3439 ( .A(w_mem_inst__abc_21378_n5818), .B(w_mem_inst__abc_21378_n5814), .Y(w_mem_inst__0w_mem_2__31_0__27_) );
  OR2X2 OR2X2_344 ( .A(_abc_15724_n1765), .B(_abc_15724_n1769), .Y(_abc_15724_n1770) );
  OR2X2 OR2X2_3440 ( .A(w_mem_inst__abc_21378_n5823), .B(w_mem_inst__abc_21378_n5821), .Y(w_mem_inst__abc_21378_n5824) );
  OR2X2 OR2X2_3441 ( .A(w_mem_inst__abc_21378_n5824), .B(w_mem_inst__abc_21378_n5820), .Y(w_mem_inst__0w_mem_2__31_0__28_) );
  OR2X2 OR2X2_3442 ( .A(w_mem_inst__abc_21378_n5829), .B(w_mem_inst__abc_21378_n5827), .Y(w_mem_inst__abc_21378_n5830) );
  OR2X2 OR2X2_3443 ( .A(w_mem_inst__abc_21378_n5830), .B(w_mem_inst__abc_21378_n5826), .Y(w_mem_inst__0w_mem_2__31_0__29_) );
  OR2X2 OR2X2_3444 ( .A(w_mem_inst__abc_21378_n5835), .B(w_mem_inst__abc_21378_n5833), .Y(w_mem_inst__abc_21378_n5836) );
  OR2X2 OR2X2_3445 ( .A(w_mem_inst__abc_21378_n5836), .B(w_mem_inst__abc_21378_n5832), .Y(w_mem_inst__0w_mem_2__31_0__30_) );
  OR2X2 OR2X2_3446 ( .A(w_mem_inst__abc_21378_n5841), .B(w_mem_inst__abc_21378_n5839), .Y(w_mem_inst__abc_21378_n5842) );
  OR2X2 OR2X2_3447 ( .A(w_mem_inst__abc_21378_n5842), .B(w_mem_inst__abc_21378_n5838), .Y(w_mem_inst__0w_mem_2__31_0__31_) );
  OR2X2 OR2X2_3448 ( .A(w_mem_inst__abc_21378_n5847), .B(w_mem_inst__abc_21378_n5845), .Y(w_mem_inst__abc_21378_n5848) );
  OR2X2 OR2X2_3449 ( .A(w_mem_inst__abc_21378_n5848), .B(w_mem_inst__abc_21378_n5844), .Y(w_mem_inst__0w_mem_1__31_0__0_) );
  OR2X2 OR2X2_345 ( .A(_abc_15724_n1764), .B(_abc_15724_n1771), .Y(_abc_15724_n1772_1) );
  OR2X2 OR2X2_3450 ( .A(w_mem_inst__abc_21378_n5853), .B(w_mem_inst__abc_21378_n5851), .Y(w_mem_inst__abc_21378_n5854) );
  OR2X2 OR2X2_3451 ( .A(w_mem_inst__abc_21378_n5854), .B(w_mem_inst__abc_21378_n5850), .Y(w_mem_inst__0w_mem_1__31_0__1_) );
  OR2X2 OR2X2_3452 ( .A(w_mem_inst__abc_21378_n5859), .B(w_mem_inst__abc_21378_n5857), .Y(w_mem_inst__abc_21378_n5860) );
  OR2X2 OR2X2_3453 ( .A(w_mem_inst__abc_21378_n5860), .B(w_mem_inst__abc_21378_n5856), .Y(w_mem_inst__0w_mem_1__31_0__2_) );
  OR2X2 OR2X2_3454 ( .A(w_mem_inst__abc_21378_n5865), .B(w_mem_inst__abc_21378_n5863), .Y(w_mem_inst__abc_21378_n5866) );
  OR2X2 OR2X2_3455 ( .A(w_mem_inst__abc_21378_n5866), .B(w_mem_inst__abc_21378_n5862), .Y(w_mem_inst__0w_mem_1__31_0__3_) );
  OR2X2 OR2X2_3456 ( .A(w_mem_inst__abc_21378_n5871), .B(w_mem_inst__abc_21378_n5869), .Y(w_mem_inst__abc_21378_n5872) );
  OR2X2 OR2X2_3457 ( .A(w_mem_inst__abc_21378_n5872), .B(w_mem_inst__abc_21378_n5868), .Y(w_mem_inst__0w_mem_1__31_0__4_) );
  OR2X2 OR2X2_3458 ( .A(w_mem_inst__abc_21378_n5877), .B(w_mem_inst__abc_21378_n5875), .Y(w_mem_inst__abc_21378_n5878) );
  OR2X2 OR2X2_3459 ( .A(w_mem_inst__abc_21378_n5878), .B(w_mem_inst__abc_21378_n5874), .Y(w_mem_inst__0w_mem_1__31_0__5_) );
  OR2X2 OR2X2_346 ( .A(_abc_15724_n851_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_81_), .Y(_abc_15724_n1775) );
  OR2X2 OR2X2_3460 ( .A(w_mem_inst__abc_21378_n5883), .B(w_mem_inst__abc_21378_n5881), .Y(w_mem_inst__abc_21378_n5884) );
  OR2X2 OR2X2_3461 ( .A(w_mem_inst__abc_21378_n5884), .B(w_mem_inst__abc_21378_n5880), .Y(w_mem_inst__0w_mem_1__31_0__6_) );
  OR2X2 OR2X2_3462 ( .A(w_mem_inst__abc_21378_n5889), .B(w_mem_inst__abc_21378_n5887), .Y(w_mem_inst__abc_21378_n5890) );
  OR2X2 OR2X2_3463 ( .A(w_mem_inst__abc_21378_n5890), .B(w_mem_inst__abc_21378_n5886), .Y(w_mem_inst__0w_mem_1__31_0__7_) );
  OR2X2 OR2X2_3464 ( .A(w_mem_inst__abc_21378_n5895), .B(w_mem_inst__abc_21378_n5893), .Y(w_mem_inst__abc_21378_n5896) );
  OR2X2 OR2X2_3465 ( .A(w_mem_inst__abc_21378_n5896), .B(w_mem_inst__abc_21378_n5892), .Y(w_mem_inst__0w_mem_1__31_0__8_) );
  OR2X2 OR2X2_3466 ( .A(w_mem_inst__abc_21378_n5901), .B(w_mem_inst__abc_21378_n5899), .Y(w_mem_inst__abc_21378_n5902) );
  OR2X2 OR2X2_3467 ( .A(w_mem_inst__abc_21378_n5902), .B(w_mem_inst__abc_21378_n5898), .Y(w_mem_inst__0w_mem_1__31_0__9_) );
  OR2X2 OR2X2_3468 ( .A(w_mem_inst__abc_21378_n5907), .B(w_mem_inst__abc_21378_n5905), .Y(w_mem_inst__abc_21378_n5908) );
  OR2X2 OR2X2_3469 ( .A(w_mem_inst__abc_21378_n5908), .B(w_mem_inst__abc_21378_n5904), .Y(w_mem_inst__0w_mem_1__31_0__10_) );
  OR2X2 OR2X2_347 ( .A(_abc_15724_n1774), .B(_abc_15724_n1776), .Y(H2_reg_17__FF_INPUT) );
  OR2X2 OR2X2_3470 ( .A(w_mem_inst__abc_21378_n5913), .B(w_mem_inst__abc_21378_n5911), .Y(w_mem_inst__abc_21378_n5914) );
  OR2X2 OR2X2_3471 ( .A(w_mem_inst__abc_21378_n5914), .B(w_mem_inst__abc_21378_n5910), .Y(w_mem_inst__0w_mem_1__31_0__11_) );
  OR2X2 OR2X2_3472 ( .A(w_mem_inst__abc_21378_n5919), .B(w_mem_inst__abc_21378_n5917), .Y(w_mem_inst__abc_21378_n5920) );
  OR2X2 OR2X2_3473 ( .A(w_mem_inst__abc_21378_n5920), .B(w_mem_inst__abc_21378_n5916), .Y(w_mem_inst__0w_mem_1__31_0__12_) );
  OR2X2 OR2X2_3474 ( .A(w_mem_inst__abc_21378_n5925), .B(w_mem_inst__abc_21378_n5923), .Y(w_mem_inst__abc_21378_n5926) );
  OR2X2 OR2X2_3475 ( .A(w_mem_inst__abc_21378_n5926), .B(w_mem_inst__abc_21378_n5922), .Y(w_mem_inst__0w_mem_1__31_0__13_) );
  OR2X2 OR2X2_3476 ( .A(w_mem_inst__abc_21378_n5931), .B(w_mem_inst__abc_21378_n5929), .Y(w_mem_inst__abc_21378_n5932) );
  OR2X2 OR2X2_3477 ( .A(w_mem_inst__abc_21378_n5932), .B(w_mem_inst__abc_21378_n5928), .Y(w_mem_inst__0w_mem_1__31_0__14_) );
  OR2X2 OR2X2_3478 ( .A(w_mem_inst__abc_21378_n5937), .B(w_mem_inst__abc_21378_n5935), .Y(w_mem_inst__abc_21378_n5938) );
  OR2X2 OR2X2_3479 ( .A(w_mem_inst__abc_21378_n5938), .B(w_mem_inst__abc_21378_n5934), .Y(w_mem_inst__0w_mem_1__31_0__15_) );
  OR2X2 OR2X2_348 ( .A(_abc_15724_n1771), .B(_abc_15724_n1756), .Y(_abc_15724_n1779) );
  OR2X2 OR2X2_3480 ( .A(w_mem_inst__abc_21378_n5943), .B(w_mem_inst__abc_21378_n5941), .Y(w_mem_inst__abc_21378_n5944) );
  OR2X2 OR2X2_3481 ( .A(w_mem_inst__abc_21378_n5944), .B(w_mem_inst__abc_21378_n5940), .Y(w_mem_inst__0w_mem_1__31_0__16_) );
  OR2X2 OR2X2_3482 ( .A(w_mem_inst__abc_21378_n5949), .B(w_mem_inst__abc_21378_n5947), .Y(w_mem_inst__abc_21378_n5950) );
  OR2X2 OR2X2_3483 ( .A(w_mem_inst__abc_21378_n5950), .B(w_mem_inst__abc_21378_n5946), .Y(w_mem_inst__0w_mem_1__31_0__17_) );
  OR2X2 OR2X2_3484 ( .A(w_mem_inst__abc_21378_n5955), .B(w_mem_inst__abc_21378_n5953), .Y(w_mem_inst__abc_21378_n5956) );
  OR2X2 OR2X2_3485 ( .A(w_mem_inst__abc_21378_n5956), .B(w_mem_inst__abc_21378_n5952), .Y(w_mem_inst__0w_mem_1__31_0__18_) );
  OR2X2 OR2X2_3486 ( .A(w_mem_inst__abc_21378_n5961), .B(w_mem_inst__abc_21378_n5959), .Y(w_mem_inst__abc_21378_n5962) );
  OR2X2 OR2X2_3487 ( .A(w_mem_inst__abc_21378_n5962), .B(w_mem_inst__abc_21378_n5958), .Y(w_mem_inst__0w_mem_1__31_0__19_) );
  OR2X2 OR2X2_3488 ( .A(w_mem_inst__abc_21378_n5967), .B(w_mem_inst__abc_21378_n5965), .Y(w_mem_inst__abc_21378_n5968) );
  OR2X2 OR2X2_3489 ( .A(w_mem_inst__abc_21378_n5968), .B(w_mem_inst__abc_21378_n5964), .Y(w_mem_inst__0w_mem_1__31_0__20_) );
  OR2X2 OR2X2_349 ( .A(_abc_15724_n1783), .B(_abc_15724_n1781_1), .Y(_abc_15724_n1784) );
  OR2X2 OR2X2_3490 ( .A(w_mem_inst__abc_21378_n5973), .B(w_mem_inst__abc_21378_n5971), .Y(w_mem_inst__abc_21378_n5974) );
  OR2X2 OR2X2_3491 ( .A(w_mem_inst__abc_21378_n5974), .B(w_mem_inst__abc_21378_n5970), .Y(w_mem_inst__0w_mem_1__31_0__21_) );
  OR2X2 OR2X2_3492 ( .A(w_mem_inst__abc_21378_n5979), .B(w_mem_inst__abc_21378_n5977), .Y(w_mem_inst__abc_21378_n5980) );
  OR2X2 OR2X2_3493 ( .A(w_mem_inst__abc_21378_n5980), .B(w_mem_inst__abc_21378_n5976), .Y(w_mem_inst__0w_mem_1__31_0__22_) );
  OR2X2 OR2X2_3494 ( .A(w_mem_inst__abc_21378_n5985), .B(w_mem_inst__abc_21378_n5983), .Y(w_mem_inst__abc_21378_n5986) );
  OR2X2 OR2X2_3495 ( .A(w_mem_inst__abc_21378_n5986), .B(w_mem_inst__abc_21378_n5982), .Y(w_mem_inst__0w_mem_1__31_0__23_) );
  OR2X2 OR2X2_3496 ( .A(w_mem_inst__abc_21378_n5991), .B(w_mem_inst__abc_21378_n5989), .Y(w_mem_inst__abc_21378_n5992) );
  OR2X2 OR2X2_3497 ( .A(w_mem_inst__abc_21378_n5992), .B(w_mem_inst__abc_21378_n5988), .Y(w_mem_inst__0w_mem_1__31_0__24_) );
  OR2X2 OR2X2_3498 ( .A(w_mem_inst__abc_21378_n5997), .B(w_mem_inst__abc_21378_n5995), .Y(w_mem_inst__abc_21378_n5998) );
  OR2X2 OR2X2_3499 ( .A(w_mem_inst__abc_21378_n5998), .B(w_mem_inst__abc_21378_n5994), .Y(w_mem_inst__0w_mem_1__31_0__25_) );
  OR2X2 OR2X2_35 ( .A(_abc_15724_n822), .B(_abc_15724_n772), .Y(_abc_15724_n823) );
  OR2X2 OR2X2_350 ( .A(_auto_iopadmap_cc_313_execute_26059_82_), .B(c_reg_18_), .Y(_abc_15724_n1785) );
  OR2X2 OR2X2_3500 ( .A(w_mem_inst__abc_21378_n6003), .B(w_mem_inst__abc_21378_n6001), .Y(w_mem_inst__abc_21378_n6004) );
  OR2X2 OR2X2_3501 ( .A(w_mem_inst__abc_21378_n6004), .B(w_mem_inst__abc_21378_n6000), .Y(w_mem_inst__0w_mem_1__31_0__26_) );
  OR2X2 OR2X2_3502 ( .A(w_mem_inst__abc_21378_n6009), .B(w_mem_inst__abc_21378_n6007), .Y(w_mem_inst__abc_21378_n6010) );
  OR2X2 OR2X2_3503 ( .A(w_mem_inst__abc_21378_n6010), .B(w_mem_inst__abc_21378_n6006), .Y(w_mem_inst__0w_mem_1__31_0__27_) );
  OR2X2 OR2X2_3504 ( .A(w_mem_inst__abc_21378_n6015), .B(w_mem_inst__abc_21378_n6013), .Y(w_mem_inst__abc_21378_n6016) );
  OR2X2 OR2X2_3505 ( .A(w_mem_inst__abc_21378_n6016), .B(w_mem_inst__abc_21378_n6012), .Y(w_mem_inst__0w_mem_1__31_0__28_) );
  OR2X2 OR2X2_3506 ( .A(w_mem_inst__abc_21378_n6021), .B(w_mem_inst__abc_21378_n6019), .Y(w_mem_inst__abc_21378_n6022) );
  OR2X2 OR2X2_3507 ( .A(w_mem_inst__abc_21378_n6022), .B(w_mem_inst__abc_21378_n6018), .Y(w_mem_inst__0w_mem_1__31_0__29_) );
  OR2X2 OR2X2_3508 ( .A(w_mem_inst__abc_21378_n6027), .B(w_mem_inst__abc_21378_n6025), .Y(w_mem_inst__abc_21378_n6028) );
  OR2X2 OR2X2_3509 ( .A(w_mem_inst__abc_21378_n6028), .B(w_mem_inst__abc_21378_n6024), .Y(w_mem_inst__0w_mem_1__31_0__30_) );
  OR2X2 OR2X2_351 ( .A(_abc_15724_n1784), .B(_abc_15724_n1788), .Y(_abc_15724_n1789) );
  OR2X2 OR2X2_3510 ( .A(w_mem_inst__abc_21378_n6033), .B(w_mem_inst__abc_21378_n6031), .Y(w_mem_inst__abc_21378_n6034) );
  OR2X2 OR2X2_3511 ( .A(w_mem_inst__abc_21378_n6034), .B(w_mem_inst__abc_21378_n6030), .Y(w_mem_inst__0w_mem_1__31_0__31_) );
  OR2X2 OR2X2_3512 ( .A(w_mem_inst__abc_21378_n6039), .B(w_mem_inst__abc_21378_n6037), .Y(w_mem_inst__abc_21378_n6040) );
  OR2X2 OR2X2_3513 ( .A(w_mem_inst__abc_21378_n6040), .B(w_mem_inst__abc_21378_n6036), .Y(w_mem_inst__0w_mem_0__31_0__0_) );
  OR2X2 OR2X2_3514 ( .A(w_mem_inst__abc_21378_n6045), .B(w_mem_inst__abc_21378_n6043), .Y(w_mem_inst__abc_21378_n6046) );
  OR2X2 OR2X2_3515 ( .A(w_mem_inst__abc_21378_n6046), .B(w_mem_inst__abc_21378_n6042), .Y(w_mem_inst__0w_mem_0__31_0__1_) );
  OR2X2 OR2X2_3516 ( .A(w_mem_inst__abc_21378_n6051), .B(w_mem_inst__abc_21378_n6049), .Y(w_mem_inst__abc_21378_n6052) );
  OR2X2 OR2X2_3517 ( .A(w_mem_inst__abc_21378_n6052), .B(w_mem_inst__abc_21378_n6048), .Y(w_mem_inst__0w_mem_0__31_0__2_) );
  OR2X2 OR2X2_3518 ( .A(w_mem_inst__abc_21378_n6057), .B(w_mem_inst__abc_21378_n6055), .Y(w_mem_inst__abc_21378_n6058) );
  OR2X2 OR2X2_3519 ( .A(w_mem_inst__abc_21378_n6058), .B(w_mem_inst__abc_21378_n6054), .Y(w_mem_inst__0w_mem_0__31_0__3_) );
  OR2X2 OR2X2_352 ( .A(_abc_15724_n1793), .B(_abc_15724_n1778), .Y(H2_reg_18__FF_INPUT) );
  OR2X2 OR2X2_3520 ( .A(w_mem_inst__abc_21378_n6063), .B(w_mem_inst__abc_21378_n6061), .Y(w_mem_inst__abc_21378_n6064) );
  OR2X2 OR2X2_3521 ( .A(w_mem_inst__abc_21378_n6064), .B(w_mem_inst__abc_21378_n6060), .Y(w_mem_inst__0w_mem_0__31_0__4_) );
  OR2X2 OR2X2_3522 ( .A(w_mem_inst__abc_21378_n6069), .B(w_mem_inst__abc_21378_n6067), .Y(w_mem_inst__abc_21378_n6070) );
  OR2X2 OR2X2_3523 ( .A(w_mem_inst__abc_21378_n6070), .B(w_mem_inst__abc_21378_n6066), .Y(w_mem_inst__0w_mem_0__31_0__5_) );
  OR2X2 OR2X2_3524 ( .A(w_mem_inst__abc_21378_n6075), .B(w_mem_inst__abc_21378_n6073), .Y(w_mem_inst__abc_21378_n6076) );
  OR2X2 OR2X2_3525 ( .A(w_mem_inst__abc_21378_n6076), .B(w_mem_inst__abc_21378_n6072), .Y(w_mem_inst__0w_mem_0__31_0__6_) );
  OR2X2 OR2X2_3526 ( .A(w_mem_inst__abc_21378_n6081), .B(w_mem_inst__abc_21378_n6079), .Y(w_mem_inst__abc_21378_n6082) );
  OR2X2 OR2X2_3527 ( .A(w_mem_inst__abc_21378_n6082), .B(w_mem_inst__abc_21378_n6078), .Y(w_mem_inst__0w_mem_0__31_0__7_) );
  OR2X2 OR2X2_3528 ( .A(w_mem_inst__abc_21378_n6087), .B(w_mem_inst__abc_21378_n6085), .Y(w_mem_inst__abc_21378_n6088) );
  OR2X2 OR2X2_3529 ( .A(w_mem_inst__abc_21378_n6088), .B(w_mem_inst__abc_21378_n6084), .Y(w_mem_inst__0w_mem_0__31_0__8_) );
  OR2X2 OR2X2_353 ( .A(_auto_iopadmap_cc_313_execute_26059_83_), .B(c_reg_19_), .Y(_abc_15724_n1797) );
  OR2X2 OR2X2_3530 ( .A(w_mem_inst__abc_21378_n6093), .B(w_mem_inst__abc_21378_n6091), .Y(w_mem_inst__abc_21378_n6094) );
  OR2X2 OR2X2_3531 ( .A(w_mem_inst__abc_21378_n6094), .B(w_mem_inst__abc_21378_n6090), .Y(w_mem_inst__0w_mem_0__31_0__9_) );
  OR2X2 OR2X2_3532 ( .A(w_mem_inst__abc_21378_n6099), .B(w_mem_inst__abc_21378_n6097), .Y(w_mem_inst__abc_21378_n6100) );
  OR2X2 OR2X2_3533 ( .A(w_mem_inst__abc_21378_n6100), .B(w_mem_inst__abc_21378_n6096), .Y(w_mem_inst__0w_mem_0__31_0__10_) );
  OR2X2 OR2X2_3534 ( .A(w_mem_inst__abc_21378_n6105), .B(w_mem_inst__abc_21378_n6103), .Y(w_mem_inst__abc_21378_n6106) );
  OR2X2 OR2X2_3535 ( .A(w_mem_inst__abc_21378_n6106), .B(w_mem_inst__abc_21378_n6102), .Y(w_mem_inst__0w_mem_0__31_0__11_) );
  OR2X2 OR2X2_3536 ( .A(w_mem_inst__abc_21378_n6111), .B(w_mem_inst__abc_21378_n6109), .Y(w_mem_inst__abc_21378_n6112) );
  OR2X2 OR2X2_3537 ( .A(w_mem_inst__abc_21378_n6112), .B(w_mem_inst__abc_21378_n6108), .Y(w_mem_inst__0w_mem_0__31_0__12_) );
  OR2X2 OR2X2_3538 ( .A(w_mem_inst__abc_21378_n6117), .B(w_mem_inst__abc_21378_n6115), .Y(w_mem_inst__abc_21378_n6118) );
  OR2X2 OR2X2_3539 ( .A(w_mem_inst__abc_21378_n6118), .B(w_mem_inst__abc_21378_n6114), .Y(w_mem_inst__0w_mem_0__31_0__13_) );
  OR2X2 OR2X2_354 ( .A(_abc_15724_n1796), .B(_abc_15724_n1800), .Y(_abc_15724_n1801) );
  OR2X2 OR2X2_3540 ( .A(w_mem_inst__abc_21378_n6123), .B(w_mem_inst__abc_21378_n6121), .Y(w_mem_inst__abc_21378_n6124) );
  OR2X2 OR2X2_3541 ( .A(w_mem_inst__abc_21378_n6124), .B(w_mem_inst__abc_21378_n6120), .Y(w_mem_inst__0w_mem_0__31_0__14_) );
  OR2X2 OR2X2_3542 ( .A(w_mem_inst__abc_21378_n6129), .B(w_mem_inst__abc_21378_n6127), .Y(w_mem_inst__abc_21378_n6130) );
  OR2X2 OR2X2_3543 ( .A(w_mem_inst__abc_21378_n6130), .B(w_mem_inst__abc_21378_n6126), .Y(w_mem_inst__0w_mem_0__31_0__15_) );
  OR2X2 OR2X2_3544 ( .A(w_mem_inst__abc_21378_n6135), .B(w_mem_inst__abc_21378_n6133), .Y(w_mem_inst__abc_21378_n6136) );
  OR2X2 OR2X2_3545 ( .A(w_mem_inst__abc_21378_n6136), .B(w_mem_inst__abc_21378_n6132), .Y(w_mem_inst__0w_mem_0__31_0__16_) );
  OR2X2 OR2X2_3546 ( .A(w_mem_inst__abc_21378_n6141), .B(w_mem_inst__abc_21378_n6139), .Y(w_mem_inst__abc_21378_n6142) );
  OR2X2 OR2X2_3547 ( .A(w_mem_inst__abc_21378_n6142), .B(w_mem_inst__abc_21378_n6138), .Y(w_mem_inst__0w_mem_0__31_0__17_) );
  OR2X2 OR2X2_3548 ( .A(w_mem_inst__abc_21378_n6147), .B(w_mem_inst__abc_21378_n6145), .Y(w_mem_inst__abc_21378_n6148) );
  OR2X2 OR2X2_3549 ( .A(w_mem_inst__abc_21378_n6148), .B(w_mem_inst__abc_21378_n6144), .Y(w_mem_inst__0w_mem_0__31_0__18_) );
  OR2X2 OR2X2_355 ( .A(_abc_15724_n1795_1), .B(_abc_15724_n1802), .Y(_abc_15724_n1803) );
  OR2X2 OR2X2_3550 ( .A(w_mem_inst__abc_21378_n6153), .B(w_mem_inst__abc_21378_n6151), .Y(w_mem_inst__abc_21378_n6154) );
  OR2X2 OR2X2_3551 ( .A(w_mem_inst__abc_21378_n6154), .B(w_mem_inst__abc_21378_n6150), .Y(w_mem_inst__0w_mem_0__31_0__19_) );
  OR2X2 OR2X2_3552 ( .A(w_mem_inst__abc_21378_n6159), .B(w_mem_inst__abc_21378_n6157), .Y(w_mem_inst__abc_21378_n6160) );
  OR2X2 OR2X2_3553 ( .A(w_mem_inst__abc_21378_n6160), .B(w_mem_inst__abc_21378_n6156), .Y(w_mem_inst__0w_mem_0__31_0__20_) );
  OR2X2 OR2X2_3554 ( .A(w_mem_inst__abc_21378_n6165), .B(w_mem_inst__abc_21378_n6163), .Y(w_mem_inst__abc_21378_n6166) );
  OR2X2 OR2X2_3555 ( .A(w_mem_inst__abc_21378_n6166), .B(w_mem_inst__abc_21378_n6162), .Y(w_mem_inst__0w_mem_0__31_0__21_) );
  OR2X2 OR2X2_3556 ( .A(w_mem_inst__abc_21378_n6171), .B(w_mem_inst__abc_21378_n6169), .Y(w_mem_inst__abc_21378_n6172) );
  OR2X2 OR2X2_3557 ( .A(w_mem_inst__abc_21378_n6172), .B(w_mem_inst__abc_21378_n6168), .Y(w_mem_inst__0w_mem_0__31_0__22_) );
  OR2X2 OR2X2_3558 ( .A(w_mem_inst__abc_21378_n6177), .B(w_mem_inst__abc_21378_n6175), .Y(w_mem_inst__abc_21378_n6178) );
  OR2X2 OR2X2_3559 ( .A(w_mem_inst__abc_21378_n6178), .B(w_mem_inst__abc_21378_n6174), .Y(w_mem_inst__0w_mem_0__31_0__23_) );
  OR2X2 OR2X2_356 ( .A(_abc_15724_n851_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_83_), .Y(_abc_15724_n1806) );
  OR2X2 OR2X2_3560 ( .A(w_mem_inst__abc_21378_n6183), .B(w_mem_inst__abc_21378_n6181), .Y(w_mem_inst__abc_21378_n6184) );
  OR2X2 OR2X2_3561 ( .A(w_mem_inst__abc_21378_n6184), .B(w_mem_inst__abc_21378_n6180), .Y(w_mem_inst__0w_mem_0__31_0__24_) );
  OR2X2 OR2X2_3562 ( .A(w_mem_inst__abc_21378_n6189), .B(w_mem_inst__abc_21378_n6187), .Y(w_mem_inst__abc_21378_n6190) );
  OR2X2 OR2X2_3563 ( .A(w_mem_inst__abc_21378_n6190), .B(w_mem_inst__abc_21378_n6186), .Y(w_mem_inst__0w_mem_0__31_0__25_) );
  OR2X2 OR2X2_3564 ( .A(w_mem_inst__abc_21378_n6195), .B(w_mem_inst__abc_21378_n6193), .Y(w_mem_inst__abc_21378_n6196) );
  OR2X2 OR2X2_3565 ( .A(w_mem_inst__abc_21378_n6196), .B(w_mem_inst__abc_21378_n6192), .Y(w_mem_inst__0w_mem_0__31_0__26_) );
  OR2X2 OR2X2_3566 ( .A(w_mem_inst__abc_21378_n6201), .B(w_mem_inst__abc_21378_n6199), .Y(w_mem_inst__abc_21378_n6202) );
  OR2X2 OR2X2_3567 ( .A(w_mem_inst__abc_21378_n6202), .B(w_mem_inst__abc_21378_n6198), .Y(w_mem_inst__0w_mem_0__31_0__27_) );
  OR2X2 OR2X2_3568 ( .A(w_mem_inst__abc_21378_n6207), .B(w_mem_inst__abc_21378_n6205), .Y(w_mem_inst__abc_21378_n6208) );
  OR2X2 OR2X2_3569 ( .A(w_mem_inst__abc_21378_n6208), .B(w_mem_inst__abc_21378_n6204), .Y(w_mem_inst__0w_mem_0__31_0__28_) );
  OR2X2 OR2X2_357 ( .A(_abc_15724_n1805), .B(_abc_15724_n1807), .Y(H2_reg_19__FF_INPUT) );
  OR2X2 OR2X2_3570 ( .A(w_mem_inst__abc_21378_n6213), .B(w_mem_inst__abc_21378_n6211), .Y(w_mem_inst__abc_21378_n6214) );
  OR2X2 OR2X2_3571 ( .A(w_mem_inst__abc_21378_n6214), .B(w_mem_inst__abc_21378_n6210), .Y(w_mem_inst__0w_mem_0__31_0__29_) );
  OR2X2 OR2X2_3572 ( .A(w_mem_inst__abc_21378_n6219), .B(w_mem_inst__abc_21378_n6217), .Y(w_mem_inst__abc_21378_n6220) );
  OR2X2 OR2X2_3573 ( .A(w_mem_inst__abc_21378_n6220), .B(w_mem_inst__abc_21378_n6216), .Y(w_mem_inst__0w_mem_0__31_0__30_) );
  OR2X2 OR2X2_3574 ( .A(w_mem_inst__abc_21378_n6225), .B(w_mem_inst__abc_21378_n6223), .Y(w_mem_inst__abc_21378_n6226) );
  OR2X2 OR2X2_3575 ( .A(w_mem_inst__abc_21378_n6226), .B(w_mem_inst__abc_21378_n6222), .Y(w_mem_inst__0w_mem_0__31_0__31_) );
  OR2X2 OR2X2_3576 ( .A(w_mem_inst_w_ctr_reg_0_), .B(round_ctr_inc_bF_buf11), .Y(w_mem_inst__abc_21378_n6228) );
  OR2X2 OR2X2_3577 ( .A(w_mem_inst__abc_21378_n6230), .B(w_mem_inst__abc_21378_n1623_1), .Y(w_mem_inst__abc_21378_n6231) );
  OR2X2 OR2X2_3578 ( .A(w_mem_inst__abc_21378_n1615_1), .B(w_mem_inst__abc_21378_n1624), .Y(w_mem_inst__abc_21378_n6234) );
  OR2X2 OR2X2_3579 ( .A(w_mem_inst__abc_21378_n6235), .B(w_mem_inst__abc_21378_n6233), .Y(w_mem_inst_w_ctr_reg_1__FF_INPUT) );
  OR2X2 OR2X2_358 ( .A(_abc_15724_n1752), .B(_abc_15724_n1811), .Y(_abc_15724_n1812) );
  OR2X2 OR2X2_3580 ( .A(w_mem_inst__abc_21378_n3156_bF_buf0), .B(round_ctr_inc_bF_buf8), .Y(w_mem_inst__abc_21378_n6237) );
  OR2X2 OR2X2_3581 ( .A(w_mem_inst__abc_21378_n6238), .B(w_mem_inst__abc_21378_n6239), .Y(w_mem_inst__abc_21378_n6240) );
  OR2X2 OR2X2_3582 ( .A(w_mem_inst__abc_21378_n6242), .B(w_mem_inst__abc_21378_n6245), .Y(w_mem_inst__abc_21378_n6246) );
  OR2X2 OR2X2_3583 ( .A(w_mem_inst__abc_21378_n6247), .B(w_mem_inst__abc_21378_n6250), .Y(w_mem_inst__abc_21378_n6251) );
  OR2X2 OR2X2_3584 ( .A(w_mem_inst__abc_21378_n6252), .B(w_mem_inst__abc_21378_n6255), .Y(w_mem_inst__abc_21378_n6256) );
  OR2X2 OR2X2_3585 ( .A(w_mem_inst__abc_21378_n6257), .B(w_mem_inst__abc_21378_n6260), .Y(w_mem_inst__abc_21378_n6261) );
  OR2X2 OR2X2_359 ( .A(_abc_15724_n1814), .B(_abc_15724_n1798), .Y(_abc_15724_n1815) );
  OR2X2 OR2X2_36 ( .A(_abc_15724_n824_1), .B(_abc_15724_n749), .Y(_abc_15724_n825_1) );
  OR2X2 OR2X2_360 ( .A(_abc_15724_n1813_1), .B(_abc_15724_n1815), .Y(_abc_15724_n1816) );
  OR2X2 OR2X2_361 ( .A(_auto_iopadmap_cc_313_execute_26059_84_), .B(c_reg_20_), .Y(_abc_15724_n1820) );
  OR2X2 OR2X2_362 ( .A(_abc_15724_n1819), .B(_abc_15724_n1823_1), .Y(_abc_15724_n1824) );
  OR2X2 OR2X2_363 ( .A(_abc_15724_n851_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_84_), .Y(_abc_15724_n1829) );
  OR2X2 OR2X2_364 ( .A(_abc_15724_n1828), .B(_abc_15724_n1830), .Y(H2_reg_20__FF_INPUT) );
  OR2X2 OR2X2_365 ( .A(_auto_iopadmap_cc_313_execute_26059_85_), .B(c_reg_21_), .Y(_abc_15724_n1834) );
  OR2X2 OR2X2_366 ( .A(_abc_15724_n1833), .B(_abc_15724_n1837), .Y(_abc_15724_n1838) );
  OR2X2 OR2X2_367 ( .A(_abc_15724_n1832), .B(_abc_15724_n1839), .Y(_abc_15724_n1840) );
  OR2X2 OR2X2_368 ( .A(_abc_15724_n851_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_85_), .Y(_abc_15724_n1843) );
  OR2X2 OR2X2_369 ( .A(_abc_15724_n1842), .B(_abc_15724_n1844), .Y(H2_reg_21__FF_INPUT) );
  OR2X2 OR2X2_37 ( .A(e_reg_16_), .B(_auto_iopadmap_cc_313_execute_26059_16_), .Y(_abc_15724_n827) );
  OR2X2 OR2X2_370 ( .A(_abc_15724_n1839), .B(_abc_15724_n1822), .Y(_abc_15724_n1847) );
  OR2X2 OR2X2_371 ( .A(_abc_15724_n1851_1), .B(_abc_15724_n1849), .Y(_abc_15724_n1852) );
  OR2X2 OR2X2_372 ( .A(_auto_iopadmap_cc_313_execute_26059_86_), .B(c_reg_22_), .Y(_abc_15724_n1853) );
  OR2X2 OR2X2_373 ( .A(_abc_15724_n1852), .B(_abc_15724_n1856_1), .Y(_abc_15724_n1859) );
  OR2X2 OR2X2_374 ( .A(_abc_15724_n1861_1), .B(_abc_15724_n1846_1), .Y(H2_reg_22__FF_INPUT) );
  OR2X2 OR2X2_375 ( .A(_auto_iopadmap_cc_313_execute_26059_87_), .B(c_reg_23_), .Y(_abc_15724_n1865_1) );
  OR2X2 OR2X2_376 ( .A(_abc_15724_n1864), .B(_abc_15724_n1868), .Y(_abc_15724_n1869) );
  OR2X2 OR2X2_377 ( .A(_abc_15724_n1863), .B(_abc_15724_n1870_1), .Y(_abc_15724_n1871) );
  OR2X2 OR2X2_378 ( .A(_abc_15724_n851_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_87_), .Y(_abc_15724_n1874) );
  OR2X2 OR2X2_379 ( .A(_abc_15724_n1873), .B(_abc_15724_n1875_1), .Y(H2_reg_23__FF_INPUT) );
  OR2X2 OR2X2_38 ( .A(_abc_15724_n826_1), .B(_abc_15724_n831), .Y(_abc_15724_n832_1) );
  OR2X2 OR2X2_380 ( .A(_abc_15724_n1880_1), .B(_abc_15724_n1866), .Y(_abc_15724_n1881) );
  OR2X2 OR2X2_381 ( .A(_abc_15724_n1879), .B(_abc_15724_n1881), .Y(_abc_15724_n1882) );
  OR2X2 OR2X2_382 ( .A(_abc_15724_n1818_1), .B(_abc_15724_n1885_1), .Y(_abc_15724_n1886) );
  OR2X2 OR2X2_383 ( .A(_auto_iopadmap_cc_313_execute_26059_88_), .B(c_reg_24_), .Y(_abc_15724_n1889_1) );
  OR2X2 OR2X2_384 ( .A(_abc_15724_n1888), .B(_abc_15724_n1892), .Y(_abc_15724_n1893_1) );
  OR2X2 OR2X2_385 ( .A(_abc_15724_n1897_1), .B(_abc_15724_n1877), .Y(H2_reg_24__FF_INPUT) );
  OR2X2 OR2X2_386 ( .A(_auto_iopadmap_cc_313_execute_26059_89_), .B(c_reg_25_), .Y(_abc_15724_n1900) );
  OR2X2 OR2X2_387 ( .A(_abc_15724_n1903), .B(_abc_15724_n1890), .Y(_abc_15724_n1904) );
  OR2X2 OR2X2_388 ( .A(_abc_15724_n1894), .B(_abc_15724_n1904), .Y(_abc_15724_n1905_1) );
  OR2X2 OR2X2_389 ( .A(_abc_15724_n1913_1), .B(_abc_15724_n1899), .Y(H2_reg_25__FF_INPUT) );
  OR2X2 OR2X2_39 ( .A(_auto_iopadmap_cc_313_execute_26059_20_), .B(e_reg_20_), .Y(_abc_15724_n836) );
  OR2X2 OR2X2_390 ( .A(_auto_iopadmap_cc_313_execute_26059_90_), .B(c_reg_26_), .Y(_abc_15724_n1919) );
  OR2X2 OR2X2_391 ( .A(_abc_15724_n1918_1), .B(_abc_15724_n1922), .Y(_abc_15724_n1923_1) );
  OR2X2 OR2X2_392 ( .A(_abc_15724_n1927_1), .B(_abc_15724_n1915), .Y(H2_reg_26__FF_INPUT) );
  OR2X2 OR2X2_393 ( .A(_abc_15724_n1924), .B(_abc_15724_n1920), .Y(_abc_15724_n1929) );
  OR2X2 OR2X2_394 ( .A(_auto_iopadmap_cc_313_execute_26059_91_), .B(c_reg_27_), .Y(_abc_15724_n1930) );
  OR2X2 OR2X2_395 ( .A(_abc_15724_n1929), .B(_abc_15724_n1933), .Y(_abc_15724_n1934) );
  OR2X2 OR2X2_396 ( .A(_abc_15724_n1935_1), .B(_abc_15724_n1936), .Y(_abc_15724_n1937) );
  OR2X2 OR2X2_397 ( .A(_abc_15724_n851_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_91_), .Y(_abc_15724_n1940_1) );
  OR2X2 OR2X2_398 ( .A(_abc_15724_n1939), .B(_abc_15724_n1941), .Y(H2_reg_27__FF_INPUT) );
  OR2X2 OR2X2_399 ( .A(_abc_15724_n1943), .B(_abc_15724_n1931_1), .Y(_abc_15724_n1944_1) );
  OR2X2 OR2X2_4 ( .A(e_reg_18_), .B(_auto_iopadmap_cc_313_execute_26059_18_), .Y(_abc_15724_n711) );
  OR2X2 OR2X2_40 ( .A(_abc_15724_n839), .B(_abc_15724_n704), .Y(_abc_15724_n840_1) );
  OR2X2 OR2X2_400 ( .A(_abc_15724_n1916), .B(_abc_15724_n1947), .Y(_abc_15724_n1948_1) );
  OR2X2 OR2X2_401 ( .A(_abc_15724_n1887), .B(_abc_15724_n1951), .Y(_abc_15724_n1952) );
  OR2X2 OR2X2_402 ( .A(_auto_iopadmap_cc_313_execute_26059_92_), .B(c_reg_28_), .Y(_abc_15724_n1955) );
  OR2X2 OR2X2_403 ( .A(_abc_15724_n1954), .B(_abc_15724_n1958), .Y(_abc_15724_n1959) );
  OR2X2 OR2X2_404 ( .A(_abc_15724_n851_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_92_), .Y(_abc_15724_n1964) );
  OR2X2 OR2X2_405 ( .A(_abc_15724_n1963), .B(_abc_15724_n1965), .Y(H2_reg_28__FF_INPUT) );
  OR2X2 OR2X2_406 ( .A(_auto_iopadmap_cc_313_execute_26059_93_), .B(c_reg_29_), .Y(_abc_15724_n1969) );
  OR2X2 OR2X2_407 ( .A(_abc_15724_n1968), .B(_abc_15724_n1973), .Y(_abc_15724_n1974_1) );
  OR2X2 OR2X2_408 ( .A(_abc_15724_n1975), .B(_abc_15724_n1972), .Y(_abc_15724_n1976) );
  OR2X2 OR2X2_409 ( .A(_abc_15724_n1978), .B(_abc_15724_n1967), .Y(H2_reg_29__FF_INPUT) );
  OR2X2 OR2X2_41 ( .A(e_reg_22_), .B(_auto_iopadmap_cc_313_execute_26059_22_), .Y(_abc_15724_n841) );
  OR2X2 OR2X2_410 ( .A(_auto_iopadmap_cc_313_execute_26059_94_), .B(c_reg_30_), .Y(_abc_15724_n1983_1) );
  OR2X2 OR2X2_411 ( .A(_abc_15724_n1986), .B(_abc_15724_n1970_1), .Y(_abc_15724_n1987) );
  OR2X2 OR2X2_412 ( .A(_abc_15724_n1953_1), .B(_abc_15724_n1990), .Y(_abc_15724_n1991) );
  OR2X2 OR2X2_413 ( .A(_abc_15724_n1992), .B(_abc_15724_n1985), .Y(_abc_15724_n1993_1) );
  OR2X2 OR2X2_414 ( .A(_abc_15724_n1994), .B(_abc_15724_n1984), .Y(_abc_15724_n1995) );
  OR2X2 OR2X2_415 ( .A(_abc_15724_n1997), .B(_abc_15724_n1980), .Y(H2_reg_30__FF_INPUT) );
  OR2X2 OR2X2_416 ( .A(_abc_15724_n2001), .B(c_reg_31_), .Y(_abc_15724_n2002_1) );
  OR2X2 OR2X2_417 ( .A(_abc_15724_n2003), .B(_auto_iopadmap_cc_313_execute_26059_95_), .Y(_abc_15724_n2004) );
  OR2X2 OR2X2_418 ( .A(_abc_15724_n2000), .B(_abc_15724_n2006_1), .Y(_abc_15724_n2007) );
  OR2X2 OR2X2_419 ( .A(_abc_15724_n1999), .B(_abc_15724_n2005), .Y(_abc_15724_n2008) );
  OR2X2 OR2X2_42 ( .A(_abc_15724_n840_1), .B(_abc_15724_n844_1), .Y(_abc_15724_n845_1) );
  OR2X2 OR2X2_420 ( .A(_abc_15724_n851_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_95_), .Y(_abc_15724_n2011_1) );
  OR2X2 OR2X2_421 ( .A(_abc_15724_n2010), .B(_abc_15724_n2012), .Y(H2_reg_31__FF_INPUT) );
  OR2X2 OR2X2_422 ( .A(_auto_iopadmap_cc_313_execute_26059_96_), .B(b_reg_0_), .Y(_abc_15724_n2014) );
  OR2X2 OR2X2_423 ( .A(_abc_15724_n851_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_96_), .Y(_abc_15724_n2019) );
  OR2X2 OR2X2_424 ( .A(_abc_15724_n2018), .B(_abc_15724_n2020_1), .Y(H1_reg_0__FF_INPUT) );
  OR2X2 OR2X2_425 ( .A(_auto_iopadmap_cc_313_execute_26059_97_), .B(b_reg_1_), .Y(_abc_15724_n2022) );
  OR2X2 OR2X2_426 ( .A(_abc_15724_n2025), .B(_abc_15724_n2015), .Y(_abc_15724_n2026) );
  OR2X2 OR2X2_427 ( .A(_abc_15724_n2030), .B(_abc_15724_n2031), .Y(H1_reg_1__FF_INPUT) );
  OR2X2 OR2X2_428 ( .A(_auto_iopadmap_cc_313_execute_26059_98_), .B(b_reg_2_), .Y(_abc_15724_n2035) );
  OR2X2 OR2X2_429 ( .A(_abc_15724_n2034_1), .B(_abc_15724_n2038_1), .Y(_abc_15724_n2041) );
  OR2X2 OR2X2_43 ( .A(_abc_15724_n851_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_22_), .Y(_abc_15724_n852) );
  OR2X2 OR2X2_430 ( .A(_abc_15724_n2043_1), .B(_abc_15724_n2044), .Y(H1_reg_2__FF_INPUT) );
  OR2X2 OR2X2_431 ( .A(_abc_15724_n2039), .B(_abc_15724_n2036), .Y(_abc_15724_n2046) );
  OR2X2 OR2X2_432 ( .A(_auto_iopadmap_cc_313_execute_26059_99_), .B(b_reg_3_), .Y(_abc_15724_n2047) );
  OR2X2 OR2X2_433 ( .A(_abc_15724_n2046), .B(_abc_15724_n2050), .Y(_abc_15724_n2051) );
  OR2X2 OR2X2_434 ( .A(_abc_15724_n2052), .B(_abc_15724_n2053_1), .Y(_abc_15724_n2054) );
  OR2X2 OR2X2_435 ( .A(_abc_15724_n851_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_99_), .Y(_abc_15724_n2057_1) );
  OR2X2 OR2X2_436 ( .A(_abc_15724_n2056), .B(_abc_15724_n2058), .Y(H1_reg_3__FF_INPUT) );
  OR2X2 OR2X2_437 ( .A(_auto_iopadmap_cc_313_execute_26059_100_), .B(b_reg_4_), .Y(_abc_15724_n2060) );
  OR2X2 OR2X2_438 ( .A(_abc_15724_n2064), .B(_abc_15724_n2048_1), .Y(_abc_15724_n2065_1) );
  OR2X2 OR2X2_439 ( .A(_abc_15724_n2065_1), .B(_abc_15724_n2063), .Y(_abc_15724_n2068) );
  OR2X2 OR2X2_44 ( .A(_abc_15724_n849), .B(_abc_15724_n853_1), .Y(H4_reg_22__FF_INPUT) );
  OR2X2 OR2X2_440 ( .A(_abc_15724_n2070_1), .B(_abc_15724_n2071), .Y(H1_reg_4__FF_INPUT) );
  OR2X2 OR2X2_441 ( .A(_abc_15724_n2066), .B(_abc_15724_n2061_1), .Y(_abc_15724_n2074_1) );
  OR2X2 OR2X2_442 ( .A(_auto_iopadmap_cc_313_execute_26059_101_), .B(b_reg_5_), .Y(_abc_15724_n2075) );
  OR2X2 OR2X2_443 ( .A(_abc_15724_n2074_1), .B(_abc_15724_n2078), .Y(_abc_15724_n2081) );
  OR2X2 OR2X2_444 ( .A(_abc_15724_n2083_1), .B(_abc_15724_n2073), .Y(H1_reg_5__FF_INPUT) );
  OR2X2 OR2X2_445 ( .A(_abc_15724_n2079_1), .B(_abc_15724_n2076), .Y(_abc_15724_n2086) );
  OR2X2 OR2X2_446 ( .A(_auto_iopadmap_cc_313_execute_26059_102_), .B(b_reg_6_), .Y(_abc_15724_n2087) );
  OR2X2 OR2X2_447 ( .A(_abc_15724_n2086), .B(_abc_15724_n2090), .Y(_abc_15724_n2091) );
  OR2X2 OR2X2_448 ( .A(_abc_15724_n2095), .B(_abc_15724_n2085), .Y(H1_reg_6__FF_INPUT) );
  OR2X2 OR2X2_449 ( .A(_abc_15724_n851_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_103_), .Y(_abc_15724_n2097) );
  OR2X2 OR2X2_45 ( .A(_abc_15724_n846), .B(_abc_15724_n842), .Y(_abc_15724_n855_1) );
  OR2X2 OR2X2_450 ( .A(_abc_15724_n2097), .B(digest_update_bF_buf1), .Y(_abc_15724_n2098) );
  OR2X2 OR2X2_451 ( .A(_abc_15724_n2092_1), .B(_abc_15724_n2088_1), .Y(_abc_15724_n2099) );
  OR2X2 OR2X2_452 ( .A(_auto_iopadmap_cc_313_execute_26059_103_), .B(b_reg_7_), .Y(_abc_15724_n2101_1) );
  OR2X2 OR2X2_453 ( .A(_abc_15724_n2107), .B(_abc_15724_n850_bF_buf8), .Y(_abc_15724_n2108) );
  OR2X2 OR2X2_454 ( .A(_abc_15724_n2108), .B(_abc_15724_n2105_1), .Y(_abc_15724_n2109_1) );
  OR2X2 OR2X2_455 ( .A(_auto_iopadmap_cc_313_execute_26059_104_), .B(b_reg_8_), .Y(_abc_15724_n2111) );
  OR2X2 OR2X2_456 ( .A(_abc_15724_n2115), .B(_abc_15724_n2102), .Y(_abc_15724_n2116) );
  OR2X2 OR2X2_457 ( .A(_abc_15724_n2116), .B(_abc_15724_n2114_1), .Y(_abc_15724_n2117) );
  OR2X2 OR2X2_458 ( .A(_abc_15724_n851_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_104_), .Y(_abc_15724_n2122) );
  OR2X2 OR2X2_459 ( .A(_abc_15724_n2121), .B(_abc_15724_n2123_1), .Y(H1_reg_8__FF_INPUT) );
  OR2X2 OR2X2_46 ( .A(e_reg_23_), .B(_auto_iopadmap_cc_313_execute_26059_23_), .Y(_abc_15724_n856) );
  OR2X2 OR2X2_460 ( .A(_auto_iopadmap_cc_313_execute_26059_105_), .B(b_reg_9_), .Y(_abc_15724_n2127_1) );
  OR2X2 OR2X2_461 ( .A(_abc_15724_n2126), .B(_abc_15724_n2130), .Y(_abc_15724_n2131_1) );
  OR2X2 OR2X2_462 ( .A(_abc_15724_n2125), .B(_abc_15724_n2132), .Y(_abc_15724_n2133) );
  OR2X2 OR2X2_463 ( .A(_abc_15724_n851_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_105_), .Y(_abc_15724_n2136) );
  OR2X2 OR2X2_464 ( .A(_abc_15724_n2135_1), .B(_abc_15724_n2137), .Y(H1_reg_9__FF_INPUT) );
  OR2X2 OR2X2_465 ( .A(_abc_15724_n2132), .B(_abc_15724_n2113), .Y(_abc_15724_n2140) );
  OR2X2 OR2X2_466 ( .A(_abc_15724_n2144), .B(_abc_15724_n2142), .Y(_abc_15724_n2145) );
  OR2X2 OR2X2_467 ( .A(_auto_iopadmap_cc_313_execute_26059_106_), .B(b_reg_10_), .Y(_abc_15724_n2146) );
  OR2X2 OR2X2_468 ( .A(_abc_15724_n2145), .B(_abc_15724_n2149), .Y(_abc_15724_n2150) );
  OR2X2 OR2X2_469 ( .A(_abc_15724_n2154), .B(_abc_15724_n2139_1), .Y(H1_reg_10__FF_INPUT) );
  OR2X2 OR2X2_47 ( .A(_abc_15724_n855_1), .B(_abc_15724_n859), .Y(_abc_15724_n860) );
  OR2X2 OR2X2_470 ( .A(_auto_iopadmap_cc_313_execute_26059_107_), .B(b_reg_11_), .Y(_abc_15724_n2158) );
  OR2X2 OR2X2_471 ( .A(_abc_15724_n2157), .B(_abc_15724_n2161), .Y(_abc_15724_n2162) );
  OR2X2 OR2X2_472 ( .A(_abc_15724_n2156_1), .B(_abc_15724_n2163_1), .Y(_abc_15724_n2164) );
  OR2X2 OR2X2_473 ( .A(_abc_15724_n851_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_107_), .Y(_abc_15724_n2167) );
  OR2X2 OR2X2_474 ( .A(_abc_15724_n2166), .B(_abc_15724_n2168_1), .Y(H1_reg_11__FF_INPUT) );
  OR2X2 OR2X2_475 ( .A(_abc_15724_n2175), .B(_abc_15724_n2159), .Y(_abc_15724_n2176) );
  OR2X2 OR2X2_476 ( .A(_abc_15724_n2174), .B(_abc_15724_n2176), .Y(_abc_15724_n2177) );
  OR2X2 OR2X2_477 ( .A(_abc_15724_n2173), .B(_abc_15724_n2177), .Y(_abc_15724_n2178) );
  OR2X2 OR2X2_478 ( .A(_auto_iopadmap_cc_313_execute_26059_108_), .B(b_reg_12_), .Y(_abc_15724_n2179) );
  OR2X2 OR2X2_479 ( .A(_abc_15724_n2178), .B(_abc_15724_n2182_1), .Y(_abc_15724_n2183) );
  OR2X2 OR2X2_48 ( .A(_abc_15724_n861), .B(_abc_15724_n862), .Y(_abc_15724_n863_1) );
  OR2X2 OR2X2_480 ( .A(_abc_15724_n2187), .B(_abc_15724_n2170), .Y(H1_reg_12__FF_INPUT) );
  OR2X2 OR2X2_481 ( .A(_auto_iopadmap_cc_313_execute_26059_109_), .B(b_reg_13_), .Y(_abc_15724_n2191) );
  OR2X2 OR2X2_482 ( .A(_abc_15724_n2190), .B(_abc_15724_n2194), .Y(_abc_15724_n2195_1) );
  OR2X2 OR2X2_483 ( .A(_abc_15724_n2189), .B(_abc_15724_n2196), .Y(_abc_15724_n2197) );
  OR2X2 OR2X2_484 ( .A(_abc_15724_n851_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_109_), .Y(_abc_15724_n2200) );
  OR2X2 OR2X2_485 ( .A(_abc_15724_n2199), .B(_abc_15724_n2201), .Y(H1_reg_13__FF_INPUT) );
  OR2X2 OR2X2_486 ( .A(_abc_15724_n2196), .B(_abc_15724_n2181), .Y(_abc_15724_n2204) );
  OR2X2 OR2X2_487 ( .A(_abc_15724_n2208), .B(_abc_15724_n2206), .Y(_abc_15724_n2209) );
  OR2X2 OR2X2_488 ( .A(_auto_iopadmap_cc_313_execute_26059_110_), .B(b_reg_14_), .Y(_abc_15724_n2210) );
  OR2X2 OR2X2_489 ( .A(_abc_15724_n2209), .B(_abc_15724_n2213), .Y(_abc_15724_n2216) );
  OR2X2 OR2X2_49 ( .A(_abc_15724_n851_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_23_), .Y(_abc_15724_n866_1) );
  OR2X2 OR2X2_490 ( .A(_abc_15724_n2218), .B(_abc_15724_n2203), .Y(H1_reg_14__FF_INPUT) );
  OR2X2 OR2X2_491 ( .A(_auto_iopadmap_cc_313_execute_26059_111_), .B(b_reg_15_), .Y(_abc_15724_n2222) );
  OR2X2 OR2X2_492 ( .A(_abc_15724_n2221), .B(_abc_15724_n2225), .Y(_abc_15724_n2226) );
  OR2X2 OR2X2_493 ( .A(_abc_15724_n2220), .B(_abc_15724_n2227), .Y(_abc_15724_n2228) );
  OR2X2 OR2X2_494 ( .A(_abc_15724_n851_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_111_), .Y(_abc_15724_n2231) );
  OR2X2 OR2X2_495 ( .A(_abc_15724_n2230), .B(_abc_15724_n2232), .Y(H1_reg_15__FF_INPUT) );
  OR2X2 OR2X2_496 ( .A(_abc_15724_n2236), .B(_abc_15724_n2223), .Y(_abc_15724_n2237) );
  OR2X2 OR2X2_497 ( .A(_abc_15724_n2235), .B(_abc_15724_n2237), .Y(_abc_15724_n2238) );
  OR2X2 OR2X2_498 ( .A(_abc_15724_n2240), .B(_abc_15724_n2238), .Y(_abc_15724_n2241) );
  OR2X2 OR2X2_499 ( .A(_auto_iopadmap_cc_313_execute_26059_112_), .B(b_reg_16_), .Y(_abc_15724_n2242) );
  OR2X2 OR2X2_5 ( .A(_auto_iopadmap_cc_313_execute_26059_17_), .B(e_reg_17_), .Y(_abc_15724_n718_1) );
  OR2X2 OR2X2_50 ( .A(_abc_15724_n865), .B(_abc_15724_n867), .Y(H4_reg_23__FF_INPUT) );
  OR2X2 OR2X2_500 ( .A(_abc_15724_n2241), .B(_abc_15724_n2245), .Y(_abc_15724_n2246_1) );
  OR2X2 OR2X2_501 ( .A(_abc_15724_n851_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_112_), .Y(_abc_15724_n2251) );
  OR2X2 OR2X2_502 ( .A(_abc_15724_n2250_1), .B(_abc_15724_n2252), .Y(H1_reg_16__FF_INPUT) );
  OR2X2 OR2X2_503 ( .A(_auto_iopadmap_cc_313_execute_26059_113_), .B(b_reg_17_), .Y(_abc_15724_n2254) );
  OR2X2 OR2X2_504 ( .A(_abc_15724_n2259), .B(_abc_15724_n2257), .Y(_abc_15724_n2260) );
  OR2X2 OR2X2_505 ( .A(_abc_15724_n2264), .B(_abc_15724_n2265), .Y(H1_reg_17__FF_INPUT) );
  OR2X2 OR2X2_506 ( .A(_auto_iopadmap_cc_313_execute_26059_114_), .B(b_reg_18_), .Y(_abc_15724_n2269) );
  OR2X2 OR2X2_507 ( .A(_abc_15724_n2268), .B(_abc_15724_n2272), .Y(_abc_15724_n2273) );
  OR2X2 OR2X2_508 ( .A(_abc_15724_n851_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_114_), .Y(_abc_15724_n2278) );
  OR2X2 OR2X2_509 ( .A(_abc_15724_n2277), .B(_abc_15724_n2279), .Y(H1_reg_18__FF_INPUT) );
  OR2X2 OR2X2_51 ( .A(_abc_15724_n875_1), .B(_abc_15724_n857), .Y(_abc_15724_n876_1) );
  OR2X2 OR2X2_510 ( .A(_abc_15724_n2274), .B(_abc_15724_n2270), .Y(_abc_15724_n2281) );
  OR2X2 OR2X2_511 ( .A(_auto_iopadmap_cc_313_execute_26059_115_), .B(b_reg_19_), .Y(_abc_15724_n2282) );
  OR2X2 OR2X2_512 ( .A(_abc_15724_n2281), .B(_abc_15724_n2285), .Y(_abc_15724_n2286) );
  OR2X2 OR2X2_513 ( .A(_abc_15724_n2287_1), .B(_abc_15724_n2288), .Y(_abc_15724_n2289) );
  OR2X2 OR2X2_514 ( .A(_abc_15724_n851_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_115_), .Y(_abc_15724_n2292) );
  OR2X2 OR2X2_515 ( .A(_abc_15724_n2291_1), .B(_abc_15724_n2293), .Y(H1_reg_19__FF_INPUT) );
  OR2X2 OR2X2_516 ( .A(_abc_15724_n2296), .B(_abc_15724_n2255), .Y(_abc_15724_n2297) );
  OR2X2 OR2X2_517 ( .A(_abc_15724_n2300), .B(_abc_15724_n2283), .Y(_abc_15724_n2301) );
  OR2X2 OR2X2_518 ( .A(_abc_15724_n2299), .B(_abc_15724_n2301), .Y(_abc_15724_n2302) );
  OR2X2 OR2X2_519 ( .A(_abc_15724_n2305), .B(_abc_15724_n2302), .Y(_abc_15724_n2306) );
  OR2X2 OR2X2_52 ( .A(_abc_15724_n874), .B(_abc_15724_n876_1), .Y(_abc_15724_n877) );
  OR2X2 OR2X2_520 ( .A(_auto_iopadmap_cc_313_execute_26059_116_), .B(b_reg_20_), .Y(_abc_15724_n2307) );
  OR2X2 OR2X2_521 ( .A(_abc_15724_n2306), .B(_abc_15724_n2310), .Y(_abc_15724_n2311) );
  OR2X2 OR2X2_522 ( .A(_abc_15724_n2315), .B(_abc_15724_n2295), .Y(H1_reg_20__FF_INPUT) );
  OR2X2 OR2X2_523 ( .A(_auto_iopadmap_cc_313_execute_26059_117_), .B(b_reg_21_), .Y(_abc_15724_n2318) );
  OR2X2 OR2X2_524 ( .A(_abc_15724_n2312), .B(_abc_15724_n2308), .Y(_abc_15724_n2322) );
  OR2X2 OR2X2_525 ( .A(_abc_15724_n2322), .B(_abc_15724_n2321), .Y(_abc_15724_n2323) );
  OR2X2 OR2X2_526 ( .A(_abc_15724_n2327), .B(_abc_15724_n2317), .Y(H1_reg_21__FF_INPUT) );
  OR2X2 OR2X2_527 ( .A(_abc_15724_n2324), .B(_abc_15724_n2319), .Y(_abc_15724_n2329) );
  OR2X2 OR2X2_528 ( .A(_auto_iopadmap_cc_313_execute_26059_118_), .B(b_reg_22_), .Y(_abc_15724_n2330_1) );
  OR2X2 OR2X2_529 ( .A(_abc_15724_n2329), .B(_abc_15724_n2333), .Y(_abc_15724_n2334) );
  OR2X2 OR2X2_53 ( .A(_abc_15724_n873), .B(_abc_15724_n877), .Y(_abc_15724_n878_1) );
  OR2X2 OR2X2_530 ( .A(_abc_15724_n851_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_118_), .Y(_abc_15724_n2339) );
  OR2X2 OR2X2_531 ( .A(_abc_15724_n2338), .B(_abc_15724_n2340), .Y(H1_reg_22__FF_INPUT) );
  OR2X2 OR2X2_532 ( .A(_abc_15724_n2335), .B(_abc_15724_n2331), .Y(_abc_15724_n2342) );
  OR2X2 OR2X2_533 ( .A(_auto_iopadmap_cc_313_execute_26059_119_), .B(b_reg_23_), .Y(_abc_15724_n2344) );
  OR2X2 OR2X2_534 ( .A(_abc_15724_n2348), .B(_abc_15724_n2350), .Y(_abc_15724_n2351) );
  OR2X2 OR2X2_535 ( .A(_abc_15724_n851_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_119_), .Y(_abc_15724_n2353) );
  OR2X2 OR2X2_536 ( .A(_abc_15724_n2352), .B(_abc_15724_n2354), .Y(H1_reg_23__FF_INPUT) );
  OR2X2 OR2X2_537 ( .A(_abc_15724_n2362), .B(_abc_15724_n2345), .Y(_abc_15724_n2363) );
  OR2X2 OR2X2_538 ( .A(_abc_15724_n2364), .B(_abc_15724_n2319), .Y(_abc_15724_n2365) );
  OR2X2 OR2X2_539 ( .A(_abc_15724_n2366_1), .B(_abc_15724_n2363), .Y(_abc_15724_n2367) );
  OR2X2 OR2X2_54 ( .A(_abc_15724_n872), .B(_abc_15724_n878_1), .Y(_abc_15724_n879) );
  OR2X2 OR2X2_540 ( .A(_abc_15724_n2361), .B(_abc_15724_n2367), .Y(_abc_15724_n2368) );
  OR2X2 OR2X2_541 ( .A(_abc_15724_n2360), .B(_abc_15724_n2368), .Y(_abc_15724_n2369) );
  OR2X2 OR2X2_542 ( .A(_auto_iopadmap_cc_313_execute_26059_120_), .B(b_reg_24_), .Y(_abc_15724_n2370_1) );
  OR2X2 OR2X2_543 ( .A(_abc_15724_n2369), .B(_abc_15724_n2373), .Y(_abc_15724_n2374) );
  OR2X2 OR2X2_544 ( .A(_abc_15724_n851_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_120_), .Y(_abc_15724_n2379) );
  OR2X2 OR2X2_545 ( .A(_abc_15724_n2378), .B(_abc_15724_n2380), .Y(H1_reg_24__FF_INPUT) );
  OR2X2 OR2X2_546 ( .A(_auto_iopadmap_cc_313_execute_26059_121_), .B(b_reg_25_), .Y(_abc_15724_n2384) );
  OR2X2 OR2X2_547 ( .A(_abc_15724_n2383), .B(_abc_15724_n2387), .Y(_abc_15724_n2388) );
  OR2X2 OR2X2_548 ( .A(_abc_15724_n2382), .B(_abc_15724_n2389), .Y(_abc_15724_n2390) );
  OR2X2 OR2X2_549 ( .A(_abc_15724_n851_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_121_), .Y(_abc_15724_n2393) );
  OR2X2 OR2X2_55 ( .A(e_reg_24_), .B(_auto_iopadmap_cc_313_execute_26059_24_), .Y(_abc_15724_n880) );
  OR2X2 OR2X2_550 ( .A(_abc_15724_n2392), .B(_abc_15724_n2394), .Y(H1_reg_25__FF_INPUT) );
  OR2X2 OR2X2_551 ( .A(_abc_15724_n2398), .B(_abc_15724_n2385), .Y(_abc_15724_n2399) );
  OR2X2 OR2X2_552 ( .A(_abc_15724_n2397), .B(_abc_15724_n2399), .Y(_abc_15724_n2400) );
  OR2X2 OR2X2_553 ( .A(_auto_iopadmap_cc_313_execute_26059_122_), .B(b_reg_26_), .Y(_abc_15724_n2401) );
  OR2X2 OR2X2_554 ( .A(_abc_15724_n2400), .B(_abc_15724_n2404), .Y(_abc_15724_n2405) );
  OR2X2 OR2X2_555 ( .A(_abc_15724_n851_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_122_), .Y(_abc_15724_n2410) );
  OR2X2 OR2X2_556 ( .A(_abc_15724_n2409), .B(_abc_15724_n2411), .Y(H1_reg_26__FF_INPUT) );
  OR2X2 OR2X2_557 ( .A(_auto_iopadmap_cc_313_execute_26059_123_), .B(b_reg_27_), .Y(_abc_15724_n2415) );
  OR2X2 OR2X2_558 ( .A(_abc_15724_n2414), .B(_abc_15724_n2418), .Y(_abc_15724_n2419) );
  OR2X2 OR2X2_559 ( .A(_abc_15724_n2413), .B(_abc_15724_n2420), .Y(_abc_15724_n2421) );
  OR2X2 OR2X2_56 ( .A(_abc_15724_n879), .B(_abc_15724_n883), .Y(_abc_15724_n884_1) );
  OR2X2 OR2X2_560 ( .A(_abc_15724_n851_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_123_), .Y(_abc_15724_n2424) );
  OR2X2 OR2X2_561 ( .A(_abc_15724_n2423), .B(_abc_15724_n2425), .Y(H1_reg_27__FF_INPUT) );
  OR2X2 OR2X2_562 ( .A(_abc_15724_n2428), .B(_abc_15724_n2416), .Y(_abc_15724_n2429) );
  OR2X2 OR2X2_563 ( .A(_abc_15724_n2431), .B(_abc_15724_n2429), .Y(_abc_15724_n2432) );
  OR2X2 OR2X2_564 ( .A(_abc_15724_n2434), .B(_abc_15724_n2432), .Y(_abc_15724_n2435) );
  OR2X2 OR2X2_565 ( .A(_auto_iopadmap_cc_313_execute_26059_124_), .B(b_reg_28_), .Y(_abc_15724_n2436) );
  OR2X2 OR2X2_566 ( .A(_abc_15724_n2435), .B(_abc_15724_n2439), .Y(_abc_15724_n2440) );
  OR2X2 OR2X2_567 ( .A(_abc_15724_n2444), .B(_abc_15724_n2427), .Y(H1_reg_28__FF_INPUT) );
  OR2X2 OR2X2_568 ( .A(_auto_iopadmap_cc_313_execute_26059_125_), .B(b_reg_29_), .Y(_abc_15724_n2447) );
  OR2X2 OR2X2_569 ( .A(_abc_15724_n2454), .B(_abc_15724_n2451), .Y(_abc_15724_n2455) );
  OR2X2 OR2X2_57 ( .A(_abc_15724_n851_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_24_), .Y(_abc_15724_n889) );
  OR2X2 OR2X2_570 ( .A(_abc_15724_n851_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_125_), .Y(_abc_15724_n2457) );
  OR2X2 OR2X2_571 ( .A(_abc_15724_n2456), .B(_abc_15724_n2458), .Y(H1_reg_29__FF_INPUT) );
  OR2X2 OR2X2_572 ( .A(_auto_iopadmap_cc_313_execute_26059_126_), .B(b_reg_30_), .Y(_abc_15724_n2460) );
  OR2X2 OR2X2_573 ( .A(_abc_15724_n2464), .B(_abc_15724_n2448), .Y(_abc_15724_n2465) );
  OR2X2 OR2X2_574 ( .A(_abc_15724_n2467), .B(_abc_15724_n2465), .Y(_abc_15724_n2468) );
  OR2X2 OR2X2_575 ( .A(_abc_15724_n2468), .B(_abc_15724_n2463), .Y(_abc_15724_n2469) );
  OR2X2 OR2X2_576 ( .A(_abc_15724_n851_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_126_), .Y(_abc_15724_n2474) );
  OR2X2 OR2X2_577 ( .A(_abc_15724_n2473), .B(_abc_15724_n2475), .Y(H1_reg_30__FF_INPUT) );
  OR2X2 OR2X2_578 ( .A(_abc_15724_n2470), .B(_abc_15724_n2461), .Y(_abc_15724_n2477) );
  OR2X2 OR2X2_579 ( .A(_abc_15724_n2478), .B(b_reg_31_), .Y(_abc_15724_n2479) );
  OR2X2 OR2X2_58 ( .A(_abc_15724_n888), .B(_abc_15724_n890), .Y(H4_reg_24__FF_INPUT) );
  OR2X2 OR2X2_580 ( .A(_abc_15724_n2480), .B(_auto_iopadmap_cc_313_execute_26059_127_), .Y(_abc_15724_n2481) );
  OR2X2 OR2X2_581 ( .A(_abc_15724_n2477), .B(_abc_15724_n2483), .Y(_abc_15724_n2484_1) );
  OR2X2 OR2X2_582 ( .A(_abc_15724_n2485), .B(_abc_15724_n2482), .Y(_abc_15724_n2486) );
  OR2X2 OR2X2_583 ( .A(_abc_15724_n851_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_127_), .Y(_abc_15724_n2489) );
  OR2X2 OR2X2_584 ( .A(_abc_15724_n2488_1), .B(_abc_15724_n2490), .Y(H1_reg_31__FF_INPUT) );
  OR2X2 OR2X2_585 ( .A(_auto_iopadmap_cc_313_execute_26059_128_), .B(a_reg_0_), .Y(_abc_15724_n2492) );
  OR2X2 OR2X2_586 ( .A(_abc_15724_n851_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_128_), .Y(_abc_15724_n2497) );
  OR2X2 OR2X2_587 ( .A(_abc_15724_n2496), .B(_abc_15724_n2498), .Y(H0_reg_0__FF_INPUT) );
  OR2X2 OR2X2_588 ( .A(_auto_iopadmap_cc_313_execute_26059_129_), .B(a_reg_1_), .Y(_abc_15724_n2500) );
  OR2X2 OR2X2_589 ( .A(_abc_15724_n2503), .B(_abc_15724_n2493), .Y(_abc_15724_n2504) );
  OR2X2 OR2X2_59 ( .A(e_reg_25_), .B(_auto_iopadmap_cc_313_execute_26059_25_), .Y(_abc_15724_n894) );
  OR2X2 OR2X2_590 ( .A(_abc_15724_n2508), .B(_abc_15724_n2509), .Y(H0_reg_1__FF_INPUT) );
  OR2X2 OR2X2_591 ( .A(_auto_iopadmap_cc_313_execute_26059_130_), .B(a_reg_2_), .Y(_abc_15724_n2512) );
  OR2X2 OR2X2_592 ( .A(_abc_15724_n2511), .B(_abc_15724_n2516), .Y(_abc_15724_n2517) );
  OR2X2 OR2X2_593 ( .A(_abc_15724_n2518), .B(_abc_15724_n2515), .Y(_abc_15724_n2519) );
  OR2X2 OR2X2_594 ( .A(_abc_15724_n2521), .B(_abc_15724_n2522), .Y(H0_reg_2__FF_INPUT) );
  OR2X2 OR2X2_595 ( .A(_auto_iopadmap_cc_313_execute_26059_131_), .B(a_reg_3_), .Y(_abc_15724_n2526) );
  OR2X2 OR2X2_596 ( .A(_abc_15724_n2525), .B(_abc_15724_n2529), .Y(_abc_15724_n2530) );
  OR2X2 OR2X2_597 ( .A(_abc_15724_n2524_1), .B(_abc_15724_n2531), .Y(_abc_15724_n2532) );
  OR2X2 OR2X2_598 ( .A(_abc_15724_n2534), .B(_abc_15724_n2535), .Y(H0_reg_3__FF_INPUT) );
  OR2X2 OR2X2_599 ( .A(_auto_iopadmap_cc_313_execute_26059_132_), .B(a_reg_4_), .Y(_abc_15724_n2537) );
  OR2X2 OR2X2_6 ( .A(_abc_15724_n720), .B(_abc_15724_n717), .Y(_abc_15724_n721_1) );
  OR2X2 OR2X2_60 ( .A(_abc_15724_n893), .B(_abc_15724_n897_1), .Y(_abc_15724_n898_1) );
  OR2X2 OR2X2_600 ( .A(_abc_15724_n2524_1), .B(_abc_15724_n2542), .Y(_abc_15724_n2543) );
  OR2X2 OR2X2_601 ( .A(_abc_15724_n2544), .B(_abc_15724_n2541), .Y(_abc_15724_n2545) );
  OR2X2 OR2X2_602 ( .A(_abc_15724_n2546), .B(_abc_15724_n2540), .Y(_abc_15724_n2547) );
  OR2X2 OR2X2_603 ( .A(_abc_15724_n2549), .B(_abc_15724_n2550), .Y(H0_reg_4__FF_INPUT) );
  OR2X2 OR2X2_604 ( .A(_auto_iopadmap_cc_313_execute_26059_133_), .B(a_reg_5_), .Y(_abc_15724_n2554) );
  OR2X2 OR2X2_605 ( .A(_abc_15724_n2553), .B(_abc_15724_n2558), .Y(_abc_15724_n2559) );
  OR2X2 OR2X2_606 ( .A(_abc_15724_n2560), .B(_abc_15724_n2557), .Y(_abc_15724_n2561) );
  OR2X2 OR2X2_607 ( .A(_abc_15724_n2563), .B(_abc_15724_n2552), .Y(H0_reg_5__FF_INPUT) );
  OR2X2 OR2X2_608 ( .A(_auto_iopadmap_cc_313_execute_26059_134_), .B(a_reg_6_), .Y(_abc_15724_n2568) );
  OR2X2 OR2X2_609 ( .A(_abc_15724_n2567), .B(_abc_15724_n2571), .Y(_abc_15724_n2572) );
  OR2X2 OR2X2_61 ( .A(_abc_15724_n892), .B(_abc_15724_n899_1), .Y(_abc_15724_n900) );
  OR2X2 OR2X2_610 ( .A(_abc_15724_n2566), .B(_abc_15724_n2573_1), .Y(_abc_15724_n2574) );
  OR2X2 OR2X2_611 ( .A(_abc_15724_n2576), .B(_abc_15724_n2565), .Y(H0_reg_6__FF_INPUT) );
  OR2X2 OR2X2_612 ( .A(_auto_iopadmap_cc_313_execute_26059_135_), .B(a_reg_7_), .Y(_abc_15724_n2580) );
  OR2X2 OR2X2_613 ( .A(_abc_15724_n2583), .B(_abc_15724_n2569), .Y(_abc_15724_n2584) );
  OR2X2 OR2X2_614 ( .A(_abc_15724_n2579), .B(_abc_15724_n2584), .Y(_abc_15724_n2585) );
  OR2X2 OR2X2_615 ( .A(_abc_15724_n2574), .B(_abc_15724_n2586), .Y(_abc_15724_n2587) );
  OR2X2 OR2X2_616 ( .A(_abc_15724_n2592), .B(_abc_15724_n2578), .Y(H0_reg_7__FF_INPUT) );
  OR2X2 OR2X2_617 ( .A(_auto_iopadmap_cc_313_execute_26059_136_), .B(a_reg_8_), .Y(_abc_15724_n2597) );
  OR2X2 OR2X2_618 ( .A(_abc_15724_n2596), .B(_abc_15724_n2600), .Y(_abc_15724_n2601) );
  OR2X2 OR2X2_619 ( .A(_abc_15724_n851_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_136_), .Y(_abc_15724_n2606) );
  OR2X2 OR2X2_62 ( .A(_abc_15724_n851_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_25_), .Y(_abc_15724_n903) );
  OR2X2 OR2X2_620 ( .A(_abc_15724_n2605), .B(_abc_15724_n2607_1), .Y(H0_reg_8__FF_INPUT) );
  OR2X2 OR2X2_621 ( .A(_auto_iopadmap_cc_313_execute_26059_137_), .B(a_reg_9_), .Y(_abc_15724_n2611) );
  OR2X2 OR2X2_622 ( .A(_abc_15724_n2610), .B(_abc_15724_n2614), .Y(_abc_15724_n2615) );
  OR2X2 OR2X2_623 ( .A(_abc_15724_n2609), .B(_abc_15724_n2616), .Y(_abc_15724_n2617) );
  OR2X2 OR2X2_624 ( .A(_abc_15724_n851_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_137_), .Y(_abc_15724_n2620) );
  OR2X2 OR2X2_625 ( .A(_abc_15724_n2619), .B(_abc_15724_n2621), .Y(H0_reg_9__FF_INPUT) );
  OR2X2 OR2X2_626 ( .A(_auto_iopadmap_cc_313_execute_26059_138_), .B(a_reg_10_), .Y(_abc_15724_n2624) );
  OR2X2 OR2X2_627 ( .A(_abc_15724_n2616), .B(_abc_15724_n2599), .Y(_abc_15724_n2628) );
  OR2X2 OR2X2_628 ( .A(_abc_15724_n2632), .B(_abc_15724_n2630), .Y(_abc_15724_n2633) );
  OR2X2 OR2X2_629 ( .A(_abc_15724_n2633), .B(_abc_15724_n2627), .Y(_abc_15724_n2634) );
  OR2X2 OR2X2_63 ( .A(_abc_15724_n902), .B(_abc_15724_n904), .Y(H4_reg_25__FF_INPUT) );
  OR2X2 OR2X2_630 ( .A(_abc_15724_n2638), .B(_abc_15724_n2623), .Y(H0_reg_10__FF_INPUT) );
  OR2X2 OR2X2_631 ( .A(_auto_iopadmap_cc_313_execute_26059_139_), .B(a_reg_11_), .Y(_abc_15724_n2641) );
  OR2X2 OR2X2_632 ( .A(_abc_15724_n2648_1), .B(_abc_15724_n2645), .Y(_abc_15724_n2649) );
  OR2X2 OR2X2_633 ( .A(_abc_15724_n2650), .B(_abc_15724_n2651), .Y(H0_reg_11__FF_INPUT) );
  OR2X2 OR2X2_634 ( .A(_abc_15724_n2595), .B(_abc_15724_n2656), .Y(_abc_15724_n2657) );
  OR2X2 OR2X2_635 ( .A(_abc_15724_n2659), .B(_abc_15724_n2642), .Y(_abc_15724_n2660) );
  OR2X2 OR2X2_636 ( .A(_abc_15724_n2658), .B(_abc_15724_n2660), .Y(_abc_15724_n2661) );
  OR2X2 OR2X2_637 ( .A(_auto_iopadmap_cc_313_execute_26059_140_), .B(a_reg_12_), .Y(_abc_15724_n2665) );
  OR2X2 OR2X2_638 ( .A(_abc_15724_n2664), .B(_abc_15724_n2668), .Y(_abc_15724_n2669) );
  OR2X2 OR2X2_639 ( .A(_abc_15724_n2673), .B(_abc_15724_n2653), .Y(H0_reg_12__FF_INPUT) );
  OR2X2 OR2X2_64 ( .A(_abc_15724_n911), .B(_abc_15724_n895), .Y(_abc_15724_n912) );
  OR2X2 OR2X2_640 ( .A(_auto_iopadmap_cc_313_execute_26059_141_), .B(a_reg_13_), .Y(_abc_15724_n2677) );
  OR2X2 OR2X2_641 ( .A(_abc_15724_n2676), .B(_abc_15724_n2680), .Y(_abc_15724_n2681) );
  OR2X2 OR2X2_642 ( .A(_abc_15724_n2675), .B(_abc_15724_n2682), .Y(_abc_15724_n2683) );
  OR2X2 OR2X2_643 ( .A(_abc_15724_n851_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_141_), .Y(_abc_15724_n2686) );
  OR2X2 OR2X2_644 ( .A(_abc_15724_n2685), .B(_abc_15724_n2687_1), .Y(H0_reg_13__FF_INPUT) );
  OR2X2 OR2X2_645 ( .A(_auto_iopadmap_cc_313_execute_26059_142_), .B(a_reg_14_), .Y(_abc_15724_n2690) );
  OR2X2 OR2X2_646 ( .A(_abc_15724_n2696), .B(_abc_15724_n2694), .Y(_abc_15724_n2697) );
  OR2X2 OR2X2_647 ( .A(_abc_15724_n2698), .B(_abc_15724_n2693), .Y(_abc_15724_n2701) );
  OR2X2 OR2X2_648 ( .A(_abc_15724_n2703), .B(_abc_15724_n2689), .Y(H0_reg_14__FF_INPUT) );
  OR2X2 OR2X2_649 ( .A(_auto_iopadmap_cc_313_execute_26059_143_), .B(a_reg_15_), .Y(_abc_15724_n2706) );
  OR2X2 OR2X2_65 ( .A(_abc_15724_n910), .B(_abc_15724_n912), .Y(_abc_15724_n913) );
  OR2X2 OR2X2_650 ( .A(_abc_15724_n2705), .B(_abc_15724_n2710), .Y(_abc_15724_n2711) );
  OR2X2 OR2X2_651 ( .A(_abc_15724_n2712), .B(_abc_15724_n2709), .Y(_abc_15724_n2713) );
  OR2X2 OR2X2_652 ( .A(_abc_15724_n2715), .B(_abc_15724_n2716), .Y(H0_reg_15__FF_INPUT) );
  OR2X2 OR2X2_653 ( .A(_abc_15724_n2718), .B(_abc_15724_n2707), .Y(_abc_15724_n2719) );
  OR2X2 OR2X2_654 ( .A(_abc_15724_n2695), .B(_abc_15724_n2694), .Y(_abc_15724_n2721) );
  OR2X2 OR2X2_655 ( .A(_abc_15724_n2723), .B(_abc_15724_n2721), .Y(_abc_15724_n2724) );
  OR2X2 OR2X2_656 ( .A(_abc_15724_n2663), .B(_abc_15724_n2728), .Y(_abc_15724_n2729) );
  OR2X2 OR2X2_657 ( .A(_auto_iopadmap_cc_313_execute_26059_144_), .B(a_reg_16_), .Y(_abc_15724_n2732) );
  OR2X2 OR2X2_658 ( .A(_abc_15724_n2731_1), .B(_abc_15724_n2735), .Y(_abc_15724_n2736) );
  OR2X2 OR2X2_659 ( .A(_abc_15724_n851_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_144_), .Y(_abc_15724_n2741) );
  OR2X2 OR2X2_66 ( .A(_auto_iopadmap_cc_313_execute_26059_26_), .B(e_reg_26_), .Y(_abc_15724_n914) );
  OR2X2 OR2X2_660 ( .A(_abc_15724_n2740), .B(_abc_15724_n2742), .Y(H0_reg_16__FF_INPUT) );
  OR2X2 OR2X2_661 ( .A(_auto_iopadmap_cc_313_execute_26059_145_), .B(a_reg_17_), .Y(_abc_15724_n2744) );
  OR2X2 OR2X2_662 ( .A(_abc_15724_n2749), .B(_abc_15724_n2747), .Y(_abc_15724_n2750) );
  OR2X2 OR2X2_663 ( .A(_abc_15724_n2754), .B(_abc_15724_n2755), .Y(H0_reg_17__FF_INPUT) );
  OR2X2 OR2X2_664 ( .A(_auto_iopadmap_cc_313_execute_26059_146_), .B(a_reg_18_), .Y(_abc_15724_n2759) );
  OR2X2 OR2X2_665 ( .A(_abc_15724_n2758), .B(_abc_15724_n2762), .Y(_abc_15724_n2763) );
  OR2X2 OR2X2_666 ( .A(_abc_15724_n851_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_146_), .Y(_abc_15724_n2768_1) );
  OR2X2 OR2X2_667 ( .A(_abc_15724_n2767), .B(_abc_15724_n2769), .Y(H0_reg_18__FF_INPUT) );
  OR2X2 OR2X2_668 ( .A(_auto_iopadmap_cc_313_execute_26059_147_), .B(a_reg_19_), .Y(_abc_15724_n2772_1) );
  OR2X2 OR2X2_669 ( .A(_abc_15724_n2779), .B(_abc_15724_n2776), .Y(_abc_15724_n2780) );
  OR2X2 OR2X2_67 ( .A(_abc_15724_n913), .B(_abc_15724_n917), .Y(_abc_15724_n918) );
  OR2X2 OR2X2_670 ( .A(_abc_15724_n2781), .B(_abc_15724_n2782), .Y(H0_reg_19__FF_INPUT) );
  OR2X2 OR2X2_671 ( .A(_abc_15724_n2730), .B(_abc_15724_n2788), .Y(_abc_15724_n2789) );
  OR2X2 OR2X2_672 ( .A(_abc_15724_n2790), .B(_abc_15724_n2745), .Y(_abc_15724_n2791) );
  OR2X2 OR2X2_673 ( .A(_abc_15724_n2793), .B(_abc_15724_n2773), .Y(_abc_15724_n2794) );
  OR2X2 OR2X2_674 ( .A(_abc_15724_n2792), .B(_abc_15724_n2794), .Y(_abc_15724_n2795) );
  OR2X2 OR2X2_675 ( .A(_auto_iopadmap_cc_313_execute_26059_148_), .B(a_reg_20_), .Y(_abc_15724_n2799) );
  OR2X2 OR2X2_676 ( .A(_abc_15724_n2798), .B(_abc_15724_n2802), .Y(_abc_15724_n2803) );
  OR2X2 OR2X2_677 ( .A(_abc_15724_n2807), .B(_abc_15724_n2784), .Y(H0_reg_20__FF_INPUT) );
  OR2X2 OR2X2_678 ( .A(_auto_iopadmap_cc_313_execute_26059_149_), .B(a_reg_21_), .Y(_abc_15724_n2809) );
  OR2X2 OR2X2_679 ( .A(_abc_15724_n2814), .B(_abc_15724_n2812_1), .Y(_abc_15724_n2815) );
  OR2X2 OR2X2_68 ( .A(_abc_15724_n922_1), .B(_abc_15724_n908_1), .Y(H4_reg_26__FF_INPUT) );
  OR2X2 OR2X2_680 ( .A(_abc_15724_n2819), .B(_abc_15724_n2820), .Y(H0_reg_21__FF_INPUT) );
  OR2X2 OR2X2_681 ( .A(_abc_15724_n2816), .B(_abc_15724_n2810), .Y(_abc_15724_n2822) );
  OR2X2 OR2X2_682 ( .A(_auto_iopadmap_cc_313_execute_26059_150_), .B(a_reg_22_), .Y(_abc_15724_n2823) );
  OR2X2 OR2X2_683 ( .A(_abc_15724_n2822), .B(_abc_15724_n2826), .Y(_abc_15724_n2827) );
  OR2X2 OR2X2_684 ( .A(_abc_15724_n851_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_150_), .Y(_abc_15724_n2832) );
  OR2X2 OR2X2_685 ( .A(_abc_15724_n2831), .B(_abc_15724_n2833), .Y(H0_reg_22__FF_INPUT) );
  OR2X2 OR2X2_686 ( .A(_abc_15724_n2828), .B(_abc_15724_n2824), .Y(_abc_15724_n2835) );
  OR2X2 OR2X2_687 ( .A(_auto_iopadmap_cc_313_execute_26059_151_), .B(a_reg_23_), .Y(_abc_15724_n2837) );
  OR2X2 OR2X2_688 ( .A(_abc_15724_n2841), .B(_abc_15724_n2843), .Y(_abc_15724_n2844) );
  OR2X2 OR2X2_689 ( .A(_abc_15724_n2845_1), .B(_abc_15724_n2846), .Y(H0_reg_23__FF_INPUT) );
  OR2X2 OR2X2_69 ( .A(_auto_iopadmap_cc_313_execute_26059_27_), .B(e_reg_27_), .Y(_abc_15724_n925) );
  OR2X2 OR2X2_690 ( .A(_abc_15724_n2848_1), .B(_abc_15724_n2810), .Y(_abc_15724_n2849) );
  OR2X2 OR2X2_691 ( .A(_abc_15724_n2852), .B(_abc_15724_n2838), .Y(_abc_15724_n2853) );
  OR2X2 OR2X2_692 ( .A(_abc_15724_n2851), .B(_abc_15724_n2853), .Y(_abc_15724_n2854) );
  OR2X2 OR2X2_693 ( .A(_abc_15724_n2797), .B(_abc_15724_n2858), .Y(_abc_15724_n2859) );
  OR2X2 OR2X2_694 ( .A(_auto_iopadmap_cc_313_execute_26059_152_), .B(a_reg_24_), .Y(_abc_15724_n2862) );
  OR2X2 OR2X2_695 ( .A(_abc_15724_n2861), .B(_abc_15724_n2865), .Y(_abc_15724_n2866) );
  OR2X2 OR2X2_696 ( .A(_abc_15724_n851_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_152_), .Y(_abc_15724_n2871) );
  OR2X2 OR2X2_697 ( .A(_abc_15724_n2870), .B(_abc_15724_n2872), .Y(H0_reg_24__FF_INPUT) );
  OR2X2 OR2X2_698 ( .A(_auto_iopadmap_cc_313_execute_26059_153_), .B(a_reg_25_), .Y(_abc_15724_n2876) );
  OR2X2 OR2X2_699 ( .A(_abc_15724_n2875), .B(_abc_15724_n2879), .Y(_abc_15724_n2880) );
  OR2X2 OR2X2_7 ( .A(_abc_15724_n725), .B(_abc_15724_n705), .Y(_abc_15724_n726) );
  OR2X2 OR2X2_70 ( .A(_abc_15724_n928), .B(_abc_15724_n915), .Y(_abc_15724_n929) );
  OR2X2 OR2X2_700 ( .A(_abc_15724_n2874), .B(_abc_15724_n2881), .Y(_abc_15724_n2882) );
  OR2X2 OR2X2_701 ( .A(_abc_15724_n851_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_153_), .Y(_abc_15724_n2885) );
  OR2X2 OR2X2_702 ( .A(_abc_15724_n2884), .B(_abc_15724_n2886), .Y(H0_reg_25__FF_INPUT) );
  OR2X2 OR2X2_703 ( .A(_abc_15724_n2890_1), .B(_abc_15724_n2877), .Y(_abc_15724_n2891) );
  OR2X2 OR2X2_704 ( .A(_abc_15724_n2889), .B(_abc_15724_n2891), .Y(_abc_15724_n2892) );
  OR2X2 OR2X2_705 ( .A(_auto_iopadmap_cc_313_execute_26059_154_), .B(a_reg_26_), .Y(_abc_15724_n2893) );
  OR2X2 OR2X2_706 ( .A(_abc_15724_n2892), .B(_abc_15724_n2896), .Y(_abc_15724_n2897) );
  OR2X2 OR2X2_707 ( .A(_abc_15724_n851_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_154_), .Y(_abc_15724_n2902) );
  OR2X2 OR2X2_708 ( .A(_abc_15724_n2901), .B(_abc_15724_n2903), .Y(H0_reg_26__FF_INPUT) );
  OR2X2 OR2X2_709 ( .A(_auto_iopadmap_cc_313_execute_26059_155_), .B(a_reg_27_), .Y(_abc_15724_n2906) );
  OR2X2 OR2X2_71 ( .A(_abc_15724_n919), .B(_abc_15724_n929), .Y(_abc_15724_n930) );
  OR2X2 OR2X2_710 ( .A(_abc_15724_n2909), .B(_abc_15724_n2894_1), .Y(_abc_15724_n2910) );
  OR2X2 OR2X2_711 ( .A(_abc_15724_n2898), .B(_abc_15724_n2910), .Y(_abc_15724_n2911) );
  OR2X2 OR2X2_712 ( .A(_abc_15724_n2913), .B(_abc_15724_n2912), .Y(_abc_15724_n2914) );
  OR2X2 OR2X2_713 ( .A(_abc_15724_n2916), .B(_abc_15724_n2905), .Y(H0_reg_27__FF_INPUT) );
  OR2X2 OR2X2_714 ( .A(_abc_15724_n2860), .B(_abc_15724_n2927_1), .Y(_abc_15724_n2928) );
  OR2X2 OR2X2_715 ( .A(_auto_iopadmap_cc_313_execute_26059_156_), .B(a_reg_28_), .Y(_abc_15724_n2931) );
  OR2X2 OR2X2_716 ( .A(_abc_15724_n2930_1), .B(_abc_15724_n2934), .Y(_abc_15724_n2935) );
  OR2X2 OR2X2_717 ( .A(_abc_15724_n2939), .B(_abc_15724_n2918), .Y(H0_reg_28__FF_INPUT) );
  OR2X2 OR2X2_718 ( .A(_auto_iopadmap_cc_313_execute_26059_157_), .B(a_reg_29_), .Y(_abc_15724_n2942) );
  OR2X2 OR2X2_719 ( .A(_abc_15724_n2941), .B(_abc_15724_n2946), .Y(_abc_15724_n2947) );
  OR2X2 OR2X2_72 ( .A(_abc_15724_n938), .B(_abc_15724_n924), .Y(H4_reg_27__FF_INPUT) );
  OR2X2 OR2X2_720 ( .A(_abc_15724_n2948), .B(_abc_15724_n2945), .Y(_abc_15724_n2949) );
  OR2X2 OR2X2_721 ( .A(_abc_15724_n851_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_157_), .Y(_abc_15724_n2952) );
  OR2X2 OR2X2_722 ( .A(_abc_15724_n2951), .B(_abc_15724_n2953), .Y(H0_reg_29__FF_INPUT) );
  OR2X2 OR2X2_723 ( .A(_auto_iopadmap_cc_313_execute_26059_158_), .B(a_reg_30_), .Y(_abc_15724_n2955) );
  OR2X2 OR2X2_724 ( .A(_abc_15724_n2959), .B(_abc_15724_n2943), .Y(_abc_15724_n2960) );
  OR2X2 OR2X2_725 ( .A(_abc_15724_n2929), .B(_abc_15724_n2963), .Y(_abc_15724_n2964_1) );
  OR2X2 OR2X2_726 ( .A(_abc_15724_n2966), .B(_abc_15724_n2958), .Y(_abc_15724_n2967) );
  OR2X2 OR2X2_727 ( .A(_abc_15724_n2965), .B(_abc_15724_n2968_1), .Y(_abc_15724_n2969) );
  OR2X2 OR2X2_728 ( .A(_abc_15724_n851_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_158_), .Y(_abc_15724_n2972) );
  OR2X2 OR2X2_729 ( .A(_abc_15724_n2971), .B(_abc_15724_n2973), .Y(H0_reg_30__FF_INPUT) );
  OR2X2 OR2X2_73 ( .A(_abc_15724_n932_1), .B(_abc_15724_n942), .Y(_abc_15724_n943_1) );
  OR2X2 OR2X2_730 ( .A(_auto_iopadmap_cc_313_execute_26059_159_), .B(a_reg_31_), .Y(_abc_15724_n2976) );
  OR2X2 OR2X2_731 ( .A(_abc_15724_n2983), .B(_abc_15724_n2980), .Y(_abc_15724_n2984) );
  OR2X2 OR2X2_732 ( .A(_abc_15724_n2985), .B(_abc_15724_n2986), .Y(H0_reg_31__FF_INPUT) );
  OR2X2 OR2X2_733 ( .A(init), .B(next), .Y(_abc_15724_n2988) );
  OR2X2 OR2X2_734 ( .A(_abc_15724_n2996), .B(_abc_15724_n2997), .Y(_abc_15724_n2998) );
  OR2X2 OR2X2_735 ( .A(_abc_15724_n2998), .B(_abc_15724_n2993), .Y(e_reg_0__FF_INPUT) );
  OR2X2 OR2X2_736 ( .A(_abc_15724_n3002), .B(_abc_15724_n3003_1), .Y(_abc_15724_n3004) );
  OR2X2 OR2X2_737 ( .A(_abc_15724_n3004), .B(_abc_15724_n3000), .Y(e_reg_1__FF_INPUT) );
  OR2X2 OR2X2_738 ( .A(_abc_15724_n3008), .B(_abc_15724_n3009), .Y(_abc_15724_n3010) );
  OR2X2 OR2X2_739 ( .A(_abc_15724_n3010), .B(_abc_15724_n3006), .Y(e_reg_2__FF_INPUT) );
  OR2X2 OR2X2_74 ( .A(_auto_iopadmap_cc_313_execute_26059_28_), .B(e_reg_28_), .Y(_abc_15724_n944_1) );
  OR2X2 OR2X2_740 ( .A(_abc_15724_n3014), .B(_abc_15724_n3015), .Y(_abc_15724_n3016) );
  OR2X2 OR2X2_741 ( .A(_abc_15724_n3016), .B(_abc_15724_n3012), .Y(e_reg_3__FF_INPUT) );
  OR2X2 OR2X2_742 ( .A(_abc_15724_n851_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_4_), .Y(_abc_15724_n3019) );
  OR2X2 OR2X2_743 ( .A(_abc_15724_n3020), .B(_abc_15724_n3021), .Y(_abc_15724_n3022) );
  OR2X2 OR2X2_744 ( .A(_abc_15724_n3022), .B(_abc_15724_n3018), .Y(e_reg_4__FF_INPUT) );
  OR2X2 OR2X2_745 ( .A(_abc_15724_n851_bF_buf8), .B(_auto_iopadmap_cc_313_execute_26059_5_), .Y(_abc_15724_n3025) );
  OR2X2 OR2X2_746 ( .A(_abc_15724_n3026), .B(_abc_15724_n3027), .Y(_abc_15724_n3028) );
  OR2X2 OR2X2_747 ( .A(_abc_15724_n3028), .B(_abc_15724_n3024), .Y(e_reg_5__FF_INPUT) );
  OR2X2 OR2X2_748 ( .A(_abc_15724_n851_bF_buf7), .B(_auto_iopadmap_cc_313_execute_26059_6_), .Y(_abc_15724_n3031) );
  OR2X2 OR2X2_749 ( .A(_abc_15724_n3032), .B(_abc_15724_n3033), .Y(_abc_15724_n3034) );
  OR2X2 OR2X2_75 ( .A(_abc_15724_n943_1), .B(_abc_15724_n947), .Y(_abc_15724_n948) );
  OR2X2 OR2X2_750 ( .A(_abc_15724_n3034), .B(_abc_15724_n3030), .Y(e_reg_6__FF_INPUT) );
  OR2X2 OR2X2_751 ( .A(_abc_15724_n851_bF_buf6), .B(_auto_iopadmap_cc_313_execute_26059_7_), .Y(_abc_15724_n3037) );
  OR2X2 OR2X2_752 ( .A(_abc_15724_n3038), .B(_abc_15724_n3039), .Y(_abc_15724_n3040_1) );
  OR2X2 OR2X2_753 ( .A(_abc_15724_n3040_1), .B(_abc_15724_n3036), .Y(e_reg_7__FF_INPUT) );
  OR2X2 OR2X2_754 ( .A(_abc_15724_n851_bF_buf5), .B(_auto_iopadmap_cc_313_execute_26059_8_), .Y(_abc_15724_n3043) );
  OR2X2 OR2X2_755 ( .A(_abc_15724_n3044_1), .B(_abc_15724_n3045), .Y(_abc_15724_n3046) );
  OR2X2 OR2X2_756 ( .A(_abc_15724_n3046), .B(_abc_15724_n3042), .Y(e_reg_8__FF_INPUT) );
  OR2X2 OR2X2_757 ( .A(_abc_15724_n3050), .B(_abc_15724_n3051), .Y(_abc_15724_n3052) );
  OR2X2 OR2X2_758 ( .A(_abc_15724_n3052), .B(_abc_15724_n3048), .Y(e_reg_9__FF_INPUT) );
  OR2X2 OR2X2_759 ( .A(_abc_15724_n3056), .B(_abc_15724_n3057), .Y(_abc_15724_n3058) );
  OR2X2 OR2X2_76 ( .A(_abc_15724_n952), .B(_abc_15724_n940), .Y(H4_reg_28__FF_INPUT) );
  OR2X2 OR2X2_760 ( .A(_abc_15724_n3058), .B(_abc_15724_n3054), .Y(e_reg_10__FF_INPUT) );
  OR2X2 OR2X2_761 ( .A(_abc_15724_n3062), .B(_abc_15724_n3063), .Y(_abc_15724_n3064) );
  OR2X2 OR2X2_762 ( .A(_abc_15724_n3064), .B(_abc_15724_n3060), .Y(e_reg_11__FF_INPUT) );
  OR2X2 OR2X2_763 ( .A(_abc_15724_n3068), .B(_abc_15724_n3069), .Y(_abc_15724_n3070) );
  OR2X2 OR2X2_764 ( .A(_abc_15724_n3070), .B(_abc_15724_n3066), .Y(e_reg_12__FF_INPUT) );
  OR2X2 OR2X2_765 ( .A(_abc_15724_n851_bF_buf4), .B(_auto_iopadmap_cc_313_execute_26059_13_), .Y(_abc_15724_n3073) );
  OR2X2 OR2X2_766 ( .A(_abc_15724_n3074), .B(_abc_15724_n3075), .Y(_abc_15724_n3076_1) );
  OR2X2 OR2X2_767 ( .A(_abc_15724_n3076_1), .B(_abc_15724_n3072), .Y(e_reg_13__FF_INPUT) );
  OR2X2 OR2X2_768 ( .A(_abc_15724_n851_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_14_), .Y(_abc_15724_n3079_1) );
  OR2X2 OR2X2_769 ( .A(_abc_15724_n3080), .B(_abc_15724_n3081), .Y(_abc_15724_n3082) );
  OR2X2 OR2X2_77 ( .A(_abc_15724_n954_1), .B(digest_update_bF_buf3), .Y(_abc_15724_n955) );
  OR2X2 OR2X2_770 ( .A(_abc_15724_n3082), .B(_abc_15724_n3078), .Y(e_reg_14__FF_INPUT) );
  OR2X2 OR2X2_771 ( .A(_abc_15724_n851_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_15_), .Y(_abc_15724_n3085) );
  OR2X2 OR2X2_772 ( .A(_abc_15724_n3086), .B(_abc_15724_n3087), .Y(_abc_15724_n3088) );
  OR2X2 OR2X2_773 ( .A(_abc_15724_n3088), .B(_abc_15724_n3084), .Y(e_reg_15__FF_INPUT) );
  OR2X2 OR2X2_774 ( .A(_abc_15724_n3092), .B(_abc_15724_n3093), .Y(_abc_15724_n3094) );
  OR2X2 OR2X2_775 ( .A(_abc_15724_n3094), .B(_abc_15724_n3090), .Y(e_reg_16__FF_INPUT) );
  OR2X2 OR2X2_776 ( .A(_abc_15724_n851_bF_buf1), .B(_auto_iopadmap_cc_313_execute_26059_17_), .Y(_abc_15724_n3097) );
  OR2X2 OR2X2_777 ( .A(_abc_15724_n3098), .B(_abc_15724_n3099), .Y(_abc_15724_n3100) );
  OR2X2 OR2X2_778 ( .A(_abc_15724_n3100), .B(_abc_15724_n3096), .Y(e_reg_17__FF_INPUT) );
  OR2X2 OR2X2_779 ( .A(_abc_15724_n3104), .B(_abc_15724_n3105), .Y(_abc_15724_n3106) );
  OR2X2 OR2X2_78 ( .A(_auto_iopadmap_cc_313_execute_26059_29_), .B(e_reg_29_), .Y(_abc_15724_n958) );
  OR2X2 OR2X2_780 ( .A(_abc_15724_n3106), .B(_abc_15724_n3102), .Y(e_reg_18__FF_INPUT) );
  OR2X2 OR2X2_781 ( .A(_abc_15724_n3110), .B(_abc_15724_n3111), .Y(_abc_15724_n3112) );
  OR2X2 OR2X2_782 ( .A(_abc_15724_n3112), .B(_abc_15724_n3108), .Y(e_reg_19__FF_INPUT) );
  OR2X2 OR2X2_783 ( .A(_abc_15724_n851_bF_buf0), .B(_auto_iopadmap_cc_313_execute_26059_20_), .Y(_abc_15724_n3115) );
  OR2X2 OR2X2_784 ( .A(_abc_15724_n3116), .B(_abc_15724_n3117), .Y(_abc_15724_n3118_1) );
  OR2X2 OR2X2_785 ( .A(_abc_15724_n3118_1), .B(_abc_15724_n3114_1), .Y(e_reg_20__FF_INPUT) );
  OR2X2 OR2X2_786 ( .A(_abc_15724_n3122), .B(_abc_15724_n3123), .Y(_abc_15724_n3124) );
  OR2X2 OR2X2_787 ( .A(_abc_15724_n3124), .B(_abc_15724_n3120), .Y(e_reg_21__FF_INPUT) );
  OR2X2 OR2X2_788 ( .A(_abc_15724_n3127), .B(_abc_15724_n3128), .Y(_abc_15724_n3129) );
  OR2X2 OR2X2_789 ( .A(_abc_15724_n3129), .B(_abc_15724_n3126), .Y(e_reg_22__FF_INPUT) );
  OR2X2 OR2X2_79 ( .A(_abc_15724_n957), .B(_abc_15724_n961), .Y(_abc_15724_n962) );
  OR2X2 OR2X2_790 ( .A(_abc_15724_n3132), .B(_abc_15724_n3133), .Y(_abc_15724_n3134) );
  OR2X2 OR2X2_791 ( .A(_abc_15724_n3134), .B(_abc_15724_n3131), .Y(e_reg_23__FF_INPUT) );
  OR2X2 OR2X2_792 ( .A(_abc_15724_n3137), .B(_abc_15724_n3138), .Y(_abc_15724_n3139) );
  OR2X2 OR2X2_793 ( .A(_abc_15724_n3139), .B(_abc_15724_n3136), .Y(e_reg_24__FF_INPUT) );
  OR2X2 OR2X2_794 ( .A(_abc_15724_n3142), .B(_abc_15724_n3143), .Y(_abc_15724_n3144) );
  OR2X2 OR2X2_795 ( .A(_abc_15724_n3144), .B(_abc_15724_n3141), .Y(e_reg_25__FF_INPUT) );
  OR2X2 OR2X2_796 ( .A(_abc_15724_n3148), .B(_abc_15724_n3149), .Y(_abc_15724_n3150_1) );
  OR2X2 OR2X2_797 ( .A(_abc_15724_n3150_1), .B(_abc_15724_n3146), .Y(e_reg_26__FF_INPUT) );
  OR2X2 OR2X2_798 ( .A(_abc_15724_n3154), .B(_abc_15724_n3155), .Y(_abc_15724_n3156) );
  OR2X2 OR2X2_799 ( .A(_abc_15724_n3156), .B(_abc_15724_n3152), .Y(e_reg_27__FF_INPUT) );
  OR2X2 OR2X2_8 ( .A(_abc_15724_n724), .B(_abc_15724_n726), .Y(_abc_15724_n727) );
  OR2X2 OR2X2_80 ( .A(_abc_15724_n956_1), .B(_abc_15724_n963), .Y(_abc_15724_n964) );
  OR2X2 OR2X2_800 ( .A(_abc_15724_n3160), .B(_abc_15724_n3161), .Y(_abc_15724_n3162) );
  OR2X2 OR2X2_801 ( .A(_abc_15724_n3162), .B(_abc_15724_n3158), .Y(e_reg_28__FF_INPUT) );
  OR2X2 OR2X2_802 ( .A(_abc_15724_n3165), .B(_abc_15724_n3166), .Y(_abc_15724_n3167) );
  OR2X2 OR2X2_803 ( .A(_abc_15724_n3167), .B(_abc_15724_n3164), .Y(e_reg_29__FF_INPUT) );
  OR2X2 OR2X2_804 ( .A(_abc_15724_n3170), .B(_abc_15724_n3171), .Y(_abc_15724_n3172) );
  OR2X2 OR2X2_805 ( .A(_abc_15724_n3172), .B(_abc_15724_n3169), .Y(e_reg_30__FF_INPUT) );
  OR2X2 OR2X2_806 ( .A(_abc_15724_n3175), .B(_abc_15724_n3176), .Y(_abc_15724_n3177) );
  OR2X2 OR2X2_807 ( .A(_abc_15724_n3177), .B(_abc_15724_n3174), .Y(e_reg_31__FF_INPUT) );
  OR2X2 OR2X2_808 ( .A(_abc_15724_n3180), .B(_abc_15724_n3181), .Y(_abc_15724_n3182) );
  OR2X2 OR2X2_809 ( .A(_abc_15724_n3182), .B(_abc_15724_n3179), .Y(d_reg_0__FF_INPUT) );
  OR2X2 OR2X2_81 ( .A(_abc_15724_n965), .B(_abc_15724_n850_bF_buf3), .Y(_abc_15724_n966_1) );
  OR2X2 OR2X2_810 ( .A(_abc_15724_n3185), .B(_abc_15724_n3186), .Y(_abc_15724_n3187) );
  OR2X2 OR2X2_811 ( .A(_abc_15724_n3187), .B(_abc_15724_n3184), .Y(d_reg_1__FF_INPUT) );
  OR2X2 OR2X2_812 ( .A(_abc_15724_n3190), .B(_abc_15724_n3191), .Y(_abc_15724_n3192) );
  OR2X2 OR2X2_813 ( .A(_abc_15724_n3192), .B(_abc_15724_n3189), .Y(d_reg_2__FF_INPUT) );
  OR2X2 OR2X2_814 ( .A(_abc_15724_n3196), .B(_abc_15724_n3197), .Y(_abc_15724_n3198_1) );
  OR2X2 OR2X2_815 ( .A(_abc_15724_n3198_1), .B(_abc_15724_n3194), .Y(d_reg_3__FF_INPUT) );
  OR2X2 OR2X2_816 ( .A(_abc_15724_n3201), .B(_abc_15724_n3202), .Y(_abc_15724_n3203) );
  OR2X2 OR2X2_817 ( .A(_abc_15724_n3203), .B(_abc_15724_n3200), .Y(d_reg_4__FF_INPUT) );
  OR2X2 OR2X2_818 ( .A(_abc_15724_n3206), .B(_abc_15724_n3207), .Y(_abc_15724_n3208) );
  OR2X2 OR2X2_819 ( .A(_abc_15724_n3208), .B(_abc_15724_n3205), .Y(d_reg_5__FF_INPUT) );
  OR2X2 OR2X2_82 ( .A(e_reg_30_), .B(_auto_iopadmap_cc_313_execute_26059_30_), .Y(_abc_15724_n968_1) );
  OR2X2 OR2X2_820 ( .A(_abc_15724_n3211), .B(_abc_15724_n3212), .Y(_abc_15724_n3213) );
  OR2X2 OR2X2_821 ( .A(_abc_15724_n3213), .B(_abc_15724_n3210), .Y(d_reg_6__FF_INPUT) );
  OR2X2 OR2X2_822 ( .A(_abc_15724_n3217), .B(_abc_15724_n3218), .Y(_abc_15724_n3219) );
  OR2X2 OR2X2_823 ( .A(_abc_15724_n3219), .B(_abc_15724_n3215), .Y(d_reg_7__FF_INPUT) );
  OR2X2 OR2X2_824 ( .A(_abc_15724_n3223), .B(_abc_15724_n3224), .Y(_abc_15724_n3225) );
  OR2X2 OR2X2_825 ( .A(_abc_15724_n3225), .B(_abc_15724_n3221), .Y(d_reg_8__FF_INPUT) );
  OR2X2 OR2X2_826 ( .A(_abc_15724_n3229), .B(_abc_15724_n3230_1), .Y(_abc_15724_n3231) );
  OR2X2 OR2X2_827 ( .A(_abc_15724_n3231), .B(_abc_15724_n3227), .Y(d_reg_9__FF_INPUT) );
  OR2X2 OR2X2_828 ( .A(_abc_15724_n3234), .B(_abc_15724_n3235), .Y(_abc_15724_n3236) );
  OR2X2 OR2X2_829 ( .A(_abc_15724_n3236), .B(_abc_15724_n3233_1), .Y(d_reg_10__FF_INPUT) );
  OR2X2 OR2X2_83 ( .A(_abc_15724_n972), .B(_abc_15724_n959), .Y(_abc_15724_n973) );
  OR2X2 OR2X2_830 ( .A(_abc_15724_n3240), .B(_abc_15724_n3241), .Y(_abc_15724_n3242) );
  OR2X2 OR2X2_831 ( .A(_abc_15724_n3242), .B(_abc_15724_n3238), .Y(d_reg_11__FF_INPUT) );
  OR2X2 OR2X2_832 ( .A(_abc_15724_n3245), .B(_abc_15724_n3246), .Y(_abc_15724_n3247) );
  OR2X2 OR2X2_833 ( .A(_abc_15724_n3247), .B(_abc_15724_n3244), .Y(d_reg_12__FF_INPUT) );
  OR2X2 OR2X2_834 ( .A(_abc_15724_n3251), .B(_abc_15724_n3252), .Y(_abc_15724_n3253) );
  OR2X2 OR2X2_835 ( .A(_abc_15724_n3253), .B(_abc_15724_n3249), .Y(d_reg_13__FF_INPUT) );
  OR2X2 OR2X2_836 ( .A(_abc_15724_n3256), .B(_abc_15724_n3257), .Y(_abc_15724_n3258) );
  OR2X2 OR2X2_837 ( .A(_abc_15724_n3258), .B(_abc_15724_n3255), .Y(d_reg_14__FF_INPUT) );
  OR2X2 OR2X2_838 ( .A(_abc_15724_n3262), .B(_abc_15724_n3263), .Y(_abc_15724_n3264) );
  OR2X2 OR2X2_839 ( .A(_abc_15724_n3264), .B(_abc_15724_n3260), .Y(d_reg_15__FF_INPUT) );
  OR2X2 OR2X2_84 ( .A(_abc_15724_n975), .B(_abc_15724_n973), .Y(_abc_15724_n976_1) );
  OR2X2 OR2X2_840 ( .A(_abc_15724_n3268), .B(_abc_15724_n3269), .Y(_abc_15724_n3270_1) );
  OR2X2 OR2X2_841 ( .A(_abc_15724_n3270_1), .B(_abc_15724_n3266), .Y(d_reg_16__FF_INPUT) );
  OR2X2 OR2X2_842 ( .A(_abc_15724_n3273), .B(_abc_15724_n3274_1), .Y(_abc_15724_n3275) );
  OR2X2 OR2X2_843 ( .A(_abc_15724_n3275), .B(_abc_15724_n3272), .Y(d_reg_17__FF_INPUT) );
  OR2X2 OR2X2_844 ( .A(_abc_15724_n3279), .B(_abc_15724_n3280), .Y(_abc_15724_n3281) );
  OR2X2 OR2X2_845 ( .A(_abc_15724_n3281), .B(_abc_15724_n3277), .Y(d_reg_18__FF_INPUT) );
  OR2X2 OR2X2_846 ( .A(_abc_15724_n3285), .B(_abc_15724_n3286), .Y(_abc_15724_n3287) );
  OR2X2 OR2X2_847 ( .A(_abc_15724_n3287), .B(_abc_15724_n3283), .Y(d_reg_19__FF_INPUT) );
  OR2X2 OR2X2_848 ( .A(_abc_15724_n3290), .B(_abc_15724_n3291), .Y(_abc_15724_n3292) );
  OR2X2 OR2X2_849 ( .A(_abc_15724_n3292), .B(_abc_15724_n3289), .Y(d_reg_20__FF_INPUT) );
  OR2X2 OR2X2_85 ( .A(_abc_15724_n976_1), .B(_abc_15724_n971), .Y(_abc_15724_n977_1) );
  OR2X2 OR2X2_850 ( .A(_abc_15724_n3295), .B(_abc_15724_n3296), .Y(_abc_15724_n3297) );
  OR2X2 OR2X2_851 ( .A(_abc_15724_n3297), .B(_abc_15724_n3294), .Y(d_reg_21__FF_INPUT) );
  OR2X2 OR2X2_852 ( .A(_abc_15724_n3301), .B(_abc_15724_n3302), .Y(_abc_15724_n3303) );
  OR2X2 OR2X2_853 ( .A(_abc_15724_n3303), .B(_abc_15724_n3299), .Y(d_reg_22__FF_INPUT) );
  OR2X2 OR2X2_854 ( .A(_abc_15724_n3307_1), .B(_abc_15724_n3308), .Y(_abc_15724_n3309) );
  OR2X2 OR2X2_855 ( .A(_abc_15724_n3309), .B(_abc_15724_n3305), .Y(d_reg_23__FF_INPUT) );
  OR2X2 OR2X2_856 ( .A(_abc_15724_n3313), .B(_abc_15724_n3314), .Y(_abc_15724_n3315) );
  OR2X2 OR2X2_857 ( .A(_abc_15724_n3315), .B(_abc_15724_n3311_1), .Y(d_reg_24__FF_INPUT) );
  OR2X2 OR2X2_858 ( .A(_abc_15724_n3319), .B(_abc_15724_n3320), .Y(_abc_15724_n3321) );
  OR2X2 OR2X2_859 ( .A(_abc_15724_n3321), .B(_abc_15724_n3317), .Y(d_reg_25__FF_INPUT) );
  OR2X2 OR2X2_86 ( .A(_abc_15724_n851_bF_buf3), .B(_auto_iopadmap_cc_313_execute_26059_30_), .Y(_abc_15724_n982) );
  OR2X2 OR2X2_860 ( .A(_abc_15724_n3325), .B(_abc_15724_n3326), .Y(_abc_15724_n3327) );
  OR2X2 OR2X2_861 ( .A(_abc_15724_n3327), .B(_abc_15724_n3323), .Y(d_reg_26__FF_INPUT) );
  OR2X2 OR2X2_862 ( .A(_abc_15724_n3331), .B(_abc_15724_n3332), .Y(_abc_15724_n3333) );
  OR2X2 OR2X2_863 ( .A(_abc_15724_n3333), .B(_abc_15724_n3329), .Y(d_reg_27__FF_INPUT) );
  OR2X2 OR2X2_864 ( .A(_abc_15724_n3336), .B(_abc_15724_n3337), .Y(_abc_15724_n3338) );
  OR2X2 OR2X2_865 ( .A(_abc_15724_n3338), .B(_abc_15724_n3335), .Y(d_reg_28__FF_INPUT) );
  OR2X2 OR2X2_866 ( .A(_abc_15724_n3341), .B(_abc_15724_n3342), .Y(_abc_15724_n3343) );
  OR2X2 OR2X2_867 ( .A(_abc_15724_n3343), .B(_abc_15724_n3340), .Y(d_reg_29__FF_INPUT) );
  OR2X2 OR2X2_868 ( .A(_abc_15724_n3347), .B(_abc_15724_n3348), .Y(_abc_15724_n3349_1) );
  OR2X2 OR2X2_869 ( .A(_abc_15724_n3349_1), .B(_abc_15724_n3345), .Y(d_reg_30__FF_INPUT) );
  OR2X2 OR2X2_87 ( .A(_abc_15724_n981), .B(_abc_15724_n983), .Y(H4_reg_30__FF_INPUT) );
  OR2X2 OR2X2_870 ( .A(_abc_15724_n3353), .B(_abc_15724_n3354), .Y(_abc_15724_n3355) );
  OR2X2 OR2X2_871 ( .A(_abc_15724_n3355), .B(_abc_15724_n3351), .Y(d_reg_31__FF_INPUT) );
  OR2X2 OR2X2_872 ( .A(_abc_15724_n3358), .B(_abc_15724_n3359), .Y(_abc_15724_n3360) );
  OR2X2 OR2X2_873 ( .A(_abc_15724_n3360), .B(_abc_15724_n3357), .Y(c_reg_0__FF_INPUT) );
  OR2X2 OR2X2_874 ( .A(_abc_15724_n3363), .B(_abc_15724_n3364), .Y(_abc_15724_n3365) );
  OR2X2 OR2X2_875 ( .A(_abc_15724_n3365), .B(_abc_15724_n3362), .Y(c_reg_1__FF_INPUT) );
  OR2X2 OR2X2_876 ( .A(_abc_15724_n3368), .B(_abc_15724_n3369), .Y(_abc_15724_n3370) );
  OR2X2 OR2X2_877 ( .A(_abc_15724_n3370), .B(_abc_15724_n3367), .Y(c_reg_2__FF_INPUT) );
  OR2X2 OR2X2_878 ( .A(_abc_15724_n3373), .B(_abc_15724_n3374), .Y(_abc_15724_n3375) );
  OR2X2 OR2X2_879 ( .A(_abc_15724_n3375), .B(_abc_15724_n3372), .Y(c_reg_3__FF_INPUT) );
  OR2X2 OR2X2_88 ( .A(_abc_15724_n978), .B(_abc_15724_n969), .Y(_abc_15724_n985) );
  OR2X2 OR2X2_880 ( .A(_abc_15724_n3378), .B(_abc_15724_n3379), .Y(_abc_15724_n3380) );
  OR2X2 OR2X2_881 ( .A(_abc_15724_n3380), .B(_abc_15724_n3377), .Y(c_reg_4__FF_INPUT) );
  OR2X2 OR2X2_882 ( .A(_abc_15724_n3383), .B(_abc_15724_n3384), .Y(_abc_15724_n3385) );
  OR2X2 OR2X2_883 ( .A(_abc_15724_n3385), .B(_abc_15724_n3382), .Y(c_reg_5__FF_INPUT) );
  OR2X2 OR2X2_884 ( .A(_abc_15724_n3388), .B(_abc_15724_n3389_1), .Y(_abc_15724_n3390) );
  OR2X2 OR2X2_885 ( .A(_abc_15724_n3390), .B(_abc_15724_n3387), .Y(c_reg_6__FF_INPUT) );
  OR2X2 OR2X2_886 ( .A(_abc_15724_n3393), .B(_abc_15724_n3394), .Y(_abc_15724_n3395) );
  OR2X2 OR2X2_887 ( .A(_abc_15724_n3395), .B(_abc_15724_n3392), .Y(c_reg_7__FF_INPUT) );
  OR2X2 OR2X2_888 ( .A(_abc_15724_n3399), .B(_abc_15724_n3400), .Y(_abc_15724_n3401) );
  OR2X2 OR2X2_889 ( .A(_abc_15724_n3401), .B(_abc_15724_n3397), .Y(c_reg_8__FF_INPUT) );
  OR2X2 OR2X2_89 ( .A(_abc_15724_n986), .B(_auto_iopadmap_cc_313_execute_26059_31_), .Y(_abc_15724_n987_1) );
  OR2X2 OR2X2_890 ( .A(_abc_15724_n3405), .B(_abc_15724_n3406), .Y(_abc_15724_n3407) );
  OR2X2 OR2X2_891 ( .A(_abc_15724_n3407), .B(_abc_15724_n3403), .Y(c_reg_9__FF_INPUT) );
  OR2X2 OR2X2_892 ( .A(_abc_15724_n3410), .B(_abc_15724_n3411), .Y(_abc_15724_n3412) );
  OR2X2 OR2X2_893 ( .A(_abc_15724_n3412), .B(_abc_15724_n3409), .Y(c_reg_10__FF_INPUT) );
  OR2X2 OR2X2_894 ( .A(_abc_15724_n3415), .B(_abc_15724_n3416), .Y(_abc_15724_n3417) );
  OR2X2 OR2X2_895 ( .A(_abc_15724_n3417), .B(_abc_15724_n3414), .Y(c_reg_11__FF_INPUT) );
  OR2X2 OR2X2_896 ( .A(_abc_15724_n3420), .B(_abc_15724_n3421), .Y(_abc_15724_n3422) );
  OR2X2 OR2X2_897 ( .A(_abc_15724_n3422), .B(_abc_15724_n3419), .Y(c_reg_12__FF_INPUT) );
  OR2X2 OR2X2_898 ( .A(_abc_15724_n3426), .B(_abc_15724_n3427), .Y(_abc_15724_n3428) );
  OR2X2 OR2X2_899 ( .A(_abc_15724_n3428), .B(_abc_15724_n3424), .Y(c_reg_13__FF_INPUT) );
  OR2X2 OR2X2_9 ( .A(_auto_iopadmap_cc_313_execute_26059_15_), .B(e_reg_15_), .Y(_abc_15724_n731_1) );
  OR2X2 OR2X2_90 ( .A(_abc_15724_n988_1), .B(e_reg_31_), .Y(_abc_15724_n989_1) );
  OR2X2 OR2X2_900 ( .A(_abc_15724_n3431), .B(_abc_15724_n3432), .Y(_abc_15724_n3433) );
  OR2X2 OR2X2_901 ( .A(_abc_15724_n3433), .B(_abc_15724_n3430), .Y(c_reg_14__FF_INPUT) );
  OR2X2 OR2X2_902 ( .A(_abc_15724_n3436), .B(_abc_15724_n3437), .Y(_abc_15724_n3438) );
  OR2X2 OR2X2_903 ( .A(_abc_15724_n3438), .B(_abc_15724_n3435), .Y(c_reg_15__FF_INPUT) );
  OR2X2 OR2X2_904 ( .A(_abc_15724_n3442), .B(_abc_15724_n3443), .Y(_abc_15724_n3444) );
  OR2X2 OR2X2_905 ( .A(_abc_15724_n3444), .B(_abc_15724_n3440), .Y(c_reg_16__FF_INPUT) );
  OR2X2 OR2X2_906 ( .A(_abc_15724_n3447), .B(_abc_15724_n3448), .Y(_abc_15724_n3449) );
  OR2X2 OR2X2_907 ( .A(_abc_15724_n3449), .B(_abc_15724_n3446), .Y(c_reg_17__FF_INPUT) );
  OR2X2 OR2X2_908 ( .A(_abc_15724_n3453), .B(_abc_15724_n3454), .Y(_abc_15724_n3455) );
  OR2X2 OR2X2_909 ( .A(_abc_15724_n3455), .B(_abc_15724_n3451), .Y(c_reg_18__FF_INPUT) );
  OR2X2 OR2X2_91 ( .A(_abc_15724_n985), .B(_abc_15724_n991), .Y(_abc_15724_n992) );
  OR2X2 OR2X2_910 ( .A(_abc_15724_n3458), .B(_abc_15724_n3459), .Y(_abc_15724_n3460) );
  OR2X2 OR2X2_911 ( .A(_abc_15724_n3460), .B(_abc_15724_n3457), .Y(c_reg_19__FF_INPUT) );
  OR2X2 OR2X2_912 ( .A(_abc_15724_n3463), .B(_abc_15724_n3464), .Y(_abc_15724_n3465_1) );
  OR2X2 OR2X2_913 ( .A(_abc_15724_n3465_1), .B(_abc_15724_n3462), .Y(c_reg_20__FF_INPUT) );
  OR2X2 OR2X2_914 ( .A(_abc_15724_n3468_1), .B(_abc_15724_n3469_1), .Y(_abc_15724_n3470) );
  OR2X2 OR2X2_915 ( .A(_abc_15724_n3470), .B(_abc_15724_n3467), .Y(c_reg_21__FF_INPUT) );
  OR2X2 OR2X2_916 ( .A(_abc_15724_n3474), .B(_abc_15724_n3475), .Y(_abc_15724_n3476) );
  OR2X2 OR2X2_917 ( .A(_abc_15724_n3476), .B(_abc_15724_n3472), .Y(c_reg_22__FF_INPUT) );
  OR2X2 OR2X2_918 ( .A(_abc_15724_n3479), .B(_abc_15724_n3480), .Y(_abc_15724_n3481) );
  OR2X2 OR2X2_919 ( .A(_abc_15724_n3481), .B(_abc_15724_n3478), .Y(c_reg_23__FF_INPUT) );
  OR2X2 OR2X2_92 ( .A(_abc_15724_n993), .B(_abc_15724_n990), .Y(_abc_15724_n994) );
  OR2X2 OR2X2_920 ( .A(_abc_15724_n3485), .B(_abc_15724_n3486), .Y(_abc_15724_n3487) );
  OR2X2 OR2X2_921 ( .A(_abc_15724_n3487), .B(_abc_15724_n3483_1), .Y(c_reg_24__FF_INPUT) );
  OR2X2 OR2X2_922 ( .A(_abc_15724_n3491_1), .B(_abc_15724_n3492_1), .Y(_abc_15724_n3493) );
  OR2X2 OR2X2_923 ( .A(_abc_15724_n3493), .B(_abc_15724_n3489_1), .Y(c_reg_25__FF_INPUT) );
  OR2X2 OR2X2_924 ( .A(_abc_15724_n3497_1), .B(_abc_15724_n3498), .Y(_abc_15724_n3499) );
  OR2X2 OR2X2_925 ( .A(_abc_15724_n3499), .B(_abc_15724_n3495), .Y(c_reg_26__FF_INPUT) );
  OR2X2 OR2X2_926 ( .A(_abc_15724_n3502), .B(_abc_15724_n3503), .Y(_abc_15724_n3504) );
  OR2X2 OR2X2_927 ( .A(_abc_15724_n3504), .B(_abc_15724_n3501_1), .Y(c_reg_27__FF_INPUT) );
  OR2X2 OR2X2_928 ( .A(_abc_15724_n3507_1), .B(_abc_15724_n3508), .Y(_abc_15724_n3509) );
  OR2X2 OR2X2_929 ( .A(_abc_15724_n3509), .B(_abc_15724_n3506), .Y(c_reg_28__FF_INPUT) );
  OR2X2 OR2X2_93 ( .A(_abc_15724_n851_bF_buf2), .B(_auto_iopadmap_cc_313_execute_26059_31_), .Y(_abc_15724_n997_1) );
  OR2X2 OR2X2_930 ( .A(_abc_15724_n3513_1), .B(_abc_15724_n3514_1), .Y(_abc_15724_n3515) );
  OR2X2 OR2X2_931 ( .A(_abc_15724_n3515), .B(_abc_15724_n3511), .Y(c_reg_29__FF_INPUT) );
  OR2X2 OR2X2_932 ( .A(_abc_15724_n3519), .B(_abc_15724_n3520), .Y(_abc_15724_n3521_1) );
  OR2X2 OR2X2_933 ( .A(_abc_15724_n3521_1), .B(_abc_15724_n3517_1), .Y(c_reg_30__FF_INPUT) );
  OR2X2 OR2X2_934 ( .A(_abc_15724_n3524), .B(_abc_15724_n3525), .Y(_abc_15724_n3526) );
  OR2X2 OR2X2_935 ( .A(_abc_15724_n3526), .B(_abc_15724_n3523), .Y(c_reg_31__FF_INPUT) );
  OR2X2 OR2X2_936 ( .A(_abc_15724_n3529_1), .B(_abc_15724_n3530), .Y(_abc_15724_n3531) );
  OR2X2 OR2X2_937 ( .A(_abc_15724_n3531), .B(_abc_15724_n3528_1), .Y(b_reg_0__FF_INPUT) );
  OR2X2 OR2X2_938 ( .A(_abc_15724_n3535_1), .B(_abc_15724_n3536), .Y(_abc_15724_n3537) );
  OR2X2 OR2X2_939 ( .A(_abc_15724_n3537), .B(_abc_15724_n3533), .Y(b_reg_1__FF_INPUT) );
  OR2X2 OR2X2_94 ( .A(_abc_15724_n996_1), .B(_abc_15724_n998_1), .Y(H4_reg_31__FF_INPUT) );
  OR2X2 OR2X2_940 ( .A(_abc_15724_n3541), .B(_abc_15724_n3542), .Y(_abc_15724_n3543) );
  OR2X2 OR2X2_941 ( .A(_abc_15724_n3543), .B(_abc_15724_n3539), .Y(b_reg_2__FF_INPUT) );
  OR2X2 OR2X2_942 ( .A(_abc_15724_n3546_1), .B(_abc_15724_n3547), .Y(_abc_15724_n3548) );
  OR2X2 OR2X2_943 ( .A(_abc_15724_n3548), .B(_abc_15724_n3545), .Y(b_reg_3__FF_INPUT) );
  OR2X2 OR2X2_944 ( .A(_abc_15724_n3552), .B(_abc_15724_n3553), .Y(_abc_15724_n3554_1) );
  OR2X2 OR2X2_945 ( .A(_abc_15724_n3554_1), .B(_abc_15724_n3550), .Y(b_reg_4__FF_INPUT) );
  OR2X2 OR2X2_946 ( .A(_abc_15724_n3558), .B(_abc_15724_n3559), .Y(_abc_15724_n3560) );
  OR2X2 OR2X2_947 ( .A(_abc_15724_n3560), .B(_abc_15724_n3556), .Y(b_reg_5__FF_INPUT) );
  OR2X2 OR2X2_948 ( .A(_abc_15724_n3564_1), .B(_abc_15724_n3565), .Y(_abc_15724_n3566) );
  OR2X2 OR2X2_949 ( .A(_abc_15724_n3566), .B(_abc_15724_n3562), .Y(b_reg_6__FF_INPUT) );
  OR2X2 OR2X2_95 ( .A(_auto_iopadmap_cc_313_execute_26059_32_), .B(d_reg_0_), .Y(_abc_15724_n1000) );
  OR2X2 OR2X2_950 ( .A(_abc_15724_n3569), .B(_abc_15724_n3570), .Y(_abc_15724_n3571) );
  OR2X2 OR2X2_951 ( .A(_abc_15724_n3571), .B(_abc_15724_n3568), .Y(b_reg_7__FF_INPUT) );
  OR2X2 OR2X2_952 ( .A(_abc_15724_n3574), .B(_abc_15724_n3575), .Y(_abc_15724_n3576) );
  OR2X2 OR2X2_953 ( .A(_abc_15724_n3576), .B(_abc_15724_n3573), .Y(b_reg_8__FF_INPUT) );
  OR2X2 OR2X2_954 ( .A(_abc_15724_n3579), .B(_abc_15724_n3580), .Y(_abc_15724_n3581) );
  OR2X2 OR2X2_955 ( .A(_abc_15724_n3581), .B(_abc_15724_n3578), .Y(b_reg_9__FF_INPUT) );
  OR2X2 OR2X2_956 ( .A(_abc_15724_n3585_1), .B(_abc_15724_n3586), .Y(_abc_15724_n3587) );
  OR2X2 OR2X2_957 ( .A(_abc_15724_n3587), .B(_abc_15724_n3583), .Y(b_reg_10__FF_INPUT) );
  OR2X2 OR2X2_958 ( .A(_abc_15724_n3590), .B(_abc_15724_n3591_1), .Y(_abc_15724_n3592_1) );
  OR2X2 OR2X2_959 ( .A(_abc_15724_n3592_1), .B(_abc_15724_n3589), .Y(b_reg_11__FF_INPUT) );
  OR2X2 OR2X2_96 ( .A(_abc_15724_n1003), .B(_abc_15724_n850_bF_buf0), .Y(_abc_15724_n1004) );
  OR2X2 OR2X2_960 ( .A(_abc_15724_n3596), .B(_abc_15724_n3597), .Y(_abc_15724_n3598) );
  OR2X2 OR2X2_961 ( .A(_abc_15724_n3598), .B(_abc_15724_n3594), .Y(b_reg_12__FF_INPUT) );
  OR2X2 OR2X2_962 ( .A(_abc_15724_n3601), .B(_abc_15724_n3602_1), .Y(_abc_15724_n3603_1) );
  OR2X2 OR2X2_963 ( .A(_abc_15724_n3603_1), .B(_abc_15724_n3600), .Y(b_reg_13__FF_INPUT) );
  OR2X2 OR2X2_964 ( .A(_abc_15724_n3607), .B(_abc_15724_n3608), .Y(_abc_15724_n3609_1) );
  OR2X2 OR2X2_965 ( .A(_abc_15724_n3609_1), .B(_abc_15724_n3605), .Y(b_reg_14__FF_INPUT) );
  OR2X2 OR2X2_966 ( .A(_abc_15724_n3612), .B(_abc_15724_n3613), .Y(_abc_15724_n3614) );
  OR2X2 OR2X2_967 ( .A(_abc_15724_n3614), .B(_abc_15724_n3611), .Y(b_reg_15__FF_INPUT) );
  OR2X2 OR2X2_968 ( .A(_abc_15724_n3617), .B(_abc_15724_n3618), .Y(_abc_15724_n3619) );
  OR2X2 OR2X2_969 ( .A(_abc_15724_n3619), .B(_abc_15724_n3616), .Y(b_reg_16__FF_INPUT) );
  OR2X2 OR2X2_97 ( .A(_abc_15724_n1005), .B(digest_update_bF_buf0), .Y(_abc_15724_n1006) );
  OR2X2 OR2X2_970 ( .A(_abc_15724_n3623), .B(_abc_15724_n3624), .Y(_abc_15724_n3625) );
  OR2X2 OR2X2_971 ( .A(_abc_15724_n3625), .B(_abc_15724_n3621_1), .Y(b_reg_17__FF_INPUT) );
  OR2X2 OR2X2_972 ( .A(_abc_15724_n3628), .B(_abc_15724_n3629_1), .Y(_abc_15724_n3630) );
  OR2X2 OR2X2_973 ( .A(_abc_15724_n3630), .B(_abc_15724_n3627), .Y(b_reg_18__FF_INPUT) );
  OR2X2 OR2X2_974 ( .A(_abc_15724_n3633), .B(_abc_15724_n3634), .Y(_abc_15724_n3635) );
  OR2X2 OR2X2_975 ( .A(_abc_15724_n3635), .B(_abc_15724_n3632), .Y(b_reg_19__FF_INPUT) );
  OR2X2 OR2X2_976 ( .A(_abc_15724_n3639_1), .B(_abc_15724_n3640), .Y(_abc_15724_n3641) );
  OR2X2 OR2X2_977 ( .A(_abc_15724_n3641), .B(_abc_15724_n3637), .Y(b_reg_20__FF_INPUT) );
  OR2X2 OR2X2_978 ( .A(_abc_15724_n3645_1), .B(_abc_15724_n3646_1), .Y(_abc_15724_n3647) );
  OR2X2 OR2X2_979 ( .A(_abc_15724_n3647), .B(_abc_15724_n3643), .Y(b_reg_21__FF_INPUT) );
  OR2X2 OR2X2_98 ( .A(_abc_15724_n1010), .B(_abc_15724_n1011), .Y(_abc_15724_n1012) );
  OR2X2 OR2X2_980 ( .A(_abc_15724_n3650), .B(_abc_15724_n3651), .Y(_abc_15724_n3652) );
  OR2X2 OR2X2_981 ( .A(_abc_15724_n3652), .B(_abc_15724_n3649), .Y(b_reg_22__FF_INPUT) );
  OR2X2 OR2X2_982 ( .A(_abc_15724_n3655), .B(_abc_15724_n3656), .Y(_abc_15724_n3657) );
  OR2X2 OR2X2_983 ( .A(_abc_15724_n3657), .B(_abc_15724_n3654), .Y(b_reg_23__FF_INPUT) );
  OR2X2 OR2X2_984 ( .A(_abc_15724_n3660), .B(_abc_15724_n3661), .Y(_abc_15724_n3662_1) );
  OR2X2 OR2X2_985 ( .A(_abc_15724_n3662_1), .B(_abc_15724_n3659), .Y(b_reg_24__FF_INPUT) );
  OR2X2 OR2X2_986 ( .A(_abc_15724_n3665), .B(_abc_15724_n3666), .Y(_abc_15724_n3667) );
  OR2X2 OR2X2_987 ( .A(_abc_15724_n3667), .B(_abc_15724_n3664), .Y(b_reg_25__FF_INPUT) );
  OR2X2 OR2X2_988 ( .A(_abc_15724_n3670_1), .B(_abc_15724_n3671_1), .Y(_abc_15724_n3672) );
  OR2X2 OR2X2_989 ( .A(_abc_15724_n3672), .B(_abc_15724_n3669), .Y(b_reg_26__FF_INPUT) );
  OR2X2 OR2X2_99 ( .A(_abc_15724_n1012), .B(_abc_15724_n1002), .Y(_abc_15724_n1013) );
  OR2X2 OR2X2_990 ( .A(_abc_15724_n3675), .B(_abc_15724_n3676), .Y(_abc_15724_n3677) );
  OR2X2 OR2X2_991 ( .A(_abc_15724_n3677), .B(_abc_15724_n3674), .Y(b_reg_27__FF_INPUT) );
  OR2X2 OR2X2_992 ( .A(_abc_15724_n3681), .B(_abc_15724_n3682), .Y(_abc_15724_n3683) );
  OR2X2 OR2X2_993 ( .A(_abc_15724_n3683), .B(_abc_15724_n3679_1), .Y(b_reg_28__FF_INPUT) );
  OR2X2 OR2X2_994 ( .A(_abc_15724_n3686_1), .B(_abc_15724_n3687), .Y(_abc_15724_n3688) );
  OR2X2 OR2X2_995 ( .A(_abc_15724_n3688), .B(_abc_15724_n3685), .Y(b_reg_29__FF_INPUT) );
  OR2X2 OR2X2_996 ( .A(_abc_15724_n3691), .B(_abc_15724_n3692), .Y(_abc_15724_n3693) );
  OR2X2 OR2X2_997 ( .A(_abc_15724_n3693), .B(_abc_15724_n3690), .Y(b_reg_30__FF_INPUT) );
  OR2X2 OR2X2_998 ( .A(_abc_15724_n3696), .B(_abc_15724_n3697), .Y(_abc_15724_n3698_1) );
  OR2X2 OR2X2_999 ( .A(_abc_15724_n3698_1), .B(_abc_15724_n3695), .Y(b_reg_31__FF_INPUT) );
endmodule
