module completogpio(\WAddress[0] , \WAddress[1] , \WAddress[2] , \WAddress[3] , \WAddress[4] , \WAddress[5] , \WAddress[6] , \WAddress[7] , \WAddress[8] , \WAddress[9] , \WAddress[10] , \WAddress[11] , \WAddress[12] , \WAddress[13] , \WAddress[14] , \WAddress[15] , \WAddress[16] , \WAddress[17] , \WAddress[18] , \WAddress[19] , \WAddress[20] , \WAddress[21] , \WAddress[22] , \WAddress[23] , \WAddress[24] , \WAddress[25] , \WAddress[26] , \WAddress[27] , \WAddress[28] , \WAddress[29] , \WAddress[30] , \WAddress[31] , \Wdata[0] , \Wdata[1] , \Wdata[2] , \Wdata[3] , \Wdata[4] , \Wdata[5] , \Wdata[6] , \Wdata[7] , \Wdata[8] , \Wdata[9] , \Wdata[10] , \Wdata[11] , \Wdata[12] , \Wdata[13] , \Wdata[14] , \Wdata[15] , \Wdata[16] , \Wdata[17] , \Wdata[18] , \Wdata[19] , \Wdata[20] , \Wdata[21] , \Wdata[22] , \Wdata[23] , \Wdata[24] , \Wdata[25] , \Wdata[26] , \Wdata[27] , \Wdata[28] , \Wdata[29] , \Wdata[30] , \Wdata[31] , AWvalid, \pindata[0] , \pindata[1] , \pindata[2] , \pindata[3] , \pindata[4] , \pindata[5] , \pindata[6] , \pindata[7] , \RAddress[0] , \RAddress[1] , \RAddress[2] , \RAddress[3] , \RAddress[4] , \RAddress[5] , \RAddress[6] , \RAddress[7] , \RAddress[8] , \RAddress[9] , \RAddress[10] , \RAddress[11] , \RAddress[12] , \RAddress[13] , \RAddress[14] , \RAddress[15] , \RAddress[16] , \RAddress[17] , \RAddress[18] , \RAddress[19] , \RAddress[20] , \RAddress[21] , \RAddress[22] , \RAddress[23] , \RAddress[24] , \RAddress[25] , \RAddress[26] , \RAddress[27] , \RAddress[28] , \RAddress[29] , \RAddress[30] , \RAddress[31] , Wvalid, clock, ARvalid, reset, Rready, Bready, ARready, Rvalid, AWready, Wready, Bvalid, \Rx[0] , \Rx[1] , \Rx[2] , \Rx[3] , \Rx[4] , \Rx[5] , \Rx[6] , \Rx[7] , \datanw[0] , \datanw[1] , \datanw[2] , \datanw[3] , \datanw[4] , \datanw[5] , \datanw[6] , \datanw[7] , \Tx[0] , \Tx[1] , \Tx[2] , \Tx[3] , \Tx[4] , \Tx[5] , \Tx[6] , \Tx[7] , \DSE[0] , \DSE[1] , \DSE[2] , \DSE[3] , \DSE[4] , \DSE[5] , \DSE[6] , \DSE[7] , \Rdata[0] , \Rdata[1] , \Rdata[2] , \Rdata[3] , \Rdata[4] , \Rdata[5] , \Rdata[6] , \Rdata[7] , \Rdata[8] , \Rdata[9] , \Rdata[10] , \Rdata[11] , \Rdata[12] , \Rdata[13] , \Rdata[14] , \Rdata[15] , \Rdata[16] , \Rdata[17] , \Rdata[18] , \Rdata[19] , \Rdata[20] , \Rdata[21] , \Rdata[22] , \Rdata[23] , \Rdata[24] , \Rdata[25] , \Rdata[26] , \Rdata[27] , \Rdata[28] , \Rdata[29] , \Rdata[30] , \Rdata[31] );
  output ARready;
  input ARvalid;
  output AWready;
  input AWvalid;
  input Bready;
  output Bvalid;
  output \DSE[0] ;
  output \DSE[1] ;
  output \DSE[2] ;
  output \DSE[3] ;
  output \DSE[4] ;
  output \DSE[5] ;
  output \DSE[6] ;
  output \DSE[7] ;
  wire LRAddress_0_;
  wire LRAddress_1_;
  wire LRAddress_2_;
  wire LWAddress_0_;
  wire LWAddress_1_;
  wire LWAddress_2_;
  input \RAddress[0] ;
  input \RAddress[10] ;
  input \RAddress[11] ;
  input \RAddress[12] ;
  input \RAddress[13] ;
  input \RAddress[14] ;
  input \RAddress[15] ;
  input \RAddress[16] ;
  input \RAddress[17] ;
  input \RAddress[18] ;
  input \RAddress[19] ;
  input \RAddress[1] ;
  input \RAddress[20] ;
  input \RAddress[21] ;
  input \RAddress[22] ;
  input \RAddress[23] ;
  input \RAddress[24] ;
  input \RAddress[25] ;
  input \RAddress[26] ;
  input \RAddress[27] ;
  input \RAddress[28] ;
  input \RAddress[29] ;
  input \RAddress[2] ;
  input \RAddress[30] ;
  input \RAddress[31] ;
  input \RAddress[3] ;
  input \RAddress[4] ;
  input \RAddress[5] ;
  input \RAddress[6] ;
  input \RAddress[7] ;
  input \RAddress[8] ;
  input \RAddress[9] ;
  output \Rdata[0] ;
  output \Rdata[10] ;
  output \Rdata[11] ;
  output \Rdata[12] ;
  output \Rdata[13] ;
  output \Rdata[14] ;
  output \Rdata[15] ;
  output \Rdata[16] ;
  output \Rdata[17] ;
  output \Rdata[18] ;
  output \Rdata[19] ;
  output \Rdata[1] ;
  output \Rdata[20] ;
  output \Rdata[21] ;
  output \Rdata[22] ;
  output \Rdata[23] ;
  output \Rdata[24] ;
  output \Rdata[25] ;
  output \Rdata[26] ;
  output \Rdata[27] ;
  output \Rdata[28] ;
  output \Rdata[29] ;
  output \Rdata[2] ;
  output \Rdata[30] ;
  output \Rdata[31] ;
  output \Rdata[3] ;
  output \Rdata[4] ;
  output \Rdata[5] ;
  output \Rdata[6] ;
  output \Rdata[7] ;
  output \Rdata[8] ;
  output \Rdata[9] ;
  wire Rdata_FF_INPUT;
  input Rready;
  output Rvalid;
  output \Rx[0] ;
  output \Rx[1] ;
  output \Rx[2] ;
  output \Rx[3] ;
  output \Rx[4] ;
  output \Rx[5] ;
  output \Rx[6] ;
  output \Rx[7] ;
  output \Tx[0] ;
  output \Tx[1] ;
  output \Tx[2] ;
  output \Tx[3] ;
  output \Tx[4] ;
  output \Tx[5] ;
  output \Tx[6] ;
  output \Tx[7] ;
  input \WAddress[0] ;
  input \WAddress[10] ;
  input \WAddress[11] ;
  input \WAddress[12] ;
  input \WAddress[13] ;
  input \WAddress[14] ;
  input \WAddress[15] ;
  input \WAddress[16] ;
  input \WAddress[17] ;
  input \WAddress[18] ;
  input \WAddress[19] ;
  input \WAddress[1] ;
  input \WAddress[20] ;
  input \WAddress[21] ;
  input \WAddress[22] ;
  input \WAddress[23] ;
  input \WAddress[24] ;
  input \WAddress[25] ;
  input \WAddress[26] ;
  input \WAddress[27] ;
  input \WAddress[28] ;
  input \WAddress[29] ;
  input \WAddress[2] ;
  input \WAddress[30] ;
  input \WAddress[31] ;
  input \WAddress[3] ;
  input \WAddress[4] ;
  input \WAddress[5] ;
  input \WAddress[6] ;
  input \WAddress[7] ;
  input \WAddress[8] ;
  input \WAddress[9] ;
  input \Wdata[0] ;
  input \Wdata[10] ;
  input \Wdata[11] ;
  input \Wdata[12] ;
  input \Wdata[13] ;
  input \Wdata[14] ;
  input \Wdata[15] ;
  input \Wdata[16] ;
  input \Wdata[17] ;
  input \Wdata[18] ;
  input \Wdata[19] ;
  input \Wdata[1] ;
  input \Wdata[20] ;
  input \Wdata[21] ;
  input \Wdata[22] ;
  input \Wdata[23] ;
  input \Wdata[24] ;
  input \Wdata[25] ;
  input \Wdata[26] ;
  input \Wdata[27] ;
  input \Wdata[28] ;
  input \Wdata[29] ;
  input \Wdata[2] ;
  input \Wdata[30] ;
  input \Wdata[31] ;
  input \Wdata[3] ;
  input \Wdata[4] ;
  input \Wdata[5] ;
  input \Wdata[6] ;
  input \Wdata[7] ;
  input \Wdata[8] ;
  input \Wdata[9] ;
  output Wready;
  input Wvalid;
  wire _abc_1206_n18;
  wire _abc_1206_n19;
  wire _abc_1206_n20;
  wire _abc_1206_n21;
  wire _abc_1206_n23;
  wire _abc_1206_n24;
  wire _abc_1206_n25_1;
  wire _abc_1206_n26;
  wire _abc_1206_n27;
  wire _abc_1206_n28;
  wire _abc_1206_n29;
  wire _abc_1206_n30_1;
  wire _abc_1206_n31_1;
  wire _abc_1206_n32;
  wire _abc_1206_n33;
  wire _abc_1206_n34_1;
  input clock;
  output \datanw[0] ;
  output \datanw[1] ;
  output \datanw[2] ;
  output \datanw[3] ;
  output \datanw[4] ;
  output \datanw[5] ;
  output \datanw[6] ;
  output \datanw[7] ;
  wire decor__abc_1225_n13;
  wire decor__abc_1225_n14_1;
  wire decor__abc_1225_n15;
  wire decor__abc_1225_n17_1;
  wire decor__abc_1225_n18_1;
  wire decor__abc_1225_n20;
  wire decor__abc_1225_n21;
  wire decor__abc_1225_n23;
  wire decor__abc_1225_n25;
  wire decow__abc_1225_n13;
  wire decow__abc_1225_n14_1;
  wire decow__abc_1225_n15;
  wire decow__abc_1225_n17_1;
  wire decow__abc_1225_n18_1;
  wire decow__abc_1225_n20;
  wire decow__abc_1225_n21;
  wire decow__abc_1225_n23;
  wire decow__abc_1225_n25;
  wire flip1_R1;
  wire flip1_Rx;
  wire flip1_Rx_FF_INPUT;
  wire flip1_Tx;
  wire flip1_Tx_FF_INPUT;
  wire flip1_W1;
  wire flip1__abc_1243_n10_1;
  wire flip1__abc_1243_n12;
  wire flip1__abc_1243_n13;
  wire flip1__abc_1243_n8;
  wire flip1__abc_1243_n9;
  wire flip2_R1;
  wire flip2_Rx;
  wire flip2_Rx_FF_INPUT;
  wire flip2_Tx;
  wire flip2_Tx_FF_INPUT;
  wire flip2_W1;
  wire flip2__abc_1243_n10_1;
  wire flip2__abc_1243_n12;
  wire flip2__abc_1243_n13;
  wire flip2__abc_1243_n8;
  wire flip2__abc_1243_n9;
  wire flip3_R1;
  wire flip3_Rx;
  wire flip3_Rx_FF_INPUT;
  wire flip3_Tx;
  wire flip3_Tx_FF_INPUT;
  wire flip3_W1;
  wire flip3__abc_1243_n10_1;
  wire flip3__abc_1243_n12;
  wire flip3__abc_1243_n13;
  wire flip3__abc_1243_n8;
  wire flip3__abc_1243_n9;
  wire flip4_R1;
  wire flip4_Rx;
  wire flip4_Rx_FF_INPUT;
  wire flip4_Tx;
  wire flip4_Tx_FF_INPUT;
  wire flip4_W1;
  wire flip4__abc_1243_n10_1;
  wire flip4__abc_1243_n12;
  wire flip4__abc_1243_n13;
  wire flip4__abc_1243_n8;
  wire flip4__abc_1243_n9;
  wire flip5_R1;
  wire flip5_Rx;
  wire flip5_Rx_FF_INPUT;
  wire flip5_Tx;
  wire flip5_Tx_FF_INPUT;
  wire flip5_W1;
  wire flip5__abc_1243_n10_1;
  wire flip5__abc_1243_n12;
  wire flip5__abc_1243_n13;
  wire flip5__abc_1243_n8;
  wire flip5__abc_1243_n9;
  wire flip6_R1;
  wire flip6_Rx;
  wire flip6_Rx_FF_INPUT;
  wire flip6_Tx;
  wire flip6_Tx_FF_INPUT;
  wire flip6_W1;
  wire flip6__abc_1243_n10_1;
  wire flip6__abc_1243_n12;
  wire flip6__abc_1243_n13;
  wire flip6__abc_1243_n8;
  wire flip6__abc_1243_n9;
  wire flip7_R1;
  wire flip7_Rx;
  wire flip7_Rx_FF_INPUT;
  wire flip7_Tx;
  wire flip7_Tx_FF_INPUT;
  wire flip7_W1;
  wire flip7__abc_1243_n10_1;
  wire flip7__abc_1243_n12;
  wire flip7__abc_1243_n13;
  wire flip7__abc_1243_n8;
  wire flip7__abc_1243_n9;
  wire flip8_R1;
  wire flip8_Rx;
  wire flip8_Rx_FF_INPUT;
  wire flip8_Tx;
  wire flip8_Tx_FF_INPUT;
  wire flip8_W1;
  wire flip8__abc_1243_n10_1;
  wire flip8__abc_1243_n12;
  wire flip8__abc_1243_n13;
  wire flip8__abc_1243_n8;
  wire flip8__abc_1243_n9;
  wire flipw1_DS;
  wire flipw1_DS_FF_INPUT;
  wire flipw1__abc_1251_n10;
  wire flipw1__abc_1251_n11;
  wire flipw1__abc_1251_n12;
  wire flipw1__abc_1251_n14;
  wire flipw1__abc_1251_n15;
  wire flipw1__abc_1251_n9_1;
  wire flipw1_outdata;
  wire flipw1_outdata_FF_INPUT;
  wire flipw2_DS;
  wire flipw2_DS_FF_INPUT;
  wire flipw2__abc_1251_n10;
  wire flipw2__abc_1251_n11;
  wire flipw2__abc_1251_n12;
  wire flipw2__abc_1251_n14;
  wire flipw2__abc_1251_n15;
  wire flipw2__abc_1251_n9_1;
  wire flipw2_outdata;
  wire flipw2_outdata_FF_INPUT;
  wire flipw3_DS;
  wire flipw3_DS_FF_INPUT;
  wire flipw3__abc_1251_n10;
  wire flipw3__abc_1251_n11;
  wire flipw3__abc_1251_n12;
  wire flipw3__abc_1251_n14;
  wire flipw3__abc_1251_n15;
  wire flipw3__abc_1251_n9_1;
  wire flipw3_outdata;
  wire flipw3_outdata_FF_INPUT;
  wire flipw4_DS;
  wire flipw4_DS_FF_INPUT;
  wire flipw4__abc_1251_n10;
  wire flipw4__abc_1251_n11;
  wire flipw4__abc_1251_n12;
  wire flipw4__abc_1251_n14;
  wire flipw4__abc_1251_n15;
  wire flipw4__abc_1251_n9_1;
  wire flipw4_outdata;
  wire flipw4_outdata_FF_INPUT;
  wire flipw5_DS;
  wire flipw5_DS_FF_INPUT;
  wire flipw5__abc_1251_n10;
  wire flipw5__abc_1251_n11;
  wire flipw5__abc_1251_n12;
  wire flipw5__abc_1251_n14;
  wire flipw5__abc_1251_n15;
  wire flipw5__abc_1251_n9_1;
  wire flipw5_outdata;
  wire flipw5_outdata_FF_INPUT;
  wire flipw6_DS;
  wire flipw6_DS_FF_INPUT;
  wire flipw6__abc_1251_n10;
  wire flipw6__abc_1251_n11;
  wire flipw6__abc_1251_n12;
  wire flipw6__abc_1251_n14;
  wire flipw6__abc_1251_n15;
  wire flipw6__abc_1251_n9_1;
  wire flipw6_outdata;
  wire flipw6_outdata_FF_INPUT;
  wire flipw7_DS;
  wire flipw7_DS_FF_INPUT;
  wire flipw7__abc_1251_n10;
  wire flipw7__abc_1251_n11;
  wire flipw7__abc_1251_n12;
  wire flipw7__abc_1251_n14;
  wire flipw7__abc_1251_n15;
  wire flipw7__abc_1251_n9_1;
  wire flipw7_outdata;
  wire flipw7_outdata_FF_INPUT;
  wire flipw8_DS;
  wire flipw8_DS_FF_INPUT;
  wire flipw8__abc_1251_n10;
  wire flipw8__abc_1251_n11;
  wire flipw8__abc_1251_n12;
  wire flipw8__abc_1251_n14;
  wire flipw8__abc_1251_n15;
  wire flipw8__abc_1251_n9_1;
  wire flipw8_outdata;
  wire flipw8_outdata_FF_INPUT;
  wire latchR_LWAddres_0__FF_INPUT;
  wire latchR_LWAddres_1__FF_INPUT;
  wire latchR_LWAddres_2__FF_INPUT;
  wire latchR__abc_1260_n12;
  wire latchR__abc_1260_n13_1;
  wire latchR__abc_1260_n14;
  wire latchR__abc_1260_n15;
  wire latchR__abc_1260_n17;
  wire latchR__abc_1260_n18;
  wire latchR__abc_1260_n20;
  wire latchR__abc_1260_n21;
  wire latchW_LWAddres_0__FF_INPUT;
  wire latchW_LWAddres_1__FF_INPUT;
  wire latchW_LWAddres_2__FF_INPUT;
  wire latchW__abc_1260_n12;
  wire latchW__abc_1260_n13_1;
  wire latchW__abc_1260_n14;
  wire latchW__abc_1260_n15;
  wire latchW__abc_1260_n17;
  wire latchW__abc_1260_n18;
  wire latchW__abc_1260_n20;
  wire latchW__abc_1260_n21;
  wire maquina__abc_1145_n107;
  wire maquina__abc_1145_n108;
  wire maquina__abc_1145_n109;
  wire maquina__abc_1145_n110;
  wire maquina__abc_1145_n111;
  wire maquina__abc_1145_n112;
  wire maquina__abc_1145_n113;
  wire maquina__abc_1145_n14;
  wire maquina__abc_1145_n35;
  wire maquina__abc_1145_n45;
  wire maquina__abc_1145_n9;
  wire maquina__abc_1272_n35_1;
  wire maquina__abc_1272_n36;
  wire maquina__abc_1272_n37_1;
  wire maquina__abc_1272_n38;
  wire maquina__abc_1272_n39;
  wire maquina__abc_1272_n40;
  wire maquina__abc_1272_n41_1;
  wire maquina__abc_1272_n43;
  wire maquina__abc_1272_n44_1;
  wire maquina__abc_1272_n46;
  wire maquina__abc_1272_n47;
  wire maquina__abc_1272_n48;
  wire maquina__abc_1272_n49_1;
  wire maquina__abc_1272_n50;
  wire maquina__abc_1272_n52;
  wire maquina__abc_1272_n53;
  wire maquina__abc_1272_n54;
  wire maquina__abc_1272_n55_1;
  wire maquina__abc_1272_n57;
  wire maquina__abc_1272_n58;
  wire maquina__abc_1272_n59;
  wire maquina__abc_1272_n60_1;
  wire maquina__abc_1272_n61;
  wire maquina__abc_1272_n62;
  wire maquina__abc_1272_n64;
  wire maquina__abc_1272_n66;
  wire maquina__abc_1272_n67_1;
  wire maquina__abc_1272_n69_1;
  wire maquina__abc_1272_n70;
  wire maquina__abc_1272_n71_1;
  wire maquina__abc_1272_n73;
  wire maquina__abc_1272_n74_1;
  wire maquina__abc_1272_n75;
  wire maquina__abc_1272_n79;
  wire maquina__abc_1272_n82;
  wire maquina__abc_1272_n84;
  wire maquina_state_0_;
  wire maquina_state_10_;
  wire maquina_state_1_;
  wire maquina_state_2_;
  wire maquina_state_3_;
  wire maquina_state_4_;
  wire maquina_state_5_;
  wire maquina_state_6_;
  wire maquina_state_7_;
  wire maquina_state_8_;
  wire maquina_state_9_;
  wire maquina_vel;
  input \pindata[0] ;
  input \pindata[1] ;
  input \pindata[2] ;
  input \pindata[3] ;
  input \pindata[4] ;
  input \pindata[5] ;
  input \pindata[6] ;
  input \pindata[7] ;
  input reset;
  wire vel_FF_INPUT;
  AND2X2 AND2X2_1 ( .A(maquina__abc_1272_n48), .B(Rready), .Y(maquina__abc_1272_n49_1) );
  AND2X2 AND2X2_2 ( .A(reset), .B(maquina_state_7_), .Y(maquina__abc_1145_n107) );
  AND2X2 AND2X2_3 ( .A(reset), .B(maquina_state_6_), .Y(maquina__abc_1145_n108) );
  AND2X2 AND2X2_4 ( .A(reset), .B(maquina_state_1_), .Y(maquina__abc_1145_n110) );
  AOI21X1 AOI21X1_1 ( .A(_abc_1206_n19), .B(maquina_vel), .C(_abc_1206_n20), .Y(_abc_1206_n21) );
  AOI21X1 AOI21X1_10 ( .A(flip8__abc_1243_n12), .B(flip8__abc_1243_n10_1), .C(flip8__abc_1243_n13), .Y(flip8_Rx_FF_INPUT) );
  AOI21X1 AOI21X1_11 ( .A(flipw1__abc_1251_n12), .B(flipw1__abc_1251_n10), .C(flipw1__abc_1251_n9_1), .Y(flipw1_outdata_FF_INPUT) );
  AOI21X1 AOI21X1_12 ( .A(flipw1__abc_1251_n15), .B(flipw1__abc_1251_n14), .C(flipw1__abc_1251_n9_1), .Y(flipw1_DS_FF_INPUT) );
  AOI21X1 AOI21X1_13 ( .A(flipw2__abc_1251_n12), .B(flipw2__abc_1251_n10), .C(flipw2__abc_1251_n9_1), .Y(flipw2_outdata_FF_INPUT) );
  AOI21X1 AOI21X1_14 ( .A(flipw2__abc_1251_n15), .B(flipw2__abc_1251_n14), .C(flipw2__abc_1251_n9_1), .Y(flipw2_DS_FF_INPUT) );
  AOI21X1 AOI21X1_15 ( .A(flipw3__abc_1251_n12), .B(flipw3__abc_1251_n10), .C(flipw3__abc_1251_n9_1), .Y(flipw3_outdata_FF_INPUT) );
  AOI21X1 AOI21X1_16 ( .A(flipw3__abc_1251_n15), .B(flipw3__abc_1251_n14), .C(flipw3__abc_1251_n9_1), .Y(flipw3_DS_FF_INPUT) );
  AOI21X1 AOI21X1_17 ( .A(flipw4__abc_1251_n12), .B(flipw4__abc_1251_n10), .C(flipw4__abc_1251_n9_1), .Y(flipw4_outdata_FF_INPUT) );
  AOI21X1 AOI21X1_18 ( .A(flipw4__abc_1251_n15), .B(flipw4__abc_1251_n14), .C(flipw4__abc_1251_n9_1), .Y(flipw4_DS_FF_INPUT) );
  AOI21X1 AOI21X1_19 ( .A(flipw5__abc_1251_n12), .B(flipw5__abc_1251_n10), .C(flipw5__abc_1251_n9_1), .Y(flipw5_outdata_FF_INPUT) );
  AOI21X1 AOI21X1_2 ( .A(_abc_1206_n28), .B(_abc_1206_n34_1), .C(_abc_1206_n20), .Y(Rdata_FF_INPUT) );
  AOI21X1 AOI21X1_20 ( .A(flipw5__abc_1251_n15), .B(flipw5__abc_1251_n14), .C(flipw5__abc_1251_n9_1), .Y(flipw5_DS_FF_INPUT) );
  AOI21X1 AOI21X1_21 ( .A(flipw6__abc_1251_n12), .B(flipw6__abc_1251_n10), .C(flipw6__abc_1251_n9_1), .Y(flipw6_outdata_FF_INPUT) );
  AOI21X1 AOI21X1_22 ( .A(flipw6__abc_1251_n15), .B(flipw6__abc_1251_n14), .C(flipw6__abc_1251_n9_1), .Y(flipw6_DS_FF_INPUT) );
  AOI21X1 AOI21X1_23 ( .A(flipw7__abc_1251_n12), .B(flipw7__abc_1251_n10), .C(flipw7__abc_1251_n9_1), .Y(flipw7_outdata_FF_INPUT) );
  AOI21X1 AOI21X1_24 ( .A(flipw7__abc_1251_n15), .B(flipw7__abc_1251_n14), .C(flipw7__abc_1251_n9_1), .Y(flipw7_DS_FF_INPUT) );
  AOI21X1 AOI21X1_25 ( .A(flipw8__abc_1251_n12), .B(flipw8__abc_1251_n10), .C(flipw8__abc_1251_n9_1), .Y(flipw8_outdata_FF_INPUT) );
  AOI21X1 AOI21X1_26 ( .A(flipw8__abc_1251_n15), .B(flipw8__abc_1251_n14), .C(flipw8__abc_1251_n9_1), .Y(flipw8_DS_FF_INPUT) );
  AOI21X1 AOI21X1_27 ( .A(latchR__abc_1260_n15), .B(latchR__abc_1260_n13_1), .C(latchR__abc_1260_n12), .Y(latchR_LWAddres_0__FF_INPUT) );
  AOI21X1 AOI21X1_28 ( .A(latchR__abc_1260_n18), .B(latchR__abc_1260_n17), .C(latchR__abc_1260_n12), .Y(latchR_LWAddres_1__FF_INPUT) );
  AOI21X1 AOI21X1_29 ( .A(latchR__abc_1260_n21), .B(latchR__abc_1260_n20), .C(latchR__abc_1260_n12), .Y(latchR_LWAddres_2__FF_INPUT) );
  AOI21X1 AOI21X1_3 ( .A(flip1__abc_1243_n12), .B(flip1__abc_1243_n10_1), .C(flip1__abc_1243_n13), .Y(flip1_Rx_FF_INPUT) );
  AOI21X1 AOI21X1_30 ( .A(latchW__abc_1260_n15), .B(latchW__abc_1260_n13_1), .C(latchW__abc_1260_n12), .Y(latchW_LWAddres_0__FF_INPUT) );
  AOI21X1 AOI21X1_31 ( .A(latchW__abc_1260_n18), .B(latchW__abc_1260_n17), .C(latchW__abc_1260_n12), .Y(latchW_LWAddres_1__FF_INPUT) );
  AOI21X1 AOI21X1_32 ( .A(latchW__abc_1260_n21), .B(latchW__abc_1260_n20), .C(latchW__abc_1260_n12), .Y(latchW_LWAddres_2__FF_INPUT) );
  AOI21X1 AOI21X1_33 ( .A(maquina_state_9_), .B(Rready), .C(maquina__abc_1272_n38), .Y(maquina__abc_1272_n39) );
  AOI21X1 AOI21X1_34 ( .A(maquina__abc_1272_n53), .B(maquina__abc_1272_n60_1), .C(maquina__abc_1272_n64), .Y(Wready) );
  AOI21X1 AOI21X1_35 ( .A(maquina__abc_1272_n67_1), .B(maquina__abc_1272_n53), .C(maquina__abc_1272_n66), .Y(AWready) );
  AOI21X1 AOI21X1_36 ( .A(maquina__abc_1272_n75), .B(maquina__abc_1272_n46), .C(maquina_state_0_), .Y(ARready) );
  AOI21X1 AOI21X1_4 ( .A(flip2__abc_1243_n12), .B(flip2__abc_1243_n10_1), .C(flip2__abc_1243_n13), .Y(flip2_Rx_FF_INPUT) );
  AOI21X1 AOI21X1_5 ( .A(flip3__abc_1243_n12), .B(flip3__abc_1243_n10_1), .C(flip3__abc_1243_n13), .Y(flip3_Rx_FF_INPUT) );
  AOI21X1 AOI21X1_6 ( .A(flip4__abc_1243_n12), .B(flip4__abc_1243_n10_1), .C(flip4__abc_1243_n13), .Y(flip4_Rx_FF_INPUT) );
  AOI21X1 AOI21X1_7 ( .A(flip5__abc_1243_n12), .B(flip5__abc_1243_n10_1), .C(flip5__abc_1243_n13), .Y(flip5_Rx_FF_INPUT) );
  AOI21X1 AOI21X1_8 ( .A(flip6__abc_1243_n12), .B(flip6__abc_1243_n10_1), .C(flip6__abc_1243_n13), .Y(flip6_Rx_FF_INPUT) );
  AOI21X1 AOI21X1_9 ( .A(flip7__abc_1243_n12), .B(flip7__abc_1243_n10_1), .C(flip7__abc_1243_n13), .Y(flip7_Rx_FF_INPUT) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(Rdata_FF_INPUT), .Q(\Rdata[0] ) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(flip4_Tx_FF_INPUT), .Q(\Tx[3] ) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(flip5_Rx_FF_INPUT), .Q(\Rx[4] ) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(flip5_Tx_FF_INPUT), .Q(\Tx[4] ) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(flip6_Rx_FF_INPUT), .Q(\Rx[5] ) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(flip6_Tx_FF_INPUT), .Q(\Tx[5] ) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(flip7_Rx_FF_INPUT), .Q(\Rx[6] ) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(flip7_Tx_FF_INPUT), .Q(\Tx[6] ) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(flip8_Rx_FF_INPUT), .Q(\Rx[7] ) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(flip8_Tx_FF_INPUT), .Q(\Tx[7] ) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(flipw1_DS_FF_INPUT), .Q(\DSE[0] ) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(vel_FF_INPUT), .Q(maquina_vel) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(flipw1_outdata_FF_INPUT), .Q(\datanw[0] ) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(flipw2_DS_FF_INPUT), .Q(\DSE[1] ) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(flipw2_outdata_FF_INPUT), .Q(\datanw[1] ) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(flipw3_DS_FF_INPUT), .Q(\DSE[2] ) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(flipw3_outdata_FF_INPUT), .Q(\datanw[2] ) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(flipw4_DS_FF_INPUT), .Q(\DSE[3] ) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(flipw4_outdata_FF_INPUT), .Q(\datanw[3] ) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(flipw5_DS_FF_INPUT), .Q(\DSE[4] ) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(flipw5_outdata_FF_INPUT), .Q(\datanw[4] ) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(clock), .D(flipw6_DS_FF_INPUT), .Q(\DSE[5] ) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(flip1_Rx_FF_INPUT), .Q(\Rx[0] ) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(clock), .D(flipw6_outdata_FF_INPUT), .Q(\datanw[5] ) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(clock), .D(flipw7_DS_FF_INPUT), .Q(\DSE[6] ) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(clock), .D(flipw7_outdata_FF_INPUT), .Q(\datanw[6] ) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(clock), .D(flipw8_DS_FF_INPUT), .Q(\DSE[7] ) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(clock), .D(flipw8_outdata_FF_INPUT), .Q(\datanw[7] ) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(clock), .D(latchR_LWAddres_0__FF_INPUT), .Q(LRAddress_0_) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(clock), .D(latchR_LWAddres_1__FF_INPUT), .Q(LRAddress_1_) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(clock), .D(latchR_LWAddres_2__FF_INPUT), .Q(LRAddress_2_) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(clock), .D(latchW_LWAddres_0__FF_INPUT), .Q(LWAddress_0_) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(clock), .D(latchW_LWAddres_1__FF_INPUT), .Q(LWAddress_1_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(flip1_Tx_FF_INPUT), .Q(\Tx[0] ) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(clock), .D(latchW_LWAddres_2__FF_INPUT), .Q(LWAddress_2_) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(clock), .D(maquina__abc_1145_n9), .Q(maquina_state_0_) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(clock), .D(maquina__abc_1145_n113), .Q(maquina_state_1_) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(clock), .D(maquina__abc_1145_n14), .Q(maquina_state_2_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(clock), .D(maquina__abc_1145_n108), .Q(maquina_state_3_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(clock), .D(maquina__abc_1145_n107), .Q(maquina_state_4_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(clock), .D(maquina__abc_1145_n109), .Q(maquina_state_5_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(clock), .D(maquina__abc_1145_n110), .Q(maquina_state_6_) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(clock), .D(maquina__abc_1145_n111), .Q(maquina_state_7_) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(clock), .D(maquina__abc_1145_n112), .Q(maquina_state_8_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(flip2_Rx_FF_INPUT), .Q(\Rx[1] ) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(clock), .D(maquina__abc_1145_n35), .Q(maquina_state_9_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(clock), .D(maquina__abc_1145_n45), .Q(maquina_state_10_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(flip2_Tx_FF_INPUT), .Q(\Tx[1] ) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(flip3_Rx_FF_INPUT), .Q(\Rx[2] ) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(flip3_Tx_FF_INPUT), .Q(\Tx[2] ) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(flip4_Rx_FF_INPUT), .Q(\Rx[3] ) );
  INVX1 INVX1_1 ( .A(\Wdata[2] ), .Y(_abc_1206_n18) );
  INVX1 INVX1_10 ( .A(LWAddress_1_), .Y(decow__abc_1225_n17_1) );
  INVX1 INVX1_11 ( .A(LWAddress_0_), .Y(decow__abc_1225_n20) );
  INVX1 INVX1_12 ( .A(flip1_W1), .Y(flip1__abc_1243_n8) );
  INVX1 INVX1_13 ( .A(\Rx[0] ), .Y(flip1__abc_1243_n12) );
  INVX1 INVX1_14 ( .A(flip2_W1), .Y(flip2__abc_1243_n8) );
  INVX1 INVX1_15 ( .A(\Rx[1] ), .Y(flip2__abc_1243_n12) );
  INVX1 INVX1_16 ( .A(flip3_W1), .Y(flip3__abc_1243_n8) );
  INVX1 INVX1_17 ( .A(\Rx[2] ), .Y(flip3__abc_1243_n12) );
  INVX1 INVX1_18 ( .A(flip4_W1), .Y(flip4__abc_1243_n8) );
  INVX1 INVX1_19 ( .A(\Rx[3] ), .Y(flip4__abc_1243_n12) );
  INVX1 INVX1_2 ( .A(Wvalid), .Y(_abc_1206_n19) );
  INVX1 INVX1_20 ( .A(flip5_W1), .Y(flip5__abc_1243_n8) );
  INVX1 INVX1_21 ( .A(\Rx[4] ), .Y(flip5__abc_1243_n12) );
  INVX1 INVX1_22 ( .A(flip6_W1), .Y(flip6__abc_1243_n8) );
  INVX1 INVX1_23 ( .A(\Rx[5] ), .Y(flip6__abc_1243_n12) );
  INVX1 INVX1_24 ( .A(flip7_W1), .Y(flip7__abc_1243_n8) );
  INVX1 INVX1_25 ( .A(\Rx[6] ), .Y(flip7__abc_1243_n12) );
  INVX1 INVX1_26 ( .A(flip8_W1), .Y(flip8__abc_1243_n8) );
  INVX1 INVX1_27 ( .A(\Rx[7] ), .Y(flip8__abc_1243_n12) );
  INVX1 INVX1_28 ( .A(reset), .Y(flipw1__abc_1251_n9_1) );
  INVX1 INVX1_29 ( .A(flip1_W1), .Y(flipw1__abc_1251_n11) );
  INVX1 INVX1_3 ( .A(reset), .Y(_abc_1206_n20) );
  INVX1 INVX1_30 ( .A(reset), .Y(flipw2__abc_1251_n9_1) );
  INVX1 INVX1_31 ( .A(flip2_W1), .Y(flipw2__abc_1251_n11) );
  INVX1 INVX1_32 ( .A(reset), .Y(flipw3__abc_1251_n9_1) );
  INVX1 INVX1_33 ( .A(flip3_W1), .Y(flipw3__abc_1251_n11) );
  INVX1 INVX1_34 ( .A(reset), .Y(flipw4__abc_1251_n9_1) );
  INVX1 INVX1_35 ( .A(flip4_W1), .Y(flipw4__abc_1251_n11) );
  INVX1 INVX1_36 ( .A(reset), .Y(flipw5__abc_1251_n9_1) );
  INVX1 INVX1_37 ( .A(flip5_W1), .Y(flipw5__abc_1251_n11) );
  INVX1 INVX1_38 ( .A(reset), .Y(flipw6__abc_1251_n9_1) );
  INVX1 INVX1_39 ( .A(flip6_W1), .Y(flipw6__abc_1251_n11) );
  INVX1 INVX1_4 ( .A(LRAddress_1_), .Y(_abc_1206_n23) );
  INVX1 INVX1_40 ( .A(reset), .Y(flipw7__abc_1251_n9_1) );
  INVX1 INVX1_41 ( .A(flip7_W1), .Y(flipw7__abc_1251_n11) );
  INVX1 INVX1_42 ( .A(reset), .Y(flipw8__abc_1251_n9_1) );
  INVX1 INVX1_43 ( .A(flip8_W1), .Y(flipw8__abc_1251_n11) );
  INVX1 INVX1_44 ( .A(reset), .Y(latchR__abc_1260_n12) );
  INVX1 INVX1_45 ( .A(ARvalid), .Y(latchR__abc_1260_n14) );
  INVX1 INVX1_46 ( .A(reset), .Y(latchW__abc_1260_n12) );
  INVX1 INVX1_47 ( .A(AWvalid), .Y(latchW__abc_1260_n14) );
  INVX1 INVX1_48 ( .A(maquina_state_0_), .Y(maquina__abc_1272_n35_1) );
  INVX1 INVX1_49 ( .A(reset), .Y(maquina__abc_1272_n38) );
  INVX1 INVX1_5 ( .A(LRAddress_2_), .Y(_abc_1206_n29) );
  INVX1 INVX1_50 ( .A(maquina__abc_1272_n40), .Y(maquina__abc_1272_n41_1) );
  INVX1 INVX1_51 ( .A(maquina_state_5_), .Y(maquina__abc_1272_n46) );
  INVX1 INVX1_52 ( .A(maquina_state_3_), .Y(maquina__abc_1272_n48) );
  INVX1 INVX1_53 ( .A(maquina_state_8_), .Y(maquina__abc_1272_n52) );
  INVX1 INVX1_54 ( .A(Bready), .Y(maquina__abc_1272_n54) );
  INVX1 INVX1_55 ( .A(maquina_state_2_), .Y(maquina__abc_1272_n57) );
  INVX1 INVX1_56 ( .A(maquina_state_4_), .Y(maquina__abc_1272_n58) );
  INVX1 INVX1_57 ( .A(maquina__abc_1272_n61), .Y(maquina__abc_1272_n66) );
  INVX1 INVX1_58 ( .A(maquina__abc_1272_n79), .Y(maquina__abc_1145_n109) );
  INVX1 INVX1_59 ( .A(maquina__abc_1272_n84), .Y(maquina__abc_1145_n112) );
  INVX1 INVX1_6 ( .A(LRAddress_2_), .Y(decor__abc_1225_n13) );
  INVX1 INVX1_7 ( .A(LRAddress_1_), .Y(decor__abc_1225_n17_1) );
  INVX1 INVX1_8 ( .A(LRAddress_0_), .Y(decor__abc_1225_n20) );
  INVX1 INVX1_9 ( .A(LWAddress_2_), .Y(decow__abc_1225_n13) );
  MUX2X1 MUX2X1_1 ( .A(\pindata[6] ), .B(\pindata[4] ), .S(LRAddress_1_), .Y(_abc_1206_n26) );
  MUX2X1 MUX2X1_2 ( .A(\pindata[2] ), .B(\pindata[0] ), .S(LRAddress_1_), .Y(_abc_1206_n32) );
  NAND2X1 NAND2X1_1 ( .A(LRAddress_2_), .B(_abc_1206_n27), .Y(_abc_1206_n28) );
  NAND2X1 NAND2X1_10 ( .A(LWAddress_1_), .B(decow__abc_1225_n20), .Y(decow__abc_1225_n21) );
  NAND2X1 NAND2X1_11 ( .A(LWAddress_0_), .B(LWAddress_1_), .Y(decow__abc_1225_n23) );
  NAND2X1 NAND2X1_12 ( .A(LWAddress_2_), .B(AWready), .Y(decow__abc_1225_n25) );
  NAND2X1 NAND2X1_13 ( .A(flip1_R1), .B(flip1__abc_1243_n8), .Y(flip1__abc_1243_n10_1) );
  NAND2X1 NAND2X1_14 ( .A(flip2_R1), .B(flip2__abc_1243_n8), .Y(flip2__abc_1243_n10_1) );
  NAND2X1 NAND2X1_15 ( .A(flip3_R1), .B(flip3__abc_1243_n8), .Y(flip3__abc_1243_n10_1) );
  NAND2X1 NAND2X1_16 ( .A(flip4_R1), .B(flip4__abc_1243_n8), .Y(flip4__abc_1243_n10_1) );
  NAND2X1 NAND2X1_17 ( .A(flip5_R1), .B(flip5__abc_1243_n8), .Y(flip5__abc_1243_n10_1) );
  NAND2X1 NAND2X1_18 ( .A(flip6_R1), .B(flip6__abc_1243_n8), .Y(flip6__abc_1243_n10_1) );
  NAND2X1 NAND2X1_19 ( .A(flip7_R1), .B(flip7__abc_1243_n8), .Y(flip7__abc_1243_n10_1) );
  NAND2X1 NAND2X1_2 ( .A(_abc_1206_n29), .B(_abc_1206_n33), .Y(_abc_1206_n34_1) );
  NAND2X1 NAND2X1_20 ( .A(flip8_R1), .B(flip8__abc_1243_n8), .Y(flip8__abc_1243_n10_1) );
  NAND2X1 NAND2X1_21 ( .A(\Wdata[0] ), .B(flip1_W1), .Y(flipw1__abc_1251_n10) );
  NAND2X1 NAND2X1_22 ( .A(\datanw[0] ), .B(flipw1__abc_1251_n11), .Y(flipw1__abc_1251_n12) );
  NAND2X1 NAND2X1_23 ( .A(flip1_W1), .B(\Wdata[1] ), .Y(flipw1__abc_1251_n14) );
  NAND2X1 NAND2X1_24 ( .A(\DSE[0] ), .B(flipw1__abc_1251_n11), .Y(flipw1__abc_1251_n15) );
  NAND2X1 NAND2X1_25 ( .A(\Wdata[0] ), .B(flip2_W1), .Y(flipw2__abc_1251_n10) );
  NAND2X1 NAND2X1_26 ( .A(\datanw[1] ), .B(flipw2__abc_1251_n11), .Y(flipw2__abc_1251_n12) );
  NAND2X1 NAND2X1_27 ( .A(flip2_W1), .B(\Wdata[1] ), .Y(flipw2__abc_1251_n14) );
  NAND2X1 NAND2X1_28 ( .A(\DSE[1] ), .B(flipw2__abc_1251_n11), .Y(flipw2__abc_1251_n15) );
  NAND2X1 NAND2X1_29 ( .A(\Wdata[0] ), .B(flip3_W1), .Y(flipw3__abc_1251_n10) );
  NAND2X1 NAND2X1_3 ( .A(ARready), .B(decor__abc_1225_n13), .Y(decor__abc_1225_n14_1) );
  NAND2X1 NAND2X1_30 ( .A(\datanw[2] ), .B(flipw3__abc_1251_n11), .Y(flipw3__abc_1251_n12) );
  NAND2X1 NAND2X1_31 ( .A(flip3_W1), .B(\Wdata[1] ), .Y(flipw3__abc_1251_n14) );
  NAND2X1 NAND2X1_32 ( .A(\DSE[2] ), .B(flipw3__abc_1251_n11), .Y(flipw3__abc_1251_n15) );
  NAND2X1 NAND2X1_33 ( .A(\Wdata[0] ), .B(flip4_W1), .Y(flipw4__abc_1251_n10) );
  NAND2X1 NAND2X1_34 ( .A(\datanw[3] ), .B(flipw4__abc_1251_n11), .Y(flipw4__abc_1251_n12) );
  NAND2X1 NAND2X1_35 ( .A(flip4_W1), .B(\Wdata[1] ), .Y(flipw4__abc_1251_n14) );
  NAND2X1 NAND2X1_36 ( .A(\DSE[3] ), .B(flipw4__abc_1251_n11), .Y(flipw4__abc_1251_n15) );
  NAND2X1 NAND2X1_37 ( .A(\Wdata[0] ), .B(flip5_W1), .Y(flipw5__abc_1251_n10) );
  NAND2X1 NAND2X1_38 ( .A(\datanw[4] ), .B(flipw5__abc_1251_n11), .Y(flipw5__abc_1251_n12) );
  NAND2X1 NAND2X1_39 ( .A(flip5_W1), .B(\Wdata[1] ), .Y(flipw5__abc_1251_n14) );
  NAND2X1 NAND2X1_4 ( .A(LRAddress_0_), .B(decor__abc_1225_n17_1), .Y(decor__abc_1225_n18_1) );
  NAND2X1 NAND2X1_40 ( .A(\DSE[4] ), .B(flipw5__abc_1251_n11), .Y(flipw5__abc_1251_n15) );
  NAND2X1 NAND2X1_41 ( .A(\Wdata[0] ), .B(flip6_W1), .Y(flipw6__abc_1251_n10) );
  NAND2X1 NAND2X1_42 ( .A(\datanw[5] ), .B(flipw6__abc_1251_n11), .Y(flipw6__abc_1251_n12) );
  NAND2X1 NAND2X1_43 ( .A(flip6_W1), .B(\Wdata[1] ), .Y(flipw6__abc_1251_n14) );
  NAND2X1 NAND2X1_44 ( .A(\DSE[5] ), .B(flipw6__abc_1251_n11), .Y(flipw6__abc_1251_n15) );
  NAND2X1 NAND2X1_45 ( .A(\Wdata[0] ), .B(flip7_W1), .Y(flipw7__abc_1251_n10) );
  NAND2X1 NAND2X1_46 ( .A(\datanw[6] ), .B(flipw7__abc_1251_n11), .Y(flipw7__abc_1251_n12) );
  NAND2X1 NAND2X1_47 ( .A(flip7_W1), .B(\Wdata[1] ), .Y(flipw7__abc_1251_n14) );
  NAND2X1 NAND2X1_48 ( .A(\DSE[6] ), .B(flipw7__abc_1251_n11), .Y(flipw7__abc_1251_n15) );
  NAND2X1 NAND2X1_49 ( .A(\Wdata[0] ), .B(flip8_W1), .Y(flipw8__abc_1251_n10) );
  NAND2X1 NAND2X1_5 ( .A(LRAddress_1_), .B(decor__abc_1225_n20), .Y(decor__abc_1225_n21) );
  NAND2X1 NAND2X1_50 ( .A(\datanw[7] ), .B(flipw8__abc_1251_n11), .Y(flipw8__abc_1251_n12) );
  NAND2X1 NAND2X1_51 ( .A(flip8_W1), .B(\Wdata[1] ), .Y(flipw8__abc_1251_n14) );
  NAND2X1 NAND2X1_52 ( .A(\DSE[7] ), .B(flipw8__abc_1251_n11), .Y(flipw8__abc_1251_n15) );
  NAND2X1 NAND2X1_53 ( .A(\RAddress[0] ), .B(ARvalid), .Y(latchR__abc_1260_n13_1) );
  NAND2X1 NAND2X1_54 ( .A(LRAddress_0_), .B(latchR__abc_1260_n14), .Y(latchR__abc_1260_n15) );
  NAND2X1 NAND2X1_55 ( .A(ARvalid), .B(\RAddress[1] ), .Y(latchR__abc_1260_n17) );
  NAND2X1 NAND2X1_56 ( .A(LRAddress_1_), .B(latchR__abc_1260_n14), .Y(latchR__abc_1260_n18) );
  NAND2X1 NAND2X1_57 ( .A(ARvalid), .B(\RAddress[2] ), .Y(latchR__abc_1260_n20) );
  NAND2X1 NAND2X1_58 ( .A(LRAddress_2_), .B(latchR__abc_1260_n14), .Y(latchR__abc_1260_n21) );
  NAND2X1 NAND2X1_59 ( .A(\WAddress[0] ), .B(AWvalid), .Y(latchW__abc_1260_n13_1) );
  NAND2X1 NAND2X1_6 ( .A(LRAddress_0_), .B(LRAddress_1_), .Y(decor__abc_1225_n23) );
  NAND2X1 NAND2X1_60 ( .A(LWAddress_0_), .B(latchW__abc_1260_n14), .Y(latchW__abc_1260_n15) );
  NAND2X1 NAND2X1_61 ( .A(AWvalid), .B(\WAddress[1] ), .Y(latchW__abc_1260_n17) );
  NAND2X1 NAND2X1_62 ( .A(LWAddress_1_), .B(latchW__abc_1260_n14), .Y(latchW__abc_1260_n18) );
  NAND2X1 NAND2X1_63 ( .A(AWvalid), .B(\WAddress[2] ), .Y(latchW__abc_1260_n20) );
  NAND2X1 NAND2X1_64 ( .A(LWAddress_2_), .B(latchW__abc_1260_n14), .Y(latchW__abc_1260_n21) );
  NAND2X1 NAND2X1_65 ( .A(maquina_state_10_), .B(Bready), .Y(maquina__abc_1272_n37_1) );
  NAND2X1 NAND2X1_66 ( .A(maquina__abc_1272_n37_1), .B(maquina__abc_1272_n39), .Y(maquina__abc_1272_n40) );
  NAND2X1 NAND2X1_67 ( .A(reset), .B(maquina_state_2_), .Y(maquina__abc_1272_n43) );
  NAND2X1 NAND2X1_68 ( .A(AWvalid), .B(reset), .Y(maquina__abc_1272_n44_1) );
  NAND2X1 NAND2X1_69 ( .A(reset), .B(maquina_vel), .Y(maquina__abc_1272_n47) );
  NAND2X1 NAND2X1_7 ( .A(LRAddress_2_), .B(ARready), .Y(decor__abc_1225_n25) );
  NAND2X1 NAND2X1_70 ( .A(maquina__abc_1272_n60_1), .B(maquina__abc_1272_n61), .Y(maquina__abc_1272_n62) );
  NAND2X1 NAND2X1_71 ( .A(maquina__abc_1272_n53), .B(maquina__abc_1272_n67_1), .Y(maquina__abc_1272_n69_1) );
  NAND2X1 NAND2X1_72 ( .A(maquina__abc_1272_n73), .B(maquina__abc_1272_n70), .Y(maquina__abc_1272_n74_1) );
  NAND2X1 NAND2X1_8 ( .A(AWready), .B(decow__abc_1225_n13), .Y(decow__abc_1225_n14_1) );
  NAND2X1 NAND2X1_9 ( .A(LWAddress_0_), .B(decow__abc_1225_n17_1), .Y(decow__abc_1225_n18_1) );
  NAND3X1 NAND3X1_1 ( .A(reset), .B(flip1__abc_1243_n10_1), .C(flip1__abc_1243_n9), .Y(flip1_Tx_FF_INPUT) );
  NAND3X1 NAND3X1_10 ( .A(maquina_state_9_), .B(maquina__abc_1272_n48), .C(maquina__abc_1272_n70), .Y(maquina__abc_1272_n71_1) );
  NAND3X1 NAND3X1_11 ( .A(maquina__abc_1272_n53), .B(maquina__abc_1272_n67_1), .C(maquina__abc_1272_n74_1), .Y(maquina__abc_1272_n75) );
  NAND3X1 NAND3X1_12 ( .A(maquina_state_0_), .B(ARvalid), .C(reset), .Y(maquina__abc_1272_n79) );
  NAND3X1 NAND3X1_13 ( .A(reset), .B(maquina_state_2_), .C(Wvalid), .Y(maquina__abc_1272_n84) );
  NAND3X1 NAND3X1_2 ( .A(reset), .B(flip2__abc_1243_n10_1), .C(flip2__abc_1243_n9), .Y(flip2_Tx_FF_INPUT) );
  NAND3X1 NAND3X1_3 ( .A(reset), .B(flip3__abc_1243_n10_1), .C(flip3__abc_1243_n9), .Y(flip3_Tx_FF_INPUT) );
  NAND3X1 NAND3X1_4 ( .A(reset), .B(flip4__abc_1243_n10_1), .C(flip4__abc_1243_n9), .Y(flip4_Tx_FF_INPUT) );
  NAND3X1 NAND3X1_5 ( .A(reset), .B(flip5__abc_1243_n10_1), .C(flip5__abc_1243_n9), .Y(flip5_Tx_FF_INPUT) );
  NAND3X1 NAND3X1_6 ( .A(reset), .B(flip6__abc_1243_n10_1), .C(flip6__abc_1243_n9), .Y(flip6_Tx_FF_INPUT) );
  NAND3X1 NAND3X1_7 ( .A(reset), .B(flip7__abc_1243_n10_1), .C(flip7__abc_1243_n9), .Y(flip7_Tx_FF_INPUT) );
  NAND3X1 NAND3X1_8 ( .A(reset), .B(flip8__abc_1243_n10_1), .C(flip8__abc_1243_n9), .Y(flip8_Tx_FF_INPUT) );
  NAND3X1 NAND3X1_9 ( .A(maquina_state_10_), .B(maquina__abc_1272_n57), .C(maquina__abc_1272_n58), .Y(maquina__abc_1272_n59) );
  NOR2X1 NOR2X1_1 ( .A(\pindata[7] ), .B(_abc_1206_n23), .Y(_abc_1206_n24) );
  NOR2X1 NOR2X1_10 ( .A(decor__abc_1225_n23), .B(decor__abc_1225_n25), .Y(flip8_R1) );
  NOR2X1 NOR2X1_11 ( .A(decow__abc_1225_n15), .B(decow__abc_1225_n14_1), .Y(flip1_W1) );
  NOR2X1 NOR2X1_12 ( .A(decow__abc_1225_n14_1), .B(decow__abc_1225_n18_1), .Y(flip2_W1) );
  NOR2X1 NOR2X1_13 ( .A(decow__abc_1225_n14_1), .B(decow__abc_1225_n21), .Y(flip3_W1) );
  NOR2X1 NOR2X1_14 ( .A(decow__abc_1225_n23), .B(decow__abc_1225_n14_1), .Y(flip4_W1) );
  NOR2X1 NOR2X1_15 ( .A(decow__abc_1225_n25), .B(decow__abc_1225_n15), .Y(flip5_W1) );
  NOR2X1 NOR2X1_16 ( .A(decow__abc_1225_n25), .B(decow__abc_1225_n18_1), .Y(flip6_W1) );
  NOR2X1 NOR2X1_17 ( .A(decow__abc_1225_n25), .B(decow__abc_1225_n21), .Y(flip7_W1) );
  NOR2X1 NOR2X1_18 ( .A(decow__abc_1225_n23), .B(decow__abc_1225_n25), .Y(flip8_W1) );
  NOR2X1 NOR2X1_19 ( .A(maquina_state_10_), .B(maquina_state_4_), .Y(maquina__abc_1272_n53) );
  NOR2X1 NOR2X1_2 ( .A(\pindata[3] ), .B(_abc_1206_n23), .Y(_abc_1206_n30_1) );
  NOR2X1 NOR2X1_20 ( .A(maquina_state_8_), .B(maquina_state_7_), .Y(maquina__abc_1272_n60_1) );
  NOR2X1 NOR2X1_21 ( .A(maquina_state_0_), .B(maquina_state_5_), .Y(maquina__abc_1272_n61) );
  NOR2X1 NOR2X1_22 ( .A(maquina__abc_1272_n59), .B(maquina__abc_1272_n62), .Y(Bvalid) );
  NOR2X1 NOR2X1_23 ( .A(maquina_state_1_), .B(maquina_state_6_), .Y(maquina__abc_1272_n70) );
  NOR2X1 NOR2X1_24 ( .A(maquina_state_9_), .B(maquina_state_3_), .Y(maquina__abc_1272_n73) );
  NOR2X1 NOR2X1_25 ( .A(maquina__abc_1272_n52), .B(maquina__abc_1272_n82), .Y(maquina__abc_1145_n111) );
  NOR2X1 NOR2X1_26 ( .A(maquina__abc_1272_n46), .B(maquina__abc_1272_n82), .Y(maquina__abc_1145_n113) );
  NOR2X1 NOR2X1_3 ( .A(decor__abc_1225_n15), .B(decor__abc_1225_n14_1), .Y(flip1_R1) );
  NOR2X1 NOR2X1_4 ( .A(decor__abc_1225_n14_1), .B(decor__abc_1225_n18_1), .Y(flip2_R1) );
  NOR2X1 NOR2X1_5 ( .A(decor__abc_1225_n14_1), .B(decor__abc_1225_n21), .Y(flip3_R1) );
  NOR2X1 NOR2X1_6 ( .A(decor__abc_1225_n23), .B(decor__abc_1225_n14_1), .Y(flip4_R1) );
  NOR2X1 NOR2X1_7 ( .A(decor__abc_1225_n25), .B(decor__abc_1225_n15), .Y(flip5_R1) );
  NOR2X1 NOR2X1_8 ( .A(decor__abc_1225_n25), .B(decor__abc_1225_n18_1), .Y(flip6_R1) );
  NOR2X1 NOR2X1_9 ( .A(decor__abc_1225_n25), .B(decor__abc_1225_n21), .Y(flip7_R1) );
  NOR3X1 NOR3X1_1 ( .A(maquina_state_2_), .B(maquina_state_8_), .C(maquina_state_7_), .Y(maquina__abc_1272_n67_1) );
  NOR3X1 NOR3X1_2 ( .A(maquina__abc_1272_n66), .B(maquina__abc_1272_n71_1), .C(maquina__abc_1272_n69_1), .Y(Rvalid) );
  OAI21X1 OAI21X1_1 ( .A(_abc_1206_n18), .B(_abc_1206_n19), .C(_abc_1206_n21), .Y(vel_FF_INPUT) );
  OAI21X1 OAI21X1_10 ( .A(flip4_R1), .B(flip4__abc_1243_n8), .C(\Tx[3] ), .Y(flip4__abc_1243_n9) );
  OAI21X1 OAI21X1_11 ( .A(flip4_R1), .B(flip4__abc_1243_n8), .C(reset), .Y(flip4__abc_1243_n13) );
  OAI21X1 OAI21X1_12 ( .A(flip5_R1), .B(flip5__abc_1243_n8), .C(\Tx[4] ), .Y(flip5__abc_1243_n9) );
  OAI21X1 OAI21X1_13 ( .A(flip5_R1), .B(flip5__abc_1243_n8), .C(reset), .Y(flip5__abc_1243_n13) );
  OAI21X1 OAI21X1_14 ( .A(flip6_R1), .B(flip6__abc_1243_n8), .C(\Tx[5] ), .Y(flip6__abc_1243_n9) );
  OAI21X1 OAI21X1_15 ( .A(flip6_R1), .B(flip6__abc_1243_n8), .C(reset), .Y(flip6__abc_1243_n13) );
  OAI21X1 OAI21X1_16 ( .A(flip7_R1), .B(flip7__abc_1243_n8), .C(\Tx[6] ), .Y(flip7__abc_1243_n9) );
  OAI21X1 OAI21X1_17 ( .A(flip7_R1), .B(flip7__abc_1243_n8), .C(reset), .Y(flip7__abc_1243_n13) );
  OAI21X1 OAI21X1_18 ( .A(flip8_R1), .B(flip8__abc_1243_n8), .C(\Tx[7] ), .Y(flip8__abc_1243_n9) );
  OAI21X1 OAI21X1_19 ( .A(flip8_R1), .B(flip8__abc_1243_n8), .C(reset), .Y(flip8__abc_1243_n13) );
  OAI21X1 OAI21X1_2 ( .A(LRAddress_1_), .B(\pindata[5] ), .C(LRAddress_0_), .Y(_abc_1206_n25_1) );
  OAI21X1 OAI21X1_20 ( .A(AWvalid), .B(maquina__abc_1272_n36), .C(maquina__abc_1272_n41_1), .Y(maquina__abc_1145_n9) );
  OAI21X1 OAI21X1_21 ( .A(maquina_state_9_), .B(maquina_state_3_), .C(reset), .Y(maquina__abc_1272_n50) );
  OAI21X1 OAI21X1_22 ( .A(maquina_state_4_), .B(maquina__abc_1272_n54), .C(reset), .Y(maquina__abc_1272_n55_1) );
  OAI21X1 OAI21X1_23 ( .A(maquina__abc_1272_n57), .B(maquina_state_8_), .C(maquina__abc_1272_n61), .Y(maquina__abc_1272_n64) );
  OAI21X1 OAI21X1_3 ( .A(LRAddress_1_), .B(\pindata[1] ), .C(LRAddress_0_), .Y(_abc_1206_n31_1) );
  OAI21X1 OAI21X1_4 ( .A(flip1_R1), .B(flip1__abc_1243_n8), .C(\Tx[0] ), .Y(flip1__abc_1243_n9) );
  OAI21X1 OAI21X1_5 ( .A(flip1_R1), .B(flip1__abc_1243_n8), .C(reset), .Y(flip1__abc_1243_n13) );
  OAI21X1 OAI21X1_6 ( .A(flip2_R1), .B(flip2__abc_1243_n8), .C(\Tx[1] ), .Y(flip2__abc_1243_n9) );
  OAI21X1 OAI21X1_7 ( .A(flip2_R1), .B(flip2__abc_1243_n8), .C(reset), .Y(flip2__abc_1243_n13) );
  OAI21X1 OAI21X1_8 ( .A(flip3_R1), .B(flip3__abc_1243_n8), .C(\Tx[2] ), .Y(flip3__abc_1243_n9) );
  OAI21X1 OAI21X1_9 ( .A(flip3_R1), .B(flip3__abc_1243_n8), .C(reset), .Y(flip3__abc_1243_n13) );
  OAI22X1 OAI22X1_1 ( .A(_abc_1206_n25_1), .B(_abc_1206_n24), .C(LRAddress_0_), .D(_abc_1206_n26), .Y(_abc_1206_n27) );
  OAI22X1 OAI22X1_2 ( .A(_abc_1206_n31_1), .B(_abc_1206_n30_1), .C(LRAddress_0_), .D(_abc_1206_n32), .Y(_abc_1206_n33) );
  OAI22X1 OAI22X1_3 ( .A(Wvalid), .B(maquina__abc_1272_n43), .C(maquina__abc_1272_n44_1), .D(maquina__abc_1272_n36), .Y(maquina__abc_1145_n14) );
  OAI22X1 OAI22X1_4 ( .A(maquina__abc_1272_n46), .B(maquina__abc_1272_n47), .C(maquina__abc_1272_n50), .D(maquina__abc_1272_n49_1), .Y(maquina__abc_1145_n35) );
  OAI22X1 OAI22X1_5 ( .A(maquina__abc_1272_n52), .B(maquina__abc_1272_n47), .C(maquina__abc_1272_n53), .D(maquina__abc_1272_n55_1), .Y(maquina__abc_1145_n45) );
  OR2X2 OR2X2_1 ( .A(LRAddress_0_), .B(LRAddress_1_), .Y(decor__abc_1225_n15) );
  OR2X2 OR2X2_2 ( .A(LWAddress_0_), .B(LWAddress_1_), .Y(decow__abc_1225_n15) );
  OR2X2 OR2X2_3 ( .A(maquina__abc_1272_n35_1), .B(ARvalid), .Y(maquina__abc_1272_n36) );
  OR2X2 OR2X2_4 ( .A(maquina__abc_1272_n38), .B(maquina_vel), .Y(maquina__abc_1272_n82) );
endmodule