module b08_reset(clock, RESET_G, nRESET_G, START, I_7_, I_6_, I_5_, I_4_, I_3_, I_2_, I_1_, I_0_, O_REG_3_, O_REG_2_, O_REG_1_, O_REG_0_);

wire IN_R_REG_0_; 
wire IN_R_REG_1_; 
wire IN_R_REG_2_; 
wire IN_R_REG_3_; 
wire IN_R_REG_4_; 
wire IN_R_REG_5_; 
wire IN_R_REG_6_; 
wire IN_R_REG_7_; 
input I_0_;
input I_1_;
input I_2_;
input I_3_;
input I_4_;
input I_5_;
input I_6_;
input I_7_;
wire MAR_REG_0_; 
wire MAR_REG_1_; 
wire MAR_REG_2_; 
wire OUT_R_REG_0_; 
wire OUT_R_REG_1_; 
wire OUT_R_REG_2_; 
wire OUT_R_REG_3_; 
output O_REG_0_;
output O_REG_1_;
output O_REG_2_;
output O_REG_3_;
input RESET_G;
input START;
wire STATO_REG_0_; 
wire STATO_REG_1_; 
wire _abc_1014_new_n100_; 
wire _abc_1014_new_n101_; 
wire _abc_1014_new_n102_; 
wire _abc_1014_new_n103_; 
wire _abc_1014_new_n104_; 
wire _abc_1014_new_n105_; 
wire _abc_1014_new_n106_; 
wire _abc_1014_new_n107_; 
wire _abc_1014_new_n108_; 
wire _abc_1014_new_n109_; 
wire _abc_1014_new_n110_; 
wire _abc_1014_new_n111_; 
wire _abc_1014_new_n112_; 
wire _abc_1014_new_n113_; 
wire _abc_1014_new_n114_; 
wire _abc_1014_new_n115_; 
wire _abc_1014_new_n116_; 
wire _abc_1014_new_n117_; 
wire _abc_1014_new_n118_; 
wire _abc_1014_new_n119_; 
wire _abc_1014_new_n120_; 
wire _abc_1014_new_n121_; 
wire _abc_1014_new_n122_; 
wire _abc_1014_new_n123_; 
wire _abc_1014_new_n124_; 
wire _abc_1014_new_n125_; 
wire _abc_1014_new_n126_; 
wire _abc_1014_new_n127_; 
wire _abc_1014_new_n128_; 
wire _abc_1014_new_n129_; 
wire _abc_1014_new_n130_; 
wire _abc_1014_new_n131_; 
wire _abc_1014_new_n132_; 
wire _abc_1014_new_n133_; 
wire _abc_1014_new_n134_; 
wire _abc_1014_new_n135_; 
wire _abc_1014_new_n136_; 
wire _abc_1014_new_n137_; 
wire _abc_1014_new_n138_; 
wire _abc_1014_new_n139_; 
wire _abc_1014_new_n140_; 
wire _abc_1014_new_n141_; 
wire _abc_1014_new_n142_; 
wire _abc_1014_new_n143_; 
wire _abc_1014_new_n144_; 
wire _abc_1014_new_n145_; 
wire _abc_1014_new_n146_; 
wire _abc_1014_new_n147_; 
wire _abc_1014_new_n148_; 
wire _abc_1014_new_n149_; 
wire _abc_1014_new_n150_; 
wire _abc_1014_new_n151_; 
wire _abc_1014_new_n152_; 
wire _abc_1014_new_n153_; 
wire _abc_1014_new_n154_; 
wire _abc_1014_new_n155_; 
wire _abc_1014_new_n156_; 
wire _abc_1014_new_n157_; 
wire _abc_1014_new_n158_; 
wire _abc_1014_new_n159_; 
wire _abc_1014_new_n160_; 
wire _abc_1014_new_n161_; 
wire _abc_1014_new_n163_; 
wire _abc_1014_new_n164_; 
wire _abc_1014_new_n165_; 
wire _abc_1014_new_n167_; 
wire _abc_1014_new_n168_; 
wire _abc_1014_new_n169_; 
wire _abc_1014_new_n170_; 
wire _abc_1014_new_n172_; 
wire _abc_1014_new_n173_; 
wire _abc_1014_new_n174_; 
wire _abc_1014_new_n176_; 
wire _abc_1014_new_n177_; 
wire _abc_1014_new_n178_; 
wire _abc_1014_new_n180_; 
wire _abc_1014_new_n181_; 
wire _abc_1014_new_n182_; 
wire _abc_1014_new_n183_; 
wire _abc_1014_new_n185_; 
wire _abc_1014_new_n186_; 
wire _abc_1014_new_n188_; 
wire _abc_1014_new_n189_; 
wire _abc_1014_new_n190_; 
wire _abc_1014_new_n192_; 
wire _abc_1014_new_n193_; 
wire _abc_1014_new_n194_; 
wire _abc_1014_new_n195_; 
wire _abc_1014_new_n196_; 
wire _abc_1014_new_n198_; 
wire _abc_1014_new_n199_; 
wire _abc_1014_new_n200_; 
wire _abc_1014_new_n202_; 
wire _abc_1014_new_n203_; 
wire _abc_1014_new_n204_; 
wire _abc_1014_new_n206_; 
wire _abc_1014_new_n207_; 
wire _abc_1014_new_n208_; 
wire _abc_1014_new_n210_; 
wire _abc_1014_new_n211_; 
wire _abc_1014_new_n212_; 
wire _abc_1014_new_n214_; 
wire _abc_1014_new_n215_; 
wire _abc_1014_new_n216_; 
wire _abc_1014_new_n218_; 
wire _abc_1014_new_n219_; 
wire _abc_1014_new_n220_; 
wire _abc_1014_new_n53_; 
wire _abc_1014_new_n54_; 
wire _abc_1014_new_n55_; 
wire _abc_1014_new_n56_; 
wire _abc_1014_new_n57_; 
wire _abc_1014_new_n58_; 
wire _abc_1014_new_n59_; 
wire _abc_1014_new_n61_; 
wire _abc_1014_new_n62_; 
wire _abc_1014_new_n63_; 
wire _abc_1014_new_n65_; 
wire _abc_1014_new_n66_; 
wire _abc_1014_new_n67_; 
wire _abc_1014_new_n68_; 
wire _abc_1014_new_n69_; 
wire _abc_1014_new_n70_; 
wire _abc_1014_new_n71_; 
wire _abc_1014_new_n72_; 
wire _abc_1014_new_n73_; 
wire _abc_1014_new_n74_; 
wire _abc_1014_new_n76_; 
wire _abc_1014_new_n77_; 
wire _abc_1014_new_n78_; 
wire _abc_1014_new_n80_; 
wire _abc_1014_new_n81_; 
wire _abc_1014_new_n82_; 
wire _abc_1014_new_n84_; 
wire _abc_1014_new_n85_; 
wire _abc_1014_new_n86_; 
wire _abc_1014_new_n88_; 
wire _abc_1014_new_n89_; 
wire _abc_1014_new_n90_; 
wire _abc_1014_new_n91_; 
wire _abc_1014_new_n92_; 
wire _abc_1014_new_n93_; 
wire _abc_1014_new_n94_; 
wire _abc_1014_new_n95_; 
wire _abc_1014_new_n96_; 
wire _abc_1014_new_n97_; 
wire _abc_1014_new_n98_; 
wire _abc_1014_new_n99_; 
input clock;
wire n101; 
wire n106; 
wire n111; 
wire n116; 
wire n121; 
wire n125; 
wire n129; 
wire n32; 
wire n36; 
wire n41; 
wire n46; 
wire n51; 
wire n56; 
wire n61; 
wire n66; 
wire n71; 
wire n76; 
wire n81; 
wire n86; 
wire n91; 
wire n96; 
input nRESET_G;
AND2X2 AND2X2_1 ( .A(_abc_1014_new_n55_), .B(I_1_), .Y(_abc_1014_new_n56_));
AND2X2 AND2X2_10 ( .A(_abc_1014_new_n71_), .B(O_REG_3_), .Y(_abc_1014_new_n72_));
AND2X2 AND2X2_11 ( .A(_abc_1014_new_n70_), .B(OUT_R_REG_3_), .Y(_abc_1014_new_n73_));
AND2X2 AND2X2_12 ( .A(_abc_1014_new_n71_), .B(O_REG_2_), .Y(_abc_1014_new_n76_));
AND2X2 AND2X2_13 ( .A(_abc_1014_new_n70_), .B(OUT_R_REG_2_), .Y(_abc_1014_new_n77_));
AND2X2 AND2X2_14 ( .A(_abc_1014_new_n71_), .B(O_REG_1_), .Y(_abc_1014_new_n80_));
AND2X2 AND2X2_15 ( .A(_abc_1014_new_n70_), .B(OUT_R_REG_1_), .Y(_abc_1014_new_n81_));
AND2X2 AND2X2_16 ( .A(_abc_1014_new_n71_), .B(O_REG_0_), .Y(_abc_1014_new_n84_));
AND2X2 AND2X2_17 ( .A(_abc_1014_new_n70_), .B(OUT_R_REG_0_), .Y(_abc_1014_new_n85_));
AND2X2 AND2X2_18 ( .A(_abc_1014_new_n54_), .B(OUT_R_REG_0_), .Y(_abc_1014_new_n88_));
AND2X2 AND2X2_19 ( .A(_abc_1014_new_n89_), .B(MAR_REG_1_), .Y(_abc_1014_new_n90_));
AND2X2 AND2X2_2 ( .A(_abc_1014_new_n54_), .B(IN_R_REG_1_), .Y(_abc_1014_new_n58_));
AND2X2 AND2X2_20 ( .A(_abc_1014_new_n91_), .B(_abc_1014_new_n92_), .Y(_abc_1014_new_n93_));
AND2X2 AND2X2_21 ( .A(_abc_1014_new_n93_), .B(_abc_1014_new_n89_), .Y(_abc_1014_new_n94_));
AND2X2 AND2X2_22 ( .A(_abc_1014_new_n92_), .B(MAR_REG_0_), .Y(_abc_1014_new_n95_));
AND2X2 AND2X2_23 ( .A(_abc_1014_new_n95_), .B(_abc_1014_new_n91_), .Y(_abc_1014_new_n96_));
AND2X2 AND2X2_24 ( .A(MAR_REG_1_), .B(MAR_REG_0_), .Y(_abc_1014_new_n98_));
AND2X2 AND2X2_25 ( .A(_abc_1014_new_n91_), .B(MAR_REG_2_), .Y(_abc_1014_new_n99_));
AND2X2 AND2X2_26 ( .A(_abc_1014_new_n103_), .B(_abc_1014_new_n104_), .Y(_abc_1014_new_n105_));
AND2X2 AND2X2_27 ( .A(_abc_1014_new_n98_), .B(_abc_1014_new_n92_), .Y(_abc_1014_new_n106_));
AND2X2 AND2X2_28 ( .A(_abc_1014_new_n109_), .B(_abc_1014_new_n101_), .Y(_abc_1014_new_n110_));
AND2X2 AND2X2_29 ( .A(_abc_1014_new_n90_), .B(MAR_REG_2_), .Y(_abc_1014_new_n115_));
AND2X2 AND2X2_3 ( .A(_abc_1014_new_n55_), .B(I_0_), .Y(_abc_1014_new_n61_));
AND2X2 AND2X2_30 ( .A(_abc_1014_new_n116_), .B(_abc_1014_new_n113_), .Y(_abc_1014_new_n117_));
AND2X2 AND2X2_31 ( .A(_abc_1014_new_n118_), .B(_abc_1014_new_n112_), .Y(_abc_1014_new_n119_));
AND2X2 AND2X2_32 ( .A(_abc_1014_new_n99_), .B(_abc_1014_new_n89_), .Y(_abc_1014_new_n120_));
AND2X2 AND2X2_33 ( .A(_abc_1014_new_n91_), .B(MAR_REG_0_), .Y(_abc_1014_new_n122_));
AND2X2 AND2X2_34 ( .A(_abc_1014_new_n125_), .B(_abc_1014_new_n123_), .Y(_abc_1014_new_n126_));
AND2X2 AND2X2_35 ( .A(_abc_1014_new_n127_), .B(_abc_1014_new_n119_), .Y(_abc_1014_new_n128_));
AND2X2 AND2X2_36 ( .A(_abc_1014_new_n128_), .B(_abc_1014_new_n111_), .Y(_abc_1014_new_n129_));
AND2X2 AND2X2_37 ( .A(_abc_1014_new_n132_), .B(_abc_1014_new_n135_), .Y(_abc_1014_new_n136_));
AND2X2 AND2X2_38 ( .A(_abc_1014_new_n140_), .B(_abc_1014_new_n139_), .Y(_abc_1014_new_n141_));
AND2X2 AND2X2_39 ( .A(_abc_1014_new_n106_), .B(_abc_1014_new_n143_), .Y(_abc_1014_new_n144_));
AND2X2 AND2X2_4 ( .A(_abc_1014_new_n54_), .B(IN_R_REG_0_), .Y(_abc_1014_new_n62_));
AND2X2 AND2X2_40 ( .A(_abc_1014_new_n146_), .B(_abc_1014_new_n145_), .Y(_abc_1014_new_n147_));
AND2X2 AND2X2_41 ( .A(_abc_1014_new_n53_), .B(STATO_REG_1_), .Y(_abc_1014_new_n148_));
AND2X2 AND2X2_42 ( .A(_abc_1014_new_n115_), .B(IN_R_REG_5_), .Y(_abc_1014_new_n149_));
AND2X2 AND2X2_43 ( .A(_abc_1014_new_n150_), .B(_abc_1014_new_n148_), .Y(_abc_1014_new_n151_));
AND2X2 AND2X2_44 ( .A(_abc_1014_new_n152_), .B(_abc_1014_new_n104_), .Y(_abc_1014_new_n153_));
AND2X2 AND2X2_45 ( .A(_abc_1014_new_n151_), .B(_abc_1014_new_n154_), .Y(_abc_1014_new_n155_));
AND2X2 AND2X2_46 ( .A(_abc_1014_new_n155_), .B(_abc_1014_new_n147_), .Y(_abc_1014_new_n156_));
AND2X2 AND2X2_47 ( .A(_abc_1014_new_n156_), .B(_abc_1014_new_n142_), .Y(_abc_1014_new_n157_));
AND2X2 AND2X2_48 ( .A(_abc_1014_new_n137_), .B(_abc_1014_new_n157_), .Y(_abc_1014_new_n158_));
AND2X2 AND2X2_49 ( .A(_abc_1014_new_n130_), .B(_abc_1014_new_n158_), .Y(_abc_1014_new_n159_));
AND2X2 AND2X2_5 ( .A(STATO_REG_1_), .B(STATO_REG_0_), .Y(_abc_1014_new_n65_));
AND2X2 AND2X2_50 ( .A(_abc_1014_new_n159_), .B(_abc_1014_new_n90_), .Y(_abc_1014_new_n160_));
AND2X2 AND2X2_51 ( .A(_abc_1014_new_n159_), .B(_abc_1014_new_n121_), .Y(_abc_1014_new_n163_));
AND2X2 AND2X2_52 ( .A(_abc_1014_new_n54_), .B(OUT_R_REG_2_), .Y(_abc_1014_new_n164_));
AND2X2 AND2X2_53 ( .A(_abc_1014_new_n159_), .B(_abc_1014_new_n167_), .Y(_abc_1014_new_n168_));
AND2X2 AND2X2_54 ( .A(_abc_1014_new_n54_), .B(OUT_R_REG_1_), .Y(_abc_1014_new_n169_));
AND2X2 AND2X2_55 ( .A(_abc_1014_new_n159_), .B(_abc_1014_new_n134_), .Y(_abc_1014_new_n172_));
AND2X2 AND2X2_56 ( .A(_abc_1014_new_n54_), .B(OUT_R_REG_3_), .Y(_abc_1014_new_n173_));
AND2X2 AND2X2_57 ( .A(_abc_1014_new_n106_), .B(_abc_1014_new_n65_), .Y(_abc_1014_new_n176_));
AND2X2 AND2X2_58 ( .A(_abc_1014_new_n54_), .B(MAR_REG_2_), .Y(_abc_1014_new_n177_));
AND2X2 AND2X2_59 ( .A(_abc_1014_new_n180_), .B(_abc_1014_new_n54_), .Y(_abc_1014_new_n181_));
AND2X2 AND2X2_6 ( .A(MAR_REG_0_), .B(MAR_REG_2_), .Y(_abc_1014_new_n67_));
AND2X2 AND2X2_60 ( .A(_abc_1014_new_n181_), .B(START), .Y(_abc_1014_new_n182_));
AND2X2 AND2X2_61 ( .A(_abc_1014_new_n71_), .B(_abc_1014_new_n185_), .Y(_abc_1014_new_n186_));
AND2X2 AND2X2_62 ( .A(_abc_1014_new_n181_), .B(MAR_REG_0_), .Y(_abc_1014_new_n188_));
AND2X2 AND2X2_63 ( .A(_abc_1014_new_n65_), .B(_abc_1014_new_n89_), .Y(_abc_1014_new_n189_));
AND2X2 AND2X2_64 ( .A(_abc_1014_new_n54_), .B(MAR_REG_1_), .Y(_abc_1014_new_n193_));
AND2X2 AND2X2_65 ( .A(_abc_1014_new_n192_), .B(_abc_1014_new_n193_), .Y(_abc_1014_new_n194_));
AND2X2 AND2X2_66 ( .A(_abc_1014_new_n122_), .B(_abc_1014_new_n65_), .Y(_abc_1014_new_n195_));
AND2X2 AND2X2_67 ( .A(_abc_1014_new_n55_), .B(I_7_), .Y(_abc_1014_new_n198_));
AND2X2 AND2X2_68 ( .A(_abc_1014_new_n54_), .B(IN_R_REG_7_), .Y(_abc_1014_new_n199_));
AND2X2 AND2X2_69 ( .A(_abc_1014_new_n55_), .B(I_6_), .Y(_abc_1014_new_n202_));
AND2X2 AND2X2_7 ( .A(_abc_1014_new_n67_), .B(MAR_REG_1_), .Y(_abc_1014_new_n68_));
AND2X2 AND2X2_70 ( .A(_abc_1014_new_n54_), .B(IN_R_REG_6_), .Y(_abc_1014_new_n203_));
AND2X2 AND2X2_71 ( .A(_abc_1014_new_n55_), .B(I_5_), .Y(_abc_1014_new_n206_));
AND2X2 AND2X2_72 ( .A(_abc_1014_new_n54_), .B(IN_R_REG_5_), .Y(_abc_1014_new_n207_));
AND2X2 AND2X2_73 ( .A(_abc_1014_new_n55_), .B(I_4_), .Y(_abc_1014_new_n210_));
AND2X2 AND2X2_74 ( .A(_abc_1014_new_n54_), .B(IN_R_REG_4_), .Y(_abc_1014_new_n211_));
AND2X2 AND2X2_75 ( .A(_abc_1014_new_n55_), .B(I_3_), .Y(_abc_1014_new_n214_));
AND2X2 AND2X2_76 ( .A(_abc_1014_new_n54_), .B(IN_R_REG_3_), .Y(_abc_1014_new_n215_));
AND2X2 AND2X2_77 ( .A(_abc_1014_new_n55_), .B(I_2_), .Y(_abc_1014_new_n218_));
AND2X2 AND2X2_78 ( .A(_abc_1014_new_n54_), .B(IN_R_REG_2_), .Y(_abc_1014_new_n219_));
AND2X2 AND2X2_8 ( .A(_abc_1014_new_n68_), .B(_abc_1014_new_n66_), .Y(_abc_1014_new_n69_));
AND2X2 AND2X2_9 ( .A(_abc_1014_new_n69_), .B(_abc_1014_new_n65_), .Y(_abc_1014_new_n70_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n121), .Q(O_REG_3_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(n61), .Q(IN_R_REG_7_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(n66), .Q(IN_R_REG_6_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(n71), .Q(IN_R_REG_5_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(n76), .Q(IN_R_REG_4_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(n81), .Q(IN_R_REG_3_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(n86), .Q(IN_R_REG_2_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(n91), .Q(IN_R_REG_1_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(n96), .Q(IN_R_REG_0_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(n101), .Q(OUT_R_REG_3_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(n106), .Q(OUT_R_REG_2_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n129), .Q(O_REG_1_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(n111), .Q(OUT_R_REG_1_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(n116), .Q(OUT_R_REG_0_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n41), .Q(STATO_REG_0_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n32), .Q(O_REG_0_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n36), .Q(STATO_REG_1_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n125), .Q(O_REG_2_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n46), .Q(MAR_REG_2_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n51), .Q(MAR_REG_1_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(n56), .Q(MAR_REG_0_));
INVX1 INVX1_1 ( .A(STATO_REG_0_), .Y(_abc_1014_new_n53_));
INVX1 INVX1_10 ( .A(_abc_1014_new_n102_), .Y(_abc_1014_new_n103_));
INVX1 INVX1_11 ( .A(IN_R_REG_2_), .Y(_abc_1014_new_n113_));
INVX1 INVX1_12 ( .A(IN_R_REG_1_), .Y(_abc_1014_new_n114_));
INVX1 INVX1_13 ( .A(IN_R_REG_6_), .Y(_abc_1014_new_n133_));
INVX1 INVX1_14 ( .A(IN_R_REG_7_), .Y(_abc_1014_new_n138_));
INVX1 INVX1_15 ( .A(IN_R_REG_4_), .Y(_abc_1014_new_n143_));
INVX1 INVX1_16 ( .A(_abc_1014_new_n144_), .Y(_abc_1014_new_n145_));
INVX1 INVX1_17 ( .A(_abc_1014_new_n149_), .Y(_abc_1014_new_n150_));
INVX1 INVX1_18 ( .A(_abc_1014_new_n93_), .Y(_abc_1014_new_n152_));
INVX1 INVX1_19 ( .A(_abc_1014_new_n67_), .Y(_abc_1014_new_n167_));
INVX1 INVX1_2 ( .A(_abc_1014_new_n54_), .Y(_abc_1014_new_n55_));
INVX1 INVX1_3 ( .A(nRESET_G), .Y(_abc_1014_new_n57_));
INVX1 INVX1_4 ( .A(START), .Y(_abc_1014_new_n66_));
INVX1 INVX1_5 ( .A(_abc_1014_new_n70_), .Y(_abc_1014_new_n71_));
INVX1 INVX1_6 ( .A(MAR_REG_0_), .Y(_abc_1014_new_n89_));
INVX1 INVX1_7 ( .A(MAR_REG_1_), .Y(_abc_1014_new_n91_));
INVX1 INVX1_8 ( .A(MAR_REG_2_), .Y(_abc_1014_new_n92_));
INVX1 INVX1_9 ( .A(IN_R_REG_0_), .Y(_abc_1014_new_n97_));
OR2X2 OR2X2_1 ( .A(_abc_1014_new_n53_), .B(STATO_REG_1_), .Y(_abc_1014_new_n54_));
OR2X2 OR2X2_10 ( .A(_abc_1014_new_n81_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n82_));
OR2X2 OR2X2_11 ( .A(_abc_1014_new_n82_), .B(_abc_1014_new_n80_), .Y(n129));
OR2X2 OR2X2_12 ( .A(_abc_1014_new_n85_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n86_));
OR2X2 OR2X2_13 ( .A(_abc_1014_new_n86_), .B(_abc_1014_new_n84_), .Y(n32));
OR2X2 OR2X2_14 ( .A(_abc_1014_new_n99_), .B(_abc_1014_new_n98_), .Y(_abc_1014_new_n100_));
OR2X2 OR2X2_15 ( .A(_abc_1014_new_n100_), .B(_abc_1014_new_n97_), .Y(_abc_1014_new_n101_));
OR2X2 OR2X2_16 ( .A(_abc_1014_new_n95_), .B(_abc_1014_new_n91_), .Y(_abc_1014_new_n102_));
OR2X2 OR2X2_17 ( .A(_abc_1014_new_n92_), .B(MAR_REG_0_), .Y(_abc_1014_new_n104_));
OR2X2 OR2X2_18 ( .A(_abc_1014_new_n106_), .B(_abc_1014_new_n99_), .Y(_abc_1014_new_n107_));
OR2X2 OR2X2_19 ( .A(_abc_1014_new_n107_), .B(IN_R_REG_1_), .Y(_abc_1014_new_n108_));
OR2X2 OR2X2_2 ( .A(_abc_1014_new_n58_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n59_));
OR2X2 OR2X2_20 ( .A(_abc_1014_new_n105_), .B(_abc_1014_new_n108_), .Y(_abc_1014_new_n109_));
OR2X2 OR2X2_21 ( .A(_abc_1014_new_n110_), .B(_abc_1014_new_n96_), .Y(_abc_1014_new_n111_));
OR2X2 OR2X2_22 ( .A(MAR_REG_1_), .B(IN_R_REG_0_), .Y(_abc_1014_new_n112_));
OR2X2 OR2X2_23 ( .A(_abc_1014_new_n115_), .B(_abc_1014_new_n114_), .Y(_abc_1014_new_n116_));
OR2X2 OR2X2_24 ( .A(_abc_1014_new_n117_), .B(_abc_1014_new_n100_), .Y(_abc_1014_new_n118_));
OR2X2 OR2X2_25 ( .A(_abc_1014_new_n105_), .B(_abc_1014_new_n120_), .Y(_abc_1014_new_n121_));
OR2X2 OR2X2_26 ( .A(_abc_1014_new_n122_), .B(IN_R_REG_7_), .Y(_abc_1014_new_n123_));
OR2X2 OR2X2_27 ( .A(_abc_1014_new_n96_), .B(IN_R_REG_2_), .Y(_abc_1014_new_n124_));
OR2X2 OR2X2_28 ( .A(_abc_1014_new_n124_), .B(_abc_1014_new_n115_), .Y(_abc_1014_new_n125_));
OR2X2 OR2X2_29 ( .A(_abc_1014_new_n126_), .B(_abc_1014_new_n121_), .Y(_abc_1014_new_n127_));
OR2X2 OR2X2_3 ( .A(_abc_1014_new_n59_), .B(_abc_1014_new_n56_), .Y(n91));
OR2X2 OR2X2_30 ( .A(_abc_1014_new_n129_), .B(_abc_1014_new_n94_), .Y(_abc_1014_new_n130_));
OR2X2 OR2X2_31 ( .A(_abc_1014_new_n95_), .B(IN_R_REG_6_), .Y(_abc_1014_new_n131_));
OR2X2 OR2X2_32 ( .A(_abc_1014_new_n121_), .B(_abc_1014_new_n131_), .Y(_abc_1014_new_n132_));
OR2X2 OR2X2_33 ( .A(_abc_1014_new_n107_), .B(_abc_1014_new_n94_), .Y(_abc_1014_new_n134_));
OR2X2 OR2X2_34 ( .A(_abc_1014_new_n134_), .B(_abc_1014_new_n133_), .Y(_abc_1014_new_n135_));
OR2X2 OR2X2_35 ( .A(_abc_1014_new_n136_), .B(_abc_1014_new_n115_), .Y(_abc_1014_new_n137_));
OR2X2 OR2X2_36 ( .A(_abc_1014_new_n90_), .B(_abc_1014_new_n138_), .Y(_abc_1014_new_n139_));
OR2X2 OR2X2_37 ( .A(_abc_1014_new_n103_), .B(IN_R_REG_5_), .Y(_abc_1014_new_n140_));
OR2X2 OR2X2_38 ( .A(_abc_1014_new_n141_), .B(_abc_1014_new_n107_), .Y(_abc_1014_new_n142_));
OR2X2 OR2X2_39 ( .A(_abc_1014_new_n102_), .B(_abc_1014_new_n143_), .Y(_abc_1014_new_n146_));
OR2X2 OR2X2_4 ( .A(_abc_1014_new_n62_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n63_));
OR2X2 OR2X2_40 ( .A(_abc_1014_new_n153_), .B(IN_R_REG_3_), .Y(_abc_1014_new_n154_));
OR2X2 OR2X2_41 ( .A(_abc_1014_new_n160_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n161_));
OR2X2 OR2X2_42 ( .A(_abc_1014_new_n161_), .B(_abc_1014_new_n88_), .Y(n116));
OR2X2 OR2X2_43 ( .A(_abc_1014_new_n164_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n165_));
OR2X2 OR2X2_44 ( .A(_abc_1014_new_n163_), .B(_abc_1014_new_n165_), .Y(n106));
OR2X2 OR2X2_45 ( .A(_abc_1014_new_n169_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n170_));
OR2X2 OR2X2_46 ( .A(_abc_1014_new_n168_), .B(_abc_1014_new_n170_), .Y(n111));
OR2X2 OR2X2_47 ( .A(_abc_1014_new_n172_), .B(_abc_1014_new_n173_), .Y(_abc_1014_new_n174_));
OR2X2 OR2X2_48 ( .A(_abc_1014_new_n161_), .B(_abc_1014_new_n174_), .Y(n101));
OR2X2 OR2X2_49 ( .A(_abc_1014_new_n177_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n178_));
OR2X2 OR2X2_5 ( .A(_abc_1014_new_n63_), .B(_abc_1014_new_n61_), .Y(n96));
OR2X2 OR2X2_50 ( .A(_abc_1014_new_n178_), .B(_abc_1014_new_n176_), .Y(n46));
OR2X2 OR2X2_51 ( .A(_abc_1014_new_n68_), .B(_abc_1014_new_n53_), .Y(_abc_1014_new_n180_));
OR2X2 OR2X2_52 ( .A(_abc_1014_new_n148_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n183_));
OR2X2 OR2X2_53 ( .A(_abc_1014_new_n182_), .B(_abc_1014_new_n183_), .Y(n41));
OR2X2 OR2X2_54 ( .A(STATO_REG_1_), .B(STATO_REG_0_), .Y(_abc_1014_new_n185_));
OR2X2 OR2X2_55 ( .A(_abc_1014_new_n186_), .B(_abc_1014_new_n57_), .Y(n36));
OR2X2 OR2X2_56 ( .A(_abc_1014_new_n189_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n190_));
OR2X2 OR2X2_57 ( .A(_abc_1014_new_n188_), .B(_abc_1014_new_n190_), .Y(n56));
OR2X2 OR2X2_58 ( .A(_abc_1014_new_n180_), .B(_abc_1014_new_n89_), .Y(_abc_1014_new_n192_));
OR2X2 OR2X2_59 ( .A(_abc_1014_new_n195_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n196_));
OR2X2 OR2X2_6 ( .A(_abc_1014_new_n73_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n74_));
OR2X2 OR2X2_60 ( .A(_abc_1014_new_n194_), .B(_abc_1014_new_n196_), .Y(n51));
OR2X2 OR2X2_61 ( .A(_abc_1014_new_n199_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n200_));
OR2X2 OR2X2_62 ( .A(_abc_1014_new_n200_), .B(_abc_1014_new_n198_), .Y(n61));
OR2X2 OR2X2_63 ( .A(_abc_1014_new_n203_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n204_));
OR2X2 OR2X2_64 ( .A(_abc_1014_new_n204_), .B(_abc_1014_new_n202_), .Y(n66));
OR2X2 OR2X2_65 ( .A(_abc_1014_new_n207_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n208_));
OR2X2 OR2X2_66 ( .A(_abc_1014_new_n208_), .B(_abc_1014_new_n206_), .Y(n71));
OR2X2 OR2X2_67 ( .A(_abc_1014_new_n211_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n212_));
OR2X2 OR2X2_68 ( .A(_abc_1014_new_n212_), .B(_abc_1014_new_n210_), .Y(n76));
OR2X2 OR2X2_69 ( .A(_abc_1014_new_n215_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n216_));
OR2X2 OR2X2_7 ( .A(_abc_1014_new_n74_), .B(_abc_1014_new_n72_), .Y(n121));
OR2X2 OR2X2_70 ( .A(_abc_1014_new_n216_), .B(_abc_1014_new_n214_), .Y(n81));
OR2X2 OR2X2_71 ( .A(_abc_1014_new_n219_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n220_));
OR2X2 OR2X2_72 ( .A(_abc_1014_new_n220_), .B(_abc_1014_new_n218_), .Y(n86));
OR2X2 OR2X2_8 ( .A(_abc_1014_new_n77_), .B(_abc_1014_new_n57_), .Y(_abc_1014_new_n78_));
OR2X2 OR2X2_9 ( .A(_abc_1014_new_n78_), .B(_abc_1014_new_n76_), .Y(n125));


endmodule