module spi_axi_master(CEB, SCLK, DATA, RST, CLK, axi_awready, axi_wready, axi_bvalid, axi_arready, axi_rvalid, \axi_rdata[0] , \axi_rdata[1] , \axi_rdata[2] , \axi_rdata[3] , \axi_rdata[4] , \axi_rdata[5] , \axi_rdata[6] , \axi_rdata[7] , \axi_rdata[8] , \axi_rdata[9] , \axi_rdata[10] , \axi_rdata[11] , \axi_rdata[12] , \axi_rdata[13] , \axi_rdata[14] , \axi_rdata[15] , \axi_rdata[16] , \axi_rdata[17] , \axi_rdata[18] , \axi_rdata[19] , \axi_rdata[20] , \axi_rdata[21] , \axi_rdata[22] , \axi_rdata[23] , \axi_rdata[24] , \axi_rdata[25] , \axi_rdata[26] , \axi_rdata[27] , \axi_rdata[28] , \axi_rdata[29] , \axi_rdata[30] , \axi_rdata[31] , DOUT, PICORV_RST, axi_awvalid, \axi_awaddr[0] , \axi_awaddr[1] , \axi_awaddr[2] , \axi_awaddr[3] , \axi_awaddr[4] , \axi_awaddr[5] , \axi_awaddr[6] , \axi_awaddr[7] , \axi_awaddr[8] , \axi_awaddr[9] , \axi_awaddr[10] , \axi_awaddr[11] , \axi_awaddr[12] , \axi_awaddr[13] , \axi_awaddr[14] , \axi_awaddr[15] , \axi_awaddr[16] , \axi_awaddr[17] , \axi_awaddr[18] , \axi_awaddr[19] , \axi_awaddr[20] , \axi_awaddr[21] , \axi_awaddr[22] , \axi_awaddr[23] , \axi_awaddr[24] , \axi_awaddr[25] , \axi_awaddr[26] , \axi_awaddr[27] , \axi_awaddr[28] , \axi_awaddr[29] , \axi_awaddr[30] , \axi_awaddr[31] , \axi_awprot[0] , \axi_awprot[1] , \axi_awprot[2] , axi_wvalid, \axi_wdata[0] , \axi_wdata[1] , \axi_wdata[2] , \axi_wdata[3] , \axi_wdata[4] , \axi_wdata[5] , \axi_wdata[6] , \axi_wdata[7] , \axi_wdata[8] , \axi_wdata[9] , \axi_wdata[10] , \axi_wdata[11] , \axi_wdata[12] , \axi_wdata[13] , \axi_wdata[14] , \axi_wdata[15] , \axi_wdata[16] , \axi_wdata[17] , \axi_wdata[18] , \axi_wdata[19] , \axi_wdata[20] , \axi_wdata[21] , \axi_wdata[22] , \axi_wdata[23] , \axi_wdata[24] , \axi_wdata[25] , \axi_wdata[26] , \axi_wdata[27] , \axi_wdata[28] , \axi_wdata[29] , \axi_wdata[30] , \axi_wdata[31] , \axi_wstrb[0] , \axi_wstrb[1] , \axi_wstrb[2] , \axi_wstrb[3] , axi_bready, axi_arvalid, \axi_araddr[0] , \axi_araddr[1] , \axi_araddr[2] , \axi_araddr[3] , \axi_araddr[4] , \axi_araddr[5] , \axi_araddr[6] , \axi_araddr[7] , \axi_araddr[8] , \axi_araddr[9] , \axi_araddr[10] , \axi_araddr[11] , \axi_araddr[12] , \axi_araddr[13] , \axi_araddr[14] , \axi_araddr[15] , \axi_araddr[16] , \axi_araddr[17] , \axi_araddr[18] , \axi_araddr[19] , \axi_araddr[20] , \axi_araddr[21] , \axi_araddr[22] , \axi_araddr[23] , \axi_araddr[24] , \axi_araddr[25] , \axi_araddr[26] , \axi_araddr[27] , \axi_araddr[28] , \axi_araddr[29] , \axi_araddr[30] , \axi_araddr[31] , \axi_arprot[0] , \axi_arprot[1] , \axi_arprot[2] , axi_rready);
  wire A_ADDR_0_;
  wire A_ADDR_0__FF_INPUT;
  wire A_ADDR_10_;
  wire A_ADDR_10__FF_INPUT;
  wire A_ADDR_11_;
  wire A_ADDR_11__FF_INPUT;
  wire A_ADDR_12_;
  wire A_ADDR_12__FF_INPUT;
  wire A_ADDR_13_;
  wire A_ADDR_13__FF_INPUT;
  wire A_ADDR_14_;
  wire A_ADDR_14__FF_INPUT;
  wire A_ADDR_15_;
  wire A_ADDR_15__FF_INPUT;
  wire A_ADDR_16_;
  wire A_ADDR_16__FF_INPUT;
  wire A_ADDR_17_;
  wire A_ADDR_17__FF_INPUT;
  wire A_ADDR_18_;
  wire A_ADDR_18__FF_INPUT;
  wire A_ADDR_19_;
  wire A_ADDR_19__FF_INPUT;
  wire A_ADDR_1_;
  wire A_ADDR_1__FF_INPUT;
  wire A_ADDR_20_;
  wire A_ADDR_20__FF_INPUT;
  wire A_ADDR_21_;
  wire A_ADDR_21__FF_INPUT;
  wire A_ADDR_22_;
  wire A_ADDR_22__FF_INPUT;
  wire A_ADDR_23_;
  wire A_ADDR_23__FF_INPUT;
  wire A_ADDR_24_;
  wire A_ADDR_24__FF_INPUT;
  wire A_ADDR_25_;
  wire A_ADDR_25__FF_INPUT;
  wire A_ADDR_26_;
  wire A_ADDR_26__FF_INPUT;
  wire A_ADDR_27_;
  wire A_ADDR_27__FF_INPUT;
  wire A_ADDR_28_;
  wire A_ADDR_28__FF_INPUT;
  wire A_ADDR_29_;
  wire A_ADDR_29__FF_INPUT;
  wire A_ADDR_2_;
  wire A_ADDR_2__FF_INPUT;
  wire A_ADDR_30_;
  wire A_ADDR_30__FF_INPUT;
  wire A_ADDR_31_;
  wire A_ADDR_31__FF_INPUT;
  wire A_ADDR_3_;
  wire A_ADDR_3__FF_INPUT;
  wire A_ADDR_4_;
  wire A_ADDR_4__FF_INPUT;
  wire A_ADDR_5_;
  wire A_ADDR_5__FF_INPUT;
  wire A_ADDR_6_;
  wire A_ADDR_6__FF_INPUT;
  wire A_ADDR_7_;
  wire A_ADDR_7__FF_INPUT;
  wire A_ADDR_8_;
  wire A_ADDR_8__FF_INPUT;
  wire A_ADDR_9_;
  wire A_ADDR_9__FF_INPUT;
  input CEB;
  input CLK;
  input DATA;
  output DOUT;
  output PICORV_RST;
  wire PICORV_RST_SPI;
  wire PICORV_RST_SPI_FF_INPUT;
  input RST;
  input SCLK;
  wire WDATA_0_;
  wire WDATA_0__FF_INPUT;
  wire WDATA_10_;
  wire WDATA_10__FF_INPUT;
  wire WDATA_11_;
  wire WDATA_11__FF_INPUT;
  wire WDATA_12_;
  wire WDATA_12__FF_INPUT;
  wire WDATA_13_;
  wire WDATA_13__FF_INPUT;
  wire WDATA_14_;
  wire WDATA_14__FF_INPUT;
  wire WDATA_15_;
  wire WDATA_15__FF_INPUT;
  wire WDATA_16_;
  wire WDATA_16__FF_INPUT;
  wire WDATA_17_;
  wire WDATA_17__FF_INPUT;
  wire WDATA_18_;
  wire WDATA_18__FF_INPUT;
  wire WDATA_19_;
  wire WDATA_19__FF_INPUT;
  wire WDATA_1_;
  wire WDATA_1__FF_INPUT;
  wire WDATA_20_;
  wire WDATA_20__FF_INPUT;
  wire WDATA_21_;
  wire WDATA_21__FF_INPUT;
  wire WDATA_22_;
  wire WDATA_22__FF_INPUT;
  wire WDATA_23_;
  wire WDATA_23__FF_INPUT;
  wire WDATA_24_;
  wire WDATA_24__FF_INPUT;
  wire WDATA_25_;
  wire WDATA_25__FF_INPUT;
  wire WDATA_26_;
  wire WDATA_26__FF_INPUT;
  wire WDATA_27_;
  wire WDATA_27__FF_INPUT;
  wire WDATA_28_;
  wire WDATA_28__FF_INPUT;
  wire WDATA_29_;
  wire WDATA_29__FF_INPUT;
  wire WDATA_2_;
  wire WDATA_2__FF_INPUT;
  wire WDATA_30_;
  wire WDATA_30__FF_INPUT;
  wire WDATA_31_;
  wire WDATA_31__FF_INPUT;
  wire WDATA_3_;
  wire WDATA_3__FF_INPUT;
  wire WDATA_4_;
  wire WDATA_4__FF_INPUT;
  wire WDATA_5_;
  wire WDATA_5__FF_INPUT;
  wire WDATA_6_;
  wire WDATA_6__FF_INPUT;
  wire WDATA_7_;
  wire WDATA_7__FF_INPUT;
  wire WDATA_8_;
  wire WDATA_8__FF_INPUT;
  wire WDATA_9_;
  wire WDATA_9__FF_INPUT;
  wire _abc_2913_n1025;
  wire _abc_2913_n1036;
  wire _abc_2913_n105;
  wire _abc_2913_n116;
  wire _abc_2913_n129;
  wire _abc_2913_n70;
  wire _abc_2913_n78;
  wire _abc_2913_n87;
  wire _abc_2913_n95;
  wire _abc_4108_n1001;
  wire _abc_4108_n1002;
  wire _abc_4108_n1004;
  wire _abc_4108_n1005;
  wire _abc_4108_n1007;
  wire _abc_4108_n1008;
  wire _abc_4108_n1010;
  wire _abc_4108_n1011;
  wire _abc_4108_n1013;
  wire _abc_4108_n1014;
  wire _abc_4108_n1016;
  wire _abc_4108_n1017;
  wire _abc_4108_n1019;
  wire _abc_4108_n1020;
  wire _abc_4108_n1022;
  wire _abc_4108_n1023;
  wire _abc_4108_n1025;
  wire _abc_4108_n1026;
  wire _abc_4108_n1028;
  wire _abc_4108_n1029;
  wire _abc_4108_n1031;
  wire _abc_4108_n1032;
  wire _abc_4108_n1034;
  wire _abc_4108_n1035;
  wire _abc_4108_n1037;
  wire _abc_4108_n1038;
  wire _abc_4108_n1040;
  wire _abc_4108_n1041;
  wire _abc_4108_n1043;
  wire _abc_4108_n1044;
  wire _abc_4108_n1046;
  wire _abc_4108_n1047;
  wire _abc_4108_n1049;
  wire _abc_4108_n1050;
  wire _abc_4108_n1052;
  wire _abc_4108_n1053;
  wire _abc_4108_n1054;
  wire _abc_4108_n1055;
  wire _abc_4108_n1056;
  wire _abc_4108_n1057;
  wire _abc_4108_n1059;
  wire _abc_4108_n1060;
  wire _abc_4108_n1062;
  wire _abc_4108_n1063;
  wire _abc_4108_n1065;
  wire _abc_4108_n1066;
  wire _abc_4108_n1068;
  wire _abc_4108_n1069;
  wire _abc_4108_n1071;
  wire _abc_4108_n1072;
  wire _abc_4108_n1074;
  wire _abc_4108_n1075;
  wire _abc_4108_n1077;
  wire _abc_4108_n1078;
  wire _abc_4108_n1080;
  wire _abc_4108_n1081;
  wire _abc_4108_n1083;
  wire _abc_4108_n1084;
  wire _abc_4108_n1086;
  wire _abc_4108_n1087;
  wire _abc_4108_n1089;
  wire _abc_4108_n1090;
  wire _abc_4108_n1092;
  wire _abc_4108_n1093;
  wire _abc_4108_n1095;
  wire _abc_4108_n1096;
  wire _abc_4108_n1098;
  wire _abc_4108_n1099;
  wire _abc_4108_n1101;
  wire _abc_4108_n1102;
  wire _abc_4108_n1104;
  wire _abc_4108_n1105;
  wire _abc_4108_n1107;
  wire _abc_4108_n1108;
  wire _abc_4108_n1110;
  wire _abc_4108_n1111;
  wire _abc_4108_n1113;
  wire _abc_4108_n1114;
  wire _abc_4108_n1116;
  wire _abc_4108_n1117;
  wire _abc_4108_n1119;
  wire _abc_4108_n1120;
  wire _abc_4108_n1122;
  wire _abc_4108_n1123;
  wire _abc_4108_n1125;
  wire _abc_4108_n1126;
  wire _abc_4108_n1128;
  wire _abc_4108_n1129;
  wire _abc_4108_n1131;
  wire _abc_4108_n1132;
  wire _abc_4108_n1134;
  wire _abc_4108_n1135;
  wire _abc_4108_n1137;
  wire _abc_4108_n1138;
  wire _abc_4108_n1140;
  wire _abc_4108_n1141;
  wire _abc_4108_n1143;
  wire _abc_4108_n1144;
  wire _abc_4108_n1146;
  wire _abc_4108_n1147;
  wire _abc_4108_n1149;
  wire _abc_4108_n1150;
  wire _abc_4108_n1152;
  wire _abc_4108_n1154;
  wire _abc_4108_n1156;
  wire _abc_4108_n1158;
  wire _abc_4108_n1160;
  wire _abc_4108_n1162;
  wire _abc_4108_n1164;
  wire _abc_4108_n1166;
  wire _abc_4108_n1168;
  wire _abc_4108_n1170;
  wire _abc_4108_n1172;
  wire _abc_4108_n1174;
  wire _abc_4108_n1176;
  wire _abc_4108_n1178;
  wire _abc_4108_n1180;
  wire _abc_4108_n1182;
  wire _abc_4108_n1184;
  wire _abc_4108_n1186;
  wire _abc_4108_n1188;
  wire _abc_4108_n1190;
  wire _abc_4108_n1192;
  wire _abc_4108_n1194;
  wire _abc_4108_n1196;
  wire _abc_4108_n1198;
  wire _abc_4108_n1200;
  wire _abc_4108_n1202;
  wire _abc_4108_n1204;
  wire _abc_4108_n1206;
  wire _abc_4108_n1208;
  wire _abc_4108_n1210;
  wire _abc_4108_n1212;
  wire _abc_4108_n1215;
  wire _abc_4108_n1221;
  wire _abc_4108_n1225;
  wire _abc_4108_n1228;
  wire _abc_4108_n1230;
  wire _abc_4108_n1232;
  wire _abc_4108_n1234;
  wire _abc_4108_n1236;
  wire _abc_4108_n1238;
  wire _abc_4108_n1240;
  wire _abc_4108_n1242;
  wire _abc_4108_n1246;
  wire _abc_4108_n1248;
  wire _abc_4108_n1250;
  wire _abc_4108_n1252;
  wire _abc_4108_n1254;
  wire _abc_4108_n1257;
  wire _abc_4108_n1259;
  wire _abc_4108_n1261;
  wire _abc_4108_n1264;
  wire _abc_4108_n1266;
  wire _abc_4108_n1268;
  wire _abc_4108_n1271;
  wire _abc_4108_n1273;
  wire _abc_4108_n1275;
  wire _abc_4108_n1277;
  wire _abc_4108_n1279;
  wire _abc_4108_n1281;
  wire _abc_4108_n1283;
  wire _abc_4108_n1285;
  wire _abc_4108_n1287;
  wire _abc_4108_n1289;
  wire _abc_4108_n1291;
  wire _abc_4108_n1293;
  wire _abc_4108_n1295;
  wire _abc_4108_n1297;
  wire _abc_4108_n1299;
  wire _abc_4108_n1301;
  wire _abc_4108_n1303;
  wire _abc_4108_n1305;
  wire _abc_4108_n1307;
  wire _abc_4108_n1309;
  wire _abc_4108_n1311;
  wire _abc_4108_n1313;
  wire _abc_4108_n1315;
  wire _abc_4108_n1317;
  wire _abc_4108_n1319;
  wire _abc_4108_n1321;
  wire _abc_4108_n1323;
  wire _abc_4108_n1325;
  wire _abc_4108_n1327;
  wire _abc_4108_n1329;
  wire _abc_4108_n1331;
  wire _abc_4108_n1333;
  wire _abc_4108_n1334;
  wire _abc_4108_n1335;
  wire _abc_4108_n1336;
  wire _abc_4108_n1338;
  wire _abc_4108_n1339;
  wire _abc_4108_n1341;
  wire _abc_4108_n1343;
  wire _abc_4108_n1345;
  wire _abc_4108_n558_1;
  wire _abc_4108_n559_1;
  wire _abc_4108_n561;
  wire _abc_4108_n562_1;
  wire _abc_4108_n563_1;
  wire _abc_4108_n565;
  wire _abc_4108_n566;
  wire _abc_4108_n568_1;
  wire _abc_4108_n569_1;
  wire _abc_4108_n570;
  wire _abc_4108_n571;
  wire _abc_4108_n572_1;
  wire _abc_4108_n573_1;
  wire _abc_4108_n575;
  wire _abc_4108_n576;
  wire _abc_4108_n577_1;
  wire _abc_4108_n579_1;
  wire _abc_4108_n580;
  wire _abc_4108_n582_1;
  wire _abc_4108_n583_1;
  wire _abc_4108_n584_1;
  wire _abc_4108_n586;
  wire _abc_4108_n587_1;
  wire _abc_4108_n590;
  wire _abc_4108_n591;
  wire _abc_4108_n593_1;
  wire _abc_4108_n595;
  wire _abc_4108_n596;
  wire _abc_4108_n597_1;
  wire _abc_4108_n598_1;
  wire _abc_4108_n599_1;
  wire _abc_4108_n600;
  wire _abc_4108_n601;
  wire _abc_4108_n602_1;
  wire _abc_4108_n603_1;
  wire _abc_4108_n604_1;
  wire _abc_4108_n605;
  wire _abc_4108_n606;
  wire _abc_4108_n607_1;
  wire _abc_4108_n608_1;
  wire _abc_4108_n609_1;
  wire _abc_4108_n610;
  wire _abc_4108_n611;
  wire _abc_4108_n612_1;
  wire _abc_4108_n613_1;
  wire _abc_4108_n614_1;
  wire _abc_4108_n615;
  wire _abc_4108_n616;
  wire _abc_4108_n617_1;
  wire _abc_4108_n618_1;
  wire _abc_4108_n619_1;
  wire _abc_4108_n620;
  wire _abc_4108_n621;
  wire _abc_4108_n622_1;
  wire _abc_4108_n623_1;
  wire _abc_4108_n624_1;
  wire _abc_4108_n625;
  wire _abc_4108_n626;
  wire _abc_4108_n627_1;
  wire _abc_4108_n628;
  wire _abc_4108_n629;
  wire _abc_4108_n630_1;
  wire _abc_4108_n631;
  wire _abc_4108_n632;
  wire _abc_4108_n633_1;
  wire _abc_4108_n634_1;
  wire _abc_4108_n635;
  wire _abc_4108_n636;
  wire _abc_4108_n637_1;
  wire _abc_4108_n638_1;
  wire _abc_4108_n639;
  wire _abc_4108_n640;
  wire _abc_4108_n641_1;
  wire _abc_4108_n642_1;
  wire _abc_4108_n643;
  wire _abc_4108_n644;
  wire _abc_4108_n646_1;
  wire _abc_4108_n647;
  wire _abc_4108_n648;
  wire _abc_4108_n649_1;
  wire _abc_4108_n650_1;
  wire _abc_4108_n652;
  wire _abc_4108_n653_1;
  wire _abc_4108_n654_1;
  wire _abc_4108_n655;
  wire _abc_4108_n656;
  wire _abc_4108_n657_1;
  wire _abc_4108_n658_1;
  wire _abc_4108_n660;
  wire _abc_4108_n661_1;
  wire _abc_4108_n662_1;
  wire _abc_4108_n663;
  wire _abc_4108_n664;
  wire _abc_4108_n665_1;
  wire _abc_4108_n666_1;
  wire _abc_4108_n667;
  wire _abc_4108_n668;
  wire _abc_4108_n669_1;
  wire _abc_4108_n670_1;
  wire _abc_4108_n671;
  wire _abc_4108_n672;
  wire _abc_4108_n673_1;
  wire _abc_4108_n674_1;
  wire _abc_4108_n675;
  wire _abc_4108_n676;
  wire _abc_4108_n677_1;
  wire _abc_4108_n678_1;
  wire _abc_4108_n679;
  wire _abc_4108_n680;
  wire _abc_4108_n681_1;
  wire _abc_4108_n682_1;
  wire _abc_4108_n683;
  wire _abc_4108_n684;
  wire _abc_4108_n685_1;
  wire _abc_4108_n686_1;
  wire _abc_4108_n687;
  wire _abc_4108_n688;
  wire _abc_4108_n690_1;
  wire _abc_4108_n691;
  wire _abc_4108_n692;
  wire _abc_4108_n693_1;
  wire _abc_4108_n694_1;
  wire _abc_4108_n696;
  wire _abc_4108_n697_1;
  wire _abc_4108_n698_1;
  wire _abc_4108_n699;
  wire _abc_4108_n700;
  wire _abc_4108_n702_1;
  wire _abc_4108_n703;
  wire _abc_4108_n704;
  wire _abc_4108_n705_1;
  wire _abc_4108_n706_1;
  wire _abc_4108_n708;
  wire _abc_4108_n709_1;
  wire _abc_4108_n710_1;
  wire _abc_4108_n711;
  wire _abc_4108_n712;
  wire _abc_4108_n714_1;
  wire _abc_4108_n715;
  wire _abc_4108_n716;
  wire _abc_4108_n717_1;
  wire _abc_4108_n718_1;
  wire _abc_4108_n720;
  wire _abc_4108_n721_1;
  wire _abc_4108_n722_1;
  wire _abc_4108_n723;
  wire _abc_4108_n724;
  wire _abc_4108_n726_1;
  wire _abc_4108_n727;
  wire _abc_4108_n728;
  wire _abc_4108_n729_1;
  wire _abc_4108_n730_1;
  wire _abc_4108_n732;
  wire _abc_4108_n733_1;
  wire _abc_4108_n734_1;
  wire _abc_4108_n735;
  wire _abc_4108_n736;
  wire _abc_4108_n738_1;
  wire _abc_4108_n739;
  wire _abc_4108_n740;
  wire _abc_4108_n741_1;
  wire _abc_4108_n742_1;
  wire _abc_4108_n744;
  wire _abc_4108_n745_1;
  wire _abc_4108_n746_1;
  wire _abc_4108_n747;
  wire _abc_4108_n748;
  wire _abc_4108_n750_1;
  wire _abc_4108_n751;
  wire _abc_4108_n752;
  wire _abc_4108_n753_1;
  wire _abc_4108_n754_1;
  wire _abc_4108_n756;
  wire _abc_4108_n757_1;
  wire _abc_4108_n758;
  wire _abc_4108_n759_1;
  wire _abc_4108_n760;
  wire _abc_4108_n762;
  wire _abc_4108_n763_1;
  wire _abc_4108_n764;
  wire _abc_4108_n765_1;
  wire _abc_4108_n766;
  wire _abc_4108_n768;
  wire _abc_4108_n769_1;
  wire _abc_4108_n770;
  wire _abc_4108_n771_1;
  wire _abc_4108_n772;
  wire _abc_4108_n774;
  wire _abc_4108_n775_1;
  wire _abc_4108_n776;
  wire _abc_4108_n777_1;
  wire _abc_4108_n778;
  wire _abc_4108_n780;
  wire _abc_4108_n781_1;
  wire _abc_4108_n782;
  wire _abc_4108_n783_1;
  wire _abc_4108_n784;
  wire _abc_4108_n786;
  wire _abc_4108_n787_1;
  wire _abc_4108_n788;
  wire _abc_4108_n789_1;
  wire _abc_4108_n790;
  wire _abc_4108_n792;
  wire _abc_4108_n793_1;
  wire _abc_4108_n794;
  wire _abc_4108_n795_1;
  wire _abc_4108_n796;
  wire _abc_4108_n798;
  wire _abc_4108_n799_1;
  wire _abc_4108_n800;
  wire _abc_4108_n801_1;
  wire _abc_4108_n802;
  wire _abc_4108_n804;
  wire _abc_4108_n805_1;
  wire _abc_4108_n806;
  wire _abc_4108_n807_1;
  wire _abc_4108_n808;
  wire _abc_4108_n810;
  wire _abc_4108_n811_1;
  wire _abc_4108_n812;
  wire _abc_4108_n813_1;
  wire _abc_4108_n814;
  wire _abc_4108_n816;
  wire _abc_4108_n817_1;
  wire _abc_4108_n818;
  wire _abc_4108_n819_1;
  wire _abc_4108_n820_1;
  wire _abc_4108_n822;
  wire _abc_4108_n823_1;
  wire _abc_4108_n824_1;
  wire _abc_4108_n825_1;
  wire _abc_4108_n826;
  wire _abc_4108_n828;
  wire _abc_4108_n829_1;
  wire _abc_4108_n830;
  wire _abc_4108_n831_1;
  wire _abc_4108_n832;
  wire _abc_4108_n834;
  wire _abc_4108_n835_1;
  wire _abc_4108_n836;
  wire _abc_4108_n837_1;
  wire _abc_4108_n838;
  wire _abc_4108_n840;
  wire _abc_4108_n841_1;
  wire _abc_4108_n842;
  wire _abc_4108_n843_1;
  wire _abc_4108_n844;
  wire _abc_4108_n846;
  wire _abc_4108_n847_1;
  wire _abc_4108_n848;
  wire _abc_4108_n849_1;
  wire _abc_4108_n850;
  wire _abc_4108_n852;
  wire _abc_4108_n853_1;
  wire _abc_4108_n854;
  wire _abc_4108_n855_1;
  wire _abc_4108_n856;
  wire _abc_4108_n858;
  wire _abc_4108_n859_1;
  wire _abc_4108_n861_1;
  wire _abc_4108_n862;
  wire _abc_4108_n864;
  wire _abc_4108_n865_1;
  wire _abc_4108_n867_1;
  wire _abc_4108_n868;
  wire _abc_4108_n870;
  wire _abc_4108_n871_1;
  wire _abc_4108_n873_1;
  wire _abc_4108_n874;
  wire _abc_4108_n876;
  wire _abc_4108_n877_1;
  wire _abc_4108_n879_1;
  wire _abc_4108_n880;
  wire _abc_4108_n882;
  wire _abc_4108_n883_1;
  wire _abc_4108_n885_1;
  wire _abc_4108_n886;
  wire _abc_4108_n888;
  wire _abc_4108_n889_1;
  wire _abc_4108_n891_1;
  wire _abc_4108_n892_1;
  wire _abc_4108_n894_1;
  wire _abc_4108_n895_1;
  wire _abc_4108_n897_1;
  wire _abc_4108_n898_1;
  wire _abc_4108_n900_1;
  wire _abc_4108_n901_1;
  wire _abc_4108_n903_1;
  wire _abc_4108_n904_1;
  wire _abc_4108_n906_1;
  wire _abc_4108_n907_1;
  wire _abc_4108_n909_1;
  wire _abc_4108_n910_1;
  wire _abc_4108_n912_1;
  wire _abc_4108_n913_1;
  wire _abc_4108_n915_1;
  wire _abc_4108_n916_1;
  wire _abc_4108_n918_1;
  wire _abc_4108_n919_1;
  wire _abc_4108_n921_1;
  wire _abc_4108_n922_1;
  wire _abc_4108_n924_1;
  wire _abc_4108_n925_1;
  wire _abc_4108_n927_1;
  wire _abc_4108_n928_1;
  wire _abc_4108_n930_1;
  wire _abc_4108_n931_1;
  wire _abc_4108_n933_1;
  wire _abc_4108_n934_1;
  wire _abc_4108_n936_1;
  wire _abc_4108_n937_1;
  wire _abc_4108_n939_1;
  wire _abc_4108_n940_1;
  wire _abc_4108_n942_1;
  wire _abc_4108_n943_1;
  wire _abc_4108_n945_1;
  wire _abc_4108_n946_1;
  wire _abc_4108_n948_1;
  wire _abc_4108_n949_1;
  wire _abc_4108_n951_1;
  wire _abc_4108_n952;
  wire _abc_4108_n954;
  wire _abc_4108_n955_1;
  wire _abc_4108_n956;
  wire _abc_4108_n957;
  wire _abc_4108_n959;
  wire _abc_4108_n960;
  wire _abc_4108_n962;
  wire _abc_4108_n963_1;
  wire _abc_4108_n965;
  wire _abc_4108_n966_1;
  wire _abc_4108_n968_1;
  wire _abc_4108_n969_1;
  wire _abc_4108_n971;
  wire _abc_4108_n972;
  wire _abc_4108_n974;
  wire _abc_4108_n975;
  wire _abc_4108_n977;
  wire _abc_4108_n978;
  wire _abc_4108_n980;
  wire _abc_4108_n981;
  wire _abc_4108_n983;
  wire _abc_4108_n984;
  wire _abc_4108_n986;
  wire _abc_4108_n987;
  wire _abc_4108_n989;
  wire _abc_4108_n990;
  wire _abc_4108_n992;
  wire _abc_4108_n993;
  wire _abc_4108_n995;
  wire _abc_4108_n996;
  wire _abc_4108_n998;
  wire _abc_4108_n999;
  output \axi_araddr[0] ;
  output \axi_araddr[10] ;
  output \axi_araddr[11] ;
  output \axi_araddr[12] ;
  output \axi_araddr[13] ;
  output \axi_araddr[14] ;
  output \axi_araddr[15] ;
  output \axi_araddr[16] ;
  output \axi_araddr[17] ;
  output \axi_araddr[18] ;
  output \axi_araddr[19] ;
  output \axi_araddr[1] ;
  output \axi_araddr[20] ;
  output \axi_araddr[21] ;
  output \axi_araddr[22] ;
  output \axi_araddr[23] ;
  output \axi_araddr[24] ;
  output \axi_araddr[25] ;
  output \axi_araddr[26] ;
  output \axi_araddr[27] ;
  output \axi_araddr[28] ;
  output \axi_araddr[29] ;
  output \axi_araddr[2] ;
  output \axi_araddr[30] ;
  output \axi_araddr[31] ;
  output \axi_araddr[3] ;
  output \axi_araddr[4] ;
  output \axi_araddr[5] ;
  output \axi_araddr[6] ;
  output \axi_araddr[7] ;
  output \axi_araddr[8] ;
  output \axi_araddr[9] ;
  output \axi_arprot[0] ;
  output \axi_arprot[1] ;
  output \axi_arprot[2] ;
  input axi_arready;
  output axi_arvalid;
  output \axi_awaddr[0] ;
  output \axi_awaddr[10] ;
  output \axi_awaddr[11] ;
  output \axi_awaddr[12] ;
  output \axi_awaddr[13] ;
  output \axi_awaddr[14] ;
  output \axi_awaddr[15] ;
  output \axi_awaddr[16] ;
  output \axi_awaddr[17] ;
  output \axi_awaddr[18] ;
  output \axi_awaddr[19] ;
  output \axi_awaddr[1] ;
  output \axi_awaddr[20] ;
  output \axi_awaddr[21] ;
  output \axi_awaddr[22] ;
  output \axi_awaddr[23] ;
  output \axi_awaddr[24] ;
  output \axi_awaddr[25] ;
  output \axi_awaddr[26] ;
  output \axi_awaddr[27] ;
  output \axi_awaddr[28] ;
  output \axi_awaddr[29] ;
  output \axi_awaddr[2] ;
  output \axi_awaddr[30] ;
  output \axi_awaddr[31] ;
  output \axi_awaddr[3] ;
  output \axi_awaddr[4] ;
  output \axi_awaddr[5] ;
  output \axi_awaddr[6] ;
  output \axi_awaddr[7] ;
  output \axi_awaddr[8] ;
  output \axi_awaddr[9] ;
  output \axi_awprot[0] ;
  output \axi_awprot[1] ;
  output \axi_awprot[2] ;
  input axi_awready;
  output axi_awvalid;
  output axi_bready;
  input axi_bvalid;
  input \axi_rdata[0] ;
  input \axi_rdata[10] ;
  input \axi_rdata[11] ;
  input \axi_rdata[12] ;
  input \axi_rdata[13] ;
  input \axi_rdata[14] ;
  input \axi_rdata[15] ;
  input \axi_rdata[16] ;
  input \axi_rdata[17] ;
  input \axi_rdata[18] ;
  input \axi_rdata[19] ;
  input \axi_rdata[1] ;
  input \axi_rdata[20] ;
  input \axi_rdata[21] ;
  input \axi_rdata[22] ;
  input \axi_rdata[23] ;
  input \axi_rdata[24] ;
  input \axi_rdata[25] ;
  input \axi_rdata[26] ;
  input \axi_rdata[27] ;
  input \axi_rdata[28] ;
  input \axi_rdata[29] ;
  input \axi_rdata[2] ;
  input \axi_rdata[30] ;
  input \axi_rdata[31] ;
  input \axi_rdata[3] ;
  input \axi_rdata[4] ;
  input \axi_rdata[5] ;
  input \axi_rdata[6] ;
  input \axi_rdata[7] ;
  input \axi_rdata[8] ;
  input \axi_rdata[9] ;
  output axi_rready;
  input axi_rvalid;
  output \axi_wdata[0] ;
  output \axi_wdata[10] ;
  output \axi_wdata[11] ;
  output \axi_wdata[12] ;
  output \axi_wdata[13] ;
  output \axi_wdata[14] ;
  output \axi_wdata[15] ;
  output \axi_wdata[16] ;
  output \axi_wdata[17] ;
  output \axi_wdata[18] ;
  output \axi_wdata[19] ;
  output \axi_wdata[1] ;
  output \axi_wdata[20] ;
  output \axi_wdata[21] ;
  output \axi_wdata[22] ;
  output \axi_wdata[23] ;
  output \axi_wdata[24] ;
  output \axi_wdata[25] ;
  output \axi_wdata[26] ;
  output \axi_wdata[27] ;
  output \axi_wdata[28] ;
  output \axi_wdata[29] ;
  output \axi_wdata[2] ;
  output \axi_wdata[30] ;
  output \axi_wdata[31] ;
  output \axi_wdata[3] ;
  output \axi_wdata[4] ;
  output \axi_wdata[5] ;
  output \axi_wdata[6] ;
  output \axi_wdata[7] ;
  output \axi_wdata[8] ;
  output \axi_wdata[9] ;
  input axi_wready;
  output \axi_wstrb[0] ;
  output \axi_wstrb[1] ;
  output \axi_wstrb[2] ;
  output \axi_wstrb[3] ;
  output axi_wvalid;
  wire bus_cap_0_;
  wire bus_cap_0__FF_INPUT;
  wire bus_cap_10_;
  wire bus_cap_10__FF_INPUT;
  wire bus_cap_11_;
  wire bus_cap_11__FF_INPUT;
  wire bus_cap_12_;
  wire bus_cap_12__FF_INPUT;
  wire bus_cap_13_;
  wire bus_cap_13__FF_INPUT;
  wire bus_cap_14_;
  wire bus_cap_14__FF_INPUT;
  wire bus_cap_15_;
  wire bus_cap_15__FF_INPUT;
  wire bus_cap_16_;
  wire bus_cap_16__FF_INPUT;
  wire bus_cap_17_;
  wire bus_cap_17__FF_INPUT;
  wire bus_cap_18_;
  wire bus_cap_18__FF_INPUT;
  wire bus_cap_19_;
  wire bus_cap_19__FF_INPUT;
  wire bus_cap_1_;
  wire bus_cap_1__FF_INPUT;
  wire bus_cap_20_;
  wire bus_cap_20__FF_INPUT;
  wire bus_cap_21_;
  wire bus_cap_21__FF_INPUT;
  wire bus_cap_22_;
  wire bus_cap_22__FF_INPUT;
  wire bus_cap_23_;
  wire bus_cap_23__FF_INPUT;
  wire bus_cap_24_;
  wire bus_cap_24__FF_INPUT;
  wire bus_cap_25_;
  wire bus_cap_25__FF_INPUT;
  wire bus_cap_26_;
  wire bus_cap_26__FF_INPUT;
  wire bus_cap_27_;
  wire bus_cap_27__FF_INPUT;
  wire bus_cap_28_;
  wire bus_cap_28__FF_INPUT;
  wire bus_cap_29_;
  wire bus_cap_29__FF_INPUT;
  wire bus_cap_2_;
  wire bus_cap_2__FF_INPUT;
  wire bus_cap_30_;
  wire bus_cap_30__FF_INPUT;
  wire bus_cap_31__FF_INPUT;
  wire bus_cap_3_;
  wire bus_cap_3__FF_INPUT;
  wire bus_cap_4_;
  wire bus_cap_4__FF_INPUT;
  wire bus_cap_5_;
  wire bus_cap_5__FF_INPUT;
  wire bus_cap_6_;
  wire bus_cap_6__FF_INPUT;
  wire bus_cap_7_;
  wire bus_cap_7__FF_INPUT;
  wire bus_cap_8_;
  wire bus_cap_8__FF_INPUT;
  wire bus_cap_9_;
  wire bus_cap_9__FF_INPUT;
  wire bus_sync_axi_bus_ECLK1;
  wire bus_sync_axi_bus_ECLK1_FF_INPUT;
  wire bus_sync_axi_bus_EECLK1;
  wire bus_sync_axi_bus_EECLK1_FF_INPUT;
  wire bus_sync_axi_bus_NCLK2;
  wire bus_sync_axi_bus__abc_3782_n457;
  wire bus_sync_axi_bus__abc_3782_n458;
  wire bus_sync_axi_bus__abc_3782_n460;
  wire bus_sync_axi_bus__abc_3782_n461;
  wire bus_sync_axi_bus__abc_3782_n462;
  wire bus_sync_axi_bus__abc_3782_n463;
  wire bus_sync_axi_bus__abc_3782_n465;
  wire bus_sync_axi_bus__abc_3782_n466;
  wire bus_sync_axi_bus__abc_3782_n468;
  wire bus_sync_axi_bus__abc_3782_n469;
  wire bus_sync_axi_bus__abc_3782_n471;
  wire bus_sync_axi_bus__abc_3782_n472;
  wire bus_sync_axi_bus__abc_3782_n474;
  wire bus_sync_axi_bus__abc_3782_n475;
  wire bus_sync_axi_bus__abc_3782_n477;
  wire bus_sync_axi_bus__abc_3782_n478;
  wire bus_sync_axi_bus__abc_3782_n480;
  wire bus_sync_axi_bus__abc_3782_n481;
  wire bus_sync_axi_bus__abc_3782_n483;
  wire bus_sync_axi_bus__abc_3782_n484;
  wire bus_sync_axi_bus__abc_3782_n486;
  wire bus_sync_axi_bus__abc_3782_n487;
  wire bus_sync_axi_bus__abc_3782_n489;
  wire bus_sync_axi_bus__abc_3782_n490;
  wire bus_sync_axi_bus__abc_3782_n492;
  wire bus_sync_axi_bus__abc_3782_n493;
  wire bus_sync_axi_bus__abc_3782_n495;
  wire bus_sync_axi_bus__abc_3782_n496;
  wire bus_sync_axi_bus__abc_3782_n498;
  wire bus_sync_axi_bus__abc_3782_n499;
  wire bus_sync_axi_bus__abc_3782_n501;
  wire bus_sync_axi_bus__abc_3782_n502;
  wire bus_sync_axi_bus__abc_3782_n504;
  wire bus_sync_axi_bus__abc_3782_n505;
  wire bus_sync_axi_bus__abc_3782_n507;
  wire bus_sync_axi_bus__abc_3782_n508;
  wire bus_sync_axi_bus__abc_3782_n510;
  wire bus_sync_axi_bus__abc_3782_n511;
  wire bus_sync_axi_bus__abc_3782_n513;
  wire bus_sync_axi_bus__abc_3782_n514;
  wire bus_sync_axi_bus__abc_3782_n516;
  wire bus_sync_axi_bus__abc_3782_n517;
  wire bus_sync_axi_bus__abc_3782_n519;
  wire bus_sync_axi_bus__abc_3782_n520;
  wire bus_sync_axi_bus__abc_3782_n522;
  wire bus_sync_axi_bus__abc_3782_n523;
  wire bus_sync_axi_bus__abc_3782_n525;
  wire bus_sync_axi_bus__abc_3782_n526;
  wire bus_sync_axi_bus__abc_3782_n528;
  wire bus_sync_axi_bus__abc_3782_n529;
  wire bus_sync_axi_bus__abc_3782_n531;
  wire bus_sync_axi_bus__abc_3782_n532;
  wire bus_sync_axi_bus__abc_3782_n534;
  wire bus_sync_axi_bus__abc_3782_n535;
  wire bus_sync_axi_bus__abc_3782_n537;
  wire bus_sync_axi_bus__abc_3782_n538;
  wire bus_sync_axi_bus__abc_3782_n540;
  wire bus_sync_axi_bus__abc_3782_n541;
  wire bus_sync_axi_bus__abc_3782_n543;
  wire bus_sync_axi_bus__abc_3782_n544;
  wire bus_sync_axi_bus__abc_3782_n546;
  wire bus_sync_axi_bus__abc_3782_n547;
  wire bus_sync_axi_bus__abc_3782_n549;
  wire bus_sync_axi_bus__abc_3782_n550;
  wire bus_sync_axi_bus__abc_3782_n552;
  wire bus_sync_axi_bus__abc_3782_n553;
  wire bus_sync_axi_bus__abc_3782_n555;
  wire bus_sync_axi_bus__abc_3782_n556;
  wire bus_sync_axi_bus__abc_3782_n558;
  wire bus_sync_axi_bus__abc_3782_n559;
  wire bus_sync_axi_bus__abc_3782_n561;
  wire bus_sync_axi_bus__abc_3782_n562;
  wire bus_sync_axi_bus__abc_3782_n564;
  wire bus_sync_axi_bus__abc_3782_n565;
  wire bus_sync_axi_bus__abc_3782_n567;
  wire bus_sync_axi_bus__abc_3782_n568;
  wire bus_sync_axi_bus__abc_3782_n570;
  wire bus_sync_axi_bus__abc_3782_n571;
  wire bus_sync_axi_bus__abc_3782_n573;
  wire bus_sync_axi_bus__abc_3782_n574;
  wire bus_sync_axi_bus__abc_3782_n576;
  wire bus_sync_axi_bus__abc_3782_n577;
  wire bus_sync_axi_bus__abc_3782_n579;
  wire bus_sync_axi_bus__abc_3782_n580;
  wire bus_sync_axi_bus__abc_3782_n582;
  wire bus_sync_axi_bus__abc_3782_n583;
  wire bus_sync_axi_bus__abc_3782_n585;
  wire bus_sync_axi_bus__abc_3782_n586;
  wire bus_sync_axi_bus__abc_3782_n588;
  wire bus_sync_axi_bus__abc_3782_n589;
  wire bus_sync_axi_bus__abc_3782_n591;
  wire bus_sync_axi_bus__abc_3782_n592;
  wire bus_sync_axi_bus__abc_3782_n594;
  wire bus_sync_axi_bus__abc_3782_n595;
  wire bus_sync_axi_bus__abc_3782_n597;
  wire bus_sync_axi_bus__abc_3782_n598;
  wire bus_sync_axi_bus__abc_3782_n600;
  wire bus_sync_axi_bus__abc_3782_n601;
  wire bus_sync_axi_bus__abc_3782_n603;
  wire bus_sync_axi_bus__abc_3782_n604;
  wire bus_sync_axi_bus__abc_3782_n606;
  wire bus_sync_axi_bus__abc_3782_n607;
  wire bus_sync_axi_bus__abc_3782_n609;
  wire bus_sync_axi_bus__abc_3782_n610;
  wire bus_sync_axi_bus__abc_3782_n612;
  wire bus_sync_axi_bus__abc_3782_n613;
  wire bus_sync_axi_bus__abc_3782_n615;
  wire bus_sync_axi_bus__abc_3782_n616;
  wire bus_sync_axi_bus__abc_3782_n618;
  wire bus_sync_axi_bus__abc_3782_n619;
  wire bus_sync_axi_bus__abc_3782_n621;
  wire bus_sync_axi_bus__abc_3782_n622;
  wire bus_sync_axi_bus__abc_3782_n624;
  wire bus_sync_axi_bus__abc_3782_n625;
  wire bus_sync_axi_bus__abc_3782_n627;
  wire bus_sync_axi_bus__abc_3782_n628;
  wire bus_sync_axi_bus__abc_3782_n630;
  wire bus_sync_axi_bus__abc_3782_n631;
  wire bus_sync_axi_bus__abc_3782_n633;
  wire bus_sync_axi_bus__abc_3782_n634;
  wire bus_sync_axi_bus__abc_3782_n636;
  wire bus_sync_axi_bus__abc_3782_n637;
  wire bus_sync_axi_bus__abc_3782_n639;
  wire bus_sync_axi_bus__abc_3782_n640;
  wire bus_sync_axi_bus__abc_3782_n642;
  wire bus_sync_axi_bus__abc_3782_n643;
  wire bus_sync_axi_bus__abc_3782_n645;
  wire bus_sync_axi_bus__abc_3782_n646;
  wire bus_sync_axi_bus__abc_3782_n648;
  wire bus_sync_axi_bus__abc_3782_n649;
  wire bus_sync_axi_bus_reg_data1_0_;
  wire bus_sync_axi_bus_reg_data1_0__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_10_;
  wire bus_sync_axi_bus_reg_data1_10__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_11_;
  wire bus_sync_axi_bus_reg_data1_11__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_12_;
  wire bus_sync_axi_bus_reg_data1_12__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_13_;
  wire bus_sync_axi_bus_reg_data1_13__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_14_;
  wire bus_sync_axi_bus_reg_data1_14__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_15_;
  wire bus_sync_axi_bus_reg_data1_15__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_16_;
  wire bus_sync_axi_bus_reg_data1_16__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_17_;
  wire bus_sync_axi_bus_reg_data1_17__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_18_;
  wire bus_sync_axi_bus_reg_data1_18__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_19_;
  wire bus_sync_axi_bus_reg_data1_19__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_1_;
  wire bus_sync_axi_bus_reg_data1_1__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_20_;
  wire bus_sync_axi_bus_reg_data1_20__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_21_;
  wire bus_sync_axi_bus_reg_data1_21__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_22_;
  wire bus_sync_axi_bus_reg_data1_22__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_23_;
  wire bus_sync_axi_bus_reg_data1_23__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_24_;
  wire bus_sync_axi_bus_reg_data1_24__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_25_;
  wire bus_sync_axi_bus_reg_data1_25__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_26_;
  wire bus_sync_axi_bus_reg_data1_26__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_27_;
  wire bus_sync_axi_bus_reg_data1_27__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_28_;
  wire bus_sync_axi_bus_reg_data1_28__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_29_;
  wire bus_sync_axi_bus_reg_data1_29__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_2_;
  wire bus_sync_axi_bus_reg_data1_2__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_30_;
  wire bus_sync_axi_bus_reg_data1_30__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_31_;
  wire bus_sync_axi_bus_reg_data1_31__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_32_;
  wire bus_sync_axi_bus_reg_data1_32__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_33_;
  wire bus_sync_axi_bus_reg_data1_33__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_34_;
  wire bus_sync_axi_bus_reg_data1_34__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_35_;
  wire bus_sync_axi_bus_reg_data1_35__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_36_;
  wire bus_sync_axi_bus_reg_data1_36__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_37_;
  wire bus_sync_axi_bus_reg_data1_37__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_38_;
  wire bus_sync_axi_bus_reg_data1_38__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_39_;
  wire bus_sync_axi_bus_reg_data1_39__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_3_;
  wire bus_sync_axi_bus_reg_data1_3__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_40_;
  wire bus_sync_axi_bus_reg_data1_40__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_41_;
  wire bus_sync_axi_bus_reg_data1_41__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_42_;
  wire bus_sync_axi_bus_reg_data1_42__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_43_;
  wire bus_sync_axi_bus_reg_data1_43__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_44_;
  wire bus_sync_axi_bus_reg_data1_44__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_45_;
  wire bus_sync_axi_bus_reg_data1_45__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_46_;
  wire bus_sync_axi_bus_reg_data1_46__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_47_;
  wire bus_sync_axi_bus_reg_data1_47__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_48_;
  wire bus_sync_axi_bus_reg_data1_48__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_49_;
  wire bus_sync_axi_bus_reg_data1_49__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_4_;
  wire bus_sync_axi_bus_reg_data1_4__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_50_;
  wire bus_sync_axi_bus_reg_data1_50__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_51_;
  wire bus_sync_axi_bus_reg_data1_51__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_52_;
  wire bus_sync_axi_bus_reg_data1_52__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_53_;
  wire bus_sync_axi_bus_reg_data1_53__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_54_;
  wire bus_sync_axi_bus_reg_data1_54__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_55_;
  wire bus_sync_axi_bus_reg_data1_55__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_56_;
  wire bus_sync_axi_bus_reg_data1_56__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_57_;
  wire bus_sync_axi_bus_reg_data1_57__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_58_;
  wire bus_sync_axi_bus_reg_data1_58__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_59_;
  wire bus_sync_axi_bus_reg_data1_59__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_5_;
  wire bus_sync_axi_bus_reg_data1_5__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_60_;
  wire bus_sync_axi_bus_reg_data1_60__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_61_;
  wire bus_sync_axi_bus_reg_data1_61__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_62_;
  wire bus_sync_axi_bus_reg_data1_62__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_63_;
  wire bus_sync_axi_bus_reg_data1_63__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_6_;
  wire bus_sync_axi_bus_reg_data1_6__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_7_;
  wire bus_sync_axi_bus_reg_data1_7__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_8_;
  wire bus_sync_axi_bus_reg_data1_8__FF_INPUT;
  wire bus_sync_axi_bus_reg_data1_9_;
  wire bus_sync_axi_bus_reg_data1_9__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_0_;
  wire bus_sync_axi_bus_reg_data2_0__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_10_;
  wire bus_sync_axi_bus_reg_data2_10__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_11_;
  wire bus_sync_axi_bus_reg_data2_11__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_12_;
  wire bus_sync_axi_bus_reg_data2_12__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_13_;
  wire bus_sync_axi_bus_reg_data2_13__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_14_;
  wire bus_sync_axi_bus_reg_data2_14__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_15_;
  wire bus_sync_axi_bus_reg_data2_15__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_16_;
  wire bus_sync_axi_bus_reg_data2_16__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_17_;
  wire bus_sync_axi_bus_reg_data2_17__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_18_;
  wire bus_sync_axi_bus_reg_data2_18__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_19_;
  wire bus_sync_axi_bus_reg_data2_19__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_1_;
  wire bus_sync_axi_bus_reg_data2_1__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_20_;
  wire bus_sync_axi_bus_reg_data2_20__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_21_;
  wire bus_sync_axi_bus_reg_data2_21__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_22_;
  wire bus_sync_axi_bus_reg_data2_22__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_23_;
  wire bus_sync_axi_bus_reg_data2_23__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_24_;
  wire bus_sync_axi_bus_reg_data2_24__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_25_;
  wire bus_sync_axi_bus_reg_data2_25__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_26_;
  wire bus_sync_axi_bus_reg_data2_26__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_27_;
  wire bus_sync_axi_bus_reg_data2_27__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_28_;
  wire bus_sync_axi_bus_reg_data2_28__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_29_;
  wire bus_sync_axi_bus_reg_data2_29__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_2_;
  wire bus_sync_axi_bus_reg_data2_2__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_30_;
  wire bus_sync_axi_bus_reg_data2_30__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_31_;
  wire bus_sync_axi_bus_reg_data2_31__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_32_;
  wire bus_sync_axi_bus_reg_data2_32__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_33_;
  wire bus_sync_axi_bus_reg_data2_33__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_34_;
  wire bus_sync_axi_bus_reg_data2_34__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_35_;
  wire bus_sync_axi_bus_reg_data2_35__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_36_;
  wire bus_sync_axi_bus_reg_data2_36__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_37_;
  wire bus_sync_axi_bus_reg_data2_37__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_38_;
  wire bus_sync_axi_bus_reg_data2_38__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_39_;
  wire bus_sync_axi_bus_reg_data2_39__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_3_;
  wire bus_sync_axi_bus_reg_data2_3__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_40_;
  wire bus_sync_axi_bus_reg_data2_40__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_41_;
  wire bus_sync_axi_bus_reg_data2_41__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_42_;
  wire bus_sync_axi_bus_reg_data2_42__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_43_;
  wire bus_sync_axi_bus_reg_data2_43__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_44_;
  wire bus_sync_axi_bus_reg_data2_44__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_45_;
  wire bus_sync_axi_bus_reg_data2_45__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_46_;
  wire bus_sync_axi_bus_reg_data2_46__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_47_;
  wire bus_sync_axi_bus_reg_data2_47__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_48_;
  wire bus_sync_axi_bus_reg_data2_48__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_49_;
  wire bus_sync_axi_bus_reg_data2_49__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_4_;
  wire bus_sync_axi_bus_reg_data2_4__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_50_;
  wire bus_sync_axi_bus_reg_data2_50__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_51_;
  wire bus_sync_axi_bus_reg_data2_51__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_52_;
  wire bus_sync_axi_bus_reg_data2_52__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_53_;
  wire bus_sync_axi_bus_reg_data2_53__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_54_;
  wire bus_sync_axi_bus_reg_data2_54__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_55_;
  wire bus_sync_axi_bus_reg_data2_55__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_56_;
  wire bus_sync_axi_bus_reg_data2_56__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_57_;
  wire bus_sync_axi_bus_reg_data2_57__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_58_;
  wire bus_sync_axi_bus_reg_data2_58__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_59_;
  wire bus_sync_axi_bus_reg_data2_59__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_5_;
  wire bus_sync_axi_bus_reg_data2_5__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_60_;
  wire bus_sync_axi_bus_reg_data2_60__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_61_;
  wire bus_sync_axi_bus_reg_data2_61__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_62_;
  wire bus_sync_axi_bus_reg_data2_62__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_63_;
  wire bus_sync_axi_bus_reg_data2_63__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_6_;
  wire bus_sync_axi_bus_reg_data2_6__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_7_;
  wire bus_sync_axi_bus_reg_data2_7__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_8_;
  wire bus_sync_axi_bus_reg_data2_8__FF_INPUT;
  wire bus_sync_axi_bus_reg_data2_9_;
  wire bus_sync_axi_bus_reg_data2_9__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_0__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_10__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_11__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_12__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_13__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_14__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_15__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_16__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_17__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_18__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_19__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_1__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_20__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_21__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_22__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_23__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_24__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_25__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_26__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_27__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_28__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_29__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_2__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_30__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_31__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_32__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_33__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_34__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_35__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_36__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_37__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_38__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_39__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_3__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_40__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_41__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_42__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_43__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_44__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_45__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_46__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_47__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_48__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_49__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_4__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_50__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_51__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_52__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_53__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_54__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_55__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_56__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_57__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_58__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_59__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_5__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_60__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_61__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_62__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_63__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_6__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_7__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_8__FF_INPUT;
  wire bus_sync_axi_bus_reg_data3_9__FF_INPUT;
  wire bus_sync_rdata_ECLK2;
  wire bus_sync_rdata_ECLK2_FF_INPUT;
  wire bus_sync_rdata_EECLK2;
  wire bus_sync_rdata_EECLK2_FF_INPUT;
  wire bus_sync_rdata_NCLK1;
  wire bus_sync_rdata__abc_3590_n201_1;
  wire bus_sync_rdata__abc_3590_n202_1;
  wire bus_sync_rdata__abc_3590_n204_1;
  wire bus_sync_rdata__abc_3590_n205_1;
  wire bus_sync_rdata__abc_3590_n206_1;
  wire bus_sync_rdata__abc_3590_n207_1;
  wire bus_sync_rdata__abc_3590_n209_1;
  wire bus_sync_rdata__abc_3590_n210_1;
  wire bus_sync_rdata__abc_3590_n212_1;
  wire bus_sync_rdata__abc_3590_n213_1;
  wire bus_sync_rdata__abc_3590_n215_1;
  wire bus_sync_rdata__abc_3590_n216_1;
  wire bus_sync_rdata__abc_3590_n218_1;
  wire bus_sync_rdata__abc_3590_n219_1;
  wire bus_sync_rdata__abc_3590_n221_1;
  wire bus_sync_rdata__abc_3590_n222_1;
  wire bus_sync_rdata__abc_3590_n224_1;
  wire bus_sync_rdata__abc_3590_n225_1;
  wire bus_sync_rdata__abc_3590_n227_1;
  wire bus_sync_rdata__abc_3590_n228_1;
  wire bus_sync_rdata__abc_3590_n230_1;
  wire bus_sync_rdata__abc_3590_n231_1;
  wire bus_sync_rdata__abc_3590_n233;
  wire bus_sync_rdata__abc_3590_n234;
  wire bus_sync_rdata__abc_3590_n236;
  wire bus_sync_rdata__abc_3590_n237;
  wire bus_sync_rdata__abc_3590_n239;
  wire bus_sync_rdata__abc_3590_n240;
  wire bus_sync_rdata__abc_3590_n242;
  wire bus_sync_rdata__abc_3590_n243;
  wire bus_sync_rdata__abc_3590_n245;
  wire bus_sync_rdata__abc_3590_n246;
  wire bus_sync_rdata__abc_3590_n248;
  wire bus_sync_rdata__abc_3590_n249;
  wire bus_sync_rdata__abc_3590_n251;
  wire bus_sync_rdata__abc_3590_n252;
  wire bus_sync_rdata__abc_3590_n254;
  wire bus_sync_rdata__abc_3590_n255;
  wire bus_sync_rdata__abc_3590_n257;
  wire bus_sync_rdata__abc_3590_n258;
  wire bus_sync_rdata__abc_3590_n260;
  wire bus_sync_rdata__abc_3590_n261;
  wire bus_sync_rdata__abc_3590_n263;
  wire bus_sync_rdata__abc_3590_n264;
  wire bus_sync_rdata__abc_3590_n266;
  wire bus_sync_rdata__abc_3590_n267;
  wire bus_sync_rdata__abc_3590_n269;
  wire bus_sync_rdata__abc_3590_n270;
  wire bus_sync_rdata__abc_3590_n272;
  wire bus_sync_rdata__abc_3590_n273;
  wire bus_sync_rdata__abc_3590_n275;
  wire bus_sync_rdata__abc_3590_n276;
  wire bus_sync_rdata__abc_3590_n278;
  wire bus_sync_rdata__abc_3590_n279;
  wire bus_sync_rdata__abc_3590_n281;
  wire bus_sync_rdata__abc_3590_n282;
  wire bus_sync_rdata__abc_3590_n284;
  wire bus_sync_rdata__abc_3590_n285;
  wire bus_sync_rdata__abc_3590_n287;
  wire bus_sync_rdata__abc_3590_n288;
  wire bus_sync_rdata__abc_3590_n290;
  wire bus_sync_rdata__abc_3590_n291;
  wire bus_sync_rdata__abc_3590_n293;
  wire bus_sync_rdata__abc_3590_n294;
  wire bus_sync_rdata__abc_3590_n296;
  wire bus_sync_rdata__abc_3590_n297;
  wire bus_sync_rdata_data_in_0_;
  wire bus_sync_rdata_data_in_10_;
  wire bus_sync_rdata_data_in_11_;
  wire bus_sync_rdata_data_in_12_;
  wire bus_sync_rdata_data_in_13_;
  wire bus_sync_rdata_data_in_14_;
  wire bus_sync_rdata_data_in_15_;
  wire bus_sync_rdata_data_in_16_;
  wire bus_sync_rdata_data_in_17_;
  wire bus_sync_rdata_data_in_18_;
  wire bus_sync_rdata_data_in_19_;
  wire bus_sync_rdata_data_in_1_;
  wire bus_sync_rdata_data_in_20_;
  wire bus_sync_rdata_data_in_21_;
  wire bus_sync_rdata_data_in_22_;
  wire bus_sync_rdata_data_in_23_;
  wire bus_sync_rdata_data_in_24_;
  wire bus_sync_rdata_data_in_25_;
  wire bus_sync_rdata_data_in_26_;
  wire bus_sync_rdata_data_in_27_;
  wire bus_sync_rdata_data_in_28_;
  wire bus_sync_rdata_data_in_29_;
  wire bus_sync_rdata_data_in_2_;
  wire bus_sync_rdata_data_in_30_;
  wire bus_sync_rdata_data_in_31_;
  wire bus_sync_rdata_data_in_3_;
  wire bus_sync_rdata_data_in_4_;
  wire bus_sync_rdata_data_in_5_;
  wire bus_sync_rdata_data_in_6_;
  wire bus_sync_rdata_data_in_7_;
  wire bus_sync_rdata_data_in_8_;
  wire bus_sync_rdata_data_in_9_;
  wire bus_sync_rdata_data_out_0_;
  wire bus_sync_rdata_data_out_10_;
  wire bus_sync_rdata_data_out_11_;
  wire bus_sync_rdata_data_out_12_;
  wire bus_sync_rdata_data_out_13_;
  wire bus_sync_rdata_data_out_14_;
  wire bus_sync_rdata_data_out_15_;
  wire bus_sync_rdata_data_out_16_;
  wire bus_sync_rdata_data_out_17_;
  wire bus_sync_rdata_data_out_18_;
  wire bus_sync_rdata_data_out_19_;
  wire bus_sync_rdata_data_out_1_;
  wire bus_sync_rdata_data_out_20_;
  wire bus_sync_rdata_data_out_21_;
  wire bus_sync_rdata_data_out_22_;
  wire bus_sync_rdata_data_out_23_;
  wire bus_sync_rdata_data_out_24_;
  wire bus_sync_rdata_data_out_25_;
  wire bus_sync_rdata_data_out_26_;
  wire bus_sync_rdata_data_out_27_;
  wire bus_sync_rdata_data_out_28_;
  wire bus_sync_rdata_data_out_29_;
  wire bus_sync_rdata_data_out_2_;
  wire bus_sync_rdata_data_out_30_;
  wire bus_sync_rdata_data_out_31_;
  wire bus_sync_rdata_data_out_3_;
  wire bus_sync_rdata_data_out_4_;
  wire bus_sync_rdata_data_out_5_;
  wire bus_sync_rdata_data_out_6_;
  wire bus_sync_rdata_data_out_7_;
  wire bus_sync_rdata_data_out_8_;
  wire bus_sync_rdata_data_out_9_;
  wire bus_sync_rdata_reg_data1_0_;
  wire bus_sync_rdata_reg_data1_0__FF_INPUT;
  wire bus_sync_rdata_reg_data1_10_;
  wire bus_sync_rdata_reg_data1_10__FF_INPUT;
  wire bus_sync_rdata_reg_data1_11_;
  wire bus_sync_rdata_reg_data1_11__FF_INPUT;
  wire bus_sync_rdata_reg_data1_12_;
  wire bus_sync_rdata_reg_data1_12__FF_INPUT;
  wire bus_sync_rdata_reg_data1_13_;
  wire bus_sync_rdata_reg_data1_13__FF_INPUT;
  wire bus_sync_rdata_reg_data1_14_;
  wire bus_sync_rdata_reg_data1_14__FF_INPUT;
  wire bus_sync_rdata_reg_data1_15_;
  wire bus_sync_rdata_reg_data1_15__FF_INPUT;
  wire bus_sync_rdata_reg_data1_16_;
  wire bus_sync_rdata_reg_data1_16__FF_INPUT;
  wire bus_sync_rdata_reg_data1_17_;
  wire bus_sync_rdata_reg_data1_17__FF_INPUT;
  wire bus_sync_rdata_reg_data1_18_;
  wire bus_sync_rdata_reg_data1_18__FF_INPUT;
  wire bus_sync_rdata_reg_data1_19_;
  wire bus_sync_rdata_reg_data1_19__FF_INPUT;
  wire bus_sync_rdata_reg_data1_1_;
  wire bus_sync_rdata_reg_data1_1__FF_INPUT;
  wire bus_sync_rdata_reg_data1_20_;
  wire bus_sync_rdata_reg_data1_20__FF_INPUT;
  wire bus_sync_rdata_reg_data1_21_;
  wire bus_sync_rdata_reg_data1_21__FF_INPUT;
  wire bus_sync_rdata_reg_data1_22_;
  wire bus_sync_rdata_reg_data1_22__FF_INPUT;
  wire bus_sync_rdata_reg_data1_23_;
  wire bus_sync_rdata_reg_data1_23__FF_INPUT;
  wire bus_sync_rdata_reg_data1_24_;
  wire bus_sync_rdata_reg_data1_24__FF_INPUT;
  wire bus_sync_rdata_reg_data1_25_;
  wire bus_sync_rdata_reg_data1_25__FF_INPUT;
  wire bus_sync_rdata_reg_data1_26_;
  wire bus_sync_rdata_reg_data1_26__FF_INPUT;
  wire bus_sync_rdata_reg_data1_27_;
  wire bus_sync_rdata_reg_data1_27__FF_INPUT;
  wire bus_sync_rdata_reg_data1_28_;
  wire bus_sync_rdata_reg_data1_28__FF_INPUT;
  wire bus_sync_rdata_reg_data1_29_;
  wire bus_sync_rdata_reg_data1_29__FF_INPUT;
  wire bus_sync_rdata_reg_data1_2_;
  wire bus_sync_rdata_reg_data1_2__FF_INPUT;
  wire bus_sync_rdata_reg_data1_30_;
  wire bus_sync_rdata_reg_data1_30__FF_INPUT;
  wire bus_sync_rdata_reg_data1_31_;
  wire bus_sync_rdata_reg_data1_31__FF_INPUT;
  wire bus_sync_rdata_reg_data1_3_;
  wire bus_sync_rdata_reg_data1_3__FF_INPUT;
  wire bus_sync_rdata_reg_data1_4_;
  wire bus_sync_rdata_reg_data1_4__FF_INPUT;
  wire bus_sync_rdata_reg_data1_5_;
  wire bus_sync_rdata_reg_data1_5__FF_INPUT;
  wire bus_sync_rdata_reg_data1_6_;
  wire bus_sync_rdata_reg_data1_6__FF_INPUT;
  wire bus_sync_rdata_reg_data1_7_;
  wire bus_sync_rdata_reg_data1_7__FF_INPUT;
  wire bus_sync_rdata_reg_data1_8_;
  wire bus_sync_rdata_reg_data1_8__FF_INPUT;
  wire bus_sync_rdata_reg_data1_9_;
  wire bus_sync_rdata_reg_data1_9__FF_INPUT;
  wire bus_sync_rdata_reg_data2_0_;
  wire bus_sync_rdata_reg_data2_0__FF_INPUT;
  wire bus_sync_rdata_reg_data2_10_;
  wire bus_sync_rdata_reg_data2_10__FF_INPUT;
  wire bus_sync_rdata_reg_data2_11_;
  wire bus_sync_rdata_reg_data2_11__FF_INPUT;
  wire bus_sync_rdata_reg_data2_12_;
  wire bus_sync_rdata_reg_data2_12__FF_INPUT;
  wire bus_sync_rdata_reg_data2_13_;
  wire bus_sync_rdata_reg_data2_13__FF_INPUT;
  wire bus_sync_rdata_reg_data2_14_;
  wire bus_sync_rdata_reg_data2_14__FF_INPUT;
  wire bus_sync_rdata_reg_data2_15_;
  wire bus_sync_rdata_reg_data2_15__FF_INPUT;
  wire bus_sync_rdata_reg_data2_16_;
  wire bus_sync_rdata_reg_data2_16__FF_INPUT;
  wire bus_sync_rdata_reg_data2_17_;
  wire bus_sync_rdata_reg_data2_17__FF_INPUT;
  wire bus_sync_rdata_reg_data2_18_;
  wire bus_sync_rdata_reg_data2_18__FF_INPUT;
  wire bus_sync_rdata_reg_data2_19_;
  wire bus_sync_rdata_reg_data2_19__FF_INPUT;
  wire bus_sync_rdata_reg_data2_1_;
  wire bus_sync_rdata_reg_data2_1__FF_INPUT;
  wire bus_sync_rdata_reg_data2_20_;
  wire bus_sync_rdata_reg_data2_20__FF_INPUT;
  wire bus_sync_rdata_reg_data2_21_;
  wire bus_sync_rdata_reg_data2_21__FF_INPUT;
  wire bus_sync_rdata_reg_data2_22_;
  wire bus_sync_rdata_reg_data2_22__FF_INPUT;
  wire bus_sync_rdata_reg_data2_23_;
  wire bus_sync_rdata_reg_data2_23__FF_INPUT;
  wire bus_sync_rdata_reg_data2_24_;
  wire bus_sync_rdata_reg_data2_24__FF_INPUT;
  wire bus_sync_rdata_reg_data2_25_;
  wire bus_sync_rdata_reg_data2_25__FF_INPUT;
  wire bus_sync_rdata_reg_data2_26_;
  wire bus_sync_rdata_reg_data2_26__FF_INPUT;
  wire bus_sync_rdata_reg_data2_27_;
  wire bus_sync_rdata_reg_data2_27__FF_INPUT;
  wire bus_sync_rdata_reg_data2_28_;
  wire bus_sync_rdata_reg_data2_28__FF_INPUT;
  wire bus_sync_rdata_reg_data2_29_;
  wire bus_sync_rdata_reg_data2_29__FF_INPUT;
  wire bus_sync_rdata_reg_data2_2_;
  wire bus_sync_rdata_reg_data2_2__FF_INPUT;
  wire bus_sync_rdata_reg_data2_30_;
  wire bus_sync_rdata_reg_data2_30__FF_INPUT;
  wire bus_sync_rdata_reg_data2_31_;
  wire bus_sync_rdata_reg_data2_31__FF_INPUT;
  wire bus_sync_rdata_reg_data2_3_;
  wire bus_sync_rdata_reg_data2_3__FF_INPUT;
  wire bus_sync_rdata_reg_data2_4_;
  wire bus_sync_rdata_reg_data2_4__FF_INPUT;
  wire bus_sync_rdata_reg_data2_5_;
  wire bus_sync_rdata_reg_data2_5__FF_INPUT;
  wire bus_sync_rdata_reg_data2_6_;
  wire bus_sync_rdata_reg_data2_6__FF_INPUT;
  wire bus_sync_rdata_reg_data2_7_;
  wire bus_sync_rdata_reg_data2_7__FF_INPUT;
  wire bus_sync_rdata_reg_data2_8_;
  wire bus_sync_rdata_reg_data2_8__FF_INPUT;
  wire bus_sync_rdata_reg_data2_9_;
  wire bus_sync_rdata_reg_data2_9__FF_INPUT;
  wire bus_sync_rdata_reg_data3_0__FF_INPUT;
  wire bus_sync_rdata_reg_data3_10__FF_INPUT;
  wire bus_sync_rdata_reg_data3_11__FF_INPUT;
  wire bus_sync_rdata_reg_data3_12__FF_INPUT;
  wire bus_sync_rdata_reg_data3_13__FF_INPUT;
  wire bus_sync_rdata_reg_data3_14__FF_INPUT;
  wire bus_sync_rdata_reg_data3_15__FF_INPUT;
  wire bus_sync_rdata_reg_data3_16__FF_INPUT;
  wire bus_sync_rdata_reg_data3_17__FF_INPUT;
  wire bus_sync_rdata_reg_data3_18__FF_INPUT;
  wire bus_sync_rdata_reg_data3_19__FF_INPUT;
  wire bus_sync_rdata_reg_data3_1__FF_INPUT;
  wire bus_sync_rdata_reg_data3_20__FF_INPUT;
  wire bus_sync_rdata_reg_data3_21__FF_INPUT;
  wire bus_sync_rdata_reg_data3_22__FF_INPUT;
  wire bus_sync_rdata_reg_data3_23__FF_INPUT;
  wire bus_sync_rdata_reg_data3_24__FF_INPUT;
  wire bus_sync_rdata_reg_data3_25__FF_INPUT;
  wire bus_sync_rdata_reg_data3_26__FF_INPUT;
  wire bus_sync_rdata_reg_data3_27__FF_INPUT;
  wire bus_sync_rdata_reg_data3_28__FF_INPUT;
  wire bus_sync_rdata_reg_data3_29__FF_INPUT;
  wire bus_sync_rdata_reg_data3_2__FF_INPUT;
  wire bus_sync_rdata_reg_data3_30__FF_INPUT;
  wire bus_sync_rdata_reg_data3_31__FF_INPUT;
  wire bus_sync_rdata_reg_data3_3__FF_INPUT;
  wire bus_sync_rdata_reg_data3_4__FF_INPUT;
  wire bus_sync_rdata_reg_data3_5__FF_INPUT;
  wire bus_sync_rdata_reg_data3_6__FF_INPUT;
  wire bus_sync_rdata_reg_data3_7__FF_INPUT;
  wire bus_sync_rdata_reg_data3_8__FF_INPUT;
  wire bus_sync_rdata_reg_data3_9__FF_INPUT;
  wire bus_sync_state_machine_ECLK1;
  wire bus_sync_state_machine_ECLK1_FF_INPUT;
  wire bus_sync_state_machine_EECLK1;
  wire bus_sync_state_machine_EECLK1_FF_INPUT;
  wire bus_sync_state_machine_NCLK2;
  wire bus_sync_state_machine__abc_3756_n37;
  wire bus_sync_state_machine__abc_3756_n38;
  wire bus_sync_state_machine__abc_3756_n40;
  wire bus_sync_state_machine__abc_3756_n41;
  wire bus_sync_state_machine__abc_3756_n42;
  wire bus_sync_state_machine__abc_3756_n43;
  wire bus_sync_state_machine__abc_3756_n45;
  wire bus_sync_state_machine__abc_3756_n46;
  wire bus_sync_state_machine__abc_3756_n48;
  wire bus_sync_state_machine__abc_3756_n49;
  wire bus_sync_state_machine_reg_data1_0_;
  wire bus_sync_state_machine_reg_data1_0__FF_INPUT;
  wire bus_sync_state_machine_reg_data1_1_;
  wire bus_sync_state_machine_reg_data1_1__FF_INPUT;
  wire bus_sync_state_machine_reg_data1_2_;
  wire bus_sync_state_machine_reg_data1_2__FF_INPUT;
  wire bus_sync_state_machine_reg_data1_3_;
  wire bus_sync_state_machine_reg_data1_3__FF_INPUT;
  wire bus_sync_state_machine_reg_data2_0_;
  wire bus_sync_state_machine_reg_data2_0__FF_INPUT;
  wire bus_sync_state_machine_reg_data2_1_;
  wire bus_sync_state_machine_reg_data2_1__FF_INPUT;
  wire bus_sync_state_machine_reg_data2_2_;
  wire bus_sync_state_machine_reg_data2_2__FF_INPUT;
  wire bus_sync_state_machine_reg_data2_3_;
  wire bus_sync_state_machine_reg_data2_3__FF_INPUT;
  wire bus_sync_state_machine_reg_data3_0__FF_INPUT;
  wire bus_sync_state_machine_reg_data3_1__FF_INPUT;
  wire bus_sync_state_machine_reg_data3_2__FF_INPUT;
  wire bus_sync_state_machine_reg_data3_3__FF_INPUT;
  wire bus_sync_status_ECLK2;
  wire bus_sync_status_ECLK2_FF_INPUT;
  wire bus_sync_status_EECLK2;
  wire bus_sync_status_EECLK2_FF_INPUT;
  wire bus_sync_status_NCLK1;
  wire bus_sync_status__abc_3569_n30;
  wire bus_sync_status__abc_3569_n31;
  wire bus_sync_status__abc_3569_n33;
  wire bus_sync_status__abc_3569_n34;
  wire bus_sync_status__abc_3569_n35;
  wire bus_sync_status__abc_3569_n36;
  wire bus_sync_status__abc_3569_n38;
  wire bus_sync_status__abc_3569_n39;
  wire bus_sync_status_data_out_0_;
  wire bus_sync_status_data_out_1_;
  wire bus_sync_status_data_out_2_;
  wire bus_sync_status_reg_data1_0_;
  wire bus_sync_status_reg_data1_0__FF_INPUT;
  wire bus_sync_status_reg_data1_1_;
  wire bus_sync_status_reg_data1_1__FF_INPUT;
  wire bus_sync_status_reg_data1_2_;
  wire bus_sync_status_reg_data1_2__FF_INPUT;
  wire bus_sync_status_reg_data2_0_;
  wire bus_sync_status_reg_data2_0__FF_INPUT;
  wire bus_sync_status_reg_data2_1_;
  wire bus_sync_status_reg_data2_1__FF_INPUT;
  wire bus_sync_status_reg_data2_2_;
  wire bus_sync_status_reg_data2_2__FF_INPUT;
  wire bus_sync_status_reg_data3_0__FF_INPUT;
  wire bus_sync_status_reg_data3_1__FF_INPUT;
  wire bus_sync_status_reg_data3_2__FF_INPUT;
  wire busy;
  wire counter_0_;
  wire counter_0__FF_INPUT;
  wire counter_10_;
  wire counter_10__FF_INPUT;
  wire counter_11_;
  wire counter_11__FF_INPUT;
  wire counter_12_;
  wire counter_12__FF_INPUT;
  wire counter_13_;
  wire counter_13__FF_INPUT;
  wire counter_14_;
  wire counter_14__FF_INPUT;
  wire counter_15_;
  wire counter_15__FF_INPUT;
  wire counter_16_;
  wire counter_16__FF_INPUT;
  wire counter_17_;
  wire counter_17__FF_INPUT;
  wire counter_18_;
  wire counter_18__FF_INPUT;
  wire counter_19_;
  wire counter_19__FF_INPUT;
  wire counter_1_;
  wire counter_1__FF_INPUT;
  wire counter_20_;
  wire counter_20__FF_INPUT;
  wire counter_21_;
  wire counter_21__FF_INPUT;
  wire counter_22_;
  wire counter_22__FF_INPUT;
  wire counter_23_;
  wire counter_23__FF_INPUT;
  wire counter_24_;
  wire counter_24__FF_INPUT;
  wire counter_25_;
  wire counter_25__FF_INPUT;
  wire counter_26_;
  wire counter_26__FF_INPUT;
  wire counter_27_;
  wire counter_27__FF_INPUT;
  wire counter_28_;
  wire counter_28__FF_INPUT;
  wire counter_29_;
  wire counter_29__FF_INPUT;
  wire counter_2_;
  wire counter_2__FF_INPUT;
  wire counter_30_;
  wire counter_30__FF_INPUT;
  wire counter_31_;
  wire counter_31__FF_INPUT;
  wire counter_32_;
  wire counter_32__FF_INPUT;
  wire counter_33_;
  wire counter_33__FF_INPUT;
  wire counter_34_;
  wire counter_34__FF_INPUT;
  wire counter_35_;
  wire counter_35__FF_INPUT;
  wire counter_36_;
  wire counter_36__FF_INPUT;
  wire counter_37_;
  wire counter_37__FF_INPUT;
  wire counter_38_;
  wire counter_38__FF_INPUT;
  wire counter_39_;
  wire counter_39__FF_INPUT;
  wire counter_3_;
  wire counter_3__FF_INPUT;
  wire counter_40_;
  wire counter_40__FF_INPUT;
  wire counter_41_;
  wire counter_41__FF_INPUT;
  wire counter_42_;
  wire counter_42__FF_INPUT;
  wire counter_43_;
  wire counter_43__FF_INPUT;
  wire counter_44_;
  wire counter_44__FF_INPUT;
  wire counter_45_;
  wire counter_45__FF_INPUT;
  wire counter_46_;
  wire counter_46__FF_INPUT;
  wire counter_47_;
  wire counter_47__FF_INPUT;
  wire counter_48_;
  wire counter_48__FF_INPUT;
  wire counter_49_;
  wire counter_49__FF_INPUT;
  wire counter_4_;
  wire counter_4__FF_INPUT;
  wire counter_50_;
  wire counter_50__FF_INPUT;
  wire counter_51_;
  wire counter_51__FF_INPUT;
  wire counter_52_;
  wire counter_52__FF_INPUT;
  wire counter_53_;
  wire counter_53__FF_INPUT;
  wire counter_54_;
  wire counter_54__FF_INPUT;
  wire counter_55_;
  wire counter_55__FF_INPUT;
  wire counter_56_;
  wire counter_56__FF_INPUT;
  wire counter_57_;
  wire counter_57__FF_INPUT;
  wire counter_58_;
  wire counter_58__FF_INPUT;
  wire counter_59_;
  wire counter_59__FF_INPUT;
  wire counter_5_;
  wire counter_5__FF_INPUT;
  wire counter_60_;
  wire counter_60__FF_INPUT;
  wire counter_61_;
  wire counter_61__FF_INPUT;
  wire counter_62_;
  wire counter_62__FF_INPUT;
  wire counter_63_;
  wire counter_63__FF_INPUT;
  wire counter_64_;
  wire counter_64__FF_INPUT;
  wire counter_65_;
  wire counter_65__FF_INPUT;
  wire counter_6_;
  wire counter_6__FF_INPUT;
  wire counter_7_;
  wire counter_7__FF_INPUT;
  wire counter_8_;
  wire counter_8__FF_INPUT;
  wire counter_9_;
  wire counter_9__FF_INPUT;
  wire fini_spi;
  wire fini_spi_FF_INPUT;
  wire fini_spi_clk;
  wire rdata_0__FF_INPUT;
  wire rdata_10__FF_INPUT;
  wire rdata_11__FF_INPUT;
  wire rdata_12__FF_INPUT;
  wire rdata_13__FF_INPUT;
  wire rdata_14__FF_INPUT;
  wire rdata_15__FF_INPUT;
  wire rdata_16__FF_INPUT;
  wire rdata_17__FF_INPUT;
  wire rdata_18__FF_INPUT;
  wire rdata_19__FF_INPUT;
  wire rdata_1__FF_INPUT;
  wire rdata_20__FF_INPUT;
  wire rdata_21__FF_INPUT;
  wire rdata_22__FF_INPUT;
  wire rdata_23__FF_INPUT;
  wire rdata_24__FF_INPUT;
  wire rdata_25__FF_INPUT;
  wire rdata_26__FF_INPUT;
  wire rdata_27__FF_INPUT;
  wire rdata_28__FF_INPUT;
  wire rdata_29__FF_INPUT;
  wire rdata_2__FF_INPUT;
  wire rdata_30__FF_INPUT;
  wire rdata_31__FF_INPUT;
  wire rdata_3__FF_INPUT;
  wire rdata_4__FF_INPUT;
  wire rdata_5__FF_INPUT;
  wire rdata_6__FF_INPUT;
  wire rdata_7__FF_INPUT;
  wire rdata_8__FF_INPUT;
  wire rdata_9__FF_INPUT;
  wire re;
  wire re_FF_INPUT;
  wire re_clk;
  wire sft_reg_0_;
  wire sft_reg_0__FF_INPUT;
  wire sft_reg_10_;
  wire sft_reg_10__FF_INPUT;
  wire sft_reg_11_;
  wire sft_reg_11__FF_INPUT;
  wire sft_reg_12_;
  wire sft_reg_12__FF_INPUT;
  wire sft_reg_13_;
  wire sft_reg_13__FF_INPUT;
  wire sft_reg_14_;
  wire sft_reg_14__FF_INPUT;
  wire sft_reg_15_;
  wire sft_reg_15__FF_INPUT;
  wire sft_reg_16_;
  wire sft_reg_16__FF_INPUT;
  wire sft_reg_17_;
  wire sft_reg_17__FF_INPUT;
  wire sft_reg_18_;
  wire sft_reg_18__FF_INPUT;
  wire sft_reg_19_;
  wire sft_reg_19__FF_INPUT;
  wire sft_reg_1_;
  wire sft_reg_1__FF_INPUT;
  wire sft_reg_20_;
  wire sft_reg_20__FF_INPUT;
  wire sft_reg_21_;
  wire sft_reg_21__FF_INPUT;
  wire sft_reg_22_;
  wire sft_reg_22__FF_INPUT;
  wire sft_reg_23_;
  wire sft_reg_23__FF_INPUT;
  wire sft_reg_24_;
  wire sft_reg_24__FF_INPUT;
  wire sft_reg_25_;
  wire sft_reg_25__FF_INPUT;
  wire sft_reg_26_;
  wire sft_reg_26__FF_INPUT;
  wire sft_reg_27_;
  wire sft_reg_27__FF_INPUT;
  wire sft_reg_28_;
  wire sft_reg_28__FF_INPUT;
  wire sft_reg_29_;
  wire sft_reg_29__FF_INPUT;
  wire sft_reg_2_;
  wire sft_reg_2__FF_INPUT;
  wire sft_reg_30_;
  wire sft_reg_30__FF_INPUT;
  wire sft_reg_3_;
  wire sft_reg_3__FF_INPUT;
  wire sft_reg_4_;
  wire sft_reg_4__FF_INPUT;
  wire sft_reg_5_;
  wire sft_reg_5__FF_INPUT;
  wire sft_reg_6_;
  wire sft_reg_6__FF_INPUT;
  wire sft_reg_7_;
  wire sft_reg_7__FF_INPUT;
  wire sft_reg_8_;
  wire sft_reg_8__FF_INPUT;
  wire sft_reg_9_;
  wire sft_reg_9__FF_INPUT;
  wire state_0_;
  wire state_1_;
  wire state_3_;
  wire state_4_;
  wire state_5_;
  wire state_6_;
  wire state_7_;
  wire we;
  wire we_FF_INPUT;
  wire we_clk;
  AND2X2 AND2X2_1 ( .A(_abc_4108_n598_1), .B(_abc_4108_n600), .Y(_abc_4108_n601) );
  AND2X2 AND2X2_10 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_7_), .Y(bus_sync_axi_bus_reg_data3_7__FF_INPUT) );
  AND2X2 AND2X2_100 ( .A(RST), .B(A_ADDR_1_), .Y(bus_sync_axi_bus_reg_data1_33__FF_INPUT) );
  AND2X2 AND2X2_101 ( .A(RST), .B(A_ADDR_2_), .Y(bus_sync_axi_bus_reg_data1_34__FF_INPUT) );
  AND2X2 AND2X2_102 ( .A(RST), .B(A_ADDR_3_), .Y(bus_sync_axi_bus_reg_data1_35__FF_INPUT) );
  AND2X2 AND2X2_103 ( .A(RST), .B(A_ADDR_4_), .Y(bus_sync_axi_bus_reg_data1_36__FF_INPUT) );
  AND2X2 AND2X2_104 ( .A(RST), .B(A_ADDR_5_), .Y(bus_sync_axi_bus_reg_data1_37__FF_INPUT) );
  AND2X2 AND2X2_105 ( .A(RST), .B(A_ADDR_6_), .Y(bus_sync_axi_bus_reg_data1_38__FF_INPUT) );
  AND2X2 AND2X2_106 ( .A(RST), .B(A_ADDR_7_), .Y(bus_sync_axi_bus_reg_data1_39__FF_INPUT) );
  AND2X2 AND2X2_107 ( .A(RST), .B(A_ADDR_8_), .Y(bus_sync_axi_bus_reg_data1_40__FF_INPUT) );
  AND2X2 AND2X2_108 ( .A(RST), .B(A_ADDR_9_), .Y(bus_sync_axi_bus_reg_data1_41__FF_INPUT) );
  AND2X2 AND2X2_109 ( .A(RST), .B(A_ADDR_10_), .Y(bus_sync_axi_bus_reg_data1_42__FF_INPUT) );
  AND2X2 AND2X2_11 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_8_), .Y(bus_sync_axi_bus_reg_data3_8__FF_INPUT) );
  AND2X2 AND2X2_110 ( .A(RST), .B(A_ADDR_11_), .Y(bus_sync_axi_bus_reg_data1_43__FF_INPUT) );
  AND2X2 AND2X2_111 ( .A(RST), .B(A_ADDR_12_), .Y(bus_sync_axi_bus_reg_data1_44__FF_INPUT) );
  AND2X2 AND2X2_112 ( .A(RST), .B(A_ADDR_13_), .Y(bus_sync_axi_bus_reg_data1_45__FF_INPUT) );
  AND2X2 AND2X2_113 ( .A(RST), .B(A_ADDR_14_), .Y(bus_sync_axi_bus_reg_data1_46__FF_INPUT) );
  AND2X2 AND2X2_114 ( .A(RST), .B(A_ADDR_15_), .Y(bus_sync_axi_bus_reg_data1_47__FF_INPUT) );
  AND2X2 AND2X2_115 ( .A(RST), .B(A_ADDR_16_), .Y(bus_sync_axi_bus_reg_data1_48__FF_INPUT) );
  AND2X2 AND2X2_116 ( .A(RST), .B(A_ADDR_17_), .Y(bus_sync_axi_bus_reg_data1_49__FF_INPUT) );
  AND2X2 AND2X2_117 ( .A(RST), .B(A_ADDR_18_), .Y(bus_sync_axi_bus_reg_data1_50__FF_INPUT) );
  AND2X2 AND2X2_118 ( .A(RST), .B(A_ADDR_19_), .Y(bus_sync_axi_bus_reg_data1_51__FF_INPUT) );
  AND2X2 AND2X2_119 ( .A(RST), .B(A_ADDR_20_), .Y(bus_sync_axi_bus_reg_data1_52__FF_INPUT) );
  AND2X2 AND2X2_12 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_9_), .Y(bus_sync_axi_bus_reg_data3_9__FF_INPUT) );
  AND2X2 AND2X2_120 ( .A(RST), .B(A_ADDR_21_), .Y(bus_sync_axi_bus_reg_data1_53__FF_INPUT) );
  AND2X2 AND2X2_121 ( .A(RST), .B(A_ADDR_22_), .Y(bus_sync_axi_bus_reg_data1_54__FF_INPUT) );
  AND2X2 AND2X2_122 ( .A(RST), .B(A_ADDR_23_), .Y(bus_sync_axi_bus_reg_data1_55__FF_INPUT) );
  AND2X2 AND2X2_123 ( .A(RST), .B(A_ADDR_24_), .Y(bus_sync_axi_bus_reg_data1_56__FF_INPUT) );
  AND2X2 AND2X2_124 ( .A(RST), .B(A_ADDR_25_), .Y(bus_sync_axi_bus_reg_data1_57__FF_INPUT) );
  AND2X2 AND2X2_125 ( .A(RST), .B(A_ADDR_26_), .Y(bus_sync_axi_bus_reg_data1_58__FF_INPUT) );
  AND2X2 AND2X2_126 ( .A(RST), .B(A_ADDR_27_), .Y(bus_sync_axi_bus_reg_data1_59__FF_INPUT) );
  AND2X2 AND2X2_127 ( .A(RST), .B(A_ADDR_28_), .Y(bus_sync_axi_bus_reg_data1_60__FF_INPUT) );
  AND2X2 AND2X2_128 ( .A(RST), .B(A_ADDR_29_), .Y(bus_sync_axi_bus_reg_data1_61__FF_INPUT) );
  AND2X2 AND2X2_129 ( .A(RST), .B(A_ADDR_30_), .Y(bus_sync_axi_bus_reg_data1_62__FF_INPUT) );
  AND2X2 AND2X2_13 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_10_), .Y(bus_sync_axi_bus_reg_data3_10__FF_INPUT) );
  AND2X2 AND2X2_130 ( .A(RST), .B(A_ADDR_31_), .Y(bus_sync_axi_bus_reg_data1_63__FF_INPUT) );
  AND2X2 AND2X2_131 ( .A(RST), .B(bus_sync_axi_bus_ECLK1), .Y(bus_sync_axi_bus_EECLK1_FF_INPUT) );
  AND2X2 AND2X2_132 ( .A(RST), .B(SCLK), .Y(bus_sync_axi_bus_ECLK1_FF_INPUT) );
  AND2X2 AND2X2_133 ( .A(RST), .B(bus_sync_rdata_data_in_0_), .Y(bus_sync_rdata_reg_data1_0__FF_INPUT) );
  AND2X2 AND2X2_134 ( .A(RST), .B(bus_sync_rdata_data_in_1_), .Y(bus_sync_rdata_reg_data1_1__FF_INPUT) );
  AND2X2 AND2X2_135 ( .A(RST), .B(bus_sync_rdata_data_in_2_), .Y(bus_sync_rdata_reg_data1_2__FF_INPUT) );
  AND2X2 AND2X2_136 ( .A(RST), .B(bus_sync_rdata_data_in_3_), .Y(bus_sync_rdata_reg_data1_3__FF_INPUT) );
  AND2X2 AND2X2_137 ( .A(RST), .B(bus_sync_rdata_data_in_4_), .Y(bus_sync_rdata_reg_data1_4__FF_INPUT) );
  AND2X2 AND2X2_138 ( .A(RST), .B(bus_sync_rdata_data_in_5_), .Y(bus_sync_rdata_reg_data1_5__FF_INPUT) );
  AND2X2 AND2X2_139 ( .A(RST), .B(bus_sync_rdata_data_in_6_), .Y(bus_sync_rdata_reg_data1_6__FF_INPUT) );
  AND2X2 AND2X2_14 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_11_), .Y(bus_sync_axi_bus_reg_data3_11__FF_INPUT) );
  AND2X2 AND2X2_140 ( .A(RST), .B(bus_sync_rdata_data_in_7_), .Y(bus_sync_rdata_reg_data1_7__FF_INPUT) );
  AND2X2 AND2X2_141 ( .A(RST), .B(bus_sync_rdata_data_in_8_), .Y(bus_sync_rdata_reg_data1_8__FF_INPUT) );
  AND2X2 AND2X2_142 ( .A(RST), .B(bus_sync_rdata_data_in_9_), .Y(bus_sync_rdata_reg_data1_9__FF_INPUT) );
  AND2X2 AND2X2_143 ( .A(RST), .B(bus_sync_rdata_data_in_10_), .Y(bus_sync_rdata_reg_data1_10__FF_INPUT) );
  AND2X2 AND2X2_144 ( .A(RST), .B(bus_sync_rdata_data_in_11_), .Y(bus_sync_rdata_reg_data1_11__FF_INPUT) );
  AND2X2 AND2X2_145 ( .A(RST), .B(bus_sync_rdata_data_in_12_), .Y(bus_sync_rdata_reg_data1_12__FF_INPUT) );
  AND2X2 AND2X2_146 ( .A(RST), .B(bus_sync_rdata_data_in_13_), .Y(bus_sync_rdata_reg_data1_13__FF_INPUT) );
  AND2X2 AND2X2_147 ( .A(RST), .B(bus_sync_rdata_data_in_14_), .Y(bus_sync_rdata_reg_data1_14__FF_INPUT) );
  AND2X2 AND2X2_148 ( .A(RST), .B(bus_sync_rdata_data_in_15_), .Y(bus_sync_rdata_reg_data1_15__FF_INPUT) );
  AND2X2 AND2X2_149 ( .A(RST), .B(bus_sync_rdata_data_in_16_), .Y(bus_sync_rdata_reg_data1_16__FF_INPUT) );
  AND2X2 AND2X2_15 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_12_), .Y(bus_sync_axi_bus_reg_data3_12__FF_INPUT) );
  AND2X2 AND2X2_150 ( .A(RST), .B(bus_sync_rdata_data_in_17_), .Y(bus_sync_rdata_reg_data1_17__FF_INPUT) );
  AND2X2 AND2X2_151 ( .A(RST), .B(bus_sync_rdata_data_in_18_), .Y(bus_sync_rdata_reg_data1_18__FF_INPUT) );
  AND2X2 AND2X2_152 ( .A(RST), .B(bus_sync_rdata_data_in_19_), .Y(bus_sync_rdata_reg_data1_19__FF_INPUT) );
  AND2X2 AND2X2_153 ( .A(RST), .B(bus_sync_rdata_data_in_20_), .Y(bus_sync_rdata_reg_data1_20__FF_INPUT) );
  AND2X2 AND2X2_154 ( .A(RST), .B(bus_sync_rdata_data_in_21_), .Y(bus_sync_rdata_reg_data1_21__FF_INPUT) );
  AND2X2 AND2X2_155 ( .A(RST), .B(bus_sync_rdata_data_in_22_), .Y(bus_sync_rdata_reg_data1_22__FF_INPUT) );
  AND2X2 AND2X2_156 ( .A(RST), .B(bus_sync_rdata_data_in_23_), .Y(bus_sync_rdata_reg_data1_23__FF_INPUT) );
  AND2X2 AND2X2_157 ( .A(RST), .B(bus_sync_rdata_data_in_24_), .Y(bus_sync_rdata_reg_data1_24__FF_INPUT) );
  AND2X2 AND2X2_158 ( .A(RST), .B(bus_sync_rdata_data_in_25_), .Y(bus_sync_rdata_reg_data1_25__FF_INPUT) );
  AND2X2 AND2X2_159 ( .A(RST), .B(bus_sync_rdata_data_in_26_), .Y(bus_sync_rdata_reg_data1_26__FF_INPUT) );
  AND2X2 AND2X2_16 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_13_), .Y(bus_sync_axi_bus_reg_data3_13__FF_INPUT) );
  AND2X2 AND2X2_160 ( .A(RST), .B(bus_sync_rdata_data_in_27_), .Y(bus_sync_rdata_reg_data1_27__FF_INPUT) );
  AND2X2 AND2X2_161 ( .A(RST), .B(bus_sync_rdata_data_in_28_), .Y(bus_sync_rdata_reg_data1_28__FF_INPUT) );
  AND2X2 AND2X2_162 ( .A(RST), .B(bus_sync_rdata_data_in_29_), .Y(bus_sync_rdata_reg_data1_29__FF_INPUT) );
  AND2X2 AND2X2_163 ( .A(RST), .B(bus_sync_rdata_data_in_30_), .Y(bus_sync_rdata_reg_data1_30__FF_INPUT) );
  AND2X2 AND2X2_164 ( .A(RST), .B(bus_sync_rdata_data_in_31_), .Y(bus_sync_rdata_reg_data1_31__FF_INPUT) );
  AND2X2 AND2X2_165 ( .A(bus_sync_rdata_reg_data2_0_), .B(RST), .Y(bus_sync_rdata_reg_data3_0__FF_INPUT) );
  AND2X2 AND2X2_166 ( .A(RST), .B(bus_sync_rdata_reg_data2_1_), .Y(bus_sync_rdata_reg_data3_1__FF_INPUT) );
  AND2X2 AND2X2_167 ( .A(RST), .B(bus_sync_rdata_reg_data2_2_), .Y(bus_sync_rdata_reg_data3_2__FF_INPUT) );
  AND2X2 AND2X2_168 ( .A(RST), .B(bus_sync_rdata_reg_data2_3_), .Y(bus_sync_rdata_reg_data3_3__FF_INPUT) );
  AND2X2 AND2X2_169 ( .A(RST), .B(bus_sync_rdata_reg_data2_4_), .Y(bus_sync_rdata_reg_data3_4__FF_INPUT) );
  AND2X2 AND2X2_17 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_14_), .Y(bus_sync_axi_bus_reg_data3_14__FF_INPUT) );
  AND2X2 AND2X2_170 ( .A(RST), .B(bus_sync_rdata_reg_data2_5_), .Y(bus_sync_rdata_reg_data3_5__FF_INPUT) );
  AND2X2 AND2X2_171 ( .A(RST), .B(bus_sync_rdata_reg_data2_6_), .Y(bus_sync_rdata_reg_data3_6__FF_INPUT) );
  AND2X2 AND2X2_172 ( .A(RST), .B(bus_sync_rdata_reg_data2_7_), .Y(bus_sync_rdata_reg_data3_7__FF_INPUT) );
  AND2X2 AND2X2_173 ( .A(RST), .B(bus_sync_rdata_reg_data2_8_), .Y(bus_sync_rdata_reg_data3_8__FF_INPUT) );
  AND2X2 AND2X2_174 ( .A(RST), .B(bus_sync_rdata_reg_data2_9_), .Y(bus_sync_rdata_reg_data3_9__FF_INPUT) );
  AND2X2 AND2X2_175 ( .A(RST), .B(bus_sync_rdata_reg_data2_10_), .Y(bus_sync_rdata_reg_data3_10__FF_INPUT) );
  AND2X2 AND2X2_176 ( .A(RST), .B(bus_sync_rdata_reg_data2_11_), .Y(bus_sync_rdata_reg_data3_11__FF_INPUT) );
  AND2X2 AND2X2_177 ( .A(RST), .B(bus_sync_rdata_reg_data2_12_), .Y(bus_sync_rdata_reg_data3_12__FF_INPUT) );
  AND2X2 AND2X2_178 ( .A(RST), .B(bus_sync_rdata_reg_data2_13_), .Y(bus_sync_rdata_reg_data3_13__FF_INPUT) );
  AND2X2 AND2X2_179 ( .A(RST), .B(bus_sync_rdata_reg_data2_14_), .Y(bus_sync_rdata_reg_data3_14__FF_INPUT) );
  AND2X2 AND2X2_18 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_15_), .Y(bus_sync_axi_bus_reg_data3_15__FF_INPUT) );
  AND2X2 AND2X2_180 ( .A(RST), .B(bus_sync_rdata_reg_data2_15_), .Y(bus_sync_rdata_reg_data3_15__FF_INPUT) );
  AND2X2 AND2X2_181 ( .A(RST), .B(bus_sync_rdata_reg_data2_16_), .Y(bus_sync_rdata_reg_data3_16__FF_INPUT) );
  AND2X2 AND2X2_182 ( .A(RST), .B(bus_sync_rdata_reg_data2_17_), .Y(bus_sync_rdata_reg_data3_17__FF_INPUT) );
  AND2X2 AND2X2_183 ( .A(RST), .B(bus_sync_rdata_reg_data2_18_), .Y(bus_sync_rdata_reg_data3_18__FF_INPUT) );
  AND2X2 AND2X2_184 ( .A(RST), .B(bus_sync_rdata_reg_data2_19_), .Y(bus_sync_rdata_reg_data3_19__FF_INPUT) );
  AND2X2 AND2X2_185 ( .A(RST), .B(bus_sync_rdata_reg_data2_20_), .Y(bus_sync_rdata_reg_data3_20__FF_INPUT) );
  AND2X2 AND2X2_186 ( .A(RST), .B(bus_sync_rdata_reg_data2_21_), .Y(bus_sync_rdata_reg_data3_21__FF_INPUT) );
  AND2X2 AND2X2_187 ( .A(RST), .B(bus_sync_rdata_reg_data2_22_), .Y(bus_sync_rdata_reg_data3_22__FF_INPUT) );
  AND2X2 AND2X2_188 ( .A(RST), .B(bus_sync_rdata_reg_data2_23_), .Y(bus_sync_rdata_reg_data3_23__FF_INPUT) );
  AND2X2 AND2X2_189 ( .A(RST), .B(bus_sync_rdata_reg_data2_24_), .Y(bus_sync_rdata_reg_data3_24__FF_INPUT) );
  AND2X2 AND2X2_19 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_16_), .Y(bus_sync_axi_bus_reg_data3_16__FF_INPUT) );
  AND2X2 AND2X2_190 ( .A(RST), .B(bus_sync_rdata_reg_data2_25_), .Y(bus_sync_rdata_reg_data3_25__FF_INPUT) );
  AND2X2 AND2X2_191 ( .A(RST), .B(bus_sync_rdata_reg_data2_26_), .Y(bus_sync_rdata_reg_data3_26__FF_INPUT) );
  AND2X2 AND2X2_192 ( .A(RST), .B(bus_sync_rdata_reg_data2_27_), .Y(bus_sync_rdata_reg_data3_27__FF_INPUT) );
  AND2X2 AND2X2_193 ( .A(RST), .B(bus_sync_rdata_reg_data2_28_), .Y(bus_sync_rdata_reg_data3_28__FF_INPUT) );
  AND2X2 AND2X2_194 ( .A(RST), .B(bus_sync_rdata_reg_data2_29_), .Y(bus_sync_rdata_reg_data3_29__FF_INPUT) );
  AND2X2 AND2X2_195 ( .A(RST), .B(bus_sync_rdata_reg_data2_30_), .Y(bus_sync_rdata_reg_data3_30__FF_INPUT) );
  AND2X2 AND2X2_196 ( .A(RST), .B(bus_sync_rdata_reg_data2_31_), .Y(bus_sync_rdata_reg_data3_31__FF_INPUT) );
  AND2X2 AND2X2_197 ( .A(RST), .B(bus_sync_rdata_ECLK2), .Y(bus_sync_rdata_EECLK2_FF_INPUT) );
  AND2X2 AND2X2_198 ( .A(RST), .B(SCLK), .Y(bus_sync_rdata_ECLK2_FF_INPUT) );
  AND2X2 AND2X2_199 ( .A(RST), .B(bus_sync_state_machine_reg_data2_0_), .Y(bus_sync_state_machine_reg_data3_0__FF_INPUT) );
  AND2X2 AND2X2_2 ( .A(RST), .B(counter_65_), .Y(fini_spi_FF_INPUT) );
  AND2X2 AND2X2_20 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_17_), .Y(bus_sync_axi_bus_reg_data3_17__FF_INPUT) );
  AND2X2 AND2X2_200 ( .A(RST), .B(bus_sync_state_machine_reg_data2_1_), .Y(bus_sync_state_machine_reg_data3_1__FF_INPUT) );
  AND2X2 AND2X2_201 ( .A(RST), .B(bus_sync_state_machine_reg_data2_2_), .Y(bus_sync_state_machine_reg_data3_2__FF_INPUT) );
  AND2X2 AND2X2_202 ( .A(RST), .B(bus_sync_state_machine_reg_data2_3_), .Y(bus_sync_state_machine_reg_data3_3__FF_INPUT) );
  AND2X2 AND2X2_203 ( .A(RST), .B(fini_spi), .Y(bus_sync_state_machine_reg_data1_0__FF_INPUT) );
  AND2X2 AND2X2_204 ( .A(RST), .B(re), .Y(bus_sync_state_machine_reg_data1_1__FF_INPUT) );
  AND2X2 AND2X2_205 ( .A(RST), .B(we), .Y(bus_sync_state_machine_reg_data1_2__FF_INPUT) );
  AND2X2 AND2X2_206 ( .A(RST), .B(PICORV_RST_SPI), .Y(bus_sync_state_machine_reg_data1_3__FF_INPUT) );
  AND2X2 AND2X2_207 ( .A(RST), .B(bus_sync_state_machine_ECLK1), .Y(bus_sync_state_machine_EECLK1_FF_INPUT) );
  AND2X2 AND2X2_208 ( .A(RST), .B(SCLK), .Y(bus_sync_state_machine_ECLK1_FF_INPUT) );
  AND2X2 AND2X2_209 ( .A(RST), .B(bus_sync_status_reg_data2_0_), .Y(bus_sync_status_reg_data3_0__FF_INPUT) );
  AND2X2 AND2X2_21 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_18_), .Y(bus_sync_axi_bus_reg_data3_18__FF_INPUT) );
  AND2X2 AND2X2_210 ( .A(RST), .B(bus_sync_status_reg_data2_1_), .Y(bus_sync_status_reg_data3_1__FF_INPUT) );
  AND2X2 AND2X2_211 ( .A(RST), .B(bus_sync_status_reg_data2_2_), .Y(bus_sync_status_reg_data3_2__FF_INPUT) );
  AND2X2 AND2X2_212 ( .A(RST), .B(busy), .Y(bus_sync_status_reg_data1_0__FF_INPUT) );
  AND2X2 AND2X2_213 ( .A(RST), .B(axi_awvalid), .Y(bus_sync_status_reg_data1_1__FF_INPUT) );
  AND2X2 AND2X2_214 ( .A(RST), .B(axi_arvalid), .Y(bus_sync_status_reg_data1_2__FF_INPUT) );
  AND2X2 AND2X2_215 ( .A(RST), .B(bus_sync_status_ECLK2), .Y(bus_sync_status_EECLK2_FF_INPUT) );
  AND2X2 AND2X2_216 ( .A(RST), .B(SCLK), .Y(bus_sync_status_ECLK2_FF_INPUT) );
  AND2X2 AND2X2_22 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_19_), .Y(bus_sync_axi_bus_reg_data3_19__FF_INPUT) );
  AND2X2 AND2X2_23 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_20_), .Y(bus_sync_axi_bus_reg_data3_20__FF_INPUT) );
  AND2X2 AND2X2_24 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_21_), .Y(bus_sync_axi_bus_reg_data3_21__FF_INPUT) );
  AND2X2 AND2X2_25 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_22_), .Y(bus_sync_axi_bus_reg_data3_22__FF_INPUT) );
  AND2X2 AND2X2_26 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_23_), .Y(bus_sync_axi_bus_reg_data3_23__FF_INPUT) );
  AND2X2 AND2X2_27 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_24_), .Y(bus_sync_axi_bus_reg_data3_24__FF_INPUT) );
  AND2X2 AND2X2_28 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_25_), .Y(bus_sync_axi_bus_reg_data3_25__FF_INPUT) );
  AND2X2 AND2X2_29 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_26_), .Y(bus_sync_axi_bus_reg_data3_26__FF_INPUT) );
  AND2X2 AND2X2_3 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_0_), .Y(bus_sync_axi_bus_reg_data3_0__FF_INPUT) );
  AND2X2 AND2X2_30 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_27_), .Y(bus_sync_axi_bus_reg_data3_27__FF_INPUT) );
  AND2X2 AND2X2_31 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_28_), .Y(bus_sync_axi_bus_reg_data3_28__FF_INPUT) );
  AND2X2 AND2X2_32 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_29_), .Y(bus_sync_axi_bus_reg_data3_29__FF_INPUT) );
  AND2X2 AND2X2_33 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_30_), .Y(bus_sync_axi_bus_reg_data3_30__FF_INPUT) );
  AND2X2 AND2X2_34 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_31_), .Y(bus_sync_axi_bus_reg_data3_31__FF_INPUT) );
  AND2X2 AND2X2_35 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_32_), .Y(bus_sync_axi_bus_reg_data3_32__FF_INPUT) );
  AND2X2 AND2X2_36 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_33_), .Y(bus_sync_axi_bus_reg_data3_33__FF_INPUT) );
  AND2X2 AND2X2_37 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_34_), .Y(bus_sync_axi_bus_reg_data3_34__FF_INPUT) );
  AND2X2 AND2X2_38 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_35_), .Y(bus_sync_axi_bus_reg_data3_35__FF_INPUT) );
  AND2X2 AND2X2_39 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_36_), .Y(bus_sync_axi_bus_reg_data3_36__FF_INPUT) );
  AND2X2 AND2X2_4 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_1_), .Y(bus_sync_axi_bus_reg_data3_1__FF_INPUT) );
  AND2X2 AND2X2_40 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_37_), .Y(bus_sync_axi_bus_reg_data3_37__FF_INPUT) );
  AND2X2 AND2X2_41 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_38_), .Y(bus_sync_axi_bus_reg_data3_38__FF_INPUT) );
  AND2X2 AND2X2_42 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_39_), .Y(bus_sync_axi_bus_reg_data3_39__FF_INPUT) );
  AND2X2 AND2X2_43 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_40_), .Y(bus_sync_axi_bus_reg_data3_40__FF_INPUT) );
  AND2X2 AND2X2_44 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_41_), .Y(bus_sync_axi_bus_reg_data3_41__FF_INPUT) );
  AND2X2 AND2X2_45 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_42_), .Y(bus_sync_axi_bus_reg_data3_42__FF_INPUT) );
  AND2X2 AND2X2_46 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_43_), .Y(bus_sync_axi_bus_reg_data3_43__FF_INPUT) );
  AND2X2 AND2X2_47 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_44_), .Y(bus_sync_axi_bus_reg_data3_44__FF_INPUT) );
  AND2X2 AND2X2_48 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_45_), .Y(bus_sync_axi_bus_reg_data3_45__FF_INPUT) );
  AND2X2 AND2X2_49 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_46_), .Y(bus_sync_axi_bus_reg_data3_46__FF_INPUT) );
  AND2X2 AND2X2_5 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_2_), .Y(bus_sync_axi_bus_reg_data3_2__FF_INPUT) );
  AND2X2 AND2X2_50 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_47_), .Y(bus_sync_axi_bus_reg_data3_47__FF_INPUT) );
  AND2X2 AND2X2_51 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_48_), .Y(bus_sync_axi_bus_reg_data3_48__FF_INPUT) );
  AND2X2 AND2X2_52 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_49_), .Y(bus_sync_axi_bus_reg_data3_49__FF_INPUT) );
  AND2X2 AND2X2_53 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_50_), .Y(bus_sync_axi_bus_reg_data3_50__FF_INPUT) );
  AND2X2 AND2X2_54 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_51_), .Y(bus_sync_axi_bus_reg_data3_51__FF_INPUT) );
  AND2X2 AND2X2_55 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_52_), .Y(bus_sync_axi_bus_reg_data3_52__FF_INPUT) );
  AND2X2 AND2X2_56 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_53_), .Y(bus_sync_axi_bus_reg_data3_53__FF_INPUT) );
  AND2X2 AND2X2_57 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_54_), .Y(bus_sync_axi_bus_reg_data3_54__FF_INPUT) );
  AND2X2 AND2X2_58 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_55_), .Y(bus_sync_axi_bus_reg_data3_55__FF_INPUT) );
  AND2X2 AND2X2_59 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_56_), .Y(bus_sync_axi_bus_reg_data3_56__FF_INPUT) );
  AND2X2 AND2X2_6 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_3_), .Y(bus_sync_axi_bus_reg_data3_3__FF_INPUT) );
  AND2X2 AND2X2_60 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_57_), .Y(bus_sync_axi_bus_reg_data3_57__FF_INPUT) );
  AND2X2 AND2X2_61 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_58_), .Y(bus_sync_axi_bus_reg_data3_58__FF_INPUT) );
  AND2X2 AND2X2_62 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_59_), .Y(bus_sync_axi_bus_reg_data3_59__FF_INPUT) );
  AND2X2 AND2X2_63 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_60_), .Y(bus_sync_axi_bus_reg_data3_60__FF_INPUT) );
  AND2X2 AND2X2_64 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_61_), .Y(bus_sync_axi_bus_reg_data3_61__FF_INPUT) );
  AND2X2 AND2X2_65 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_62_), .Y(bus_sync_axi_bus_reg_data3_62__FF_INPUT) );
  AND2X2 AND2X2_66 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_63_), .Y(bus_sync_axi_bus_reg_data3_63__FF_INPUT) );
  AND2X2 AND2X2_67 ( .A(RST), .B(WDATA_0_), .Y(bus_sync_axi_bus_reg_data1_0__FF_INPUT) );
  AND2X2 AND2X2_68 ( .A(RST), .B(WDATA_1_), .Y(bus_sync_axi_bus_reg_data1_1__FF_INPUT) );
  AND2X2 AND2X2_69 ( .A(RST), .B(WDATA_2_), .Y(bus_sync_axi_bus_reg_data1_2__FF_INPUT) );
  AND2X2 AND2X2_7 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_4_), .Y(bus_sync_axi_bus_reg_data3_4__FF_INPUT) );
  AND2X2 AND2X2_70 ( .A(RST), .B(WDATA_3_), .Y(bus_sync_axi_bus_reg_data1_3__FF_INPUT) );
  AND2X2 AND2X2_71 ( .A(RST), .B(WDATA_4_), .Y(bus_sync_axi_bus_reg_data1_4__FF_INPUT) );
  AND2X2 AND2X2_72 ( .A(RST), .B(WDATA_5_), .Y(bus_sync_axi_bus_reg_data1_5__FF_INPUT) );
  AND2X2 AND2X2_73 ( .A(RST), .B(WDATA_6_), .Y(bus_sync_axi_bus_reg_data1_6__FF_INPUT) );
  AND2X2 AND2X2_74 ( .A(RST), .B(WDATA_7_), .Y(bus_sync_axi_bus_reg_data1_7__FF_INPUT) );
  AND2X2 AND2X2_75 ( .A(RST), .B(WDATA_8_), .Y(bus_sync_axi_bus_reg_data1_8__FF_INPUT) );
  AND2X2 AND2X2_76 ( .A(RST), .B(WDATA_9_), .Y(bus_sync_axi_bus_reg_data1_9__FF_INPUT) );
  AND2X2 AND2X2_77 ( .A(RST), .B(WDATA_10_), .Y(bus_sync_axi_bus_reg_data1_10__FF_INPUT) );
  AND2X2 AND2X2_78 ( .A(RST), .B(WDATA_11_), .Y(bus_sync_axi_bus_reg_data1_11__FF_INPUT) );
  AND2X2 AND2X2_79 ( .A(RST), .B(WDATA_12_), .Y(bus_sync_axi_bus_reg_data1_12__FF_INPUT) );
  AND2X2 AND2X2_8 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_5_), .Y(bus_sync_axi_bus_reg_data3_5__FF_INPUT) );
  AND2X2 AND2X2_80 ( .A(RST), .B(WDATA_13_), .Y(bus_sync_axi_bus_reg_data1_13__FF_INPUT) );
  AND2X2 AND2X2_81 ( .A(RST), .B(WDATA_14_), .Y(bus_sync_axi_bus_reg_data1_14__FF_INPUT) );
  AND2X2 AND2X2_82 ( .A(RST), .B(WDATA_15_), .Y(bus_sync_axi_bus_reg_data1_15__FF_INPUT) );
  AND2X2 AND2X2_83 ( .A(RST), .B(WDATA_16_), .Y(bus_sync_axi_bus_reg_data1_16__FF_INPUT) );
  AND2X2 AND2X2_84 ( .A(RST), .B(WDATA_17_), .Y(bus_sync_axi_bus_reg_data1_17__FF_INPUT) );
  AND2X2 AND2X2_85 ( .A(RST), .B(WDATA_18_), .Y(bus_sync_axi_bus_reg_data1_18__FF_INPUT) );
  AND2X2 AND2X2_86 ( .A(RST), .B(WDATA_19_), .Y(bus_sync_axi_bus_reg_data1_19__FF_INPUT) );
  AND2X2 AND2X2_87 ( .A(RST), .B(WDATA_20_), .Y(bus_sync_axi_bus_reg_data1_20__FF_INPUT) );
  AND2X2 AND2X2_88 ( .A(RST), .B(WDATA_21_), .Y(bus_sync_axi_bus_reg_data1_21__FF_INPUT) );
  AND2X2 AND2X2_89 ( .A(RST), .B(WDATA_22_), .Y(bus_sync_axi_bus_reg_data1_22__FF_INPUT) );
  AND2X2 AND2X2_9 ( .A(RST), .B(bus_sync_axi_bus_reg_data2_6_), .Y(bus_sync_axi_bus_reg_data3_6__FF_INPUT) );
  AND2X2 AND2X2_90 ( .A(RST), .B(WDATA_23_), .Y(bus_sync_axi_bus_reg_data1_23__FF_INPUT) );
  AND2X2 AND2X2_91 ( .A(RST), .B(WDATA_24_), .Y(bus_sync_axi_bus_reg_data1_24__FF_INPUT) );
  AND2X2 AND2X2_92 ( .A(RST), .B(WDATA_25_), .Y(bus_sync_axi_bus_reg_data1_25__FF_INPUT) );
  AND2X2 AND2X2_93 ( .A(RST), .B(WDATA_26_), .Y(bus_sync_axi_bus_reg_data1_26__FF_INPUT) );
  AND2X2 AND2X2_94 ( .A(RST), .B(WDATA_27_), .Y(bus_sync_axi_bus_reg_data1_27__FF_INPUT) );
  AND2X2 AND2X2_95 ( .A(RST), .B(WDATA_28_), .Y(bus_sync_axi_bus_reg_data1_28__FF_INPUT) );
  AND2X2 AND2X2_96 ( .A(RST), .B(WDATA_29_), .Y(bus_sync_axi_bus_reg_data1_29__FF_INPUT) );
  AND2X2 AND2X2_97 ( .A(RST), .B(WDATA_30_), .Y(bus_sync_axi_bus_reg_data1_30__FF_INPUT) );
  AND2X2 AND2X2_98 ( .A(RST), .B(WDATA_31_), .Y(bus_sync_axi_bus_reg_data1_31__FF_INPUT) );
  AND2X2 AND2X2_99 ( .A(RST), .B(A_ADDR_0_), .Y(bus_sync_axi_bus_reg_data1_32__FF_INPUT) );
  AOI21X1 AOI21X1_1 ( .A(_abc_4108_n566), .B(_abc_4108_n565), .C(_abc_4108_n561), .Y(_abc_2913_n87) );
  AOI21X1 AOI21X1_10 ( .A(_abc_4108_n712), .B(_abc_4108_n708), .C(_abc_4108_n561), .Y(bus_cap_7__FF_INPUT) );
  AOI21X1 AOI21X1_100 ( .A(CEB), .B(_abc_4108_n1152), .C(_abc_4108_n1056), .Y(sft_reg_0__FF_INPUT) );
  AOI21X1 AOI21X1_101 ( .A(CEB), .B(_abc_4108_n1154), .C(_abc_4108_n1060), .Y(sft_reg_1__FF_INPUT) );
  AOI21X1 AOI21X1_102 ( .A(CEB), .B(_abc_4108_n1156), .C(_abc_4108_n1063), .Y(sft_reg_2__FF_INPUT) );
  AOI21X1 AOI21X1_103 ( .A(CEB), .B(_abc_4108_n1158), .C(_abc_4108_n1066), .Y(sft_reg_3__FF_INPUT) );
  AOI21X1 AOI21X1_104 ( .A(CEB), .B(_abc_4108_n1160), .C(_abc_4108_n1069), .Y(sft_reg_4__FF_INPUT) );
  AOI21X1 AOI21X1_105 ( .A(CEB), .B(_abc_4108_n1162), .C(_abc_4108_n1072), .Y(sft_reg_5__FF_INPUT) );
  AOI21X1 AOI21X1_106 ( .A(CEB), .B(_abc_4108_n1164), .C(_abc_4108_n1075), .Y(sft_reg_6__FF_INPUT) );
  AOI21X1 AOI21X1_107 ( .A(CEB), .B(_abc_4108_n1166), .C(_abc_4108_n1078), .Y(sft_reg_7__FF_INPUT) );
  AOI21X1 AOI21X1_108 ( .A(CEB), .B(_abc_4108_n1168), .C(_abc_4108_n1081), .Y(sft_reg_8__FF_INPUT) );
  AOI21X1 AOI21X1_109 ( .A(CEB), .B(_abc_4108_n1170), .C(_abc_4108_n1084), .Y(sft_reg_9__FF_INPUT) );
  AOI21X1 AOI21X1_11 ( .A(_abc_4108_n718_1), .B(_abc_4108_n714_1), .C(_abc_4108_n561), .Y(bus_cap_8__FF_INPUT) );
  AOI21X1 AOI21X1_110 ( .A(CEB), .B(_abc_4108_n1172), .C(_abc_4108_n1087), .Y(sft_reg_10__FF_INPUT) );
  AOI21X1 AOI21X1_111 ( .A(CEB), .B(_abc_4108_n1174), .C(_abc_4108_n1090), .Y(sft_reg_11__FF_INPUT) );
  AOI21X1 AOI21X1_112 ( .A(CEB), .B(_abc_4108_n1176), .C(_abc_4108_n1093), .Y(sft_reg_12__FF_INPUT) );
  AOI21X1 AOI21X1_113 ( .A(CEB), .B(_abc_4108_n1178), .C(_abc_4108_n1096), .Y(sft_reg_13__FF_INPUT) );
  AOI21X1 AOI21X1_114 ( .A(CEB), .B(_abc_4108_n1180), .C(_abc_4108_n1099), .Y(sft_reg_14__FF_INPUT) );
  AOI21X1 AOI21X1_115 ( .A(CEB), .B(_abc_4108_n1182), .C(_abc_4108_n1102), .Y(sft_reg_15__FF_INPUT) );
  AOI21X1 AOI21X1_116 ( .A(CEB), .B(_abc_4108_n1184), .C(_abc_4108_n1105), .Y(sft_reg_16__FF_INPUT) );
  AOI21X1 AOI21X1_117 ( .A(CEB), .B(_abc_4108_n1186), .C(_abc_4108_n1108), .Y(sft_reg_17__FF_INPUT) );
  AOI21X1 AOI21X1_118 ( .A(CEB), .B(_abc_4108_n1188), .C(_abc_4108_n1111), .Y(sft_reg_18__FF_INPUT) );
  AOI21X1 AOI21X1_119 ( .A(CEB), .B(_abc_4108_n1190), .C(_abc_4108_n1114), .Y(sft_reg_19__FF_INPUT) );
  AOI21X1 AOI21X1_12 ( .A(_abc_4108_n724), .B(_abc_4108_n720), .C(_abc_4108_n561), .Y(bus_cap_9__FF_INPUT) );
  AOI21X1 AOI21X1_120 ( .A(CEB), .B(_abc_4108_n1192), .C(_abc_4108_n1117), .Y(sft_reg_20__FF_INPUT) );
  AOI21X1 AOI21X1_121 ( .A(CEB), .B(_abc_4108_n1194), .C(_abc_4108_n1120), .Y(sft_reg_21__FF_INPUT) );
  AOI21X1 AOI21X1_122 ( .A(CEB), .B(_abc_4108_n1196), .C(_abc_4108_n1123), .Y(sft_reg_22__FF_INPUT) );
  AOI21X1 AOI21X1_123 ( .A(CEB), .B(_abc_4108_n1198), .C(_abc_4108_n1126), .Y(sft_reg_23__FF_INPUT) );
  AOI21X1 AOI21X1_124 ( .A(CEB), .B(_abc_4108_n1200), .C(_abc_4108_n1129), .Y(sft_reg_24__FF_INPUT) );
  AOI21X1 AOI21X1_125 ( .A(CEB), .B(_abc_4108_n1202), .C(_abc_4108_n1132), .Y(sft_reg_25__FF_INPUT) );
  AOI21X1 AOI21X1_126 ( .A(CEB), .B(_abc_4108_n1204), .C(_abc_4108_n1135), .Y(sft_reg_26__FF_INPUT) );
  AOI21X1 AOI21X1_127 ( .A(CEB), .B(_abc_4108_n1206), .C(_abc_4108_n1138), .Y(sft_reg_27__FF_INPUT) );
  AOI21X1 AOI21X1_128 ( .A(CEB), .B(_abc_4108_n1208), .C(_abc_4108_n1141), .Y(sft_reg_28__FF_INPUT) );
  AOI21X1 AOI21X1_129 ( .A(CEB), .B(_abc_4108_n1210), .C(_abc_4108_n1144), .Y(sft_reg_29__FF_INPUT) );
  AOI21X1 AOI21X1_13 ( .A(_abc_4108_n730_1), .B(_abc_4108_n726_1), .C(_abc_4108_n561), .Y(bus_cap_10__FF_INPUT) );
  AOI21X1 AOI21X1_130 ( .A(CEB), .B(_abc_4108_n1212), .C(_abc_4108_n1147), .Y(sft_reg_30__FF_INPUT) );
  AOI21X1 AOI21X1_131 ( .A(_abc_4108_n1333), .B(_abc_4108_n1335), .C(_abc_4108_n1336), .Y(PICORV_RST_SPI_FF_INPUT) );
  AOI21X1 AOI21X1_132 ( .A(_abc_4108_n599_1), .B(_abc_4108_n1338), .C(_abc_4108_n1339), .Y(re_FF_INPUT) );
  AOI21X1 AOI21X1_133 ( .A(_abc_4108_n595), .B(_abc_4108_n1215), .C(_abc_4108_n1343), .Y(we_FF_INPUT) );
  AOI21X1 AOI21X1_134 ( .A(bus_sync_axi_bus__abc_3782_n457), .B(bus_sync_axi_bus_EECLK1), .C(bus_sync_axi_bus__abc_3782_n458), .Y(bus_sync_axi_bus_reg_data2_0__FF_INPUT) );
  AOI21X1 AOI21X1_135 ( .A(bus_sync_axi_bus__abc_3782_n462), .B(bus_sync_axi_bus__abc_3782_n463), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_1__FF_INPUT) );
  AOI21X1 AOI21X1_136 ( .A(bus_sync_axi_bus__abc_3782_n465), .B(bus_sync_axi_bus__abc_3782_n466), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_2__FF_INPUT) );
  AOI21X1 AOI21X1_137 ( .A(bus_sync_axi_bus__abc_3782_n468), .B(bus_sync_axi_bus__abc_3782_n469), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_3__FF_INPUT) );
  AOI21X1 AOI21X1_138 ( .A(bus_sync_axi_bus__abc_3782_n471), .B(bus_sync_axi_bus__abc_3782_n472), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_4__FF_INPUT) );
  AOI21X1 AOI21X1_139 ( .A(bus_sync_axi_bus__abc_3782_n474), .B(bus_sync_axi_bus__abc_3782_n475), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_5__FF_INPUT) );
  AOI21X1 AOI21X1_14 ( .A(_abc_4108_n736), .B(_abc_4108_n732), .C(_abc_4108_n561), .Y(bus_cap_11__FF_INPUT) );
  AOI21X1 AOI21X1_140 ( .A(bus_sync_axi_bus__abc_3782_n477), .B(bus_sync_axi_bus__abc_3782_n478), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_6__FF_INPUT) );
  AOI21X1 AOI21X1_141 ( .A(bus_sync_axi_bus__abc_3782_n480), .B(bus_sync_axi_bus__abc_3782_n481), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_7__FF_INPUT) );
  AOI21X1 AOI21X1_142 ( .A(bus_sync_axi_bus__abc_3782_n483), .B(bus_sync_axi_bus__abc_3782_n484), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_8__FF_INPUT) );
  AOI21X1 AOI21X1_143 ( .A(bus_sync_axi_bus__abc_3782_n486), .B(bus_sync_axi_bus__abc_3782_n487), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_9__FF_INPUT) );
  AOI21X1 AOI21X1_144 ( .A(bus_sync_axi_bus__abc_3782_n489), .B(bus_sync_axi_bus__abc_3782_n490), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_10__FF_INPUT) );
  AOI21X1 AOI21X1_145 ( .A(bus_sync_axi_bus__abc_3782_n492), .B(bus_sync_axi_bus__abc_3782_n493), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_11__FF_INPUT) );
  AOI21X1 AOI21X1_146 ( .A(bus_sync_axi_bus__abc_3782_n495), .B(bus_sync_axi_bus__abc_3782_n496), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_12__FF_INPUT) );
  AOI21X1 AOI21X1_147 ( .A(bus_sync_axi_bus__abc_3782_n498), .B(bus_sync_axi_bus__abc_3782_n499), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_13__FF_INPUT) );
  AOI21X1 AOI21X1_148 ( .A(bus_sync_axi_bus__abc_3782_n501), .B(bus_sync_axi_bus__abc_3782_n502), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_14__FF_INPUT) );
  AOI21X1 AOI21X1_149 ( .A(bus_sync_axi_bus__abc_3782_n504), .B(bus_sync_axi_bus__abc_3782_n505), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_15__FF_INPUT) );
  AOI21X1 AOI21X1_15 ( .A(_abc_4108_n742_1), .B(_abc_4108_n738_1), .C(_abc_4108_n561), .Y(bus_cap_12__FF_INPUT) );
  AOI21X1 AOI21X1_150 ( .A(bus_sync_axi_bus__abc_3782_n507), .B(bus_sync_axi_bus__abc_3782_n508), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_16__FF_INPUT) );
  AOI21X1 AOI21X1_151 ( .A(bus_sync_axi_bus__abc_3782_n510), .B(bus_sync_axi_bus__abc_3782_n511), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_17__FF_INPUT) );
  AOI21X1 AOI21X1_152 ( .A(bus_sync_axi_bus__abc_3782_n513), .B(bus_sync_axi_bus__abc_3782_n514), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_18__FF_INPUT) );
  AOI21X1 AOI21X1_153 ( .A(bus_sync_axi_bus__abc_3782_n516), .B(bus_sync_axi_bus__abc_3782_n517), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_19__FF_INPUT) );
  AOI21X1 AOI21X1_154 ( .A(bus_sync_axi_bus__abc_3782_n519), .B(bus_sync_axi_bus__abc_3782_n520), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_20__FF_INPUT) );
  AOI21X1 AOI21X1_155 ( .A(bus_sync_axi_bus__abc_3782_n522), .B(bus_sync_axi_bus__abc_3782_n523), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_21__FF_INPUT) );
  AOI21X1 AOI21X1_156 ( .A(bus_sync_axi_bus__abc_3782_n525), .B(bus_sync_axi_bus__abc_3782_n526), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_22__FF_INPUT) );
  AOI21X1 AOI21X1_157 ( .A(bus_sync_axi_bus__abc_3782_n528), .B(bus_sync_axi_bus__abc_3782_n529), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_23__FF_INPUT) );
  AOI21X1 AOI21X1_158 ( .A(bus_sync_axi_bus__abc_3782_n531), .B(bus_sync_axi_bus__abc_3782_n532), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_24__FF_INPUT) );
  AOI21X1 AOI21X1_159 ( .A(bus_sync_axi_bus__abc_3782_n534), .B(bus_sync_axi_bus__abc_3782_n535), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_25__FF_INPUT) );
  AOI21X1 AOI21X1_16 ( .A(_abc_4108_n748), .B(_abc_4108_n744), .C(_abc_4108_n561), .Y(bus_cap_13__FF_INPUT) );
  AOI21X1 AOI21X1_160 ( .A(bus_sync_axi_bus__abc_3782_n537), .B(bus_sync_axi_bus__abc_3782_n538), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_26__FF_INPUT) );
  AOI21X1 AOI21X1_161 ( .A(bus_sync_axi_bus__abc_3782_n540), .B(bus_sync_axi_bus__abc_3782_n541), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_27__FF_INPUT) );
  AOI21X1 AOI21X1_162 ( .A(bus_sync_axi_bus__abc_3782_n543), .B(bus_sync_axi_bus__abc_3782_n544), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_28__FF_INPUT) );
  AOI21X1 AOI21X1_163 ( .A(bus_sync_axi_bus__abc_3782_n546), .B(bus_sync_axi_bus__abc_3782_n547), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_29__FF_INPUT) );
  AOI21X1 AOI21X1_164 ( .A(bus_sync_axi_bus__abc_3782_n549), .B(bus_sync_axi_bus__abc_3782_n550), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_30__FF_INPUT) );
  AOI21X1 AOI21X1_165 ( .A(bus_sync_axi_bus__abc_3782_n552), .B(bus_sync_axi_bus__abc_3782_n553), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_31__FF_INPUT) );
  AOI21X1 AOI21X1_166 ( .A(bus_sync_axi_bus__abc_3782_n555), .B(bus_sync_axi_bus__abc_3782_n556), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_32__FF_INPUT) );
  AOI21X1 AOI21X1_167 ( .A(bus_sync_axi_bus__abc_3782_n558), .B(bus_sync_axi_bus__abc_3782_n559), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_33__FF_INPUT) );
  AOI21X1 AOI21X1_168 ( .A(bus_sync_axi_bus__abc_3782_n561), .B(bus_sync_axi_bus__abc_3782_n562), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_34__FF_INPUT) );
  AOI21X1 AOI21X1_169 ( .A(bus_sync_axi_bus__abc_3782_n564), .B(bus_sync_axi_bus__abc_3782_n565), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_35__FF_INPUT) );
  AOI21X1 AOI21X1_17 ( .A(_abc_4108_n754_1), .B(_abc_4108_n750_1), .C(_abc_4108_n561), .Y(bus_cap_14__FF_INPUT) );
  AOI21X1 AOI21X1_170 ( .A(bus_sync_axi_bus__abc_3782_n567), .B(bus_sync_axi_bus__abc_3782_n568), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_36__FF_INPUT) );
  AOI21X1 AOI21X1_171 ( .A(bus_sync_axi_bus__abc_3782_n570), .B(bus_sync_axi_bus__abc_3782_n571), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_37__FF_INPUT) );
  AOI21X1 AOI21X1_172 ( .A(bus_sync_axi_bus__abc_3782_n573), .B(bus_sync_axi_bus__abc_3782_n574), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_38__FF_INPUT) );
  AOI21X1 AOI21X1_173 ( .A(bus_sync_axi_bus__abc_3782_n576), .B(bus_sync_axi_bus__abc_3782_n577), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_39__FF_INPUT) );
  AOI21X1 AOI21X1_174 ( .A(bus_sync_axi_bus__abc_3782_n579), .B(bus_sync_axi_bus__abc_3782_n580), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_40__FF_INPUT) );
  AOI21X1 AOI21X1_175 ( .A(bus_sync_axi_bus__abc_3782_n582), .B(bus_sync_axi_bus__abc_3782_n583), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_41__FF_INPUT) );
  AOI21X1 AOI21X1_176 ( .A(bus_sync_axi_bus__abc_3782_n585), .B(bus_sync_axi_bus__abc_3782_n586), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_42__FF_INPUT) );
  AOI21X1 AOI21X1_177 ( .A(bus_sync_axi_bus__abc_3782_n588), .B(bus_sync_axi_bus__abc_3782_n589), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_43__FF_INPUT) );
  AOI21X1 AOI21X1_178 ( .A(bus_sync_axi_bus__abc_3782_n591), .B(bus_sync_axi_bus__abc_3782_n592), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_44__FF_INPUT) );
  AOI21X1 AOI21X1_179 ( .A(bus_sync_axi_bus__abc_3782_n594), .B(bus_sync_axi_bus__abc_3782_n595), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_45__FF_INPUT) );
  AOI21X1 AOI21X1_18 ( .A(_abc_4108_n760), .B(_abc_4108_n756), .C(_abc_4108_n561), .Y(bus_cap_15__FF_INPUT) );
  AOI21X1 AOI21X1_180 ( .A(bus_sync_axi_bus__abc_3782_n597), .B(bus_sync_axi_bus__abc_3782_n598), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_46__FF_INPUT) );
  AOI21X1 AOI21X1_181 ( .A(bus_sync_axi_bus__abc_3782_n600), .B(bus_sync_axi_bus__abc_3782_n601), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_47__FF_INPUT) );
  AOI21X1 AOI21X1_182 ( .A(bus_sync_axi_bus__abc_3782_n603), .B(bus_sync_axi_bus__abc_3782_n604), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_48__FF_INPUT) );
  AOI21X1 AOI21X1_183 ( .A(bus_sync_axi_bus__abc_3782_n606), .B(bus_sync_axi_bus__abc_3782_n607), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_49__FF_INPUT) );
  AOI21X1 AOI21X1_184 ( .A(bus_sync_axi_bus__abc_3782_n609), .B(bus_sync_axi_bus__abc_3782_n610), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_50__FF_INPUT) );
  AOI21X1 AOI21X1_185 ( .A(bus_sync_axi_bus__abc_3782_n612), .B(bus_sync_axi_bus__abc_3782_n613), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_51__FF_INPUT) );
  AOI21X1 AOI21X1_186 ( .A(bus_sync_axi_bus__abc_3782_n615), .B(bus_sync_axi_bus__abc_3782_n616), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_52__FF_INPUT) );
  AOI21X1 AOI21X1_187 ( .A(bus_sync_axi_bus__abc_3782_n618), .B(bus_sync_axi_bus__abc_3782_n619), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_53__FF_INPUT) );
  AOI21X1 AOI21X1_188 ( .A(bus_sync_axi_bus__abc_3782_n621), .B(bus_sync_axi_bus__abc_3782_n622), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_54__FF_INPUT) );
  AOI21X1 AOI21X1_189 ( .A(bus_sync_axi_bus__abc_3782_n624), .B(bus_sync_axi_bus__abc_3782_n625), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_55__FF_INPUT) );
  AOI21X1 AOI21X1_19 ( .A(_abc_4108_n766), .B(_abc_4108_n762), .C(_abc_4108_n561), .Y(bus_cap_16__FF_INPUT) );
  AOI21X1 AOI21X1_190 ( .A(bus_sync_axi_bus__abc_3782_n627), .B(bus_sync_axi_bus__abc_3782_n628), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_56__FF_INPUT) );
  AOI21X1 AOI21X1_191 ( .A(bus_sync_axi_bus__abc_3782_n630), .B(bus_sync_axi_bus__abc_3782_n631), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_57__FF_INPUT) );
  AOI21X1 AOI21X1_192 ( .A(bus_sync_axi_bus__abc_3782_n633), .B(bus_sync_axi_bus__abc_3782_n634), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_58__FF_INPUT) );
  AOI21X1 AOI21X1_193 ( .A(bus_sync_axi_bus__abc_3782_n636), .B(bus_sync_axi_bus__abc_3782_n637), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_59__FF_INPUT) );
  AOI21X1 AOI21X1_194 ( .A(bus_sync_axi_bus__abc_3782_n639), .B(bus_sync_axi_bus__abc_3782_n640), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_60__FF_INPUT) );
  AOI21X1 AOI21X1_195 ( .A(bus_sync_axi_bus__abc_3782_n642), .B(bus_sync_axi_bus__abc_3782_n643), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_61__FF_INPUT) );
  AOI21X1 AOI21X1_196 ( .A(bus_sync_axi_bus__abc_3782_n645), .B(bus_sync_axi_bus__abc_3782_n646), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_62__FF_INPUT) );
  AOI21X1 AOI21X1_197 ( .A(bus_sync_axi_bus__abc_3782_n648), .B(bus_sync_axi_bus__abc_3782_n649), .C(bus_sync_axi_bus__abc_3782_n460), .Y(bus_sync_axi_bus_reg_data2_63__FF_INPUT) );
  AOI21X1 AOI21X1_198 ( .A(bus_sync_rdata__abc_3590_n201_1), .B(bus_sync_rdata_EECLK2), .C(bus_sync_rdata__abc_3590_n202_1), .Y(bus_sync_rdata_reg_data2_0__FF_INPUT) );
  AOI21X1 AOI21X1_199 ( .A(bus_sync_rdata__abc_3590_n206_1), .B(bus_sync_rdata__abc_3590_n207_1), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_1__FF_INPUT) );
  AOI21X1 AOI21X1_2 ( .A(_abc_4108_n583_1), .B(state_1_), .C(_abc_4108_n561), .Y(_abc_4108_n584_1) );
  AOI21X1 AOI21X1_20 ( .A(_abc_4108_n772), .B(_abc_4108_n768), .C(_abc_4108_n561), .Y(bus_cap_17__FF_INPUT) );
  AOI21X1 AOI21X1_200 ( .A(bus_sync_rdata__abc_3590_n209_1), .B(bus_sync_rdata__abc_3590_n210_1), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_2__FF_INPUT) );
  AOI21X1 AOI21X1_201 ( .A(bus_sync_rdata__abc_3590_n212_1), .B(bus_sync_rdata__abc_3590_n213_1), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_3__FF_INPUT) );
  AOI21X1 AOI21X1_202 ( .A(bus_sync_rdata__abc_3590_n215_1), .B(bus_sync_rdata__abc_3590_n216_1), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_4__FF_INPUT) );
  AOI21X1 AOI21X1_203 ( .A(bus_sync_rdata__abc_3590_n218_1), .B(bus_sync_rdata__abc_3590_n219_1), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_5__FF_INPUT) );
  AOI21X1 AOI21X1_204 ( .A(bus_sync_rdata__abc_3590_n221_1), .B(bus_sync_rdata__abc_3590_n222_1), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_6__FF_INPUT) );
  AOI21X1 AOI21X1_205 ( .A(bus_sync_rdata__abc_3590_n224_1), .B(bus_sync_rdata__abc_3590_n225_1), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_7__FF_INPUT) );
  AOI21X1 AOI21X1_206 ( .A(bus_sync_rdata__abc_3590_n227_1), .B(bus_sync_rdata__abc_3590_n228_1), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_8__FF_INPUT) );
  AOI21X1 AOI21X1_207 ( .A(bus_sync_rdata__abc_3590_n230_1), .B(bus_sync_rdata__abc_3590_n231_1), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_9__FF_INPUT) );
  AOI21X1 AOI21X1_208 ( .A(bus_sync_rdata__abc_3590_n233), .B(bus_sync_rdata__abc_3590_n234), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_10__FF_INPUT) );
  AOI21X1 AOI21X1_209 ( .A(bus_sync_rdata__abc_3590_n236), .B(bus_sync_rdata__abc_3590_n237), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_11__FF_INPUT) );
  AOI21X1 AOI21X1_21 ( .A(_abc_4108_n778), .B(_abc_4108_n774), .C(_abc_4108_n561), .Y(bus_cap_18__FF_INPUT) );
  AOI21X1 AOI21X1_210 ( .A(bus_sync_rdata__abc_3590_n239), .B(bus_sync_rdata__abc_3590_n240), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_12__FF_INPUT) );
  AOI21X1 AOI21X1_211 ( .A(bus_sync_rdata__abc_3590_n242), .B(bus_sync_rdata__abc_3590_n243), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_13__FF_INPUT) );
  AOI21X1 AOI21X1_212 ( .A(bus_sync_rdata__abc_3590_n245), .B(bus_sync_rdata__abc_3590_n246), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_14__FF_INPUT) );
  AOI21X1 AOI21X1_213 ( .A(bus_sync_rdata__abc_3590_n248), .B(bus_sync_rdata__abc_3590_n249), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_15__FF_INPUT) );
  AOI21X1 AOI21X1_214 ( .A(bus_sync_rdata__abc_3590_n251), .B(bus_sync_rdata__abc_3590_n252), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_16__FF_INPUT) );
  AOI21X1 AOI21X1_215 ( .A(bus_sync_rdata__abc_3590_n254), .B(bus_sync_rdata__abc_3590_n255), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_17__FF_INPUT) );
  AOI21X1 AOI21X1_216 ( .A(bus_sync_rdata__abc_3590_n257), .B(bus_sync_rdata__abc_3590_n258), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_18__FF_INPUT) );
  AOI21X1 AOI21X1_217 ( .A(bus_sync_rdata__abc_3590_n260), .B(bus_sync_rdata__abc_3590_n261), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_19__FF_INPUT) );
  AOI21X1 AOI21X1_218 ( .A(bus_sync_rdata__abc_3590_n263), .B(bus_sync_rdata__abc_3590_n264), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_20__FF_INPUT) );
  AOI21X1 AOI21X1_219 ( .A(bus_sync_rdata__abc_3590_n266), .B(bus_sync_rdata__abc_3590_n267), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_21__FF_INPUT) );
  AOI21X1 AOI21X1_22 ( .A(_abc_4108_n784), .B(_abc_4108_n780), .C(_abc_4108_n561), .Y(bus_cap_19__FF_INPUT) );
  AOI21X1 AOI21X1_220 ( .A(bus_sync_rdata__abc_3590_n269), .B(bus_sync_rdata__abc_3590_n270), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_22__FF_INPUT) );
  AOI21X1 AOI21X1_221 ( .A(bus_sync_rdata__abc_3590_n272), .B(bus_sync_rdata__abc_3590_n273), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_23__FF_INPUT) );
  AOI21X1 AOI21X1_222 ( .A(bus_sync_rdata__abc_3590_n275), .B(bus_sync_rdata__abc_3590_n276), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_24__FF_INPUT) );
  AOI21X1 AOI21X1_223 ( .A(bus_sync_rdata__abc_3590_n278), .B(bus_sync_rdata__abc_3590_n279), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_25__FF_INPUT) );
  AOI21X1 AOI21X1_224 ( .A(bus_sync_rdata__abc_3590_n281), .B(bus_sync_rdata__abc_3590_n282), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_26__FF_INPUT) );
  AOI21X1 AOI21X1_225 ( .A(bus_sync_rdata__abc_3590_n284), .B(bus_sync_rdata__abc_3590_n285), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_27__FF_INPUT) );
  AOI21X1 AOI21X1_226 ( .A(bus_sync_rdata__abc_3590_n287), .B(bus_sync_rdata__abc_3590_n288), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_28__FF_INPUT) );
  AOI21X1 AOI21X1_227 ( .A(bus_sync_rdata__abc_3590_n290), .B(bus_sync_rdata__abc_3590_n291), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_29__FF_INPUT) );
  AOI21X1 AOI21X1_228 ( .A(bus_sync_rdata__abc_3590_n293), .B(bus_sync_rdata__abc_3590_n294), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_30__FF_INPUT) );
  AOI21X1 AOI21X1_229 ( .A(bus_sync_rdata__abc_3590_n296), .B(bus_sync_rdata__abc_3590_n297), .C(bus_sync_rdata__abc_3590_n204_1), .Y(bus_sync_rdata_reg_data2_31__FF_INPUT) );
  AOI21X1 AOI21X1_23 ( .A(_abc_4108_n790), .B(_abc_4108_n786), .C(_abc_4108_n561), .Y(bus_cap_20__FF_INPUT) );
  AOI21X1 AOI21X1_230 ( .A(bus_sync_state_machine__abc_3756_n37), .B(bus_sync_state_machine_EECLK1), .C(bus_sync_state_machine__abc_3756_n38), .Y(bus_sync_state_machine_reg_data2_0__FF_INPUT) );
  AOI21X1 AOI21X1_231 ( .A(bus_sync_state_machine__abc_3756_n42), .B(bus_sync_state_machine__abc_3756_n43), .C(bus_sync_state_machine__abc_3756_n40), .Y(bus_sync_state_machine_reg_data2_1__FF_INPUT) );
  AOI21X1 AOI21X1_232 ( .A(bus_sync_state_machine__abc_3756_n45), .B(bus_sync_state_machine__abc_3756_n46), .C(bus_sync_state_machine__abc_3756_n40), .Y(bus_sync_state_machine_reg_data2_2__FF_INPUT) );
  AOI21X1 AOI21X1_233 ( .A(bus_sync_state_machine__abc_3756_n48), .B(bus_sync_state_machine__abc_3756_n49), .C(bus_sync_state_machine__abc_3756_n40), .Y(bus_sync_state_machine_reg_data2_3__FF_INPUT) );
  AOI21X1 AOI21X1_234 ( .A(bus_sync_status__abc_3569_n30), .B(bus_sync_status_EECLK2), .C(bus_sync_status__abc_3569_n31), .Y(bus_sync_status_reg_data2_0__FF_INPUT) );
  AOI21X1 AOI21X1_235 ( .A(bus_sync_status__abc_3569_n35), .B(bus_sync_status__abc_3569_n36), .C(bus_sync_status__abc_3569_n33), .Y(bus_sync_status_reg_data2_1__FF_INPUT) );
  AOI21X1 AOI21X1_236 ( .A(bus_sync_status__abc_3569_n38), .B(bus_sync_status__abc_3569_n39), .C(bus_sync_status__abc_3569_n33), .Y(bus_sync_status_reg_data2_2__FF_INPUT) );
  AOI21X1 AOI21X1_24 ( .A(_abc_4108_n796), .B(_abc_4108_n792), .C(_abc_4108_n561), .Y(bus_cap_21__FF_INPUT) );
  AOI21X1 AOI21X1_25 ( .A(_abc_4108_n802), .B(_abc_4108_n798), .C(_abc_4108_n561), .Y(bus_cap_22__FF_INPUT) );
  AOI21X1 AOI21X1_26 ( .A(_abc_4108_n808), .B(_abc_4108_n804), .C(_abc_4108_n561), .Y(bus_cap_23__FF_INPUT) );
  AOI21X1 AOI21X1_27 ( .A(_abc_4108_n814), .B(_abc_4108_n810), .C(_abc_4108_n561), .Y(bus_cap_24__FF_INPUT) );
  AOI21X1 AOI21X1_28 ( .A(_abc_4108_n820_1), .B(_abc_4108_n816), .C(_abc_4108_n561), .Y(bus_cap_25__FF_INPUT) );
  AOI21X1 AOI21X1_29 ( .A(_abc_4108_n826), .B(_abc_4108_n822), .C(_abc_4108_n561), .Y(bus_cap_26__FF_INPUT) );
  AOI21X1 AOI21X1_3 ( .A(_abc_4108_n639), .B(_abc_4108_n601), .C(_abc_4108_n644), .Y(bus_cap_0__FF_INPUT) );
  AOI21X1 AOI21X1_30 ( .A(_abc_4108_n832), .B(_abc_4108_n828), .C(_abc_4108_n561), .Y(bus_cap_27__FF_INPUT) );
  AOI21X1 AOI21X1_31 ( .A(_abc_4108_n838), .B(_abc_4108_n834), .C(_abc_4108_n561), .Y(bus_cap_28__FF_INPUT) );
  AOI21X1 AOI21X1_32 ( .A(_abc_4108_n844), .B(_abc_4108_n840), .C(_abc_4108_n561), .Y(bus_cap_29__FF_INPUT) );
  AOI21X1 AOI21X1_33 ( .A(_abc_4108_n850), .B(_abc_4108_n846), .C(_abc_4108_n561), .Y(bus_cap_30__FF_INPUT) );
  AOI21X1 AOI21X1_34 ( .A(_abc_4108_n856), .B(_abc_4108_n852), .C(_abc_4108_n561), .Y(bus_cap_31__FF_INPUT) );
  AOI21X1 AOI21X1_35 ( .A(_abc_4108_n579_1), .B(_abc_4108_n858), .C(_abc_4108_n859_1), .Y(rdata_0__FF_INPUT) );
  AOI21X1 AOI21X1_36 ( .A(_abc_4108_n579_1), .B(_abc_4108_n861_1), .C(_abc_4108_n862), .Y(rdata_1__FF_INPUT) );
  AOI21X1 AOI21X1_37 ( .A(_abc_4108_n579_1), .B(_abc_4108_n864), .C(_abc_4108_n865_1), .Y(rdata_2__FF_INPUT) );
  AOI21X1 AOI21X1_38 ( .A(_abc_4108_n579_1), .B(_abc_4108_n867_1), .C(_abc_4108_n868), .Y(rdata_3__FF_INPUT) );
  AOI21X1 AOI21X1_39 ( .A(_abc_4108_n579_1), .B(_abc_4108_n870), .C(_abc_4108_n871_1), .Y(rdata_4__FF_INPUT) );
  AOI21X1 AOI21X1_4 ( .A(_abc_4108_n646_1), .B(_abc_4108_n601), .C(_abc_4108_n650_1), .Y(bus_cap_1__FF_INPUT) );
  AOI21X1 AOI21X1_40 ( .A(_abc_4108_n579_1), .B(_abc_4108_n873_1), .C(_abc_4108_n874), .Y(rdata_5__FF_INPUT) );
  AOI21X1 AOI21X1_41 ( .A(_abc_4108_n579_1), .B(_abc_4108_n876), .C(_abc_4108_n877_1), .Y(rdata_6__FF_INPUT) );
  AOI21X1 AOI21X1_42 ( .A(_abc_4108_n579_1), .B(_abc_4108_n879_1), .C(_abc_4108_n880), .Y(rdata_7__FF_INPUT) );
  AOI21X1 AOI21X1_43 ( .A(_abc_4108_n579_1), .B(_abc_4108_n882), .C(_abc_4108_n883_1), .Y(rdata_8__FF_INPUT) );
  AOI21X1 AOI21X1_44 ( .A(_abc_4108_n579_1), .B(_abc_4108_n885_1), .C(_abc_4108_n886), .Y(rdata_9__FF_INPUT) );
  AOI21X1 AOI21X1_45 ( .A(_abc_4108_n579_1), .B(_abc_4108_n888), .C(_abc_4108_n889_1), .Y(rdata_10__FF_INPUT) );
  AOI21X1 AOI21X1_46 ( .A(_abc_4108_n579_1), .B(_abc_4108_n891_1), .C(_abc_4108_n892_1), .Y(rdata_11__FF_INPUT) );
  AOI21X1 AOI21X1_47 ( .A(_abc_4108_n579_1), .B(_abc_4108_n894_1), .C(_abc_4108_n895_1), .Y(rdata_12__FF_INPUT) );
  AOI21X1 AOI21X1_48 ( .A(_abc_4108_n579_1), .B(_abc_4108_n897_1), .C(_abc_4108_n898_1), .Y(rdata_13__FF_INPUT) );
  AOI21X1 AOI21X1_49 ( .A(_abc_4108_n579_1), .B(_abc_4108_n900_1), .C(_abc_4108_n901_1), .Y(rdata_14__FF_INPUT) );
  AOI21X1 AOI21X1_5 ( .A(_abc_4108_n654_1), .B(_abc_4108_n601), .C(_abc_4108_n658_1), .Y(bus_cap_2__FF_INPUT) );
  AOI21X1 AOI21X1_50 ( .A(_abc_4108_n579_1), .B(_abc_4108_n903_1), .C(_abc_4108_n904_1), .Y(rdata_15__FF_INPUT) );
  AOI21X1 AOI21X1_51 ( .A(_abc_4108_n579_1), .B(_abc_4108_n906_1), .C(_abc_4108_n907_1), .Y(rdata_16__FF_INPUT) );
  AOI21X1 AOI21X1_52 ( .A(_abc_4108_n579_1), .B(_abc_4108_n909_1), .C(_abc_4108_n910_1), .Y(rdata_17__FF_INPUT) );
  AOI21X1 AOI21X1_53 ( .A(_abc_4108_n579_1), .B(_abc_4108_n912_1), .C(_abc_4108_n913_1), .Y(rdata_18__FF_INPUT) );
  AOI21X1 AOI21X1_54 ( .A(_abc_4108_n579_1), .B(_abc_4108_n915_1), .C(_abc_4108_n916_1), .Y(rdata_19__FF_INPUT) );
  AOI21X1 AOI21X1_55 ( .A(_abc_4108_n579_1), .B(_abc_4108_n918_1), .C(_abc_4108_n919_1), .Y(rdata_20__FF_INPUT) );
  AOI21X1 AOI21X1_56 ( .A(_abc_4108_n579_1), .B(_abc_4108_n921_1), .C(_abc_4108_n922_1), .Y(rdata_21__FF_INPUT) );
  AOI21X1 AOI21X1_57 ( .A(_abc_4108_n579_1), .B(_abc_4108_n924_1), .C(_abc_4108_n925_1), .Y(rdata_22__FF_INPUT) );
  AOI21X1 AOI21X1_58 ( .A(_abc_4108_n579_1), .B(_abc_4108_n927_1), .C(_abc_4108_n928_1), .Y(rdata_23__FF_INPUT) );
  AOI21X1 AOI21X1_59 ( .A(_abc_4108_n579_1), .B(_abc_4108_n930_1), .C(_abc_4108_n931_1), .Y(rdata_24__FF_INPUT) );
  AOI21X1 AOI21X1_6 ( .A(_abc_4108_n688), .B(_abc_4108_n660), .C(_abc_4108_n561), .Y(bus_cap_3__FF_INPUT) );
  AOI21X1 AOI21X1_60 ( .A(_abc_4108_n579_1), .B(_abc_4108_n933_1), .C(_abc_4108_n934_1), .Y(rdata_25__FF_INPUT) );
  AOI21X1 AOI21X1_61 ( .A(_abc_4108_n579_1), .B(_abc_4108_n936_1), .C(_abc_4108_n937_1), .Y(rdata_26__FF_INPUT) );
  AOI21X1 AOI21X1_62 ( .A(_abc_4108_n579_1), .B(_abc_4108_n939_1), .C(_abc_4108_n940_1), .Y(rdata_27__FF_INPUT) );
  AOI21X1 AOI21X1_63 ( .A(_abc_4108_n579_1), .B(_abc_4108_n942_1), .C(_abc_4108_n943_1), .Y(rdata_28__FF_INPUT) );
  AOI21X1 AOI21X1_64 ( .A(_abc_4108_n579_1), .B(_abc_4108_n945_1), .C(_abc_4108_n946_1), .Y(rdata_29__FF_INPUT) );
  AOI21X1 AOI21X1_65 ( .A(_abc_4108_n579_1), .B(_abc_4108_n948_1), .C(_abc_4108_n949_1), .Y(rdata_30__FF_INPUT) );
  AOI21X1 AOI21X1_66 ( .A(_abc_4108_n579_1), .B(_abc_4108_n951_1), .C(_abc_4108_n952), .Y(rdata_31__FF_INPUT) );
  AOI21X1 AOI21X1_67 ( .A(_abc_4108_n954), .B(_abc_4108_n956), .C(_abc_4108_n957), .Y(WDATA_0__FF_INPUT) );
  AOI21X1 AOI21X1_68 ( .A(_abc_4108_n959), .B(_abc_4108_n956), .C(_abc_4108_n960), .Y(WDATA_1__FF_INPUT) );
  AOI21X1 AOI21X1_69 ( .A(_abc_4108_n962), .B(_abc_4108_n956), .C(_abc_4108_n963_1), .Y(WDATA_2__FF_INPUT) );
  AOI21X1 AOI21X1_7 ( .A(_abc_4108_n694_1), .B(_abc_4108_n690_1), .C(_abc_4108_n561), .Y(bus_cap_4__FF_INPUT) );
  AOI21X1 AOI21X1_70 ( .A(_abc_4108_n965), .B(_abc_4108_n956), .C(_abc_4108_n966_1), .Y(WDATA_3__FF_INPUT) );
  AOI21X1 AOI21X1_71 ( .A(_abc_4108_n968_1), .B(_abc_4108_n956), .C(_abc_4108_n969_1), .Y(WDATA_4__FF_INPUT) );
  AOI21X1 AOI21X1_72 ( .A(_abc_4108_n971), .B(_abc_4108_n956), .C(_abc_4108_n972), .Y(WDATA_5__FF_INPUT) );
  AOI21X1 AOI21X1_73 ( .A(_abc_4108_n974), .B(_abc_4108_n956), .C(_abc_4108_n975), .Y(WDATA_6__FF_INPUT) );
  AOI21X1 AOI21X1_74 ( .A(_abc_4108_n977), .B(_abc_4108_n956), .C(_abc_4108_n978), .Y(WDATA_7__FF_INPUT) );
  AOI21X1 AOI21X1_75 ( .A(_abc_4108_n980), .B(_abc_4108_n956), .C(_abc_4108_n981), .Y(WDATA_8__FF_INPUT) );
  AOI21X1 AOI21X1_76 ( .A(_abc_4108_n983), .B(_abc_4108_n956), .C(_abc_4108_n984), .Y(WDATA_9__FF_INPUT) );
  AOI21X1 AOI21X1_77 ( .A(_abc_4108_n986), .B(_abc_4108_n956), .C(_abc_4108_n987), .Y(WDATA_10__FF_INPUT) );
  AOI21X1 AOI21X1_78 ( .A(_abc_4108_n989), .B(_abc_4108_n956), .C(_abc_4108_n990), .Y(WDATA_11__FF_INPUT) );
  AOI21X1 AOI21X1_79 ( .A(_abc_4108_n992), .B(_abc_4108_n956), .C(_abc_4108_n993), .Y(WDATA_12__FF_INPUT) );
  AOI21X1 AOI21X1_8 ( .A(_abc_4108_n700), .B(_abc_4108_n696), .C(_abc_4108_n561), .Y(bus_cap_5__FF_INPUT) );
  AOI21X1 AOI21X1_80 ( .A(_abc_4108_n995), .B(_abc_4108_n956), .C(_abc_4108_n996), .Y(WDATA_13__FF_INPUT) );
  AOI21X1 AOI21X1_81 ( .A(_abc_4108_n998), .B(_abc_4108_n956), .C(_abc_4108_n999), .Y(WDATA_14__FF_INPUT) );
  AOI21X1 AOI21X1_82 ( .A(_abc_4108_n1001), .B(_abc_4108_n956), .C(_abc_4108_n1002), .Y(WDATA_15__FF_INPUT) );
  AOI21X1 AOI21X1_83 ( .A(_abc_4108_n1004), .B(_abc_4108_n956), .C(_abc_4108_n1005), .Y(WDATA_16__FF_INPUT) );
  AOI21X1 AOI21X1_84 ( .A(_abc_4108_n1007), .B(_abc_4108_n956), .C(_abc_4108_n1008), .Y(WDATA_17__FF_INPUT) );
  AOI21X1 AOI21X1_85 ( .A(_abc_4108_n1010), .B(_abc_4108_n956), .C(_abc_4108_n1011), .Y(WDATA_18__FF_INPUT) );
  AOI21X1 AOI21X1_86 ( .A(_abc_4108_n1013), .B(_abc_4108_n956), .C(_abc_4108_n1014), .Y(WDATA_19__FF_INPUT) );
  AOI21X1 AOI21X1_87 ( .A(_abc_4108_n1016), .B(_abc_4108_n956), .C(_abc_4108_n1017), .Y(WDATA_20__FF_INPUT) );
  AOI21X1 AOI21X1_88 ( .A(_abc_4108_n1019), .B(_abc_4108_n956), .C(_abc_4108_n1020), .Y(WDATA_21__FF_INPUT) );
  AOI21X1 AOI21X1_89 ( .A(_abc_4108_n1022), .B(_abc_4108_n956), .C(_abc_4108_n1023), .Y(WDATA_22__FF_INPUT) );
  AOI21X1 AOI21X1_9 ( .A(_abc_4108_n706_1), .B(_abc_4108_n702_1), .C(_abc_4108_n561), .Y(bus_cap_6__FF_INPUT) );
  AOI21X1 AOI21X1_90 ( .A(_abc_4108_n1025), .B(_abc_4108_n956), .C(_abc_4108_n1026), .Y(WDATA_23__FF_INPUT) );
  AOI21X1 AOI21X1_91 ( .A(_abc_4108_n1028), .B(_abc_4108_n956), .C(_abc_4108_n1029), .Y(WDATA_24__FF_INPUT) );
  AOI21X1 AOI21X1_92 ( .A(_abc_4108_n1031), .B(_abc_4108_n956), .C(_abc_4108_n1032), .Y(WDATA_25__FF_INPUT) );
  AOI21X1 AOI21X1_93 ( .A(_abc_4108_n1034), .B(_abc_4108_n956), .C(_abc_4108_n1035), .Y(WDATA_26__FF_INPUT) );
  AOI21X1 AOI21X1_94 ( .A(_abc_4108_n1037), .B(_abc_4108_n956), .C(_abc_4108_n1038), .Y(WDATA_27__FF_INPUT) );
  AOI21X1 AOI21X1_95 ( .A(_abc_4108_n1040), .B(_abc_4108_n956), .C(_abc_4108_n1041), .Y(WDATA_28__FF_INPUT) );
  AOI21X1 AOI21X1_96 ( .A(_abc_4108_n1043), .B(_abc_4108_n956), .C(_abc_4108_n1044), .Y(WDATA_29__FF_INPUT) );
  AOI21X1 AOI21X1_97 ( .A(_abc_4108_n1046), .B(_abc_4108_n956), .C(_abc_4108_n1047), .Y(WDATA_30__FF_INPUT) );
  AOI21X1 AOI21X1_98 ( .A(_abc_4108_n1049), .B(_abc_4108_n956), .C(_abc_4108_n1050), .Y(WDATA_31__FF_INPUT) );
  AOI21X1 AOI21X1_99 ( .A(_abc_4108_n1149), .B(_abc_4108_n1055), .C(_abc_4108_n1150), .Y(A_ADDR_31__FF_INPUT) );
  AOI22X1 AOI22X1_1 ( .A(axi_awready), .B(state_5_), .C(state_3_), .D(_abc_4108_n562_1), .Y(_abc_4108_n563_1) );
  AOI22X1 AOI22X1_10 ( .A(_abc_4108_n1057), .B(_abc_4108_n1078), .C(_abc_4108_n1077), .D(_abc_4108_n1055), .Y(A_ADDR_7__FF_INPUT) );
  AOI22X1 AOI22X1_11 ( .A(_abc_4108_n1057), .B(_abc_4108_n1081), .C(_abc_4108_n1080), .D(_abc_4108_n1055), .Y(A_ADDR_8__FF_INPUT) );
  AOI22X1 AOI22X1_12 ( .A(_abc_4108_n1057), .B(_abc_4108_n1084), .C(_abc_4108_n1083), .D(_abc_4108_n1055), .Y(A_ADDR_9__FF_INPUT) );
  AOI22X1 AOI22X1_13 ( .A(_abc_4108_n1057), .B(_abc_4108_n1087), .C(_abc_4108_n1086), .D(_abc_4108_n1055), .Y(A_ADDR_10__FF_INPUT) );
  AOI22X1 AOI22X1_14 ( .A(_abc_4108_n1057), .B(_abc_4108_n1090), .C(_abc_4108_n1089), .D(_abc_4108_n1055), .Y(A_ADDR_11__FF_INPUT) );
  AOI22X1 AOI22X1_15 ( .A(_abc_4108_n1057), .B(_abc_4108_n1093), .C(_abc_4108_n1092), .D(_abc_4108_n1055), .Y(A_ADDR_12__FF_INPUT) );
  AOI22X1 AOI22X1_16 ( .A(_abc_4108_n1057), .B(_abc_4108_n1096), .C(_abc_4108_n1095), .D(_abc_4108_n1055), .Y(A_ADDR_13__FF_INPUT) );
  AOI22X1 AOI22X1_17 ( .A(_abc_4108_n1057), .B(_abc_4108_n1099), .C(_abc_4108_n1098), .D(_abc_4108_n1055), .Y(A_ADDR_14__FF_INPUT) );
  AOI22X1 AOI22X1_18 ( .A(_abc_4108_n1057), .B(_abc_4108_n1102), .C(_abc_4108_n1101), .D(_abc_4108_n1055), .Y(A_ADDR_15__FF_INPUT) );
  AOI22X1 AOI22X1_19 ( .A(_abc_4108_n1057), .B(_abc_4108_n1105), .C(_abc_4108_n1104), .D(_abc_4108_n1055), .Y(A_ADDR_16__FF_INPUT) );
  AOI22X1 AOI22X1_2 ( .A(_abc_4108_n575), .B(state_5_), .C(state_0_), .D(_abc_4108_n576), .Y(_abc_4108_n577_1) );
  AOI22X1 AOI22X1_20 ( .A(_abc_4108_n1057), .B(_abc_4108_n1108), .C(_abc_4108_n1107), .D(_abc_4108_n1055), .Y(A_ADDR_17__FF_INPUT) );
  AOI22X1 AOI22X1_21 ( .A(_abc_4108_n1057), .B(_abc_4108_n1111), .C(_abc_4108_n1110), .D(_abc_4108_n1055), .Y(A_ADDR_18__FF_INPUT) );
  AOI22X1 AOI22X1_22 ( .A(_abc_4108_n1057), .B(_abc_4108_n1114), .C(_abc_4108_n1113), .D(_abc_4108_n1055), .Y(A_ADDR_19__FF_INPUT) );
  AOI22X1 AOI22X1_23 ( .A(_abc_4108_n1057), .B(_abc_4108_n1117), .C(_abc_4108_n1116), .D(_abc_4108_n1055), .Y(A_ADDR_20__FF_INPUT) );
  AOI22X1 AOI22X1_24 ( .A(_abc_4108_n1057), .B(_abc_4108_n1120), .C(_abc_4108_n1119), .D(_abc_4108_n1055), .Y(A_ADDR_21__FF_INPUT) );
  AOI22X1 AOI22X1_25 ( .A(_abc_4108_n1057), .B(_abc_4108_n1123), .C(_abc_4108_n1122), .D(_abc_4108_n1055), .Y(A_ADDR_22__FF_INPUT) );
  AOI22X1 AOI22X1_26 ( .A(_abc_4108_n1057), .B(_abc_4108_n1126), .C(_abc_4108_n1125), .D(_abc_4108_n1055), .Y(A_ADDR_23__FF_INPUT) );
  AOI22X1 AOI22X1_27 ( .A(_abc_4108_n1057), .B(_abc_4108_n1129), .C(_abc_4108_n1128), .D(_abc_4108_n1055), .Y(A_ADDR_24__FF_INPUT) );
  AOI22X1 AOI22X1_28 ( .A(_abc_4108_n1057), .B(_abc_4108_n1132), .C(_abc_4108_n1131), .D(_abc_4108_n1055), .Y(A_ADDR_25__FF_INPUT) );
  AOI22X1 AOI22X1_29 ( .A(_abc_4108_n1057), .B(_abc_4108_n1135), .C(_abc_4108_n1134), .D(_abc_4108_n1055), .Y(A_ADDR_26__FF_INPUT) );
  AOI22X1 AOI22X1_3 ( .A(_abc_4108_n1056), .B(_abc_4108_n1057), .C(_abc_4108_n1052), .D(_abc_4108_n1055), .Y(A_ADDR_0__FF_INPUT) );
  AOI22X1 AOI22X1_30 ( .A(_abc_4108_n1057), .B(_abc_4108_n1138), .C(_abc_4108_n1137), .D(_abc_4108_n1055), .Y(A_ADDR_27__FF_INPUT) );
  AOI22X1 AOI22X1_31 ( .A(_abc_4108_n1057), .B(_abc_4108_n1141), .C(_abc_4108_n1140), .D(_abc_4108_n1055), .Y(A_ADDR_28__FF_INPUT) );
  AOI22X1 AOI22X1_32 ( .A(_abc_4108_n1057), .B(_abc_4108_n1144), .C(_abc_4108_n1143), .D(_abc_4108_n1055), .Y(A_ADDR_29__FF_INPUT) );
  AOI22X1 AOI22X1_33 ( .A(_abc_4108_n1057), .B(_abc_4108_n1147), .C(_abc_4108_n1146), .D(_abc_4108_n1055), .Y(A_ADDR_30__FF_INPUT) );
  AOI22X1 AOI22X1_4 ( .A(_abc_4108_n1057), .B(_abc_4108_n1060), .C(_abc_4108_n1059), .D(_abc_4108_n1055), .Y(A_ADDR_1__FF_INPUT) );
  AOI22X1 AOI22X1_5 ( .A(_abc_4108_n1057), .B(_abc_4108_n1063), .C(_abc_4108_n1062), .D(_abc_4108_n1055), .Y(A_ADDR_2__FF_INPUT) );
  AOI22X1 AOI22X1_6 ( .A(_abc_4108_n1057), .B(_abc_4108_n1066), .C(_abc_4108_n1065), .D(_abc_4108_n1055), .Y(A_ADDR_3__FF_INPUT) );
  AOI22X1 AOI22X1_7 ( .A(_abc_4108_n1057), .B(_abc_4108_n1069), .C(_abc_4108_n1068), .D(_abc_4108_n1055), .Y(A_ADDR_4__FF_INPUT) );
  AOI22X1 AOI22X1_8 ( .A(_abc_4108_n1057), .B(_abc_4108_n1072), .C(_abc_4108_n1071), .D(_abc_4108_n1055), .Y(A_ADDR_5__FF_INPUT) );
  AOI22X1 AOI22X1_9 ( .A(_abc_4108_n1057), .B(_abc_4108_n1075), .C(_abc_4108_n1074), .D(_abc_4108_n1055), .Y(A_ADDR_6__FF_INPUT) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(SCLK), .D(counter_0__FF_INPUT), .Q(counter_0_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(SCLK), .D(counter_9__FF_INPUT), .Q(counter_9_) );
  DFFPOSX1 DFFPOSX1_100 ( .CLK(CLK), .D(rdata_0__FF_INPUT), .Q(bus_sync_rdata_data_in_0_) );
  DFFPOSX1 DFFPOSX1_101 ( .CLK(CLK), .D(rdata_1__FF_INPUT), .Q(bus_sync_rdata_data_in_1_) );
  DFFPOSX1 DFFPOSX1_102 ( .CLK(CLK), .D(rdata_2__FF_INPUT), .Q(bus_sync_rdata_data_in_2_) );
  DFFPOSX1 DFFPOSX1_103 ( .CLK(CLK), .D(rdata_3__FF_INPUT), .Q(bus_sync_rdata_data_in_3_) );
  DFFPOSX1 DFFPOSX1_104 ( .CLK(CLK), .D(rdata_4__FF_INPUT), .Q(bus_sync_rdata_data_in_4_) );
  DFFPOSX1 DFFPOSX1_105 ( .CLK(CLK), .D(rdata_5__FF_INPUT), .Q(bus_sync_rdata_data_in_5_) );
  DFFPOSX1 DFFPOSX1_106 ( .CLK(CLK), .D(rdata_6__FF_INPUT), .Q(bus_sync_rdata_data_in_6_) );
  DFFPOSX1 DFFPOSX1_107 ( .CLK(CLK), .D(rdata_7__FF_INPUT), .Q(bus_sync_rdata_data_in_7_) );
  DFFPOSX1 DFFPOSX1_108 ( .CLK(CLK), .D(rdata_8__FF_INPUT), .Q(bus_sync_rdata_data_in_8_) );
  DFFPOSX1 DFFPOSX1_109 ( .CLK(CLK), .D(rdata_9__FF_INPUT), .Q(bus_sync_rdata_data_in_9_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(SCLK), .D(counter_10__FF_INPUT), .Q(counter_10_) );
  DFFPOSX1 DFFPOSX1_110 ( .CLK(CLK), .D(rdata_10__FF_INPUT), .Q(bus_sync_rdata_data_in_10_) );
  DFFPOSX1 DFFPOSX1_111 ( .CLK(CLK), .D(rdata_11__FF_INPUT), .Q(bus_sync_rdata_data_in_11_) );
  DFFPOSX1 DFFPOSX1_112 ( .CLK(CLK), .D(rdata_12__FF_INPUT), .Q(bus_sync_rdata_data_in_12_) );
  DFFPOSX1 DFFPOSX1_113 ( .CLK(CLK), .D(rdata_13__FF_INPUT), .Q(bus_sync_rdata_data_in_13_) );
  DFFPOSX1 DFFPOSX1_114 ( .CLK(CLK), .D(rdata_14__FF_INPUT), .Q(bus_sync_rdata_data_in_14_) );
  DFFPOSX1 DFFPOSX1_115 ( .CLK(CLK), .D(rdata_15__FF_INPUT), .Q(bus_sync_rdata_data_in_15_) );
  DFFPOSX1 DFFPOSX1_116 ( .CLK(CLK), .D(rdata_16__FF_INPUT), .Q(bus_sync_rdata_data_in_16_) );
  DFFPOSX1 DFFPOSX1_117 ( .CLK(CLK), .D(rdata_17__FF_INPUT), .Q(bus_sync_rdata_data_in_17_) );
  DFFPOSX1 DFFPOSX1_118 ( .CLK(CLK), .D(rdata_18__FF_INPUT), .Q(bus_sync_rdata_data_in_18_) );
  DFFPOSX1 DFFPOSX1_119 ( .CLK(CLK), .D(rdata_19__FF_INPUT), .Q(bus_sync_rdata_data_in_19_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(SCLK), .D(counter_11__FF_INPUT), .Q(counter_11_) );
  DFFPOSX1 DFFPOSX1_120 ( .CLK(CLK), .D(rdata_20__FF_INPUT), .Q(bus_sync_rdata_data_in_20_) );
  DFFPOSX1 DFFPOSX1_121 ( .CLK(CLK), .D(rdata_21__FF_INPUT), .Q(bus_sync_rdata_data_in_21_) );
  DFFPOSX1 DFFPOSX1_122 ( .CLK(CLK), .D(rdata_22__FF_INPUT), .Q(bus_sync_rdata_data_in_22_) );
  DFFPOSX1 DFFPOSX1_123 ( .CLK(CLK), .D(rdata_23__FF_INPUT), .Q(bus_sync_rdata_data_in_23_) );
  DFFPOSX1 DFFPOSX1_124 ( .CLK(CLK), .D(rdata_24__FF_INPUT), .Q(bus_sync_rdata_data_in_24_) );
  DFFPOSX1 DFFPOSX1_125 ( .CLK(CLK), .D(rdata_25__FF_INPUT), .Q(bus_sync_rdata_data_in_25_) );
  DFFPOSX1 DFFPOSX1_126 ( .CLK(CLK), .D(rdata_26__FF_INPUT), .Q(bus_sync_rdata_data_in_26_) );
  DFFPOSX1 DFFPOSX1_127 ( .CLK(CLK), .D(rdata_27__FF_INPUT), .Q(bus_sync_rdata_data_in_27_) );
  DFFPOSX1 DFFPOSX1_128 ( .CLK(CLK), .D(rdata_28__FF_INPUT), .Q(bus_sync_rdata_data_in_28_) );
  DFFPOSX1 DFFPOSX1_129 ( .CLK(CLK), .D(rdata_29__FF_INPUT), .Q(bus_sync_rdata_data_in_29_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(SCLK), .D(counter_12__FF_INPUT), .Q(counter_12_) );
  DFFPOSX1 DFFPOSX1_130 ( .CLK(CLK), .D(rdata_30__FF_INPUT), .Q(bus_sync_rdata_data_in_30_) );
  DFFPOSX1 DFFPOSX1_131 ( .CLK(CLK), .D(rdata_31__FF_INPUT), .Q(bus_sync_rdata_data_in_31_) );
  DFFPOSX1 DFFPOSX1_132 ( .CLK(SCLK), .D(A_ADDR_0__FF_INPUT), .Q(A_ADDR_0_) );
  DFFPOSX1 DFFPOSX1_133 ( .CLK(SCLK), .D(A_ADDR_1__FF_INPUT), .Q(A_ADDR_1_) );
  DFFPOSX1 DFFPOSX1_134 ( .CLK(SCLK), .D(A_ADDR_2__FF_INPUT), .Q(A_ADDR_2_) );
  DFFPOSX1 DFFPOSX1_135 ( .CLK(SCLK), .D(A_ADDR_3__FF_INPUT), .Q(A_ADDR_3_) );
  DFFPOSX1 DFFPOSX1_136 ( .CLK(SCLK), .D(A_ADDR_4__FF_INPUT), .Q(A_ADDR_4_) );
  DFFPOSX1 DFFPOSX1_137 ( .CLK(SCLK), .D(A_ADDR_5__FF_INPUT), .Q(A_ADDR_5_) );
  DFFPOSX1 DFFPOSX1_138 ( .CLK(SCLK), .D(A_ADDR_6__FF_INPUT), .Q(A_ADDR_6_) );
  DFFPOSX1 DFFPOSX1_139 ( .CLK(SCLK), .D(A_ADDR_7__FF_INPUT), .Q(A_ADDR_7_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(SCLK), .D(counter_13__FF_INPUT), .Q(counter_13_) );
  DFFPOSX1 DFFPOSX1_140 ( .CLK(SCLK), .D(A_ADDR_8__FF_INPUT), .Q(A_ADDR_8_) );
  DFFPOSX1 DFFPOSX1_141 ( .CLK(SCLK), .D(A_ADDR_9__FF_INPUT), .Q(A_ADDR_9_) );
  DFFPOSX1 DFFPOSX1_142 ( .CLK(SCLK), .D(A_ADDR_10__FF_INPUT), .Q(A_ADDR_10_) );
  DFFPOSX1 DFFPOSX1_143 ( .CLK(SCLK), .D(A_ADDR_11__FF_INPUT), .Q(A_ADDR_11_) );
  DFFPOSX1 DFFPOSX1_144 ( .CLK(SCLK), .D(A_ADDR_12__FF_INPUT), .Q(A_ADDR_12_) );
  DFFPOSX1 DFFPOSX1_145 ( .CLK(SCLK), .D(A_ADDR_13__FF_INPUT), .Q(A_ADDR_13_) );
  DFFPOSX1 DFFPOSX1_146 ( .CLK(SCLK), .D(A_ADDR_14__FF_INPUT), .Q(A_ADDR_14_) );
  DFFPOSX1 DFFPOSX1_147 ( .CLK(SCLK), .D(A_ADDR_15__FF_INPUT), .Q(A_ADDR_15_) );
  DFFPOSX1 DFFPOSX1_148 ( .CLK(SCLK), .D(A_ADDR_16__FF_INPUT), .Q(A_ADDR_16_) );
  DFFPOSX1 DFFPOSX1_149 ( .CLK(SCLK), .D(A_ADDR_17__FF_INPUT), .Q(A_ADDR_17_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(SCLK), .D(counter_14__FF_INPUT), .Q(counter_14_) );
  DFFPOSX1 DFFPOSX1_150 ( .CLK(SCLK), .D(A_ADDR_18__FF_INPUT), .Q(A_ADDR_18_) );
  DFFPOSX1 DFFPOSX1_151 ( .CLK(SCLK), .D(A_ADDR_19__FF_INPUT), .Q(A_ADDR_19_) );
  DFFPOSX1 DFFPOSX1_152 ( .CLK(SCLK), .D(A_ADDR_20__FF_INPUT), .Q(A_ADDR_20_) );
  DFFPOSX1 DFFPOSX1_153 ( .CLK(SCLK), .D(A_ADDR_21__FF_INPUT), .Q(A_ADDR_21_) );
  DFFPOSX1 DFFPOSX1_154 ( .CLK(SCLK), .D(A_ADDR_22__FF_INPUT), .Q(A_ADDR_22_) );
  DFFPOSX1 DFFPOSX1_155 ( .CLK(SCLK), .D(A_ADDR_23__FF_INPUT), .Q(A_ADDR_23_) );
  DFFPOSX1 DFFPOSX1_156 ( .CLK(SCLK), .D(A_ADDR_24__FF_INPUT), .Q(A_ADDR_24_) );
  DFFPOSX1 DFFPOSX1_157 ( .CLK(SCLK), .D(A_ADDR_25__FF_INPUT), .Q(A_ADDR_25_) );
  DFFPOSX1 DFFPOSX1_158 ( .CLK(SCLK), .D(A_ADDR_26__FF_INPUT), .Q(A_ADDR_26_) );
  DFFPOSX1 DFFPOSX1_159 ( .CLK(SCLK), .D(A_ADDR_27__FF_INPUT), .Q(A_ADDR_27_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(SCLK), .D(counter_15__FF_INPUT), .Q(counter_15_) );
  DFFPOSX1 DFFPOSX1_160 ( .CLK(SCLK), .D(A_ADDR_28__FF_INPUT), .Q(A_ADDR_28_) );
  DFFPOSX1 DFFPOSX1_161 ( .CLK(SCLK), .D(A_ADDR_29__FF_INPUT), .Q(A_ADDR_29_) );
  DFFPOSX1 DFFPOSX1_162 ( .CLK(SCLK), .D(A_ADDR_30__FF_INPUT), .Q(A_ADDR_30_) );
  DFFPOSX1 DFFPOSX1_163 ( .CLK(SCLK), .D(A_ADDR_31__FF_INPUT), .Q(A_ADDR_31_) );
  DFFPOSX1 DFFPOSX1_164 ( .CLK(SCLK), .D(WDATA_0__FF_INPUT), .Q(WDATA_0_) );
  DFFPOSX1 DFFPOSX1_165 ( .CLK(SCLK), .D(WDATA_1__FF_INPUT), .Q(WDATA_1_) );
  DFFPOSX1 DFFPOSX1_166 ( .CLK(SCLK), .D(WDATA_2__FF_INPUT), .Q(WDATA_2_) );
  DFFPOSX1 DFFPOSX1_167 ( .CLK(SCLK), .D(WDATA_3__FF_INPUT), .Q(WDATA_3_) );
  DFFPOSX1 DFFPOSX1_168 ( .CLK(SCLK), .D(WDATA_4__FF_INPUT), .Q(WDATA_4_) );
  DFFPOSX1 DFFPOSX1_169 ( .CLK(SCLK), .D(WDATA_5__FF_INPUT), .Q(WDATA_5_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(SCLK), .D(counter_16__FF_INPUT), .Q(counter_16_) );
  DFFPOSX1 DFFPOSX1_170 ( .CLK(SCLK), .D(WDATA_6__FF_INPUT), .Q(WDATA_6_) );
  DFFPOSX1 DFFPOSX1_171 ( .CLK(SCLK), .D(WDATA_7__FF_INPUT), .Q(WDATA_7_) );
  DFFPOSX1 DFFPOSX1_172 ( .CLK(SCLK), .D(WDATA_8__FF_INPUT), .Q(WDATA_8_) );
  DFFPOSX1 DFFPOSX1_173 ( .CLK(SCLK), .D(WDATA_9__FF_INPUT), .Q(WDATA_9_) );
  DFFPOSX1 DFFPOSX1_174 ( .CLK(SCLK), .D(WDATA_10__FF_INPUT), .Q(WDATA_10_) );
  DFFPOSX1 DFFPOSX1_175 ( .CLK(SCLK), .D(WDATA_11__FF_INPUT), .Q(WDATA_11_) );
  DFFPOSX1 DFFPOSX1_176 ( .CLK(SCLK), .D(WDATA_12__FF_INPUT), .Q(WDATA_12_) );
  DFFPOSX1 DFFPOSX1_177 ( .CLK(SCLK), .D(WDATA_13__FF_INPUT), .Q(WDATA_13_) );
  DFFPOSX1 DFFPOSX1_178 ( .CLK(SCLK), .D(WDATA_14__FF_INPUT), .Q(WDATA_14_) );
  DFFPOSX1 DFFPOSX1_179 ( .CLK(SCLK), .D(WDATA_15__FF_INPUT), .Q(WDATA_15_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(SCLK), .D(counter_17__FF_INPUT), .Q(counter_17_) );
  DFFPOSX1 DFFPOSX1_180 ( .CLK(SCLK), .D(WDATA_16__FF_INPUT), .Q(WDATA_16_) );
  DFFPOSX1 DFFPOSX1_181 ( .CLK(SCLK), .D(WDATA_17__FF_INPUT), .Q(WDATA_17_) );
  DFFPOSX1 DFFPOSX1_182 ( .CLK(SCLK), .D(WDATA_18__FF_INPUT), .Q(WDATA_18_) );
  DFFPOSX1 DFFPOSX1_183 ( .CLK(SCLK), .D(WDATA_19__FF_INPUT), .Q(WDATA_19_) );
  DFFPOSX1 DFFPOSX1_184 ( .CLK(SCLK), .D(WDATA_20__FF_INPUT), .Q(WDATA_20_) );
  DFFPOSX1 DFFPOSX1_185 ( .CLK(SCLK), .D(WDATA_21__FF_INPUT), .Q(WDATA_21_) );
  DFFPOSX1 DFFPOSX1_186 ( .CLK(SCLK), .D(WDATA_22__FF_INPUT), .Q(WDATA_22_) );
  DFFPOSX1 DFFPOSX1_187 ( .CLK(SCLK), .D(WDATA_23__FF_INPUT), .Q(WDATA_23_) );
  DFFPOSX1 DFFPOSX1_188 ( .CLK(SCLK), .D(WDATA_24__FF_INPUT), .Q(WDATA_24_) );
  DFFPOSX1 DFFPOSX1_189 ( .CLK(SCLK), .D(WDATA_25__FF_INPUT), .Q(WDATA_25_) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(SCLK), .D(counter_18__FF_INPUT), .Q(counter_18_) );
  DFFPOSX1 DFFPOSX1_190 ( .CLK(SCLK), .D(WDATA_26__FF_INPUT), .Q(WDATA_26_) );
  DFFPOSX1 DFFPOSX1_191 ( .CLK(SCLK), .D(WDATA_27__FF_INPUT), .Q(WDATA_27_) );
  DFFPOSX1 DFFPOSX1_192 ( .CLK(SCLK), .D(WDATA_28__FF_INPUT), .Q(WDATA_28_) );
  DFFPOSX1 DFFPOSX1_193 ( .CLK(SCLK), .D(WDATA_29__FF_INPUT), .Q(WDATA_29_) );
  DFFPOSX1 DFFPOSX1_194 ( .CLK(SCLK), .D(WDATA_30__FF_INPUT), .Q(WDATA_30_) );
  DFFPOSX1 DFFPOSX1_195 ( .CLK(SCLK), .D(WDATA_31__FF_INPUT), .Q(WDATA_31_) );
  DFFPOSX1 DFFPOSX1_196 ( .CLK(SCLK), .D(PICORV_RST_SPI_FF_INPUT), .Q(PICORV_RST_SPI) );
  DFFPOSX1 DFFPOSX1_197 ( .CLK(SCLK), .D(we_FF_INPUT), .Q(we) );
  DFFPOSX1 DFFPOSX1_198 ( .CLK(SCLK), .D(re_FF_INPUT), .Q(re) );
  DFFPOSX1 DFFPOSX1_199 ( .CLK(SCLK), .D(sft_reg_0__FF_INPUT), .Q(sft_reg_0_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(SCLK), .D(counter_1__FF_INPUT), .Q(counter_1_) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(SCLK), .D(counter_19__FF_INPUT), .Q(counter_19_) );
  DFFPOSX1 DFFPOSX1_200 ( .CLK(SCLK), .D(sft_reg_1__FF_INPUT), .Q(sft_reg_1_) );
  DFFPOSX1 DFFPOSX1_201 ( .CLK(SCLK), .D(sft_reg_2__FF_INPUT), .Q(sft_reg_2_) );
  DFFPOSX1 DFFPOSX1_202 ( .CLK(SCLK), .D(sft_reg_3__FF_INPUT), .Q(sft_reg_3_) );
  DFFPOSX1 DFFPOSX1_203 ( .CLK(SCLK), .D(sft_reg_4__FF_INPUT), .Q(sft_reg_4_) );
  DFFPOSX1 DFFPOSX1_204 ( .CLK(SCLK), .D(sft_reg_5__FF_INPUT), .Q(sft_reg_5_) );
  DFFPOSX1 DFFPOSX1_205 ( .CLK(SCLK), .D(sft_reg_6__FF_INPUT), .Q(sft_reg_6_) );
  DFFPOSX1 DFFPOSX1_206 ( .CLK(SCLK), .D(sft_reg_7__FF_INPUT), .Q(sft_reg_7_) );
  DFFPOSX1 DFFPOSX1_207 ( .CLK(SCLK), .D(sft_reg_8__FF_INPUT), .Q(sft_reg_8_) );
  DFFPOSX1 DFFPOSX1_208 ( .CLK(SCLK), .D(sft_reg_9__FF_INPUT), .Q(sft_reg_9_) );
  DFFPOSX1 DFFPOSX1_209 ( .CLK(SCLK), .D(sft_reg_10__FF_INPUT), .Q(sft_reg_10_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(SCLK), .D(counter_20__FF_INPUT), .Q(counter_20_) );
  DFFPOSX1 DFFPOSX1_210 ( .CLK(SCLK), .D(sft_reg_11__FF_INPUT), .Q(sft_reg_11_) );
  DFFPOSX1 DFFPOSX1_211 ( .CLK(SCLK), .D(sft_reg_12__FF_INPUT), .Q(sft_reg_12_) );
  DFFPOSX1 DFFPOSX1_212 ( .CLK(SCLK), .D(sft_reg_13__FF_INPUT), .Q(sft_reg_13_) );
  DFFPOSX1 DFFPOSX1_213 ( .CLK(SCLK), .D(sft_reg_14__FF_INPUT), .Q(sft_reg_14_) );
  DFFPOSX1 DFFPOSX1_214 ( .CLK(SCLK), .D(sft_reg_15__FF_INPUT), .Q(sft_reg_15_) );
  DFFPOSX1 DFFPOSX1_215 ( .CLK(SCLK), .D(sft_reg_16__FF_INPUT), .Q(sft_reg_16_) );
  DFFPOSX1 DFFPOSX1_216 ( .CLK(SCLK), .D(sft_reg_17__FF_INPUT), .Q(sft_reg_17_) );
  DFFPOSX1 DFFPOSX1_217 ( .CLK(SCLK), .D(sft_reg_18__FF_INPUT), .Q(sft_reg_18_) );
  DFFPOSX1 DFFPOSX1_218 ( .CLK(SCLK), .D(sft_reg_19__FF_INPUT), .Q(sft_reg_19_) );
  DFFPOSX1 DFFPOSX1_219 ( .CLK(SCLK), .D(sft_reg_20__FF_INPUT), .Q(sft_reg_20_) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(SCLK), .D(counter_21__FF_INPUT), .Q(counter_21_) );
  DFFPOSX1 DFFPOSX1_220 ( .CLK(SCLK), .D(sft_reg_21__FF_INPUT), .Q(sft_reg_21_) );
  DFFPOSX1 DFFPOSX1_221 ( .CLK(SCLK), .D(sft_reg_22__FF_INPUT), .Q(sft_reg_22_) );
  DFFPOSX1 DFFPOSX1_222 ( .CLK(SCLK), .D(sft_reg_23__FF_INPUT), .Q(sft_reg_23_) );
  DFFPOSX1 DFFPOSX1_223 ( .CLK(SCLK), .D(sft_reg_24__FF_INPUT), .Q(sft_reg_24_) );
  DFFPOSX1 DFFPOSX1_224 ( .CLK(SCLK), .D(sft_reg_25__FF_INPUT), .Q(sft_reg_25_) );
  DFFPOSX1 DFFPOSX1_225 ( .CLK(SCLK), .D(sft_reg_26__FF_INPUT), .Q(sft_reg_26_) );
  DFFPOSX1 DFFPOSX1_226 ( .CLK(SCLK), .D(sft_reg_27__FF_INPUT), .Q(sft_reg_27_) );
  DFFPOSX1 DFFPOSX1_227 ( .CLK(SCLK), .D(sft_reg_28__FF_INPUT), .Q(sft_reg_28_) );
  DFFPOSX1 DFFPOSX1_228 ( .CLK(SCLK), .D(sft_reg_29__FF_INPUT), .Q(sft_reg_29_) );
  DFFPOSX1 DFFPOSX1_229 ( .CLK(SCLK), .D(sft_reg_30__FF_INPUT), .Q(sft_reg_30_) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(SCLK), .D(counter_22__FF_INPUT), .Q(counter_22_) );
  DFFPOSX1 DFFPOSX1_230 ( .CLK(CLK), .D(_abc_2913_n116), .Q(state_0_) );
  DFFPOSX1 DFFPOSX1_231 ( .CLK(CLK), .D(_abc_2913_n87), .Q(state_1_) );
  DFFPOSX1 DFFPOSX1_232 ( .CLK(CLK), .D(_abc_2913_n1036), .Q(axi_bready) );
  DFFPOSX1 DFFPOSX1_233 ( .CLK(CLK), .D(_abc_2913_n78), .Q(state_3_) );
  DFFPOSX1 DFFPOSX1_234 ( .CLK(CLK), .D(_abc_2913_n129), .Q(state_4_) );
  DFFPOSX1 DFFPOSX1_235 ( .CLK(CLK), .D(_abc_2913_n105), .Q(state_5_) );
  DFFPOSX1 DFFPOSX1_236 ( .CLK(CLK), .D(_abc_2913_n95), .Q(state_6_) );
  DFFPOSX1 DFFPOSX1_237 ( .CLK(CLK), .D(_abc_2913_n70), .Q(state_7_) );
  DFFPOSX1 DFFPOSX1_238 ( .CLK(CLK), .D(_abc_2913_n1025), .Q(axi_rready) );
  DFFPOSX1 DFFPOSX1_239 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_0__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_0_) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(SCLK), .D(counter_23__FF_INPUT), .Q(counter_23_) );
  DFFPOSX1 DFFPOSX1_240 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_1__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_1_) );
  DFFPOSX1 DFFPOSX1_241 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_2__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_2_) );
  DFFPOSX1 DFFPOSX1_242 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_3__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_3_) );
  DFFPOSX1 DFFPOSX1_243 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_4__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_4_) );
  DFFPOSX1 DFFPOSX1_244 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_5__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_5_) );
  DFFPOSX1 DFFPOSX1_245 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_6__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_6_) );
  DFFPOSX1 DFFPOSX1_246 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_7__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_7_) );
  DFFPOSX1 DFFPOSX1_247 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_8__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_8_) );
  DFFPOSX1 DFFPOSX1_248 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_9__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_9_) );
  DFFPOSX1 DFFPOSX1_249 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_10__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_10_) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(SCLK), .D(counter_24__FF_INPUT), .Q(counter_24_) );
  DFFPOSX1 DFFPOSX1_250 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_11__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_11_) );
  DFFPOSX1 DFFPOSX1_251 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_12__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_12_) );
  DFFPOSX1 DFFPOSX1_252 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_13__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_13_) );
  DFFPOSX1 DFFPOSX1_253 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_14__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_14_) );
  DFFPOSX1 DFFPOSX1_254 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_15__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_15_) );
  DFFPOSX1 DFFPOSX1_255 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_16__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_16_) );
  DFFPOSX1 DFFPOSX1_256 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_17__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_17_) );
  DFFPOSX1 DFFPOSX1_257 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_18__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_18_) );
  DFFPOSX1 DFFPOSX1_258 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_19__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_19_) );
  DFFPOSX1 DFFPOSX1_259 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_20__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_20_) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(SCLK), .D(counter_25__FF_INPUT), .Q(counter_25_) );
  DFFPOSX1 DFFPOSX1_260 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_21__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_21_) );
  DFFPOSX1 DFFPOSX1_261 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_22__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_22_) );
  DFFPOSX1 DFFPOSX1_262 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_23__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_23_) );
  DFFPOSX1 DFFPOSX1_263 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_24__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_24_) );
  DFFPOSX1 DFFPOSX1_264 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_25__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_25_) );
  DFFPOSX1 DFFPOSX1_265 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_26__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_26_) );
  DFFPOSX1 DFFPOSX1_266 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_27__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_27_) );
  DFFPOSX1 DFFPOSX1_267 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_28__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_28_) );
  DFFPOSX1 DFFPOSX1_268 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_29__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_29_) );
  DFFPOSX1 DFFPOSX1_269 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_30__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_30_) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(SCLK), .D(counter_26__FF_INPUT), .Q(counter_26_) );
  DFFPOSX1 DFFPOSX1_270 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_31__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_31_) );
  DFFPOSX1 DFFPOSX1_271 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_32__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_32_) );
  DFFPOSX1 DFFPOSX1_272 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_33__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_33_) );
  DFFPOSX1 DFFPOSX1_273 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_34__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_34_) );
  DFFPOSX1 DFFPOSX1_274 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_35__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_35_) );
  DFFPOSX1 DFFPOSX1_275 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_36__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_36_) );
  DFFPOSX1 DFFPOSX1_276 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_37__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_37_) );
  DFFPOSX1 DFFPOSX1_277 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_38__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_38_) );
  DFFPOSX1 DFFPOSX1_278 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_39__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_39_) );
  DFFPOSX1 DFFPOSX1_279 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_40__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_40_) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(SCLK), .D(counter_27__FF_INPUT), .Q(counter_27_) );
  DFFPOSX1 DFFPOSX1_280 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_41__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_41_) );
  DFFPOSX1 DFFPOSX1_281 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_42__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_42_) );
  DFFPOSX1 DFFPOSX1_282 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_43__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_43_) );
  DFFPOSX1 DFFPOSX1_283 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_44__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_44_) );
  DFFPOSX1 DFFPOSX1_284 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_45__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_45_) );
  DFFPOSX1 DFFPOSX1_285 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_46__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_46_) );
  DFFPOSX1 DFFPOSX1_286 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_47__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_47_) );
  DFFPOSX1 DFFPOSX1_287 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_48__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_48_) );
  DFFPOSX1 DFFPOSX1_288 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_49__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_49_) );
  DFFPOSX1 DFFPOSX1_289 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_50__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_50_) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(SCLK), .D(counter_28__FF_INPUT), .Q(counter_28_) );
  DFFPOSX1 DFFPOSX1_290 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_51__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_51_) );
  DFFPOSX1 DFFPOSX1_291 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_52__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_52_) );
  DFFPOSX1 DFFPOSX1_292 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_53__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_53_) );
  DFFPOSX1 DFFPOSX1_293 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_54__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_54_) );
  DFFPOSX1 DFFPOSX1_294 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_55__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_55_) );
  DFFPOSX1 DFFPOSX1_295 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_56__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_56_) );
  DFFPOSX1 DFFPOSX1_296 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_57__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_57_) );
  DFFPOSX1 DFFPOSX1_297 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_58__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_58_) );
  DFFPOSX1 DFFPOSX1_298 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_59__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_59_) );
  DFFPOSX1 DFFPOSX1_299 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_60__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_60_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(SCLK), .D(counter_2__FF_INPUT), .Q(counter_2_) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(SCLK), .D(counter_29__FF_INPUT), .Q(counter_29_) );
  DFFPOSX1 DFFPOSX1_300 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_61__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_61_) );
  DFFPOSX1 DFFPOSX1_301 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_62__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_62_) );
  DFFPOSX1 DFFPOSX1_302 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data2_63__FF_INPUT), .Q(bus_sync_axi_bus_reg_data2_63_) );
  DFFPOSX1 DFFPOSX1_303 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_0__FF_INPUT), .Q(\axi_wdata[0] ) );
  DFFPOSX1 DFFPOSX1_304 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_1__FF_INPUT), .Q(\axi_wdata[1] ) );
  DFFPOSX1 DFFPOSX1_305 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_2__FF_INPUT), .Q(\axi_wdata[2] ) );
  DFFPOSX1 DFFPOSX1_306 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_3__FF_INPUT), .Q(\axi_wdata[3] ) );
  DFFPOSX1 DFFPOSX1_307 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_4__FF_INPUT), .Q(\axi_wdata[4] ) );
  DFFPOSX1 DFFPOSX1_308 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_5__FF_INPUT), .Q(\axi_wdata[5] ) );
  DFFPOSX1 DFFPOSX1_309 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_6__FF_INPUT), .Q(\axi_wdata[6] ) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(SCLK), .D(counter_30__FF_INPUT), .Q(counter_30_) );
  DFFPOSX1 DFFPOSX1_310 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_7__FF_INPUT), .Q(\axi_wdata[7] ) );
  DFFPOSX1 DFFPOSX1_311 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_8__FF_INPUT), .Q(\axi_wdata[8] ) );
  DFFPOSX1 DFFPOSX1_312 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_9__FF_INPUT), .Q(\axi_wdata[9] ) );
  DFFPOSX1 DFFPOSX1_313 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_10__FF_INPUT), .Q(\axi_wdata[10] ) );
  DFFPOSX1 DFFPOSX1_314 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_11__FF_INPUT), .Q(\axi_wdata[11] ) );
  DFFPOSX1 DFFPOSX1_315 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_12__FF_INPUT), .Q(\axi_wdata[12] ) );
  DFFPOSX1 DFFPOSX1_316 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_13__FF_INPUT), .Q(\axi_wdata[13] ) );
  DFFPOSX1 DFFPOSX1_317 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_14__FF_INPUT), .Q(\axi_wdata[14] ) );
  DFFPOSX1 DFFPOSX1_318 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_15__FF_INPUT), .Q(\axi_wdata[15] ) );
  DFFPOSX1 DFFPOSX1_319 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_16__FF_INPUT), .Q(\axi_wdata[16] ) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(SCLK), .D(counter_31__FF_INPUT), .Q(counter_31_) );
  DFFPOSX1 DFFPOSX1_320 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_17__FF_INPUT), .Q(\axi_wdata[17] ) );
  DFFPOSX1 DFFPOSX1_321 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_18__FF_INPUT), .Q(\axi_wdata[18] ) );
  DFFPOSX1 DFFPOSX1_322 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_19__FF_INPUT), .Q(\axi_wdata[19] ) );
  DFFPOSX1 DFFPOSX1_323 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_20__FF_INPUT), .Q(\axi_wdata[20] ) );
  DFFPOSX1 DFFPOSX1_324 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_21__FF_INPUT), .Q(\axi_wdata[21] ) );
  DFFPOSX1 DFFPOSX1_325 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_22__FF_INPUT), .Q(\axi_wdata[22] ) );
  DFFPOSX1 DFFPOSX1_326 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_23__FF_INPUT), .Q(\axi_wdata[23] ) );
  DFFPOSX1 DFFPOSX1_327 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_24__FF_INPUT), .Q(\axi_wdata[24] ) );
  DFFPOSX1 DFFPOSX1_328 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_25__FF_INPUT), .Q(\axi_wdata[25] ) );
  DFFPOSX1 DFFPOSX1_329 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_26__FF_INPUT), .Q(\axi_wdata[26] ) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(SCLK), .D(counter_32__FF_INPUT), .Q(counter_32_) );
  DFFPOSX1 DFFPOSX1_330 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_27__FF_INPUT), .Q(\axi_wdata[27] ) );
  DFFPOSX1 DFFPOSX1_331 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_28__FF_INPUT), .Q(\axi_wdata[28] ) );
  DFFPOSX1 DFFPOSX1_332 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_29__FF_INPUT), .Q(\axi_wdata[29] ) );
  DFFPOSX1 DFFPOSX1_333 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_30__FF_INPUT), .Q(\axi_wdata[30] ) );
  DFFPOSX1 DFFPOSX1_334 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_31__FF_INPUT), .Q(\axi_wdata[31] ) );
  DFFPOSX1 DFFPOSX1_335 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_32__FF_INPUT), .Q(\axi_awaddr[0] ) );
  DFFPOSX1 DFFPOSX1_336 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_33__FF_INPUT), .Q(\axi_awaddr[1] ) );
  DFFPOSX1 DFFPOSX1_337 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_34__FF_INPUT), .Q(\axi_awaddr[2] ) );
  DFFPOSX1 DFFPOSX1_338 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_35__FF_INPUT), .Q(\axi_awaddr[3] ) );
  DFFPOSX1 DFFPOSX1_339 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_36__FF_INPUT), .Q(\axi_awaddr[4] ) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(SCLK), .D(counter_33__FF_INPUT), .Q(counter_33_) );
  DFFPOSX1 DFFPOSX1_340 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_37__FF_INPUT), .Q(\axi_awaddr[5] ) );
  DFFPOSX1 DFFPOSX1_341 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_38__FF_INPUT), .Q(\axi_awaddr[6] ) );
  DFFPOSX1 DFFPOSX1_342 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_39__FF_INPUT), .Q(\axi_awaddr[7] ) );
  DFFPOSX1 DFFPOSX1_343 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_40__FF_INPUT), .Q(\axi_awaddr[8] ) );
  DFFPOSX1 DFFPOSX1_344 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_41__FF_INPUT), .Q(\axi_awaddr[9] ) );
  DFFPOSX1 DFFPOSX1_345 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_42__FF_INPUT), .Q(\axi_awaddr[10] ) );
  DFFPOSX1 DFFPOSX1_346 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_43__FF_INPUT), .Q(\axi_awaddr[11] ) );
  DFFPOSX1 DFFPOSX1_347 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_44__FF_INPUT), .Q(\axi_awaddr[12] ) );
  DFFPOSX1 DFFPOSX1_348 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_45__FF_INPUT), .Q(\axi_awaddr[13] ) );
  DFFPOSX1 DFFPOSX1_349 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_46__FF_INPUT), .Q(\axi_awaddr[14] ) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(SCLK), .D(counter_34__FF_INPUT), .Q(counter_34_) );
  DFFPOSX1 DFFPOSX1_350 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_47__FF_INPUT), .Q(\axi_awaddr[15] ) );
  DFFPOSX1 DFFPOSX1_351 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_48__FF_INPUT), .Q(\axi_awaddr[16] ) );
  DFFPOSX1 DFFPOSX1_352 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_49__FF_INPUT), .Q(\axi_awaddr[17] ) );
  DFFPOSX1 DFFPOSX1_353 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_50__FF_INPUT), .Q(\axi_awaddr[18] ) );
  DFFPOSX1 DFFPOSX1_354 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_51__FF_INPUT), .Q(\axi_awaddr[19] ) );
  DFFPOSX1 DFFPOSX1_355 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_52__FF_INPUT), .Q(\axi_awaddr[20] ) );
  DFFPOSX1 DFFPOSX1_356 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_53__FF_INPUT), .Q(\axi_awaddr[21] ) );
  DFFPOSX1 DFFPOSX1_357 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_54__FF_INPUT), .Q(\axi_awaddr[22] ) );
  DFFPOSX1 DFFPOSX1_358 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_55__FF_INPUT), .Q(\axi_awaddr[23] ) );
  DFFPOSX1 DFFPOSX1_359 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_56__FF_INPUT), .Q(\axi_awaddr[24] ) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(SCLK), .D(counter_35__FF_INPUT), .Q(counter_35_) );
  DFFPOSX1 DFFPOSX1_360 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_57__FF_INPUT), .Q(\axi_awaddr[25] ) );
  DFFPOSX1 DFFPOSX1_361 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_58__FF_INPUT), .Q(\axi_awaddr[26] ) );
  DFFPOSX1 DFFPOSX1_362 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_59__FF_INPUT), .Q(\axi_awaddr[27] ) );
  DFFPOSX1 DFFPOSX1_363 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_60__FF_INPUT), .Q(\axi_awaddr[28] ) );
  DFFPOSX1 DFFPOSX1_364 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_61__FF_INPUT), .Q(\axi_awaddr[29] ) );
  DFFPOSX1 DFFPOSX1_365 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_62__FF_INPUT), .Q(\axi_awaddr[30] ) );
  DFFPOSX1 DFFPOSX1_366 ( .CLK(CLK), .D(bus_sync_axi_bus_reg_data3_63__FF_INPUT), .Q(\axi_awaddr[31] ) );
  DFFPOSX1 DFFPOSX1_367 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_0__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_0_) );
  DFFPOSX1 DFFPOSX1_368 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_1__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_1_) );
  DFFPOSX1 DFFPOSX1_369 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_2__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_2_) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(SCLK), .D(counter_36__FF_INPUT), .Q(counter_36_) );
  DFFPOSX1 DFFPOSX1_370 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_3__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_3_) );
  DFFPOSX1 DFFPOSX1_371 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_4__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_4_) );
  DFFPOSX1 DFFPOSX1_372 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_5__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_5_) );
  DFFPOSX1 DFFPOSX1_373 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_6__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_6_) );
  DFFPOSX1 DFFPOSX1_374 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_7__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_7_) );
  DFFPOSX1 DFFPOSX1_375 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_8__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_8_) );
  DFFPOSX1 DFFPOSX1_376 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_9__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_9_) );
  DFFPOSX1 DFFPOSX1_377 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_10__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_10_) );
  DFFPOSX1 DFFPOSX1_378 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_11__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_11_) );
  DFFPOSX1 DFFPOSX1_379 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_12__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_12_) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(SCLK), .D(counter_37__FF_INPUT), .Q(counter_37_) );
  DFFPOSX1 DFFPOSX1_380 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_13__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_13_) );
  DFFPOSX1 DFFPOSX1_381 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_14__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_14_) );
  DFFPOSX1 DFFPOSX1_382 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_15__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_15_) );
  DFFPOSX1 DFFPOSX1_383 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_16__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_16_) );
  DFFPOSX1 DFFPOSX1_384 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_17__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_17_) );
  DFFPOSX1 DFFPOSX1_385 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_18__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_18_) );
  DFFPOSX1 DFFPOSX1_386 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_19__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_19_) );
  DFFPOSX1 DFFPOSX1_387 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_20__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_20_) );
  DFFPOSX1 DFFPOSX1_388 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_21__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_21_) );
  DFFPOSX1 DFFPOSX1_389 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_22__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_22_) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(SCLK), .D(counter_38__FF_INPUT), .Q(counter_38_) );
  DFFPOSX1 DFFPOSX1_390 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_23__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_23_) );
  DFFPOSX1 DFFPOSX1_391 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_24__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_24_) );
  DFFPOSX1 DFFPOSX1_392 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_25__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_25_) );
  DFFPOSX1 DFFPOSX1_393 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_26__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_26_) );
  DFFPOSX1 DFFPOSX1_394 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_27__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_27_) );
  DFFPOSX1 DFFPOSX1_395 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_28__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_28_) );
  DFFPOSX1 DFFPOSX1_396 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_29__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_29_) );
  DFFPOSX1 DFFPOSX1_397 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_30__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_30_) );
  DFFPOSX1 DFFPOSX1_398 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_31__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_31_) );
  DFFPOSX1 DFFPOSX1_399 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_32__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_32_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(SCLK), .D(counter_3__FF_INPUT), .Q(counter_3_) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(SCLK), .D(counter_39__FF_INPUT), .Q(counter_39_) );
  DFFPOSX1 DFFPOSX1_400 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_33__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_33_) );
  DFFPOSX1 DFFPOSX1_401 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_34__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_34_) );
  DFFPOSX1 DFFPOSX1_402 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_35__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_35_) );
  DFFPOSX1 DFFPOSX1_403 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_36__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_36_) );
  DFFPOSX1 DFFPOSX1_404 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_37__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_37_) );
  DFFPOSX1 DFFPOSX1_405 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_38__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_38_) );
  DFFPOSX1 DFFPOSX1_406 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_39__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_39_) );
  DFFPOSX1 DFFPOSX1_407 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_40__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_40_) );
  DFFPOSX1 DFFPOSX1_408 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_41__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_41_) );
  DFFPOSX1 DFFPOSX1_409 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_42__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_42_) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(SCLK), .D(counter_40__FF_INPUT), .Q(counter_40_) );
  DFFPOSX1 DFFPOSX1_410 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_43__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_43_) );
  DFFPOSX1 DFFPOSX1_411 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_44__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_44_) );
  DFFPOSX1 DFFPOSX1_412 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_45__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_45_) );
  DFFPOSX1 DFFPOSX1_413 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_46__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_46_) );
  DFFPOSX1 DFFPOSX1_414 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_47__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_47_) );
  DFFPOSX1 DFFPOSX1_415 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_48__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_48_) );
  DFFPOSX1 DFFPOSX1_416 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_49__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_49_) );
  DFFPOSX1 DFFPOSX1_417 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_50__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_50_) );
  DFFPOSX1 DFFPOSX1_418 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_51__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_51_) );
  DFFPOSX1 DFFPOSX1_419 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_52__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_52_) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(SCLK), .D(counter_41__FF_INPUT), .Q(counter_41_) );
  DFFPOSX1 DFFPOSX1_420 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_53__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_53_) );
  DFFPOSX1 DFFPOSX1_421 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_54__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_54_) );
  DFFPOSX1 DFFPOSX1_422 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_55__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_55_) );
  DFFPOSX1 DFFPOSX1_423 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_56__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_56_) );
  DFFPOSX1 DFFPOSX1_424 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_57__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_57_) );
  DFFPOSX1 DFFPOSX1_425 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_58__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_58_) );
  DFFPOSX1 DFFPOSX1_426 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_59__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_59_) );
  DFFPOSX1 DFFPOSX1_427 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_60__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_60_) );
  DFFPOSX1 DFFPOSX1_428 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_61__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_61_) );
  DFFPOSX1 DFFPOSX1_429 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_62__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_62_) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(SCLK), .D(counter_42__FF_INPUT), .Q(counter_42_) );
  DFFPOSX1 DFFPOSX1_430 ( .CLK(SCLK), .D(bus_sync_axi_bus_reg_data1_63__FF_INPUT), .Q(bus_sync_axi_bus_reg_data1_63_) );
  DFFPOSX1 DFFPOSX1_431 ( .CLK(bus_sync_axi_bus_NCLK2), .D(bus_sync_axi_bus_ECLK1_FF_INPUT), .Q(bus_sync_axi_bus_ECLK1) );
  DFFPOSX1 DFFPOSX1_432 ( .CLK(bus_sync_axi_bus_NCLK2), .D(bus_sync_axi_bus_EECLK1_FF_INPUT), .Q(bus_sync_axi_bus_EECLK1) );
  DFFPOSX1 DFFPOSX1_433 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_0__FF_INPUT), .Q(bus_sync_rdata_data_out_0_) );
  DFFPOSX1 DFFPOSX1_434 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_1__FF_INPUT), .Q(bus_sync_rdata_data_out_1_) );
  DFFPOSX1 DFFPOSX1_435 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_2__FF_INPUT), .Q(bus_sync_rdata_data_out_2_) );
  DFFPOSX1 DFFPOSX1_436 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_3__FF_INPUT), .Q(bus_sync_rdata_data_out_3_) );
  DFFPOSX1 DFFPOSX1_437 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_4__FF_INPUT), .Q(bus_sync_rdata_data_out_4_) );
  DFFPOSX1 DFFPOSX1_438 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_5__FF_INPUT), .Q(bus_sync_rdata_data_out_5_) );
  DFFPOSX1 DFFPOSX1_439 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_6__FF_INPUT), .Q(bus_sync_rdata_data_out_6_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(SCLK), .D(counter_43__FF_INPUT), .Q(counter_43_) );
  DFFPOSX1 DFFPOSX1_440 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_7__FF_INPUT), .Q(bus_sync_rdata_data_out_7_) );
  DFFPOSX1 DFFPOSX1_441 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_8__FF_INPUT), .Q(bus_sync_rdata_data_out_8_) );
  DFFPOSX1 DFFPOSX1_442 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_9__FF_INPUT), .Q(bus_sync_rdata_data_out_9_) );
  DFFPOSX1 DFFPOSX1_443 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_10__FF_INPUT), .Q(bus_sync_rdata_data_out_10_) );
  DFFPOSX1 DFFPOSX1_444 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_11__FF_INPUT), .Q(bus_sync_rdata_data_out_11_) );
  DFFPOSX1 DFFPOSX1_445 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_12__FF_INPUT), .Q(bus_sync_rdata_data_out_12_) );
  DFFPOSX1 DFFPOSX1_446 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_13__FF_INPUT), .Q(bus_sync_rdata_data_out_13_) );
  DFFPOSX1 DFFPOSX1_447 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_14__FF_INPUT), .Q(bus_sync_rdata_data_out_14_) );
  DFFPOSX1 DFFPOSX1_448 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_15__FF_INPUT), .Q(bus_sync_rdata_data_out_15_) );
  DFFPOSX1 DFFPOSX1_449 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_16__FF_INPUT), .Q(bus_sync_rdata_data_out_16_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(SCLK), .D(counter_44__FF_INPUT), .Q(counter_44_) );
  DFFPOSX1 DFFPOSX1_450 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_17__FF_INPUT), .Q(bus_sync_rdata_data_out_17_) );
  DFFPOSX1 DFFPOSX1_451 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_18__FF_INPUT), .Q(bus_sync_rdata_data_out_18_) );
  DFFPOSX1 DFFPOSX1_452 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_19__FF_INPUT), .Q(bus_sync_rdata_data_out_19_) );
  DFFPOSX1 DFFPOSX1_453 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_20__FF_INPUT), .Q(bus_sync_rdata_data_out_20_) );
  DFFPOSX1 DFFPOSX1_454 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_21__FF_INPUT), .Q(bus_sync_rdata_data_out_21_) );
  DFFPOSX1 DFFPOSX1_455 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_22__FF_INPUT), .Q(bus_sync_rdata_data_out_22_) );
  DFFPOSX1 DFFPOSX1_456 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_23__FF_INPUT), .Q(bus_sync_rdata_data_out_23_) );
  DFFPOSX1 DFFPOSX1_457 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_24__FF_INPUT), .Q(bus_sync_rdata_data_out_24_) );
  DFFPOSX1 DFFPOSX1_458 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_25__FF_INPUT), .Q(bus_sync_rdata_data_out_25_) );
  DFFPOSX1 DFFPOSX1_459 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_26__FF_INPUT), .Q(bus_sync_rdata_data_out_26_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(SCLK), .D(counter_45__FF_INPUT), .Q(counter_45_) );
  DFFPOSX1 DFFPOSX1_460 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_27__FF_INPUT), .Q(bus_sync_rdata_data_out_27_) );
  DFFPOSX1 DFFPOSX1_461 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_28__FF_INPUT), .Q(bus_sync_rdata_data_out_28_) );
  DFFPOSX1 DFFPOSX1_462 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_29__FF_INPUT), .Q(bus_sync_rdata_data_out_29_) );
  DFFPOSX1 DFFPOSX1_463 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_30__FF_INPUT), .Q(bus_sync_rdata_data_out_30_) );
  DFFPOSX1 DFFPOSX1_464 ( .CLK(SCLK), .D(bus_sync_rdata_reg_data3_31__FF_INPUT), .Q(bus_sync_rdata_data_out_31_) );
  DFFPOSX1 DFFPOSX1_465 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_0__FF_INPUT), .Q(bus_sync_rdata_reg_data1_0_) );
  DFFPOSX1 DFFPOSX1_466 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_1__FF_INPUT), .Q(bus_sync_rdata_reg_data1_1_) );
  DFFPOSX1 DFFPOSX1_467 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_2__FF_INPUT), .Q(bus_sync_rdata_reg_data1_2_) );
  DFFPOSX1 DFFPOSX1_468 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_3__FF_INPUT), .Q(bus_sync_rdata_reg_data1_3_) );
  DFFPOSX1 DFFPOSX1_469 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_4__FF_INPUT), .Q(bus_sync_rdata_reg_data1_4_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(SCLK), .D(counter_46__FF_INPUT), .Q(counter_46_) );
  DFFPOSX1 DFFPOSX1_470 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_5__FF_INPUT), .Q(bus_sync_rdata_reg_data1_5_) );
  DFFPOSX1 DFFPOSX1_471 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_6__FF_INPUT), .Q(bus_sync_rdata_reg_data1_6_) );
  DFFPOSX1 DFFPOSX1_472 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_7__FF_INPUT), .Q(bus_sync_rdata_reg_data1_7_) );
  DFFPOSX1 DFFPOSX1_473 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_8__FF_INPUT), .Q(bus_sync_rdata_reg_data1_8_) );
  DFFPOSX1 DFFPOSX1_474 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_9__FF_INPUT), .Q(bus_sync_rdata_reg_data1_9_) );
  DFFPOSX1 DFFPOSX1_475 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_10__FF_INPUT), .Q(bus_sync_rdata_reg_data1_10_) );
  DFFPOSX1 DFFPOSX1_476 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_11__FF_INPUT), .Q(bus_sync_rdata_reg_data1_11_) );
  DFFPOSX1 DFFPOSX1_477 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_12__FF_INPUT), .Q(bus_sync_rdata_reg_data1_12_) );
  DFFPOSX1 DFFPOSX1_478 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_13__FF_INPUT), .Q(bus_sync_rdata_reg_data1_13_) );
  DFFPOSX1 DFFPOSX1_479 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_14__FF_INPUT), .Q(bus_sync_rdata_reg_data1_14_) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(SCLK), .D(counter_47__FF_INPUT), .Q(counter_47_) );
  DFFPOSX1 DFFPOSX1_480 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_15__FF_INPUT), .Q(bus_sync_rdata_reg_data1_15_) );
  DFFPOSX1 DFFPOSX1_481 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_16__FF_INPUT), .Q(bus_sync_rdata_reg_data1_16_) );
  DFFPOSX1 DFFPOSX1_482 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_17__FF_INPUT), .Q(bus_sync_rdata_reg_data1_17_) );
  DFFPOSX1 DFFPOSX1_483 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_18__FF_INPUT), .Q(bus_sync_rdata_reg_data1_18_) );
  DFFPOSX1 DFFPOSX1_484 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_19__FF_INPUT), .Q(bus_sync_rdata_reg_data1_19_) );
  DFFPOSX1 DFFPOSX1_485 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_20__FF_INPUT), .Q(bus_sync_rdata_reg_data1_20_) );
  DFFPOSX1 DFFPOSX1_486 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_21__FF_INPUT), .Q(bus_sync_rdata_reg_data1_21_) );
  DFFPOSX1 DFFPOSX1_487 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_22__FF_INPUT), .Q(bus_sync_rdata_reg_data1_22_) );
  DFFPOSX1 DFFPOSX1_488 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_23__FF_INPUT), .Q(bus_sync_rdata_reg_data1_23_) );
  DFFPOSX1 DFFPOSX1_489 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_24__FF_INPUT), .Q(bus_sync_rdata_reg_data1_24_) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(SCLK), .D(counter_48__FF_INPUT), .Q(counter_48_) );
  DFFPOSX1 DFFPOSX1_490 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_25__FF_INPUT), .Q(bus_sync_rdata_reg_data1_25_) );
  DFFPOSX1 DFFPOSX1_491 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_26__FF_INPUT), .Q(bus_sync_rdata_reg_data1_26_) );
  DFFPOSX1 DFFPOSX1_492 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_27__FF_INPUT), .Q(bus_sync_rdata_reg_data1_27_) );
  DFFPOSX1 DFFPOSX1_493 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_28__FF_INPUT), .Q(bus_sync_rdata_reg_data1_28_) );
  DFFPOSX1 DFFPOSX1_494 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_29__FF_INPUT), .Q(bus_sync_rdata_reg_data1_29_) );
  DFFPOSX1 DFFPOSX1_495 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_30__FF_INPUT), .Q(bus_sync_rdata_reg_data1_30_) );
  DFFPOSX1 DFFPOSX1_496 ( .CLK(CLK), .D(bus_sync_rdata_reg_data1_31__FF_INPUT), .Q(bus_sync_rdata_reg_data1_31_) );
  DFFPOSX1 DFFPOSX1_497 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_0__FF_INPUT), .Q(bus_sync_rdata_reg_data2_0_) );
  DFFPOSX1 DFFPOSX1_498 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_1__FF_INPUT), .Q(bus_sync_rdata_reg_data2_1_) );
  DFFPOSX1 DFFPOSX1_499 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_2__FF_INPUT), .Q(bus_sync_rdata_reg_data2_2_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(SCLK), .D(counter_4__FF_INPUT), .Q(counter_4_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(SCLK), .D(counter_49__FF_INPUT), .Q(counter_49_) );
  DFFPOSX1 DFFPOSX1_500 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_3__FF_INPUT), .Q(bus_sync_rdata_reg_data2_3_) );
  DFFPOSX1 DFFPOSX1_501 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_4__FF_INPUT), .Q(bus_sync_rdata_reg_data2_4_) );
  DFFPOSX1 DFFPOSX1_502 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_5__FF_INPUT), .Q(bus_sync_rdata_reg_data2_5_) );
  DFFPOSX1 DFFPOSX1_503 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_6__FF_INPUT), .Q(bus_sync_rdata_reg_data2_6_) );
  DFFPOSX1 DFFPOSX1_504 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_7__FF_INPUT), .Q(bus_sync_rdata_reg_data2_7_) );
  DFFPOSX1 DFFPOSX1_505 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_8__FF_INPUT), .Q(bus_sync_rdata_reg_data2_8_) );
  DFFPOSX1 DFFPOSX1_506 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_9__FF_INPUT), .Q(bus_sync_rdata_reg_data2_9_) );
  DFFPOSX1 DFFPOSX1_507 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_10__FF_INPUT), .Q(bus_sync_rdata_reg_data2_10_) );
  DFFPOSX1 DFFPOSX1_508 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_11__FF_INPUT), .Q(bus_sync_rdata_reg_data2_11_) );
  DFFPOSX1 DFFPOSX1_509 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_12__FF_INPUT), .Q(bus_sync_rdata_reg_data2_12_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(SCLK), .D(counter_50__FF_INPUT), .Q(counter_50_) );
  DFFPOSX1 DFFPOSX1_510 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_13__FF_INPUT), .Q(bus_sync_rdata_reg_data2_13_) );
  DFFPOSX1 DFFPOSX1_511 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_14__FF_INPUT), .Q(bus_sync_rdata_reg_data2_14_) );
  DFFPOSX1 DFFPOSX1_512 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_15__FF_INPUT), .Q(bus_sync_rdata_reg_data2_15_) );
  DFFPOSX1 DFFPOSX1_513 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_16__FF_INPUT), .Q(bus_sync_rdata_reg_data2_16_) );
  DFFPOSX1 DFFPOSX1_514 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_17__FF_INPUT), .Q(bus_sync_rdata_reg_data2_17_) );
  DFFPOSX1 DFFPOSX1_515 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_18__FF_INPUT), .Q(bus_sync_rdata_reg_data2_18_) );
  DFFPOSX1 DFFPOSX1_516 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_19__FF_INPUT), .Q(bus_sync_rdata_reg_data2_19_) );
  DFFPOSX1 DFFPOSX1_517 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_20__FF_INPUT), .Q(bus_sync_rdata_reg_data2_20_) );
  DFFPOSX1 DFFPOSX1_518 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_21__FF_INPUT), .Q(bus_sync_rdata_reg_data2_21_) );
  DFFPOSX1 DFFPOSX1_519 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_22__FF_INPUT), .Q(bus_sync_rdata_reg_data2_22_) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(SCLK), .D(counter_51__FF_INPUT), .Q(counter_51_) );
  DFFPOSX1 DFFPOSX1_520 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_23__FF_INPUT), .Q(bus_sync_rdata_reg_data2_23_) );
  DFFPOSX1 DFFPOSX1_521 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_24__FF_INPUT), .Q(bus_sync_rdata_reg_data2_24_) );
  DFFPOSX1 DFFPOSX1_522 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_25__FF_INPUT), .Q(bus_sync_rdata_reg_data2_25_) );
  DFFPOSX1 DFFPOSX1_523 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_26__FF_INPUT), .Q(bus_sync_rdata_reg_data2_26_) );
  DFFPOSX1 DFFPOSX1_524 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_27__FF_INPUT), .Q(bus_sync_rdata_reg_data2_27_) );
  DFFPOSX1 DFFPOSX1_525 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_28__FF_INPUT), .Q(bus_sync_rdata_reg_data2_28_) );
  DFFPOSX1 DFFPOSX1_526 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_29__FF_INPUT), .Q(bus_sync_rdata_reg_data2_29_) );
  DFFPOSX1 DFFPOSX1_527 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_30__FF_INPUT), .Q(bus_sync_rdata_reg_data2_30_) );
  DFFPOSX1 DFFPOSX1_528 ( .CLK(CLK), .D(bus_sync_rdata_reg_data2_31__FF_INPUT), .Q(bus_sync_rdata_reg_data2_31_) );
  DFFPOSX1 DFFPOSX1_529 ( .CLK(bus_sync_rdata_NCLK1), .D(bus_sync_rdata_ECLK2_FF_INPUT), .Q(bus_sync_rdata_ECLK2) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(SCLK), .D(counter_52__FF_INPUT), .Q(counter_52_) );
  DFFPOSX1 DFFPOSX1_530 ( .CLK(bus_sync_rdata_NCLK1), .D(bus_sync_rdata_EECLK2_FF_INPUT), .Q(bus_sync_rdata_EECLK2) );
  DFFPOSX1 DFFPOSX1_531 ( .CLK(CLK), .D(bus_sync_state_machine_reg_data2_0__FF_INPUT), .Q(bus_sync_state_machine_reg_data2_0_) );
  DFFPOSX1 DFFPOSX1_532 ( .CLK(CLK), .D(bus_sync_state_machine_reg_data2_1__FF_INPUT), .Q(bus_sync_state_machine_reg_data2_1_) );
  DFFPOSX1 DFFPOSX1_533 ( .CLK(CLK), .D(bus_sync_state_machine_reg_data2_2__FF_INPUT), .Q(bus_sync_state_machine_reg_data2_2_) );
  DFFPOSX1 DFFPOSX1_534 ( .CLK(CLK), .D(bus_sync_state_machine_reg_data2_3__FF_INPUT), .Q(bus_sync_state_machine_reg_data2_3_) );
  DFFPOSX1 DFFPOSX1_535 ( .CLK(CLK), .D(bus_sync_state_machine_reg_data3_0__FF_INPUT), .Q(fini_spi_clk) );
  DFFPOSX1 DFFPOSX1_536 ( .CLK(CLK), .D(bus_sync_state_machine_reg_data3_1__FF_INPUT), .Q(re_clk) );
  DFFPOSX1 DFFPOSX1_537 ( .CLK(CLK), .D(bus_sync_state_machine_reg_data3_2__FF_INPUT), .Q(we_clk) );
  DFFPOSX1 DFFPOSX1_538 ( .CLK(CLK), .D(bus_sync_state_machine_reg_data3_3__FF_INPUT), .Q(PICORV_RST) );
  DFFPOSX1 DFFPOSX1_539 ( .CLK(SCLK), .D(bus_sync_state_machine_reg_data1_0__FF_INPUT), .Q(bus_sync_state_machine_reg_data1_0_) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(SCLK), .D(counter_53__FF_INPUT), .Q(counter_53_) );
  DFFPOSX1 DFFPOSX1_540 ( .CLK(SCLK), .D(bus_sync_state_machine_reg_data1_1__FF_INPUT), .Q(bus_sync_state_machine_reg_data1_1_) );
  DFFPOSX1 DFFPOSX1_541 ( .CLK(SCLK), .D(bus_sync_state_machine_reg_data1_2__FF_INPUT), .Q(bus_sync_state_machine_reg_data1_2_) );
  DFFPOSX1 DFFPOSX1_542 ( .CLK(SCLK), .D(bus_sync_state_machine_reg_data1_3__FF_INPUT), .Q(bus_sync_state_machine_reg_data1_3_) );
  DFFPOSX1 DFFPOSX1_543 ( .CLK(bus_sync_state_machine_NCLK2), .D(bus_sync_state_machine_ECLK1_FF_INPUT), .Q(bus_sync_state_machine_ECLK1) );
  DFFPOSX1 DFFPOSX1_544 ( .CLK(bus_sync_state_machine_NCLK2), .D(bus_sync_state_machine_EECLK1_FF_INPUT), .Q(bus_sync_state_machine_EECLK1) );
  DFFPOSX1 DFFPOSX1_545 ( .CLK(SCLK), .D(bus_sync_status_reg_data3_0__FF_INPUT), .Q(bus_sync_status_data_out_0_) );
  DFFPOSX1 DFFPOSX1_546 ( .CLK(SCLK), .D(bus_sync_status_reg_data3_1__FF_INPUT), .Q(bus_sync_status_data_out_1_) );
  DFFPOSX1 DFFPOSX1_547 ( .CLK(SCLK), .D(bus_sync_status_reg_data3_2__FF_INPUT), .Q(bus_sync_status_data_out_2_) );
  DFFPOSX1 DFFPOSX1_548 ( .CLK(CLK), .D(bus_sync_status_reg_data1_0__FF_INPUT), .Q(bus_sync_status_reg_data1_0_) );
  DFFPOSX1 DFFPOSX1_549 ( .CLK(CLK), .D(bus_sync_status_reg_data1_1__FF_INPUT), .Q(bus_sync_status_reg_data1_1_) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(SCLK), .D(counter_54__FF_INPUT), .Q(counter_54_) );
  DFFPOSX1 DFFPOSX1_550 ( .CLK(CLK), .D(bus_sync_status_reg_data1_2__FF_INPUT), .Q(bus_sync_status_reg_data1_2_) );
  DFFPOSX1 DFFPOSX1_551 ( .CLK(CLK), .D(bus_sync_status_reg_data2_0__FF_INPUT), .Q(bus_sync_status_reg_data2_0_) );
  DFFPOSX1 DFFPOSX1_552 ( .CLK(CLK), .D(bus_sync_status_reg_data2_1__FF_INPUT), .Q(bus_sync_status_reg_data2_1_) );
  DFFPOSX1 DFFPOSX1_553 ( .CLK(CLK), .D(bus_sync_status_reg_data2_2__FF_INPUT), .Q(bus_sync_status_reg_data2_2_) );
  DFFPOSX1 DFFPOSX1_554 ( .CLK(bus_sync_status_NCLK1), .D(bus_sync_status_ECLK2_FF_INPUT), .Q(bus_sync_status_ECLK2) );
  DFFPOSX1 DFFPOSX1_555 ( .CLK(bus_sync_status_NCLK1), .D(bus_sync_status_EECLK2_FF_INPUT), .Q(bus_sync_status_EECLK2) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(SCLK), .D(counter_55__FF_INPUT), .Q(counter_55_) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(SCLK), .D(counter_56__FF_INPUT), .Q(counter_56_) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(SCLK), .D(counter_57__FF_INPUT), .Q(counter_57_) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(SCLK), .D(counter_58__FF_INPUT), .Q(counter_58_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(SCLK), .D(counter_5__FF_INPUT), .Q(counter_5_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(SCLK), .D(counter_59__FF_INPUT), .Q(counter_59_) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(SCLK), .D(counter_60__FF_INPUT), .Q(counter_60_) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(SCLK), .D(counter_61__FF_INPUT), .Q(counter_61_) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(SCLK), .D(counter_62__FF_INPUT), .Q(counter_62_) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(SCLK), .D(counter_63__FF_INPUT), .Q(counter_63_) );
  DFFPOSX1 DFFPOSX1_65 ( .CLK(SCLK), .D(counter_64__FF_INPUT), .Q(counter_64_) );
  DFFPOSX1 DFFPOSX1_66 ( .CLK(SCLK), .D(counter_65__FF_INPUT), .Q(counter_65_) );
  DFFPOSX1 DFFPOSX1_67 ( .CLK(SCLK), .D(fini_spi_FF_INPUT), .Q(fini_spi) );
  DFFPOSX1 DFFPOSX1_68 ( .CLK(SCLK), .D(bus_cap_0__FF_INPUT), .Q(bus_cap_0_) );
  DFFPOSX1 DFFPOSX1_69 ( .CLK(SCLK), .D(bus_cap_1__FF_INPUT), .Q(bus_cap_1_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(SCLK), .D(counter_6__FF_INPUT), .Q(counter_6_) );
  DFFPOSX1 DFFPOSX1_70 ( .CLK(SCLK), .D(bus_cap_2__FF_INPUT), .Q(bus_cap_2_) );
  DFFPOSX1 DFFPOSX1_71 ( .CLK(SCLK), .D(bus_cap_3__FF_INPUT), .Q(bus_cap_3_) );
  DFFPOSX1 DFFPOSX1_72 ( .CLK(SCLK), .D(bus_cap_4__FF_INPUT), .Q(bus_cap_4_) );
  DFFPOSX1 DFFPOSX1_73 ( .CLK(SCLK), .D(bus_cap_5__FF_INPUT), .Q(bus_cap_5_) );
  DFFPOSX1 DFFPOSX1_74 ( .CLK(SCLK), .D(bus_cap_6__FF_INPUT), .Q(bus_cap_6_) );
  DFFPOSX1 DFFPOSX1_75 ( .CLK(SCLK), .D(bus_cap_7__FF_INPUT), .Q(bus_cap_7_) );
  DFFPOSX1 DFFPOSX1_76 ( .CLK(SCLK), .D(bus_cap_8__FF_INPUT), .Q(bus_cap_8_) );
  DFFPOSX1 DFFPOSX1_77 ( .CLK(SCLK), .D(bus_cap_9__FF_INPUT), .Q(bus_cap_9_) );
  DFFPOSX1 DFFPOSX1_78 ( .CLK(SCLK), .D(bus_cap_10__FF_INPUT), .Q(bus_cap_10_) );
  DFFPOSX1 DFFPOSX1_79 ( .CLK(SCLK), .D(bus_cap_11__FF_INPUT), .Q(bus_cap_11_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(SCLK), .D(counter_7__FF_INPUT), .Q(counter_7_) );
  DFFPOSX1 DFFPOSX1_80 ( .CLK(SCLK), .D(bus_cap_12__FF_INPUT), .Q(bus_cap_12_) );
  DFFPOSX1 DFFPOSX1_81 ( .CLK(SCLK), .D(bus_cap_13__FF_INPUT), .Q(bus_cap_13_) );
  DFFPOSX1 DFFPOSX1_82 ( .CLK(SCLK), .D(bus_cap_14__FF_INPUT), .Q(bus_cap_14_) );
  DFFPOSX1 DFFPOSX1_83 ( .CLK(SCLK), .D(bus_cap_15__FF_INPUT), .Q(bus_cap_15_) );
  DFFPOSX1 DFFPOSX1_84 ( .CLK(SCLK), .D(bus_cap_16__FF_INPUT), .Q(bus_cap_16_) );
  DFFPOSX1 DFFPOSX1_85 ( .CLK(SCLK), .D(bus_cap_17__FF_INPUT), .Q(bus_cap_17_) );
  DFFPOSX1 DFFPOSX1_86 ( .CLK(SCLK), .D(bus_cap_18__FF_INPUT), .Q(bus_cap_18_) );
  DFFPOSX1 DFFPOSX1_87 ( .CLK(SCLK), .D(bus_cap_19__FF_INPUT), .Q(bus_cap_19_) );
  DFFPOSX1 DFFPOSX1_88 ( .CLK(SCLK), .D(bus_cap_20__FF_INPUT), .Q(bus_cap_20_) );
  DFFPOSX1 DFFPOSX1_89 ( .CLK(SCLK), .D(bus_cap_21__FF_INPUT), .Q(bus_cap_21_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(SCLK), .D(counter_8__FF_INPUT), .Q(counter_8_) );
  DFFPOSX1 DFFPOSX1_90 ( .CLK(SCLK), .D(bus_cap_22__FF_INPUT), .Q(bus_cap_22_) );
  DFFPOSX1 DFFPOSX1_91 ( .CLK(SCLK), .D(bus_cap_23__FF_INPUT), .Q(bus_cap_23_) );
  DFFPOSX1 DFFPOSX1_92 ( .CLK(SCLK), .D(bus_cap_24__FF_INPUT), .Q(bus_cap_24_) );
  DFFPOSX1 DFFPOSX1_93 ( .CLK(SCLK), .D(bus_cap_25__FF_INPUT), .Q(bus_cap_25_) );
  DFFPOSX1 DFFPOSX1_94 ( .CLK(SCLK), .D(bus_cap_26__FF_INPUT), .Q(bus_cap_26_) );
  DFFPOSX1 DFFPOSX1_95 ( .CLK(SCLK), .D(bus_cap_27__FF_INPUT), .Q(bus_cap_27_) );
  DFFPOSX1 DFFPOSX1_96 ( .CLK(SCLK), .D(bus_cap_28__FF_INPUT), .Q(bus_cap_28_) );
  DFFPOSX1 DFFPOSX1_97 ( .CLK(SCLK), .D(bus_cap_29__FF_INPUT), .Q(bus_cap_29_) );
  DFFPOSX1 DFFPOSX1_98 ( .CLK(SCLK), .D(bus_cap_30__FF_INPUT), .Q(bus_cap_30_) );
  DFFPOSX1 DFFPOSX1_99 ( .CLK(SCLK), .D(bus_cap_31__FF_INPUT), .Q(DOUT) );
  INVX1 INVX1_1 ( .A(RST), .Y(_abc_4108_n561) );
  INVX1 INVX1_10 ( .A(DATA), .Y(_abc_4108_n599_1) );
  INVX1 INVX1_100 ( .A(WDATA_12_), .Y(_abc_4108_n992) );
  INVX1 INVX1_101 ( .A(WDATA_13_), .Y(_abc_4108_n995) );
  INVX1 INVX1_102 ( .A(WDATA_14_), .Y(_abc_4108_n998) );
  INVX1 INVX1_103 ( .A(WDATA_15_), .Y(_abc_4108_n1001) );
  INVX1 INVX1_104 ( .A(WDATA_16_), .Y(_abc_4108_n1004) );
  INVX1 INVX1_105 ( .A(WDATA_17_), .Y(_abc_4108_n1007) );
  INVX1 INVX1_106 ( .A(WDATA_18_), .Y(_abc_4108_n1010) );
  INVX1 INVX1_107 ( .A(WDATA_19_), .Y(_abc_4108_n1013) );
  INVX1 INVX1_108 ( .A(WDATA_20_), .Y(_abc_4108_n1016) );
  INVX1 INVX1_109 ( .A(WDATA_21_), .Y(_abc_4108_n1019) );
  INVX1 INVX1_11 ( .A(counter_2_), .Y(_abc_4108_n615) );
  INVX1 INVX1_110 ( .A(WDATA_22_), .Y(_abc_4108_n1022) );
  INVX1 INVX1_111 ( .A(WDATA_23_), .Y(_abc_4108_n1025) );
  INVX1 INVX1_112 ( .A(WDATA_24_), .Y(_abc_4108_n1028) );
  INVX1 INVX1_113 ( .A(WDATA_25_), .Y(_abc_4108_n1031) );
  INVX1 INVX1_114 ( .A(WDATA_26_), .Y(_abc_4108_n1034) );
  INVX1 INVX1_115 ( .A(WDATA_27_), .Y(_abc_4108_n1037) );
  INVX1 INVX1_116 ( .A(WDATA_28_), .Y(_abc_4108_n1040) );
  INVX1 INVX1_117 ( .A(WDATA_29_), .Y(_abc_4108_n1043) );
  INVX1 INVX1_118 ( .A(WDATA_30_), .Y(_abc_4108_n1046) );
  INVX1 INVX1_119 ( .A(WDATA_31_), .Y(_abc_4108_n1049) );
  INVX1 INVX1_12 ( .A(counter_3_), .Y(_abc_4108_n616) );
  INVX1 INVX1_120 ( .A(A_ADDR_0_), .Y(_abc_4108_n1052) );
  INVX1 INVX1_121 ( .A(counter_33_), .Y(_abc_4108_n1053) );
  INVX1 INVX1_122 ( .A(A_ADDR_1_), .Y(_abc_4108_n1059) );
  INVX1 INVX1_123 ( .A(A_ADDR_2_), .Y(_abc_4108_n1062) );
  INVX1 INVX1_124 ( .A(A_ADDR_3_), .Y(_abc_4108_n1065) );
  INVX1 INVX1_125 ( .A(A_ADDR_4_), .Y(_abc_4108_n1068) );
  INVX1 INVX1_126 ( .A(A_ADDR_5_), .Y(_abc_4108_n1071) );
  INVX1 INVX1_127 ( .A(A_ADDR_6_), .Y(_abc_4108_n1074) );
  INVX1 INVX1_128 ( .A(A_ADDR_7_), .Y(_abc_4108_n1077) );
  INVX1 INVX1_129 ( .A(A_ADDR_8_), .Y(_abc_4108_n1080) );
  INVX1 INVX1_13 ( .A(counter_18_), .Y(_abc_4108_n624_1) );
  INVX1 INVX1_130 ( .A(A_ADDR_9_), .Y(_abc_4108_n1083) );
  INVX1 INVX1_131 ( .A(A_ADDR_10_), .Y(_abc_4108_n1086) );
  INVX1 INVX1_132 ( .A(A_ADDR_11_), .Y(_abc_4108_n1089) );
  INVX1 INVX1_133 ( .A(A_ADDR_12_), .Y(_abc_4108_n1092) );
  INVX1 INVX1_134 ( .A(A_ADDR_13_), .Y(_abc_4108_n1095) );
  INVX1 INVX1_135 ( .A(A_ADDR_14_), .Y(_abc_4108_n1098) );
  INVX1 INVX1_136 ( .A(A_ADDR_15_), .Y(_abc_4108_n1101) );
  INVX1 INVX1_137 ( .A(A_ADDR_16_), .Y(_abc_4108_n1104) );
  INVX1 INVX1_138 ( .A(A_ADDR_17_), .Y(_abc_4108_n1107) );
  INVX1 INVX1_139 ( .A(A_ADDR_18_), .Y(_abc_4108_n1110) );
  INVX1 INVX1_14 ( .A(counter_19_), .Y(_abc_4108_n625) );
  INVX1 INVX1_140 ( .A(A_ADDR_19_), .Y(_abc_4108_n1113) );
  INVX1 INVX1_141 ( .A(A_ADDR_20_), .Y(_abc_4108_n1116) );
  INVX1 INVX1_142 ( .A(A_ADDR_21_), .Y(_abc_4108_n1119) );
  INVX1 INVX1_143 ( .A(A_ADDR_22_), .Y(_abc_4108_n1122) );
  INVX1 INVX1_144 ( .A(A_ADDR_23_), .Y(_abc_4108_n1125) );
  INVX1 INVX1_145 ( .A(A_ADDR_24_), .Y(_abc_4108_n1128) );
  INVX1 INVX1_146 ( .A(A_ADDR_25_), .Y(_abc_4108_n1131) );
  INVX1 INVX1_147 ( .A(A_ADDR_26_), .Y(_abc_4108_n1134) );
  INVX1 INVX1_148 ( .A(A_ADDR_27_), .Y(_abc_4108_n1137) );
  INVX1 INVX1_149 ( .A(A_ADDR_28_), .Y(_abc_4108_n1140) );
  INVX1 INVX1_15 ( .A(counter_6_), .Y(_abc_4108_n632) );
  INVX1 INVX1_150 ( .A(A_ADDR_29_), .Y(_abc_4108_n1143) );
  INVX1 INVX1_151 ( .A(A_ADDR_30_), .Y(_abc_4108_n1146) );
  INVX1 INVX1_152 ( .A(A_ADDR_31_), .Y(_abc_4108_n1149) );
  INVX1 INVX1_153 ( .A(sft_reg_0_), .Y(_abc_4108_n1152) );
  INVX1 INVX1_154 ( .A(sft_reg_1_), .Y(_abc_4108_n1154) );
  INVX1 INVX1_155 ( .A(sft_reg_2_), .Y(_abc_4108_n1156) );
  INVX1 INVX1_156 ( .A(sft_reg_3_), .Y(_abc_4108_n1158) );
  INVX1 INVX1_157 ( .A(sft_reg_4_), .Y(_abc_4108_n1160) );
  INVX1 INVX1_158 ( .A(sft_reg_5_), .Y(_abc_4108_n1162) );
  INVX1 INVX1_159 ( .A(sft_reg_6_), .Y(_abc_4108_n1164) );
  INVX1 INVX1_16 ( .A(counter_7_), .Y(_abc_4108_n633_1) );
  INVX1 INVX1_160 ( .A(sft_reg_7_), .Y(_abc_4108_n1166) );
  INVX1 INVX1_161 ( .A(sft_reg_8_), .Y(_abc_4108_n1168) );
  INVX1 INVX1_162 ( .A(sft_reg_9_), .Y(_abc_4108_n1170) );
  INVX1 INVX1_163 ( .A(sft_reg_10_), .Y(_abc_4108_n1172) );
  INVX1 INVX1_164 ( .A(sft_reg_11_), .Y(_abc_4108_n1174) );
  INVX1 INVX1_165 ( .A(sft_reg_12_), .Y(_abc_4108_n1176) );
  INVX1 INVX1_166 ( .A(sft_reg_13_), .Y(_abc_4108_n1178) );
  INVX1 INVX1_167 ( .A(sft_reg_14_), .Y(_abc_4108_n1180) );
  INVX1 INVX1_168 ( .A(sft_reg_15_), .Y(_abc_4108_n1182) );
  INVX1 INVX1_169 ( .A(sft_reg_16_), .Y(_abc_4108_n1184) );
  INVX1 INVX1_17 ( .A(_abc_4108_n598_1), .Y(_abc_4108_n640) );
  INVX1 INVX1_170 ( .A(sft_reg_17_), .Y(_abc_4108_n1186) );
  INVX1 INVX1_171 ( .A(sft_reg_18_), .Y(_abc_4108_n1188) );
  INVX1 INVX1_172 ( .A(sft_reg_19_), .Y(_abc_4108_n1190) );
  INVX1 INVX1_173 ( .A(sft_reg_20_), .Y(_abc_4108_n1192) );
  INVX1 INVX1_174 ( .A(sft_reg_21_), .Y(_abc_4108_n1194) );
  INVX1 INVX1_175 ( .A(sft_reg_22_), .Y(_abc_4108_n1196) );
  INVX1 INVX1_176 ( .A(sft_reg_23_), .Y(_abc_4108_n1198) );
  INVX1 INVX1_177 ( .A(sft_reg_24_), .Y(_abc_4108_n1200) );
  INVX1 INVX1_178 ( .A(sft_reg_25_), .Y(_abc_4108_n1202) );
  INVX1 INVX1_179 ( .A(sft_reg_26_), .Y(_abc_4108_n1204) );
  INVX1 INVX1_18 ( .A(_abc_4108_n642_1), .Y(_abc_4108_n643) );
  INVX1 INVX1_180 ( .A(sft_reg_27_), .Y(_abc_4108_n1206) );
  INVX1 INVX1_181 ( .A(sft_reg_28_), .Y(_abc_4108_n1208) );
  INVX1 INVX1_182 ( .A(sft_reg_29_), .Y(_abc_4108_n1210) );
  INVX1 INVX1_183 ( .A(sft_reg_30_), .Y(_abc_4108_n1212) );
  INVX1 INVX1_184 ( .A(counter_5_), .Y(_abc_4108_n1221) );
  INVX1 INVX1_185 ( .A(counter_8_), .Y(_abc_4108_n1225) );
  INVX1 INVX1_186 ( .A(counter_10_), .Y(_abc_4108_n1228) );
  INVX1 INVX1_187 ( .A(counter_11_), .Y(_abc_4108_n1230) );
  INVX1 INVX1_188 ( .A(counter_12_), .Y(_abc_4108_n1232) );
  INVX1 INVX1_189 ( .A(counter_13_), .Y(_abc_4108_n1234) );
  INVX1 INVX1_19 ( .A(_abc_4108_n648), .Y(_abc_4108_n649_1) );
  INVX1 INVX1_190 ( .A(counter_14_), .Y(_abc_4108_n1236) );
  INVX1 INVX1_191 ( .A(counter_15_), .Y(_abc_4108_n1238) );
  INVX1 INVX1_192 ( .A(counter_16_), .Y(_abc_4108_n1240) );
  INVX1 INVX1_193 ( .A(counter_17_), .Y(_abc_4108_n1242) );
  INVX1 INVX1_194 ( .A(counter_20_), .Y(_abc_4108_n1246) );
  INVX1 INVX1_195 ( .A(counter_21_), .Y(_abc_4108_n1248) );
  INVX1 INVX1_196 ( .A(counter_22_), .Y(_abc_4108_n1250) );
  INVX1 INVX1_197 ( .A(counter_23_), .Y(_abc_4108_n1252) );
  INVX1 INVX1_198 ( .A(counter_24_), .Y(_abc_4108_n1254) );
  INVX1 INVX1_199 ( .A(counter_26_), .Y(_abc_4108_n1257) );
  INVX1 INVX1_2 ( .A(axi_wready), .Y(_abc_4108_n562_1) );
  INVX1 INVX1_20 ( .A(bus_cap_2_), .Y(_abc_4108_n652) );
  INVX1 INVX1_200 ( .A(counter_27_), .Y(_abc_4108_n1259) );
  INVX1 INVX1_201 ( .A(counter_28_), .Y(_abc_4108_n1261) );
  INVX1 INVX1_202 ( .A(counter_30_), .Y(_abc_4108_n1264) );
  INVX1 INVX1_203 ( .A(counter_31_), .Y(_abc_4108_n1266) );
  INVX1 INVX1_204 ( .A(counter_32_), .Y(_abc_4108_n1268) );
  INVX1 INVX1_205 ( .A(counter_34_), .Y(_abc_4108_n1271) );
  INVX1 INVX1_206 ( .A(counter_35_), .Y(_abc_4108_n1273) );
  INVX1 INVX1_207 ( .A(counter_36_), .Y(_abc_4108_n1275) );
  INVX1 INVX1_208 ( .A(counter_37_), .Y(_abc_4108_n1277) );
  INVX1 INVX1_209 ( .A(counter_38_), .Y(_abc_4108_n1279) );
  INVX1 INVX1_21 ( .A(_abc_4108_n656), .Y(_abc_4108_n657_1) );
  INVX1 INVX1_210 ( .A(counter_39_), .Y(_abc_4108_n1281) );
  INVX1 INVX1_211 ( .A(counter_40_), .Y(_abc_4108_n1283) );
  INVX1 INVX1_212 ( .A(counter_41_), .Y(_abc_4108_n1285) );
  INVX1 INVX1_213 ( .A(counter_42_), .Y(_abc_4108_n1287) );
  INVX1 INVX1_214 ( .A(counter_43_), .Y(_abc_4108_n1289) );
  INVX1 INVX1_215 ( .A(counter_44_), .Y(_abc_4108_n1291) );
  INVX1 INVX1_216 ( .A(counter_45_), .Y(_abc_4108_n1293) );
  INVX1 INVX1_217 ( .A(counter_46_), .Y(_abc_4108_n1295) );
  INVX1 INVX1_218 ( .A(counter_47_), .Y(_abc_4108_n1297) );
  INVX1 INVX1_219 ( .A(counter_48_), .Y(_abc_4108_n1299) );
  INVX1 INVX1_22 ( .A(counter_29_), .Y(_abc_4108_n661_1) );
  INVX1 INVX1_220 ( .A(counter_49_), .Y(_abc_4108_n1301) );
  INVX1 INVX1_221 ( .A(counter_50_), .Y(_abc_4108_n1303) );
  INVX1 INVX1_222 ( .A(counter_51_), .Y(_abc_4108_n1305) );
  INVX1 INVX1_223 ( .A(counter_52_), .Y(_abc_4108_n1307) );
  INVX1 INVX1_224 ( .A(counter_53_), .Y(_abc_4108_n1309) );
  INVX1 INVX1_225 ( .A(counter_54_), .Y(_abc_4108_n1311) );
  INVX1 INVX1_226 ( .A(counter_55_), .Y(_abc_4108_n1313) );
  INVX1 INVX1_227 ( .A(counter_56_), .Y(_abc_4108_n1315) );
  INVX1 INVX1_228 ( .A(counter_57_), .Y(_abc_4108_n1317) );
  INVX1 INVX1_229 ( .A(counter_58_), .Y(_abc_4108_n1319) );
  INVX1 INVX1_23 ( .A(counter_25_), .Y(_abc_4108_n662_1) );
  INVX1 INVX1_230 ( .A(counter_59_), .Y(_abc_4108_n1321) );
  INVX1 INVX1_231 ( .A(counter_60_), .Y(_abc_4108_n1323) );
  INVX1 INVX1_232 ( .A(counter_61_), .Y(_abc_4108_n1325) );
  INVX1 INVX1_233 ( .A(counter_62_), .Y(_abc_4108_n1327) );
  INVX1 INVX1_234 ( .A(counter_63_), .Y(_abc_4108_n1329) );
  INVX1 INVX1_235 ( .A(counter_64_), .Y(_abc_4108_n1331) );
  INVX1 INVX1_236 ( .A(PICORV_RST_SPI), .Y(_abc_4108_n1333) );
  INVX1 INVX1_237 ( .A(_abc_4108_n602_1), .Y(_abc_4108_n1334) );
  INVX1 INVX1_238 ( .A(_abc_4108_n1341), .Y(_abc_2913_n1025) );
  INVX1 INVX1_239 ( .A(_abc_4108_n1345), .Y(_abc_2913_n1036) );
  INVX1 INVX1_24 ( .A(counter_4_), .Y(_abc_4108_n676) );
  INVX1 INVX1_240 ( .A(bus_sync_axi_bus_reg_data1_0_), .Y(bus_sync_axi_bus__abc_3782_n457) );
  INVX1 INVX1_241 ( .A(RST), .Y(bus_sync_axi_bus__abc_3782_n460) );
  INVX1 INVX1_242 ( .A(bus_sync_axi_bus_EECLK1), .Y(bus_sync_axi_bus__abc_3782_n461) );
  INVX1 INVX1_243 ( .A(CLK), .Y(bus_sync_axi_bus_NCLK2) );
  INVX1 INVX1_244 ( .A(bus_sync_rdata_reg_data1_0_), .Y(bus_sync_rdata__abc_3590_n201_1) );
  INVX1 INVX1_245 ( .A(RST), .Y(bus_sync_rdata__abc_3590_n204_1) );
  INVX1 INVX1_246 ( .A(bus_sync_rdata_EECLK2), .Y(bus_sync_rdata__abc_3590_n205_1) );
  INVX1 INVX1_247 ( .A(CLK), .Y(bus_sync_rdata_NCLK1) );
  INVX1 INVX1_248 ( .A(bus_sync_state_machine_reg_data1_0_), .Y(bus_sync_state_machine__abc_3756_n37) );
  INVX1 INVX1_249 ( .A(RST), .Y(bus_sync_state_machine__abc_3756_n40) );
  INVX1 INVX1_25 ( .A(counter_9_), .Y(_abc_4108_n677_1) );
  INVX1 INVX1_250 ( .A(bus_sync_state_machine_EECLK1), .Y(bus_sync_state_machine__abc_3756_n41) );
  INVX1 INVX1_251 ( .A(CLK), .Y(bus_sync_state_machine_NCLK2) );
  INVX1 INVX1_252 ( .A(bus_sync_status_reg_data1_0_), .Y(bus_sync_status__abc_3569_n30) );
  INVX1 INVX1_253 ( .A(RST), .Y(bus_sync_status__abc_3569_n33) );
  INVX1 INVX1_254 ( .A(bus_sync_status_EECLK2), .Y(bus_sync_status__abc_3569_n34) );
  INVX1 INVX1_255 ( .A(CLK), .Y(bus_sync_status_NCLK1) );
  INVX1 INVX1_26 ( .A(bus_cap_3_), .Y(_abc_4108_n686_1) );
  INVX1 INVX1_27 ( .A(bus_cap_4_), .Y(_abc_4108_n692) );
  INVX1 INVX1_28 ( .A(bus_cap_5_), .Y(_abc_4108_n698_1) );
  INVX1 INVX1_29 ( .A(bus_cap_6_), .Y(_abc_4108_n704) );
  INVX1 INVX1_3 ( .A(axi_awready), .Y(_abc_4108_n575) );
  INVX1 INVX1_30 ( .A(bus_cap_7_), .Y(_abc_4108_n710_1) );
  INVX1 INVX1_31 ( .A(bus_cap_8_), .Y(_abc_4108_n716) );
  INVX1 INVX1_32 ( .A(bus_cap_9_), .Y(_abc_4108_n722_1) );
  INVX1 INVX1_33 ( .A(bus_cap_10_), .Y(_abc_4108_n728) );
  INVX1 INVX1_34 ( .A(bus_cap_11_), .Y(_abc_4108_n734_1) );
  INVX1 INVX1_35 ( .A(bus_cap_12_), .Y(_abc_4108_n740) );
  INVX1 INVX1_36 ( .A(bus_cap_13_), .Y(_abc_4108_n746_1) );
  INVX1 INVX1_37 ( .A(bus_cap_14_), .Y(_abc_4108_n752) );
  INVX1 INVX1_38 ( .A(bus_cap_15_), .Y(_abc_4108_n758) );
  INVX1 INVX1_39 ( .A(bus_cap_16_), .Y(_abc_4108_n764) );
  INVX1 INVX1_4 ( .A(axi_rready), .Y(_abc_4108_n579_1) );
  INVX1 INVX1_40 ( .A(bus_cap_17_), .Y(_abc_4108_n770) );
  INVX1 INVX1_41 ( .A(bus_cap_18_), .Y(_abc_4108_n776) );
  INVX1 INVX1_42 ( .A(bus_cap_19_), .Y(_abc_4108_n782) );
  INVX1 INVX1_43 ( .A(bus_cap_20_), .Y(_abc_4108_n788) );
  INVX1 INVX1_44 ( .A(bus_cap_21_), .Y(_abc_4108_n794) );
  INVX1 INVX1_45 ( .A(bus_cap_22_), .Y(_abc_4108_n800) );
  INVX1 INVX1_46 ( .A(bus_cap_23_), .Y(_abc_4108_n806) );
  INVX1 INVX1_47 ( .A(bus_cap_24_), .Y(_abc_4108_n812) );
  INVX1 INVX1_48 ( .A(bus_cap_25_), .Y(_abc_4108_n818) );
  INVX1 INVX1_49 ( .A(bus_cap_26_), .Y(_abc_4108_n824_1) );
  INVX1 INVX1_5 ( .A(fini_spi_clk), .Y(_abc_4108_n583_1) );
  INVX1 INVX1_50 ( .A(bus_cap_27_), .Y(_abc_4108_n830) );
  INVX1 INVX1_51 ( .A(bus_cap_28_), .Y(_abc_4108_n836) );
  INVX1 INVX1_52 ( .A(bus_cap_29_), .Y(_abc_4108_n842) );
  INVX1 INVX1_53 ( .A(bus_cap_30_), .Y(_abc_4108_n848) );
  INVX1 INVX1_54 ( .A(DOUT), .Y(_abc_4108_n854) );
  INVX1 INVX1_55 ( .A(bus_sync_rdata_data_in_0_), .Y(_abc_4108_n858) );
  INVX1 INVX1_56 ( .A(bus_sync_rdata_data_in_1_), .Y(_abc_4108_n861_1) );
  INVX1 INVX1_57 ( .A(bus_sync_rdata_data_in_2_), .Y(_abc_4108_n864) );
  INVX1 INVX1_58 ( .A(bus_sync_rdata_data_in_3_), .Y(_abc_4108_n867_1) );
  INVX1 INVX1_59 ( .A(bus_sync_rdata_data_in_4_), .Y(_abc_4108_n870) );
  INVX1 INVX1_6 ( .A(axi_bready), .Y(_abc_4108_n586) );
  INVX1 INVX1_60 ( .A(bus_sync_rdata_data_in_5_), .Y(_abc_4108_n873_1) );
  INVX1 INVX1_61 ( .A(bus_sync_rdata_data_in_6_), .Y(_abc_4108_n876) );
  INVX1 INVX1_62 ( .A(bus_sync_rdata_data_in_7_), .Y(_abc_4108_n879_1) );
  INVX1 INVX1_63 ( .A(bus_sync_rdata_data_in_8_), .Y(_abc_4108_n882) );
  INVX1 INVX1_64 ( .A(bus_sync_rdata_data_in_9_), .Y(_abc_4108_n885_1) );
  INVX1 INVX1_65 ( .A(bus_sync_rdata_data_in_10_), .Y(_abc_4108_n888) );
  INVX1 INVX1_66 ( .A(bus_sync_rdata_data_in_11_), .Y(_abc_4108_n891_1) );
  INVX1 INVX1_67 ( .A(bus_sync_rdata_data_in_12_), .Y(_abc_4108_n894_1) );
  INVX1 INVX1_68 ( .A(bus_sync_rdata_data_in_13_), .Y(_abc_4108_n897_1) );
  INVX1 INVX1_69 ( .A(bus_sync_rdata_data_in_14_), .Y(_abc_4108_n900_1) );
  INVX1 INVX1_7 ( .A(axi_arready), .Y(_abc_4108_n590) );
  INVX1 INVX1_70 ( .A(bus_sync_rdata_data_in_15_), .Y(_abc_4108_n903_1) );
  INVX1 INVX1_71 ( .A(bus_sync_rdata_data_in_16_), .Y(_abc_4108_n906_1) );
  INVX1 INVX1_72 ( .A(bus_sync_rdata_data_in_17_), .Y(_abc_4108_n909_1) );
  INVX1 INVX1_73 ( .A(bus_sync_rdata_data_in_18_), .Y(_abc_4108_n912_1) );
  INVX1 INVX1_74 ( .A(bus_sync_rdata_data_in_19_), .Y(_abc_4108_n915_1) );
  INVX1 INVX1_75 ( .A(bus_sync_rdata_data_in_20_), .Y(_abc_4108_n918_1) );
  INVX1 INVX1_76 ( .A(bus_sync_rdata_data_in_21_), .Y(_abc_4108_n921_1) );
  INVX1 INVX1_77 ( .A(bus_sync_rdata_data_in_22_), .Y(_abc_4108_n924_1) );
  INVX1 INVX1_78 ( .A(bus_sync_rdata_data_in_23_), .Y(_abc_4108_n927_1) );
  INVX1 INVX1_79 ( .A(bus_sync_rdata_data_in_24_), .Y(_abc_4108_n930_1) );
  INVX1 INVX1_8 ( .A(we), .Y(_abc_4108_n595) );
  INVX1 INVX1_80 ( .A(bus_sync_rdata_data_in_25_), .Y(_abc_4108_n933_1) );
  INVX1 INVX1_81 ( .A(bus_sync_rdata_data_in_26_), .Y(_abc_4108_n936_1) );
  INVX1 INVX1_82 ( .A(bus_sync_rdata_data_in_27_), .Y(_abc_4108_n939_1) );
  INVX1 INVX1_83 ( .A(bus_sync_rdata_data_in_28_), .Y(_abc_4108_n942_1) );
  INVX1 INVX1_84 ( .A(bus_sync_rdata_data_in_29_), .Y(_abc_4108_n945_1) );
  INVX1 INVX1_85 ( .A(bus_sync_rdata_data_in_30_), .Y(_abc_4108_n948_1) );
  INVX1 INVX1_86 ( .A(bus_sync_rdata_data_in_31_), .Y(_abc_4108_n951_1) );
  INVX1 INVX1_87 ( .A(WDATA_0_), .Y(_abc_4108_n954) );
  INVX1 INVX1_88 ( .A(CEB), .Y(_abc_4108_n955_1) );
  INVX1 INVX1_89 ( .A(WDATA_1_), .Y(_abc_4108_n959) );
  INVX1 INVX1_9 ( .A(counter_1_), .Y(_abc_4108_n596) );
  INVX1 INVX1_90 ( .A(WDATA_2_), .Y(_abc_4108_n962) );
  INVX1 INVX1_91 ( .A(WDATA_3_), .Y(_abc_4108_n965) );
  INVX1 INVX1_92 ( .A(WDATA_4_), .Y(_abc_4108_n968_1) );
  INVX1 INVX1_93 ( .A(WDATA_5_), .Y(_abc_4108_n971) );
  INVX1 INVX1_94 ( .A(WDATA_6_), .Y(_abc_4108_n974) );
  INVX1 INVX1_95 ( .A(WDATA_7_), .Y(_abc_4108_n977) );
  INVX1 INVX1_96 ( .A(WDATA_8_), .Y(_abc_4108_n980) );
  INVX1 INVX1_97 ( .A(WDATA_9_), .Y(_abc_4108_n983) );
  INVX1 INVX1_98 ( .A(WDATA_10_), .Y(_abc_4108_n986) );
  INVX1 INVX1_99 ( .A(WDATA_11_), .Y(_abc_4108_n989) );
  MUX2X1 MUX2X1_1 ( .A(bus_cap_1_), .B(bus_cap_0_), .S(_abc_4108_n638_1), .Y(_abc_4108_n646_1) );
  NAND2X1 NAND2X1_1 ( .A(RST), .B(state_7_), .Y(_abc_4108_n558_1) );
  NAND2X1 NAND2X1_10 ( .A(DATA), .B(_abc_4108_n597_1), .Y(_abc_4108_n598_1) );
  NAND2X1 NAND2X1_100 ( .A(bus_sync_axi_bus_reg_data2_9_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n486) );
  NAND2X1 NAND2X1_101 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_9_), .Y(bus_sync_axi_bus__abc_3782_n487) );
  NAND2X1 NAND2X1_102 ( .A(bus_sync_axi_bus_reg_data2_10_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n489) );
  NAND2X1 NAND2X1_103 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_10_), .Y(bus_sync_axi_bus__abc_3782_n490) );
  NAND2X1 NAND2X1_104 ( .A(bus_sync_axi_bus_reg_data2_11_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n492) );
  NAND2X1 NAND2X1_105 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_11_), .Y(bus_sync_axi_bus__abc_3782_n493) );
  NAND2X1 NAND2X1_106 ( .A(bus_sync_axi_bus_reg_data2_12_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n495) );
  NAND2X1 NAND2X1_107 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_12_), .Y(bus_sync_axi_bus__abc_3782_n496) );
  NAND2X1 NAND2X1_108 ( .A(bus_sync_axi_bus_reg_data2_13_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n498) );
  NAND2X1 NAND2X1_109 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_13_), .Y(bus_sync_axi_bus__abc_3782_n499) );
  NAND2X1 NAND2X1_11 ( .A(re), .B(we), .Y(_abc_4108_n603_1) );
  NAND2X1 NAND2X1_110 ( .A(bus_sync_axi_bus_reg_data2_14_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n501) );
  NAND2X1 NAND2X1_111 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_14_), .Y(bus_sync_axi_bus__abc_3782_n502) );
  NAND2X1 NAND2X1_112 ( .A(bus_sync_axi_bus_reg_data2_15_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n504) );
  NAND2X1 NAND2X1_113 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_15_), .Y(bus_sync_axi_bus__abc_3782_n505) );
  NAND2X1 NAND2X1_114 ( .A(bus_sync_axi_bus_reg_data2_16_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n507) );
  NAND2X1 NAND2X1_115 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_16_), .Y(bus_sync_axi_bus__abc_3782_n508) );
  NAND2X1 NAND2X1_116 ( .A(bus_sync_axi_bus_reg_data2_17_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n510) );
  NAND2X1 NAND2X1_117 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_17_), .Y(bus_sync_axi_bus__abc_3782_n511) );
  NAND2X1 NAND2X1_118 ( .A(bus_sync_axi_bus_reg_data2_18_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n513) );
  NAND2X1 NAND2X1_119 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_18_), .Y(bus_sync_axi_bus__abc_3782_n514) );
  NAND2X1 NAND2X1_12 ( .A(_abc_4108_n603_1), .B(_abc_4108_n602_1), .Y(_abc_4108_n604_1) );
  NAND2X1 NAND2X1_120 ( .A(bus_sync_axi_bus_reg_data2_19_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n516) );
  NAND2X1 NAND2X1_121 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_19_), .Y(bus_sync_axi_bus__abc_3782_n517) );
  NAND2X1 NAND2X1_122 ( .A(bus_sync_axi_bus_reg_data2_20_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n519) );
  NAND2X1 NAND2X1_123 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_20_), .Y(bus_sync_axi_bus__abc_3782_n520) );
  NAND2X1 NAND2X1_124 ( .A(bus_sync_axi_bus_reg_data2_21_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n522) );
  NAND2X1 NAND2X1_125 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_21_), .Y(bus_sync_axi_bus__abc_3782_n523) );
  NAND2X1 NAND2X1_126 ( .A(bus_sync_axi_bus_reg_data2_22_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n525) );
  NAND2X1 NAND2X1_127 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_22_), .Y(bus_sync_axi_bus__abc_3782_n526) );
  NAND2X1 NAND2X1_128 ( .A(bus_sync_axi_bus_reg_data2_23_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n528) );
  NAND2X1 NAND2X1_129 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_23_), .Y(bus_sync_axi_bus__abc_3782_n529) );
  NAND2X1 NAND2X1_13 ( .A(_abc_4108_n605), .B(_abc_4108_n606), .Y(_abc_4108_n607_1) );
  NAND2X1 NAND2X1_130 ( .A(bus_sync_axi_bus_reg_data2_24_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n531) );
  NAND2X1 NAND2X1_131 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_24_), .Y(bus_sync_axi_bus__abc_3782_n532) );
  NAND2X1 NAND2X1_132 ( .A(bus_sync_axi_bus_reg_data2_25_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n534) );
  NAND2X1 NAND2X1_133 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_25_), .Y(bus_sync_axi_bus__abc_3782_n535) );
  NAND2X1 NAND2X1_134 ( .A(bus_sync_axi_bus_reg_data2_26_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n537) );
  NAND2X1 NAND2X1_135 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_26_), .Y(bus_sync_axi_bus__abc_3782_n538) );
  NAND2X1 NAND2X1_136 ( .A(bus_sync_axi_bus_reg_data2_27_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n540) );
  NAND2X1 NAND2X1_137 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_27_), .Y(bus_sync_axi_bus__abc_3782_n541) );
  NAND2X1 NAND2X1_138 ( .A(bus_sync_axi_bus_reg_data2_28_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n543) );
  NAND2X1 NAND2X1_139 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_28_), .Y(bus_sync_axi_bus__abc_3782_n544) );
  NAND2X1 NAND2X1_14 ( .A(_abc_4108_n608_1), .B(_abc_4108_n609_1), .Y(_abc_4108_n610) );
  NAND2X1 NAND2X1_140 ( .A(bus_sync_axi_bus_reg_data2_29_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n546) );
  NAND2X1 NAND2X1_141 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_29_), .Y(bus_sync_axi_bus__abc_3782_n547) );
  NAND2X1 NAND2X1_142 ( .A(bus_sync_axi_bus_reg_data2_30_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n549) );
  NAND2X1 NAND2X1_143 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_30_), .Y(bus_sync_axi_bus__abc_3782_n550) );
  NAND2X1 NAND2X1_144 ( .A(bus_sync_axi_bus_reg_data2_31_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n552) );
  NAND2X1 NAND2X1_145 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_31_), .Y(bus_sync_axi_bus__abc_3782_n553) );
  NAND2X1 NAND2X1_146 ( .A(bus_sync_axi_bus_reg_data2_32_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n555) );
  NAND2X1 NAND2X1_147 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_32_), .Y(bus_sync_axi_bus__abc_3782_n556) );
  NAND2X1 NAND2X1_148 ( .A(bus_sync_axi_bus_reg_data2_33_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n558) );
  NAND2X1 NAND2X1_149 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_33_), .Y(bus_sync_axi_bus__abc_3782_n559) );
  NAND2X1 NAND2X1_15 ( .A(_abc_4108_n612_1), .B(_abc_4108_n613_1), .Y(_abc_4108_n614_1) );
  NAND2X1 NAND2X1_150 ( .A(bus_sync_axi_bus_reg_data2_34_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n561) );
  NAND2X1 NAND2X1_151 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_34_), .Y(bus_sync_axi_bus__abc_3782_n562) );
  NAND2X1 NAND2X1_152 ( .A(bus_sync_axi_bus_reg_data2_35_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n564) );
  NAND2X1 NAND2X1_153 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_35_), .Y(bus_sync_axi_bus__abc_3782_n565) );
  NAND2X1 NAND2X1_154 ( .A(bus_sync_axi_bus_reg_data2_36_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n567) );
  NAND2X1 NAND2X1_155 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_36_), .Y(bus_sync_axi_bus__abc_3782_n568) );
  NAND2X1 NAND2X1_156 ( .A(bus_sync_axi_bus_reg_data2_37_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n570) );
  NAND2X1 NAND2X1_157 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_37_), .Y(bus_sync_axi_bus__abc_3782_n571) );
  NAND2X1 NAND2X1_158 ( .A(bus_sync_axi_bus_reg_data2_38_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n573) );
  NAND2X1 NAND2X1_159 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_38_), .Y(bus_sync_axi_bus__abc_3782_n574) );
  NAND2X1 NAND2X1_16 ( .A(_abc_4108_n611), .B(_abc_4108_n619_1), .Y(_abc_4108_n620) );
  NAND2X1 NAND2X1_160 ( .A(bus_sync_axi_bus_reg_data2_39_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n576) );
  NAND2X1 NAND2X1_161 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_39_), .Y(bus_sync_axi_bus__abc_3782_n577) );
  NAND2X1 NAND2X1_162 ( .A(bus_sync_axi_bus_reg_data2_40_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n579) );
  NAND2X1 NAND2X1_163 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_40_), .Y(bus_sync_axi_bus__abc_3782_n580) );
  NAND2X1 NAND2X1_164 ( .A(bus_sync_axi_bus_reg_data2_41_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n582) );
  NAND2X1 NAND2X1_165 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_41_), .Y(bus_sync_axi_bus__abc_3782_n583) );
  NAND2X1 NAND2X1_166 ( .A(bus_sync_axi_bus_reg_data2_42_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n585) );
  NAND2X1 NAND2X1_167 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_42_), .Y(bus_sync_axi_bus__abc_3782_n586) );
  NAND2X1 NAND2X1_168 ( .A(bus_sync_axi_bus_reg_data2_43_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n588) );
  NAND2X1 NAND2X1_169 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_43_), .Y(bus_sync_axi_bus__abc_3782_n589) );
  NAND2X1 NAND2X1_17 ( .A(_abc_4108_n621), .B(_abc_4108_n622_1), .Y(_abc_4108_n623_1) );
  NAND2X1 NAND2X1_170 ( .A(bus_sync_axi_bus_reg_data2_44_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n591) );
  NAND2X1 NAND2X1_171 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_44_), .Y(bus_sync_axi_bus__abc_3782_n592) );
  NAND2X1 NAND2X1_172 ( .A(bus_sync_axi_bus_reg_data2_45_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n594) );
  NAND2X1 NAND2X1_173 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_45_), .Y(bus_sync_axi_bus__abc_3782_n595) );
  NAND2X1 NAND2X1_174 ( .A(bus_sync_axi_bus_reg_data2_46_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n597) );
  NAND2X1 NAND2X1_175 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_46_), .Y(bus_sync_axi_bus__abc_3782_n598) );
  NAND2X1 NAND2X1_176 ( .A(bus_sync_axi_bus_reg_data2_47_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n600) );
  NAND2X1 NAND2X1_177 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_47_), .Y(bus_sync_axi_bus__abc_3782_n601) );
  NAND2X1 NAND2X1_178 ( .A(bus_sync_axi_bus_reg_data2_48_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n603) );
  NAND2X1 NAND2X1_179 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_48_), .Y(bus_sync_axi_bus__abc_3782_n604) );
  NAND2X1 NAND2X1_18 ( .A(_abc_4108_n629), .B(_abc_4108_n630_1), .Y(_abc_4108_n631) );
  NAND2X1 NAND2X1_180 ( .A(bus_sync_axi_bus_reg_data2_49_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n606) );
  NAND2X1 NAND2X1_181 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_49_), .Y(bus_sync_axi_bus__abc_3782_n607) );
  NAND2X1 NAND2X1_182 ( .A(bus_sync_axi_bus_reg_data2_50_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n609) );
  NAND2X1 NAND2X1_183 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_50_), .Y(bus_sync_axi_bus__abc_3782_n610) );
  NAND2X1 NAND2X1_184 ( .A(bus_sync_axi_bus_reg_data2_51_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n612) );
  NAND2X1 NAND2X1_185 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_51_), .Y(bus_sync_axi_bus__abc_3782_n613) );
  NAND2X1 NAND2X1_186 ( .A(bus_sync_axi_bus_reg_data2_52_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n615) );
  NAND2X1 NAND2X1_187 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_52_), .Y(bus_sync_axi_bus__abc_3782_n616) );
  NAND2X1 NAND2X1_188 ( .A(bus_sync_axi_bus_reg_data2_53_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n618) );
  NAND2X1 NAND2X1_189 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_53_), .Y(bus_sync_axi_bus__abc_3782_n619) );
  NAND2X1 NAND2X1_19 ( .A(_abc_4108_n628), .B(_abc_4108_n636), .Y(_abc_4108_n637_1) );
  NAND2X1 NAND2X1_190 ( .A(bus_sync_axi_bus_reg_data2_54_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n621) );
  NAND2X1 NAND2X1_191 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_54_), .Y(bus_sync_axi_bus__abc_3782_n622) );
  NAND2X1 NAND2X1_192 ( .A(bus_sync_axi_bus_reg_data2_55_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n624) );
  NAND2X1 NAND2X1_193 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_55_), .Y(bus_sync_axi_bus__abc_3782_n625) );
  NAND2X1 NAND2X1_194 ( .A(bus_sync_axi_bus_reg_data2_56_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n627) );
  NAND2X1 NAND2X1_195 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_56_), .Y(bus_sync_axi_bus__abc_3782_n628) );
  NAND2X1 NAND2X1_196 ( .A(bus_sync_axi_bus_reg_data2_57_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n630) );
  NAND2X1 NAND2X1_197 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_57_), .Y(bus_sync_axi_bus__abc_3782_n631) );
  NAND2X1 NAND2X1_198 ( .A(bus_sync_axi_bus_reg_data2_58_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n633) );
  NAND2X1 NAND2X1_199 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_58_), .Y(bus_sync_axi_bus__abc_3782_n634) );
  NAND2X1 NAND2X1_2 ( .A(state_1_), .B(fini_spi_clk), .Y(_abc_4108_n565) );
  NAND2X1 NAND2X1_20 ( .A(bus_cap_0_), .B(_abc_4108_n638_1), .Y(_abc_4108_n639) );
  NAND2X1 NAND2X1_200 ( .A(bus_sync_axi_bus_reg_data2_59_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n636) );
  NAND2X1 NAND2X1_201 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_59_), .Y(bus_sync_axi_bus__abc_3782_n637) );
  NAND2X1 NAND2X1_202 ( .A(bus_sync_axi_bus_reg_data2_60_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n639) );
  NAND2X1 NAND2X1_203 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_60_), .Y(bus_sync_axi_bus__abc_3782_n640) );
  NAND2X1 NAND2X1_204 ( .A(bus_sync_axi_bus_reg_data2_61_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n642) );
  NAND2X1 NAND2X1_205 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_61_), .Y(bus_sync_axi_bus__abc_3782_n643) );
  NAND2X1 NAND2X1_206 ( .A(bus_sync_axi_bus_reg_data2_62_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n645) );
  NAND2X1 NAND2X1_207 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_62_), .Y(bus_sync_axi_bus__abc_3782_n646) );
  NAND2X1 NAND2X1_208 ( .A(bus_sync_axi_bus_reg_data2_63_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n648) );
  NAND2X1 NAND2X1_209 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_63_), .Y(bus_sync_axi_bus__abc_3782_n649) );
  NAND2X1 NAND2X1_21 ( .A(_abc_4108_n652), .B(_abc_4108_n638_1), .Y(_abc_4108_n653_1) );
  NAND2X1 NAND2X1_210 ( .A(bus_sync_rdata_reg_data2_1_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n206_1) );
  NAND2X1 NAND2X1_211 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_1_), .Y(bus_sync_rdata__abc_3590_n207_1) );
  NAND2X1 NAND2X1_212 ( .A(bus_sync_rdata_reg_data2_2_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n209_1) );
  NAND2X1 NAND2X1_213 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_2_), .Y(bus_sync_rdata__abc_3590_n210_1) );
  NAND2X1 NAND2X1_214 ( .A(bus_sync_rdata_reg_data2_3_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n212_1) );
  NAND2X1 NAND2X1_215 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_3_), .Y(bus_sync_rdata__abc_3590_n213_1) );
  NAND2X1 NAND2X1_216 ( .A(bus_sync_rdata_reg_data2_4_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n215_1) );
  NAND2X1 NAND2X1_217 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_4_), .Y(bus_sync_rdata__abc_3590_n216_1) );
  NAND2X1 NAND2X1_218 ( .A(bus_sync_rdata_reg_data2_5_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n218_1) );
  NAND2X1 NAND2X1_219 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_5_), .Y(bus_sync_rdata__abc_3590_n219_1) );
  NAND2X1 NAND2X1_22 ( .A(bus_sync_rdata_data_out_3_), .B(_abc_4108_n640), .Y(_abc_4108_n660) );
  NAND2X1 NAND2X1_220 ( .A(bus_sync_rdata_reg_data2_6_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n221_1) );
  NAND2X1 NAND2X1_221 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_6_), .Y(bus_sync_rdata__abc_3590_n222_1) );
  NAND2X1 NAND2X1_222 ( .A(bus_sync_rdata_reg_data2_7_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n224_1) );
  NAND2X1 NAND2X1_223 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_7_), .Y(bus_sync_rdata__abc_3590_n225_1) );
  NAND2X1 NAND2X1_224 ( .A(bus_sync_rdata_reg_data2_8_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n227_1) );
  NAND2X1 NAND2X1_225 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_8_), .Y(bus_sync_rdata__abc_3590_n228_1) );
  NAND2X1 NAND2X1_226 ( .A(bus_sync_rdata_reg_data2_9_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n230_1) );
  NAND2X1 NAND2X1_227 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_9_), .Y(bus_sync_rdata__abc_3590_n231_1) );
  NAND2X1 NAND2X1_228 ( .A(bus_sync_rdata_reg_data2_10_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n233) );
  NAND2X1 NAND2X1_229 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_10_), .Y(bus_sync_rdata__abc_3590_n234) );
  NAND2X1 NAND2X1_23 ( .A(_abc_4108_n676), .B(_abc_4108_n677_1), .Y(_abc_4108_n678_1) );
  NAND2X1 NAND2X1_230 ( .A(bus_sync_rdata_reg_data2_11_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n236) );
  NAND2X1 NAND2X1_231 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_11_), .Y(bus_sync_rdata__abc_3590_n237) );
  NAND2X1 NAND2X1_232 ( .A(bus_sync_rdata_reg_data2_12_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n239) );
  NAND2X1 NAND2X1_233 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_12_), .Y(bus_sync_rdata__abc_3590_n240) );
  NAND2X1 NAND2X1_234 ( .A(bus_sync_rdata_reg_data2_13_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n242) );
  NAND2X1 NAND2X1_235 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_13_), .Y(bus_sync_rdata__abc_3590_n243) );
  NAND2X1 NAND2X1_236 ( .A(bus_sync_rdata_reg_data2_14_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n245) );
  NAND2X1 NAND2X1_237 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_14_), .Y(bus_sync_rdata__abc_3590_n246) );
  NAND2X1 NAND2X1_238 ( .A(bus_sync_rdata_reg_data2_15_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n248) );
  NAND2X1 NAND2X1_239 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_15_), .Y(bus_sync_rdata__abc_3590_n249) );
  NAND2X1 NAND2X1_24 ( .A(_abc_4108_n686_1), .B(_abc_4108_n638_1), .Y(_abc_4108_n687) );
  NAND2X1 NAND2X1_240 ( .A(bus_sync_rdata_reg_data2_16_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n251) );
  NAND2X1 NAND2X1_241 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_16_), .Y(bus_sync_rdata__abc_3590_n252) );
  NAND2X1 NAND2X1_242 ( .A(bus_sync_rdata_reg_data2_17_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n254) );
  NAND2X1 NAND2X1_243 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_17_), .Y(bus_sync_rdata__abc_3590_n255) );
  NAND2X1 NAND2X1_244 ( .A(bus_sync_rdata_reg_data2_18_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n257) );
  NAND2X1 NAND2X1_245 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_18_), .Y(bus_sync_rdata__abc_3590_n258) );
  NAND2X1 NAND2X1_246 ( .A(bus_sync_rdata_reg_data2_19_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n260) );
  NAND2X1 NAND2X1_247 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_19_), .Y(bus_sync_rdata__abc_3590_n261) );
  NAND2X1 NAND2X1_248 ( .A(bus_sync_rdata_reg_data2_20_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n263) );
  NAND2X1 NAND2X1_249 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_20_), .Y(bus_sync_rdata__abc_3590_n264) );
  NAND2X1 NAND2X1_25 ( .A(bus_sync_rdata_data_out_4_), .B(_abc_4108_n640), .Y(_abc_4108_n690_1) );
  NAND2X1 NAND2X1_250 ( .A(bus_sync_rdata_reg_data2_21_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n266) );
  NAND2X1 NAND2X1_251 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_21_), .Y(bus_sync_rdata__abc_3590_n267) );
  NAND2X1 NAND2X1_252 ( .A(bus_sync_rdata_reg_data2_22_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n269) );
  NAND2X1 NAND2X1_253 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_22_), .Y(bus_sync_rdata__abc_3590_n270) );
  NAND2X1 NAND2X1_254 ( .A(bus_sync_rdata_reg_data2_23_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n272) );
  NAND2X1 NAND2X1_255 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_23_), .Y(bus_sync_rdata__abc_3590_n273) );
  NAND2X1 NAND2X1_256 ( .A(bus_sync_rdata_reg_data2_24_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n275) );
  NAND2X1 NAND2X1_257 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_24_), .Y(bus_sync_rdata__abc_3590_n276) );
  NAND2X1 NAND2X1_258 ( .A(bus_sync_rdata_reg_data2_25_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n278) );
  NAND2X1 NAND2X1_259 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_25_), .Y(bus_sync_rdata__abc_3590_n279) );
  NAND2X1 NAND2X1_26 ( .A(_abc_4108_n692), .B(_abc_4108_n638_1), .Y(_abc_4108_n693_1) );
  NAND2X1 NAND2X1_260 ( .A(bus_sync_rdata_reg_data2_26_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n281) );
  NAND2X1 NAND2X1_261 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_26_), .Y(bus_sync_rdata__abc_3590_n282) );
  NAND2X1 NAND2X1_262 ( .A(bus_sync_rdata_reg_data2_27_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n284) );
  NAND2X1 NAND2X1_263 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_27_), .Y(bus_sync_rdata__abc_3590_n285) );
  NAND2X1 NAND2X1_264 ( .A(bus_sync_rdata_reg_data2_28_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n287) );
  NAND2X1 NAND2X1_265 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_28_), .Y(bus_sync_rdata__abc_3590_n288) );
  NAND2X1 NAND2X1_266 ( .A(bus_sync_rdata_reg_data2_29_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n290) );
  NAND2X1 NAND2X1_267 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_29_), .Y(bus_sync_rdata__abc_3590_n291) );
  NAND2X1 NAND2X1_268 ( .A(bus_sync_rdata_reg_data2_30_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n293) );
  NAND2X1 NAND2X1_269 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_30_), .Y(bus_sync_rdata__abc_3590_n294) );
  NAND2X1 NAND2X1_27 ( .A(bus_sync_rdata_data_out_5_), .B(_abc_4108_n640), .Y(_abc_4108_n696) );
  NAND2X1 NAND2X1_270 ( .A(bus_sync_rdata_reg_data2_31_), .B(bus_sync_rdata__abc_3590_n205_1), .Y(bus_sync_rdata__abc_3590_n296) );
  NAND2X1 NAND2X1_271 ( .A(bus_sync_rdata_EECLK2), .B(bus_sync_rdata_reg_data1_31_), .Y(bus_sync_rdata__abc_3590_n297) );
  NAND2X1 NAND2X1_272 ( .A(bus_sync_state_machine_reg_data2_1_), .B(bus_sync_state_machine__abc_3756_n41), .Y(bus_sync_state_machine__abc_3756_n42) );
  NAND2X1 NAND2X1_273 ( .A(bus_sync_state_machine_EECLK1), .B(bus_sync_state_machine_reg_data1_1_), .Y(bus_sync_state_machine__abc_3756_n43) );
  NAND2X1 NAND2X1_274 ( .A(bus_sync_state_machine_reg_data2_2_), .B(bus_sync_state_machine__abc_3756_n41), .Y(bus_sync_state_machine__abc_3756_n45) );
  NAND2X1 NAND2X1_275 ( .A(bus_sync_state_machine_EECLK1), .B(bus_sync_state_machine_reg_data1_2_), .Y(bus_sync_state_machine__abc_3756_n46) );
  NAND2X1 NAND2X1_276 ( .A(bus_sync_state_machine_reg_data2_3_), .B(bus_sync_state_machine__abc_3756_n41), .Y(bus_sync_state_machine__abc_3756_n48) );
  NAND2X1 NAND2X1_277 ( .A(bus_sync_state_machine_EECLK1), .B(bus_sync_state_machine_reg_data1_3_), .Y(bus_sync_state_machine__abc_3756_n49) );
  NAND2X1 NAND2X1_278 ( .A(bus_sync_status_reg_data2_1_), .B(bus_sync_status__abc_3569_n34), .Y(bus_sync_status__abc_3569_n35) );
  NAND2X1 NAND2X1_279 ( .A(bus_sync_status_EECLK2), .B(bus_sync_status_reg_data1_1_), .Y(bus_sync_status__abc_3569_n36) );
  NAND2X1 NAND2X1_28 ( .A(_abc_4108_n698_1), .B(_abc_4108_n638_1), .Y(_abc_4108_n699) );
  NAND2X1 NAND2X1_280 ( .A(bus_sync_status_reg_data2_2_), .B(bus_sync_status__abc_3569_n34), .Y(bus_sync_status__abc_3569_n38) );
  NAND2X1 NAND2X1_281 ( .A(bus_sync_status_EECLK2), .B(bus_sync_status_reg_data1_2_), .Y(bus_sync_status__abc_3569_n39) );
  NAND2X1 NAND2X1_29 ( .A(bus_sync_rdata_data_out_6_), .B(_abc_4108_n640), .Y(_abc_4108_n702_1) );
  NAND2X1 NAND2X1_3 ( .A(RST), .B(state_6_), .Y(_abc_4108_n568_1) );
  NAND2X1 NAND2X1_30 ( .A(_abc_4108_n704), .B(_abc_4108_n638_1), .Y(_abc_4108_n705_1) );
  NAND2X1 NAND2X1_31 ( .A(bus_sync_rdata_data_out_7_), .B(_abc_4108_n640), .Y(_abc_4108_n708) );
  NAND2X1 NAND2X1_32 ( .A(_abc_4108_n710_1), .B(_abc_4108_n638_1), .Y(_abc_4108_n711) );
  NAND2X1 NAND2X1_33 ( .A(bus_sync_rdata_data_out_8_), .B(_abc_4108_n640), .Y(_abc_4108_n714_1) );
  NAND2X1 NAND2X1_34 ( .A(_abc_4108_n716), .B(_abc_4108_n638_1), .Y(_abc_4108_n717_1) );
  NAND2X1 NAND2X1_35 ( .A(bus_sync_rdata_data_out_9_), .B(_abc_4108_n640), .Y(_abc_4108_n720) );
  NAND2X1 NAND2X1_36 ( .A(_abc_4108_n722_1), .B(_abc_4108_n638_1), .Y(_abc_4108_n723) );
  NAND2X1 NAND2X1_37 ( .A(bus_sync_rdata_data_out_10_), .B(_abc_4108_n640), .Y(_abc_4108_n726_1) );
  NAND2X1 NAND2X1_38 ( .A(_abc_4108_n728), .B(_abc_4108_n638_1), .Y(_abc_4108_n729_1) );
  NAND2X1 NAND2X1_39 ( .A(bus_sync_rdata_data_out_11_), .B(_abc_4108_n640), .Y(_abc_4108_n732) );
  NAND2X1 NAND2X1_4 ( .A(fini_spi_clk), .B(we_clk), .Y(_abc_4108_n569_1) );
  NAND2X1 NAND2X1_40 ( .A(_abc_4108_n734_1), .B(_abc_4108_n638_1), .Y(_abc_4108_n735) );
  NAND2X1 NAND2X1_41 ( .A(bus_sync_rdata_data_out_12_), .B(_abc_4108_n640), .Y(_abc_4108_n738_1) );
  NAND2X1 NAND2X1_42 ( .A(_abc_4108_n740), .B(_abc_4108_n638_1), .Y(_abc_4108_n741_1) );
  NAND2X1 NAND2X1_43 ( .A(bus_sync_rdata_data_out_13_), .B(_abc_4108_n640), .Y(_abc_4108_n744) );
  NAND2X1 NAND2X1_44 ( .A(_abc_4108_n746_1), .B(_abc_4108_n638_1), .Y(_abc_4108_n747) );
  NAND2X1 NAND2X1_45 ( .A(bus_sync_rdata_data_out_14_), .B(_abc_4108_n640), .Y(_abc_4108_n750_1) );
  NAND2X1 NAND2X1_46 ( .A(_abc_4108_n752), .B(_abc_4108_n638_1), .Y(_abc_4108_n753_1) );
  NAND2X1 NAND2X1_47 ( .A(bus_sync_rdata_data_out_15_), .B(_abc_4108_n640), .Y(_abc_4108_n756) );
  NAND2X1 NAND2X1_48 ( .A(_abc_4108_n758), .B(_abc_4108_n638_1), .Y(_abc_4108_n759_1) );
  NAND2X1 NAND2X1_49 ( .A(bus_sync_rdata_data_out_16_), .B(_abc_4108_n640), .Y(_abc_4108_n762) );
  NAND2X1 NAND2X1_5 ( .A(fini_spi_clk), .B(re_clk), .Y(_abc_4108_n571) );
  NAND2X1 NAND2X1_50 ( .A(_abc_4108_n764), .B(_abc_4108_n638_1), .Y(_abc_4108_n765_1) );
  NAND2X1 NAND2X1_51 ( .A(bus_sync_rdata_data_out_17_), .B(_abc_4108_n640), .Y(_abc_4108_n768) );
  NAND2X1 NAND2X1_52 ( .A(_abc_4108_n770), .B(_abc_4108_n638_1), .Y(_abc_4108_n771_1) );
  NAND2X1 NAND2X1_53 ( .A(bus_sync_rdata_data_out_18_), .B(_abc_4108_n640), .Y(_abc_4108_n774) );
  NAND2X1 NAND2X1_54 ( .A(_abc_4108_n776), .B(_abc_4108_n638_1), .Y(_abc_4108_n777_1) );
  NAND2X1 NAND2X1_55 ( .A(bus_sync_rdata_data_out_19_), .B(_abc_4108_n640), .Y(_abc_4108_n780) );
  NAND2X1 NAND2X1_56 ( .A(_abc_4108_n782), .B(_abc_4108_n638_1), .Y(_abc_4108_n783_1) );
  NAND2X1 NAND2X1_57 ( .A(bus_sync_rdata_data_out_20_), .B(_abc_4108_n640), .Y(_abc_4108_n786) );
  NAND2X1 NAND2X1_58 ( .A(_abc_4108_n788), .B(_abc_4108_n638_1), .Y(_abc_4108_n789_1) );
  NAND2X1 NAND2X1_59 ( .A(bus_sync_rdata_data_out_21_), .B(_abc_4108_n640), .Y(_abc_4108_n792) );
  NAND2X1 NAND2X1_6 ( .A(state_0_), .B(_abc_4108_n572_1), .Y(_abc_4108_n573_1) );
  NAND2X1 NAND2X1_60 ( .A(_abc_4108_n794), .B(_abc_4108_n638_1), .Y(_abc_4108_n795_1) );
  NAND2X1 NAND2X1_61 ( .A(bus_sync_rdata_data_out_22_), .B(_abc_4108_n640), .Y(_abc_4108_n798) );
  NAND2X1 NAND2X1_62 ( .A(_abc_4108_n800), .B(_abc_4108_n638_1), .Y(_abc_4108_n801_1) );
  NAND2X1 NAND2X1_63 ( .A(bus_sync_rdata_data_out_23_), .B(_abc_4108_n640), .Y(_abc_4108_n804) );
  NAND2X1 NAND2X1_64 ( .A(_abc_4108_n806), .B(_abc_4108_n638_1), .Y(_abc_4108_n807_1) );
  NAND2X1 NAND2X1_65 ( .A(bus_sync_rdata_data_out_24_), .B(_abc_4108_n640), .Y(_abc_4108_n810) );
  NAND2X1 NAND2X1_66 ( .A(_abc_4108_n812), .B(_abc_4108_n638_1), .Y(_abc_4108_n813_1) );
  NAND2X1 NAND2X1_67 ( .A(bus_sync_rdata_data_out_25_), .B(_abc_4108_n640), .Y(_abc_4108_n816) );
  NAND2X1 NAND2X1_68 ( .A(_abc_4108_n818), .B(_abc_4108_n638_1), .Y(_abc_4108_n819_1) );
  NAND2X1 NAND2X1_69 ( .A(bus_sync_rdata_data_out_26_), .B(_abc_4108_n640), .Y(_abc_4108_n822) );
  NAND2X1 NAND2X1_7 ( .A(_abc_4108_n579_1), .B(_abc_4108_n580), .Y(axi_arvalid) );
  NAND2X1 NAND2X1_70 ( .A(_abc_4108_n824_1), .B(_abc_4108_n638_1), .Y(_abc_4108_n825_1) );
  NAND2X1 NAND2X1_71 ( .A(bus_sync_rdata_data_out_27_), .B(_abc_4108_n640), .Y(_abc_4108_n828) );
  NAND2X1 NAND2X1_72 ( .A(_abc_4108_n830), .B(_abc_4108_n638_1), .Y(_abc_4108_n831_1) );
  NAND2X1 NAND2X1_73 ( .A(bus_sync_rdata_data_out_28_), .B(_abc_4108_n640), .Y(_abc_4108_n834) );
  NAND2X1 NAND2X1_74 ( .A(_abc_4108_n836), .B(_abc_4108_n638_1), .Y(_abc_4108_n837_1) );
  NAND2X1 NAND2X1_75 ( .A(bus_sync_rdata_data_out_29_), .B(_abc_4108_n640), .Y(_abc_4108_n840) );
  NAND2X1 NAND2X1_76 ( .A(_abc_4108_n842), .B(_abc_4108_n638_1), .Y(_abc_4108_n843_1) );
  NAND2X1 NAND2X1_77 ( .A(bus_sync_rdata_data_out_30_), .B(_abc_4108_n640), .Y(_abc_4108_n846) );
  NAND2X1 NAND2X1_78 ( .A(_abc_4108_n848), .B(_abc_4108_n638_1), .Y(_abc_4108_n849_1) );
  NAND2X1 NAND2X1_79 ( .A(bus_sync_rdata_data_out_31_), .B(_abc_4108_n640), .Y(_abc_4108_n852) );
  NAND2X1 NAND2X1_8 ( .A(_abc_4108_n586), .B(_abc_4108_n587_1), .Y(axi_wvalid) );
  NAND2X1 NAND2X1_80 ( .A(_abc_4108_n854), .B(_abc_4108_n638_1), .Y(_abc_4108_n855_1) );
  NAND2X1 NAND2X1_81 ( .A(_abc_4108_n955_1), .B(_abc_4108_n1054), .Y(_abc_4108_n1055) );
  NAND2X1 NAND2X1_82 ( .A(RST), .B(_abc_4108_n955_1), .Y(counter_0__FF_INPUT) );
  NAND2X1 NAND2X1_83 ( .A(counter_0_), .B(_abc_4108_n955_1), .Y(_abc_4108_n1215) );
  NAND2X1 NAND2X1_84 ( .A(bus_sync_axi_bus_reg_data2_1_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n462) );
  NAND2X1 NAND2X1_85 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_1_), .Y(bus_sync_axi_bus__abc_3782_n463) );
  NAND2X1 NAND2X1_86 ( .A(bus_sync_axi_bus_reg_data2_2_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n465) );
  NAND2X1 NAND2X1_87 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_2_), .Y(bus_sync_axi_bus__abc_3782_n466) );
  NAND2X1 NAND2X1_88 ( .A(bus_sync_axi_bus_reg_data2_3_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n468) );
  NAND2X1 NAND2X1_89 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_3_), .Y(bus_sync_axi_bus__abc_3782_n469) );
  NAND2X1 NAND2X1_9 ( .A(RST), .B(state_4_), .Y(_abc_4108_n591) );
  NAND2X1 NAND2X1_90 ( .A(bus_sync_axi_bus_reg_data2_4_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n471) );
  NAND2X1 NAND2X1_91 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_4_), .Y(bus_sync_axi_bus__abc_3782_n472) );
  NAND2X1 NAND2X1_92 ( .A(bus_sync_axi_bus_reg_data2_5_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n474) );
  NAND2X1 NAND2X1_93 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_5_), .Y(bus_sync_axi_bus__abc_3782_n475) );
  NAND2X1 NAND2X1_94 ( .A(bus_sync_axi_bus_reg_data2_6_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n477) );
  NAND2X1 NAND2X1_95 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_6_), .Y(bus_sync_axi_bus__abc_3782_n478) );
  NAND2X1 NAND2X1_96 ( .A(bus_sync_axi_bus_reg_data2_7_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n480) );
  NAND2X1 NAND2X1_97 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_7_), .Y(bus_sync_axi_bus__abc_3782_n481) );
  NAND2X1 NAND2X1_98 ( .A(bus_sync_axi_bus_reg_data2_8_), .B(bus_sync_axi_bus__abc_3782_n461), .Y(bus_sync_axi_bus__abc_3782_n483) );
  NAND2X1 NAND2X1_99 ( .A(bus_sync_axi_bus_EECLK1), .B(bus_sync_axi_bus_reg_data1_8_), .Y(bus_sync_axi_bus__abc_3782_n484) );
  NAND3X1 NAND3X1_1 ( .A(RST), .B(state_3_), .C(axi_wready), .Y(_abc_4108_n559_1) );
  NAND3X1 NAND3X1_10 ( .A(_abc_4108_n679), .B(_abc_4108_n680), .C(_abc_4108_n681_1), .Y(_abc_4108_n682_1) );
  NAND3X1 NAND3X1_11 ( .A(_abc_4108_n669_1), .B(_abc_4108_n683), .C(_abc_4108_n675), .Y(_abc_4108_n684) );
  NAND3X1 NAND3X1_12 ( .A(_abc_4108_n652), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n685_1) );
  NAND3X1 NAND3X1_13 ( .A(_abc_4108_n601), .B(_abc_4108_n685_1), .C(_abc_4108_n687), .Y(_abc_4108_n688) );
  NAND3X1 NAND3X1_14 ( .A(_abc_4108_n686_1), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n691) );
  NAND3X1 NAND3X1_15 ( .A(_abc_4108_n601), .B(_abc_4108_n691), .C(_abc_4108_n693_1), .Y(_abc_4108_n694_1) );
  NAND3X1 NAND3X1_16 ( .A(_abc_4108_n692), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n697_1) );
  NAND3X1 NAND3X1_17 ( .A(_abc_4108_n601), .B(_abc_4108_n697_1), .C(_abc_4108_n699), .Y(_abc_4108_n700) );
  NAND3X1 NAND3X1_18 ( .A(_abc_4108_n698_1), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n703) );
  NAND3X1 NAND3X1_19 ( .A(_abc_4108_n601), .B(_abc_4108_n703), .C(_abc_4108_n705_1), .Y(_abc_4108_n706_1) );
  NAND3X1 NAND3X1_2 ( .A(counter_1_), .B(_abc_4108_n595), .C(_abc_4108_n599_1), .Y(_abc_4108_n600) );
  NAND3X1 NAND3X1_20 ( .A(_abc_4108_n704), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n709_1) );
  NAND3X1 NAND3X1_21 ( .A(_abc_4108_n601), .B(_abc_4108_n709_1), .C(_abc_4108_n711), .Y(_abc_4108_n712) );
  NAND3X1 NAND3X1_22 ( .A(_abc_4108_n710_1), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n715) );
  NAND3X1 NAND3X1_23 ( .A(_abc_4108_n601), .B(_abc_4108_n715), .C(_abc_4108_n717_1), .Y(_abc_4108_n718_1) );
  NAND3X1 NAND3X1_24 ( .A(_abc_4108_n716), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n721_1) );
  NAND3X1 NAND3X1_25 ( .A(_abc_4108_n601), .B(_abc_4108_n721_1), .C(_abc_4108_n723), .Y(_abc_4108_n724) );
  NAND3X1 NAND3X1_26 ( .A(_abc_4108_n722_1), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n727) );
  NAND3X1 NAND3X1_27 ( .A(_abc_4108_n601), .B(_abc_4108_n727), .C(_abc_4108_n729_1), .Y(_abc_4108_n730_1) );
  NAND3X1 NAND3X1_28 ( .A(_abc_4108_n728), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n733_1) );
  NAND3X1 NAND3X1_29 ( .A(_abc_4108_n601), .B(_abc_4108_n733_1), .C(_abc_4108_n735), .Y(_abc_4108_n736) );
  NAND3X1 NAND3X1_3 ( .A(_abc_4108_n615), .B(_abc_4108_n616), .C(_abc_4108_n617_1), .Y(_abc_4108_n618_1) );
  NAND3X1 NAND3X1_30 ( .A(_abc_4108_n734_1), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n739) );
  NAND3X1 NAND3X1_31 ( .A(_abc_4108_n601), .B(_abc_4108_n739), .C(_abc_4108_n741_1), .Y(_abc_4108_n742_1) );
  NAND3X1 NAND3X1_32 ( .A(_abc_4108_n740), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n745_1) );
  NAND3X1 NAND3X1_33 ( .A(_abc_4108_n601), .B(_abc_4108_n745_1), .C(_abc_4108_n747), .Y(_abc_4108_n748) );
  NAND3X1 NAND3X1_34 ( .A(_abc_4108_n746_1), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n751) );
  NAND3X1 NAND3X1_35 ( .A(_abc_4108_n601), .B(_abc_4108_n751), .C(_abc_4108_n753_1), .Y(_abc_4108_n754_1) );
  NAND3X1 NAND3X1_36 ( .A(_abc_4108_n752), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n757_1) );
  NAND3X1 NAND3X1_37 ( .A(_abc_4108_n601), .B(_abc_4108_n757_1), .C(_abc_4108_n759_1), .Y(_abc_4108_n760) );
  NAND3X1 NAND3X1_38 ( .A(_abc_4108_n758), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n763_1) );
  NAND3X1 NAND3X1_39 ( .A(_abc_4108_n601), .B(_abc_4108_n763_1), .C(_abc_4108_n765_1), .Y(_abc_4108_n766) );
  NAND3X1 NAND3X1_4 ( .A(_abc_4108_n624_1), .B(_abc_4108_n625), .C(_abc_4108_n626), .Y(_abc_4108_n627_1) );
  NAND3X1 NAND3X1_40 ( .A(_abc_4108_n764), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n769_1) );
  NAND3X1 NAND3X1_41 ( .A(_abc_4108_n601), .B(_abc_4108_n769_1), .C(_abc_4108_n771_1), .Y(_abc_4108_n772) );
  NAND3X1 NAND3X1_42 ( .A(_abc_4108_n770), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n775_1) );
  NAND3X1 NAND3X1_43 ( .A(_abc_4108_n601), .B(_abc_4108_n775_1), .C(_abc_4108_n777_1), .Y(_abc_4108_n778) );
  NAND3X1 NAND3X1_44 ( .A(_abc_4108_n776), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n781_1) );
  NAND3X1 NAND3X1_45 ( .A(_abc_4108_n601), .B(_abc_4108_n781_1), .C(_abc_4108_n783_1), .Y(_abc_4108_n784) );
  NAND3X1 NAND3X1_46 ( .A(_abc_4108_n782), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n787_1) );
  NAND3X1 NAND3X1_47 ( .A(_abc_4108_n601), .B(_abc_4108_n787_1), .C(_abc_4108_n789_1), .Y(_abc_4108_n790) );
  NAND3X1 NAND3X1_48 ( .A(_abc_4108_n788), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n793_1) );
  NAND3X1 NAND3X1_49 ( .A(_abc_4108_n601), .B(_abc_4108_n793_1), .C(_abc_4108_n795_1), .Y(_abc_4108_n796) );
  NAND3X1 NAND3X1_5 ( .A(_abc_4108_n632), .B(_abc_4108_n633_1), .C(_abc_4108_n634_1), .Y(_abc_4108_n635) );
  NAND3X1 NAND3X1_50 ( .A(_abc_4108_n794), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n799_1) );
  NAND3X1 NAND3X1_51 ( .A(_abc_4108_n601), .B(_abc_4108_n799_1), .C(_abc_4108_n801_1), .Y(_abc_4108_n802) );
  NAND3X1 NAND3X1_52 ( .A(_abc_4108_n800), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n805_1) );
  NAND3X1 NAND3X1_53 ( .A(_abc_4108_n601), .B(_abc_4108_n805_1), .C(_abc_4108_n807_1), .Y(_abc_4108_n808) );
  NAND3X1 NAND3X1_54 ( .A(_abc_4108_n806), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n811_1) );
  NAND3X1 NAND3X1_55 ( .A(_abc_4108_n601), .B(_abc_4108_n811_1), .C(_abc_4108_n813_1), .Y(_abc_4108_n814) );
  NAND3X1 NAND3X1_56 ( .A(_abc_4108_n812), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n817_1) );
  NAND3X1 NAND3X1_57 ( .A(_abc_4108_n601), .B(_abc_4108_n817_1), .C(_abc_4108_n819_1), .Y(_abc_4108_n820_1) );
  NAND3X1 NAND3X1_58 ( .A(_abc_4108_n818), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n823_1) );
  NAND3X1 NAND3X1_59 ( .A(_abc_4108_n601), .B(_abc_4108_n823_1), .C(_abc_4108_n825_1), .Y(_abc_4108_n826) );
  NAND3X1 NAND3X1_6 ( .A(_abc_4108_n661_1), .B(_abc_4108_n662_1), .C(_abc_4108_n663), .Y(_abc_4108_n664) );
  NAND3X1 NAND3X1_60 ( .A(_abc_4108_n824_1), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n829_1) );
  NAND3X1 NAND3X1_61 ( .A(_abc_4108_n601), .B(_abc_4108_n829_1), .C(_abc_4108_n831_1), .Y(_abc_4108_n832) );
  NAND3X1 NAND3X1_62 ( .A(_abc_4108_n830), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n835_1) );
  NAND3X1 NAND3X1_63 ( .A(_abc_4108_n601), .B(_abc_4108_n835_1), .C(_abc_4108_n837_1), .Y(_abc_4108_n838) );
  NAND3X1 NAND3X1_64 ( .A(_abc_4108_n836), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n841_1) );
  NAND3X1 NAND3X1_65 ( .A(_abc_4108_n601), .B(_abc_4108_n841_1), .C(_abc_4108_n843_1), .Y(_abc_4108_n844) );
  NAND3X1 NAND3X1_66 ( .A(_abc_4108_n842), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n847_1) );
  NAND3X1 NAND3X1_67 ( .A(_abc_4108_n601), .B(_abc_4108_n847_1), .C(_abc_4108_n849_1), .Y(_abc_4108_n850) );
  NAND3X1 NAND3X1_68 ( .A(_abc_4108_n848), .B(_abc_4108_n604_1), .C(_abc_4108_n684), .Y(_abc_4108_n853_1) );
  NAND3X1 NAND3X1_69 ( .A(_abc_4108_n601), .B(_abc_4108_n853_1), .C(_abc_4108_n855_1), .Y(_abc_4108_n856) );
  NAND3X1 NAND3X1_7 ( .A(_abc_4108_n665_1), .B(_abc_4108_n666_1), .C(_abc_4108_n667), .Y(_abc_4108_n668) );
  NAND3X1 NAND3X1_70 ( .A(we), .B(counter_65_), .C(_abc_4108_n955_1), .Y(_abc_4108_n956) );
  NAND3X1 NAND3X1_71 ( .A(counter_65_), .B(_abc_4108_n955_1), .C(_abc_4108_n1334), .Y(_abc_4108_n1335) );
  NAND3X1 NAND3X1_72 ( .A(RST), .B(state_4_), .C(axi_rvalid), .Y(_abc_4108_n1341) );
  NAND3X1 NAND3X1_73 ( .A(RST), .B(state_7_), .C(axi_bvalid), .Y(_abc_4108_n1345) );
  NAND3X1 NAND3X1_8 ( .A(_abc_4108_n612_1), .B(_abc_4108_n629), .C(_abc_4108_n670_1), .Y(_abc_4108_n671) );
  NAND3X1 NAND3X1_9 ( .A(_abc_4108_n613_1), .B(_abc_4108_n673_1), .C(_abc_4108_n672), .Y(_abc_4108_n674_1) );
  NOR2X1 NOR2X1_1 ( .A(_abc_4108_n561), .B(_abc_4108_n563_1), .Y(_abc_2913_n78) );
  NOR2X1 NOR2X1_10 ( .A(counter_26_), .B(counter_27_), .Y(_abc_4108_n606) );
  NOR2X1 NOR2X1_100 ( .A(_abc_4108_n1327), .B(counter_0__FF_INPUT), .Y(counter_63__FF_INPUT) );
  NOR2X1 NOR2X1_101 ( .A(_abc_4108_n1329), .B(counter_0__FF_INPUT), .Y(counter_64__FF_INPUT) );
  NOR2X1 NOR2X1_102 ( .A(_abc_4108_n1331), .B(counter_0__FF_INPUT), .Y(counter_65__FF_INPUT) );
  NOR2X1 NOR2X1_103 ( .A(CEB), .B(_abc_4108_n596), .Y(_abc_4108_n1338) );
  NOR2X1 NOR2X1_11 ( .A(counter_24_), .B(counter_25_), .Y(_abc_4108_n608_1) );
  NOR2X1 NOR2X1_12 ( .A(counter_22_), .B(counter_23_), .Y(_abc_4108_n609_1) );
  NOR2X1 NOR2X1_13 ( .A(_abc_4108_n607_1), .B(_abc_4108_n610), .Y(_abc_4108_n611) );
  NOR2X1 NOR2X1_14 ( .A(counter_16_), .B(counter_15_), .Y(_abc_4108_n612_1) );
  NOR2X1 NOR2X1_15 ( .A(counter_17_), .B(counter_14_), .Y(_abc_4108_n613_1) );
  NOR2X1 NOR2X1_16 ( .A(counter_4_), .B(counter_5_), .Y(_abc_4108_n617_1) );
  NOR2X1 NOR2X1_17 ( .A(_abc_4108_n614_1), .B(_abc_4108_n618_1), .Y(_abc_4108_n619_1) );
  NOR2X1 NOR2X1_18 ( .A(counter_32_), .B(counter_33_), .Y(_abc_4108_n621) );
  NOR2X1 NOR2X1_19 ( .A(counter_30_), .B(counter_31_), .Y(_abc_4108_n622_1) );
  NOR2X1 NOR2X1_2 ( .A(axi_bready), .B(axi_rready), .Y(_abc_4108_n566) );
  NOR2X1 NOR2X1_20 ( .A(counter_20_), .B(counter_21_), .Y(_abc_4108_n626) );
  NOR2X1 NOR2X1_21 ( .A(_abc_4108_n623_1), .B(_abc_4108_n627_1), .Y(_abc_4108_n628) );
  NOR2X1 NOR2X1_22 ( .A(counter_12_), .B(counter_11_), .Y(_abc_4108_n629) );
  NOR2X1 NOR2X1_23 ( .A(counter_13_), .B(counter_10_), .Y(_abc_4108_n630_1) );
  NOR2X1 NOR2X1_24 ( .A(counter_8_), .B(counter_9_), .Y(_abc_4108_n634_1) );
  NOR2X1 NOR2X1_25 ( .A(_abc_4108_n631), .B(_abc_4108_n635), .Y(_abc_4108_n636) );
  NOR2X1 NOR2X1_26 ( .A(counter_26_), .B(counter_24_), .Y(_abc_4108_n663) );
  NOR2X1 NOR2X1_27 ( .A(counter_10_), .B(counter_6_), .Y(_abc_4108_n665_1) );
  NOR2X1 NOR2X1_28 ( .A(counter_28_), .B(counter_31_), .Y(_abc_4108_n666_1) );
  NOR2X1 NOR2X1_29 ( .A(counter_13_), .B(counter_7_), .Y(_abc_4108_n667) );
  NOR2X1 NOR2X1_3 ( .A(we_clk), .B(_abc_4108_n571), .Y(_abc_4108_n572_1) );
  NOR2X1 NOR2X1_30 ( .A(_abc_4108_n664), .B(_abc_4108_n668), .Y(_abc_4108_n669_1) );
  NOR2X1 NOR2X1_31 ( .A(counter_27_), .B(counter_18_), .Y(_abc_4108_n673_1) );
  NOR2X1 NOR2X1_32 ( .A(_abc_4108_n671), .B(_abc_4108_n674_1), .Y(_abc_4108_n675) );
  NOR2X1 NOR2X1_33 ( .A(counter_19_), .B(counter_22_), .Y(_abc_4108_n679) );
  NOR2X1 NOR2X1_34 ( .A(counter_20_), .B(counter_23_), .Y(_abc_4108_n680) );
  NOR2X1 NOR2X1_35 ( .A(counter_3_), .B(counter_8_), .Y(_abc_4108_n681_1) );
  NOR2X1 NOR2X1_36 ( .A(_abc_4108_n678_1), .B(_abc_4108_n682_1), .Y(_abc_4108_n683) );
  NOR2X1 NOR2X1_37 ( .A(_abc_4108_n1053), .B(_abc_4108_n604_1), .Y(_abc_4108_n1054) );
  NOR2X1 NOR2X1_38 ( .A(_abc_4108_n561), .B(_abc_4108_n1215), .Y(counter_1__FF_INPUT) );
  NOR2X1 NOR2X1_39 ( .A(_abc_4108_n596), .B(counter_0__FF_INPUT), .Y(counter_2__FF_INPUT) );
  NOR2X1 NOR2X1_4 ( .A(re_clk), .B(_abc_4108_n569_1), .Y(_abc_4108_n576) );
  NOR2X1 NOR2X1_40 ( .A(_abc_4108_n615), .B(counter_0__FF_INPUT), .Y(counter_3__FF_INPUT) );
  NOR2X1 NOR2X1_41 ( .A(_abc_4108_n616), .B(counter_0__FF_INPUT), .Y(counter_4__FF_INPUT) );
  NOR2X1 NOR2X1_42 ( .A(_abc_4108_n676), .B(counter_0__FF_INPUT), .Y(counter_5__FF_INPUT) );
  NOR2X1 NOR2X1_43 ( .A(_abc_4108_n1221), .B(counter_0__FF_INPUT), .Y(counter_6__FF_INPUT) );
  NOR2X1 NOR2X1_44 ( .A(_abc_4108_n632), .B(counter_0__FF_INPUT), .Y(counter_7__FF_INPUT) );
  NOR2X1 NOR2X1_45 ( .A(_abc_4108_n633_1), .B(counter_0__FF_INPUT), .Y(counter_8__FF_INPUT) );
  NOR2X1 NOR2X1_46 ( .A(_abc_4108_n1225), .B(counter_0__FF_INPUT), .Y(counter_9__FF_INPUT) );
  NOR2X1 NOR2X1_47 ( .A(_abc_4108_n677_1), .B(counter_0__FF_INPUT), .Y(counter_10__FF_INPUT) );
  NOR2X1 NOR2X1_48 ( .A(_abc_4108_n1228), .B(counter_0__FF_INPUT), .Y(counter_11__FF_INPUT) );
  NOR2X1 NOR2X1_49 ( .A(_abc_4108_n1230), .B(counter_0__FF_INPUT), .Y(counter_12__FF_INPUT) );
  NOR2X1 NOR2X1_5 ( .A(_abc_4108_n561), .B(_abc_4108_n577_1), .Y(_abc_2913_n105) );
  NOR2X1 NOR2X1_50 ( .A(_abc_4108_n1232), .B(counter_0__FF_INPUT), .Y(counter_13__FF_INPUT) );
  NOR2X1 NOR2X1_51 ( .A(_abc_4108_n1234), .B(counter_0__FF_INPUT), .Y(counter_14__FF_INPUT) );
  NOR2X1 NOR2X1_52 ( .A(_abc_4108_n1236), .B(counter_0__FF_INPUT), .Y(counter_15__FF_INPUT) );
  NOR2X1 NOR2X1_53 ( .A(_abc_4108_n1238), .B(counter_0__FF_INPUT), .Y(counter_16__FF_INPUT) );
  NOR2X1 NOR2X1_54 ( .A(_abc_4108_n1240), .B(counter_0__FF_INPUT), .Y(counter_17__FF_INPUT) );
  NOR2X1 NOR2X1_55 ( .A(_abc_4108_n1242), .B(counter_0__FF_INPUT), .Y(counter_18__FF_INPUT) );
  NOR2X1 NOR2X1_56 ( .A(_abc_4108_n624_1), .B(counter_0__FF_INPUT), .Y(counter_19__FF_INPUT) );
  NOR2X1 NOR2X1_57 ( .A(_abc_4108_n625), .B(counter_0__FF_INPUT), .Y(counter_20__FF_INPUT) );
  NOR2X1 NOR2X1_58 ( .A(_abc_4108_n1246), .B(counter_0__FF_INPUT), .Y(counter_21__FF_INPUT) );
  NOR2X1 NOR2X1_59 ( .A(_abc_4108_n1248), .B(counter_0__FF_INPUT), .Y(counter_22__FF_INPUT) );
  NOR2X1 NOR2X1_6 ( .A(state_6_), .B(state_4_), .Y(_abc_4108_n580) );
  NOR2X1 NOR2X1_60 ( .A(_abc_4108_n1250), .B(counter_0__FF_INPUT), .Y(counter_23__FF_INPUT) );
  NOR2X1 NOR2X1_61 ( .A(_abc_4108_n1252), .B(counter_0__FF_INPUT), .Y(counter_24__FF_INPUT) );
  NOR2X1 NOR2X1_62 ( .A(_abc_4108_n1254), .B(counter_0__FF_INPUT), .Y(counter_25__FF_INPUT) );
  NOR2X1 NOR2X1_63 ( .A(_abc_4108_n662_1), .B(counter_0__FF_INPUT), .Y(counter_26__FF_INPUT) );
  NOR2X1 NOR2X1_64 ( .A(_abc_4108_n1257), .B(counter_0__FF_INPUT), .Y(counter_27__FF_INPUT) );
  NOR2X1 NOR2X1_65 ( .A(_abc_4108_n1259), .B(counter_0__FF_INPUT), .Y(counter_28__FF_INPUT) );
  NOR2X1 NOR2X1_66 ( .A(_abc_4108_n1261), .B(counter_0__FF_INPUT), .Y(counter_29__FF_INPUT) );
  NOR2X1 NOR2X1_67 ( .A(_abc_4108_n661_1), .B(counter_0__FF_INPUT), .Y(counter_30__FF_INPUT) );
  NOR2X1 NOR2X1_68 ( .A(_abc_4108_n1264), .B(counter_0__FF_INPUT), .Y(counter_31__FF_INPUT) );
  NOR2X1 NOR2X1_69 ( .A(_abc_4108_n1266), .B(counter_0__FF_INPUT), .Y(counter_32__FF_INPUT) );
  NOR2X1 NOR2X1_7 ( .A(state_3_), .B(state_7_), .Y(_abc_4108_n587_1) );
  NOR2X1 NOR2X1_70 ( .A(_abc_4108_n1268), .B(counter_0__FF_INPUT), .Y(counter_33__FF_INPUT) );
  NOR2X1 NOR2X1_71 ( .A(_abc_4108_n1053), .B(counter_0__FF_INPUT), .Y(counter_34__FF_INPUT) );
  NOR2X1 NOR2X1_72 ( .A(_abc_4108_n1271), .B(counter_0__FF_INPUT), .Y(counter_35__FF_INPUT) );
  NOR2X1 NOR2X1_73 ( .A(_abc_4108_n1273), .B(counter_0__FF_INPUT), .Y(counter_36__FF_INPUT) );
  NOR2X1 NOR2X1_74 ( .A(_abc_4108_n1275), .B(counter_0__FF_INPUT), .Y(counter_37__FF_INPUT) );
  NOR2X1 NOR2X1_75 ( .A(_abc_4108_n1277), .B(counter_0__FF_INPUT), .Y(counter_38__FF_INPUT) );
  NOR2X1 NOR2X1_76 ( .A(_abc_4108_n1279), .B(counter_0__FF_INPUT), .Y(counter_39__FF_INPUT) );
  NOR2X1 NOR2X1_77 ( .A(_abc_4108_n1281), .B(counter_0__FF_INPUT), .Y(counter_40__FF_INPUT) );
  NOR2X1 NOR2X1_78 ( .A(_abc_4108_n1283), .B(counter_0__FF_INPUT), .Y(counter_41__FF_INPUT) );
  NOR2X1 NOR2X1_79 ( .A(_abc_4108_n1285), .B(counter_0__FF_INPUT), .Y(counter_42__FF_INPUT) );
  NOR2X1 NOR2X1_8 ( .A(_abc_4108_n595), .B(_abc_4108_n596), .Y(_abc_4108_n597_1) );
  NOR2X1 NOR2X1_80 ( .A(_abc_4108_n1287), .B(counter_0__FF_INPUT), .Y(counter_43__FF_INPUT) );
  NOR2X1 NOR2X1_81 ( .A(_abc_4108_n1289), .B(counter_0__FF_INPUT), .Y(counter_44__FF_INPUT) );
  NOR2X1 NOR2X1_82 ( .A(_abc_4108_n1291), .B(counter_0__FF_INPUT), .Y(counter_45__FF_INPUT) );
  NOR2X1 NOR2X1_83 ( .A(_abc_4108_n1293), .B(counter_0__FF_INPUT), .Y(counter_46__FF_INPUT) );
  NOR2X1 NOR2X1_84 ( .A(_abc_4108_n1295), .B(counter_0__FF_INPUT), .Y(counter_47__FF_INPUT) );
  NOR2X1 NOR2X1_85 ( .A(_abc_4108_n1297), .B(counter_0__FF_INPUT), .Y(counter_48__FF_INPUT) );
  NOR2X1 NOR2X1_86 ( .A(_abc_4108_n1299), .B(counter_0__FF_INPUT), .Y(counter_49__FF_INPUT) );
  NOR2X1 NOR2X1_87 ( .A(_abc_4108_n1301), .B(counter_0__FF_INPUT), .Y(counter_50__FF_INPUT) );
  NOR2X1 NOR2X1_88 ( .A(_abc_4108_n1303), .B(counter_0__FF_INPUT), .Y(counter_51__FF_INPUT) );
  NOR2X1 NOR2X1_89 ( .A(_abc_4108_n1305), .B(counter_0__FF_INPUT), .Y(counter_52__FF_INPUT) );
  NOR2X1 NOR2X1_9 ( .A(counter_28_), .B(counter_29_), .Y(_abc_4108_n605) );
  NOR2X1 NOR2X1_90 ( .A(_abc_4108_n1307), .B(counter_0__FF_INPUT), .Y(counter_53__FF_INPUT) );
  NOR2X1 NOR2X1_91 ( .A(_abc_4108_n1309), .B(counter_0__FF_INPUT), .Y(counter_54__FF_INPUT) );
  NOR2X1 NOR2X1_92 ( .A(_abc_4108_n1311), .B(counter_0__FF_INPUT), .Y(counter_55__FF_INPUT) );
  NOR2X1 NOR2X1_93 ( .A(_abc_4108_n1313), .B(counter_0__FF_INPUT), .Y(counter_56__FF_INPUT) );
  NOR2X1 NOR2X1_94 ( .A(_abc_4108_n1315), .B(counter_0__FF_INPUT), .Y(counter_57__FF_INPUT) );
  NOR2X1 NOR2X1_95 ( .A(_abc_4108_n1317), .B(counter_0__FF_INPUT), .Y(counter_58__FF_INPUT) );
  NOR2X1 NOR2X1_96 ( .A(_abc_4108_n1319), .B(counter_0__FF_INPUT), .Y(counter_59__FF_INPUT) );
  NOR2X1 NOR2X1_97 ( .A(_abc_4108_n1321), .B(counter_0__FF_INPUT), .Y(counter_60__FF_INPUT) );
  NOR2X1 NOR2X1_98 ( .A(_abc_4108_n1323), .B(counter_0__FF_INPUT), .Y(counter_61__FF_INPUT) );
  NOR2X1 NOR2X1_99 ( .A(_abc_4108_n1325), .B(counter_0__FF_INPUT), .Y(counter_62__FF_INPUT) );
  NOR3X1 NOR3X1_1 ( .A(counter_5_), .B(counter_2_), .C(counter_30_), .Y(_abc_4108_n670_1) );
  NOR3X1 NOR3X1_2 ( .A(counter_32_), .B(counter_33_), .C(counter_21_), .Y(_abc_4108_n672) );
  OAI21X1 OAI21X1_1 ( .A(axi_bvalid), .B(_abc_4108_n558_1), .C(_abc_4108_n559_1), .Y(_abc_2913_n70) );
  OAI21X1 OAI21X1_10 ( .A(bus_cap_1_), .B(_abc_4108_n638_1), .C(_abc_4108_n653_1), .Y(_abc_4108_n654_1) );
  OAI21X1 OAI21X1_100 ( .A(CEB), .B(sft_reg_21_), .C(RST), .Y(_abc_4108_n1123) );
  OAI21X1 OAI21X1_101 ( .A(CEB), .B(sft_reg_22_), .C(RST), .Y(_abc_4108_n1126) );
  OAI21X1 OAI21X1_102 ( .A(CEB), .B(sft_reg_23_), .C(RST), .Y(_abc_4108_n1129) );
  OAI21X1 OAI21X1_103 ( .A(CEB), .B(sft_reg_24_), .C(RST), .Y(_abc_4108_n1132) );
  OAI21X1 OAI21X1_104 ( .A(CEB), .B(sft_reg_25_), .C(RST), .Y(_abc_4108_n1135) );
  OAI21X1 OAI21X1_105 ( .A(CEB), .B(sft_reg_26_), .C(RST), .Y(_abc_4108_n1138) );
  OAI21X1 OAI21X1_106 ( .A(CEB), .B(sft_reg_27_), .C(RST), .Y(_abc_4108_n1141) );
  OAI21X1 OAI21X1_107 ( .A(CEB), .B(sft_reg_28_), .C(RST), .Y(_abc_4108_n1144) );
  OAI21X1 OAI21X1_108 ( .A(CEB), .B(sft_reg_29_), .C(RST), .Y(_abc_4108_n1147) );
  OAI21X1 OAI21X1_109 ( .A(sft_reg_30_), .B(_abc_4108_n1055), .C(RST), .Y(_abc_4108_n1150) );
  OAI21X1 OAI21X1_11 ( .A(bus_sync_rdata_data_out_2_), .B(_abc_4108_n598_1), .C(RST), .Y(_abc_4108_n656) );
  OAI21X1 OAI21X1_110 ( .A(DATA), .B(_abc_4108_n1335), .C(RST), .Y(_abc_4108_n1336) );
  OAI21X1 OAI21X1_111 ( .A(re), .B(_abc_4108_n1338), .C(RST), .Y(_abc_4108_n1339) );
  OAI21X1 OAI21X1_112 ( .A(DATA), .B(_abc_4108_n1215), .C(RST), .Y(_abc_4108_n1343) );
  OAI21X1 OAI21X1_113 ( .A(bus_sync_axi_bus_reg_data2_0_), .B(bus_sync_axi_bus_EECLK1), .C(RST), .Y(bus_sync_axi_bus__abc_3782_n458) );
  OAI21X1 OAI21X1_114 ( .A(bus_sync_rdata_reg_data2_0_), .B(bus_sync_rdata_EECLK2), .C(RST), .Y(bus_sync_rdata__abc_3590_n202_1) );
  OAI21X1 OAI21X1_115 ( .A(bus_sync_state_machine_reg_data2_0_), .B(bus_sync_state_machine_EECLK1), .C(RST), .Y(bus_sync_state_machine__abc_3756_n38) );
  OAI21X1 OAI21X1_116 ( .A(bus_sync_status_reg_data2_0_), .B(bus_sync_status_EECLK2), .C(RST), .Y(bus_sync_status__abc_3569_n31) );
  OAI21X1 OAI21X1_12 ( .A(_abc_4108_n600), .B(_abc_4108_n655), .C(_abc_4108_n657_1), .Y(_abc_4108_n658_1) );
  OAI21X1 OAI21X1_13 ( .A(\axi_rdata[0] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n859_1) );
  OAI21X1 OAI21X1_14 ( .A(\axi_rdata[1] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n862) );
  OAI21X1 OAI21X1_15 ( .A(\axi_rdata[2] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n865_1) );
  OAI21X1 OAI21X1_16 ( .A(\axi_rdata[3] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n868) );
  OAI21X1 OAI21X1_17 ( .A(\axi_rdata[4] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n871_1) );
  OAI21X1 OAI21X1_18 ( .A(\axi_rdata[5] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n874) );
  OAI21X1 OAI21X1_19 ( .A(\axi_rdata[6] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n877_1) );
  OAI21X1 OAI21X1_2 ( .A(re_clk), .B(_abc_4108_n569_1), .C(RST), .Y(_abc_4108_n570) );
  OAI21X1 OAI21X1_20 ( .A(\axi_rdata[7] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n880) );
  OAI21X1 OAI21X1_21 ( .A(\axi_rdata[8] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n883_1) );
  OAI21X1 OAI21X1_22 ( .A(\axi_rdata[9] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n886) );
  OAI21X1 OAI21X1_23 ( .A(\axi_rdata[10] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n889_1) );
  OAI21X1 OAI21X1_24 ( .A(\axi_rdata[11] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n892_1) );
  OAI21X1 OAI21X1_25 ( .A(\axi_rdata[12] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n895_1) );
  OAI21X1 OAI21X1_26 ( .A(\axi_rdata[13] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n898_1) );
  OAI21X1 OAI21X1_27 ( .A(\axi_rdata[14] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n901_1) );
  OAI21X1 OAI21X1_28 ( .A(\axi_rdata[15] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n904_1) );
  OAI21X1 OAI21X1_29 ( .A(\axi_rdata[16] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n907_1) );
  OAI21X1 OAI21X1_3 ( .A(we_clk), .B(_abc_4108_n571), .C(state_0_), .Y(_abc_4108_n582_1) );
  OAI21X1 OAI21X1_30 ( .A(\axi_rdata[17] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n910_1) );
  OAI21X1 OAI21X1_31 ( .A(\axi_rdata[18] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n913_1) );
  OAI21X1 OAI21X1_32 ( .A(\axi_rdata[19] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n916_1) );
  OAI21X1 OAI21X1_33 ( .A(\axi_rdata[20] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n919_1) );
  OAI21X1 OAI21X1_34 ( .A(\axi_rdata[21] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n922_1) );
  OAI21X1 OAI21X1_35 ( .A(\axi_rdata[22] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n925_1) );
  OAI21X1 OAI21X1_36 ( .A(\axi_rdata[23] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n928_1) );
  OAI21X1 OAI21X1_37 ( .A(\axi_rdata[24] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n931_1) );
  OAI21X1 OAI21X1_38 ( .A(\axi_rdata[25] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n934_1) );
  OAI21X1 OAI21X1_39 ( .A(\axi_rdata[26] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n937_1) );
  OAI21X1 OAI21X1_4 ( .A(_abc_4108_n570), .B(_abc_4108_n582_1), .C(_abc_4108_n584_1), .Y(_abc_2913_n116) );
  OAI21X1 OAI21X1_40 ( .A(\axi_rdata[27] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n940_1) );
  OAI21X1 OAI21X1_41 ( .A(\axi_rdata[28] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n943_1) );
  OAI21X1 OAI21X1_42 ( .A(\axi_rdata[29] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n946_1) );
  OAI21X1 OAI21X1_43 ( .A(\axi_rdata[30] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n949_1) );
  OAI21X1 OAI21X1_44 ( .A(\axi_rdata[31] ), .B(_abc_4108_n579_1), .C(RST), .Y(_abc_4108_n952) );
  OAI21X1 OAI21X1_45 ( .A(DATA), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n957) );
  OAI21X1 OAI21X1_46 ( .A(sft_reg_0_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n960) );
  OAI21X1 OAI21X1_47 ( .A(sft_reg_1_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n963_1) );
  OAI21X1 OAI21X1_48 ( .A(sft_reg_2_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n966_1) );
  OAI21X1 OAI21X1_49 ( .A(sft_reg_3_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n969_1) );
  OAI21X1 OAI21X1_5 ( .A(_abc_4108_n620), .B(_abc_4108_n637_1), .C(_abc_4108_n604_1), .Y(_abc_4108_n638_1) );
  OAI21X1 OAI21X1_50 ( .A(sft_reg_4_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n972) );
  OAI21X1 OAI21X1_51 ( .A(sft_reg_5_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n975) );
  OAI21X1 OAI21X1_52 ( .A(sft_reg_6_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n978) );
  OAI21X1 OAI21X1_53 ( .A(sft_reg_7_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n981) );
  OAI21X1 OAI21X1_54 ( .A(sft_reg_8_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n984) );
  OAI21X1 OAI21X1_55 ( .A(sft_reg_9_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n987) );
  OAI21X1 OAI21X1_56 ( .A(sft_reg_10_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n990) );
  OAI21X1 OAI21X1_57 ( .A(sft_reg_11_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n993) );
  OAI21X1 OAI21X1_58 ( .A(sft_reg_12_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n996) );
  OAI21X1 OAI21X1_59 ( .A(sft_reg_13_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n999) );
  OAI21X1 OAI21X1_6 ( .A(bus_sync_rdata_data_out_0_), .B(_abc_4108_n598_1), .C(RST), .Y(_abc_4108_n642_1) );
  OAI21X1 OAI21X1_60 ( .A(sft_reg_14_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1002) );
  OAI21X1 OAI21X1_61 ( .A(sft_reg_15_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1005) );
  OAI21X1 OAI21X1_62 ( .A(sft_reg_16_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1008) );
  OAI21X1 OAI21X1_63 ( .A(sft_reg_17_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1011) );
  OAI21X1 OAI21X1_64 ( .A(sft_reg_18_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1014) );
  OAI21X1 OAI21X1_65 ( .A(sft_reg_19_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1017) );
  OAI21X1 OAI21X1_66 ( .A(sft_reg_20_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1020) );
  OAI21X1 OAI21X1_67 ( .A(sft_reg_21_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1023) );
  OAI21X1 OAI21X1_68 ( .A(sft_reg_22_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1026) );
  OAI21X1 OAI21X1_69 ( .A(sft_reg_23_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1029) );
  OAI21X1 OAI21X1_7 ( .A(_abc_4108_n600), .B(_abc_4108_n641_1), .C(_abc_4108_n643), .Y(_abc_4108_n644) );
  OAI21X1 OAI21X1_70 ( .A(sft_reg_24_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1032) );
  OAI21X1 OAI21X1_71 ( .A(sft_reg_25_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1035) );
  OAI21X1 OAI21X1_72 ( .A(sft_reg_26_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1038) );
  OAI21X1 OAI21X1_73 ( .A(sft_reg_27_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1041) );
  OAI21X1 OAI21X1_74 ( .A(sft_reg_28_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1044) );
  OAI21X1 OAI21X1_75 ( .A(sft_reg_29_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1047) );
  OAI21X1 OAI21X1_76 ( .A(sft_reg_30_), .B(_abc_4108_n956), .C(RST), .Y(_abc_4108_n1050) );
  OAI21X1 OAI21X1_77 ( .A(DATA), .B(CEB), .C(RST), .Y(_abc_4108_n1056) );
  OAI21X1 OAI21X1_78 ( .A(_abc_4108_n1053), .B(_abc_4108_n604_1), .C(RST), .Y(_abc_4108_n1057) );
  OAI21X1 OAI21X1_79 ( .A(CEB), .B(sft_reg_0_), .C(RST), .Y(_abc_4108_n1060) );
  OAI21X1 OAI21X1_8 ( .A(bus_sync_rdata_data_out_1_), .B(_abc_4108_n598_1), .C(RST), .Y(_abc_4108_n648) );
  OAI21X1 OAI21X1_80 ( .A(CEB), .B(sft_reg_1_), .C(RST), .Y(_abc_4108_n1063) );
  OAI21X1 OAI21X1_81 ( .A(CEB), .B(sft_reg_2_), .C(RST), .Y(_abc_4108_n1066) );
  OAI21X1 OAI21X1_82 ( .A(CEB), .B(sft_reg_3_), .C(RST), .Y(_abc_4108_n1069) );
  OAI21X1 OAI21X1_83 ( .A(CEB), .B(sft_reg_4_), .C(RST), .Y(_abc_4108_n1072) );
  OAI21X1 OAI21X1_84 ( .A(CEB), .B(sft_reg_5_), .C(RST), .Y(_abc_4108_n1075) );
  OAI21X1 OAI21X1_85 ( .A(CEB), .B(sft_reg_6_), .C(RST), .Y(_abc_4108_n1078) );
  OAI21X1 OAI21X1_86 ( .A(CEB), .B(sft_reg_7_), .C(RST), .Y(_abc_4108_n1081) );
  OAI21X1 OAI21X1_87 ( .A(CEB), .B(sft_reg_8_), .C(RST), .Y(_abc_4108_n1084) );
  OAI21X1 OAI21X1_88 ( .A(CEB), .B(sft_reg_9_), .C(RST), .Y(_abc_4108_n1087) );
  OAI21X1 OAI21X1_89 ( .A(CEB), .B(sft_reg_10_), .C(RST), .Y(_abc_4108_n1090) );
  OAI21X1 OAI21X1_9 ( .A(_abc_4108_n600), .B(_abc_4108_n647), .C(_abc_4108_n649_1), .Y(_abc_4108_n650_1) );
  OAI21X1 OAI21X1_90 ( .A(CEB), .B(sft_reg_11_), .C(RST), .Y(_abc_4108_n1093) );
  OAI21X1 OAI21X1_91 ( .A(CEB), .B(sft_reg_12_), .C(RST), .Y(_abc_4108_n1096) );
  OAI21X1 OAI21X1_92 ( .A(CEB), .B(sft_reg_13_), .C(RST), .Y(_abc_4108_n1099) );
  OAI21X1 OAI21X1_93 ( .A(CEB), .B(sft_reg_14_), .C(RST), .Y(_abc_4108_n1102) );
  OAI21X1 OAI21X1_94 ( .A(CEB), .B(sft_reg_15_), .C(RST), .Y(_abc_4108_n1105) );
  OAI21X1 OAI21X1_95 ( .A(CEB), .B(sft_reg_16_), .C(RST), .Y(_abc_4108_n1108) );
  OAI21X1 OAI21X1_96 ( .A(CEB), .B(sft_reg_17_), .C(RST), .Y(_abc_4108_n1111) );
  OAI21X1 OAI21X1_97 ( .A(CEB), .B(sft_reg_18_), .C(RST), .Y(_abc_4108_n1114) );
  OAI21X1 OAI21X1_98 ( .A(CEB), .B(sft_reg_19_), .C(RST), .Y(_abc_4108_n1117) );
  OAI21X1 OAI21X1_99 ( .A(CEB), .B(sft_reg_20_), .C(RST), .Y(_abc_4108_n1120) );
  OAI22X1 OAI22X1_1 ( .A(axi_arready), .B(_abc_4108_n568_1), .C(_abc_4108_n570), .D(_abc_4108_n573_1), .Y(_abc_2913_n95) );
  OAI22X1 OAI22X1_2 ( .A(_abc_4108_n590), .B(_abc_4108_n568_1), .C(axi_rvalid), .D(_abc_4108_n591), .Y(_abc_2913_n129) );
  OR2X2 OR2X2_1 ( .A(axi_wvalid), .B(state_5_), .Y(axi_awvalid) );
  OR2X2 OR2X2_2 ( .A(axi_arvalid), .B(state_1_), .Y(_abc_4108_n593_1) );
  OR2X2 OR2X2_3 ( .A(_abc_4108_n593_1), .B(axi_awvalid), .Y(busy) );
  OR2X2 OR2X2_4 ( .A(re), .B(we), .Y(_abc_4108_n602_1) );
  OR2X2 OR2X2_5 ( .A(_abc_4108_n640), .B(bus_sync_status_data_out_0_), .Y(_abc_4108_n641_1) );
  OR2X2 OR2X2_6 ( .A(_abc_4108_n640), .B(bus_sync_status_data_out_1_), .Y(_abc_4108_n647) );
  OR2X2 OR2X2_7 ( .A(_abc_4108_n640), .B(bus_sync_status_data_out_2_), .Y(_abc_4108_n655) );
endmodule