module b08_reset(clock, RESET_G, nRESET_G, START, I_7_, I_6_, I_5_, I_4_, I_3_, I_2_, I_1_, I_0_, O_REG_3_, O_REG_2_, O_REG_1_, O_REG_0_);

wire IN_R_REG_0_; 
wire IN_R_REG_1_; 
wire IN_R_REG_2_; 
wire IN_R_REG_3_; 
wire IN_R_REG_4_; 
wire IN_R_REG_5_; 
wire IN_R_REG_6_; 
wire IN_R_REG_7_; 
input I_0_;
input I_1_;
input I_2_;
input I_3_;
input I_4_;
input I_5_;
input I_6_;
input I_7_;
wire MAR_REG_0_; 
wire MAR_REG_1_; 
wire MAR_REG_2_; 
wire OUT_R_REG_0_; 
wire OUT_R_REG_1_; 
wire OUT_R_REG_2_; 
wire OUT_R_REG_3_; 
output O_REG_0_;
output O_REG_1_;
output O_REG_2_;
output O_REG_3_;
input RESET_G;
input START;
wire STATO_REG_0_; 
wire STATO_REG_1_; 
wire _abc_1014_new_n100_; 
wire _abc_1014_new_n101_; 
wire _abc_1014_new_n102_; 
wire _abc_1014_new_n103_; 
wire _abc_1014_new_n104_; 
wire _abc_1014_new_n105_; 
wire _abc_1014_new_n106_; 
wire _abc_1014_new_n107_; 
wire _abc_1014_new_n108_; 
wire _abc_1014_new_n109_; 
wire _abc_1014_new_n110_; 
wire _abc_1014_new_n111_; 
wire _abc_1014_new_n112_; 
wire _abc_1014_new_n113_; 
wire _abc_1014_new_n114_; 
wire _abc_1014_new_n115_; 
wire _abc_1014_new_n116_; 
wire _abc_1014_new_n117_; 
wire _abc_1014_new_n118_; 
wire _abc_1014_new_n119_; 
wire _abc_1014_new_n120_; 
wire _abc_1014_new_n121_; 
wire _abc_1014_new_n122_; 
wire _abc_1014_new_n123_; 
wire _abc_1014_new_n124_; 
wire _abc_1014_new_n125_; 
wire _abc_1014_new_n126_; 
wire _abc_1014_new_n127_; 
wire _abc_1014_new_n128_; 
wire _abc_1014_new_n129_; 
wire _abc_1014_new_n130_; 
wire _abc_1014_new_n131_; 
wire _abc_1014_new_n132_; 
wire _abc_1014_new_n133_; 
wire _abc_1014_new_n135_; 
wire _abc_1014_new_n136_; 
wire _abc_1014_new_n138_; 
wire _abc_1014_new_n139_; 
wire _abc_1014_new_n141_; 
wire _abc_1014_new_n143_; 
wire _abc_1014_new_n144_; 
wire _abc_1014_new_n146_; 
wire _abc_1014_new_n147_; 
wire _abc_1014_new_n149_; 
wire _abc_1014_new_n151_; 
wire _abc_1014_new_n152_; 
wire _abc_1014_new_n154_; 
wire _abc_1014_new_n155_; 
wire _abc_1014_new_n156_; 
wire _abc_1014_new_n158_; 
wire _abc_1014_new_n159_; 
wire _abc_1014_new_n161_; 
wire _abc_1014_new_n163_; 
wire _abc_1014_new_n164_; 
wire _abc_1014_new_n166_; 
wire _abc_1014_new_n167_; 
wire _abc_1014_new_n169_; 
wire _abc_1014_new_n170_; 
wire _abc_1014_new_n172_; 
wire _abc_1014_new_n173_; 
wire _abc_1014_new_n53_; 
wire _abc_1014_new_n54_; 
wire _abc_1014_new_n55_; 
wire _abc_1014_new_n56_; 
wire _abc_1014_new_n57_; 
wire _abc_1014_new_n58_; 
wire _abc_1014_new_n60_; 
wire _abc_1014_new_n61_; 
wire _abc_1014_new_n62_; 
wire _abc_1014_new_n64_; 
wire _abc_1014_new_n65_; 
wire _abc_1014_new_n66_; 
wire _abc_1014_new_n67_; 
wire _abc_1014_new_n68_; 
wire _abc_1014_new_n69_; 
wire _abc_1014_new_n70_; 
wire _abc_1014_new_n72_; 
wire _abc_1014_new_n73_; 
wire _abc_1014_new_n75_; 
wire _abc_1014_new_n76_; 
wire _abc_1014_new_n78_; 
wire _abc_1014_new_n79_; 
wire _abc_1014_new_n81_; 
wire _abc_1014_new_n82_; 
wire _abc_1014_new_n83_; 
wire _abc_1014_new_n84_; 
wire _abc_1014_new_n85_; 
wire _abc_1014_new_n86_; 
wire _abc_1014_new_n87_; 
wire _abc_1014_new_n88_; 
wire _abc_1014_new_n89_; 
wire _abc_1014_new_n90_; 
wire _abc_1014_new_n91_; 
wire _abc_1014_new_n92_; 
wire _abc_1014_new_n93_; 
wire _abc_1014_new_n94_; 
wire _abc_1014_new_n95_; 
wire _abc_1014_new_n96_; 
wire _abc_1014_new_n97_; 
wire _abc_1014_new_n98_; 
wire _abc_1014_new_n99_; 
input clock;
wire n101; 
wire n106; 
wire n111; 
wire n116; 
wire n121; 
wire n125; 
wire n129; 
wire n32; 
wire n36; 
wire n41; 
wire n46; 
wire n51; 
wire n56; 
wire n61; 
wire n66; 
wire n71; 
wire n76; 
wire n81; 
wire n86; 
wire n91; 
wire n96; 
input nRESET_G;
AOI21X1 AOI21X1_1 ( .A(_abc_1014_new_n54_), .B(I_0_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n62_));
AOI21X1 AOI21X1_10 ( .A(_abc_1014_new_n132_), .B(_abc_1014_new_n83_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n133_));
AOI21X1 AOI21X1_11 ( .A(_abc_1014_new_n55_), .B(OUT_R_REG_2_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n136_));
AOI21X1 AOI21X1_12 ( .A(_abc_1014_new_n55_), .B(OUT_R_REG_1_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n139_));
AOI21X1 AOI21X1_13 ( .A(_abc_1014_new_n143_), .B(_abc_1014_new_n66_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n144_));
AOI21X1 AOI21X1_14 ( .A(_abc_1014_new_n146_), .B(START), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n147_));
AOI21X1 AOI21X1_15 ( .A(_abc_1014_new_n66_), .B(_abc_1014_new_n84_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n152_));
AOI21X1 AOI21X1_16 ( .A(_abc_1014_new_n54_), .B(I_6_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n161_));
AOI21X1 AOI21X1_17 ( .A(_abc_1014_new_n55_), .B(IN_R_REG_4_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n167_));
AOI21X1 AOI21X1_18 ( .A(_abc_1014_new_n55_), .B(IN_R_REG_3_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n170_));
AOI21X1 AOI21X1_2 ( .A(_abc_1014_new_n69_), .B(O_REG_3_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n70_));
AOI21X1 AOI21X1_3 ( .A(_abc_1014_new_n69_), .B(O_REG_2_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n73_));
AOI21X1 AOI21X1_4 ( .A(_abc_1014_new_n69_), .B(O_REG_1_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n76_));
AOI21X1 AOI21X1_5 ( .A(_abc_1014_new_n69_), .B(O_REG_0_), .C(_abc_1014_new_n61_), .Y(_abc_1014_new_n79_));
AOI21X1 AOI21X1_6 ( .A(_abc_1014_new_n111_), .B(_abc_1014_new_n106_), .C(_abc_1014_new_n103_), .Y(_abc_1014_new_n112_));
AOI21X1 AOI21X1_7 ( .A(_abc_1014_new_n85_), .B(MAR_REG_0_), .C(_abc_1014_new_n82_), .Y(_abc_1014_new_n119_));
AOI21X1 AOI21X1_8 ( .A(_abc_1014_new_n125_), .B(_abc_1014_new_n126_), .C(IN_R_REG_3_), .Y(_abc_1014_new_n127_));
AOI21X1 AOI21X1_9 ( .A(_abc_1014_new_n86_), .B(_abc_1014_new_n113_), .C(_abc_1014_new_n131_), .Y(_abc_1014_new_n132_));
AOI22X1 AOI22X1_1 ( .A(OUT_R_REG_3_), .B(_abc_1014_new_n55_), .C(_abc_1014_new_n116_), .D(_abc_1014_new_n132_), .Y(_abc_1014_new_n141_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n121), .Q(O_REG_3_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(n61), .Q(IN_R_REG_7_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(n66), .Q(IN_R_REG_6_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(n71), .Q(IN_R_REG_5_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(n76), .Q(IN_R_REG_4_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(n81), .Q(IN_R_REG_3_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(n86), .Q(IN_R_REG_2_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(n91), .Q(IN_R_REG_1_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(n96), .Q(IN_R_REG_0_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(n101), .Q(OUT_R_REG_3_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(n106), .Q(OUT_R_REG_2_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n129), .Q(O_REG_1_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(n111), .Q(OUT_R_REG_1_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(n116), .Q(OUT_R_REG_0_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n41), .Q(STATO_REG_0_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n32), .Q(O_REG_0_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n36), .Q(STATO_REG_1_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n125), .Q(O_REG_2_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n46), .Q(MAR_REG_2_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n51), .Q(MAR_REG_1_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(n56), .Q(MAR_REG_0_));
INVX1 INVX1_1 ( .A(STATO_REG_0_), .Y(_abc_1014_new_n53_));
INVX1 INVX1_10 ( .A(OUT_R_REG_0_), .Y(_abc_1014_new_n78_));
INVX1 INVX1_11 ( .A(MAR_REG_1_), .Y(_abc_1014_new_n82_));
INVX1 INVX1_12 ( .A(MAR_REG_0_), .Y(_abc_1014_new_n84_));
INVX1 INVX1_13 ( .A(MAR_REG_2_), .Y(_abc_1014_new_n85_));
INVX1 INVX1_14 ( .A(_abc_1014_new_n105_), .Y(_abc_1014_new_n106_));
INVX1 INVX1_15 ( .A(IN_R_REG_7_), .Y(_abc_1014_new_n107_));
INVX1 INVX1_16 ( .A(IN_R_REG_2_), .Y(_abc_1014_new_n109_));
INVX1 INVX1_17 ( .A(IN_R_REG_6_), .Y(_abc_1014_new_n114_));
INVX1 INVX1_18 ( .A(IN_R_REG_5_), .Y(_abc_1014_new_n122_));
INVX1 INVX1_19 ( .A(_abc_1014_new_n88_), .Y(_abc_1014_new_n125_));
INVX1 INVX1_2 ( .A(_abc_1014_new_n54_), .Y(_abc_1014_new_n55_));
INVX1 INVX1_20 ( .A(_abc_1014_new_n132_), .Y(_abc_1014_new_n135_));
INVX1 INVX1_21 ( .A(_abc_1014_new_n90_), .Y(_abc_1014_new_n138_));
INVX1 INVX1_22 ( .A(_abc_1014_new_n94_), .Y(_abc_1014_new_n143_));
INVX1 INVX1_23 ( .A(_abc_1014_new_n146_), .Y(_abc_1014_new_n151_));
INVX1 INVX1_24 ( .A(I_4_), .Y(_abc_1014_new_n166_));
INVX1 INVX1_25 ( .A(I_3_), .Y(_abc_1014_new_n169_));
INVX1 INVX1_3 ( .A(IN_R_REG_1_), .Y(_abc_1014_new_n56_));
INVX1 INVX1_4 ( .A(IN_R_REG_0_), .Y(_abc_1014_new_n60_));
INVX1 INVX1_5 ( .A(nRESET_G), .Y(_abc_1014_new_n61_));
INVX1 INVX1_6 ( .A(OUT_R_REG_3_), .Y(_abc_1014_new_n64_));
INVX1 INVX1_7 ( .A(STATO_REG_1_), .Y(_abc_1014_new_n65_));
INVX1 INVX1_8 ( .A(OUT_R_REG_2_), .Y(_abc_1014_new_n72_));
INVX1 INVX1_9 ( .A(OUT_R_REG_1_), .Y(_abc_1014_new_n75_));
MUX2X1 MUX2X1_1 ( .A(MAR_REG_0_), .B(MAR_REG_2_), .S(MAR_REG_1_), .Y(_abc_1014_new_n99_));
MUX2X1 MUX2X1_2 ( .A(_abc_1014_new_n128_), .B(_abc_1014_new_n94_), .S(IN_R_REG_4_), .Y(_abc_1014_new_n129_));
NAND2X1 NAND2X1_1 ( .A(nRESET_G), .B(_abc_1014_new_n58_), .Y(n91));
NAND2X1 NAND2X1_10 ( .A(_abc_1014_new_n101_), .B(_abc_1014_new_n117_), .Y(_abc_1014_new_n118_));
NAND2X1 NAND2X1_11 ( .A(MAR_REG_2_), .B(_abc_1014_new_n84_), .Y(_abc_1014_new_n126_));
NAND2X1 NAND2X1_12 ( .A(_abc_1014_new_n81_), .B(_abc_1014_new_n133_), .Y(n116));
NAND2X1 NAND2X1_13 ( .A(_abc_1014_new_n141_), .B(_abc_1014_new_n133_), .Y(n101));
NAND2X1 NAND2X1_14 ( .A(nRESET_G), .B(_abc_1014_new_n149_), .Y(n36));
NAND2X1 NAND2X1_15 ( .A(nRESET_G), .B(_abc_1014_new_n159_), .Y(n61));
NAND2X1 NAND2X1_16 ( .A(nRESET_G), .B(_abc_1014_new_n164_), .Y(n71));
NAND2X1 NAND2X1_17 ( .A(nRESET_G), .B(_abc_1014_new_n173_), .Y(n86));
NAND2X1 NAND2X1_2 ( .A(_abc_1014_new_n66_), .B(_abc_1014_new_n68_), .Y(_abc_1014_new_n69_));
NAND2X1 NAND2X1_3 ( .A(MAR_REG_0_), .B(MAR_REG_2_), .Y(_abc_1014_new_n90_));
NAND2X1 NAND2X1_4 ( .A(MAR_REG_2_), .B(_abc_1014_new_n82_), .Y(_abc_1014_new_n93_));
NAND2X1 NAND2X1_5 ( .A(_abc_1014_new_n87_), .B(_abc_1014_new_n96_), .Y(_abc_1014_new_n97_));
NAND2X1 NAND2X1_6 ( .A(_abc_1014_new_n82_), .B(_abc_1014_new_n60_), .Y(_abc_1014_new_n98_));
NAND2X1 NAND2X1_7 ( .A(IN_R_REG_2_), .B(_abc_1014_new_n99_), .Y(_abc_1014_new_n100_));
NAND2X1 NAND2X1_8 ( .A(_abc_1014_new_n108_), .B(_abc_1014_new_n110_), .Y(_abc_1014_new_n111_));
NAND2X1 NAND2X1_9 ( .A(_abc_1014_new_n97_), .B(_abc_1014_new_n112_), .Y(_abc_1014_new_n113_));
NAND3X1 NAND3X1_1 ( .A(MAR_REG_1_), .B(MAR_REG_0_), .C(MAR_REG_2_), .Y(_abc_1014_new_n67_));
NAND3X1 NAND3X1_10 ( .A(MAR_REG_2_), .B(_abc_1014_new_n82_), .C(_abc_1014_new_n84_), .Y(_abc_1014_new_n104_));
NAND3X1 NAND3X1_11 ( .A(_abc_1014_new_n67_), .B(_abc_1014_new_n91_), .C(_abc_1014_new_n104_), .Y(_abc_1014_new_n105_));
NAND3X1 NAND3X1_12 ( .A(_abc_1014_new_n109_), .B(_abc_1014_new_n101_), .C(_abc_1014_new_n87_), .Y(_abc_1014_new_n110_));
NAND3X1 NAND3X1_13 ( .A(_abc_1014_new_n93_), .B(_abc_1014_new_n94_), .C(_abc_1014_new_n86_), .Y(_abc_1014_new_n116_));
NAND3X1 NAND3X1_14 ( .A(_abc_1014_new_n121_), .B(_abc_1014_new_n130_), .C(_abc_1014_new_n118_), .Y(_abc_1014_new_n131_));
NAND3X1 NAND3X1_15 ( .A(_abc_1014_new_n82_), .B(MAR_REG_0_), .C(_abc_1014_new_n66_), .Y(_abc_1014_new_n156_));
NAND3X1 NAND3X1_16 ( .A(nRESET_G), .B(_abc_1014_new_n156_), .C(_abc_1014_new_n155_), .Y(n51));
NAND3X1 NAND3X1_2 ( .A(_abc_1014_new_n82_), .B(_abc_1014_new_n84_), .C(_abc_1014_new_n85_), .Y(_abc_1014_new_n86_));
NAND3X1 NAND3X1_3 ( .A(MAR_REG_0_), .B(_abc_1014_new_n82_), .C(_abc_1014_new_n85_), .Y(_abc_1014_new_n87_));
NAND3X1 NAND3X1_4 ( .A(MAR_REG_1_), .B(_abc_1014_new_n84_), .C(_abc_1014_new_n85_), .Y(_abc_1014_new_n91_));
NAND3X1 NAND3X1_5 ( .A(MAR_REG_1_), .B(MAR_REG_0_), .C(_abc_1014_new_n85_), .Y(_abc_1014_new_n94_));
NAND3X1 NAND3X1_6 ( .A(_abc_1014_new_n56_), .B(_abc_1014_new_n93_), .C(_abc_1014_new_n94_), .Y(_abc_1014_new_n95_));
NAND3X1 NAND3X1_7 ( .A(MAR_REG_1_), .B(MAR_REG_2_), .C(_abc_1014_new_n84_), .Y(_abc_1014_new_n101_));
NAND3X1 NAND3X1_8 ( .A(IN_R_REG_1_), .B(_abc_1014_new_n101_), .C(_abc_1014_new_n99_), .Y(_abc_1014_new_n102_));
NAND3X1 NAND3X1_9 ( .A(_abc_1014_new_n98_), .B(_abc_1014_new_n100_), .C(_abc_1014_new_n102_), .Y(_abc_1014_new_n103_));
NOR2X1 NOR2X1_1 ( .A(STATO_REG_1_), .B(_abc_1014_new_n53_), .Y(_abc_1014_new_n54_));
NOR2X1 NOR2X1_2 ( .A(_abc_1014_new_n65_), .B(_abc_1014_new_n53_), .Y(_abc_1014_new_n66_));
NOR2X1 NOR2X1_3 ( .A(START), .B(_abc_1014_new_n67_), .Y(_abc_1014_new_n68_));
NOR2X1 NOR2X1_4 ( .A(MAR_REG_0_), .B(_abc_1014_new_n82_), .Y(_abc_1014_new_n83_));
NOR2X1 NOR2X1_5 ( .A(MAR_REG_1_), .B(MAR_REG_2_), .Y(_abc_1014_new_n88_));
NOR2X1 NOR2X1_6 ( .A(STATO_REG_0_), .B(_abc_1014_new_n65_), .Y(_abc_1014_new_n123_));
NOR2X1 NOR2X1_7 ( .A(MAR_REG_0_), .B(_abc_1014_new_n65_), .Y(_abc_1014_new_n154_));
NOR3X1 NOR3X1_1 ( .A(_abc_1014_new_n124_), .B(_abc_1014_new_n127_), .C(_abc_1014_new_n129_), .Y(_abc_1014_new_n130_));
OAI21X1 OAI21X1_1 ( .A(STATO_REG_1_), .B(_abc_1014_new_n53_), .C(_abc_1014_new_n56_), .Y(_abc_1014_new_n57_));
OAI21X1 OAI21X1_10 ( .A(_abc_1014_new_n82_), .B(_abc_1014_new_n90_), .C(_abc_1014_new_n91_), .Y(_abc_1014_new_n92_));
OAI21X1 OAI21X1_11 ( .A(_abc_1014_new_n95_), .B(_abc_1014_new_n92_), .C(_abc_1014_new_n89_), .Y(_abc_1014_new_n96_));
OAI21X1 OAI21X1_12 ( .A(MAR_REG_1_), .B(_abc_1014_new_n84_), .C(_abc_1014_new_n107_), .Y(_abc_1014_new_n108_));
OAI21X1 OAI21X1_13 ( .A(MAR_REG_2_), .B(_abc_1014_new_n84_), .C(_abc_1014_new_n114_), .Y(_abc_1014_new_n115_));
OAI21X1 OAI21X1_14 ( .A(_abc_1014_new_n88_), .B(_abc_1014_new_n119_), .C(_abc_1014_new_n120_), .Y(_abc_1014_new_n121_));
OAI21X1 OAI21X1_15 ( .A(_abc_1014_new_n122_), .B(_abc_1014_new_n101_), .C(_abc_1014_new_n123_), .Y(_abc_1014_new_n124_));
OAI21X1 OAI21X1_16 ( .A(MAR_REG_2_), .B(_abc_1014_new_n84_), .C(MAR_REG_1_), .Y(_abc_1014_new_n128_));
OAI21X1 OAI21X1_17 ( .A(_abc_1014_new_n106_), .B(_abc_1014_new_n135_), .C(_abc_1014_new_n136_), .Y(n106));
OAI21X1 OAI21X1_18 ( .A(_abc_1014_new_n138_), .B(_abc_1014_new_n135_), .C(_abc_1014_new_n139_), .Y(n111));
OAI21X1 OAI21X1_19 ( .A(_abc_1014_new_n85_), .B(_abc_1014_new_n54_), .C(_abc_1014_new_n144_), .Y(n46));
OAI21X1 OAI21X1_2 ( .A(I_1_), .B(_abc_1014_new_n55_), .C(_abc_1014_new_n57_), .Y(_abc_1014_new_n58_));
OAI21X1 OAI21X1_20 ( .A(_abc_1014_new_n65_), .B(_abc_1014_new_n67_), .C(STATO_REG_0_), .Y(_abc_1014_new_n146_));
OAI21X1 OAI21X1_21 ( .A(_abc_1014_new_n65_), .B(STATO_REG_0_), .C(_abc_1014_new_n147_), .Y(n41));
OAI21X1 OAI21X1_22 ( .A(STATO_REG_1_), .B(STATO_REG_0_), .C(_abc_1014_new_n69_), .Y(_abc_1014_new_n149_));
OAI21X1 OAI21X1_23 ( .A(_abc_1014_new_n84_), .B(_abc_1014_new_n151_), .C(_abc_1014_new_n152_), .Y(n56));
OAI21X1 OAI21X1_24 ( .A(_abc_1014_new_n154_), .B(_abc_1014_new_n146_), .C(MAR_REG_1_), .Y(_abc_1014_new_n155_));
OAI21X1 OAI21X1_25 ( .A(STATO_REG_1_), .B(_abc_1014_new_n53_), .C(_abc_1014_new_n107_), .Y(_abc_1014_new_n158_));
OAI21X1 OAI21X1_26 ( .A(I_7_), .B(_abc_1014_new_n55_), .C(_abc_1014_new_n158_), .Y(_abc_1014_new_n159_));
OAI21X1 OAI21X1_27 ( .A(_abc_1014_new_n114_), .B(_abc_1014_new_n54_), .C(_abc_1014_new_n161_), .Y(n66));
OAI21X1 OAI21X1_28 ( .A(STATO_REG_1_), .B(_abc_1014_new_n53_), .C(_abc_1014_new_n122_), .Y(_abc_1014_new_n163_));
OAI21X1 OAI21X1_29 ( .A(I_5_), .B(_abc_1014_new_n55_), .C(_abc_1014_new_n163_), .Y(_abc_1014_new_n164_));
OAI21X1 OAI21X1_3 ( .A(_abc_1014_new_n60_), .B(_abc_1014_new_n54_), .C(_abc_1014_new_n62_), .Y(n96));
OAI21X1 OAI21X1_30 ( .A(_abc_1014_new_n166_), .B(_abc_1014_new_n55_), .C(_abc_1014_new_n167_), .Y(n76));
OAI21X1 OAI21X1_31 ( .A(_abc_1014_new_n169_), .B(_abc_1014_new_n55_), .C(_abc_1014_new_n170_), .Y(n81));
OAI21X1 OAI21X1_32 ( .A(STATO_REG_1_), .B(_abc_1014_new_n53_), .C(_abc_1014_new_n109_), .Y(_abc_1014_new_n172_));
OAI21X1 OAI21X1_33 ( .A(I_2_), .B(_abc_1014_new_n55_), .C(_abc_1014_new_n172_), .Y(_abc_1014_new_n173_));
OAI21X1 OAI21X1_4 ( .A(_abc_1014_new_n64_), .B(_abc_1014_new_n69_), .C(_abc_1014_new_n70_), .Y(n121));
OAI21X1 OAI21X1_5 ( .A(_abc_1014_new_n72_), .B(_abc_1014_new_n69_), .C(_abc_1014_new_n73_), .Y(n125));
OAI21X1 OAI21X1_6 ( .A(_abc_1014_new_n75_), .B(_abc_1014_new_n69_), .C(_abc_1014_new_n76_), .Y(n129));
OAI21X1 OAI21X1_7 ( .A(_abc_1014_new_n78_), .B(_abc_1014_new_n69_), .C(_abc_1014_new_n79_), .Y(n32));
OAI21X1 OAI21X1_8 ( .A(STATO_REG_1_), .B(_abc_1014_new_n53_), .C(OUT_R_REG_0_), .Y(_abc_1014_new_n81_));
OAI21X1 OAI21X1_9 ( .A(_abc_1014_new_n88_), .B(_abc_1014_new_n83_), .C(IN_R_REG_0_), .Y(_abc_1014_new_n89_));
OAI22X1 OAI22X1_1 ( .A(_abc_1014_new_n114_), .B(_abc_1014_new_n116_), .C(_abc_1014_new_n115_), .D(_abc_1014_new_n105_), .Y(_abc_1014_new_n117_));
OAI22X1 OAI22X1_2 ( .A(_abc_1014_new_n107_), .B(_abc_1014_new_n83_), .C(IN_R_REG_5_), .D(_abc_1014_new_n119_), .Y(_abc_1014_new_n120_));


endmodule