module mc_top(clk_i, rst_i, \wb_data_i[0] , \wb_data_i[1] , \wb_data_i[2] , \wb_data_i[3] , \wb_data_i[4] , \wb_data_i[5] , \wb_data_i[6] , \wb_data_i[7] , \wb_data_i[8] , \wb_data_i[9] , \wb_data_i[10] , \wb_data_i[11] , \wb_data_i[12] , \wb_data_i[13] , \wb_data_i[14] , \wb_data_i[15] , \wb_data_i[16] , \wb_data_i[17] , \wb_data_i[18] , \wb_data_i[19] , \wb_data_i[20] , \wb_data_i[21] , \wb_data_i[22] , \wb_data_i[23] , \wb_data_i[24] , \wb_data_i[25] , \wb_data_i[26] , \wb_data_i[27] , \wb_data_i[28] , \wb_data_i[29] , \wb_data_i[30] , \wb_data_i[31] , \wb_addr_i[0] , \wb_addr_i[1] , \wb_addr_i[2] , \wb_addr_i[3] , \wb_addr_i[4] , \wb_addr_i[5] , \wb_addr_i[6] , \wb_addr_i[7] , \wb_addr_i[8] , \wb_addr_i[9] , \wb_addr_i[10] , \wb_addr_i[11] , \wb_addr_i[12] , \wb_addr_i[13] , \wb_addr_i[14] , \wb_addr_i[15] , \wb_addr_i[16] , \wb_addr_i[17] , \wb_addr_i[18] , \wb_addr_i[19] , \wb_addr_i[20] , \wb_addr_i[21] , \wb_addr_i[22] , \wb_addr_i[23] , \wb_addr_i[24] , \wb_addr_i[25] , \wb_addr_i[26] , \wb_addr_i[27] , \wb_addr_i[28] , \wb_addr_i[29] , \wb_addr_i[30] , \wb_addr_i[31] , \wb_sel_i[0] , \wb_sel_i[1] , \wb_sel_i[2] , \wb_sel_i[3] , wb_we_i, wb_cyc_i, wb_stb_i, susp_req_i, resume_req_i, mc_clk_i, mc_br_pad_i, mc_ack_pad_i, \mc_data_pad_i[0] , \mc_data_pad_i[1] , \mc_data_pad_i[2] , \mc_data_pad_i[3] , \mc_data_pad_i[4] , \mc_data_pad_i[5] , \mc_data_pad_i[6] , \mc_data_pad_i[7] , \mc_data_pad_i[8] , \mc_data_pad_i[9] , \mc_data_pad_i[10] , \mc_data_pad_i[11] , \mc_data_pad_i[12] , \mc_data_pad_i[13] , \mc_data_pad_i[14] , \mc_data_pad_i[15] , \mc_data_pad_i[16] , \mc_data_pad_i[17] , \mc_data_pad_i[18] , \mc_data_pad_i[19] , \mc_data_pad_i[20] , \mc_data_pad_i[21] , \mc_data_pad_i[22] , \mc_data_pad_i[23] , \mc_data_pad_i[24] , \mc_data_pad_i[25] , \mc_data_pad_i[26] , \mc_data_pad_i[27] , \mc_data_pad_i[28] , \mc_data_pad_i[29] , \mc_data_pad_i[30] , \mc_data_pad_i[31] , \mc_dp_pad_i[0] , \mc_dp_pad_i[1] , \mc_dp_pad_i[2] , \mc_dp_pad_i[3] , mc_sts_pad_i, \wb_data_o[0] , \wb_data_o[1] , \wb_data_o[2] , \wb_data_o[3] , \wb_data_o[4] , \wb_data_o[5] , \wb_data_o[6] , \wb_data_o[7] , \wb_data_o[8] , \wb_data_o[9] , \wb_data_o[10] , \wb_data_o[11] , \wb_data_o[12] , \wb_data_o[13] , \wb_data_o[14] , \wb_data_o[15] , \wb_data_o[16] , \wb_data_o[17] , \wb_data_o[18] , \wb_data_o[19] , \wb_data_o[20] , \wb_data_o[21] , \wb_data_o[22] , \wb_data_o[23] , \wb_data_o[24] , \wb_data_o[25] , \wb_data_o[26] , \wb_data_o[27] , \wb_data_o[28] , \wb_data_o[29] , \wb_data_o[30] , \wb_data_o[31] , wb_ack_o, wb_err_o, suspended_o, \poc_o[0] , \poc_o[1] , \poc_o[2] , \poc_o[3] , \poc_o[4] , \poc_o[5] , \poc_o[6] , \poc_o[7] , \poc_o[8] , \poc_o[9] , \poc_o[10] , \poc_o[11] , \poc_o[12] , \poc_o[13] , \poc_o[14] , \poc_o[15] , \poc_o[16] , \poc_o[17] , \poc_o[18] , \poc_o[19] , \poc_o[20] , \poc_o[21] , \poc_o[22] , \poc_o[23] , \poc_o[24] , \poc_o[25] , \poc_o[26] , \poc_o[27] , \poc_o[28] , \poc_o[29] , \poc_o[30] , \poc_o[31] , mc_bg_pad_o, \mc_addr_pad_o[0] , \mc_addr_pad_o[1] , \mc_addr_pad_o[2] , \mc_addr_pad_o[3] , \mc_addr_pad_o[4] , \mc_addr_pad_o[5] , \mc_addr_pad_o[6] , \mc_addr_pad_o[7] , \mc_addr_pad_o[8] , \mc_addr_pad_o[9] , \mc_addr_pad_o[10] , \mc_addr_pad_o[11] , \mc_addr_pad_o[12] , \mc_addr_pad_o[13] , \mc_addr_pad_o[14] , \mc_addr_pad_o[15] , \mc_addr_pad_o[16] , \mc_addr_pad_o[17] , \mc_addr_pad_o[18] , \mc_addr_pad_o[19] , \mc_addr_pad_o[20] , \mc_addr_pad_o[21] , \mc_addr_pad_o[22] , \mc_addr_pad_o[23] , \mc_data_pad_o[0] , \mc_data_pad_o[1] , \mc_data_pad_o[2] , \mc_data_pad_o[3] , \mc_data_pad_o[4] , \mc_data_pad_o[5] , \mc_data_pad_o[6] , \mc_data_pad_o[7] , \mc_data_pad_o[8] , \mc_data_pad_o[9] , \mc_data_pad_o[10] , \mc_data_pad_o[11] , \mc_data_pad_o[12] , \mc_data_pad_o[13] , \mc_data_pad_o[14] , \mc_data_pad_o[15] , \mc_data_pad_o[16] , \mc_data_pad_o[17] , \mc_data_pad_o[18] , \mc_data_pad_o[19] , \mc_data_pad_o[20] , \mc_data_pad_o[21] , \mc_data_pad_o[22] , \mc_data_pad_o[23] , \mc_data_pad_o[24] , \mc_data_pad_o[25] , \mc_data_pad_o[26] , \mc_data_pad_o[27] , \mc_data_pad_o[28] , \mc_data_pad_o[29] , \mc_data_pad_o[30] , \mc_data_pad_o[31] , \mc_dp_pad_o[0] , \mc_dp_pad_o[1] , \mc_dp_pad_o[2] , \mc_dp_pad_o[3] , mc_doe_pad_doe_o, \mc_dqm_pad_o[0] , \mc_dqm_pad_o[1] , \mc_dqm_pad_o[2] , \mc_dqm_pad_o[3] , mc_oe_pad_o_, mc_we_pad_o_, mc_cas_pad_o_, mc_ras_pad_o_, mc_cke_pad_o_, \mc_cs_pad_o_[0] , \mc_cs_pad_o_[1] , \mc_cs_pad_o_[2] , \mc_cs_pad_o_[3] , \mc_cs_pad_o_[4] , \mc_cs_pad_o_[5] , \mc_cs_pad_o_[6] , \mc_cs_pad_o_[7] , mc_rp_pad_o_, mc_vpen_pad_o, mc_adsc_pad_o_, mc_adv_pad_o_, mc_zz_pad_o, mc_coe_pad_coe_o);

wire _abc_85006_new_n237_; 
wire _abc_85006_new_n238_; 
wire _abc_85006_new_n239_; 
wire _abc_85006_new_n240_; 
wire _abc_85006_new_n240__bF_buf0; 
wire _abc_85006_new_n240__bF_buf1; 
wire _abc_85006_new_n240__bF_buf2; 
wire _abc_85006_new_n240__bF_buf3; 
wire _abc_85006_new_n240__bF_buf4; 
wire _abc_85006_new_n240__bF_buf5; 
wire _abc_85006_new_n241_; 
wire _abc_85006_new_n242_; 
wire _abc_85006_new_n243_; 
wire _abc_85006_new_n244_; 
wire _abc_85006_new_n245_; 
wire _abc_85006_new_n246_; 
wire _abc_85006_new_n248_; 
wire _abc_85006_new_n249_; 
wire _abc_85006_new_n250_; 
wire _abc_85006_new_n251_; 
wire _abc_85006_new_n252_; 
wire _abc_85006_new_n254_; 
wire _abc_85006_new_n255_; 
wire _abc_85006_new_n256_; 
wire _abc_85006_new_n257_; 
wire _abc_85006_new_n258_; 
wire _abc_85006_new_n260_; 
wire _abc_85006_new_n261_; 
wire _abc_85006_new_n262_; 
wire _abc_85006_new_n263_; 
wire _abc_85006_new_n264_; 
wire _abc_85006_new_n266_; 
wire _abc_85006_new_n267_; 
wire _abc_85006_new_n268_; 
wire _abc_85006_new_n269_; 
wire _abc_85006_new_n270_; 
wire _abc_85006_new_n272_; 
wire _abc_85006_new_n273_; 
wire _abc_85006_new_n274_; 
wire _abc_85006_new_n275_; 
wire _abc_85006_new_n276_; 
wire _abc_85006_new_n278_; 
wire _abc_85006_new_n279_; 
wire _abc_85006_new_n280_; 
wire _abc_85006_new_n281_; 
wire _abc_85006_new_n282_; 
wire _abc_85006_new_n284_; 
wire _abc_85006_new_n285_; 
wire _abc_85006_new_n286_; 
wire _abc_85006_new_n287_; 
wire _abc_85006_new_n288_; 
wire _abc_85006_new_n290_; 
wire _abc_85006_new_n291_; 
wire _abc_85006_new_n293_; 
wire _abc_85006_new_n294_; 
wire _abc_85006_new_n296_; 
wire _abc_85006_new_n297_; 
wire _abc_85006_new_n299_; 
wire _abc_85006_new_n300_; 
wire _abc_85006_new_n302_; 
wire _abc_85006_new_n303_; 
wire _abc_85006_new_n305_; 
wire _abc_85006_new_n306_; 
wire _abc_85006_new_n308_; 
wire _abc_85006_new_n309_; 
wire _abc_85006_new_n311_; 
wire _abc_85006_new_n312_; 
wire _abc_85006_new_n314_; 
wire _abc_85006_new_n315_; 
wire _abc_85006_new_n317_; 
wire _abc_85006_new_n318_; 
wire _abc_85006_new_n320_; 
wire _abc_85006_new_n321_; 
wire _abc_85006_new_n323_; 
wire _abc_85006_new_n324_; 
wire _abc_85006_new_n326_; 
wire _abc_85006_new_n327_; 
wire _abc_85006_new_n329_; 
wire _abc_85006_new_n330_; 
wire _abc_85006_new_n332_; 
wire _abc_85006_new_n333_; 
wire _abc_85006_new_n335_; 
wire _abc_85006_new_n336_; 
wire _abc_85006_new_n338_; 
wire _abc_85006_new_n339_; 
wire _abc_85006_new_n341_; 
wire _abc_85006_new_n342_; 
wire _abc_85006_new_n344_; 
wire _abc_85006_new_n345_; 
wire _abc_85006_new_n347_; 
wire _abc_85006_new_n348_; 
wire _abc_85006_new_n350_; 
wire _abc_85006_new_n351_; 
wire _abc_85006_new_n353_; 
wire _abc_85006_new_n354_; 
wire _abc_85006_new_n356_; 
wire _abc_85006_new_n357_; 
wire _abc_85006_new_n359_; 
wire _abc_85006_new_n360_; 
wire _abc_85006_new_n362_; 
wire _abc_85006_new_n363_; 
wire _abc_85006_new_n365_; 
wire _abc_85006_new_n366_; 
wire _abc_85006_new_n368_; 
wire _abc_85006_new_n369_; 
wire _abc_85006_new_n371_; 
wire _abc_85006_new_n372_; 
wire _abc_85006_new_n389_; 
wire _abc_85006_new_n390_; 
wire _abc_85006_new_n392_; 
wire _abc_85006_new_n393_; 
wire _abc_85006_new_n395_; 
wire _abc_85006_new_n396_; 
wire _abc_85006_new_n398_; 
wire _abc_85006_new_n399_; 
wire _abc_85006_new_n401_; 
wire _abc_85006_new_n402_; 
wire _abc_85006_new_n404_; 
wire _abc_85006_new_n405_; 
wire _abc_85006_new_n407_; 
wire _abc_85006_new_n408_; 
wire _abc_85006_new_n413_; 
wire _abc_85006_new_n414_; 
wire _abc_85006_new_n416_; 
wire _abc_85006_new_n417_; 
wire _abc_85006_new_n482_; 
wire _abc_85006_new_n483_; 
wire _abc_85006_new_n484_; 
wire _auto_iopadmap_cc_368_execute_85420_0_; 
wire _auto_iopadmap_cc_368_execute_85420_10_; 
wire _auto_iopadmap_cc_368_execute_85420_11_; 
wire _auto_iopadmap_cc_368_execute_85420_12_; 
wire _auto_iopadmap_cc_368_execute_85420_13_; 
wire _auto_iopadmap_cc_368_execute_85420_14_; 
wire _auto_iopadmap_cc_368_execute_85420_15_; 
wire _auto_iopadmap_cc_368_execute_85420_16_; 
wire _auto_iopadmap_cc_368_execute_85420_17_; 
wire _auto_iopadmap_cc_368_execute_85420_18_; 
wire _auto_iopadmap_cc_368_execute_85420_19_; 
wire _auto_iopadmap_cc_368_execute_85420_1_; 
wire _auto_iopadmap_cc_368_execute_85420_20_; 
wire _auto_iopadmap_cc_368_execute_85420_21_; 
wire _auto_iopadmap_cc_368_execute_85420_22_; 
wire _auto_iopadmap_cc_368_execute_85420_23_; 
wire _auto_iopadmap_cc_368_execute_85420_2_; 
wire _auto_iopadmap_cc_368_execute_85420_3_; 
wire _auto_iopadmap_cc_368_execute_85420_4_; 
wire _auto_iopadmap_cc_368_execute_85420_5_; 
wire _auto_iopadmap_cc_368_execute_85420_6_; 
wire _auto_iopadmap_cc_368_execute_85420_7_; 
wire _auto_iopadmap_cc_368_execute_85420_8_; 
wire _auto_iopadmap_cc_368_execute_85420_9_; 
wire _auto_iopadmap_cc_368_execute_85445; 
wire _auto_iopadmap_cc_368_execute_85447; 
wire _auto_iopadmap_cc_368_execute_85449; 
wire _auto_iopadmap_cc_368_execute_85451; 
wire _auto_iopadmap_cc_368_execute_85453; 
wire _auto_iopadmap_cc_368_execute_85455; 
wire _auto_iopadmap_cc_368_execute_85457_0_; 
wire _auto_iopadmap_cc_368_execute_85457_1_; 
wire _auto_iopadmap_cc_368_execute_85457_2_; 
wire _auto_iopadmap_cc_368_execute_85457_3_; 
wire _auto_iopadmap_cc_368_execute_85457_4_; 
wire _auto_iopadmap_cc_368_execute_85457_5_; 
wire _auto_iopadmap_cc_368_execute_85457_6_; 
wire _auto_iopadmap_cc_368_execute_85457_7_; 
wire _auto_iopadmap_cc_368_execute_85466_0_; 
wire _auto_iopadmap_cc_368_execute_85466_10_; 
wire _auto_iopadmap_cc_368_execute_85466_11_; 
wire _auto_iopadmap_cc_368_execute_85466_12_; 
wire _auto_iopadmap_cc_368_execute_85466_13_; 
wire _auto_iopadmap_cc_368_execute_85466_14_; 
wire _auto_iopadmap_cc_368_execute_85466_15_; 
wire _auto_iopadmap_cc_368_execute_85466_16_; 
wire _auto_iopadmap_cc_368_execute_85466_17_; 
wire _auto_iopadmap_cc_368_execute_85466_18_; 
wire _auto_iopadmap_cc_368_execute_85466_19_; 
wire _auto_iopadmap_cc_368_execute_85466_1_; 
wire _auto_iopadmap_cc_368_execute_85466_20_; 
wire _auto_iopadmap_cc_368_execute_85466_21_; 
wire _auto_iopadmap_cc_368_execute_85466_22_; 
wire _auto_iopadmap_cc_368_execute_85466_23_; 
wire _auto_iopadmap_cc_368_execute_85466_24_; 
wire _auto_iopadmap_cc_368_execute_85466_25_; 
wire _auto_iopadmap_cc_368_execute_85466_26_; 
wire _auto_iopadmap_cc_368_execute_85466_27_; 
wire _auto_iopadmap_cc_368_execute_85466_28_; 
wire _auto_iopadmap_cc_368_execute_85466_29_; 
wire _auto_iopadmap_cc_368_execute_85466_2_; 
wire _auto_iopadmap_cc_368_execute_85466_30_; 
wire _auto_iopadmap_cc_368_execute_85466_31_; 
wire _auto_iopadmap_cc_368_execute_85466_3_; 
wire _auto_iopadmap_cc_368_execute_85466_4_; 
wire _auto_iopadmap_cc_368_execute_85466_5_; 
wire _auto_iopadmap_cc_368_execute_85466_6_; 
wire _auto_iopadmap_cc_368_execute_85466_7_; 
wire _auto_iopadmap_cc_368_execute_85466_8_; 
wire _auto_iopadmap_cc_368_execute_85466_9_; 
wire _auto_iopadmap_cc_368_execute_85499; 
wire _auto_iopadmap_cc_368_execute_85501_0_; 
wire _auto_iopadmap_cc_368_execute_85501_1_; 
wire _auto_iopadmap_cc_368_execute_85501_2_; 
wire _auto_iopadmap_cc_368_execute_85501_3_; 
wire _auto_iopadmap_cc_368_execute_85506_0_; 
wire _auto_iopadmap_cc_368_execute_85506_1_; 
wire _auto_iopadmap_cc_368_execute_85506_2_; 
wire _auto_iopadmap_cc_368_execute_85506_3_; 
wire _auto_iopadmap_cc_368_execute_85511; 
wire _auto_iopadmap_cc_368_execute_85513; 
wire _auto_iopadmap_cc_368_execute_85515; 
wire _auto_iopadmap_cc_368_execute_85519; 
wire _auto_iopadmap_cc_368_execute_85521; 
wire _auto_iopadmap_cc_368_execute_85523_0_; 
wire _auto_iopadmap_cc_368_execute_85523_10_; 
wire _auto_iopadmap_cc_368_execute_85523_11_; 
wire _auto_iopadmap_cc_368_execute_85523_12_; 
wire _auto_iopadmap_cc_368_execute_85523_13_; 
wire _auto_iopadmap_cc_368_execute_85523_14_; 
wire _auto_iopadmap_cc_368_execute_85523_15_; 
wire _auto_iopadmap_cc_368_execute_85523_16_; 
wire _auto_iopadmap_cc_368_execute_85523_17_; 
wire _auto_iopadmap_cc_368_execute_85523_18_; 
wire _auto_iopadmap_cc_368_execute_85523_19_; 
wire _auto_iopadmap_cc_368_execute_85523_1_; 
wire _auto_iopadmap_cc_368_execute_85523_20_; 
wire _auto_iopadmap_cc_368_execute_85523_21_; 
wire _auto_iopadmap_cc_368_execute_85523_22_; 
wire _auto_iopadmap_cc_368_execute_85523_23_; 
wire _auto_iopadmap_cc_368_execute_85523_24_; 
wire _auto_iopadmap_cc_368_execute_85523_25_; 
wire _auto_iopadmap_cc_368_execute_85523_26_; 
wire _auto_iopadmap_cc_368_execute_85523_27_; 
wire _auto_iopadmap_cc_368_execute_85523_28_; 
wire _auto_iopadmap_cc_368_execute_85523_29_; 
wire _auto_iopadmap_cc_368_execute_85523_2_; 
wire _auto_iopadmap_cc_368_execute_85523_30_; 
wire _auto_iopadmap_cc_368_execute_85523_31_; 
wire _auto_iopadmap_cc_368_execute_85523_3_; 
wire _auto_iopadmap_cc_368_execute_85523_4_; 
wire _auto_iopadmap_cc_368_execute_85523_5_; 
wire _auto_iopadmap_cc_368_execute_85523_6_; 
wire _auto_iopadmap_cc_368_execute_85523_7_; 
wire _auto_iopadmap_cc_368_execute_85523_8_; 
wire _auto_iopadmap_cc_368_execute_85523_9_; 
wire _auto_iopadmap_cc_368_execute_85556; 
wire _auto_iopadmap_cc_368_execute_85558; 
wire _auto_iopadmap_cc_368_execute_85560_0_; 
wire _auto_iopadmap_cc_368_execute_85560_10_; 
wire _auto_iopadmap_cc_368_execute_85560_11_; 
wire _auto_iopadmap_cc_368_execute_85560_12_; 
wire _auto_iopadmap_cc_368_execute_85560_13_; 
wire _auto_iopadmap_cc_368_execute_85560_14_; 
wire _auto_iopadmap_cc_368_execute_85560_15_; 
wire _auto_iopadmap_cc_368_execute_85560_16_; 
wire _auto_iopadmap_cc_368_execute_85560_17_; 
wire _auto_iopadmap_cc_368_execute_85560_18_; 
wire _auto_iopadmap_cc_368_execute_85560_19_; 
wire _auto_iopadmap_cc_368_execute_85560_1_; 
wire _auto_iopadmap_cc_368_execute_85560_20_; 
wire _auto_iopadmap_cc_368_execute_85560_21_; 
wire _auto_iopadmap_cc_368_execute_85560_22_; 
wire _auto_iopadmap_cc_368_execute_85560_23_; 
wire _auto_iopadmap_cc_368_execute_85560_24_; 
wire _auto_iopadmap_cc_368_execute_85560_25_; 
wire _auto_iopadmap_cc_368_execute_85560_26_; 
wire _auto_iopadmap_cc_368_execute_85560_27_; 
wire _auto_iopadmap_cc_368_execute_85560_28_; 
wire _auto_iopadmap_cc_368_execute_85560_29_; 
wire _auto_iopadmap_cc_368_execute_85560_2_; 
wire _auto_iopadmap_cc_368_execute_85560_30_; 
wire _auto_iopadmap_cc_368_execute_85560_31_; 
wire _auto_iopadmap_cc_368_execute_85560_3_; 
wire _auto_iopadmap_cc_368_execute_85560_4_; 
wire _auto_iopadmap_cc_368_execute_85560_5_; 
wire _auto_iopadmap_cc_368_execute_85560_6_; 
wire _auto_iopadmap_cc_368_execute_85560_7_; 
wire _auto_iopadmap_cc_368_execute_85560_8_; 
wire _auto_iopadmap_cc_368_execute_85560_9_; 
wire _auto_iopadmap_cc_368_execute_85593; 
wire bank_adr_0_; 
wire bank_adr_1_; 
wire bank_clr; 
wire bank_clr_all; 
wire bank_open; 
wire bank_set; 
wire cas_; 
input clk_i;
wire clk_i_bF_buf0; 
wire clk_i_bF_buf1; 
wire clk_i_bF_buf10; 
wire clk_i_bF_buf11; 
wire clk_i_bF_buf12; 
wire clk_i_bF_buf13; 
wire clk_i_bF_buf14; 
wire clk_i_bF_buf15; 
wire clk_i_bF_buf16; 
wire clk_i_bF_buf17; 
wire clk_i_bF_buf18; 
wire clk_i_bF_buf19; 
wire clk_i_bF_buf2; 
wire clk_i_bF_buf20; 
wire clk_i_bF_buf21; 
wire clk_i_bF_buf22; 
wire clk_i_bF_buf23; 
wire clk_i_bF_buf24; 
wire clk_i_bF_buf25; 
wire clk_i_bF_buf26; 
wire clk_i_bF_buf27; 
wire clk_i_bF_buf28; 
wire clk_i_bF_buf29; 
wire clk_i_bF_buf3; 
wire clk_i_bF_buf30; 
wire clk_i_bF_buf31; 
wire clk_i_bF_buf32; 
wire clk_i_bF_buf33; 
wire clk_i_bF_buf34; 
wire clk_i_bF_buf35; 
wire clk_i_bF_buf36; 
wire clk_i_bF_buf37; 
wire clk_i_bF_buf38; 
wire clk_i_bF_buf39; 
wire clk_i_bF_buf4; 
wire clk_i_bF_buf40; 
wire clk_i_bF_buf41; 
wire clk_i_bF_buf42; 
wire clk_i_bF_buf43; 
wire clk_i_bF_buf44; 
wire clk_i_bF_buf45; 
wire clk_i_bF_buf46; 
wire clk_i_bF_buf47; 
wire clk_i_bF_buf48; 
wire clk_i_bF_buf49; 
wire clk_i_bF_buf5; 
wire clk_i_bF_buf50; 
wire clk_i_bF_buf51; 
wire clk_i_bF_buf52; 
wire clk_i_bF_buf53; 
wire clk_i_bF_buf54; 
wire clk_i_bF_buf55; 
wire clk_i_bF_buf56; 
wire clk_i_bF_buf57; 
wire clk_i_bF_buf58; 
wire clk_i_bF_buf59; 
wire clk_i_bF_buf6; 
wire clk_i_bF_buf60; 
wire clk_i_bF_buf61; 
wire clk_i_bF_buf62; 
wire clk_i_bF_buf63; 
wire clk_i_bF_buf64; 
wire clk_i_bF_buf65; 
wire clk_i_bF_buf66; 
wire clk_i_bF_buf67; 
wire clk_i_bF_buf68; 
wire clk_i_bF_buf69; 
wire clk_i_bF_buf7; 
wire clk_i_bF_buf70; 
wire clk_i_bF_buf71; 
wire clk_i_bF_buf72; 
wire clk_i_bF_buf73; 
wire clk_i_bF_buf74; 
wire clk_i_bF_buf75; 
wire clk_i_bF_buf76; 
wire clk_i_bF_buf77; 
wire clk_i_bF_buf78; 
wire clk_i_bF_buf79; 
wire clk_i_bF_buf8; 
wire clk_i_bF_buf80; 
wire clk_i_bF_buf81; 
wire clk_i_bF_buf82; 
wire clk_i_bF_buf83; 
wire clk_i_bF_buf84; 
wire clk_i_bF_buf85; 
wire clk_i_bF_buf86; 
wire clk_i_bF_buf87; 
wire clk_i_bF_buf88; 
wire clk_i_bF_buf89; 
wire clk_i_bF_buf9; 
wire clk_i_bF_buf90; 
wire clk_i_bF_buf91; 
wire clk_i_bF_buf92; 
wire clk_i_bF_buf93; 
wire clk_i_bF_buf94; 
wire clk_i_bF_buf95; 
wire clk_i_bF_buf96; 
wire clk_i_hier0_bF_buf0; 
wire clk_i_hier0_bF_buf1; 
wire clk_i_hier0_bF_buf2; 
wire clk_i_hier0_bF_buf3; 
wire clk_i_hier0_bF_buf4; 
wire clk_i_hier0_bF_buf5; 
wire clk_i_hier0_bF_buf6; 
wire clk_i_hier0_bF_buf7; 
wire clk_i_hier0_bF_buf8; 
wire cmd_a10; 
wire cs_0_; 
wire cs_1_; 
wire cs_2_; 
wire cs_3_; 
wire cs_4_; 
wire cs_5_; 
wire cs_6_; 
wire cs_7_; 
wire cs_en; 
wire cs_le; 
wire cs_le_bF_buf0; 
wire cs_le_bF_buf1; 
wire cs_le_bF_buf2; 
wire cs_le_bF_buf3; 
wire cs_le_bF_buf4; 
wire cs_le_d; 
wire cs_need_rfr_0_; 
wire cs_need_rfr_1_; 
wire cs_need_rfr_2_; 
wire cs_need_rfr_3_; 
wire cs_need_rfr_4_; 
wire cs_need_rfr_5_; 
wire cs_need_rfr_6_; 
wire cs_need_rfr_7_; 
wire csc_10_; 
wire csc_1_; 
wire csc_2_; 
wire csc_3_; 
wire csc_4_; 
wire csc_5_; 
wire csc_5_bF_buf0_; 
wire csc_5_bF_buf1_; 
wire csc_5_bF_buf2_; 
wire csc_5_bF_buf3_; 
wire csc_5_bF_buf4_; 
wire csc_6_; 
wire csc_7_; 
wire csc_9_; 
wire csc_s_1_; 
wire csc_s_2_; 
wire csc_s_3_; 
wire csc_s_4_; 
wire csc_s_5_; 
wire csc_s_6_; 
wire csc_s_7_; 
wire data_oe; 
wire dv; 
wire err; 
wire fs; 
wire init_ack; 
wire init_req; 
wire lmr_ack; 
wire lmr_req; 
wire lmr_sel; 
wire lmr_sel_bF_buf0; 
wire lmr_sel_bF_buf1; 
wire lmr_sel_bF_buf2; 
wire lmr_sel_bF_buf3; 
wire lmr_sel_bF_buf4; 
wire lmr_sel_bF_buf5; 
wire lmr_sel_bF_buf6; 
input mc_ack_pad_i;
wire mc_ack_r; 
wire mc_addr_d_0_; 
wire mc_addr_d_10_; 
wire mc_addr_d_11_; 
wire mc_addr_d_12_; 
wire mc_addr_d_13_; 
wire mc_addr_d_14_; 
wire mc_addr_d_15_; 
wire mc_addr_d_16_; 
wire mc_addr_d_17_; 
wire mc_addr_d_18_; 
wire mc_addr_d_19_; 
wire mc_addr_d_1_; 
wire mc_addr_d_20_; 
wire mc_addr_d_21_; 
wire mc_addr_d_22_; 
wire mc_addr_d_23_; 
wire mc_addr_d_2_; 
wire mc_addr_d_3_; 
wire mc_addr_d_4_; 
wire mc_addr_d_5_; 
wire mc_addr_d_6_; 
wire mc_addr_d_7_; 
wire mc_addr_d_8_; 
wire mc_addr_d_9_; 
output \mc_addr_pad_o[0] ;
output \mc_addr_pad_o[10] ;
output \mc_addr_pad_o[11] ;
output \mc_addr_pad_o[12] ;
output \mc_addr_pad_o[13] ;
output \mc_addr_pad_o[14] ;
output \mc_addr_pad_o[15] ;
output \mc_addr_pad_o[16] ;
output \mc_addr_pad_o[17] ;
output \mc_addr_pad_o[18] ;
output \mc_addr_pad_o[19] ;
output \mc_addr_pad_o[1] ;
output \mc_addr_pad_o[20] ;
output \mc_addr_pad_o[21] ;
output \mc_addr_pad_o[22] ;
output \mc_addr_pad_o[23] ;
output \mc_addr_pad_o[2] ;
output \mc_addr_pad_o[3] ;
output \mc_addr_pad_o[4] ;
output \mc_addr_pad_o[5] ;
output \mc_addr_pad_o[6] ;
output \mc_addr_pad_o[7] ;
output \mc_addr_pad_o[8] ;
output \mc_addr_pad_o[9] ;
wire mc_adsc_d; 
output mc_adsc_pad_o_;
wire mc_adv_d; 
output mc_adv_pad_o_;
wire mc_bg_d; 
output mc_bg_pad_o;
input mc_br_pad_i;
wire mc_br_r; 
wire mc_c_oe_d; 
output mc_cas_pad_o_;
output mc_cke_pad_o_;
input mc_clk_i;
wire mc_clk_i_bF_buf0; 
wire mc_clk_i_bF_buf1; 
wire mc_clk_i_bF_buf10; 
wire mc_clk_i_bF_buf2; 
wire mc_clk_i_bF_buf3; 
wire mc_clk_i_bF_buf4; 
wire mc_clk_i_bF_buf5; 
wire mc_clk_i_bF_buf6; 
wire mc_clk_i_bF_buf7; 
wire mc_clk_i_bF_buf8; 
wire mc_clk_i_bF_buf9; 
output mc_coe_pad_coe_o;
output \mc_cs_pad_o_[0] ;
output \mc_cs_pad_o_[1] ;
output \mc_cs_pad_o_[2] ;
output \mc_cs_pad_o_[3] ;
output \mc_cs_pad_o_[4] ;
output \mc_cs_pad_o_[5] ;
output \mc_cs_pad_o_[6] ;
output \mc_cs_pad_o_[7] ;
wire mc_data_ir_0_; 
wire mc_data_ir_10_; 
wire mc_data_ir_11_; 
wire mc_data_ir_12_; 
wire mc_data_ir_13_; 
wire mc_data_ir_14_; 
wire mc_data_ir_15_; 
wire mc_data_ir_16_; 
wire mc_data_ir_17_; 
wire mc_data_ir_18_; 
wire mc_data_ir_19_; 
wire mc_data_ir_1_; 
wire mc_data_ir_20_; 
wire mc_data_ir_21_; 
wire mc_data_ir_22_; 
wire mc_data_ir_23_; 
wire mc_data_ir_24_; 
wire mc_data_ir_25_; 
wire mc_data_ir_26_; 
wire mc_data_ir_27_; 
wire mc_data_ir_28_; 
wire mc_data_ir_29_; 
wire mc_data_ir_2_; 
wire mc_data_ir_30_; 
wire mc_data_ir_31_; 
wire mc_data_ir_32_; 
wire mc_data_ir_33_; 
wire mc_data_ir_34_; 
wire mc_data_ir_35_; 
wire mc_data_ir_3_; 
wire mc_data_ir_4_; 
wire mc_data_ir_5_; 
wire mc_data_ir_6_; 
wire mc_data_ir_7_; 
wire mc_data_ir_8_; 
wire mc_data_ir_9_; 
wire mc_data_od_0_; 
wire mc_data_od_10_; 
wire mc_data_od_11_; 
wire mc_data_od_12_; 
wire mc_data_od_13_; 
wire mc_data_od_14_; 
wire mc_data_od_15_; 
wire mc_data_od_16_; 
wire mc_data_od_17_; 
wire mc_data_od_18_; 
wire mc_data_od_19_; 
wire mc_data_od_1_; 
wire mc_data_od_20_; 
wire mc_data_od_21_; 
wire mc_data_od_22_; 
wire mc_data_od_23_; 
wire mc_data_od_24_; 
wire mc_data_od_25_; 
wire mc_data_od_26_; 
wire mc_data_od_27_; 
wire mc_data_od_28_; 
wire mc_data_od_29_; 
wire mc_data_od_2_; 
wire mc_data_od_30_; 
wire mc_data_od_31_; 
wire mc_data_od_3_; 
wire mc_data_od_4_; 
wire mc_data_od_5_; 
wire mc_data_od_6_; 
wire mc_data_od_7_; 
wire mc_data_od_8_; 
wire mc_data_od_9_; 
input \mc_data_pad_i[0] ;
input \mc_data_pad_i[10] ;
input \mc_data_pad_i[11] ;
input \mc_data_pad_i[12] ;
input \mc_data_pad_i[13] ;
input \mc_data_pad_i[14] ;
input \mc_data_pad_i[15] ;
input \mc_data_pad_i[16] ;
input \mc_data_pad_i[17] ;
input \mc_data_pad_i[18] ;
input \mc_data_pad_i[19] ;
input \mc_data_pad_i[1] ;
input \mc_data_pad_i[20] ;
input \mc_data_pad_i[21] ;
input \mc_data_pad_i[22] ;
input \mc_data_pad_i[23] ;
input \mc_data_pad_i[24] ;
input \mc_data_pad_i[25] ;
input \mc_data_pad_i[26] ;
input \mc_data_pad_i[27] ;
input \mc_data_pad_i[28] ;
input \mc_data_pad_i[29] ;
input \mc_data_pad_i[2] ;
input \mc_data_pad_i[30] ;
input \mc_data_pad_i[31] ;
input \mc_data_pad_i[3] ;
input \mc_data_pad_i[4] ;
input \mc_data_pad_i[5] ;
input \mc_data_pad_i[6] ;
input \mc_data_pad_i[7] ;
input \mc_data_pad_i[8] ;
input \mc_data_pad_i[9] ;
output \mc_data_pad_o[0] ;
output \mc_data_pad_o[10] ;
output \mc_data_pad_o[11] ;
output \mc_data_pad_o[12] ;
output \mc_data_pad_o[13] ;
output \mc_data_pad_o[14] ;
output \mc_data_pad_o[15] ;
output \mc_data_pad_o[16] ;
output \mc_data_pad_o[17] ;
output \mc_data_pad_o[18] ;
output \mc_data_pad_o[19] ;
output \mc_data_pad_o[1] ;
output \mc_data_pad_o[20] ;
output \mc_data_pad_o[21] ;
output \mc_data_pad_o[22] ;
output \mc_data_pad_o[23] ;
output \mc_data_pad_o[24] ;
output \mc_data_pad_o[25] ;
output \mc_data_pad_o[26] ;
output \mc_data_pad_o[27] ;
output \mc_data_pad_o[28] ;
output \mc_data_pad_o[29] ;
output \mc_data_pad_o[2] ;
output \mc_data_pad_o[30] ;
output \mc_data_pad_o[31] ;
output \mc_data_pad_o[3] ;
output \mc_data_pad_o[4] ;
output \mc_data_pad_o[5] ;
output \mc_data_pad_o[6] ;
output \mc_data_pad_o[7] ;
output \mc_data_pad_o[8] ;
output \mc_data_pad_o[9] ;
output mc_doe_pad_doe_o;
wire mc_dp_od_0_; 
wire mc_dp_od_1_; 
wire mc_dp_od_2_; 
wire mc_dp_od_3_; 
input \mc_dp_pad_i[0] ;
input \mc_dp_pad_i[1] ;
input \mc_dp_pad_i[2] ;
input \mc_dp_pad_i[3] ;
output \mc_dp_pad_o[0] ;
output \mc_dp_pad_o[1] ;
output \mc_dp_pad_o[2] ;
output \mc_dp_pad_o[3] ;
output \mc_dqm_pad_o[0] ;
output \mc_dqm_pad_o[1] ;
output \mc_dqm_pad_o[2] ;
output \mc_dqm_pad_o[3] ;
output mc_oe_pad_o_;
output mc_ras_pad_o_;
output mc_rp_pad_o_;
wire mc_sts_ir; 
input mc_sts_pad_i;
output mc_vpen_pad_o;
output mc_we_pad_o_;
output mc_zz_pad_o;
wire mem_ack; 
wire mem_ack_r; 
wire mem_dout_0_; 
wire mem_dout_10_; 
wire mem_dout_11_; 
wire mem_dout_12_; 
wire mem_dout_13_; 
wire mem_dout_14_; 
wire mem_dout_15_; 
wire mem_dout_16_; 
wire mem_dout_17_; 
wire mem_dout_18_; 
wire mem_dout_19_; 
wire mem_dout_1_; 
wire mem_dout_20_; 
wire mem_dout_21_; 
wire mem_dout_22_; 
wire mem_dout_23_; 
wire mem_dout_24_; 
wire mem_dout_25_; 
wire mem_dout_26_; 
wire mem_dout_27_; 
wire mem_dout_28_; 
wire mem_dout_29_; 
wire mem_dout_2_; 
wire mem_dout_30_; 
wire mem_dout_31_; 
wire mem_dout_3_; 
wire mem_dout_4_; 
wire mem_dout_5_; 
wire mem_dout_6_; 
wire mem_dout_7_; 
wire mem_dout_8_; 
wire mem_dout_9_; 
wire next_adr; 
wire next_adr_bF_buf0; 
wire next_adr_bF_buf1; 
wire next_adr_bF_buf2; 
wire next_adr_bF_buf3; 
wire next_adr_bF_buf4; 
wire not_mem_cyc; 
wire obct_cs_0_; 
wire obct_cs_1_; 
wire obct_cs_2_; 
wire obct_cs_3_; 
wire obct_cs_4_; 
wire obct_cs_5_; 
wire obct_cs_6_; 
wire obct_cs_7_; 
wire oe_; 
wire pack_le0; 
wire pack_le1; 
wire pack_le2; 
wire page_size_10_; 
wire page_size_8_; 
wire page_size_9_; 
wire par_err; 
output \poc_o[0] ;
output \poc_o[10] ;
output \poc_o[11] ;
output \poc_o[12] ;
output \poc_o[13] ;
output \poc_o[14] ;
output \poc_o[15] ;
output \poc_o[16] ;
output \poc_o[17] ;
output \poc_o[18] ;
output \poc_o[19] ;
output \poc_o[1] ;
output \poc_o[20] ;
output \poc_o[21] ;
output \poc_o[22] ;
output \poc_o[23] ;
output \poc_o[24] ;
output \poc_o[25] ;
output \poc_o[26] ;
output \poc_o[27] ;
output \poc_o[28] ;
output \poc_o[29] ;
output \poc_o[2] ;
output \poc_o[30] ;
output \poc_o[31] ;
output \poc_o[3] ;
output \poc_o[4] ;
output \poc_o[5] ;
output \poc_o[6] ;
output \poc_o[7] ;
output \poc_o[8] ;
output \poc_o[9] ;
wire ras_; 
wire ref_int_0_; 
wire ref_int_1_; 
wire ref_int_2_; 
input resume_req_i;
wire rf_dout_0_; 
wire rf_dout_10_; 
wire rf_dout_11_; 
wire rf_dout_12_; 
wire rf_dout_13_; 
wire rf_dout_14_; 
wire rf_dout_15_; 
wire rf_dout_16_; 
wire rf_dout_17_; 
wire rf_dout_18_; 
wire rf_dout_19_; 
wire rf_dout_1_; 
wire rf_dout_20_; 
wire rf_dout_21_; 
wire rf_dout_22_; 
wire rf_dout_23_; 
wire rf_dout_24_; 
wire rf_dout_25_; 
wire rf_dout_26_; 
wire rf_dout_27_; 
wire rf_dout_28_; 
wire rf_dout_29_; 
wire rf_dout_2_; 
wire rf_dout_30_; 
wire rf_dout_31_; 
wire rf_dout_3_; 
wire rf_dout_4_; 
wire rf_dout_5_; 
wire rf_dout_6_; 
wire rf_dout_7_; 
wire rf_dout_8_; 
wire rf_dout_9_; 
wire rfr_ack; 
wire rfr_ps_val_0_; 
wire rfr_ps_val_1_; 
wire rfr_ps_val_2_; 
wire rfr_ps_val_3_; 
wire rfr_ps_val_4_; 
wire rfr_ps_val_5_; 
wire rfr_ps_val_6_; 
wire rfr_ps_val_7_; 
wire rfr_req; 
wire row_adr_0_; 
wire row_adr_0_bF_buf0_; 
wire row_adr_0_bF_buf1_; 
wire row_adr_0_bF_buf2_; 
wire row_adr_0_bF_buf3_; 
wire row_adr_10_; 
wire row_adr_10_bF_buf0_; 
wire row_adr_10_bF_buf1_; 
wire row_adr_10_bF_buf2_; 
wire row_adr_10_bF_buf3_; 
wire row_adr_11_; 
wire row_adr_11_bF_buf0_; 
wire row_adr_11_bF_buf1_; 
wire row_adr_11_bF_buf2_; 
wire row_adr_11_bF_buf3_; 
wire row_adr_12_; 
wire row_adr_12_bF_buf0_; 
wire row_adr_12_bF_buf1_; 
wire row_adr_12_bF_buf2_; 
wire row_adr_12_bF_buf3_; 
wire row_adr_1_; 
wire row_adr_1_bF_buf0_; 
wire row_adr_1_bF_buf1_; 
wire row_adr_1_bF_buf2_; 
wire row_adr_1_bF_buf3_; 
wire row_adr_2_; 
wire row_adr_2_bF_buf0_; 
wire row_adr_2_bF_buf1_; 
wire row_adr_2_bF_buf2_; 
wire row_adr_2_bF_buf3_; 
wire row_adr_3_; 
wire row_adr_3_bF_buf0_; 
wire row_adr_3_bF_buf1_; 
wire row_adr_3_bF_buf2_; 
wire row_adr_3_bF_buf3_; 
wire row_adr_4_; 
wire row_adr_4_bF_buf0_; 
wire row_adr_4_bF_buf1_; 
wire row_adr_4_bF_buf2_; 
wire row_adr_4_bF_buf3_; 
wire row_adr_5_; 
wire row_adr_5_bF_buf0_; 
wire row_adr_5_bF_buf1_; 
wire row_adr_5_bF_buf2_; 
wire row_adr_5_bF_buf3_; 
wire row_adr_6_; 
wire row_adr_6_bF_buf0_; 
wire row_adr_6_bF_buf1_; 
wire row_adr_6_bF_buf2_; 
wire row_adr_6_bF_buf3_; 
wire row_adr_7_; 
wire row_adr_7_bF_buf0_; 
wire row_adr_7_bF_buf1_; 
wire row_adr_7_bF_buf2_; 
wire row_adr_7_bF_buf3_; 
wire row_adr_8_; 
wire row_adr_8_bF_buf0_; 
wire row_adr_8_bF_buf1_; 
wire row_adr_8_bF_buf2_; 
wire row_adr_8_bF_buf3_; 
wire row_adr_9_; 
wire row_adr_9_bF_buf0_; 
wire row_adr_9_bF_buf1_; 
wire row_adr_9_bF_buf2_; 
wire row_adr_9_bF_buf3_; 
wire row_same; 
wire row_sel; 
input rst_i;
wire sp_csc_10_; 
wire sp_csc_1_; 
wire sp_csc_2_; 
wire sp_csc_3_; 
wire sp_csc_4_; 
wire sp_csc_5_; 
wire sp_csc_6_; 
wire sp_csc_7_; 
wire sp_csc_9_; 
wire sp_tms_0_; 
wire sp_tms_10_; 
wire sp_tms_11_; 
wire sp_tms_12_; 
wire sp_tms_13_; 
wire sp_tms_14_; 
wire sp_tms_15_; 
wire sp_tms_16_; 
wire sp_tms_17_; 
wire sp_tms_18_; 
wire sp_tms_19_; 
wire sp_tms_1_; 
wire sp_tms_20_; 
wire sp_tms_21_; 
wire sp_tms_22_; 
wire sp_tms_23_; 
wire sp_tms_24_; 
wire sp_tms_25_; 
wire sp_tms_26_; 
wire sp_tms_27_; 
wire sp_tms_2_; 
wire sp_tms_3_; 
wire sp_tms_4_; 
wire sp_tms_5_; 
wire sp_tms_6_; 
wire sp_tms_7_; 
wire sp_tms_8_; 
wire sp_tms_9_; 
wire spec_req_cs_0_; 
wire spec_req_cs_0_bF_buf0_; 
wire spec_req_cs_0_bF_buf1_; 
wire spec_req_cs_0_bF_buf2_; 
wire spec_req_cs_0_bF_buf3_; 
wire spec_req_cs_0_bF_buf4_; 
wire spec_req_cs_0_bF_buf5_; 
wire spec_req_cs_1_; 
wire spec_req_cs_1_bF_buf0_; 
wire spec_req_cs_1_bF_buf1_; 
wire spec_req_cs_1_bF_buf2_; 
wire spec_req_cs_1_bF_buf3_; 
wire spec_req_cs_1_bF_buf4_; 
wire spec_req_cs_1_bF_buf5_; 
wire spec_req_cs_2_; 
wire spec_req_cs_2_bF_buf0_; 
wire spec_req_cs_2_bF_buf1_; 
wire spec_req_cs_2_bF_buf2_; 
wire spec_req_cs_2_bF_buf3_; 
wire spec_req_cs_2_bF_buf4_; 
wire spec_req_cs_2_bF_buf5_; 
wire spec_req_cs_3_; 
wire spec_req_cs_3_bF_buf0_; 
wire spec_req_cs_3_bF_buf1_; 
wire spec_req_cs_3_bF_buf2_; 
wire spec_req_cs_3_bF_buf3_; 
wire spec_req_cs_3_bF_buf4_; 
wire spec_req_cs_3_bF_buf5_; 
wire spec_req_cs_4_; 
wire spec_req_cs_4_bF_buf0_; 
wire spec_req_cs_4_bF_buf1_; 
wire spec_req_cs_4_bF_buf2_; 
wire spec_req_cs_4_bF_buf3_; 
wire spec_req_cs_4_bF_buf4_; 
wire spec_req_cs_4_bF_buf5_; 
wire spec_req_cs_5_; 
wire spec_req_cs_5_bF_buf0_; 
wire spec_req_cs_5_bF_buf1_; 
wire spec_req_cs_5_bF_buf2_; 
wire spec_req_cs_5_bF_buf3_; 
wire spec_req_cs_5_bF_buf4_; 
wire spec_req_cs_5_bF_buf5_; 
wire spec_req_cs_6_; 
wire spec_req_cs_6_bF_buf0_; 
wire spec_req_cs_6_bF_buf1_; 
wire spec_req_cs_6_bF_buf2_; 
wire spec_req_cs_6_bF_buf3_; 
wire spec_req_cs_6_bF_buf4_; 
wire spec_req_cs_6_bF_buf5_; 
wire spec_req_cs_7_; 
input susp_req_i;
wire susp_sel; 
output suspended_o;
wire tms_0_; 
wire tms_10_; 
wire tms_11_; 
wire tms_12_; 
wire tms_13_; 
wire tms_14_; 
wire tms_15_; 
wire tms_16_; 
wire tms_17_; 
wire tms_18_; 
wire tms_19_; 
wire tms_1_; 
wire tms_20_; 
wire tms_21_; 
wire tms_22_; 
wire tms_23_; 
wire tms_24_; 
wire tms_25_; 
wire tms_26_; 
wire tms_27_; 
wire tms_2_; 
wire tms_3_; 
wire tms_4_; 
wire tms_5_; 
wire tms_6_; 
wire tms_7_; 
wire tms_8_; 
wire tms_9_; 
wire tms_s_0_; 
wire tms_s_10_; 
wire tms_s_11_; 
wire tms_s_12_; 
wire tms_s_13_; 
wire tms_s_14_; 
wire tms_s_15_; 
wire tms_s_16_; 
wire tms_s_17_; 
wire tms_s_18_; 
wire tms_s_19_; 
wire tms_s_1_; 
wire tms_s_20_; 
wire tms_s_21_; 
wire tms_s_22_; 
wire tms_s_23_; 
wire tms_s_24_; 
wire tms_s_25_; 
wire tms_s_26_; 
wire tms_s_27_; 
wire tms_s_2_; 
wire tms_s_3_; 
wire tms_s_4_; 
wire tms_s_5_; 
wire tms_s_6_; 
wire tms_s_7_; 
wire tms_s_8_; 
wire tms_s_9_; 
wire u0__0cs_7_0__0_; 
wire u0__0cs_7_0__1_; 
wire u0__0cs_7_0__2_; 
wire u0__0cs_7_0__3_; 
wire u0__0cs_7_0__4_; 
wire u0__0cs_7_0__5_; 
wire u0__0cs_7_0__6_; 
wire u0__0cs_7_0__7_; 
wire u0__0csc_31_0__10_; 
wire u0__0csc_31_0__11_; 
wire u0__0csc_31_0__1_; 
wire u0__0csc_31_0__2_; 
wire u0__0csc_31_0__3_; 
wire u0__0csc_31_0__4_; 
wire u0__0csc_31_0__5_; 
wire u0__0csc_31_0__6_; 
wire u0__0csc_31_0__7_; 
wire u0__0csc_31_0__9_; 
wire u0__0csc_mask_r_10_0__0_; 
wire u0__0csc_mask_r_10_0__10_; 
wire u0__0csc_mask_r_10_0__1_; 
wire u0__0csc_mask_r_10_0__2_; 
wire u0__0csc_mask_r_10_0__3_; 
wire u0__0csc_mask_r_10_0__4_; 
wire u0__0csc_mask_r_10_0__5_; 
wire u0__0csc_mask_r_10_0__6_; 
wire u0__0csc_mask_r_10_0__7_; 
wire u0__0csc_mask_r_10_0__8_; 
wire u0__0csc_mask_r_10_0__9_; 
wire u0__0csr_r2_7_0__0_; 
wire u0__0csr_r2_7_0__1_; 
wire u0__0csr_r2_7_0__2_; 
wire u0__0csr_r2_7_0__3_; 
wire u0__0csr_r2_7_0__4_; 
wire u0__0csr_r2_7_0__5_; 
wire u0__0csr_r2_7_0__6_; 
wire u0__0csr_r2_7_0__7_; 
wire u0__0csr_r_10_1__0_; 
wire u0__0csr_r_10_1__1_; 
wire u0__0csr_r_10_1__2_; 
wire u0__0csr_r_10_1__3_; 
wire u0__0csr_r_10_1__4_; 
wire u0__0csr_r_10_1__5_; 
wire u0__0csr_r_10_1__6_; 
wire u0__0csr_r_10_1__7_; 
wire u0__0csr_r_10_1__8_; 
wire u0__0csr_r_10_1__9_; 
wire u0__0init_req_0_0_; 
wire u0__0lmr_req_0_0_; 
wire u0__0poc_31_0__0_; 
wire u0__0poc_31_0__10_; 
wire u0__0poc_31_0__11_; 
wire u0__0poc_31_0__12_; 
wire u0__0poc_31_0__13_; 
wire u0__0poc_31_0__14_; 
wire u0__0poc_31_0__15_; 
wire u0__0poc_31_0__16_; 
wire u0__0poc_31_0__17_; 
wire u0__0poc_31_0__18_; 
wire u0__0poc_31_0__19_; 
wire u0__0poc_31_0__1_; 
wire u0__0poc_31_0__20_; 
wire u0__0poc_31_0__21_; 
wire u0__0poc_31_0__22_; 
wire u0__0poc_31_0__23_; 
wire u0__0poc_31_0__24_; 
wire u0__0poc_31_0__25_; 
wire u0__0poc_31_0__26_; 
wire u0__0poc_31_0__27_; 
wire u0__0poc_31_0__28_; 
wire u0__0poc_31_0__29_; 
wire u0__0poc_31_0__2_; 
wire u0__0poc_31_0__30_; 
wire u0__0poc_31_0__31_; 
wire u0__0poc_31_0__3_; 
wire u0__0poc_31_0__4_; 
wire u0__0poc_31_0__5_; 
wire u0__0poc_31_0__6_; 
wire u0__0poc_31_0__7_; 
wire u0__0poc_31_0__8_; 
wire u0__0poc_31_0__9_; 
wire u0__0rf_we_0_0_; 
wire u0__0sp_csc_31_0__10_; 
wire u0__0sp_csc_31_0__1_; 
wire u0__0sp_csc_31_0__2_; 
wire u0__0sp_csc_31_0__3_; 
wire u0__0sp_csc_31_0__4_; 
wire u0__0sp_csc_31_0__5_; 
wire u0__0sp_csc_31_0__6_; 
wire u0__0sp_csc_31_0__7_; 
wire u0__0sp_csc_31_0__9_; 
wire u0__0sp_tms_31_0__0_; 
wire u0__0sp_tms_31_0__10_; 
wire u0__0sp_tms_31_0__11_; 
wire u0__0sp_tms_31_0__12_; 
wire u0__0sp_tms_31_0__13_; 
wire u0__0sp_tms_31_0__14_; 
wire u0__0sp_tms_31_0__15_; 
wire u0__0sp_tms_31_0__16_; 
wire u0__0sp_tms_31_0__17_; 
wire u0__0sp_tms_31_0__18_; 
wire u0__0sp_tms_31_0__19_; 
wire u0__0sp_tms_31_0__1_; 
wire u0__0sp_tms_31_0__20_; 
wire u0__0sp_tms_31_0__21_; 
wire u0__0sp_tms_31_0__22_; 
wire u0__0sp_tms_31_0__23_; 
wire u0__0sp_tms_31_0__24_; 
wire u0__0sp_tms_31_0__25_; 
wire u0__0sp_tms_31_0__26_; 
wire u0__0sp_tms_31_0__27_; 
wire u0__0sp_tms_31_0__2_; 
wire u0__0sp_tms_31_0__3_; 
wire u0__0sp_tms_31_0__4_; 
wire u0__0sp_tms_31_0__5_; 
wire u0__0sp_tms_31_0__6_; 
wire u0__0sp_tms_31_0__7_; 
wire u0__0sp_tms_31_0__8_; 
wire u0__0sp_tms_31_0__9_; 
wire u0__0spec_req_cs_7_0__0_; 
wire u0__0spec_req_cs_7_0__1_; 
wire u0__0spec_req_cs_7_0__2_; 
wire u0__0spec_req_cs_7_0__3_; 
wire u0__0spec_req_cs_7_0__4_; 
wire u0__0spec_req_cs_7_0__5_; 
wire u0__0spec_req_cs_7_0__6_; 
wire u0__0spec_req_cs_7_0__7_; 
wire u0__0sreq_cs_le_0_0_; 
wire u0__0tms_31_0__0_; 
wire u0__0tms_31_0__10_; 
wire u0__0tms_31_0__11_; 
wire u0__0tms_31_0__12_; 
wire u0__0tms_31_0__13_; 
wire u0__0tms_31_0__14_; 
wire u0__0tms_31_0__15_; 
wire u0__0tms_31_0__16_; 
wire u0__0tms_31_0__17_; 
wire u0__0tms_31_0__18_; 
wire u0__0tms_31_0__19_; 
wire u0__0tms_31_0__1_; 
wire u0__0tms_31_0__20_; 
wire u0__0tms_31_0__21_; 
wire u0__0tms_31_0__22_; 
wire u0__0tms_31_0__23_; 
wire u0__0tms_31_0__24_; 
wire u0__0tms_31_0__25_; 
wire u0__0tms_31_0__26_; 
wire u0__0tms_31_0__27_; 
wire u0__0tms_31_0__2_; 
wire u0__0tms_31_0__3_; 
wire u0__0tms_31_0__4_; 
wire u0__0tms_31_0__5_; 
wire u0__0tms_31_0__6_; 
wire u0__0tms_31_0__7_; 
wire u0__0tms_31_0__8_; 
wire u0__0tms_31_0__9_; 
wire u0__0wp_err_0_0_; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8; 
wire u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9; 
wire u0__abc_76628_new_n1100_; 
wire u0__abc_76628_new_n1101_; 
wire u0__abc_76628_new_n1102_; 
wire u0__abc_76628_new_n1103_; 
wire u0__abc_76628_new_n1104_; 
wire u0__abc_76628_new_n1105_; 
wire u0__abc_76628_new_n1106_; 
wire u0__abc_76628_new_n1107_; 
wire u0__abc_76628_new_n1109_; 
wire u0__abc_76628_new_n1110_; 
wire u0__abc_76628_new_n1111_; 
wire u0__abc_76628_new_n1112_; 
wire u0__abc_76628_new_n1113_; 
wire u0__abc_76628_new_n1114_; 
wire u0__abc_76628_new_n1116_; 
wire u0__abc_76628_new_n1117_; 
wire u0__abc_76628_new_n1118_; 
wire u0__abc_76628_new_n1119_; 
wire u0__abc_76628_new_n1120_; 
wire u0__abc_76628_new_n1121_; 
wire u0__abc_76628_new_n1122_; 
wire u0__abc_76628_new_n1124_; 
wire u0__abc_76628_new_n1125_; 
wire u0__abc_76628_new_n1126_; 
wire u0__abc_76628_new_n1127_; 
wire u0__abc_76628_new_n1128_; 
wire u0__abc_76628_new_n1129_; 
wire u0__abc_76628_new_n1130_; 
wire u0__abc_76628_new_n1132_; 
wire u0__abc_76628_new_n1133_; 
wire u0__abc_76628_new_n1134_; 
wire u0__abc_76628_new_n1135_; 
wire u0__abc_76628_new_n1136_; 
wire u0__abc_76628_new_n1137_; 
wire u0__abc_76628_new_n1138_; 
wire u0__abc_76628_new_n1139_; 
wire u0__abc_76628_new_n1141_; 
wire u0__abc_76628_new_n1142_; 
wire u0__abc_76628_new_n1143_; 
wire u0__abc_76628_new_n1144_; 
wire u0__abc_76628_new_n1145_; 
wire u0__abc_76628_new_n1146_; 
wire u0__abc_76628_new_n1147_; 
wire u0__abc_76628_new_n1149_; 
wire u0__abc_76628_new_n1150_; 
wire u0__abc_76628_new_n1151_; 
wire u0__abc_76628_new_n1152_; 
wire u0__abc_76628_new_n1153_; 
wire u0__abc_76628_new_n1154_; 
wire u0__abc_76628_new_n1155_; 
wire u0__abc_76628_new_n1156_; 
wire u0__abc_76628_new_n1158_; 
wire u0__abc_76628_new_n1159_; 
wire u0__abc_76628_new_n1160_; 
wire u0__abc_76628_new_n1161_; 
wire u0__abc_76628_new_n1162_; 
wire u0__abc_76628_new_n1163_; 
wire u0__abc_76628_new_n1164_; 
wire u0__abc_76628_new_n1165_; 
wire u0__abc_76628_new_n1167_; 
wire u0__abc_76628_new_n1168_; 
wire u0__abc_76628_new_n1169_; 
wire u0__abc_76628_new_n1169__bF_buf0; 
wire u0__abc_76628_new_n1169__bF_buf1; 
wire u0__abc_76628_new_n1169__bF_buf2; 
wire u0__abc_76628_new_n1169__bF_buf3; 
wire u0__abc_76628_new_n1169__bF_buf4; 
wire u0__abc_76628_new_n1169__bF_buf5; 
wire u0__abc_76628_new_n1169__bF_buf6; 
wire u0__abc_76628_new_n1170_; 
wire u0__abc_76628_new_n1170__bF_buf0; 
wire u0__abc_76628_new_n1170__bF_buf1; 
wire u0__abc_76628_new_n1170__bF_buf2; 
wire u0__abc_76628_new_n1170__bF_buf3; 
wire u0__abc_76628_new_n1170__bF_buf4; 
wire u0__abc_76628_new_n1170__bF_buf5; 
wire u0__abc_76628_new_n1170__bF_buf6; 
wire u0__abc_76628_new_n1171_; 
wire u0__abc_76628_new_n1172_; 
wire u0__abc_76628_new_n1172__bF_buf0; 
wire u0__abc_76628_new_n1172__bF_buf1; 
wire u0__abc_76628_new_n1172__bF_buf2; 
wire u0__abc_76628_new_n1172__bF_buf3; 
wire u0__abc_76628_new_n1172__bF_buf4; 
wire u0__abc_76628_new_n1172__bF_buf5; 
wire u0__abc_76628_new_n1173_; 
wire u0__abc_76628_new_n1173__bF_buf0; 
wire u0__abc_76628_new_n1173__bF_buf1; 
wire u0__abc_76628_new_n1173__bF_buf2; 
wire u0__abc_76628_new_n1173__bF_buf3; 
wire u0__abc_76628_new_n1173__bF_buf4; 
wire u0__abc_76628_new_n1173__bF_buf5; 
wire u0__abc_76628_new_n1174_; 
wire u0__abc_76628_new_n1174__bF_buf0; 
wire u0__abc_76628_new_n1174__bF_buf1; 
wire u0__abc_76628_new_n1174__bF_buf2; 
wire u0__abc_76628_new_n1174__bF_buf3; 
wire u0__abc_76628_new_n1174__bF_buf4; 
wire u0__abc_76628_new_n1174__bF_buf5; 
wire u0__abc_76628_new_n1175_; 
wire u0__abc_76628_new_n1175__bF_buf0; 
wire u0__abc_76628_new_n1175__bF_buf1; 
wire u0__abc_76628_new_n1175__bF_buf2; 
wire u0__abc_76628_new_n1175__bF_buf3; 
wire u0__abc_76628_new_n1175__bF_buf4; 
wire u0__abc_76628_new_n1175__bF_buf5; 
wire u0__abc_76628_new_n1176_; 
wire u0__abc_76628_new_n1177_; 
wire u0__abc_76628_new_n1177__bF_buf0; 
wire u0__abc_76628_new_n1177__bF_buf1; 
wire u0__abc_76628_new_n1177__bF_buf2; 
wire u0__abc_76628_new_n1177__bF_buf3; 
wire u0__abc_76628_new_n1177__bF_buf4; 
wire u0__abc_76628_new_n1177__bF_buf5; 
wire u0__abc_76628_new_n1178_; 
wire u0__abc_76628_new_n1179_; 
wire u0__abc_76628_new_n1179__bF_buf0; 
wire u0__abc_76628_new_n1179__bF_buf1; 
wire u0__abc_76628_new_n1179__bF_buf2; 
wire u0__abc_76628_new_n1179__bF_buf3; 
wire u0__abc_76628_new_n1179__bF_buf4; 
wire u0__abc_76628_new_n1179__bF_buf5; 
wire u0__abc_76628_new_n1180_; 
wire u0__abc_76628_new_n1181_; 
wire u0__abc_76628_new_n1182_; 
wire u0__abc_76628_new_n1183_; 
wire u0__abc_76628_new_n1184_; 
wire u0__abc_76628_new_n1185_; 
wire u0__abc_76628_new_n1186_; 
wire u0__abc_76628_new_n1187_; 
wire u0__abc_76628_new_n1188_; 
wire u0__abc_76628_new_n1189_; 
wire u0__abc_76628_new_n1190_; 
wire u0__abc_76628_new_n1191_; 
wire u0__abc_76628_new_n1192_; 
wire u0__abc_76628_new_n1193_; 
wire u0__abc_76628_new_n1194_; 
wire u0__abc_76628_new_n1195_; 
wire u0__abc_76628_new_n1196_; 
wire u0__abc_76628_new_n1197_; 
wire u0__abc_76628_new_n1197__bF_buf0; 
wire u0__abc_76628_new_n1197__bF_buf1; 
wire u0__abc_76628_new_n1197__bF_buf2; 
wire u0__abc_76628_new_n1197__bF_buf3; 
wire u0__abc_76628_new_n1197__bF_buf4; 
wire u0__abc_76628_new_n1197__bF_buf5; 
wire u0__abc_76628_new_n1198_; 
wire u0__abc_76628_new_n1199_; 
wire u0__abc_76628_new_n1200_; 
wire u0__abc_76628_new_n1202_; 
wire u0__abc_76628_new_n1203_; 
wire u0__abc_76628_new_n1204_; 
wire u0__abc_76628_new_n1205_; 
wire u0__abc_76628_new_n1206_; 
wire u0__abc_76628_new_n1207_; 
wire u0__abc_76628_new_n1208_; 
wire u0__abc_76628_new_n1209_; 
wire u0__abc_76628_new_n1210_; 
wire u0__abc_76628_new_n1211_; 
wire u0__abc_76628_new_n1212_; 
wire u0__abc_76628_new_n1213_; 
wire u0__abc_76628_new_n1214_; 
wire u0__abc_76628_new_n1215_; 
wire u0__abc_76628_new_n1216_; 
wire u0__abc_76628_new_n1217_; 
wire u0__abc_76628_new_n1218_; 
wire u0__abc_76628_new_n1219_; 
wire u0__abc_76628_new_n1220_; 
wire u0__abc_76628_new_n1221_; 
wire u0__abc_76628_new_n1222_; 
wire u0__abc_76628_new_n1223_; 
wire u0__abc_76628_new_n1224_; 
wire u0__abc_76628_new_n1226_; 
wire u0__abc_76628_new_n1227_; 
wire u0__abc_76628_new_n1228_; 
wire u0__abc_76628_new_n1229_; 
wire u0__abc_76628_new_n1230_; 
wire u0__abc_76628_new_n1231_; 
wire u0__abc_76628_new_n1232_; 
wire u0__abc_76628_new_n1233_; 
wire u0__abc_76628_new_n1234_; 
wire u0__abc_76628_new_n1235_; 
wire u0__abc_76628_new_n1236_; 
wire u0__abc_76628_new_n1237_; 
wire u0__abc_76628_new_n1238_; 
wire u0__abc_76628_new_n1239_; 
wire u0__abc_76628_new_n1240_; 
wire u0__abc_76628_new_n1241_; 
wire u0__abc_76628_new_n1242_; 
wire u0__abc_76628_new_n1243_; 
wire u0__abc_76628_new_n1244_; 
wire u0__abc_76628_new_n1245_; 
wire u0__abc_76628_new_n1246_; 
wire u0__abc_76628_new_n1247_; 
wire u0__abc_76628_new_n1248_; 
wire u0__abc_76628_new_n1250_; 
wire u0__abc_76628_new_n1251_; 
wire u0__abc_76628_new_n1252_; 
wire u0__abc_76628_new_n1253_; 
wire u0__abc_76628_new_n1254_; 
wire u0__abc_76628_new_n1255_; 
wire u0__abc_76628_new_n1256_; 
wire u0__abc_76628_new_n1257_; 
wire u0__abc_76628_new_n1258_; 
wire u0__abc_76628_new_n1259_; 
wire u0__abc_76628_new_n1260_; 
wire u0__abc_76628_new_n1261_; 
wire u0__abc_76628_new_n1262_; 
wire u0__abc_76628_new_n1263_; 
wire u0__abc_76628_new_n1264_; 
wire u0__abc_76628_new_n1265_; 
wire u0__abc_76628_new_n1266_; 
wire u0__abc_76628_new_n1267_; 
wire u0__abc_76628_new_n1268_; 
wire u0__abc_76628_new_n1269_; 
wire u0__abc_76628_new_n1270_; 
wire u0__abc_76628_new_n1271_; 
wire u0__abc_76628_new_n1272_; 
wire u0__abc_76628_new_n1274_; 
wire u0__abc_76628_new_n1275_; 
wire u0__abc_76628_new_n1276_; 
wire u0__abc_76628_new_n1277_; 
wire u0__abc_76628_new_n1278_; 
wire u0__abc_76628_new_n1279_; 
wire u0__abc_76628_new_n1280_; 
wire u0__abc_76628_new_n1281_; 
wire u0__abc_76628_new_n1282_; 
wire u0__abc_76628_new_n1283_; 
wire u0__abc_76628_new_n1284_; 
wire u0__abc_76628_new_n1285_; 
wire u0__abc_76628_new_n1286_; 
wire u0__abc_76628_new_n1287_; 
wire u0__abc_76628_new_n1288_; 
wire u0__abc_76628_new_n1289_; 
wire u0__abc_76628_new_n1290_; 
wire u0__abc_76628_new_n1291_; 
wire u0__abc_76628_new_n1292_; 
wire u0__abc_76628_new_n1293_; 
wire u0__abc_76628_new_n1294_; 
wire u0__abc_76628_new_n1295_; 
wire u0__abc_76628_new_n1296_; 
wire u0__abc_76628_new_n1298_; 
wire u0__abc_76628_new_n1299_; 
wire u0__abc_76628_new_n1300_; 
wire u0__abc_76628_new_n1301_; 
wire u0__abc_76628_new_n1302_; 
wire u0__abc_76628_new_n1303_; 
wire u0__abc_76628_new_n1304_; 
wire u0__abc_76628_new_n1305_; 
wire u0__abc_76628_new_n1306_; 
wire u0__abc_76628_new_n1307_; 
wire u0__abc_76628_new_n1308_; 
wire u0__abc_76628_new_n1309_; 
wire u0__abc_76628_new_n1310_; 
wire u0__abc_76628_new_n1311_; 
wire u0__abc_76628_new_n1312_; 
wire u0__abc_76628_new_n1313_; 
wire u0__abc_76628_new_n1314_; 
wire u0__abc_76628_new_n1315_; 
wire u0__abc_76628_new_n1316_; 
wire u0__abc_76628_new_n1317_; 
wire u0__abc_76628_new_n1318_; 
wire u0__abc_76628_new_n1319_; 
wire u0__abc_76628_new_n1320_; 
wire u0__abc_76628_new_n1322_; 
wire u0__abc_76628_new_n1323_; 
wire u0__abc_76628_new_n1324_; 
wire u0__abc_76628_new_n1325_; 
wire u0__abc_76628_new_n1326_; 
wire u0__abc_76628_new_n1327_; 
wire u0__abc_76628_new_n1328_; 
wire u0__abc_76628_new_n1329_; 
wire u0__abc_76628_new_n1330_; 
wire u0__abc_76628_new_n1331_; 
wire u0__abc_76628_new_n1332_; 
wire u0__abc_76628_new_n1333_; 
wire u0__abc_76628_new_n1334_; 
wire u0__abc_76628_new_n1335_; 
wire u0__abc_76628_new_n1336_; 
wire u0__abc_76628_new_n1337_; 
wire u0__abc_76628_new_n1338_; 
wire u0__abc_76628_new_n1339_; 
wire u0__abc_76628_new_n1340_; 
wire u0__abc_76628_new_n1341_; 
wire u0__abc_76628_new_n1342_; 
wire u0__abc_76628_new_n1343_; 
wire u0__abc_76628_new_n1344_; 
wire u0__abc_76628_new_n1346_; 
wire u0__abc_76628_new_n1347_; 
wire u0__abc_76628_new_n1348_; 
wire u0__abc_76628_new_n1349_; 
wire u0__abc_76628_new_n1350_; 
wire u0__abc_76628_new_n1351_; 
wire u0__abc_76628_new_n1352_; 
wire u0__abc_76628_new_n1353_; 
wire u0__abc_76628_new_n1354_; 
wire u0__abc_76628_new_n1355_; 
wire u0__abc_76628_new_n1356_; 
wire u0__abc_76628_new_n1357_; 
wire u0__abc_76628_new_n1358_; 
wire u0__abc_76628_new_n1359_; 
wire u0__abc_76628_new_n1360_; 
wire u0__abc_76628_new_n1361_; 
wire u0__abc_76628_new_n1362_; 
wire u0__abc_76628_new_n1363_; 
wire u0__abc_76628_new_n1364_; 
wire u0__abc_76628_new_n1365_; 
wire u0__abc_76628_new_n1366_; 
wire u0__abc_76628_new_n1367_; 
wire u0__abc_76628_new_n1368_; 
wire u0__abc_76628_new_n1370_; 
wire u0__abc_76628_new_n1371_; 
wire u0__abc_76628_new_n1372_; 
wire u0__abc_76628_new_n1373_; 
wire u0__abc_76628_new_n1374_; 
wire u0__abc_76628_new_n1375_; 
wire u0__abc_76628_new_n1376_; 
wire u0__abc_76628_new_n1377_; 
wire u0__abc_76628_new_n1378_; 
wire u0__abc_76628_new_n1379_; 
wire u0__abc_76628_new_n1380_; 
wire u0__abc_76628_new_n1381_; 
wire u0__abc_76628_new_n1382_; 
wire u0__abc_76628_new_n1383_; 
wire u0__abc_76628_new_n1384_; 
wire u0__abc_76628_new_n1385_; 
wire u0__abc_76628_new_n1386_; 
wire u0__abc_76628_new_n1387_; 
wire u0__abc_76628_new_n1388_; 
wire u0__abc_76628_new_n1389_; 
wire u0__abc_76628_new_n1390_; 
wire u0__abc_76628_new_n1391_; 
wire u0__abc_76628_new_n1392_; 
wire u0__abc_76628_new_n1394_; 
wire u0__abc_76628_new_n1395_; 
wire u0__abc_76628_new_n1396_; 
wire u0__abc_76628_new_n1397_; 
wire u0__abc_76628_new_n1398_; 
wire u0__abc_76628_new_n1399_; 
wire u0__abc_76628_new_n1400_; 
wire u0__abc_76628_new_n1401_; 
wire u0__abc_76628_new_n1402_; 
wire u0__abc_76628_new_n1403_; 
wire u0__abc_76628_new_n1404_; 
wire u0__abc_76628_new_n1405_; 
wire u0__abc_76628_new_n1406_; 
wire u0__abc_76628_new_n1407_; 
wire u0__abc_76628_new_n1408_; 
wire u0__abc_76628_new_n1409_; 
wire u0__abc_76628_new_n1410_; 
wire u0__abc_76628_new_n1411_; 
wire u0__abc_76628_new_n1412_; 
wire u0__abc_76628_new_n1413_; 
wire u0__abc_76628_new_n1414_; 
wire u0__abc_76628_new_n1415_; 
wire u0__abc_76628_new_n1416_; 
wire u0__abc_76628_new_n1418_; 
wire u0__abc_76628_new_n1419_; 
wire u0__abc_76628_new_n1420_; 
wire u0__abc_76628_new_n1421_; 
wire u0__abc_76628_new_n1422_; 
wire u0__abc_76628_new_n1423_; 
wire u0__abc_76628_new_n1424_; 
wire u0__abc_76628_new_n1425_; 
wire u0__abc_76628_new_n1426_; 
wire u0__abc_76628_new_n1427_; 
wire u0__abc_76628_new_n1428_; 
wire u0__abc_76628_new_n1429_; 
wire u0__abc_76628_new_n1430_; 
wire u0__abc_76628_new_n1431_; 
wire u0__abc_76628_new_n1432_; 
wire u0__abc_76628_new_n1433_; 
wire u0__abc_76628_new_n1434_; 
wire u0__abc_76628_new_n1435_; 
wire u0__abc_76628_new_n1436_; 
wire u0__abc_76628_new_n1437_; 
wire u0__abc_76628_new_n1438_; 
wire u0__abc_76628_new_n1439_; 
wire u0__abc_76628_new_n1440_; 
wire u0__abc_76628_new_n1442_; 
wire u0__abc_76628_new_n1443_; 
wire u0__abc_76628_new_n1444_; 
wire u0__abc_76628_new_n1445_; 
wire u0__abc_76628_new_n1446_; 
wire u0__abc_76628_new_n1447_; 
wire u0__abc_76628_new_n1448_; 
wire u0__abc_76628_new_n1449_; 
wire u0__abc_76628_new_n1450_; 
wire u0__abc_76628_new_n1451_; 
wire u0__abc_76628_new_n1452_; 
wire u0__abc_76628_new_n1453_; 
wire u0__abc_76628_new_n1454_; 
wire u0__abc_76628_new_n1455_; 
wire u0__abc_76628_new_n1456_; 
wire u0__abc_76628_new_n1457_; 
wire u0__abc_76628_new_n1458_; 
wire u0__abc_76628_new_n1459_; 
wire u0__abc_76628_new_n1460_; 
wire u0__abc_76628_new_n1461_; 
wire u0__abc_76628_new_n1462_; 
wire u0__abc_76628_new_n1463_; 
wire u0__abc_76628_new_n1464_; 
wire u0__abc_76628_new_n1466_; 
wire u0__abc_76628_new_n1467_; 
wire u0__abc_76628_new_n1468_; 
wire u0__abc_76628_new_n1469_; 
wire u0__abc_76628_new_n1470_; 
wire u0__abc_76628_new_n1471_; 
wire u0__abc_76628_new_n1472_; 
wire u0__abc_76628_new_n1473_; 
wire u0__abc_76628_new_n1474_; 
wire u0__abc_76628_new_n1475_; 
wire u0__abc_76628_new_n1476_; 
wire u0__abc_76628_new_n1477_; 
wire u0__abc_76628_new_n1478_; 
wire u0__abc_76628_new_n1479_; 
wire u0__abc_76628_new_n1480_; 
wire u0__abc_76628_new_n1481_; 
wire u0__abc_76628_new_n1482_; 
wire u0__abc_76628_new_n1483_; 
wire u0__abc_76628_new_n1484_; 
wire u0__abc_76628_new_n1485_; 
wire u0__abc_76628_new_n1486_; 
wire u0__abc_76628_new_n1487_; 
wire u0__abc_76628_new_n1488_; 
wire u0__abc_76628_new_n1490_; 
wire u0__abc_76628_new_n1491_; 
wire u0__abc_76628_new_n1492_; 
wire u0__abc_76628_new_n1493_; 
wire u0__abc_76628_new_n1494_; 
wire u0__abc_76628_new_n1495_; 
wire u0__abc_76628_new_n1496_; 
wire u0__abc_76628_new_n1497_; 
wire u0__abc_76628_new_n1498_; 
wire u0__abc_76628_new_n1499_; 
wire u0__abc_76628_new_n1500_; 
wire u0__abc_76628_new_n1501_; 
wire u0__abc_76628_new_n1502_; 
wire u0__abc_76628_new_n1503_; 
wire u0__abc_76628_new_n1504_; 
wire u0__abc_76628_new_n1505_; 
wire u0__abc_76628_new_n1506_; 
wire u0__abc_76628_new_n1507_; 
wire u0__abc_76628_new_n1508_; 
wire u0__abc_76628_new_n1509_; 
wire u0__abc_76628_new_n1510_; 
wire u0__abc_76628_new_n1511_; 
wire u0__abc_76628_new_n1512_; 
wire u0__abc_76628_new_n1514_; 
wire u0__abc_76628_new_n1515_; 
wire u0__abc_76628_new_n1516_; 
wire u0__abc_76628_new_n1517_; 
wire u0__abc_76628_new_n1518_; 
wire u0__abc_76628_new_n1519_; 
wire u0__abc_76628_new_n1520_; 
wire u0__abc_76628_new_n1521_; 
wire u0__abc_76628_new_n1522_; 
wire u0__abc_76628_new_n1523_; 
wire u0__abc_76628_new_n1524_; 
wire u0__abc_76628_new_n1525_; 
wire u0__abc_76628_new_n1526_; 
wire u0__abc_76628_new_n1527_; 
wire u0__abc_76628_new_n1528_; 
wire u0__abc_76628_new_n1529_; 
wire u0__abc_76628_new_n1530_; 
wire u0__abc_76628_new_n1531_; 
wire u0__abc_76628_new_n1532_; 
wire u0__abc_76628_new_n1533_; 
wire u0__abc_76628_new_n1534_; 
wire u0__abc_76628_new_n1535_; 
wire u0__abc_76628_new_n1536_; 
wire u0__abc_76628_new_n1538_; 
wire u0__abc_76628_new_n1539_; 
wire u0__abc_76628_new_n1540_; 
wire u0__abc_76628_new_n1541_; 
wire u0__abc_76628_new_n1542_; 
wire u0__abc_76628_new_n1543_; 
wire u0__abc_76628_new_n1544_; 
wire u0__abc_76628_new_n1545_; 
wire u0__abc_76628_new_n1546_; 
wire u0__abc_76628_new_n1547_; 
wire u0__abc_76628_new_n1548_; 
wire u0__abc_76628_new_n1549_; 
wire u0__abc_76628_new_n1550_; 
wire u0__abc_76628_new_n1551_; 
wire u0__abc_76628_new_n1552_; 
wire u0__abc_76628_new_n1553_; 
wire u0__abc_76628_new_n1554_; 
wire u0__abc_76628_new_n1555_; 
wire u0__abc_76628_new_n1556_; 
wire u0__abc_76628_new_n1557_; 
wire u0__abc_76628_new_n1558_; 
wire u0__abc_76628_new_n1559_; 
wire u0__abc_76628_new_n1560_; 
wire u0__abc_76628_new_n1562_; 
wire u0__abc_76628_new_n1563_; 
wire u0__abc_76628_new_n1564_; 
wire u0__abc_76628_new_n1565_; 
wire u0__abc_76628_new_n1566_; 
wire u0__abc_76628_new_n1567_; 
wire u0__abc_76628_new_n1568_; 
wire u0__abc_76628_new_n1569_; 
wire u0__abc_76628_new_n1570_; 
wire u0__abc_76628_new_n1571_; 
wire u0__abc_76628_new_n1572_; 
wire u0__abc_76628_new_n1573_; 
wire u0__abc_76628_new_n1574_; 
wire u0__abc_76628_new_n1575_; 
wire u0__abc_76628_new_n1576_; 
wire u0__abc_76628_new_n1577_; 
wire u0__abc_76628_new_n1578_; 
wire u0__abc_76628_new_n1579_; 
wire u0__abc_76628_new_n1580_; 
wire u0__abc_76628_new_n1581_; 
wire u0__abc_76628_new_n1582_; 
wire u0__abc_76628_new_n1583_; 
wire u0__abc_76628_new_n1584_; 
wire u0__abc_76628_new_n1586_; 
wire u0__abc_76628_new_n1587_; 
wire u0__abc_76628_new_n1588_; 
wire u0__abc_76628_new_n1589_; 
wire u0__abc_76628_new_n1590_; 
wire u0__abc_76628_new_n1591_; 
wire u0__abc_76628_new_n1592_; 
wire u0__abc_76628_new_n1593_; 
wire u0__abc_76628_new_n1594_; 
wire u0__abc_76628_new_n1595_; 
wire u0__abc_76628_new_n1596_; 
wire u0__abc_76628_new_n1597_; 
wire u0__abc_76628_new_n1598_; 
wire u0__abc_76628_new_n1599_; 
wire u0__abc_76628_new_n1600_; 
wire u0__abc_76628_new_n1601_; 
wire u0__abc_76628_new_n1602_; 
wire u0__abc_76628_new_n1603_; 
wire u0__abc_76628_new_n1604_; 
wire u0__abc_76628_new_n1605_; 
wire u0__abc_76628_new_n1606_; 
wire u0__abc_76628_new_n1607_; 
wire u0__abc_76628_new_n1608_; 
wire u0__abc_76628_new_n1610_; 
wire u0__abc_76628_new_n1611_; 
wire u0__abc_76628_new_n1612_; 
wire u0__abc_76628_new_n1613_; 
wire u0__abc_76628_new_n1614_; 
wire u0__abc_76628_new_n1615_; 
wire u0__abc_76628_new_n1616_; 
wire u0__abc_76628_new_n1617_; 
wire u0__abc_76628_new_n1618_; 
wire u0__abc_76628_new_n1619_; 
wire u0__abc_76628_new_n1620_; 
wire u0__abc_76628_new_n1621_; 
wire u0__abc_76628_new_n1622_; 
wire u0__abc_76628_new_n1623_; 
wire u0__abc_76628_new_n1624_; 
wire u0__abc_76628_new_n1625_; 
wire u0__abc_76628_new_n1626_; 
wire u0__abc_76628_new_n1627_; 
wire u0__abc_76628_new_n1628_; 
wire u0__abc_76628_new_n1629_; 
wire u0__abc_76628_new_n1630_; 
wire u0__abc_76628_new_n1631_; 
wire u0__abc_76628_new_n1632_; 
wire u0__abc_76628_new_n1634_; 
wire u0__abc_76628_new_n1635_; 
wire u0__abc_76628_new_n1636_; 
wire u0__abc_76628_new_n1637_; 
wire u0__abc_76628_new_n1638_; 
wire u0__abc_76628_new_n1639_; 
wire u0__abc_76628_new_n1640_; 
wire u0__abc_76628_new_n1641_; 
wire u0__abc_76628_new_n1642_; 
wire u0__abc_76628_new_n1643_; 
wire u0__abc_76628_new_n1644_; 
wire u0__abc_76628_new_n1645_; 
wire u0__abc_76628_new_n1646_; 
wire u0__abc_76628_new_n1647_; 
wire u0__abc_76628_new_n1648_; 
wire u0__abc_76628_new_n1649_; 
wire u0__abc_76628_new_n1650_; 
wire u0__abc_76628_new_n1651_; 
wire u0__abc_76628_new_n1652_; 
wire u0__abc_76628_new_n1653_; 
wire u0__abc_76628_new_n1654_; 
wire u0__abc_76628_new_n1655_; 
wire u0__abc_76628_new_n1656_; 
wire u0__abc_76628_new_n1658_; 
wire u0__abc_76628_new_n1659_; 
wire u0__abc_76628_new_n1660_; 
wire u0__abc_76628_new_n1661_; 
wire u0__abc_76628_new_n1662_; 
wire u0__abc_76628_new_n1663_; 
wire u0__abc_76628_new_n1664_; 
wire u0__abc_76628_new_n1665_; 
wire u0__abc_76628_new_n1666_; 
wire u0__abc_76628_new_n1667_; 
wire u0__abc_76628_new_n1668_; 
wire u0__abc_76628_new_n1669_; 
wire u0__abc_76628_new_n1670_; 
wire u0__abc_76628_new_n1671_; 
wire u0__abc_76628_new_n1672_; 
wire u0__abc_76628_new_n1673_; 
wire u0__abc_76628_new_n1674_; 
wire u0__abc_76628_new_n1675_; 
wire u0__abc_76628_new_n1676_; 
wire u0__abc_76628_new_n1677_; 
wire u0__abc_76628_new_n1678_; 
wire u0__abc_76628_new_n1679_; 
wire u0__abc_76628_new_n1680_; 
wire u0__abc_76628_new_n1682_; 
wire u0__abc_76628_new_n1683_; 
wire u0__abc_76628_new_n1684_; 
wire u0__abc_76628_new_n1685_; 
wire u0__abc_76628_new_n1686_; 
wire u0__abc_76628_new_n1687_; 
wire u0__abc_76628_new_n1688_; 
wire u0__abc_76628_new_n1689_; 
wire u0__abc_76628_new_n1690_; 
wire u0__abc_76628_new_n1691_; 
wire u0__abc_76628_new_n1692_; 
wire u0__abc_76628_new_n1693_; 
wire u0__abc_76628_new_n1694_; 
wire u0__abc_76628_new_n1695_; 
wire u0__abc_76628_new_n1696_; 
wire u0__abc_76628_new_n1697_; 
wire u0__abc_76628_new_n1698_; 
wire u0__abc_76628_new_n1699_; 
wire u0__abc_76628_new_n1700_; 
wire u0__abc_76628_new_n1701_; 
wire u0__abc_76628_new_n1702_; 
wire u0__abc_76628_new_n1703_; 
wire u0__abc_76628_new_n1704_; 
wire u0__abc_76628_new_n1706_; 
wire u0__abc_76628_new_n1707_; 
wire u0__abc_76628_new_n1708_; 
wire u0__abc_76628_new_n1709_; 
wire u0__abc_76628_new_n1710_; 
wire u0__abc_76628_new_n1711_; 
wire u0__abc_76628_new_n1712_; 
wire u0__abc_76628_new_n1713_; 
wire u0__abc_76628_new_n1714_; 
wire u0__abc_76628_new_n1715_; 
wire u0__abc_76628_new_n1716_; 
wire u0__abc_76628_new_n1717_; 
wire u0__abc_76628_new_n1718_; 
wire u0__abc_76628_new_n1719_; 
wire u0__abc_76628_new_n1720_; 
wire u0__abc_76628_new_n1721_; 
wire u0__abc_76628_new_n1722_; 
wire u0__abc_76628_new_n1723_; 
wire u0__abc_76628_new_n1724_; 
wire u0__abc_76628_new_n1725_; 
wire u0__abc_76628_new_n1726_; 
wire u0__abc_76628_new_n1727_; 
wire u0__abc_76628_new_n1728_; 
wire u0__abc_76628_new_n1730_; 
wire u0__abc_76628_new_n1731_; 
wire u0__abc_76628_new_n1732_; 
wire u0__abc_76628_new_n1733_; 
wire u0__abc_76628_new_n1734_; 
wire u0__abc_76628_new_n1735_; 
wire u0__abc_76628_new_n1736_; 
wire u0__abc_76628_new_n1737_; 
wire u0__abc_76628_new_n1738_; 
wire u0__abc_76628_new_n1739_; 
wire u0__abc_76628_new_n1740_; 
wire u0__abc_76628_new_n1741_; 
wire u0__abc_76628_new_n1742_; 
wire u0__abc_76628_new_n1743_; 
wire u0__abc_76628_new_n1744_; 
wire u0__abc_76628_new_n1745_; 
wire u0__abc_76628_new_n1746_; 
wire u0__abc_76628_new_n1747_; 
wire u0__abc_76628_new_n1748_; 
wire u0__abc_76628_new_n1749_; 
wire u0__abc_76628_new_n1750_; 
wire u0__abc_76628_new_n1751_; 
wire u0__abc_76628_new_n1752_; 
wire u0__abc_76628_new_n1754_; 
wire u0__abc_76628_new_n1755_; 
wire u0__abc_76628_new_n1756_; 
wire u0__abc_76628_new_n1757_; 
wire u0__abc_76628_new_n1758_; 
wire u0__abc_76628_new_n1759_; 
wire u0__abc_76628_new_n1760_; 
wire u0__abc_76628_new_n1761_; 
wire u0__abc_76628_new_n1762_; 
wire u0__abc_76628_new_n1763_; 
wire u0__abc_76628_new_n1764_; 
wire u0__abc_76628_new_n1765_; 
wire u0__abc_76628_new_n1766_; 
wire u0__abc_76628_new_n1767_; 
wire u0__abc_76628_new_n1768_; 
wire u0__abc_76628_new_n1769_; 
wire u0__abc_76628_new_n1770_; 
wire u0__abc_76628_new_n1771_; 
wire u0__abc_76628_new_n1772_; 
wire u0__abc_76628_new_n1773_; 
wire u0__abc_76628_new_n1774_; 
wire u0__abc_76628_new_n1775_; 
wire u0__abc_76628_new_n1776_; 
wire u0__abc_76628_new_n1778_; 
wire u0__abc_76628_new_n1779_; 
wire u0__abc_76628_new_n1780_; 
wire u0__abc_76628_new_n1781_; 
wire u0__abc_76628_new_n1782_; 
wire u0__abc_76628_new_n1783_; 
wire u0__abc_76628_new_n1784_; 
wire u0__abc_76628_new_n1785_; 
wire u0__abc_76628_new_n1786_; 
wire u0__abc_76628_new_n1787_; 
wire u0__abc_76628_new_n1788_; 
wire u0__abc_76628_new_n1789_; 
wire u0__abc_76628_new_n1790_; 
wire u0__abc_76628_new_n1791_; 
wire u0__abc_76628_new_n1792_; 
wire u0__abc_76628_new_n1793_; 
wire u0__abc_76628_new_n1794_; 
wire u0__abc_76628_new_n1795_; 
wire u0__abc_76628_new_n1796_; 
wire u0__abc_76628_new_n1797_; 
wire u0__abc_76628_new_n1798_; 
wire u0__abc_76628_new_n1799_; 
wire u0__abc_76628_new_n1800_; 
wire u0__abc_76628_new_n1802_; 
wire u0__abc_76628_new_n1803_; 
wire u0__abc_76628_new_n1804_; 
wire u0__abc_76628_new_n1805_; 
wire u0__abc_76628_new_n1806_; 
wire u0__abc_76628_new_n1807_; 
wire u0__abc_76628_new_n1808_; 
wire u0__abc_76628_new_n1809_; 
wire u0__abc_76628_new_n1810_; 
wire u0__abc_76628_new_n1811_; 
wire u0__abc_76628_new_n1812_; 
wire u0__abc_76628_new_n1813_; 
wire u0__abc_76628_new_n1814_; 
wire u0__abc_76628_new_n1815_; 
wire u0__abc_76628_new_n1816_; 
wire u0__abc_76628_new_n1817_; 
wire u0__abc_76628_new_n1818_; 
wire u0__abc_76628_new_n1819_; 
wire u0__abc_76628_new_n1820_; 
wire u0__abc_76628_new_n1821_; 
wire u0__abc_76628_new_n1822_; 
wire u0__abc_76628_new_n1823_; 
wire u0__abc_76628_new_n1824_; 
wire u0__abc_76628_new_n1826_; 
wire u0__abc_76628_new_n1827_; 
wire u0__abc_76628_new_n1828_; 
wire u0__abc_76628_new_n1829_; 
wire u0__abc_76628_new_n1830_; 
wire u0__abc_76628_new_n1831_; 
wire u0__abc_76628_new_n1832_; 
wire u0__abc_76628_new_n1833_; 
wire u0__abc_76628_new_n1834_; 
wire u0__abc_76628_new_n1835_; 
wire u0__abc_76628_new_n1836_; 
wire u0__abc_76628_new_n1837_; 
wire u0__abc_76628_new_n1838_; 
wire u0__abc_76628_new_n1839_; 
wire u0__abc_76628_new_n1840_; 
wire u0__abc_76628_new_n1841_; 
wire u0__abc_76628_new_n1842_; 
wire u0__abc_76628_new_n1843_; 
wire u0__abc_76628_new_n1844_; 
wire u0__abc_76628_new_n1845_; 
wire u0__abc_76628_new_n1846_; 
wire u0__abc_76628_new_n1847_; 
wire u0__abc_76628_new_n1848_; 
wire u0__abc_76628_new_n1946_; 
wire u0__abc_76628_new_n1946__bF_buf0; 
wire u0__abc_76628_new_n1946__bF_buf1; 
wire u0__abc_76628_new_n1946__bF_buf2; 
wire u0__abc_76628_new_n1946__bF_buf3; 
wire u0__abc_76628_new_n1947_; 
wire u0__abc_76628_new_n1947__bF_buf0; 
wire u0__abc_76628_new_n1947__bF_buf1; 
wire u0__abc_76628_new_n1947__bF_buf2; 
wire u0__abc_76628_new_n1947__bF_buf3; 
wire u0__abc_76628_new_n1972_; 
wire u0__abc_76628_new_n1973_; 
wire u0__abc_76628_new_n1974_; 
wire u0__abc_76628_new_n1975_; 
wire u0__abc_76628_new_n1976_; 
wire u0__abc_76628_new_n1977_; 
wire u0__abc_76628_new_n1978_; 
wire u0__abc_76628_new_n1979_; 
wire u0__abc_76628_new_n1980_; 
wire u0__abc_76628_new_n1981_; 
wire u0__abc_76628_new_n1982_; 
wire u0__abc_76628_new_n1983_; 
wire u0__abc_76628_new_n1984_; 
wire u0__abc_76628_new_n1985_; 
wire u0__abc_76628_new_n1986_; 
wire u0__abc_76628_new_n1987_; 
wire u0__abc_76628_new_n1988_; 
wire u0__abc_76628_new_n1989_; 
wire u0__abc_76628_new_n1990_; 
wire u0__abc_76628_new_n1991_; 
wire u0__abc_76628_new_n1992_; 
wire u0__abc_76628_new_n1993_; 
wire u0__abc_76628_new_n1994_; 
wire u0__abc_76628_new_n1996_; 
wire u0__abc_76628_new_n1997_; 
wire u0__abc_76628_new_n1998_; 
wire u0__abc_76628_new_n1999_; 
wire u0__abc_76628_new_n2000_; 
wire u0__abc_76628_new_n2001_; 
wire u0__abc_76628_new_n2002_; 
wire u0__abc_76628_new_n2003_; 
wire u0__abc_76628_new_n2004_; 
wire u0__abc_76628_new_n2005_; 
wire u0__abc_76628_new_n2006_; 
wire u0__abc_76628_new_n2007_; 
wire u0__abc_76628_new_n2008_; 
wire u0__abc_76628_new_n2009_; 
wire u0__abc_76628_new_n2010_; 
wire u0__abc_76628_new_n2011_; 
wire u0__abc_76628_new_n2012_; 
wire u0__abc_76628_new_n2013_; 
wire u0__abc_76628_new_n2014_; 
wire u0__abc_76628_new_n2015_; 
wire u0__abc_76628_new_n2016_; 
wire u0__abc_76628_new_n2017_; 
wire u0__abc_76628_new_n2018_; 
wire u0__abc_76628_new_n2020_; 
wire u0__abc_76628_new_n2021_; 
wire u0__abc_76628_new_n2022_; 
wire u0__abc_76628_new_n2023_; 
wire u0__abc_76628_new_n2024_; 
wire u0__abc_76628_new_n2025_; 
wire u0__abc_76628_new_n2026_; 
wire u0__abc_76628_new_n2027_; 
wire u0__abc_76628_new_n2028_; 
wire u0__abc_76628_new_n2029_; 
wire u0__abc_76628_new_n2030_; 
wire u0__abc_76628_new_n2031_; 
wire u0__abc_76628_new_n2032_; 
wire u0__abc_76628_new_n2033_; 
wire u0__abc_76628_new_n2034_; 
wire u0__abc_76628_new_n2035_; 
wire u0__abc_76628_new_n2036_; 
wire u0__abc_76628_new_n2037_; 
wire u0__abc_76628_new_n2038_; 
wire u0__abc_76628_new_n2039_; 
wire u0__abc_76628_new_n2040_; 
wire u0__abc_76628_new_n2041_; 
wire u0__abc_76628_new_n2042_; 
wire u0__abc_76628_new_n2044_; 
wire u0__abc_76628_new_n2045_; 
wire u0__abc_76628_new_n2046_; 
wire u0__abc_76628_new_n2047_; 
wire u0__abc_76628_new_n2048_; 
wire u0__abc_76628_new_n2049_; 
wire u0__abc_76628_new_n2050_; 
wire u0__abc_76628_new_n2051_; 
wire u0__abc_76628_new_n2052_; 
wire u0__abc_76628_new_n2053_; 
wire u0__abc_76628_new_n2054_; 
wire u0__abc_76628_new_n2055_; 
wire u0__abc_76628_new_n2056_; 
wire u0__abc_76628_new_n2057_; 
wire u0__abc_76628_new_n2058_; 
wire u0__abc_76628_new_n2059_; 
wire u0__abc_76628_new_n2060_; 
wire u0__abc_76628_new_n2061_; 
wire u0__abc_76628_new_n2062_; 
wire u0__abc_76628_new_n2063_; 
wire u0__abc_76628_new_n2064_; 
wire u0__abc_76628_new_n2065_; 
wire u0__abc_76628_new_n2066_; 
wire u0__abc_76628_new_n2068_; 
wire u0__abc_76628_new_n2069_; 
wire u0__abc_76628_new_n2070_; 
wire u0__abc_76628_new_n2071_; 
wire u0__abc_76628_new_n2072_; 
wire u0__abc_76628_new_n2073_; 
wire u0__abc_76628_new_n2074_; 
wire u0__abc_76628_new_n2075_; 
wire u0__abc_76628_new_n2076_; 
wire u0__abc_76628_new_n2077_; 
wire u0__abc_76628_new_n2078_; 
wire u0__abc_76628_new_n2079_; 
wire u0__abc_76628_new_n2080_; 
wire u0__abc_76628_new_n2081_; 
wire u0__abc_76628_new_n2082_; 
wire u0__abc_76628_new_n2083_; 
wire u0__abc_76628_new_n2084_; 
wire u0__abc_76628_new_n2085_; 
wire u0__abc_76628_new_n2086_; 
wire u0__abc_76628_new_n2087_; 
wire u0__abc_76628_new_n2088_; 
wire u0__abc_76628_new_n2089_; 
wire u0__abc_76628_new_n2090_; 
wire u0__abc_76628_new_n2092_; 
wire u0__abc_76628_new_n2093_; 
wire u0__abc_76628_new_n2094_; 
wire u0__abc_76628_new_n2095_; 
wire u0__abc_76628_new_n2096_; 
wire u0__abc_76628_new_n2097_; 
wire u0__abc_76628_new_n2098_; 
wire u0__abc_76628_new_n2099_; 
wire u0__abc_76628_new_n2100_; 
wire u0__abc_76628_new_n2101_; 
wire u0__abc_76628_new_n2102_; 
wire u0__abc_76628_new_n2103_; 
wire u0__abc_76628_new_n2104_; 
wire u0__abc_76628_new_n2105_; 
wire u0__abc_76628_new_n2106_; 
wire u0__abc_76628_new_n2107_; 
wire u0__abc_76628_new_n2108_; 
wire u0__abc_76628_new_n2109_; 
wire u0__abc_76628_new_n2110_; 
wire u0__abc_76628_new_n2111_; 
wire u0__abc_76628_new_n2112_; 
wire u0__abc_76628_new_n2113_; 
wire u0__abc_76628_new_n2114_; 
wire u0__abc_76628_new_n2116_; 
wire u0__abc_76628_new_n2117_; 
wire u0__abc_76628_new_n2118_; 
wire u0__abc_76628_new_n2119_; 
wire u0__abc_76628_new_n2120_; 
wire u0__abc_76628_new_n2121_; 
wire u0__abc_76628_new_n2122_; 
wire u0__abc_76628_new_n2123_; 
wire u0__abc_76628_new_n2124_; 
wire u0__abc_76628_new_n2125_; 
wire u0__abc_76628_new_n2126_; 
wire u0__abc_76628_new_n2127_; 
wire u0__abc_76628_new_n2128_; 
wire u0__abc_76628_new_n2129_; 
wire u0__abc_76628_new_n2130_; 
wire u0__abc_76628_new_n2131_; 
wire u0__abc_76628_new_n2132_; 
wire u0__abc_76628_new_n2133_; 
wire u0__abc_76628_new_n2134_; 
wire u0__abc_76628_new_n2135_; 
wire u0__abc_76628_new_n2136_; 
wire u0__abc_76628_new_n2137_; 
wire u0__abc_76628_new_n2138_; 
wire u0__abc_76628_new_n2164_; 
wire u0__abc_76628_new_n2165_; 
wire u0__abc_76628_new_n2166_; 
wire u0__abc_76628_new_n2167_; 
wire u0__abc_76628_new_n2168_; 
wire u0__abc_76628_new_n2169_; 
wire u0__abc_76628_new_n2170_; 
wire u0__abc_76628_new_n2171_; 
wire u0__abc_76628_new_n2172_; 
wire u0__abc_76628_new_n2173_; 
wire u0__abc_76628_new_n2174_; 
wire u0__abc_76628_new_n2175_; 
wire u0__abc_76628_new_n2176_; 
wire u0__abc_76628_new_n2177_; 
wire u0__abc_76628_new_n2178_; 
wire u0__abc_76628_new_n2179_; 
wire u0__abc_76628_new_n2180_; 
wire u0__abc_76628_new_n2181_; 
wire u0__abc_76628_new_n2182_; 
wire u0__abc_76628_new_n2183_; 
wire u0__abc_76628_new_n2184_; 
wire u0__abc_76628_new_n2185_; 
wire u0__abc_76628_new_n2186_; 
wire u0__abc_76628_new_n2188_; 
wire u0__abc_76628_new_n2189_; 
wire u0__abc_76628_new_n2190_; 
wire u0__abc_76628_new_n2191_; 
wire u0__abc_76628_new_n2192_; 
wire u0__abc_76628_new_n2193_; 
wire u0__abc_76628_new_n2194_; 
wire u0__abc_76628_new_n2195_; 
wire u0__abc_76628_new_n2196_; 
wire u0__abc_76628_new_n2197_; 
wire u0__abc_76628_new_n2198_; 
wire u0__abc_76628_new_n2199_; 
wire u0__abc_76628_new_n2200_; 
wire u0__abc_76628_new_n2201_; 
wire u0__abc_76628_new_n2202_; 
wire u0__abc_76628_new_n2203_; 
wire u0__abc_76628_new_n2204_; 
wire u0__abc_76628_new_n2205_; 
wire u0__abc_76628_new_n2206_; 
wire u0__abc_76628_new_n2207_; 
wire u0__abc_76628_new_n2208_; 
wire u0__abc_76628_new_n2209_; 
wire u0__abc_76628_new_n2210_; 
wire u0__abc_76628_new_n2716_; 
wire u0__abc_76628_new_n2717_; 
wire u0__abc_76628_new_n2717__bF_buf0; 
wire u0__abc_76628_new_n2717__bF_buf1; 
wire u0__abc_76628_new_n2717__bF_buf2; 
wire u0__abc_76628_new_n2717__bF_buf3; 
wire u0__abc_76628_new_n2717__bF_buf4; 
wire u0__abc_76628_new_n2717__bF_buf5; 
wire u0__abc_76628_new_n2718_; 
wire u0__abc_76628_new_n2718__bF_buf0; 
wire u0__abc_76628_new_n2718__bF_buf1; 
wire u0__abc_76628_new_n2718__bF_buf2; 
wire u0__abc_76628_new_n2718__bF_buf3; 
wire u0__abc_76628_new_n2718__bF_buf4; 
wire u0__abc_76628_new_n2718__bF_buf5; 
wire u0__abc_76628_new_n2719_; 
wire u0__abc_76628_new_n2719__bF_buf0; 
wire u0__abc_76628_new_n2719__bF_buf1; 
wire u0__abc_76628_new_n2719__bF_buf2; 
wire u0__abc_76628_new_n2719__bF_buf3; 
wire u0__abc_76628_new_n2719__bF_buf4; 
wire u0__abc_76628_new_n2719__bF_buf5; 
wire u0__abc_76628_new_n2720_; 
wire u0__abc_76628_new_n2720__bF_buf0; 
wire u0__abc_76628_new_n2720__bF_buf1; 
wire u0__abc_76628_new_n2720__bF_buf2; 
wire u0__abc_76628_new_n2720__bF_buf3; 
wire u0__abc_76628_new_n2720__bF_buf4; 
wire u0__abc_76628_new_n2720__bF_buf5; 
wire u0__abc_76628_new_n2721_; 
wire u0__abc_76628_new_n2722_; 
wire u0__abc_76628_new_n2722__bF_buf0; 
wire u0__abc_76628_new_n2722__bF_buf1; 
wire u0__abc_76628_new_n2722__bF_buf2; 
wire u0__abc_76628_new_n2722__bF_buf3; 
wire u0__abc_76628_new_n2722__bF_buf4; 
wire u0__abc_76628_new_n2722__bF_buf5; 
wire u0__abc_76628_new_n2723_; 
wire u0__abc_76628_new_n2724_; 
wire u0__abc_76628_new_n2724__bF_buf0; 
wire u0__abc_76628_new_n2724__bF_buf1; 
wire u0__abc_76628_new_n2724__bF_buf2; 
wire u0__abc_76628_new_n2724__bF_buf3; 
wire u0__abc_76628_new_n2724__bF_buf4; 
wire u0__abc_76628_new_n2724__bF_buf5; 
wire u0__abc_76628_new_n2725_; 
wire u0__abc_76628_new_n2726_; 
wire u0__abc_76628_new_n2727_; 
wire u0__abc_76628_new_n2728_; 
wire u0__abc_76628_new_n2729_; 
wire u0__abc_76628_new_n2730_; 
wire u0__abc_76628_new_n2731_; 
wire u0__abc_76628_new_n2732_; 
wire u0__abc_76628_new_n2733_; 
wire u0__abc_76628_new_n2734_; 
wire u0__abc_76628_new_n2735_; 
wire u0__abc_76628_new_n2736_; 
wire u0__abc_76628_new_n2737_; 
wire u0__abc_76628_new_n2738_; 
wire u0__abc_76628_new_n2739_; 
wire u0__abc_76628_new_n2740_; 
wire u0__abc_76628_new_n2741_; 
wire u0__abc_76628_new_n2742_; 
wire u0__abc_76628_new_n2742__bF_buf0; 
wire u0__abc_76628_new_n2742__bF_buf1; 
wire u0__abc_76628_new_n2742__bF_buf2; 
wire u0__abc_76628_new_n2742__bF_buf3; 
wire u0__abc_76628_new_n2742__bF_buf4; 
wire u0__abc_76628_new_n2742__bF_buf5; 
wire u0__abc_76628_new_n2743_; 
wire u0__abc_76628_new_n2744_; 
wire u0__abc_76628_new_n2745_; 
wire u0__abc_76628_new_n2747_; 
wire u0__abc_76628_new_n2748_; 
wire u0__abc_76628_new_n2749_; 
wire u0__abc_76628_new_n2750_; 
wire u0__abc_76628_new_n2751_; 
wire u0__abc_76628_new_n2752_; 
wire u0__abc_76628_new_n2753_; 
wire u0__abc_76628_new_n2754_; 
wire u0__abc_76628_new_n2755_; 
wire u0__abc_76628_new_n2756_; 
wire u0__abc_76628_new_n2757_; 
wire u0__abc_76628_new_n2758_; 
wire u0__abc_76628_new_n2759_; 
wire u0__abc_76628_new_n2760_; 
wire u0__abc_76628_new_n2761_; 
wire u0__abc_76628_new_n2762_; 
wire u0__abc_76628_new_n2763_; 
wire u0__abc_76628_new_n2764_; 
wire u0__abc_76628_new_n2765_; 
wire u0__abc_76628_new_n2766_; 
wire u0__abc_76628_new_n2767_; 
wire u0__abc_76628_new_n2768_; 
wire u0__abc_76628_new_n2769_; 
wire u0__abc_76628_new_n2771_; 
wire u0__abc_76628_new_n2772_; 
wire u0__abc_76628_new_n2773_; 
wire u0__abc_76628_new_n2774_; 
wire u0__abc_76628_new_n2775_; 
wire u0__abc_76628_new_n2776_; 
wire u0__abc_76628_new_n2777_; 
wire u0__abc_76628_new_n2778_; 
wire u0__abc_76628_new_n2779_; 
wire u0__abc_76628_new_n2780_; 
wire u0__abc_76628_new_n2781_; 
wire u0__abc_76628_new_n2782_; 
wire u0__abc_76628_new_n2783_; 
wire u0__abc_76628_new_n2784_; 
wire u0__abc_76628_new_n2785_; 
wire u0__abc_76628_new_n2786_; 
wire u0__abc_76628_new_n2787_; 
wire u0__abc_76628_new_n2788_; 
wire u0__abc_76628_new_n2789_; 
wire u0__abc_76628_new_n2790_; 
wire u0__abc_76628_new_n2791_; 
wire u0__abc_76628_new_n2792_; 
wire u0__abc_76628_new_n2793_; 
wire u0__abc_76628_new_n2795_; 
wire u0__abc_76628_new_n2796_; 
wire u0__abc_76628_new_n2797_; 
wire u0__abc_76628_new_n2798_; 
wire u0__abc_76628_new_n2799_; 
wire u0__abc_76628_new_n2800_; 
wire u0__abc_76628_new_n2801_; 
wire u0__abc_76628_new_n2802_; 
wire u0__abc_76628_new_n2803_; 
wire u0__abc_76628_new_n2804_; 
wire u0__abc_76628_new_n2805_; 
wire u0__abc_76628_new_n2806_; 
wire u0__abc_76628_new_n2807_; 
wire u0__abc_76628_new_n2808_; 
wire u0__abc_76628_new_n2809_; 
wire u0__abc_76628_new_n2810_; 
wire u0__abc_76628_new_n2811_; 
wire u0__abc_76628_new_n2812_; 
wire u0__abc_76628_new_n2813_; 
wire u0__abc_76628_new_n2814_; 
wire u0__abc_76628_new_n2815_; 
wire u0__abc_76628_new_n2816_; 
wire u0__abc_76628_new_n2817_; 
wire u0__abc_76628_new_n2819_; 
wire u0__abc_76628_new_n2820_; 
wire u0__abc_76628_new_n2821_; 
wire u0__abc_76628_new_n2822_; 
wire u0__abc_76628_new_n2823_; 
wire u0__abc_76628_new_n2824_; 
wire u0__abc_76628_new_n2825_; 
wire u0__abc_76628_new_n2826_; 
wire u0__abc_76628_new_n2827_; 
wire u0__abc_76628_new_n2828_; 
wire u0__abc_76628_new_n2829_; 
wire u0__abc_76628_new_n2830_; 
wire u0__abc_76628_new_n2831_; 
wire u0__abc_76628_new_n2832_; 
wire u0__abc_76628_new_n2833_; 
wire u0__abc_76628_new_n2834_; 
wire u0__abc_76628_new_n2835_; 
wire u0__abc_76628_new_n2836_; 
wire u0__abc_76628_new_n2837_; 
wire u0__abc_76628_new_n2838_; 
wire u0__abc_76628_new_n2839_; 
wire u0__abc_76628_new_n2840_; 
wire u0__abc_76628_new_n2841_; 
wire u0__abc_76628_new_n2843_; 
wire u0__abc_76628_new_n2844_; 
wire u0__abc_76628_new_n2845_; 
wire u0__abc_76628_new_n2846_; 
wire u0__abc_76628_new_n2847_; 
wire u0__abc_76628_new_n2848_; 
wire u0__abc_76628_new_n2849_; 
wire u0__abc_76628_new_n2850_; 
wire u0__abc_76628_new_n2851_; 
wire u0__abc_76628_new_n2852_; 
wire u0__abc_76628_new_n2853_; 
wire u0__abc_76628_new_n2854_; 
wire u0__abc_76628_new_n2855_; 
wire u0__abc_76628_new_n2856_; 
wire u0__abc_76628_new_n2857_; 
wire u0__abc_76628_new_n2858_; 
wire u0__abc_76628_new_n2859_; 
wire u0__abc_76628_new_n2860_; 
wire u0__abc_76628_new_n2861_; 
wire u0__abc_76628_new_n2862_; 
wire u0__abc_76628_new_n2863_; 
wire u0__abc_76628_new_n2864_; 
wire u0__abc_76628_new_n2865_; 
wire u0__abc_76628_new_n2867_; 
wire u0__abc_76628_new_n2868_; 
wire u0__abc_76628_new_n2869_; 
wire u0__abc_76628_new_n2870_; 
wire u0__abc_76628_new_n2871_; 
wire u0__abc_76628_new_n2872_; 
wire u0__abc_76628_new_n2873_; 
wire u0__abc_76628_new_n2874_; 
wire u0__abc_76628_new_n2875_; 
wire u0__abc_76628_new_n2876_; 
wire u0__abc_76628_new_n2877_; 
wire u0__abc_76628_new_n2878_; 
wire u0__abc_76628_new_n2879_; 
wire u0__abc_76628_new_n2880_; 
wire u0__abc_76628_new_n2881_; 
wire u0__abc_76628_new_n2882_; 
wire u0__abc_76628_new_n2883_; 
wire u0__abc_76628_new_n2884_; 
wire u0__abc_76628_new_n2885_; 
wire u0__abc_76628_new_n2886_; 
wire u0__abc_76628_new_n2887_; 
wire u0__abc_76628_new_n2888_; 
wire u0__abc_76628_new_n2889_; 
wire u0__abc_76628_new_n2891_; 
wire u0__abc_76628_new_n2892_; 
wire u0__abc_76628_new_n2893_; 
wire u0__abc_76628_new_n2894_; 
wire u0__abc_76628_new_n2895_; 
wire u0__abc_76628_new_n2896_; 
wire u0__abc_76628_new_n2897_; 
wire u0__abc_76628_new_n2898_; 
wire u0__abc_76628_new_n2899_; 
wire u0__abc_76628_new_n2900_; 
wire u0__abc_76628_new_n2901_; 
wire u0__abc_76628_new_n2902_; 
wire u0__abc_76628_new_n2903_; 
wire u0__abc_76628_new_n2904_; 
wire u0__abc_76628_new_n2905_; 
wire u0__abc_76628_new_n2906_; 
wire u0__abc_76628_new_n2907_; 
wire u0__abc_76628_new_n2908_; 
wire u0__abc_76628_new_n2909_; 
wire u0__abc_76628_new_n2910_; 
wire u0__abc_76628_new_n2911_; 
wire u0__abc_76628_new_n2912_; 
wire u0__abc_76628_new_n2913_; 
wire u0__abc_76628_new_n2915_; 
wire u0__abc_76628_new_n2916_; 
wire u0__abc_76628_new_n2917_; 
wire u0__abc_76628_new_n2918_; 
wire u0__abc_76628_new_n2919_; 
wire u0__abc_76628_new_n2920_; 
wire u0__abc_76628_new_n2921_; 
wire u0__abc_76628_new_n2922_; 
wire u0__abc_76628_new_n2923_; 
wire u0__abc_76628_new_n2924_; 
wire u0__abc_76628_new_n2925_; 
wire u0__abc_76628_new_n2926_; 
wire u0__abc_76628_new_n2927_; 
wire u0__abc_76628_new_n2928_; 
wire u0__abc_76628_new_n2929_; 
wire u0__abc_76628_new_n2930_; 
wire u0__abc_76628_new_n2931_; 
wire u0__abc_76628_new_n2932_; 
wire u0__abc_76628_new_n2933_; 
wire u0__abc_76628_new_n2934_; 
wire u0__abc_76628_new_n2935_; 
wire u0__abc_76628_new_n2936_; 
wire u0__abc_76628_new_n2937_; 
wire u0__abc_76628_new_n2939_; 
wire u0__abc_76628_new_n2940_; 
wire u0__abc_76628_new_n2941_; 
wire u0__abc_76628_new_n2942_; 
wire u0__abc_76628_new_n2943_; 
wire u0__abc_76628_new_n2944_; 
wire u0__abc_76628_new_n2945_; 
wire u0__abc_76628_new_n2946_; 
wire u0__abc_76628_new_n2947_; 
wire u0__abc_76628_new_n2948_; 
wire u0__abc_76628_new_n2949_; 
wire u0__abc_76628_new_n2950_; 
wire u0__abc_76628_new_n2951_; 
wire u0__abc_76628_new_n2952_; 
wire u0__abc_76628_new_n2953_; 
wire u0__abc_76628_new_n2954_; 
wire u0__abc_76628_new_n2955_; 
wire u0__abc_76628_new_n2956_; 
wire u0__abc_76628_new_n2957_; 
wire u0__abc_76628_new_n2958_; 
wire u0__abc_76628_new_n2959_; 
wire u0__abc_76628_new_n2960_; 
wire u0__abc_76628_new_n2961_; 
wire u0__abc_76628_new_n2963_; 
wire u0__abc_76628_new_n2964_; 
wire u0__abc_76628_new_n2965_; 
wire u0__abc_76628_new_n2966_; 
wire u0__abc_76628_new_n2967_; 
wire u0__abc_76628_new_n2968_; 
wire u0__abc_76628_new_n2969_; 
wire u0__abc_76628_new_n2970_; 
wire u0__abc_76628_new_n2971_; 
wire u0__abc_76628_new_n2972_; 
wire u0__abc_76628_new_n2973_; 
wire u0__abc_76628_new_n2974_; 
wire u0__abc_76628_new_n2975_; 
wire u0__abc_76628_new_n2976_; 
wire u0__abc_76628_new_n2977_; 
wire u0__abc_76628_new_n2978_; 
wire u0__abc_76628_new_n2979_; 
wire u0__abc_76628_new_n2980_; 
wire u0__abc_76628_new_n2981_; 
wire u0__abc_76628_new_n2982_; 
wire u0__abc_76628_new_n2983_; 
wire u0__abc_76628_new_n2984_; 
wire u0__abc_76628_new_n2985_; 
wire u0__abc_76628_new_n2987_; 
wire u0__abc_76628_new_n2988_; 
wire u0__abc_76628_new_n2989_; 
wire u0__abc_76628_new_n2990_; 
wire u0__abc_76628_new_n2991_; 
wire u0__abc_76628_new_n2992_; 
wire u0__abc_76628_new_n2993_; 
wire u0__abc_76628_new_n2994_; 
wire u0__abc_76628_new_n2995_; 
wire u0__abc_76628_new_n2996_; 
wire u0__abc_76628_new_n2997_; 
wire u0__abc_76628_new_n2998_; 
wire u0__abc_76628_new_n2999_; 
wire u0__abc_76628_new_n3000_; 
wire u0__abc_76628_new_n3001_; 
wire u0__abc_76628_new_n3002_; 
wire u0__abc_76628_new_n3003_; 
wire u0__abc_76628_new_n3004_; 
wire u0__abc_76628_new_n3005_; 
wire u0__abc_76628_new_n3006_; 
wire u0__abc_76628_new_n3007_; 
wire u0__abc_76628_new_n3008_; 
wire u0__abc_76628_new_n3009_; 
wire u0__abc_76628_new_n3011_; 
wire u0__abc_76628_new_n3012_; 
wire u0__abc_76628_new_n3013_; 
wire u0__abc_76628_new_n3014_; 
wire u0__abc_76628_new_n3015_; 
wire u0__abc_76628_new_n3016_; 
wire u0__abc_76628_new_n3017_; 
wire u0__abc_76628_new_n3018_; 
wire u0__abc_76628_new_n3019_; 
wire u0__abc_76628_new_n3020_; 
wire u0__abc_76628_new_n3021_; 
wire u0__abc_76628_new_n3022_; 
wire u0__abc_76628_new_n3023_; 
wire u0__abc_76628_new_n3024_; 
wire u0__abc_76628_new_n3025_; 
wire u0__abc_76628_new_n3026_; 
wire u0__abc_76628_new_n3027_; 
wire u0__abc_76628_new_n3028_; 
wire u0__abc_76628_new_n3029_; 
wire u0__abc_76628_new_n3030_; 
wire u0__abc_76628_new_n3031_; 
wire u0__abc_76628_new_n3032_; 
wire u0__abc_76628_new_n3033_; 
wire u0__abc_76628_new_n3035_; 
wire u0__abc_76628_new_n3036_; 
wire u0__abc_76628_new_n3037_; 
wire u0__abc_76628_new_n3038_; 
wire u0__abc_76628_new_n3039_; 
wire u0__abc_76628_new_n3040_; 
wire u0__abc_76628_new_n3041_; 
wire u0__abc_76628_new_n3042_; 
wire u0__abc_76628_new_n3043_; 
wire u0__abc_76628_new_n3044_; 
wire u0__abc_76628_new_n3045_; 
wire u0__abc_76628_new_n3046_; 
wire u0__abc_76628_new_n3047_; 
wire u0__abc_76628_new_n3048_; 
wire u0__abc_76628_new_n3049_; 
wire u0__abc_76628_new_n3050_; 
wire u0__abc_76628_new_n3051_; 
wire u0__abc_76628_new_n3052_; 
wire u0__abc_76628_new_n3053_; 
wire u0__abc_76628_new_n3054_; 
wire u0__abc_76628_new_n3055_; 
wire u0__abc_76628_new_n3056_; 
wire u0__abc_76628_new_n3057_; 
wire u0__abc_76628_new_n3059_; 
wire u0__abc_76628_new_n3060_; 
wire u0__abc_76628_new_n3061_; 
wire u0__abc_76628_new_n3062_; 
wire u0__abc_76628_new_n3063_; 
wire u0__abc_76628_new_n3064_; 
wire u0__abc_76628_new_n3065_; 
wire u0__abc_76628_new_n3066_; 
wire u0__abc_76628_new_n3067_; 
wire u0__abc_76628_new_n3068_; 
wire u0__abc_76628_new_n3069_; 
wire u0__abc_76628_new_n3070_; 
wire u0__abc_76628_new_n3071_; 
wire u0__abc_76628_new_n3072_; 
wire u0__abc_76628_new_n3073_; 
wire u0__abc_76628_new_n3074_; 
wire u0__abc_76628_new_n3075_; 
wire u0__abc_76628_new_n3076_; 
wire u0__abc_76628_new_n3077_; 
wire u0__abc_76628_new_n3078_; 
wire u0__abc_76628_new_n3079_; 
wire u0__abc_76628_new_n3080_; 
wire u0__abc_76628_new_n3081_; 
wire u0__abc_76628_new_n3083_; 
wire u0__abc_76628_new_n3084_; 
wire u0__abc_76628_new_n3085_; 
wire u0__abc_76628_new_n3086_; 
wire u0__abc_76628_new_n3087_; 
wire u0__abc_76628_new_n3088_; 
wire u0__abc_76628_new_n3089_; 
wire u0__abc_76628_new_n3090_; 
wire u0__abc_76628_new_n3091_; 
wire u0__abc_76628_new_n3092_; 
wire u0__abc_76628_new_n3093_; 
wire u0__abc_76628_new_n3094_; 
wire u0__abc_76628_new_n3095_; 
wire u0__abc_76628_new_n3096_; 
wire u0__abc_76628_new_n3097_; 
wire u0__abc_76628_new_n3098_; 
wire u0__abc_76628_new_n3099_; 
wire u0__abc_76628_new_n3100_; 
wire u0__abc_76628_new_n3101_; 
wire u0__abc_76628_new_n3102_; 
wire u0__abc_76628_new_n3103_; 
wire u0__abc_76628_new_n3104_; 
wire u0__abc_76628_new_n3105_; 
wire u0__abc_76628_new_n3107_; 
wire u0__abc_76628_new_n3108_; 
wire u0__abc_76628_new_n3109_; 
wire u0__abc_76628_new_n3110_; 
wire u0__abc_76628_new_n3111_; 
wire u0__abc_76628_new_n3112_; 
wire u0__abc_76628_new_n3113_; 
wire u0__abc_76628_new_n3114_; 
wire u0__abc_76628_new_n3115_; 
wire u0__abc_76628_new_n3116_; 
wire u0__abc_76628_new_n3117_; 
wire u0__abc_76628_new_n3118_; 
wire u0__abc_76628_new_n3119_; 
wire u0__abc_76628_new_n3120_; 
wire u0__abc_76628_new_n3121_; 
wire u0__abc_76628_new_n3122_; 
wire u0__abc_76628_new_n3123_; 
wire u0__abc_76628_new_n3124_; 
wire u0__abc_76628_new_n3125_; 
wire u0__abc_76628_new_n3126_; 
wire u0__abc_76628_new_n3127_; 
wire u0__abc_76628_new_n3128_; 
wire u0__abc_76628_new_n3129_; 
wire u0__abc_76628_new_n3131_; 
wire u0__abc_76628_new_n3132_; 
wire u0__abc_76628_new_n3133_; 
wire u0__abc_76628_new_n3134_; 
wire u0__abc_76628_new_n3135_; 
wire u0__abc_76628_new_n3136_; 
wire u0__abc_76628_new_n3137_; 
wire u0__abc_76628_new_n3138_; 
wire u0__abc_76628_new_n3139_; 
wire u0__abc_76628_new_n3140_; 
wire u0__abc_76628_new_n3141_; 
wire u0__abc_76628_new_n3142_; 
wire u0__abc_76628_new_n3143_; 
wire u0__abc_76628_new_n3144_; 
wire u0__abc_76628_new_n3145_; 
wire u0__abc_76628_new_n3146_; 
wire u0__abc_76628_new_n3147_; 
wire u0__abc_76628_new_n3148_; 
wire u0__abc_76628_new_n3149_; 
wire u0__abc_76628_new_n3150_; 
wire u0__abc_76628_new_n3151_; 
wire u0__abc_76628_new_n3152_; 
wire u0__abc_76628_new_n3153_; 
wire u0__abc_76628_new_n3155_; 
wire u0__abc_76628_new_n3156_; 
wire u0__abc_76628_new_n3157_; 
wire u0__abc_76628_new_n3158_; 
wire u0__abc_76628_new_n3159_; 
wire u0__abc_76628_new_n3160_; 
wire u0__abc_76628_new_n3161_; 
wire u0__abc_76628_new_n3162_; 
wire u0__abc_76628_new_n3163_; 
wire u0__abc_76628_new_n3164_; 
wire u0__abc_76628_new_n3165_; 
wire u0__abc_76628_new_n3166_; 
wire u0__abc_76628_new_n3167_; 
wire u0__abc_76628_new_n3168_; 
wire u0__abc_76628_new_n3169_; 
wire u0__abc_76628_new_n3170_; 
wire u0__abc_76628_new_n3171_; 
wire u0__abc_76628_new_n3172_; 
wire u0__abc_76628_new_n3173_; 
wire u0__abc_76628_new_n3174_; 
wire u0__abc_76628_new_n3175_; 
wire u0__abc_76628_new_n3176_; 
wire u0__abc_76628_new_n3177_; 
wire u0__abc_76628_new_n3179_; 
wire u0__abc_76628_new_n3180_; 
wire u0__abc_76628_new_n3181_; 
wire u0__abc_76628_new_n3182_; 
wire u0__abc_76628_new_n3183_; 
wire u0__abc_76628_new_n3184_; 
wire u0__abc_76628_new_n3185_; 
wire u0__abc_76628_new_n3186_; 
wire u0__abc_76628_new_n3187_; 
wire u0__abc_76628_new_n3188_; 
wire u0__abc_76628_new_n3189_; 
wire u0__abc_76628_new_n3190_; 
wire u0__abc_76628_new_n3191_; 
wire u0__abc_76628_new_n3192_; 
wire u0__abc_76628_new_n3193_; 
wire u0__abc_76628_new_n3194_; 
wire u0__abc_76628_new_n3195_; 
wire u0__abc_76628_new_n3196_; 
wire u0__abc_76628_new_n3197_; 
wire u0__abc_76628_new_n3198_; 
wire u0__abc_76628_new_n3199_; 
wire u0__abc_76628_new_n3200_; 
wire u0__abc_76628_new_n3201_; 
wire u0__abc_76628_new_n3203_; 
wire u0__abc_76628_new_n3204_; 
wire u0__abc_76628_new_n3205_; 
wire u0__abc_76628_new_n3206_; 
wire u0__abc_76628_new_n3207_; 
wire u0__abc_76628_new_n3208_; 
wire u0__abc_76628_new_n3209_; 
wire u0__abc_76628_new_n3210_; 
wire u0__abc_76628_new_n3211_; 
wire u0__abc_76628_new_n3212_; 
wire u0__abc_76628_new_n3213_; 
wire u0__abc_76628_new_n3214_; 
wire u0__abc_76628_new_n3215_; 
wire u0__abc_76628_new_n3216_; 
wire u0__abc_76628_new_n3217_; 
wire u0__abc_76628_new_n3218_; 
wire u0__abc_76628_new_n3219_; 
wire u0__abc_76628_new_n3220_; 
wire u0__abc_76628_new_n3221_; 
wire u0__abc_76628_new_n3222_; 
wire u0__abc_76628_new_n3223_; 
wire u0__abc_76628_new_n3224_; 
wire u0__abc_76628_new_n3225_; 
wire u0__abc_76628_new_n3227_; 
wire u0__abc_76628_new_n3228_; 
wire u0__abc_76628_new_n3229_; 
wire u0__abc_76628_new_n3230_; 
wire u0__abc_76628_new_n3231_; 
wire u0__abc_76628_new_n3232_; 
wire u0__abc_76628_new_n3233_; 
wire u0__abc_76628_new_n3234_; 
wire u0__abc_76628_new_n3235_; 
wire u0__abc_76628_new_n3236_; 
wire u0__abc_76628_new_n3237_; 
wire u0__abc_76628_new_n3238_; 
wire u0__abc_76628_new_n3239_; 
wire u0__abc_76628_new_n3240_; 
wire u0__abc_76628_new_n3241_; 
wire u0__abc_76628_new_n3242_; 
wire u0__abc_76628_new_n3243_; 
wire u0__abc_76628_new_n3244_; 
wire u0__abc_76628_new_n3245_; 
wire u0__abc_76628_new_n3246_; 
wire u0__abc_76628_new_n3247_; 
wire u0__abc_76628_new_n3248_; 
wire u0__abc_76628_new_n3249_; 
wire u0__abc_76628_new_n3251_; 
wire u0__abc_76628_new_n3252_; 
wire u0__abc_76628_new_n3253_; 
wire u0__abc_76628_new_n3254_; 
wire u0__abc_76628_new_n3255_; 
wire u0__abc_76628_new_n3256_; 
wire u0__abc_76628_new_n3257_; 
wire u0__abc_76628_new_n3258_; 
wire u0__abc_76628_new_n3259_; 
wire u0__abc_76628_new_n3260_; 
wire u0__abc_76628_new_n3261_; 
wire u0__abc_76628_new_n3262_; 
wire u0__abc_76628_new_n3263_; 
wire u0__abc_76628_new_n3264_; 
wire u0__abc_76628_new_n3265_; 
wire u0__abc_76628_new_n3266_; 
wire u0__abc_76628_new_n3267_; 
wire u0__abc_76628_new_n3268_; 
wire u0__abc_76628_new_n3269_; 
wire u0__abc_76628_new_n3270_; 
wire u0__abc_76628_new_n3271_; 
wire u0__abc_76628_new_n3272_; 
wire u0__abc_76628_new_n3273_; 
wire u0__abc_76628_new_n3275_; 
wire u0__abc_76628_new_n3276_; 
wire u0__abc_76628_new_n3277_; 
wire u0__abc_76628_new_n3278_; 
wire u0__abc_76628_new_n3279_; 
wire u0__abc_76628_new_n3280_; 
wire u0__abc_76628_new_n3281_; 
wire u0__abc_76628_new_n3282_; 
wire u0__abc_76628_new_n3283_; 
wire u0__abc_76628_new_n3284_; 
wire u0__abc_76628_new_n3285_; 
wire u0__abc_76628_new_n3286_; 
wire u0__abc_76628_new_n3287_; 
wire u0__abc_76628_new_n3288_; 
wire u0__abc_76628_new_n3289_; 
wire u0__abc_76628_new_n3290_; 
wire u0__abc_76628_new_n3291_; 
wire u0__abc_76628_new_n3292_; 
wire u0__abc_76628_new_n3293_; 
wire u0__abc_76628_new_n3294_; 
wire u0__abc_76628_new_n3295_; 
wire u0__abc_76628_new_n3296_; 
wire u0__abc_76628_new_n3297_; 
wire u0__abc_76628_new_n3299_; 
wire u0__abc_76628_new_n3300_; 
wire u0__abc_76628_new_n3301_; 
wire u0__abc_76628_new_n3302_; 
wire u0__abc_76628_new_n3303_; 
wire u0__abc_76628_new_n3304_; 
wire u0__abc_76628_new_n3305_; 
wire u0__abc_76628_new_n3306_; 
wire u0__abc_76628_new_n3307_; 
wire u0__abc_76628_new_n3308_; 
wire u0__abc_76628_new_n3309_; 
wire u0__abc_76628_new_n3310_; 
wire u0__abc_76628_new_n3311_; 
wire u0__abc_76628_new_n3312_; 
wire u0__abc_76628_new_n3313_; 
wire u0__abc_76628_new_n3314_; 
wire u0__abc_76628_new_n3315_; 
wire u0__abc_76628_new_n3316_; 
wire u0__abc_76628_new_n3317_; 
wire u0__abc_76628_new_n3318_; 
wire u0__abc_76628_new_n3319_; 
wire u0__abc_76628_new_n3320_; 
wire u0__abc_76628_new_n3321_; 
wire u0__abc_76628_new_n3323_; 
wire u0__abc_76628_new_n3324_; 
wire u0__abc_76628_new_n3325_; 
wire u0__abc_76628_new_n3326_; 
wire u0__abc_76628_new_n3327_; 
wire u0__abc_76628_new_n3328_; 
wire u0__abc_76628_new_n3329_; 
wire u0__abc_76628_new_n3330_; 
wire u0__abc_76628_new_n3331_; 
wire u0__abc_76628_new_n3332_; 
wire u0__abc_76628_new_n3333_; 
wire u0__abc_76628_new_n3334_; 
wire u0__abc_76628_new_n3335_; 
wire u0__abc_76628_new_n3336_; 
wire u0__abc_76628_new_n3337_; 
wire u0__abc_76628_new_n3338_; 
wire u0__abc_76628_new_n3339_; 
wire u0__abc_76628_new_n3340_; 
wire u0__abc_76628_new_n3341_; 
wire u0__abc_76628_new_n3342_; 
wire u0__abc_76628_new_n3343_; 
wire u0__abc_76628_new_n3344_; 
wire u0__abc_76628_new_n3345_; 
wire u0__abc_76628_new_n3347_; 
wire u0__abc_76628_new_n3348_; 
wire u0__abc_76628_new_n3349_; 
wire u0__abc_76628_new_n3350_; 
wire u0__abc_76628_new_n3351_; 
wire u0__abc_76628_new_n3352_; 
wire u0__abc_76628_new_n3353_; 
wire u0__abc_76628_new_n3354_; 
wire u0__abc_76628_new_n3355_; 
wire u0__abc_76628_new_n3356_; 
wire u0__abc_76628_new_n3357_; 
wire u0__abc_76628_new_n3358_; 
wire u0__abc_76628_new_n3359_; 
wire u0__abc_76628_new_n3360_; 
wire u0__abc_76628_new_n3361_; 
wire u0__abc_76628_new_n3362_; 
wire u0__abc_76628_new_n3363_; 
wire u0__abc_76628_new_n3364_; 
wire u0__abc_76628_new_n3365_; 
wire u0__abc_76628_new_n3366_; 
wire u0__abc_76628_new_n3367_; 
wire u0__abc_76628_new_n3368_; 
wire u0__abc_76628_new_n3369_; 
wire u0__abc_76628_new_n3371_; 
wire u0__abc_76628_new_n3372_; 
wire u0__abc_76628_new_n3373_; 
wire u0__abc_76628_new_n3374_; 
wire u0__abc_76628_new_n3375_; 
wire u0__abc_76628_new_n3376_; 
wire u0__abc_76628_new_n3377_; 
wire u0__abc_76628_new_n3378_; 
wire u0__abc_76628_new_n3379_; 
wire u0__abc_76628_new_n3380_; 
wire u0__abc_76628_new_n3381_; 
wire u0__abc_76628_new_n3382_; 
wire u0__abc_76628_new_n3383_; 
wire u0__abc_76628_new_n3384_; 
wire u0__abc_76628_new_n3385_; 
wire u0__abc_76628_new_n3386_; 
wire u0__abc_76628_new_n3387_; 
wire u0__abc_76628_new_n3388_; 
wire u0__abc_76628_new_n3389_; 
wire u0__abc_76628_new_n3390_; 
wire u0__abc_76628_new_n3391_; 
wire u0__abc_76628_new_n3392_; 
wire u0__abc_76628_new_n3393_; 
wire u0__abc_76628_new_n3515_; 
wire u0__abc_76628_new_n3516_; 
wire u0__abc_76628_new_n3517_; 
wire u0__abc_76628_new_n3518_; 
wire u0__abc_76628_new_n3519_; 
wire u0__abc_76628_new_n3520_; 
wire u0__abc_76628_new_n3521_; 
wire u0__abc_76628_new_n3522_; 
wire u0__abc_76628_new_n3523_; 
wire u0__abc_76628_new_n3524_; 
wire u0__abc_76628_new_n3525_; 
wire u0__abc_76628_new_n3526_; 
wire u0__abc_76628_new_n3527_; 
wire u0__abc_76628_new_n3528_; 
wire u0__abc_76628_new_n3529_; 
wire u0__abc_76628_new_n3530_; 
wire u0__abc_76628_new_n3531_; 
wire u0__abc_76628_new_n3532_; 
wire u0__abc_76628_new_n3533_; 
wire u0__abc_76628_new_n3534_; 
wire u0__abc_76628_new_n3535_; 
wire u0__abc_76628_new_n3536_; 
wire u0__abc_76628_new_n3537_; 
wire u0__abc_76628_new_n3539_; 
wire u0__abc_76628_new_n3540_; 
wire u0__abc_76628_new_n3541_; 
wire u0__abc_76628_new_n3542_; 
wire u0__abc_76628_new_n3543_; 
wire u0__abc_76628_new_n3544_; 
wire u0__abc_76628_new_n3545_; 
wire u0__abc_76628_new_n3546_; 
wire u0__abc_76628_new_n3547_; 
wire u0__abc_76628_new_n3548_; 
wire u0__abc_76628_new_n3549_; 
wire u0__abc_76628_new_n3550_; 
wire u0__abc_76628_new_n3551_; 
wire u0__abc_76628_new_n3552_; 
wire u0__abc_76628_new_n3553_; 
wire u0__abc_76628_new_n3554_; 
wire u0__abc_76628_new_n3555_; 
wire u0__abc_76628_new_n3556_; 
wire u0__abc_76628_new_n3557_; 
wire u0__abc_76628_new_n3558_; 
wire u0__abc_76628_new_n3559_; 
wire u0__abc_76628_new_n3560_; 
wire u0__abc_76628_new_n3561_; 
wire u0__abc_76628_new_n3563_; 
wire u0__abc_76628_new_n3564_; 
wire u0__abc_76628_new_n3565_; 
wire u0__abc_76628_new_n3566_; 
wire u0__abc_76628_new_n3567_; 
wire u0__abc_76628_new_n3568_; 
wire u0__abc_76628_new_n3569_; 
wire u0__abc_76628_new_n3570_; 
wire u0__abc_76628_new_n3571_; 
wire u0__abc_76628_new_n3572_; 
wire u0__abc_76628_new_n3573_; 
wire u0__abc_76628_new_n3574_; 
wire u0__abc_76628_new_n3575_; 
wire u0__abc_76628_new_n3576_; 
wire u0__abc_76628_new_n3577_; 
wire u0__abc_76628_new_n3578_; 
wire u0__abc_76628_new_n3579_; 
wire u0__abc_76628_new_n3580_; 
wire u0__abc_76628_new_n3581_; 
wire u0__abc_76628_new_n3582_; 
wire u0__abc_76628_new_n3583_; 
wire u0__abc_76628_new_n3584_; 
wire u0__abc_76628_new_n3585_; 
wire u0__abc_76628_new_n3587_; 
wire u0__abc_76628_new_n3588_; 
wire u0__abc_76628_new_n3589_; 
wire u0__abc_76628_new_n3590_; 
wire u0__abc_76628_new_n3591_; 
wire u0__abc_76628_new_n3592_; 
wire u0__abc_76628_new_n3593_; 
wire u0__abc_76628_new_n3594_; 
wire u0__abc_76628_new_n3595_; 
wire u0__abc_76628_new_n3596_; 
wire u0__abc_76628_new_n3597_; 
wire u0__abc_76628_new_n3598_; 
wire u0__abc_76628_new_n3599_; 
wire u0__abc_76628_new_n3600_; 
wire u0__abc_76628_new_n3601_; 
wire u0__abc_76628_new_n3602_; 
wire u0__abc_76628_new_n3603_; 
wire u0__abc_76628_new_n3604_; 
wire u0__abc_76628_new_n3605_; 
wire u0__abc_76628_new_n3606_; 
wire u0__abc_76628_new_n3607_; 
wire u0__abc_76628_new_n3608_; 
wire u0__abc_76628_new_n3609_; 
wire u0__abc_76628_new_n3611_; 
wire u0__abc_76628_new_n3612_; 
wire u0__abc_76628_new_n3613_; 
wire u0__abc_76628_new_n3614_; 
wire u0__abc_76628_new_n3615_; 
wire u0__abc_76628_new_n3616_; 
wire u0__abc_76628_new_n3617_; 
wire u0__abc_76628_new_n3618_; 
wire u0__abc_76628_new_n3619_; 
wire u0__abc_76628_new_n3620_; 
wire u0__abc_76628_new_n3621_; 
wire u0__abc_76628_new_n3622_; 
wire u0__abc_76628_new_n3623_; 
wire u0__abc_76628_new_n3624_; 
wire u0__abc_76628_new_n3625_; 
wire u0__abc_76628_new_n3626_; 
wire u0__abc_76628_new_n3627_; 
wire u0__abc_76628_new_n3628_; 
wire u0__abc_76628_new_n3629_; 
wire u0__abc_76628_new_n3630_; 
wire u0__abc_76628_new_n3631_; 
wire u0__abc_76628_new_n3632_; 
wire u0__abc_76628_new_n3633_; 
wire u0__abc_76628_new_n3635_; 
wire u0__abc_76628_new_n3636_; 
wire u0__abc_76628_new_n3637_; 
wire u0__abc_76628_new_n3638_; 
wire u0__abc_76628_new_n3639_; 
wire u0__abc_76628_new_n3640_; 
wire u0__abc_76628_new_n3641_; 
wire u0__abc_76628_new_n3642_; 
wire u0__abc_76628_new_n3643_; 
wire u0__abc_76628_new_n3644_; 
wire u0__abc_76628_new_n3645_; 
wire u0__abc_76628_new_n3646_; 
wire u0__abc_76628_new_n3647_; 
wire u0__abc_76628_new_n3648_; 
wire u0__abc_76628_new_n3649_; 
wire u0__abc_76628_new_n3650_; 
wire u0__abc_76628_new_n3651_; 
wire u0__abc_76628_new_n3652_; 
wire u0__abc_76628_new_n3653_; 
wire u0__abc_76628_new_n3654_; 
wire u0__abc_76628_new_n3655_; 
wire u0__abc_76628_new_n3656_; 
wire u0__abc_76628_new_n3657_; 
wire u0__abc_76628_new_n3659_; 
wire u0__abc_76628_new_n3660_; 
wire u0__abc_76628_new_n3661_; 
wire u0__abc_76628_new_n3662_; 
wire u0__abc_76628_new_n3663_; 
wire u0__abc_76628_new_n3664_; 
wire u0__abc_76628_new_n3665_; 
wire u0__abc_76628_new_n3666_; 
wire u0__abc_76628_new_n3667_; 
wire u0__abc_76628_new_n3668_; 
wire u0__abc_76628_new_n3669_; 
wire u0__abc_76628_new_n3670_; 
wire u0__abc_76628_new_n3671_; 
wire u0__abc_76628_new_n3672_; 
wire u0__abc_76628_new_n3673_; 
wire u0__abc_76628_new_n3674_; 
wire u0__abc_76628_new_n3675_; 
wire u0__abc_76628_new_n3676_; 
wire u0__abc_76628_new_n3677_; 
wire u0__abc_76628_new_n3678_; 
wire u0__abc_76628_new_n3679_; 
wire u0__abc_76628_new_n3680_; 
wire u0__abc_76628_new_n3681_; 
wire u0__abc_76628_new_n3707_; 
wire u0__abc_76628_new_n3708_; 
wire u0__abc_76628_new_n3709_; 
wire u0__abc_76628_new_n3710_; 
wire u0__abc_76628_new_n3711_; 
wire u0__abc_76628_new_n3712_; 
wire u0__abc_76628_new_n3713_; 
wire u0__abc_76628_new_n3714_; 
wire u0__abc_76628_new_n3715_; 
wire u0__abc_76628_new_n3716_; 
wire u0__abc_76628_new_n3717_; 
wire u0__abc_76628_new_n3718_; 
wire u0__abc_76628_new_n3719_; 
wire u0__abc_76628_new_n3720_; 
wire u0__abc_76628_new_n3721_; 
wire u0__abc_76628_new_n3722_; 
wire u0__abc_76628_new_n3723_; 
wire u0__abc_76628_new_n3724_; 
wire u0__abc_76628_new_n3725_; 
wire u0__abc_76628_new_n3726_; 
wire u0__abc_76628_new_n3727_; 
wire u0__abc_76628_new_n3728_; 
wire u0__abc_76628_new_n3729_; 
wire u0__abc_76628_new_n3731_; 
wire u0__abc_76628_new_n3732_; 
wire u0__abc_76628_new_n3733_; 
wire u0__abc_76628_new_n3734_; 
wire u0__abc_76628_new_n3735_; 
wire u0__abc_76628_new_n3736_; 
wire u0__abc_76628_new_n3737_; 
wire u0__abc_76628_new_n3738_; 
wire u0__abc_76628_new_n3739_; 
wire u0__abc_76628_new_n3740_; 
wire u0__abc_76628_new_n3741_; 
wire u0__abc_76628_new_n3742_; 
wire u0__abc_76628_new_n3743_; 
wire u0__abc_76628_new_n3744_; 
wire u0__abc_76628_new_n3745_; 
wire u0__abc_76628_new_n3746_; 
wire u0__abc_76628_new_n3747_; 
wire u0__abc_76628_new_n3748_; 
wire u0__abc_76628_new_n3749_; 
wire u0__abc_76628_new_n3750_; 
wire u0__abc_76628_new_n3751_; 
wire u0__abc_76628_new_n3752_; 
wire u0__abc_76628_new_n3753_; 
wire u0__abc_76628_new_n3755_; 
wire u0__abc_76628_new_n3756_; 
wire u0__abc_76628_new_n3757_; 
wire u0__abc_76628_new_n3758_; 
wire u0__abc_76628_new_n3759_; 
wire u0__abc_76628_new_n3760_; 
wire u0__abc_76628_new_n3761_; 
wire u0__abc_76628_new_n3762_; 
wire u0__abc_76628_new_n3763_; 
wire u0__abc_76628_new_n3764_; 
wire u0__abc_76628_new_n3765_; 
wire u0__abc_76628_new_n3766_; 
wire u0__abc_76628_new_n3767_; 
wire u0__abc_76628_new_n3768_; 
wire u0__abc_76628_new_n3769_; 
wire u0__abc_76628_new_n3770_; 
wire u0__abc_76628_new_n3771_; 
wire u0__abc_76628_new_n3772_; 
wire u0__abc_76628_new_n3773_; 
wire u0__abc_76628_new_n3774_; 
wire u0__abc_76628_new_n3775_; 
wire u0__abc_76628_new_n3776_; 
wire u0__abc_76628_new_n3777_; 
wire u0__abc_76628_new_n4259_; 
wire u0__abc_76628_new_n4260_; 
wire u0__abc_76628_new_n4261_; 
wire u0__abc_76628_new_n4262_; 
wire u0__abc_76628_new_n4263_; 
wire u0__abc_76628_new_n4264_; 
wire u0__abc_76628_new_n4265_; 
wire u0__abc_76628_new_n4266_; 
wire u0__abc_76628_new_n4267_; 
wire u0__abc_76628_new_n4268_; 
wire u0__abc_76628_new_n4269_; 
wire u0__abc_76628_new_n4270_; 
wire u0__abc_76628_new_n4272_; 
wire u0__abc_76628_new_n4273_; 
wire u0__abc_76628_new_n4274_; 
wire u0__abc_76628_new_n4276_; 
wire u0__abc_76628_new_n4277_; 
wire u0__abc_76628_new_n4279_; 
wire u0__abc_76628_new_n4280_; 
wire u0__abc_76628_new_n4282_; 
wire u0__abc_76628_new_n4283_; 
wire u0__abc_76628_new_n4285_; 
wire u0__abc_76628_new_n4286_; 
wire u0__abc_76628_new_n4288_; 
wire u0__abc_76628_new_n4289_; 
wire u0__abc_76628_new_n4291_; 
wire u0__abc_76628_new_n4292_; 
wire u0__abc_76628_new_n4294_; 
wire u0__abc_76628_new_n4295_; 
wire u0__abc_76628_new_n4297_; 
wire u0__abc_76628_new_n4298_; 
wire u0__abc_76628_new_n4298__bF_buf0; 
wire u0__abc_76628_new_n4298__bF_buf1; 
wire u0__abc_76628_new_n4298__bF_buf2; 
wire u0__abc_76628_new_n4298__bF_buf3; 
wire u0__abc_76628_new_n4298__bF_buf4; 
wire u0__abc_76628_new_n4299_; 
wire u0__abc_76628_new_n4301_; 
wire u0__abc_76628_new_n4302_; 
wire u0__abc_76628_new_n4304_; 
wire u0__abc_76628_new_n4305_; 
wire u0__abc_76628_new_n4307_; 
wire u0__abc_76628_new_n4308_; 
wire u0__abc_76628_new_n4310_; 
wire u0__abc_76628_new_n4311_; 
wire u0__abc_76628_new_n4313_; 
wire u0__abc_76628_new_n4314_; 
wire u0__abc_76628_new_n4316_; 
wire u0__abc_76628_new_n4317_; 
wire u0__abc_76628_new_n4319_; 
wire u0__abc_76628_new_n4320_; 
wire u0__abc_76628_new_n4322_; 
wire u0__abc_76628_new_n4323_; 
wire u0__abc_76628_new_n4325_; 
wire u0__abc_76628_new_n4326_; 
wire u0__abc_76628_new_n4328_; 
wire u0__abc_76628_new_n4329_; 
wire u0__abc_76628_new_n4331_; 
wire u0__abc_76628_new_n4332_; 
wire u0__abc_76628_new_n4334_; 
wire u0__abc_76628_new_n4335_; 
wire u0__abc_76628_new_n4337_; 
wire u0__abc_76628_new_n4338_; 
wire u0__abc_76628_new_n4340_; 
wire u0__abc_76628_new_n4341_; 
wire u0__abc_76628_new_n4343_; 
wire u0__abc_76628_new_n4344_; 
wire u0__abc_76628_new_n4346_; 
wire u0__abc_76628_new_n4347_; 
wire u0__abc_76628_new_n4349_; 
wire u0__abc_76628_new_n4350_; 
wire u0__abc_76628_new_n4352_; 
wire u0__abc_76628_new_n4353_; 
wire u0__abc_76628_new_n4355_; 
wire u0__abc_76628_new_n4356_; 
wire u0__abc_76628_new_n4358_; 
wire u0__abc_76628_new_n4359_; 
wire u0__abc_76628_new_n4361_; 
wire u0__abc_76628_new_n4362_; 
wire u0__abc_76628_new_n4364_; 
wire u0__abc_76628_new_n4365_; 
wire u0__abc_76628_new_n4367_; 
wire u0__abc_76628_new_n4368_; 
wire u0__abc_76628_new_n4370_; 
wire u0__abc_76628_new_n4371_; 
wire u0__abc_76628_new_n4373_; 
wire u0__abc_76628_new_n4374_; 
wire u0__abc_76628_new_n4376_; 
wire u0__abc_76628_new_n4377_; 
wire u0__abc_76628_new_n4379_; 
wire u0__abc_76628_new_n4380_; 
wire u0__abc_76628_new_n4382_; 
wire u0__abc_76628_new_n4383_; 
wire u0__abc_76628_new_n4385_; 
wire u0__abc_76628_new_n4386_; 
wire u0__abc_76628_new_n4388_; 
wire u0__abc_76628_new_n4389_; 
wire u0__abc_76628_new_n4391_; 
wire u0__abc_76628_new_n4392_; 
wire u0__abc_76628_new_n4394_; 
wire u0__abc_76628_new_n4395_; 
wire u0__abc_76628_new_n4396_; 
wire u0__abc_76628_new_n4397_; 
wire u0__abc_76628_new_n4398_; 
wire u0__abc_76628_new_n4399_; 
wire u0__abc_76628_new_n4400_; 
wire u0__abc_76628_new_n4401_; 
wire u0__abc_76628_new_n4402_; 
wire u0__abc_76628_new_n4403_; 
wire u0__abc_76628_new_n4404_; 
wire u0__abc_76628_new_n4406_; 
wire u0__abc_76628_new_n4407_; 
wire u0__abc_76628_new_n4409_; 
wire u0__abc_76628_new_n4410_; 
wire u0__abc_76628_new_n4412_; 
wire u0__abc_76628_new_n4413_; 
wire u0__abc_76628_new_n4415_; 
wire u0__abc_76628_new_n4416_; 
wire u0__abc_76628_new_n4418_; 
wire u0__abc_76628_new_n4419_; 
wire u0__abc_76628_new_n4421_; 
wire u0__abc_76628_new_n4422_; 
wire u0__abc_76628_new_n4424_; 
wire u0__abc_76628_new_n4425_; 
wire u0__abc_76628_new_n4427_; 
wire u0__abc_76628_new_n4428_; 
wire u0__abc_76628_new_n4430_; 
wire u0__abc_76628_new_n4431_; 
wire u0__abc_76628_new_n4433_; 
wire u0__abc_76628_new_n4434_; 
wire u0__abc_76628_new_n4436_; 
wire u0__abc_76628_new_n4437_; 
wire u0__abc_76628_new_n4437__bF_buf0; 
wire u0__abc_76628_new_n4437__bF_buf1; 
wire u0__abc_76628_new_n4437__bF_buf2; 
wire u0__abc_76628_new_n4437__bF_buf3; 
wire u0__abc_76628_new_n4438_; 
wire u0__abc_76628_new_n4438__bF_buf0; 
wire u0__abc_76628_new_n4438__bF_buf1; 
wire u0__abc_76628_new_n4438__bF_buf2; 
wire u0__abc_76628_new_n4438__bF_buf3; 
wire u0__abc_76628_new_n4439_; 
wire u0__abc_76628_new_n4440_; 
wire u0__abc_76628_new_n4442_; 
wire u0__abc_76628_new_n4443_; 
wire u0__abc_76628_new_n4445_; 
wire u0__abc_76628_new_n4446_; 
wire u0__abc_76628_new_n4448_; 
wire u0__abc_76628_new_n4449_; 
wire u0__abc_76628_new_n4451_; 
wire u0__abc_76628_new_n4452_; 
wire u0__abc_76628_new_n4454_; 
wire u0__abc_76628_new_n4455_; 
wire u0__abc_76628_new_n4457_; 
wire u0__abc_76628_new_n4458_; 
wire u0__abc_76628_new_n4460_; 
wire u0__abc_76628_new_n4461_; 
wire u0__abc_76628_new_n4463_; 
wire u0__abc_76628_new_n4464_; 
wire u0__abc_76628_new_n4466_; 
wire u0__abc_76628_new_n4467_; 
wire u0__abc_76628_new_n4469_; 
wire u0__abc_76628_new_n4470_; 
wire u0__abc_76628_new_n4472_; 
wire u0__abc_76628_new_n4473_; 
wire u0__abc_76628_new_n4475_; 
wire u0__abc_76628_new_n4476_; 
wire u0__abc_76628_new_n4478_; 
wire u0__abc_76628_new_n4479_; 
wire u0__abc_76628_new_n4481_; 
wire u0__abc_76628_new_n4482_; 
wire u0__abc_76628_new_n4484_; 
wire u0__abc_76628_new_n4485_; 
wire u0__abc_76628_new_n4487_; 
wire u0__abc_76628_new_n4488_; 
wire u0__abc_76628_new_n4490_; 
wire u0__abc_76628_new_n4491_; 
wire u0__abc_76628_new_n4493_; 
wire u0__abc_76628_new_n4494_; 
wire u0__abc_76628_new_n4495_; 
wire u0__abc_76628_new_n4496_; 
wire u0__abc_76628_new_n4497_; 
wire u0__abc_76628_new_n4498_; 
wire u0__abc_76628_new_n4499_; 
wire u0__abc_76628_new_n4500_; 
wire u0__abc_76628_new_n4500__bF_buf0; 
wire u0__abc_76628_new_n4500__bF_buf1; 
wire u0__abc_76628_new_n4500__bF_buf2; 
wire u0__abc_76628_new_n4500__bF_buf3; 
wire u0__abc_76628_new_n4500__bF_buf4; 
wire u0__abc_76628_new_n4501_; 
wire u0__abc_76628_new_n4502_; 
wire u0__abc_76628_new_n4503_; 
wire u0__abc_76628_new_n4503__bF_buf0; 
wire u0__abc_76628_new_n4503__bF_buf1; 
wire u0__abc_76628_new_n4503__bF_buf2; 
wire u0__abc_76628_new_n4503__bF_buf3; 
wire u0__abc_76628_new_n4503__bF_buf4; 
wire u0__abc_76628_new_n4504_; 
wire u0__abc_76628_new_n4505_; 
wire u0__abc_76628_new_n4506_; 
wire u0__abc_76628_new_n4507_; 
wire u0__abc_76628_new_n4507__bF_buf0; 
wire u0__abc_76628_new_n4507__bF_buf1; 
wire u0__abc_76628_new_n4507__bF_buf2; 
wire u0__abc_76628_new_n4507__bF_buf3; 
wire u0__abc_76628_new_n4507__bF_buf4; 
wire u0__abc_76628_new_n4508_; 
wire u0__abc_76628_new_n4509_; 
wire u0__abc_76628_new_n4510_; 
wire u0__abc_76628_new_n4510__bF_buf0; 
wire u0__abc_76628_new_n4510__bF_buf1; 
wire u0__abc_76628_new_n4510__bF_buf2; 
wire u0__abc_76628_new_n4510__bF_buf3; 
wire u0__abc_76628_new_n4510__bF_buf4; 
wire u0__abc_76628_new_n4511_; 
wire u0__abc_76628_new_n4512_; 
wire u0__abc_76628_new_n4513_; 
wire u0__abc_76628_new_n4514_; 
wire u0__abc_76628_new_n4515_; 
wire u0__abc_76628_new_n4516_; 
wire u0__abc_76628_new_n4517_; 
wire u0__abc_76628_new_n4517__bF_buf0; 
wire u0__abc_76628_new_n4517__bF_buf1; 
wire u0__abc_76628_new_n4517__bF_buf2; 
wire u0__abc_76628_new_n4517__bF_buf3; 
wire u0__abc_76628_new_n4517__bF_buf4; 
wire u0__abc_76628_new_n4518_; 
wire u0__abc_76628_new_n4519_; 
wire u0__abc_76628_new_n4520_; 
wire u0__abc_76628_new_n4520__bF_buf0; 
wire u0__abc_76628_new_n4520__bF_buf1; 
wire u0__abc_76628_new_n4520__bF_buf2; 
wire u0__abc_76628_new_n4520__bF_buf3; 
wire u0__abc_76628_new_n4520__bF_buf4; 
wire u0__abc_76628_new_n4521_; 
wire u0__abc_76628_new_n4522_; 
wire u0__abc_76628_new_n4523_; 
wire u0__abc_76628_new_n4523__bF_buf0; 
wire u0__abc_76628_new_n4523__bF_buf1; 
wire u0__abc_76628_new_n4523__bF_buf2; 
wire u0__abc_76628_new_n4523__bF_buf3; 
wire u0__abc_76628_new_n4523__bF_buf4; 
wire u0__abc_76628_new_n4524_; 
wire u0__abc_76628_new_n4525_; 
wire u0__abc_76628_new_n4526_; 
wire u0__abc_76628_new_n4527_; 
wire u0__abc_76628_new_n4528_; 
wire u0__abc_76628_new_n4528__bF_buf0; 
wire u0__abc_76628_new_n4528__bF_buf1; 
wire u0__abc_76628_new_n4528__bF_buf2; 
wire u0__abc_76628_new_n4528__bF_buf3; 
wire u0__abc_76628_new_n4528__bF_buf4; 
wire u0__abc_76628_new_n4529_; 
wire u0__abc_76628_new_n4530_; 
wire u0__abc_76628_new_n4531_; 
wire u0__abc_76628_new_n4531__bF_buf0; 
wire u0__abc_76628_new_n4531__bF_buf1; 
wire u0__abc_76628_new_n4531__bF_buf2; 
wire u0__abc_76628_new_n4531__bF_buf3; 
wire u0__abc_76628_new_n4531__bF_buf4; 
wire u0__abc_76628_new_n4532_; 
wire u0__abc_76628_new_n4533_; 
wire u0__abc_76628_new_n4534_; 
wire u0__abc_76628_new_n4535_; 
wire u0__abc_76628_new_n4536_; 
wire u0__abc_76628_new_n4537_; 
wire u0__abc_76628_new_n4538_; 
wire u0__abc_76628_new_n4539_; 
wire u0__abc_76628_new_n4540_; 
wire u0__abc_76628_new_n4541_; 
wire u0__abc_76628_new_n4541__bF_buf0; 
wire u0__abc_76628_new_n4541__bF_buf1; 
wire u0__abc_76628_new_n4541__bF_buf2; 
wire u0__abc_76628_new_n4541__bF_buf3; 
wire u0__abc_76628_new_n4542_; 
wire u0__abc_76628_new_n4543_; 
wire u0__abc_76628_new_n4544_; 
wire u0__abc_76628_new_n4545_; 
wire u0__abc_76628_new_n4545__bF_buf0; 
wire u0__abc_76628_new_n4545__bF_buf1; 
wire u0__abc_76628_new_n4545__bF_buf2; 
wire u0__abc_76628_new_n4545__bF_buf3; 
wire u0__abc_76628_new_n4545__bF_buf4; 
wire u0__abc_76628_new_n4546_; 
wire u0__abc_76628_new_n4547_; 
wire u0__abc_76628_new_n4547__bF_buf0; 
wire u0__abc_76628_new_n4547__bF_buf1; 
wire u0__abc_76628_new_n4547__bF_buf2; 
wire u0__abc_76628_new_n4547__bF_buf3; 
wire u0__abc_76628_new_n4547__bF_buf4; 
wire u0__abc_76628_new_n4548_; 
wire u0__abc_76628_new_n4549_; 
wire u0__abc_76628_new_n4549__bF_buf0; 
wire u0__abc_76628_new_n4549__bF_buf1; 
wire u0__abc_76628_new_n4549__bF_buf2; 
wire u0__abc_76628_new_n4549__bF_buf3; 
wire u0__abc_76628_new_n4549__bF_buf4; 
wire u0__abc_76628_new_n4550_; 
wire u0__abc_76628_new_n4551_; 
wire u0__abc_76628_new_n4552_; 
wire u0__abc_76628_new_n4553_; 
wire u0__abc_76628_new_n4554_; 
wire u0__abc_76628_new_n4554__bF_buf0; 
wire u0__abc_76628_new_n4554__bF_buf1; 
wire u0__abc_76628_new_n4554__bF_buf2; 
wire u0__abc_76628_new_n4554__bF_buf3; 
wire u0__abc_76628_new_n4554__bF_buf4; 
wire u0__abc_76628_new_n4555_; 
wire u0__abc_76628_new_n4556_; 
wire u0__abc_76628_new_n4556__bF_buf0; 
wire u0__abc_76628_new_n4556__bF_buf1; 
wire u0__abc_76628_new_n4556__bF_buf2; 
wire u0__abc_76628_new_n4556__bF_buf3; 
wire u0__abc_76628_new_n4556__bF_buf4; 
wire u0__abc_76628_new_n4557_; 
wire u0__abc_76628_new_n4558_; 
wire u0__abc_76628_new_n4558__bF_buf0; 
wire u0__abc_76628_new_n4558__bF_buf1; 
wire u0__abc_76628_new_n4558__bF_buf2; 
wire u0__abc_76628_new_n4558__bF_buf3; 
wire u0__abc_76628_new_n4558__bF_buf4; 
wire u0__abc_76628_new_n4559_; 
wire u0__abc_76628_new_n4560_; 
wire u0__abc_76628_new_n4561_; 
wire u0__abc_76628_new_n4562_; 
wire u0__abc_76628_new_n4562__bF_buf0; 
wire u0__abc_76628_new_n4562__bF_buf1; 
wire u0__abc_76628_new_n4562__bF_buf2; 
wire u0__abc_76628_new_n4562__bF_buf3; 
wire u0__abc_76628_new_n4562__bF_buf4; 
wire u0__abc_76628_new_n4563_; 
wire u0__abc_76628_new_n4564_; 
wire u0__abc_76628_new_n4565_; 
wire u0__abc_76628_new_n4566_; 
wire u0__abc_76628_new_n4566__bF_buf0; 
wire u0__abc_76628_new_n4566__bF_buf1; 
wire u0__abc_76628_new_n4566__bF_buf2; 
wire u0__abc_76628_new_n4566__bF_buf3; 
wire u0__abc_76628_new_n4566__bF_buf4; 
wire u0__abc_76628_new_n4567_; 
wire u0__abc_76628_new_n4568_; 
wire u0__abc_76628_new_n4569_; 
wire u0__abc_76628_new_n4570_; 
wire u0__abc_76628_new_n4571_; 
wire u0__abc_76628_new_n4573_; 
wire u0__abc_76628_new_n4574_; 
wire u0__abc_76628_new_n4575_; 
wire u0__abc_76628_new_n4576_; 
wire u0__abc_76628_new_n4577_; 
wire u0__abc_76628_new_n4578_; 
wire u0__abc_76628_new_n4579_; 
wire u0__abc_76628_new_n4580_; 
wire u0__abc_76628_new_n4581_; 
wire u0__abc_76628_new_n4582_; 
wire u0__abc_76628_new_n4583_; 
wire u0__abc_76628_new_n4584_; 
wire u0__abc_76628_new_n4585_; 
wire u0__abc_76628_new_n4586_; 
wire u0__abc_76628_new_n4587_; 
wire u0__abc_76628_new_n4588_; 
wire u0__abc_76628_new_n4589_; 
wire u0__abc_76628_new_n4590_; 
wire u0__abc_76628_new_n4591_; 
wire u0__abc_76628_new_n4592_; 
wire u0__abc_76628_new_n4593_; 
wire u0__abc_76628_new_n4594_; 
wire u0__abc_76628_new_n4595_; 
wire u0__abc_76628_new_n4596_; 
wire u0__abc_76628_new_n4597_; 
wire u0__abc_76628_new_n4598_; 
wire u0__abc_76628_new_n4599_; 
wire u0__abc_76628_new_n4600_; 
wire u0__abc_76628_new_n4601_; 
wire u0__abc_76628_new_n4602_; 
wire u0__abc_76628_new_n4603_; 
wire u0__abc_76628_new_n4604_; 
wire u0__abc_76628_new_n4605_; 
wire u0__abc_76628_new_n4606_; 
wire u0__abc_76628_new_n4607_; 
wire u0__abc_76628_new_n4608_; 
wire u0__abc_76628_new_n4610_; 
wire u0__abc_76628_new_n4611_; 
wire u0__abc_76628_new_n4612_; 
wire u0__abc_76628_new_n4613_; 
wire u0__abc_76628_new_n4614_; 
wire u0__abc_76628_new_n4615_; 
wire u0__abc_76628_new_n4616_; 
wire u0__abc_76628_new_n4617_; 
wire u0__abc_76628_new_n4618_; 
wire u0__abc_76628_new_n4619_; 
wire u0__abc_76628_new_n4620_; 
wire u0__abc_76628_new_n4621_; 
wire u0__abc_76628_new_n4622_; 
wire u0__abc_76628_new_n4623_; 
wire u0__abc_76628_new_n4624_; 
wire u0__abc_76628_new_n4625_; 
wire u0__abc_76628_new_n4626_; 
wire u0__abc_76628_new_n4627_; 
wire u0__abc_76628_new_n4628_; 
wire u0__abc_76628_new_n4629_; 
wire u0__abc_76628_new_n4630_; 
wire u0__abc_76628_new_n4631_; 
wire u0__abc_76628_new_n4632_; 
wire u0__abc_76628_new_n4633_; 
wire u0__abc_76628_new_n4634_; 
wire u0__abc_76628_new_n4635_; 
wire u0__abc_76628_new_n4636_; 
wire u0__abc_76628_new_n4637_; 
wire u0__abc_76628_new_n4638_; 
wire u0__abc_76628_new_n4639_; 
wire u0__abc_76628_new_n4640_; 
wire u0__abc_76628_new_n4641_; 
wire u0__abc_76628_new_n4642_; 
wire u0__abc_76628_new_n4643_; 
wire u0__abc_76628_new_n4644_; 
wire u0__abc_76628_new_n4645_; 
wire u0__abc_76628_new_n4647_; 
wire u0__abc_76628_new_n4648_; 
wire u0__abc_76628_new_n4649_; 
wire u0__abc_76628_new_n4650_; 
wire u0__abc_76628_new_n4651_; 
wire u0__abc_76628_new_n4652_; 
wire u0__abc_76628_new_n4653_; 
wire u0__abc_76628_new_n4654_; 
wire u0__abc_76628_new_n4655_; 
wire u0__abc_76628_new_n4656_; 
wire u0__abc_76628_new_n4657_; 
wire u0__abc_76628_new_n4658_; 
wire u0__abc_76628_new_n4659_; 
wire u0__abc_76628_new_n4660_; 
wire u0__abc_76628_new_n4661_; 
wire u0__abc_76628_new_n4662_; 
wire u0__abc_76628_new_n4663_; 
wire u0__abc_76628_new_n4664_; 
wire u0__abc_76628_new_n4665_; 
wire u0__abc_76628_new_n4666_; 
wire u0__abc_76628_new_n4667_; 
wire u0__abc_76628_new_n4668_; 
wire u0__abc_76628_new_n4669_; 
wire u0__abc_76628_new_n4670_; 
wire u0__abc_76628_new_n4671_; 
wire u0__abc_76628_new_n4672_; 
wire u0__abc_76628_new_n4673_; 
wire u0__abc_76628_new_n4674_; 
wire u0__abc_76628_new_n4675_; 
wire u0__abc_76628_new_n4676_; 
wire u0__abc_76628_new_n4677_; 
wire u0__abc_76628_new_n4678_; 
wire u0__abc_76628_new_n4679_; 
wire u0__abc_76628_new_n4680_; 
wire u0__abc_76628_new_n4681_; 
wire u0__abc_76628_new_n4682_; 
wire u0__abc_76628_new_n4684_; 
wire u0__abc_76628_new_n4685_; 
wire u0__abc_76628_new_n4686_; 
wire u0__abc_76628_new_n4687_; 
wire u0__abc_76628_new_n4688_; 
wire u0__abc_76628_new_n4689_; 
wire u0__abc_76628_new_n4690_; 
wire u0__abc_76628_new_n4691_; 
wire u0__abc_76628_new_n4692_; 
wire u0__abc_76628_new_n4693_; 
wire u0__abc_76628_new_n4694_; 
wire u0__abc_76628_new_n4695_; 
wire u0__abc_76628_new_n4696_; 
wire u0__abc_76628_new_n4697_; 
wire u0__abc_76628_new_n4698_; 
wire u0__abc_76628_new_n4699_; 
wire u0__abc_76628_new_n4700_; 
wire u0__abc_76628_new_n4701_; 
wire u0__abc_76628_new_n4702_; 
wire u0__abc_76628_new_n4703_; 
wire u0__abc_76628_new_n4704_; 
wire u0__abc_76628_new_n4705_; 
wire u0__abc_76628_new_n4706_; 
wire u0__abc_76628_new_n4707_; 
wire u0__abc_76628_new_n4708_; 
wire u0__abc_76628_new_n4709_; 
wire u0__abc_76628_new_n4710_; 
wire u0__abc_76628_new_n4711_; 
wire u0__abc_76628_new_n4712_; 
wire u0__abc_76628_new_n4713_; 
wire u0__abc_76628_new_n4714_; 
wire u0__abc_76628_new_n4715_; 
wire u0__abc_76628_new_n4716_; 
wire u0__abc_76628_new_n4717_; 
wire u0__abc_76628_new_n4718_; 
wire u0__abc_76628_new_n4719_; 
wire u0__abc_76628_new_n4721_; 
wire u0__abc_76628_new_n4722_; 
wire u0__abc_76628_new_n4723_; 
wire u0__abc_76628_new_n4724_; 
wire u0__abc_76628_new_n4725_; 
wire u0__abc_76628_new_n4726_; 
wire u0__abc_76628_new_n4727_; 
wire u0__abc_76628_new_n4728_; 
wire u0__abc_76628_new_n4729_; 
wire u0__abc_76628_new_n4730_; 
wire u0__abc_76628_new_n4731_; 
wire u0__abc_76628_new_n4732_; 
wire u0__abc_76628_new_n4733_; 
wire u0__abc_76628_new_n4734_; 
wire u0__abc_76628_new_n4735_; 
wire u0__abc_76628_new_n4736_; 
wire u0__abc_76628_new_n4737_; 
wire u0__abc_76628_new_n4738_; 
wire u0__abc_76628_new_n4739_; 
wire u0__abc_76628_new_n4740_; 
wire u0__abc_76628_new_n4741_; 
wire u0__abc_76628_new_n4742_; 
wire u0__abc_76628_new_n4743_; 
wire u0__abc_76628_new_n4744_; 
wire u0__abc_76628_new_n4745_; 
wire u0__abc_76628_new_n4746_; 
wire u0__abc_76628_new_n4747_; 
wire u0__abc_76628_new_n4748_; 
wire u0__abc_76628_new_n4749_; 
wire u0__abc_76628_new_n4750_; 
wire u0__abc_76628_new_n4751_; 
wire u0__abc_76628_new_n4752_; 
wire u0__abc_76628_new_n4753_; 
wire u0__abc_76628_new_n4754_; 
wire u0__abc_76628_new_n4755_; 
wire u0__abc_76628_new_n4756_; 
wire u0__abc_76628_new_n4758_; 
wire u0__abc_76628_new_n4759_; 
wire u0__abc_76628_new_n4760_; 
wire u0__abc_76628_new_n4761_; 
wire u0__abc_76628_new_n4762_; 
wire u0__abc_76628_new_n4763_; 
wire u0__abc_76628_new_n4764_; 
wire u0__abc_76628_new_n4765_; 
wire u0__abc_76628_new_n4766_; 
wire u0__abc_76628_new_n4767_; 
wire u0__abc_76628_new_n4768_; 
wire u0__abc_76628_new_n4769_; 
wire u0__abc_76628_new_n4770_; 
wire u0__abc_76628_new_n4771_; 
wire u0__abc_76628_new_n4772_; 
wire u0__abc_76628_new_n4773_; 
wire u0__abc_76628_new_n4774_; 
wire u0__abc_76628_new_n4775_; 
wire u0__abc_76628_new_n4776_; 
wire u0__abc_76628_new_n4777_; 
wire u0__abc_76628_new_n4778_; 
wire u0__abc_76628_new_n4779_; 
wire u0__abc_76628_new_n4780_; 
wire u0__abc_76628_new_n4781_; 
wire u0__abc_76628_new_n4782_; 
wire u0__abc_76628_new_n4783_; 
wire u0__abc_76628_new_n4784_; 
wire u0__abc_76628_new_n4785_; 
wire u0__abc_76628_new_n4786_; 
wire u0__abc_76628_new_n4787_; 
wire u0__abc_76628_new_n4788_; 
wire u0__abc_76628_new_n4789_; 
wire u0__abc_76628_new_n4790_; 
wire u0__abc_76628_new_n4791_; 
wire u0__abc_76628_new_n4792_; 
wire u0__abc_76628_new_n4793_; 
wire u0__abc_76628_new_n4795_; 
wire u0__abc_76628_new_n4796_; 
wire u0__abc_76628_new_n4797_; 
wire u0__abc_76628_new_n4798_; 
wire u0__abc_76628_new_n4799_; 
wire u0__abc_76628_new_n4800_; 
wire u0__abc_76628_new_n4801_; 
wire u0__abc_76628_new_n4802_; 
wire u0__abc_76628_new_n4803_; 
wire u0__abc_76628_new_n4804_; 
wire u0__abc_76628_new_n4805_; 
wire u0__abc_76628_new_n4806_; 
wire u0__abc_76628_new_n4807_; 
wire u0__abc_76628_new_n4808_; 
wire u0__abc_76628_new_n4809_; 
wire u0__abc_76628_new_n4810_; 
wire u0__abc_76628_new_n4811_; 
wire u0__abc_76628_new_n4812_; 
wire u0__abc_76628_new_n4813_; 
wire u0__abc_76628_new_n4814_; 
wire u0__abc_76628_new_n4815_; 
wire u0__abc_76628_new_n4816_; 
wire u0__abc_76628_new_n4817_; 
wire u0__abc_76628_new_n4818_; 
wire u0__abc_76628_new_n4819_; 
wire u0__abc_76628_new_n4820_; 
wire u0__abc_76628_new_n4821_; 
wire u0__abc_76628_new_n4822_; 
wire u0__abc_76628_new_n4823_; 
wire u0__abc_76628_new_n4824_; 
wire u0__abc_76628_new_n4825_; 
wire u0__abc_76628_new_n4826_; 
wire u0__abc_76628_new_n4827_; 
wire u0__abc_76628_new_n4828_; 
wire u0__abc_76628_new_n4829_; 
wire u0__abc_76628_new_n4830_; 
wire u0__abc_76628_new_n4832_; 
wire u0__abc_76628_new_n4833_; 
wire u0__abc_76628_new_n4834_; 
wire u0__abc_76628_new_n4835_; 
wire u0__abc_76628_new_n4836_; 
wire u0__abc_76628_new_n4837_; 
wire u0__abc_76628_new_n4838_; 
wire u0__abc_76628_new_n4839_; 
wire u0__abc_76628_new_n4840_; 
wire u0__abc_76628_new_n4841_; 
wire u0__abc_76628_new_n4842_; 
wire u0__abc_76628_new_n4843_; 
wire u0__abc_76628_new_n4844_; 
wire u0__abc_76628_new_n4845_; 
wire u0__abc_76628_new_n4846_; 
wire u0__abc_76628_new_n4847_; 
wire u0__abc_76628_new_n4848_; 
wire u0__abc_76628_new_n4849_; 
wire u0__abc_76628_new_n4850_; 
wire u0__abc_76628_new_n4851_; 
wire u0__abc_76628_new_n4852_; 
wire u0__abc_76628_new_n4853_; 
wire u0__abc_76628_new_n4854_; 
wire u0__abc_76628_new_n4855_; 
wire u0__abc_76628_new_n4856_; 
wire u0__abc_76628_new_n4857_; 
wire u0__abc_76628_new_n4858_; 
wire u0__abc_76628_new_n4859_; 
wire u0__abc_76628_new_n4860_; 
wire u0__abc_76628_new_n4861_; 
wire u0__abc_76628_new_n4862_; 
wire u0__abc_76628_new_n4863_; 
wire u0__abc_76628_new_n4864_; 
wire u0__abc_76628_new_n4865_; 
wire u0__abc_76628_new_n4866_; 
wire u0__abc_76628_new_n4867_; 
wire u0__abc_76628_new_n4869_; 
wire u0__abc_76628_new_n4870_; 
wire u0__abc_76628_new_n4871_; 
wire u0__abc_76628_new_n4872_; 
wire u0__abc_76628_new_n4873_; 
wire u0__abc_76628_new_n4874_; 
wire u0__abc_76628_new_n4875_; 
wire u0__abc_76628_new_n4876_; 
wire u0__abc_76628_new_n4877_; 
wire u0__abc_76628_new_n4878_; 
wire u0__abc_76628_new_n4879_; 
wire u0__abc_76628_new_n4880_; 
wire u0__abc_76628_new_n4881_; 
wire u0__abc_76628_new_n4882_; 
wire u0__abc_76628_new_n4883_; 
wire u0__abc_76628_new_n4884_; 
wire u0__abc_76628_new_n4885_; 
wire u0__abc_76628_new_n4886_; 
wire u0__abc_76628_new_n4887_; 
wire u0__abc_76628_new_n4888_; 
wire u0__abc_76628_new_n4889_; 
wire u0__abc_76628_new_n4890_; 
wire u0__abc_76628_new_n4891_; 
wire u0__abc_76628_new_n4892_; 
wire u0__abc_76628_new_n4893_; 
wire u0__abc_76628_new_n4894_; 
wire u0__abc_76628_new_n4895_; 
wire u0__abc_76628_new_n4896_; 
wire u0__abc_76628_new_n4897_; 
wire u0__abc_76628_new_n4898_; 
wire u0__abc_76628_new_n4899_; 
wire u0__abc_76628_new_n4900_; 
wire u0__abc_76628_new_n4901_; 
wire u0__abc_76628_new_n4902_; 
wire u0__abc_76628_new_n4903_; 
wire u0__abc_76628_new_n4904_; 
wire u0__abc_76628_new_n4906_; 
wire u0__abc_76628_new_n4907_; 
wire u0__abc_76628_new_n4908_; 
wire u0__abc_76628_new_n4909_; 
wire u0__abc_76628_new_n4910_; 
wire u0__abc_76628_new_n4911_; 
wire u0__abc_76628_new_n4912_; 
wire u0__abc_76628_new_n4913_; 
wire u0__abc_76628_new_n4914_; 
wire u0__abc_76628_new_n4915_; 
wire u0__abc_76628_new_n4916_; 
wire u0__abc_76628_new_n4917_; 
wire u0__abc_76628_new_n4918_; 
wire u0__abc_76628_new_n4919_; 
wire u0__abc_76628_new_n4920_; 
wire u0__abc_76628_new_n4921_; 
wire u0__abc_76628_new_n4922_; 
wire u0__abc_76628_new_n4923_; 
wire u0__abc_76628_new_n4924_; 
wire u0__abc_76628_new_n4925_; 
wire u0__abc_76628_new_n4926_; 
wire u0__abc_76628_new_n4927_; 
wire u0__abc_76628_new_n4928_; 
wire u0__abc_76628_new_n4929_; 
wire u0__abc_76628_new_n4930_; 
wire u0__abc_76628_new_n4931_; 
wire u0__abc_76628_new_n4932_; 
wire u0__abc_76628_new_n4933_; 
wire u0__abc_76628_new_n4934_; 
wire u0__abc_76628_new_n4935_; 
wire u0__abc_76628_new_n4936_; 
wire u0__abc_76628_new_n4937_; 
wire u0__abc_76628_new_n4938_; 
wire u0__abc_76628_new_n4939_; 
wire u0__abc_76628_new_n4940_; 
wire u0__abc_76628_new_n4941_; 
wire u0__abc_76628_new_n4943_; 
wire u0__abc_76628_new_n4944_; 
wire u0__abc_76628_new_n4945_; 
wire u0__abc_76628_new_n4946_; 
wire u0__abc_76628_new_n4947_; 
wire u0__abc_76628_new_n4948_; 
wire u0__abc_76628_new_n4949_; 
wire u0__abc_76628_new_n4950_; 
wire u0__abc_76628_new_n4951_; 
wire u0__abc_76628_new_n4952_; 
wire u0__abc_76628_new_n4953_; 
wire u0__abc_76628_new_n4954_; 
wire u0__abc_76628_new_n4955_; 
wire u0__abc_76628_new_n4956_; 
wire u0__abc_76628_new_n4957_; 
wire u0__abc_76628_new_n4958_; 
wire u0__abc_76628_new_n4959_; 
wire u0__abc_76628_new_n4960_; 
wire u0__abc_76628_new_n4961_; 
wire u0__abc_76628_new_n4962_; 
wire u0__abc_76628_new_n4963_; 
wire u0__abc_76628_new_n4964_; 
wire u0__abc_76628_new_n4965_; 
wire u0__abc_76628_new_n4966_; 
wire u0__abc_76628_new_n4967_; 
wire u0__abc_76628_new_n4968_; 
wire u0__abc_76628_new_n4969_; 
wire u0__abc_76628_new_n4970_; 
wire u0__abc_76628_new_n4971_; 
wire u0__abc_76628_new_n4972_; 
wire u0__abc_76628_new_n4973_; 
wire u0__abc_76628_new_n4974_; 
wire u0__abc_76628_new_n4976_; 
wire u0__abc_76628_new_n4977_; 
wire u0__abc_76628_new_n4978_; 
wire u0__abc_76628_new_n4979_; 
wire u0__abc_76628_new_n4980_; 
wire u0__abc_76628_new_n4981_; 
wire u0__abc_76628_new_n4982_; 
wire u0__abc_76628_new_n4983_; 
wire u0__abc_76628_new_n4984_; 
wire u0__abc_76628_new_n4985_; 
wire u0__abc_76628_new_n4986_; 
wire u0__abc_76628_new_n4987_; 
wire u0__abc_76628_new_n4988_; 
wire u0__abc_76628_new_n4989_; 
wire u0__abc_76628_new_n4990_; 
wire u0__abc_76628_new_n4991_; 
wire u0__abc_76628_new_n4992_; 
wire u0__abc_76628_new_n4993_; 
wire u0__abc_76628_new_n4994_; 
wire u0__abc_76628_new_n4995_; 
wire u0__abc_76628_new_n4996_; 
wire u0__abc_76628_new_n4997_; 
wire u0__abc_76628_new_n4998_; 
wire u0__abc_76628_new_n4999_; 
wire u0__abc_76628_new_n5000_; 
wire u0__abc_76628_new_n5001_; 
wire u0__abc_76628_new_n5002_; 
wire u0__abc_76628_new_n5003_; 
wire u0__abc_76628_new_n5004_; 
wire u0__abc_76628_new_n5005_; 
wire u0__abc_76628_new_n5006_; 
wire u0__abc_76628_new_n5007_; 
wire u0__abc_76628_new_n5009_; 
wire u0__abc_76628_new_n5010_; 
wire u0__abc_76628_new_n5011_; 
wire u0__abc_76628_new_n5012_; 
wire u0__abc_76628_new_n5013_; 
wire u0__abc_76628_new_n5014_; 
wire u0__abc_76628_new_n5015_; 
wire u0__abc_76628_new_n5016_; 
wire u0__abc_76628_new_n5017_; 
wire u0__abc_76628_new_n5018_; 
wire u0__abc_76628_new_n5019_; 
wire u0__abc_76628_new_n5020_; 
wire u0__abc_76628_new_n5021_; 
wire u0__abc_76628_new_n5022_; 
wire u0__abc_76628_new_n5023_; 
wire u0__abc_76628_new_n5024_; 
wire u0__abc_76628_new_n5025_; 
wire u0__abc_76628_new_n5026_; 
wire u0__abc_76628_new_n5027_; 
wire u0__abc_76628_new_n5028_; 
wire u0__abc_76628_new_n5029_; 
wire u0__abc_76628_new_n5030_; 
wire u0__abc_76628_new_n5031_; 
wire u0__abc_76628_new_n5032_; 
wire u0__abc_76628_new_n5033_; 
wire u0__abc_76628_new_n5034_; 
wire u0__abc_76628_new_n5035_; 
wire u0__abc_76628_new_n5036_; 
wire u0__abc_76628_new_n5037_; 
wire u0__abc_76628_new_n5038_; 
wire u0__abc_76628_new_n5039_; 
wire u0__abc_76628_new_n5040_; 
wire u0__abc_76628_new_n5042_; 
wire u0__abc_76628_new_n5043_; 
wire u0__abc_76628_new_n5044_; 
wire u0__abc_76628_new_n5045_; 
wire u0__abc_76628_new_n5046_; 
wire u0__abc_76628_new_n5047_; 
wire u0__abc_76628_new_n5048_; 
wire u0__abc_76628_new_n5049_; 
wire u0__abc_76628_new_n5050_; 
wire u0__abc_76628_new_n5051_; 
wire u0__abc_76628_new_n5052_; 
wire u0__abc_76628_new_n5053_; 
wire u0__abc_76628_new_n5054_; 
wire u0__abc_76628_new_n5055_; 
wire u0__abc_76628_new_n5056_; 
wire u0__abc_76628_new_n5057_; 
wire u0__abc_76628_new_n5058_; 
wire u0__abc_76628_new_n5059_; 
wire u0__abc_76628_new_n5060_; 
wire u0__abc_76628_new_n5061_; 
wire u0__abc_76628_new_n5062_; 
wire u0__abc_76628_new_n5063_; 
wire u0__abc_76628_new_n5064_; 
wire u0__abc_76628_new_n5065_; 
wire u0__abc_76628_new_n5066_; 
wire u0__abc_76628_new_n5067_; 
wire u0__abc_76628_new_n5068_; 
wire u0__abc_76628_new_n5069_; 
wire u0__abc_76628_new_n5070_; 
wire u0__abc_76628_new_n5071_; 
wire u0__abc_76628_new_n5072_; 
wire u0__abc_76628_new_n5073_; 
wire u0__abc_76628_new_n5075_; 
wire u0__abc_76628_new_n5076_; 
wire u0__abc_76628_new_n5077_; 
wire u0__abc_76628_new_n5078_; 
wire u0__abc_76628_new_n5079_; 
wire u0__abc_76628_new_n5080_; 
wire u0__abc_76628_new_n5081_; 
wire u0__abc_76628_new_n5082_; 
wire u0__abc_76628_new_n5083_; 
wire u0__abc_76628_new_n5084_; 
wire u0__abc_76628_new_n5085_; 
wire u0__abc_76628_new_n5086_; 
wire u0__abc_76628_new_n5087_; 
wire u0__abc_76628_new_n5088_; 
wire u0__abc_76628_new_n5089_; 
wire u0__abc_76628_new_n5090_; 
wire u0__abc_76628_new_n5091_; 
wire u0__abc_76628_new_n5092_; 
wire u0__abc_76628_new_n5093_; 
wire u0__abc_76628_new_n5094_; 
wire u0__abc_76628_new_n5095_; 
wire u0__abc_76628_new_n5096_; 
wire u0__abc_76628_new_n5097_; 
wire u0__abc_76628_new_n5098_; 
wire u0__abc_76628_new_n5099_; 
wire u0__abc_76628_new_n5100_; 
wire u0__abc_76628_new_n5101_; 
wire u0__abc_76628_new_n5102_; 
wire u0__abc_76628_new_n5103_; 
wire u0__abc_76628_new_n5104_; 
wire u0__abc_76628_new_n5105_; 
wire u0__abc_76628_new_n5106_; 
wire u0__abc_76628_new_n5108_; 
wire u0__abc_76628_new_n5109_; 
wire u0__abc_76628_new_n5110_; 
wire u0__abc_76628_new_n5111_; 
wire u0__abc_76628_new_n5112_; 
wire u0__abc_76628_new_n5113_; 
wire u0__abc_76628_new_n5114_; 
wire u0__abc_76628_new_n5115_; 
wire u0__abc_76628_new_n5116_; 
wire u0__abc_76628_new_n5117_; 
wire u0__abc_76628_new_n5118_; 
wire u0__abc_76628_new_n5119_; 
wire u0__abc_76628_new_n5120_; 
wire u0__abc_76628_new_n5121_; 
wire u0__abc_76628_new_n5122_; 
wire u0__abc_76628_new_n5123_; 
wire u0__abc_76628_new_n5124_; 
wire u0__abc_76628_new_n5125_; 
wire u0__abc_76628_new_n5126_; 
wire u0__abc_76628_new_n5127_; 
wire u0__abc_76628_new_n5128_; 
wire u0__abc_76628_new_n5129_; 
wire u0__abc_76628_new_n5130_; 
wire u0__abc_76628_new_n5131_; 
wire u0__abc_76628_new_n5132_; 
wire u0__abc_76628_new_n5133_; 
wire u0__abc_76628_new_n5134_; 
wire u0__abc_76628_new_n5135_; 
wire u0__abc_76628_new_n5136_; 
wire u0__abc_76628_new_n5137_; 
wire u0__abc_76628_new_n5138_; 
wire u0__abc_76628_new_n5139_; 
wire u0__abc_76628_new_n5141_; 
wire u0__abc_76628_new_n5142_; 
wire u0__abc_76628_new_n5143_; 
wire u0__abc_76628_new_n5144_; 
wire u0__abc_76628_new_n5145_; 
wire u0__abc_76628_new_n5146_; 
wire u0__abc_76628_new_n5147_; 
wire u0__abc_76628_new_n5148_; 
wire u0__abc_76628_new_n5149_; 
wire u0__abc_76628_new_n5150_; 
wire u0__abc_76628_new_n5151_; 
wire u0__abc_76628_new_n5152_; 
wire u0__abc_76628_new_n5153_; 
wire u0__abc_76628_new_n5154_; 
wire u0__abc_76628_new_n5155_; 
wire u0__abc_76628_new_n5156_; 
wire u0__abc_76628_new_n5157_; 
wire u0__abc_76628_new_n5158_; 
wire u0__abc_76628_new_n5159_; 
wire u0__abc_76628_new_n5160_; 
wire u0__abc_76628_new_n5161_; 
wire u0__abc_76628_new_n5162_; 
wire u0__abc_76628_new_n5163_; 
wire u0__abc_76628_new_n5164_; 
wire u0__abc_76628_new_n5165_; 
wire u0__abc_76628_new_n5166_; 
wire u0__abc_76628_new_n5167_; 
wire u0__abc_76628_new_n5168_; 
wire u0__abc_76628_new_n5169_; 
wire u0__abc_76628_new_n5170_; 
wire u0__abc_76628_new_n5171_; 
wire u0__abc_76628_new_n5172_; 
wire u0__abc_76628_new_n5174_; 
wire u0__abc_76628_new_n5175_; 
wire u0__abc_76628_new_n5176_; 
wire u0__abc_76628_new_n5177_; 
wire u0__abc_76628_new_n5178_; 
wire u0__abc_76628_new_n5179_; 
wire u0__abc_76628_new_n5180_; 
wire u0__abc_76628_new_n5181_; 
wire u0__abc_76628_new_n5182_; 
wire u0__abc_76628_new_n5183_; 
wire u0__abc_76628_new_n5184_; 
wire u0__abc_76628_new_n5185_; 
wire u0__abc_76628_new_n5186_; 
wire u0__abc_76628_new_n5187_; 
wire u0__abc_76628_new_n5188_; 
wire u0__abc_76628_new_n5189_; 
wire u0__abc_76628_new_n5190_; 
wire u0__abc_76628_new_n5191_; 
wire u0__abc_76628_new_n5192_; 
wire u0__abc_76628_new_n5193_; 
wire u0__abc_76628_new_n5194_; 
wire u0__abc_76628_new_n5195_; 
wire u0__abc_76628_new_n5196_; 
wire u0__abc_76628_new_n5197_; 
wire u0__abc_76628_new_n5198_; 
wire u0__abc_76628_new_n5199_; 
wire u0__abc_76628_new_n5200_; 
wire u0__abc_76628_new_n5201_; 
wire u0__abc_76628_new_n5202_; 
wire u0__abc_76628_new_n5203_; 
wire u0__abc_76628_new_n5204_; 
wire u0__abc_76628_new_n5205_; 
wire u0__abc_76628_new_n5207_; 
wire u0__abc_76628_new_n5208_; 
wire u0__abc_76628_new_n5209_; 
wire u0__abc_76628_new_n5210_; 
wire u0__abc_76628_new_n5211_; 
wire u0__abc_76628_new_n5212_; 
wire u0__abc_76628_new_n5213_; 
wire u0__abc_76628_new_n5214_; 
wire u0__abc_76628_new_n5215_; 
wire u0__abc_76628_new_n5216_; 
wire u0__abc_76628_new_n5217_; 
wire u0__abc_76628_new_n5218_; 
wire u0__abc_76628_new_n5219_; 
wire u0__abc_76628_new_n5220_; 
wire u0__abc_76628_new_n5221_; 
wire u0__abc_76628_new_n5222_; 
wire u0__abc_76628_new_n5223_; 
wire u0__abc_76628_new_n5224_; 
wire u0__abc_76628_new_n5225_; 
wire u0__abc_76628_new_n5226_; 
wire u0__abc_76628_new_n5227_; 
wire u0__abc_76628_new_n5228_; 
wire u0__abc_76628_new_n5229_; 
wire u0__abc_76628_new_n5230_; 
wire u0__abc_76628_new_n5231_; 
wire u0__abc_76628_new_n5232_; 
wire u0__abc_76628_new_n5233_; 
wire u0__abc_76628_new_n5234_; 
wire u0__abc_76628_new_n5235_; 
wire u0__abc_76628_new_n5236_; 
wire u0__abc_76628_new_n5237_; 
wire u0__abc_76628_new_n5238_; 
wire u0__abc_76628_new_n5240_; 
wire u0__abc_76628_new_n5241_; 
wire u0__abc_76628_new_n5242_; 
wire u0__abc_76628_new_n5243_; 
wire u0__abc_76628_new_n5244_; 
wire u0__abc_76628_new_n5245_; 
wire u0__abc_76628_new_n5246_; 
wire u0__abc_76628_new_n5247_; 
wire u0__abc_76628_new_n5248_; 
wire u0__abc_76628_new_n5249_; 
wire u0__abc_76628_new_n5250_; 
wire u0__abc_76628_new_n5251_; 
wire u0__abc_76628_new_n5252_; 
wire u0__abc_76628_new_n5253_; 
wire u0__abc_76628_new_n5254_; 
wire u0__abc_76628_new_n5255_; 
wire u0__abc_76628_new_n5256_; 
wire u0__abc_76628_new_n5257_; 
wire u0__abc_76628_new_n5258_; 
wire u0__abc_76628_new_n5259_; 
wire u0__abc_76628_new_n5260_; 
wire u0__abc_76628_new_n5261_; 
wire u0__abc_76628_new_n5262_; 
wire u0__abc_76628_new_n5263_; 
wire u0__abc_76628_new_n5264_; 
wire u0__abc_76628_new_n5265_; 
wire u0__abc_76628_new_n5266_; 
wire u0__abc_76628_new_n5267_; 
wire u0__abc_76628_new_n5268_; 
wire u0__abc_76628_new_n5269_; 
wire u0__abc_76628_new_n5270_; 
wire u0__abc_76628_new_n5271_; 
wire u0__abc_76628_new_n5273_; 
wire u0__abc_76628_new_n5274_; 
wire u0__abc_76628_new_n5275_; 
wire u0__abc_76628_new_n5276_; 
wire u0__abc_76628_new_n5277_; 
wire u0__abc_76628_new_n5278_; 
wire u0__abc_76628_new_n5279_; 
wire u0__abc_76628_new_n5280_; 
wire u0__abc_76628_new_n5281_; 
wire u0__abc_76628_new_n5282_; 
wire u0__abc_76628_new_n5283_; 
wire u0__abc_76628_new_n5284_; 
wire u0__abc_76628_new_n5285_; 
wire u0__abc_76628_new_n5286_; 
wire u0__abc_76628_new_n5287_; 
wire u0__abc_76628_new_n5288_; 
wire u0__abc_76628_new_n5289_; 
wire u0__abc_76628_new_n5290_; 
wire u0__abc_76628_new_n5291_; 
wire u0__abc_76628_new_n5292_; 
wire u0__abc_76628_new_n5293_; 
wire u0__abc_76628_new_n5294_; 
wire u0__abc_76628_new_n5295_; 
wire u0__abc_76628_new_n5296_; 
wire u0__abc_76628_new_n5297_; 
wire u0__abc_76628_new_n5298_; 
wire u0__abc_76628_new_n5299_; 
wire u0__abc_76628_new_n5300_; 
wire u0__abc_76628_new_n5301_; 
wire u0__abc_76628_new_n5302_; 
wire u0__abc_76628_new_n5303_; 
wire u0__abc_76628_new_n5304_; 
wire u0__abc_76628_new_n5306_; 
wire u0__abc_76628_new_n5307_; 
wire u0__abc_76628_new_n5308_; 
wire u0__abc_76628_new_n5309_; 
wire u0__abc_76628_new_n5310_; 
wire u0__abc_76628_new_n5311_; 
wire u0__abc_76628_new_n5312_; 
wire u0__abc_76628_new_n5313_; 
wire u0__abc_76628_new_n5314_; 
wire u0__abc_76628_new_n5315_; 
wire u0__abc_76628_new_n5316_; 
wire u0__abc_76628_new_n5317_; 
wire u0__abc_76628_new_n5318_; 
wire u0__abc_76628_new_n5319_; 
wire u0__abc_76628_new_n5320_; 
wire u0__abc_76628_new_n5321_; 
wire u0__abc_76628_new_n5322_; 
wire u0__abc_76628_new_n5323_; 
wire u0__abc_76628_new_n5324_; 
wire u0__abc_76628_new_n5325_; 
wire u0__abc_76628_new_n5326_; 
wire u0__abc_76628_new_n5327_; 
wire u0__abc_76628_new_n5328_; 
wire u0__abc_76628_new_n5329_; 
wire u0__abc_76628_new_n5330_; 
wire u0__abc_76628_new_n5331_; 
wire u0__abc_76628_new_n5332_; 
wire u0__abc_76628_new_n5333_; 
wire u0__abc_76628_new_n5334_; 
wire u0__abc_76628_new_n5335_; 
wire u0__abc_76628_new_n5336_; 
wire u0__abc_76628_new_n5337_; 
wire u0__abc_76628_new_n5339_; 
wire u0__abc_76628_new_n5340_; 
wire u0__abc_76628_new_n5341_; 
wire u0__abc_76628_new_n5342_; 
wire u0__abc_76628_new_n5343_; 
wire u0__abc_76628_new_n5344_; 
wire u0__abc_76628_new_n5345_; 
wire u0__abc_76628_new_n5346_; 
wire u0__abc_76628_new_n5347_; 
wire u0__abc_76628_new_n5348_; 
wire u0__abc_76628_new_n5349_; 
wire u0__abc_76628_new_n5350_; 
wire u0__abc_76628_new_n5351_; 
wire u0__abc_76628_new_n5352_; 
wire u0__abc_76628_new_n5353_; 
wire u0__abc_76628_new_n5354_; 
wire u0__abc_76628_new_n5355_; 
wire u0__abc_76628_new_n5356_; 
wire u0__abc_76628_new_n5357_; 
wire u0__abc_76628_new_n5358_; 
wire u0__abc_76628_new_n5359_; 
wire u0__abc_76628_new_n5360_; 
wire u0__abc_76628_new_n5361_; 
wire u0__abc_76628_new_n5362_; 
wire u0__abc_76628_new_n5363_; 
wire u0__abc_76628_new_n5364_; 
wire u0__abc_76628_new_n5365_; 
wire u0__abc_76628_new_n5366_; 
wire u0__abc_76628_new_n5367_; 
wire u0__abc_76628_new_n5368_; 
wire u0__abc_76628_new_n5369_; 
wire u0__abc_76628_new_n5370_; 
wire u0__abc_76628_new_n5372_; 
wire u0__abc_76628_new_n5373_; 
wire u0__abc_76628_new_n5374_; 
wire u0__abc_76628_new_n5375_; 
wire u0__abc_76628_new_n5376_; 
wire u0__abc_76628_new_n5377_; 
wire u0__abc_76628_new_n5378_; 
wire u0__abc_76628_new_n5379_; 
wire u0__abc_76628_new_n5380_; 
wire u0__abc_76628_new_n5381_; 
wire u0__abc_76628_new_n5382_; 
wire u0__abc_76628_new_n5383_; 
wire u0__abc_76628_new_n5384_; 
wire u0__abc_76628_new_n5385_; 
wire u0__abc_76628_new_n5386_; 
wire u0__abc_76628_new_n5387_; 
wire u0__abc_76628_new_n5388_; 
wire u0__abc_76628_new_n5389_; 
wire u0__abc_76628_new_n5390_; 
wire u0__abc_76628_new_n5391_; 
wire u0__abc_76628_new_n5392_; 
wire u0__abc_76628_new_n5393_; 
wire u0__abc_76628_new_n5394_; 
wire u0__abc_76628_new_n5395_; 
wire u0__abc_76628_new_n5396_; 
wire u0__abc_76628_new_n5397_; 
wire u0__abc_76628_new_n5398_; 
wire u0__abc_76628_new_n5399_; 
wire u0__abc_76628_new_n5400_; 
wire u0__abc_76628_new_n5401_; 
wire u0__abc_76628_new_n5402_; 
wire u0__abc_76628_new_n5403_; 
wire u0__abc_76628_new_n5404_; 
wire u0__abc_76628_new_n5405_; 
wire u0__abc_76628_new_n5407_; 
wire u0__abc_76628_new_n5408_; 
wire u0__abc_76628_new_n5409_; 
wire u0__abc_76628_new_n5410_; 
wire u0__abc_76628_new_n5411_; 
wire u0__abc_76628_new_n5412_; 
wire u0__abc_76628_new_n5413_; 
wire u0__abc_76628_new_n5414_; 
wire u0__abc_76628_new_n5415_; 
wire u0__abc_76628_new_n5416_; 
wire u0__abc_76628_new_n5417_; 
wire u0__abc_76628_new_n5418_; 
wire u0__abc_76628_new_n5419_; 
wire u0__abc_76628_new_n5420_; 
wire u0__abc_76628_new_n5421_; 
wire u0__abc_76628_new_n5422_; 
wire u0__abc_76628_new_n5423_; 
wire u0__abc_76628_new_n5424_; 
wire u0__abc_76628_new_n5425_; 
wire u0__abc_76628_new_n5426_; 
wire u0__abc_76628_new_n5427_; 
wire u0__abc_76628_new_n5428_; 
wire u0__abc_76628_new_n5429_; 
wire u0__abc_76628_new_n5430_; 
wire u0__abc_76628_new_n5431_; 
wire u0__abc_76628_new_n5432_; 
wire u0__abc_76628_new_n5433_; 
wire u0__abc_76628_new_n5434_; 
wire u0__abc_76628_new_n5435_; 
wire u0__abc_76628_new_n5436_; 
wire u0__abc_76628_new_n5437_; 
wire u0__abc_76628_new_n5438_; 
wire u0__abc_76628_new_n5439_; 
wire u0__abc_76628_new_n5440_; 
wire u0__abc_76628_new_n5442_; 
wire u0__abc_76628_new_n5443_; 
wire u0__abc_76628_new_n5444_; 
wire u0__abc_76628_new_n5445_; 
wire u0__abc_76628_new_n5446_; 
wire u0__abc_76628_new_n5447_; 
wire u0__abc_76628_new_n5448_; 
wire u0__abc_76628_new_n5449_; 
wire u0__abc_76628_new_n5450_; 
wire u0__abc_76628_new_n5451_; 
wire u0__abc_76628_new_n5452_; 
wire u0__abc_76628_new_n5453_; 
wire u0__abc_76628_new_n5454_; 
wire u0__abc_76628_new_n5455_; 
wire u0__abc_76628_new_n5456_; 
wire u0__abc_76628_new_n5457_; 
wire u0__abc_76628_new_n5458_; 
wire u0__abc_76628_new_n5459_; 
wire u0__abc_76628_new_n5460_; 
wire u0__abc_76628_new_n5461_; 
wire u0__abc_76628_new_n5462_; 
wire u0__abc_76628_new_n5463_; 
wire u0__abc_76628_new_n5464_; 
wire u0__abc_76628_new_n5465_; 
wire u0__abc_76628_new_n5466_; 
wire u0__abc_76628_new_n5467_; 
wire u0__abc_76628_new_n5468_; 
wire u0__abc_76628_new_n5469_; 
wire u0__abc_76628_new_n5470_; 
wire u0__abc_76628_new_n5471_; 
wire u0__abc_76628_new_n5472_; 
wire u0__abc_76628_new_n5473_; 
wire u0__abc_76628_new_n5474_; 
wire u0__abc_76628_new_n5475_; 
wire u0__abc_76628_new_n5477_; 
wire u0__abc_76628_new_n5478_; 
wire u0__abc_76628_new_n5479_; 
wire u0__abc_76628_new_n5480_; 
wire u0__abc_76628_new_n5481_; 
wire u0__abc_76628_new_n5482_; 
wire u0__abc_76628_new_n5483_; 
wire u0__abc_76628_new_n5484_; 
wire u0__abc_76628_new_n5485_; 
wire u0__abc_76628_new_n5486_; 
wire u0__abc_76628_new_n5487_; 
wire u0__abc_76628_new_n5488_; 
wire u0__abc_76628_new_n5489_; 
wire u0__abc_76628_new_n5490_; 
wire u0__abc_76628_new_n5491_; 
wire u0__abc_76628_new_n5492_; 
wire u0__abc_76628_new_n5493_; 
wire u0__abc_76628_new_n5494_; 
wire u0__abc_76628_new_n5495_; 
wire u0__abc_76628_new_n5496_; 
wire u0__abc_76628_new_n5497_; 
wire u0__abc_76628_new_n5498_; 
wire u0__abc_76628_new_n5499_; 
wire u0__abc_76628_new_n5500_; 
wire u0__abc_76628_new_n5501_; 
wire u0__abc_76628_new_n5502_; 
wire u0__abc_76628_new_n5503_; 
wire u0__abc_76628_new_n5504_; 
wire u0__abc_76628_new_n5505_; 
wire u0__abc_76628_new_n5506_; 
wire u0__abc_76628_new_n5507_; 
wire u0__abc_76628_new_n5508_; 
wire u0__abc_76628_new_n5509_; 
wire u0__abc_76628_new_n5510_; 
wire u0__abc_76628_new_n5512_; 
wire u0__abc_76628_new_n5513_; 
wire u0__abc_76628_new_n5514_; 
wire u0__abc_76628_new_n5515_; 
wire u0__abc_76628_new_n5516_; 
wire u0__abc_76628_new_n5517_; 
wire u0__abc_76628_new_n5518_; 
wire u0__abc_76628_new_n5519_; 
wire u0__abc_76628_new_n5520_; 
wire u0__abc_76628_new_n5521_; 
wire u0__abc_76628_new_n5522_; 
wire u0__abc_76628_new_n5523_; 
wire u0__abc_76628_new_n5524_; 
wire u0__abc_76628_new_n5525_; 
wire u0__abc_76628_new_n5526_; 
wire u0__abc_76628_new_n5527_; 
wire u0__abc_76628_new_n5528_; 
wire u0__abc_76628_new_n5529_; 
wire u0__abc_76628_new_n5530_; 
wire u0__abc_76628_new_n5531_; 
wire u0__abc_76628_new_n5532_; 
wire u0__abc_76628_new_n5533_; 
wire u0__abc_76628_new_n5534_; 
wire u0__abc_76628_new_n5535_; 
wire u0__abc_76628_new_n5536_; 
wire u0__abc_76628_new_n5537_; 
wire u0__abc_76628_new_n5538_; 
wire u0__abc_76628_new_n5539_; 
wire u0__abc_76628_new_n5540_; 
wire u0__abc_76628_new_n5541_; 
wire u0__abc_76628_new_n5542_; 
wire u0__abc_76628_new_n5543_; 
wire u0__abc_76628_new_n5544_; 
wire u0__abc_76628_new_n5545_; 
wire u0__abc_76628_new_n5547_; 
wire u0__abc_76628_new_n5548_; 
wire u0__abc_76628_new_n5549_; 
wire u0__abc_76628_new_n5550_; 
wire u0__abc_76628_new_n5551_; 
wire u0__abc_76628_new_n5552_; 
wire u0__abc_76628_new_n5553_; 
wire u0__abc_76628_new_n5554_; 
wire u0__abc_76628_new_n5555_; 
wire u0__abc_76628_new_n5556_; 
wire u0__abc_76628_new_n5557_; 
wire u0__abc_76628_new_n5558_; 
wire u0__abc_76628_new_n5559_; 
wire u0__abc_76628_new_n5560_; 
wire u0__abc_76628_new_n5561_; 
wire u0__abc_76628_new_n5562_; 
wire u0__abc_76628_new_n5563_; 
wire u0__abc_76628_new_n5564_; 
wire u0__abc_76628_new_n5565_; 
wire u0__abc_76628_new_n5566_; 
wire u0__abc_76628_new_n5567_; 
wire u0__abc_76628_new_n5568_; 
wire u0__abc_76628_new_n5569_; 
wire u0__abc_76628_new_n5570_; 
wire u0__abc_76628_new_n5571_; 
wire u0__abc_76628_new_n5572_; 
wire u0__abc_76628_new_n5573_; 
wire u0__abc_76628_new_n5574_; 
wire u0__abc_76628_new_n5575_; 
wire u0__abc_76628_new_n5576_; 
wire u0__abc_76628_new_n5577_; 
wire u0__abc_76628_new_n5578_; 
wire u0__abc_76628_new_n5579_; 
wire u0__abc_76628_new_n5580_; 
wire u0__abc_76628_new_n5582_; 
wire u0__abc_76628_new_n5583_; 
wire u0__abc_76628_new_n5584_; 
wire u0__abc_76628_new_n5585_; 
wire u0__abc_76628_new_n5586_; 
wire u0__abc_76628_new_n5587_; 
wire u0__abc_76628_new_n5588_; 
wire u0__abc_76628_new_n5589_; 
wire u0__abc_76628_new_n5590_; 
wire u0__abc_76628_new_n5591_; 
wire u0__abc_76628_new_n5592_; 
wire u0__abc_76628_new_n5593_; 
wire u0__abc_76628_new_n5594_; 
wire u0__abc_76628_new_n5595_; 
wire u0__abc_76628_new_n5596_; 
wire u0__abc_76628_new_n5597_; 
wire u0__abc_76628_new_n5598_; 
wire u0__abc_76628_new_n5599_; 
wire u0__abc_76628_new_n5600_; 
wire u0__abc_76628_new_n5601_; 
wire u0__abc_76628_new_n5602_; 
wire u0__abc_76628_new_n5603_; 
wire u0__abc_76628_new_n5604_; 
wire u0__abc_76628_new_n5605_; 
wire u0__abc_76628_new_n5606_; 
wire u0__abc_76628_new_n5607_; 
wire u0__abc_76628_new_n5608_; 
wire u0__abc_76628_new_n5609_; 
wire u0__abc_76628_new_n5610_; 
wire u0__abc_76628_new_n5611_; 
wire u0__abc_76628_new_n5612_; 
wire u0__abc_76628_new_n5613_; 
wire u0__abc_76628_new_n5614_; 
wire u0__abc_76628_new_n5615_; 
wire u0__abc_76628_new_n5617_; 
wire u0__abc_76628_new_n5618_; 
wire u0__abc_76628_new_n5619_; 
wire u0__abc_76628_new_n5620_; 
wire u0__abc_76628_new_n5621_; 
wire u0__abc_76628_new_n5622_; 
wire u0__abc_76628_new_n5623_; 
wire u0__abc_76628_new_n5624_; 
wire u0__abc_76628_new_n5625_; 
wire u0__abc_76628_new_n5626_; 
wire u0__abc_76628_new_n5627_; 
wire u0__abc_76628_new_n5628_; 
wire u0__abc_76628_new_n5629_; 
wire u0__abc_76628_new_n5630_; 
wire u0__abc_76628_new_n5631_; 
wire u0__abc_76628_new_n5632_; 
wire u0__abc_76628_new_n5633_; 
wire u0__abc_76628_new_n5634_; 
wire u0__abc_76628_new_n5635_; 
wire u0__abc_76628_new_n5636_; 
wire u0__abc_76628_new_n5637_; 
wire u0__abc_76628_new_n5638_; 
wire u0__abc_76628_new_n5639_; 
wire u0__abc_76628_new_n5640_; 
wire u0__abc_76628_new_n5641_; 
wire u0__abc_76628_new_n5642_; 
wire u0__abc_76628_new_n5643_; 
wire u0__abc_76628_new_n5644_; 
wire u0__abc_76628_new_n5645_; 
wire u0__abc_76628_new_n5646_; 
wire u0__abc_76628_new_n5647_; 
wire u0__abc_76628_new_n5648_; 
wire u0__abc_76628_new_n5649_; 
wire u0__abc_76628_new_n5650_; 
wire u0__abc_76628_new_n5652_; 
wire u0__abc_76628_new_n5653_; 
wire u0__abc_76628_new_n5654_; 
wire u0__abc_76628_new_n5655_; 
wire u0__abc_76628_new_n5656_; 
wire u0__abc_76628_new_n5660_; 
wire u0__abc_76628_new_n5661_; 
wire u0__abc_76628_new_n5662_; 
wire u0__abc_76628_new_n5663_; 
wire u0__abc_76628_new_n5664_; 
wire u0__abc_76628_new_n5666_; 
wire u0__abc_76628_new_n5667_; 
wire u0__abc_76628_new_n5668_; 
wire u0__abc_76628_new_n5669_; 
wire u0__abc_76628_new_n5670_; 
wire u0__abc_76628_new_n5672_; 
wire u0__abc_76628_new_n5673_; 
wire u0__abc_76628_new_n5674_; 
wire u0__abc_76628_new_n5675_; 
wire u0__abc_76628_new_n5676_; 
wire u0__abc_76628_new_n5678_; 
wire u0__abc_76628_new_n5679_; 
wire u0__abc_76628_new_n5680_; 
wire u0__abc_76628_new_n5681_; 
wire u0__abc_76628_new_n5682_; 
wire u0__abc_76628_new_n5684_; 
wire u0__abc_76628_new_n5685_; 
wire u0__abc_76628_new_n5686_; 
wire u0__abc_76628_new_n5687_; 
wire u0__abc_76628_new_n5688_; 
wire u0__abc_76628_new_n5690_; 
wire u0__abc_76628_new_n5691_; 
wire u0__abc_76628_new_n5692_; 
wire u0__abc_76628_new_n5693_; 
wire u0__abc_76628_new_n5694_; 
wire u0__abc_76628_new_n5696_; 
wire u0__abc_76628_new_n5697_; 
wire u0__abc_76628_new_n5698_; 
wire u0__abc_76628_new_n5699_; 
wire u0__abc_76628_new_n5700_; 
wire u0__abc_76628_new_n5702_; 
wire u0__abc_76628_new_n5703_; 
wire u0__abc_76628_new_n5704_; 
wire u0__abc_76628_new_n5705_; 
wire u0__abc_76628_new_n5706_; 
wire u0__abc_76628_new_n5708_; 
wire u0__abc_76628_new_n5709_; 
wire u0__abc_76628_new_n5710_; 
wire u0__abc_76628_new_n5711_; 
wire u0__abc_76628_new_n5712_; 
wire u0__abc_76628_new_n5713_; 
wire u0__abc_76628_new_n5714_; 
wire u0__abc_76628_new_n5716_; 
wire u0__abc_76628_new_n5717_; 
wire u0__abc_76628_new_n5718_; 
wire u0__abc_76628_new_n5719_; 
wire u0__abc_76628_new_n5720_; 
wire u0__abc_76628_new_n5721_; 
wire u0__abc_76628_new_n5723_; 
wire u0__abc_76628_new_n5724_; 
wire u0__abc_76628_new_n5725_; 
wire u0__abc_76628_new_n5726_; 
wire u0__abc_76628_new_n5727_; 
wire u0__abc_76628_new_n5728_; 
wire u0_cs0; 
wire u0_cs0_bF_buf0; 
wire u0_cs0_bF_buf1; 
wire u0_cs0_bF_buf2; 
wire u0_cs0_bF_buf3; 
wire u0_cs0_bF_buf4; 
wire u0_cs0_bF_buf5; 
wire u0_cs1; 
wire u0_cs1_bF_buf0; 
wire u0_cs1_bF_buf1; 
wire u0_cs1_bF_buf2; 
wire u0_cs1_bF_buf3; 
wire u0_cs1_bF_buf4; 
wire u0_cs1_bF_buf5; 
wire u0_csc0_0_; 
wire u0_csc0_10_; 
wire u0_csc0_11_; 
wire u0_csc0_12_; 
wire u0_csc0_13_; 
wire u0_csc0_14_; 
wire u0_csc0_15_; 
wire u0_csc0_16_; 
wire u0_csc0_17_; 
wire u0_csc0_18_; 
wire u0_csc0_19_; 
wire u0_csc0_1_; 
wire u0_csc0_20_; 
wire u0_csc0_21_; 
wire u0_csc0_22_; 
wire u0_csc0_23_; 
wire u0_csc0_24_; 
wire u0_csc0_25_; 
wire u0_csc0_26_; 
wire u0_csc0_27_; 
wire u0_csc0_28_; 
wire u0_csc0_29_; 
wire u0_csc0_2_; 
wire u0_csc0_30_; 
wire u0_csc0_31_; 
wire u0_csc0_3_; 
wire u0_csc0_4_; 
wire u0_csc0_5_; 
wire u0_csc0_6_; 
wire u0_csc0_7_; 
wire u0_csc0_8_; 
wire u0_csc0_9_; 
wire u0_csc1_0_; 
wire u0_csc1_10_; 
wire u0_csc1_11_; 
wire u0_csc1_12_; 
wire u0_csc1_13_; 
wire u0_csc1_14_; 
wire u0_csc1_15_; 
wire u0_csc1_16_; 
wire u0_csc1_17_; 
wire u0_csc1_18_; 
wire u0_csc1_19_; 
wire u0_csc1_1_; 
wire u0_csc1_20_; 
wire u0_csc1_21_; 
wire u0_csc1_22_; 
wire u0_csc1_23_; 
wire u0_csc1_24_; 
wire u0_csc1_25_; 
wire u0_csc1_26_; 
wire u0_csc1_27_; 
wire u0_csc1_28_; 
wire u0_csc1_29_; 
wire u0_csc1_2_; 
wire u0_csc1_30_; 
wire u0_csc1_31_; 
wire u0_csc1_3_; 
wire u0_csc1_4_; 
wire u0_csc1_5_; 
wire u0_csc1_6_; 
wire u0_csc1_7_; 
wire u0_csc1_8_; 
wire u0_csc1_9_; 
wire u0_csc_mask_0_; 
wire u0_csc_mask_10_; 
wire u0_csc_mask_1_; 
wire u0_csc_mask_2_; 
wire u0_csc_mask_3_; 
wire u0_csc_mask_4_; 
wire u0_csc_mask_5_; 
wire u0_csc_mask_6_; 
wire u0_csc_mask_7_; 
wire u0_csc_mask_8_; 
wire u0_csc_mask_9_; 
wire u0_csr_0_; 
wire u0_csr_1_; 
wire u0_csr_3_; 
wire u0_csr_4_; 
wire u0_csr_5_; 
wire u0_csr_6_; 
wire u0_csr_7_; 
wire u0_init_ack0; 
wire u0_init_ack1; 
wire u0_init_ack_r; 
wire u0_init_req0; 
wire u0_init_req1; 
wire u0_lmr_ack0; 
wire u0_lmr_ack1; 
wire u0_lmr_ack_r; 
wire u0_lmr_req0; 
wire u0_lmr_req1; 
wire u0_rf_we; 
wire u0_rst_r2; 
wire u0_rst_r3; 
wire u0_rst_r3_bF_buf0; 
wire u0_rst_r3_bF_buf1; 
wire u0_rst_r3_bF_buf2; 
wire u0_rst_r3_bF_buf3; 
wire u0_rst_r3_bF_buf4; 
wire u0_sreq_cs_le; 
wire u0_tms0_0_; 
wire u0_tms0_10_; 
wire u0_tms0_11_; 
wire u0_tms0_12_; 
wire u0_tms0_13_; 
wire u0_tms0_14_; 
wire u0_tms0_15_; 
wire u0_tms0_16_; 
wire u0_tms0_17_; 
wire u0_tms0_18_; 
wire u0_tms0_19_; 
wire u0_tms0_1_; 
wire u0_tms0_20_; 
wire u0_tms0_21_; 
wire u0_tms0_22_; 
wire u0_tms0_23_; 
wire u0_tms0_24_; 
wire u0_tms0_25_; 
wire u0_tms0_26_; 
wire u0_tms0_27_; 
wire u0_tms0_28_; 
wire u0_tms0_29_; 
wire u0_tms0_2_; 
wire u0_tms0_30_; 
wire u0_tms0_31_; 
wire u0_tms0_3_; 
wire u0_tms0_4_; 
wire u0_tms0_5_; 
wire u0_tms0_6_; 
wire u0_tms0_7_; 
wire u0_tms0_8_; 
wire u0_tms0_9_; 
wire u0_tms1_0_; 
wire u0_tms1_10_; 
wire u0_tms1_11_; 
wire u0_tms1_12_; 
wire u0_tms1_13_; 
wire u0_tms1_14_; 
wire u0_tms1_15_; 
wire u0_tms1_16_; 
wire u0_tms1_17_; 
wire u0_tms1_18_; 
wire u0_tms1_19_; 
wire u0_tms1_1_; 
wire u0_tms1_20_; 
wire u0_tms1_21_; 
wire u0_tms1_22_; 
wire u0_tms1_23_; 
wire u0_tms1_24_; 
wire u0_tms1_25_; 
wire u0_tms1_26_; 
wire u0_tms1_27_; 
wire u0_tms1_28_; 
wire u0_tms1_29_; 
wire u0_tms1_2_; 
wire u0_tms1_30_; 
wire u0_tms1_31_; 
wire u0_tms1_3_; 
wire u0_tms1_4_; 
wire u0_tms1_5_; 
wire u0_tms1_6_; 
wire u0_tms1_7_; 
wire u0_tms1_8_; 
wire u0_tms1_9_; 
wire u0_u0__0csc_31_0__0_; 
wire u0_u0__0csc_31_0__10_; 
wire u0_u0__0csc_31_0__11_; 
wire u0_u0__0csc_31_0__12_; 
wire u0_u0__0csc_31_0__13_; 
wire u0_u0__0csc_31_0__14_; 
wire u0_u0__0csc_31_0__15_; 
wire u0_u0__0csc_31_0__16_; 
wire u0_u0__0csc_31_0__17_; 
wire u0_u0__0csc_31_0__18_; 
wire u0_u0__0csc_31_0__19_; 
wire u0_u0__0csc_31_0__1_; 
wire u0_u0__0csc_31_0__20_; 
wire u0_u0__0csc_31_0__21_; 
wire u0_u0__0csc_31_0__22_; 
wire u0_u0__0csc_31_0__23_; 
wire u0_u0__0csc_31_0__24_; 
wire u0_u0__0csc_31_0__25_; 
wire u0_u0__0csc_31_0__26_; 
wire u0_u0__0csc_31_0__27_; 
wire u0_u0__0csc_31_0__28_; 
wire u0_u0__0csc_31_0__29_; 
wire u0_u0__0csc_31_0__2_; 
wire u0_u0__0csc_31_0__30_; 
wire u0_u0__0csc_31_0__31_; 
wire u0_u0__0csc_31_0__3_; 
wire u0_u0__0csc_31_0__4_; 
wire u0_u0__0csc_31_0__5_; 
wire u0_u0__0csc_31_0__6_; 
wire u0_u0__0csc_31_0__7_; 
wire u0_u0__0csc_31_0__8_; 
wire u0_u0__0csc_31_0__9_; 
wire u0_u0__0init_req_0_0_; 
wire u0_u0__0init_req_we_0_0_; 
wire u0_u0__0init_req_we_0_0_bF_buf0_; 
wire u0_u0__0init_req_we_0_0_bF_buf1_; 
wire u0_u0__0init_req_we_0_0_bF_buf2_; 
wire u0_u0__0init_req_we_0_0_bF_buf3_; 
wire u0_u0__0init_req_we_0_0_bF_buf4_; 
wire u0_u0__0inited_0_0_; 
wire u0_u0__0lmr_req_0_0_; 
wire u0_u0__0lmr_req_we_0_0_; 
wire u0_u0__0lmr_req_we_0_0_bF_buf0_; 
wire u0_u0__0lmr_req_we_0_0_bF_buf1_; 
wire u0_u0__0lmr_req_we_0_0_bF_buf2_; 
wire u0_u0__0lmr_req_we_0_0_bF_buf3_; 
wire u0_u0__0lmr_req_we_0_0_bF_buf4_; 
wire u0_u0__0tms_31_0__0_; 
wire u0_u0__0tms_31_0__10_; 
wire u0_u0__0tms_31_0__11_; 
wire u0_u0__0tms_31_0__12_; 
wire u0_u0__0tms_31_0__13_; 
wire u0_u0__0tms_31_0__14_; 
wire u0_u0__0tms_31_0__15_; 
wire u0_u0__0tms_31_0__16_; 
wire u0_u0__0tms_31_0__17_; 
wire u0_u0__0tms_31_0__18_; 
wire u0_u0__0tms_31_0__19_; 
wire u0_u0__0tms_31_0__1_; 
wire u0_u0__0tms_31_0__20_; 
wire u0_u0__0tms_31_0__21_; 
wire u0_u0__0tms_31_0__22_; 
wire u0_u0__0tms_31_0__23_; 
wire u0_u0__0tms_31_0__24_; 
wire u0_u0__0tms_31_0__25_; 
wire u0_u0__0tms_31_0__26_; 
wire u0_u0__0tms_31_0__27_; 
wire u0_u0__0tms_31_0__28_; 
wire u0_u0__0tms_31_0__29_; 
wire u0_u0__0tms_31_0__2_; 
wire u0_u0__0tms_31_0__30_; 
wire u0_u0__0tms_31_0__31_; 
wire u0_u0__0tms_31_0__3_; 
wire u0_u0__0tms_31_0__4_; 
wire u0_u0__0tms_31_0__5_; 
wire u0_u0__0tms_31_0__6_; 
wire u0_u0__0tms_31_0__7_; 
wire u0_u0__0tms_31_0__8_; 
wire u0_u0__0tms_31_0__9_; 
wire u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494; 
wire u0_u0__abc_72207_new_n205_; 
wire u0_u0__abc_72207_new_n206_; 
wire u0_u0__abc_72207_new_n207_; 
wire u0_u0__abc_72207_new_n208_; 
wire u0_u0__abc_72207_new_n209_; 
wire u0_u0__abc_72207_new_n210_; 
wire u0_u0__abc_72207_new_n211_; 
wire u0_u0__abc_72207_new_n212_; 
wire u0_u0__abc_72207_new_n213_; 
wire u0_u0__abc_72207_new_n215_; 
wire u0_u0__abc_72207_new_n216_; 
wire u0_u0__abc_72207_new_n217_; 
wire u0_u0__abc_72207_new_n218_; 
wire u0_u0__abc_72207_new_n219_; 
wire u0_u0__abc_72207_new_n220_; 
wire u0_u0__abc_72207_new_n221_; 
wire u0_u0__abc_72207_new_n223_; 
wire u0_u0__abc_72207_new_n224_; 
wire u0_u0__abc_72207_new_n224__bF_buf0; 
wire u0_u0__abc_72207_new_n224__bF_buf1; 
wire u0_u0__abc_72207_new_n224__bF_buf2; 
wire u0_u0__abc_72207_new_n224__bF_buf3; 
wire u0_u0__abc_72207_new_n224__bF_buf4; 
wire u0_u0__abc_72207_new_n225_; 
wire u0_u0__abc_72207_new_n226_; 
wire u0_u0__abc_72207_new_n228_; 
wire u0_u0__abc_72207_new_n229_; 
wire u0_u0__abc_72207_new_n230_; 
wire u0_u0__abc_72207_new_n232_; 
wire u0_u0__abc_72207_new_n233_; 
wire u0_u0__abc_72207_new_n234_; 
wire u0_u0__abc_72207_new_n236_; 
wire u0_u0__abc_72207_new_n237_; 
wire u0_u0__abc_72207_new_n238_; 
wire u0_u0__abc_72207_new_n240_; 
wire u0_u0__abc_72207_new_n241_; 
wire u0_u0__abc_72207_new_n242_; 
wire u0_u0__abc_72207_new_n244_; 
wire u0_u0__abc_72207_new_n245_; 
wire u0_u0__abc_72207_new_n246_; 
wire u0_u0__abc_72207_new_n248_; 
wire u0_u0__abc_72207_new_n249_; 
wire u0_u0__abc_72207_new_n250_; 
wire u0_u0__abc_72207_new_n252_; 
wire u0_u0__abc_72207_new_n253_; 
wire u0_u0__abc_72207_new_n254_; 
wire u0_u0__abc_72207_new_n256_; 
wire u0_u0__abc_72207_new_n257_; 
wire u0_u0__abc_72207_new_n258_; 
wire u0_u0__abc_72207_new_n260_; 
wire u0_u0__abc_72207_new_n261_; 
wire u0_u0__abc_72207_new_n262_; 
wire u0_u0__abc_72207_new_n264_; 
wire u0_u0__abc_72207_new_n265_; 
wire u0_u0__abc_72207_new_n266_; 
wire u0_u0__abc_72207_new_n268_; 
wire u0_u0__abc_72207_new_n269_; 
wire u0_u0__abc_72207_new_n270_; 
wire u0_u0__abc_72207_new_n272_; 
wire u0_u0__abc_72207_new_n273_; 
wire u0_u0__abc_72207_new_n274_; 
wire u0_u0__abc_72207_new_n276_; 
wire u0_u0__abc_72207_new_n277_; 
wire u0_u0__abc_72207_new_n278_; 
wire u0_u0__abc_72207_new_n280_; 
wire u0_u0__abc_72207_new_n281_; 
wire u0_u0__abc_72207_new_n282_; 
wire u0_u0__abc_72207_new_n284_; 
wire u0_u0__abc_72207_new_n285_; 
wire u0_u0__abc_72207_new_n286_; 
wire u0_u0__abc_72207_new_n288_; 
wire u0_u0__abc_72207_new_n289_; 
wire u0_u0__abc_72207_new_n290_; 
wire u0_u0__abc_72207_new_n292_; 
wire u0_u0__abc_72207_new_n293_; 
wire u0_u0__abc_72207_new_n294_; 
wire u0_u0__abc_72207_new_n296_; 
wire u0_u0__abc_72207_new_n297_; 
wire u0_u0__abc_72207_new_n298_; 
wire u0_u0__abc_72207_new_n300_; 
wire u0_u0__abc_72207_new_n301_; 
wire u0_u0__abc_72207_new_n302_; 
wire u0_u0__abc_72207_new_n304_; 
wire u0_u0__abc_72207_new_n305_; 
wire u0_u0__abc_72207_new_n306_; 
wire u0_u0__abc_72207_new_n308_; 
wire u0_u0__abc_72207_new_n309_; 
wire u0_u0__abc_72207_new_n310_; 
wire u0_u0__abc_72207_new_n312_; 
wire u0_u0__abc_72207_new_n313_; 
wire u0_u0__abc_72207_new_n314_; 
wire u0_u0__abc_72207_new_n316_; 
wire u0_u0__abc_72207_new_n317_; 
wire u0_u0__abc_72207_new_n318_; 
wire u0_u0__abc_72207_new_n320_; 
wire u0_u0__abc_72207_new_n321_; 
wire u0_u0__abc_72207_new_n322_; 
wire u0_u0__abc_72207_new_n324_; 
wire u0_u0__abc_72207_new_n325_; 
wire u0_u0__abc_72207_new_n326_; 
wire u0_u0__abc_72207_new_n328_; 
wire u0_u0__abc_72207_new_n329_; 
wire u0_u0__abc_72207_new_n330_; 
wire u0_u0__abc_72207_new_n332_; 
wire u0_u0__abc_72207_new_n333_; 
wire u0_u0__abc_72207_new_n334_; 
wire u0_u0__abc_72207_new_n336_; 
wire u0_u0__abc_72207_new_n337_; 
wire u0_u0__abc_72207_new_n338_; 
wire u0_u0__abc_72207_new_n340_; 
wire u0_u0__abc_72207_new_n341_; 
wire u0_u0__abc_72207_new_n342_; 
wire u0_u0__abc_72207_new_n344_; 
wire u0_u0__abc_72207_new_n345_; 
wire u0_u0__abc_72207_new_n346_; 
wire u0_u0__abc_72207_new_n348_; 
wire u0_u0__abc_72207_new_n349_; 
wire u0_u0__abc_72207_new_n350_; 
wire u0_u0__abc_72207_new_n352_; 
wire u0_u0__abc_72207_new_n354_; 
wire u0_u0__abc_72207_new_n354__bF_buf0; 
wire u0_u0__abc_72207_new_n354__bF_buf1; 
wire u0_u0__abc_72207_new_n354__bF_buf2; 
wire u0_u0__abc_72207_new_n354__bF_buf3; 
wire u0_u0__abc_72207_new_n354__bF_buf4; 
wire u0_u0__abc_72207_new_n355_; 
wire u0_u0__abc_72207_new_n356_; 
wire u0_u0__abc_72207_new_n357_; 
wire u0_u0__abc_72207_new_n358_; 
wire u0_u0__abc_72207_new_n359_; 
wire u0_u0__abc_72207_new_n360_; 
wire u0_u0__abc_72207_new_n361_; 
wire u0_u0__abc_72207_new_n361__bF_buf0; 
wire u0_u0__abc_72207_new_n361__bF_buf1; 
wire u0_u0__abc_72207_new_n361__bF_buf2; 
wire u0_u0__abc_72207_new_n361__bF_buf3; 
wire u0_u0__abc_72207_new_n361__bF_buf4; 
wire u0_u0__abc_72207_new_n362_; 
wire u0_u0__abc_72207_new_n363_; 
wire u0_u0__abc_72207_new_n364_; 
wire u0_u0__abc_72207_new_n365_; 
wire u0_u0__abc_72207_new_n366_; 
wire u0_u0__abc_72207_new_n367_; 
wire u0_u0__abc_72207_new_n369_; 
wire u0_u0__abc_72207_new_n370_; 
wire u0_u0__abc_72207_new_n371_; 
wire u0_u0__abc_72207_new_n372_; 
wire u0_u0__abc_72207_new_n374_; 
wire u0_u0__abc_72207_new_n375_; 
wire u0_u0__abc_72207_new_n376_; 
wire u0_u0__abc_72207_new_n377_; 
wire u0_u0__abc_72207_new_n379_; 
wire u0_u0__abc_72207_new_n380_; 
wire u0_u0__abc_72207_new_n381_; 
wire u0_u0__abc_72207_new_n383_; 
wire u0_u0__abc_72207_new_n384_; 
wire u0_u0__abc_72207_new_n385_; 
wire u0_u0__abc_72207_new_n386_; 
wire u0_u0__abc_72207_new_n387_; 
wire u0_u0__abc_72207_new_n389_; 
wire u0_u0__abc_72207_new_n390_; 
wire u0_u0__abc_72207_new_n391_; 
wire u0_u0__abc_72207_new_n392_; 
wire u0_u0__abc_72207_new_n393_; 
wire u0_u0__abc_72207_new_n395_; 
wire u0_u0__abc_72207_new_n396_; 
wire u0_u0__abc_72207_new_n397_; 
wire u0_u0__abc_72207_new_n399_; 
wire u0_u0__abc_72207_new_n400_; 
wire u0_u0__abc_72207_new_n401_; 
wire u0_u0__abc_72207_new_n403_; 
wire u0_u0__abc_72207_new_n404_; 
wire u0_u0__abc_72207_new_n405_; 
wire u0_u0__abc_72207_new_n407_; 
wire u0_u0__abc_72207_new_n408_; 
wire u0_u0__abc_72207_new_n409_; 
wire u0_u0__abc_72207_new_n411_; 
wire u0_u0__abc_72207_new_n412_; 
wire u0_u0__abc_72207_new_n413_; 
wire u0_u0__abc_72207_new_n415_; 
wire u0_u0__abc_72207_new_n416_; 
wire u0_u0__abc_72207_new_n417_; 
wire u0_u0__abc_72207_new_n419_; 
wire u0_u0__abc_72207_new_n420_; 
wire u0_u0__abc_72207_new_n421_; 
wire u0_u0__abc_72207_new_n423_; 
wire u0_u0__abc_72207_new_n424_; 
wire u0_u0__abc_72207_new_n425_; 
wire u0_u0__abc_72207_new_n427_; 
wire u0_u0__abc_72207_new_n428_; 
wire u0_u0__abc_72207_new_n429_; 
wire u0_u0__abc_72207_new_n431_; 
wire u0_u0__abc_72207_new_n432_; 
wire u0_u0__abc_72207_new_n433_; 
wire u0_u0__abc_72207_new_n435_; 
wire u0_u0__abc_72207_new_n436_; 
wire u0_u0__abc_72207_new_n437_; 
wire u0_u0__abc_72207_new_n439_; 
wire u0_u0__abc_72207_new_n440_; 
wire u0_u0__abc_72207_new_n441_; 
wire u0_u0__abc_72207_new_n443_; 
wire u0_u0__abc_72207_new_n444_; 
wire u0_u0__abc_72207_new_n445_; 
wire u0_u0__abc_72207_new_n447_; 
wire u0_u0__abc_72207_new_n448_; 
wire u0_u0__abc_72207_new_n449_; 
wire u0_u0__abc_72207_new_n451_; 
wire u0_u0__abc_72207_new_n452_; 
wire u0_u0__abc_72207_new_n453_; 
wire u0_u0__abc_72207_new_n455_; 
wire u0_u0__abc_72207_new_n456_; 
wire u0_u0__abc_72207_new_n457_; 
wire u0_u0__abc_72207_new_n459_; 
wire u0_u0__abc_72207_new_n460_; 
wire u0_u0__abc_72207_new_n461_; 
wire u0_u0__abc_72207_new_n463_; 
wire u0_u0__abc_72207_new_n464_; 
wire u0_u0__abc_72207_new_n465_; 
wire u0_u0__abc_72207_new_n467_; 
wire u0_u0__abc_72207_new_n468_; 
wire u0_u0__abc_72207_new_n469_; 
wire u0_u0__abc_72207_new_n471_; 
wire u0_u0__abc_72207_new_n472_; 
wire u0_u0__abc_72207_new_n473_; 
wire u0_u0__abc_72207_new_n475_; 
wire u0_u0__abc_72207_new_n476_; 
wire u0_u0__abc_72207_new_n477_; 
wire u0_u0__abc_72207_new_n479_; 
wire u0_u0__abc_72207_new_n480_; 
wire u0_u0__abc_72207_new_n481_; 
wire u0_u0__abc_72207_new_n483_; 
wire u0_u0__abc_72207_new_n484_; 
wire u0_u0__abc_72207_new_n485_; 
wire u0_u0__abc_72207_new_n487_; 
wire u0_u0__abc_72207_new_n488_; 
wire u0_u0__abc_72207_new_n489_; 
wire u0_u0__abc_72207_new_n491_; 
wire u0_u0__abc_72207_new_n492_; 
wire u0_u0__abc_72207_new_n493_; 
wire u0_u0__abc_72207_new_n495_; 
wire u0_u0__abc_72207_new_n496_; 
wire u0_u0__abc_72207_new_n497_; 
wire u0_u0__abc_72207_new_n499_; 
wire u0_u0__abc_72207_new_n500_; 
wire u0_u0__abc_72207_new_n501_; 
wire u0_u0__abc_72207_new_n502_; 
wire u0_u0__abc_72207_new_n503_; 
wire u0_u0__abc_72207_new_n504_; 
wire u0_u0__abc_72207_new_n505_; 
wire u0_u0__abc_72207_new_n506_; 
wire u0_u0__abc_72207_new_n507_; 
wire u0_u0__abc_72207_new_n508_; 
wire u0_u0__abc_72207_new_n509_; 
wire u0_u0__abc_72207_new_n510_; 
wire u0_u0__abc_72207_new_n511_; 
wire u0_u0__abc_72207_new_n512_; 
wire u0_u0__abc_72207_new_n513_; 
wire u0_u0__abc_72207_new_n514_; 
wire u0_u0__abc_72207_new_n515_; 
wire u0_u0__abc_72207_new_n516_; 
wire u0_u0__abc_72207_new_n517_; 
wire u0_u0__abc_72207_new_n518_; 
wire u0_u0__abc_72207_new_n519_; 
wire u0_u0__abc_72207_new_n520_; 
wire u0_u0__abc_72207_new_n521_; 
wire u0_u0__abc_72207_new_n522_; 
wire u0_u0__abc_72207_new_n523_; 
wire u0_u0__abc_72207_new_n524_; 
wire u0_u0__abc_72207_new_n525_; 
wire u0_u0__abc_72207_new_n526_; 
wire u0_u0__abc_72207_new_n527_; 
wire u0_u0__abc_72207_new_n528_; 
wire u0_u0__abc_72207_new_n529_; 
wire u0_u0__abc_72207_new_n530_; 
wire u0_u0__abc_72207_new_n531_; 
wire u0_u0__abc_72207_new_n532_; 
wire u0_u0__abc_72207_new_n533_; 
wire u0_u0__abc_72207_new_n534_; 
wire u0_u0__abc_72207_new_n535_; 
wire u0_u0__abc_72207_new_n536_; 
wire u0_u0__abc_72207_new_n537_; 
wire u0_u0__abc_72207_new_n538_; 
wire u0_u0__abc_72207_new_n539_; 
wire u0_u0__abc_72207_new_n540_; 
wire u0_u0__abc_72207_new_n541_; 
wire u0_u0__abc_72207_new_n542_; 
wire u0_u0__abc_72207_new_n543_; 
wire u0_u0__abc_72207_new_n544_; 
wire u0_u0__abc_72207_new_n545_; 
wire u0_u0__abc_72207_new_n546_; 
wire u0_u0__abc_72207_new_n547_; 
wire u0_u0__abc_72207_new_n548_; 
wire u0_u0__abc_72207_new_n549_; 
wire u0_u0__abc_72207_new_n550_; 
wire u0_u0__abc_72207_new_n551_; 
wire u0_u0__abc_72207_new_n552_; 
wire u0_u0__abc_72207_new_n553_; 
wire u0_u0__abc_72207_new_n554_; 
wire u0_u0__abc_72207_new_n555_; 
wire u0_u0__abc_72207_new_n556_; 
wire u0_u0__abc_72207_new_n557_; 
wire u0_u0__abc_72207_new_n558_; 
wire u0_u0__abc_72207_new_n559_; 
wire u0_u0__abc_72207_new_n560_; 
wire u0_u0__abc_72207_new_n561_; 
wire u0_u0__abc_72207_new_n562_; 
wire u0_u0__abc_72207_new_n563_; 
wire u0_u0__abc_72207_new_n565_; 
wire u0_u0__abc_72207_new_n568_; 
wire u0_u0__abc_72207_new_n569_; 
wire u0_u0__abc_72207_new_n570_; 
wire u0_u0__abc_72207_new_n571_; 
wire u0_u0__abc_72207_new_n572_; 
wire u0_u0__abc_72207_new_n573_; 
wire u0_u0_addr_r_2_; 
wire u0_u0_addr_r_3_; 
wire u0_u0_addr_r_4_; 
wire u0_u0_addr_r_5_; 
wire u0_u0_addr_r_6_; 
wire u0_u0_init_req_we; 
wire u0_u0_inited; 
wire u0_u0_lmr_req_we; 
wire u0_u0_rst_r2; 
wire u0_u0_rst_r2_bF_buf0; 
wire u0_u0_rst_r2_bF_buf1; 
wire u0_u0_rst_r2_bF_buf2; 
wire u0_u0_rst_r2_bF_buf3; 
wire u0_u0_rst_r2_bF_buf4; 
wire u0_u0_rst_r2_bF_buf5; 
wire u0_u0_wp_err; 
wire u0_u1__0csc_31_0__0_; 
wire u0_u1__0csc_31_0__10_; 
wire u0_u1__0csc_31_0__11_; 
wire u0_u1__0csc_31_0__12_; 
wire u0_u1__0csc_31_0__13_; 
wire u0_u1__0csc_31_0__14_; 
wire u0_u1__0csc_31_0__15_; 
wire u0_u1__0csc_31_0__16_; 
wire u0_u1__0csc_31_0__17_; 
wire u0_u1__0csc_31_0__18_; 
wire u0_u1__0csc_31_0__19_; 
wire u0_u1__0csc_31_0__1_; 
wire u0_u1__0csc_31_0__20_; 
wire u0_u1__0csc_31_0__21_; 
wire u0_u1__0csc_31_0__22_; 
wire u0_u1__0csc_31_0__23_; 
wire u0_u1__0csc_31_0__24_; 
wire u0_u1__0csc_31_0__25_; 
wire u0_u1__0csc_31_0__26_; 
wire u0_u1__0csc_31_0__27_; 
wire u0_u1__0csc_31_0__28_; 
wire u0_u1__0csc_31_0__29_; 
wire u0_u1__0csc_31_0__2_; 
wire u0_u1__0csc_31_0__30_; 
wire u0_u1__0csc_31_0__31_; 
wire u0_u1__0csc_31_0__3_; 
wire u0_u1__0csc_31_0__4_; 
wire u0_u1__0csc_31_0__5_; 
wire u0_u1__0csc_31_0__6_; 
wire u0_u1__0csc_31_0__7_; 
wire u0_u1__0csc_31_0__8_; 
wire u0_u1__0csc_31_0__9_; 
wire u0_u1__0init_req_0_0_; 
wire u0_u1__0init_req_we_0_0_; 
wire u0_u1__0init_req_we_0_0_bF_buf0_; 
wire u0_u1__0init_req_we_0_0_bF_buf1_; 
wire u0_u1__0init_req_we_0_0_bF_buf2_; 
wire u0_u1__0init_req_we_0_0_bF_buf3_; 
wire u0_u1__0init_req_we_0_0_bF_buf4_; 
wire u0_u1__0init_req_we_0_0_bF_buf5_; 
wire u0_u1__0init_req_we_0_0_bF_buf6_; 
wire u0_u1__0init_req_we_0_0_bF_buf7_; 
wire u0_u1__0inited_0_0_; 
wire u0_u1__0lmr_req_0_0_; 
wire u0_u1__0lmr_req_we_0_0_; 
wire u0_u1__0lmr_req_we_0_0_bF_buf0_; 
wire u0_u1__0lmr_req_we_0_0_bF_buf1_; 
wire u0_u1__0lmr_req_we_0_0_bF_buf2_; 
wire u0_u1__0lmr_req_we_0_0_bF_buf3_; 
wire u0_u1__0lmr_req_we_0_0_bF_buf4_; 
wire u0_u1__0lmr_req_we_0_0_bF_buf5_; 
wire u0_u1__0lmr_req_we_0_0_bF_buf6_; 
wire u0_u1__0lmr_req_we_0_0_bF_buf7_; 
wire u0_u1__0tms_31_0__0_; 
wire u0_u1__0tms_31_0__10_; 
wire u0_u1__0tms_31_0__11_; 
wire u0_u1__0tms_31_0__12_; 
wire u0_u1__0tms_31_0__13_; 
wire u0_u1__0tms_31_0__14_; 
wire u0_u1__0tms_31_0__15_; 
wire u0_u1__0tms_31_0__16_; 
wire u0_u1__0tms_31_0__17_; 
wire u0_u1__0tms_31_0__18_; 
wire u0_u1__0tms_31_0__19_; 
wire u0_u1__0tms_31_0__1_; 
wire u0_u1__0tms_31_0__20_; 
wire u0_u1__0tms_31_0__21_; 
wire u0_u1__0tms_31_0__22_; 
wire u0_u1__0tms_31_0__23_; 
wire u0_u1__0tms_31_0__24_; 
wire u0_u1__0tms_31_0__25_; 
wire u0_u1__0tms_31_0__26_; 
wire u0_u1__0tms_31_0__27_; 
wire u0_u1__0tms_31_0__28_; 
wire u0_u1__0tms_31_0__29_; 
wire u0_u1__0tms_31_0__2_; 
wire u0_u1__0tms_31_0__30_; 
wire u0_u1__0tms_31_0__31_; 
wire u0_u1__0tms_31_0__3_; 
wire u0_u1__0tms_31_0__4_; 
wire u0_u1__0tms_31_0__5_; 
wire u0_u1__0tms_31_0__6_; 
wire u0_u1__0tms_31_0__7_; 
wire u0_u1__0tms_31_0__8_; 
wire u0_u1__0tms_31_0__9_; 
wire u0_u1__abc_72579_auto_rtlil_cc_1942_NotGate_71506; 
wire u0_u1__abc_72579_new_n201_; 
wire u0_u1__abc_72579_new_n202_; 
wire u0_u1__abc_72579_new_n203_; 
wire u0_u1__abc_72579_new_n204_; 
wire u0_u1__abc_72579_new_n205_; 
wire u0_u1__abc_72579_new_n206_; 
wire u0_u1__abc_72579_new_n207_; 
wire u0_u1__abc_72579_new_n208_; 
wire u0_u1__abc_72579_new_n209_; 
wire u0_u1__abc_72579_new_n211_; 
wire u0_u1__abc_72579_new_n212_; 
wire u0_u1__abc_72579_new_n213_; 
wire u0_u1__abc_72579_new_n214_; 
wire u0_u1__abc_72579_new_n215_; 
wire u0_u1__abc_72579_new_n216_; 
wire u0_u1__abc_72579_new_n218_; 
wire u0_u1__abc_72579_new_n219_; 
wire u0_u1__abc_72579_new_n219__bF_buf0; 
wire u0_u1__abc_72579_new_n219__bF_buf1; 
wire u0_u1__abc_72579_new_n219__bF_buf2; 
wire u0_u1__abc_72579_new_n219__bF_buf3; 
wire u0_u1__abc_72579_new_n219__bF_buf4; 
wire u0_u1__abc_72579_new_n219__bF_buf5; 
wire u0_u1__abc_72579_new_n219__bF_buf6; 
wire u0_u1__abc_72579_new_n219__bF_buf7; 
wire u0_u1__abc_72579_new_n220_; 
wire u0_u1__abc_72579_new_n221_; 
wire u0_u1__abc_72579_new_n222_; 
wire u0_u1__abc_72579_new_n223_; 
wire u0_u1__abc_72579_new_n225_; 
wire u0_u1__abc_72579_new_n226_; 
wire u0_u1__abc_72579_new_n227_; 
wire u0_u1__abc_72579_new_n228_; 
wire u0_u1__abc_72579_new_n229_; 
wire u0_u1__abc_72579_new_n231_; 
wire u0_u1__abc_72579_new_n232_; 
wire u0_u1__abc_72579_new_n233_; 
wire u0_u1__abc_72579_new_n234_; 
wire u0_u1__abc_72579_new_n235_; 
wire u0_u1__abc_72579_new_n237_; 
wire u0_u1__abc_72579_new_n238_; 
wire u0_u1__abc_72579_new_n239_; 
wire u0_u1__abc_72579_new_n240_; 
wire u0_u1__abc_72579_new_n241_; 
wire u0_u1__abc_72579_new_n243_; 
wire u0_u1__abc_72579_new_n244_; 
wire u0_u1__abc_72579_new_n245_; 
wire u0_u1__abc_72579_new_n246_; 
wire u0_u1__abc_72579_new_n247_; 
wire u0_u1__abc_72579_new_n249_; 
wire u0_u1__abc_72579_new_n250_; 
wire u0_u1__abc_72579_new_n251_; 
wire u0_u1__abc_72579_new_n252_; 
wire u0_u1__abc_72579_new_n253_; 
wire u0_u1__abc_72579_new_n255_; 
wire u0_u1__abc_72579_new_n256_; 
wire u0_u1__abc_72579_new_n257_; 
wire u0_u1__abc_72579_new_n258_; 
wire u0_u1__abc_72579_new_n259_; 
wire u0_u1__abc_72579_new_n261_; 
wire u0_u1__abc_72579_new_n262_; 
wire u0_u1__abc_72579_new_n263_; 
wire u0_u1__abc_72579_new_n264_; 
wire u0_u1__abc_72579_new_n265_; 
wire u0_u1__abc_72579_new_n267_; 
wire u0_u1__abc_72579_new_n268_; 
wire u0_u1__abc_72579_new_n269_; 
wire u0_u1__abc_72579_new_n270_; 
wire u0_u1__abc_72579_new_n271_; 
wire u0_u1__abc_72579_new_n273_; 
wire u0_u1__abc_72579_new_n274_; 
wire u0_u1__abc_72579_new_n275_; 
wire u0_u1__abc_72579_new_n276_; 
wire u0_u1__abc_72579_new_n277_; 
wire u0_u1__abc_72579_new_n279_; 
wire u0_u1__abc_72579_new_n280_; 
wire u0_u1__abc_72579_new_n281_; 
wire u0_u1__abc_72579_new_n282_; 
wire u0_u1__abc_72579_new_n283_; 
wire u0_u1__abc_72579_new_n285_; 
wire u0_u1__abc_72579_new_n286_; 
wire u0_u1__abc_72579_new_n287_; 
wire u0_u1__abc_72579_new_n288_; 
wire u0_u1__abc_72579_new_n289_; 
wire u0_u1__abc_72579_new_n291_; 
wire u0_u1__abc_72579_new_n292_; 
wire u0_u1__abc_72579_new_n293_; 
wire u0_u1__abc_72579_new_n294_; 
wire u0_u1__abc_72579_new_n295_; 
wire u0_u1__abc_72579_new_n297_; 
wire u0_u1__abc_72579_new_n298_; 
wire u0_u1__abc_72579_new_n299_; 
wire u0_u1__abc_72579_new_n300_; 
wire u0_u1__abc_72579_new_n301_; 
wire u0_u1__abc_72579_new_n303_; 
wire u0_u1__abc_72579_new_n304_; 
wire u0_u1__abc_72579_new_n305_; 
wire u0_u1__abc_72579_new_n306_; 
wire u0_u1__abc_72579_new_n307_; 
wire u0_u1__abc_72579_new_n309_; 
wire u0_u1__abc_72579_new_n310_; 
wire u0_u1__abc_72579_new_n311_; 
wire u0_u1__abc_72579_new_n312_; 
wire u0_u1__abc_72579_new_n313_; 
wire u0_u1__abc_72579_new_n315_; 
wire u0_u1__abc_72579_new_n316_; 
wire u0_u1__abc_72579_new_n317_; 
wire u0_u1__abc_72579_new_n318_; 
wire u0_u1__abc_72579_new_n319_; 
wire u0_u1__abc_72579_new_n321_; 
wire u0_u1__abc_72579_new_n322_; 
wire u0_u1__abc_72579_new_n323_; 
wire u0_u1__abc_72579_new_n324_; 
wire u0_u1__abc_72579_new_n325_; 
wire u0_u1__abc_72579_new_n327_; 
wire u0_u1__abc_72579_new_n328_; 
wire u0_u1__abc_72579_new_n329_; 
wire u0_u1__abc_72579_new_n330_; 
wire u0_u1__abc_72579_new_n331_; 
wire u0_u1__abc_72579_new_n333_; 
wire u0_u1__abc_72579_new_n334_; 
wire u0_u1__abc_72579_new_n335_; 
wire u0_u1__abc_72579_new_n336_; 
wire u0_u1__abc_72579_new_n337_; 
wire u0_u1__abc_72579_new_n339_; 
wire u0_u1__abc_72579_new_n340_; 
wire u0_u1__abc_72579_new_n341_; 
wire u0_u1__abc_72579_new_n342_; 
wire u0_u1__abc_72579_new_n343_; 
wire u0_u1__abc_72579_new_n345_; 
wire u0_u1__abc_72579_new_n346_; 
wire u0_u1__abc_72579_new_n347_; 
wire u0_u1__abc_72579_new_n348_; 
wire u0_u1__abc_72579_new_n349_; 
wire u0_u1__abc_72579_new_n351_; 
wire u0_u1__abc_72579_new_n352_; 
wire u0_u1__abc_72579_new_n353_; 
wire u0_u1__abc_72579_new_n354_; 
wire u0_u1__abc_72579_new_n355_; 
wire u0_u1__abc_72579_new_n357_; 
wire u0_u1__abc_72579_new_n358_; 
wire u0_u1__abc_72579_new_n359_; 
wire u0_u1__abc_72579_new_n360_; 
wire u0_u1__abc_72579_new_n361_; 
wire u0_u1__abc_72579_new_n363_; 
wire u0_u1__abc_72579_new_n364_; 
wire u0_u1__abc_72579_new_n365_; 
wire u0_u1__abc_72579_new_n366_; 
wire u0_u1__abc_72579_new_n367_; 
wire u0_u1__abc_72579_new_n369_; 
wire u0_u1__abc_72579_new_n370_; 
wire u0_u1__abc_72579_new_n371_; 
wire u0_u1__abc_72579_new_n372_; 
wire u0_u1__abc_72579_new_n373_; 
wire u0_u1__abc_72579_new_n375_; 
wire u0_u1__abc_72579_new_n376_; 
wire u0_u1__abc_72579_new_n377_; 
wire u0_u1__abc_72579_new_n378_; 
wire u0_u1__abc_72579_new_n379_; 
wire u0_u1__abc_72579_new_n381_; 
wire u0_u1__abc_72579_new_n382_; 
wire u0_u1__abc_72579_new_n383_; 
wire u0_u1__abc_72579_new_n384_; 
wire u0_u1__abc_72579_new_n385_; 
wire u0_u1__abc_72579_new_n387_; 
wire u0_u1__abc_72579_new_n388_; 
wire u0_u1__abc_72579_new_n389_; 
wire u0_u1__abc_72579_new_n390_; 
wire u0_u1__abc_72579_new_n391_; 
wire u0_u1__abc_72579_new_n393_; 
wire u0_u1__abc_72579_new_n394_; 
wire u0_u1__abc_72579_new_n395_; 
wire u0_u1__abc_72579_new_n396_; 
wire u0_u1__abc_72579_new_n397_; 
wire u0_u1__abc_72579_new_n399_; 
wire u0_u1__abc_72579_new_n400_; 
wire u0_u1__abc_72579_new_n401_; 
wire u0_u1__abc_72579_new_n402_; 
wire u0_u1__abc_72579_new_n403_; 
wire u0_u1__abc_72579_new_n405_; 
wire u0_u1__abc_72579_new_n406_; 
wire u0_u1__abc_72579_new_n407_; 
wire u0_u1__abc_72579_new_n408_; 
wire u0_u1__abc_72579_new_n409_; 
wire u0_u1__abc_72579_new_n411_; 
wire u0_u1__abc_72579_new_n413_; 
wire u0_u1__abc_72579_new_n414_; 
wire u0_u1__abc_72579_new_n415_; 
wire u0_u1__abc_72579_new_n416_; 
wire u0_u1__abc_72579_new_n418_; 
wire u0_u1__abc_72579_new_n419_; 
wire u0_u1__abc_72579_new_n420_; 
wire u0_u1__abc_72579_new_n421_; 
wire u0_u1__abc_72579_new_n423_; 
wire u0_u1__abc_72579_new_n424_; 
wire u0_u1__abc_72579_new_n425_; 
wire u0_u1__abc_72579_new_n426_; 
wire u0_u1__abc_72579_new_n428_; 
wire u0_u1__abc_72579_new_n429_; 
wire u0_u1__abc_72579_new_n430_; 
wire u0_u1__abc_72579_new_n431_; 
wire u0_u1__abc_72579_new_n433_; 
wire u0_u1__abc_72579_new_n434_; 
wire u0_u1__abc_72579_new_n435_; 
wire u0_u1__abc_72579_new_n436_; 
wire u0_u1__abc_72579_new_n438_; 
wire u0_u1__abc_72579_new_n439_; 
wire u0_u1__abc_72579_new_n440_; 
wire u0_u1__abc_72579_new_n441_; 
wire u0_u1__abc_72579_new_n443_; 
wire u0_u1__abc_72579_new_n444_; 
wire u0_u1__abc_72579_new_n445_; 
wire u0_u1__abc_72579_new_n446_; 
wire u0_u1__abc_72579_new_n448_; 
wire u0_u1__abc_72579_new_n449_; 
wire u0_u1__abc_72579_new_n450_; 
wire u0_u1__abc_72579_new_n451_; 
wire u0_u1__abc_72579_new_n453_; 
wire u0_u1__abc_72579_new_n454_; 
wire u0_u1__abc_72579_new_n455_; 
wire u0_u1__abc_72579_new_n456_; 
wire u0_u1__abc_72579_new_n458_; 
wire u0_u1__abc_72579_new_n459_; 
wire u0_u1__abc_72579_new_n460_; 
wire u0_u1__abc_72579_new_n461_; 
wire u0_u1__abc_72579_new_n463_; 
wire u0_u1__abc_72579_new_n464_; 
wire u0_u1__abc_72579_new_n465_; 
wire u0_u1__abc_72579_new_n466_; 
wire u0_u1__abc_72579_new_n468_; 
wire u0_u1__abc_72579_new_n469_; 
wire u0_u1__abc_72579_new_n470_; 
wire u0_u1__abc_72579_new_n471_; 
wire u0_u1__abc_72579_new_n473_; 
wire u0_u1__abc_72579_new_n474_; 
wire u0_u1__abc_72579_new_n475_; 
wire u0_u1__abc_72579_new_n476_; 
wire u0_u1__abc_72579_new_n478_; 
wire u0_u1__abc_72579_new_n479_; 
wire u0_u1__abc_72579_new_n480_; 
wire u0_u1__abc_72579_new_n481_; 
wire u0_u1__abc_72579_new_n483_; 
wire u0_u1__abc_72579_new_n484_; 
wire u0_u1__abc_72579_new_n485_; 
wire u0_u1__abc_72579_new_n486_; 
wire u0_u1__abc_72579_new_n488_; 
wire u0_u1__abc_72579_new_n489_; 
wire u0_u1__abc_72579_new_n490_; 
wire u0_u1__abc_72579_new_n491_; 
wire u0_u1__abc_72579_new_n493_; 
wire u0_u1__abc_72579_new_n494_; 
wire u0_u1__abc_72579_new_n495_; 
wire u0_u1__abc_72579_new_n496_; 
wire u0_u1__abc_72579_new_n498_; 
wire u0_u1__abc_72579_new_n499_; 
wire u0_u1__abc_72579_new_n500_; 
wire u0_u1__abc_72579_new_n501_; 
wire u0_u1__abc_72579_new_n503_; 
wire u0_u1__abc_72579_new_n504_; 
wire u0_u1__abc_72579_new_n505_; 
wire u0_u1__abc_72579_new_n506_; 
wire u0_u1__abc_72579_new_n508_; 
wire u0_u1__abc_72579_new_n509_; 
wire u0_u1__abc_72579_new_n510_; 
wire u0_u1__abc_72579_new_n511_; 
wire u0_u1__abc_72579_new_n513_; 
wire u0_u1__abc_72579_new_n514_; 
wire u0_u1__abc_72579_new_n515_; 
wire u0_u1__abc_72579_new_n516_; 
wire u0_u1__abc_72579_new_n518_; 
wire u0_u1__abc_72579_new_n519_; 
wire u0_u1__abc_72579_new_n520_; 
wire u0_u1__abc_72579_new_n521_; 
wire u0_u1__abc_72579_new_n523_; 
wire u0_u1__abc_72579_new_n524_; 
wire u0_u1__abc_72579_new_n525_; 
wire u0_u1__abc_72579_new_n526_; 
wire u0_u1__abc_72579_new_n528_; 
wire u0_u1__abc_72579_new_n529_; 
wire u0_u1__abc_72579_new_n530_; 
wire u0_u1__abc_72579_new_n531_; 
wire u0_u1__abc_72579_new_n533_; 
wire u0_u1__abc_72579_new_n534_; 
wire u0_u1__abc_72579_new_n535_; 
wire u0_u1__abc_72579_new_n536_; 
wire u0_u1__abc_72579_new_n538_; 
wire u0_u1__abc_72579_new_n539_; 
wire u0_u1__abc_72579_new_n540_; 
wire u0_u1__abc_72579_new_n541_; 
wire u0_u1__abc_72579_new_n543_; 
wire u0_u1__abc_72579_new_n544_; 
wire u0_u1__abc_72579_new_n545_; 
wire u0_u1__abc_72579_new_n546_; 
wire u0_u1__abc_72579_new_n548_; 
wire u0_u1__abc_72579_new_n549_; 
wire u0_u1__abc_72579_new_n550_; 
wire u0_u1__abc_72579_new_n551_; 
wire u0_u1__abc_72579_new_n553_; 
wire u0_u1__abc_72579_new_n554_; 
wire u0_u1__abc_72579_new_n555_; 
wire u0_u1__abc_72579_new_n556_; 
wire u0_u1__abc_72579_new_n558_; 
wire u0_u1__abc_72579_new_n559_; 
wire u0_u1__abc_72579_new_n560_; 
wire u0_u1__abc_72579_new_n561_; 
wire u0_u1__abc_72579_new_n563_; 
wire u0_u1__abc_72579_new_n564_; 
wire u0_u1__abc_72579_new_n565_; 
wire u0_u1__abc_72579_new_n566_; 
wire u0_u1__abc_72579_new_n568_; 
wire u0_u1__abc_72579_new_n569_; 
wire u0_u1__abc_72579_new_n570_; 
wire u0_u1__abc_72579_new_n571_; 
wire u0_u1__abc_72579_new_n573_; 
wire u0_u1__abc_72579_new_n574_; 
wire u0_u1__abc_72579_new_n575_; 
wire u0_u1__abc_72579_new_n576_; 
wire u0_u1__abc_72579_new_n577_; 
wire u0_u1__abc_72579_new_n578_; 
wire u0_u1__abc_72579_new_n579_; 
wire u0_u1__abc_72579_new_n580_; 
wire u0_u1__abc_72579_new_n581_; 
wire u0_u1__abc_72579_new_n582_; 
wire u0_u1__abc_72579_new_n583_; 
wire u0_u1__abc_72579_new_n584_; 
wire u0_u1__abc_72579_new_n585_; 
wire u0_u1__abc_72579_new_n586_; 
wire u0_u1__abc_72579_new_n587_; 
wire u0_u1__abc_72579_new_n588_; 
wire u0_u1__abc_72579_new_n589_; 
wire u0_u1__abc_72579_new_n590_; 
wire u0_u1__abc_72579_new_n591_; 
wire u0_u1__abc_72579_new_n592_; 
wire u0_u1__abc_72579_new_n593_; 
wire u0_u1__abc_72579_new_n594_; 
wire u0_u1__abc_72579_new_n595_; 
wire u0_u1__abc_72579_new_n596_; 
wire u0_u1__abc_72579_new_n597_; 
wire u0_u1__abc_72579_new_n598_; 
wire u0_u1__abc_72579_new_n599_; 
wire u0_u1__abc_72579_new_n600_; 
wire u0_u1__abc_72579_new_n601_; 
wire u0_u1__abc_72579_new_n602_; 
wire u0_u1__abc_72579_new_n603_; 
wire u0_u1__abc_72579_new_n604_; 
wire u0_u1__abc_72579_new_n605_; 
wire u0_u1__abc_72579_new_n606_; 
wire u0_u1__abc_72579_new_n607_; 
wire u0_u1__abc_72579_new_n608_; 
wire u0_u1__abc_72579_new_n609_; 
wire u0_u1__abc_72579_new_n610_; 
wire u0_u1__abc_72579_new_n611_; 
wire u0_u1__abc_72579_new_n612_; 
wire u0_u1__abc_72579_new_n613_; 
wire u0_u1__abc_72579_new_n614_; 
wire u0_u1__abc_72579_new_n615_; 
wire u0_u1__abc_72579_new_n616_; 
wire u0_u1__abc_72579_new_n617_; 
wire u0_u1__abc_72579_new_n618_; 
wire u0_u1__abc_72579_new_n619_; 
wire u0_u1__abc_72579_new_n620_; 
wire u0_u1__abc_72579_new_n621_; 
wire u0_u1__abc_72579_new_n622_; 
wire u0_u1__abc_72579_new_n623_; 
wire u0_u1__abc_72579_new_n624_; 
wire u0_u1__abc_72579_new_n625_; 
wire u0_u1__abc_72579_new_n626_; 
wire u0_u1__abc_72579_new_n627_; 
wire u0_u1__abc_72579_new_n628_; 
wire u0_u1__abc_72579_new_n629_; 
wire u0_u1__abc_72579_new_n630_; 
wire u0_u1__abc_72579_new_n631_; 
wire u0_u1__abc_72579_new_n632_; 
wire u0_u1__abc_72579_new_n633_; 
wire u0_u1__abc_72579_new_n634_; 
wire u0_u1__abc_72579_new_n635_; 
wire u0_u1__abc_72579_new_n636_; 
wire u0_u1__abc_72579_new_n637_; 
wire u0_u1__abc_72579_new_n639_; 
wire u0_u1__abc_72579_new_n642_; 
wire u0_u1__abc_72579_new_n643_; 
wire u0_u1__abc_72579_new_n644_; 
wire u0_u1__abc_72579_new_n645_; 
wire u0_u1__abc_72579_new_n646_; 
wire u0_u1__abc_72579_new_n647_; 
wire u0_u1_addr_r_2_; 
wire u0_u1_addr_r_3_; 
wire u0_u1_addr_r_4_; 
wire u0_u1_addr_r_5_; 
wire u0_u1_addr_r_6_; 
wire u0_u1_init_req_we; 
wire u0_u1_inited; 
wire u0_u1_lmr_req_we; 
wire u0_u1_rst_r2; 
wire u0_u1_wp_err; 
wire u0_wb_addr_r_2_; 
wire u0_wb_addr_r_3_; 
wire u0_wb_addr_r_4_; 
wire u0_wb_addr_r_5_; 
wire u0_wb_addr_r_6_; 
wire u0_wp_err; 
wire u1__0acs_addr_23_0__0_; 
wire u1__0acs_addr_23_0__10_; 
wire u1__0acs_addr_23_0__11_; 
wire u1__0acs_addr_23_0__12_; 
wire u1__0acs_addr_23_0__13_; 
wire u1__0acs_addr_23_0__14_; 
wire u1__0acs_addr_23_0__15_; 
wire u1__0acs_addr_23_0__16_; 
wire u1__0acs_addr_23_0__17_; 
wire u1__0acs_addr_23_0__18_; 
wire u1__0acs_addr_23_0__19_; 
wire u1__0acs_addr_23_0__1_; 
wire u1__0acs_addr_23_0__20_; 
wire u1__0acs_addr_23_0__21_; 
wire u1__0acs_addr_23_0__22_; 
wire u1__0acs_addr_23_0__23_; 
wire u1__0acs_addr_23_0__2_; 
wire u1__0acs_addr_23_0__3_; 
wire u1__0acs_addr_23_0__4_; 
wire u1__0acs_addr_23_0__5_; 
wire u1__0acs_addr_23_0__6_; 
wire u1__0acs_addr_23_0__7_; 
wire u1__0acs_addr_23_0__8_; 
wire u1__0acs_addr_23_0__9_; 
wire u1__0bank_adr_1_0__0_; 
wire u1__0bank_adr_1_0__1_; 
wire u1__0col_adr_9_0__0_; 
wire u1__0col_adr_9_0__1_; 
wire u1__0col_adr_9_0__2_; 
wire u1__0col_adr_9_0__3_; 
wire u1__0col_adr_9_0__4_; 
wire u1__0col_adr_9_0__5_; 
wire u1__0col_adr_9_0__6_; 
wire u1__0col_adr_9_0__7_; 
wire u1__0col_adr_9_0__8_; 
wire u1__0col_adr_9_0__9_; 
wire u1__0row_adr_12_0__0_; 
wire u1__0row_adr_12_0__10_; 
wire u1__0row_adr_12_0__11_; 
wire u1__0row_adr_12_0__12_; 
wire u1__0row_adr_12_0__1_; 
wire u1__0row_adr_12_0__2_; 
wire u1__0row_adr_12_0__3_; 
wire u1__0row_adr_12_0__4_; 
wire u1__0row_adr_12_0__5_; 
wire u1__0row_adr_12_0__6_; 
wire u1__0row_adr_12_0__7_; 
wire u1__0row_adr_12_0__8_; 
wire u1__0row_adr_12_0__9_; 
wire u1__0sram_addr_23_0__0_; 
wire u1__0sram_addr_23_0__10_; 
wire u1__0sram_addr_23_0__11_; 
wire u1__0sram_addr_23_0__12_; 
wire u1__0sram_addr_23_0__13_; 
wire u1__0sram_addr_23_0__14_; 
wire u1__0sram_addr_23_0__15_; 
wire u1__0sram_addr_23_0__16_; 
wire u1__0sram_addr_23_0__17_; 
wire u1__0sram_addr_23_0__18_; 
wire u1__0sram_addr_23_0__19_; 
wire u1__0sram_addr_23_0__1_; 
wire u1__0sram_addr_23_0__20_; 
wire u1__0sram_addr_23_0__21_; 
wire u1__0sram_addr_23_0__22_; 
wire u1__0sram_addr_23_0__23_; 
wire u1__0sram_addr_23_0__2_; 
wire u1__0sram_addr_23_0__3_; 
wire u1__0sram_addr_23_0__4_; 
wire u1__0sram_addr_23_0__5_; 
wire u1__0sram_addr_23_0__6_; 
wire u1__0sram_addr_23_0__7_; 
wire u1__0sram_addr_23_0__8_; 
wire u1__0sram_addr_23_0__9_; 
wire u1__abc_73140_new_n1000_; 
wire u1__abc_73140_new_n1001_; 
wire u1__abc_73140_new_n1002_; 
wire u1__abc_73140_new_n1004_; 
wire u1__abc_73140_new_n1005_; 
wire u1__abc_73140_new_n1006_; 
wire u1__abc_73140_new_n1007_; 
wire u1__abc_73140_new_n1008_; 
wire u1__abc_73140_new_n1009_; 
wire u1__abc_73140_new_n1010_; 
wire u1__abc_73140_new_n1011_; 
wire u1__abc_73140_new_n1012_; 
wire u1__abc_73140_new_n1013_; 
wire u1__abc_73140_new_n1014_; 
wire u1__abc_73140_new_n1015_; 
wire u1__abc_73140_new_n1016_; 
wire u1__abc_73140_new_n1017_; 
wire u1__abc_73140_new_n1019_; 
wire u1__abc_73140_new_n1020_; 
wire u1__abc_73140_new_n1021_; 
wire u1__abc_73140_new_n1022_; 
wire u1__abc_73140_new_n1023_; 
wire u1__abc_73140_new_n1024_; 
wire u1__abc_73140_new_n1025_; 
wire u1__abc_73140_new_n1026_; 
wire u1__abc_73140_new_n1027_; 
wire u1__abc_73140_new_n1028_; 
wire u1__abc_73140_new_n1029_; 
wire u1__abc_73140_new_n1030_; 
wire u1__abc_73140_new_n1031_; 
wire u1__abc_73140_new_n1032_; 
wire u1__abc_73140_new_n1034_; 
wire u1__abc_73140_new_n1035_; 
wire u1__abc_73140_new_n1036_; 
wire u1__abc_73140_new_n1037_; 
wire u1__abc_73140_new_n1038_; 
wire u1__abc_73140_new_n1039_; 
wire u1__abc_73140_new_n1040_; 
wire u1__abc_73140_new_n1041_; 
wire u1__abc_73140_new_n1042_; 
wire u1__abc_73140_new_n1043_; 
wire u1__abc_73140_new_n1044_; 
wire u1__abc_73140_new_n1045_; 
wire u1__abc_73140_new_n1046_; 
wire u1__abc_73140_new_n1047_; 
wire u1__abc_73140_new_n1049_; 
wire u1__abc_73140_new_n1050_; 
wire u1__abc_73140_new_n1051_; 
wire u1__abc_73140_new_n1052_; 
wire u1__abc_73140_new_n1053_; 
wire u1__abc_73140_new_n1054_; 
wire u1__abc_73140_new_n1055_; 
wire u1__abc_73140_new_n1056_; 
wire u1__abc_73140_new_n1057_; 
wire u1__abc_73140_new_n1058_; 
wire u1__abc_73140_new_n1059_; 
wire u1__abc_73140_new_n1060_; 
wire u1__abc_73140_new_n1061_; 
wire u1__abc_73140_new_n1062_; 
wire u1__abc_73140_new_n1064_; 
wire u1__abc_73140_new_n1065_; 
wire u1__abc_73140_new_n1066_; 
wire u1__abc_73140_new_n1067_; 
wire u1__abc_73140_new_n1068_; 
wire u1__abc_73140_new_n1069_; 
wire u1__abc_73140_new_n1070_; 
wire u1__abc_73140_new_n1071_; 
wire u1__abc_73140_new_n1072_; 
wire u1__abc_73140_new_n1073_; 
wire u1__abc_73140_new_n1074_; 
wire u1__abc_73140_new_n1075_; 
wire u1__abc_73140_new_n1077_; 
wire u1__abc_73140_new_n1078_; 
wire u1__abc_73140_new_n1079_; 
wire u1__abc_73140_new_n1080_; 
wire u1__abc_73140_new_n1081_; 
wire u1__abc_73140_new_n1082_; 
wire u1__abc_73140_new_n1083_; 
wire u1__abc_73140_new_n1084_; 
wire u1__abc_73140_new_n1085_; 
wire u1__abc_73140_new_n1086_; 
wire u1__abc_73140_new_n1087_; 
wire u1__abc_73140_new_n1088_; 
wire u1__abc_73140_new_n1090_; 
wire u1__abc_73140_new_n1091_; 
wire u1__abc_73140_new_n1092_; 
wire u1__abc_73140_new_n1093_; 
wire u1__abc_73140_new_n1094_; 
wire u1__abc_73140_new_n1095_; 
wire u1__abc_73140_new_n1096_; 
wire u1__abc_73140_new_n1097_; 
wire u1__abc_73140_new_n1099_; 
wire u1__abc_73140_new_n1100_; 
wire u1__abc_73140_new_n1101_; 
wire u1__abc_73140_new_n1102_; 
wire u1__abc_73140_new_n1103_; 
wire u1__abc_73140_new_n1104_; 
wire u1__abc_73140_new_n1105_; 
wire u1__abc_73140_new_n1106_; 
wire u1__abc_73140_new_n1108_; 
wire u1__abc_73140_new_n1109_; 
wire u1__abc_73140_new_n1110_; 
wire u1__abc_73140_new_n1111_; 
wire u1__abc_73140_new_n1112_; 
wire u1__abc_73140_new_n1113_; 
wire u1__abc_73140_new_n1115_; 
wire u1__abc_73140_new_n1116_; 
wire u1__abc_73140_new_n1117_; 
wire u1__abc_73140_new_n1118_; 
wire u1__abc_73140_new_n1119_; 
wire u1__abc_73140_new_n1120_; 
wire u1__abc_73140_new_n1122_; 
wire u1__abc_73140_new_n1123_; 
wire u1__abc_73140_new_n1124_; 
wire u1__abc_73140_new_n1125_; 
wire u1__abc_73140_new_n1126_; 
wire u1__abc_73140_new_n1127_; 
wire u1__abc_73140_new_n1129_; 
wire u1__abc_73140_new_n1130_; 
wire u1__abc_73140_new_n1131_; 
wire u1__abc_73140_new_n1132_; 
wire u1__abc_73140_new_n1133_; 
wire u1__abc_73140_new_n1134_; 
wire u1__abc_73140_new_n1136_; 
wire u1__abc_73140_new_n1137_; 
wire u1__abc_73140_new_n1138_; 
wire u1__abc_73140_new_n1139_; 
wire u1__abc_73140_new_n1140_; 
wire u1__abc_73140_new_n1141_; 
wire u1__abc_73140_new_n1143_; 
wire u1__abc_73140_new_n1144_; 
wire u1__abc_73140_new_n1145_; 
wire u1__abc_73140_new_n1146_; 
wire u1__abc_73140_new_n1147_; 
wire u1__abc_73140_new_n1148_; 
wire u1__abc_73140_new_n1150_; 
wire u1__abc_73140_new_n1151_; 
wire u1__abc_73140_new_n1152_; 
wire u1__abc_73140_new_n1153_; 
wire u1__abc_73140_new_n1154_; 
wire u1__abc_73140_new_n1155_; 
wire u1__abc_73140_new_n1157_; 
wire u1__abc_73140_new_n1158_; 
wire u1__abc_73140_new_n1159_; 
wire u1__abc_73140_new_n1160_; 
wire u1__abc_73140_new_n1161_; 
wire u1__abc_73140_new_n1162_; 
wire u1__abc_73140_new_n1164_; 
wire u1__abc_73140_new_n1165_; 
wire u1__abc_73140_new_n1166_; 
wire u1__abc_73140_new_n1167_; 
wire u1__abc_73140_new_n1168_; 
wire u1__abc_73140_new_n1169_; 
wire u1__abc_73140_new_n1171_; 
wire u1__abc_73140_new_n1172_; 
wire u1__abc_73140_new_n1173_; 
wire u1__abc_73140_new_n1174_; 
wire u1__abc_73140_new_n1175_; 
wire u1__abc_73140_new_n1176_; 
wire u1__abc_73140_new_n1177_; 
wire u1__abc_73140_new_n1178_; 
wire u1__abc_73140_new_n1179_; 
wire u1__abc_73140_new_n1180_; 
wire u1__abc_73140_new_n1181_; 
wire u1__abc_73140_new_n1182_; 
wire u1__abc_73140_new_n1183_; 
wire u1__abc_73140_new_n1184_; 
wire u1__abc_73140_new_n1185_; 
wire u1__abc_73140_new_n258_; 
wire u1__abc_73140_new_n259_; 
wire u1__abc_73140_new_n260_; 
wire u1__abc_73140_new_n261_; 
wire u1__abc_73140_new_n262_; 
wire u1__abc_73140_new_n263_; 
wire u1__abc_73140_new_n264_; 
wire u1__abc_73140_new_n265_; 
wire u1__abc_73140_new_n266_; 
wire u1__abc_73140_new_n267_; 
wire u1__abc_73140_new_n268_; 
wire u1__abc_73140_new_n268__bF_buf0; 
wire u1__abc_73140_new_n268__bF_buf1; 
wire u1__abc_73140_new_n268__bF_buf2; 
wire u1__abc_73140_new_n268__bF_buf3; 
wire u1__abc_73140_new_n268__bF_buf4; 
wire u1__abc_73140_new_n269_; 
wire u1__abc_73140_new_n270_; 
wire u1__abc_73140_new_n271_; 
wire u1__abc_73140_new_n272_; 
wire u1__abc_73140_new_n273_; 
wire u1__abc_73140_new_n274_; 
wire u1__abc_73140_new_n275_; 
wire u1__abc_73140_new_n275__bF_buf0; 
wire u1__abc_73140_new_n275__bF_buf1; 
wire u1__abc_73140_new_n275__bF_buf2; 
wire u1__abc_73140_new_n275__bF_buf3; 
wire u1__abc_73140_new_n275__bF_buf4; 
wire u1__abc_73140_new_n276_; 
wire u1__abc_73140_new_n277_; 
wire u1__abc_73140_new_n278_; 
wire u1__abc_73140_new_n280_; 
wire u1__abc_73140_new_n282_; 
wire u1__abc_73140_new_n283_; 
wire u1__abc_73140_new_n284_; 
wire u1__abc_73140_new_n285_; 
wire u1__abc_73140_new_n287_; 
wire u1__abc_73140_new_n288_; 
wire u1__abc_73140_new_n289_; 
wire u1__abc_73140_new_n290_; 
wire u1__abc_73140_new_n291_; 
wire u1__abc_73140_new_n292_; 
wire u1__abc_73140_new_n293_; 
wire u1__abc_73140_new_n294_; 
wire u1__abc_73140_new_n295_; 
wire u1__abc_73140_new_n296_; 
wire u1__abc_73140_new_n297_; 
wire u1__abc_73140_new_n298_; 
wire u1__abc_73140_new_n299_; 
wire u1__abc_73140_new_n300_; 
wire u1__abc_73140_new_n301_; 
wire u1__abc_73140_new_n302_; 
wire u1__abc_73140_new_n303_; 
wire u1__abc_73140_new_n304_; 
wire u1__abc_73140_new_n305_; 
wire u1__abc_73140_new_n306_; 
wire u1__abc_73140_new_n307_; 
wire u1__abc_73140_new_n308_; 
wire u1__abc_73140_new_n309_; 
wire u1__abc_73140_new_n310_; 
wire u1__abc_73140_new_n311_; 
wire u1__abc_73140_new_n312_; 
wire u1__abc_73140_new_n313_; 
wire u1__abc_73140_new_n314_; 
wire u1__abc_73140_new_n315_; 
wire u1__abc_73140_new_n316_; 
wire u1__abc_73140_new_n317_; 
wire u1__abc_73140_new_n318_; 
wire u1__abc_73140_new_n319_; 
wire u1__abc_73140_new_n320_; 
wire u1__abc_73140_new_n321_; 
wire u1__abc_73140_new_n322_; 
wire u1__abc_73140_new_n323_; 
wire u1__abc_73140_new_n325_; 
wire u1__abc_73140_new_n326_; 
wire u1__abc_73140_new_n327_; 
wire u1__abc_73140_new_n328_; 
wire u1__abc_73140_new_n329_; 
wire u1__abc_73140_new_n330_; 
wire u1__abc_73140_new_n331_; 
wire u1__abc_73140_new_n332_; 
wire u1__abc_73140_new_n333_; 
wire u1__abc_73140_new_n334_; 
wire u1__abc_73140_new_n335_; 
wire u1__abc_73140_new_n336_; 
wire u1__abc_73140_new_n337_; 
wire u1__abc_73140_new_n338_; 
wire u1__abc_73140_new_n339_; 
wire u1__abc_73140_new_n340_; 
wire u1__abc_73140_new_n341_; 
wire u1__abc_73140_new_n342_; 
wire u1__abc_73140_new_n343_; 
wire u1__abc_73140_new_n344_; 
wire u1__abc_73140_new_n346_; 
wire u1__abc_73140_new_n347_; 
wire u1__abc_73140_new_n348_; 
wire u1__abc_73140_new_n349_; 
wire u1__abc_73140_new_n350_; 
wire u1__abc_73140_new_n351_; 
wire u1__abc_73140_new_n352_; 
wire u1__abc_73140_new_n353_; 
wire u1__abc_73140_new_n354_; 
wire u1__abc_73140_new_n355_; 
wire u1__abc_73140_new_n357_; 
wire u1__abc_73140_new_n358_; 
wire u1__abc_73140_new_n359_; 
wire u1__abc_73140_new_n360_; 
wire u1__abc_73140_new_n361_; 
wire u1__abc_73140_new_n362_; 
wire u1__abc_73140_new_n363_; 
wire u1__abc_73140_new_n364_; 
wire u1__abc_73140_new_n365_; 
wire u1__abc_73140_new_n366_; 
wire u1__abc_73140_new_n367_; 
wire u1__abc_73140_new_n368_; 
wire u1__abc_73140_new_n369_; 
wire u1__abc_73140_new_n370_; 
wire u1__abc_73140_new_n371_; 
wire u1__abc_73140_new_n372_; 
wire u1__abc_73140_new_n373_; 
wire u1__abc_73140_new_n374_; 
wire u1__abc_73140_new_n375_; 
wire u1__abc_73140_new_n377_; 
wire u1__abc_73140_new_n378_; 
wire u1__abc_73140_new_n379_; 
wire u1__abc_73140_new_n380_; 
wire u1__abc_73140_new_n381_; 
wire u1__abc_73140_new_n382_; 
wire u1__abc_73140_new_n383_; 
wire u1__abc_73140_new_n384_; 
wire u1__abc_73140_new_n385_; 
wire u1__abc_73140_new_n386_; 
wire u1__abc_73140_new_n387_; 
wire u1__abc_73140_new_n388_; 
wire u1__abc_73140_new_n390_; 
wire u1__abc_73140_new_n391_; 
wire u1__abc_73140_new_n392_; 
wire u1__abc_73140_new_n393_; 
wire u1__abc_73140_new_n394_; 
wire u1__abc_73140_new_n395_; 
wire u1__abc_73140_new_n396_; 
wire u1__abc_73140_new_n397_; 
wire u1__abc_73140_new_n398_; 
wire u1__abc_73140_new_n399_; 
wire u1__abc_73140_new_n400_; 
wire u1__abc_73140_new_n401_; 
wire u1__abc_73140_new_n403_; 
wire u1__abc_73140_new_n404_; 
wire u1__abc_73140_new_n405_; 
wire u1__abc_73140_new_n406_; 
wire u1__abc_73140_new_n407_; 
wire u1__abc_73140_new_n408_; 
wire u1__abc_73140_new_n409_; 
wire u1__abc_73140_new_n410_; 
wire u1__abc_73140_new_n411_; 
wire u1__abc_73140_new_n412_; 
wire u1__abc_73140_new_n413_; 
wire u1__abc_73140_new_n414_; 
wire u1__abc_73140_new_n416_; 
wire u1__abc_73140_new_n417_; 
wire u1__abc_73140_new_n418_; 
wire u1__abc_73140_new_n419_; 
wire u1__abc_73140_new_n420_; 
wire u1__abc_73140_new_n421_; 
wire u1__abc_73140_new_n422_; 
wire u1__abc_73140_new_n423_; 
wire u1__abc_73140_new_n424_; 
wire u1__abc_73140_new_n425_; 
wire u1__abc_73140_new_n426_; 
wire u1__abc_73140_new_n427_; 
wire u1__abc_73140_new_n429_; 
wire u1__abc_73140_new_n430_; 
wire u1__abc_73140_new_n431_; 
wire u1__abc_73140_new_n432_; 
wire u1__abc_73140_new_n433_; 
wire u1__abc_73140_new_n434_; 
wire u1__abc_73140_new_n435_; 
wire u1__abc_73140_new_n436_; 
wire u1__abc_73140_new_n437_; 
wire u1__abc_73140_new_n438_; 
wire u1__abc_73140_new_n439_; 
wire u1__abc_73140_new_n440_; 
wire u1__abc_73140_new_n442_; 
wire u1__abc_73140_new_n443_; 
wire u1__abc_73140_new_n444_; 
wire u1__abc_73140_new_n445_; 
wire u1__abc_73140_new_n446_; 
wire u1__abc_73140_new_n447_; 
wire u1__abc_73140_new_n448_; 
wire u1__abc_73140_new_n449_; 
wire u1__abc_73140_new_n450_; 
wire u1__abc_73140_new_n451_; 
wire u1__abc_73140_new_n453_; 
wire u1__abc_73140_new_n454_; 
wire u1__abc_73140_new_n455_; 
wire u1__abc_73140_new_n456_; 
wire u1__abc_73140_new_n457_; 
wire u1__abc_73140_new_n458_; 
wire u1__abc_73140_new_n459_; 
wire u1__abc_73140_new_n460_; 
wire u1__abc_73140_new_n461_; 
wire u1__abc_73140_new_n462_; 
wire u1__abc_73140_new_n464_; 
wire u1__abc_73140_new_n465_; 
wire u1__abc_73140_new_n466_; 
wire u1__abc_73140_new_n467_; 
wire u1__abc_73140_new_n468_; 
wire u1__abc_73140_new_n469_; 
wire u1__abc_73140_new_n470_; 
wire u1__abc_73140_new_n471_; 
wire u1__abc_73140_new_n472_; 
wire u1__abc_73140_new_n473_; 
wire u1__abc_73140_new_n474_; 
wire u1__abc_73140_new_n475_; 
wire u1__abc_73140_new_n476_; 
wire u1__abc_73140_new_n477_; 
wire u1__abc_73140_new_n478_; 
wire u1__abc_73140_new_n480_; 
wire u1__abc_73140_new_n481_; 
wire u1__abc_73140_new_n482_; 
wire u1__abc_73140_new_n483_; 
wire u1__abc_73140_new_n484_; 
wire u1__abc_73140_new_n485_; 
wire u1__abc_73140_new_n486_; 
wire u1__abc_73140_new_n487_; 
wire u1__abc_73140_new_n488_; 
wire u1__abc_73140_new_n489_; 
wire u1__abc_73140_new_n490_; 
wire u1__abc_73140_new_n491_; 
wire u1__abc_73140_new_n492_; 
wire u1__abc_73140_new_n493_; 
wire u1__abc_73140_new_n494_; 
wire u1__abc_73140_new_n495_; 
wire u1__abc_73140_new_n496_; 
wire u1__abc_73140_new_n498_; 
wire u1__abc_73140_new_n499_; 
wire u1__abc_73140_new_n500_; 
wire u1__abc_73140_new_n501_; 
wire u1__abc_73140_new_n502_; 
wire u1__abc_73140_new_n503_; 
wire u1__abc_73140_new_n504_; 
wire u1__abc_73140_new_n505_; 
wire u1__abc_73140_new_n506_; 
wire u1__abc_73140_new_n507_; 
wire u1__abc_73140_new_n508_; 
wire u1__abc_73140_new_n509_; 
wire u1__abc_73140_new_n511_; 
wire u1__abc_73140_new_n512_; 
wire u1__abc_73140_new_n513_; 
wire u1__abc_73140_new_n514_; 
wire u1__abc_73140_new_n515_; 
wire u1__abc_73140_new_n516_; 
wire u1__abc_73140_new_n517_; 
wire u1__abc_73140_new_n518_; 
wire u1__abc_73140_new_n519_; 
wire u1__abc_73140_new_n520_; 
wire u1__abc_73140_new_n521_; 
wire u1__abc_73140_new_n522_; 
wire u1__abc_73140_new_n524_; 
wire u1__abc_73140_new_n525_; 
wire u1__abc_73140_new_n526_; 
wire u1__abc_73140_new_n527_; 
wire u1__abc_73140_new_n528_; 
wire u1__abc_73140_new_n529_; 
wire u1__abc_73140_new_n530_; 
wire u1__abc_73140_new_n532_; 
wire u1__abc_73140_new_n533_; 
wire u1__abc_73140_new_n535_; 
wire u1__abc_73140_new_n536_; 
wire u1__abc_73140_new_n538_; 
wire u1__abc_73140_new_n539_; 
wire u1__abc_73140_new_n541_; 
wire u1__abc_73140_new_n542_; 
wire u1__abc_73140_new_n544_; 
wire u1__abc_73140_new_n545_; 
wire u1__abc_73140_new_n547_; 
wire u1__abc_73140_new_n548_; 
wire u1__abc_73140_new_n550_; 
wire u1__abc_73140_new_n551_; 
wire u1__abc_73140_new_n553_; 
wire u1__abc_73140_new_n554_; 
wire u1__abc_73140_new_n555_; 
wire u1__abc_73140_new_n557_; 
wire u1__abc_73140_new_n558_; 
wire u1__abc_73140_new_n559_; 
wire u1__abc_73140_new_n561_; 
wire u1__abc_73140_new_n561__bF_buf0; 
wire u1__abc_73140_new_n561__bF_buf1; 
wire u1__abc_73140_new_n561__bF_buf2; 
wire u1__abc_73140_new_n561__bF_buf3; 
wire u1__abc_73140_new_n561__bF_buf4; 
wire u1__abc_73140_new_n562_; 
wire u1__abc_73140_new_n563_; 
wire u1__abc_73140_new_n563__bF_buf0; 
wire u1__abc_73140_new_n563__bF_buf1; 
wire u1__abc_73140_new_n563__bF_buf2; 
wire u1__abc_73140_new_n563__bF_buf3; 
wire u1__abc_73140_new_n564_; 
wire u1__abc_73140_new_n565_; 
wire u1__abc_73140_new_n566_; 
wire u1__abc_73140_new_n567_; 
wire u1__abc_73140_new_n567__bF_buf0; 
wire u1__abc_73140_new_n567__bF_buf1; 
wire u1__abc_73140_new_n567__bF_buf2; 
wire u1__abc_73140_new_n567__bF_buf3; 
wire u1__abc_73140_new_n568_; 
wire u1__abc_73140_new_n569_; 
wire u1__abc_73140_new_n570_; 
wire u1__abc_73140_new_n570__bF_buf0; 
wire u1__abc_73140_new_n570__bF_buf1; 
wire u1__abc_73140_new_n570__bF_buf2; 
wire u1__abc_73140_new_n570__bF_buf3; 
wire u1__abc_73140_new_n571_; 
wire u1__abc_73140_new_n572_; 
wire u1__abc_73140_new_n573_; 
wire u1__abc_73140_new_n574_; 
wire u1__abc_73140_new_n576_; 
wire u1__abc_73140_new_n577_; 
wire u1__abc_73140_new_n578_; 
wire u1__abc_73140_new_n579_; 
wire u1__abc_73140_new_n580_; 
wire u1__abc_73140_new_n581_; 
wire u1__abc_73140_new_n582_; 
wire u1__abc_73140_new_n583_; 
wire u1__abc_73140_new_n584_; 
wire u1__abc_73140_new_n585_; 
wire u1__abc_73140_new_n587_; 
wire u1__abc_73140_new_n588_; 
wire u1__abc_73140_new_n589_; 
wire u1__abc_73140_new_n590_; 
wire u1__abc_73140_new_n591_; 
wire u1__abc_73140_new_n592_; 
wire u1__abc_73140_new_n593_; 
wire u1__abc_73140_new_n594_; 
wire u1__abc_73140_new_n595_; 
wire u1__abc_73140_new_n596_; 
wire u1__abc_73140_new_n598_; 
wire u1__abc_73140_new_n599_; 
wire u1__abc_73140_new_n600_; 
wire u1__abc_73140_new_n601_; 
wire u1__abc_73140_new_n602_; 
wire u1__abc_73140_new_n603_; 
wire u1__abc_73140_new_n604_; 
wire u1__abc_73140_new_n605_; 
wire u1__abc_73140_new_n606_; 
wire u1__abc_73140_new_n607_; 
wire u1__abc_73140_new_n609_; 
wire u1__abc_73140_new_n610_; 
wire u1__abc_73140_new_n611_; 
wire u1__abc_73140_new_n612_; 
wire u1__abc_73140_new_n613_; 
wire u1__abc_73140_new_n614_; 
wire u1__abc_73140_new_n615_; 
wire u1__abc_73140_new_n616_; 
wire u1__abc_73140_new_n617_; 
wire u1__abc_73140_new_n618_; 
wire u1__abc_73140_new_n620_; 
wire u1__abc_73140_new_n621_; 
wire u1__abc_73140_new_n622_; 
wire u1__abc_73140_new_n623_; 
wire u1__abc_73140_new_n624_; 
wire u1__abc_73140_new_n625_; 
wire u1__abc_73140_new_n626_; 
wire u1__abc_73140_new_n627_; 
wire u1__abc_73140_new_n628_; 
wire u1__abc_73140_new_n629_; 
wire u1__abc_73140_new_n631_; 
wire u1__abc_73140_new_n632_; 
wire u1__abc_73140_new_n633_; 
wire u1__abc_73140_new_n634_; 
wire u1__abc_73140_new_n635_; 
wire u1__abc_73140_new_n636_; 
wire u1__abc_73140_new_n637_; 
wire u1__abc_73140_new_n638_; 
wire u1__abc_73140_new_n639_; 
wire u1__abc_73140_new_n640_; 
wire u1__abc_73140_new_n642_; 
wire u1__abc_73140_new_n643_; 
wire u1__abc_73140_new_n644_; 
wire u1__abc_73140_new_n645_; 
wire u1__abc_73140_new_n646_; 
wire u1__abc_73140_new_n647_; 
wire u1__abc_73140_new_n648_; 
wire u1__abc_73140_new_n649_; 
wire u1__abc_73140_new_n650_; 
wire u1__abc_73140_new_n651_; 
wire u1__abc_73140_new_n653_; 
wire u1__abc_73140_new_n654_; 
wire u1__abc_73140_new_n655_; 
wire u1__abc_73140_new_n656_; 
wire u1__abc_73140_new_n657_; 
wire u1__abc_73140_new_n658_; 
wire u1__abc_73140_new_n659_; 
wire u1__abc_73140_new_n660_; 
wire u1__abc_73140_new_n661_; 
wire u1__abc_73140_new_n662_; 
wire u1__abc_73140_new_n664_; 
wire u1__abc_73140_new_n665_; 
wire u1__abc_73140_new_n666_; 
wire u1__abc_73140_new_n667_; 
wire u1__abc_73140_new_n668_; 
wire u1__abc_73140_new_n669_; 
wire u1__abc_73140_new_n670_; 
wire u1__abc_73140_new_n671_; 
wire u1__abc_73140_new_n672_; 
wire u1__abc_73140_new_n673_; 
wire u1__abc_73140_new_n675_; 
wire u1__abc_73140_new_n676_; 
wire u1__abc_73140_new_n677_; 
wire u1__abc_73140_new_n678_; 
wire u1__abc_73140_new_n679_; 
wire u1__abc_73140_new_n680_; 
wire u1__abc_73140_new_n681_; 
wire u1__abc_73140_new_n682_; 
wire u1__abc_73140_new_n683_; 
wire u1__abc_73140_new_n684_; 
wire u1__abc_73140_new_n686_; 
wire u1__abc_73140_new_n687_; 
wire u1__abc_73140_new_n688_; 
wire u1__abc_73140_new_n689_; 
wire u1__abc_73140_new_n690_; 
wire u1__abc_73140_new_n691_; 
wire u1__abc_73140_new_n692_; 
wire u1__abc_73140_new_n693_; 
wire u1__abc_73140_new_n694_; 
wire u1__abc_73140_new_n695_; 
wire u1__abc_73140_new_n697_; 
wire u1__abc_73140_new_n698_; 
wire u1__abc_73140_new_n699_; 
wire u1__abc_73140_new_n700_; 
wire u1__abc_73140_new_n701_; 
wire u1__abc_73140_new_n702_; 
wire u1__abc_73140_new_n703_; 
wire u1__abc_73140_new_n704_; 
wire u1__abc_73140_new_n705_; 
wire u1__abc_73140_new_n706_; 
wire u1__abc_73140_new_n708_; 
wire u1__abc_73140_new_n709_; 
wire u1__abc_73140_new_n710_; 
wire u1__abc_73140_new_n711_; 
wire u1__abc_73140_new_n712_; 
wire u1__abc_73140_new_n713_; 
wire u1__abc_73140_new_n714_; 
wire u1__abc_73140_new_n715_; 
wire u1__abc_73140_new_n716_; 
wire u1__abc_73140_new_n717_; 
wire u1__abc_73140_new_n719_; 
wire u1__abc_73140_new_n720_; 
wire u1__abc_73140_new_n721_; 
wire u1__abc_73140_new_n722_; 
wire u1__abc_73140_new_n723_; 
wire u1__abc_73140_new_n724_; 
wire u1__abc_73140_new_n725_; 
wire u1__abc_73140_new_n726_; 
wire u1__abc_73140_new_n727_; 
wire u1__abc_73140_new_n728_; 
wire u1__abc_73140_new_n730_; 
wire u1__abc_73140_new_n731_; 
wire u1__abc_73140_new_n732_; 
wire u1__abc_73140_new_n733_; 
wire u1__abc_73140_new_n734_; 
wire u1__abc_73140_new_n735_; 
wire u1__abc_73140_new_n736_; 
wire u1__abc_73140_new_n737_; 
wire u1__abc_73140_new_n738_; 
wire u1__abc_73140_new_n739_; 
wire u1__abc_73140_new_n741_; 
wire u1__abc_73140_new_n742_; 
wire u1__abc_73140_new_n743_; 
wire u1__abc_73140_new_n744_; 
wire u1__abc_73140_new_n745_; 
wire u1__abc_73140_new_n746_; 
wire u1__abc_73140_new_n747_; 
wire u1__abc_73140_new_n748_; 
wire u1__abc_73140_new_n749_; 
wire u1__abc_73140_new_n750_; 
wire u1__abc_73140_new_n752_; 
wire u1__abc_73140_new_n753_; 
wire u1__abc_73140_new_n754_; 
wire u1__abc_73140_new_n755_; 
wire u1__abc_73140_new_n756_; 
wire u1__abc_73140_new_n757_; 
wire u1__abc_73140_new_n758_; 
wire u1__abc_73140_new_n759_; 
wire u1__abc_73140_new_n760_; 
wire u1__abc_73140_new_n761_; 
wire u1__abc_73140_new_n763_; 
wire u1__abc_73140_new_n764_; 
wire u1__abc_73140_new_n765_; 
wire u1__abc_73140_new_n766_; 
wire u1__abc_73140_new_n767_; 
wire u1__abc_73140_new_n768_; 
wire u1__abc_73140_new_n769_; 
wire u1__abc_73140_new_n770_; 
wire u1__abc_73140_new_n771_; 
wire u1__abc_73140_new_n772_; 
wire u1__abc_73140_new_n774_; 
wire u1__abc_73140_new_n775_; 
wire u1__abc_73140_new_n776_; 
wire u1__abc_73140_new_n777_; 
wire u1__abc_73140_new_n778_; 
wire u1__abc_73140_new_n779_; 
wire u1__abc_73140_new_n780_; 
wire u1__abc_73140_new_n781_; 
wire u1__abc_73140_new_n782_; 
wire u1__abc_73140_new_n784_; 
wire u1__abc_73140_new_n785_; 
wire u1__abc_73140_new_n786_; 
wire u1__abc_73140_new_n787_; 
wire u1__abc_73140_new_n788_; 
wire u1__abc_73140_new_n789_; 
wire u1__abc_73140_new_n790_; 
wire u1__abc_73140_new_n791_; 
wire u1__abc_73140_new_n792_; 
wire u1__abc_73140_new_n794_; 
wire u1__abc_73140_new_n795_; 
wire u1__abc_73140_new_n796_; 
wire u1__abc_73140_new_n797_; 
wire u1__abc_73140_new_n798_; 
wire u1__abc_73140_new_n799_; 
wire u1__abc_73140_new_n800_; 
wire u1__abc_73140_new_n801_; 
wire u1__abc_73140_new_n802_; 
wire u1__abc_73140_new_n803_; 
wire u1__abc_73140_new_n805_; 
wire u1__abc_73140_new_n806_; 
wire u1__abc_73140_new_n807_; 
wire u1__abc_73140_new_n808_; 
wire u1__abc_73140_new_n809_; 
wire u1__abc_73140_new_n810_; 
wire u1__abc_73140_new_n811_; 
wire u1__abc_73140_new_n812_; 
wire u1__abc_73140_new_n814_; 
wire u1__abc_73140_new_n815_; 
wire u1__abc_73140_new_n816_; 
wire u1__abc_73140_new_n817_; 
wire u1__abc_73140_new_n818_; 
wire u1__abc_73140_new_n819_; 
wire u1__abc_73140_new_n820_; 
wire u1__abc_73140_new_n821_; 
wire u1__abc_73140_new_n822_; 
wire u1__abc_73140_new_n823_; 
wire u1__abc_73140_new_n825_; 
wire u1__abc_73140_new_n826_; 
wire u1__abc_73140_new_n826__bF_buf0; 
wire u1__abc_73140_new_n826__bF_buf1; 
wire u1__abc_73140_new_n826__bF_buf2; 
wire u1__abc_73140_new_n826__bF_buf3; 
wire u1__abc_73140_new_n827_; 
wire u1__abc_73140_new_n829_; 
wire u1__abc_73140_new_n830_; 
wire u1__abc_73140_new_n832_; 
wire u1__abc_73140_new_n833_; 
wire u1__abc_73140_new_n835_; 
wire u1__abc_73140_new_n836_; 
wire u1__abc_73140_new_n838_; 
wire u1__abc_73140_new_n839_; 
wire u1__abc_73140_new_n841_; 
wire u1__abc_73140_new_n842_; 
wire u1__abc_73140_new_n844_; 
wire u1__abc_73140_new_n845_; 
wire u1__abc_73140_new_n847_; 
wire u1__abc_73140_new_n848_; 
wire u1__abc_73140_new_n850_; 
wire u1__abc_73140_new_n851_; 
wire u1__abc_73140_new_n853_; 
wire u1__abc_73140_new_n854_; 
wire u1__abc_73140_new_n856_; 
wire u1__abc_73140_new_n857_; 
wire u1__abc_73140_new_n859_; 
wire u1__abc_73140_new_n860_; 
wire u1__abc_73140_new_n862_; 
wire u1__abc_73140_new_n863_; 
wire u1__abc_73140_new_n865_; 
wire u1__abc_73140_new_n866_; 
wire u1__abc_73140_new_n868_; 
wire u1__abc_73140_new_n869_; 
wire u1__abc_73140_new_n871_; 
wire u1__abc_73140_new_n872_; 
wire u1__abc_73140_new_n874_; 
wire u1__abc_73140_new_n875_; 
wire u1__abc_73140_new_n877_; 
wire u1__abc_73140_new_n878_; 
wire u1__abc_73140_new_n880_; 
wire u1__abc_73140_new_n881_; 
wire u1__abc_73140_new_n883_; 
wire u1__abc_73140_new_n884_; 
wire u1__abc_73140_new_n886_; 
wire u1__abc_73140_new_n887_; 
wire u1__abc_73140_new_n889_; 
wire u1__abc_73140_new_n890_; 
wire u1__abc_73140_new_n892_; 
wire u1__abc_73140_new_n893_; 
wire u1__abc_73140_new_n895_; 
wire u1__abc_73140_new_n896_; 
wire u1__abc_73140_new_n898_; 
wire u1__abc_73140_new_n899_; 
wire u1__abc_73140_new_n900_; 
wire u1__abc_73140_new_n900__bF_buf0; 
wire u1__abc_73140_new_n900__bF_buf1; 
wire u1__abc_73140_new_n900__bF_buf2; 
wire u1__abc_73140_new_n900__bF_buf3; 
wire u1__abc_73140_new_n900__bF_buf4; 
wire u1__abc_73140_new_n901_; 
wire u1__abc_73140_new_n902_; 
wire u1__abc_73140_new_n903_; 
wire u1__abc_73140_new_n904_; 
wire u1__abc_73140_new_n904__bF_buf0; 
wire u1__abc_73140_new_n904__bF_buf1; 
wire u1__abc_73140_new_n904__bF_buf2; 
wire u1__abc_73140_new_n904__bF_buf3; 
wire u1__abc_73140_new_n904__bF_buf4; 
wire u1__abc_73140_new_n905_; 
wire u1__abc_73140_new_n906_; 
wire u1__abc_73140_new_n906__bF_buf0; 
wire u1__abc_73140_new_n906__bF_buf1; 
wire u1__abc_73140_new_n906__bF_buf2; 
wire u1__abc_73140_new_n906__bF_buf3; 
wire u1__abc_73140_new_n907_; 
wire u1__abc_73140_new_n908_; 
wire u1__abc_73140_new_n909_; 
wire u1__abc_73140_new_n910_; 
wire u1__abc_73140_new_n911_; 
wire u1__abc_73140_new_n912_; 
wire u1__abc_73140_new_n912__bF_buf0; 
wire u1__abc_73140_new_n912__bF_buf1; 
wire u1__abc_73140_new_n912__bF_buf2; 
wire u1__abc_73140_new_n912__bF_buf3; 
wire u1__abc_73140_new_n913_; 
wire u1__abc_73140_new_n914_; 
wire u1__abc_73140_new_n915_; 
wire u1__abc_73140_new_n916_; 
wire u1__abc_73140_new_n917_; 
wire u1__abc_73140_new_n918_; 
wire u1__abc_73140_new_n919_; 
wire u1__abc_73140_new_n920_; 
wire u1__abc_73140_new_n921_; 
wire u1__abc_73140_new_n922_; 
wire u1__abc_73140_new_n923_; 
wire u1__abc_73140_new_n924_; 
wire u1__abc_73140_new_n925_; 
wire u1__abc_73140_new_n926_; 
wire u1__abc_73140_new_n927_; 
wire u1__abc_73140_new_n929_; 
wire u1__abc_73140_new_n930_; 
wire u1__abc_73140_new_n931_; 
wire u1__abc_73140_new_n932_; 
wire u1__abc_73140_new_n933_; 
wire u1__abc_73140_new_n934_; 
wire u1__abc_73140_new_n935_; 
wire u1__abc_73140_new_n936_; 
wire u1__abc_73140_new_n937_; 
wire u1__abc_73140_new_n938_; 
wire u1__abc_73140_new_n939_; 
wire u1__abc_73140_new_n940_; 
wire u1__abc_73140_new_n941_; 
wire u1__abc_73140_new_n942_; 
wire u1__abc_73140_new_n944_; 
wire u1__abc_73140_new_n945_; 
wire u1__abc_73140_new_n946_; 
wire u1__abc_73140_new_n947_; 
wire u1__abc_73140_new_n948_; 
wire u1__abc_73140_new_n949_; 
wire u1__abc_73140_new_n950_; 
wire u1__abc_73140_new_n951_; 
wire u1__abc_73140_new_n952_; 
wire u1__abc_73140_new_n953_; 
wire u1__abc_73140_new_n954_; 
wire u1__abc_73140_new_n955_; 
wire u1__abc_73140_new_n956_; 
wire u1__abc_73140_new_n957_; 
wire u1__abc_73140_new_n959_; 
wire u1__abc_73140_new_n960_; 
wire u1__abc_73140_new_n961_; 
wire u1__abc_73140_new_n962_; 
wire u1__abc_73140_new_n963_; 
wire u1__abc_73140_new_n964_; 
wire u1__abc_73140_new_n965_; 
wire u1__abc_73140_new_n966_; 
wire u1__abc_73140_new_n967_; 
wire u1__abc_73140_new_n968_; 
wire u1__abc_73140_new_n969_; 
wire u1__abc_73140_new_n970_; 
wire u1__abc_73140_new_n971_; 
wire u1__abc_73140_new_n972_; 
wire u1__abc_73140_new_n974_; 
wire u1__abc_73140_new_n975_; 
wire u1__abc_73140_new_n976_; 
wire u1__abc_73140_new_n977_; 
wire u1__abc_73140_new_n978_; 
wire u1__abc_73140_new_n979_; 
wire u1__abc_73140_new_n980_; 
wire u1__abc_73140_new_n981_; 
wire u1__abc_73140_new_n982_; 
wire u1__abc_73140_new_n983_; 
wire u1__abc_73140_new_n984_; 
wire u1__abc_73140_new_n985_; 
wire u1__abc_73140_new_n986_; 
wire u1__abc_73140_new_n987_; 
wire u1__abc_73140_new_n989_; 
wire u1__abc_73140_new_n990_; 
wire u1__abc_73140_new_n991_; 
wire u1__abc_73140_new_n992_; 
wire u1__abc_73140_new_n993_; 
wire u1__abc_73140_new_n994_; 
wire u1__abc_73140_new_n995_; 
wire u1__abc_73140_new_n996_; 
wire u1__abc_73140_new_n997_; 
wire u1__abc_73140_new_n998_; 
wire u1__abc_73140_new_n999_; 
wire u1_acs_addr_0_; 
wire u1_acs_addr_10_; 
wire u1_acs_addr_11_; 
wire u1_acs_addr_12_; 
wire u1_acs_addr_13_; 
wire u1_acs_addr_14_; 
wire u1_acs_addr_15_; 
wire u1_acs_addr_16_; 
wire u1_acs_addr_17_; 
wire u1_acs_addr_18_; 
wire u1_acs_addr_19_; 
wire u1_acs_addr_1_; 
wire u1_acs_addr_20_; 
wire u1_acs_addr_21_; 
wire u1_acs_addr_22_; 
wire u1_acs_addr_23_; 
wire u1_acs_addr_2_; 
wire u1_acs_addr_3_; 
wire u1_acs_addr_4_; 
wire u1_acs_addr_5_; 
wire u1_acs_addr_6_; 
wire u1_acs_addr_7_; 
wire u1_acs_addr_8_; 
wire u1_acs_addr_9_; 
wire u1_acs_addr_pl1_0_; 
wire u1_acs_addr_pl1_10_; 
wire u1_acs_addr_pl1_11_; 
wire u1_acs_addr_pl1_12_; 
wire u1_acs_addr_pl1_13_; 
wire u1_acs_addr_pl1_14_; 
wire u1_acs_addr_pl1_15_; 
wire u1_acs_addr_pl1_16_; 
wire u1_acs_addr_pl1_17_; 
wire u1_acs_addr_pl1_18_; 
wire u1_acs_addr_pl1_19_; 
wire u1_acs_addr_pl1_1_; 
wire u1_acs_addr_pl1_20_; 
wire u1_acs_addr_pl1_21_; 
wire u1_acs_addr_pl1_22_; 
wire u1_acs_addr_pl1_23_; 
wire u1_acs_addr_pl1_2_; 
wire u1_acs_addr_pl1_3_; 
wire u1_acs_addr_pl1_4_; 
wire u1_acs_addr_pl1_5_; 
wire u1_acs_addr_pl1_6_; 
wire u1_acs_addr_pl1_7_; 
wire u1_acs_addr_pl1_8_; 
wire u1_acs_addr_pl1_9_; 
wire u1_bas; 
wire u1_bas_bF_buf0; 
wire u1_bas_bF_buf1; 
wire u1_bas_bF_buf2; 
wire u1_bas_bF_buf3; 
wire u1_col_adr_0_; 
wire u1_col_adr_1_; 
wire u1_col_adr_2_; 
wire u1_col_adr_3_; 
wire u1_col_adr_4_; 
wire u1_col_adr_5_; 
wire u1_col_adr_6_; 
wire u1_col_adr_7_; 
wire u1_col_adr_8_; 
wire u1_col_adr_9_; 
wire u1_sram_addr_0_; 
wire u1_sram_addr_10_; 
wire u1_sram_addr_11_; 
wire u1_sram_addr_12_; 
wire u1_sram_addr_13_; 
wire u1_sram_addr_14_; 
wire u1_sram_addr_15_; 
wire u1_sram_addr_16_; 
wire u1_sram_addr_17_; 
wire u1_sram_addr_18_; 
wire u1_sram_addr_19_; 
wire u1_sram_addr_1_; 
wire u1_sram_addr_20_; 
wire u1_sram_addr_21_; 
wire u1_sram_addr_22_; 
wire u1_sram_addr_23_; 
wire u1_sram_addr_2_; 
wire u1_sram_addr_3_; 
wire u1_sram_addr_4_; 
wire u1_sram_addr_5_; 
wire u1_sram_addr_6_; 
wire u1_sram_addr_7_; 
wire u1_sram_addr_8_; 
wire u1_sram_addr_9_; 
wire u1_u0__0out_r_12_0__0_; 
wire u1_u0__0out_r_12_0__10_; 
wire u1_u0__0out_r_12_0__11_; 
wire u1_u0__0out_r_12_0__12_; 
wire u1_u0__0out_r_12_0__1_; 
wire u1_u0__0out_r_12_0__2_; 
wire u1_u0__0out_r_12_0__3_; 
wire u1_u0__0out_r_12_0__4_; 
wire u1_u0__0out_r_12_0__5_; 
wire u1_u0__0out_r_12_0__6_; 
wire u1_u0__0out_r_12_0__7_; 
wire u1_u0__0out_r_12_0__8_; 
wire u1_u0__0out_r_12_0__9_; 
wire u1_u0__abc_73035_new_n102_; 
wire u1_u0__abc_73035_new_n103_; 
wire u1_u0__abc_73035_new_n104_; 
wire u1_u0__abc_73035_new_n105_; 
wire u1_u0__abc_73035_new_n107_; 
wire u1_u0__abc_73035_new_n108_; 
wire u1_u0__abc_73035_new_n109_; 
wire u1_u0__abc_73035_new_n111_; 
wire u1_u0__abc_73035_new_n112_; 
wire u1_u0__abc_73035_new_n113_; 
wire u1_u0__abc_73035_new_n114_; 
wire u1_u0__abc_73035_new_n116_; 
wire u1_u0__abc_73035_new_n117_; 
wire u1_u0__abc_73035_new_n118_; 
wire u1_u0__abc_73035_new_n120_; 
wire u1_u0__abc_73035_new_n121_; 
wire u1_u0__abc_73035_new_n122_; 
wire u1_u0__abc_73035_new_n123_; 
wire u1_u0__abc_73035_new_n125_; 
wire u1_u0__abc_73035_new_n126_; 
wire u1_u0__abc_73035_new_n127_; 
wire u1_u0__abc_73035_new_n129_; 
wire u1_u0__abc_73035_new_n130_; 
wire u1_u0__abc_73035_new_n131_; 
wire u1_u0__abc_73035_new_n132_; 
wire u1_u0__abc_73035_new_n133_; 
wire u1_u0__abc_73035_new_n135_; 
wire u1_u0__abc_73035_new_n136_; 
wire u1_u0__abc_73035_new_n137_; 
wire u1_u0__abc_73035_new_n139_; 
wire u1_u0__abc_73035_new_n140_; 
wire u1_u0__abc_73035_new_n141_; 
wire u1_u0__abc_73035_new_n142_; 
wire u1_u0__abc_73035_new_n144_; 
wire u1_u0__abc_73035_new_n145_; 
wire u1_u0__abc_73035_new_n146_; 
wire u1_u0__abc_73035_new_n148_; 
wire u1_u0__abc_73035_new_n149_; 
wire u1_u0__abc_73035_new_n150_; 
wire u1_u0__abc_73035_new_n152_; 
wire u1_u0__abc_73035_new_n153_; 
wire u1_u0__abc_73035_new_n51_; 
wire u1_u0__abc_73035_new_n52_; 
wire u1_u0__abc_73035_new_n53_; 
wire u1_u0__abc_73035_new_n55_; 
wire u1_u0__abc_73035_new_n56_; 
wire u1_u0__abc_73035_new_n57_; 
wire u1_u0__abc_73035_new_n59_; 
wire u1_u0__abc_73035_new_n60_; 
wire u1_u0__abc_73035_new_n61_; 
wire u1_u0__abc_73035_new_n63_; 
wire u1_u0__abc_73035_new_n64_; 
wire u1_u0__abc_73035_new_n65_; 
wire u1_u0__abc_73035_new_n67_; 
wire u1_u0__abc_73035_new_n68_; 
wire u1_u0__abc_73035_new_n69_; 
wire u1_u0__abc_73035_new_n70_; 
wire u1_u0__abc_73035_new_n72_; 
wire u1_u0__abc_73035_new_n73_; 
wire u1_u0__abc_73035_new_n74_; 
wire u1_u0__abc_73035_new_n76_; 
wire u1_u0__abc_73035_new_n77_; 
wire u1_u0__abc_73035_new_n78_; 
wire u1_u0__abc_73035_new_n79_; 
wire u1_u0__abc_73035_new_n80_; 
wire u1_u0__abc_73035_new_n82_; 
wire u1_u0__abc_73035_new_n83_; 
wire u1_u0__abc_73035_new_n84_; 
wire u1_u0__abc_73035_new_n86_; 
wire u1_u0__abc_73035_new_n87_; 
wire u1_u0__abc_73035_new_n88_; 
wire u1_u0__abc_73035_new_n89_; 
wire u1_u0__abc_73035_new_n91_; 
wire u1_u0__abc_73035_new_n92_; 
wire u1_u0__abc_73035_new_n93_; 
wire u1_u0__abc_73035_new_n95_; 
wire u1_u0__abc_73035_new_n96_; 
wire u1_u0__abc_73035_new_n98_; 
wire u1_u0__abc_73035_new_n99_; 
wire u1_u0_inc_next; 
wire u1_wb_write_go; 
wire u1_wr_cycle; 
wire u1_wr_hold; 
wire u2__0bank_open_0_0_; 
wire u2__0row_same_0_0_; 
wire u2__abc_75448_new_n100_; 
wire u2__abc_75448_new_n101_; 
wire u2__abc_75448_new_n102_; 
wire u2__abc_75448_new_n103_; 
wire u2__abc_75448_new_n104_; 
wire u2__abc_75448_new_n105_; 
wire u2__abc_75448_new_n106_; 
wire u2__abc_75448_new_n107_; 
wire u2__abc_75448_new_n108_; 
wire u2__abc_75448_new_n109_; 
wire u2__abc_75448_new_n111_; 
wire u2__abc_75448_new_n112_; 
wire u2__abc_75448_new_n113_; 
wire u2__abc_75448_new_n114_; 
wire u2__abc_75448_new_n115_; 
wire u2__abc_75448_new_n116_; 
wire u2__abc_75448_new_n117_; 
wire u2__abc_75448_new_n118_; 
wire u2__abc_75448_new_n119_; 
wire u2__abc_75448_new_n120_; 
wire u2__abc_75448_new_n121_; 
wire u2__abc_75448_new_n122_; 
wire u2__abc_75448_new_n123_; 
wire u2__abc_75448_new_n124_; 
wire u2__abc_75448_new_n80_; 
wire u2__abc_75448_new_n82_; 
wire u2__abc_75448_new_n96_; 
wire u2__abc_75448_new_n97_; 
wire u2__abc_75448_new_n98_; 
wire u2__abc_75448_new_n99_; 
wire u2_bank_clr_0; 
wire u2_bank_clr_1; 
wire u2_bank_clr_all_0; 
wire u2_bank_clr_all_1; 
wire u2_bank_open_0; 
wire u2_bank_open_1; 
wire u2_bank_set_0; 
wire u2_bank_set_1; 
wire u2_row_same_0; 
wire u2_row_same_1; 
wire u2_u0__0b0_last_row_12_0__0_; 
wire u2_u0__0b0_last_row_12_0__10_; 
wire u2_u0__0b0_last_row_12_0__11_; 
wire u2_u0__0b0_last_row_12_0__12_; 
wire u2_u0__0b0_last_row_12_0__1_; 
wire u2_u0__0b0_last_row_12_0__2_; 
wire u2_u0__0b0_last_row_12_0__3_; 
wire u2_u0__0b0_last_row_12_0__4_; 
wire u2_u0__0b0_last_row_12_0__5_; 
wire u2_u0__0b0_last_row_12_0__6_; 
wire u2_u0__0b0_last_row_12_0__7_; 
wire u2_u0__0b0_last_row_12_0__8_; 
wire u2_u0__0b0_last_row_12_0__9_; 
wire u2_u0__0b1_last_row_12_0__0_; 
wire u2_u0__0b1_last_row_12_0__10_; 
wire u2_u0__0b1_last_row_12_0__11_; 
wire u2_u0__0b1_last_row_12_0__12_; 
wire u2_u0__0b1_last_row_12_0__1_; 
wire u2_u0__0b1_last_row_12_0__2_; 
wire u2_u0__0b1_last_row_12_0__3_; 
wire u2_u0__0b1_last_row_12_0__4_; 
wire u2_u0__0b1_last_row_12_0__5_; 
wire u2_u0__0b1_last_row_12_0__6_; 
wire u2_u0__0b1_last_row_12_0__7_; 
wire u2_u0__0b1_last_row_12_0__8_; 
wire u2_u0__0b1_last_row_12_0__9_; 
wire u2_u0__0b2_last_row_12_0__0_; 
wire u2_u0__0b2_last_row_12_0__10_; 
wire u2_u0__0b2_last_row_12_0__11_; 
wire u2_u0__0b2_last_row_12_0__12_; 
wire u2_u0__0b2_last_row_12_0__1_; 
wire u2_u0__0b2_last_row_12_0__2_; 
wire u2_u0__0b2_last_row_12_0__3_; 
wire u2_u0__0b2_last_row_12_0__4_; 
wire u2_u0__0b2_last_row_12_0__5_; 
wire u2_u0__0b2_last_row_12_0__6_; 
wire u2_u0__0b2_last_row_12_0__7_; 
wire u2_u0__0b2_last_row_12_0__8_; 
wire u2_u0__0b2_last_row_12_0__9_; 
wire u2_u0__0b3_last_row_12_0__0_; 
wire u2_u0__0b3_last_row_12_0__10_; 
wire u2_u0__0b3_last_row_12_0__11_; 
wire u2_u0__0b3_last_row_12_0__12_; 
wire u2_u0__0b3_last_row_12_0__1_; 
wire u2_u0__0b3_last_row_12_0__2_; 
wire u2_u0__0b3_last_row_12_0__3_; 
wire u2_u0__0b3_last_row_12_0__4_; 
wire u2_u0__0b3_last_row_12_0__5_; 
wire u2_u0__0b3_last_row_12_0__6_; 
wire u2_u0__0b3_last_row_12_0__7_; 
wire u2_u0__0b3_last_row_12_0__8_; 
wire u2_u0__0b3_last_row_12_0__9_; 
wire u2_u0__0bank0_open_0_0_; 
wire u2_u0__0bank1_open_0_0_; 
wire u2_u0__0bank2_open_0_0_; 
wire u2_u0__0bank3_open_0_0_; 
wire u2_u0__abc_74955_auto_rtlil_cc_1942_NotGate_71538; 
wire u2_u0__abc_74955_new_n136_; 
wire u2_u0__abc_74955_new_n137_; 
wire u2_u0__abc_74955_new_n137__bF_buf0; 
wire u2_u0__abc_74955_new_n137__bF_buf1; 
wire u2_u0__abc_74955_new_n137__bF_buf2; 
wire u2_u0__abc_74955_new_n137__bF_buf3; 
wire u2_u0__abc_74955_new_n137__bF_buf4; 
wire u2_u0__abc_74955_new_n138_; 
wire u2_u0__abc_74955_new_n139_; 
wire u2_u0__abc_74955_new_n140_; 
wire u2_u0__abc_74955_new_n141_; 
wire u2_u0__abc_74955_new_n143_; 
wire u2_u0__abc_74955_new_n144_; 
wire u2_u0__abc_74955_new_n145_; 
wire u2_u0__abc_74955_new_n146_; 
wire u2_u0__abc_74955_new_n148_; 
wire u2_u0__abc_74955_new_n149_; 
wire u2_u0__abc_74955_new_n150_; 
wire u2_u0__abc_74955_new_n151_; 
wire u2_u0__abc_74955_new_n153_; 
wire u2_u0__abc_74955_new_n154_; 
wire u2_u0__abc_74955_new_n155_; 
wire u2_u0__abc_74955_new_n156_; 
wire u2_u0__abc_74955_new_n158_; 
wire u2_u0__abc_74955_new_n159_; 
wire u2_u0__abc_74955_new_n160_; 
wire u2_u0__abc_74955_new_n161_; 
wire u2_u0__abc_74955_new_n163_; 
wire u2_u0__abc_74955_new_n164_; 
wire u2_u0__abc_74955_new_n165_; 
wire u2_u0__abc_74955_new_n166_; 
wire u2_u0__abc_74955_new_n168_; 
wire u2_u0__abc_74955_new_n169_; 
wire u2_u0__abc_74955_new_n170_; 
wire u2_u0__abc_74955_new_n171_; 
wire u2_u0__abc_74955_new_n173_; 
wire u2_u0__abc_74955_new_n174_; 
wire u2_u0__abc_74955_new_n175_; 
wire u2_u0__abc_74955_new_n176_; 
wire u2_u0__abc_74955_new_n178_; 
wire u2_u0__abc_74955_new_n179_; 
wire u2_u0__abc_74955_new_n180_; 
wire u2_u0__abc_74955_new_n181_; 
wire u2_u0__abc_74955_new_n183_; 
wire u2_u0__abc_74955_new_n184_; 
wire u2_u0__abc_74955_new_n185_; 
wire u2_u0__abc_74955_new_n186_; 
wire u2_u0__abc_74955_new_n188_; 
wire u2_u0__abc_74955_new_n189_; 
wire u2_u0__abc_74955_new_n190_; 
wire u2_u0__abc_74955_new_n191_; 
wire u2_u0__abc_74955_new_n193_; 
wire u2_u0__abc_74955_new_n194_; 
wire u2_u0__abc_74955_new_n195_; 
wire u2_u0__abc_74955_new_n196_; 
wire u2_u0__abc_74955_new_n198_; 
wire u2_u0__abc_74955_new_n199_; 
wire u2_u0__abc_74955_new_n200_; 
wire u2_u0__abc_74955_new_n201_; 
wire u2_u0__abc_74955_new_n203_; 
wire u2_u0__abc_74955_new_n204_; 
wire u2_u0__abc_74955_new_n205_; 
wire u2_u0__abc_74955_new_n206_; 
wire u2_u0__abc_74955_new_n207_; 
wire u2_u0__abc_74955_new_n208_; 
wire u2_u0__abc_74955_new_n209_; 
wire u2_u0__abc_74955_new_n211_; 
wire u2_u0__abc_74955_new_n212_; 
wire u2_u0__abc_74955_new_n214_; 
wire u2_u0__abc_74955_new_n215_; 
wire u2_u0__abc_74955_new_n217_; 
wire u2_u0__abc_74955_new_n218_; 
wire u2_u0__abc_74955_new_n220_; 
wire u2_u0__abc_74955_new_n221_; 
wire u2_u0__abc_74955_new_n223_; 
wire u2_u0__abc_74955_new_n224_; 
wire u2_u0__abc_74955_new_n226_; 
wire u2_u0__abc_74955_new_n227_; 
wire u2_u0__abc_74955_new_n229_; 
wire u2_u0__abc_74955_new_n230_; 
wire u2_u0__abc_74955_new_n232_; 
wire u2_u0__abc_74955_new_n233_; 
wire u2_u0__abc_74955_new_n235_; 
wire u2_u0__abc_74955_new_n236_; 
wire u2_u0__abc_74955_new_n238_; 
wire u2_u0__abc_74955_new_n239_; 
wire u2_u0__abc_74955_new_n241_; 
wire u2_u0__abc_74955_new_n242_; 
wire u2_u0__abc_74955_new_n244_; 
wire u2_u0__abc_74955_new_n245_; 
wire u2_u0__abc_74955_new_n247_; 
wire u2_u0__abc_74955_new_n248_; 
wire u2_u0__abc_74955_new_n249_; 
wire u2_u0__abc_74955_new_n250_; 
wire u2_u0__abc_74955_new_n251_; 
wire u2_u0__abc_74955_new_n253_; 
wire u2_u0__abc_74955_new_n254_; 
wire u2_u0__abc_74955_new_n256_; 
wire u2_u0__abc_74955_new_n257_; 
wire u2_u0__abc_74955_new_n259_; 
wire u2_u0__abc_74955_new_n260_; 
wire u2_u0__abc_74955_new_n262_; 
wire u2_u0__abc_74955_new_n263_; 
wire u2_u0__abc_74955_new_n265_; 
wire u2_u0__abc_74955_new_n266_; 
wire u2_u0__abc_74955_new_n268_; 
wire u2_u0__abc_74955_new_n269_; 
wire u2_u0__abc_74955_new_n271_; 
wire u2_u0__abc_74955_new_n272_; 
wire u2_u0__abc_74955_new_n274_; 
wire u2_u0__abc_74955_new_n275_; 
wire u2_u0__abc_74955_new_n277_; 
wire u2_u0__abc_74955_new_n278_; 
wire u2_u0__abc_74955_new_n280_; 
wire u2_u0__abc_74955_new_n281_; 
wire u2_u0__abc_74955_new_n283_; 
wire u2_u0__abc_74955_new_n284_; 
wire u2_u0__abc_74955_new_n286_; 
wire u2_u0__abc_74955_new_n287_; 
wire u2_u0__abc_74955_new_n289_; 
wire u2_u0__abc_74955_new_n290_; 
wire u2_u0__abc_74955_new_n291_; 
wire u2_u0__abc_74955_new_n292_; 
wire u2_u0__abc_74955_new_n293_; 
wire u2_u0__abc_74955_new_n295_; 
wire u2_u0__abc_74955_new_n296_; 
wire u2_u0__abc_74955_new_n298_; 
wire u2_u0__abc_74955_new_n299_; 
wire u2_u0__abc_74955_new_n301_; 
wire u2_u0__abc_74955_new_n302_; 
wire u2_u0__abc_74955_new_n304_; 
wire u2_u0__abc_74955_new_n305_; 
wire u2_u0__abc_74955_new_n307_; 
wire u2_u0__abc_74955_new_n308_; 
wire u2_u0__abc_74955_new_n310_; 
wire u2_u0__abc_74955_new_n311_; 
wire u2_u0__abc_74955_new_n313_; 
wire u2_u0__abc_74955_new_n314_; 
wire u2_u0__abc_74955_new_n316_; 
wire u2_u0__abc_74955_new_n317_; 
wire u2_u0__abc_74955_new_n319_; 
wire u2_u0__abc_74955_new_n320_; 
wire u2_u0__abc_74955_new_n322_; 
wire u2_u0__abc_74955_new_n323_; 
wire u2_u0__abc_74955_new_n325_; 
wire u2_u0__abc_74955_new_n326_; 
wire u2_u0__abc_74955_new_n328_; 
wire u2_u0__abc_74955_new_n329_; 
wire u2_u0__abc_74955_new_n331_; 
wire u2_u0__abc_74955_new_n332_; 
wire u2_u0__abc_74955_new_n333_; 
wire u2_u0__abc_74955_new_n334_; 
wire u2_u0__abc_74955_new_n335_; 
wire u2_u0__abc_74955_new_n336_; 
wire u2_u0__abc_74955_new_n337_; 
wire u2_u0__abc_74955_new_n338_; 
wire u2_u0__abc_74955_new_n339_; 
wire u2_u0__abc_74955_new_n340_; 
wire u2_u0__abc_74955_new_n341_; 
wire u2_u0__abc_74955_new_n342_; 
wire u2_u0__abc_74955_new_n343_; 
wire u2_u0__abc_74955_new_n344_; 
wire u2_u0__abc_74955_new_n345_; 
wire u2_u0__abc_74955_new_n346_; 
wire u2_u0__abc_74955_new_n347_; 
wire u2_u0__abc_74955_new_n348_; 
wire u2_u0__abc_74955_new_n349_; 
wire u2_u0__abc_74955_new_n350_; 
wire u2_u0__abc_74955_new_n351_; 
wire u2_u0__abc_74955_new_n352_; 
wire u2_u0__abc_74955_new_n353_; 
wire u2_u0__abc_74955_new_n354_; 
wire u2_u0__abc_74955_new_n355_; 
wire u2_u0__abc_74955_new_n356_; 
wire u2_u0__abc_74955_new_n357_; 
wire u2_u0__abc_74955_new_n358_; 
wire u2_u0__abc_74955_new_n359_; 
wire u2_u0__abc_74955_new_n360_; 
wire u2_u0__abc_74955_new_n361_; 
wire u2_u0__abc_74955_new_n362_; 
wire u2_u0__abc_74955_new_n363_; 
wire u2_u0__abc_74955_new_n364_; 
wire u2_u0__abc_74955_new_n365_; 
wire u2_u0__abc_74955_new_n366_; 
wire u2_u0__abc_74955_new_n367_; 
wire u2_u0__abc_74955_new_n368_; 
wire u2_u0__abc_74955_new_n369_; 
wire u2_u0__abc_74955_new_n370_; 
wire u2_u0__abc_74955_new_n371_; 
wire u2_u0__abc_74955_new_n372_; 
wire u2_u0__abc_74955_new_n373_; 
wire u2_u0__abc_74955_new_n374_; 
wire u2_u0__abc_74955_new_n375_; 
wire u2_u0__abc_74955_new_n376_; 
wire u2_u0__abc_74955_new_n377_; 
wire u2_u0__abc_74955_new_n378_; 
wire u2_u0__abc_74955_new_n379_; 
wire u2_u0__abc_74955_new_n380_; 
wire u2_u0__abc_74955_new_n381_; 
wire u2_u0__abc_74955_new_n382_; 
wire u2_u0__abc_74955_new_n383_; 
wire u2_u0__abc_74955_new_n384_; 
wire u2_u0__abc_74955_new_n385_; 
wire u2_u0__abc_74955_new_n386_; 
wire u2_u0__abc_74955_new_n387_; 
wire u2_u0__abc_74955_new_n388_; 
wire u2_u0__abc_74955_new_n389_; 
wire u2_u0__abc_74955_new_n390_; 
wire u2_u0__abc_74955_new_n391_; 
wire u2_u0__abc_74955_new_n392_; 
wire u2_u0__abc_74955_new_n393_; 
wire u2_u0__abc_74955_new_n394_; 
wire u2_u0__abc_74955_new_n395_; 
wire u2_u0__abc_74955_new_n396_; 
wire u2_u0__abc_74955_new_n397_; 
wire u2_u0__abc_74955_new_n398_; 
wire u2_u0__abc_74955_new_n399_; 
wire u2_u0__abc_74955_new_n400_; 
wire u2_u0__abc_74955_new_n401_; 
wire u2_u0__abc_74955_new_n402_; 
wire u2_u0__abc_74955_new_n403_; 
wire u2_u0__abc_74955_new_n404_; 
wire u2_u0__abc_74955_new_n405_; 
wire u2_u0__abc_74955_new_n406_; 
wire u2_u0__abc_74955_new_n407_; 
wire u2_u0__abc_74955_new_n408_; 
wire u2_u0__abc_74955_new_n409_; 
wire u2_u0__abc_74955_new_n410_; 
wire u2_u0__abc_74955_new_n411_; 
wire u2_u0__abc_74955_new_n412_; 
wire u2_u0__abc_74955_new_n413_; 
wire u2_u0__abc_74955_new_n414_; 
wire u2_u0__abc_74955_new_n415_; 
wire u2_u0__abc_74955_new_n416_; 
wire u2_u0__abc_74955_new_n417_; 
wire u2_u0__abc_74955_new_n418_; 
wire u2_u0__abc_74955_new_n419_; 
wire u2_u0__abc_74955_new_n420_; 
wire u2_u0__abc_74955_new_n421_; 
wire u2_u0__abc_74955_new_n422_; 
wire u2_u0__abc_74955_new_n423_; 
wire u2_u0__abc_74955_new_n424_; 
wire u2_u0__abc_74955_new_n425_; 
wire u2_u0__abc_74955_new_n426_; 
wire u2_u0__abc_74955_new_n427_; 
wire u2_u0__abc_74955_new_n428_; 
wire u2_u0__abc_74955_new_n429_; 
wire u2_u0__abc_74955_new_n430_; 
wire u2_u0__abc_74955_new_n431_; 
wire u2_u0__abc_74955_new_n432_; 
wire u2_u0__abc_74955_new_n433_; 
wire u2_u0__abc_74955_new_n434_; 
wire u2_u0__abc_74955_new_n435_; 
wire u2_u0__abc_74955_new_n436_; 
wire u2_u0__abc_74955_new_n437_; 
wire u2_u0__abc_74955_new_n438_; 
wire u2_u0__abc_74955_new_n439_; 
wire u2_u0__abc_74955_new_n440_; 
wire u2_u0__abc_74955_new_n441_; 
wire u2_u0__abc_74955_new_n442_; 
wire u2_u0__abc_74955_new_n443_; 
wire u2_u0__abc_74955_new_n444_; 
wire u2_u0__abc_74955_new_n445_; 
wire u2_u0__abc_74955_new_n446_; 
wire u2_u0__abc_74955_new_n447_; 
wire u2_u0__abc_74955_new_n448_; 
wire u2_u0__abc_74955_new_n449_; 
wire u2_u0__abc_74955_new_n450_; 
wire u2_u0__abc_74955_new_n451_; 
wire u2_u0__abc_74955_new_n452_; 
wire u2_u0__abc_74955_new_n453_; 
wire u2_u0__abc_74955_new_n454_; 
wire u2_u0__abc_74955_new_n455_; 
wire u2_u0__abc_74955_new_n456_; 
wire u2_u0__abc_74955_new_n457_; 
wire u2_u0__abc_74955_new_n458_; 
wire u2_u0__abc_74955_new_n459_; 
wire u2_u0__abc_74955_new_n460_; 
wire u2_u0__abc_74955_new_n461_; 
wire u2_u0__abc_74955_new_n462_; 
wire u2_u0__abc_74955_new_n463_; 
wire u2_u0__abc_74955_new_n464_; 
wire u2_u0__abc_74955_new_n465_; 
wire u2_u0__abc_74955_new_n466_; 
wire u2_u0__abc_74955_new_n467_; 
wire u2_u0__abc_74955_new_n468_; 
wire u2_u0__abc_74955_new_n469_; 
wire u2_u0__abc_74955_new_n470_; 
wire u2_u0__abc_74955_new_n471_; 
wire u2_u0__abc_74955_new_n472_; 
wire u2_u0__abc_74955_new_n473_; 
wire u2_u0__abc_74955_new_n474_; 
wire u2_u0__abc_74955_new_n475_; 
wire u2_u0__abc_74955_new_n476_; 
wire u2_u0__abc_74955_new_n477_; 
wire u2_u0__abc_74955_new_n478_; 
wire u2_u0__abc_74955_new_n479_; 
wire u2_u0__abc_74955_new_n480_; 
wire u2_u0__abc_74955_new_n481_; 
wire u2_u0__abc_74955_new_n482_; 
wire u2_u0__abc_74955_new_n483_; 
wire u2_u0__abc_74955_new_n484_; 
wire u2_u0__abc_74955_new_n485_; 
wire u2_u0__abc_74955_new_n486_; 
wire u2_u0__abc_74955_new_n487_; 
wire u2_u0__abc_74955_new_n488_; 
wire u2_u0__abc_74955_new_n489_; 
wire u2_u0__abc_74955_new_n490_; 
wire u2_u0__abc_74955_new_n491_; 
wire u2_u0__abc_74955_new_n492_; 
wire u2_u0__abc_74955_new_n493_; 
wire u2_u0__abc_74955_new_n494_; 
wire u2_u0__abc_74955_new_n495_; 
wire u2_u0__abc_74955_new_n496_; 
wire u2_u0__abc_74955_new_n497_; 
wire u2_u0__abc_74955_new_n498_; 
wire u2_u0__abc_74955_new_n499_; 
wire u2_u0__abc_74955_new_n500_; 
wire u2_u0__abc_74955_new_n501_; 
wire u2_u0__abc_74955_new_n502_; 
wire u2_u0__abc_74955_new_n503_; 
wire u2_u0__abc_74955_new_n504_; 
wire u2_u0__abc_74955_new_n505_; 
wire u2_u0__abc_74955_new_n506_; 
wire u2_u0__abc_74955_new_n507_; 
wire u2_u0__abc_74955_new_n508_; 
wire u2_u0__abc_74955_new_n509_; 
wire u2_u0__abc_74955_new_n510_; 
wire u2_u0__abc_74955_new_n511_; 
wire u2_u0__abc_74955_new_n512_; 
wire u2_u0__abc_74955_new_n513_; 
wire u2_u0__abc_74955_new_n514_; 
wire u2_u0__abc_74955_new_n515_; 
wire u2_u0__abc_74955_new_n516_; 
wire u2_u0__abc_74955_new_n517_; 
wire u2_u0__abc_74955_new_n518_; 
wire u2_u0__abc_74955_new_n519_; 
wire u2_u0__abc_74955_new_n520_; 
wire u2_u0__abc_74955_new_n521_; 
wire u2_u0__abc_74955_new_n522_; 
wire u2_u0__abc_74955_new_n523_; 
wire u2_u0__abc_74955_new_n524_; 
wire u2_u0__abc_74955_new_n525_; 
wire u2_u0__abc_74955_new_n526_; 
wire u2_u0__abc_74955_new_n527_; 
wire u2_u0__abc_74955_new_n528_; 
wire u2_u0__abc_74955_new_n529_; 
wire u2_u0__abc_74955_new_n530_; 
wire u2_u0__abc_74955_new_n531_; 
wire u2_u0__abc_74955_new_n532_; 
wire u2_u0__abc_74955_new_n533_; 
wire u2_u0__abc_74955_new_n534_; 
wire u2_u0__abc_74955_new_n535_; 
wire u2_u0__abc_74955_new_n536_; 
wire u2_u0__abc_74955_new_n537_; 
wire u2_u0__abc_74955_new_n538_; 
wire u2_u0__abc_74955_new_n539_; 
wire u2_u0__abc_74955_new_n540_; 
wire u2_u0__abc_74955_new_n541_; 
wire u2_u0__abc_74955_new_n542_; 
wire u2_u0__abc_74955_new_n543_; 
wire u2_u0__abc_74955_new_n544_; 
wire u2_u0__abc_74955_new_n545_; 
wire u2_u0__abc_74955_new_n546_; 
wire u2_u0__abc_74955_new_n547_; 
wire u2_u0__abc_74955_new_n548_; 
wire u2_u0__abc_74955_new_n549_; 
wire u2_u0__abc_74955_new_n550_; 
wire u2_u0__abc_74955_new_n551_; 
wire u2_u0__abc_74955_new_n552_; 
wire u2_u0__abc_74955_new_n553_; 
wire u2_u0__abc_74955_new_n554_; 
wire u2_u0__abc_74955_new_n555_; 
wire u2_u0__abc_74955_new_n556_; 
wire u2_u0__abc_74955_new_n557_; 
wire u2_u0__abc_74955_new_n558_; 
wire u2_u0__abc_74955_new_n559_; 
wire u2_u0__abc_74955_new_n560_; 
wire u2_u0__abc_74955_new_n561_; 
wire u2_u0__abc_74955_new_n562_; 
wire u2_u0__abc_74955_new_n563_; 
wire u2_u0__abc_74955_new_n564_; 
wire u2_u0__abc_74955_new_n565_; 
wire u2_u0__abc_74955_new_n566_; 
wire u2_u0__abc_74955_new_n567_; 
wire u2_u0__abc_74955_new_n568_; 
wire u2_u0__abc_74955_new_n569_; 
wire u2_u0__abc_74955_new_n570_; 
wire u2_u0__abc_74955_new_n571_; 
wire u2_u0__abc_74955_new_n572_; 
wire u2_u0__abc_74955_new_n573_; 
wire u2_u0__abc_74955_new_n574_; 
wire u2_u0__abc_74955_new_n575_; 
wire u2_u0__abc_74955_new_n576_; 
wire u2_u0__abc_74955_new_n577_; 
wire u2_u0__abc_74955_new_n578_; 
wire u2_u0__abc_74955_new_n579_; 
wire u2_u0__abc_74955_new_n580_; 
wire u2_u0__abc_74955_new_n581_; 
wire u2_u0__abc_74955_new_n582_; 
wire u2_u0__abc_74955_new_n583_; 
wire u2_u0__abc_74955_new_n584_; 
wire u2_u0__abc_74955_new_n585_; 
wire u2_u0__abc_74955_new_n586_; 
wire u2_u0__abc_74955_new_n587_; 
wire u2_u0__abc_74955_new_n588_; 
wire u2_u0__abc_74955_new_n589_; 
wire u2_u0__abc_74955_new_n590_; 
wire u2_u0__abc_74955_new_n591_; 
wire u2_u0__abc_74955_new_n592_; 
wire u2_u0__abc_74955_new_n594_; 
wire u2_u0__abc_74955_new_n595_; 
wire u2_u0__abc_74955_new_n596_; 
wire u2_u0__abc_74955_new_n597_; 
wire u2_u0__abc_74955_new_n598_; 
wire u2_u0__abc_74955_new_n599_; 
wire u2_u0__abc_74955_new_n601_; 
wire u2_u0__abc_74955_new_n602_; 
wire u2_u0__abc_74955_new_n603_; 
wire u2_u0__abc_74955_new_n604_; 
wire u2_u0__abc_74955_new_n605_; 
wire u2_u0__abc_74955_new_n606_; 
wire u2_u0__abc_74955_new_n608_; 
wire u2_u0__abc_74955_new_n609_; 
wire u2_u0__abc_74955_new_n610_; 
wire u2_u0__abc_74955_new_n611_; 
wire u2_u0__abc_74955_new_n616_; 
wire u2_u0__abc_74955_new_n617_; 
wire u2_u0__abc_74955_new_n618_; 
wire u2_u0__abc_74955_new_n619_; 
wire u2_u0__abc_74955_new_n621_; 
wire u2_u0__abc_74955_new_n622_; 
wire u2_u0__abc_74955_new_n623_; 
wire u2_u0__abc_74955_new_n624_; 
wire u2_u0_b0_last_row_0_; 
wire u2_u0_b0_last_row_10_; 
wire u2_u0_b0_last_row_11_; 
wire u2_u0_b0_last_row_12_; 
wire u2_u0_b0_last_row_1_; 
wire u2_u0_b0_last_row_2_; 
wire u2_u0_b0_last_row_3_; 
wire u2_u0_b0_last_row_4_; 
wire u2_u0_b0_last_row_5_; 
wire u2_u0_b0_last_row_6_; 
wire u2_u0_b0_last_row_7_; 
wire u2_u0_b0_last_row_8_; 
wire u2_u0_b0_last_row_9_; 
wire u2_u0_b1_last_row_0_; 
wire u2_u0_b1_last_row_10_; 
wire u2_u0_b1_last_row_11_; 
wire u2_u0_b1_last_row_12_; 
wire u2_u0_b1_last_row_1_; 
wire u2_u0_b1_last_row_2_; 
wire u2_u0_b1_last_row_3_; 
wire u2_u0_b1_last_row_4_; 
wire u2_u0_b1_last_row_5_; 
wire u2_u0_b1_last_row_6_; 
wire u2_u0_b1_last_row_7_; 
wire u2_u0_b1_last_row_8_; 
wire u2_u0_b1_last_row_9_; 
wire u2_u0_b2_last_row_0_; 
wire u2_u0_b2_last_row_10_; 
wire u2_u0_b2_last_row_11_; 
wire u2_u0_b2_last_row_12_; 
wire u2_u0_b2_last_row_1_; 
wire u2_u0_b2_last_row_2_; 
wire u2_u0_b2_last_row_3_; 
wire u2_u0_b2_last_row_4_; 
wire u2_u0_b2_last_row_5_; 
wire u2_u0_b2_last_row_6_; 
wire u2_u0_b2_last_row_7_; 
wire u2_u0_b2_last_row_8_; 
wire u2_u0_b2_last_row_9_; 
wire u2_u0_b3_last_row_0_; 
wire u2_u0_b3_last_row_10_; 
wire u2_u0_b3_last_row_11_; 
wire u2_u0_b3_last_row_12_; 
wire u2_u0_b3_last_row_1_; 
wire u2_u0_b3_last_row_2_; 
wire u2_u0_b3_last_row_3_; 
wire u2_u0_b3_last_row_4_; 
wire u2_u0_b3_last_row_5_; 
wire u2_u0_b3_last_row_6_; 
wire u2_u0_b3_last_row_7_; 
wire u2_u0_b3_last_row_8_; 
wire u2_u0_b3_last_row_9_; 
wire u2_u0_bank0_open; 
wire u2_u0_bank1_open; 
wire u2_u0_bank2_open; 
wire u2_u0_bank3_open; 
wire u2_u1__0b0_last_row_12_0__0_; 
wire u2_u1__0b0_last_row_12_0__10_; 
wire u2_u1__0b0_last_row_12_0__11_; 
wire u2_u1__0b0_last_row_12_0__12_; 
wire u2_u1__0b0_last_row_12_0__1_; 
wire u2_u1__0b0_last_row_12_0__2_; 
wire u2_u1__0b0_last_row_12_0__3_; 
wire u2_u1__0b0_last_row_12_0__4_; 
wire u2_u1__0b0_last_row_12_0__5_; 
wire u2_u1__0b0_last_row_12_0__6_; 
wire u2_u1__0b0_last_row_12_0__7_; 
wire u2_u1__0b0_last_row_12_0__8_; 
wire u2_u1__0b0_last_row_12_0__9_; 
wire u2_u1__0b1_last_row_12_0__0_; 
wire u2_u1__0b1_last_row_12_0__10_; 
wire u2_u1__0b1_last_row_12_0__11_; 
wire u2_u1__0b1_last_row_12_0__12_; 
wire u2_u1__0b1_last_row_12_0__1_; 
wire u2_u1__0b1_last_row_12_0__2_; 
wire u2_u1__0b1_last_row_12_0__3_; 
wire u2_u1__0b1_last_row_12_0__4_; 
wire u2_u1__0b1_last_row_12_0__5_; 
wire u2_u1__0b1_last_row_12_0__6_; 
wire u2_u1__0b1_last_row_12_0__7_; 
wire u2_u1__0b1_last_row_12_0__8_; 
wire u2_u1__0b1_last_row_12_0__9_; 
wire u2_u1__0b2_last_row_12_0__0_; 
wire u2_u1__0b2_last_row_12_0__10_; 
wire u2_u1__0b2_last_row_12_0__11_; 
wire u2_u1__0b2_last_row_12_0__12_; 
wire u2_u1__0b2_last_row_12_0__1_; 
wire u2_u1__0b2_last_row_12_0__2_; 
wire u2_u1__0b2_last_row_12_0__3_; 
wire u2_u1__0b2_last_row_12_0__4_; 
wire u2_u1__0b2_last_row_12_0__5_; 
wire u2_u1__0b2_last_row_12_0__6_; 
wire u2_u1__0b2_last_row_12_0__7_; 
wire u2_u1__0b2_last_row_12_0__8_; 
wire u2_u1__0b2_last_row_12_0__9_; 
wire u2_u1__0b3_last_row_12_0__0_; 
wire u2_u1__0b3_last_row_12_0__10_; 
wire u2_u1__0b3_last_row_12_0__11_; 
wire u2_u1__0b3_last_row_12_0__12_; 
wire u2_u1__0b3_last_row_12_0__1_; 
wire u2_u1__0b3_last_row_12_0__2_; 
wire u2_u1__0b3_last_row_12_0__3_; 
wire u2_u1__0b3_last_row_12_0__4_; 
wire u2_u1__0b3_last_row_12_0__5_; 
wire u2_u1__0b3_last_row_12_0__6_; 
wire u2_u1__0b3_last_row_12_0__7_; 
wire u2_u1__0b3_last_row_12_0__8_; 
wire u2_u1__0b3_last_row_12_0__9_; 
wire u2_u1__0bank0_open_0_0_; 
wire u2_u1__0bank1_open_0_0_; 
wire u2_u1__0bank2_open_0_0_; 
wire u2_u1__0bank3_open_0_0_; 
wire u2_u1__abc_74955_auto_rtlil_cc_1942_NotGate_71538; 
wire u2_u1__abc_74955_new_n136_; 
wire u2_u1__abc_74955_new_n137_; 
wire u2_u1__abc_74955_new_n137__bF_buf0; 
wire u2_u1__abc_74955_new_n137__bF_buf1; 
wire u2_u1__abc_74955_new_n137__bF_buf2; 
wire u2_u1__abc_74955_new_n137__bF_buf3; 
wire u2_u1__abc_74955_new_n137__bF_buf4; 
wire u2_u1__abc_74955_new_n138_; 
wire u2_u1__abc_74955_new_n139_; 
wire u2_u1__abc_74955_new_n140_; 
wire u2_u1__abc_74955_new_n141_; 
wire u2_u1__abc_74955_new_n143_; 
wire u2_u1__abc_74955_new_n144_; 
wire u2_u1__abc_74955_new_n145_; 
wire u2_u1__abc_74955_new_n146_; 
wire u2_u1__abc_74955_new_n148_; 
wire u2_u1__abc_74955_new_n149_; 
wire u2_u1__abc_74955_new_n150_; 
wire u2_u1__abc_74955_new_n151_; 
wire u2_u1__abc_74955_new_n153_; 
wire u2_u1__abc_74955_new_n154_; 
wire u2_u1__abc_74955_new_n155_; 
wire u2_u1__abc_74955_new_n156_; 
wire u2_u1__abc_74955_new_n158_; 
wire u2_u1__abc_74955_new_n159_; 
wire u2_u1__abc_74955_new_n160_; 
wire u2_u1__abc_74955_new_n161_; 
wire u2_u1__abc_74955_new_n163_; 
wire u2_u1__abc_74955_new_n164_; 
wire u2_u1__abc_74955_new_n165_; 
wire u2_u1__abc_74955_new_n166_; 
wire u2_u1__abc_74955_new_n168_; 
wire u2_u1__abc_74955_new_n169_; 
wire u2_u1__abc_74955_new_n170_; 
wire u2_u1__abc_74955_new_n171_; 
wire u2_u1__abc_74955_new_n173_; 
wire u2_u1__abc_74955_new_n174_; 
wire u2_u1__abc_74955_new_n175_; 
wire u2_u1__abc_74955_new_n176_; 
wire u2_u1__abc_74955_new_n178_; 
wire u2_u1__abc_74955_new_n179_; 
wire u2_u1__abc_74955_new_n180_; 
wire u2_u1__abc_74955_new_n181_; 
wire u2_u1__abc_74955_new_n183_; 
wire u2_u1__abc_74955_new_n184_; 
wire u2_u1__abc_74955_new_n185_; 
wire u2_u1__abc_74955_new_n186_; 
wire u2_u1__abc_74955_new_n188_; 
wire u2_u1__abc_74955_new_n189_; 
wire u2_u1__abc_74955_new_n190_; 
wire u2_u1__abc_74955_new_n191_; 
wire u2_u1__abc_74955_new_n193_; 
wire u2_u1__abc_74955_new_n194_; 
wire u2_u1__abc_74955_new_n195_; 
wire u2_u1__abc_74955_new_n196_; 
wire u2_u1__abc_74955_new_n198_; 
wire u2_u1__abc_74955_new_n199_; 
wire u2_u1__abc_74955_new_n200_; 
wire u2_u1__abc_74955_new_n201_; 
wire u2_u1__abc_74955_new_n203_; 
wire u2_u1__abc_74955_new_n204_; 
wire u2_u1__abc_74955_new_n205_; 
wire u2_u1__abc_74955_new_n206_; 
wire u2_u1__abc_74955_new_n207_; 
wire u2_u1__abc_74955_new_n208_; 
wire u2_u1__abc_74955_new_n209_; 
wire u2_u1__abc_74955_new_n211_; 
wire u2_u1__abc_74955_new_n212_; 
wire u2_u1__abc_74955_new_n214_; 
wire u2_u1__abc_74955_new_n215_; 
wire u2_u1__abc_74955_new_n217_; 
wire u2_u1__abc_74955_new_n218_; 
wire u2_u1__abc_74955_new_n220_; 
wire u2_u1__abc_74955_new_n221_; 
wire u2_u1__abc_74955_new_n223_; 
wire u2_u1__abc_74955_new_n224_; 
wire u2_u1__abc_74955_new_n226_; 
wire u2_u1__abc_74955_new_n227_; 
wire u2_u1__abc_74955_new_n229_; 
wire u2_u1__abc_74955_new_n230_; 
wire u2_u1__abc_74955_new_n232_; 
wire u2_u1__abc_74955_new_n233_; 
wire u2_u1__abc_74955_new_n235_; 
wire u2_u1__abc_74955_new_n236_; 
wire u2_u1__abc_74955_new_n238_; 
wire u2_u1__abc_74955_new_n239_; 
wire u2_u1__abc_74955_new_n241_; 
wire u2_u1__abc_74955_new_n242_; 
wire u2_u1__abc_74955_new_n244_; 
wire u2_u1__abc_74955_new_n245_; 
wire u2_u1__abc_74955_new_n247_; 
wire u2_u1__abc_74955_new_n248_; 
wire u2_u1__abc_74955_new_n249_; 
wire u2_u1__abc_74955_new_n250_; 
wire u2_u1__abc_74955_new_n251_; 
wire u2_u1__abc_74955_new_n253_; 
wire u2_u1__abc_74955_new_n254_; 
wire u2_u1__abc_74955_new_n256_; 
wire u2_u1__abc_74955_new_n257_; 
wire u2_u1__abc_74955_new_n259_; 
wire u2_u1__abc_74955_new_n260_; 
wire u2_u1__abc_74955_new_n262_; 
wire u2_u1__abc_74955_new_n263_; 
wire u2_u1__abc_74955_new_n265_; 
wire u2_u1__abc_74955_new_n266_; 
wire u2_u1__abc_74955_new_n268_; 
wire u2_u1__abc_74955_new_n269_; 
wire u2_u1__abc_74955_new_n271_; 
wire u2_u1__abc_74955_new_n272_; 
wire u2_u1__abc_74955_new_n274_; 
wire u2_u1__abc_74955_new_n275_; 
wire u2_u1__abc_74955_new_n277_; 
wire u2_u1__abc_74955_new_n278_; 
wire u2_u1__abc_74955_new_n280_; 
wire u2_u1__abc_74955_new_n281_; 
wire u2_u1__abc_74955_new_n283_; 
wire u2_u1__abc_74955_new_n284_; 
wire u2_u1__abc_74955_new_n286_; 
wire u2_u1__abc_74955_new_n287_; 
wire u2_u1__abc_74955_new_n289_; 
wire u2_u1__abc_74955_new_n290_; 
wire u2_u1__abc_74955_new_n291_; 
wire u2_u1__abc_74955_new_n292_; 
wire u2_u1__abc_74955_new_n293_; 
wire u2_u1__abc_74955_new_n295_; 
wire u2_u1__abc_74955_new_n296_; 
wire u2_u1__abc_74955_new_n298_; 
wire u2_u1__abc_74955_new_n299_; 
wire u2_u1__abc_74955_new_n301_; 
wire u2_u1__abc_74955_new_n302_; 
wire u2_u1__abc_74955_new_n304_; 
wire u2_u1__abc_74955_new_n305_; 
wire u2_u1__abc_74955_new_n307_; 
wire u2_u1__abc_74955_new_n308_; 
wire u2_u1__abc_74955_new_n310_; 
wire u2_u1__abc_74955_new_n311_; 
wire u2_u1__abc_74955_new_n313_; 
wire u2_u1__abc_74955_new_n314_; 
wire u2_u1__abc_74955_new_n316_; 
wire u2_u1__abc_74955_new_n317_; 
wire u2_u1__abc_74955_new_n319_; 
wire u2_u1__abc_74955_new_n320_; 
wire u2_u1__abc_74955_new_n322_; 
wire u2_u1__abc_74955_new_n323_; 
wire u2_u1__abc_74955_new_n325_; 
wire u2_u1__abc_74955_new_n326_; 
wire u2_u1__abc_74955_new_n328_; 
wire u2_u1__abc_74955_new_n329_; 
wire u2_u1__abc_74955_new_n331_; 
wire u2_u1__abc_74955_new_n332_; 
wire u2_u1__abc_74955_new_n333_; 
wire u2_u1__abc_74955_new_n334_; 
wire u2_u1__abc_74955_new_n335_; 
wire u2_u1__abc_74955_new_n336_; 
wire u2_u1__abc_74955_new_n337_; 
wire u2_u1__abc_74955_new_n338_; 
wire u2_u1__abc_74955_new_n339_; 
wire u2_u1__abc_74955_new_n340_; 
wire u2_u1__abc_74955_new_n341_; 
wire u2_u1__abc_74955_new_n342_; 
wire u2_u1__abc_74955_new_n343_; 
wire u2_u1__abc_74955_new_n344_; 
wire u2_u1__abc_74955_new_n345_; 
wire u2_u1__abc_74955_new_n346_; 
wire u2_u1__abc_74955_new_n347_; 
wire u2_u1__abc_74955_new_n348_; 
wire u2_u1__abc_74955_new_n349_; 
wire u2_u1__abc_74955_new_n350_; 
wire u2_u1__abc_74955_new_n351_; 
wire u2_u1__abc_74955_new_n352_; 
wire u2_u1__abc_74955_new_n353_; 
wire u2_u1__abc_74955_new_n354_; 
wire u2_u1__abc_74955_new_n355_; 
wire u2_u1__abc_74955_new_n356_; 
wire u2_u1__abc_74955_new_n357_; 
wire u2_u1__abc_74955_new_n358_; 
wire u2_u1__abc_74955_new_n359_; 
wire u2_u1__abc_74955_new_n360_; 
wire u2_u1__abc_74955_new_n361_; 
wire u2_u1__abc_74955_new_n362_; 
wire u2_u1__abc_74955_new_n363_; 
wire u2_u1__abc_74955_new_n364_; 
wire u2_u1__abc_74955_new_n365_; 
wire u2_u1__abc_74955_new_n366_; 
wire u2_u1__abc_74955_new_n367_; 
wire u2_u1__abc_74955_new_n368_; 
wire u2_u1__abc_74955_new_n369_; 
wire u2_u1__abc_74955_new_n370_; 
wire u2_u1__abc_74955_new_n371_; 
wire u2_u1__abc_74955_new_n372_; 
wire u2_u1__abc_74955_new_n373_; 
wire u2_u1__abc_74955_new_n374_; 
wire u2_u1__abc_74955_new_n375_; 
wire u2_u1__abc_74955_new_n376_; 
wire u2_u1__abc_74955_new_n377_; 
wire u2_u1__abc_74955_new_n378_; 
wire u2_u1__abc_74955_new_n379_; 
wire u2_u1__abc_74955_new_n380_; 
wire u2_u1__abc_74955_new_n381_; 
wire u2_u1__abc_74955_new_n382_; 
wire u2_u1__abc_74955_new_n383_; 
wire u2_u1__abc_74955_new_n384_; 
wire u2_u1__abc_74955_new_n385_; 
wire u2_u1__abc_74955_new_n386_; 
wire u2_u1__abc_74955_new_n387_; 
wire u2_u1__abc_74955_new_n388_; 
wire u2_u1__abc_74955_new_n389_; 
wire u2_u1__abc_74955_new_n390_; 
wire u2_u1__abc_74955_new_n391_; 
wire u2_u1__abc_74955_new_n392_; 
wire u2_u1__abc_74955_new_n393_; 
wire u2_u1__abc_74955_new_n394_; 
wire u2_u1__abc_74955_new_n395_; 
wire u2_u1__abc_74955_new_n396_; 
wire u2_u1__abc_74955_new_n397_; 
wire u2_u1__abc_74955_new_n398_; 
wire u2_u1__abc_74955_new_n399_; 
wire u2_u1__abc_74955_new_n400_; 
wire u2_u1__abc_74955_new_n401_; 
wire u2_u1__abc_74955_new_n402_; 
wire u2_u1__abc_74955_new_n403_; 
wire u2_u1__abc_74955_new_n404_; 
wire u2_u1__abc_74955_new_n405_; 
wire u2_u1__abc_74955_new_n406_; 
wire u2_u1__abc_74955_new_n407_; 
wire u2_u1__abc_74955_new_n408_; 
wire u2_u1__abc_74955_new_n409_; 
wire u2_u1__abc_74955_new_n410_; 
wire u2_u1__abc_74955_new_n411_; 
wire u2_u1__abc_74955_new_n412_; 
wire u2_u1__abc_74955_new_n413_; 
wire u2_u1__abc_74955_new_n414_; 
wire u2_u1__abc_74955_new_n415_; 
wire u2_u1__abc_74955_new_n416_; 
wire u2_u1__abc_74955_new_n417_; 
wire u2_u1__abc_74955_new_n418_; 
wire u2_u1__abc_74955_new_n419_; 
wire u2_u1__abc_74955_new_n420_; 
wire u2_u1__abc_74955_new_n421_; 
wire u2_u1__abc_74955_new_n422_; 
wire u2_u1__abc_74955_new_n423_; 
wire u2_u1__abc_74955_new_n424_; 
wire u2_u1__abc_74955_new_n425_; 
wire u2_u1__abc_74955_new_n426_; 
wire u2_u1__abc_74955_new_n427_; 
wire u2_u1__abc_74955_new_n428_; 
wire u2_u1__abc_74955_new_n429_; 
wire u2_u1__abc_74955_new_n430_; 
wire u2_u1__abc_74955_new_n431_; 
wire u2_u1__abc_74955_new_n432_; 
wire u2_u1__abc_74955_new_n433_; 
wire u2_u1__abc_74955_new_n434_; 
wire u2_u1__abc_74955_new_n435_; 
wire u2_u1__abc_74955_new_n436_; 
wire u2_u1__abc_74955_new_n437_; 
wire u2_u1__abc_74955_new_n438_; 
wire u2_u1__abc_74955_new_n439_; 
wire u2_u1__abc_74955_new_n440_; 
wire u2_u1__abc_74955_new_n441_; 
wire u2_u1__abc_74955_new_n442_; 
wire u2_u1__abc_74955_new_n443_; 
wire u2_u1__abc_74955_new_n444_; 
wire u2_u1__abc_74955_new_n445_; 
wire u2_u1__abc_74955_new_n446_; 
wire u2_u1__abc_74955_new_n447_; 
wire u2_u1__abc_74955_new_n448_; 
wire u2_u1__abc_74955_new_n449_; 
wire u2_u1__abc_74955_new_n450_; 
wire u2_u1__abc_74955_new_n451_; 
wire u2_u1__abc_74955_new_n452_; 
wire u2_u1__abc_74955_new_n453_; 
wire u2_u1__abc_74955_new_n454_; 
wire u2_u1__abc_74955_new_n455_; 
wire u2_u1__abc_74955_new_n456_; 
wire u2_u1__abc_74955_new_n457_; 
wire u2_u1__abc_74955_new_n458_; 
wire u2_u1__abc_74955_new_n459_; 
wire u2_u1__abc_74955_new_n460_; 
wire u2_u1__abc_74955_new_n461_; 
wire u2_u1__abc_74955_new_n462_; 
wire u2_u1__abc_74955_new_n463_; 
wire u2_u1__abc_74955_new_n464_; 
wire u2_u1__abc_74955_new_n465_; 
wire u2_u1__abc_74955_new_n466_; 
wire u2_u1__abc_74955_new_n467_; 
wire u2_u1__abc_74955_new_n468_; 
wire u2_u1__abc_74955_new_n469_; 
wire u2_u1__abc_74955_new_n470_; 
wire u2_u1__abc_74955_new_n471_; 
wire u2_u1__abc_74955_new_n472_; 
wire u2_u1__abc_74955_new_n473_; 
wire u2_u1__abc_74955_new_n474_; 
wire u2_u1__abc_74955_new_n475_; 
wire u2_u1__abc_74955_new_n476_; 
wire u2_u1__abc_74955_new_n477_; 
wire u2_u1__abc_74955_new_n478_; 
wire u2_u1__abc_74955_new_n479_; 
wire u2_u1__abc_74955_new_n480_; 
wire u2_u1__abc_74955_new_n481_; 
wire u2_u1__abc_74955_new_n482_; 
wire u2_u1__abc_74955_new_n483_; 
wire u2_u1__abc_74955_new_n484_; 
wire u2_u1__abc_74955_new_n485_; 
wire u2_u1__abc_74955_new_n486_; 
wire u2_u1__abc_74955_new_n487_; 
wire u2_u1__abc_74955_new_n488_; 
wire u2_u1__abc_74955_new_n489_; 
wire u2_u1__abc_74955_new_n490_; 
wire u2_u1__abc_74955_new_n491_; 
wire u2_u1__abc_74955_new_n492_; 
wire u2_u1__abc_74955_new_n493_; 
wire u2_u1__abc_74955_new_n494_; 
wire u2_u1__abc_74955_new_n495_; 
wire u2_u1__abc_74955_new_n496_; 
wire u2_u1__abc_74955_new_n497_; 
wire u2_u1__abc_74955_new_n498_; 
wire u2_u1__abc_74955_new_n499_; 
wire u2_u1__abc_74955_new_n500_; 
wire u2_u1__abc_74955_new_n501_; 
wire u2_u1__abc_74955_new_n502_; 
wire u2_u1__abc_74955_new_n503_; 
wire u2_u1__abc_74955_new_n504_; 
wire u2_u1__abc_74955_new_n505_; 
wire u2_u1__abc_74955_new_n506_; 
wire u2_u1__abc_74955_new_n507_; 
wire u2_u1__abc_74955_new_n508_; 
wire u2_u1__abc_74955_new_n509_; 
wire u2_u1__abc_74955_new_n510_; 
wire u2_u1__abc_74955_new_n511_; 
wire u2_u1__abc_74955_new_n512_; 
wire u2_u1__abc_74955_new_n513_; 
wire u2_u1__abc_74955_new_n514_; 
wire u2_u1__abc_74955_new_n515_; 
wire u2_u1__abc_74955_new_n516_; 
wire u2_u1__abc_74955_new_n517_; 
wire u2_u1__abc_74955_new_n518_; 
wire u2_u1__abc_74955_new_n519_; 
wire u2_u1__abc_74955_new_n520_; 
wire u2_u1__abc_74955_new_n521_; 
wire u2_u1__abc_74955_new_n522_; 
wire u2_u1__abc_74955_new_n523_; 
wire u2_u1__abc_74955_new_n524_; 
wire u2_u1__abc_74955_new_n525_; 
wire u2_u1__abc_74955_new_n526_; 
wire u2_u1__abc_74955_new_n527_; 
wire u2_u1__abc_74955_new_n528_; 
wire u2_u1__abc_74955_new_n529_; 
wire u2_u1__abc_74955_new_n530_; 
wire u2_u1__abc_74955_new_n531_; 
wire u2_u1__abc_74955_new_n532_; 
wire u2_u1__abc_74955_new_n533_; 
wire u2_u1__abc_74955_new_n534_; 
wire u2_u1__abc_74955_new_n535_; 
wire u2_u1__abc_74955_new_n536_; 
wire u2_u1__abc_74955_new_n537_; 
wire u2_u1__abc_74955_new_n538_; 
wire u2_u1__abc_74955_new_n539_; 
wire u2_u1__abc_74955_new_n540_; 
wire u2_u1__abc_74955_new_n541_; 
wire u2_u1__abc_74955_new_n542_; 
wire u2_u1__abc_74955_new_n543_; 
wire u2_u1__abc_74955_new_n544_; 
wire u2_u1__abc_74955_new_n545_; 
wire u2_u1__abc_74955_new_n546_; 
wire u2_u1__abc_74955_new_n547_; 
wire u2_u1__abc_74955_new_n548_; 
wire u2_u1__abc_74955_new_n549_; 
wire u2_u1__abc_74955_new_n550_; 
wire u2_u1__abc_74955_new_n551_; 
wire u2_u1__abc_74955_new_n552_; 
wire u2_u1__abc_74955_new_n553_; 
wire u2_u1__abc_74955_new_n554_; 
wire u2_u1__abc_74955_new_n555_; 
wire u2_u1__abc_74955_new_n556_; 
wire u2_u1__abc_74955_new_n557_; 
wire u2_u1__abc_74955_new_n558_; 
wire u2_u1__abc_74955_new_n559_; 
wire u2_u1__abc_74955_new_n560_; 
wire u2_u1__abc_74955_new_n561_; 
wire u2_u1__abc_74955_new_n562_; 
wire u2_u1__abc_74955_new_n563_; 
wire u2_u1__abc_74955_new_n564_; 
wire u2_u1__abc_74955_new_n565_; 
wire u2_u1__abc_74955_new_n566_; 
wire u2_u1__abc_74955_new_n567_; 
wire u2_u1__abc_74955_new_n568_; 
wire u2_u1__abc_74955_new_n569_; 
wire u2_u1__abc_74955_new_n570_; 
wire u2_u1__abc_74955_new_n571_; 
wire u2_u1__abc_74955_new_n572_; 
wire u2_u1__abc_74955_new_n573_; 
wire u2_u1__abc_74955_new_n574_; 
wire u2_u1__abc_74955_new_n575_; 
wire u2_u1__abc_74955_new_n576_; 
wire u2_u1__abc_74955_new_n577_; 
wire u2_u1__abc_74955_new_n578_; 
wire u2_u1__abc_74955_new_n579_; 
wire u2_u1__abc_74955_new_n580_; 
wire u2_u1__abc_74955_new_n581_; 
wire u2_u1__abc_74955_new_n582_; 
wire u2_u1__abc_74955_new_n583_; 
wire u2_u1__abc_74955_new_n584_; 
wire u2_u1__abc_74955_new_n585_; 
wire u2_u1__abc_74955_new_n586_; 
wire u2_u1__abc_74955_new_n587_; 
wire u2_u1__abc_74955_new_n588_; 
wire u2_u1__abc_74955_new_n589_; 
wire u2_u1__abc_74955_new_n590_; 
wire u2_u1__abc_74955_new_n591_; 
wire u2_u1__abc_74955_new_n592_; 
wire u2_u1__abc_74955_new_n594_; 
wire u2_u1__abc_74955_new_n595_; 
wire u2_u1__abc_74955_new_n596_; 
wire u2_u1__abc_74955_new_n597_; 
wire u2_u1__abc_74955_new_n598_; 
wire u2_u1__abc_74955_new_n599_; 
wire u2_u1__abc_74955_new_n601_; 
wire u2_u1__abc_74955_new_n602_; 
wire u2_u1__abc_74955_new_n603_; 
wire u2_u1__abc_74955_new_n604_; 
wire u2_u1__abc_74955_new_n605_; 
wire u2_u1__abc_74955_new_n606_; 
wire u2_u1__abc_74955_new_n608_; 
wire u2_u1__abc_74955_new_n609_; 
wire u2_u1__abc_74955_new_n610_; 
wire u2_u1__abc_74955_new_n611_; 
wire u2_u1__abc_74955_new_n616_; 
wire u2_u1__abc_74955_new_n617_; 
wire u2_u1__abc_74955_new_n618_; 
wire u2_u1__abc_74955_new_n619_; 
wire u2_u1__abc_74955_new_n621_; 
wire u2_u1__abc_74955_new_n622_; 
wire u2_u1__abc_74955_new_n623_; 
wire u2_u1__abc_74955_new_n624_; 
wire u2_u1_b0_last_row_0_; 
wire u2_u1_b0_last_row_10_; 
wire u2_u1_b0_last_row_11_; 
wire u2_u1_b0_last_row_12_; 
wire u2_u1_b0_last_row_1_; 
wire u2_u1_b0_last_row_2_; 
wire u2_u1_b0_last_row_3_; 
wire u2_u1_b0_last_row_4_; 
wire u2_u1_b0_last_row_5_; 
wire u2_u1_b0_last_row_6_; 
wire u2_u1_b0_last_row_7_; 
wire u2_u1_b0_last_row_8_; 
wire u2_u1_b0_last_row_9_; 
wire u2_u1_b1_last_row_0_; 
wire u2_u1_b1_last_row_10_; 
wire u2_u1_b1_last_row_11_; 
wire u2_u1_b1_last_row_12_; 
wire u2_u1_b1_last_row_1_; 
wire u2_u1_b1_last_row_2_; 
wire u2_u1_b1_last_row_3_; 
wire u2_u1_b1_last_row_4_; 
wire u2_u1_b1_last_row_5_; 
wire u2_u1_b1_last_row_6_; 
wire u2_u1_b1_last_row_7_; 
wire u2_u1_b1_last_row_8_; 
wire u2_u1_b1_last_row_9_; 
wire u2_u1_b2_last_row_0_; 
wire u2_u1_b2_last_row_10_; 
wire u2_u1_b2_last_row_11_; 
wire u2_u1_b2_last_row_12_; 
wire u2_u1_b2_last_row_1_; 
wire u2_u1_b2_last_row_2_; 
wire u2_u1_b2_last_row_3_; 
wire u2_u1_b2_last_row_4_; 
wire u2_u1_b2_last_row_5_; 
wire u2_u1_b2_last_row_6_; 
wire u2_u1_b2_last_row_7_; 
wire u2_u1_b2_last_row_8_; 
wire u2_u1_b2_last_row_9_; 
wire u2_u1_b3_last_row_0_; 
wire u2_u1_b3_last_row_10_; 
wire u2_u1_b3_last_row_11_; 
wire u2_u1_b3_last_row_12_; 
wire u2_u1_b3_last_row_1_; 
wire u2_u1_b3_last_row_2_; 
wire u2_u1_b3_last_row_3_; 
wire u2_u1_b3_last_row_4_; 
wire u2_u1_b3_last_row_5_; 
wire u2_u1_b3_last_row_6_; 
wire u2_u1_b3_last_row_7_; 
wire u2_u1_b3_last_row_8_; 
wire u2_u1_b3_last_row_9_; 
wire u2_u1_bank0_open; 
wire u2_u1_bank1_open; 
wire u2_u1_bank2_open; 
wire u2_u1_bank3_open; 
wire u3__0byte0_7_0__0_; 
wire u3__0byte0_7_0__1_; 
wire u3__0byte0_7_0__2_; 
wire u3__0byte0_7_0__3_; 
wire u3__0byte0_7_0__4_; 
wire u3__0byte0_7_0__5_; 
wire u3__0byte0_7_0__6_; 
wire u3__0byte0_7_0__7_; 
wire u3__0byte1_7_0__0_; 
wire u3__0byte1_7_0__1_; 
wire u3__0byte1_7_0__2_; 
wire u3__0byte1_7_0__3_; 
wire u3__0byte1_7_0__4_; 
wire u3__0byte1_7_0__5_; 
wire u3__0byte1_7_0__6_; 
wire u3__0byte1_7_0__7_; 
wire u3__0byte2_7_0__0_; 
wire u3__0byte2_7_0__1_; 
wire u3__0byte2_7_0__2_; 
wire u3__0byte2_7_0__3_; 
wire u3__0byte2_7_0__4_; 
wire u3__0byte2_7_0__5_; 
wire u3__0byte2_7_0__6_; 
wire u3__0byte2_7_0__7_; 
wire u3__0mc_data_o_31_0__0_; 
wire u3__0mc_data_o_31_0__10_; 
wire u3__0mc_data_o_31_0__11_; 
wire u3__0mc_data_o_31_0__12_; 
wire u3__0mc_data_o_31_0__13_; 
wire u3__0mc_data_o_31_0__14_; 
wire u3__0mc_data_o_31_0__15_; 
wire u3__0mc_data_o_31_0__16_; 
wire u3__0mc_data_o_31_0__17_; 
wire u3__0mc_data_o_31_0__18_; 
wire u3__0mc_data_o_31_0__19_; 
wire u3__0mc_data_o_31_0__1_; 
wire u3__0mc_data_o_31_0__20_; 
wire u3__0mc_data_o_31_0__21_; 
wire u3__0mc_data_o_31_0__22_; 
wire u3__0mc_data_o_31_0__23_; 
wire u3__0mc_data_o_31_0__24_; 
wire u3__0mc_data_o_31_0__25_; 
wire u3__0mc_data_o_31_0__26_; 
wire u3__0mc_data_o_31_0__27_; 
wire u3__0mc_data_o_31_0__28_; 
wire u3__0mc_data_o_31_0__29_; 
wire u3__0mc_data_o_31_0__2_; 
wire u3__0mc_data_o_31_0__30_; 
wire u3__0mc_data_o_31_0__31_; 
wire u3__0mc_data_o_31_0__3_; 
wire u3__0mc_data_o_31_0__4_; 
wire u3__0mc_data_o_31_0__5_; 
wire u3__0mc_data_o_31_0__6_; 
wire u3__0mc_data_o_31_0__7_; 
wire u3__0mc_data_o_31_0__8_; 
wire u3__0mc_data_o_31_0__9_; 
wire u3__0mc_dp_o_3_0__0_; 
wire u3__0mc_dp_o_3_0__1_; 
wire u3__0mc_dp_o_3_0__2_; 
wire u3__0mc_dp_o_3_0__3_; 
wire u3__abc_74070_new_n1000_; 
wire u3__abc_74070_new_n1001_; 
wire u3__abc_74070_new_n1002_; 
wire u3__abc_74070_new_n1003_; 
wire u3__abc_74070_new_n1004_; 
wire u3__abc_74070_new_n1005_; 
wire u3__abc_74070_new_n1006_; 
wire u3__abc_74070_new_n1007_; 
wire u3__abc_74070_new_n1008_; 
wire u3__abc_74070_new_n1009_; 
wire u3__abc_74070_new_n1010_; 
wire u3__abc_74070_new_n1011_; 
wire u3__abc_74070_new_n1012_; 
wire u3__abc_74070_new_n1013_; 
wire u3__abc_74070_new_n1014_; 
wire u3__abc_74070_new_n1015_; 
wire u3__abc_74070_new_n1016_; 
wire u3__abc_74070_new_n1017_; 
wire u3__abc_74070_new_n1018_; 
wire u3__abc_74070_new_n1019_; 
wire u3__abc_74070_new_n1020_; 
wire u3__abc_74070_new_n1021_; 
wire u3__abc_74070_new_n1022_; 
wire u3__abc_74070_new_n1023_; 
wire u3__abc_74070_new_n1024_; 
wire u3__abc_74070_new_n1025_; 
wire u3__abc_74070_new_n1026_; 
wire u3__abc_74070_new_n1027_; 
wire u3__abc_74070_new_n1028_; 
wire u3__abc_74070_new_n1029_; 
wire u3__abc_74070_new_n1030_; 
wire u3__abc_74070_new_n1031_; 
wire u3__abc_74070_new_n1032_; 
wire u3__abc_74070_new_n275_; 
wire u3__abc_74070_new_n275__bF_buf0; 
wire u3__abc_74070_new_n275__bF_buf1; 
wire u3__abc_74070_new_n275__bF_buf2; 
wire u3__abc_74070_new_n275__bF_buf3; 
wire u3__abc_74070_new_n275__bF_buf4; 
wire u3__abc_74070_new_n276_; 
wire u3__abc_74070_new_n277_; 
wire u3__abc_74070_new_n277__bF_buf0; 
wire u3__abc_74070_new_n277__bF_buf1; 
wire u3__abc_74070_new_n277__bF_buf2; 
wire u3__abc_74070_new_n277__bF_buf3; 
wire u3__abc_74070_new_n277__bF_buf4; 
wire u3__abc_74070_new_n277__bF_buf5; 
wire u3__abc_74070_new_n278_; 
wire u3__abc_74070_new_n279_; 
wire u3__abc_74070_new_n279__bF_buf0; 
wire u3__abc_74070_new_n279__bF_buf1; 
wire u3__abc_74070_new_n279__bF_buf2; 
wire u3__abc_74070_new_n279__bF_buf3; 
wire u3__abc_74070_new_n279__bF_buf4; 
wire u3__abc_74070_new_n279__bF_buf5; 
wire u3__abc_74070_new_n280_; 
wire u3__abc_74070_new_n281_; 
wire u3__abc_74070_new_n282_; 
wire u3__abc_74070_new_n283_; 
wire u3__abc_74070_new_n284_; 
wire u3__abc_74070_new_n285_; 
wire u3__abc_74070_new_n286_; 
wire u3__abc_74070_new_n287_; 
wire u3__abc_74070_new_n288_; 
wire u3__abc_74070_new_n289_; 
wire u3__abc_74070_new_n290_; 
wire u3__abc_74070_new_n291_; 
wire u3__abc_74070_new_n292_; 
wire u3__abc_74070_new_n293_; 
wire u3__abc_74070_new_n294_; 
wire u3__abc_74070_new_n295_; 
wire u3__abc_74070_new_n296_; 
wire u3__abc_74070_new_n297_; 
wire u3__abc_74070_new_n298_; 
wire u3__abc_74070_new_n299_; 
wire u3__abc_74070_new_n300_; 
wire u3__abc_74070_new_n301_; 
wire u3__abc_74070_new_n302_; 
wire u3__abc_74070_new_n303_; 
wire u3__abc_74070_new_n304_; 
wire u3__abc_74070_new_n305_; 
wire u3__abc_74070_new_n306_; 
wire u3__abc_74070_new_n307_; 
wire u3__abc_74070_new_n308_; 
wire u3__abc_74070_new_n309_; 
wire u3__abc_74070_new_n310_; 
wire u3__abc_74070_new_n311_; 
wire u3__abc_74070_new_n312_; 
wire u3__abc_74070_new_n313_; 
wire u3__abc_74070_new_n315_; 
wire u3__abc_74070_new_n316_; 
wire u3__abc_74070_new_n317_; 
wire u3__abc_74070_new_n318_; 
wire u3__abc_74070_new_n319_; 
wire u3__abc_74070_new_n320_; 
wire u3__abc_74070_new_n321_; 
wire u3__abc_74070_new_n322_; 
wire u3__abc_74070_new_n323_; 
wire u3__abc_74070_new_n324_; 
wire u3__abc_74070_new_n325_; 
wire u3__abc_74070_new_n326_; 
wire u3__abc_74070_new_n327_; 
wire u3__abc_74070_new_n328_; 
wire u3__abc_74070_new_n329_; 
wire u3__abc_74070_new_n330_; 
wire u3__abc_74070_new_n331_; 
wire u3__abc_74070_new_n332_; 
wire u3__abc_74070_new_n333_; 
wire u3__abc_74070_new_n334_; 
wire u3__abc_74070_new_n335_; 
wire u3__abc_74070_new_n336_; 
wire u3__abc_74070_new_n337_; 
wire u3__abc_74070_new_n338_; 
wire u3__abc_74070_new_n339_; 
wire u3__abc_74070_new_n340_; 
wire u3__abc_74070_new_n341_; 
wire u3__abc_74070_new_n342_; 
wire u3__abc_74070_new_n343_; 
wire u3__abc_74070_new_n344_; 
wire u3__abc_74070_new_n345_; 
wire u3__abc_74070_new_n346_; 
wire u3__abc_74070_new_n347_; 
wire u3__abc_74070_new_n348_; 
wire u3__abc_74070_new_n349_; 
wire u3__abc_74070_new_n351_; 
wire u3__abc_74070_new_n352_; 
wire u3__abc_74070_new_n353_; 
wire u3__abc_74070_new_n354_; 
wire u3__abc_74070_new_n355_; 
wire u3__abc_74070_new_n356_; 
wire u3__abc_74070_new_n357_; 
wire u3__abc_74070_new_n358_; 
wire u3__abc_74070_new_n359_; 
wire u3__abc_74070_new_n360_; 
wire u3__abc_74070_new_n361_; 
wire u3__abc_74070_new_n362_; 
wire u3__abc_74070_new_n363_; 
wire u3__abc_74070_new_n364_; 
wire u3__abc_74070_new_n365_; 
wire u3__abc_74070_new_n366_; 
wire u3__abc_74070_new_n367_; 
wire u3__abc_74070_new_n368_; 
wire u3__abc_74070_new_n369_; 
wire u3__abc_74070_new_n370_; 
wire u3__abc_74070_new_n371_; 
wire u3__abc_74070_new_n372_; 
wire u3__abc_74070_new_n373_; 
wire u3__abc_74070_new_n374_; 
wire u3__abc_74070_new_n375_; 
wire u3__abc_74070_new_n376_; 
wire u3__abc_74070_new_n377_; 
wire u3__abc_74070_new_n378_; 
wire u3__abc_74070_new_n379_; 
wire u3__abc_74070_new_n380_; 
wire u3__abc_74070_new_n381_; 
wire u3__abc_74070_new_n382_; 
wire u3__abc_74070_new_n383_; 
wire u3__abc_74070_new_n384_; 
wire u3__abc_74070_new_n385_; 
wire u3__abc_74070_new_n387_; 
wire u3__abc_74070_new_n388_; 
wire u3__abc_74070_new_n389_; 
wire u3__abc_74070_new_n390_; 
wire u3__abc_74070_new_n391_; 
wire u3__abc_74070_new_n392_; 
wire u3__abc_74070_new_n393_; 
wire u3__abc_74070_new_n394_; 
wire u3__abc_74070_new_n395_; 
wire u3__abc_74070_new_n396_; 
wire u3__abc_74070_new_n397_; 
wire u3__abc_74070_new_n398_; 
wire u3__abc_74070_new_n399_; 
wire u3__abc_74070_new_n400_; 
wire u3__abc_74070_new_n401_; 
wire u3__abc_74070_new_n402_; 
wire u3__abc_74070_new_n403_; 
wire u3__abc_74070_new_n404_; 
wire u3__abc_74070_new_n405_; 
wire u3__abc_74070_new_n406_; 
wire u3__abc_74070_new_n407_; 
wire u3__abc_74070_new_n408_; 
wire u3__abc_74070_new_n409_; 
wire u3__abc_74070_new_n410_; 
wire u3__abc_74070_new_n411_; 
wire u3__abc_74070_new_n412_; 
wire u3__abc_74070_new_n413_; 
wire u3__abc_74070_new_n414_; 
wire u3__abc_74070_new_n415_; 
wire u3__abc_74070_new_n416_; 
wire u3__abc_74070_new_n417_; 
wire u3__abc_74070_new_n418_; 
wire u3__abc_74070_new_n419_; 
wire u3__abc_74070_new_n420_; 
wire u3__abc_74070_new_n421_; 
wire u3__abc_74070_new_n423_; 
wire u3__abc_74070_new_n424_; 
wire u3__abc_74070_new_n425_; 
wire u3__abc_74070_new_n427_; 
wire u3__abc_74070_new_n428_; 
wire u3__abc_74070_new_n430_; 
wire u3__abc_74070_new_n431_; 
wire u3__abc_74070_new_n433_; 
wire u3__abc_74070_new_n434_; 
wire u3__abc_74070_new_n436_; 
wire u3__abc_74070_new_n437_; 
wire u3__abc_74070_new_n439_; 
wire u3__abc_74070_new_n440_; 
wire u3__abc_74070_new_n442_; 
wire u3__abc_74070_new_n443_; 
wire u3__abc_74070_new_n445_; 
wire u3__abc_74070_new_n446_; 
wire u3__abc_74070_new_n448_; 
wire u3__abc_74070_new_n449_; 
wire u3__abc_74070_new_n449__bF_buf0; 
wire u3__abc_74070_new_n449__bF_buf1; 
wire u3__abc_74070_new_n449__bF_buf2; 
wire u3__abc_74070_new_n449__bF_buf3; 
wire u3__abc_74070_new_n450_; 
wire u3__abc_74070_new_n450__bF_buf0; 
wire u3__abc_74070_new_n450__bF_buf1; 
wire u3__abc_74070_new_n450__bF_buf2; 
wire u3__abc_74070_new_n450__bF_buf3; 
wire u3__abc_74070_new_n451_; 
wire u3__abc_74070_new_n452_; 
wire u3__abc_74070_new_n452__bF_buf0; 
wire u3__abc_74070_new_n452__bF_buf1; 
wire u3__abc_74070_new_n452__bF_buf2; 
wire u3__abc_74070_new_n452__bF_buf3; 
wire u3__abc_74070_new_n453_; 
wire u3__abc_74070_new_n454_; 
wire u3__abc_74070_new_n455_; 
wire u3__abc_74070_new_n456_; 
wire u3__abc_74070_new_n457_; 
wire u3__abc_74070_new_n458_; 
wire u3__abc_74070_new_n459_; 
wire u3__abc_74070_new_n460_; 
wire u3__abc_74070_new_n462_; 
wire u3__abc_74070_new_n463_; 
wire u3__abc_74070_new_n464_; 
wire u3__abc_74070_new_n465_; 
wire u3__abc_74070_new_n466_; 
wire u3__abc_74070_new_n468_; 
wire u3__abc_74070_new_n469_; 
wire u3__abc_74070_new_n470_; 
wire u3__abc_74070_new_n471_; 
wire u3__abc_74070_new_n472_; 
wire u3__abc_74070_new_n474_; 
wire u3__abc_74070_new_n475_; 
wire u3__abc_74070_new_n476_; 
wire u3__abc_74070_new_n477_; 
wire u3__abc_74070_new_n478_; 
wire u3__abc_74070_new_n480_; 
wire u3__abc_74070_new_n481_; 
wire u3__abc_74070_new_n482_; 
wire u3__abc_74070_new_n483_; 
wire u3__abc_74070_new_n484_; 
wire u3__abc_74070_new_n486_; 
wire u3__abc_74070_new_n487_; 
wire u3__abc_74070_new_n488_; 
wire u3__abc_74070_new_n489_; 
wire u3__abc_74070_new_n490_; 
wire u3__abc_74070_new_n492_; 
wire u3__abc_74070_new_n493_; 
wire u3__abc_74070_new_n494_; 
wire u3__abc_74070_new_n495_; 
wire u3__abc_74070_new_n496_; 
wire u3__abc_74070_new_n498_; 
wire u3__abc_74070_new_n499_; 
wire u3__abc_74070_new_n500_; 
wire u3__abc_74070_new_n501_; 
wire u3__abc_74070_new_n502_; 
wire u3__abc_74070_new_n504_; 
wire u3__abc_74070_new_n505_; 
wire u3__abc_74070_new_n506_; 
wire u3__abc_74070_new_n508_; 
wire u3__abc_74070_new_n509_; 
wire u3__abc_74070_new_n511_; 
wire u3__abc_74070_new_n512_; 
wire u3__abc_74070_new_n514_; 
wire u3__abc_74070_new_n515_; 
wire u3__abc_74070_new_n517_; 
wire u3__abc_74070_new_n518_; 
wire u3__abc_74070_new_n520_; 
wire u3__abc_74070_new_n521_; 
wire u3__abc_74070_new_n523_; 
wire u3__abc_74070_new_n524_; 
wire u3__abc_74070_new_n526_; 
wire u3__abc_74070_new_n527_; 
wire u3__abc_74070_new_n529_; 
wire u3__abc_74070_new_n530_; 
wire u3__abc_74070_new_n532_; 
wire u3__abc_74070_new_n533_; 
wire u3__abc_74070_new_n535_; 
wire u3__abc_74070_new_n536_; 
wire u3__abc_74070_new_n538_; 
wire u3__abc_74070_new_n539_; 
wire u3__abc_74070_new_n541_; 
wire u3__abc_74070_new_n542_; 
wire u3__abc_74070_new_n544_; 
wire u3__abc_74070_new_n545_; 
wire u3__abc_74070_new_n547_; 
wire u3__abc_74070_new_n548_; 
wire u3__abc_74070_new_n550_; 
wire u3__abc_74070_new_n551_; 
wire u3__abc_74070_new_n553_; 
wire u3__abc_74070_new_n554_; 
wire u3__abc_74070_new_n556_; 
wire u3__abc_74070_new_n557_; 
wire u3__abc_74070_new_n559_; 
wire u3__abc_74070_new_n560_; 
wire u3__abc_74070_new_n562_; 
wire u3__abc_74070_new_n563_; 
wire u3__abc_74070_new_n565_; 
wire u3__abc_74070_new_n566_; 
wire u3__abc_74070_new_n568_; 
wire u3__abc_74070_new_n569_; 
wire u3__abc_74070_new_n571_; 
wire u3__abc_74070_new_n572_; 
wire u3__abc_74070_new_n574_; 
wire u3__abc_74070_new_n575_; 
wire u3__abc_74070_new_n577_; 
wire u3__abc_74070_new_n578_; 
wire u3__abc_74070_new_n580_; 
wire u3__abc_74070_new_n581_; 
wire u3__abc_74070_new_n583_; 
wire u3__abc_74070_new_n584_; 
wire u3__abc_74070_new_n586_; 
wire u3__abc_74070_new_n587_; 
wire u3__abc_74070_new_n589_; 
wire u3__abc_74070_new_n590_; 
wire u3__abc_74070_new_n592_; 
wire u3__abc_74070_new_n593_; 
wire u3__abc_74070_new_n595_; 
wire u3__abc_74070_new_n596_; 
wire u3__abc_74070_new_n598_; 
wire u3__abc_74070_new_n599_; 
wire u3__abc_74070_new_n601_; 
wire u3__abc_74070_new_n602_; 
wire u3__abc_74070_new_n604_; 
wire u3__abc_74070_new_n605_; 
wire u3__abc_74070_new_n607_; 
wire u3__abc_74070_new_n608_; 
wire u3__abc_74070_new_n610_; 
wire u3__abc_74070_new_n611_; 
wire u3__abc_74070_new_n613_; 
wire u3__abc_74070_new_n614_; 
wire u3__abc_74070_new_n616_; 
wire u3__abc_74070_new_n617_; 
wire u3__abc_74070_new_n619_; 
wire u3__abc_74070_new_n620_; 
wire u3__abc_74070_new_n622_; 
wire u3__abc_74070_new_n623_; 
wire u3__abc_74070_new_n625_; 
wire u3__abc_74070_new_n625__bF_buf0; 
wire u3__abc_74070_new_n625__bF_buf1; 
wire u3__abc_74070_new_n625__bF_buf2; 
wire u3__abc_74070_new_n625__bF_buf3; 
wire u3__abc_74070_new_n625__bF_buf4; 
wire u3__abc_74070_new_n626_; 
wire u3__abc_74070_new_n627_; 
wire u3__abc_74070_new_n628_; 
wire u3__abc_74070_new_n629_; 
wire u3__abc_74070_new_n630_; 
wire u3__abc_74070_new_n632_; 
wire u3__abc_74070_new_n633_; 
wire u3__abc_74070_new_n634_; 
wire u3__abc_74070_new_n635_; 
wire u3__abc_74070_new_n636_; 
wire u3__abc_74070_new_n638_; 
wire u3__abc_74070_new_n639_; 
wire u3__abc_74070_new_n640_; 
wire u3__abc_74070_new_n641_; 
wire u3__abc_74070_new_n642_; 
wire u3__abc_74070_new_n644_; 
wire u3__abc_74070_new_n645_; 
wire u3__abc_74070_new_n646_; 
wire u3__abc_74070_new_n647_; 
wire u3__abc_74070_new_n648_; 
wire u3__abc_74070_new_n650_; 
wire u3__abc_74070_new_n651_; 
wire u3__abc_74070_new_n652_; 
wire u3__abc_74070_new_n653_; 
wire u3__abc_74070_new_n654_; 
wire u3__abc_74070_new_n656_; 
wire u3__abc_74070_new_n657_; 
wire u3__abc_74070_new_n658_; 
wire u3__abc_74070_new_n659_; 
wire u3__abc_74070_new_n660_; 
wire u3__abc_74070_new_n662_; 
wire u3__abc_74070_new_n663_; 
wire u3__abc_74070_new_n664_; 
wire u3__abc_74070_new_n665_; 
wire u3__abc_74070_new_n666_; 
wire u3__abc_74070_new_n668_; 
wire u3__abc_74070_new_n669_; 
wire u3__abc_74070_new_n670_; 
wire u3__abc_74070_new_n671_; 
wire u3__abc_74070_new_n672_; 
wire u3__abc_74070_new_n674_; 
wire u3__abc_74070_new_n675_; 
wire u3__abc_74070_new_n676_; 
wire u3__abc_74070_new_n677_; 
wire u3__abc_74070_new_n678_; 
wire u3__abc_74070_new_n680_; 
wire u3__abc_74070_new_n681_; 
wire u3__abc_74070_new_n682_; 
wire u3__abc_74070_new_n683_; 
wire u3__abc_74070_new_n684_; 
wire u3__abc_74070_new_n686_; 
wire u3__abc_74070_new_n687_; 
wire u3__abc_74070_new_n688_; 
wire u3__abc_74070_new_n689_; 
wire u3__abc_74070_new_n690_; 
wire u3__abc_74070_new_n692_; 
wire u3__abc_74070_new_n693_; 
wire u3__abc_74070_new_n694_; 
wire u3__abc_74070_new_n695_; 
wire u3__abc_74070_new_n696_; 
wire u3__abc_74070_new_n698_; 
wire u3__abc_74070_new_n699_; 
wire u3__abc_74070_new_n700_; 
wire u3__abc_74070_new_n701_; 
wire u3__abc_74070_new_n702_; 
wire u3__abc_74070_new_n704_; 
wire u3__abc_74070_new_n705_; 
wire u3__abc_74070_new_n706_; 
wire u3__abc_74070_new_n707_; 
wire u3__abc_74070_new_n708_; 
wire u3__abc_74070_new_n710_; 
wire u3__abc_74070_new_n711_; 
wire u3__abc_74070_new_n712_; 
wire u3__abc_74070_new_n713_; 
wire u3__abc_74070_new_n714_; 
wire u3__abc_74070_new_n716_; 
wire u3__abc_74070_new_n717_; 
wire u3__abc_74070_new_n718_; 
wire u3__abc_74070_new_n719_; 
wire u3__abc_74070_new_n720_; 
wire u3__abc_74070_new_n722_; 
wire u3__abc_74070_new_n723_; 
wire u3__abc_74070_new_n724_; 
wire u3__abc_74070_new_n725_; 
wire u3__abc_74070_new_n726_; 
wire u3__abc_74070_new_n727_; 
wire u3__abc_74070_new_n728_; 
wire u3__abc_74070_new_n730_; 
wire u3__abc_74070_new_n731_; 
wire u3__abc_74070_new_n732_; 
wire u3__abc_74070_new_n733_; 
wire u3__abc_74070_new_n734_; 
wire u3__abc_74070_new_n735_; 
wire u3__abc_74070_new_n736_; 
wire u3__abc_74070_new_n738_; 
wire u3__abc_74070_new_n739_; 
wire u3__abc_74070_new_n740_; 
wire u3__abc_74070_new_n741_; 
wire u3__abc_74070_new_n742_; 
wire u3__abc_74070_new_n743_; 
wire u3__abc_74070_new_n744_; 
wire u3__abc_74070_new_n746_; 
wire u3__abc_74070_new_n747_; 
wire u3__abc_74070_new_n748_; 
wire u3__abc_74070_new_n749_; 
wire u3__abc_74070_new_n750_; 
wire u3__abc_74070_new_n751_; 
wire u3__abc_74070_new_n752_; 
wire u3__abc_74070_new_n754_; 
wire u3__abc_74070_new_n755_; 
wire u3__abc_74070_new_n756_; 
wire u3__abc_74070_new_n757_; 
wire u3__abc_74070_new_n758_; 
wire u3__abc_74070_new_n759_; 
wire u3__abc_74070_new_n760_; 
wire u3__abc_74070_new_n762_; 
wire u3__abc_74070_new_n763_; 
wire u3__abc_74070_new_n764_; 
wire u3__abc_74070_new_n765_; 
wire u3__abc_74070_new_n766_; 
wire u3__abc_74070_new_n767_; 
wire u3__abc_74070_new_n768_; 
wire u3__abc_74070_new_n770_; 
wire u3__abc_74070_new_n771_; 
wire u3__abc_74070_new_n772_; 
wire u3__abc_74070_new_n773_; 
wire u3__abc_74070_new_n774_; 
wire u3__abc_74070_new_n775_; 
wire u3__abc_74070_new_n776_; 
wire u3__abc_74070_new_n778_; 
wire u3__abc_74070_new_n779_; 
wire u3__abc_74070_new_n780_; 
wire u3__abc_74070_new_n781_; 
wire u3__abc_74070_new_n782_; 
wire u3__abc_74070_new_n783_; 
wire u3__abc_74070_new_n784_; 
wire u3__abc_74070_new_n786_; 
wire u3__abc_74070_new_n787_; 
wire u3__abc_74070_new_n788_; 
wire u3__abc_74070_new_n789_; 
wire u3__abc_74070_new_n790_; 
wire u3__abc_74070_new_n791_; 
wire u3__abc_74070_new_n792_; 
wire u3__abc_74070_new_n794_; 
wire u3__abc_74070_new_n795_; 
wire u3__abc_74070_new_n796_; 
wire u3__abc_74070_new_n797_; 
wire u3__abc_74070_new_n798_; 
wire u3__abc_74070_new_n799_; 
wire u3__abc_74070_new_n800_; 
wire u3__abc_74070_new_n802_; 
wire u3__abc_74070_new_n803_; 
wire u3__abc_74070_new_n804_; 
wire u3__abc_74070_new_n805_; 
wire u3__abc_74070_new_n806_; 
wire u3__abc_74070_new_n807_; 
wire u3__abc_74070_new_n808_; 
wire u3__abc_74070_new_n810_; 
wire u3__abc_74070_new_n811_; 
wire u3__abc_74070_new_n812_; 
wire u3__abc_74070_new_n813_; 
wire u3__abc_74070_new_n814_; 
wire u3__abc_74070_new_n815_; 
wire u3__abc_74070_new_n816_; 
wire u3__abc_74070_new_n818_; 
wire u3__abc_74070_new_n819_; 
wire u3__abc_74070_new_n820_; 
wire u3__abc_74070_new_n821_; 
wire u3__abc_74070_new_n822_; 
wire u3__abc_74070_new_n823_; 
wire u3__abc_74070_new_n824_; 
wire u3__abc_74070_new_n826_; 
wire u3__abc_74070_new_n827_; 
wire u3__abc_74070_new_n828_; 
wire u3__abc_74070_new_n829_; 
wire u3__abc_74070_new_n830_; 
wire u3__abc_74070_new_n831_; 
wire u3__abc_74070_new_n832_; 
wire u3__abc_74070_new_n834_; 
wire u3__abc_74070_new_n835_; 
wire u3__abc_74070_new_n836_; 
wire u3__abc_74070_new_n837_; 
wire u3__abc_74070_new_n838_; 
wire u3__abc_74070_new_n839_; 
wire u3__abc_74070_new_n840_; 
wire u3__abc_74070_new_n842_; 
wire u3__abc_74070_new_n843_; 
wire u3__abc_74070_new_n844_; 
wire u3__abc_74070_new_n845_; 
wire u3__abc_74070_new_n846_; 
wire u3__abc_74070_new_n847_; 
wire u3__abc_74070_new_n848_; 
wire u3__abc_74070_new_n850_; 
wire u3__abc_74070_new_n851_; 
wire u3__abc_74070_new_n854_; 
wire u3__abc_74070_new_n855_; 
wire u3__abc_74070_new_n856_; 
wire u3__abc_74070_new_n857_; 
wire u3__abc_74070_new_n858_; 
wire u3__abc_74070_new_n859_; 
wire u3__abc_74070_new_n860_; 
wire u3__abc_74070_new_n861_; 
wire u3__abc_74070_new_n862_; 
wire u3__abc_74070_new_n863_; 
wire u3__abc_74070_new_n864_; 
wire u3__abc_74070_new_n865_; 
wire u3__abc_74070_new_n866_; 
wire u3__abc_74070_new_n867_; 
wire u3__abc_74070_new_n868_; 
wire u3__abc_74070_new_n869_; 
wire u3__abc_74070_new_n870_; 
wire u3__abc_74070_new_n871_; 
wire u3__abc_74070_new_n872_; 
wire u3__abc_74070_new_n873_; 
wire u3__abc_74070_new_n874_; 
wire u3__abc_74070_new_n875_; 
wire u3__abc_74070_new_n876_; 
wire u3__abc_74070_new_n877_; 
wire u3__abc_74070_new_n878_; 
wire u3__abc_74070_new_n879_; 
wire u3__abc_74070_new_n880_; 
wire u3__abc_74070_new_n881_; 
wire u3__abc_74070_new_n882_; 
wire u3__abc_74070_new_n883_; 
wire u3__abc_74070_new_n884_; 
wire u3__abc_74070_new_n885_; 
wire u3__abc_74070_new_n886_; 
wire u3__abc_74070_new_n887_; 
wire u3__abc_74070_new_n888_; 
wire u3__abc_74070_new_n889_; 
wire u3__abc_74070_new_n890_; 
wire u3__abc_74070_new_n891_; 
wire u3__abc_74070_new_n892_; 
wire u3__abc_74070_new_n893_; 
wire u3__abc_74070_new_n894_; 
wire u3__abc_74070_new_n895_; 
wire u3__abc_74070_new_n896_; 
wire u3__abc_74070_new_n897_; 
wire u3__abc_74070_new_n898_; 
wire u3__abc_74070_new_n899_; 
wire u3__abc_74070_new_n900_; 
wire u3__abc_74070_new_n901_; 
wire u3__abc_74070_new_n902_; 
wire u3__abc_74070_new_n903_; 
wire u3__abc_74070_new_n904_; 
wire u3__abc_74070_new_n905_; 
wire u3__abc_74070_new_n906_; 
wire u3__abc_74070_new_n907_; 
wire u3__abc_74070_new_n908_; 
wire u3__abc_74070_new_n909_; 
wire u3__abc_74070_new_n910_; 
wire u3__abc_74070_new_n911_; 
wire u3__abc_74070_new_n912_; 
wire u3__abc_74070_new_n913_; 
wire u3__abc_74070_new_n914_; 
wire u3__abc_74070_new_n915_; 
wire u3__abc_74070_new_n916_; 
wire u3__abc_74070_new_n917_; 
wire u3__abc_74070_new_n918_; 
wire u3__abc_74070_new_n919_; 
wire u3__abc_74070_new_n920_; 
wire u3__abc_74070_new_n921_; 
wire u3__abc_74070_new_n922_; 
wire u3__abc_74070_new_n923_; 
wire u3__abc_74070_new_n924_; 
wire u3__abc_74070_new_n925_; 
wire u3__abc_74070_new_n926_; 
wire u3__abc_74070_new_n927_; 
wire u3__abc_74070_new_n928_; 
wire u3__abc_74070_new_n929_; 
wire u3__abc_74070_new_n930_; 
wire u3__abc_74070_new_n931_; 
wire u3__abc_74070_new_n932_; 
wire u3__abc_74070_new_n933_; 
wire u3__abc_74070_new_n934_; 
wire u3__abc_74070_new_n935_; 
wire u3__abc_74070_new_n936_; 
wire u3__abc_74070_new_n937_; 
wire u3__abc_74070_new_n938_; 
wire u3__abc_74070_new_n939_; 
wire u3__abc_74070_new_n940_; 
wire u3__abc_74070_new_n941_; 
wire u3__abc_74070_new_n942_; 
wire u3__abc_74070_new_n943_; 
wire u3__abc_74070_new_n944_; 
wire u3__abc_74070_new_n945_; 
wire u3__abc_74070_new_n946_; 
wire u3__abc_74070_new_n947_; 
wire u3__abc_74070_new_n948_; 
wire u3__abc_74070_new_n949_; 
wire u3__abc_74070_new_n950_; 
wire u3__abc_74070_new_n951_; 
wire u3__abc_74070_new_n952_; 
wire u3__abc_74070_new_n953_; 
wire u3__abc_74070_new_n954_; 
wire u3__abc_74070_new_n955_; 
wire u3__abc_74070_new_n956_; 
wire u3__abc_74070_new_n957_; 
wire u3__abc_74070_new_n958_; 
wire u3__abc_74070_new_n959_; 
wire u3__abc_74070_new_n960_; 
wire u3__abc_74070_new_n961_; 
wire u3__abc_74070_new_n962_; 
wire u3__abc_74070_new_n963_; 
wire u3__abc_74070_new_n964_; 
wire u3__abc_74070_new_n965_; 
wire u3__abc_74070_new_n966_; 
wire u3__abc_74070_new_n967_; 
wire u3__abc_74070_new_n968_; 
wire u3__abc_74070_new_n969_; 
wire u3__abc_74070_new_n970_; 
wire u3__abc_74070_new_n971_; 
wire u3__abc_74070_new_n972_; 
wire u3__abc_74070_new_n973_; 
wire u3__abc_74070_new_n974_; 
wire u3__abc_74070_new_n975_; 
wire u3__abc_74070_new_n976_; 
wire u3__abc_74070_new_n977_; 
wire u3__abc_74070_new_n978_; 
wire u3__abc_74070_new_n979_; 
wire u3__abc_74070_new_n980_; 
wire u3__abc_74070_new_n981_; 
wire u3__abc_74070_new_n982_; 
wire u3__abc_74070_new_n983_; 
wire u3__abc_74070_new_n984_; 
wire u3__abc_74070_new_n985_; 
wire u3__abc_74070_new_n986_; 
wire u3__abc_74070_new_n987_; 
wire u3__abc_74070_new_n988_; 
wire u3__abc_74070_new_n989_; 
wire u3__abc_74070_new_n990_; 
wire u3__abc_74070_new_n991_; 
wire u3__abc_74070_new_n992_; 
wire u3__abc_74070_new_n993_; 
wire u3__abc_74070_new_n994_; 
wire u3__abc_74070_new_n995_; 
wire u3__abc_74070_new_n996_; 
wire u3__abc_74070_new_n997_; 
wire u3__abc_74070_new_n998_; 
wire u3__abc_74070_new_n999_; 
wire u3_byte0_0_; 
wire u3_byte0_1_; 
wire u3_byte0_2_; 
wire u3_byte0_3_; 
wire u3_byte0_4_; 
wire u3_byte0_5_; 
wire u3_byte0_6_; 
wire u3_byte0_7_; 
wire u3_byte1_0_; 
wire u3_byte1_1_; 
wire u3_byte1_2_; 
wire u3_byte1_3_; 
wire u3_byte1_4_; 
wire u3_byte1_5_; 
wire u3_byte1_6_; 
wire u3_byte1_7_; 
wire u3_byte2_0_; 
wire u3_byte2_1_; 
wire u3_byte2_2_; 
wire u3_byte2_3_; 
wire u3_byte2_4_; 
wire u3_byte2_5_; 
wire u3_byte2_6_; 
wire u3_byte2_7_; 
wire u3_pen; 
wire u3_rd_fifo_clr; 
wire u3_rd_fifo_out_0_; 
wire u3_rd_fifo_out_10_; 
wire u3_rd_fifo_out_11_; 
wire u3_rd_fifo_out_12_; 
wire u3_rd_fifo_out_13_; 
wire u3_rd_fifo_out_14_; 
wire u3_rd_fifo_out_15_; 
wire u3_rd_fifo_out_16_; 
wire u3_rd_fifo_out_17_; 
wire u3_rd_fifo_out_18_; 
wire u3_rd_fifo_out_19_; 
wire u3_rd_fifo_out_1_; 
wire u3_rd_fifo_out_20_; 
wire u3_rd_fifo_out_21_; 
wire u3_rd_fifo_out_22_; 
wire u3_rd_fifo_out_23_; 
wire u3_rd_fifo_out_24_; 
wire u3_rd_fifo_out_25_; 
wire u3_rd_fifo_out_26_; 
wire u3_rd_fifo_out_27_; 
wire u3_rd_fifo_out_28_; 
wire u3_rd_fifo_out_29_; 
wire u3_rd_fifo_out_2_; 
wire u3_rd_fifo_out_30_; 
wire u3_rd_fifo_out_31_; 
wire u3_rd_fifo_out_32_; 
wire u3_rd_fifo_out_33_; 
wire u3_rd_fifo_out_34_; 
wire u3_rd_fifo_out_35_; 
wire u3_rd_fifo_out_3_; 
wire u3_rd_fifo_out_4_; 
wire u3_rd_fifo_out_5_; 
wire u3_rd_fifo_out_6_; 
wire u3_rd_fifo_out_7_; 
wire u3_rd_fifo_out_8_; 
wire u3_rd_fifo_out_9_; 
wire u3_re; 
wire u3_u0__0r0_35_0__0_; 
wire u3_u0__0r0_35_0__10_; 
wire u3_u0__0r0_35_0__11_; 
wire u3_u0__0r0_35_0__12_; 
wire u3_u0__0r0_35_0__13_; 
wire u3_u0__0r0_35_0__14_; 
wire u3_u0__0r0_35_0__15_; 
wire u3_u0__0r0_35_0__16_; 
wire u3_u0__0r0_35_0__17_; 
wire u3_u0__0r0_35_0__18_; 
wire u3_u0__0r0_35_0__19_; 
wire u3_u0__0r0_35_0__1_; 
wire u3_u0__0r0_35_0__20_; 
wire u3_u0__0r0_35_0__21_; 
wire u3_u0__0r0_35_0__22_; 
wire u3_u0__0r0_35_0__23_; 
wire u3_u0__0r0_35_0__24_; 
wire u3_u0__0r0_35_0__25_; 
wire u3_u0__0r0_35_0__26_; 
wire u3_u0__0r0_35_0__27_; 
wire u3_u0__0r0_35_0__28_; 
wire u3_u0__0r0_35_0__29_; 
wire u3_u0__0r0_35_0__2_; 
wire u3_u0__0r0_35_0__30_; 
wire u3_u0__0r0_35_0__31_; 
wire u3_u0__0r0_35_0__32_; 
wire u3_u0__0r0_35_0__33_; 
wire u3_u0__0r0_35_0__34_; 
wire u3_u0__0r0_35_0__35_; 
wire u3_u0__0r0_35_0__3_; 
wire u3_u0__0r0_35_0__4_; 
wire u3_u0__0r0_35_0__5_; 
wire u3_u0__0r0_35_0__6_; 
wire u3_u0__0r0_35_0__7_; 
wire u3_u0__0r0_35_0__8_; 
wire u3_u0__0r0_35_0__9_; 
wire u3_u0__0r1_35_0__0_; 
wire u3_u0__0r1_35_0__10_; 
wire u3_u0__0r1_35_0__11_; 
wire u3_u0__0r1_35_0__12_; 
wire u3_u0__0r1_35_0__13_; 
wire u3_u0__0r1_35_0__14_; 
wire u3_u0__0r1_35_0__15_; 
wire u3_u0__0r1_35_0__16_; 
wire u3_u0__0r1_35_0__17_; 
wire u3_u0__0r1_35_0__18_; 
wire u3_u0__0r1_35_0__19_; 
wire u3_u0__0r1_35_0__1_; 
wire u3_u0__0r1_35_0__20_; 
wire u3_u0__0r1_35_0__21_; 
wire u3_u0__0r1_35_0__22_; 
wire u3_u0__0r1_35_0__23_; 
wire u3_u0__0r1_35_0__24_; 
wire u3_u0__0r1_35_0__25_; 
wire u3_u0__0r1_35_0__26_; 
wire u3_u0__0r1_35_0__27_; 
wire u3_u0__0r1_35_0__28_; 
wire u3_u0__0r1_35_0__29_; 
wire u3_u0__0r1_35_0__2_; 
wire u3_u0__0r1_35_0__30_; 
wire u3_u0__0r1_35_0__31_; 
wire u3_u0__0r1_35_0__32_; 
wire u3_u0__0r1_35_0__33_; 
wire u3_u0__0r1_35_0__34_; 
wire u3_u0__0r1_35_0__35_; 
wire u3_u0__0r1_35_0__3_; 
wire u3_u0__0r1_35_0__4_; 
wire u3_u0__0r1_35_0__5_; 
wire u3_u0__0r1_35_0__6_; 
wire u3_u0__0r1_35_0__7_; 
wire u3_u0__0r1_35_0__8_; 
wire u3_u0__0r1_35_0__9_; 
wire u3_u0__0r2_35_0__0_; 
wire u3_u0__0r2_35_0__10_; 
wire u3_u0__0r2_35_0__11_; 
wire u3_u0__0r2_35_0__12_; 
wire u3_u0__0r2_35_0__13_; 
wire u3_u0__0r2_35_0__14_; 
wire u3_u0__0r2_35_0__15_; 
wire u3_u0__0r2_35_0__16_; 
wire u3_u0__0r2_35_0__17_; 
wire u3_u0__0r2_35_0__18_; 
wire u3_u0__0r2_35_0__19_; 
wire u3_u0__0r2_35_0__1_; 
wire u3_u0__0r2_35_0__20_; 
wire u3_u0__0r2_35_0__21_; 
wire u3_u0__0r2_35_0__22_; 
wire u3_u0__0r2_35_0__23_; 
wire u3_u0__0r2_35_0__24_; 
wire u3_u0__0r2_35_0__25_; 
wire u3_u0__0r2_35_0__26_; 
wire u3_u0__0r2_35_0__27_; 
wire u3_u0__0r2_35_0__28_; 
wire u3_u0__0r2_35_0__29_; 
wire u3_u0__0r2_35_0__2_; 
wire u3_u0__0r2_35_0__30_; 
wire u3_u0__0r2_35_0__31_; 
wire u3_u0__0r2_35_0__32_; 
wire u3_u0__0r2_35_0__33_; 
wire u3_u0__0r2_35_0__34_; 
wire u3_u0__0r2_35_0__35_; 
wire u3_u0__0r2_35_0__3_; 
wire u3_u0__0r2_35_0__4_; 
wire u3_u0__0r2_35_0__5_; 
wire u3_u0__0r2_35_0__6_; 
wire u3_u0__0r2_35_0__7_; 
wire u3_u0__0r2_35_0__8_; 
wire u3_u0__0r2_35_0__9_; 
wire u3_u0__0r3_35_0__0_; 
wire u3_u0__0r3_35_0__10_; 
wire u3_u0__0r3_35_0__11_; 
wire u3_u0__0r3_35_0__12_; 
wire u3_u0__0r3_35_0__13_; 
wire u3_u0__0r3_35_0__14_; 
wire u3_u0__0r3_35_0__15_; 
wire u3_u0__0r3_35_0__16_; 
wire u3_u0__0r3_35_0__17_; 
wire u3_u0__0r3_35_0__18_; 
wire u3_u0__0r3_35_0__19_; 
wire u3_u0__0r3_35_0__1_; 
wire u3_u0__0r3_35_0__20_; 
wire u3_u0__0r3_35_0__21_; 
wire u3_u0__0r3_35_0__22_; 
wire u3_u0__0r3_35_0__23_; 
wire u3_u0__0r3_35_0__24_; 
wire u3_u0__0r3_35_0__25_; 
wire u3_u0__0r3_35_0__26_; 
wire u3_u0__0r3_35_0__27_; 
wire u3_u0__0r3_35_0__28_; 
wire u3_u0__0r3_35_0__29_; 
wire u3_u0__0r3_35_0__2_; 
wire u3_u0__0r3_35_0__30_; 
wire u3_u0__0r3_35_0__31_; 
wire u3_u0__0r3_35_0__32_; 
wire u3_u0__0r3_35_0__33_; 
wire u3_u0__0r3_35_0__34_; 
wire u3_u0__0r3_35_0__35_; 
wire u3_u0__0r3_35_0__3_; 
wire u3_u0__0r3_35_0__4_; 
wire u3_u0__0r3_35_0__5_; 
wire u3_u0__0r3_35_0__6_; 
wire u3_u0__0r3_35_0__7_; 
wire u3_u0__0r3_35_0__8_; 
wire u3_u0__0r3_35_0__9_; 
wire u3_u0__0rd_adr_3_0__0_; 
wire u3_u0__0rd_adr_3_0__1_; 
wire u3_u0__0rd_adr_3_0__2_; 
wire u3_u0__0rd_adr_3_0__3_; 
wire u3_u0__0wr_adr_3_0__0_; 
wire u3_u0__0wr_adr_3_0__1_; 
wire u3_u0__0wr_adr_3_0__2_; 
wire u3_u0__0wr_adr_3_0__3_; 
wire u3_u0__abc_75526_auto_rtlil_cc_1942_NotGate_71546; 
wire u3_u0__abc_75526_new_n1001_; 
wire u3_u0__abc_75526_new_n1002_; 
wire u3_u0__abc_75526_new_n1003_; 
wire u3_u0__abc_75526_new_n1005_; 
wire u3_u0__abc_75526_new_n1006_; 
wire u3_u0__abc_75526_new_n1007_; 
wire u3_u0__abc_75526_new_n1009_; 
wire u3_u0__abc_75526_new_n1010_; 
wire u3_u0__abc_75526_new_n1011_; 
wire u3_u0__abc_75526_new_n1013_; 
wire u3_u0__abc_75526_new_n1014_; 
wire u3_u0__abc_75526_new_n1015_; 
wire u3_u0__abc_75526_new_n1017_; 
wire u3_u0__abc_75526_new_n1018_; 
wire u3_u0__abc_75526_new_n1019_; 
wire u3_u0__abc_75526_new_n1021_; 
wire u3_u0__abc_75526_new_n1022_; 
wire u3_u0__abc_75526_new_n1023_; 
wire u3_u0__abc_75526_new_n1025_; 
wire u3_u0__abc_75526_new_n1026_; 
wire u3_u0__abc_75526_new_n1027_; 
wire u3_u0__abc_75526_new_n1029_; 
wire u3_u0__abc_75526_new_n1030_; 
wire u3_u0__abc_75526_new_n1031_; 
wire u3_u0__abc_75526_new_n1032_; 
wire u3_u0__abc_75526_new_n1033_; 
wire u3_u0__abc_75526_new_n1034_; 
wire u3_u0__abc_75526_new_n1034__bF_buf0; 
wire u3_u0__abc_75526_new_n1034__bF_buf1; 
wire u3_u0__abc_75526_new_n1034__bF_buf2; 
wire u3_u0__abc_75526_new_n1034__bF_buf3; 
wire u3_u0__abc_75526_new_n1034__bF_buf4; 
wire u3_u0__abc_75526_new_n1034__bF_buf5; 
wire u3_u0__abc_75526_new_n1035_; 
wire u3_u0__abc_75526_new_n1036_; 
wire u3_u0__abc_75526_new_n1037_; 
wire u3_u0__abc_75526_new_n1038_; 
wire u3_u0__abc_75526_new_n1039_; 
wire u3_u0__abc_75526_new_n1040_; 
wire u3_u0__abc_75526_new_n1041_; 
wire u3_u0__abc_75526_new_n1042_; 
wire u3_u0__abc_75526_new_n1043_; 
wire u3_u0__abc_75526_new_n1043__bF_buf0; 
wire u3_u0__abc_75526_new_n1043__bF_buf1; 
wire u3_u0__abc_75526_new_n1043__bF_buf2; 
wire u3_u0__abc_75526_new_n1043__bF_buf3; 
wire u3_u0__abc_75526_new_n1043__bF_buf4; 
wire u3_u0__abc_75526_new_n1043__bF_buf5; 
wire u3_u0__abc_75526_new_n1044_; 
wire u3_u0__abc_75526_new_n1045_; 
wire u3_u0__abc_75526_new_n1046_; 
wire u3_u0__abc_75526_new_n1047_; 
wire u3_u0__abc_75526_new_n1048_; 
wire u3_u0__abc_75526_new_n1049_; 
wire u3_u0__abc_75526_new_n1049__bF_buf0; 
wire u3_u0__abc_75526_new_n1049__bF_buf1; 
wire u3_u0__abc_75526_new_n1049__bF_buf2; 
wire u3_u0__abc_75526_new_n1049__bF_buf3; 
wire u3_u0__abc_75526_new_n1049__bF_buf4; 
wire u3_u0__abc_75526_new_n1049__bF_buf5; 
wire u3_u0__abc_75526_new_n1050_; 
wire u3_u0__abc_75526_new_n1051_; 
wire u3_u0__abc_75526_new_n1052_; 
wire u3_u0__abc_75526_new_n1052__bF_buf0; 
wire u3_u0__abc_75526_new_n1052__bF_buf1; 
wire u3_u0__abc_75526_new_n1052__bF_buf2; 
wire u3_u0__abc_75526_new_n1052__bF_buf3; 
wire u3_u0__abc_75526_new_n1052__bF_buf4; 
wire u3_u0__abc_75526_new_n1052__bF_buf5; 
wire u3_u0__abc_75526_new_n1053_; 
wire u3_u0__abc_75526_new_n1054_; 
wire u3_u0__abc_75526_new_n1055_; 
wire u3_u0__abc_75526_new_n1057_; 
wire u3_u0__abc_75526_new_n1058_; 
wire u3_u0__abc_75526_new_n1059_; 
wire u3_u0__abc_75526_new_n1060_; 
wire u3_u0__abc_75526_new_n1061_; 
wire u3_u0__abc_75526_new_n1062_; 
wire u3_u0__abc_75526_new_n1064_; 
wire u3_u0__abc_75526_new_n1065_; 
wire u3_u0__abc_75526_new_n1066_; 
wire u3_u0__abc_75526_new_n1067_; 
wire u3_u0__abc_75526_new_n1068_; 
wire u3_u0__abc_75526_new_n1069_; 
wire u3_u0__abc_75526_new_n1071_; 
wire u3_u0__abc_75526_new_n1072_; 
wire u3_u0__abc_75526_new_n1073_; 
wire u3_u0__abc_75526_new_n1074_; 
wire u3_u0__abc_75526_new_n1075_; 
wire u3_u0__abc_75526_new_n1076_; 
wire u3_u0__abc_75526_new_n1078_; 
wire u3_u0__abc_75526_new_n1079_; 
wire u3_u0__abc_75526_new_n1080_; 
wire u3_u0__abc_75526_new_n1081_; 
wire u3_u0__abc_75526_new_n1082_; 
wire u3_u0__abc_75526_new_n1083_; 
wire u3_u0__abc_75526_new_n1085_; 
wire u3_u0__abc_75526_new_n1086_; 
wire u3_u0__abc_75526_new_n1087_; 
wire u3_u0__abc_75526_new_n1088_; 
wire u3_u0__abc_75526_new_n1089_; 
wire u3_u0__abc_75526_new_n1090_; 
wire u3_u0__abc_75526_new_n1092_; 
wire u3_u0__abc_75526_new_n1093_; 
wire u3_u0__abc_75526_new_n1094_; 
wire u3_u0__abc_75526_new_n1095_; 
wire u3_u0__abc_75526_new_n1096_; 
wire u3_u0__abc_75526_new_n1097_; 
wire u3_u0__abc_75526_new_n1099_; 
wire u3_u0__abc_75526_new_n1100_; 
wire u3_u0__abc_75526_new_n1101_; 
wire u3_u0__abc_75526_new_n1102_; 
wire u3_u0__abc_75526_new_n1103_; 
wire u3_u0__abc_75526_new_n1104_; 
wire u3_u0__abc_75526_new_n1106_; 
wire u3_u0__abc_75526_new_n1107_; 
wire u3_u0__abc_75526_new_n1108_; 
wire u3_u0__abc_75526_new_n1109_; 
wire u3_u0__abc_75526_new_n1110_; 
wire u3_u0__abc_75526_new_n1111_; 
wire u3_u0__abc_75526_new_n1113_; 
wire u3_u0__abc_75526_new_n1114_; 
wire u3_u0__abc_75526_new_n1115_; 
wire u3_u0__abc_75526_new_n1116_; 
wire u3_u0__abc_75526_new_n1117_; 
wire u3_u0__abc_75526_new_n1118_; 
wire u3_u0__abc_75526_new_n1120_; 
wire u3_u0__abc_75526_new_n1121_; 
wire u3_u0__abc_75526_new_n1122_; 
wire u3_u0__abc_75526_new_n1123_; 
wire u3_u0__abc_75526_new_n1124_; 
wire u3_u0__abc_75526_new_n1125_; 
wire u3_u0__abc_75526_new_n1127_; 
wire u3_u0__abc_75526_new_n1128_; 
wire u3_u0__abc_75526_new_n1129_; 
wire u3_u0__abc_75526_new_n1130_; 
wire u3_u0__abc_75526_new_n1131_; 
wire u3_u0__abc_75526_new_n1132_; 
wire u3_u0__abc_75526_new_n1134_; 
wire u3_u0__abc_75526_new_n1135_; 
wire u3_u0__abc_75526_new_n1136_; 
wire u3_u0__abc_75526_new_n1137_; 
wire u3_u0__abc_75526_new_n1138_; 
wire u3_u0__abc_75526_new_n1139_; 
wire u3_u0__abc_75526_new_n1141_; 
wire u3_u0__abc_75526_new_n1142_; 
wire u3_u0__abc_75526_new_n1143_; 
wire u3_u0__abc_75526_new_n1144_; 
wire u3_u0__abc_75526_new_n1145_; 
wire u3_u0__abc_75526_new_n1146_; 
wire u3_u0__abc_75526_new_n1148_; 
wire u3_u0__abc_75526_new_n1149_; 
wire u3_u0__abc_75526_new_n1150_; 
wire u3_u0__abc_75526_new_n1151_; 
wire u3_u0__abc_75526_new_n1152_; 
wire u3_u0__abc_75526_new_n1153_; 
wire u3_u0__abc_75526_new_n1155_; 
wire u3_u0__abc_75526_new_n1156_; 
wire u3_u0__abc_75526_new_n1157_; 
wire u3_u0__abc_75526_new_n1158_; 
wire u3_u0__abc_75526_new_n1159_; 
wire u3_u0__abc_75526_new_n1160_; 
wire u3_u0__abc_75526_new_n1162_; 
wire u3_u0__abc_75526_new_n1163_; 
wire u3_u0__abc_75526_new_n1164_; 
wire u3_u0__abc_75526_new_n1165_; 
wire u3_u0__abc_75526_new_n1166_; 
wire u3_u0__abc_75526_new_n1167_; 
wire u3_u0__abc_75526_new_n1169_; 
wire u3_u0__abc_75526_new_n1170_; 
wire u3_u0__abc_75526_new_n1171_; 
wire u3_u0__abc_75526_new_n1172_; 
wire u3_u0__abc_75526_new_n1173_; 
wire u3_u0__abc_75526_new_n1174_; 
wire u3_u0__abc_75526_new_n1176_; 
wire u3_u0__abc_75526_new_n1177_; 
wire u3_u0__abc_75526_new_n1178_; 
wire u3_u0__abc_75526_new_n1179_; 
wire u3_u0__abc_75526_new_n1180_; 
wire u3_u0__abc_75526_new_n1181_; 
wire u3_u0__abc_75526_new_n1183_; 
wire u3_u0__abc_75526_new_n1184_; 
wire u3_u0__abc_75526_new_n1185_; 
wire u3_u0__abc_75526_new_n1186_; 
wire u3_u0__abc_75526_new_n1187_; 
wire u3_u0__abc_75526_new_n1188_; 
wire u3_u0__abc_75526_new_n1190_; 
wire u3_u0__abc_75526_new_n1191_; 
wire u3_u0__abc_75526_new_n1192_; 
wire u3_u0__abc_75526_new_n1193_; 
wire u3_u0__abc_75526_new_n1194_; 
wire u3_u0__abc_75526_new_n1195_; 
wire u3_u0__abc_75526_new_n1197_; 
wire u3_u0__abc_75526_new_n1198_; 
wire u3_u0__abc_75526_new_n1199_; 
wire u3_u0__abc_75526_new_n1200_; 
wire u3_u0__abc_75526_new_n1201_; 
wire u3_u0__abc_75526_new_n1202_; 
wire u3_u0__abc_75526_new_n1204_; 
wire u3_u0__abc_75526_new_n1205_; 
wire u3_u0__abc_75526_new_n1206_; 
wire u3_u0__abc_75526_new_n1207_; 
wire u3_u0__abc_75526_new_n1208_; 
wire u3_u0__abc_75526_new_n1209_; 
wire u3_u0__abc_75526_new_n1211_; 
wire u3_u0__abc_75526_new_n1212_; 
wire u3_u0__abc_75526_new_n1213_; 
wire u3_u0__abc_75526_new_n1214_; 
wire u3_u0__abc_75526_new_n1215_; 
wire u3_u0__abc_75526_new_n1216_; 
wire u3_u0__abc_75526_new_n1218_; 
wire u3_u0__abc_75526_new_n1219_; 
wire u3_u0__abc_75526_new_n1220_; 
wire u3_u0__abc_75526_new_n1221_; 
wire u3_u0__abc_75526_new_n1222_; 
wire u3_u0__abc_75526_new_n1223_; 
wire u3_u0__abc_75526_new_n1225_; 
wire u3_u0__abc_75526_new_n1226_; 
wire u3_u0__abc_75526_new_n1227_; 
wire u3_u0__abc_75526_new_n1228_; 
wire u3_u0__abc_75526_new_n1229_; 
wire u3_u0__abc_75526_new_n1230_; 
wire u3_u0__abc_75526_new_n1232_; 
wire u3_u0__abc_75526_new_n1233_; 
wire u3_u0__abc_75526_new_n1234_; 
wire u3_u0__abc_75526_new_n1235_; 
wire u3_u0__abc_75526_new_n1236_; 
wire u3_u0__abc_75526_new_n1237_; 
wire u3_u0__abc_75526_new_n1239_; 
wire u3_u0__abc_75526_new_n1240_; 
wire u3_u0__abc_75526_new_n1241_; 
wire u3_u0__abc_75526_new_n1242_; 
wire u3_u0__abc_75526_new_n1243_; 
wire u3_u0__abc_75526_new_n1244_; 
wire u3_u0__abc_75526_new_n1246_; 
wire u3_u0__abc_75526_new_n1247_; 
wire u3_u0__abc_75526_new_n1248_; 
wire u3_u0__abc_75526_new_n1249_; 
wire u3_u0__abc_75526_new_n1250_; 
wire u3_u0__abc_75526_new_n1251_; 
wire u3_u0__abc_75526_new_n1253_; 
wire u3_u0__abc_75526_new_n1254_; 
wire u3_u0__abc_75526_new_n1255_; 
wire u3_u0__abc_75526_new_n1256_; 
wire u3_u0__abc_75526_new_n1257_; 
wire u3_u0__abc_75526_new_n1258_; 
wire u3_u0__abc_75526_new_n1260_; 
wire u3_u0__abc_75526_new_n1261_; 
wire u3_u0__abc_75526_new_n1262_; 
wire u3_u0__abc_75526_new_n1263_; 
wire u3_u0__abc_75526_new_n1264_; 
wire u3_u0__abc_75526_new_n1265_; 
wire u3_u0__abc_75526_new_n1267_; 
wire u3_u0__abc_75526_new_n1268_; 
wire u3_u0__abc_75526_new_n1269_; 
wire u3_u0__abc_75526_new_n1270_; 
wire u3_u0__abc_75526_new_n1271_; 
wire u3_u0__abc_75526_new_n1272_; 
wire u3_u0__abc_75526_new_n1274_; 
wire u3_u0__abc_75526_new_n1275_; 
wire u3_u0__abc_75526_new_n1276_; 
wire u3_u0__abc_75526_new_n1277_; 
wire u3_u0__abc_75526_new_n1278_; 
wire u3_u0__abc_75526_new_n1279_; 
wire u3_u0__abc_75526_new_n1281_; 
wire u3_u0__abc_75526_new_n1282_; 
wire u3_u0__abc_75526_new_n1283_; 
wire u3_u0__abc_75526_new_n1284_; 
wire u3_u0__abc_75526_new_n1285_; 
wire u3_u0__abc_75526_new_n1286_; 
wire u3_u0__abc_75526_new_n1288_; 
wire u3_u0__abc_75526_new_n1289_; 
wire u3_u0__abc_75526_new_n1290_; 
wire u3_u0__abc_75526_new_n1291_; 
wire u3_u0__abc_75526_new_n1292_; 
wire u3_u0__abc_75526_new_n1293_; 
wire u3_u0__abc_75526_new_n1295_; 
wire u3_u0__abc_75526_new_n1296_; 
wire u3_u0__abc_75526_new_n1297_; 
wire u3_u0__abc_75526_new_n1298_; 
wire u3_u0__abc_75526_new_n1299_; 
wire u3_u0__abc_75526_new_n1300_; 
wire u3_u0__abc_75526_new_n382_; 
wire u3_u0__abc_75526_new_n382__bF_buf0; 
wire u3_u0__abc_75526_new_n382__bF_buf1; 
wire u3_u0__abc_75526_new_n382__bF_buf2; 
wire u3_u0__abc_75526_new_n382__bF_buf3; 
wire u3_u0__abc_75526_new_n382__bF_buf4; 
wire u3_u0__abc_75526_new_n382__bF_buf5; 
wire u3_u0__abc_75526_new_n382__bF_buf6; 
wire u3_u0__abc_75526_new_n382__bF_buf7; 
wire u3_u0__abc_75526_new_n383_; 
wire u3_u0__abc_75526_new_n384_; 
wire u3_u0__abc_75526_new_n385_; 
wire u3_u0__abc_75526_new_n386_; 
wire u3_u0__abc_75526_new_n388_; 
wire u3_u0__abc_75526_new_n389_; 
wire u3_u0__abc_75526_new_n390_; 
wire u3_u0__abc_75526_new_n391_; 
wire u3_u0__abc_75526_new_n393_; 
wire u3_u0__abc_75526_new_n394_; 
wire u3_u0__abc_75526_new_n395_; 
wire u3_u0__abc_75526_new_n396_; 
wire u3_u0__abc_75526_new_n398_; 
wire u3_u0__abc_75526_new_n399_; 
wire u3_u0__abc_75526_new_n400_; 
wire u3_u0__abc_75526_new_n401_; 
wire u3_u0__abc_75526_new_n403_; 
wire u3_u0__abc_75526_new_n404_; 
wire u3_u0__abc_75526_new_n405_; 
wire u3_u0__abc_75526_new_n406_; 
wire u3_u0__abc_75526_new_n408_; 
wire u3_u0__abc_75526_new_n409_; 
wire u3_u0__abc_75526_new_n410_; 
wire u3_u0__abc_75526_new_n411_; 
wire u3_u0__abc_75526_new_n413_; 
wire u3_u0__abc_75526_new_n414_; 
wire u3_u0__abc_75526_new_n415_; 
wire u3_u0__abc_75526_new_n416_; 
wire u3_u0__abc_75526_new_n418_; 
wire u3_u0__abc_75526_new_n419_; 
wire u3_u0__abc_75526_new_n420_; 
wire u3_u0__abc_75526_new_n421_; 
wire u3_u0__abc_75526_new_n423_; 
wire u3_u0__abc_75526_new_n424_; 
wire u3_u0__abc_75526_new_n425_; 
wire u3_u0__abc_75526_new_n426_; 
wire u3_u0__abc_75526_new_n428_; 
wire u3_u0__abc_75526_new_n429_; 
wire u3_u0__abc_75526_new_n430_; 
wire u3_u0__abc_75526_new_n431_; 
wire u3_u0__abc_75526_new_n433_; 
wire u3_u0__abc_75526_new_n434_; 
wire u3_u0__abc_75526_new_n435_; 
wire u3_u0__abc_75526_new_n436_; 
wire u3_u0__abc_75526_new_n438_; 
wire u3_u0__abc_75526_new_n439_; 
wire u3_u0__abc_75526_new_n440_; 
wire u3_u0__abc_75526_new_n441_; 
wire u3_u0__abc_75526_new_n443_; 
wire u3_u0__abc_75526_new_n444_; 
wire u3_u0__abc_75526_new_n445_; 
wire u3_u0__abc_75526_new_n446_; 
wire u3_u0__abc_75526_new_n448_; 
wire u3_u0__abc_75526_new_n449_; 
wire u3_u0__abc_75526_new_n450_; 
wire u3_u0__abc_75526_new_n451_; 
wire u3_u0__abc_75526_new_n453_; 
wire u3_u0__abc_75526_new_n454_; 
wire u3_u0__abc_75526_new_n455_; 
wire u3_u0__abc_75526_new_n456_; 
wire u3_u0__abc_75526_new_n458_; 
wire u3_u0__abc_75526_new_n459_; 
wire u3_u0__abc_75526_new_n460_; 
wire u3_u0__abc_75526_new_n461_; 
wire u3_u0__abc_75526_new_n463_; 
wire u3_u0__abc_75526_new_n464_; 
wire u3_u0__abc_75526_new_n465_; 
wire u3_u0__abc_75526_new_n466_; 
wire u3_u0__abc_75526_new_n468_; 
wire u3_u0__abc_75526_new_n469_; 
wire u3_u0__abc_75526_new_n470_; 
wire u3_u0__abc_75526_new_n471_; 
wire u3_u0__abc_75526_new_n473_; 
wire u3_u0__abc_75526_new_n474_; 
wire u3_u0__abc_75526_new_n475_; 
wire u3_u0__abc_75526_new_n476_; 
wire u3_u0__abc_75526_new_n478_; 
wire u3_u0__abc_75526_new_n479_; 
wire u3_u0__abc_75526_new_n480_; 
wire u3_u0__abc_75526_new_n481_; 
wire u3_u0__abc_75526_new_n483_; 
wire u3_u0__abc_75526_new_n484_; 
wire u3_u0__abc_75526_new_n485_; 
wire u3_u0__abc_75526_new_n486_; 
wire u3_u0__abc_75526_new_n488_; 
wire u3_u0__abc_75526_new_n489_; 
wire u3_u0__abc_75526_new_n490_; 
wire u3_u0__abc_75526_new_n491_; 
wire u3_u0__abc_75526_new_n493_; 
wire u3_u0__abc_75526_new_n494_; 
wire u3_u0__abc_75526_new_n495_; 
wire u3_u0__abc_75526_new_n496_; 
wire u3_u0__abc_75526_new_n498_; 
wire u3_u0__abc_75526_new_n499_; 
wire u3_u0__abc_75526_new_n500_; 
wire u3_u0__abc_75526_new_n501_; 
wire u3_u0__abc_75526_new_n503_; 
wire u3_u0__abc_75526_new_n504_; 
wire u3_u0__abc_75526_new_n505_; 
wire u3_u0__abc_75526_new_n506_; 
wire u3_u0__abc_75526_new_n508_; 
wire u3_u0__abc_75526_new_n509_; 
wire u3_u0__abc_75526_new_n510_; 
wire u3_u0__abc_75526_new_n511_; 
wire u3_u0__abc_75526_new_n513_; 
wire u3_u0__abc_75526_new_n514_; 
wire u3_u0__abc_75526_new_n515_; 
wire u3_u0__abc_75526_new_n516_; 
wire u3_u0__abc_75526_new_n518_; 
wire u3_u0__abc_75526_new_n519_; 
wire u3_u0__abc_75526_new_n520_; 
wire u3_u0__abc_75526_new_n521_; 
wire u3_u0__abc_75526_new_n523_; 
wire u3_u0__abc_75526_new_n524_; 
wire u3_u0__abc_75526_new_n525_; 
wire u3_u0__abc_75526_new_n526_; 
wire u3_u0__abc_75526_new_n528_; 
wire u3_u0__abc_75526_new_n529_; 
wire u3_u0__abc_75526_new_n530_; 
wire u3_u0__abc_75526_new_n531_; 
wire u3_u0__abc_75526_new_n533_; 
wire u3_u0__abc_75526_new_n534_; 
wire u3_u0__abc_75526_new_n535_; 
wire u3_u0__abc_75526_new_n536_; 
wire u3_u0__abc_75526_new_n538_; 
wire u3_u0__abc_75526_new_n539_; 
wire u3_u0__abc_75526_new_n540_; 
wire u3_u0__abc_75526_new_n541_; 
wire u3_u0__abc_75526_new_n543_; 
wire u3_u0__abc_75526_new_n544_; 
wire u3_u0__abc_75526_new_n545_; 
wire u3_u0__abc_75526_new_n546_; 
wire u3_u0__abc_75526_new_n548_; 
wire u3_u0__abc_75526_new_n549_; 
wire u3_u0__abc_75526_new_n550_; 
wire u3_u0__abc_75526_new_n551_; 
wire u3_u0__abc_75526_new_n553_; 
wire u3_u0__abc_75526_new_n554_; 
wire u3_u0__abc_75526_new_n555_; 
wire u3_u0__abc_75526_new_n556_; 
wire u3_u0__abc_75526_new_n558_; 
wire u3_u0__abc_75526_new_n559_; 
wire u3_u0__abc_75526_new_n560_; 
wire u3_u0__abc_75526_new_n561_; 
wire u3_u0__abc_75526_new_n563_; 
wire u3_u0__abc_75526_new_n563__bF_buf0; 
wire u3_u0__abc_75526_new_n563__bF_buf1; 
wire u3_u0__abc_75526_new_n563__bF_buf2; 
wire u3_u0__abc_75526_new_n563__bF_buf3; 
wire u3_u0__abc_75526_new_n563__bF_buf4; 
wire u3_u0__abc_75526_new_n563__bF_buf5; 
wire u3_u0__abc_75526_new_n563__bF_buf6; 
wire u3_u0__abc_75526_new_n563__bF_buf7; 
wire u3_u0__abc_75526_new_n564_; 
wire u3_u0__abc_75526_new_n565_; 
wire u3_u0__abc_75526_new_n566_; 
wire u3_u0__abc_75526_new_n568_; 
wire u3_u0__abc_75526_new_n569_; 
wire u3_u0__abc_75526_new_n570_; 
wire u3_u0__abc_75526_new_n572_; 
wire u3_u0__abc_75526_new_n573_; 
wire u3_u0__abc_75526_new_n574_; 
wire u3_u0__abc_75526_new_n576_; 
wire u3_u0__abc_75526_new_n577_; 
wire u3_u0__abc_75526_new_n578_; 
wire u3_u0__abc_75526_new_n580_; 
wire u3_u0__abc_75526_new_n581_; 
wire u3_u0__abc_75526_new_n582_; 
wire u3_u0__abc_75526_new_n584_; 
wire u3_u0__abc_75526_new_n585_; 
wire u3_u0__abc_75526_new_n586_; 
wire u3_u0__abc_75526_new_n588_; 
wire u3_u0__abc_75526_new_n589_; 
wire u3_u0__abc_75526_new_n590_; 
wire u3_u0__abc_75526_new_n592_; 
wire u3_u0__abc_75526_new_n593_; 
wire u3_u0__abc_75526_new_n594_; 
wire u3_u0__abc_75526_new_n596_; 
wire u3_u0__abc_75526_new_n597_; 
wire u3_u0__abc_75526_new_n598_; 
wire u3_u0__abc_75526_new_n600_; 
wire u3_u0__abc_75526_new_n601_; 
wire u3_u0__abc_75526_new_n602_; 
wire u3_u0__abc_75526_new_n604_; 
wire u3_u0__abc_75526_new_n605_; 
wire u3_u0__abc_75526_new_n606_; 
wire u3_u0__abc_75526_new_n608_; 
wire u3_u0__abc_75526_new_n609_; 
wire u3_u0__abc_75526_new_n610_; 
wire u3_u0__abc_75526_new_n612_; 
wire u3_u0__abc_75526_new_n613_; 
wire u3_u0__abc_75526_new_n614_; 
wire u3_u0__abc_75526_new_n616_; 
wire u3_u0__abc_75526_new_n617_; 
wire u3_u0__abc_75526_new_n618_; 
wire u3_u0__abc_75526_new_n620_; 
wire u3_u0__abc_75526_new_n621_; 
wire u3_u0__abc_75526_new_n622_; 
wire u3_u0__abc_75526_new_n624_; 
wire u3_u0__abc_75526_new_n625_; 
wire u3_u0__abc_75526_new_n626_; 
wire u3_u0__abc_75526_new_n628_; 
wire u3_u0__abc_75526_new_n629_; 
wire u3_u0__abc_75526_new_n630_; 
wire u3_u0__abc_75526_new_n632_; 
wire u3_u0__abc_75526_new_n633_; 
wire u3_u0__abc_75526_new_n634_; 
wire u3_u0__abc_75526_new_n636_; 
wire u3_u0__abc_75526_new_n637_; 
wire u3_u0__abc_75526_new_n638_; 
wire u3_u0__abc_75526_new_n640_; 
wire u3_u0__abc_75526_new_n641_; 
wire u3_u0__abc_75526_new_n642_; 
wire u3_u0__abc_75526_new_n644_; 
wire u3_u0__abc_75526_new_n645_; 
wire u3_u0__abc_75526_new_n646_; 
wire u3_u0__abc_75526_new_n648_; 
wire u3_u0__abc_75526_new_n649_; 
wire u3_u0__abc_75526_new_n650_; 
wire u3_u0__abc_75526_new_n652_; 
wire u3_u0__abc_75526_new_n653_; 
wire u3_u0__abc_75526_new_n654_; 
wire u3_u0__abc_75526_new_n656_; 
wire u3_u0__abc_75526_new_n657_; 
wire u3_u0__abc_75526_new_n658_; 
wire u3_u0__abc_75526_new_n660_; 
wire u3_u0__abc_75526_new_n661_; 
wire u3_u0__abc_75526_new_n662_; 
wire u3_u0__abc_75526_new_n664_; 
wire u3_u0__abc_75526_new_n665_; 
wire u3_u0__abc_75526_new_n666_; 
wire u3_u0__abc_75526_new_n668_; 
wire u3_u0__abc_75526_new_n669_; 
wire u3_u0__abc_75526_new_n670_; 
wire u3_u0__abc_75526_new_n672_; 
wire u3_u0__abc_75526_new_n673_; 
wire u3_u0__abc_75526_new_n674_; 
wire u3_u0__abc_75526_new_n676_; 
wire u3_u0__abc_75526_new_n677_; 
wire u3_u0__abc_75526_new_n678_; 
wire u3_u0__abc_75526_new_n680_; 
wire u3_u0__abc_75526_new_n681_; 
wire u3_u0__abc_75526_new_n682_; 
wire u3_u0__abc_75526_new_n684_; 
wire u3_u0__abc_75526_new_n685_; 
wire u3_u0__abc_75526_new_n686_; 
wire u3_u0__abc_75526_new_n688_; 
wire u3_u0__abc_75526_new_n689_; 
wire u3_u0__abc_75526_new_n690_; 
wire u3_u0__abc_75526_new_n692_; 
wire u3_u0__abc_75526_new_n693_; 
wire u3_u0__abc_75526_new_n694_; 
wire u3_u0__abc_75526_new_n696_; 
wire u3_u0__abc_75526_new_n697_; 
wire u3_u0__abc_75526_new_n698_; 
wire u3_u0__abc_75526_new_n700_; 
wire u3_u0__abc_75526_new_n701_; 
wire u3_u0__abc_75526_new_n702_; 
wire u3_u0__abc_75526_new_n704_; 
wire u3_u0__abc_75526_new_n705_; 
wire u3_u0__abc_75526_new_n706_; 
wire u3_u0__abc_75526_new_n708_; 
wire u3_u0__abc_75526_new_n708__bF_buf0; 
wire u3_u0__abc_75526_new_n708__bF_buf1; 
wire u3_u0__abc_75526_new_n708__bF_buf2; 
wire u3_u0__abc_75526_new_n708__bF_buf3; 
wire u3_u0__abc_75526_new_n708__bF_buf4; 
wire u3_u0__abc_75526_new_n708__bF_buf5; 
wire u3_u0__abc_75526_new_n708__bF_buf6; 
wire u3_u0__abc_75526_new_n708__bF_buf7; 
wire u3_u0__abc_75526_new_n709_; 
wire u3_u0__abc_75526_new_n710_; 
wire u3_u0__abc_75526_new_n711_; 
wire u3_u0__abc_75526_new_n713_; 
wire u3_u0__abc_75526_new_n714_; 
wire u3_u0__abc_75526_new_n715_; 
wire u3_u0__abc_75526_new_n717_; 
wire u3_u0__abc_75526_new_n718_; 
wire u3_u0__abc_75526_new_n719_; 
wire u3_u0__abc_75526_new_n721_; 
wire u3_u0__abc_75526_new_n722_; 
wire u3_u0__abc_75526_new_n723_; 
wire u3_u0__abc_75526_new_n725_; 
wire u3_u0__abc_75526_new_n726_; 
wire u3_u0__abc_75526_new_n727_; 
wire u3_u0__abc_75526_new_n729_; 
wire u3_u0__abc_75526_new_n730_; 
wire u3_u0__abc_75526_new_n731_; 
wire u3_u0__abc_75526_new_n733_; 
wire u3_u0__abc_75526_new_n734_; 
wire u3_u0__abc_75526_new_n735_; 
wire u3_u0__abc_75526_new_n737_; 
wire u3_u0__abc_75526_new_n738_; 
wire u3_u0__abc_75526_new_n739_; 
wire u3_u0__abc_75526_new_n741_; 
wire u3_u0__abc_75526_new_n742_; 
wire u3_u0__abc_75526_new_n743_; 
wire u3_u0__abc_75526_new_n745_; 
wire u3_u0__abc_75526_new_n746_; 
wire u3_u0__abc_75526_new_n747_; 
wire u3_u0__abc_75526_new_n749_; 
wire u3_u0__abc_75526_new_n750_; 
wire u3_u0__abc_75526_new_n751_; 
wire u3_u0__abc_75526_new_n753_; 
wire u3_u0__abc_75526_new_n754_; 
wire u3_u0__abc_75526_new_n755_; 
wire u3_u0__abc_75526_new_n757_; 
wire u3_u0__abc_75526_new_n758_; 
wire u3_u0__abc_75526_new_n759_; 
wire u3_u0__abc_75526_new_n761_; 
wire u3_u0__abc_75526_new_n762_; 
wire u3_u0__abc_75526_new_n763_; 
wire u3_u0__abc_75526_new_n765_; 
wire u3_u0__abc_75526_new_n766_; 
wire u3_u0__abc_75526_new_n767_; 
wire u3_u0__abc_75526_new_n769_; 
wire u3_u0__abc_75526_new_n770_; 
wire u3_u0__abc_75526_new_n771_; 
wire u3_u0__abc_75526_new_n773_; 
wire u3_u0__abc_75526_new_n774_; 
wire u3_u0__abc_75526_new_n775_; 
wire u3_u0__abc_75526_new_n777_; 
wire u3_u0__abc_75526_new_n778_; 
wire u3_u0__abc_75526_new_n779_; 
wire u3_u0__abc_75526_new_n781_; 
wire u3_u0__abc_75526_new_n782_; 
wire u3_u0__abc_75526_new_n783_; 
wire u3_u0__abc_75526_new_n785_; 
wire u3_u0__abc_75526_new_n786_; 
wire u3_u0__abc_75526_new_n787_; 
wire u3_u0__abc_75526_new_n789_; 
wire u3_u0__abc_75526_new_n790_; 
wire u3_u0__abc_75526_new_n791_; 
wire u3_u0__abc_75526_new_n793_; 
wire u3_u0__abc_75526_new_n794_; 
wire u3_u0__abc_75526_new_n795_; 
wire u3_u0__abc_75526_new_n797_; 
wire u3_u0__abc_75526_new_n798_; 
wire u3_u0__abc_75526_new_n799_; 
wire u3_u0__abc_75526_new_n801_; 
wire u3_u0__abc_75526_new_n802_; 
wire u3_u0__abc_75526_new_n803_; 
wire u3_u0__abc_75526_new_n805_; 
wire u3_u0__abc_75526_new_n806_; 
wire u3_u0__abc_75526_new_n807_; 
wire u3_u0__abc_75526_new_n809_; 
wire u3_u0__abc_75526_new_n810_; 
wire u3_u0__abc_75526_new_n811_; 
wire u3_u0__abc_75526_new_n813_; 
wire u3_u0__abc_75526_new_n814_; 
wire u3_u0__abc_75526_new_n815_; 
wire u3_u0__abc_75526_new_n817_; 
wire u3_u0__abc_75526_new_n818_; 
wire u3_u0__abc_75526_new_n819_; 
wire u3_u0__abc_75526_new_n821_; 
wire u3_u0__abc_75526_new_n822_; 
wire u3_u0__abc_75526_new_n823_; 
wire u3_u0__abc_75526_new_n825_; 
wire u3_u0__abc_75526_new_n826_; 
wire u3_u0__abc_75526_new_n827_; 
wire u3_u0__abc_75526_new_n829_; 
wire u3_u0__abc_75526_new_n830_; 
wire u3_u0__abc_75526_new_n831_; 
wire u3_u0__abc_75526_new_n833_; 
wire u3_u0__abc_75526_new_n834_; 
wire u3_u0__abc_75526_new_n835_; 
wire u3_u0__abc_75526_new_n837_; 
wire u3_u0__abc_75526_new_n838_; 
wire u3_u0__abc_75526_new_n839_; 
wire u3_u0__abc_75526_new_n841_; 
wire u3_u0__abc_75526_new_n842_; 
wire u3_u0__abc_75526_new_n843_; 
wire u3_u0__abc_75526_new_n845_; 
wire u3_u0__abc_75526_new_n846_; 
wire u3_u0__abc_75526_new_n847_; 
wire u3_u0__abc_75526_new_n849_; 
wire u3_u0__abc_75526_new_n850_; 
wire u3_u0__abc_75526_new_n851_; 
wire u3_u0__abc_75526_new_n853_; 
wire u3_u0__abc_75526_new_n854_; 
wire u3_u0__abc_75526_new_n855_; 
wire u3_u0__abc_75526_new_n856_; 
wire u3_u0__abc_75526_new_n858_; 
wire u3_u0__abc_75526_new_n859_; 
wire u3_u0__abc_75526_new_n860_; 
wire u3_u0__abc_75526_new_n861_; 
wire u3_u0__abc_75526_new_n863_; 
wire u3_u0__abc_75526_new_n864_; 
wire u3_u0__abc_75526_new_n865_; 
wire u3_u0__abc_75526_new_n867_; 
wire u3_u0__abc_75526_new_n868_; 
wire u3_u0__abc_75526_new_n869_; 
wire u3_u0__abc_75526_new_n871_; 
wire u3_u0__abc_75526_new_n872_; 
wire u3_u0__abc_75526_new_n873_; 
wire u3_u0__abc_75526_new_n875_; 
wire u3_u0__abc_75526_new_n876_; 
wire u3_u0__abc_75526_new_n876__bF_buf0; 
wire u3_u0__abc_75526_new_n876__bF_buf1; 
wire u3_u0__abc_75526_new_n876__bF_buf2; 
wire u3_u0__abc_75526_new_n876__bF_buf3; 
wire u3_u0__abc_75526_new_n876__bF_buf4; 
wire u3_u0__abc_75526_new_n876__bF_buf5; 
wire u3_u0__abc_75526_new_n876__bF_buf6; 
wire u3_u0__abc_75526_new_n876__bF_buf7; 
wire u3_u0__abc_75526_new_n877_; 
wire u3_u0__abc_75526_new_n879_; 
wire u3_u0__abc_75526_new_n880_; 
wire u3_u0__abc_75526_new_n882_; 
wire u3_u0__abc_75526_new_n883_; 
wire u3_u0__abc_75526_new_n885_; 
wire u3_u0__abc_75526_new_n886_; 
wire u3_u0__abc_75526_new_n887_; 
wire u3_u0__abc_75526_new_n889_; 
wire u3_u0__abc_75526_new_n890_; 
wire u3_u0__abc_75526_new_n891_; 
wire u3_u0__abc_75526_new_n893_; 
wire u3_u0__abc_75526_new_n894_; 
wire u3_u0__abc_75526_new_n895_; 
wire u3_u0__abc_75526_new_n897_; 
wire u3_u0__abc_75526_new_n898_; 
wire u3_u0__abc_75526_new_n899_; 
wire u3_u0__abc_75526_new_n901_; 
wire u3_u0__abc_75526_new_n902_; 
wire u3_u0__abc_75526_new_n903_; 
wire u3_u0__abc_75526_new_n905_; 
wire u3_u0__abc_75526_new_n906_; 
wire u3_u0__abc_75526_new_n907_; 
wire u3_u0__abc_75526_new_n909_; 
wire u3_u0__abc_75526_new_n910_; 
wire u3_u0__abc_75526_new_n911_; 
wire u3_u0__abc_75526_new_n913_; 
wire u3_u0__abc_75526_new_n914_; 
wire u3_u0__abc_75526_new_n915_; 
wire u3_u0__abc_75526_new_n917_; 
wire u3_u0__abc_75526_new_n918_; 
wire u3_u0__abc_75526_new_n919_; 
wire u3_u0__abc_75526_new_n921_; 
wire u3_u0__abc_75526_new_n922_; 
wire u3_u0__abc_75526_new_n923_; 
wire u3_u0__abc_75526_new_n925_; 
wire u3_u0__abc_75526_new_n926_; 
wire u3_u0__abc_75526_new_n927_; 
wire u3_u0__abc_75526_new_n929_; 
wire u3_u0__abc_75526_new_n930_; 
wire u3_u0__abc_75526_new_n931_; 
wire u3_u0__abc_75526_new_n933_; 
wire u3_u0__abc_75526_new_n934_; 
wire u3_u0__abc_75526_new_n935_; 
wire u3_u0__abc_75526_new_n937_; 
wire u3_u0__abc_75526_new_n938_; 
wire u3_u0__abc_75526_new_n939_; 
wire u3_u0__abc_75526_new_n941_; 
wire u3_u0__abc_75526_new_n942_; 
wire u3_u0__abc_75526_new_n943_; 
wire u3_u0__abc_75526_new_n945_; 
wire u3_u0__abc_75526_new_n946_; 
wire u3_u0__abc_75526_new_n947_; 
wire u3_u0__abc_75526_new_n949_; 
wire u3_u0__abc_75526_new_n950_; 
wire u3_u0__abc_75526_new_n951_; 
wire u3_u0__abc_75526_new_n953_; 
wire u3_u0__abc_75526_new_n954_; 
wire u3_u0__abc_75526_new_n955_; 
wire u3_u0__abc_75526_new_n957_; 
wire u3_u0__abc_75526_new_n958_; 
wire u3_u0__abc_75526_new_n959_; 
wire u3_u0__abc_75526_new_n961_; 
wire u3_u0__abc_75526_new_n962_; 
wire u3_u0__abc_75526_new_n963_; 
wire u3_u0__abc_75526_new_n965_; 
wire u3_u0__abc_75526_new_n966_; 
wire u3_u0__abc_75526_new_n967_; 
wire u3_u0__abc_75526_new_n969_; 
wire u3_u0__abc_75526_new_n970_; 
wire u3_u0__abc_75526_new_n971_; 
wire u3_u0__abc_75526_new_n973_; 
wire u3_u0__abc_75526_new_n974_; 
wire u3_u0__abc_75526_new_n975_; 
wire u3_u0__abc_75526_new_n977_; 
wire u3_u0__abc_75526_new_n978_; 
wire u3_u0__abc_75526_new_n979_; 
wire u3_u0__abc_75526_new_n981_; 
wire u3_u0__abc_75526_new_n982_; 
wire u3_u0__abc_75526_new_n983_; 
wire u3_u0__abc_75526_new_n985_; 
wire u3_u0__abc_75526_new_n986_; 
wire u3_u0__abc_75526_new_n987_; 
wire u3_u0__abc_75526_new_n989_; 
wire u3_u0__abc_75526_new_n990_; 
wire u3_u0__abc_75526_new_n991_; 
wire u3_u0__abc_75526_new_n993_; 
wire u3_u0__abc_75526_new_n994_; 
wire u3_u0__abc_75526_new_n995_; 
wire u3_u0__abc_75526_new_n997_; 
wire u3_u0__abc_75526_new_n998_; 
wire u3_u0__abc_75526_new_n999_; 
wire u3_u0_r0_0_; 
wire u3_u0_r0_10_; 
wire u3_u0_r0_11_; 
wire u3_u0_r0_12_; 
wire u3_u0_r0_13_; 
wire u3_u0_r0_14_; 
wire u3_u0_r0_15_; 
wire u3_u0_r0_16_; 
wire u3_u0_r0_17_; 
wire u3_u0_r0_18_; 
wire u3_u0_r0_19_; 
wire u3_u0_r0_1_; 
wire u3_u0_r0_20_; 
wire u3_u0_r0_21_; 
wire u3_u0_r0_22_; 
wire u3_u0_r0_23_; 
wire u3_u0_r0_24_; 
wire u3_u0_r0_25_; 
wire u3_u0_r0_26_; 
wire u3_u0_r0_27_; 
wire u3_u0_r0_28_; 
wire u3_u0_r0_29_; 
wire u3_u0_r0_2_; 
wire u3_u0_r0_30_; 
wire u3_u0_r0_31_; 
wire u3_u0_r0_32_; 
wire u3_u0_r0_33_; 
wire u3_u0_r0_34_; 
wire u3_u0_r0_35_; 
wire u3_u0_r0_3_; 
wire u3_u0_r0_4_; 
wire u3_u0_r0_5_; 
wire u3_u0_r0_6_; 
wire u3_u0_r0_7_; 
wire u3_u0_r0_8_; 
wire u3_u0_r0_9_; 
wire u3_u0_r1_0_; 
wire u3_u0_r1_10_; 
wire u3_u0_r1_11_; 
wire u3_u0_r1_12_; 
wire u3_u0_r1_13_; 
wire u3_u0_r1_14_; 
wire u3_u0_r1_15_; 
wire u3_u0_r1_16_; 
wire u3_u0_r1_17_; 
wire u3_u0_r1_18_; 
wire u3_u0_r1_19_; 
wire u3_u0_r1_1_; 
wire u3_u0_r1_20_; 
wire u3_u0_r1_21_; 
wire u3_u0_r1_22_; 
wire u3_u0_r1_23_; 
wire u3_u0_r1_24_; 
wire u3_u0_r1_25_; 
wire u3_u0_r1_26_; 
wire u3_u0_r1_27_; 
wire u3_u0_r1_28_; 
wire u3_u0_r1_29_; 
wire u3_u0_r1_2_; 
wire u3_u0_r1_30_; 
wire u3_u0_r1_31_; 
wire u3_u0_r1_32_; 
wire u3_u0_r1_33_; 
wire u3_u0_r1_34_; 
wire u3_u0_r1_35_; 
wire u3_u0_r1_3_; 
wire u3_u0_r1_4_; 
wire u3_u0_r1_5_; 
wire u3_u0_r1_6_; 
wire u3_u0_r1_7_; 
wire u3_u0_r1_8_; 
wire u3_u0_r1_9_; 
wire u3_u0_r2_0_; 
wire u3_u0_r2_10_; 
wire u3_u0_r2_11_; 
wire u3_u0_r2_12_; 
wire u3_u0_r2_13_; 
wire u3_u0_r2_14_; 
wire u3_u0_r2_15_; 
wire u3_u0_r2_16_; 
wire u3_u0_r2_17_; 
wire u3_u0_r2_18_; 
wire u3_u0_r2_19_; 
wire u3_u0_r2_1_; 
wire u3_u0_r2_20_; 
wire u3_u0_r2_21_; 
wire u3_u0_r2_22_; 
wire u3_u0_r2_23_; 
wire u3_u0_r2_24_; 
wire u3_u0_r2_25_; 
wire u3_u0_r2_26_; 
wire u3_u0_r2_27_; 
wire u3_u0_r2_28_; 
wire u3_u0_r2_29_; 
wire u3_u0_r2_2_; 
wire u3_u0_r2_30_; 
wire u3_u0_r2_31_; 
wire u3_u0_r2_32_; 
wire u3_u0_r2_33_; 
wire u3_u0_r2_34_; 
wire u3_u0_r2_35_; 
wire u3_u0_r2_3_; 
wire u3_u0_r2_4_; 
wire u3_u0_r2_5_; 
wire u3_u0_r2_6_; 
wire u3_u0_r2_7_; 
wire u3_u0_r2_8_; 
wire u3_u0_r2_9_; 
wire u3_u0_r3_0_; 
wire u3_u0_r3_10_; 
wire u3_u0_r3_11_; 
wire u3_u0_r3_12_; 
wire u3_u0_r3_13_; 
wire u3_u0_r3_14_; 
wire u3_u0_r3_15_; 
wire u3_u0_r3_16_; 
wire u3_u0_r3_17_; 
wire u3_u0_r3_18_; 
wire u3_u0_r3_19_; 
wire u3_u0_r3_1_; 
wire u3_u0_r3_20_; 
wire u3_u0_r3_21_; 
wire u3_u0_r3_22_; 
wire u3_u0_r3_23_; 
wire u3_u0_r3_24_; 
wire u3_u0_r3_25_; 
wire u3_u0_r3_26_; 
wire u3_u0_r3_27_; 
wire u3_u0_r3_28_; 
wire u3_u0_r3_29_; 
wire u3_u0_r3_2_; 
wire u3_u0_r3_30_; 
wire u3_u0_r3_31_; 
wire u3_u0_r3_32_; 
wire u3_u0_r3_33_; 
wire u3_u0_r3_34_; 
wire u3_u0_r3_35_; 
wire u3_u0_r3_3_; 
wire u3_u0_r3_4_; 
wire u3_u0_r3_5_; 
wire u3_u0_r3_6_; 
wire u3_u0_r3_7_; 
wire u3_u0_r3_8_; 
wire u3_u0_r3_9_; 
wire u3_u0_rd_adr_0_; 
wire u3_u0_rd_adr_1_; 
wire u3_u0_rd_adr_2_; 
wire u3_u0_rd_adr_3_; 
wire u3_u0_wr_adr_0_; 
wire u3_u0_wr_adr_1_; 
wire u3_u0_wr_adr_2_; 
wire u3_u0_wr_adr_3_; 
wire u3_wb_read_go; 
wire u4__0ps_cnt_7_0__0_; 
wire u4__0ps_cnt_7_0__1_; 
wire u4__0ps_cnt_7_0__2_; 
wire u4__0ps_cnt_7_0__3_; 
wire u4__0ps_cnt_7_0__4_; 
wire u4__0ps_cnt_7_0__5_; 
wire u4__0ps_cnt_7_0__6_; 
wire u4__0ps_cnt_7_0__7_; 
wire u4__0rfr_clr_0_0_; 
wire u4__0rfr_cnt_7_0__0_; 
wire u4__0rfr_cnt_7_0__1_; 
wire u4__0rfr_cnt_7_0__2_; 
wire u4__0rfr_cnt_7_0__3_; 
wire u4__0rfr_cnt_7_0__4_; 
wire u4__0rfr_cnt_7_0__5_; 
wire u4__0rfr_cnt_7_0__6_; 
wire u4__0rfr_cnt_7_0__7_; 
wire u4__0rfr_early_0_0_; 
wire u4__0rfr_en_0_0_; 
wire u4__0rfr_req_0_0_; 
wire u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562; 
wire u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf0; 
wire u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf1; 
wire u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf2; 
wire u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf3; 
wire u4__abc_76448_new_n100_; 
wire u4__abc_76448_new_n101_; 
wire u4__abc_76448_new_n102_; 
wire u4__abc_76448_new_n103_; 
wire u4__abc_76448_new_n104_; 
wire u4__abc_76448_new_n105_; 
wire u4__abc_76448_new_n106_; 
wire u4__abc_76448_new_n107_; 
wire u4__abc_76448_new_n108_; 
wire u4__abc_76448_new_n109_; 
wire u4__abc_76448_new_n110_; 
wire u4__abc_76448_new_n111_; 
wire u4__abc_76448_new_n112_; 
wire u4__abc_76448_new_n113_; 
wire u4__abc_76448_new_n114_; 
wire u4__abc_76448_new_n116_; 
wire u4__abc_76448_new_n117_; 
wire u4__abc_76448_new_n119_; 
wire u4__abc_76448_new_n120_; 
wire u4__abc_76448_new_n121_; 
wire u4__abc_76448_new_n122_; 
wire u4__abc_76448_new_n124_; 
wire u4__abc_76448_new_n125_; 
wire u4__abc_76448_new_n126_; 
wire u4__abc_76448_new_n127_; 
wire u4__abc_76448_new_n129_; 
wire u4__abc_76448_new_n130_; 
wire u4__abc_76448_new_n131_; 
wire u4__abc_76448_new_n132_; 
wire u4__abc_76448_new_n133_; 
wire u4__abc_76448_new_n134_; 
wire u4__abc_76448_new_n136_; 
wire u4__abc_76448_new_n137_; 
wire u4__abc_76448_new_n138_; 
wire u4__abc_76448_new_n139_; 
wire u4__abc_76448_new_n140_; 
wire u4__abc_76448_new_n142_; 
wire u4__abc_76448_new_n143_; 
wire u4__abc_76448_new_n144_; 
wire u4__abc_76448_new_n145_; 
wire u4__abc_76448_new_n146_; 
wire u4__abc_76448_new_n147_; 
wire u4__abc_76448_new_n149_; 
wire u4__abc_76448_new_n150_; 
wire u4__abc_76448_new_n151_; 
wire u4__abc_76448_new_n152_; 
wire u4__abc_76448_new_n153_; 
wire u4__abc_76448_new_n155_; 
wire u4__abc_76448_new_n156_; 
wire u4__abc_76448_new_n157_; 
wire u4__abc_76448_new_n158_; 
wire u4__abc_76448_new_n159_; 
wire u4__abc_76448_new_n161_; 
wire u4__abc_76448_new_n162_; 
wire u4__abc_76448_new_n163_; 
wire u4__abc_76448_new_n164_; 
wire u4__abc_76448_new_n166_; 
wire u4__abc_76448_new_n167_; 
wire u4__abc_76448_new_n168_; 
wire u4__abc_76448_new_n169_; 
wire u4__abc_76448_new_n170_; 
wire u4__abc_76448_new_n171_; 
wire u4__abc_76448_new_n172_; 
wire u4__abc_76448_new_n173_; 
wire u4__abc_76448_new_n174_; 
wire u4__abc_76448_new_n175_; 
wire u4__abc_76448_new_n176_; 
wire u4__abc_76448_new_n177_; 
wire u4__abc_76448_new_n179_; 
wire u4__abc_76448_new_n180_; 
wire u4__abc_76448_new_n181_; 
wire u4__abc_76448_new_n182_; 
wire u4__abc_76448_new_n184_; 
wire u4__abc_76448_new_n185_; 
wire u4__abc_76448_new_n186_; 
wire u4__abc_76448_new_n187_; 
wire u4__abc_76448_new_n189_; 
wire u4__abc_76448_new_n190_; 
wire u4__abc_76448_new_n191_; 
wire u4__abc_76448_new_n192_; 
wire u4__abc_76448_new_n194_; 
wire u4__abc_76448_new_n195_; 
wire u4__abc_76448_new_n196_; 
wire u4__abc_76448_new_n197_; 
wire u4__abc_76448_new_n199_; 
wire u4__abc_76448_new_n200_; 
wire u4__abc_76448_new_n201_; 
wire u4__abc_76448_new_n202_; 
wire u4__abc_76448_new_n204_; 
wire u4__abc_76448_new_n205_; 
wire u4__abc_76448_new_n206_; 
wire u4__abc_76448_new_n207_; 
wire u4__abc_76448_new_n208_; 
wire u4__abc_76448_new_n209_; 
wire u4__abc_76448_new_n211_; 
wire u4__abc_76448_new_n212_; 
wire u4__abc_76448_new_n213_; 
wire u4__abc_76448_new_n214_; 
wire u4__abc_76448_new_n216_; 
wire u4__abc_76448_new_n217_; 
wire u4__abc_76448_new_n218_; 
wire u4__abc_76448_new_n219_; 
wire u4__abc_76448_new_n220_; 
wire u4__abc_76448_new_n222_; 
wire u4__abc_76448_new_n223_; 
wire u4__abc_76448_new_n224_; 
wire u4__abc_76448_new_n225_; 
wire u4__abc_76448_new_n226_; 
wire u4__abc_76448_new_n227_; 
wire u4__abc_76448_new_n228_; 
wire u4__abc_76448_new_n229_; 
wire u4__abc_76448_new_n230_; 
wire u4__abc_76448_new_n231_; 
wire u4__abc_76448_new_n232_; 
wire u4__abc_76448_new_n233_; 
wire u4__abc_76448_new_n234_; 
wire u4__abc_76448_new_n235_; 
wire u4__abc_76448_new_n236_; 
wire u4__abc_76448_new_n237_; 
wire u4__abc_76448_new_n238_; 
wire u4__abc_76448_new_n239_; 
wire u4__abc_76448_new_n240_; 
wire u4__abc_76448_new_n241_; 
wire u4__abc_76448_new_n65_; 
wire u4__abc_76448_new_n66_; 
wire u4__abc_76448_new_n67_; 
wire u4__abc_76448_new_n68_; 
wire u4__abc_76448_new_n69_; 
wire u4__abc_76448_new_n70_; 
wire u4__abc_76448_new_n72_; 
wire u4__abc_76448_new_n73_; 
wire u4__abc_76448_new_n74_; 
wire u4__abc_76448_new_n75_; 
wire u4__abc_76448_new_n76_; 
wire u4__abc_76448_new_n77_; 
wire u4__abc_76448_new_n78_; 
wire u4__abc_76448_new_n79_; 
wire u4__abc_76448_new_n80_; 
wire u4__abc_76448_new_n81_; 
wire u4__abc_76448_new_n82_; 
wire u4__abc_76448_new_n83_; 
wire u4__abc_76448_new_n84_; 
wire u4__abc_76448_new_n85_; 
wire u4__abc_76448_new_n86_; 
wire u4__abc_76448_new_n87_; 
wire u4__abc_76448_new_n88_; 
wire u4__abc_76448_new_n89_; 
wire u4__abc_76448_new_n90_; 
wire u4__abc_76448_new_n91_; 
wire u4__abc_76448_new_n92_; 
wire u4__abc_76448_new_n93_; 
wire u4__abc_76448_new_n94_; 
wire u4__abc_76448_new_n95_; 
wire u4__abc_76448_new_n96_; 
wire u4__abc_76448_new_n97_; 
wire u4__abc_76448_new_n98_; 
wire u4__abc_76448_new_n99_; 
wire u4_ps_cnt_0_; 
wire u4_ps_cnt_1_; 
wire u4_ps_cnt_2_; 
wire u4_ps_cnt_3_; 
wire u4_ps_cnt_4_; 
wire u4_ps_cnt_5_; 
wire u4_ps_cnt_6_; 
wire u4_ps_cnt_7_; 
wire u4_ps_cnt_clr; 
wire u4_rfr_ce; 
wire u4_rfr_clr; 
wire u4_rfr_cnt_0_; 
wire u4_rfr_cnt_1_; 
wire u4_rfr_cnt_2_; 
wire u4_rfr_cnt_3_; 
wire u4_rfr_cnt_4_; 
wire u4_rfr_cnt_5_; 
wire u4_rfr_cnt_6_; 
wire u4_rfr_cnt_7_; 
wire u4_rfr_early; 
wire u4_rfr_en; 
wire u5__0ack_cnt_3_0__0_; 
wire u5__0ack_cnt_3_0__1_; 
wire u5__0ack_cnt_3_0__2_; 
wire u5__0ack_cnt_3_0__3_; 
wire u5__0ap_en_0_0_; 
wire u5__0burst_act_rd_0_0_; 
wire u5__0burst_cnt_10_0__0_; 
wire u5__0burst_cnt_10_0__10_; 
wire u5__0burst_cnt_10_0__1_; 
wire u5__0burst_cnt_10_0__2_; 
wire u5__0burst_cnt_10_0__3_; 
wire u5__0burst_cnt_10_0__4_; 
wire u5__0burst_cnt_10_0__5_; 
wire u5__0burst_cnt_10_0__6_; 
wire u5__0burst_cnt_10_0__7_; 
wire u5__0burst_cnt_10_0__8_; 
wire u5__0burst_cnt_10_0__9_; 
wire u5__0cke__0_0_; 
wire u5__0cmd_asserted2_0_0_; 
wire u5__0cmd_asserted_0_0_; 
wire u5__0data_oe_0_0_; 
wire u5__0ir_cnt_3_0__0_; 
wire u5__0ir_cnt_3_0__1_; 
wire u5__0ir_cnt_3_0__2_; 
wire u5__0ir_cnt_3_0__3_; 
wire u5__0ir_cnt_done_0_0_; 
wire u5__0lookup_ready1_0_0_; 
wire u5__0lookup_ready2_0_0_; 
wire u5__0mc_adv_r1_0_0_; 
wire u5__0mc_adv_r_0_0_; 
wire u5__0mc_le_0_0_; 
wire u5__0no_wb_cycle_0_0_; 
wire u5__0oe__0_0_; 
wire u5__0susp_sel_r_0_0_; 
wire u5__0timer2_8_0__0_; 
wire u5__0timer2_8_0__1_; 
wire u5__0timer2_8_0__2_; 
wire u5__0timer2_8_0__3_; 
wire u5__0timer2_8_0__4_; 
wire u5__0timer2_8_0__5_; 
wire u5__0timer2_8_0__6_; 
wire u5__0timer2_8_0__7_; 
wire u5__0timer2_8_0__8_; 
wire u5__0timer_7_0__0_; 
wire u5__0timer_7_0__1_; 
wire u5__0timer_7_0__2_; 
wire u5__0timer_7_0__3_; 
wire u5__0timer_7_0__4_; 
wire u5__0timer_7_0__5_; 
wire u5__0timer_7_0__6_; 
wire u5__0timer_7_0__7_; 
wire u5__0tmr2_done_0_0_; 
wire u5__0wb_cycle_0_0_; 
wire u5__0wb_stb_first_0_0_; 
wire u5__0wr_cycle_0_0_; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9; 
wire u5__abc_81276_auto_rtlil_cc_1942_NotGate_72182; 
wire u5__abc_81276_new_n1000_; 
wire u5__abc_81276_new_n1001_; 
wire u5__abc_81276_new_n1002_; 
wire u5__abc_81276_new_n1003_; 
wire u5__abc_81276_new_n1004_; 
wire u5__abc_81276_new_n1005_; 
wire u5__abc_81276_new_n1006_; 
wire u5__abc_81276_new_n1007_; 
wire u5__abc_81276_new_n1008_; 
wire u5__abc_81276_new_n1009_; 
wire u5__abc_81276_new_n1010_; 
wire u5__abc_81276_new_n1011_; 
wire u5__abc_81276_new_n1012_; 
wire u5__abc_81276_new_n1013_; 
wire u5__abc_81276_new_n1014_; 
wire u5__abc_81276_new_n1015_; 
wire u5__abc_81276_new_n1016_; 
wire u5__abc_81276_new_n1017_; 
wire u5__abc_81276_new_n1018_; 
wire u5__abc_81276_new_n1019_; 
wire u5__abc_81276_new_n1020_; 
wire u5__abc_81276_new_n1021_; 
wire u5__abc_81276_new_n1022_; 
wire u5__abc_81276_new_n1023_; 
wire u5__abc_81276_new_n1024_; 
wire u5__abc_81276_new_n1025_; 
wire u5__abc_81276_new_n1026_; 
wire u5__abc_81276_new_n1027_; 
wire u5__abc_81276_new_n1028_; 
wire u5__abc_81276_new_n1029_; 
wire u5__abc_81276_new_n1030_; 
wire u5__abc_81276_new_n1031_; 
wire u5__abc_81276_new_n1032_; 
wire u5__abc_81276_new_n1033_; 
wire u5__abc_81276_new_n1034_; 
wire u5__abc_81276_new_n1035_; 
wire u5__abc_81276_new_n1036_; 
wire u5__abc_81276_new_n1037_; 
wire u5__abc_81276_new_n1038_; 
wire u5__abc_81276_new_n1039_; 
wire u5__abc_81276_new_n1040_; 
wire u5__abc_81276_new_n1041_; 
wire u5__abc_81276_new_n1042_; 
wire u5__abc_81276_new_n1043_; 
wire u5__abc_81276_new_n1044_; 
wire u5__abc_81276_new_n1045_; 
wire u5__abc_81276_new_n1046_; 
wire u5__abc_81276_new_n1047_; 
wire u5__abc_81276_new_n1048_; 
wire u5__abc_81276_new_n1049_; 
wire u5__abc_81276_new_n1050_; 
wire u5__abc_81276_new_n1051_; 
wire u5__abc_81276_new_n1052_; 
wire u5__abc_81276_new_n1053_; 
wire u5__abc_81276_new_n1054_; 
wire u5__abc_81276_new_n1055_; 
wire u5__abc_81276_new_n1056_; 
wire u5__abc_81276_new_n1057_; 
wire u5__abc_81276_new_n1058_; 
wire u5__abc_81276_new_n1059_; 
wire u5__abc_81276_new_n1060_; 
wire u5__abc_81276_new_n1061_; 
wire u5__abc_81276_new_n1062_; 
wire u5__abc_81276_new_n1063_; 
wire u5__abc_81276_new_n1064_; 
wire u5__abc_81276_new_n1065_; 
wire u5__abc_81276_new_n1066_; 
wire u5__abc_81276_new_n1067_; 
wire u5__abc_81276_new_n1068_; 
wire u5__abc_81276_new_n1069_; 
wire u5__abc_81276_new_n1070_; 
wire u5__abc_81276_new_n1071_; 
wire u5__abc_81276_new_n1072_; 
wire u5__abc_81276_new_n1073_; 
wire u5__abc_81276_new_n1074_; 
wire u5__abc_81276_new_n1075_; 
wire u5__abc_81276_new_n1076_; 
wire u5__abc_81276_new_n1077_; 
wire u5__abc_81276_new_n1078_; 
wire u5__abc_81276_new_n1079_; 
wire u5__abc_81276_new_n1080_; 
wire u5__abc_81276_new_n1081_; 
wire u5__abc_81276_new_n1082_; 
wire u5__abc_81276_new_n1083_; 
wire u5__abc_81276_new_n1084_; 
wire u5__abc_81276_new_n1085_; 
wire u5__abc_81276_new_n1086_; 
wire u5__abc_81276_new_n1087_; 
wire u5__abc_81276_new_n1088_; 
wire u5__abc_81276_new_n1089_; 
wire u5__abc_81276_new_n1090_; 
wire u5__abc_81276_new_n1091_; 
wire u5__abc_81276_new_n1092_; 
wire u5__abc_81276_new_n1093_; 
wire u5__abc_81276_new_n1094_; 
wire u5__abc_81276_new_n1095_; 
wire u5__abc_81276_new_n1096_; 
wire u5__abc_81276_new_n1097_; 
wire u5__abc_81276_new_n1098_; 
wire u5__abc_81276_new_n1101_; 
wire u5__abc_81276_new_n1102_; 
wire u5__abc_81276_new_n1103_; 
wire u5__abc_81276_new_n1104_; 
wire u5__abc_81276_new_n1105_; 
wire u5__abc_81276_new_n1106_; 
wire u5__abc_81276_new_n1107_; 
wire u5__abc_81276_new_n1108_; 
wire u5__abc_81276_new_n1109_; 
wire u5__abc_81276_new_n1110_; 
wire u5__abc_81276_new_n1111_; 
wire u5__abc_81276_new_n1112_; 
wire u5__abc_81276_new_n1113_; 
wire u5__abc_81276_new_n1114_; 
wire u5__abc_81276_new_n1116_; 
wire u5__abc_81276_new_n1117_; 
wire u5__abc_81276_new_n1118_; 
wire u5__abc_81276_new_n1119_; 
wire u5__abc_81276_new_n1120_; 
wire u5__abc_81276_new_n1121_; 
wire u5__abc_81276_new_n1123_; 
wire u5__abc_81276_new_n1124_; 
wire u5__abc_81276_new_n1126_; 
wire u5__abc_81276_new_n1126__bF_buf0; 
wire u5__abc_81276_new_n1126__bF_buf1; 
wire u5__abc_81276_new_n1126__bF_buf2; 
wire u5__abc_81276_new_n1126__bF_buf3; 
wire u5__abc_81276_new_n1127_; 
wire u5__abc_81276_new_n1128_; 
wire u5__abc_81276_new_n1129_; 
wire u5__abc_81276_new_n1130_; 
wire u5__abc_81276_new_n1131_; 
wire u5__abc_81276_new_n1132_; 
wire u5__abc_81276_new_n1133_; 
wire u5__abc_81276_new_n1134_; 
wire u5__abc_81276_new_n1135_; 
wire u5__abc_81276_new_n1136_; 
wire u5__abc_81276_new_n1137_; 
wire u5__abc_81276_new_n1138_; 
wire u5__abc_81276_new_n1139_; 
wire u5__abc_81276_new_n1140_; 
wire u5__abc_81276_new_n1141_; 
wire u5__abc_81276_new_n1142_; 
wire u5__abc_81276_new_n1143_; 
wire u5__abc_81276_new_n1144_; 
wire u5__abc_81276_new_n1145_; 
wire u5__abc_81276_new_n1146_; 
wire u5__abc_81276_new_n1147_; 
wire u5__abc_81276_new_n1148_; 
wire u5__abc_81276_new_n1149_; 
wire u5__abc_81276_new_n1150_; 
wire u5__abc_81276_new_n1151_; 
wire u5__abc_81276_new_n1152_; 
wire u5__abc_81276_new_n1153_; 
wire u5__abc_81276_new_n1154_; 
wire u5__abc_81276_new_n1155_; 
wire u5__abc_81276_new_n1156_; 
wire u5__abc_81276_new_n1157_; 
wire u5__abc_81276_new_n1158_; 
wire u5__abc_81276_new_n1159_; 
wire u5__abc_81276_new_n1160_; 
wire u5__abc_81276_new_n1161_; 
wire u5__abc_81276_new_n1162_; 
wire u5__abc_81276_new_n1163_; 
wire u5__abc_81276_new_n1164_; 
wire u5__abc_81276_new_n1165_; 
wire u5__abc_81276_new_n1166_; 
wire u5__abc_81276_new_n1167_; 
wire u5__abc_81276_new_n1168_; 
wire u5__abc_81276_new_n1169_; 
wire u5__abc_81276_new_n1170_; 
wire u5__abc_81276_new_n1171_; 
wire u5__abc_81276_new_n1172_; 
wire u5__abc_81276_new_n1173_; 
wire u5__abc_81276_new_n1174_; 
wire u5__abc_81276_new_n1175_; 
wire u5__abc_81276_new_n1176_; 
wire u5__abc_81276_new_n1177_; 
wire u5__abc_81276_new_n1178_; 
wire u5__abc_81276_new_n1179_; 
wire u5__abc_81276_new_n1180_; 
wire u5__abc_81276_new_n1181_; 
wire u5__abc_81276_new_n1182_; 
wire u5__abc_81276_new_n1183_; 
wire u5__abc_81276_new_n1184_; 
wire u5__abc_81276_new_n1185_; 
wire u5__abc_81276_new_n1186_; 
wire u5__abc_81276_new_n1187_; 
wire u5__abc_81276_new_n1188_; 
wire u5__abc_81276_new_n1189_; 
wire u5__abc_81276_new_n1190_; 
wire u5__abc_81276_new_n1191_; 
wire u5__abc_81276_new_n1192_; 
wire u5__abc_81276_new_n1193_; 
wire u5__abc_81276_new_n1194_; 
wire u5__abc_81276_new_n1195_; 
wire u5__abc_81276_new_n1196_; 
wire u5__abc_81276_new_n1197_; 
wire u5__abc_81276_new_n1198_; 
wire u5__abc_81276_new_n1199_; 
wire u5__abc_81276_new_n1200_; 
wire u5__abc_81276_new_n1201_; 
wire u5__abc_81276_new_n1202_; 
wire u5__abc_81276_new_n1203_; 
wire u5__abc_81276_new_n1204_; 
wire u5__abc_81276_new_n1205_; 
wire u5__abc_81276_new_n1206_; 
wire u5__abc_81276_new_n1207_; 
wire u5__abc_81276_new_n1208_; 
wire u5__abc_81276_new_n1209_; 
wire u5__abc_81276_new_n1210_; 
wire u5__abc_81276_new_n1211_; 
wire u5__abc_81276_new_n1212_; 
wire u5__abc_81276_new_n1213_; 
wire u5__abc_81276_new_n1214_; 
wire u5__abc_81276_new_n1215_; 
wire u5__abc_81276_new_n1216_; 
wire u5__abc_81276_new_n1217_; 
wire u5__abc_81276_new_n1218_; 
wire u5__abc_81276_new_n1219_; 
wire u5__abc_81276_new_n1220_; 
wire u5__abc_81276_new_n1221_; 
wire u5__abc_81276_new_n1222_; 
wire u5__abc_81276_new_n1223_; 
wire u5__abc_81276_new_n1224_; 
wire u5__abc_81276_new_n1225_; 
wire u5__abc_81276_new_n1226_; 
wire u5__abc_81276_new_n1227_; 
wire u5__abc_81276_new_n1228_; 
wire u5__abc_81276_new_n1229_; 
wire u5__abc_81276_new_n1230_; 
wire u5__abc_81276_new_n1231_; 
wire u5__abc_81276_new_n1232_; 
wire u5__abc_81276_new_n1233_; 
wire u5__abc_81276_new_n1234_; 
wire u5__abc_81276_new_n1235_; 
wire u5__abc_81276_new_n1236_; 
wire u5__abc_81276_new_n1237_; 
wire u5__abc_81276_new_n1238_; 
wire u5__abc_81276_new_n1239_; 
wire u5__abc_81276_new_n1240_; 
wire u5__abc_81276_new_n1241_; 
wire u5__abc_81276_new_n1242_; 
wire u5__abc_81276_new_n1243_; 
wire u5__abc_81276_new_n1244_; 
wire u5__abc_81276_new_n1245_; 
wire u5__abc_81276_new_n1246_; 
wire u5__abc_81276_new_n1247_; 
wire u5__abc_81276_new_n1248_; 
wire u5__abc_81276_new_n1249_; 
wire u5__abc_81276_new_n1250_; 
wire u5__abc_81276_new_n1251_; 
wire u5__abc_81276_new_n1252_; 
wire u5__abc_81276_new_n1253_; 
wire u5__abc_81276_new_n1254_; 
wire u5__abc_81276_new_n1255_; 
wire u5__abc_81276_new_n1256_; 
wire u5__abc_81276_new_n1257_; 
wire u5__abc_81276_new_n1258_; 
wire u5__abc_81276_new_n1259_; 
wire u5__abc_81276_new_n1260_; 
wire u5__abc_81276_new_n1261_; 
wire u5__abc_81276_new_n1262_; 
wire u5__abc_81276_new_n1263_; 
wire u5__abc_81276_new_n1264_; 
wire u5__abc_81276_new_n1265_; 
wire u5__abc_81276_new_n1266_; 
wire u5__abc_81276_new_n1267_; 
wire u5__abc_81276_new_n1268_; 
wire u5__abc_81276_new_n1269_; 
wire u5__abc_81276_new_n1270_; 
wire u5__abc_81276_new_n1271_; 
wire u5__abc_81276_new_n1272_; 
wire u5__abc_81276_new_n1273_; 
wire u5__abc_81276_new_n1274_; 
wire u5__abc_81276_new_n1275_; 
wire u5__abc_81276_new_n1276_; 
wire u5__abc_81276_new_n1277_; 
wire u5__abc_81276_new_n1278_; 
wire u5__abc_81276_new_n1279_; 
wire u5__abc_81276_new_n1280_; 
wire u5__abc_81276_new_n1281_; 
wire u5__abc_81276_new_n1282_; 
wire u5__abc_81276_new_n1283_; 
wire u5__abc_81276_new_n1284_; 
wire u5__abc_81276_new_n1285_; 
wire u5__abc_81276_new_n1286_; 
wire u5__abc_81276_new_n1287_; 
wire u5__abc_81276_new_n1288_; 
wire u5__abc_81276_new_n1289_; 
wire u5__abc_81276_new_n1290_; 
wire u5__abc_81276_new_n1291_; 
wire u5__abc_81276_new_n1292_; 
wire u5__abc_81276_new_n1293_; 
wire u5__abc_81276_new_n1294_; 
wire u5__abc_81276_new_n1295_; 
wire u5__abc_81276_new_n1296_; 
wire u5__abc_81276_new_n1297_; 
wire u5__abc_81276_new_n1298_; 
wire u5__abc_81276_new_n1299_; 
wire u5__abc_81276_new_n1300_; 
wire u5__abc_81276_new_n1301_; 
wire u5__abc_81276_new_n1302_; 
wire u5__abc_81276_new_n1303_; 
wire u5__abc_81276_new_n1304_; 
wire u5__abc_81276_new_n1305_; 
wire u5__abc_81276_new_n1306_; 
wire u5__abc_81276_new_n1307_; 
wire u5__abc_81276_new_n1308_; 
wire u5__abc_81276_new_n1309_; 
wire u5__abc_81276_new_n1310_; 
wire u5__abc_81276_new_n1311_; 
wire u5__abc_81276_new_n1312_; 
wire u5__abc_81276_new_n1313_; 
wire u5__abc_81276_new_n1314_; 
wire u5__abc_81276_new_n1315_; 
wire u5__abc_81276_new_n1316_; 
wire u5__abc_81276_new_n1317_; 
wire u5__abc_81276_new_n1318_; 
wire u5__abc_81276_new_n1319_; 
wire u5__abc_81276_new_n1320_; 
wire u5__abc_81276_new_n1321_; 
wire u5__abc_81276_new_n1322_; 
wire u5__abc_81276_new_n1323_; 
wire u5__abc_81276_new_n1324_; 
wire u5__abc_81276_new_n1325_; 
wire u5__abc_81276_new_n1326_; 
wire u5__abc_81276_new_n1327_; 
wire u5__abc_81276_new_n1328_; 
wire u5__abc_81276_new_n1329_; 
wire u5__abc_81276_new_n1330_; 
wire u5__abc_81276_new_n1331_; 
wire u5__abc_81276_new_n1332_; 
wire u5__abc_81276_new_n1333_; 
wire u5__abc_81276_new_n1334_; 
wire u5__abc_81276_new_n1335_; 
wire u5__abc_81276_new_n1336_; 
wire u5__abc_81276_new_n1337_; 
wire u5__abc_81276_new_n1338_; 
wire u5__abc_81276_new_n1339_; 
wire u5__abc_81276_new_n1340_; 
wire u5__abc_81276_new_n1341_; 
wire u5__abc_81276_new_n1342_; 
wire u5__abc_81276_new_n1343_; 
wire u5__abc_81276_new_n1344_; 
wire u5__abc_81276_new_n1345_; 
wire u5__abc_81276_new_n1346_; 
wire u5__abc_81276_new_n1347_; 
wire u5__abc_81276_new_n1348_; 
wire u5__abc_81276_new_n1349_; 
wire u5__abc_81276_new_n1350_; 
wire u5__abc_81276_new_n1351_; 
wire u5__abc_81276_new_n1352_; 
wire u5__abc_81276_new_n1353_; 
wire u5__abc_81276_new_n1354_; 
wire u5__abc_81276_new_n1355_; 
wire u5__abc_81276_new_n1356_; 
wire u5__abc_81276_new_n1357_; 
wire u5__abc_81276_new_n1358_; 
wire u5__abc_81276_new_n1359_; 
wire u5__abc_81276_new_n1360_; 
wire u5__abc_81276_new_n1361_; 
wire u5__abc_81276_new_n1362_; 
wire u5__abc_81276_new_n1363_; 
wire u5__abc_81276_new_n1364_; 
wire u5__abc_81276_new_n1365_; 
wire u5__abc_81276_new_n1366_; 
wire u5__abc_81276_new_n1367_; 
wire u5__abc_81276_new_n1368_; 
wire u5__abc_81276_new_n1369_; 
wire u5__abc_81276_new_n1370_; 
wire u5__abc_81276_new_n1371_; 
wire u5__abc_81276_new_n1372_; 
wire u5__abc_81276_new_n1373_; 
wire u5__abc_81276_new_n1374_; 
wire u5__abc_81276_new_n1375_; 
wire u5__abc_81276_new_n1376_; 
wire u5__abc_81276_new_n1377_; 
wire u5__abc_81276_new_n1378_; 
wire u5__abc_81276_new_n1379_; 
wire u5__abc_81276_new_n1380_; 
wire u5__abc_81276_new_n1381_; 
wire u5__abc_81276_new_n1382_; 
wire u5__abc_81276_new_n1383_; 
wire u5__abc_81276_new_n1384_; 
wire u5__abc_81276_new_n1385_; 
wire u5__abc_81276_new_n1386_; 
wire u5__abc_81276_new_n1387_; 
wire u5__abc_81276_new_n1388_; 
wire u5__abc_81276_new_n1389_; 
wire u5__abc_81276_new_n1390_; 
wire u5__abc_81276_new_n1391_; 
wire u5__abc_81276_new_n1392_; 
wire u5__abc_81276_new_n1393_; 
wire u5__abc_81276_new_n1394_; 
wire u5__abc_81276_new_n1395_; 
wire u5__abc_81276_new_n1396_; 
wire u5__abc_81276_new_n1397_; 
wire u5__abc_81276_new_n1398_; 
wire u5__abc_81276_new_n1399_; 
wire u5__abc_81276_new_n1400_; 
wire u5__abc_81276_new_n1401_; 
wire u5__abc_81276_new_n1402_; 
wire u5__abc_81276_new_n1403_; 
wire u5__abc_81276_new_n1404_; 
wire u5__abc_81276_new_n1405_; 
wire u5__abc_81276_new_n1406_; 
wire u5__abc_81276_new_n1407_; 
wire u5__abc_81276_new_n1408_; 
wire u5__abc_81276_new_n1409_; 
wire u5__abc_81276_new_n1410_; 
wire u5__abc_81276_new_n1411_; 
wire u5__abc_81276_new_n1412_; 
wire u5__abc_81276_new_n1413_; 
wire u5__abc_81276_new_n1414_; 
wire u5__abc_81276_new_n1415_; 
wire u5__abc_81276_new_n1416_; 
wire u5__abc_81276_new_n1417_; 
wire u5__abc_81276_new_n1418_; 
wire u5__abc_81276_new_n1419_; 
wire u5__abc_81276_new_n1420_; 
wire u5__abc_81276_new_n1421_; 
wire u5__abc_81276_new_n1422_; 
wire u5__abc_81276_new_n1423_; 
wire u5__abc_81276_new_n1424_; 
wire u5__abc_81276_new_n1425_; 
wire u5__abc_81276_new_n1426_; 
wire u5__abc_81276_new_n1427_; 
wire u5__abc_81276_new_n1428_; 
wire u5__abc_81276_new_n1429_; 
wire u5__abc_81276_new_n1430_; 
wire u5__abc_81276_new_n1431_; 
wire u5__abc_81276_new_n1432_; 
wire u5__abc_81276_new_n1433_; 
wire u5__abc_81276_new_n1434_; 
wire u5__abc_81276_new_n1435_; 
wire u5__abc_81276_new_n1436_; 
wire u5__abc_81276_new_n1437_; 
wire u5__abc_81276_new_n1438_; 
wire u5__abc_81276_new_n1439_; 
wire u5__abc_81276_new_n1440_; 
wire u5__abc_81276_new_n1441_; 
wire u5__abc_81276_new_n1442_; 
wire u5__abc_81276_new_n1443_; 
wire u5__abc_81276_new_n1444_; 
wire u5__abc_81276_new_n1445_; 
wire u5__abc_81276_new_n1446_; 
wire u5__abc_81276_new_n1447_; 
wire u5__abc_81276_new_n1448_; 
wire u5__abc_81276_new_n1449_; 
wire u5__abc_81276_new_n1450_; 
wire u5__abc_81276_new_n1451_; 
wire u5__abc_81276_new_n1452_; 
wire u5__abc_81276_new_n1453_; 
wire u5__abc_81276_new_n1454_; 
wire u5__abc_81276_new_n1455_; 
wire u5__abc_81276_new_n1456_; 
wire u5__abc_81276_new_n1457_; 
wire u5__abc_81276_new_n1458_; 
wire u5__abc_81276_new_n1459_; 
wire u5__abc_81276_new_n1460_; 
wire u5__abc_81276_new_n1461_; 
wire u5__abc_81276_new_n1462_; 
wire u5__abc_81276_new_n1463_; 
wire u5__abc_81276_new_n1464_; 
wire u5__abc_81276_new_n1465_; 
wire u5__abc_81276_new_n1466_; 
wire u5__abc_81276_new_n1467_; 
wire u5__abc_81276_new_n1468_; 
wire u5__abc_81276_new_n1469_; 
wire u5__abc_81276_new_n1470_; 
wire u5__abc_81276_new_n1471_; 
wire u5__abc_81276_new_n1472_; 
wire u5__abc_81276_new_n1473_; 
wire u5__abc_81276_new_n1474_; 
wire u5__abc_81276_new_n1475_; 
wire u5__abc_81276_new_n1476_; 
wire u5__abc_81276_new_n1477_; 
wire u5__abc_81276_new_n1478_; 
wire u5__abc_81276_new_n1479_; 
wire u5__abc_81276_new_n1480_; 
wire u5__abc_81276_new_n1481_; 
wire u5__abc_81276_new_n1482_; 
wire u5__abc_81276_new_n1483_; 
wire u5__abc_81276_new_n1484_; 
wire u5__abc_81276_new_n1485_; 
wire u5__abc_81276_new_n1486_; 
wire u5__abc_81276_new_n1487_; 
wire u5__abc_81276_new_n1488_; 
wire u5__abc_81276_new_n1489_; 
wire u5__abc_81276_new_n1490_; 
wire u5__abc_81276_new_n1491_; 
wire u5__abc_81276_new_n1492_; 
wire u5__abc_81276_new_n1493_; 
wire u5__abc_81276_new_n1494_; 
wire u5__abc_81276_new_n1495_; 
wire u5__abc_81276_new_n1496_; 
wire u5__abc_81276_new_n1497_; 
wire u5__abc_81276_new_n1498_; 
wire u5__abc_81276_new_n1499_; 
wire u5__abc_81276_new_n1500_; 
wire u5__abc_81276_new_n1501_; 
wire u5__abc_81276_new_n1502_; 
wire u5__abc_81276_new_n1503_; 
wire u5__abc_81276_new_n1504_; 
wire u5__abc_81276_new_n1505_; 
wire u5__abc_81276_new_n1506_; 
wire u5__abc_81276_new_n1507_; 
wire u5__abc_81276_new_n1508_; 
wire u5__abc_81276_new_n1509_; 
wire u5__abc_81276_new_n1510_; 
wire u5__abc_81276_new_n1511_; 
wire u5__abc_81276_new_n1512_; 
wire u5__abc_81276_new_n1513_; 
wire u5__abc_81276_new_n1514_; 
wire u5__abc_81276_new_n1515_; 
wire u5__abc_81276_new_n1516_; 
wire u5__abc_81276_new_n1517_; 
wire u5__abc_81276_new_n1518_; 
wire u5__abc_81276_new_n1519_; 
wire u5__abc_81276_new_n1520_; 
wire u5__abc_81276_new_n1521_; 
wire u5__abc_81276_new_n1522_; 
wire u5__abc_81276_new_n1523_; 
wire u5__abc_81276_new_n1524_; 
wire u5__abc_81276_new_n1525_; 
wire u5__abc_81276_new_n1526_; 
wire u5__abc_81276_new_n1526__bF_buf0; 
wire u5__abc_81276_new_n1526__bF_buf1; 
wire u5__abc_81276_new_n1526__bF_buf2; 
wire u5__abc_81276_new_n1526__bF_buf3; 
wire u5__abc_81276_new_n1527_; 
wire u5__abc_81276_new_n1528_; 
wire u5__abc_81276_new_n1529_; 
wire u5__abc_81276_new_n1530_; 
wire u5__abc_81276_new_n1531_; 
wire u5__abc_81276_new_n1533_; 
wire u5__abc_81276_new_n1534_; 
wire u5__abc_81276_new_n1535_; 
wire u5__abc_81276_new_n1536_; 
wire u5__abc_81276_new_n1537_; 
wire u5__abc_81276_new_n1538_; 
wire u5__abc_81276_new_n1539_; 
wire u5__abc_81276_new_n1540_; 
wire u5__abc_81276_new_n1541_; 
wire u5__abc_81276_new_n1542_; 
wire u5__abc_81276_new_n1543_; 
wire u5__abc_81276_new_n1544_; 
wire u5__abc_81276_new_n1545_; 
wire u5__abc_81276_new_n1546_; 
wire u5__abc_81276_new_n1547_; 
wire u5__abc_81276_new_n1548_; 
wire u5__abc_81276_new_n1549_; 
wire u5__abc_81276_new_n1550_; 
wire u5__abc_81276_new_n1551_; 
wire u5__abc_81276_new_n1552_; 
wire u5__abc_81276_new_n1553_; 
wire u5__abc_81276_new_n1554_; 
wire u5__abc_81276_new_n1555_; 
wire u5__abc_81276_new_n1556_; 
wire u5__abc_81276_new_n1557_; 
wire u5__abc_81276_new_n1558_; 
wire u5__abc_81276_new_n1559_; 
wire u5__abc_81276_new_n1560_; 
wire u5__abc_81276_new_n1561_; 
wire u5__abc_81276_new_n1562_; 
wire u5__abc_81276_new_n1563_; 
wire u5__abc_81276_new_n1564_; 
wire u5__abc_81276_new_n1565_; 
wire u5__abc_81276_new_n1566_; 
wire u5__abc_81276_new_n1567_; 
wire u5__abc_81276_new_n1568_; 
wire u5__abc_81276_new_n1569_; 
wire u5__abc_81276_new_n1570_; 
wire u5__abc_81276_new_n1571_; 
wire u5__abc_81276_new_n1572_; 
wire u5__abc_81276_new_n1573_; 
wire u5__abc_81276_new_n1574_; 
wire u5__abc_81276_new_n1575_; 
wire u5__abc_81276_new_n1576_; 
wire u5__abc_81276_new_n1577_; 
wire u5__abc_81276_new_n1578_; 
wire u5__abc_81276_new_n1579_; 
wire u5__abc_81276_new_n1580_; 
wire u5__abc_81276_new_n1581_; 
wire u5__abc_81276_new_n1582_; 
wire u5__abc_81276_new_n1583_; 
wire u5__abc_81276_new_n1584_; 
wire u5__abc_81276_new_n1585_; 
wire u5__abc_81276_new_n1586_; 
wire u5__abc_81276_new_n1587_; 
wire u5__abc_81276_new_n1588_; 
wire u5__abc_81276_new_n1589_; 
wire u5__abc_81276_new_n1590_; 
wire u5__abc_81276_new_n1591_; 
wire u5__abc_81276_new_n1592_; 
wire u5__abc_81276_new_n1593_; 
wire u5__abc_81276_new_n1594_; 
wire u5__abc_81276_new_n1595_; 
wire u5__abc_81276_new_n1596_; 
wire u5__abc_81276_new_n1597_; 
wire u5__abc_81276_new_n1598_; 
wire u5__abc_81276_new_n1599_; 
wire u5__abc_81276_new_n1600_; 
wire u5__abc_81276_new_n1601_; 
wire u5__abc_81276_new_n1602_; 
wire u5__abc_81276_new_n1603_; 
wire u5__abc_81276_new_n1604_; 
wire u5__abc_81276_new_n1605_; 
wire u5__abc_81276_new_n1606_; 
wire u5__abc_81276_new_n1607_; 
wire u5__abc_81276_new_n1608_; 
wire u5__abc_81276_new_n1609_; 
wire u5__abc_81276_new_n1610_; 
wire u5__abc_81276_new_n1611_; 
wire u5__abc_81276_new_n1612_; 
wire u5__abc_81276_new_n1613_; 
wire u5__abc_81276_new_n1614_; 
wire u5__abc_81276_new_n1615_; 
wire u5__abc_81276_new_n1616_; 
wire u5__abc_81276_new_n1617_; 
wire u5__abc_81276_new_n1618_; 
wire u5__abc_81276_new_n1619_; 
wire u5__abc_81276_new_n1620_; 
wire u5__abc_81276_new_n1621_; 
wire u5__abc_81276_new_n1622_; 
wire u5__abc_81276_new_n1623_; 
wire u5__abc_81276_new_n1624_; 
wire u5__abc_81276_new_n1625_; 
wire u5__abc_81276_new_n1626_; 
wire u5__abc_81276_new_n1627_; 
wire u5__abc_81276_new_n1628_; 
wire u5__abc_81276_new_n1629_; 
wire u5__abc_81276_new_n1630_; 
wire u5__abc_81276_new_n1631_; 
wire u5__abc_81276_new_n1632_; 
wire u5__abc_81276_new_n1633_; 
wire u5__abc_81276_new_n1634_; 
wire u5__abc_81276_new_n1636_; 
wire u5__abc_81276_new_n1637_; 
wire u5__abc_81276_new_n1638_; 
wire u5__abc_81276_new_n1640_; 
wire u5__abc_81276_new_n1641_; 
wire u5__abc_81276_new_n1642_; 
wire u5__abc_81276_new_n1643_; 
wire u5__abc_81276_new_n1644_; 
wire u5__abc_81276_new_n1645_; 
wire u5__abc_81276_new_n1646_; 
wire u5__abc_81276_new_n1647_; 
wire u5__abc_81276_new_n1648_; 
wire u5__abc_81276_new_n1649_; 
wire u5__abc_81276_new_n1650_; 
wire u5__abc_81276_new_n1651_; 
wire u5__abc_81276_new_n1652_; 
wire u5__abc_81276_new_n1653_; 
wire u5__abc_81276_new_n1654_; 
wire u5__abc_81276_new_n1655_; 
wire u5__abc_81276_new_n1656_; 
wire u5__abc_81276_new_n1657_; 
wire u5__abc_81276_new_n1658_; 
wire u5__abc_81276_new_n1659_; 
wire u5__abc_81276_new_n1660_; 
wire u5__abc_81276_new_n1662_; 
wire u5__abc_81276_new_n1663_; 
wire u5__abc_81276_new_n1665_; 
wire u5__abc_81276_new_n1666_; 
wire u5__abc_81276_new_n1667_; 
wire u5__abc_81276_new_n1668_; 
wire u5__abc_81276_new_n1669_; 
wire u5__abc_81276_new_n1670_; 
wire u5__abc_81276_new_n1671_; 
wire u5__abc_81276_new_n1672_; 
wire u5__abc_81276_new_n1673_; 
wire u5__abc_81276_new_n1675_; 
wire u5__abc_81276_new_n1676_; 
wire u5__abc_81276_new_n1678_; 
wire u5__abc_81276_new_n1679_; 
wire u5__abc_81276_new_n1680_; 
wire u5__abc_81276_new_n1681_; 
wire u5__abc_81276_new_n1682_; 
wire u5__abc_81276_new_n1682__bF_buf0; 
wire u5__abc_81276_new_n1682__bF_buf1; 
wire u5__abc_81276_new_n1682__bF_buf2; 
wire u5__abc_81276_new_n1682__bF_buf3; 
wire u5__abc_81276_new_n1682__bF_buf4; 
wire u5__abc_81276_new_n1683_; 
wire u5__abc_81276_new_n1684_; 
wire u5__abc_81276_new_n1685_; 
wire u5__abc_81276_new_n1686_; 
wire u5__abc_81276_new_n1687_; 
wire u5__abc_81276_new_n1688_; 
wire u5__abc_81276_new_n1689_; 
wire u5__abc_81276_new_n1690_; 
wire u5__abc_81276_new_n1691_; 
wire u5__abc_81276_new_n1692_; 
wire u5__abc_81276_new_n1693_; 
wire u5__abc_81276_new_n1694_; 
wire u5__abc_81276_new_n1695_; 
wire u5__abc_81276_new_n1696_; 
wire u5__abc_81276_new_n1697_; 
wire u5__abc_81276_new_n1698_; 
wire u5__abc_81276_new_n1699_; 
wire u5__abc_81276_new_n1700_; 
wire u5__abc_81276_new_n1701_; 
wire u5__abc_81276_new_n1702_; 
wire u5__abc_81276_new_n1703_; 
wire u5__abc_81276_new_n1704_; 
wire u5__abc_81276_new_n1705_; 
wire u5__abc_81276_new_n1706_; 
wire u5__abc_81276_new_n1707_; 
wire u5__abc_81276_new_n1708_; 
wire u5__abc_81276_new_n1709_; 
wire u5__abc_81276_new_n1710_; 
wire u5__abc_81276_new_n1711_; 
wire u5__abc_81276_new_n1712_; 
wire u5__abc_81276_new_n1713_; 
wire u5__abc_81276_new_n1714_; 
wire u5__abc_81276_new_n1715_; 
wire u5__abc_81276_new_n1716_; 
wire u5__abc_81276_new_n1717_; 
wire u5__abc_81276_new_n1718_; 
wire u5__abc_81276_new_n1719_; 
wire u5__abc_81276_new_n1720_; 
wire u5__abc_81276_new_n1721_; 
wire u5__abc_81276_new_n1722_; 
wire u5__abc_81276_new_n1724_; 
wire u5__abc_81276_new_n1725_; 
wire u5__abc_81276_new_n1727_; 
wire u5__abc_81276_new_n1728_; 
wire u5__abc_81276_new_n1729_; 
wire u5__abc_81276_new_n1730_; 
wire u5__abc_81276_new_n1731_; 
wire u5__abc_81276_new_n1732_; 
wire u5__abc_81276_new_n1733_; 
wire u5__abc_81276_new_n1734_; 
wire u5__abc_81276_new_n1735_; 
wire u5__abc_81276_new_n1736_; 
wire u5__abc_81276_new_n1737_; 
wire u5__abc_81276_new_n1738_; 
wire u5__abc_81276_new_n1740_; 
wire u5__abc_81276_new_n1741_; 
wire u5__abc_81276_new_n1743_; 
wire u5__abc_81276_new_n1744_; 
wire u5__abc_81276_new_n1745_; 
wire u5__abc_81276_new_n1746_; 
wire u5__abc_81276_new_n1747_; 
wire u5__abc_81276_new_n1748_; 
wire u5__abc_81276_new_n1749_; 
wire u5__abc_81276_new_n1750_; 
wire u5__abc_81276_new_n1751_; 
wire u5__abc_81276_new_n1752_; 
wire u5__abc_81276_new_n1753_; 
wire u5__abc_81276_new_n1754_; 
wire u5__abc_81276_new_n1755_; 
wire u5__abc_81276_new_n1756_; 
wire u5__abc_81276_new_n1757_; 
wire u5__abc_81276_new_n1758_; 
wire u5__abc_81276_new_n1759_; 
wire u5__abc_81276_new_n1760_; 
wire u5__abc_81276_new_n1761_; 
wire u5__abc_81276_new_n1762_; 
wire u5__abc_81276_new_n1763_; 
wire u5__abc_81276_new_n1764_; 
wire u5__abc_81276_new_n1765_; 
wire u5__abc_81276_new_n1766_; 
wire u5__abc_81276_new_n1767_; 
wire u5__abc_81276_new_n1768_; 
wire u5__abc_81276_new_n1769_; 
wire u5__abc_81276_new_n1770_; 
wire u5__abc_81276_new_n1771_; 
wire u5__abc_81276_new_n1772_; 
wire u5__abc_81276_new_n1773_; 
wire u5__abc_81276_new_n1774_; 
wire u5__abc_81276_new_n1775_; 
wire u5__abc_81276_new_n1776_; 
wire u5__abc_81276_new_n1777_; 
wire u5__abc_81276_new_n1778_; 
wire u5__abc_81276_new_n1779_; 
wire u5__abc_81276_new_n1780_; 
wire u5__abc_81276_new_n1781_; 
wire u5__abc_81276_new_n1782_; 
wire u5__abc_81276_new_n1783_; 
wire u5__abc_81276_new_n1784_; 
wire u5__abc_81276_new_n1785_; 
wire u5__abc_81276_new_n1786_; 
wire u5__abc_81276_new_n1787_; 
wire u5__abc_81276_new_n1788_; 
wire u5__abc_81276_new_n1789_; 
wire u5__abc_81276_new_n1790_; 
wire u5__abc_81276_new_n1791_; 
wire u5__abc_81276_new_n1793_; 
wire u5__abc_81276_new_n1794_; 
wire u5__abc_81276_new_n1795_; 
wire u5__abc_81276_new_n1796_; 
wire u5__abc_81276_new_n1797_; 
wire u5__abc_81276_new_n1798_; 
wire u5__abc_81276_new_n1799_; 
wire u5__abc_81276_new_n1800_; 
wire u5__abc_81276_new_n1801_; 
wire u5__abc_81276_new_n1802_; 
wire u5__abc_81276_new_n1803_; 
wire u5__abc_81276_new_n1804_; 
wire u5__abc_81276_new_n1805_; 
wire u5__abc_81276_new_n1807_; 
wire u5__abc_81276_new_n1808_; 
wire u5__abc_81276_new_n1809_; 
wire u5__abc_81276_new_n1810_; 
wire u5__abc_81276_new_n1811_; 
wire u5__abc_81276_new_n1812_; 
wire u5__abc_81276_new_n1813_; 
wire u5__abc_81276_new_n1815_; 
wire u5__abc_81276_new_n1816_; 
wire u5__abc_81276_new_n1817_; 
wire u5__abc_81276_new_n1818_; 
wire u5__abc_81276_new_n1819_; 
wire u5__abc_81276_new_n1820_; 
wire u5__abc_81276_new_n1821_; 
wire u5__abc_81276_new_n1822_; 
wire u5__abc_81276_new_n1823_; 
wire u5__abc_81276_new_n1824_; 
wire u5__abc_81276_new_n1825_; 
wire u5__abc_81276_new_n1826_; 
wire u5__abc_81276_new_n1827_; 
wire u5__abc_81276_new_n1828_; 
wire u5__abc_81276_new_n1829_; 
wire u5__abc_81276_new_n1830_; 
wire u5__abc_81276_new_n1831_; 
wire u5__abc_81276_new_n1832_; 
wire u5__abc_81276_new_n1833_; 
wire u5__abc_81276_new_n1834_; 
wire u5__abc_81276_new_n1835_; 
wire u5__abc_81276_new_n1836_; 
wire u5__abc_81276_new_n1837_; 
wire u5__abc_81276_new_n1838_; 
wire u5__abc_81276_new_n1839_; 
wire u5__abc_81276_new_n1840_; 
wire u5__abc_81276_new_n1841_; 
wire u5__abc_81276_new_n1842_; 
wire u5__abc_81276_new_n1843_; 
wire u5__abc_81276_new_n1844_; 
wire u5__abc_81276_new_n1845_; 
wire u5__abc_81276_new_n1846_; 
wire u5__abc_81276_new_n1847_; 
wire u5__abc_81276_new_n1848_; 
wire u5__abc_81276_new_n1849_; 
wire u5__abc_81276_new_n1850_; 
wire u5__abc_81276_new_n1851_; 
wire u5__abc_81276_new_n1852_; 
wire u5__abc_81276_new_n1853_; 
wire u5__abc_81276_new_n1854_; 
wire u5__abc_81276_new_n1855_; 
wire u5__abc_81276_new_n1856_; 
wire u5__abc_81276_new_n1857_; 
wire u5__abc_81276_new_n1858_; 
wire u5__abc_81276_new_n1859_; 
wire u5__abc_81276_new_n1860_; 
wire u5__abc_81276_new_n1861_; 
wire u5__abc_81276_new_n1862_; 
wire u5__abc_81276_new_n1863_; 
wire u5__abc_81276_new_n1864_; 
wire u5__abc_81276_new_n1865_; 
wire u5__abc_81276_new_n1867_; 
wire u5__abc_81276_new_n1868_; 
wire u5__abc_81276_new_n1870_; 
wire u5__abc_81276_new_n1871_; 
wire u5__abc_81276_new_n1872_; 
wire u5__abc_81276_new_n1873_; 
wire u5__abc_81276_new_n1874_; 
wire u5__abc_81276_new_n1875_; 
wire u5__abc_81276_new_n1876_; 
wire u5__abc_81276_new_n1877_; 
wire u5__abc_81276_new_n1878_; 
wire u5__abc_81276_new_n1879_; 
wire u5__abc_81276_new_n1880_; 
wire u5__abc_81276_new_n1881_; 
wire u5__abc_81276_new_n1882_; 
wire u5__abc_81276_new_n1883_; 
wire u5__abc_81276_new_n1884_; 
wire u5__abc_81276_new_n1885_; 
wire u5__abc_81276_new_n1886_; 
wire u5__abc_81276_new_n1887_; 
wire u5__abc_81276_new_n1888_; 
wire u5__abc_81276_new_n1889_; 
wire u5__abc_81276_new_n1890_; 
wire u5__abc_81276_new_n1891_; 
wire u5__abc_81276_new_n1892_; 
wire u5__abc_81276_new_n1893_; 
wire u5__abc_81276_new_n1894_; 
wire u5__abc_81276_new_n1895_; 
wire u5__abc_81276_new_n1896_; 
wire u5__abc_81276_new_n1897_; 
wire u5__abc_81276_new_n1898_; 
wire u5__abc_81276_new_n1899_; 
wire u5__abc_81276_new_n1900_; 
wire u5__abc_81276_new_n1901_; 
wire u5__abc_81276_new_n1902_; 
wire u5__abc_81276_new_n1903_; 
wire u5__abc_81276_new_n1904_; 
wire u5__abc_81276_new_n1905_; 
wire u5__abc_81276_new_n1906_; 
wire u5__abc_81276_new_n1907_; 
wire u5__abc_81276_new_n1908_; 
wire u5__abc_81276_new_n1909_; 
wire u5__abc_81276_new_n1910_; 
wire u5__abc_81276_new_n1911_; 
wire u5__abc_81276_new_n1912_; 
wire u5__abc_81276_new_n1913_; 
wire u5__abc_81276_new_n1914_; 
wire u5__abc_81276_new_n1915_; 
wire u5__abc_81276_new_n1916_; 
wire u5__abc_81276_new_n1917_; 
wire u5__abc_81276_new_n1918_; 
wire u5__abc_81276_new_n1919_; 
wire u5__abc_81276_new_n1920_; 
wire u5__abc_81276_new_n1921_; 
wire u5__abc_81276_new_n1922_; 
wire u5__abc_81276_new_n1923_; 
wire u5__abc_81276_new_n1924_; 
wire u5__abc_81276_new_n1925_; 
wire u5__abc_81276_new_n1926_; 
wire u5__abc_81276_new_n1927_; 
wire u5__abc_81276_new_n1928_; 
wire u5__abc_81276_new_n1929_; 
wire u5__abc_81276_new_n1930_; 
wire u5__abc_81276_new_n1931_; 
wire u5__abc_81276_new_n1932_; 
wire u5__abc_81276_new_n1933_; 
wire u5__abc_81276_new_n1934_; 
wire u5__abc_81276_new_n1935_; 
wire u5__abc_81276_new_n1936_; 
wire u5__abc_81276_new_n1937_; 
wire u5__abc_81276_new_n1938_; 
wire u5__abc_81276_new_n1939_; 
wire u5__abc_81276_new_n1940_; 
wire u5__abc_81276_new_n1941_; 
wire u5__abc_81276_new_n1942_; 
wire u5__abc_81276_new_n1943_; 
wire u5__abc_81276_new_n1944_; 
wire u5__abc_81276_new_n1945_; 
wire u5__abc_81276_new_n1946_; 
wire u5__abc_81276_new_n1947_; 
wire u5__abc_81276_new_n1948_; 
wire u5__abc_81276_new_n1949_; 
wire u5__abc_81276_new_n1950_; 
wire u5__abc_81276_new_n1951_; 
wire u5__abc_81276_new_n1952_; 
wire u5__abc_81276_new_n1953_; 
wire u5__abc_81276_new_n1954_; 
wire u5__abc_81276_new_n1955_; 
wire u5__abc_81276_new_n1956_; 
wire u5__abc_81276_new_n1957_; 
wire u5__abc_81276_new_n1958_; 
wire u5__abc_81276_new_n1959_; 
wire u5__abc_81276_new_n1960_; 
wire u5__abc_81276_new_n1961_; 
wire u5__abc_81276_new_n1962_; 
wire u5__abc_81276_new_n1963_; 
wire u5__abc_81276_new_n1964_; 
wire u5__abc_81276_new_n1965_; 
wire u5__abc_81276_new_n1966_; 
wire u5__abc_81276_new_n1967_; 
wire u5__abc_81276_new_n1968_; 
wire u5__abc_81276_new_n1969_; 
wire u5__abc_81276_new_n1970_; 
wire u5__abc_81276_new_n1971_; 
wire u5__abc_81276_new_n1972_; 
wire u5__abc_81276_new_n1973_; 
wire u5__abc_81276_new_n1974_; 
wire u5__abc_81276_new_n1975_; 
wire u5__abc_81276_new_n1976_; 
wire u5__abc_81276_new_n1977_; 
wire u5__abc_81276_new_n1978_; 
wire u5__abc_81276_new_n1979_; 
wire u5__abc_81276_new_n1980_; 
wire u5__abc_81276_new_n1981_; 
wire u5__abc_81276_new_n1982_; 
wire u5__abc_81276_new_n1983_; 
wire u5__abc_81276_new_n1984_; 
wire u5__abc_81276_new_n1985_; 
wire u5__abc_81276_new_n1986_; 
wire u5__abc_81276_new_n1987_; 
wire u5__abc_81276_new_n1988_; 
wire u5__abc_81276_new_n1989_; 
wire u5__abc_81276_new_n1990_; 
wire u5__abc_81276_new_n1991_; 
wire u5__abc_81276_new_n1992_; 
wire u5__abc_81276_new_n1993_; 
wire u5__abc_81276_new_n1994_; 
wire u5__abc_81276_new_n1995_; 
wire u5__abc_81276_new_n1996_; 
wire u5__abc_81276_new_n1997_; 
wire u5__abc_81276_new_n1998_; 
wire u5__abc_81276_new_n1999_; 
wire u5__abc_81276_new_n2000_; 
wire u5__abc_81276_new_n2001_; 
wire u5__abc_81276_new_n2002_; 
wire u5__abc_81276_new_n2003_; 
wire u5__abc_81276_new_n2004_; 
wire u5__abc_81276_new_n2005_; 
wire u5__abc_81276_new_n2006_; 
wire u5__abc_81276_new_n2007_; 
wire u5__abc_81276_new_n2008_; 
wire u5__abc_81276_new_n2009_; 
wire u5__abc_81276_new_n2010_; 
wire u5__abc_81276_new_n2011_; 
wire u5__abc_81276_new_n2012_; 
wire u5__abc_81276_new_n2013_; 
wire u5__abc_81276_new_n2014_; 
wire u5__abc_81276_new_n2015_; 
wire u5__abc_81276_new_n2016_; 
wire u5__abc_81276_new_n2017_; 
wire u5__abc_81276_new_n2018_; 
wire u5__abc_81276_new_n2019_; 
wire u5__abc_81276_new_n2020_; 
wire u5__abc_81276_new_n2021_; 
wire u5__abc_81276_new_n2022_; 
wire u5__abc_81276_new_n2023_; 
wire u5__abc_81276_new_n2024_; 
wire u5__abc_81276_new_n2025_; 
wire u5__abc_81276_new_n2026_; 
wire u5__abc_81276_new_n2027_; 
wire u5__abc_81276_new_n2028_; 
wire u5__abc_81276_new_n2029_; 
wire u5__abc_81276_new_n2030_; 
wire u5__abc_81276_new_n2031_; 
wire u5__abc_81276_new_n2032_; 
wire u5__abc_81276_new_n2033_; 
wire u5__abc_81276_new_n2034_; 
wire u5__abc_81276_new_n2035_; 
wire u5__abc_81276_new_n2036_; 
wire u5__abc_81276_new_n2037_; 
wire u5__abc_81276_new_n2038_; 
wire u5__abc_81276_new_n2039_; 
wire u5__abc_81276_new_n2040_; 
wire u5__abc_81276_new_n2041_; 
wire u5__abc_81276_new_n2042_; 
wire u5__abc_81276_new_n2043_; 
wire u5__abc_81276_new_n2044_; 
wire u5__abc_81276_new_n2045_; 
wire u5__abc_81276_new_n2046_; 
wire u5__abc_81276_new_n2047_; 
wire u5__abc_81276_new_n2048_; 
wire u5__abc_81276_new_n2049_; 
wire u5__abc_81276_new_n2050_; 
wire u5__abc_81276_new_n2051_; 
wire u5__abc_81276_new_n2052_; 
wire u5__abc_81276_new_n2053_; 
wire u5__abc_81276_new_n2054_; 
wire u5__abc_81276_new_n2055_; 
wire u5__abc_81276_new_n2056_; 
wire u5__abc_81276_new_n2057_; 
wire u5__abc_81276_new_n2058_; 
wire u5__abc_81276_new_n2059_; 
wire u5__abc_81276_new_n2060_; 
wire u5__abc_81276_new_n2061_; 
wire u5__abc_81276_new_n2062_; 
wire u5__abc_81276_new_n2063_; 
wire u5__abc_81276_new_n2064_; 
wire u5__abc_81276_new_n2065_; 
wire u5__abc_81276_new_n2066_; 
wire u5__abc_81276_new_n2067_; 
wire u5__abc_81276_new_n2068_; 
wire u5__abc_81276_new_n2069_; 
wire u5__abc_81276_new_n2070_; 
wire u5__abc_81276_new_n2071_; 
wire u5__abc_81276_new_n2072_; 
wire u5__abc_81276_new_n2073_; 
wire u5__abc_81276_new_n2074_; 
wire u5__abc_81276_new_n2075_; 
wire u5__abc_81276_new_n2076_; 
wire u5__abc_81276_new_n2077_; 
wire u5__abc_81276_new_n2078_; 
wire u5__abc_81276_new_n2079_; 
wire u5__abc_81276_new_n2080_; 
wire u5__abc_81276_new_n2081_; 
wire u5__abc_81276_new_n2082_; 
wire u5__abc_81276_new_n2083_; 
wire u5__abc_81276_new_n2084_; 
wire u5__abc_81276_new_n2085_; 
wire u5__abc_81276_new_n2086_; 
wire u5__abc_81276_new_n2087_; 
wire u5__abc_81276_new_n2088_; 
wire u5__abc_81276_new_n2089_; 
wire u5__abc_81276_new_n2090_; 
wire u5__abc_81276_new_n2091_; 
wire u5__abc_81276_new_n2092_; 
wire u5__abc_81276_new_n2093_; 
wire u5__abc_81276_new_n2094_; 
wire u5__abc_81276_new_n2095_; 
wire u5__abc_81276_new_n2096_; 
wire u5__abc_81276_new_n2097_; 
wire u5__abc_81276_new_n2098_; 
wire u5__abc_81276_new_n2099_; 
wire u5__abc_81276_new_n2100_; 
wire u5__abc_81276_new_n2101_; 
wire u5__abc_81276_new_n2102_; 
wire u5__abc_81276_new_n2103_; 
wire u5__abc_81276_new_n2104_; 
wire u5__abc_81276_new_n2105_; 
wire u5__abc_81276_new_n2106_; 
wire u5__abc_81276_new_n2107_; 
wire u5__abc_81276_new_n2108_; 
wire u5__abc_81276_new_n2109_; 
wire u5__abc_81276_new_n2110_; 
wire u5__abc_81276_new_n2111_; 
wire u5__abc_81276_new_n2112_; 
wire u5__abc_81276_new_n2113_; 
wire u5__abc_81276_new_n2114_; 
wire u5__abc_81276_new_n2115_; 
wire u5__abc_81276_new_n2116_; 
wire u5__abc_81276_new_n2117_; 
wire u5__abc_81276_new_n2118_; 
wire u5__abc_81276_new_n2119_; 
wire u5__abc_81276_new_n2120_; 
wire u5__abc_81276_new_n2121_; 
wire u5__abc_81276_new_n2122_; 
wire u5__abc_81276_new_n2123_; 
wire u5__abc_81276_new_n2124_; 
wire u5__abc_81276_new_n2125_; 
wire u5__abc_81276_new_n2126_; 
wire u5__abc_81276_new_n2127_; 
wire u5__abc_81276_new_n2128_; 
wire u5__abc_81276_new_n2129_; 
wire u5__abc_81276_new_n2130_; 
wire u5__abc_81276_new_n2131_; 
wire u5__abc_81276_new_n2132_; 
wire u5__abc_81276_new_n2133_; 
wire u5__abc_81276_new_n2134_; 
wire u5__abc_81276_new_n2135_; 
wire u5__abc_81276_new_n2136_; 
wire u5__abc_81276_new_n2137_; 
wire u5__abc_81276_new_n2138_; 
wire u5__abc_81276_new_n2139_; 
wire u5__abc_81276_new_n2140_; 
wire u5__abc_81276_new_n2141_; 
wire u5__abc_81276_new_n2142_; 
wire u5__abc_81276_new_n2143_; 
wire u5__abc_81276_new_n2144_; 
wire u5__abc_81276_new_n2145_; 
wire u5__abc_81276_new_n2146_; 
wire u5__abc_81276_new_n2147_; 
wire u5__abc_81276_new_n2148_; 
wire u5__abc_81276_new_n2149_; 
wire u5__abc_81276_new_n2150_; 
wire u5__abc_81276_new_n2151_; 
wire u5__abc_81276_new_n2152_; 
wire u5__abc_81276_new_n2153_; 
wire u5__abc_81276_new_n2154_; 
wire u5__abc_81276_new_n2155_; 
wire u5__abc_81276_new_n2156_; 
wire u5__abc_81276_new_n2157_; 
wire u5__abc_81276_new_n2158_; 
wire u5__abc_81276_new_n2159_; 
wire u5__abc_81276_new_n2160_; 
wire u5__abc_81276_new_n2161_; 
wire u5__abc_81276_new_n2162_; 
wire u5__abc_81276_new_n2163_; 
wire u5__abc_81276_new_n2164_; 
wire u5__abc_81276_new_n2165_; 
wire u5__abc_81276_new_n2166_; 
wire u5__abc_81276_new_n2167_; 
wire u5__abc_81276_new_n2168_; 
wire u5__abc_81276_new_n2169_; 
wire u5__abc_81276_new_n2170_; 
wire u5__abc_81276_new_n2171_; 
wire u5__abc_81276_new_n2172_; 
wire u5__abc_81276_new_n2173_; 
wire u5__abc_81276_new_n2174_; 
wire u5__abc_81276_new_n2175_; 
wire u5__abc_81276_new_n2176_; 
wire u5__abc_81276_new_n2177_; 
wire u5__abc_81276_new_n2178_; 
wire u5__abc_81276_new_n2179_; 
wire u5__abc_81276_new_n2180_; 
wire u5__abc_81276_new_n2181_; 
wire u5__abc_81276_new_n2182_; 
wire u5__abc_81276_new_n2183_; 
wire u5__abc_81276_new_n2184_; 
wire u5__abc_81276_new_n2185_; 
wire u5__abc_81276_new_n2186_; 
wire u5__abc_81276_new_n2187_; 
wire u5__abc_81276_new_n2188_; 
wire u5__abc_81276_new_n2189_; 
wire u5__abc_81276_new_n2190_; 
wire u5__abc_81276_new_n2191_; 
wire u5__abc_81276_new_n2192_; 
wire u5__abc_81276_new_n2193_; 
wire u5__abc_81276_new_n2194_; 
wire u5__abc_81276_new_n2195_; 
wire u5__abc_81276_new_n2196_; 
wire u5__abc_81276_new_n2197_; 
wire u5__abc_81276_new_n2198_; 
wire u5__abc_81276_new_n2199_; 
wire u5__abc_81276_new_n2200_; 
wire u5__abc_81276_new_n2201_; 
wire u5__abc_81276_new_n2202_; 
wire u5__abc_81276_new_n2203_; 
wire u5__abc_81276_new_n2204_; 
wire u5__abc_81276_new_n2205_; 
wire u5__abc_81276_new_n2206_; 
wire u5__abc_81276_new_n2207_; 
wire u5__abc_81276_new_n2208_; 
wire u5__abc_81276_new_n2209_; 
wire u5__abc_81276_new_n2210_; 
wire u5__abc_81276_new_n2211_; 
wire u5__abc_81276_new_n2212_; 
wire u5__abc_81276_new_n2213_; 
wire u5__abc_81276_new_n2214_; 
wire u5__abc_81276_new_n2215_; 
wire u5__abc_81276_new_n2216_; 
wire u5__abc_81276_new_n2217_; 
wire u5__abc_81276_new_n2218_; 
wire u5__abc_81276_new_n2219_; 
wire u5__abc_81276_new_n2220_; 
wire u5__abc_81276_new_n2221_; 
wire u5__abc_81276_new_n2222_; 
wire u5__abc_81276_new_n2223_; 
wire u5__abc_81276_new_n2224_; 
wire u5__abc_81276_new_n2225_; 
wire u5__abc_81276_new_n2226_; 
wire u5__abc_81276_new_n2227_; 
wire u5__abc_81276_new_n2228_; 
wire u5__abc_81276_new_n2229_; 
wire u5__abc_81276_new_n2230_; 
wire u5__abc_81276_new_n2231_; 
wire u5__abc_81276_new_n2232_; 
wire u5__abc_81276_new_n2233_; 
wire u5__abc_81276_new_n2234_; 
wire u5__abc_81276_new_n2235_; 
wire u5__abc_81276_new_n2236_; 
wire u5__abc_81276_new_n2237_; 
wire u5__abc_81276_new_n2238_; 
wire u5__abc_81276_new_n2239_; 
wire u5__abc_81276_new_n2240_; 
wire u5__abc_81276_new_n2241_; 
wire u5__abc_81276_new_n2242_; 
wire u5__abc_81276_new_n2243_; 
wire u5__abc_81276_new_n2244_; 
wire u5__abc_81276_new_n2245_; 
wire u5__abc_81276_new_n2246_; 
wire u5__abc_81276_new_n2247_; 
wire u5__abc_81276_new_n2248_; 
wire u5__abc_81276_new_n2249_; 
wire u5__abc_81276_new_n2250_; 
wire u5__abc_81276_new_n2251_; 
wire u5__abc_81276_new_n2252_; 
wire u5__abc_81276_new_n2253_; 
wire u5__abc_81276_new_n2254_; 
wire u5__abc_81276_new_n2255_; 
wire u5__abc_81276_new_n2256_; 
wire u5__abc_81276_new_n2257_; 
wire u5__abc_81276_new_n2258_; 
wire u5__abc_81276_new_n2259_; 
wire u5__abc_81276_new_n2260_; 
wire u5__abc_81276_new_n2261_; 
wire u5__abc_81276_new_n2262_; 
wire u5__abc_81276_new_n2263_; 
wire u5__abc_81276_new_n2264_; 
wire u5__abc_81276_new_n2265_; 
wire u5__abc_81276_new_n2266_; 
wire u5__abc_81276_new_n2267_; 
wire u5__abc_81276_new_n2268_; 
wire u5__abc_81276_new_n2269_; 
wire u5__abc_81276_new_n2270_; 
wire u5__abc_81276_new_n2271_; 
wire u5__abc_81276_new_n2272_; 
wire u5__abc_81276_new_n2273_; 
wire u5__abc_81276_new_n2274_; 
wire u5__abc_81276_new_n2275_; 
wire u5__abc_81276_new_n2276_; 
wire u5__abc_81276_new_n2277_; 
wire u5__abc_81276_new_n2278_; 
wire u5__abc_81276_new_n2279_; 
wire u5__abc_81276_new_n2280_; 
wire u5__abc_81276_new_n2281_; 
wire u5__abc_81276_new_n2282_; 
wire u5__abc_81276_new_n2283_; 
wire u5__abc_81276_new_n2284_; 
wire u5__abc_81276_new_n2285_; 
wire u5__abc_81276_new_n2286_; 
wire u5__abc_81276_new_n2287_; 
wire u5__abc_81276_new_n2288_; 
wire u5__abc_81276_new_n2289_; 
wire u5__abc_81276_new_n2290_; 
wire u5__abc_81276_new_n2291_; 
wire u5__abc_81276_new_n2292_; 
wire u5__abc_81276_new_n2293_; 
wire u5__abc_81276_new_n2294_; 
wire u5__abc_81276_new_n2295_; 
wire u5__abc_81276_new_n2296_; 
wire u5__abc_81276_new_n2297_; 
wire u5__abc_81276_new_n2298_; 
wire u5__abc_81276_new_n2299_; 
wire u5__abc_81276_new_n2300_; 
wire u5__abc_81276_new_n2302_; 
wire u5__abc_81276_new_n2303_; 
wire u5__abc_81276_new_n2304_; 
wire u5__abc_81276_new_n2305_; 
wire u5__abc_81276_new_n2306_; 
wire u5__abc_81276_new_n2307_; 
wire u5__abc_81276_new_n2308_; 
wire u5__abc_81276_new_n2309_; 
wire u5__abc_81276_new_n2310_; 
wire u5__abc_81276_new_n2311_; 
wire u5__abc_81276_new_n2312_; 
wire u5__abc_81276_new_n2313_; 
wire u5__abc_81276_new_n2314_; 
wire u5__abc_81276_new_n2315_; 
wire u5__abc_81276_new_n2316_; 
wire u5__abc_81276_new_n2317_; 
wire u5__abc_81276_new_n2318_; 
wire u5__abc_81276_new_n2319_; 
wire u5__abc_81276_new_n2320_; 
wire u5__abc_81276_new_n2321_; 
wire u5__abc_81276_new_n2322_; 
wire u5__abc_81276_new_n2323_; 
wire u5__abc_81276_new_n2324_; 
wire u5__abc_81276_new_n2325_; 
wire u5__abc_81276_new_n2326_; 
wire u5__abc_81276_new_n2327_; 
wire u5__abc_81276_new_n2328_; 
wire u5__abc_81276_new_n2329_; 
wire u5__abc_81276_new_n2330_; 
wire u5__abc_81276_new_n2331_; 
wire u5__abc_81276_new_n2332_; 
wire u5__abc_81276_new_n2333_; 
wire u5__abc_81276_new_n2334_; 
wire u5__abc_81276_new_n2335_; 
wire u5__abc_81276_new_n2336_; 
wire u5__abc_81276_new_n2337_; 
wire u5__abc_81276_new_n2338_; 
wire u5__abc_81276_new_n2339_; 
wire u5__abc_81276_new_n2340_; 
wire u5__abc_81276_new_n2342_; 
wire u5__abc_81276_new_n2343_; 
wire u5__abc_81276_new_n2344_; 
wire u5__abc_81276_new_n2345_; 
wire u5__abc_81276_new_n2346_; 
wire u5__abc_81276_new_n2347_; 
wire u5__abc_81276_new_n2348_; 
wire u5__abc_81276_new_n2349_; 
wire u5__abc_81276_new_n2351_; 
wire u5__abc_81276_new_n2352_; 
wire u5__abc_81276_new_n2353_; 
wire u5__abc_81276_new_n2354_; 
wire u5__abc_81276_new_n2355_; 
wire u5__abc_81276_new_n2356_; 
wire u5__abc_81276_new_n2357_; 
wire u5__abc_81276_new_n2358_; 
wire u5__abc_81276_new_n2359_; 
wire u5__abc_81276_new_n2361_; 
wire u5__abc_81276_new_n2362_; 
wire u5__abc_81276_new_n2363_; 
wire u5__abc_81276_new_n2364_; 
wire u5__abc_81276_new_n2365_; 
wire u5__abc_81276_new_n2366_; 
wire u5__abc_81276_new_n2367_; 
wire u5__abc_81276_new_n2368_; 
wire u5__abc_81276_new_n2369_; 
wire u5__abc_81276_new_n2371_; 
wire u5__abc_81276_new_n2372_; 
wire u5__abc_81276_new_n2373_; 
wire u5__abc_81276_new_n2374_; 
wire u5__abc_81276_new_n2375_; 
wire u5__abc_81276_new_n2376_; 
wire u5__abc_81276_new_n2377_; 
wire u5__abc_81276_new_n2378_; 
wire u5__abc_81276_new_n2380_; 
wire u5__abc_81276_new_n2381_; 
wire u5__abc_81276_new_n2382_; 
wire u5__abc_81276_new_n2383_; 
wire u5__abc_81276_new_n2384_; 
wire u5__abc_81276_new_n2385_; 
wire u5__abc_81276_new_n2386_; 
wire u5__abc_81276_new_n2387_; 
wire u5__abc_81276_new_n2389_; 
wire u5__abc_81276_new_n2390_; 
wire u5__abc_81276_new_n2391_; 
wire u5__abc_81276_new_n2392_; 
wire u5__abc_81276_new_n2393_; 
wire u5__abc_81276_new_n2394_; 
wire u5__abc_81276_new_n2395_; 
wire u5__abc_81276_new_n2396_; 
wire u5__abc_81276_new_n2398_; 
wire u5__abc_81276_new_n2399_; 
wire u5__abc_81276_new_n2400_; 
wire u5__abc_81276_new_n2401_; 
wire u5__abc_81276_new_n2402_; 
wire u5__abc_81276_new_n2403_; 
wire u5__abc_81276_new_n2404_; 
wire u5__abc_81276_new_n2405_; 
wire u5__abc_81276_new_n2406_; 
wire u5__abc_81276_new_n2407_; 
wire u5__abc_81276_new_n2408_; 
wire u5__abc_81276_new_n2409_; 
wire u5__abc_81276_new_n2410_; 
wire u5__abc_81276_new_n2412_; 
wire u5__abc_81276_new_n2413_; 
wire u5__abc_81276_new_n2414_; 
wire u5__abc_81276_new_n2415_; 
wire u5__abc_81276_new_n2416_; 
wire u5__abc_81276_new_n2417_; 
wire u5__abc_81276_new_n2418_; 
wire u5__abc_81276_new_n2419_; 
wire u5__abc_81276_new_n2420_; 
wire u5__abc_81276_new_n2421_; 
wire u5__abc_81276_new_n2423_; 
wire u5__abc_81276_new_n2424_; 
wire u5__abc_81276_new_n2425_; 
wire u5__abc_81276_new_n2426_; 
wire u5__abc_81276_new_n2427_; 
wire u5__abc_81276_new_n2428_; 
wire u5__abc_81276_new_n2429_; 
wire u5__abc_81276_new_n2430_; 
wire u5__abc_81276_new_n2432_; 
wire u5__abc_81276_new_n2433_; 
wire u5__abc_81276_new_n2434_; 
wire u5__abc_81276_new_n2435_; 
wire u5__abc_81276_new_n2436_; 
wire u5__abc_81276_new_n2437_; 
wire u5__abc_81276_new_n2438_; 
wire u5__abc_81276_new_n2439_; 
wire u5__abc_81276_new_n2440_; 
wire u5__abc_81276_new_n2441_; 
wire u5__abc_81276_new_n2442_; 
wire u5__abc_81276_new_n2443_; 
wire u5__abc_81276_new_n2444_; 
wire u5__abc_81276_new_n2446_; 
wire u5__abc_81276_new_n2447_; 
wire u5__abc_81276_new_n2448_; 
wire u5__abc_81276_new_n2449_; 
wire u5__abc_81276_new_n2450_; 
wire u5__abc_81276_new_n2451_; 
wire u5__abc_81276_new_n2452_; 
wire u5__abc_81276_new_n2453_; 
wire u5__abc_81276_new_n2454_; 
wire u5__abc_81276_new_n2455_; 
wire u5__abc_81276_new_n2456_; 
wire u5__abc_81276_new_n2457_; 
wire u5__abc_81276_new_n2458_; 
wire u5__abc_81276_new_n2459_; 
wire u5__abc_81276_new_n2460_; 
wire u5__abc_81276_new_n2461_; 
wire u5__abc_81276_new_n2462_; 
wire u5__abc_81276_new_n2463_; 
wire u5__abc_81276_new_n2464_; 
wire u5__abc_81276_new_n2465_; 
wire u5__abc_81276_new_n2466_; 
wire u5__abc_81276_new_n2467_; 
wire u5__abc_81276_new_n2468_; 
wire u5__abc_81276_new_n2469_; 
wire u5__abc_81276_new_n2470_; 
wire u5__abc_81276_new_n2471_; 
wire u5__abc_81276_new_n2472_; 
wire u5__abc_81276_new_n2473_; 
wire u5__abc_81276_new_n2475_; 
wire u5__abc_81276_new_n2476_; 
wire u5__abc_81276_new_n2477_; 
wire u5__abc_81276_new_n2478_; 
wire u5__abc_81276_new_n2479_; 
wire u5__abc_81276_new_n2481_; 
wire u5__abc_81276_new_n2482_; 
wire u5__abc_81276_new_n2483_; 
wire u5__abc_81276_new_n2485_; 
wire u5__abc_81276_new_n2486_; 
wire u5__abc_81276_new_n2487_; 
wire u5__abc_81276_new_n2488_; 
wire u5__abc_81276_new_n2490_; 
wire u5__abc_81276_new_n2491_; 
wire u5__abc_81276_new_n2492_; 
wire u5__abc_81276_new_n2493_; 
wire u5__abc_81276_new_n2494_; 
wire u5__abc_81276_new_n2495_; 
wire u5__abc_81276_new_n2496_; 
wire u5__abc_81276_new_n2497_; 
wire u5__abc_81276_new_n2498_; 
wire u5__abc_81276_new_n2499_; 
wire u5__abc_81276_new_n2500_; 
wire u5__abc_81276_new_n2501_; 
wire u5__abc_81276_new_n2502_; 
wire u5__abc_81276_new_n2503_; 
wire u5__abc_81276_new_n2504_; 
wire u5__abc_81276_new_n2505_; 
wire u5__abc_81276_new_n2506_; 
wire u5__abc_81276_new_n2507_; 
wire u5__abc_81276_new_n2508_; 
wire u5__abc_81276_new_n2509_; 
wire u5__abc_81276_new_n2510_; 
wire u5__abc_81276_new_n2511_; 
wire u5__abc_81276_new_n2512_; 
wire u5__abc_81276_new_n2513_; 
wire u5__abc_81276_new_n2514_; 
wire u5__abc_81276_new_n2515_; 
wire u5__abc_81276_new_n2516_; 
wire u5__abc_81276_new_n2517_; 
wire u5__abc_81276_new_n2518_; 
wire u5__abc_81276_new_n2519_; 
wire u5__abc_81276_new_n2520_; 
wire u5__abc_81276_new_n2521_; 
wire u5__abc_81276_new_n2522_; 
wire u5__abc_81276_new_n2523_; 
wire u5__abc_81276_new_n2524_; 
wire u5__abc_81276_new_n2525_; 
wire u5__abc_81276_new_n2526_; 
wire u5__abc_81276_new_n2527_; 
wire u5__abc_81276_new_n2528_; 
wire u5__abc_81276_new_n2529_; 
wire u5__abc_81276_new_n2530_; 
wire u5__abc_81276_new_n2531_; 
wire u5__abc_81276_new_n2532_; 
wire u5__abc_81276_new_n2533_; 
wire u5__abc_81276_new_n2534_; 
wire u5__abc_81276_new_n2535_; 
wire u5__abc_81276_new_n2536_; 
wire u5__abc_81276_new_n2537_; 
wire u5__abc_81276_new_n2538_; 
wire u5__abc_81276_new_n2539_; 
wire u5__abc_81276_new_n2540_; 
wire u5__abc_81276_new_n2541_; 
wire u5__abc_81276_new_n2542_; 
wire u5__abc_81276_new_n2543_; 
wire u5__abc_81276_new_n2544_; 
wire u5__abc_81276_new_n2545_; 
wire u5__abc_81276_new_n2546_; 
wire u5__abc_81276_new_n2547_; 
wire u5__abc_81276_new_n2548_; 
wire u5__abc_81276_new_n2549_; 
wire u5__abc_81276_new_n2550_; 
wire u5__abc_81276_new_n2551_; 
wire u5__abc_81276_new_n2552_; 
wire u5__abc_81276_new_n2553_; 
wire u5__abc_81276_new_n2554_; 
wire u5__abc_81276_new_n2555_; 
wire u5__abc_81276_new_n2556_; 
wire u5__abc_81276_new_n2557_; 
wire u5__abc_81276_new_n2558_; 
wire u5__abc_81276_new_n2559_; 
wire u5__abc_81276_new_n2560_; 
wire u5__abc_81276_new_n2561_; 
wire u5__abc_81276_new_n2562_; 
wire u5__abc_81276_new_n2563_; 
wire u5__abc_81276_new_n2564_; 
wire u5__abc_81276_new_n2565_; 
wire u5__abc_81276_new_n2566_; 
wire u5__abc_81276_new_n2567_; 
wire u5__abc_81276_new_n2568_; 
wire u5__abc_81276_new_n2569_; 
wire u5__abc_81276_new_n2570_; 
wire u5__abc_81276_new_n2571_; 
wire u5__abc_81276_new_n2572_; 
wire u5__abc_81276_new_n2573_; 
wire u5__abc_81276_new_n2574_; 
wire u5__abc_81276_new_n2575_; 
wire u5__abc_81276_new_n2576_; 
wire u5__abc_81276_new_n2577_; 
wire u5__abc_81276_new_n2578_; 
wire u5__abc_81276_new_n2579_; 
wire u5__abc_81276_new_n2580_; 
wire u5__abc_81276_new_n2581_; 
wire u5__abc_81276_new_n2582_; 
wire u5__abc_81276_new_n2583_; 
wire u5__abc_81276_new_n2584_; 
wire u5__abc_81276_new_n2585_; 
wire u5__abc_81276_new_n2586_; 
wire u5__abc_81276_new_n2587_; 
wire u5__abc_81276_new_n2588_; 
wire u5__abc_81276_new_n2589_; 
wire u5__abc_81276_new_n2590_; 
wire u5__abc_81276_new_n2591_; 
wire u5__abc_81276_new_n2592_; 
wire u5__abc_81276_new_n2593_; 
wire u5__abc_81276_new_n2594_; 
wire u5__abc_81276_new_n2595_; 
wire u5__abc_81276_new_n2596_; 
wire u5__abc_81276_new_n2597_; 
wire u5__abc_81276_new_n2598_; 
wire u5__abc_81276_new_n2599_; 
wire u5__abc_81276_new_n2600_; 
wire u5__abc_81276_new_n2601_; 
wire u5__abc_81276_new_n2602_; 
wire u5__abc_81276_new_n2603_; 
wire u5__abc_81276_new_n2604_; 
wire u5__abc_81276_new_n2605_; 
wire u5__abc_81276_new_n2606_; 
wire u5__abc_81276_new_n2607_; 
wire u5__abc_81276_new_n2608_; 
wire u5__abc_81276_new_n2609_; 
wire u5__abc_81276_new_n2610_; 
wire u5__abc_81276_new_n2611_; 
wire u5__abc_81276_new_n2612_; 
wire u5__abc_81276_new_n2613_; 
wire u5__abc_81276_new_n2614_; 
wire u5__abc_81276_new_n2615_; 
wire u5__abc_81276_new_n2616_; 
wire u5__abc_81276_new_n2617_; 
wire u5__abc_81276_new_n2618_; 
wire u5__abc_81276_new_n2619_; 
wire u5__abc_81276_new_n2620_; 
wire u5__abc_81276_new_n2621_; 
wire u5__abc_81276_new_n2622_; 
wire u5__abc_81276_new_n2623_; 
wire u5__abc_81276_new_n2624_; 
wire u5__abc_81276_new_n2625_; 
wire u5__abc_81276_new_n2626_; 
wire u5__abc_81276_new_n2627_; 
wire u5__abc_81276_new_n2628_; 
wire u5__abc_81276_new_n2629_; 
wire u5__abc_81276_new_n2630_; 
wire u5__abc_81276_new_n2631_; 
wire u5__abc_81276_new_n2632_; 
wire u5__abc_81276_new_n2633_; 
wire u5__abc_81276_new_n2634_; 
wire u5__abc_81276_new_n2635_; 
wire u5__abc_81276_new_n2636_; 
wire u5__abc_81276_new_n2637_; 
wire u5__abc_81276_new_n2638_; 
wire u5__abc_81276_new_n2639_; 
wire u5__abc_81276_new_n2640_; 
wire u5__abc_81276_new_n2641_; 
wire u5__abc_81276_new_n2642_; 
wire u5__abc_81276_new_n2643_; 
wire u5__abc_81276_new_n2644_; 
wire u5__abc_81276_new_n2645_; 
wire u5__abc_81276_new_n2646_; 
wire u5__abc_81276_new_n2647_; 
wire u5__abc_81276_new_n2648_; 
wire u5__abc_81276_new_n2649_; 
wire u5__abc_81276_new_n2650_; 
wire u5__abc_81276_new_n2651_; 
wire u5__abc_81276_new_n2652_; 
wire u5__abc_81276_new_n2653_; 
wire u5__abc_81276_new_n2654_; 
wire u5__abc_81276_new_n2655_; 
wire u5__abc_81276_new_n2656_; 
wire u5__abc_81276_new_n2657_; 
wire u5__abc_81276_new_n2658_; 
wire u5__abc_81276_new_n2659_; 
wire u5__abc_81276_new_n2660_; 
wire u5__abc_81276_new_n2661_; 
wire u5__abc_81276_new_n2662_; 
wire u5__abc_81276_new_n2663_; 
wire u5__abc_81276_new_n2664_; 
wire u5__abc_81276_new_n2665_; 
wire u5__abc_81276_new_n2666_; 
wire u5__abc_81276_new_n2667_; 
wire u5__abc_81276_new_n2668_; 
wire u5__abc_81276_new_n2669_; 
wire u5__abc_81276_new_n2670_; 
wire u5__abc_81276_new_n2671_; 
wire u5__abc_81276_new_n2672_; 
wire u5__abc_81276_new_n2673_; 
wire u5__abc_81276_new_n2674_; 
wire u5__abc_81276_new_n2675_; 
wire u5__abc_81276_new_n2677_; 
wire u5__abc_81276_new_n2678_; 
wire u5__abc_81276_new_n2679_; 
wire u5__abc_81276_new_n2680_; 
wire u5__abc_81276_new_n2681_; 
wire u5__abc_81276_new_n2682_; 
wire u5__abc_81276_new_n2683_; 
wire u5__abc_81276_new_n2684_; 
wire u5__abc_81276_new_n2685_; 
wire u5__abc_81276_new_n2686_; 
wire u5__abc_81276_new_n2687_; 
wire u5__abc_81276_new_n2688_; 
wire u5__abc_81276_new_n2689_; 
wire u5__abc_81276_new_n2690_; 
wire u5__abc_81276_new_n2691_; 
wire u5__abc_81276_new_n2692_; 
wire u5__abc_81276_new_n2693_; 
wire u5__abc_81276_new_n2694_; 
wire u5__abc_81276_new_n2695_; 
wire u5__abc_81276_new_n2696_; 
wire u5__abc_81276_new_n2697_; 
wire u5__abc_81276_new_n2698_; 
wire u5__abc_81276_new_n2699_; 
wire u5__abc_81276_new_n2700_; 
wire u5__abc_81276_new_n2701_; 
wire u5__abc_81276_new_n2702_; 
wire u5__abc_81276_new_n2703_; 
wire u5__abc_81276_new_n2704_; 
wire u5__abc_81276_new_n2705_; 
wire u5__abc_81276_new_n2706_; 
wire u5__abc_81276_new_n2707_; 
wire u5__abc_81276_new_n2708_; 
wire u5__abc_81276_new_n2709_; 
wire u5__abc_81276_new_n2710_; 
wire u5__abc_81276_new_n2711_; 
wire u5__abc_81276_new_n2712_; 
wire u5__abc_81276_new_n2713_; 
wire u5__abc_81276_new_n2714_; 
wire u5__abc_81276_new_n2715_; 
wire u5__abc_81276_new_n2716_; 
wire u5__abc_81276_new_n2717_; 
wire u5__abc_81276_new_n2718_; 
wire u5__abc_81276_new_n2719_; 
wire u5__abc_81276_new_n2720_; 
wire u5__abc_81276_new_n2721_; 
wire u5__abc_81276_new_n2722_; 
wire u5__abc_81276_new_n2724_; 
wire u5__abc_81276_new_n2725_; 
wire u5__abc_81276_new_n2726_; 
wire u5__abc_81276_new_n2727_; 
wire u5__abc_81276_new_n2728_; 
wire u5__abc_81276_new_n2729_; 
wire u5__abc_81276_new_n2730_; 
wire u5__abc_81276_new_n2731_; 
wire u5__abc_81276_new_n2732_; 
wire u5__abc_81276_new_n2733_; 
wire u5__abc_81276_new_n2734_; 
wire u5__abc_81276_new_n2735_; 
wire u5__abc_81276_new_n2736_; 
wire u5__abc_81276_new_n2737_; 
wire u5__abc_81276_new_n2738_; 
wire u5__abc_81276_new_n2739_; 
wire u5__abc_81276_new_n2740_; 
wire u5__abc_81276_new_n2741_; 
wire u5__abc_81276_new_n2742_; 
wire u5__abc_81276_new_n2743_; 
wire u5__abc_81276_new_n2744_; 
wire u5__abc_81276_new_n2745_; 
wire u5__abc_81276_new_n2746_; 
wire u5__abc_81276_new_n2747_; 
wire u5__abc_81276_new_n2748_; 
wire u5__abc_81276_new_n2749_; 
wire u5__abc_81276_new_n2750_; 
wire u5__abc_81276_new_n2751_; 
wire u5__abc_81276_new_n2752_; 
wire u5__abc_81276_new_n2753_; 
wire u5__abc_81276_new_n2754_; 
wire u5__abc_81276_new_n2755_; 
wire u5__abc_81276_new_n2756_; 
wire u5__abc_81276_new_n2757_; 
wire u5__abc_81276_new_n2758_; 
wire u5__abc_81276_new_n2759_; 
wire u5__abc_81276_new_n2760_; 
wire u5__abc_81276_new_n2761_; 
wire u5__abc_81276_new_n2762_; 
wire u5__abc_81276_new_n2763_; 
wire u5__abc_81276_new_n2764_; 
wire u5__abc_81276_new_n2765_; 
wire u5__abc_81276_new_n2766_; 
wire u5__abc_81276_new_n2767_; 
wire u5__abc_81276_new_n2768_; 
wire u5__abc_81276_new_n2769_; 
wire u5__abc_81276_new_n2770_; 
wire u5__abc_81276_new_n2771_; 
wire u5__abc_81276_new_n2772_; 
wire u5__abc_81276_new_n2773_; 
wire u5__abc_81276_new_n2774_; 
wire u5__abc_81276_new_n2775_; 
wire u5__abc_81276_new_n2776_; 
wire u5__abc_81276_new_n2777_; 
wire u5__abc_81276_new_n2778_; 
wire u5__abc_81276_new_n2779_; 
wire u5__abc_81276_new_n2780_; 
wire u5__abc_81276_new_n2781_; 
wire u5__abc_81276_new_n2782_; 
wire u5__abc_81276_new_n2783_; 
wire u5__abc_81276_new_n2784_; 
wire u5__abc_81276_new_n2785_; 
wire u5__abc_81276_new_n2786_; 
wire u5__abc_81276_new_n2787_; 
wire u5__abc_81276_new_n2788_; 
wire u5__abc_81276_new_n2789_; 
wire u5__abc_81276_new_n2790_; 
wire u5__abc_81276_new_n2791_; 
wire u5__abc_81276_new_n2792_; 
wire u5__abc_81276_new_n2793_; 
wire u5__abc_81276_new_n2794_; 
wire u5__abc_81276_new_n2795_; 
wire u5__abc_81276_new_n2796_; 
wire u5__abc_81276_new_n2797_; 
wire u5__abc_81276_new_n2798_; 
wire u5__abc_81276_new_n2799_; 
wire u5__abc_81276_new_n2800_; 
wire u5__abc_81276_new_n2801_; 
wire u5__abc_81276_new_n2802_; 
wire u5__abc_81276_new_n2803_; 
wire u5__abc_81276_new_n2804_; 
wire u5__abc_81276_new_n2805_; 
wire u5__abc_81276_new_n2807_; 
wire u5__abc_81276_new_n2808_; 
wire u5__abc_81276_new_n2809_; 
wire u5__abc_81276_new_n2810_; 
wire u5__abc_81276_new_n2811_; 
wire u5__abc_81276_new_n2812_; 
wire u5__abc_81276_new_n2813_; 
wire u5__abc_81276_new_n2814_; 
wire u5__abc_81276_new_n2815_; 
wire u5__abc_81276_new_n2816_; 
wire u5__abc_81276_new_n2817_; 
wire u5__abc_81276_new_n2818_; 
wire u5__abc_81276_new_n2819_; 
wire u5__abc_81276_new_n2820_; 
wire u5__abc_81276_new_n2821_; 
wire u5__abc_81276_new_n2822_; 
wire u5__abc_81276_new_n2823_; 
wire u5__abc_81276_new_n2824_; 
wire u5__abc_81276_new_n2825_; 
wire u5__abc_81276_new_n2826_; 
wire u5__abc_81276_new_n2827_; 
wire u5__abc_81276_new_n2828_; 
wire u5__abc_81276_new_n2829_; 
wire u5__abc_81276_new_n2830_; 
wire u5__abc_81276_new_n2831_; 
wire u5__abc_81276_new_n2832_; 
wire u5__abc_81276_new_n2833_; 
wire u5__abc_81276_new_n2834_; 
wire u5__abc_81276_new_n2835_; 
wire u5__abc_81276_new_n2836_; 
wire u5__abc_81276_new_n2837_; 
wire u5__abc_81276_new_n2838_; 
wire u5__abc_81276_new_n2839_; 
wire u5__abc_81276_new_n2840_; 
wire u5__abc_81276_new_n2841_; 
wire u5__abc_81276_new_n2842_; 
wire u5__abc_81276_new_n2843_; 
wire u5__abc_81276_new_n2844_; 
wire u5__abc_81276_new_n2845_; 
wire u5__abc_81276_new_n2846_; 
wire u5__abc_81276_new_n2847_; 
wire u5__abc_81276_new_n2848_; 
wire u5__abc_81276_new_n2849_; 
wire u5__abc_81276_new_n2850_; 
wire u5__abc_81276_new_n2851_; 
wire u5__abc_81276_new_n2852_; 
wire u5__abc_81276_new_n2853_; 
wire u5__abc_81276_new_n2854_; 
wire u5__abc_81276_new_n2855_; 
wire u5__abc_81276_new_n2856_; 
wire u5__abc_81276_new_n2857_; 
wire u5__abc_81276_new_n2858_; 
wire u5__abc_81276_new_n2859_; 
wire u5__abc_81276_new_n2860_; 
wire u5__abc_81276_new_n2861_; 
wire u5__abc_81276_new_n2863_; 
wire u5__abc_81276_new_n2864_; 
wire u5__abc_81276_new_n2865_; 
wire u5__abc_81276_new_n2866_; 
wire u5__abc_81276_new_n2867_; 
wire u5__abc_81276_new_n2868_; 
wire u5__abc_81276_new_n2869_; 
wire u5__abc_81276_new_n2870_; 
wire u5__abc_81276_new_n2871_; 
wire u5__abc_81276_new_n2872_; 
wire u5__abc_81276_new_n2873_; 
wire u5__abc_81276_new_n2874_; 
wire u5__abc_81276_new_n2875_; 
wire u5__abc_81276_new_n2876_; 
wire u5__abc_81276_new_n2877_; 
wire u5__abc_81276_new_n2878_; 
wire u5__abc_81276_new_n2879_; 
wire u5__abc_81276_new_n2880_; 
wire u5__abc_81276_new_n2881_; 
wire u5__abc_81276_new_n2883_; 
wire u5__abc_81276_new_n2884_; 
wire u5__abc_81276_new_n2885_; 
wire u5__abc_81276_new_n2886_; 
wire u5__abc_81276_new_n2887_; 
wire u5__abc_81276_new_n2888_; 
wire u5__abc_81276_new_n2889_; 
wire u5__abc_81276_new_n2890_; 
wire u5__abc_81276_new_n2891_; 
wire u5__abc_81276_new_n2893_; 
wire u5__abc_81276_new_n2894_; 
wire u5__abc_81276_new_n2895_; 
wire u5__abc_81276_new_n2896_; 
wire u5__abc_81276_new_n2897_; 
wire u5__abc_81276_new_n2898_; 
wire u5__abc_81276_new_n2899_; 
wire u5__abc_81276_new_n2900_; 
wire u5__abc_81276_new_n2901_; 
wire u5__abc_81276_new_n2902_; 
wire u5__abc_81276_new_n2904_; 
wire u5__abc_81276_new_n2905_; 
wire u5__abc_81276_new_n2906_; 
wire u5__abc_81276_new_n2907_; 
wire u5__abc_81276_new_n2908_; 
wire u5__abc_81276_new_n2909_; 
wire u5__abc_81276_new_n2910_; 
wire u5__abc_81276_new_n2912_; 
wire u5__abc_81276_new_n2913_; 
wire u5__abc_81276_new_n2914_; 
wire u5__abc_81276_new_n2915_; 
wire u5__abc_81276_new_n2916_; 
wire u5__abc_81276_new_n2917_; 
wire u5__abc_81276_new_n2918_; 
wire u5__abc_81276_new_n2919_; 
wire u5__abc_81276_new_n2920_; 
wire u5__abc_81276_new_n2921_; 
wire u5__abc_81276_new_n2922_; 
wire u5__abc_81276_new_n2923_; 
wire u5__abc_81276_new_n2924_; 
wire u5__abc_81276_new_n2925_; 
wire u5__abc_81276_new_n2926_; 
wire u5__abc_81276_new_n2927_; 
wire u5__abc_81276_new_n2928_; 
wire u5__abc_81276_new_n2929_; 
wire u5__abc_81276_new_n2930_; 
wire u5__abc_81276_new_n2931_; 
wire u5__abc_81276_new_n2932_; 
wire u5__abc_81276_new_n2933_; 
wire u5__abc_81276_new_n2934_; 
wire u5__abc_81276_new_n2935_; 
wire u5__abc_81276_new_n2936_; 
wire u5__abc_81276_new_n2937_; 
wire u5__abc_81276_new_n2938_; 
wire u5__abc_81276_new_n2939_; 
wire u5__abc_81276_new_n2940_; 
wire u5__abc_81276_new_n2941_; 
wire u5__abc_81276_new_n2942_; 
wire u5__abc_81276_new_n2943_; 
wire u5__abc_81276_new_n2944_; 
wire u5__abc_81276_new_n2945_; 
wire u5__abc_81276_new_n2946_; 
wire u5__abc_81276_new_n2947_; 
wire u5__abc_81276_new_n2948_; 
wire u5__abc_81276_new_n2949_; 
wire u5__abc_81276_new_n2950_; 
wire u5__abc_81276_new_n2951_; 
wire u5__abc_81276_new_n2952_; 
wire u5__abc_81276_new_n2953_; 
wire u5__abc_81276_new_n2953__bF_buf0; 
wire u5__abc_81276_new_n2953__bF_buf1; 
wire u5__abc_81276_new_n2953__bF_buf2; 
wire u5__abc_81276_new_n2953__bF_buf3; 
wire u5__abc_81276_new_n2954_; 
wire u5__abc_81276_new_n2955_; 
wire u5__abc_81276_new_n2956_; 
wire u5__abc_81276_new_n2957_; 
wire u5__abc_81276_new_n2958_; 
wire u5__abc_81276_new_n2959_; 
wire u5__abc_81276_new_n2960_; 
wire u5__abc_81276_new_n2961_; 
wire u5__abc_81276_new_n2962_; 
wire u5__abc_81276_new_n2963_; 
wire u5__abc_81276_new_n2964_; 
wire u5__abc_81276_new_n2965_; 
wire u5__abc_81276_new_n2966_; 
wire u5__abc_81276_new_n2967_; 
wire u5__abc_81276_new_n2968_; 
wire u5__abc_81276_new_n2969_; 
wire u5__abc_81276_new_n2970_; 
wire u5__abc_81276_new_n2971_; 
wire u5__abc_81276_new_n2972_; 
wire u5__abc_81276_new_n2973_; 
wire u5__abc_81276_new_n2975_; 
wire u5__abc_81276_new_n2976_; 
wire u5__abc_81276_new_n2977_; 
wire u5__abc_81276_new_n2978_; 
wire u5__abc_81276_new_n2979_; 
wire u5__abc_81276_new_n2980_; 
wire u5__abc_81276_new_n2981_; 
wire u5__abc_81276_new_n2982_; 
wire u5__abc_81276_new_n2983_; 
wire u5__abc_81276_new_n2984_; 
wire u5__abc_81276_new_n2985_; 
wire u5__abc_81276_new_n2986_; 
wire u5__abc_81276_new_n2987_; 
wire u5__abc_81276_new_n2988_; 
wire u5__abc_81276_new_n2989_; 
wire u5__abc_81276_new_n2990_; 
wire u5__abc_81276_new_n2991_; 
wire u5__abc_81276_new_n2992_; 
wire u5__abc_81276_new_n2993_; 
wire u5__abc_81276_new_n2994_; 
wire u5__abc_81276_new_n2995_; 
wire u5__abc_81276_new_n2996_; 
wire u5__abc_81276_new_n2997_; 
wire u5__abc_81276_new_n2998_; 
wire u5__abc_81276_new_n2999_; 
wire u5__abc_81276_new_n3000_; 
wire u5__abc_81276_new_n3001_; 
wire u5__abc_81276_new_n3002_; 
wire u5__abc_81276_new_n3003_; 
wire u5__abc_81276_new_n3004_; 
wire u5__abc_81276_new_n3005_; 
wire u5__abc_81276_new_n3006_; 
wire u5__abc_81276_new_n3007_; 
wire u5__abc_81276_new_n3008_; 
wire u5__abc_81276_new_n3009_; 
wire u5__abc_81276_new_n3010_; 
wire u5__abc_81276_new_n3011_; 
wire u5__abc_81276_new_n3012_; 
wire u5__abc_81276_new_n3013_; 
wire u5__abc_81276_new_n3014_; 
wire u5__abc_81276_new_n3015_; 
wire u5__abc_81276_new_n3016_; 
wire u5__abc_81276_new_n3017_; 
wire u5__abc_81276_new_n3018_; 
wire u5__abc_81276_new_n3019_; 
wire u5__abc_81276_new_n3020_; 
wire u5__abc_81276_new_n3021_; 
wire u5__abc_81276_new_n3022_; 
wire u5__abc_81276_new_n3023_; 
wire u5__abc_81276_new_n3024_; 
wire u5__abc_81276_new_n3025_; 
wire u5__abc_81276_new_n3026_; 
wire u5__abc_81276_new_n3027_; 
wire u5__abc_81276_new_n3028_; 
wire u5__abc_81276_new_n3029_; 
wire u5__abc_81276_new_n3030_; 
wire u5__abc_81276_new_n3031_; 
wire u5__abc_81276_new_n3032_; 
wire u5__abc_81276_new_n3034_; 
wire u5__abc_81276_new_n3035_; 
wire u5__abc_81276_new_n3036_; 
wire u5__abc_81276_new_n3037_; 
wire u5__abc_81276_new_n3038_; 
wire u5__abc_81276_new_n3039_; 
wire u5__abc_81276_new_n3040_; 
wire u5__abc_81276_new_n3041_; 
wire u5__abc_81276_new_n3042_; 
wire u5__abc_81276_new_n3043_; 
wire u5__abc_81276_new_n3044_; 
wire u5__abc_81276_new_n3045_; 
wire u5__abc_81276_new_n3046_; 
wire u5__abc_81276_new_n3047_; 
wire u5__abc_81276_new_n3048_; 
wire u5__abc_81276_new_n3049_; 
wire u5__abc_81276_new_n3050_; 
wire u5__abc_81276_new_n3051_; 
wire u5__abc_81276_new_n3052_; 
wire u5__abc_81276_new_n3053_; 
wire u5__abc_81276_new_n3054_; 
wire u5__abc_81276_new_n3055_; 
wire u5__abc_81276_new_n3056_; 
wire u5__abc_81276_new_n3058_; 
wire u5__abc_81276_new_n3059_; 
wire u5__abc_81276_new_n3060_; 
wire u5__abc_81276_new_n3061_; 
wire u5__abc_81276_new_n3062_; 
wire u5__abc_81276_new_n3063_; 
wire u5__abc_81276_new_n3064_; 
wire u5__abc_81276_new_n3065_; 
wire u5__abc_81276_new_n3066_; 
wire u5__abc_81276_new_n3067_; 
wire u5__abc_81276_new_n3068_; 
wire u5__abc_81276_new_n3069_; 
wire u5__abc_81276_new_n3070_; 
wire u5__abc_81276_new_n3071_; 
wire u5__abc_81276_new_n3072_; 
wire u5__abc_81276_new_n3073_; 
wire u5__abc_81276_new_n3074_; 
wire u5__abc_81276_new_n3075_; 
wire u5__abc_81276_new_n3076_; 
wire u5__abc_81276_new_n3077_; 
wire u5__abc_81276_new_n3078_; 
wire u5__abc_81276_new_n3080_; 
wire u5__abc_81276_new_n3081_; 
wire u5__abc_81276_new_n3082_; 
wire u5__abc_81276_new_n3083_; 
wire u5__abc_81276_new_n3084_; 
wire u5__abc_81276_new_n3085_; 
wire u5__abc_81276_new_n3086_; 
wire u5__abc_81276_new_n3087_; 
wire u5__abc_81276_new_n3088_; 
wire u5__abc_81276_new_n3089_; 
wire u5__abc_81276_new_n3090_; 
wire u5__abc_81276_new_n3091_; 
wire u5__abc_81276_new_n3092_; 
wire u5__abc_81276_new_n3093_; 
wire u5__abc_81276_new_n3094_; 
wire u5__abc_81276_new_n3095_; 
wire u5__abc_81276_new_n3096_; 
wire u5__abc_81276_new_n3097_; 
wire u5__abc_81276_new_n3099_; 
wire u5__abc_81276_new_n3100_; 
wire u5__abc_81276_new_n3101_; 
wire u5__abc_81276_new_n3102_; 
wire u5__abc_81276_new_n3103_; 
wire u5__abc_81276_new_n3104_; 
wire u5__abc_81276_new_n3105_; 
wire u5__abc_81276_new_n3106_; 
wire u5__abc_81276_new_n3107_; 
wire u5__abc_81276_new_n3108_; 
wire u5__abc_81276_new_n3109_; 
wire u5__abc_81276_new_n3110_; 
wire u5__abc_81276_new_n3111_; 
wire u5__abc_81276_new_n3112_; 
wire u5__abc_81276_new_n3113_; 
wire u5__abc_81276_new_n3115_; 
wire u5__abc_81276_new_n3116_; 
wire u5__abc_81276_new_n3117_; 
wire u5__abc_81276_new_n3118_; 
wire u5__abc_81276_new_n3119_; 
wire u5__abc_81276_new_n3120_; 
wire u5__abc_81276_new_n3121_; 
wire u5__abc_81276_new_n3122_; 
wire u5__abc_81276_new_n3123_; 
wire u5__abc_81276_new_n3124_; 
wire u5__abc_81276_new_n3126_; 
wire u5__abc_81276_new_n3127_; 
wire u5__abc_81276_new_n3128_; 
wire u5__abc_81276_new_n3129_; 
wire u5__abc_81276_new_n3130_; 
wire u5__abc_81276_new_n3131_; 
wire u5__abc_81276_new_n3132_; 
wire u5__abc_81276_new_n3133_; 
wire u5__abc_81276_new_n3134_; 
wire u5__abc_81276_new_n3136_; 
wire u5__abc_81276_new_n3137_; 
wire u5__abc_81276_new_n3138_; 
wire u5__abc_81276_new_n3139_; 
wire u5__abc_81276_new_n3140_; 
wire u5__abc_81276_new_n3141_; 
wire u5__abc_81276_new_n3143_; 
wire u5__abc_81276_new_n3144_; 
wire u5__abc_81276_new_n3145_; 
wire u5__abc_81276_new_n3146_; 
wire u5__abc_81276_new_n3147_; 
wire u5__abc_81276_new_n3148_; 
wire u5__abc_81276_new_n3149_; 
wire u5__abc_81276_new_n3150_; 
wire u5__abc_81276_new_n3151_; 
wire u5__abc_81276_new_n3152_; 
wire u5__abc_81276_new_n3154_; 
wire u5__abc_81276_new_n3155_; 
wire u5__abc_81276_new_n3156_; 
wire u5__abc_81276_new_n3157_; 
wire u5__abc_81276_new_n3158_; 
wire u5__abc_81276_new_n3159_; 
wire u5__abc_81276_new_n3160_; 
wire u5__abc_81276_new_n3161_; 
wire u5__abc_81276_new_n3162_; 
wire u5__abc_81276_new_n3164_; 
wire u5__abc_81276_new_n3165_; 
wire u5__abc_81276_new_n3166_; 
wire u5__abc_81276_new_n3167_; 
wire u5__abc_81276_new_n3168_; 
wire u5__abc_81276_new_n3169_; 
wire u5__abc_81276_new_n3170_; 
wire u5__abc_81276_new_n3172_; 
wire u5__abc_81276_new_n3173_; 
wire u5__abc_81276_new_n3174_; 
wire u5__abc_81276_new_n3175_; 
wire u5__abc_81276_new_n3176_; 
wire u5__abc_81276_new_n3177_; 
wire u5__abc_81276_new_n3178_; 
wire u5__abc_81276_new_n3179_; 
wire u5__abc_81276_new_n3180_; 
wire u5__abc_81276_new_n3181_; 
wire u5__abc_81276_new_n3182_; 
wire u5__abc_81276_new_n3183_; 
wire u5__abc_81276_new_n3185_; 
wire u5__abc_81276_new_n3186_; 
wire u5__abc_81276_new_n3188_; 
wire u5__abc_81276_new_n3189_; 
wire u5__abc_81276_new_n3191_; 
wire u5__abc_81276_new_n3192_; 
wire u5__abc_81276_new_n3194_; 
wire u5__abc_81276_new_n3195_; 
wire u5__abc_81276_new_n3196_; 
wire u5__abc_81276_new_n3197_; 
wire u5__abc_81276_new_n3198_; 
wire u5__abc_81276_new_n3199_; 
wire u5__abc_81276_new_n3200_; 
wire u5__abc_81276_new_n3201_; 
wire u5__abc_81276_new_n3203_; 
wire u5__abc_81276_new_n3204_; 
wire u5__abc_81276_new_n3206_; 
wire u5__abc_81276_new_n3207_; 
wire u5__abc_81276_new_n3208_; 
wire u5__abc_81276_new_n3209_; 
wire u5__abc_81276_new_n3210_; 
wire u5__abc_81276_new_n3211_; 
wire u5__abc_81276_new_n3212_; 
wire u5__abc_81276_new_n3213_; 
wire u5__abc_81276_new_n3214_; 
wire u5__abc_81276_new_n3215_; 
wire u5__abc_81276_new_n3215__bF_buf0; 
wire u5__abc_81276_new_n3215__bF_buf1; 
wire u5__abc_81276_new_n3215__bF_buf2; 
wire u5__abc_81276_new_n3215__bF_buf3; 
wire u5__abc_81276_new_n3215__bF_buf4; 
wire u5__abc_81276_new_n3216_; 
wire u5__abc_81276_new_n3218_; 
wire u5__abc_81276_new_n3219_; 
wire u5__abc_81276_new_n3220_; 
wire u5__abc_81276_new_n3221_; 
wire u5__abc_81276_new_n3222_; 
wire u5__abc_81276_new_n3223_; 
wire u5__abc_81276_new_n3224_; 
wire u5__abc_81276_new_n3225_; 
wire u5__abc_81276_new_n3226_; 
wire u5__abc_81276_new_n3227_; 
wire u5__abc_81276_new_n3228_; 
wire u5__abc_81276_new_n3229_; 
wire u5__abc_81276_new_n3230_; 
wire u5__abc_81276_new_n3231_; 
wire u5__abc_81276_new_n3232_; 
wire u5__abc_81276_new_n3233_; 
wire u5__abc_81276_new_n3234_; 
wire u5__abc_81276_new_n3235_; 
wire u5__abc_81276_new_n3236_; 
wire u5__abc_81276_new_n3238_; 
wire u5__abc_81276_new_n3239_; 
wire u5__abc_81276_new_n3240_; 
wire u5__abc_81276_new_n3241_; 
wire u5__abc_81276_new_n3242_; 
wire u5__abc_81276_new_n3243_; 
wire u5__abc_81276_new_n3244_; 
wire u5__abc_81276_new_n3245_; 
wire u5__abc_81276_new_n3246_; 
wire u5__abc_81276_new_n3247_; 
wire u5__abc_81276_new_n3248_; 
wire u5__abc_81276_new_n3249_; 
wire u5__abc_81276_new_n3250_; 
wire u5__abc_81276_new_n3251_; 
wire u5__abc_81276_new_n3252_; 
wire u5__abc_81276_new_n3253_; 
wire u5__abc_81276_new_n3254_; 
wire u5__abc_81276_new_n3255_; 
wire u5__abc_81276_new_n3256_; 
wire u5__abc_81276_new_n3257_; 
wire u5__abc_81276_new_n3258_; 
wire u5__abc_81276_new_n3259_; 
wire u5__abc_81276_new_n3260_; 
wire u5__abc_81276_new_n3261_; 
wire u5__abc_81276_new_n3262_; 
wire u5__abc_81276_new_n3263_; 
wire u5__abc_81276_new_n3264_; 
wire u5__abc_81276_new_n3265_; 
wire u5__abc_81276_new_n3266_; 
wire u5__abc_81276_new_n3267_; 
wire u5__abc_81276_new_n3268_; 
wire u5__abc_81276_new_n3269_; 
wire u5__abc_81276_new_n3270_; 
wire u5__abc_81276_new_n3271_; 
wire u5__abc_81276_new_n3272_; 
wire u5__abc_81276_new_n3273_; 
wire u5__abc_81276_new_n3274_; 
wire u5__abc_81276_new_n3275_; 
wire u5__abc_81276_new_n3276_; 
wire u5__abc_81276_new_n3277_; 
wire u5__abc_81276_new_n3278_; 
wire u5__abc_81276_new_n3279_; 
wire u5__abc_81276_new_n3280_; 
wire u5__abc_81276_new_n3281_; 
wire u5__abc_81276_new_n3282_; 
wire u5__abc_81276_new_n3283_; 
wire u5__abc_81276_new_n3284_; 
wire u5__abc_81276_new_n3285_; 
wire u5__abc_81276_new_n3286_; 
wire u5__abc_81276_new_n3287_; 
wire u5__abc_81276_new_n3288_; 
wire u5__abc_81276_new_n3289_; 
wire u5__abc_81276_new_n3290_; 
wire u5__abc_81276_new_n3292_; 
wire u5__abc_81276_new_n3293_; 
wire u5__abc_81276_new_n3294_; 
wire u5__abc_81276_new_n3295_; 
wire u5__abc_81276_new_n3296_; 
wire u5__abc_81276_new_n3297_; 
wire u5__abc_81276_new_n3299_; 
wire u5__abc_81276_new_n3300_; 
wire u5__abc_81276_new_n3301_; 
wire u5__abc_81276_new_n3302_; 
wire u5__abc_81276_new_n3303_; 
wire u5__abc_81276_new_n3304_; 
wire u5__abc_81276_new_n3305_; 
wire u5__abc_81276_new_n3306_; 
wire u5__abc_81276_new_n3307_; 
wire u5__abc_81276_new_n3308_; 
wire u5__abc_81276_new_n3309_; 
wire u5__abc_81276_new_n3310_; 
wire u5__abc_81276_new_n3311_; 
wire u5__abc_81276_new_n3312_; 
wire u5__abc_81276_new_n3313_; 
wire u5__abc_81276_new_n3314_; 
wire u5__abc_81276_new_n3315_; 
wire u5__abc_81276_new_n3317_; 
wire u5__abc_81276_new_n3318_; 
wire u5__abc_81276_new_n3319_; 
wire u5__abc_81276_new_n3320_; 
wire u5__abc_81276_new_n3321_; 
wire u5__abc_81276_new_n3323_; 
wire u5__abc_81276_new_n3323__bF_buf0; 
wire u5__abc_81276_new_n3323__bF_buf1; 
wire u5__abc_81276_new_n3323__bF_buf2; 
wire u5__abc_81276_new_n3323__bF_buf3; 
wire u5__abc_81276_new_n3324_; 
wire u5__abc_81276_new_n3325_; 
wire u5__abc_81276_new_n3326_; 
wire u5__abc_81276_new_n3327_; 
wire u5__abc_81276_new_n3328_; 
wire u5__abc_81276_new_n3329_; 
wire u5__abc_81276_new_n3330_; 
wire u5__abc_81276_new_n3331_; 
wire u5__abc_81276_new_n3332_; 
wire u5__abc_81276_new_n3333_; 
wire u5__abc_81276_new_n3334_; 
wire u5__abc_81276_new_n3335_; 
wire u5__abc_81276_new_n3336_; 
wire u5__abc_81276_new_n3337_; 
wire u5__abc_81276_new_n3338_; 
wire u5__abc_81276_new_n3339_; 
wire u5__abc_81276_new_n3340_; 
wire u5__abc_81276_new_n3341_; 
wire u5__abc_81276_new_n3342_; 
wire u5__abc_81276_new_n3343_; 
wire u5__abc_81276_new_n3344_; 
wire u5__abc_81276_new_n3346_; 
wire u5__abc_81276_new_n3347_; 
wire u5__abc_81276_new_n3348_; 
wire u5__abc_81276_new_n3349_; 
wire u5__abc_81276_new_n3350_; 
wire u5__abc_81276_new_n3351_; 
wire u5__abc_81276_new_n3352_; 
wire u5__abc_81276_new_n3353_; 
wire u5__abc_81276_new_n3354_; 
wire u5__abc_81276_new_n3355_; 
wire u5__abc_81276_new_n3356_; 
wire u5__abc_81276_new_n3357_; 
wire u5__abc_81276_new_n3358_; 
wire u5__abc_81276_new_n3359_; 
wire u5__abc_81276_new_n3361_; 
wire u5__abc_81276_new_n3362_; 
wire u5__abc_81276_new_n3363_; 
wire u5__abc_81276_new_n3364_; 
wire u5__abc_81276_new_n3365_; 
wire u5__abc_81276_new_n3366_; 
wire u5__abc_81276_new_n3367_; 
wire u5__abc_81276_new_n3368_; 
wire u5__abc_81276_new_n3369_; 
wire u5__abc_81276_new_n3370_; 
wire u5__abc_81276_new_n3371_; 
wire u5__abc_81276_new_n3372_; 
wire u5__abc_81276_new_n3373_; 
wire u5__abc_81276_new_n3374_; 
wire u5__abc_81276_new_n3375_; 
wire u5__abc_81276_new_n3376_; 
wire u5__abc_81276_new_n3377_; 
wire u5__abc_81276_new_n3378_; 
wire u5__abc_81276_new_n3379_; 
wire u5__abc_81276_new_n3381_; 
wire u5__abc_81276_new_n3382_; 
wire u5__abc_81276_new_n3383_; 
wire u5__abc_81276_new_n3384_; 
wire u5__abc_81276_new_n3385_; 
wire u5__abc_81276_new_n3386_; 
wire u5__abc_81276_new_n3387_; 
wire u5__abc_81276_new_n3388_; 
wire u5__abc_81276_new_n3389_; 
wire u5__abc_81276_new_n3390_; 
wire u5__abc_81276_new_n3391_; 
wire u5__abc_81276_new_n3392_; 
wire u5__abc_81276_new_n3393_; 
wire u5__abc_81276_new_n3394_; 
wire u5__abc_81276_new_n3395_; 
wire u5__abc_81276_new_n3396_; 
wire u5__abc_81276_new_n3397_; 
wire u5__abc_81276_new_n3398_; 
wire u5__abc_81276_new_n3399_; 
wire u5__abc_81276_new_n3400_; 
wire u5__abc_81276_new_n3402_; 
wire u5__abc_81276_new_n3403_; 
wire u5__abc_81276_new_n3404_; 
wire u5__abc_81276_new_n3405_; 
wire u5__abc_81276_new_n3406_; 
wire u5__abc_81276_new_n3408_; 
wire u5__abc_81276_new_n3409_; 
wire u5__abc_81276_new_n3410_; 
wire u5__abc_81276_new_n3411_; 
wire u5__abc_81276_new_n3412_; 
wire u5__abc_81276_new_n3413_; 
wire u5__abc_81276_new_n3414_; 
wire u5__abc_81276_new_n3415_; 
wire u5__abc_81276_new_n3416_; 
wire u5__abc_81276_new_n3417_; 
wire u5__abc_81276_new_n3418_; 
wire u5__abc_81276_new_n3419_; 
wire u5__abc_81276_new_n3421_; 
wire u5__abc_81276_new_n3422_; 
wire u5__abc_81276_new_n3423_; 
wire u5__abc_81276_new_n3424_; 
wire u5__abc_81276_new_n3425_; 
wire u5__abc_81276_new_n3426_; 
wire u5__abc_81276_new_n3427_; 
wire u5__abc_81276_new_n3428_; 
wire u5__abc_81276_new_n3430_; 
wire u5__abc_81276_new_n3431_; 
wire u5__abc_81276_new_n3432_; 
wire u5__abc_81276_new_n3433_; 
wire u5__abc_81276_new_n3434_; 
wire u5__abc_81276_new_n3435_; 
wire u5__abc_81276_new_n3437_; 
wire u5__abc_81276_new_n3438_; 
wire u5__abc_81276_new_n3439_; 
wire u5__abc_81276_new_n3440_; 
wire u5__abc_81276_new_n3441_; 
wire u5__abc_81276_new_n3442_; 
wire u5__abc_81276_new_n3443_; 
wire u5__abc_81276_new_n3444_; 
wire u5__abc_81276_new_n3445_; 
wire u5__abc_81276_new_n3446_; 
wire u5__abc_81276_new_n3447_; 
wire u5__abc_81276_new_n3448_; 
wire u5__abc_81276_new_n3449_; 
wire u5__abc_81276_new_n3450_; 
wire u5__abc_81276_new_n3451_; 
wire u5__abc_81276_new_n3452_; 
wire u5__abc_81276_new_n3454_; 
wire u5__abc_81276_new_n3455_; 
wire u5__abc_81276_new_n3456_; 
wire u5__abc_81276_new_n3457_; 
wire u5__abc_81276_new_n3458_; 
wire u5__abc_81276_new_n3459_; 
wire u5__abc_81276_new_n3460_; 
wire u5__abc_81276_new_n3461_; 
wire u5__abc_81276_new_n3462_; 
wire u5__abc_81276_new_n3463_; 
wire u5__abc_81276_new_n3464_; 
wire u5__abc_81276_new_n3465_; 
wire u5__abc_81276_new_n3466_; 
wire u5__abc_81276_new_n3467_; 
wire u5__abc_81276_new_n3468_; 
wire u5__abc_81276_new_n3469_; 
wire u5__abc_81276_new_n3470_; 
wire u5__abc_81276_new_n3471_; 
wire u5__abc_81276_new_n3472_; 
wire u5__abc_81276_new_n3473_; 
wire u5__abc_81276_new_n3474_; 
wire u5__abc_81276_new_n3475_; 
wire u5__abc_81276_new_n3476_; 
wire u5__abc_81276_new_n3478_; 
wire u5__abc_81276_new_n3479_; 
wire u5__abc_81276_new_n3480_; 
wire u5__abc_81276_new_n3481_; 
wire u5__abc_81276_new_n3482_; 
wire u5__abc_81276_new_n3483_; 
wire u5__abc_81276_new_n3484_; 
wire u5__abc_81276_new_n3485_; 
wire u5__abc_81276_new_n3486_; 
wire u5__abc_81276_new_n3487_; 
wire u5__abc_81276_new_n3488_; 
wire u5__abc_81276_new_n3489_; 
wire u5__abc_81276_new_n3490_; 
wire u5__abc_81276_new_n3491_; 
wire u5__abc_81276_new_n3492_; 
wire u5__abc_81276_new_n3493_; 
wire u5__abc_81276_new_n3494_; 
wire u5__abc_81276_new_n3495_; 
wire u5__abc_81276_new_n3496_; 
wire u5__abc_81276_new_n3497_; 
wire u5__abc_81276_new_n3498_; 
wire u5__abc_81276_new_n3499_; 
wire u5__abc_81276_new_n3500_; 
wire u5__abc_81276_new_n3501_; 
wire u5__abc_81276_new_n3502_; 
wire u5__abc_81276_new_n3504_; 
wire u5__abc_81276_new_n3505_; 
wire u5__abc_81276_new_n3506_; 
wire u5__abc_81276_new_n3507_; 
wire u5__abc_81276_new_n3508_; 
wire u5__abc_81276_new_n3509_; 
wire u5__abc_81276_new_n3510_; 
wire u5__abc_81276_new_n3511_; 
wire u5__abc_81276_new_n3512_; 
wire u5__abc_81276_new_n3513_; 
wire u5__abc_81276_new_n3514_; 
wire u5__abc_81276_new_n3515_; 
wire u5__abc_81276_new_n3516_; 
wire u5__abc_81276_new_n3517_; 
wire u5__abc_81276_new_n3518_; 
wire u5__abc_81276_new_n3520_; 
wire u5__abc_81276_new_n3521_; 
wire u5__abc_81276_new_n3522_; 
wire u5__abc_81276_new_n3523_; 
wire u5__abc_81276_new_n3524_; 
wire u5__abc_81276_new_n3526_; 
wire u5__abc_81276_new_n3527_; 
wire u5__abc_81276_new_n3528_; 
wire u5__abc_81276_new_n3529_; 
wire u5__abc_81276_new_n3530_; 
wire u5__abc_81276_new_n3531_; 
wire u5__abc_81276_new_n3532_; 
wire u5__abc_81276_new_n3533_; 
wire u5__abc_81276_new_n3535_; 
wire u5__abc_81276_new_n3536_; 
wire u5__abc_81276_new_n3537_; 
wire u5__abc_81276_new_n3538_; 
wire u5__abc_81276_new_n3539_; 
wire u5__abc_81276_new_n3540_; 
wire u5__abc_81276_new_n3541_; 
wire u5__abc_81276_new_n3542_; 
wire u5__abc_81276_new_n3543_; 
wire u5__abc_81276_new_n3545_; 
wire u5__abc_81276_new_n3546_; 
wire u5__abc_81276_new_n3548_; 
wire u5__abc_81276_new_n3549_; 
wire u5__abc_81276_new_n3550_; 
wire u5__abc_81276_new_n3551_; 
wire u5__abc_81276_new_n3552_; 
wire u5__abc_81276_new_n3553_; 
wire u5__abc_81276_new_n3555_; 
wire u5__abc_81276_new_n3556_; 
wire u5__abc_81276_new_n3557_; 
wire u5__abc_81276_new_n3558_; 
wire u5__abc_81276_new_n3559_; 
wire u5__abc_81276_new_n3560_; 
wire u5__abc_81276_new_n3561_; 
wire u5__abc_81276_new_n3563_; 
wire u5__abc_81276_new_n3564_; 
wire u5__abc_81276_new_n3565_; 
wire u5__abc_81276_new_n3566_; 
wire u5__abc_81276_new_n3567_; 
wire u5__abc_81276_new_n3568_; 
wire u5__abc_81276_new_n3569_; 
wire u5__abc_81276_new_n3570_; 
wire u5__abc_81276_new_n3571_; 
wire u5__abc_81276_new_n3572_; 
wire u5__abc_81276_new_n3573_; 
wire u5__abc_81276_new_n3575_; 
wire u5__abc_81276_new_n3576_; 
wire u5__abc_81276_new_n3577_; 
wire u5__abc_81276_new_n3578_; 
wire u5__abc_81276_new_n3579_; 
wire u5__abc_81276_new_n3580_; 
wire u5__abc_81276_new_n3581_; 
wire u5__abc_81276_new_n3583_; 
wire u5__abc_81276_new_n3584_; 
wire u5__abc_81276_new_n3585_; 
wire u5__abc_81276_new_n3586_; 
wire u5__abc_81276_new_n3587_; 
wire u5__abc_81276_new_n3588_; 
wire u5__abc_81276_new_n3589_; 
wire u5__abc_81276_new_n3590_; 
wire u5__abc_81276_new_n3592_; 
wire u5__abc_81276_new_n3593_; 
wire u5__abc_81276_new_n3594_; 
wire u5__abc_81276_new_n3595_; 
wire u5__abc_81276_new_n3596_; 
wire u5__abc_81276_new_n3598_; 
wire u5__abc_81276_new_n3599_; 
wire u5__abc_81276_new_n3600_; 
wire u5__abc_81276_new_n3601_; 
wire u5__abc_81276_new_n3602_; 
wire u5__abc_81276_new_n3604_; 
wire u5__abc_81276_new_n3605_; 
wire u5__abc_81276_new_n3606_; 
wire u5__abc_81276_new_n3607_; 
wire u5__abc_81276_new_n3608_; 
wire u5__abc_81276_new_n3609_; 
wire u5__abc_81276_new_n3610_; 
wire u5__abc_81276_new_n3612_; 
wire u5__abc_81276_new_n3613_; 
wire u5__abc_81276_new_n3614_; 
wire u5__abc_81276_new_n3615_; 
wire u5__abc_81276_new_n3616_; 
wire u5__abc_81276_new_n3617_; 
wire u5__abc_81276_new_n3618_; 
wire u5__abc_81276_new_n3619_; 
wire u5__abc_81276_new_n3621_; 
wire u5__abc_81276_new_n3622_; 
wire u5__abc_81276_new_n3623_; 
wire u5__abc_81276_new_n3624_; 
wire u5__abc_81276_new_n3626_; 
wire u5__abc_81276_new_n3627_; 
wire u5__abc_81276_new_n3628_; 
wire u5__abc_81276_new_n3629_; 
wire u5__abc_81276_new_n3630_; 
wire u5__abc_81276_new_n3632_; 
wire u5__abc_81276_new_n3633_; 
wire u5__abc_81276_new_n3634_; 
wire u5__abc_81276_new_n3636_; 
wire u5__abc_81276_new_n3638_; 
wire u5__abc_81276_new_n3639_; 
wire u5__abc_81276_new_n3640_; 
wire u5__abc_81276_new_n3642_; 
wire u5__abc_81276_new_n3643_; 
wire u5__abc_81276_new_n3644_; 
wire u5__abc_81276_new_n3645_; 
wire u5__abc_81276_new_n3646_; 
wire u5__abc_81276_new_n3647_; 
wire u5__abc_81276_new_n3648_; 
wire u5__abc_81276_new_n3649_; 
wire u5__abc_81276_new_n3650_; 
wire u5__abc_81276_new_n3652_; 
wire u5__abc_81276_new_n3653_; 
wire u5__abc_81276_new_n3654_; 
wire u5__abc_81276_new_n3655_; 
wire u5__abc_81276_new_n3656_; 
wire u5__abc_81276_new_n3658_; 
wire u5__abc_81276_new_n3659_; 
wire u5__abc_81276_new_n3660_; 
wire u5__abc_81276_new_n3661_; 
wire u5__abc_81276_new_n3662_; 
wire u5__abc_81276_new_n3663_; 
wire u5__abc_81276_new_n3664_; 
wire u5__abc_81276_new_n3666_; 
wire u5__abc_81276_new_n3667_; 
wire u5__abc_81276_new_n3668_; 
wire u5__abc_81276_new_n3669_; 
wire u5__abc_81276_new_n366_; 
wire u5__abc_81276_new_n3671_; 
wire u5__abc_81276_new_n3673_; 
wire u5__abc_81276_new_n3674_; 
wire u5__abc_81276_new_n3675_; 
wire u5__abc_81276_new_n3676_; 
wire u5__abc_81276_new_n3677_; 
wire u5__abc_81276_new_n3679_; 
wire u5__abc_81276_new_n367_; 
wire u5__abc_81276_new_n3680_; 
wire u5__abc_81276_new_n3681_; 
wire u5__abc_81276_new_n3682_; 
wire u5__abc_81276_new_n3684_; 
wire u5__abc_81276_new_n3685_; 
wire u5__abc_81276_new_n3686_; 
wire u5__abc_81276_new_n3688_; 
wire u5__abc_81276_new_n3689_; 
wire u5__abc_81276_new_n368_; 
wire u5__abc_81276_new_n3690_; 
wire u5__abc_81276_new_n3691_; 
wire u5__abc_81276_new_n3693_; 
wire u5__abc_81276_new_n3694_; 
wire u5__abc_81276_new_n3695_; 
wire u5__abc_81276_new_n3696_; 
wire u5__abc_81276_new_n3697_; 
wire u5__abc_81276_new_n3698_; 
wire u5__abc_81276_new_n3699_; 
wire u5__abc_81276_new_n369_; 
wire u5__abc_81276_new_n3701_; 
wire u5__abc_81276_new_n3702_; 
wire u5__abc_81276_new_n3703_; 
wire u5__abc_81276_new_n3704_; 
wire u5__abc_81276_new_n3706_; 
wire u5__abc_81276_new_n3707_; 
wire u5__abc_81276_new_n3708_; 
wire u5__abc_81276_new_n3709_; 
wire u5__abc_81276_new_n370_; 
wire u5__abc_81276_new_n3711_; 
wire u5__abc_81276_new_n3712_; 
wire u5__abc_81276_new_n3713_; 
wire u5__abc_81276_new_n3714_; 
wire u5__abc_81276_new_n3716_; 
wire u5__abc_81276_new_n3717_; 
wire u5__abc_81276_new_n3718_; 
wire u5__abc_81276_new_n371_; 
wire u5__abc_81276_new_n3720_; 
wire u5__abc_81276_new_n3721_; 
wire u5__abc_81276_new_n3723_; 
wire u5__abc_81276_new_n3724_; 
wire u5__abc_81276_new_n3725_; 
wire u5__abc_81276_new_n3727_; 
wire u5__abc_81276_new_n3728_; 
wire u5__abc_81276_new_n3729_; 
wire u5__abc_81276_new_n372_; 
wire u5__abc_81276_new_n3730_; 
wire u5__abc_81276_new_n3731_; 
wire u5__abc_81276_new_n3732_; 
wire u5__abc_81276_new_n3733_; 
wire u5__abc_81276_new_n3734_; 
wire u5__abc_81276_new_n3735_; 
wire u5__abc_81276_new_n3736_; 
wire u5__abc_81276_new_n3737_; 
wire u5__abc_81276_new_n3739_; 
wire u5__abc_81276_new_n373_; 
wire u5__abc_81276_new_n3740_; 
wire u5__abc_81276_new_n3741_; 
wire u5__abc_81276_new_n3742_; 
wire u5__abc_81276_new_n3743_; 
wire u5__abc_81276_new_n3745_; 
wire u5__abc_81276_new_n3746_; 
wire u5__abc_81276_new_n3747_; 
wire u5__abc_81276_new_n3748_; 
wire u5__abc_81276_new_n3749_; 
wire u5__abc_81276_new_n374_; 
wire u5__abc_81276_new_n3750_; 
wire u5__abc_81276_new_n3752_; 
wire u5__abc_81276_new_n3753_; 
wire u5__abc_81276_new_n3754_; 
wire u5__abc_81276_new_n3755_; 
wire u5__abc_81276_new_n3756_; 
wire u5__abc_81276_new_n3757_; 
wire u5__abc_81276_new_n3758_; 
wire u5__abc_81276_new_n3759_; 
wire u5__abc_81276_new_n375_; 
wire u5__abc_81276_new_n3760_; 
wire u5__abc_81276_new_n3761_; 
wire u5__abc_81276_new_n3762_; 
wire u5__abc_81276_new_n3763_; 
wire u5__abc_81276_new_n3765_; 
wire u5__abc_81276_new_n3766_; 
wire u5__abc_81276_new_n3767_; 
wire u5__abc_81276_new_n3768_; 
wire u5__abc_81276_new_n3769_; 
wire u5__abc_81276_new_n376_; 
wire u5__abc_81276_new_n3770_; 
wire u5__abc_81276_new_n3771_; 
wire u5__abc_81276_new_n3772_; 
wire u5__abc_81276_new_n3773_; 
wire u5__abc_81276_new_n3774_; 
wire u5__abc_81276_new_n3776_; 
wire u5__abc_81276_new_n3777_; 
wire u5__abc_81276_new_n3778_; 
wire u5__abc_81276_new_n3779_; 
wire u5__abc_81276_new_n377_; 
wire u5__abc_81276_new_n3780_; 
wire u5__abc_81276_new_n3781_; 
wire u5__abc_81276_new_n3782_; 
wire u5__abc_81276_new_n3783_; 
wire u5__abc_81276_new_n3784_; 
wire u5__abc_81276_new_n3785_; 
wire u5__abc_81276_new_n3786_; 
wire u5__abc_81276_new_n3788_; 
wire u5__abc_81276_new_n3789_; 
wire u5__abc_81276_new_n378_; 
wire u5__abc_81276_new_n3790_; 
wire u5__abc_81276_new_n3791_; 
wire u5__abc_81276_new_n3792_; 
wire u5__abc_81276_new_n3793_; 
wire u5__abc_81276_new_n3794_; 
wire u5__abc_81276_new_n3795_; 
wire u5__abc_81276_new_n3797_; 
wire u5__abc_81276_new_n3798_; 
wire u5__abc_81276_new_n3799_; 
wire u5__abc_81276_new_n379_; 
wire u5__abc_81276_new_n3800_; 
wire u5__abc_81276_new_n3801_; 
wire u5__abc_81276_new_n3802_; 
wire u5__abc_81276_new_n3804_; 
wire u5__abc_81276_new_n3805_; 
wire u5__abc_81276_new_n3806_; 
wire u5__abc_81276_new_n3807_; 
wire u5__abc_81276_new_n3808_; 
wire u5__abc_81276_new_n3809_; 
wire u5__abc_81276_new_n380_; 
wire u5__abc_81276_new_n3810_; 
wire u5__abc_81276_new_n3811_; 
wire u5__abc_81276_new_n3812_; 
wire u5__abc_81276_new_n3814_; 
wire u5__abc_81276_new_n3815_; 
wire u5__abc_81276_new_n3816_; 
wire u5__abc_81276_new_n3817_; 
wire u5__abc_81276_new_n3818_; 
wire u5__abc_81276_new_n3819_; 
wire u5__abc_81276_new_n381_; 
wire u5__abc_81276_new_n3820_; 
wire u5__abc_81276_new_n3822_; 
wire u5__abc_81276_new_n3823_; 
wire u5__abc_81276_new_n3824_; 
wire u5__abc_81276_new_n3826_; 
wire u5__abc_81276_new_n3827_; 
wire u5__abc_81276_new_n3828_; 
wire u5__abc_81276_new_n3829_; 
wire u5__abc_81276_new_n382_; 
wire u5__abc_81276_new_n3830_; 
wire u5__abc_81276_new_n3832_; 
wire u5__abc_81276_new_n3833_; 
wire u5__abc_81276_new_n3834_; 
wire u5__abc_81276_new_n3835_; 
wire u5__abc_81276_new_n3836_; 
wire u5__abc_81276_new_n3838_; 
wire u5__abc_81276_new_n3839_; 
wire u5__abc_81276_new_n383_; 
wire u5__abc_81276_new_n3840_; 
wire u5__abc_81276_new_n3841_; 
wire u5__abc_81276_new_n3842_; 
wire u5__abc_81276_new_n3844_; 
wire u5__abc_81276_new_n3845_; 
wire u5__abc_81276_new_n3846_; 
wire u5__abc_81276_new_n3847_; 
wire u5__abc_81276_new_n3848_; 
wire u5__abc_81276_new_n3849_; 
wire u5__abc_81276_new_n384_; 
wire u5__abc_81276_new_n3850_; 
wire u5__abc_81276_new_n3851_; 
wire u5__abc_81276_new_n3852_; 
wire u5__abc_81276_new_n3853_; 
wire u5__abc_81276_new_n3855_; 
wire u5__abc_81276_new_n3856_; 
wire u5__abc_81276_new_n3857_; 
wire u5__abc_81276_new_n3858_; 
wire u5__abc_81276_new_n3859_; 
wire u5__abc_81276_new_n385_; 
wire u5__abc_81276_new_n3860_; 
wire u5__abc_81276_new_n3861_; 
wire u5__abc_81276_new_n3862_; 
wire u5__abc_81276_new_n3863_; 
wire u5__abc_81276_new_n3864_; 
wire u5__abc_81276_new_n3865_; 
wire u5__abc_81276_new_n3866_; 
wire u5__abc_81276_new_n3867_; 
wire u5__abc_81276_new_n3868_; 
wire u5__abc_81276_new_n3869_; 
wire u5__abc_81276_new_n3870_; 
wire u5__abc_81276_new_n3871_; 
wire u5__abc_81276_new_n3872_; 
wire u5__abc_81276_new_n3873_; 
wire u5__abc_81276_new_n3875_; 
wire u5__abc_81276_new_n3876_; 
wire u5__abc_81276_new_n3877_; 
wire u5__abc_81276_new_n3878_; 
wire u5__abc_81276_new_n3879_; 
wire u5__abc_81276_new_n387_; 
wire u5__abc_81276_new_n3880_; 
wire u5__abc_81276_new_n3881_; 
wire u5__abc_81276_new_n3882_; 
wire u5__abc_81276_new_n3883_; 
wire u5__abc_81276_new_n3885_; 
wire u5__abc_81276_new_n3886_; 
wire u5__abc_81276_new_n3887_; 
wire u5__abc_81276_new_n3888_; 
wire u5__abc_81276_new_n388_; 
wire u5__abc_81276_new_n3890_; 
wire u5__abc_81276_new_n3891_; 
wire u5__abc_81276_new_n3892_; 
wire u5__abc_81276_new_n3893_; 
wire u5__abc_81276_new_n3894_; 
wire u5__abc_81276_new_n3895_; 
wire u5__abc_81276_new_n3896_; 
wire u5__abc_81276_new_n3897_; 
wire u5__abc_81276_new_n3898_; 
wire u5__abc_81276_new_n3899_; 
wire u5__abc_81276_new_n389_; 
wire u5__abc_81276_new_n3900_; 
wire u5__abc_81276_new_n3901_; 
wire u5__abc_81276_new_n3902_; 
wire u5__abc_81276_new_n3903_; 
wire u5__abc_81276_new_n3905_; 
wire u5__abc_81276_new_n3906_; 
wire u5__abc_81276_new_n3907_; 
wire u5__abc_81276_new_n3908_; 
wire u5__abc_81276_new_n3909_; 
wire u5__abc_81276_new_n390_; 
wire u5__abc_81276_new_n3910_; 
wire u5__abc_81276_new_n3911_; 
wire u5__abc_81276_new_n3912_; 
wire u5__abc_81276_new_n3913_; 
wire u5__abc_81276_new_n3914_; 
wire u5__abc_81276_new_n3915_; 
wire u5__abc_81276_new_n3916_; 
wire u5__abc_81276_new_n3917_; 
wire u5__abc_81276_new_n3918_; 
wire u5__abc_81276_new_n3919_; 
wire u5__abc_81276_new_n391_; 
wire u5__abc_81276_new_n3920_; 
wire u5__abc_81276_new_n3921_; 
wire u5__abc_81276_new_n3922_; 
wire u5__abc_81276_new_n3923_; 
wire u5__abc_81276_new_n3924_; 
wire u5__abc_81276_new_n3925_; 
wire u5__abc_81276_new_n3927_; 
wire u5__abc_81276_new_n3928_; 
wire u5__abc_81276_new_n3929_; 
wire u5__abc_81276_new_n392_; 
wire u5__abc_81276_new_n3930_; 
wire u5__abc_81276_new_n3931_; 
wire u5__abc_81276_new_n3932_; 
wire u5__abc_81276_new_n3933_; 
wire u5__abc_81276_new_n3934_; 
wire u5__abc_81276_new_n3935_; 
wire u5__abc_81276_new_n3936_; 
wire u5__abc_81276_new_n3937_; 
wire u5__abc_81276_new_n3938_; 
wire u5__abc_81276_new_n3939_; 
wire u5__abc_81276_new_n393_; 
wire u5__abc_81276_new_n3940_; 
wire u5__abc_81276_new_n3941_; 
wire u5__abc_81276_new_n3942_; 
wire u5__abc_81276_new_n3943_; 
wire u5__abc_81276_new_n3944_; 
wire u5__abc_81276_new_n3945_; 
wire u5__abc_81276_new_n3947_; 
wire u5__abc_81276_new_n3948_; 
wire u5__abc_81276_new_n3949_; 
wire u5__abc_81276_new_n394_; 
wire u5__abc_81276_new_n3950_; 
wire u5__abc_81276_new_n3951_; 
wire u5__abc_81276_new_n3952_; 
wire u5__abc_81276_new_n3953_; 
wire u5__abc_81276_new_n3954_; 
wire u5__abc_81276_new_n3955_; 
wire u5__abc_81276_new_n3957_; 
wire u5__abc_81276_new_n3958_; 
wire u5__abc_81276_new_n3959_; 
wire u5__abc_81276_new_n395_; 
wire u5__abc_81276_new_n3960_; 
wire u5__abc_81276_new_n3961_; 
wire u5__abc_81276_new_n3962_; 
wire u5__abc_81276_new_n3963_; 
wire u5__abc_81276_new_n3965_; 
wire u5__abc_81276_new_n3966_; 
wire u5__abc_81276_new_n3967_; 
wire u5__abc_81276_new_n3968_; 
wire u5__abc_81276_new_n3969_; 
wire u5__abc_81276_new_n396_; 
wire u5__abc_81276_new_n3970_; 
wire u5__abc_81276_new_n3971_; 
wire u5__abc_81276_new_n3972_; 
wire u5__abc_81276_new_n3973_; 
wire u5__abc_81276_new_n3974_; 
wire u5__abc_81276_new_n3975_; 
wire u5__abc_81276_new_n3976_; 
wire u5__abc_81276_new_n3977_; 
wire u5__abc_81276_new_n3979_; 
wire u5__abc_81276_new_n397_; 
wire u5__abc_81276_new_n3980_; 
wire u5__abc_81276_new_n3981_; 
wire u5__abc_81276_new_n3982_; 
wire u5__abc_81276_new_n3984_; 
wire u5__abc_81276_new_n3985_; 
wire u5__abc_81276_new_n3986_; 
wire u5__abc_81276_new_n3987_; 
wire u5__abc_81276_new_n3988_; 
wire u5__abc_81276_new_n3989_; 
wire u5__abc_81276_new_n398_; 
wire u5__abc_81276_new_n3990_; 
wire u5__abc_81276_new_n3991_; 
wire u5__abc_81276_new_n3992_; 
wire u5__abc_81276_new_n3993_; 
wire u5__abc_81276_new_n3994_; 
wire u5__abc_81276_new_n3995_; 
wire u5__abc_81276_new_n3996_; 
wire u5__abc_81276_new_n3997_; 
wire u5__abc_81276_new_n3998_; 
wire u5__abc_81276_new_n3999_; 
wire u5__abc_81276_new_n399_; 
wire u5__abc_81276_new_n4000_; 
wire u5__abc_81276_new_n4001_; 
wire u5__abc_81276_new_n4002_; 
wire u5__abc_81276_new_n4003_; 
wire u5__abc_81276_new_n4004_; 
wire u5__abc_81276_new_n4005_; 
wire u5__abc_81276_new_n4006_; 
wire u5__abc_81276_new_n4007_; 
wire u5__abc_81276_new_n4008_; 
wire u5__abc_81276_new_n4009_; 
wire u5__abc_81276_new_n400_; 
wire u5__abc_81276_new_n4010_; 
wire u5__abc_81276_new_n4011_; 
wire u5__abc_81276_new_n4012_; 
wire u5__abc_81276_new_n4013_; 
wire u5__abc_81276_new_n4014_; 
wire u5__abc_81276_new_n4015_; 
wire u5__abc_81276_new_n4016_; 
wire u5__abc_81276_new_n4017_; 
wire u5__abc_81276_new_n4018_; 
wire u5__abc_81276_new_n4019_; 
wire u5__abc_81276_new_n401_; 
wire u5__abc_81276_new_n401__bF_buf0; 
wire u5__abc_81276_new_n401__bF_buf1; 
wire u5__abc_81276_new_n401__bF_buf2; 
wire u5__abc_81276_new_n401__bF_buf3; 
wire u5__abc_81276_new_n4020_; 
wire u5__abc_81276_new_n4021_; 
wire u5__abc_81276_new_n4022_; 
wire u5__abc_81276_new_n4023_; 
wire u5__abc_81276_new_n4024_; 
wire u5__abc_81276_new_n4026_; 
wire u5__abc_81276_new_n4027_; 
wire u5__abc_81276_new_n4028_; 
wire u5__abc_81276_new_n4029_; 
wire u5__abc_81276_new_n402_; 
wire u5__abc_81276_new_n4030_; 
wire u5__abc_81276_new_n4031_; 
wire u5__abc_81276_new_n4033_; 
wire u5__abc_81276_new_n4034_; 
wire u5__abc_81276_new_n4035_; 
wire u5__abc_81276_new_n4036_; 
wire u5__abc_81276_new_n4037_; 
wire u5__abc_81276_new_n4039_; 
wire u5__abc_81276_new_n403_; 
wire u5__abc_81276_new_n4040_; 
wire u5__abc_81276_new_n4042_; 
wire u5__abc_81276_new_n4043_; 
wire u5__abc_81276_new_n4045_; 
wire u5__abc_81276_new_n4046_; 
wire u5__abc_81276_new_n4047_; 
wire u5__abc_81276_new_n4048_; 
wire u5__abc_81276_new_n4049_; 
wire u5__abc_81276_new_n404_; 
wire u5__abc_81276_new_n4050_; 
wire u5__abc_81276_new_n4051_; 
wire u5__abc_81276_new_n4052_; 
wire u5__abc_81276_new_n4053_; 
wire u5__abc_81276_new_n4054_; 
wire u5__abc_81276_new_n4055_; 
wire u5__abc_81276_new_n4056_; 
wire u5__abc_81276_new_n4057_; 
wire u5__abc_81276_new_n4058_; 
wire u5__abc_81276_new_n4059_; 
wire u5__abc_81276_new_n405_; 
wire u5__abc_81276_new_n4061_; 
wire u5__abc_81276_new_n4064_; 
wire u5__abc_81276_new_n4065_; 
wire u5__abc_81276_new_n4066_; 
wire u5__abc_81276_new_n4067_; 
wire u5__abc_81276_new_n4068_; 
wire u5__abc_81276_new_n406_; 
wire u5__abc_81276_new_n4070_; 
wire u5__abc_81276_new_n4071_; 
wire u5__abc_81276_new_n4072_; 
wire u5__abc_81276_new_n4073_; 
wire u5__abc_81276_new_n4074_; 
wire u5__abc_81276_new_n4075_; 
wire u5__abc_81276_new_n4076_; 
wire u5__abc_81276_new_n4077_; 
wire u5__abc_81276_new_n4078_; 
wire u5__abc_81276_new_n4079_; 
wire u5__abc_81276_new_n407_; 
wire u5__abc_81276_new_n4080_; 
wire u5__abc_81276_new_n4082_; 
wire u5__abc_81276_new_n4083_; 
wire u5__abc_81276_new_n4084_; 
wire u5__abc_81276_new_n4086_; 
wire u5__abc_81276_new_n4087_; 
wire u5__abc_81276_new_n4088_; 
wire u5__abc_81276_new_n4089_; 
wire u5__abc_81276_new_n408_; 
wire u5__abc_81276_new_n4090_; 
wire u5__abc_81276_new_n4091_; 
wire u5__abc_81276_new_n409_; 
wire u5__abc_81276_new_n410_; 
wire u5__abc_81276_new_n411_; 
wire u5__abc_81276_new_n412_; 
wire u5__abc_81276_new_n413_; 
wire u5__abc_81276_new_n414_; 
wire u5__abc_81276_new_n415_; 
wire u5__abc_81276_new_n416_; 
wire u5__abc_81276_new_n416__bF_buf0; 
wire u5__abc_81276_new_n416__bF_buf1; 
wire u5__abc_81276_new_n416__bF_buf2; 
wire u5__abc_81276_new_n416__bF_buf3; 
wire u5__abc_81276_new_n417_; 
wire u5__abc_81276_new_n417__bF_buf0; 
wire u5__abc_81276_new_n417__bF_buf1; 
wire u5__abc_81276_new_n417__bF_buf2; 
wire u5__abc_81276_new_n417__bF_buf3; 
wire u5__abc_81276_new_n418_; 
wire u5__abc_81276_new_n419_; 
wire u5__abc_81276_new_n420_; 
wire u5__abc_81276_new_n421_; 
wire u5__abc_81276_new_n422_; 
wire u5__abc_81276_new_n423_; 
wire u5__abc_81276_new_n424_; 
wire u5__abc_81276_new_n425_; 
wire u5__abc_81276_new_n426_; 
wire u5__abc_81276_new_n427_; 
wire u5__abc_81276_new_n428_; 
wire u5__abc_81276_new_n429_; 
wire u5__abc_81276_new_n430_; 
wire u5__abc_81276_new_n431_; 
wire u5__abc_81276_new_n432_; 
wire u5__abc_81276_new_n433_; 
wire u5__abc_81276_new_n434_; 
wire u5__abc_81276_new_n435_; 
wire u5__abc_81276_new_n436_; 
wire u5__abc_81276_new_n437_; 
wire u5__abc_81276_new_n438_; 
wire u5__abc_81276_new_n439_; 
wire u5__abc_81276_new_n440_; 
wire u5__abc_81276_new_n441_; 
wire u5__abc_81276_new_n442_; 
wire u5__abc_81276_new_n443_; 
wire u5__abc_81276_new_n444_; 
wire u5__abc_81276_new_n445_; 
wire u5__abc_81276_new_n446_; 
wire u5__abc_81276_new_n447_; 
wire u5__abc_81276_new_n448_; 
wire u5__abc_81276_new_n448__bF_buf0; 
wire u5__abc_81276_new_n448__bF_buf1; 
wire u5__abc_81276_new_n448__bF_buf2; 
wire u5__abc_81276_new_n448__bF_buf3; 
wire u5__abc_81276_new_n448__bF_buf4; 
wire u5__abc_81276_new_n448__bF_buf5; 
wire u5__abc_81276_new_n449_; 
wire u5__abc_81276_new_n449__bF_buf0; 
wire u5__abc_81276_new_n449__bF_buf1; 
wire u5__abc_81276_new_n449__bF_buf2; 
wire u5__abc_81276_new_n449__bF_buf3; 
wire u5__abc_81276_new_n449__bF_buf4; 
wire u5__abc_81276_new_n449__bF_buf5; 
wire u5__abc_81276_new_n449__bF_buf6; 
wire u5__abc_81276_new_n449__bF_buf7; 
wire u5__abc_81276_new_n450_; 
wire u5__abc_81276_new_n451_; 
wire u5__abc_81276_new_n452_; 
wire u5__abc_81276_new_n453_; 
wire u5__abc_81276_new_n454_; 
wire u5__abc_81276_new_n455_; 
wire u5__abc_81276_new_n456_; 
wire u5__abc_81276_new_n457_; 
wire u5__abc_81276_new_n458_; 
wire u5__abc_81276_new_n459_; 
wire u5__abc_81276_new_n460_; 
wire u5__abc_81276_new_n461_; 
wire u5__abc_81276_new_n462_; 
wire u5__abc_81276_new_n463_; 
wire u5__abc_81276_new_n464_; 
wire u5__abc_81276_new_n464__bF_buf0; 
wire u5__abc_81276_new_n464__bF_buf1; 
wire u5__abc_81276_new_n464__bF_buf2; 
wire u5__abc_81276_new_n464__bF_buf3; 
wire u5__abc_81276_new_n465_; 
wire u5__abc_81276_new_n466_; 
wire u5__abc_81276_new_n467_; 
wire u5__abc_81276_new_n468_; 
wire u5__abc_81276_new_n469_; 
wire u5__abc_81276_new_n470_; 
wire u5__abc_81276_new_n471_; 
wire u5__abc_81276_new_n472_; 
wire u5__abc_81276_new_n473_; 
wire u5__abc_81276_new_n474_; 
wire u5__abc_81276_new_n475_; 
wire u5__abc_81276_new_n476_; 
wire u5__abc_81276_new_n477_; 
wire u5__abc_81276_new_n478_; 
wire u5__abc_81276_new_n479_; 
wire u5__abc_81276_new_n479__bF_buf0; 
wire u5__abc_81276_new_n479__bF_buf1; 
wire u5__abc_81276_new_n479__bF_buf2; 
wire u5__abc_81276_new_n479__bF_buf3; 
wire u5__abc_81276_new_n480_; 
wire u5__abc_81276_new_n480__bF_buf0; 
wire u5__abc_81276_new_n480__bF_buf1; 
wire u5__abc_81276_new_n480__bF_buf2; 
wire u5__abc_81276_new_n480__bF_buf3; 
wire u5__abc_81276_new_n480__bF_buf4; 
wire u5__abc_81276_new_n481_; 
wire u5__abc_81276_new_n482_; 
wire u5__abc_81276_new_n483_; 
wire u5__abc_81276_new_n484_; 
wire u5__abc_81276_new_n485_; 
wire u5__abc_81276_new_n486_; 
wire u5__abc_81276_new_n487_; 
wire u5__abc_81276_new_n488_; 
wire u5__abc_81276_new_n489_; 
wire u5__abc_81276_new_n490_; 
wire u5__abc_81276_new_n490__bF_buf0; 
wire u5__abc_81276_new_n490__bF_buf1; 
wire u5__abc_81276_new_n490__bF_buf10; 
wire u5__abc_81276_new_n490__bF_buf2; 
wire u5__abc_81276_new_n490__bF_buf3; 
wire u5__abc_81276_new_n490__bF_buf4; 
wire u5__abc_81276_new_n490__bF_buf5; 
wire u5__abc_81276_new_n490__bF_buf6; 
wire u5__abc_81276_new_n490__bF_buf7; 
wire u5__abc_81276_new_n490__bF_buf8; 
wire u5__abc_81276_new_n490__bF_buf9; 
wire u5__abc_81276_new_n491_; 
wire u5__abc_81276_new_n492_; 
wire u5__abc_81276_new_n493_; 
wire u5__abc_81276_new_n494_; 
wire u5__abc_81276_new_n495_; 
wire u5__abc_81276_new_n496_; 
wire u5__abc_81276_new_n497_; 
wire u5__abc_81276_new_n498_; 
wire u5__abc_81276_new_n499_; 
wire u5__abc_81276_new_n500_; 
wire u5__abc_81276_new_n501_; 
wire u5__abc_81276_new_n502_; 
wire u5__abc_81276_new_n503_; 
wire u5__abc_81276_new_n504_; 
wire u5__abc_81276_new_n505_; 
wire u5__abc_81276_new_n506_; 
wire u5__abc_81276_new_n507_; 
wire u5__abc_81276_new_n508_; 
wire u5__abc_81276_new_n509_; 
wire u5__abc_81276_new_n510_; 
wire u5__abc_81276_new_n511_; 
wire u5__abc_81276_new_n512_; 
wire u5__abc_81276_new_n513_; 
wire u5__abc_81276_new_n514_; 
wire u5__abc_81276_new_n515_; 
wire u5__abc_81276_new_n516_; 
wire u5__abc_81276_new_n517_; 
wire u5__abc_81276_new_n518_; 
wire u5__abc_81276_new_n519_; 
wire u5__abc_81276_new_n520_; 
wire u5__abc_81276_new_n521_; 
wire u5__abc_81276_new_n521__bF_buf0; 
wire u5__abc_81276_new_n521__bF_buf1; 
wire u5__abc_81276_new_n521__bF_buf2; 
wire u5__abc_81276_new_n521__bF_buf3; 
wire u5__abc_81276_new_n522_; 
wire u5__abc_81276_new_n522__bF_buf0; 
wire u5__abc_81276_new_n522__bF_buf1; 
wire u5__abc_81276_new_n522__bF_buf2; 
wire u5__abc_81276_new_n522__bF_buf3; 
wire u5__abc_81276_new_n522__bF_buf4; 
wire u5__abc_81276_new_n523_; 
wire u5__abc_81276_new_n523__bF_buf0; 
wire u5__abc_81276_new_n523__bF_buf1; 
wire u5__abc_81276_new_n523__bF_buf2; 
wire u5__abc_81276_new_n523__bF_buf3; 
wire u5__abc_81276_new_n523__bF_buf4; 
wire u5__abc_81276_new_n523__bF_buf5; 
wire u5__abc_81276_new_n523__bF_buf6; 
wire u5__abc_81276_new_n523__bF_buf7; 
wire u5__abc_81276_new_n524_; 
wire u5__abc_81276_new_n525_; 
wire u5__abc_81276_new_n526_; 
wire u5__abc_81276_new_n527_; 
wire u5__abc_81276_new_n528_; 
wire u5__abc_81276_new_n529_; 
wire u5__abc_81276_new_n530_; 
wire u5__abc_81276_new_n531_; 
wire u5__abc_81276_new_n532_; 
wire u5__abc_81276_new_n533_; 
wire u5__abc_81276_new_n534_; 
wire u5__abc_81276_new_n535_; 
wire u5__abc_81276_new_n536_; 
wire u5__abc_81276_new_n537_; 
wire u5__abc_81276_new_n538_; 
wire u5__abc_81276_new_n540_; 
wire u5__abc_81276_new_n541_; 
wire u5__abc_81276_new_n542_; 
wire u5__abc_81276_new_n543_; 
wire u5__abc_81276_new_n544_; 
wire u5__abc_81276_new_n545_; 
wire u5__abc_81276_new_n546_; 
wire u5__abc_81276_new_n547_; 
wire u5__abc_81276_new_n548_; 
wire u5__abc_81276_new_n549_; 
wire u5__abc_81276_new_n550_; 
wire u5__abc_81276_new_n551_; 
wire u5__abc_81276_new_n552_; 
wire u5__abc_81276_new_n553_; 
wire u5__abc_81276_new_n554_; 
wire u5__abc_81276_new_n555_; 
wire u5__abc_81276_new_n556_; 
wire u5__abc_81276_new_n557_; 
wire u5__abc_81276_new_n558_; 
wire u5__abc_81276_new_n559_; 
wire u5__abc_81276_new_n560_; 
wire u5__abc_81276_new_n561_; 
wire u5__abc_81276_new_n562_; 
wire u5__abc_81276_new_n563_; 
wire u5__abc_81276_new_n564_; 
wire u5__abc_81276_new_n565_; 
wire u5__abc_81276_new_n566_; 
wire u5__abc_81276_new_n567_; 
wire u5__abc_81276_new_n568_; 
wire u5__abc_81276_new_n569_; 
wire u5__abc_81276_new_n570_; 
wire u5__abc_81276_new_n571_; 
wire u5__abc_81276_new_n572_; 
wire u5__abc_81276_new_n573_; 
wire u5__abc_81276_new_n574_; 
wire u5__abc_81276_new_n575_; 
wire u5__abc_81276_new_n576_; 
wire u5__abc_81276_new_n577_; 
wire u5__abc_81276_new_n578_; 
wire u5__abc_81276_new_n579_; 
wire u5__abc_81276_new_n580_; 
wire u5__abc_81276_new_n581_; 
wire u5__abc_81276_new_n582_; 
wire u5__abc_81276_new_n583_; 
wire u5__abc_81276_new_n584_; 
wire u5__abc_81276_new_n585_; 
wire u5__abc_81276_new_n586_; 
wire u5__abc_81276_new_n587_; 
wire u5__abc_81276_new_n588_; 
wire u5__abc_81276_new_n589_; 
wire u5__abc_81276_new_n590_; 
wire u5__abc_81276_new_n591_; 
wire u5__abc_81276_new_n592_; 
wire u5__abc_81276_new_n593_; 
wire u5__abc_81276_new_n594_; 
wire u5__abc_81276_new_n595_; 
wire u5__abc_81276_new_n596_; 
wire u5__abc_81276_new_n597_; 
wire u5__abc_81276_new_n598_; 
wire u5__abc_81276_new_n599_; 
wire u5__abc_81276_new_n600_; 
wire u5__abc_81276_new_n601_; 
wire u5__abc_81276_new_n602_; 
wire u5__abc_81276_new_n603_; 
wire u5__abc_81276_new_n604_; 
wire u5__abc_81276_new_n605_; 
wire u5__abc_81276_new_n606_; 
wire u5__abc_81276_new_n607_; 
wire u5__abc_81276_new_n608_; 
wire u5__abc_81276_new_n609_; 
wire u5__abc_81276_new_n610_; 
wire u5__abc_81276_new_n611_; 
wire u5__abc_81276_new_n612_; 
wire u5__abc_81276_new_n613_; 
wire u5__abc_81276_new_n614_; 
wire u5__abc_81276_new_n615_; 
wire u5__abc_81276_new_n616_; 
wire u5__abc_81276_new_n617_; 
wire u5__abc_81276_new_n618_; 
wire u5__abc_81276_new_n619_; 
wire u5__abc_81276_new_n620_; 
wire u5__abc_81276_new_n621_; 
wire u5__abc_81276_new_n622_; 
wire u5__abc_81276_new_n623_; 
wire u5__abc_81276_new_n624_; 
wire u5__abc_81276_new_n625_; 
wire u5__abc_81276_new_n626_; 
wire u5__abc_81276_new_n627_; 
wire u5__abc_81276_new_n628_; 
wire u5__abc_81276_new_n629_; 
wire u5__abc_81276_new_n630_; 
wire u5__abc_81276_new_n631_; 
wire u5__abc_81276_new_n632_; 
wire u5__abc_81276_new_n633_; 
wire u5__abc_81276_new_n634_; 
wire u5__abc_81276_new_n635_; 
wire u5__abc_81276_new_n636_; 
wire u5__abc_81276_new_n637_; 
wire u5__abc_81276_new_n638_; 
wire u5__abc_81276_new_n639_; 
wire u5__abc_81276_new_n640_; 
wire u5__abc_81276_new_n641_; 
wire u5__abc_81276_new_n642_; 
wire u5__abc_81276_new_n643_; 
wire u5__abc_81276_new_n644_; 
wire u5__abc_81276_new_n645_; 
wire u5__abc_81276_new_n646_; 
wire u5__abc_81276_new_n647_; 
wire u5__abc_81276_new_n648_; 
wire u5__abc_81276_new_n649_; 
wire u5__abc_81276_new_n650_; 
wire u5__abc_81276_new_n651_; 
wire u5__abc_81276_new_n652_; 
wire u5__abc_81276_new_n653_; 
wire u5__abc_81276_new_n654_; 
wire u5__abc_81276_new_n655_; 
wire u5__abc_81276_new_n656_; 
wire u5__abc_81276_new_n657_; 
wire u5__abc_81276_new_n658_; 
wire u5__abc_81276_new_n659_; 
wire u5__abc_81276_new_n660_; 
wire u5__abc_81276_new_n661_; 
wire u5__abc_81276_new_n662_; 
wire u5__abc_81276_new_n663_; 
wire u5__abc_81276_new_n664_; 
wire u5__abc_81276_new_n665_; 
wire u5__abc_81276_new_n666_; 
wire u5__abc_81276_new_n667_; 
wire u5__abc_81276_new_n668_; 
wire u5__abc_81276_new_n669_; 
wire u5__abc_81276_new_n670_; 
wire u5__abc_81276_new_n671_; 
wire u5__abc_81276_new_n672_; 
wire u5__abc_81276_new_n673_; 
wire u5__abc_81276_new_n674_; 
wire u5__abc_81276_new_n675_; 
wire u5__abc_81276_new_n676_; 
wire u5__abc_81276_new_n677_; 
wire u5__abc_81276_new_n678_; 
wire u5__abc_81276_new_n679_; 
wire u5__abc_81276_new_n680_; 
wire u5__abc_81276_new_n681_; 
wire u5__abc_81276_new_n682_; 
wire u5__abc_81276_new_n683_; 
wire u5__abc_81276_new_n684_; 
wire u5__abc_81276_new_n685_; 
wire u5__abc_81276_new_n686_; 
wire u5__abc_81276_new_n687_; 
wire u5__abc_81276_new_n688_; 
wire u5__abc_81276_new_n689_; 
wire u5__abc_81276_new_n690_; 
wire u5__abc_81276_new_n691_; 
wire u5__abc_81276_new_n692_; 
wire u5__abc_81276_new_n693_; 
wire u5__abc_81276_new_n694_; 
wire u5__abc_81276_new_n695_; 
wire u5__abc_81276_new_n696_; 
wire u5__abc_81276_new_n697_; 
wire u5__abc_81276_new_n698_; 
wire u5__abc_81276_new_n699_; 
wire u5__abc_81276_new_n700_; 
wire u5__abc_81276_new_n701_; 
wire u5__abc_81276_new_n702_; 
wire u5__abc_81276_new_n703_; 
wire u5__abc_81276_new_n704_; 
wire u5__abc_81276_new_n705_; 
wire u5__abc_81276_new_n706_; 
wire u5__abc_81276_new_n707_; 
wire u5__abc_81276_new_n708_; 
wire u5__abc_81276_new_n709_; 
wire u5__abc_81276_new_n710_; 
wire u5__abc_81276_new_n711_; 
wire u5__abc_81276_new_n712_; 
wire u5__abc_81276_new_n713_; 
wire u5__abc_81276_new_n714_; 
wire u5__abc_81276_new_n715_; 
wire u5__abc_81276_new_n716_; 
wire u5__abc_81276_new_n717_; 
wire u5__abc_81276_new_n718_; 
wire u5__abc_81276_new_n719_; 
wire u5__abc_81276_new_n720_; 
wire u5__abc_81276_new_n721_; 
wire u5__abc_81276_new_n722_; 
wire u5__abc_81276_new_n723_; 
wire u5__abc_81276_new_n724_; 
wire u5__abc_81276_new_n725_; 
wire u5__abc_81276_new_n726_; 
wire u5__abc_81276_new_n727_; 
wire u5__abc_81276_new_n728_; 
wire u5__abc_81276_new_n729_; 
wire u5__abc_81276_new_n730_; 
wire u5__abc_81276_new_n731_; 
wire u5__abc_81276_new_n732_; 
wire u5__abc_81276_new_n733_; 
wire u5__abc_81276_new_n734_; 
wire u5__abc_81276_new_n735_; 
wire u5__abc_81276_new_n736_; 
wire u5__abc_81276_new_n737_; 
wire u5__abc_81276_new_n738_; 
wire u5__abc_81276_new_n739_; 
wire u5__abc_81276_new_n740_; 
wire u5__abc_81276_new_n741_; 
wire u5__abc_81276_new_n742_; 
wire u5__abc_81276_new_n743_; 
wire u5__abc_81276_new_n744_; 
wire u5__abc_81276_new_n745_; 
wire u5__abc_81276_new_n746_; 
wire u5__abc_81276_new_n747_; 
wire u5__abc_81276_new_n748_; 
wire u5__abc_81276_new_n749_; 
wire u5__abc_81276_new_n750_; 
wire u5__abc_81276_new_n751_; 
wire u5__abc_81276_new_n752_; 
wire u5__abc_81276_new_n753_; 
wire u5__abc_81276_new_n754_; 
wire u5__abc_81276_new_n755_; 
wire u5__abc_81276_new_n756_; 
wire u5__abc_81276_new_n757_; 
wire u5__abc_81276_new_n758_; 
wire u5__abc_81276_new_n759_; 
wire u5__abc_81276_new_n760_; 
wire u5__abc_81276_new_n761_; 
wire u5__abc_81276_new_n762_; 
wire u5__abc_81276_new_n763_; 
wire u5__abc_81276_new_n764_; 
wire u5__abc_81276_new_n765_; 
wire u5__abc_81276_new_n766_; 
wire u5__abc_81276_new_n767_; 
wire u5__abc_81276_new_n768_; 
wire u5__abc_81276_new_n769_; 
wire u5__abc_81276_new_n770_; 
wire u5__abc_81276_new_n771_; 
wire u5__abc_81276_new_n772_; 
wire u5__abc_81276_new_n773_; 
wire u5__abc_81276_new_n774_; 
wire u5__abc_81276_new_n775_; 
wire u5__abc_81276_new_n776_; 
wire u5__abc_81276_new_n777_; 
wire u5__abc_81276_new_n778_; 
wire u5__abc_81276_new_n779_; 
wire u5__abc_81276_new_n780_; 
wire u5__abc_81276_new_n781_; 
wire u5__abc_81276_new_n782_; 
wire u5__abc_81276_new_n783_; 
wire u5__abc_81276_new_n784_; 
wire u5__abc_81276_new_n785_; 
wire u5__abc_81276_new_n786_; 
wire u5__abc_81276_new_n787_; 
wire u5__abc_81276_new_n788_; 
wire u5__abc_81276_new_n789_; 
wire u5__abc_81276_new_n790_; 
wire u5__abc_81276_new_n791_; 
wire u5__abc_81276_new_n792_; 
wire u5__abc_81276_new_n793_; 
wire u5__abc_81276_new_n794_; 
wire u5__abc_81276_new_n795_; 
wire u5__abc_81276_new_n796_; 
wire u5__abc_81276_new_n797_; 
wire u5__abc_81276_new_n798_; 
wire u5__abc_81276_new_n799_; 
wire u5__abc_81276_new_n800_; 
wire u5__abc_81276_new_n801_; 
wire u5__abc_81276_new_n802_; 
wire u5__abc_81276_new_n803_; 
wire u5__abc_81276_new_n804_; 
wire u5__abc_81276_new_n805_; 
wire u5__abc_81276_new_n806_; 
wire u5__abc_81276_new_n807_; 
wire u5__abc_81276_new_n808_; 
wire u5__abc_81276_new_n809_; 
wire u5__abc_81276_new_n810_; 
wire u5__abc_81276_new_n811_; 
wire u5__abc_81276_new_n812_; 
wire u5__abc_81276_new_n813_; 
wire u5__abc_81276_new_n814_; 
wire u5__abc_81276_new_n815_; 
wire u5__abc_81276_new_n816_; 
wire u5__abc_81276_new_n817_; 
wire u5__abc_81276_new_n818_; 
wire u5__abc_81276_new_n819_; 
wire u5__abc_81276_new_n820_; 
wire u5__abc_81276_new_n821_; 
wire u5__abc_81276_new_n822_; 
wire u5__abc_81276_new_n823_; 
wire u5__abc_81276_new_n824_; 
wire u5__abc_81276_new_n825_; 
wire u5__abc_81276_new_n826_; 
wire u5__abc_81276_new_n827_; 
wire u5__abc_81276_new_n828_; 
wire u5__abc_81276_new_n829_; 
wire u5__abc_81276_new_n830_; 
wire u5__abc_81276_new_n831_; 
wire u5__abc_81276_new_n832_; 
wire u5__abc_81276_new_n833_; 
wire u5__abc_81276_new_n834_; 
wire u5__abc_81276_new_n835_; 
wire u5__abc_81276_new_n836_; 
wire u5__abc_81276_new_n837_; 
wire u5__abc_81276_new_n838_; 
wire u5__abc_81276_new_n839_; 
wire u5__abc_81276_new_n840_; 
wire u5__abc_81276_new_n841_; 
wire u5__abc_81276_new_n842_; 
wire u5__abc_81276_new_n843_; 
wire u5__abc_81276_new_n844_; 
wire u5__abc_81276_new_n845_; 
wire u5__abc_81276_new_n846_; 
wire u5__abc_81276_new_n847_; 
wire u5__abc_81276_new_n848_; 
wire u5__abc_81276_new_n849_; 
wire u5__abc_81276_new_n850_; 
wire u5__abc_81276_new_n851_; 
wire u5__abc_81276_new_n852_; 
wire u5__abc_81276_new_n853_; 
wire u5__abc_81276_new_n854_; 
wire u5__abc_81276_new_n855_; 
wire u5__abc_81276_new_n856_; 
wire u5__abc_81276_new_n857_; 
wire u5__abc_81276_new_n858_; 
wire u5__abc_81276_new_n859_; 
wire u5__abc_81276_new_n860_; 
wire u5__abc_81276_new_n861_; 
wire u5__abc_81276_new_n862_; 
wire u5__abc_81276_new_n863_; 
wire u5__abc_81276_new_n864_; 
wire u5__abc_81276_new_n865_; 
wire u5__abc_81276_new_n866_; 
wire u5__abc_81276_new_n867_; 
wire u5__abc_81276_new_n868_; 
wire u5__abc_81276_new_n869_; 
wire u5__abc_81276_new_n870_; 
wire u5__abc_81276_new_n871_; 
wire u5__abc_81276_new_n872_; 
wire u5__abc_81276_new_n873_; 
wire u5__abc_81276_new_n874_; 
wire u5__abc_81276_new_n875_; 
wire u5__abc_81276_new_n876_; 
wire u5__abc_81276_new_n877_; 
wire u5__abc_81276_new_n878_; 
wire u5__abc_81276_new_n879_; 
wire u5__abc_81276_new_n880_; 
wire u5__abc_81276_new_n881_; 
wire u5__abc_81276_new_n882_; 
wire u5__abc_81276_new_n883_; 
wire u5__abc_81276_new_n884_; 
wire u5__abc_81276_new_n885_; 
wire u5__abc_81276_new_n886_; 
wire u5__abc_81276_new_n887_; 
wire u5__abc_81276_new_n888_; 
wire u5__abc_81276_new_n889_; 
wire u5__abc_81276_new_n890_; 
wire u5__abc_81276_new_n891_; 
wire u5__abc_81276_new_n892_; 
wire u5__abc_81276_new_n893_; 
wire u5__abc_81276_new_n894_; 
wire u5__abc_81276_new_n895_; 
wire u5__abc_81276_new_n896_; 
wire u5__abc_81276_new_n897_; 
wire u5__abc_81276_new_n898_; 
wire u5__abc_81276_new_n899_; 
wire u5__abc_81276_new_n900_; 
wire u5__abc_81276_new_n901_; 
wire u5__abc_81276_new_n902_; 
wire u5__abc_81276_new_n903_; 
wire u5__abc_81276_new_n904_; 
wire u5__abc_81276_new_n905_; 
wire u5__abc_81276_new_n906_; 
wire u5__abc_81276_new_n907_; 
wire u5__abc_81276_new_n908_; 
wire u5__abc_81276_new_n909_; 
wire u5__abc_81276_new_n910_; 
wire u5__abc_81276_new_n911_; 
wire u5__abc_81276_new_n912_; 
wire u5__abc_81276_new_n913_; 
wire u5__abc_81276_new_n914_; 
wire u5__abc_81276_new_n915_; 
wire u5__abc_81276_new_n916_; 
wire u5__abc_81276_new_n917_; 
wire u5__abc_81276_new_n918_; 
wire u5__abc_81276_new_n919_; 
wire u5__abc_81276_new_n920_; 
wire u5__abc_81276_new_n921_; 
wire u5__abc_81276_new_n922_; 
wire u5__abc_81276_new_n923_; 
wire u5__abc_81276_new_n924_; 
wire u5__abc_81276_new_n925_; 
wire u5__abc_81276_new_n926_; 
wire u5__abc_81276_new_n927_; 
wire u5__abc_81276_new_n928_; 
wire u5__abc_81276_new_n929_; 
wire u5__abc_81276_new_n930_; 
wire u5__abc_81276_new_n931_; 
wire u5__abc_81276_new_n932_; 
wire u5__abc_81276_new_n933_; 
wire u5__abc_81276_new_n934_; 
wire u5__abc_81276_new_n935_; 
wire u5__abc_81276_new_n936_; 
wire u5__abc_81276_new_n937_; 
wire u5__abc_81276_new_n938_; 
wire u5__abc_81276_new_n939_; 
wire u5__abc_81276_new_n940_; 
wire u5__abc_81276_new_n941_; 
wire u5__abc_81276_new_n942_; 
wire u5__abc_81276_new_n943_; 
wire u5__abc_81276_new_n944_; 
wire u5__abc_81276_new_n945_; 
wire u5__abc_81276_new_n946_; 
wire u5__abc_81276_new_n947_; 
wire u5__abc_81276_new_n948_; 
wire u5__abc_81276_new_n949_; 
wire u5__abc_81276_new_n950_; 
wire u5__abc_81276_new_n951_; 
wire u5__abc_81276_new_n952_; 
wire u5__abc_81276_new_n953_; 
wire u5__abc_81276_new_n954_; 
wire u5__abc_81276_new_n955_; 
wire u5__abc_81276_new_n956_; 
wire u5__abc_81276_new_n957_; 
wire u5__abc_81276_new_n958_; 
wire u5__abc_81276_new_n959_; 
wire u5__abc_81276_new_n960_; 
wire u5__abc_81276_new_n961_; 
wire u5__abc_81276_new_n962_; 
wire u5__abc_81276_new_n963_; 
wire u5__abc_81276_new_n964_; 
wire u5__abc_81276_new_n965_; 
wire u5__abc_81276_new_n966_; 
wire u5__abc_81276_new_n967_; 
wire u5__abc_81276_new_n968_; 
wire u5__abc_81276_new_n969_; 
wire u5__abc_81276_new_n970_; 
wire u5__abc_81276_new_n971_; 
wire u5__abc_81276_new_n972_; 
wire u5__abc_81276_new_n973_; 
wire u5__abc_81276_new_n974_; 
wire u5__abc_81276_new_n975_; 
wire u5__abc_81276_new_n976_; 
wire u5__abc_81276_new_n977_; 
wire u5__abc_81276_new_n978_; 
wire u5__abc_81276_new_n979_; 
wire u5__abc_81276_new_n980_; 
wire u5__abc_81276_new_n981_; 
wire u5__abc_81276_new_n982_; 
wire u5__abc_81276_new_n983_; 
wire u5__abc_81276_new_n984_; 
wire u5__abc_81276_new_n985_; 
wire u5__abc_81276_new_n986_; 
wire u5__abc_81276_new_n987_; 
wire u5__abc_81276_new_n988_; 
wire u5__abc_81276_new_n989_; 
wire u5__abc_81276_new_n990_; 
wire u5__abc_81276_new_n991_; 
wire u5__abc_81276_new_n992_; 
wire u5__abc_81276_new_n993_; 
wire u5__abc_81276_new_n994_; 
wire u5__abc_81276_new_n995_; 
wire u5__abc_81276_new_n996_; 
wire u5__abc_81276_new_n997_; 
wire u5__abc_81276_new_n998_; 
wire u5__abc_81276_new_n999_; 
wire u5_ack_cnt_0_; 
wire u5_ack_cnt_1_; 
wire u5_ack_cnt_2_; 
wire u5_ack_cnt_3_; 
wire u5_ap_en; 
wire u5_burst_act_rd; 
wire u5_burst_cnt_0_; 
wire u5_burst_cnt_10_; 
wire u5_burst_cnt_1_; 
wire u5_burst_cnt_2_; 
wire u5_burst_cnt_3_; 
wire u5_burst_cnt_4_; 
wire u5_burst_cnt_5_; 
wire u5_burst_cnt_6_; 
wire u5_burst_cnt_7_; 
wire u5_burst_cnt_8_; 
wire u5_burst_cnt_9_; 
wire u5_cke_d; 
wire u5_cke_o_del; 
wire u5_cke_o_r1; 
wire u5_cke_o_r2; 
wire u5_cke_r; 
wire u5_cmd_0_; 
wire u5_cmd_1_; 
wire u5_cmd_2_; 
wire u5_cmd_3_; 
wire u5_cmd_a10_r; 
wire u5_cmd_asserted; 
wire u5_cmd_asserted2; 
wire u5_cmd_asserted_bF_buf0; 
wire u5_cmd_asserted_bF_buf1; 
wire u5_cmd_asserted_bF_buf2; 
wire u5_cmd_asserted_bF_buf3; 
wire u5_cmd_del_0_; 
wire u5_cmd_del_1_; 
wire u5_cmd_del_2_; 
wire u5_cmd_del_3_; 
wire u5_cmd_r_0_; 
wire u5_cmd_r_1_; 
wire u5_cmd_r_2_; 
wire u5_cmd_r_3_; 
wire u5_cnt; 
wire u5_cnt_next; 
wire u5_cs_le_r; 
wire u5_cs_le_r1; 
wire u5_data_oe_d; 
wire u5_data_oe_r; 
wire u5_data_oe_r2; 
wire u5_dv_r; 
wire u5_ir_cnt_0_; 
wire u5_ir_cnt_1_; 
wire u5_ir_cnt_2_; 
wire u5_ir_cnt_3_; 
wire u5_ir_cnt_done; 
wire u5_kro; 
wire u5_lmr_ack_d; 
wire u5_lookup_ready1; 
wire u5_lookup_ready2; 
wire u5_mc_adv_r; 
wire u5_mc_adv_r1; 
wire u5_mc_c_oe_d; 
wire u5_mc_le; 
wire u5_mem_ack_r; 
wire u5_next_state_0_; 
wire u5_next_state_10_; 
wire u5_next_state_11_; 
wire u5_next_state_12_; 
wire u5_next_state_13_; 
wire u5_next_state_14_; 
wire u5_next_state_15_; 
wire u5_next_state_16_; 
wire u5_next_state_17_; 
wire u5_next_state_18_; 
wire u5_next_state_19_; 
wire u5_next_state_1_; 
wire u5_next_state_20_; 
wire u5_next_state_21_; 
wire u5_next_state_22_; 
wire u5_next_state_23_; 
wire u5_next_state_24_; 
wire u5_next_state_25_; 
wire u5_next_state_26_; 
wire u5_next_state_27_; 
wire u5_next_state_28_; 
wire u5_next_state_29_; 
wire u5_next_state_2_; 
wire u5_next_state_30_; 
wire u5_next_state_31_; 
wire u5_next_state_32_; 
wire u5_next_state_33_; 
wire u5_next_state_34_; 
wire u5_next_state_35_; 
wire u5_next_state_36_; 
wire u5_next_state_37_; 
wire u5_next_state_38_; 
wire u5_next_state_39_; 
wire u5_next_state_3_; 
wire u5_next_state_40_; 
wire u5_next_state_41_; 
wire u5_next_state_42_; 
wire u5_next_state_43_; 
wire u5_next_state_44_; 
wire u5_next_state_45_; 
wire u5_next_state_46_; 
wire u5_next_state_47_; 
wire u5_next_state_48_; 
wire u5_next_state_49_; 
wire u5_next_state_4_; 
wire u5_next_state_50_; 
wire u5_next_state_51_; 
wire u5_next_state_52_; 
wire u5_next_state_53_; 
wire u5_next_state_54_; 
wire u5_next_state_55_; 
wire u5_next_state_56_; 
wire u5_next_state_57_; 
wire u5_next_state_58_; 
wire u5_next_state_59_; 
wire u5_next_state_5_; 
wire u5_next_state_60_; 
wire u5_next_state_61_; 
wire u5_next_state_62_; 
wire u5_next_state_63_; 
wire u5_next_state_64_; 
wire u5_next_state_65_; 
wire u5_next_state_6_; 
wire u5_next_state_7_; 
wire u5_next_state_8_; 
wire u5_next_state_9_; 
wire u5_no_wb_cycle; 
wire u5_pack_le0_d; 
wire u5_pack_le1_d; 
wire u5_pack_le2_d; 
wire u5_resume_req_r; 
wire u5_rfr_ack_d; 
wire u5_rsts; 
wire u5_state_0_; 
wire u5_state_10_; 
wire u5_state_11_; 
wire u5_state_12_; 
wire u5_state_13_; 
wire u5_state_14_; 
wire u5_state_15_; 
wire u5_state_16_; 
wire u5_state_17_; 
wire u5_state_18_; 
wire u5_state_19_; 
wire u5_state_1_; 
wire u5_state_20_; 
wire u5_state_21_; 
wire u5_state_22_; 
wire u5_state_23_; 
wire u5_state_24_; 
wire u5_state_25_; 
wire u5_state_26_; 
wire u5_state_27_; 
wire u5_state_28_; 
wire u5_state_29_; 
wire u5_state_2_; 
wire u5_state_30_; 
wire u5_state_31_; 
wire u5_state_32_; 
wire u5_state_33_; 
wire u5_state_34_; 
wire u5_state_35_; 
wire u5_state_36_; 
wire u5_state_37_; 
wire u5_state_38_; 
wire u5_state_39_; 
wire u5_state_3_; 
wire u5_state_40_; 
wire u5_state_41_; 
wire u5_state_42_; 
wire u5_state_43_; 
wire u5_state_44_; 
wire u5_state_45_; 
wire u5_state_46_; 
wire u5_state_47_; 
wire u5_state_48_; 
wire u5_state_49_; 
wire u5_state_4_; 
wire u5_state_50_; 
wire u5_state_51_; 
wire u5_state_52_; 
wire u5_state_53_; 
wire u5_state_54_; 
wire u5_state_55_; 
wire u5_state_56_; 
wire u5_state_57_; 
wire u5_state_58_; 
wire u5_state_59_; 
wire u5_state_5_; 
wire u5_state_60_; 
wire u5_state_61_; 
wire u5_state_62_; 
wire u5_state_63_; 
wire u5_state_64_; 
wire u5_state_65_; 
wire u5_state_6_; 
wire u5_state_7_; 
wire u5_state_8_; 
wire u5_state_9_; 
wire u5_susp_req_r; 
wire u5_suspended_d; 
wire u5_timer2_0_; 
wire u5_timer2_1_; 
wire u5_timer2_2_; 
wire u5_timer2_3_; 
wire u5_timer2_4_; 
wire u5_timer2_5_; 
wire u5_timer2_6_; 
wire u5_timer2_7_; 
wire u5_timer2_8_; 
wire u5_timer_0_; 
wire u5_timer_1_; 
wire u5_timer_2_; 
wire u5_timer_3_; 
wire u5_timer_4_; 
wire u5_timer_5_; 
wire u5_timer_6_; 
wire u5_timer_7_; 
wire u5_timer_is_zero; 
wire u5_tmr2_done; 
wire u5_tmr_done; 
wire u5_tmr_done_bF_buf0; 
wire u5_tmr_done_bF_buf1; 
wire u5_tmr_done_bF_buf2; 
wire u5_tmr_done_bF_buf3; 
wire u5_wb_cycle; 
wire u5_wb_first; 
wire u5_wb_stb_first; 
wire u5_wb_wait; 
wire u5_wb_wait_r; 
wire u5_wb_wait_r2; 
wire u5_wb_write_go_r; 
wire u5_we_; 
wire u6__0read_go_r1_0_0_; 
wire u6__0read_go_r_0_0_; 
wire u6__0rmw_en_0_0_; 
wire u6__0rmw_r_0_0_; 
wire u6__0wb_ack_o_0_0_; 
wire u6__0wb_data_o_31_0__0_; 
wire u6__0wb_data_o_31_0__10_; 
wire u6__0wb_data_o_31_0__11_; 
wire u6__0wb_data_o_31_0__12_; 
wire u6__0wb_data_o_31_0__13_; 
wire u6__0wb_data_o_31_0__14_; 
wire u6__0wb_data_o_31_0__15_; 
wire u6__0wb_data_o_31_0__16_; 
wire u6__0wb_data_o_31_0__17_; 
wire u6__0wb_data_o_31_0__18_; 
wire u6__0wb_data_o_31_0__19_; 
wire u6__0wb_data_o_31_0__1_; 
wire u6__0wb_data_o_31_0__20_; 
wire u6__0wb_data_o_31_0__21_; 
wire u6__0wb_data_o_31_0__22_; 
wire u6__0wb_data_o_31_0__23_; 
wire u6__0wb_data_o_31_0__24_; 
wire u6__0wb_data_o_31_0__25_; 
wire u6__0wb_data_o_31_0__26_; 
wire u6__0wb_data_o_31_0__27_; 
wire u6__0wb_data_o_31_0__28_; 
wire u6__0wb_data_o_31_0__29_; 
wire u6__0wb_data_o_31_0__2_; 
wire u6__0wb_data_o_31_0__30_; 
wire u6__0wb_data_o_31_0__31_; 
wire u6__0wb_data_o_31_0__3_; 
wire u6__0wb_data_o_31_0__4_; 
wire u6__0wb_data_o_31_0__5_; 
wire u6__0wb_data_o_31_0__6_; 
wire u6__0wb_data_o_31_0__7_; 
wire u6__0wb_data_o_31_0__8_; 
wire u6__0wb_data_o_31_0__9_; 
wire u6__0wb_err_0_0_; 
wire u6__0wb_first_r_0_0_; 
wire u6__0wr_hold_0_0_; 
wire u6__0write_go_r1_0_0_; 
wire u6__0write_go_r_0_0_; 
wire u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188; 
wire u6__abc_85257_new_n133_; 
wire u6__abc_85257_new_n134_; 
wire u6__abc_85257_new_n135_; 
wire u6__abc_85257_new_n136_; 
wire u6__abc_85257_new_n137_; 
wire u6__abc_85257_new_n138_; 
wire u6__abc_85257_new_n139_; 
wire u6__abc_85257_new_n140_; 
wire u6__abc_85257_new_n141_; 
wire u6__abc_85257_new_n142_; 
wire u6__abc_85257_new_n143_; 
wire u6__abc_85257_new_n144_; 
wire u6__abc_85257_new_n145_; 
wire u6__abc_85257_new_n145__bF_buf0; 
wire u6__abc_85257_new_n145__bF_buf1; 
wire u6__abc_85257_new_n145__bF_buf2; 
wire u6__abc_85257_new_n145__bF_buf3; 
wire u6__abc_85257_new_n145__bF_buf4; 
wire u6__abc_85257_new_n145__bF_buf5; 
wire u6__abc_85257_new_n146_; 
wire u6__abc_85257_new_n147_; 
wire u6__abc_85257_new_n148_; 
wire u6__abc_85257_new_n149_; 
wire u6__abc_85257_new_n150_; 
wire u6__abc_85257_new_n151_; 
wire u6__abc_85257_new_n152_; 
wire u6__abc_85257_new_n154_; 
wire u6__abc_85257_new_n155_; 
wire u6__abc_85257_new_n155__bF_buf0; 
wire u6__abc_85257_new_n155__bF_buf1; 
wire u6__abc_85257_new_n155__bF_buf2; 
wire u6__abc_85257_new_n155__bF_buf3; 
wire u6__abc_85257_new_n155__bF_buf4; 
wire u6__abc_85257_new_n156_; 
wire u6__abc_85257_new_n158_; 
wire u6__abc_85257_new_n159_; 
wire u6__abc_85257_new_n161_; 
wire u6__abc_85257_new_n162_; 
wire u6__abc_85257_new_n164_; 
wire u6__abc_85257_new_n165_; 
wire u6__abc_85257_new_n167_; 
wire u6__abc_85257_new_n168_; 
wire u6__abc_85257_new_n170_; 
wire u6__abc_85257_new_n171_; 
wire u6__abc_85257_new_n173_; 
wire u6__abc_85257_new_n174_; 
wire u6__abc_85257_new_n176_; 
wire u6__abc_85257_new_n177_; 
wire u6__abc_85257_new_n179_; 
wire u6__abc_85257_new_n180_; 
wire u6__abc_85257_new_n182_; 
wire u6__abc_85257_new_n183_; 
wire u6__abc_85257_new_n185_; 
wire u6__abc_85257_new_n186_; 
wire u6__abc_85257_new_n188_; 
wire u6__abc_85257_new_n189_; 
wire u6__abc_85257_new_n191_; 
wire u6__abc_85257_new_n192_; 
wire u6__abc_85257_new_n194_; 
wire u6__abc_85257_new_n195_; 
wire u6__abc_85257_new_n197_; 
wire u6__abc_85257_new_n198_; 
wire u6__abc_85257_new_n200_; 
wire u6__abc_85257_new_n201_; 
wire u6__abc_85257_new_n203_; 
wire u6__abc_85257_new_n204_; 
wire u6__abc_85257_new_n206_; 
wire u6__abc_85257_new_n207_; 
wire u6__abc_85257_new_n209_; 
wire u6__abc_85257_new_n210_; 
wire u6__abc_85257_new_n212_; 
wire u6__abc_85257_new_n213_; 
wire u6__abc_85257_new_n215_; 
wire u6__abc_85257_new_n216_; 
wire u6__abc_85257_new_n218_; 
wire u6__abc_85257_new_n219_; 
wire u6__abc_85257_new_n221_; 
wire u6__abc_85257_new_n222_; 
wire u6__abc_85257_new_n224_; 
wire u6__abc_85257_new_n225_; 
wire u6__abc_85257_new_n227_; 
wire u6__abc_85257_new_n228_; 
wire u6__abc_85257_new_n230_; 
wire u6__abc_85257_new_n231_; 
wire u6__abc_85257_new_n233_; 
wire u6__abc_85257_new_n234_; 
wire u6__abc_85257_new_n236_; 
wire u6__abc_85257_new_n237_; 
wire u6__abc_85257_new_n239_; 
wire u6__abc_85257_new_n240_; 
wire u6__abc_85257_new_n242_; 
wire u6__abc_85257_new_n243_; 
wire u6__abc_85257_new_n245_; 
wire u6__abc_85257_new_n246_; 
wire u6__abc_85257_new_n248_; 
wire u6__abc_85257_new_n249_; 
wire u6__abc_85257_new_n251_; 
wire u6__abc_85257_new_n252_; 
wire u6__abc_85257_new_n254_; 
wire u6__abc_85257_new_n255_; 
wire u6__abc_85257_new_n257_; 
wire u6__abc_85257_new_n258_; 
wire u6__abc_85257_new_n259_; 
wire u6__abc_85257_new_n260_; 
wire u6__abc_85257_new_n261_; 
wire u6__abc_85257_new_n262_; 
wire u6__abc_85257_new_n263_; 
wire u6__abc_85257_new_n264_; 
wire u6__abc_85257_new_n268_; 
wire u6__abc_85257_new_n269_; 
wire u6__abc_85257_new_n271_; 
wire u6__abc_85257_new_n272_; 
wire u6__abc_85257_new_n273_; 
wire u6__abc_85257_new_n276_; 
wire u6__abc_85257_new_n277_; 
wire u6__abc_85257_new_n278_; 
wire u6__abc_85257_new_n279_; 
wire u6__abc_85257_new_n280_; 
wire u6__abc_85257_new_n281_; 
wire u6__abc_85257_new_n282_; 
wire u6__abc_85257_new_n283_; 
wire u6__abc_85257_new_n285_; 
wire u6__abc_85257_new_n286_; 
wire u6__abc_85257_new_n288_; 
wire u6__abc_85257_new_n289_; 
wire u6__abc_85257_new_n291_; 
wire u6_read_go_r; 
wire u6_read_go_r1; 
wire u6_rmw_en; 
wire u6_rmw_r; 
wire u6_wb_first_r; 
wire u6_write_go_r; 
wire u6_write_go_r1; 
wire u7__0mc_adsc__0_0_; 
wire u7__0mc_adv__0_0_; 
wire u7__0mc_cs__0_0_; 
wire u7__0mc_cs__1_1_; 
wire u7__0mc_cs__2_2_; 
wire u7__0mc_cs__3_3_; 
wire u7__0mc_cs__4_4_; 
wire u7__0mc_cs__5_5_; 
wire u7__0mc_cs__6_6_; 
wire u7__0mc_cs__7_7_; 
wire u7__0mc_data_oe_0_0_; 
wire u7__0mc_dqm_3_0__0_; 
wire u7__0mc_dqm_3_0__1_; 
wire u7__0mc_dqm_3_0__2_; 
wire u7__0mc_dqm_3_0__3_; 
wire u7__0mc_dqm_r_3_0__0_; 
wire u7__0mc_dqm_r_3_0__1_; 
wire u7__0mc_dqm_r_3_0__2_; 
wire u7__0mc_dqm_r_3_0__3_; 
wire u7__0mc_oe__0_0_; 
wire u7__0mc_rp_0_0_; 
wire u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518; 
wire u7__abc_74830_new_n100_; 
wire u7__abc_74830_new_n101_; 
wire u7__abc_74830_new_n103_; 
wire u7__abc_74830_new_n104_; 
wire u7__abc_74830_new_n106_; 
wire u7__abc_74830_new_n107_; 
wire u7__abc_74830_new_n108_; 
wire u7__abc_74830_new_n109_; 
wire u7__abc_74830_new_n110_; 
wire u7__abc_74830_new_n111_; 
wire u7__abc_74830_new_n112_; 
wire u7__abc_74830_new_n113_; 
wire u7__abc_74830_new_n114_; 
wire u7__abc_74830_new_n115_; 
wire u7__abc_74830_new_n116_; 
wire u7__abc_74830_new_n117_; 
wire u7__abc_74830_new_n119_; 
wire u7__abc_74830_new_n120_; 
wire u7__abc_74830_new_n121_; 
wire u7__abc_74830_new_n122_; 
wire u7__abc_74830_new_n123_; 
wire u7__abc_74830_new_n124_; 
wire u7__abc_74830_new_n125_; 
wire u7__abc_74830_new_n126_; 
wire u7__abc_74830_new_n127_; 
wire u7__abc_74830_new_n129_; 
wire u7__abc_74830_new_n130_; 
wire u7__abc_74830_new_n131_; 
wire u7__abc_74830_new_n132_; 
wire u7__abc_74830_new_n133_; 
wire u7__abc_74830_new_n134_; 
wire u7__abc_74830_new_n135_; 
wire u7__abc_74830_new_n136_; 
wire u7__abc_74830_new_n137_; 
wire u7__abc_74830_new_n139_; 
wire u7__abc_74830_new_n140_; 
wire u7__abc_74830_new_n141_; 
wire u7__abc_74830_new_n142_; 
wire u7__abc_74830_new_n143_; 
wire u7__abc_74830_new_n144_; 
wire u7__abc_74830_new_n145_; 
wire u7__abc_74830_new_n146_; 
wire u7__abc_74830_new_n147_; 
wire u7__abc_74830_new_n149_; 
wire u7__abc_74830_new_n150_; 
wire u7__abc_74830_new_n151_; 
wire u7__abc_74830_new_n152_; 
wire u7__abc_74830_new_n153_; 
wire u7__abc_74830_new_n154_; 
wire u7__abc_74830_new_n155_; 
wire u7__abc_74830_new_n156_; 
wire u7__abc_74830_new_n157_; 
wire u7__abc_74830_new_n159_; 
wire u7__abc_74830_new_n160_; 
wire u7__abc_74830_new_n161_; 
wire u7__abc_74830_new_n162_; 
wire u7__abc_74830_new_n163_; 
wire u7__abc_74830_new_n164_; 
wire u7__abc_74830_new_n165_; 
wire u7__abc_74830_new_n166_; 
wire u7__abc_74830_new_n167_; 
wire u7__abc_74830_new_n169_; 
wire u7__abc_74830_new_n170_; 
wire u7__abc_74830_new_n171_; 
wire u7__abc_74830_new_n172_; 
wire u7__abc_74830_new_n173_; 
wire u7__abc_74830_new_n174_; 
wire u7__abc_74830_new_n175_; 
wire u7__abc_74830_new_n176_; 
wire u7__abc_74830_new_n177_; 
wire u7__abc_74830_new_n179_; 
wire u7__abc_74830_new_n180_; 
wire u7__abc_74830_new_n181_; 
wire u7__abc_74830_new_n182_; 
wire u7__abc_74830_new_n183_; 
wire u7__abc_74830_new_n184_; 
wire u7__abc_74830_new_n185_; 
wire u7__abc_74830_new_n186_; 
wire u7__abc_74830_new_n187_; 
wire u7__abc_74830_new_n191_; 
wire u7__abc_74830_new_n192_; 
wire u7__abc_74830_new_n194_; 
wire u7__abc_74830_new_n195_; 
wire u7__abc_74830_new_n75_; 
wire u7__abc_74830_new_n76_; 
wire u7__abc_74830_new_n77_; 
wire u7__abc_74830_new_n78_; 
wire u7__abc_74830_new_n79_; 
wire u7__abc_74830_new_n80_; 
wire u7__abc_74830_new_n81_; 
wire u7__abc_74830_new_n83_; 
wire u7__abc_74830_new_n84_; 
wire u7__abc_74830_new_n86_; 
wire u7__abc_74830_new_n87_; 
wire u7__abc_74830_new_n89_; 
wire u7__abc_74830_new_n90_; 
wire u7__abc_74830_new_n92_; 
wire u7__abc_74830_new_n93_; 
wire u7__abc_74830_new_n94_; 
wire u7__abc_74830_new_n95_; 
wire u7__abc_74830_new_n97_; 
wire u7__abc_74830_new_n98_; 
wire u7_mc_dqm_r2_0_; 
wire u7_mc_dqm_r2_1_; 
wire u7_mc_dqm_r2_2_; 
wire u7_mc_dqm_r2_3_; 
wire u7_mc_dqm_r_0_; 
wire u7_mc_dqm_r_1_; 
wire u7_mc_dqm_r_2_; 
wire u7_mc_dqm_r_3_; 
output wb_ack_o;
input \wb_addr_i[0] ;
input \wb_addr_i[10] ;
input \wb_addr_i[11] ;
input \wb_addr_i[12] ;
input \wb_addr_i[13] ;
input \wb_addr_i[14] ;
input \wb_addr_i[15] ;
input \wb_addr_i[16] ;
input \wb_addr_i[17] ;
input \wb_addr_i[18] ;
input \wb_addr_i[19] ;
input \wb_addr_i[1] ;
input \wb_addr_i[20] ;
input \wb_addr_i[21] ;
input \wb_addr_i[22] ;
input \wb_addr_i[23] ;
input \wb_addr_i[24] ;
input \wb_addr_i[25] ;
input \wb_addr_i[26] ;
input \wb_addr_i[27] ;
input \wb_addr_i[28] ;
input \wb_addr_i[29] ;
input \wb_addr_i[2] ;
input \wb_addr_i[30] ;
input \wb_addr_i[31] ;
input \wb_addr_i[3] ;
input \wb_addr_i[4] ;
input \wb_addr_i[5] ;
input \wb_addr_i[6] ;
input \wb_addr_i[7] ;
input \wb_addr_i[8] ;
input \wb_addr_i[9] ;
input wb_cyc_i;
input \wb_data_i[0] ;
input \wb_data_i[10] ;
input \wb_data_i[11] ;
input \wb_data_i[12] ;
input \wb_data_i[13] ;
input \wb_data_i[14] ;
input \wb_data_i[15] ;
input \wb_data_i[16] ;
input \wb_data_i[17] ;
input \wb_data_i[18] ;
input \wb_data_i[19] ;
input \wb_data_i[1] ;
input \wb_data_i[20] ;
input \wb_data_i[21] ;
input \wb_data_i[22] ;
input \wb_data_i[23] ;
input \wb_data_i[24] ;
input \wb_data_i[25] ;
input \wb_data_i[26] ;
input \wb_data_i[27] ;
input \wb_data_i[28] ;
input \wb_data_i[29] ;
input \wb_data_i[2] ;
input \wb_data_i[30] ;
input \wb_data_i[31] ;
input \wb_data_i[3] ;
input \wb_data_i[4] ;
input \wb_data_i[5] ;
input \wb_data_i[6] ;
input \wb_data_i[7] ;
input \wb_data_i[8] ;
input \wb_data_i[9] ;
output \wb_data_o[0] ;
output \wb_data_o[10] ;
output \wb_data_o[11] ;
output \wb_data_o[12] ;
output \wb_data_o[13] ;
output \wb_data_o[14] ;
output \wb_data_o[15] ;
output \wb_data_o[16] ;
output \wb_data_o[17] ;
output \wb_data_o[18] ;
output \wb_data_o[19] ;
output \wb_data_o[1] ;
output \wb_data_o[20] ;
output \wb_data_o[21] ;
output \wb_data_o[22] ;
output \wb_data_o[23] ;
output \wb_data_o[24] ;
output \wb_data_o[25] ;
output \wb_data_o[26] ;
output \wb_data_o[27] ;
output \wb_data_o[28] ;
output \wb_data_o[29] ;
output \wb_data_o[2] ;
output \wb_data_o[30] ;
output \wb_data_o[31] ;
output \wb_data_o[3] ;
output \wb_data_o[4] ;
output \wb_data_o[5] ;
output \wb_data_o[6] ;
output \wb_data_o[7] ;
output \wb_data_o[8] ;
output \wb_data_o[9] ;
output wb_err_o;
input \wb_sel_i[0] ;
input \wb_sel_i[1] ;
input \wb_sel_i[2] ;
input \wb_sel_i[3] ;
input wb_stb_i;
wire wb_stb_i_bF_buf0; 
wire wb_stb_i_bF_buf1; 
wire wb_stb_i_bF_buf2; 
wire wb_stb_i_bF_buf3; 
wire wb_stb_i_bF_buf4; 
wire wb_stb_i_bF_buf5; 
input wb_we_i;
AND2X2 AND2X2_1 ( .A(_abc_85006_new_n238_), .B(_abc_85006_new_n239_), .Y(_abc_85006_new_n240_));
AND2X2 AND2X2_10 ( .A(_abc_85006_new_n266_), .B(_abc_85006_new_n267_), .Y(_abc_85006_new_n268_));
AND2X2 AND2X2_100 ( .A(spec_req_cs_5_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1176_));
AND2X2 AND2X2_1000 ( .A(u0__abc_76628_new_n3377_), .B(u0__abc_76628_new_n2720__bF_buf2), .Y(u0__abc_76628_new_n3378_));
AND2X2 AND2X2_1001 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3379_));
AND2X2 AND2X2_1002 ( .A(u0__abc_76628_new_n3380_), .B(u0__abc_76628_new_n2719__bF_buf2), .Y(u0__abc_76628_new_n3381_));
AND2X2 AND2X2_1003 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3382_));
AND2X2 AND2X2_1004 ( .A(u0__abc_76628_new_n3383_), .B(u0__abc_76628_new_n2718__bF_buf2), .Y(u0__abc_76628_new_n3384_));
AND2X2 AND2X2_1005 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3385_));
AND2X2 AND2X2_1006 ( .A(u0__abc_76628_new_n3386_), .B(u0__abc_76628_new_n2717__bF_buf2), .Y(u0__abc_76628_new_n3387_));
AND2X2 AND2X2_1007 ( .A(u0_tms1_27_), .B(u0_cs1_bF_buf1), .Y(u0__abc_76628_new_n3388_));
AND2X2 AND2X2_1008 ( .A(u0__abc_76628_new_n1169__bF_buf6), .B(u0__abc_76628_new_n3391_), .Y(u0__abc_76628_new_n3392_));
AND2X2 AND2X2_1009 ( .A(u0__abc_76628_new_n3390_), .B(u0__abc_76628_new_n3392_), .Y(u0__abc_76628_new_n3393_));
AND2X2 AND2X2_101 ( .A(u0__abc_76628_new_n1180_), .B(u0__abc_76628_new_n1179__bF_buf5), .Y(u0__abc_76628_new_n1181_));
AND2X2 AND2X2_1010 ( .A(u0__abc_76628_new_n1947__bF_buf2), .B(csc_1_), .Y(u0__abc_76628_new_n3515_));
AND2X2 AND2X2_1011 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3516_));
AND2X2 AND2X2_1012 ( .A(u0__abc_76628_new_n3518_), .B(u0__abc_76628_new_n2724__bF_buf1), .Y(u0__abc_76628_new_n3519_));
AND2X2 AND2X2_1013 ( .A(u0__abc_76628_new_n3519_), .B(u0__abc_76628_new_n3517_), .Y(u0__abc_76628_new_n3520_));
AND2X2 AND2X2_1014 ( .A(u0__abc_76628_new_n3521_), .B(u0__abc_76628_new_n2720__bF_buf1), .Y(u0__abc_76628_new_n3522_));
AND2X2 AND2X2_1015 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3523_));
AND2X2 AND2X2_1016 ( .A(u0__abc_76628_new_n3524_), .B(u0__abc_76628_new_n2719__bF_buf1), .Y(u0__abc_76628_new_n3525_));
AND2X2 AND2X2_1017 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3526_));
AND2X2 AND2X2_1018 ( .A(u0__abc_76628_new_n3527_), .B(u0__abc_76628_new_n2718__bF_buf1), .Y(u0__abc_76628_new_n3528_));
AND2X2 AND2X2_1019 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3529_));
AND2X2 AND2X2_102 ( .A(u0__abc_76628_new_n1181_), .B(u0__abc_76628_new_n1178_), .Y(u0__abc_76628_new_n1182_));
AND2X2 AND2X2_1020 ( .A(u0__abc_76628_new_n3530_), .B(u0__abc_76628_new_n2717__bF_buf1), .Y(u0__abc_76628_new_n3531_));
AND2X2 AND2X2_1021 ( .A(u0_csc1_1_), .B(u0_cs1_bF_buf0), .Y(u0__abc_76628_new_n3532_));
AND2X2 AND2X2_1022 ( .A(u0__abc_76628_new_n1946__bF_buf1), .B(u0__abc_76628_new_n3535_), .Y(u0__abc_76628_new_n3536_));
AND2X2 AND2X2_1023 ( .A(u0__abc_76628_new_n3534_), .B(u0__abc_76628_new_n3536_), .Y(u0__abc_76628_new_n3537_));
AND2X2 AND2X2_1024 ( .A(u0__abc_76628_new_n1947__bF_buf1), .B(csc_2_), .Y(u0__abc_76628_new_n3539_));
AND2X2 AND2X2_1025 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3540_));
AND2X2 AND2X2_1026 ( .A(u0__abc_76628_new_n3542_), .B(u0__abc_76628_new_n2724__bF_buf0), .Y(u0__abc_76628_new_n3543_));
AND2X2 AND2X2_1027 ( .A(u0__abc_76628_new_n3543_), .B(u0__abc_76628_new_n3541_), .Y(u0__abc_76628_new_n3544_));
AND2X2 AND2X2_1028 ( .A(u0__abc_76628_new_n3545_), .B(u0__abc_76628_new_n2720__bF_buf0), .Y(u0__abc_76628_new_n3546_));
AND2X2 AND2X2_1029 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3547_));
AND2X2 AND2X2_103 ( .A(u0__abc_76628_new_n1183_), .B(u0__abc_76628_new_n1175__bF_buf5), .Y(u0__abc_76628_new_n1184_));
AND2X2 AND2X2_1030 ( .A(u0__abc_76628_new_n3548_), .B(u0__abc_76628_new_n2719__bF_buf0), .Y(u0__abc_76628_new_n3549_));
AND2X2 AND2X2_1031 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3550_));
AND2X2 AND2X2_1032 ( .A(u0__abc_76628_new_n3551_), .B(u0__abc_76628_new_n2718__bF_buf0), .Y(u0__abc_76628_new_n3552_));
AND2X2 AND2X2_1033 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3553_));
AND2X2 AND2X2_1034 ( .A(u0__abc_76628_new_n3554_), .B(u0__abc_76628_new_n2717__bF_buf0), .Y(u0__abc_76628_new_n3555_));
AND2X2 AND2X2_1035 ( .A(u0_csc1_2_), .B(u0_cs1_bF_buf5), .Y(u0__abc_76628_new_n3556_));
AND2X2 AND2X2_1036 ( .A(u0__abc_76628_new_n1946__bF_buf0), .B(u0__abc_76628_new_n3559_), .Y(u0__abc_76628_new_n3560_));
AND2X2 AND2X2_1037 ( .A(u0__abc_76628_new_n3558_), .B(u0__abc_76628_new_n3560_), .Y(u0__abc_76628_new_n3561_));
AND2X2 AND2X2_1038 ( .A(u0__abc_76628_new_n1947__bF_buf0), .B(csc_3_), .Y(u0__abc_76628_new_n3563_));
AND2X2 AND2X2_1039 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3564_));
AND2X2 AND2X2_104 ( .A(spec_req_cs_4_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1185_));
AND2X2 AND2X2_1040 ( .A(u0__abc_76628_new_n3566_), .B(u0__abc_76628_new_n2724__bF_buf5), .Y(u0__abc_76628_new_n3567_));
AND2X2 AND2X2_1041 ( .A(u0__abc_76628_new_n3567_), .B(u0__abc_76628_new_n3565_), .Y(u0__abc_76628_new_n3568_));
AND2X2 AND2X2_1042 ( .A(u0__abc_76628_new_n3569_), .B(u0__abc_76628_new_n2720__bF_buf5), .Y(u0__abc_76628_new_n3570_));
AND2X2 AND2X2_1043 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3571_));
AND2X2 AND2X2_1044 ( .A(u0__abc_76628_new_n3572_), .B(u0__abc_76628_new_n2719__bF_buf5), .Y(u0__abc_76628_new_n3573_));
AND2X2 AND2X2_1045 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3574_));
AND2X2 AND2X2_1046 ( .A(u0__abc_76628_new_n3575_), .B(u0__abc_76628_new_n2718__bF_buf5), .Y(u0__abc_76628_new_n3576_));
AND2X2 AND2X2_1047 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3577_));
AND2X2 AND2X2_1048 ( .A(u0__abc_76628_new_n3578_), .B(u0__abc_76628_new_n2717__bF_buf5), .Y(u0__abc_76628_new_n3579_));
AND2X2 AND2X2_1049 ( .A(u0_csc1_3_), .B(u0_cs1_bF_buf4), .Y(u0__abc_76628_new_n3580_));
AND2X2 AND2X2_105 ( .A(u0__abc_76628_new_n1186_), .B(u0__abc_76628_new_n1174__bF_buf5), .Y(u0__abc_76628_new_n1187_));
AND2X2 AND2X2_1050 ( .A(u0__abc_76628_new_n1946__bF_buf3), .B(u0__abc_76628_new_n3583_), .Y(u0__abc_76628_new_n3584_));
AND2X2 AND2X2_1051 ( .A(u0__abc_76628_new_n3582_), .B(u0__abc_76628_new_n3584_), .Y(u0__abc_76628_new_n3585_));
AND2X2 AND2X2_1052 ( .A(u0__abc_76628_new_n1947__bF_buf3), .B(csc_4_), .Y(u0__abc_76628_new_n3587_));
AND2X2 AND2X2_1053 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3588_));
AND2X2 AND2X2_1054 ( .A(u0__abc_76628_new_n3590_), .B(u0__abc_76628_new_n2724__bF_buf4), .Y(u0__abc_76628_new_n3591_));
AND2X2 AND2X2_1055 ( .A(u0__abc_76628_new_n3591_), .B(u0__abc_76628_new_n3589_), .Y(u0__abc_76628_new_n3592_));
AND2X2 AND2X2_1056 ( .A(u0__abc_76628_new_n3593_), .B(u0__abc_76628_new_n2720__bF_buf4), .Y(u0__abc_76628_new_n3594_));
AND2X2 AND2X2_1057 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3595_));
AND2X2 AND2X2_1058 ( .A(u0__abc_76628_new_n3596_), .B(u0__abc_76628_new_n2719__bF_buf4), .Y(u0__abc_76628_new_n3597_));
AND2X2 AND2X2_1059 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3598_));
AND2X2 AND2X2_106 ( .A(spec_req_cs_3_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1188_));
AND2X2 AND2X2_1060 ( .A(u0__abc_76628_new_n3599_), .B(u0__abc_76628_new_n2718__bF_buf4), .Y(u0__abc_76628_new_n3600_));
AND2X2 AND2X2_1061 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3601_));
AND2X2 AND2X2_1062 ( .A(u0__abc_76628_new_n3602_), .B(u0__abc_76628_new_n2717__bF_buf4), .Y(u0__abc_76628_new_n3603_));
AND2X2 AND2X2_1063 ( .A(u0_csc1_4_), .B(u0_cs1_bF_buf3), .Y(u0__abc_76628_new_n3604_));
AND2X2 AND2X2_1064 ( .A(u0__abc_76628_new_n1946__bF_buf2), .B(u0__abc_76628_new_n3607_), .Y(u0__abc_76628_new_n3608_));
AND2X2 AND2X2_1065 ( .A(u0__abc_76628_new_n3606_), .B(u0__abc_76628_new_n3608_), .Y(u0__abc_76628_new_n3609_));
AND2X2 AND2X2_1066 ( .A(u0__abc_76628_new_n1947__bF_buf2), .B(csc_5_bF_buf3_), .Y(u0__abc_76628_new_n3611_));
AND2X2 AND2X2_1067 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3612_));
AND2X2 AND2X2_1068 ( .A(u0__abc_76628_new_n3614_), .B(u0__abc_76628_new_n2724__bF_buf3), .Y(u0__abc_76628_new_n3615_));
AND2X2 AND2X2_1069 ( .A(u0__abc_76628_new_n3615_), .B(u0__abc_76628_new_n3613_), .Y(u0__abc_76628_new_n3616_));
AND2X2 AND2X2_107 ( .A(u0__abc_76628_new_n1189_), .B(u0__abc_76628_new_n1173__bF_buf5), .Y(u0__abc_76628_new_n1190_));
AND2X2 AND2X2_1070 ( .A(u0__abc_76628_new_n3617_), .B(u0__abc_76628_new_n2720__bF_buf3), .Y(u0__abc_76628_new_n3618_));
AND2X2 AND2X2_1071 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3619_));
AND2X2 AND2X2_1072 ( .A(u0__abc_76628_new_n3620_), .B(u0__abc_76628_new_n2719__bF_buf3), .Y(u0__abc_76628_new_n3621_));
AND2X2 AND2X2_1073 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3622_));
AND2X2 AND2X2_1074 ( .A(u0__abc_76628_new_n3623_), .B(u0__abc_76628_new_n2718__bF_buf3), .Y(u0__abc_76628_new_n3624_));
AND2X2 AND2X2_1075 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3625_));
AND2X2 AND2X2_1076 ( .A(u0__abc_76628_new_n3626_), .B(u0__abc_76628_new_n2717__bF_buf3), .Y(u0__abc_76628_new_n3627_));
AND2X2 AND2X2_1077 ( .A(u0_csc1_5_), .B(u0_cs1_bF_buf2), .Y(u0__abc_76628_new_n3628_));
AND2X2 AND2X2_1078 ( .A(u0__abc_76628_new_n1946__bF_buf1), .B(u0__abc_76628_new_n3631_), .Y(u0__abc_76628_new_n3632_));
AND2X2 AND2X2_1079 ( .A(u0__abc_76628_new_n3630_), .B(u0__abc_76628_new_n3632_), .Y(u0__abc_76628_new_n3633_));
AND2X2 AND2X2_108 ( .A(spec_req_cs_2_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1191_));
AND2X2 AND2X2_1080 ( .A(u0__abc_76628_new_n1947__bF_buf1), .B(csc_6_), .Y(u0__abc_76628_new_n3635_));
AND2X2 AND2X2_1081 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3636_));
AND2X2 AND2X2_1082 ( .A(u0__abc_76628_new_n3638_), .B(u0__abc_76628_new_n2724__bF_buf2), .Y(u0__abc_76628_new_n3639_));
AND2X2 AND2X2_1083 ( .A(u0__abc_76628_new_n3639_), .B(u0__abc_76628_new_n3637_), .Y(u0__abc_76628_new_n3640_));
AND2X2 AND2X2_1084 ( .A(u0__abc_76628_new_n3641_), .B(u0__abc_76628_new_n2720__bF_buf2), .Y(u0__abc_76628_new_n3642_));
AND2X2 AND2X2_1085 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3643_));
AND2X2 AND2X2_1086 ( .A(u0__abc_76628_new_n3644_), .B(u0__abc_76628_new_n2719__bF_buf2), .Y(u0__abc_76628_new_n3645_));
AND2X2 AND2X2_1087 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3646_));
AND2X2 AND2X2_1088 ( .A(u0__abc_76628_new_n3647_), .B(u0__abc_76628_new_n2718__bF_buf2), .Y(u0__abc_76628_new_n3648_));
AND2X2 AND2X2_1089 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3649_));
AND2X2 AND2X2_109 ( .A(u0__abc_76628_new_n1192_), .B(u0__abc_76628_new_n1172__bF_buf5), .Y(u0__abc_76628_new_n1193_));
AND2X2 AND2X2_1090 ( .A(u0__abc_76628_new_n3650_), .B(u0__abc_76628_new_n2717__bF_buf2), .Y(u0__abc_76628_new_n3651_));
AND2X2 AND2X2_1091 ( .A(u0_csc1_6_), .B(u0_cs1_bF_buf1), .Y(u0__abc_76628_new_n3652_));
AND2X2 AND2X2_1092 ( .A(u0__abc_76628_new_n1946__bF_buf0), .B(u0__abc_76628_new_n3655_), .Y(u0__abc_76628_new_n3656_));
AND2X2 AND2X2_1093 ( .A(u0__abc_76628_new_n3654_), .B(u0__abc_76628_new_n3656_), .Y(u0__abc_76628_new_n3657_));
AND2X2 AND2X2_1094 ( .A(u0__abc_76628_new_n1947__bF_buf0), .B(csc_7_), .Y(u0__abc_76628_new_n3659_));
AND2X2 AND2X2_1095 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3660_));
AND2X2 AND2X2_1096 ( .A(u0__abc_76628_new_n3662_), .B(u0__abc_76628_new_n2724__bF_buf1), .Y(u0__abc_76628_new_n3663_));
AND2X2 AND2X2_1097 ( .A(u0__abc_76628_new_n3663_), .B(u0__abc_76628_new_n3661_), .Y(u0__abc_76628_new_n3664_));
AND2X2 AND2X2_1098 ( .A(u0__abc_76628_new_n3665_), .B(u0__abc_76628_new_n2720__bF_buf1), .Y(u0__abc_76628_new_n3666_));
AND2X2 AND2X2_1099 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3667_));
AND2X2 AND2X2_11 ( .A(_abc_85006_new_n269_), .B(_abc_85006_new_n270_), .Y(obct_cs_4_));
AND2X2 AND2X2_110 ( .A(spec_req_cs_1_bF_buf2_), .B(u0_tms1_0_), .Y(u0__abc_76628_new_n1194_));
AND2X2 AND2X2_1100 ( .A(u0__abc_76628_new_n3668_), .B(u0__abc_76628_new_n2719__bF_buf1), .Y(u0__abc_76628_new_n3669_));
AND2X2 AND2X2_1101 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3670_));
AND2X2 AND2X2_1102 ( .A(u0__abc_76628_new_n3671_), .B(u0__abc_76628_new_n2718__bF_buf1), .Y(u0__abc_76628_new_n3672_));
AND2X2 AND2X2_1103 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3673_));
AND2X2 AND2X2_1104 ( .A(u0__abc_76628_new_n3674_), .B(u0__abc_76628_new_n2717__bF_buf1), .Y(u0__abc_76628_new_n3675_));
AND2X2 AND2X2_1105 ( .A(u0_csc1_7_), .B(u0_cs1_bF_buf0), .Y(u0__abc_76628_new_n3676_));
AND2X2 AND2X2_1106 ( .A(u0__abc_76628_new_n1946__bF_buf3), .B(u0__abc_76628_new_n3679_), .Y(u0__abc_76628_new_n3680_));
AND2X2 AND2X2_1107 ( .A(u0__abc_76628_new_n3678_), .B(u0__abc_76628_new_n3680_), .Y(u0__abc_76628_new_n3681_));
AND2X2 AND2X2_1108 ( .A(u0__abc_76628_new_n1947__bF_buf3), .B(csc_9_), .Y(u0__abc_76628_new_n3707_));
AND2X2 AND2X2_1109 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3708_));
AND2X2 AND2X2_111 ( .A(u0__abc_76628_new_n1169__bF_buf5), .B(u0__abc_76628_new_n1198_), .Y(u0__abc_76628_new_n1199_));
AND2X2 AND2X2_1110 ( .A(u0__abc_76628_new_n3710_), .B(u0__abc_76628_new_n2724__bF_buf0), .Y(u0__abc_76628_new_n3711_));
AND2X2 AND2X2_1111 ( .A(u0__abc_76628_new_n3711_), .B(u0__abc_76628_new_n3709_), .Y(u0__abc_76628_new_n3712_));
AND2X2 AND2X2_1112 ( .A(u0__abc_76628_new_n3713_), .B(u0__abc_76628_new_n2720__bF_buf0), .Y(u0__abc_76628_new_n3714_));
AND2X2 AND2X2_1113 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3715_));
AND2X2 AND2X2_1114 ( .A(u0__abc_76628_new_n3716_), .B(u0__abc_76628_new_n2719__bF_buf0), .Y(u0__abc_76628_new_n3717_));
AND2X2 AND2X2_1115 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3718_));
AND2X2 AND2X2_1116 ( .A(u0__abc_76628_new_n3719_), .B(u0__abc_76628_new_n2718__bF_buf0), .Y(u0__abc_76628_new_n3720_));
AND2X2 AND2X2_1117 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3721_));
AND2X2 AND2X2_1118 ( .A(u0__abc_76628_new_n3722_), .B(u0__abc_76628_new_n2717__bF_buf0), .Y(u0__abc_76628_new_n3723_));
AND2X2 AND2X2_1119 ( .A(u0_csc1_9_), .B(u0_cs1_bF_buf5), .Y(u0__abc_76628_new_n3724_));
AND2X2 AND2X2_112 ( .A(u0__abc_76628_new_n1196_), .B(u0__abc_76628_new_n1199_), .Y(u0__abc_76628_new_n1200_));
AND2X2 AND2X2_1120 ( .A(u0__abc_76628_new_n1946__bF_buf2), .B(u0__abc_76628_new_n3727_), .Y(u0__abc_76628_new_n3728_));
AND2X2 AND2X2_1121 ( .A(u0__abc_76628_new_n3726_), .B(u0__abc_76628_new_n3728_), .Y(u0__abc_76628_new_n3729_));
AND2X2 AND2X2_1122 ( .A(u0__abc_76628_new_n1947__bF_buf2), .B(csc_10_), .Y(u0__abc_76628_new_n3731_));
AND2X2 AND2X2_1123 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3732_));
AND2X2 AND2X2_1124 ( .A(u0__abc_76628_new_n3734_), .B(u0__abc_76628_new_n2724__bF_buf5), .Y(u0__abc_76628_new_n3735_));
AND2X2 AND2X2_1125 ( .A(u0__abc_76628_new_n3735_), .B(u0__abc_76628_new_n3733_), .Y(u0__abc_76628_new_n3736_));
AND2X2 AND2X2_1126 ( .A(u0__abc_76628_new_n3737_), .B(u0__abc_76628_new_n2720__bF_buf5), .Y(u0__abc_76628_new_n3738_));
AND2X2 AND2X2_1127 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3739_));
AND2X2 AND2X2_1128 ( .A(u0__abc_76628_new_n3740_), .B(u0__abc_76628_new_n2719__bF_buf5), .Y(u0__abc_76628_new_n3741_));
AND2X2 AND2X2_1129 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3742_));
AND2X2 AND2X2_113 ( .A(u0__abc_76628_new_n1170__bF_buf5), .B(sp_tms_1_), .Y(u0__abc_76628_new_n1202_));
AND2X2 AND2X2_1130 ( .A(u0__abc_76628_new_n3743_), .B(u0__abc_76628_new_n2718__bF_buf5), .Y(u0__abc_76628_new_n3744_));
AND2X2 AND2X2_1131 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3745_));
AND2X2 AND2X2_1132 ( .A(u0__abc_76628_new_n3746_), .B(u0__abc_76628_new_n2717__bF_buf5), .Y(u0__abc_76628_new_n3747_));
AND2X2 AND2X2_1133 ( .A(u0_csc1_10_), .B(u0_cs1_bF_buf4), .Y(u0__abc_76628_new_n3748_));
AND2X2 AND2X2_1134 ( .A(u0__abc_76628_new_n1946__bF_buf1), .B(u0__abc_76628_new_n3751_), .Y(u0__abc_76628_new_n3752_));
AND2X2 AND2X2_1135 ( .A(u0__abc_76628_new_n3750_), .B(u0__abc_76628_new_n3752_), .Y(u0__abc_76628_new_n3753_));
AND2X2 AND2X2_1136 ( .A(u0__abc_76628_new_n1947__bF_buf1), .B(u3_pen), .Y(u0__abc_76628_new_n3755_));
AND2X2 AND2X2_1137 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3756_));
AND2X2 AND2X2_1138 ( .A(u0__abc_76628_new_n3758_), .B(u0__abc_76628_new_n2724__bF_buf4), .Y(u0__abc_76628_new_n3759_));
AND2X2 AND2X2_1139 ( .A(u0__abc_76628_new_n3759_), .B(u0__abc_76628_new_n3757_), .Y(u0__abc_76628_new_n3760_));
AND2X2 AND2X2_114 ( .A(spec_req_cs_5_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1203_));
AND2X2 AND2X2_1140 ( .A(u0__abc_76628_new_n3761_), .B(u0__abc_76628_new_n2720__bF_buf4), .Y(u0__abc_76628_new_n3762_));
AND2X2 AND2X2_1141 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3763_));
AND2X2 AND2X2_1142 ( .A(u0__abc_76628_new_n3764_), .B(u0__abc_76628_new_n2719__bF_buf4), .Y(u0__abc_76628_new_n3765_));
AND2X2 AND2X2_1143 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3766_));
AND2X2 AND2X2_1144 ( .A(u0__abc_76628_new_n3767_), .B(u0__abc_76628_new_n2718__bF_buf4), .Y(u0__abc_76628_new_n3768_));
AND2X2 AND2X2_1145 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3769_));
AND2X2 AND2X2_1146 ( .A(u0__abc_76628_new_n3770_), .B(u0__abc_76628_new_n2717__bF_buf4), .Y(u0__abc_76628_new_n3771_));
AND2X2 AND2X2_1147 ( .A(u0_csc1_11_), .B(u0_cs1_bF_buf3), .Y(u0__abc_76628_new_n3772_));
AND2X2 AND2X2_1148 ( .A(u0__abc_76628_new_n1946__bF_buf0), .B(u0__abc_76628_new_n3775_), .Y(u0__abc_76628_new_n3776_));
AND2X2 AND2X2_1149 ( .A(u0__abc_76628_new_n3774_), .B(u0__abc_76628_new_n3776_), .Y(u0__abc_76628_new_n3777_));
AND2X2 AND2X2_115 ( .A(u0__abc_76628_new_n1205_), .B(u0__abc_76628_new_n1179__bF_buf4), .Y(u0__abc_76628_new_n1206_));
AND2X2 AND2X2_1150 ( .A(u0__abc_76628_new_n1168_), .B(cs_le_bF_buf4), .Y(u0__abc_76628_new_n4259_));
AND2X2 AND2X2_1151 ( .A(u0__abc_76628_new_n4266_), .B(u0__abc_76628_new_n4259_), .Y(u0__abc_76628_new_n4267_));
AND2X2 AND2X2_1152 ( .A(wb_cyc_i), .B(u0_wp_err), .Y(u0__abc_76628_new_n4269_));
AND2X2 AND2X2_1153 ( .A(u0__abc_76628_new_n4268_), .B(u0__abc_76628_new_n4269_), .Y(u0__abc_76628_new_n4270_));
AND2X2 AND2X2_1154 ( .A(u0__abc_76628_new_n4274_), .B(u0__abc_76628_new_n4272_), .Y(u0__0cs_7_0__0_));
AND2X2 AND2X2_1155 ( .A(u0__abc_76628_new_n4277_), .B(u0__abc_76628_new_n4276_), .Y(u0__0cs_7_0__1_));
AND2X2 AND2X2_1156 ( .A(u0__abc_76628_new_n4280_), .B(u0__abc_76628_new_n4279_), .Y(u0__0cs_7_0__2_));
AND2X2 AND2X2_1157 ( .A(u0__abc_76628_new_n4283_), .B(u0__abc_76628_new_n4282_), .Y(u0__0cs_7_0__3_));
AND2X2 AND2X2_1158 ( .A(u0__abc_76628_new_n4286_), .B(u0__abc_76628_new_n4285_), .Y(u0__0cs_7_0__4_));
AND2X2 AND2X2_1159 ( .A(u0__abc_76628_new_n4289_), .B(u0__abc_76628_new_n4288_), .Y(u0__0cs_7_0__5_));
AND2X2 AND2X2_116 ( .A(u0__abc_76628_new_n1206_), .B(u0__abc_76628_new_n1204_), .Y(u0__abc_76628_new_n1207_));
AND2X2 AND2X2_1160 ( .A(u0__abc_76628_new_n4292_), .B(u0__abc_76628_new_n4291_), .Y(u0__0cs_7_0__6_));
AND2X2 AND2X2_1161 ( .A(u0__abc_76628_new_n4295_), .B(u0__abc_76628_new_n4294_), .Y(u0__0cs_7_0__7_));
AND2X2 AND2X2_1162 ( .A(u0__abc_76628_new_n4299_), .B(u0__abc_76628_new_n4297_), .Y(u0__0poc_31_0__0_));
AND2X2 AND2X2_1163 ( .A(u0__abc_76628_new_n4302_), .B(u0__abc_76628_new_n4301_), .Y(u0__0poc_31_0__1_));
AND2X2 AND2X2_1164 ( .A(u0__abc_76628_new_n4305_), .B(u0__abc_76628_new_n4304_), .Y(u0__0poc_31_0__2_));
AND2X2 AND2X2_1165 ( .A(u0__abc_76628_new_n4308_), .B(u0__abc_76628_new_n4307_), .Y(u0__0poc_31_0__3_));
AND2X2 AND2X2_1166 ( .A(u0__abc_76628_new_n4311_), .B(u0__abc_76628_new_n4310_), .Y(u0__0poc_31_0__4_));
AND2X2 AND2X2_1167 ( .A(u0__abc_76628_new_n4314_), .B(u0__abc_76628_new_n4313_), .Y(u0__0poc_31_0__5_));
AND2X2 AND2X2_1168 ( .A(u0__abc_76628_new_n4317_), .B(u0__abc_76628_new_n4316_), .Y(u0__0poc_31_0__6_));
AND2X2 AND2X2_1169 ( .A(u0__abc_76628_new_n4320_), .B(u0__abc_76628_new_n4319_), .Y(u0__0poc_31_0__7_));
AND2X2 AND2X2_117 ( .A(u0__abc_76628_new_n1208_), .B(u0__abc_76628_new_n1175__bF_buf4), .Y(u0__abc_76628_new_n1209_));
AND2X2 AND2X2_1170 ( .A(u0__abc_76628_new_n4323_), .B(u0__abc_76628_new_n4322_), .Y(u0__0poc_31_0__8_));
AND2X2 AND2X2_1171 ( .A(u0__abc_76628_new_n4326_), .B(u0__abc_76628_new_n4325_), .Y(u0__0poc_31_0__9_));
AND2X2 AND2X2_1172 ( .A(u0__abc_76628_new_n4329_), .B(u0__abc_76628_new_n4328_), .Y(u0__0poc_31_0__10_));
AND2X2 AND2X2_1173 ( .A(u0__abc_76628_new_n4332_), .B(u0__abc_76628_new_n4331_), .Y(u0__0poc_31_0__11_));
AND2X2 AND2X2_1174 ( .A(u0__abc_76628_new_n4335_), .B(u0__abc_76628_new_n4334_), .Y(u0__0poc_31_0__12_));
AND2X2 AND2X2_1175 ( .A(u0__abc_76628_new_n4338_), .B(u0__abc_76628_new_n4337_), .Y(u0__0poc_31_0__13_));
AND2X2 AND2X2_1176 ( .A(u0__abc_76628_new_n4341_), .B(u0__abc_76628_new_n4340_), .Y(u0__0poc_31_0__14_));
AND2X2 AND2X2_1177 ( .A(u0__abc_76628_new_n4344_), .B(u0__abc_76628_new_n4343_), .Y(u0__0poc_31_0__15_));
AND2X2 AND2X2_1178 ( .A(u0__abc_76628_new_n4347_), .B(u0__abc_76628_new_n4346_), .Y(u0__0poc_31_0__16_));
AND2X2 AND2X2_1179 ( .A(u0__abc_76628_new_n4350_), .B(u0__abc_76628_new_n4349_), .Y(u0__0poc_31_0__17_));
AND2X2 AND2X2_118 ( .A(spec_req_cs_4_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1210_));
AND2X2 AND2X2_1180 ( .A(u0__abc_76628_new_n4353_), .B(u0__abc_76628_new_n4352_), .Y(u0__0poc_31_0__18_));
AND2X2 AND2X2_1181 ( .A(u0__abc_76628_new_n4356_), .B(u0__abc_76628_new_n4355_), .Y(u0__0poc_31_0__19_));
AND2X2 AND2X2_1182 ( .A(u0__abc_76628_new_n4359_), .B(u0__abc_76628_new_n4358_), .Y(u0__0poc_31_0__20_));
AND2X2 AND2X2_1183 ( .A(u0__abc_76628_new_n4362_), .B(u0__abc_76628_new_n4361_), .Y(u0__0poc_31_0__21_));
AND2X2 AND2X2_1184 ( .A(u0__abc_76628_new_n4365_), .B(u0__abc_76628_new_n4364_), .Y(u0__0poc_31_0__22_));
AND2X2 AND2X2_1185 ( .A(u0__abc_76628_new_n4368_), .B(u0__abc_76628_new_n4367_), .Y(u0__0poc_31_0__23_));
AND2X2 AND2X2_1186 ( .A(u0__abc_76628_new_n4371_), .B(u0__abc_76628_new_n4370_), .Y(u0__0poc_31_0__24_));
AND2X2 AND2X2_1187 ( .A(u0__abc_76628_new_n4374_), .B(u0__abc_76628_new_n4373_), .Y(u0__0poc_31_0__25_));
AND2X2 AND2X2_1188 ( .A(u0__abc_76628_new_n4377_), .B(u0__abc_76628_new_n4376_), .Y(u0__0poc_31_0__26_));
AND2X2 AND2X2_1189 ( .A(u0__abc_76628_new_n4380_), .B(u0__abc_76628_new_n4379_), .Y(u0__0poc_31_0__27_));
AND2X2 AND2X2_119 ( .A(u0__abc_76628_new_n1211_), .B(u0__abc_76628_new_n1174__bF_buf4), .Y(u0__abc_76628_new_n1212_));
AND2X2 AND2X2_1190 ( .A(u0__abc_76628_new_n4383_), .B(u0__abc_76628_new_n4382_), .Y(u0__0poc_31_0__28_));
AND2X2 AND2X2_1191 ( .A(u0__abc_76628_new_n4386_), .B(u0__abc_76628_new_n4385_), .Y(u0__0poc_31_0__29_));
AND2X2 AND2X2_1192 ( .A(u0__abc_76628_new_n4389_), .B(u0__abc_76628_new_n4388_), .Y(u0__0poc_31_0__30_));
AND2X2 AND2X2_1193 ( .A(u0__abc_76628_new_n4392_), .B(u0__abc_76628_new_n4391_), .Y(u0__0poc_31_0__31_));
AND2X2 AND2X2_1194 ( .A(u0__abc_76628_new_n4399_), .B(u0_wb_addr_r_3_), .Y(u0__abc_76628_new_n4400_));
AND2X2 AND2X2_1195 ( .A(u0__abc_76628_new_n4400_), .B(u0__abc_76628_new_n4396_), .Y(u0__abc_76628_new_n4401_));
AND2X2 AND2X2_1196 ( .A(u0__abc_76628_new_n4404_), .B(u0__abc_76628_new_n4402_), .Y(u0__0csc_mask_r_10_0__0_));
AND2X2 AND2X2_1197 ( .A(u0__abc_76628_new_n4407_), .B(u0__abc_76628_new_n4406_), .Y(u0__0csc_mask_r_10_0__1_));
AND2X2 AND2X2_1198 ( .A(u0__abc_76628_new_n4410_), .B(u0__abc_76628_new_n4409_), .Y(u0__0csc_mask_r_10_0__2_));
AND2X2 AND2X2_1199 ( .A(u0__abc_76628_new_n4413_), .B(u0__abc_76628_new_n4412_), .Y(u0__0csc_mask_r_10_0__3_));
AND2X2 AND2X2_12 ( .A(_abc_85006_new_n272_), .B(_abc_85006_new_n273_), .Y(_abc_85006_new_n274_));
AND2X2 AND2X2_120 ( .A(spec_req_cs_3_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1213_));
AND2X2 AND2X2_1200 ( .A(u0__abc_76628_new_n4416_), .B(u0__abc_76628_new_n4415_), .Y(u0__0csc_mask_r_10_0__4_));
AND2X2 AND2X2_1201 ( .A(u0__abc_76628_new_n4419_), .B(u0__abc_76628_new_n4418_), .Y(u0__0csc_mask_r_10_0__5_));
AND2X2 AND2X2_1202 ( .A(u0__abc_76628_new_n4422_), .B(u0__abc_76628_new_n4421_), .Y(u0__0csc_mask_r_10_0__6_));
AND2X2 AND2X2_1203 ( .A(u0__abc_76628_new_n4425_), .B(u0__abc_76628_new_n4424_), .Y(u0__0csc_mask_r_10_0__7_));
AND2X2 AND2X2_1204 ( .A(u0__abc_76628_new_n4428_), .B(u0__abc_76628_new_n4427_), .Y(u0__0csc_mask_r_10_0__8_));
AND2X2 AND2X2_1205 ( .A(u0__abc_76628_new_n4431_), .B(u0__abc_76628_new_n4430_), .Y(u0__0csc_mask_r_10_0__9_));
AND2X2 AND2X2_1206 ( .A(u0__abc_76628_new_n4434_), .B(u0__abc_76628_new_n4433_), .Y(u0__0csc_mask_r_10_0__10_));
AND2X2 AND2X2_1207 ( .A(u0__abc_76628_new_n4439_), .B(u0__abc_76628_new_n4440_), .Y(u0__0csr_r_10_1__0_));
AND2X2 AND2X2_1208 ( .A(u0__abc_76628_new_n4442_), .B(u0__abc_76628_new_n4443_), .Y(u0__0csr_r_10_1__1_));
AND2X2 AND2X2_1209 ( .A(u0__abc_76628_new_n4445_), .B(u0__abc_76628_new_n4446_), .Y(u0__0csr_r_10_1__2_));
AND2X2 AND2X2_121 ( .A(u0__abc_76628_new_n1214_), .B(u0__abc_76628_new_n1173__bF_buf4), .Y(u0__abc_76628_new_n1215_));
AND2X2 AND2X2_1210 ( .A(u0__abc_76628_new_n4448_), .B(u0__abc_76628_new_n4449_), .Y(u0__0csr_r_10_1__3_));
AND2X2 AND2X2_1211 ( .A(u0__abc_76628_new_n4451_), .B(u0__abc_76628_new_n4452_), .Y(u0__0csr_r_10_1__4_));
AND2X2 AND2X2_1212 ( .A(u0__abc_76628_new_n4454_), .B(u0__abc_76628_new_n4455_), .Y(u0__0csr_r_10_1__5_));
AND2X2 AND2X2_1213 ( .A(u0__abc_76628_new_n4457_), .B(u0__abc_76628_new_n4458_), .Y(u0__0csr_r_10_1__6_));
AND2X2 AND2X2_1214 ( .A(u0__abc_76628_new_n4460_), .B(u0__abc_76628_new_n4461_), .Y(u0__0csr_r_10_1__7_));
AND2X2 AND2X2_1215 ( .A(u0__abc_76628_new_n4463_), .B(u0__abc_76628_new_n4464_), .Y(u0__0csr_r_10_1__8_));
AND2X2 AND2X2_1216 ( .A(u0__abc_76628_new_n4466_), .B(u0__abc_76628_new_n4467_), .Y(u0__0csr_r_10_1__9_));
AND2X2 AND2X2_1217 ( .A(u0__abc_76628_new_n4469_), .B(u0__abc_76628_new_n4470_), .Y(u0__0csr_r2_7_0__0_));
AND2X2 AND2X2_1218 ( .A(u0__abc_76628_new_n4472_), .B(u0__abc_76628_new_n4473_), .Y(u0__0csr_r2_7_0__1_));
AND2X2 AND2X2_1219 ( .A(u0__abc_76628_new_n4475_), .B(u0__abc_76628_new_n4476_), .Y(u0__0csr_r2_7_0__2_));
AND2X2 AND2X2_122 ( .A(spec_req_cs_2_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1216_));
AND2X2 AND2X2_1220 ( .A(u0__abc_76628_new_n4478_), .B(u0__abc_76628_new_n4479_), .Y(u0__0csr_r2_7_0__3_));
AND2X2 AND2X2_1221 ( .A(u0__abc_76628_new_n4481_), .B(u0__abc_76628_new_n4482_), .Y(u0__0csr_r2_7_0__4_));
AND2X2 AND2X2_1222 ( .A(u0__abc_76628_new_n4484_), .B(u0__abc_76628_new_n4485_), .Y(u0__0csr_r2_7_0__5_));
AND2X2 AND2X2_1223 ( .A(u0__abc_76628_new_n4487_), .B(u0__abc_76628_new_n4488_), .Y(u0__0csr_r2_7_0__6_));
AND2X2 AND2X2_1224 ( .A(u0__abc_76628_new_n4490_), .B(u0__abc_76628_new_n4491_), .Y(u0__0csr_r2_7_0__7_));
AND2X2 AND2X2_1225 ( .A(u0__abc_76628_new_n4493_), .B(u0__abc_76628_new_n4494_), .Y(u0__abc_76628_new_n4495_));
AND2X2 AND2X2_1226 ( .A(u0__abc_76628_new_n4495_), .B(\wb_addr_i[6] ), .Y(u0__abc_76628_new_n4496_));
AND2X2 AND2X2_1227 ( .A(u0__abc_76628_new_n4497_), .B(u0__abc_76628_new_n4498_), .Y(u0__abc_76628_new_n4499_));
AND2X2 AND2X2_1228 ( .A(u0__abc_76628_new_n4496_), .B(u0__abc_76628_new_n4499_), .Y(u0__abc_76628_new_n4500_));
AND2X2 AND2X2_1229 ( .A(u0__abc_76628_new_n4500__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4501_));
AND2X2 AND2X2_123 ( .A(u0__abc_76628_new_n1217_), .B(u0__abc_76628_new_n1172__bF_buf4), .Y(u0__abc_76628_new_n1218_));
AND2X2 AND2X2_1230 ( .A(u0__abc_76628_new_n4497_), .B(\wb_addr_i[2] ), .Y(u0__abc_76628_new_n4502_));
AND2X2 AND2X2_1231 ( .A(u0__abc_76628_new_n4496_), .B(u0__abc_76628_new_n4502_), .Y(u0__abc_76628_new_n4503_));
AND2X2 AND2X2_1232 ( .A(u0__abc_76628_new_n4503__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4504_));
AND2X2 AND2X2_1233 ( .A(\wb_addr_i[3] ), .B(\wb_addr_i[2] ), .Y(u0__abc_76628_new_n4506_));
AND2X2 AND2X2_1234 ( .A(u0__abc_76628_new_n4496_), .B(u0__abc_76628_new_n4506_), .Y(u0__abc_76628_new_n4507_));
AND2X2 AND2X2_1235 ( .A(u0__abc_76628_new_n4507__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4508_));
AND2X2 AND2X2_1236 ( .A(u0__abc_76628_new_n4498_), .B(\wb_addr_i[3] ), .Y(u0__abc_76628_new_n4509_));
AND2X2 AND2X2_1237 ( .A(u0__abc_76628_new_n4496_), .B(u0__abc_76628_new_n4509_), .Y(u0__abc_76628_new_n4510_));
AND2X2 AND2X2_1238 ( .A(u0__abc_76628_new_n4510__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4511_));
AND2X2 AND2X2_1239 ( .A(u0__abc_76628_new_n4494_), .B(\wb_addr_i[5] ), .Y(u0__abc_76628_new_n4514_));
AND2X2 AND2X2_124 ( .A(spec_req_cs_1_bF_buf1_), .B(u0_tms1_1_), .Y(u0__abc_76628_new_n1219_));
AND2X2 AND2X2_1240 ( .A(u0__abc_76628_new_n4509_), .B(u0__abc_76628_new_n4515_), .Y(u0__abc_76628_new_n4516_));
AND2X2 AND2X2_1241 ( .A(u0__abc_76628_new_n4516_), .B(u0__abc_76628_new_n4514_), .Y(u0__abc_76628_new_n4517_));
AND2X2 AND2X2_1242 ( .A(u0__abc_76628_new_n4517__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4518_));
AND2X2 AND2X2_1243 ( .A(u0__abc_76628_new_n4499_), .B(u0__abc_76628_new_n4515_), .Y(u0__abc_76628_new_n4519_));
AND2X2 AND2X2_1244 ( .A(u0__abc_76628_new_n4519_), .B(u0__abc_76628_new_n4514_), .Y(u0__abc_76628_new_n4520_));
AND2X2 AND2X2_1245 ( .A(u0__abc_76628_new_n4520__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4521_));
AND2X2 AND2X2_1246 ( .A(u0__abc_76628_new_n4502_), .B(u0__abc_76628_new_n4515_), .Y(u0__abc_76628_new_n4522_));
AND2X2 AND2X2_1247 ( .A(u0__abc_76628_new_n4522_), .B(u0__abc_76628_new_n4514_), .Y(u0__abc_76628_new_n4523_));
AND2X2 AND2X2_1248 ( .A(u0__abc_76628_new_n4523__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4524_));
AND2X2 AND2X2_1249 ( .A(u0__abc_76628_new_n4506_), .B(u0__abc_76628_new_n4515_), .Y(u0__abc_76628_new_n4527_));
AND2X2 AND2X2_125 ( .A(u0__abc_76628_new_n1169__bF_buf4), .B(u0__abc_76628_new_n1222_), .Y(u0__abc_76628_new_n1223_));
AND2X2 AND2X2_1250 ( .A(u0__abc_76628_new_n4527_), .B(u0__abc_76628_new_n4514_), .Y(u0__abc_76628_new_n4528_));
AND2X2 AND2X2_1251 ( .A(u0__abc_76628_new_n4528__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4529_));
AND2X2 AND2X2_1252 ( .A(\wb_addr_i[5] ), .B(\wb_addr_i[4] ), .Y(u0__abc_76628_new_n4530_));
AND2X2 AND2X2_1253 ( .A(u0__abc_76628_new_n4527_), .B(u0__abc_76628_new_n4530_), .Y(u0__abc_76628_new_n4531_));
AND2X2 AND2X2_1254 ( .A(u0__abc_76628_new_n4531__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4532_));
AND2X2 AND2X2_1255 ( .A(u0__abc_76628_new_n4536_), .B(\wb_addr_i[6] ), .Y(u0__abc_76628_new_n4537_));
AND2X2 AND2X2_1256 ( .A(u0__abc_76628_new_n4495_), .B(u0__abc_76628_new_n4515_), .Y(u0__abc_76628_new_n4538_));
AND2X2 AND2X2_1257 ( .A(u0__abc_76628_new_n4539_), .B(u0__abc_76628_new_n4538_), .Y(u0__abc_76628_new_n4540_));
AND2X2 AND2X2_1258 ( .A(u0__abc_76628_new_n4541__bF_buf3), .B(u0_csr_0_), .Y(u0__abc_76628_new_n4542_));
AND2X2 AND2X2_1259 ( .A(u0__abc_76628_new_n4493_), .B(\wb_addr_i[4] ), .Y(u0__abc_76628_new_n4543_));
AND2X2 AND2X2_126 ( .A(u0__abc_76628_new_n1221_), .B(u0__abc_76628_new_n1223_), .Y(u0__abc_76628_new_n1224_));
AND2X2 AND2X2_1260 ( .A(u0__abc_76628_new_n4543_), .B(u0__abc_76628_new_n4515_), .Y(u0__abc_76628_new_n4544_));
AND2X2 AND2X2_1261 ( .A(u0__abc_76628_new_n4544_), .B(u0__abc_76628_new_n4509_), .Y(u0__abc_76628_new_n4545_));
AND2X2 AND2X2_1262 ( .A(u0__abc_76628_new_n4545__bF_buf4), .B(u0_csc1_0_), .Y(u0__abc_76628_new_n4546_));
AND2X2 AND2X2_1263 ( .A(u0__abc_76628_new_n4544_), .B(u0__abc_76628_new_n4499_), .Y(u0__abc_76628_new_n4547_));
AND2X2 AND2X2_1264 ( .A(u0__abc_76628_new_n4547__bF_buf4), .B(u0_csc0_0_), .Y(u0__abc_76628_new_n4548_));
AND2X2 AND2X2_1265 ( .A(u0__abc_76628_new_n4544_), .B(u0__abc_76628_new_n4502_), .Y(u0__abc_76628_new_n4549_));
AND2X2 AND2X2_1266 ( .A(u0__abc_76628_new_n4549__bF_buf4), .B(u0_tms0_0_), .Y(u0__abc_76628_new_n4550_));
AND2X2 AND2X2_1267 ( .A(u0__abc_76628_new_n4516_), .B(u0__abc_76628_new_n4530_), .Y(u0__abc_76628_new_n4554_));
AND2X2 AND2X2_1268 ( .A(u0__abc_76628_new_n4554__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4555_));
AND2X2 AND2X2_1269 ( .A(u0__abc_76628_new_n4522_), .B(u0__abc_76628_new_n4530_), .Y(u0__abc_76628_new_n4556_));
AND2X2 AND2X2_127 ( .A(u0__abc_76628_new_n1170__bF_buf4), .B(sp_tms_2_), .Y(u0__abc_76628_new_n1226_));
AND2X2 AND2X2_1270 ( .A(u0__abc_76628_new_n4556__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4557_));
AND2X2 AND2X2_1271 ( .A(u0__abc_76628_new_n4519_), .B(u0__abc_76628_new_n4530_), .Y(u0__abc_76628_new_n4558_));
AND2X2 AND2X2_1272 ( .A(u0__abc_76628_new_n4558__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4559_));
AND2X2 AND2X2_1273 ( .A(u0__abc_76628_new_n4544_), .B(u0__abc_76628_new_n4506_), .Y(u0__abc_76628_new_n4562_));
AND2X2 AND2X2_1274 ( .A(u0__abc_76628_new_n4562__bF_buf4), .B(u0_tms1_0_), .Y(u0__abc_76628_new_n4563_));
AND2X2 AND2X2_1275 ( .A(u0__abc_76628_new_n4516_), .B(u0__abc_76628_new_n4495_), .Y(u0__abc_76628_new_n4564_));
AND2X2 AND2X2_1276 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_0_), .Y(u0__abc_76628_new_n4565_));
AND2X2 AND2X2_1277 ( .A(u0__abc_76628_new_n4522_), .B(u0__abc_76628_new_n4495_), .Y(u0__abc_76628_new_n4566_));
AND2X2 AND2X2_1278 ( .A(u0__abc_76628_new_n4566__bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_0_), .Y(u0__abc_76628_new_n4567_));
AND2X2 AND2X2_1279 ( .A(u0__abc_76628_new_n4500__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4573_));
AND2X2 AND2X2_128 ( .A(spec_req_cs_5_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1227_));
AND2X2 AND2X2_1280 ( .A(u0__abc_76628_new_n4531__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4574_));
AND2X2 AND2X2_1281 ( .A(u0__abc_76628_new_n4507__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4576_));
AND2X2 AND2X2_1282 ( .A(u0__abc_76628_new_n4556__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4577_));
AND2X2 AND2X2_1283 ( .A(u0__abc_76628_new_n4549__bF_buf3), .B(u0_tms0_1_), .Y(u0__abc_76628_new_n4579_));
AND2X2 AND2X2_1284 ( .A(u0__abc_76628_new_n4545__bF_buf3), .B(u0_csc1_1_), .Y(u0__abc_76628_new_n4580_));
AND2X2 AND2X2_1285 ( .A(u0__abc_76628_new_n4510__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4584_));
AND2X2 AND2X2_1286 ( .A(u0__abc_76628_new_n4547__bF_buf3), .B(u0_csc0_1_), .Y(u0__abc_76628_new_n4585_));
AND2X2 AND2X2_1287 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_1_), .Y(u0__abc_76628_new_n4587_));
AND2X2 AND2X2_1288 ( .A(u0__abc_76628_new_n4558__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4588_));
AND2X2 AND2X2_1289 ( .A(u0__abc_76628_new_n4517__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4591_));
AND2X2 AND2X2_129 ( .A(u0__abc_76628_new_n1229_), .B(u0__abc_76628_new_n1179__bF_buf3), .Y(u0__abc_76628_new_n1230_));
AND2X2 AND2X2_1290 ( .A(u0__abc_76628_new_n4528__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4592_));
AND2X2 AND2X2_1291 ( .A(u0__abc_76628_new_n4503__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4594_));
AND2X2 AND2X2_1292 ( .A(u0__abc_76628_new_n4554__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4595_));
AND2X2 AND2X2_1293 ( .A(u0__abc_76628_new_n4541__bF_buf2), .B(u0_csr_1_), .Y(u0__abc_76628_new_n4599_));
AND2X2 AND2X2_1294 ( .A(u0__abc_76628_new_n4520__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4600_));
AND2X2 AND2X2_1295 ( .A(u0__abc_76628_new_n4562__bF_buf3), .B(u0_tms1_1_), .Y(u0__abc_76628_new_n4601_));
AND2X2 AND2X2_1296 ( .A(u0__abc_76628_new_n4566__bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_1_), .Y(u0__abc_76628_new_n4603_));
AND2X2 AND2X2_1297 ( .A(u0__abc_76628_new_n4523__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4604_));
AND2X2 AND2X2_1298 ( .A(u0__abc_76628_new_n4500__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4610_));
AND2X2 AND2X2_1299 ( .A(u0__abc_76628_new_n4507__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4611_));
AND2X2 AND2X2_13 ( .A(_abc_85006_new_n275_), .B(_abc_85006_new_n276_), .Y(obct_cs_5_));
AND2X2 AND2X2_130 ( .A(u0__abc_76628_new_n1230_), .B(u0__abc_76628_new_n1228_), .Y(u0__abc_76628_new_n1231_));
AND2X2 AND2X2_1300 ( .A(u0__abc_76628_new_n4520__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4613_));
AND2X2 AND2X2_1301 ( .A(u0__abc_76628_new_n4523__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4614_));
AND2X2 AND2X2_1302 ( .A(u0__abc_76628_new_n4549__bF_buf2), .B(u0_tms0_2_), .Y(u0__abc_76628_new_n4616_));
AND2X2 AND2X2_1303 ( .A(u0__abc_76628_new_n4545__bF_buf2), .B(u0_csc1_2_), .Y(u0__abc_76628_new_n4617_));
AND2X2 AND2X2_1304 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_2_), .Y(u0__abc_76628_new_n4621_));
AND2X2 AND2X2_1305 ( .A(u0__abc_76628_new_n4547__bF_buf2), .B(u0_csc0_2_), .Y(u0__abc_76628_new_n4622_));
AND2X2 AND2X2_1306 ( .A(u0__abc_76628_new_n4554__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4624_));
AND2X2 AND2X2_1307 ( .A(u0__abc_76628_new_n4528__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4625_));
AND2X2 AND2X2_1308 ( .A(u0__abc_76628_new_n4503__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4628_));
AND2X2 AND2X2_1309 ( .A(u0__abc_76628_new_n4558__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4629_));
AND2X2 AND2X2_131 ( .A(u0__abc_76628_new_n1232_), .B(u0__abc_76628_new_n1175__bF_buf3), .Y(u0__abc_76628_new_n1233_));
AND2X2 AND2X2_1310 ( .A(u0__abc_76628_new_n4566__bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_2_), .Y(u0__abc_76628_new_n4631_));
AND2X2 AND2X2_1311 ( .A(u0__abc_76628_new_n4562__bF_buf2), .B(u0_tms1_2_), .Y(u0__abc_76628_new_n4632_));
AND2X2 AND2X2_1312 ( .A(u0__abc_76628_new_n4541__bF_buf1), .B(fs), .Y(u0__abc_76628_new_n4636_));
AND2X2 AND2X2_1313 ( .A(u0__abc_76628_new_n4531__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4637_));
AND2X2 AND2X2_1314 ( .A(u0__abc_76628_new_n4517__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4638_));
AND2X2 AND2X2_1315 ( .A(u0__abc_76628_new_n4510__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4640_));
AND2X2 AND2X2_1316 ( .A(u0__abc_76628_new_n4556__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4641_));
AND2X2 AND2X2_1317 ( .A(u0__abc_76628_new_n4500__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4647_));
AND2X2 AND2X2_1318 ( .A(u0__abc_76628_new_n4503__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4648_));
AND2X2 AND2X2_1319 ( .A(u0__abc_76628_new_n4507__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4650_));
AND2X2 AND2X2_132 ( .A(spec_req_cs_4_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1234_));
AND2X2 AND2X2_1320 ( .A(u0__abc_76628_new_n4510__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4651_));
AND2X2 AND2X2_1321 ( .A(u0__abc_76628_new_n4517__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4654_));
AND2X2 AND2X2_1322 ( .A(u0__abc_76628_new_n4523__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4655_));
AND2X2 AND2X2_1323 ( .A(u0__abc_76628_new_n4520__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4656_));
AND2X2 AND2X2_1324 ( .A(u0__abc_76628_new_n4531__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4659_));
AND2X2 AND2X2_1325 ( .A(u0__abc_76628_new_n4528__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4660_));
AND2X2 AND2X2_1326 ( .A(u0__abc_76628_new_n4541__bF_buf0), .B(u0_csr_3_), .Y(u0__abc_76628_new_n4664_));
AND2X2 AND2X2_1327 ( .A(u0__abc_76628_new_n4547__bF_buf1), .B(u0_csc0_3_), .Y(u0__abc_76628_new_n4665_));
AND2X2 AND2X2_1328 ( .A(u0__abc_76628_new_n4549__bF_buf1), .B(u0_tms0_3_), .Y(u0__abc_76628_new_n4666_));
AND2X2 AND2X2_1329 ( .A(u0__abc_76628_new_n4545__bF_buf1), .B(u0_csc1_3_), .Y(u0__abc_76628_new_n4668_));
AND2X2 AND2X2_133 ( .A(u0__abc_76628_new_n1235_), .B(u0__abc_76628_new_n1174__bF_buf3), .Y(u0__abc_76628_new_n1236_));
AND2X2 AND2X2_1330 ( .A(u0__abc_76628_new_n4554__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4671_));
AND2X2 AND2X2_1331 ( .A(u0__abc_76628_new_n4556__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4672_));
AND2X2 AND2X2_1332 ( .A(u0__abc_76628_new_n4558__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4673_));
AND2X2 AND2X2_1333 ( .A(u0__abc_76628_new_n4562__bF_buf1), .B(u0_tms1_3_), .Y(u0__abc_76628_new_n4676_));
AND2X2 AND2X2_1334 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_3_), .Y(u0__abc_76628_new_n4677_));
AND2X2 AND2X2_1335 ( .A(u0__abc_76628_new_n4566__bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_3_), .Y(u0__abc_76628_new_n4678_));
AND2X2 AND2X2_1336 ( .A(u0__abc_76628_new_n4510__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4684_));
AND2X2 AND2X2_1337 ( .A(u0__abc_76628_new_n4556__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4685_));
AND2X2 AND2X2_1338 ( .A(u0__abc_76628_new_n4500__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4687_));
AND2X2 AND2X2_1339 ( .A(u0__abc_76628_new_n4517__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4688_));
AND2X2 AND2X2_134 ( .A(spec_req_cs_3_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1237_));
AND2X2 AND2X2_1340 ( .A(u0__abc_76628_new_n4566__bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_4_), .Y(u0__abc_76628_new_n4690_));
AND2X2 AND2X2_1341 ( .A(u0__abc_76628_new_n4547__bF_buf0), .B(u0_csc0_4_), .Y(u0__abc_76628_new_n4691_));
AND2X2 AND2X2_1342 ( .A(u0__abc_76628_new_n4507__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4695_));
AND2X2 AND2X2_1343 ( .A(u0__abc_76628_new_n4562__bF_buf0), .B(u0_tms1_4_), .Y(u0__abc_76628_new_n4696_));
AND2X2 AND2X2_1344 ( .A(u0__abc_76628_new_n4520__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4698_));
AND2X2 AND2X2_1345 ( .A(u0__abc_76628_new_n4545__bF_buf0), .B(u0_csc1_4_), .Y(u0__abc_76628_new_n4699_));
AND2X2 AND2X2_1346 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_4_), .Y(u0__abc_76628_new_n4702_));
AND2X2 AND2X2_1347 ( .A(u0__abc_76628_new_n4554__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4703_));
AND2X2 AND2X2_1348 ( .A(u0__abc_76628_new_n4531__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4705_));
AND2X2 AND2X2_1349 ( .A(u0__abc_76628_new_n4523__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4706_));
AND2X2 AND2X2_135 ( .A(u0__abc_76628_new_n1238_), .B(u0__abc_76628_new_n1173__bF_buf3), .Y(u0__abc_76628_new_n1239_));
AND2X2 AND2X2_1350 ( .A(u0__abc_76628_new_n4541__bF_buf3), .B(u0_csr_4_), .Y(u0__abc_76628_new_n4710_));
AND2X2 AND2X2_1351 ( .A(u0__abc_76628_new_n4528__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4711_));
AND2X2 AND2X2_1352 ( .A(u0__abc_76628_new_n4549__bF_buf0), .B(u0_tms0_4_), .Y(u0__abc_76628_new_n4712_));
AND2X2 AND2X2_1353 ( .A(u0__abc_76628_new_n4503__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4714_));
AND2X2 AND2X2_1354 ( .A(u0__abc_76628_new_n4558__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4715_));
AND2X2 AND2X2_1355 ( .A(u0__abc_76628_new_n4500__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4721_));
AND2X2 AND2X2_1356 ( .A(u0__abc_76628_new_n4503__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4722_));
AND2X2 AND2X2_1357 ( .A(u0__abc_76628_new_n4510__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4724_));
AND2X2 AND2X2_1358 ( .A(u0__abc_76628_new_n4507__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4725_));
AND2X2 AND2X2_1359 ( .A(u0__abc_76628_new_n4517__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4728_));
AND2X2 AND2X2_136 ( .A(spec_req_cs_2_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1240_));
AND2X2 AND2X2_1360 ( .A(u0__abc_76628_new_n4520__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4729_));
AND2X2 AND2X2_1361 ( .A(u0__abc_76628_new_n4523__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4730_));
AND2X2 AND2X2_1362 ( .A(u0__abc_76628_new_n4531__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4733_));
AND2X2 AND2X2_1363 ( .A(u0__abc_76628_new_n4528__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4734_));
AND2X2 AND2X2_1364 ( .A(u0__abc_76628_new_n4541__bF_buf2), .B(u0_csr_5_), .Y(u0__abc_76628_new_n4738_));
AND2X2 AND2X2_1365 ( .A(u0__abc_76628_new_n4545__bF_buf4), .B(u0_csc1_5_), .Y(u0__abc_76628_new_n4739_));
AND2X2 AND2X2_1366 ( .A(u0__abc_76628_new_n4547__bF_buf4), .B(u0_csc0_5_), .Y(u0__abc_76628_new_n4740_));
AND2X2 AND2X2_1367 ( .A(u0__abc_76628_new_n4549__bF_buf4), .B(u0_tms0_5_), .Y(u0__abc_76628_new_n4741_));
AND2X2 AND2X2_1368 ( .A(u0__abc_76628_new_n4554__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4745_));
AND2X2 AND2X2_1369 ( .A(u0__abc_76628_new_n4558__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4746_));
AND2X2 AND2X2_137 ( .A(u0__abc_76628_new_n1241_), .B(u0__abc_76628_new_n1172__bF_buf3), .Y(u0__abc_76628_new_n1242_));
AND2X2 AND2X2_1370 ( .A(u0__abc_76628_new_n4556__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4747_));
AND2X2 AND2X2_1371 ( .A(u0__abc_76628_new_n4562__bF_buf4), .B(u0_tms1_5_), .Y(u0__abc_76628_new_n4750_));
AND2X2 AND2X2_1372 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_5_), .Y(u0__abc_76628_new_n4751_));
AND2X2 AND2X2_1373 ( .A(u0__abc_76628_new_n4566__bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_5_), .Y(u0__abc_76628_new_n4752_));
AND2X2 AND2X2_1374 ( .A(u0__abc_76628_new_n4510__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4758_));
AND2X2 AND2X2_1375 ( .A(u0__abc_76628_new_n4556__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4759_));
AND2X2 AND2X2_1376 ( .A(u0__abc_76628_new_n4500__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4761_));
AND2X2 AND2X2_1377 ( .A(u0__abc_76628_new_n4517__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4762_));
AND2X2 AND2X2_1378 ( .A(u0__abc_76628_new_n4566__bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_6_), .Y(u0__abc_76628_new_n4764_));
AND2X2 AND2X2_1379 ( .A(u0__abc_76628_new_n4549__bF_buf3), .B(u0_tms0_6_), .Y(u0__abc_76628_new_n4765_));
AND2X2 AND2X2_138 ( .A(spec_req_cs_1_bF_buf0_), .B(u0_tms1_2_), .Y(u0__abc_76628_new_n1243_));
AND2X2 AND2X2_1380 ( .A(u0__abc_76628_new_n4507__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4769_));
AND2X2 AND2X2_1381 ( .A(u0__abc_76628_new_n4562__bF_buf3), .B(u0_tms1_6_), .Y(u0__abc_76628_new_n4770_));
AND2X2 AND2X2_1382 ( .A(u0__abc_76628_new_n4520__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4772_));
AND2X2 AND2X2_1383 ( .A(u0__abc_76628_new_n4545__bF_buf3), .B(u0_csc1_6_), .Y(u0__abc_76628_new_n4773_));
AND2X2 AND2X2_1384 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_6_), .Y(u0__abc_76628_new_n4776_));
AND2X2 AND2X2_1385 ( .A(u0__abc_76628_new_n4554__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4777_));
AND2X2 AND2X2_1386 ( .A(u0__abc_76628_new_n4531__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4779_));
AND2X2 AND2X2_1387 ( .A(u0__abc_76628_new_n4523__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4780_));
AND2X2 AND2X2_1388 ( .A(u0__abc_76628_new_n4541__bF_buf1), .B(u0_csr_6_), .Y(u0__abc_76628_new_n4784_));
AND2X2 AND2X2_1389 ( .A(u0__abc_76628_new_n4528__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4785_));
AND2X2 AND2X2_139 ( .A(u0__abc_76628_new_n1169__bF_buf3), .B(u0__abc_76628_new_n1246_), .Y(u0__abc_76628_new_n1247_));
AND2X2 AND2X2_1390 ( .A(u0__abc_76628_new_n4547__bF_buf3), .B(u0_csc0_6_), .Y(u0__abc_76628_new_n4786_));
AND2X2 AND2X2_1391 ( .A(u0__abc_76628_new_n4503__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4788_));
AND2X2 AND2X2_1392 ( .A(u0__abc_76628_new_n4558__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4789_));
AND2X2 AND2X2_1393 ( .A(u0__abc_76628_new_n4500__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4795_));
AND2X2 AND2X2_1394 ( .A(u0__abc_76628_new_n4503__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4796_));
AND2X2 AND2X2_1395 ( .A(u0__abc_76628_new_n4510__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4798_));
AND2X2 AND2X2_1396 ( .A(u0__abc_76628_new_n4507__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4799_));
AND2X2 AND2X2_1397 ( .A(u0__abc_76628_new_n4528__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4802_));
AND2X2 AND2X2_1398 ( .A(u0__abc_76628_new_n4531__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4803_));
AND2X2 AND2X2_1399 ( .A(u0__abc_76628_new_n4517__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4805_));
AND2X2 AND2X2_14 ( .A(_abc_85006_new_n278_), .B(_abc_85006_new_n279_), .Y(_abc_85006_new_n280_));
AND2X2 AND2X2_140 ( .A(u0__abc_76628_new_n1245_), .B(u0__abc_76628_new_n1247_), .Y(u0__abc_76628_new_n1248_));
AND2X2 AND2X2_1400 ( .A(u0__abc_76628_new_n4523__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4806_));
AND2X2 AND2X2_1401 ( .A(u0__abc_76628_new_n4520__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4807_));
AND2X2 AND2X2_1402 ( .A(u0__abc_76628_new_n4541__bF_buf0), .B(u0_csr_7_), .Y(u0__abc_76628_new_n4812_));
AND2X2 AND2X2_1403 ( .A(u0__abc_76628_new_n4545__bF_buf2), .B(u0_csc1_7_), .Y(u0__abc_76628_new_n4813_));
AND2X2 AND2X2_1404 ( .A(u0__abc_76628_new_n4547__bF_buf2), .B(u0_csc0_7_), .Y(u0__abc_76628_new_n4814_));
AND2X2 AND2X2_1405 ( .A(u0__abc_76628_new_n4549__bF_buf2), .B(u0_tms0_7_), .Y(u0__abc_76628_new_n4815_));
AND2X2 AND2X2_1406 ( .A(u0__abc_76628_new_n4554__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4819_));
AND2X2 AND2X2_1407 ( .A(u0__abc_76628_new_n4558__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4820_));
AND2X2 AND2X2_1408 ( .A(u0__abc_76628_new_n4556__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4821_));
AND2X2 AND2X2_1409 ( .A(u0__abc_76628_new_n4562__bF_buf2), .B(u0_tms1_7_), .Y(u0__abc_76628_new_n4824_));
AND2X2 AND2X2_141 ( .A(u0__abc_76628_new_n1170__bF_buf3), .B(sp_tms_3_), .Y(u0__abc_76628_new_n1250_));
AND2X2 AND2X2_1410 ( .A(u0__abc_76628_new_n4566__bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_7_), .Y(u0__abc_76628_new_n4825_));
AND2X2 AND2X2_1411 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_7_), .Y(u0__abc_76628_new_n4826_));
AND2X2 AND2X2_1412 ( .A(u0__abc_76628_new_n4503__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4832_));
AND2X2 AND2X2_1413 ( .A(u0__abc_76628_new_n4520__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4833_));
AND2X2 AND2X2_1414 ( .A(u0__abc_76628_new_n4510__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4835_));
AND2X2 AND2X2_1415 ( .A(u0__abc_76628_new_n4528__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4836_));
AND2X2 AND2X2_1416 ( .A(u0__abc_76628_new_n4547__bF_buf1), .B(u0_csc0_8_), .Y(u0__abc_76628_new_n4838_));
AND2X2 AND2X2_1417 ( .A(u0__abc_76628_new_n4545__bF_buf1), .B(u0_csc1_8_), .Y(u0__abc_76628_new_n4839_));
AND2X2 AND2X2_1418 ( .A(u0__abc_76628_new_n4517__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4843_));
AND2X2 AND2X2_1419 ( .A(u0__abc_76628_new_n4549__bF_buf1), .B(u0_tms0_8_), .Y(u0__abc_76628_new_n4844_));
AND2X2 AND2X2_142 ( .A(spec_req_cs_5_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1251_));
AND2X2 AND2X2_1420 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_8_), .Y(u0__abc_76628_new_n4846_));
AND2X2 AND2X2_1421 ( .A(u0__abc_76628_new_n4507__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4847_));
AND2X2 AND2X2_1422 ( .A(u0__abc_76628_new_n4556__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4850_));
AND2X2 AND2X2_1423 ( .A(u0__abc_76628_new_n4558__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4851_));
AND2X2 AND2X2_1424 ( .A(u0__abc_76628_new_n4500__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4853_));
AND2X2 AND2X2_1425 ( .A(u0__abc_76628_new_n4523__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4854_));
AND2X2 AND2X2_1426 ( .A(u0__abc_76628_new_n4541__bF_buf3), .B(ref_int_0_), .Y(u0__abc_76628_new_n4858_));
AND2X2 AND2X2_1427 ( .A(u0__abc_76628_new_n4554__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4859_));
AND2X2 AND2X2_1428 ( .A(u0__abc_76628_new_n4562__bF_buf1), .B(u0_tms1_8_), .Y(u0__abc_76628_new_n4860_));
AND2X2 AND2X2_1429 ( .A(u0__abc_76628_new_n4566__bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_8_), .Y(u0__abc_76628_new_n4862_));
AND2X2 AND2X2_143 ( .A(u0__abc_76628_new_n1253_), .B(u0__abc_76628_new_n1179__bF_buf2), .Y(u0__abc_76628_new_n1254_));
AND2X2 AND2X2_1430 ( .A(u0__abc_76628_new_n4531__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n4863_));
AND2X2 AND2X2_1431 ( .A(u0__abc_76628_new_n4500__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4869_));
AND2X2 AND2X2_1432 ( .A(u0__abc_76628_new_n4503__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4870_));
AND2X2 AND2X2_1433 ( .A(u0__abc_76628_new_n4507__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4872_));
AND2X2 AND2X2_1434 ( .A(u0__abc_76628_new_n4510__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4873_));
AND2X2 AND2X2_1435 ( .A(u0__abc_76628_new_n4517__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4876_));
AND2X2 AND2X2_1436 ( .A(u0__abc_76628_new_n4523__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4877_));
AND2X2 AND2X2_1437 ( .A(u0__abc_76628_new_n4520__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4878_));
AND2X2 AND2X2_1438 ( .A(u0__abc_76628_new_n4531__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4881_));
AND2X2 AND2X2_1439 ( .A(u0__abc_76628_new_n4528__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4882_));
AND2X2 AND2X2_144 ( .A(u0__abc_76628_new_n1254_), .B(u0__abc_76628_new_n1252_), .Y(u0__abc_76628_new_n1255_));
AND2X2 AND2X2_1440 ( .A(u0__abc_76628_new_n4541__bF_buf2), .B(ref_int_1_), .Y(u0__abc_76628_new_n4886_));
AND2X2 AND2X2_1441 ( .A(u0__abc_76628_new_n4547__bF_buf0), .B(u0_csc0_9_), .Y(u0__abc_76628_new_n4887_));
AND2X2 AND2X2_1442 ( .A(u0__abc_76628_new_n4549__bF_buf0), .B(u0_tms0_9_), .Y(u0__abc_76628_new_n4888_));
AND2X2 AND2X2_1443 ( .A(u0__abc_76628_new_n4545__bF_buf0), .B(u0_csc1_9_), .Y(u0__abc_76628_new_n4890_));
AND2X2 AND2X2_1444 ( .A(u0__abc_76628_new_n4554__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4893_));
AND2X2 AND2X2_1445 ( .A(u0__abc_76628_new_n4556__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4894_));
AND2X2 AND2X2_1446 ( .A(u0__abc_76628_new_n4558__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n4895_));
AND2X2 AND2X2_1447 ( .A(u0__abc_76628_new_n4562__bF_buf0), .B(u0_tms1_9_), .Y(u0__abc_76628_new_n4898_));
AND2X2 AND2X2_1448 ( .A(u0__abc_76628_new_n4566__bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_9_), .Y(u0__abc_76628_new_n4899_));
AND2X2 AND2X2_1449 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_9_), .Y(u0__abc_76628_new_n4900_));
AND2X2 AND2X2_145 ( .A(u0__abc_76628_new_n1256_), .B(u0__abc_76628_new_n1175__bF_buf2), .Y(u0__abc_76628_new_n1257_));
AND2X2 AND2X2_1450 ( .A(u0__abc_76628_new_n4510__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4906_));
AND2X2 AND2X2_1451 ( .A(u0__abc_76628_new_n4556__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4907_));
AND2X2 AND2X2_1452 ( .A(u0__abc_76628_new_n4500__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4909_));
AND2X2 AND2X2_1453 ( .A(u0__abc_76628_new_n4517__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4910_));
AND2X2 AND2X2_1454 ( .A(u0__abc_76628_new_n4566__bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_10_), .Y(u0__abc_76628_new_n4912_));
AND2X2 AND2X2_1455 ( .A(u0__abc_76628_new_n4549__bF_buf4), .B(u0_tms0_10_), .Y(u0__abc_76628_new_n4913_));
AND2X2 AND2X2_1456 ( .A(u0__abc_76628_new_n4507__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4917_));
AND2X2 AND2X2_1457 ( .A(u0__abc_76628_new_n4562__bF_buf4), .B(u0_tms1_10_), .Y(u0__abc_76628_new_n4918_));
AND2X2 AND2X2_1458 ( .A(u0__abc_76628_new_n4520__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4920_));
AND2X2 AND2X2_1459 ( .A(u0__abc_76628_new_n4545__bF_buf4), .B(u0_csc1_10_), .Y(u0__abc_76628_new_n4921_));
AND2X2 AND2X2_146 ( .A(spec_req_cs_4_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1258_));
AND2X2 AND2X2_1460 ( .A(u0__abc_76628_new_n4564_), .B(u0_csc_mask_10_), .Y(u0__abc_76628_new_n4924_));
AND2X2 AND2X2_1461 ( .A(u0__abc_76628_new_n4554__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4925_));
AND2X2 AND2X2_1462 ( .A(u0__abc_76628_new_n4531__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4927_));
AND2X2 AND2X2_1463 ( .A(u0__abc_76628_new_n4523__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4928_));
AND2X2 AND2X2_1464 ( .A(u0__abc_76628_new_n4541__bF_buf1), .B(ref_int_2_), .Y(u0__abc_76628_new_n4932_));
AND2X2 AND2X2_1465 ( .A(u0__abc_76628_new_n4528__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4933_));
AND2X2 AND2X2_1466 ( .A(u0__abc_76628_new_n4547__bF_buf4), .B(u0_csc0_10_), .Y(u0__abc_76628_new_n4934_));
AND2X2 AND2X2_1467 ( .A(u0__abc_76628_new_n4503__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4936_));
AND2X2 AND2X2_1468 ( .A(u0__abc_76628_new_n4558__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n4937_));
AND2X2 AND2X2_1469 ( .A(u0__abc_76628_new_n4558__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4943_));
AND2X2 AND2X2_147 ( .A(u0__abc_76628_new_n1259_), .B(u0__abc_76628_new_n1174__bF_buf2), .Y(u0__abc_76628_new_n1260_));
AND2X2 AND2X2_1470 ( .A(u0__abc_76628_new_n4554__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4944_));
AND2X2 AND2X2_1471 ( .A(u0__abc_76628_new_n4507__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4946_));
AND2X2 AND2X2_1472 ( .A(u0__abc_76628_new_n4510__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4947_));
AND2X2 AND2X2_1473 ( .A(u0__abc_76628_new_n4566__bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_11_), .Y(u0__abc_76628_new_n4949_));
AND2X2 AND2X2_1474 ( .A(u0__abc_76628_new_n4503__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4950_));
AND2X2 AND2X2_1475 ( .A(u0__abc_76628_new_n4562__bF_buf3), .B(u0_tms1_11_), .Y(u0__abc_76628_new_n4954_));
AND2X2 AND2X2_1476 ( .A(u0__abc_76628_new_n4547__bF_buf3), .B(u0_csc0_11_), .Y(u0__abc_76628_new_n4955_));
AND2X2 AND2X2_1477 ( .A(u0__abc_76628_new_n4517__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4956_));
AND2X2 AND2X2_1478 ( .A(u0__abc_76628_new_n4556__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4959_));
AND2X2 AND2X2_1479 ( .A(u0__abc_76628_new_n4528__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4960_));
AND2X2 AND2X2_148 ( .A(spec_req_cs_3_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1261_));
AND2X2 AND2X2_1480 ( .A(u0__abc_76628_new_n4531__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4962_));
AND2X2 AND2X2_1481 ( .A(u0__abc_76628_new_n4520__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4963_));
AND2X2 AND2X2_1482 ( .A(u0__abc_76628_new_n4500__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4966_));
AND2X2 AND2X2_1483 ( .A(u0__abc_76628_new_n4549__bF_buf3), .B(u0_tms0_11_), .Y(u0__abc_76628_new_n4967_));
AND2X2 AND2X2_1484 ( .A(u0__abc_76628_new_n4545__bF_buf3), .B(u0_csc1_11_), .Y(u0__abc_76628_new_n4969_));
AND2X2 AND2X2_1485 ( .A(u0__abc_76628_new_n4523__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n4970_));
AND2X2 AND2X2_1486 ( .A(u0__abc_76628_new_n4558__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4976_));
AND2X2 AND2X2_1487 ( .A(u0__abc_76628_new_n4554__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4977_));
AND2X2 AND2X2_1488 ( .A(u0__abc_76628_new_n4507__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4979_));
AND2X2 AND2X2_1489 ( .A(u0__abc_76628_new_n4510__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4980_));
AND2X2 AND2X2_149 ( .A(u0__abc_76628_new_n1262_), .B(u0__abc_76628_new_n1173__bF_buf2), .Y(u0__abc_76628_new_n1263_));
AND2X2 AND2X2_1490 ( .A(u0__abc_76628_new_n4566__bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_12_), .Y(u0__abc_76628_new_n4982_));
AND2X2 AND2X2_1491 ( .A(u0__abc_76628_new_n4503__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4983_));
AND2X2 AND2X2_1492 ( .A(u0__abc_76628_new_n4545__bF_buf2), .B(u0_csc1_12_), .Y(u0__abc_76628_new_n4987_));
AND2X2 AND2X2_1493 ( .A(u0__abc_76628_new_n4547__bF_buf2), .B(u0_csc0_12_), .Y(u0__abc_76628_new_n4988_));
AND2X2 AND2X2_1494 ( .A(u0__abc_76628_new_n4517__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4989_));
AND2X2 AND2X2_1495 ( .A(u0__abc_76628_new_n4531__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4992_));
AND2X2 AND2X2_1496 ( .A(u0__abc_76628_new_n4528__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4993_));
AND2X2 AND2X2_1497 ( .A(u0__abc_76628_new_n4556__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4995_));
AND2X2 AND2X2_1498 ( .A(u0__abc_76628_new_n4520__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4996_));
AND2X2 AND2X2_1499 ( .A(u0__abc_76628_new_n4500__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n4999_));
AND2X2 AND2X2_15 ( .A(_abc_85006_new_n281_), .B(_abc_85006_new_n282_), .Y(obct_cs_6_));
AND2X2 AND2X2_150 ( .A(spec_req_cs_2_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1264_));
AND2X2 AND2X2_1500 ( .A(u0__abc_76628_new_n4549__bF_buf2), .B(u0_tms0_12_), .Y(u0__abc_76628_new_n5000_));
AND2X2 AND2X2_1501 ( .A(u0__abc_76628_new_n4562__bF_buf2), .B(u0_tms1_12_), .Y(u0__abc_76628_new_n5002_));
AND2X2 AND2X2_1502 ( .A(u0__abc_76628_new_n4523__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5003_));
AND2X2 AND2X2_1503 ( .A(u0__abc_76628_new_n4510__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5009_));
AND2X2 AND2X2_1504 ( .A(u0__abc_76628_new_n4520__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5010_));
AND2X2 AND2X2_1505 ( .A(u0__abc_76628_new_n4549__bF_buf1), .B(u0_tms0_13_), .Y(u0__abc_76628_new_n5012_));
AND2X2 AND2X2_1506 ( .A(u0__abc_76628_new_n4517__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5013_));
AND2X2 AND2X2_1507 ( .A(u0__abc_76628_new_n4545__bF_buf1), .B(u0_csc1_13_), .Y(u0__abc_76628_new_n5015_));
AND2X2 AND2X2_1508 ( .A(u0__abc_76628_new_n4523__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5016_));
AND2X2 AND2X2_1509 ( .A(u0__abc_76628_new_n4562__bF_buf1), .B(u0_tms1_13_), .Y(u0__abc_76628_new_n5020_));
AND2X2 AND2X2_151 ( .A(u0__abc_76628_new_n1265_), .B(u0__abc_76628_new_n1172__bF_buf2), .Y(u0__abc_76628_new_n1266_));
AND2X2 AND2X2_1510 ( .A(u0__abc_76628_new_n4500__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5021_));
AND2X2 AND2X2_1511 ( .A(u0__abc_76628_new_n4531__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5022_));
AND2X2 AND2X2_1512 ( .A(u0__abc_76628_new_n4566__bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_13_), .Y(u0__abc_76628_new_n5025_));
AND2X2 AND2X2_1513 ( .A(u0__abc_76628_new_n4554__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5026_));
AND2X2 AND2X2_1514 ( .A(u0__abc_76628_new_n4507__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5028_));
AND2X2 AND2X2_1515 ( .A(u0__abc_76628_new_n4558__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5029_));
AND2X2 AND2X2_1516 ( .A(u0__abc_76628_new_n4547__bF_buf1), .B(u0_csc0_13_), .Y(u0__abc_76628_new_n5032_));
AND2X2 AND2X2_1517 ( .A(u0__abc_76628_new_n4528__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5033_));
AND2X2 AND2X2_1518 ( .A(u0__abc_76628_new_n4503__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5035_));
AND2X2 AND2X2_1519 ( .A(u0__abc_76628_new_n4556__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5036_));
AND2X2 AND2X2_152 ( .A(spec_req_cs_1_bF_buf5_), .B(u0_tms1_3_), .Y(u0__abc_76628_new_n1267_));
AND2X2 AND2X2_1520 ( .A(u0__abc_76628_new_n4510__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5042_));
AND2X2 AND2X2_1521 ( .A(u0__abc_76628_new_n4520__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5043_));
AND2X2 AND2X2_1522 ( .A(u0__abc_76628_new_n4549__bF_buf0), .B(u0_tms0_14_), .Y(u0__abc_76628_new_n5045_));
AND2X2 AND2X2_1523 ( .A(u0__abc_76628_new_n4517__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5046_));
AND2X2 AND2X2_1524 ( .A(u0__abc_76628_new_n4545__bF_buf0), .B(u0_csc1_14_), .Y(u0__abc_76628_new_n5048_));
AND2X2 AND2X2_1525 ( .A(u0__abc_76628_new_n4523__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5049_));
AND2X2 AND2X2_1526 ( .A(u0__abc_76628_new_n4503__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5053_));
AND2X2 AND2X2_1527 ( .A(u0__abc_76628_new_n4500__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5054_));
AND2X2 AND2X2_1528 ( .A(u0__abc_76628_new_n4547__bF_buf0), .B(u0_csc0_14_), .Y(u0__abc_76628_new_n5055_));
AND2X2 AND2X2_1529 ( .A(u0__abc_76628_new_n4566__bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_14_), .Y(u0__abc_76628_new_n5058_));
AND2X2 AND2X2_153 ( .A(u0__abc_76628_new_n1169__bF_buf2), .B(u0__abc_76628_new_n1270_), .Y(u0__abc_76628_new_n1271_));
AND2X2 AND2X2_1530 ( .A(u0__abc_76628_new_n4554__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5059_));
AND2X2 AND2X2_1531 ( .A(u0__abc_76628_new_n4507__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5061_));
AND2X2 AND2X2_1532 ( .A(u0__abc_76628_new_n4558__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5062_));
AND2X2 AND2X2_1533 ( .A(u0__abc_76628_new_n4531__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5065_));
AND2X2 AND2X2_1534 ( .A(u0__abc_76628_new_n4528__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5066_));
AND2X2 AND2X2_1535 ( .A(u0__abc_76628_new_n4556__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5068_));
AND2X2 AND2X2_1536 ( .A(u0__abc_76628_new_n4562__bF_buf0), .B(u0_tms1_14_), .Y(u0__abc_76628_new_n5069_));
AND2X2 AND2X2_1537 ( .A(u0__abc_76628_new_n4517__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5075_));
AND2X2 AND2X2_1538 ( .A(u0__abc_76628_new_n4528__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5076_));
AND2X2 AND2X2_1539 ( .A(u0__abc_76628_new_n4523__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5077_));
AND2X2 AND2X2_154 ( .A(u0__abc_76628_new_n1269_), .B(u0__abc_76628_new_n1271_), .Y(u0__abc_76628_new_n1272_));
AND2X2 AND2X2_1540 ( .A(u0__abc_76628_new_n4549__bF_buf4), .B(u0_tms0_15_), .Y(u0__abc_76628_new_n5080_));
AND2X2 AND2X2_1541 ( .A(u0__abc_76628_new_n4545__bF_buf4), .B(u0_csc1_15_), .Y(u0__abc_76628_new_n5081_));
AND2X2 AND2X2_1542 ( .A(u0__abc_76628_new_n4520__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5083_));
AND2X2 AND2X2_1543 ( .A(u0__abc_76628_new_n4562__bF_buf4), .B(u0_tms1_15_), .Y(u0__abc_76628_new_n5084_));
AND2X2 AND2X2_1544 ( .A(u0__abc_76628_new_n4531__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5088_));
AND2X2 AND2X2_1545 ( .A(u0__abc_76628_new_n4547__bF_buf4), .B(u0_csc0_15_), .Y(u0__abc_76628_new_n5089_));
AND2X2 AND2X2_1546 ( .A(u0__abc_76628_new_n4556__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5090_));
AND2X2 AND2X2_1547 ( .A(u0__abc_76628_new_n4554__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5091_));
AND2X2 AND2X2_1548 ( .A(u0__abc_76628_new_n4558__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5095_));
AND2X2 AND2X2_1549 ( .A(u0__abc_76628_new_n4507__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5096_));
AND2X2 AND2X2_155 ( .A(u0__abc_76628_new_n1170__bF_buf2), .B(sp_tms_4_), .Y(u0__abc_76628_new_n1274_));
AND2X2 AND2X2_1550 ( .A(u0__abc_76628_new_n4500__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5097_));
AND2X2 AND2X2_1551 ( .A(u0__abc_76628_new_n4503__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5100_));
AND2X2 AND2X2_1552 ( .A(u0__abc_76628_new_n4510__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5101_));
AND2X2 AND2X2_1553 ( .A(u0__abc_76628_new_n4566__bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_15_), .Y(u0__abc_76628_new_n5102_));
AND2X2 AND2X2_1554 ( .A(u0__abc_76628_new_n4507__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5108_));
AND2X2 AND2X2_1555 ( .A(u0__abc_76628_new_n4547__bF_buf3), .B(u0_csc0_16_), .Y(u0__abc_76628_new_n5109_));
AND2X2 AND2X2_1556 ( .A(u0__abc_76628_new_n4566__bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_16_), .Y(u0__abc_76628_new_n5111_));
AND2X2 AND2X2_1557 ( .A(u0__abc_76628_new_n4500__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5112_));
AND2X2 AND2X2_1558 ( .A(u0__abc_76628_new_n4510__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5114_));
AND2X2 AND2X2_1559 ( .A(u0__abc_76628_new_n4554__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5115_));
AND2X2 AND2X2_156 ( .A(spec_req_cs_5_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1275_));
AND2X2 AND2X2_1560 ( .A(u0__abc_76628_new_n4545__bF_buf3), .B(u0_csc1_16_), .Y(u0__abc_76628_new_n5119_));
AND2X2 AND2X2_1561 ( .A(u0__abc_76628_new_n4549__bF_buf3), .B(u0_tms0_16_), .Y(u0__abc_76628_new_n5120_));
AND2X2 AND2X2_1562 ( .A(u0__abc_76628_new_n4523__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5121_));
AND2X2 AND2X2_1563 ( .A(u0__abc_76628_new_n4531__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5124_));
AND2X2 AND2X2_1564 ( .A(u0__abc_76628_new_n4517__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5125_));
AND2X2 AND2X2_1565 ( .A(u0__abc_76628_new_n4503__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5127_));
AND2X2 AND2X2_1566 ( .A(u0__abc_76628_new_n4528__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5128_));
AND2X2 AND2X2_1567 ( .A(u0__abc_76628_new_n4558__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5131_));
AND2X2 AND2X2_1568 ( .A(u0__abc_76628_new_n4562__bF_buf3), .B(u0_tms1_16_), .Y(u0__abc_76628_new_n5132_));
AND2X2 AND2X2_1569 ( .A(u0__abc_76628_new_n4556__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5134_));
AND2X2 AND2X2_157 ( .A(u0__abc_76628_new_n1277_), .B(u0__abc_76628_new_n1179__bF_buf1), .Y(u0__abc_76628_new_n1278_));
AND2X2 AND2X2_1570 ( .A(u0__abc_76628_new_n4520__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5135_));
AND2X2 AND2X2_1571 ( .A(u0__abc_76628_new_n4503__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5141_));
AND2X2 AND2X2_1572 ( .A(u0__abc_76628_new_n4554__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5142_));
AND2X2 AND2X2_1573 ( .A(u0__abc_76628_new_n4507__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5144_));
AND2X2 AND2X2_1574 ( .A(u0__abc_76628_new_n4510__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5145_));
AND2X2 AND2X2_1575 ( .A(u0__abc_76628_new_n4566__bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_17_), .Y(u0__abc_76628_new_n5147_));
AND2X2 AND2X2_1576 ( .A(u0__abc_76628_new_n4558__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5148_));
AND2X2 AND2X2_1577 ( .A(u0__abc_76628_new_n4545__bF_buf2), .B(u0_csc1_17_), .Y(u0__abc_76628_new_n5152_));
AND2X2 AND2X2_1578 ( .A(u0__abc_76628_new_n4531__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5153_));
AND2X2 AND2X2_1579 ( .A(u0__abc_76628_new_n4517__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5154_));
AND2X2 AND2X2_158 ( .A(u0__abc_76628_new_n1278_), .B(u0__abc_76628_new_n1276_), .Y(u0__abc_76628_new_n1279_));
AND2X2 AND2X2_1580 ( .A(u0__abc_76628_new_n4547__bF_buf2), .B(u0_csc0_17_), .Y(u0__abc_76628_new_n5157_));
AND2X2 AND2X2_1581 ( .A(u0__abc_76628_new_n4528__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5158_));
AND2X2 AND2X2_1582 ( .A(u0__abc_76628_new_n4556__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5160_));
AND2X2 AND2X2_1583 ( .A(u0__abc_76628_new_n4520__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5161_));
AND2X2 AND2X2_1584 ( .A(u0__abc_76628_new_n4500__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5164_));
AND2X2 AND2X2_1585 ( .A(u0__abc_76628_new_n4549__bF_buf2), .B(u0_tms0_17_), .Y(u0__abc_76628_new_n5165_));
AND2X2 AND2X2_1586 ( .A(u0__abc_76628_new_n4562__bF_buf2), .B(u0_tms1_17_), .Y(u0__abc_76628_new_n5167_));
AND2X2 AND2X2_1587 ( .A(u0__abc_76628_new_n4523__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5168_));
AND2X2 AND2X2_1588 ( .A(u0__abc_76628_new_n4517__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5174_));
AND2X2 AND2X2_1589 ( .A(u0__abc_76628_new_n4528__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5175_));
AND2X2 AND2X2_159 ( .A(u0__abc_76628_new_n1280_), .B(u0__abc_76628_new_n1175__bF_buf1), .Y(u0__abc_76628_new_n1281_));
AND2X2 AND2X2_1590 ( .A(u0__abc_76628_new_n4523__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5176_));
AND2X2 AND2X2_1591 ( .A(u0__abc_76628_new_n4549__bF_buf1), .B(u0_tms0_18_), .Y(u0__abc_76628_new_n5179_));
AND2X2 AND2X2_1592 ( .A(u0__abc_76628_new_n4545__bF_buf1), .B(u0_csc1_18_), .Y(u0__abc_76628_new_n5180_));
AND2X2 AND2X2_1593 ( .A(u0__abc_76628_new_n4520__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5182_));
AND2X2 AND2X2_1594 ( .A(u0__abc_76628_new_n4562__bF_buf1), .B(u0_tms1_18_), .Y(u0__abc_76628_new_n5183_));
AND2X2 AND2X2_1595 ( .A(u0__abc_76628_new_n4531__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5187_));
AND2X2 AND2X2_1596 ( .A(u0__abc_76628_new_n4547__bF_buf1), .B(u0_csc0_18_), .Y(u0__abc_76628_new_n5188_));
AND2X2 AND2X2_1597 ( .A(u0__abc_76628_new_n4554__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5189_));
AND2X2 AND2X2_1598 ( .A(u0__abc_76628_new_n4556__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5190_));
AND2X2 AND2X2_1599 ( .A(u0__abc_76628_new_n4503__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5194_));
AND2X2 AND2X2_16 ( .A(_abc_85006_new_n284_), .B(_abc_85006_new_n285_), .Y(_abc_85006_new_n286_));
AND2X2 AND2X2_160 ( .A(spec_req_cs_4_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1282_));
AND2X2 AND2X2_1600 ( .A(u0__abc_76628_new_n4500__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5195_));
AND2X2 AND2X2_1601 ( .A(u0__abc_76628_new_n4507__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5196_));
AND2X2 AND2X2_1602 ( .A(u0__abc_76628_new_n4558__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5199_));
AND2X2 AND2X2_1603 ( .A(u0__abc_76628_new_n4510__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5200_));
AND2X2 AND2X2_1604 ( .A(u0__abc_76628_new_n4566__bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_18_), .Y(u0__abc_76628_new_n5201_));
AND2X2 AND2X2_1605 ( .A(u0__abc_76628_new_n4531__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5207_));
AND2X2 AND2X2_1606 ( .A(u0__abc_76628_new_n4554__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5208_));
AND2X2 AND2X2_1607 ( .A(u0__abc_76628_new_n4556__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5209_));
AND2X2 AND2X2_1608 ( .A(u0__abc_76628_new_n4547__bF_buf0), .B(u0_csc0_19_), .Y(u0__abc_76628_new_n5212_));
AND2X2 AND2X2_1609 ( .A(u0__abc_76628_new_n4562__bF_buf0), .B(u0_tms1_19_), .Y(u0__abc_76628_new_n5213_));
AND2X2 AND2X2_161 ( .A(u0__abc_76628_new_n1283_), .B(u0__abc_76628_new_n1174__bF_buf1), .Y(u0__abc_76628_new_n1284_));
AND2X2 AND2X2_1610 ( .A(u0__abc_76628_new_n4558__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5216_));
AND2X2 AND2X2_1611 ( .A(u0__abc_76628_new_n4507__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5217_));
AND2X2 AND2X2_1612 ( .A(u0__abc_76628_new_n4500__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5218_));
AND2X2 AND2X2_1613 ( .A(u0__abc_76628_new_n4503__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5221_));
AND2X2 AND2X2_1614 ( .A(u0__abc_76628_new_n4566__bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_19_), .Y(u0__abc_76628_new_n5222_));
AND2X2 AND2X2_1615 ( .A(u0__abc_76628_new_n4510__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5223_));
AND2X2 AND2X2_1616 ( .A(u0__abc_76628_new_n4517__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5227_));
AND2X2 AND2X2_1617 ( .A(u0__abc_76628_new_n4528__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5228_));
AND2X2 AND2X2_1618 ( .A(u0__abc_76628_new_n4523__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5229_));
AND2X2 AND2X2_1619 ( .A(u0__abc_76628_new_n4520__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5232_));
AND2X2 AND2X2_162 ( .A(spec_req_cs_3_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1285_));
AND2X2 AND2X2_1620 ( .A(u0__abc_76628_new_n4545__bF_buf0), .B(u0_csc1_19_), .Y(u0__abc_76628_new_n5233_));
AND2X2 AND2X2_1621 ( .A(u0__abc_76628_new_n4549__bF_buf0), .B(u0_tms0_19_), .Y(u0__abc_76628_new_n5234_));
AND2X2 AND2X2_1622 ( .A(u0__abc_76628_new_n4517__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5240_));
AND2X2 AND2X2_1623 ( .A(u0__abc_76628_new_n4528__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5241_));
AND2X2 AND2X2_1624 ( .A(u0__abc_76628_new_n4523__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5242_));
AND2X2 AND2X2_1625 ( .A(u0__abc_76628_new_n4549__bF_buf4), .B(u0_tms0_20_), .Y(u0__abc_76628_new_n5245_));
AND2X2 AND2X2_1626 ( .A(u0__abc_76628_new_n4545__bF_buf4), .B(u0_csc1_20_), .Y(u0__abc_76628_new_n5246_));
AND2X2 AND2X2_1627 ( .A(u0__abc_76628_new_n4520__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5248_));
AND2X2 AND2X2_1628 ( .A(u0__abc_76628_new_n4562__bF_buf4), .B(u0_tms1_20_), .Y(u0__abc_76628_new_n5249_));
AND2X2 AND2X2_1629 ( .A(u0__abc_76628_new_n4547__bF_buf4), .B(u0_csc0_20_), .Y(u0__abc_76628_new_n5253_));
AND2X2 AND2X2_163 ( .A(u0__abc_76628_new_n1286_), .B(u0__abc_76628_new_n1173__bF_buf1), .Y(u0__abc_76628_new_n1287_));
AND2X2 AND2X2_1630 ( .A(u0__abc_76628_new_n4531__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5254_));
AND2X2 AND2X2_1631 ( .A(u0__abc_76628_new_n4554__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5255_));
AND2X2 AND2X2_1632 ( .A(u0__abc_76628_new_n4556__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5256_));
AND2X2 AND2X2_1633 ( .A(u0__abc_76628_new_n4503__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5260_));
AND2X2 AND2X2_1634 ( .A(u0__abc_76628_new_n4500__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5261_));
AND2X2 AND2X2_1635 ( .A(u0__abc_76628_new_n4507__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5262_));
AND2X2 AND2X2_1636 ( .A(u0__abc_76628_new_n4558__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5265_));
AND2X2 AND2X2_1637 ( .A(u0__abc_76628_new_n4510__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5266_));
AND2X2 AND2X2_1638 ( .A(u0__abc_76628_new_n4566__bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_20_), .Y(u0__abc_76628_new_n5267_));
AND2X2 AND2X2_1639 ( .A(u0__abc_76628_new_n4510__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5273_));
AND2X2 AND2X2_164 ( .A(spec_req_cs_2_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1288_));
AND2X2 AND2X2_1640 ( .A(u0__abc_76628_new_n4562__bF_buf3), .B(u0_tms1_21_), .Y(u0__abc_76628_new_n5274_));
AND2X2 AND2X2_1641 ( .A(u0__abc_76628_new_n4549__bF_buf3), .B(u0_tms0_21_), .Y(u0__abc_76628_new_n5276_));
AND2X2 AND2X2_1642 ( .A(u0__abc_76628_new_n4517__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5277_));
AND2X2 AND2X2_1643 ( .A(u0__abc_76628_new_n4545__bF_buf3), .B(u0_csc1_21_), .Y(u0__abc_76628_new_n5279_));
AND2X2 AND2X2_1644 ( .A(u0__abc_76628_new_n4523__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5280_));
AND2X2 AND2X2_1645 ( .A(u0__abc_76628_new_n4503__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5284_));
AND2X2 AND2X2_1646 ( .A(u0__abc_76628_new_n4500__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5285_));
AND2X2 AND2X2_1647 ( .A(u0__abc_76628_new_n4547__bF_buf3), .B(u0_csc0_21_), .Y(u0__abc_76628_new_n5286_));
AND2X2 AND2X2_1648 ( .A(u0__abc_76628_new_n4566__bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_21_), .Y(u0__abc_76628_new_n5289_));
AND2X2 AND2X2_1649 ( .A(u0__abc_76628_new_n4554__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5290_));
AND2X2 AND2X2_165 ( .A(u0__abc_76628_new_n1289_), .B(u0__abc_76628_new_n1172__bF_buf1), .Y(u0__abc_76628_new_n1290_));
AND2X2 AND2X2_1650 ( .A(u0__abc_76628_new_n4507__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5292_));
AND2X2 AND2X2_1651 ( .A(u0__abc_76628_new_n4558__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5293_));
AND2X2 AND2X2_1652 ( .A(u0__abc_76628_new_n4531__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5296_));
AND2X2 AND2X2_1653 ( .A(u0__abc_76628_new_n4528__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5297_));
AND2X2 AND2X2_1654 ( .A(u0__abc_76628_new_n4556__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5299_));
AND2X2 AND2X2_1655 ( .A(u0__abc_76628_new_n4520__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5300_));
AND2X2 AND2X2_1656 ( .A(u0__abc_76628_new_n4558__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5306_));
AND2X2 AND2X2_1657 ( .A(u0__abc_76628_new_n4554__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5307_));
AND2X2 AND2X2_1658 ( .A(u0__abc_76628_new_n4507__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5309_));
AND2X2 AND2X2_1659 ( .A(u0__abc_76628_new_n4510__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5310_));
AND2X2 AND2X2_166 ( .A(spec_req_cs_1_bF_buf4_), .B(u0_tms1_4_), .Y(u0__abc_76628_new_n1291_));
AND2X2 AND2X2_1660 ( .A(u0__abc_76628_new_n4566__bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_22_), .Y(u0__abc_76628_new_n5312_));
AND2X2 AND2X2_1661 ( .A(u0__abc_76628_new_n4503__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5313_));
AND2X2 AND2X2_1662 ( .A(u0__abc_76628_new_n4562__bF_buf2), .B(u0_tms1_22_), .Y(u0__abc_76628_new_n5317_));
AND2X2 AND2X2_1663 ( .A(u0__abc_76628_new_n4547__bF_buf2), .B(u0_csc0_22_), .Y(u0__abc_76628_new_n5318_));
AND2X2 AND2X2_1664 ( .A(u0__abc_76628_new_n4517__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5319_));
AND2X2 AND2X2_1665 ( .A(u0__abc_76628_new_n4556__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5322_));
AND2X2 AND2X2_1666 ( .A(u0__abc_76628_new_n4528__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5323_));
AND2X2 AND2X2_1667 ( .A(u0__abc_76628_new_n4531__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5325_));
AND2X2 AND2X2_1668 ( .A(u0__abc_76628_new_n4520__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5326_));
AND2X2 AND2X2_1669 ( .A(u0__abc_76628_new_n4500__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5329_));
AND2X2 AND2X2_167 ( .A(u0__abc_76628_new_n1169__bF_buf1), .B(u0__abc_76628_new_n1294_), .Y(u0__abc_76628_new_n1295_));
AND2X2 AND2X2_1670 ( .A(u0__abc_76628_new_n4549__bF_buf2), .B(u0_tms0_22_), .Y(u0__abc_76628_new_n5330_));
AND2X2 AND2X2_1671 ( .A(u0__abc_76628_new_n4545__bF_buf2), .B(u0_csc1_22_), .Y(u0__abc_76628_new_n5332_));
AND2X2 AND2X2_1672 ( .A(u0__abc_76628_new_n4523__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5333_));
AND2X2 AND2X2_1673 ( .A(u0__abc_76628_new_n4507__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5339_));
AND2X2 AND2X2_1674 ( .A(u0__abc_76628_new_n4547__bF_buf1), .B(u0_csc0_23_), .Y(u0__abc_76628_new_n5340_));
AND2X2 AND2X2_1675 ( .A(u0__abc_76628_new_n4566__bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_23_), .Y(u0__abc_76628_new_n5342_));
AND2X2 AND2X2_1676 ( .A(u0__abc_76628_new_n4500__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5343_));
AND2X2 AND2X2_1677 ( .A(u0__abc_76628_new_n4510__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5345_));
AND2X2 AND2X2_1678 ( .A(u0__abc_76628_new_n4554__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5346_));
AND2X2 AND2X2_1679 ( .A(u0__abc_76628_new_n4545__bF_buf1), .B(u0_csc1_23_), .Y(u0__abc_76628_new_n5350_));
AND2X2 AND2X2_168 ( .A(u0__abc_76628_new_n1293_), .B(u0__abc_76628_new_n1295_), .Y(u0__abc_76628_new_n1296_));
AND2X2 AND2X2_1680 ( .A(u0__abc_76628_new_n4549__bF_buf1), .B(u0_tms0_23_), .Y(u0__abc_76628_new_n5351_));
AND2X2 AND2X2_1681 ( .A(u0__abc_76628_new_n4523__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5352_));
AND2X2 AND2X2_1682 ( .A(u0__abc_76628_new_n4531__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5355_));
AND2X2 AND2X2_1683 ( .A(u0__abc_76628_new_n4517__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5356_));
AND2X2 AND2X2_1684 ( .A(u0__abc_76628_new_n4503__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5358_));
AND2X2 AND2X2_1685 ( .A(u0__abc_76628_new_n4528__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5359_));
AND2X2 AND2X2_1686 ( .A(u0__abc_76628_new_n4558__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5362_));
AND2X2 AND2X2_1687 ( .A(u0__abc_76628_new_n4562__bF_buf1), .B(u0_tms1_23_), .Y(u0__abc_76628_new_n5363_));
AND2X2 AND2X2_1688 ( .A(u0__abc_76628_new_n4556__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5365_));
AND2X2 AND2X2_1689 ( .A(u0__abc_76628_new_n4520__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5366_));
AND2X2 AND2X2_169 ( .A(u0__abc_76628_new_n1170__bF_buf1), .B(sp_tms_5_), .Y(u0__abc_76628_new_n1298_));
AND2X2 AND2X2_1690 ( .A(u0__abc_76628_new_n4545__bF_buf0), .B(u0_csc1_24_), .Y(u0__abc_76628_new_n5372_));
AND2X2 AND2X2_1691 ( .A(u0__abc_76628_new_n4556__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5373_));
AND2X2 AND2X2_1692 ( .A(u0__abc_76628_new_n4549__bF_buf0), .B(u0_tms0_24_), .Y(u0__abc_76628_new_n5375_));
AND2X2 AND2X2_1693 ( .A(u0__abc_76628_new_n4507__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5376_));
AND2X2 AND2X2_1694 ( .A(u0__abc_76628_new_n4562__bF_buf0), .B(u0_tms1_24_), .Y(u0__abc_76628_new_n5378_));
AND2X2 AND2X2_1695 ( .A(u0__abc_76628_new_n4503__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5379_));
AND2X2 AND2X2_1696 ( .A(u0__abc_76628_new_n4500__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5383_));
AND2X2 AND2X2_1697 ( .A(u0__abc_76628_new_n4558__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5384_));
AND2X2 AND2X2_1698 ( .A(u0__abc_76628_new_n4510__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5386_));
AND2X2 AND2X2_1699 ( .A(u0__abc_76628_new_n4531__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5387_));
AND2X2 AND2X2_17 ( .A(_abc_85006_new_n287_), .B(_abc_85006_new_n288_), .Y(obct_cs_7_));
AND2X2 AND2X2_170 ( .A(spec_req_cs_5_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1299_));
AND2X2 AND2X2_1700 ( .A(u0__abc_76628_new_n4517__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5390_));
AND2X2 AND2X2_1701 ( .A(u0__abc_76628_new_n4528__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5391_));
AND2X2 AND2X2_1702 ( .A(u0__abc_76628_new_n4566__bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_24_), .Y(u0__abc_76628_new_n5393_));
AND2X2 AND2X2_1703 ( .A(u0__abc_76628_new_n4554__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5394_));
AND2X2 AND2X2_1704 ( .A(u0__abc_76628_new_n4541__bF_buf0), .B(rfr_ps_val_0_), .Y(u0__abc_76628_new_n5398_));
AND2X2 AND2X2_1705 ( .A(u0__abc_76628_new_n4547__bF_buf0), .B(u0_csc0_24_), .Y(u0__abc_76628_new_n5399_));
AND2X2 AND2X2_1706 ( .A(u0__abc_76628_new_n4520__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5400_));
AND2X2 AND2X2_1707 ( .A(u0__abc_76628_new_n4523__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5401_));
AND2X2 AND2X2_1708 ( .A(u0__abc_76628_new_n4566__bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_25_), .Y(u0__abc_76628_new_n5407_));
AND2X2 AND2X2_1709 ( .A(u0__abc_76628_new_n4510__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5408_));
AND2X2 AND2X2_171 ( .A(u0__abc_76628_new_n1301_), .B(u0__abc_76628_new_n1179__bF_buf0), .Y(u0__abc_76628_new_n1302_));
AND2X2 AND2X2_1710 ( .A(u0__abc_76628_new_n4523__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5410_));
AND2X2 AND2X2_1711 ( .A(u0__abc_76628_new_n4517__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5411_));
AND2X2 AND2X2_1712 ( .A(u0__abc_76628_new_n4547__bF_buf4), .B(u0_csc0_25_), .Y(u0__abc_76628_new_n5413_));
AND2X2 AND2X2_1713 ( .A(u0__abc_76628_new_n4528__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5414_));
AND2X2 AND2X2_1714 ( .A(u0__abc_76628_new_n4562__bF_buf4), .B(u0_tms1_25_), .Y(u0__abc_76628_new_n5418_));
AND2X2 AND2X2_1715 ( .A(u0__abc_76628_new_n4520__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5419_));
AND2X2 AND2X2_1716 ( .A(u0__abc_76628_new_n4549__bF_buf4), .B(u0_tms0_25_), .Y(u0__abc_76628_new_n5421_));
AND2X2 AND2X2_1717 ( .A(u0__abc_76628_new_n4503__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5422_));
AND2X2 AND2X2_1718 ( .A(u0__abc_76628_new_n4500__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5425_));
AND2X2 AND2X2_1719 ( .A(u0__abc_76628_new_n4556__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5426_));
AND2X2 AND2X2_172 ( .A(u0__abc_76628_new_n1302_), .B(u0__abc_76628_new_n1300_), .Y(u0__abc_76628_new_n1303_));
AND2X2 AND2X2_1720 ( .A(u0__abc_76628_new_n4545__bF_buf4), .B(u0_csc1_25_), .Y(u0__abc_76628_new_n5428_));
AND2X2 AND2X2_1721 ( .A(u0__abc_76628_new_n4531__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5429_));
AND2X2 AND2X2_1722 ( .A(u0__abc_76628_new_n4541__bF_buf3), .B(rfr_ps_val_1_), .Y(u0__abc_76628_new_n5433_));
AND2X2 AND2X2_1723 ( .A(u0__abc_76628_new_n4558__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5434_));
AND2X2 AND2X2_1724 ( .A(u0__abc_76628_new_n4507__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5435_));
AND2X2 AND2X2_1725 ( .A(u0__abc_76628_new_n4554__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5436_));
AND2X2 AND2X2_1726 ( .A(u0__abc_76628_new_n4554__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5442_));
AND2X2 AND2X2_1727 ( .A(u0__abc_76628_new_n4531__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5443_));
AND2X2 AND2X2_1728 ( .A(u0__abc_76628_new_n4556__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5444_));
AND2X2 AND2X2_1729 ( .A(u0__abc_76628_new_n4558__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5447_));
AND2X2 AND2X2_173 ( .A(u0__abc_76628_new_n1304_), .B(u0__abc_76628_new_n1175__bF_buf0), .Y(u0__abc_76628_new_n1305_));
AND2X2 AND2X2_1730 ( .A(u0__abc_76628_new_n4507__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5448_));
AND2X2 AND2X2_1731 ( .A(u0__abc_76628_new_n4500__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5449_));
AND2X2 AND2X2_1732 ( .A(u0__abc_76628_new_n4541__bF_buf2), .B(rfr_ps_val_2_), .Y(u0__abc_76628_new_n5453_));
AND2X2 AND2X2_1733 ( .A(u0__abc_76628_new_n4520__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5454_));
AND2X2 AND2X2_1734 ( .A(u0__abc_76628_new_n4549__bF_buf3), .B(u0_tms0_26_), .Y(u0__abc_76628_new_n5455_));
AND2X2 AND2X2_1735 ( .A(u0__abc_76628_new_n4545__bF_buf3), .B(u0_csc1_26_), .Y(u0__abc_76628_new_n5456_));
AND2X2 AND2X2_1736 ( .A(u0__abc_76628_new_n4562__bF_buf3), .B(u0_tms1_26_), .Y(u0__abc_76628_new_n5461_));
AND2X2 AND2X2_1737 ( .A(u0__abc_76628_new_n4566__bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_26_), .Y(u0__abc_76628_new_n5462_));
AND2X2 AND2X2_1738 ( .A(u0__abc_76628_new_n4547__bF_buf3), .B(u0_csc0_26_), .Y(u0__abc_76628_new_n5463_));
AND2X2 AND2X2_1739 ( .A(u0__abc_76628_new_n4510__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5466_));
AND2X2 AND2X2_174 ( .A(spec_req_cs_4_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1306_));
AND2X2 AND2X2_1740 ( .A(u0__abc_76628_new_n4517__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5467_));
AND2X2 AND2X2_1741 ( .A(u0__abc_76628_new_n4523__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5468_));
AND2X2 AND2X2_1742 ( .A(u0__abc_76628_new_n4528__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5471_));
AND2X2 AND2X2_1743 ( .A(u0__abc_76628_new_n4503__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5472_));
AND2X2 AND2X2_1744 ( .A(u0__abc_76628_new_n4510__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5477_));
AND2X2 AND2X2_1745 ( .A(u0__abc_76628_new_n4556__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5478_));
AND2X2 AND2X2_1746 ( .A(u0__abc_76628_new_n4500__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5480_));
AND2X2 AND2X2_1747 ( .A(u0__abc_76628_new_n4558__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5481_));
AND2X2 AND2X2_1748 ( .A(u0__abc_76628_new_n4520__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5483_));
AND2X2 AND2X2_1749 ( .A(u0__abc_76628_new_n4503__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5484_));
AND2X2 AND2X2_175 ( .A(u0__abc_76628_new_n1307_), .B(u0__abc_76628_new_n1174__bF_buf0), .Y(u0__abc_76628_new_n1308_));
AND2X2 AND2X2_1750 ( .A(u0__abc_76628_new_n4549__bF_buf2), .B(u0_tms0_27_), .Y(u0__abc_76628_new_n5488_));
AND2X2 AND2X2_1751 ( .A(u0__abc_76628_new_n4562__bF_buf2), .B(u0_tms1_27_), .Y(u0__abc_76628_new_n5489_));
AND2X2 AND2X2_1752 ( .A(u0__abc_76628_new_n4523__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5491_));
AND2X2 AND2X2_1753 ( .A(u0__abc_76628_new_n4528__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5492_));
AND2X2 AND2X2_1754 ( .A(u0__abc_76628_new_n4517__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5495_));
AND2X2 AND2X2_1755 ( .A(u0__abc_76628_new_n4507__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5496_));
AND2X2 AND2X2_1756 ( .A(u0__abc_76628_new_n4566__bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_27_), .Y(u0__abc_76628_new_n5498_));
AND2X2 AND2X2_1757 ( .A(u0__abc_76628_new_n4545__bF_buf2), .B(u0_csc1_27_), .Y(u0__abc_76628_new_n5499_));
AND2X2 AND2X2_1758 ( .A(u0__abc_76628_new_n4541__bF_buf1), .B(rfr_ps_val_3_), .Y(u0__abc_76628_new_n5503_));
AND2X2 AND2X2_1759 ( .A(u0__abc_76628_new_n4531__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5504_));
AND2X2 AND2X2_176 ( .A(spec_req_cs_3_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1309_));
AND2X2 AND2X2_1760 ( .A(u0__abc_76628_new_n4547__bF_buf2), .B(u0_csc0_27_), .Y(u0__abc_76628_new_n5505_));
AND2X2 AND2X2_1761 ( .A(u0__abc_76628_new_n4554__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n5506_));
AND2X2 AND2X2_1762 ( .A(u0__abc_76628_new_n4554__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5512_));
AND2X2 AND2X2_1763 ( .A(u0__abc_76628_new_n4531__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5513_));
AND2X2 AND2X2_1764 ( .A(u0__abc_76628_new_n4556__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5514_));
AND2X2 AND2X2_1765 ( .A(u0__abc_76628_new_n4558__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5517_));
AND2X2 AND2X2_1766 ( .A(u0__abc_76628_new_n4507__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5518_));
AND2X2 AND2X2_1767 ( .A(u0__abc_76628_new_n4500__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5519_));
AND2X2 AND2X2_1768 ( .A(u0__abc_76628_new_n4541__bF_buf0), .B(rfr_ps_val_4_), .Y(u0__abc_76628_new_n5523_));
AND2X2 AND2X2_1769 ( .A(u0__abc_76628_new_n4562__bF_buf1), .B(u0_tms1_28_), .Y(u0__abc_76628_new_n5524_));
AND2X2 AND2X2_177 ( .A(u0__abc_76628_new_n1310_), .B(u0__abc_76628_new_n1173__bF_buf0), .Y(u0__abc_76628_new_n1311_));
AND2X2 AND2X2_1770 ( .A(u0__abc_76628_new_n4549__bF_buf1), .B(u0_tms0_28_), .Y(u0__abc_76628_new_n5525_));
AND2X2 AND2X2_1771 ( .A(u0__abc_76628_new_n4545__bF_buf1), .B(u0_csc1_28_), .Y(u0__abc_76628_new_n5526_));
AND2X2 AND2X2_1772 ( .A(u0__abc_76628_new_n4520__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5531_));
AND2X2 AND2X2_1773 ( .A(u0__abc_76628_new_n4566__bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_28_), .Y(u0__abc_76628_new_n5532_));
AND2X2 AND2X2_1774 ( .A(u0__abc_76628_new_n4547__bF_buf1), .B(u0_csc0_28_), .Y(u0__abc_76628_new_n5533_));
AND2X2 AND2X2_1775 ( .A(u0__abc_76628_new_n4510__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5536_));
AND2X2 AND2X2_1776 ( .A(u0__abc_76628_new_n4517__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5537_));
AND2X2 AND2X2_1777 ( .A(u0__abc_76628_new_n4523__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5538_));
AND2X2 AND2X2_1778 ( .A(u0__abc_76628_new_n4528__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5541_));
AND2X2 AND2X2_1779 ( .A(u0__abc_76628_new_n4503__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n5542_));
AND2X2 AND2X2_178 ( .A(spec_req_cs_2_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1312_));
AND2X2 AND2X2_1780 ( .A(u0__abc_76628_new_n4547__bF_buf0), .B(u0_csc0_29_), .Y(u0__abc_76628_new_n5547_));
AND2X2 AND2X2_1781 ( .A(u0__abc_76628_new_n4517__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5548_));
AND2X2 AND2X2_1782 ( .A(u0__abc_76628_new_n4566__bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_29_), .Y(u0__abc_76628_new_n5550_));
AND2X2 AND2X2_1783 ( .A(u0__abc_76628_new_n4510__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5551_));
AND2X2 AND2X2_1784 ( .A(u0__abc_76628_new_n4549__bF_buf0), .B(u0_tms0_29_), .Y(u0__abc_76628_new_n5553_));
AND2X2 AND2X2_1785 ( .A(u0__abc_76628_new_n4523__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5554_));
AND2X2 AND2X2_1786 ( .A(u0__abc_76628_new_n4545__bF_buf0), .B(u0_csc1_29_), .Y(u0__abc_76628_new_n5558_));
AND2X2 AND2X2_1787 ( .A(u0__abc_76628_new_n4558__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5559_));
AND2X2 AND2X2_1788 ( .A(u0__abc_76628_new_n4562__bF_buf0), .B(u0_tms1_29_), .Y(u0__abc_76628_new_n5561_));
AND2X2 AND2X2_1789 ( .A(u0__abc_76628_new_n4520__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5562_));
AND2X2 AND2X2_179 ( .A(u0__abc_76628_new_n1313_), .B(u0__abc_76628_new_n1172__bF_buf0), .Y(u0__abc_76628_new_n1314_));
AND2X2 AND2X2_1790 ( .A(u0__abc_76628_new_n4500__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5565_));
AND2X2 AND2X2_1791 ( .A(u0__abc_76628_new_n4556__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5566_));
AND2X2 AND2X2_1792 ( .A(u0__abc_76628_new_n4528__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5568_));
AND2X2 AND2X2_1793 ( .A(u0__abc_76628_new_n4531__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5569_));
AND2X2 AND2X2_1794 ( .A(u0__abc_76628_new_n4541__bF_buf3), .B(rfr_ps_val_5_), .Y(u0__abc_76628_new_n5573_));
AND2X2 AND2X2_1795 ( .A(u0__abc_76628_new_n4507__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5574_));
AND2X2 AND2X2_1796 ( .A(u0__abc_76628_new_n4503__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5575_));
AND2X2 AND2X2_1797 ( .A(u0__abc_76628_new_n4554__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n5576_));
AND2X2 AND2X2_1798 ( .A(u0__abc_76628_new_n4547__bF_buf4), .B(u0_csc0_30_), .Y(u0__abc_76628_new_n5582_));
AND2X2 AND2X2_1799 ( .A(u0__abc_76628_new_n4517__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5583_));
AND2X2 AND2X2_18 ( .A(_abc_85006_new_n290_), .B(_abc_85006_new_n291_), .Y(tms_s_0_));
AND2X2 AND2X2_180 ( .A(spec_req_cs_1_bF_buf3_), .B(u0_tms1_5_), .Y(u0__abc_76628_new_n1315_));
AND2X2 AND2X2_1800 ( .A(u0__abc_76628_new_n4566__bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_30_), .Y(u0__abc_76628_new_n5585_));
AND2X2 AND2X2_1801 ( .A(u0__abc_76628_new_n4510__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5586_));
AND2X2 AND2X2_1802 ( .A(u0__abc_76628_new_n4549__bF_buf4), .B(u0_tms0_30_), .Y(u0__abc_76628_new_n5588_));
AND2X2 AND2X2_1803 ( .A(u0__abc_76628_new_n4523__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5589_));
AND2X2 AND2X2_1804 ( .A(u0__abc_76628_new_n4545__bF_buf4), .B(u0_csc1_30_), .Y(u0__abc_76628_new_n5593_));
AND2X2 AND2X2_1805 ( .A(u0__abc_76628_new_n4558__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5594_));
AND2X2 AND2X2_1806 ( .A(u0__abc_76628_new_n4562__bF_buf4), .B(u0_tms1_30_), .Y(u0__abc_76628_new_n5596_));
AND2X2 AND2X2_1807 ( .A(u0__abc_76628_new_n4520__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5597_));
AND2X2 AND2X2_1808 ( .A(u0__abc_76628_new_n4500__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5600_));
AND2X2 AND2X2_1809 ( .A(u0__abc_76628_new_n4556__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5601_));
AND2X2 AND2X2_181 ( .A(u0__abc_76628_new_n1169__bF_buf0), .B(u0__abc_76628_new_n1318_), .Y(u0__abc_76628_new_n1319_));
AND2X2 AND2X2_1810 ( .A(u0__abc_76628_new_n4528__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5603_));
AND2X2 AND2X2_1811 ( .A(u0__abc_76628_new_n4531__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5604_));
AND2X2 AND2X2_1812 ( .A(u0__abc_76628_new_n4541__bF_buf2), .B(rfr_ps_val_6_), .Y(u0__abc_76628_new_n5608_));
AND2X2 AND2X2_1813 ( .A(u0__abc_76628_new_n4507__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5609_));
AND2X2 AND2X2_1814 ( .A(u0__abc_76628_new_n4503__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5610_));
AND2X2 AND2X2_1815 ( .A(u0__abc_76628_new_n4554__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n5611_));
AND2X2 AND2X2_1816 ( .A(u0__abc_76628_new_n4547__bF_buf3), .B(u0_csc0_31_), .Y(u0__abc_76628_new_n5617_));
AND2X2 AND2X2_1817 ( .A(u0__abc_76628_new_n4517__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5618_));
AND2X2 AND2X2_1818 ( .A(u0__abc_76628_new_n4566__bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_31_), .Y(u0__abc_76628_new_n5620_));
AND2X2 AND2X2_1819 ( .A(u0__abc_76628_new_n4528__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5621_));
AND2X2 AND2X2_182 ( .A(u0__abc_76628_new_n1317_), .B(u0__abc_76628_new_n1319_), .Y(u0__abc_76628_new_n1320_));
AND2X2 AND2X2_1820 ( .A(u0__abc_76628_new_n4549__bF_buf3), .B(u0_tms0_31_), .Y(u0__abc_76628_new_n5623_));
AND2X2 AND2X2_1821 ( .A(u0__abc_76628_new_n4523__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5624_));
AND2X2 AND2X2_1822 ( .A(u0__abc_76628_new_n4545__bF_buf3), .B(u0_csc1_31_), .Y(u0__abc_76628_new_n5628_));
AND2X2 AND2X2_1823 ( .A(u0__abc_76628_new_n4558__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5629_));
AND2X2 AND2X2_1824 ( .A(u0__abc_76628_new_n4562__bF_buf3), .B(u0_tms1_31_), .Y(u0__abc_76628_new_n5631_));
AND2X2 AND2X2_1825 ( .A(u0__abc_76628_new_n4520__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5632_));
AND2X2 AND2X2_1826 ( .A(u0__abc_76628_new_n4503__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5635_));
AND2X2 AND2X2_1827 ( .A(u0__abc_76628_new_n4556__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5636_));
AND2X2 AND2X2_1828 ( .A(u0__abc_76628_new_n4510__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5638_));
AND2X2 AND2X2_1829 ( .A(u0__abc_76628_new_n4531__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5639_));
AND2X2 AND2X2_183 ( .A(u0__abc_76628_new_n1170__bF_buf0), .B(sp_tms_6_), .Y(u0__abc_76628_new_n1322_));
AND2X2 AND2X2_1830 ( .A(u0__abc_76628_new_n4541__bF_buf1), .B(rfr_ps_val_7_), .Y(u0__abc_76628_new_n5643_));
AND2X2 AND2X2_1831 ( .A(u0__abc_76628_new_n4507__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5644_));
AND2X2 AND2X2_1832 ( .A(u0__abc_76628_new_n4500__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5645_));
AND2X2 AND2X2_1833 ( .A(u0__abc_76628_new_n4554__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n5646_));
AND2X2 AND2X2_1834 ( .A(\wb_addr_i[30] ), .B(\wb_addr_i[29] ), .Y(u0__abc_76628_new_n5653_));
AND2X2 AND2X2_1835 ( .A(u0__abc_76628_new_n5653_), .B(u0__abc_76628_new_n5652_), .Y(u0__abc_76628_new_n5654_));
AND2X2 AND2X2_1836 ( .A(u0__abc_76628_new_n5654_), .B(u0__abc_76628_new_n1168_), .Y(u0__abc_76628_new_n5655_));
AND2X2 AND2X2_1837 ( .A(u0__abc_76628_new_n4397_), .B(wb_we_i), .Y(u0__abc_76628_new_n5656_));
AND2X2 AND2X2_1838 ( .A(u0__abc_76628_new_n5655_), .B(u0__abc_76628_new_n5656_), .Y(u0__0rf_we_0_0_));
AND2X2 AND2X2_1839 ( .A(u0__abc_76628_new_n5660_), .B(u0__abc_76628_new_n5661_), .Y(u0__abc_76628_new_n5662_));
AND2X2 AND2X2_184 ( .A(spec_req_cs_5_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1323_));
AND2X2 AND2X2_1840 ( .A(u0__abc_76628_new_n5663_), .B(u0_csc0_0_), .Y(u0__abc_76628_new_n5664_));
AND2X2 AND2X2_1841 ( .A(u0__abc_76628_new_n5662_), .B(u0__abc_76628_new_n5664_), .Y(cs_need_rfr_0_));
AND2X2 AND2X2_1842 ( .A(u0__abc_76628_new_n5666_), .B(u0__abc_76628_new_n5667_), .Y(u0__abc_76628_new_n5668_));
AND2X2 AND2X2_1843 ( .A(u0__abc_76628_new_n5669_), .B(u0_csc1_0_), .Y(u0__abc_76628_new_n5670_));
AND2X2 AND2X2_1844 ( .A(u0__abc_76628_new_n5668_), .B(u0__abc_76628_new_n5670_), .Y(cs_need_rfr_1_));
AND2X2 AND2X2_1845 ( .A(u0__abc_76628_new_n5672_), .B(u0__abc_76628_new_n5673_), .Y(u0__abc_76628_new_n5674_));
AND2X2 AND2X2_1846 ( .A(u0__abc_76628_new_n5675_), .B(1'h0), .Y(u0__abc_76628_new_n5676_));
AND2X2 AND2X2_1847 ( .A(u0__abc_76628_new_n5674_), .B(u0__abc_76628_new_n5676_), .Y(cs_need_rfr_2_));
AND2X2 AND2X2_1848 ( .A(u0__abc_76628_new_n5678_), .B(u0__abc_76628_new_n5679_), .Y(u0__abc_76628_new_n5680_));
AND2X2 AND2X2_1849 ( .A(u0__abc_76628_new_n5681_), .B(1'h0), .Y(u0__abc_76628_new_n5682_));
AND2X2 AND2X2_185 ( .A(u0__abc_76628_new_n1325_), .B(u0__abc_76628_new_n1179__bF_buf5), .Y(u0__abc_76628_new_n1326_));
AND2X2 AND2X2_1850 ( .A(u0__abc_76628_new_n5680_), .B(u0__abc_76628_new_n5682_), .Y(cs_need_rfr_3_));
AND2X2 AND2X2_1851 ( .A(u0__abc_76628_new_n5684_), .B(u0__abc_76628_new_n5685_), .Y(u0__abc_76628_new_n5686_));
AND2X2 AND2X2_1852 ( .A(u0__abc_76628_new_n5687_), .B(1'h0), .Y(u0__abc_76628_new_n5688_));
AND2X2 AND2X2_1853 ( .A(u0__abc_76628_new_n5686_), .B(u0__abc_76628_new_n5688_), .Y(cs_need_rfr_4_));
AND2X2 AND2X2_1854 ( .A(u0__abc_76628_new_n5690_), .B(u0__abc_76628_new_n5691_), .Y(u0__abc_76628_new_n5692_));
AND2X2 AND2X2_1855 ( .A(u0__abc_76628_new_n5693_), .B(1'h0), .Y(u0__abc_76628_new_n5694_));
AND2X2 AND2X2_1856 ( .A(u0__abc_76628_new_n5692_), .B(u0__abc_76628_new_n5694_), .Y(cs_need_rfr_5_));
AND2X2 AND2X2_1857 ( .A(u0__abc_76628_new_n5696_), .B(u0__abc_76628_new_n5697_), .Y(u0__abc_76628_new_n5698_));
AND2X2 AND2X2_1858 ( .A(u0__abc_76628_new_n5699_), .B(1'h0), .Y(u0__abc_76628_new_n5700_));
AND2X2 AND2X2_1859 ( .A(u0__abc_76628_new_n5698_), .B(u0__abc_76628_new_n5700_), .Y(cs_need_rfr_6_));
AND2X2 AND2X2_186 ( .A(u0__abc_76628_new_n1326_), .B(u0__abc_76628_new_n1324_), .Y(u0__abc_76628_new_n1327_));
AND2X2 AND2X2_1860 ( .A(u0__abc_76628_new_n5702_), .B(u0__abc_76628_new_n5703_), .Y(u0__abc_76628_new_n5704_));
AND2X2 AND2X2_1861 ( .A(u0__abc_76628_new_n5705_), .B(1'h0), .Y(u0__abc_76628_new_n5706_));
AND2X2 AND2X2_1862 ( .A(u0__abc_76628_new_n5704_), .B(u0__abc_76628_new_n5706_), .Y(cs_need_rfr_7_));
AND2X2 AND2X2_1863 ( .A(u0__abc_76628_new_n5708_), .B(u0_lmr_ack_r), .Y(u0__abc_76628_new_n5709_));
AND2X2 AND2X2_1864 ( .A(u0__abc_76628_new_n5710_), .B(u0_init_ack_r), .Y(u0__abc_76628_new_n5711_));
AND2X2 AND2X2_1865 ( .A(u0__abc_76628_new_n1100_), .B(u0__abc_76628_new_n5712_), .Y(u0__abc_76628_new_n5713_));
AND2X2 AND2X2_1866 ( .A(u0__abc_76628_new_n5709_), .B(spec_req_cs_0_bF_buf1_), .Y(u0_lmr_ack0));
AND2X2 AND2X2_1867 ( .A(u0__abc_76628_new_n5709_), .B(spec_req_cs_1_bF_buf1_), .Y(u0_lmr_ack1));
AND2X2 AND2X2_1868 ( .A(u0__abc_76628_new_n5711_), .B(spec_req_cs_0_bF_buf0_), .Y(u0_init_ack0));
AND2X2 AND2X2_1869 ( .A(u0__abc_76628_new_n5711_), .B(spec_req_cs_1_bF_buf0_), .Y(u0_init_ack1));
AND2X2 AND2X2_187 ( .A(u0__abc_76628_new_n1328_), .B(u0__abc_76628_new_n1175__bF_buf5), .Y(u0__abc_76628_new_n1329_));
AND2X2 AND2X2_1870 ( .A(u0_u0__abc_72207_new_n207_), .B(u0_u0_lmr_req_we), .Y(u0_u0__abc_72207_new_n208_));
AND2X2 AND2X2_1871 ( .A(u0_u0__abc_72207_new_n208_), .B(u0_u0_inited), .Y(u0_u0__abc_72207_new_n209_));
AND2X2 AND2X2_1872 ( .A(u0_u0__abc_72207_new_n211_), .B(u0_lmr_req0), .Y(u0_u0__abc_72207_new_n212_));
AND2X2 AND2X2_1873 ( .A(u0_u0__abc_72207_new_n210_), .B(u0_u0__abc_72207_new_n212_), .Y(u0_u0__abc_72207_new_n213_));
AND2X2 AND2X2_1874 ( .A(u0_u0__abc_72207_new_n215_), .B(u0_rf_we), .Y(u0_u0__abc_72207_new_n216_));
AND2X2 AND2X2_1875 ( .A(u0_u0__abc_72207_new_n218_), .B(u0_u0_addr_r_4_), .Y(u0_u0__abc_72207_new_n219_));
AND2X2 AND2X2_1876 ( .A(u0_u0__abc_72207_new_n219_), .B(u0_u0__abc_72207_new_n217_), .Y(u0_u0__abc_72207_new_n220_));
AND2X2 AND2X2_1877 ( .A(u0_u0__abc_72207_new_n220_), .B(u0_u0__abc_72207_new_n216_), .Y(u0_u0__abc_72207_new_n221_));
AND2X2 AND2X2_1878 ( .A(u0_u0__abc_72207_new_n221_), .B(u0_u0_addr_r_2_), .Y(u0_u0__0lmr_req_we_0_0_));
AND2X2 AND2X2_1879 ( .A(u0_u0__abc_72207_new_n225_), .B(u0_u0__abc_72207_new_n223_), .Y(u0_u0__abc_72207_new_n226_));
AND2X2 AND2X2_188 ( .A(spec_req_cs_4_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1330_));
AND2X2 AND2X2_1880 ( .A(u0_u0__abc_72207_new_n229_), .B(u0_u0__abc_72207_new_n228_), .Y(u0_u0__abc_72207_new_n230_));
AND2X2 AND2X2_1881 ( .A(u0_u0__abc_72207_new_n233_), .B(u0_u0__abc_72207_new_n232_), .Y(u0_u0__abc_72207_new_n234_));
AND2X2 AND2X2_1882 ( .A(u0_u0__abc_72207_new_n237_), .B(u0_u0__abc_72207_new_n236_), .Y(u0_u0__abc_72207_new_n238_));
AND2X2 AND2X2_1883 ( .A(u0_u0__abc_72207_new_n241_), .B(u0_u0__abc_72207_new_n240_), .Y(u0_u0__abc_72207_new_n242_));
AND2X2 AND2X2_1884 ( .A(u0_u0__abc_72207_new_n245_), .B(u0_u0__abc_72207_new_n244_), .Y(u0_u0__abc_72207_new_n246_));
AND2X2 AND2X2_1885 ( .A(u0_u0__abc_72207_new_n249_), .B(u0_u0__abc_72207_new_n248_), .Y(u0_u0__abc_72207_new_n250_));
AND2X2 AND2X2_1886 ( .A(u0_u0__abc_72207_new_n253_), .B(u0_u0__abc_72207_new_n252_), .Y(u0_u0__abc_72207_new_n254_));
AND2X2 AND2X2_1887 ( .A(u0_u0__abc_72207_new_n257_), .B(u0_u0__abc_72207_new_n256_), .Y(u0_u0__abc_72207_new_n258_));
AND2X2 AND2X2_1888 ( .A(u0_u0__abc_72207_new_n261_), .B(u0_u0__abc_72207_new_n260_), .Y(u0_u0__abc_72207_new_n262_));
AND2X2 AND2X2_1889 ( .A(u0_u0__abc_72207_new_n265_), .B(u0_u0__abc_72207_new_n264_), .Y(u0_u0__abc_72207_new_n266_));
AND2X2 AND2X2_189 ( .A(u0__abc_76628_new_n1331_), .B(u0__abc_76628_new_n1174__bF_buf5), .Y(u0__abc_76628_new_n1332_));
AND2X2 AND2X2_1890 ( .A(u0_u0__abc_72207_new_n269_), .B(u0_u0__abc_72207_new_n268_), .Y(u0_u0__abc_72207_new_n270_));
AND2X2 AND2X2_1891 ( .A(u0_u0__abc_72207_new_n273_), .B(u0_u0__abc_72207_new_n272_), .Y(u0_u0__abc_72207_new_n274_));
AND2X2 AND2X2_1892 ( .A(u0_u0__abc_72207_new_n277_), .B(u0_u0__abc_72207_new_n276_), .Y(u0_u0__abc_72207_new_n278_));
AND2X2 AND2X2_1893 ( .A(u0_u0__abc_72207_new_n281_), .B(u0_u0__abc_72207_new_n280_), .Y(u0_u0__abc_72207_new_n282_));
AND2X2 AND2X2_1894 ( .A(u0_u0__abc_72207_new_n285_), .B(u0_u0__abc_72207_new_n284_), .Y(u0_u0__abc_72207_new_n286_));
AND2X2 AND2X2_1895 ( .A(u0_u0__abc_72207_new_n289_), .B(u0_u0__abc_72207_new_n288_), .Y(u0_u0__abc_72207_new_n290_));
AND2X2 AND2X2_1896 ( .A(u0_u0__abc_72207_new_n293_), .B(u0_u0__abc_72207_new_n292_), .Y(u0_u0__abc_72207_new_n294_));
AND2X2 AND2X2_1897 ( .A(u0_u0__abc_72207_new_n297_), .B(u0_u0__abc_72207_new_n296_), .Y(u0_u0__abc_72207_new_n298_));
AND2X2 AND2X2_1898 ( .A(u0_u0__abc_72207_new_n301_), .B(u0_u0__abc_72207_new_n300_), .Y(u0_u0__abc_72207_new_n302_));
AND2X2 AND2X2_1899 ( .A(u0_u0__abc_72207_new_n305_), .B(u0_u0__abc_72207_new_n304_), .Y(u0_u0__abc_72207_new_n306_));
AND2X2 AND2X2_19 ( .A(_abc_85006_new_n293_), .B(_abc_85006_new_n294_), .Y(tms_s_1_));
AND2X2 AND2X2_190 ( .A(spec_req_cs_3_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1333_));
AND2X2 AND2X2_1900 ( .A(u0_u0__abc_72207_new_n309_), .B(u0_u0__abc_72207_new_n308_), .Y(u0_u0__abc_72207_new_n310_));
AND2X2 AND2X2_1901 ( .A(u0_u0__abc_72207_new_n313_), .B(u0_u0__abc_72207_new_n312_), .Y(u0_u0__abc_72207_new_n314_));
AND2X2 AND2X2_1902 ( .A(u0_u0__abc_72207_new_n317_), .B(u0_u0__abc_72207_new_n316_), .Y(u0_u0__abc_72207_new_n318_));
AND2X2 AND2X2_1903 ( .A(u0_u0__abc_72207_new_n321_), .B(u0_u0__abc_72207_new_n320_), .Y(u0_u0__abc_72207_new_n322_));
AND2X2 AND2X2_1904 ( .A(u0_u0__abc_72207_new_n325_), .B(u0_u0__abc_72207_new_n324_), .Y(u0_u0__abc_72207_new_n326_));
AND2X2 AND2X2_1905 ( .A(u0_u0__abc_72207_new_n329_), .B(u0_u0__abc_72207_new_n328_), .Y(u0_u0__abc_72207_new_n330_));
AND2X2 AND2X2_1906 ( .A(u0_u0__abc_72207_new_n333_), .B(u0_u0__abc_72207_new_n332_), .Y(u0_u0__abc_72207_new_n334_));
AND2X2 AND2X2_1907 ( .A(u0_u0__abc_72207_new_n337_), .B(u0_u0__abc_72207_new_n336_), .Y(u0_u0__abc_72207_new_n338_));
AND2X2 AND2X2_1908 ( .A(u0_u0__abc_72207_new_n341_), .B(u0_u0__abc_72207_new_n340_), .Y(u0_u0__abc_72207_new_n342_));
AND2X2 AND2X2_1909 ( .A(u0_u0__abc_72207_new_n345_), .B(u0_u0__abc_72207_new_n344_), .Y(u0_u0__abc_72207_new_n346_));
AND2X2 AND2X2_191 ( .A(u0__abc_76628_new_n1334_), .B(u0__abc_76628_new_n1173__bF_buf5), .Y(u0__abc_76628_new_n1335_));
AND2X2 AND2X2_1910 ( .A(u0_u0__abc_72207_new_n349_), .B(u0_u0__abc_72207_new_n348_), .Y(u0_u0__abc_72207_new_n350_));
AND2X2 AND2X2_1911 ( .A(u0_u0__abc_72207_new_n221_), .B(u0_u0__abc_72207_new_n352_), .Y(u0_u0__0init_req_we_0_0_));
AND2X2 AND2X2_1912 ( .A(u0_u0__abc_72207_new_n362_), .B(u0_u0__abc_72207_new_n355_), .Y(u0_u0__abc_72207_new_n363_));
AND2X2 AND2X2_1913 ( .A(u0_u0__abc_72207_new_n363_), .B(u0_u0__abc_72207_new_n354__bF_buf4), .Y(u0_u0__abc_72207_new_n364_));
AND2X2 AND2X2_1914 ( .A(u0_u0_rst_r2_bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_2_), .Y(u0_u0__abc_72207_new_n365_));
AND2X2 AND2X2_1915 ( .A(u0_u0_rst_r2_bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_3_), .Y(u0_u0__abc_72207_new_n366_));
AND2X2 AND2X2_1916 ( .A(u0_u0__abc_72207_new_n370_), .B(u0_u0__abc_72207_new_n354__bF_buf3), .Y(u0_u0__abc_72207_new_n371_));
AND2X2 AND2X2_1917 ( .A(u0_u0__abc_72207_new_n371_), .B(u0_u0__abc_72207_new_n369_), .Y(u0_u0__abc_72207_new_n372_));
AND2X2 AND2X2_1918 ( .A(u0_u0__abc_72207_new_n375_), .B(u0_u0__abc_72207_new_n354__bF_buf2), .Y(u0_u0__abc_72207_new_n376_));
AND2X2 AND2X2_1919 ( .A(u0_u0__abc_72207_new_n376_), .B(u0_u0__abc_72207_new_n374_), .Y(u0_u0__abc_72207_new_n377_));
AND2X2 AND2X2_192 ( .A(spec_req_cs_2_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1336_));
AND2X2 AND2X2_1920 ( .A(u0_u0__abc_72207_new_n380_), .B(u0_u0__abc_72207_new_n354__bF_buf1), .Y(u0_u0__abc_72207_new_n381_));
AND2X2 AND2X2_1921 ( .A(u0_u0__abc_72207_new_n381_), .B(u0_u0__abc_72207_new_n379_), .Y(u0_u0__0csc_31_0__3_));
AND2X2 AND2X2_1922 ( .A(u0_u0__abc_72207_new_n384_), .B(u0_u0__abc_72207_new_n383_), .Y(u0_u0__abc_72207_new_n385_));
AND2X2 AND2X2_1923 ( .A(u0_u0__abc_72207_new_n386_), .B(u0_u0__abc_72207_new_n387_), .Y(u0_u0__0csc_31_0__4_));
AND2X2 AND2X2_1924 ( .A(u0_u0__abc_72207_new_n390_), .B(u0_u0__abc_72207_new_n389_), .Y(u0_u0__abc_72207_new_n391_));
AND2X2 AND2X2_1925 ( .A(u0_u0__abc_72207_new_n392_), .B(u0_u0__abc_72207_new_n393_), .Y(u0_u0__0csc_31_0__5_));
AND2X2 AND2X2_1926 ( .A(u0_u0__abc_72207_new_n396_), .B(u0_u0__abc_72207_new_n354__bF_buf3), .Y(u0_u0__abc_72207_new_n397_));
AND2X2 AND2X2_1927 ( .A(u0_u0__abc_72207_new_n397_), .B(u0_u0__abc_72207_new_n395_), .Y(u0_u0__0csc_31_0__6_));
AND2X2 AND2X2_1928 ( .A(u0_u0__abc_72207_new_n400_), .B(u0_u0__abc_72207_new_n354__bF_buf2), .Y(u0_u0__abc_72207_new_n401_));
AND2X2 AND2X2_1929 ( .A(u0_u0__abc_72207_new_n401_), .B(u0_u0__abc_72207_new_n399_), .Y(u0_u0__0csc_31_0__7_));
AND2X2 AND2X2_193 ( .A(u0__abc_76628_new_n1337_), .B(u0__abc_76628_new_n1172__bF_buf5), .Y(u0__abc_76628_new_n1338_));
AND2X2 AND2X2_1930 ( .A(u0_u0__abc_72207_new_n404_), .B(u0_u0__abc_72207_new_n354__bF_buf1), .Y(u0_u0__abc_72207_new_n405_));
AND2X2 AND2X2_1931 ( .A(u0_u0__abc_72207_new_n405_), .B(u0_u0__abc_72207_new_n403_), .Y(u0_u0__0csc_31_0__8_));
AND2X2 AND2X2_1932 ( .A(u0_u0__abc_72207_new_n408_), .B(u0_u0__abc_72207_new_n354__bF_buf0), .Y(u0_u0__abc_72207_new_n409_));
AND2X2 AND2X2_1933 ( .A(u0_u0__abc_72207_new_n409_), .B(u0_u0__abc_72207_new_n407_), .Y(u0_u0__0csc_31_0__9_));
AND2X2 AND2X2_1934 ( .A(u0_u0__abc_72207_new_n412_), .B(u0_u0__abc_72207_new_n354__bF_buf4), .Y(u0_u0__abc_72207_new_n413_));
AND2X2 AND2X2_1935 ( .A(u0_u0__abc_72207_new_n413_), .B(u0_u0__abc_72207_new_n411_), .Y(u0_u0__0csc_31_0__10_));
AND2X2 AND2X2_1936 ( .A(u0_u0__abc_72207_new_n416_), .B(u0_u0__abc_72207_new_n354__bF_buf3), .Y(u0_u0__abc_72207_new_n417_));
AND2X2 AND2X2_1937 ( .A(u0_u0__abc_72207_new_n417_), .B(u0_u0__abc_72207_new_n415_), .Y(u0_u0__0csc_31_0__11_));
AND2X2 AND2X2_1938 ( .A(u0_u0__abc_72207_new_n420_), .B(u0_u0__abc_72207_new_n354__bF_buf2), .Y(u0_u0__abc_72207_new_n421_));
AND2X2 AND2X2_1939 ( .A(u0_u0__abc_72207_new_n421_), .B(u0_u0__abc_72207_new_n419_), .Y(u0_u0__0csc_31_0__12_));
AND2X2 AND2X2_194 ( .A(spec_req_cs_1_bF_buf2_), .B(u0_tms1_6_), .Y(u0__abc_76628_new_n1339_));
AND2X2 AND2X2_1940 ( .A(u0_u0__abc_72207_new_n424_), .B(u0_u0__abc_72207_new_n354__bF_buf1), .Y(u0_u0__abc_72207_new_n425_));
AND2X2 AND2X2_1941 ( .A(u0_u0__abc_72207_new_n425_), .B(u0_u0__abc_72207_new_n423_), .Y(u0_u0__0csc_31_0__13_));
AND2X2 AND2X2_1942 ( .A(u0_u0__abc_72207_new_n428_), .B(u0_u0__abc_72207_new_n354__bF_buf0), .Y(u0_u0__abc_72207_new_n429_));
AND2X2 AND2X2_1943 ( .A(u0_u0__abc_72207_new_n429_), .B(u0_u0__abc_72207_new_n427_), .Y(u0_u0__0csc_31_0__14_));
AND2X2 AND2X2_1944 ( .A(u0_u0__abc_72207_new_n432_), .B(u0_u0__abc_72207_new_n354__bF_buf4), .Y(u0_u0__abc_72207_new_n433_));
AND2X2 AND2X2_1945 ( .A(u0_u0__abc_72207_new_n433_), .B(u0_u0__abc_72207_new_n431_), .Y(u0_u0__0csc_31_0__15_));
AND2X2 AND2X2_1946 ( .A(u0_u0__abc_72207_new_n436_), .B(u0_u0__abc_72207_new_n354__bF_buf3), .Y(u0_u0__abc_72207_new_n437_));
AND2X2 AND2X2_1947 ( .A(u0_u0__abc_72207_new_n437_), .B(u0_u0__abc_72207_new_n435_), .Y(u0_u0__0csc_31_0__16_));
AND2X2 AND2X2_1948 ( .A(u0_u0__abc_72207_new_n440_), .B(u0_u0__abc_72207_new_n354__bF_buf2), .Y(u0_u0__abc_72207_new_n441_));
AND2X2 AND2X2_1949 ( .A(u0_u0__abc_72207_new_n441_), .B(u0_u0__abc_72207_new_n439_), .Y(u0_u0__0csc_31_0__17_));
AND2X2 AND2X2_195 ( .A(u0__abc_76628_new_n1169__bF_buf6), .B(u0__abc_76628_new_n1342_), .Y(u0__abc_76628_new_n1343_));
AND2X2 AND2X2_1950 ( .A(u0_u0__abc_72207_new_n444_), .B(u0_u0__abc_72207_new_n354__bF_buf1), .Y(u0_u0__abc_72207_new_n445_));
AND2X2 AND2X2_1951 ( .A(u0_u0__abc_72207_new_n445_), .B(u0_u0__abc_72207_new_n443_), .Y(u0_u0__0csc_31_0__18_));
AND2X2 AND2X2_1952 ( .A(u0_u0__abc_72207_new_n448_), .B(u0_u0__abc_72207_new_n354__bF_buf0), .Y(u0_u0__abc_72207_new_n449_));
AND2X2 AND2X2_1953 ( .A(u0_u0__abc_72207_new_n449_), .B(u0_u0__abc_72207_new_n447_), .Y(u0_u0__0csc_31_0__19_));
AND2X2 AND2X2_1954 ( .A(u0_u0__abc_72207_new_n452_), .B(u0_u0__abc_72207_new_n354__bF_buf4), .Y(u0_u0__abc_72207_new_n453_));
AND2X2 AND2X2_1955 ( .A(u0_u0__abc_72207_new_n453_), .B(u0_u0__abc_72207_new_n451_), .Y(u0_u0__0csc_31_0__20_));
AND2X2 AND2X2_1956 ( .A(u0_u0__abc_72207_new_n456_), .B(u0_u0__abc_72207_new_n354__bF_buf3), .Y(u0_u0__abc_72207_new_n457_));
AND2X2 AND2X2_1957 ( .A(u0_u0__abc_72207_new_n457_), .B(u0_u0__abc_72207_new_n455_), .Y(u0_u0__0csc_31_0__21_));
AND2X2 AND2X2_1958 ( .A(u0_u0__abc_72207_new_n460_), .B(u0_u0__abc_72207_new_n354__bF_buf2), .Y(u0_u0__abc_72207_new_n461_));
AND2X2 AND2X2_1959 ( .A(u0_u0__abc_72207_new_n461_), .B(u0_u0__abc_72207_new_n459_), .Y(u0_u0__0csc_31_0__22_));
AND2X2 AND2X2_196 ( .A(u0__abc_76628_new_n1341_), .B(u0__abc_76628_new_n1343_), .Y(u0__abc_76628_new_n1344_));
AND2X2 AND2X2_1960 ( .A(u0_u0__abc_72207_new_n464_), .B(u0_u0__abc_72207_new_n354__bF_buf1), .Y(u0_u0__abc_72207_new_n465_));
AND2X2 AND2X2_1961 ( .A(u0_u0__abc_72207_new_n465_), .B(u0_u0__abc_72207_new_n463_), .Y(u0_u0__0csc_31_0__23_));
AND2X2 AND2X2_1962 ( .A(u0_u0__abc_72207_new_n468_), .B(u0_u0__abc_72207_new_n354__bF_buf0), .Y(u0_u0__abc_72207_new_n469_));
AND2X2 AND2X2_1963 ( .A(u0_u0__abc_72207_new_n469_), .B(u0_u0__abc_72207_new_n467_), .Y(u0_u0__0csc_31_0__24_));
AND2X2 AND2X2_1964 ( .A(u0_u0__abc_72207_new_n472_), .B(u0_u0__abc_72207_new_n354__bF_buf4), .Y(u0_u0__abc_72207_new_n473_));
AND2X2 AND2X2_1965 ( .A(u0_u0__abc_72207_new_n473_), .B(u0_u0__abc_72207_new_n471_), .Y(u0_u0__0csc_31_0__25_));
AND2X2 AND2X2_1966 ( .A(u0_u0__abc_72207_new_n476_), .B(u0_u0__abc_72207_new_n354__bF_buf3), .Y(u0_u0__abc_72207_new_n477_));
AND2X2 AND2X2_1967 ( .A(u0_u0__abc_72207_new_n477_), .B(u0_u0__abc_72207_new_n475_), .Y(u0_u0__0csc_31_0__26_));
AND2X2 AND2X2_1968 ( .A(u0_u0__abc_72207_new_n480_), .B(u0_u0__abc_72207_new_n354__bF_buf2), .Y(u0_u0__abc_72207_new_n481_));
AND2X2 AND2X2_1969 ( .A(u0_u0__abc_72207_new_n481_), .B(u0_u0__abc_72207_new_n479_), .Y(u0_u0__0csc_31_0__27_));
AND2X2 AND2X2_197 ( .A(u0__abc_76628_new_n1170__bF_buf6), .B(sp_tms_7_), .Y(u0__abc_76628_new_n1346_));
AND2X2 AND2X2_1970 ( .A(u0_u0__abc_72207_new_n484_), .B(u0_u0__abc_72207_new_n354__bF_buf1), .Y(u0_u0__abc_72207_new_n485_));
AND2X2 AND2X2_1971 ( .A(u0_u0__abc_72207_new_n485_), .B(u0_u0__abc_72207_new_n483_), .Y(u0_u0__0csc_31_0__28_));
AND2X2 AND2X2_1972 ( .A(u0_u0__abc_72207_new_n488_), .B(u0_u0__abc_72207_new_n354__bF_buf0), .Y(u0_u0__abc_72207_new_n489_));
AND2X2 AND2X2_1973 ( .A(u0_u0__abc_72207_new_n489_), .B(u0_u0__abc_72207_new_n487_), .Y(u0_u0__0csc_31_0__29_));
AND2X2 AND2X2_1974 ( .A(u0_u0__abc_72207_new_n492_), .B(u0_u0__abc_72207_new_n354__bF_buf4), .Y(u0_u0__abc_72207_new_n493_));
AND2X2 AND2X2_1975 ( .A(u0_u0__abc_72207_new_n493_), .B(u0_u0__abc_72207_new_n491_), .Y(u0_u0__0csc_31_0__30_));
AND2X2 AND2X2_1976 ( .A(u0_u0__abc_72207_new_n496_), .B(u0_u0__abc_72207_new_n354__bF_buf3), .Y(u0_u0__abc_72207_new_n497_));
AND2X2 AND2X2_1977 ( .A(u0_u0__abc_72207_new_n497_), .B(u0_u0__abc_72207_new_n495_), .Y(u0_u0__0csc_31_0__31_));
AND2X2 AND2X2_1978 ( .A(u0_csc0_8_), .B(wb_we_i), .Y(u0_u0__abc_72207_new_n499_));
AND2X2 AND2X2_1979 ( .A(u0_u0__abc_72207_new_n500_), .B(u0_u0__abc_72207_new_n501_), .Y(u0_u0__abc_72207_new_n502_));
AND2X2 AND2X2_198 ( .A(spec_req_cs_5_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1347_));
AND2X2 AND2X2_1980 ( .A(u0_csc0_23_), .B(\wb_addr_i[28] ), .Y(u0_u0__abc_72207_new_n504_));
AND2X2 AND2X2_1981 ( .A(u0_csc0_22_), .B(\wb_addr_i[27] ), .Y(u0_u0__abc_72207_new_n507_));
AND2X2 AND2X2_1982 ( .A(u0_u0__abc_72207_new_n509_), .B(u0_u0__abc_72207_new_n510_), .Y(u0_u0__abc_72207_new_n511_));
AND2X2 AND2X2_1983 ( .A(u0_u0__abc_72207_new_n513_), .B(u0_u0__abc_72207_new_n506_), .Y(u0_u0__abc_72207_new_n514_));
AND2X2 AND2X2_1984 ( .A(u0_csc0_21_), .B(\wb_addr_i[26] ), .Y(u0_u0__abc_72207_new_n515_));
AND2X2 AND2X2_1985 ( .A(u0_u0__abc_72207_new_n517_), .B(u0_u0__abc_72207_new_n518_), .Y(u0_u0__abc_72207_new_n519_));
AND2X2 AND2X2_1986 ( .A(u0_u0__abc_72207_new_n514_), .B(u0_u0__abc_72207_new_n521_), .Y(u0_u0__abc_72207_new_n522_));
AND2X2 AND2X2_1987 ( .A(u0_csc0_16_), .B(\wb_addr_i[21] ), .Y(u0_u0__abc_72207_new_n523_));
AND2X2 AND2X2_1988 ( .A(u0_u0__abc_72207_new_n525_), .B(u0_u0__abc_72207_new_n526_), .Y(u0_u0__abc_72207_new_n527_));
AND2X2 AND2X2_1989 ( .A(u0_u0__abc_72207_new_n529_), .B(u0_csc0_0_), .Y(u0_u0__abc_72207_new_n530_));
AND2X2 AND2X2_199 ( .A(u0__abc_76628_new_n1349_), .B(u0__abc_76628_new_n1179__bF_buf4), .Y(u0__abc_76628_new_n1350_));
AND2X2 AND2X2_1990 ( .A(u0_csc0_18_), .B(\wb_addr_i[23] ), .Y(u0_u0__abc_72207_new_n531_));
AND2X2 AND2X2_1991 ( .A(u0_u0__abc_72207_new_n533_), .B(u0_u0__abc_72207_new_n534_), .Y(u0_u0__abc_72207_new_n535_));
AND2X2 AND2X2_1992 ( .A(u0_csc_mask_1_), .B(\wb_addr_i[22] ), .Y(u0_u0__abc_72207_new_n538_));
AND2X2 AND2X2_1993 ( .A(u0_csc0_17_), .B(u0_csc_mask_1_), .Y(u0_u0__abc_72207_new_n540_));
AND2X2 AND2X2_1994 ( .A(u0_u0__abc_72207_new_n541_), .B(u0_u0__abc_72207_new_n543_), .Y(u0_u0__abc_72207_new_n544_));
AND2X2 AND2X2_1995 ( .A(u0_u0__abc_72207_new_n537_), .B(u0_u0__abc_72207_new_n544_), .Y(u0_u0__abc_72207_new_n545_));
AND2X2 AND2X2_1996 ( .A(u0_csc_mask_4_), .B(\wb_addr_i[25] ), .Y(u0_u0__abc_72207_new_n546_));
AND2X2 AND2X2_1997 ( .A(u0_csc0_20_), .B(u0_csc_mask_4_), .Y(u0_u0__abc_72207_new_n548_));
AND2X2 AND2X2_1998 ( .A(u0_u0__abc_72207_new_n549_), .B(u0_u0__abc_72207_new_n551_), .Y(u0_u0__abc_72207_new_n552_));
AND2X2 AND2X2_1999 ( .A(u0_csc_mask_3_), .B(\wb_addr_i[24] ), .Y(u0_u0__abc_72207_new_n553_));
AND2X2 AND2X2_2 ( .A(_abc_85006_new_n241_), .B(_abc_85006_new_n242_), .Y(_abc_85006_new_n243_));
AND2X2 AND2X2_20 ( .A(_abc_85006_new_n296_), .B(_abc_85006_new_n297_), .Y(tms_s_2_));
AND2X2 AND2X2_200 ( .A(u0__abc_76628_new_n1350_), .B(u0__abc_76628_new_n1348_), .Y(u0__abc_76628_new_n1351_));
AND2X2 AND2X2_2000 ( .A(u0_csc0_19_), .B(u0_csc_mask_3_), .Y(u0_u0__abc_72207_new_n555_));
AND2X2 AND2X2_2001 ( .A(u0_u0__abc_72207_new_n556_), .B(u0_u0__abc_72207_new_n558_), .Y(u0_u0__abc_72207_new_n559_));
AND2X2 AND2X2_2002 ( .A(u0_u0__abc_72207_new_n552_), .B(u0_u0__abc_72207_new_n559_), .Y(u0_u0__abc_72207_new_n560_));
AND2X2 AND2X2_2003 ( .A(u0_u0__abc_72207_new_n545_), .B(u0_u0__abc_72207_new_n560_), .Y(u0_u0__abc_72207_new_n561_));
AND2X2 AND2X2_2004 ( .A(u0_u0__abc_72207_new_n561_), .B(u0_u0__abc_72207_new_n530_), .Y(u0_u0__abc_72207_new_n562_));
AND2X2 AND2X2_2005 ( .A(u0_u0__abc_72207_new_n562_), .B(u0_u0__abc_72207_new_n522_), .Y(u0_u0__abc_72207_new_n563_));
AND2X2 AND2X2_2006 ( .A(u0_u0__abc_72207_new_n563_), .B(u0_u0__abc_72207_new_n499_), .Y(u0_u0_wp_err));
AND2X2 AND2X2_2007 ( .A(u0_u0__abc_72207_new_n563_), .B(u0_u0__abc_72207_new_n565_), .Y(u0_cs0));
AND2X2 AND2X2_2008 ( .A(u0_u0__abc_72207_new_n568_), .B(u0_init_req0), .Y(u0_u0__abc_72207_new_n569_));
AND2X2 AND2X2_2009 ( .A(u0_u0__abc_72207_new_n570_), .B(u0_csc0_0_), .Y(u0_u0__abc_72207_new_n571_));
AND2X2 AND2X2_201 ( .A(u0__abc_76628_new_n1352_), .B(u0__abc_76628_new_n1175__bF_buf4), .Y(u0__abc_76628_new_n1353_));
AND2X2 AND2X2_2010 ( .A(u0_u0__abc_72207_new_n571_), .B(u0_u0_init_req_we), .Y(u0_u0__abc_72207_new_n572_));
AND2X2 AND2X2_2011 ( .A(u0_u0__abc_72207_new_n207_), .B(u0_u0__abc_72207_new_n572_), .Y(u0_u0__abc_72207_new_n573_));
AND2X2 AND2X2_2012 ( .A(u0_u1__abc_72579_new_n203_), .B(u0_u1_lmr_req_we), .Y(u0_u1__abc_72579_new_n204_));
AND2X2 AND2X2_2013 ( .A(u0_u1__abc_72579_new_n204_), .B(u0_u1_inited), .Y(u0_u1__abc_72579_new_n205_));
AND2X2 AND2X2_2014 ( .A(u0_u1__abc_72579_new_n207_), .B(u0_lmr_req1), .Y(u0_u1__abc_72579_new_n208_));
AND2X2 AND2X2_2015 ( .A(u0_u1__abc_72579_new_n206_), .B(u0_u1__abc_72579_new_n208_), .Y(u0_u1__abc_72579_new_n209_));
AND2X2 AND2X2_2016 ( .A(u0_u1__abc_72579_new_n211_), .B(u0_rf_we), .Y(u0_u1__abc_72579_new_n212_));
AND2X2 AND2X2_2017 ( .A(u0_u1_addr_r_4_), .B(u0_u1_addr_r_3_), .Y(u0_u1__abc_72579_new_n214_));
AND2X2 AND2X2_2018 ( .A(u0_u1__abc_72579_new_n214_), .B(u0_u1__abc_72579_new_n213_), .Y(u0_u1__abc_72579_new_n215_));
AND2X2 AND2X2_2019 ( .A(u0_u1__abc_72579_new_n215_), .B(u0_u1__abc_72579_new_n212_), .Y(u0_u1__abc_72579_new_n216_));
AND2X2 AND2X2_202 ( .A(spec_req_cs_4_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1354_));
AND2X2 AND2X2_2020 ( .A(u0_u1__abc_72579_new_n216_), .B(u0_u1_addr_r_2_), .Y(u0_u1__0lmr_req_we_0_0_));
AND2X2 AND2X2_2021 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n220_), .Y(u0_u1__abc_72579_new_n221_));
AND2X2 AND2X2_2022 ( .A(u0_u1__abc_72579_new_n222_), .B(u0_u1__abc_72579_new_n219__bF_buf7), .Y(u0_u1__abc_72579_new_n223_));
AND2X2 AND2X2_2023 ( .A(u0_u1__abc_72579_new_n223_), .B(u0_u1__abc_72579_new_n218_), .Y(u0_u1__0tms_31_0__0_));
AND2X2 AND2X2_2024 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n226_), .Y(u0_u1__abc_72579_new_n227_));
AND2X2 AND2X2_2025 ( .A(u0_u1__abc_72579_new_n228_), .B(u0_u1__abc_72579_new_n219__bF_buf6), .Y(u0_u1__abc_72579_new_n229_));
AND2X2 AND2X2_2026 ( .A(u0_u1__abc_72579_new_n229_), .B(u0_u1__abc_72579_new_n225_), .Y(u0_u1__0tms_31_0__1_));
AND2X2 AND2X2_2027 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n232_), .Y(u0_u1__abc_72579_new_n233_));
AND2X2 AND2X2_2028 ( .A(u0_u1__abc_72579_new_n234_), .B(u0_u1__abc_72579_new_n219__bF_buf5), .Y(u0_u1__abc_72579_new_n235_));
AND2X2 AND2X2_2029 ( .A(u0_u1__abc_72579_new_n235_), .B(u0_u1__abc_72579_new_n231_), .Y(u0_u1__0tms_31_0__2_));
AND2X2 AND2X2_203 ( .A(u0__abc_76628_new_n1355_), .B(u0__abc_76628_new_n1174__bF_buf4), .Y(u0__abc_76628_new_n1356_));
AND2X2 AND2X2_2030 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n238_), .Y(u0_u1__abc_72579_new_n239_));
AND2X2 AND2X2_2031 ( .A(u0_u1__abc_72579_new_n240_), .B(u0_u1__abc_72579_new_n219__bF_buf4), .Y(u0_u1__abc_72579_new_n241_));
AND2X2 AND2X2_2032 ( .A(u0_u1__abc_72579_new_n241_), .B(u0_u1__abc_72579_new_n237_), .Y(u0_u1__0tms_31_0__3_));
AND2X2 AND2X2_2033 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n244_), .Y(u0_u1__abc_72579_new_n245_));
AND2X2 AND2X2_2034 ( .A(u0_u1__abc_72579_new_n246_), .B(u0_u1__abc_72579_new_n219__bF_buf3), .Y(u0_u1__abc_72579_new_n247_));
AND2X2 AND2X2_2035 ( .A(u0_u1__abc_72579_new_n247_), .B(u0_u1__abc_72579_new_n243_), .Y(u0_u1__0tms_31_0__4_));
AND2X2 AND2X2_2036 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n250_), .Y(u0_u1__abc_72579_new_n251_));
AND2X2 AND2X2_2037 ( .A(u0_u1__abc_72579_new_n252_), .B(u0_u1__abc_72579_new_n219__bF_buf2), .Y(u0_u1__abc_72579_new_n253_));
AND2X2 AND2X2_2038 ( .A(u0_u1__abc_72579_new_n253_), .B(u0_u1__abc_72579_new_n249_), .Y(u0_u1__0tms_31_0__5_));
AND2X2 AND2X2_2039 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n256_), .Y(u0_u1__abc_72579_new_n257_));
AND2X2 AND2X2_204 ( .A(spec_req_cs_3_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1357_));
AND2X2 AND2X2_2040 ( .A(u0_u1__abc_72579_new_n258_), .B(u0_u1__abc_72579_new_n219__bF_buf1), .Y(u0_u1__abc_72579_new_n259_));
AND2X2 AND2X2_2041 ( .A(u0_u1__abc_72579_new_n259_), .B(u0_u1__abc_72579_new_n255_), .Y(u0_u1__0tms_31_0__6_));
AND2X2 AND2X2_2042 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n262_), .Y(u0_u1__abc_72579_new_n263_));
AND2X2 AND2X2_2043 ( .A(u0_u1__abc_72579_new_n264_), .B(u0_u1__abc_72579_new_n219__bF_buf0), .Y(u0_u1__abc_72579_new_n265_));
AND2X2 AND2X2_2044 ( .A(u0_u1__abc_72579_new_n265_), .B(u0_u1__abc_72579_new_n261_), .Y(u0_u1__0tms_31_0__7_));
AND2X2 AND2X2_2045 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n268_), .Y(u0_u1__abc_72579_new_n269_));
AND2X2 AND2X2_2046 ( .A(u0_u1__abc_72579_new_n270_), .B(u0_u1__abc_72579_new_n219__bF_buf7), .Y(u0_u1__abc_72579_new_n271_));
AND2X2 AND2X2_2047 ( .A(u0_u1__abc_72579_new_n271_), .B(u0_u1__abc_72579_new_n267_), .Y(u0_u1__0tms_31_0__8_));
AND2X2 AND2X2_2048 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n274_), .Y(u0_u1__abc_72579_new_n275_));
AND2X2 AND2X2_2049 ( .A(u0_u1__abc_72579_new_n276_), .B(u0_u1__abc_72579_new_n219__bF_buf6), .Y(u0_u1__abc_72579_new_n277_));
AND2X2 AND2X2_205 ( .A(u0__abc_76628_new_n1358_), .B(u0__abc_76628_new_n1173__bF_buf4), .Y(u0__abc_76628_new_n1359_));
AND2X2 AND2X2_2050 ( .A(u0_u1__abc_72579_new_n277_), .B(u0_u1__abc_72579_new_n273_), .Y(u0_u1__0tms_31_0__9_));
AND2X2 AND2X2_2051 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n280_), .Y(u0_u1__abc_72579_new_n281_));
AND2X2 AND2X2_2052 ( .A(u0_u1__abc_72579_new_n282_), .B(u0_u1__abc_72579_new_n219__bF_buf5), .Y(u0_u1__abc_72579_new_n283_));
AND2X2 AND2X2_2053 ( .A(u0_u1__abc_72579_new_n283_), .B(u0_u1__abc_72579_new_n279_), .Y(u0_u1__0tms_31_0__10_));
AND2X2 AND2X2_2054 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n286_), .Y(u0_u1__abc_72579_new_n287_));
AND2X2 AND2X2_2055 ( .A(u0_u1__abc_72579_new_n288_), .B(u0_u1__abc_72579_new_n219__bF_buf4), .Y(u0_u1__abc_72579_new_n289_));
AND2X2 AND2X2_2056 ( .A(u0_u1__abc_72579_new_n289_), .B(u0_u1__abc_72579_new_n285_), .Y(u0_u1__0tms_31_0__11_));
AND2X2 AND2X2_2057 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n292_), .Y(u0_u1__abc_72579_new_n293_));
AND2X2 AND2X2_2058 ( .A(u0_u1__abc_72579_new_n294_), .B(u0_u1__abc_72579_new_n219__bF_buf3), .Y(u0_u1__abc_72579_new_n295_));
AND2X2 AND2X2_2059 ( .A(u0_u1__abc_72579_new_n295_), .B(u0_u1__abc_72579_new_n291_), .Y(u0_u1__0tms_31_0__12_));
AND2X2 AND2X2_206 ( .A(spec_req_cs_2_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1360_));
AND2X2 AND2X2_2060 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n298_), .Y(u0_u1__abc_72579_new_n299_));
AND2X2 AND2X2_2061 ( .A(u0_u1__abc_72579_new_n300_), .B(u0_u1__abc_72579_new_n219__bF_buf2), .Y(u0_u1__abc_72579_new_n301_));
AND2X2 AND2X2_2062 ( .A(u0_u1__abc_72579_new_n301_), .B(u0_u1__abc_72579_new_n297_), .Y(u0_u1__0tms_31_0__13_));
AND2X2 AND2X2_2063 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n304_), .Y(u0_u1__abc_72579_new_n305_));
AND2X2 AND2X2_2064 ( .A(u0_u1__abc_72579_new_n306_), .B(u0_u1__abc_72579_new_n219__bF_buf1), .Y(u0_u1__abc_72579_new_n307_));
AND2X2 AND2X2_2065 ( .A(u0_u1__abc_72579_new_n307_), .B(u0_u1__abc_72579_new_n303_), .Y(u0_u1__0tms_31_0__14_));
AND2X2 AND2X2_2066 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n310_), .Y(u0_u1__abc_72579_new_n311_));
AND2X2 AND2X2_2067 ( .A(u0_u1__abc_72579_new_n312_), .B(u0_u1__abc_72579_new_n219__bF_buf0), .Y(u0_u1__abc_72579_new_n313_));
AND2X2 AND2X2_2068 ( .A(u0_u1__abc_72579_new_n313_), .B(u0_u1__abc_72579_new_n309_), .Y(u0_u1__0tms_31_0__15_));
AND2X2 AND2X2_2069 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n316_), .Y(u0_u1__abc_72579_new_n317_));
AND2X2 AND2X2_207 ( .A(u0__abc_76628_new_n1361_), .B(u0__abc_76628_new_n1172__bF_buf4), .Y(u0__abc_76628_new_n1362_));
AND2X2 AND2X2_2070 ( .A(u0_u1__abc_72579_new_n318_), .B(u0_u1__abc_72579_new_n219__bF_buf7), .Y(u0_u1__abc_72579_new_n319_));
AND2X2 AND2X2_2071 ( .A(u0_u1__abc_72579_new_n319_), .B(u0_u1__abc_72579_new_n315_), .Y(u0_u1__0tms_31_0__16_));
AND2X2 AND2X2_2072 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n322_), .Y(u0_u1__abc_72579_new_n323_));
AND2X2 AND2X2_2073 ( .A(u0_u1__abc_72579_new_n324_), .B(u0_u1__abc_72579_new_n219__bF_buf6), .Y(u0_u1__abc_72579_new_n325_));
AND2X2 AND2X2_2074 ( .A(u0_u1__abc_72579_new_n325_), .B(u0_u1__abc_72579_new_n321_), .Y(u0_u1__0tms_31_0__17_));
AND2X2 AND2X2_2075 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n328_), .Y(u0_u1__abc_72579_new_n329_));
AND2X2 AND2X2_2076 ( .A(u0_u1__abc_72579_new_n330_), .B(u0_u1__abc_72579_new_n219__bF_buf5), .Y(u0_u1__abc_72579_new_n331_));
AND2X2 AND2X2_2077 ( .A(u0_u1__abc_72579_new_n331_), .B(u0_u1__abc_72579_new_n327_), .Y(u0_u1__0tms_31_0__18_));
AND2X2 AND2X2_2078 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n334_), .Y(u0_u1__abc_72579_new_n335_));
AND2X2 AND2X2_2079 ( .A(u0_u1__abc_72579_new_n336_), .B(u0_u1__abc_72579_new_n219__bF_buf4), .Y(u0_u1__abc_72579_new_n337_));
AND2X2 AND2X2_208 ( .A(spec_req_cs_1_bF_buf1_), .B(u0_tms1_7_), .Y(u0__abc_76628_new_n1363_));
AND2X2 AND2X2_2080 ( .A(u0_u1__abc_72579_new_n337_), .B(u0_u1__abc_72579_new_n333_), .Y(u0_u1__0tms_31_0__19_));
AND2X2 AND2X2_2081 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n340_), .Y(u0_u1__abc_72579_new_n341_));
AND2X2 AND2X2_2082 ( .A(u0_u1__abc_72579_new_n342_), .B(u0_u1__abc_72579_new_n219__bF_buf3), .Y(u0_u1__abc_72579_new_n343_));
AND2X2 AND2X2_2083 ( .A(u0_u1__abc_72579_new_n343_), .B(u0_u1__abc_72579_new_n339_), .Y(u0_u1__0tms_31_0__20_));
AND2X2 AND2X2_2084 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n346_), .Y(u0_u1__abc_72579_new_n347_));
AND2X2 AND2X2_2085 ( .A(u0_u1__abc_72579_new_n348_), .B(u0_u1__abc_72579_new_n219__bF_buf2), .Y(u0_u1__abc_72579_new_n349_));
AND2X2 AND2X2_2086 ( .A(u0_u1__abc_72579_new_n349_), .B(u0_u1__abc_72579_new_n345_), .Y(u0_u1__0tms_31_0__21_));
AND2X2 AND2X2_2087 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n352_), .Y(u0_u1__abc_72579_new_n353_));
AND2X2 AND2X2_2088 ( .A(u0_u1__abc_72579_new_n354_), .B(u0_u1__abc_72579_new_n219__bF_buf1), .Y(u0_u1__abc_72579_new_n355_));
AND2X2 AND2X2_2089 ( .A(u0_u1__abc_72579_new_n355_), .B(u0_u1__abc_72579_new_n351_), .Y(u0_u1__0tms_31_0__22_));
AND2X2 AND2X2_209 ( .A(u0__abc_76628_new_n1169__bF_buf5), .B(u0__abc_76628_new_n1366_), .Y(u0__abc_76628_new_n1367_));
AND2X2 AND2X2_2090 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n358_), .Y(u0_u1__abc_72579_new_n359_));
AND2X2 AND2X2_2091 ( .A(u0_u1__abc_72579_new_n360_), .B(u0_u1__abc_72579_new_n219__bF_buf0), .Y(u0_u1__abc_72579_new_n361_));
AND2X2 AND2X2_2092 ( .A(u0_u1__abc_72579_new_n361_), .B(u0_u1__abc_72579_new_n357_), .Y(u0_u1__0tms_31_0__23_));
AND2X2 AND2X2_2093 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n364_), .Y(u0_u1__abc_72579_new_n365_));
AND2X2 AND2X2_2094 ( .A(u0_u1__abc_72579_new_n366_), .B(u0_u1__abc_72579_new_n219__bF_buf7), .Y(u0_u1__abc_72579_new_n367_));
AND2X2 AND2X2_2095 ( .A(u0_u1__abc_72579_new_n367_), .B(u0_u1__abc_72579_new_n363_), .Y(u0_u1__0tms_31_0__24_));
AND2X2 AND2X2_2096 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n370_), .Y(u0_u1__abc_72579_new_n371_));
AND2X2 AND2X2_2097 ( .A(u0_u1__abc_72579_new_n372_), .B(u0_u1__abc_72579_new_n219__bF_buf6), .Y(u0_u1__abc_72579_new_n373_));
AND2X2 AND2X2_2098 ( .A(u0_u1__abc_72579_new_n373_), .B(u0_u1__abc_72579_new_n369_), .Y(u0_u1__0tms_31_0__25_));
AND2X2 AND2X2_2099 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n376_), .Y(u0_u1__abc_72579_new_n377_));
AND2X2 AND2X2_21 ( .A(_abc_85006_new_n299_), .B(_abc_85006_new_n300_), .Y(tms_s_3_));
AND2X2 AND2X2_210 ( .A(u0__abc_76628_new_n1365_), .B(u0__abc_76628_new_n1367_), .Y(u0__abc_76628_new_n1368_));
AND2X2 AND2X2_2100 ( .A(u0_u1__abc_72579_new_n378_), .B(u0_u1__abc_72579_new_n219__bF_buf5), .Y(u0_u1__abc_72579_new_n379_));
AND2X2 AND2X2_2101 ( .A(u0_u1__abc_72579_new_n379_), .B(u0_u1__abc_72579_new_n375_), .Y(u0_u1__0tms_31_0__26_));
AND2X2 AND2X2_2102 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n382_), .Y(u0_u1__abc_72579_new_n383_));
AND2X2 AND2X2_2103 ( .A(u0_u1__abc_72579_new_n384_), .B(u0_u1__abc_72579_new_n219__bF_buf4), .Y(u0_u1__abc_72579_new_n385_));
AND2X2 AND2X2_2104 ( .A(u0_u1__abc_72579_new_n385_), .B(u0_u1__abc_72579_new_n381_), .Y(u0_u1__0tms_31_0__27_));
AND2X2 AND2X2_2105 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n388_), .Y(u0_u1__abc_72579_new_n389_));
AND2X2 AND2X2_2106 ( .A(u0_u1__abc_72579_new_n390_), .B(u0_u1__abc_72579_new_n219__bF_buf3), .Y(u0_u1__abc_72579_new_n391_));
AND2X2 AND2X2_2107 ( .A(u0_u1__abc_72579_new_n391_), .B(u0_u1__abc_72579_new_n387_), .Y(u0_u1__0tms_31_0__28_));
AND2X2 AND2X2_2108 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n394_), .Y(u0_u1__abc_72579_new_n395_));
AND2X2 AND2X2_2109 ( .A(u0_u1__abc_72579_new_n396_), .B(u0_u1__abc_72579_new_n219__bF_buf2), .Y(u0_u1__abc_72579_new_n397_));
AND2X2 AND2X2_211 ( .A(u0__abc_76628_new_n1170__bF_buf5), .B(sp_tms_8_), .Y(u0__abc_76628_new_n1370_));
AND2X2 AND2X2_2110 ( .A(u0_u1__abc_72579_new_n397_), .B(u0_u1__abc_72579_new_n393_), .Y(u0_u1__0tms_31_0__29_));
AND2X2 AND2X2_2111 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n400_), .Y(u0_u1__abc_72579_new_n401_));
AND2X2 AND2X2_2112 ( .A(u0_u1__abc_72579_new_n402_), .B(u0_u1__abc_72579_new_n219__bF_buf1), .Y(u0_u1__abc_72579_new_n403_));
AND2X2 AND2X2_2113 ( .A(u0_u1__abc_72579_new_n403_), .B(u0_u1__abc_72579_new_n399_), .Y(u0_u1__0tms_31_0__30_));
AND2X2 AND2X2_2114 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n406_), .Y(u0_u1__abc_72579_new_n407_));
AND2X2 AND2X2_2115 ( .A(u0_u1__abc_72579_new_n408_), .B(u0_u1__abc_72579_new_n219__bF_buf0), .Y(u0_u1__abc_72579_new_n409_));
AND2X2 AND2X2_2116 ( .A(u0_u1__abc_72579_new_n409_), .B(u0_u1__abc_72579_new_n405_), .Y(u0_u1__0tms_31_0__31_));
AND2X2 AND2X2_2117 ( .A(u0_u1__abc_72579_new_n216_), .B(u0_u1__abc_72579_new_n411_), .Y(u0_u1__0init_req_we_0_0_));
AND2X2 AND2X2_2118 ( .A(u0_u1__0init_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n220_), .Y(u0_u1__abc_72579_new_n414_));
AND2X2 AND2X2_2119 ( .A(u0_u1__abc_72579_new_n415_), .B(u0_u1__abc_72579_new_n219__bF_buf7), .Y(u0_u1__abc_72579_new_n416_));
AND2X2 AND2X2_212 ( .A(spec_req_cs_5_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1371_));
AND2X2 AND2X2_2120 ( .A(u0_u1__abc_72579_new_n416_), .B(u0_u1__abc_72579_new_n413_), .Y(u0_u1__0csc_31_0__0_));
AND2X2 AND2X2_2121 ( .A(u0_u1__0init_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n226_), .Y(u0_u1__abc_72579_new_n419_));
AND2X2 AND2X2_2122 ( .A(u0_u1__abc_72579_new_n420_), .B(u0_u1__abc_72579_new_n219__bF_buf6), .Y(u0_u1__abc_72579_new_n421_));
AND2X2 AND2X2_2123 ( .A(u0_u1__abc_72579_new_n421_), .B(u0_u1__abc_72579_new_n418_), .Y(u0_u1__0csc_31_0__1_));
AND2X2 AND2X2_2124 ( .A(u0_u1__0init_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n232_), .Y(u0_u1__abc_72579_new_n424_));
AND2X2 AND2X2_2125 ( .A(u0_u1__abc_72579_new_n425_), .B(u0_u1__abc_72579_new_n219__bF_buf5), .Y(u0_u1__abc_72579_new_n426_));
AND2X2 AND2X2_2126 ( .A(u0_u1__abc_72579_new_n426_), .B(u0_u1__abc_72579_new_n423_), .Y(u0_u1__0csc_31_0__2_));
AND2X2 AND2X2_2127 ( .A(u0_u1__0init_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n238_), .Y(u0_u1__abc_72579_new_n429_));
AND2X2 AND2X2_2128 ( .A(u0_u1__abc_72579_new_n430_), .B(u0_u1__abc_72579_new_n219__bF_buf4), .Y(u0_u1__abc_72579_new_n431_));
AND2X2 AND2X2_2129 ( .A(u0_u1__abc_72579_new_n431_), .B(u0_u1__abc_72579_new_n428_), .Y(u0_u1__0csc_31_0__3_));
AND2X2 AND2X2_213 ( .A(u0__abc_76628_new_n1373_), .B(u0__abc_76628_new_n1179__bF_buf3), .Y(u0__abc_76628_new_n1374_));
AND2X2 AND2X2_2130 ( .A(u0_u1__0init_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n244_), .Y(u0_u1__abc_72579_new_n434_));
AND2X2 AND2X2_2131 ( .A(u0_u1__abc_72579_new_n435_), .B(u0_u1__abc_72579_new_n219__bF_buf3), .Y(u0_u1__abc_72579_new_n436_));
AND2X2 AND2X2_2132 ( .A(u0_u1__abc_72579_new_n436_), .B(u0_u1__abc_72579_new_n433_), .Y(u0_u1__0csc_31_0__4_));
AND2X2 AND2X2_2133 ( .A(u0_u1__0init_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n250_), .Y(u0_u1__abc_72579_new_n439_));
AND2X2 AND2X2_2134 ( .A(u0_u1__abc_72579_new_n440_), .B(u0_u1__abc_72579_new_n219__bF_buf2), .Y(u0_u1__abc_72579_new_n441_));
AND2X2 AND2X2_2135 ( .A(u0_u1__abc_72579_new_n441_), .B(u0_u1__abc_72579_new_n438_), .Y(u0_u1__0csc_31_0__5_));
AND2X2 AND2X2_2136 ( .A(u0_u1__0init_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n256_), .Y(u0_u1__abc_72579_new_n444_));
AND2X2 AND2X2_2137 ( .A(u0_u1__abc_72579_new_n445_), .B(u0_u1__abc_72579_new_n219__bF_buf1), .Y(u0_u1__abc_72579_new_n446_));
AND2X2 AND2X2_2138 ( .A(u0_u1__abc_72579_new_n446_), .B(u0_u1__abc_72579_new_n443_), .Y(u0_u1__0csc_31_0__6_));
AND2X2 AND2X2_2139 ( .A(u0_u1__0init_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n262_), .Y(u0_u1__abc_72579_new_n449_));
AND2X2 AND2X2_214 ( .A(u0__abc_76628_new_n1374_), .B(u0__abc_76628_new_n1372_), .Y(u0__abc_76628_new_n1375_));
AND2X2 AND2X2_2140 ( .A(u0_u1__abc_72579_new_n450_), .B(u0_u1__abc_72579_new_n219__bF_buf0), .Y(u0_u1__abc_72579_new_n451_));
AND2X2 AND2X2_2141 ( .A(u0_u1__abc_72579_new_n451_), .B(u0_u1__abc_72579_new_n448_), .Y(u0_u1__0csc_31_0__7_));
AND2X2 AND2X2_2142 ( .A(u0_u1__0init_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n268_), .Y(u0_u1__abc_72579_new_n454_));
AND2X2 AND2X2_2143 ( .A(u0_u1__abc_72579_new_n455_), .B(u0_u1__abc_72579_new_n219__bF_buf7), .Y(u0_u1__abc_72579_new_n456_));
AND2X2 AND2X2_2144 ( .A(u0_u1__abc_72579_new_n456_), .B(u0_u1__abc_72579_new_n453_), .Y(u0_u1__0csc_31_0__8_));
AND2X2 AND2X2_2145 ( .A(u0_u1__0init_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n274_), .Y(u0_u1__abc_72579_new_n459_));
AND2X2 AND2X2_2146 ( .A(u0_u1__abc_72579_new_n460_), .B(u0_u1__abc_72579_new_n219__bF_buf6), .Y(u0_u1__abc_72579_new_n461_));
AND2X2 AND2X2_2147 ( .A(u0_u1__abc_72579_new_n461_), .B(u0_u1__abc_72579_new_n458_), .Y(u0_u1__0csc_31_0__9_));
AND2X2 AND2X2_2148 ( .A(u0_u1__0init_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n280_), .Y(u0_u1__abc_72579_new_n464_));
AND2X2 AND2X2_2149 ( .A(u0_u1__abc_72579_new_n465_), .B(u0_u1__abc_72579_new_n219__bF_buf5), .Y(u0_u1__abc_72579_new_n466_));
AND2X2 AND2X2_215 ( .A(u0__abc_76628_new_n1376_), .B(u0__abc_76628_new_n1175__bF_buf3), .Y(u0__abc_76628_new_n1377_));
AND2X2 AND2X2_2150 ( .A(u0_u1__abc_72579_new_n466_), .B(u0_u1__abc_72579_new_n463_), .Y(u0_u1__0csc_31_0__10_));
AND2X2 AND2X2_2151 ( .A(u0_u1__0init_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n286_), .Y(u0_u1__abc_72579_new_n469_));
AND2X2 AND2X2_2152 ( .A(u0_u1__abc_72579_new_n470_), .B(u0_u1__abc_72579_new_n219__bF_buf4), .Y(u0_u1__abc_72579_new_n471_));
AND2X2 AND2X2_2153 ( .A(u0_u1__abc_72579_new_n471_), .B(u0_u1__abc_72579_new_n468_), .Y(u0_u1__0csc_31_0__11_));
AND2X2 AND2X2_2154 ( .A(u0_u1__0init_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n292_), .Y(u0_u1__abc_72579_new_n474_));
AND2X2 AND2X2_2155 ( .A(u0_u1__abc_72579_new_n475_), .B(u0_u1__abc_72579_new_n219__bF_buf3), .Y(u0_u1__abc_72579_new_n476_));
AND2X2 AND2X2_2156 ( .A(u0_u1__abc_72579_new_n476_), .B(u0_u1__abc_72579_new_n473_), .Y(u0_u1__0csc_31_0__12_));
AND2X2 AND2X2_2157 ( .A(u0_u1__0init_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n298_), .Y(u0_u1__abc_72579_new_n479_));
AND2X2 AND2X2_2158 ( .A(u0_u1__abc_72579_new_n480_), .B(u0_u1__abc_72579_new_n219__bF_buf2), .Y(u0_u1__abc_72579_new_n481_));
AND2X2 AND2X2_2159 ( .A(u0_u1__abc_72579_new_n481_), .B(u0_u1__abc_72579_new_n478_), .Y(u0_u1__0csc_31_0__13_));
AND2X2 AND2X2_216 ( .A(spec_req_cs_4_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1378_));
AND2X2 AND2X2_2160 ( .A(u0_u1__0init_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n304_), .Y(u0_u1__abc_72579_new_n484_));
AND2X2 AND2X2_2161 ( .A(u0_u1__abc_72579_new_n485_), .B(u0_u1__abc_72579_new_n219__bF_buf1), .Y(u0_u1__abc_72579_new_n486_));
AND2X2 AND2X2_2162 ( .A(u0_u1__abc_72579_new_n486_), .B(u0_u1__abc_72579_new_n483_), .Y(u0_u1__0csc_31_0__14_));
AND2X2 AND2X2_2163 ( .A(u0_u1__0init_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n310_), .Y(u0_u1__abc_72579_new_n489_));
AND2X2 AND2X2_2164 ( .A(u0_u1__abc_72579_new_n490_), .B(u0_u1__abc_72579_new_n219__bF_buf0), .Y(u0_u1__abc_72579_new_n491_));
AND2X2 AND2X2_2165 ( .A(u0_u1__abc_72579_new_n491_), .B(u0_u1__abc_72579_new_n488_), .Y(u0_u1__0csc_31_0__15_));
AND2X2 AND2X2_2166 ( .A(u0_u1__0init_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n316_), .Y(u0_u1__abc_72579_new_n494_));
AND2X2 AND2X2_2167 ( .A(u0_u1__abc_72579_new_n495_), .B(u0_u1__abc_72579_new_n219__bF_buf7), .Y(u0_u1__abc_72579_new_n496_));
AND2X2 AND2X2_2168 ( .A(u0_u1__abc_72579_new_n496_), .B(u0_u1__abc_72579_new_n493_), .Y(u0_u1__0csc_31_0__16_));
AND2X2 AND2X2_2169 ( .A(u0_u1__0init_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n322_), .Y(u0_u1__abc_72579_new_n499_));
AND2X2 AND2X2_217 ( .A(u0__abc_76628_new_n1379_), .B(u0__abc_76628_new_n1174__bF_buf3), .Y(u0__abc_76628_new_n1380_));
AND2X2 AND2X2_2170 ( .A(u0_u1__abc_72579_new_n500_), .B(u0_u1__abc_72579_new_n219__bF_buf6), .Y(u0_u1__abc_72579_new_n501_));
AND2X2 AND2X2_2171 ( .A(u0_u1__abc_72579_new_n501_), .B(u0_u1__abc_72579_new_n498_), .Y(u0_u1__0csc_31_0__17_));
AND2X2 AND2X2_2172 ( .A(u0_u1__0init_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n328_), .Y(u0_u1__abc_72579_new_n504_));
AND2X2 AND2X2_2173 ( .A(u0_u1__abc_72579_new_n505_), .B(u0_u1__abc_72579_new_n219__bF_buf5), .Y(u0_u1__abc_72579_new_n506_));
AND2X2 AND2X2_2174 ( .A(u0_u1__abc_72579_new_n506_), .B(u0_u1__abc_72579_new_n503_), .Y(u0_u1__0csc_31_0__18_));
AND2X2 AND2X2_2175 ( .A(u0_u1__0init_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n334_), .Y(u0_u1__abc_72579_new_n509_));
AND2X2 AND2X2_2176 ( .A(u0_u1__abc_72579_new_n510_), .B(u0_u1__abc_72579_new_n219__bF_buf4), .Y(u0_u1__abc_72579_new_n511_));
AND2X2 AND2X2_2177 ( .A(u0_u1__abc_72579_new_n511_), .B(u0_u1__abc_72579_new_n508_), .Y(u0_u1__0csc_31_0__19_));
AND2X2 AND2X2_2178 ( .A(u0_u1__0init_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n340_), .Y(u0_u1__abc_72579_new_n514_));
AND2X2 AND2X2_2179 ( .A(u0_u1__abc_72579_new_n515_), .B(u0_u1__abc_72579_new_n219__bF_buf3), .Y(u0_u1__abc_72579_new_n516_));
AND2X2 AND2X2_218 ( .A(spec_req_cs_3_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1381_));
AND2X2 AND2X2_2180 ( .A(u0_u1__abc_72579_new_n516_), .B(u0_u1__abc_72579_new_n513_), .Y(u0_u1__0csc_31_0__20_));
AND2X2 AND2X2_2181 ( .A(u0_u1__0init_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n346_), .Y(u0_u1__abc_72579_new_n519_));
AND2X2 AND2X2_2182 ( .A(u0_u1__abc_72579_new_n520_), .B(u0_u1__abc_72579_new_n219__bF_buf2), .Y(u0_u1__abc_72579_new_n521_));
AND2X2 AND2X2_2183 ( .A(u0_u1__abc_72579_new_n521_), .B(u0_u1__abc_72579_new_n518_), .Y(u0_u1__0csc_31_0__21_));
AND2X2 AND2X2_2184 ( .A(u0_u1__0init_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n352_), .Y(u0_u1__abc_72579_new_n524_));
AND2X2 AND2X2_2185 ( .A(u0_u1__abc_72579_new_n525_), .B(u0_u1__abc_72579_new_n219__bF_buf1), .Y(u0_u1__abc_72579_new_n526_));
AND2X2 AND2X2_2186 ( .A(u0_u1__abc_72579_new_n526_), .B(u0_u1__abc_72579_new_n523_), .Y(u0_u1__0csc_31_0__22_));
AND2X2 AND2X2_2187 ( .A(u0_u1__0init_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n358_), .Y(u0_u1__abc_72579_new_n529_));
AND2X2 AND2X2_2188 ( .A(u0_u1__abc_72579_new_n530_), .B(u0_u1__abc_72579_new_n219__bF_buf0), .Y(u0_u1__abc_72579_new_n531_));
AND2X2 AND2X2_2189 ( .A(u0_u1__abc_72579_new_n531_), .B(u0_u1__abc_72579_new_n528_), .Y(u0_u1__0csc_31_0__23_));
AND2X2 AND2X2_219 ( .A(u0__abc_76628_new_n1382_), .B(u0__abc_76628_new_n1173__bF_buf3), .Y(u0__abc_76628_new_n1383_));
AND2X2 AND2X2_2190 ( .A(u0_u1__0init_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n364_), .Y(u0_u1__abc_72579_new_n534_));
AND2X2 AND2X2_2191 ( .A(u0_u1__abc_72579_new_n535_), .B(u0_u1__abc_72579_new_n219__bF_buf7), .Y(u0_u1__abc_72579_new_n536_));
AND2X2 AND2X2_2192 ( .A(u0_u1__abc_72579_new_n536_), .B(u0_u1__abc_72579_new_n533_), .Y(u0_u1__0csc_31_0__24_));
AND2X2 AND2X2_2193 ( .A(u0_u1__0init_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n370_), .Y(u0_u1__abc_72579_new_n539_));
AND2X2 AND2X2_2194 ( .A(u0_u1__abc_72579_new_n540_), .B(u0_u1__abc_72579_new_n219__bF_buf6), .Y(u0_u1__abc_72579_new_n541_));
AND2X2 AND2X2_2195 ( .A(u0_u1__abc_72579_new_n541_), .B(u0_u1__abc_72579_new_n538_), .Y(u0_u1__0csc_31_0__25_));
AND2X2 AND2X2_2196 ( .A(u0_u1__0init_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n376_), .Y(u0_u1__abc_72579_new_n544_));
AND2X2 AND2X2_2197 ( .A(u0_u1__abc_72579_new_n545_), .B(u0_u1__abc_72579_new_n219__bF_buf5), .Y(u0_u1__abc_72579_new_n546_));
AND2X2 AND2X2_2198 ( .A(u0_u1__abc_72579_new_n546_), .B(u0_u1__abc_72579_new_n543_), .Y(u0_u1__0csc_31_0__26_));
AND2X2 AND2X2_2199 ( .A(u0_u1__0init_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n382_), .Y(u0_u1__abc_72579_new_n549_));
AND2X2 AND2X2_22 ( .A(_abc_85006_new_n302_), .B(_abc_85006_new_n303_), .Y(tms_s_4_));
AND2X2 AND2X2_220 ( .A(spec_req_cs_2_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1384_));
AND2X2 AND2X2_2200 ( .A(u0_u1__abc_72579_new_n550_), .B(u0_u1__abc_72579_new_n219__bF_buf4), .Y(u0_u1__abc_72579_new_n551_));
AND2X2 AND2X2_2201 ( .A(u0_u1__abc_72579_new_n551_), .B(u0_u1__abc_72579_new_n548_), .Y(u0_u1__0csc_31_0__27_));
AND2X2 AND2X2_2202 ( .A(u0_u1__0init_req_we_0_0_bF_buf6_), .B(u0_u1__abc_72579_new_n388_), .Y(u0_u1__abc_72579_new_n554_));
AND2X2 AND2X2_2203 ( .A(u0_u1__abc_72579_new_n555_), .B(u0_u1__abc_72579_new_n219__bF_buf3), .Y(u0_u1__abc_72579_new_n556_));
AND2X2 AND2X2_2204 ( .A(u0_u1__abc_72579_new_n556_), .B(u0_u1__abc_72579_new_n553_), .Y(u0_u1__0csc_31_0__28_));
AND2X2 AND2X2_2205 ( .A(u0_u1__0init_req_we_0_0_bF_buf4_), .B(u0_u1__abc_72579_new_n394_), .Y(u0_u1__abc_72579_new_n559_));
AND2X2 AND2X2_2206 ( .A(u0_u1__abc_72579_new_n560_), .B(u0_u1__abc_72579_new_n219__bF_buf2), .Y(u0_u1__abc_72579_new_n561_));
AND2X2 AND2X2_2207 ( .A(u0_u1__abc_72579_new_n561_), .B(u0_u1__abc_72579_new_n558_), .Y(u0_u1__0csc_31_0__29_));
AND2X2 AND2X2_2208 ( .A(u0_u1__0init_req_we_0_0_bF_buf2_), .B(u0_u1__abc_72579_new_n400_), .Y(u0_u1__abc_72579_new_n564_));
AND2X2 AND2X2_2209 ( .A(u0_u1__abc_72579_new_n565_), .B(u0_u1__abc_72579_new_n219__bF_buf1), .Y(u0_u1__abc_72579_new_n566_));
AND2X2 AND2X2_221 ( .A(u0__abc_76628_new_n1385_), .B(u0__abc_76628_new_n1172__bF_buf3), .Y(u0__abc_76628_new_n1386_));
AND2X2 AND2X2_2210 ( .A(u0_u1__abc_72579_new_n566_), .B(u0_u1__abc_72579_new_n563_), .Y(u0_u1__0csc_31_0__30_));
AND2X2 AND2X2_2211 ( .A(u0_u1__0init_req_we_0_0_bF_buf0_), .B(u0_u1__abc_72579_new_n406_), .Y(u0_u1__abc_72579_new_n569_));
AND2X2 AND2X2_2212 ( .A(u0_u1__abc_72579_new_n570_), .B(u0_u1__abc_72579_new_n219__bF_buf0), .Y(u0_u1__abc_72579_new_n571_));
AND2X2 AND2X2_2213 ( .A(u0_u1__abc_72579_new_n571_), .B(u0_u1__abc_72579_new_n568_), .Y(u0_u1__0csc_31_0__31_));
AND2X2 AND2X2_2214 ( .A(u0_csc1_8_), .B(wb_we_i), .Y(u0_u1__abc_72579_new_n573_));
AND2X2 AND2X2_2215 ( .A(u0_u1__abc_72579_new_n574_), .B(u0_u1__abc_72579_new_n575_), .Y(u0_u1__abc_72579_new_n576_));
AND2X2 AND2X2_2216 ( .A(u0_csc1_23_), .B(\wb_addr_i[28] ), .Y(u0_u1__abc_72579_new_n578_));
AND2X2 AND2X2_2217 ( .A(u0_csc1_22_), .B(\wb_addr_i[27] ), .Y(u0_u1__abc_72579_new_n581_));
AND2X2 AND2X2_2218 ( .A(u0_u1__abc_72579_new_n583_), .B(u0_u1__abc_72579_new_n584_), .Y(u0_u1__abc_72579_new_n585_));
AND2X2 AND2X2_2219 ( .A(u0_u1__abc_72579_new_n587_), .B(u0_u1__abc_72579_new_n580_), .Y(u0_u1__abc_72579_new_n588_));
AND2X2 AND2X2_222 ( .A(spec_req_cs_1_bF_buf0_), .B(u0_tms1_8_), .Y(u0__abc_76628_new_n1387_));
AND2X2 AND2X2_2220 ( .A(u0_csc1_21_), .B(\wb_addr_i[26] ), .Y(u0_u1__abc_72579_new_n589_));
AND2X2 AND2X2_2221 ( .A(u0_u1__abc_72579_new_n591_), .B(u0_u1__abc_72579_new_n592_), .Y(u0_u1__abc_72579_new_n593_));
AND2X2 AND2X2_2222 ( .A(u0_u1__abc_72579_new_n588_), .B(u0_u1__abc_72579_new_n595_), .Y(u0_u1__abc_72579_new_n596_));
AND2X2 AND2X2_2223 ( .A(u0_csc1_16_), .B(\wb_addr_i[21] ), .Y(u0_u1__abc_72579_new_n597_));
AND2X2 AND2X2_2224 ( .A(u0_u1__abc_72579_new_n599_), .B(u0_u1__abc_72579_new_n600_), .Y(u0_u1__abc_72579_new_n601_));
AND2X2 AND2X2_2225 ( .A(u0_u1__abc_72579_new_n603_), .B(u0_csc1_0_), .Y(u0_u1__abc_72579_new_n604_));
AND2X2 AND2X2_2226 ( .A(u0_csc_mask_2_), .B(\wb_addr_i[23] ), .Y(u0_u1__abc_72579_new_n605_));
AND2X2 AND2X2_2227 ( .A(u0_csc1_18_), .B(u0_csc_mask_2_), .Y(u0_u1__abc_72579_new_n607_));
AND2X2 AND2X2_2228 ( .A(u0_u1__abc_72579_new_n608_), .B(u0_u1__abc_72579_new_n610_), .Y(u0_u1__abc_72579_new_n611_));
AND2X2 AND2X2_2229 ( .A(u0_csc_mask_1_), .B(\wb_addr_i[22] ), .Y(u0_u1__abc_72579_new_n612_));
AND2X2 AND2X2_223 ( .A(u0__abc_76628_new_n1169__bF_buf4), .B(u0__abc_76628_new_n1390_), .Y(u0__abc_76628_new_n1391_));
AND2X2 AND2X2_2230 ( .A(u0_csc1_17_), .B(u0_csc_mask_1_), .Y(u0_u1__abc_72579_new_n614_));
AND2X2 AND2X2_2231 ( .A(u0_u1__abc_72579_new_n615_), .B(u0_u1__abc_72579_new_n617_), .Y(u0_u1__abc_72579_new_n618_));
AND2X2 AND2X2_2232 ( .A(u0_u1__abc_72579_new_n611_), .B(u0_u1__abc_72579_new_n618_), .Y(u0_u1__abc_72579_new_n619_));
AND2X2 AND2X2_2233 ( .A(u0_csc_mask_4_), .B(\wb_addr_i[25] ), .Y(u0_u1__abc_72579_new_n620_));
AND2X2 AND2X2_2234 ( .A(u0_csc1_20_), .B(u0_csc_mask_4_), .Y(u0_u1__abc_72579_new_n622_));
AND2X2 AND2X2_2235 ( .A(u0_u1__abc_72579_new_n623_), .B(u0_u1__abc_72579_new_n625_), .Y(u0_u1__abc_72579_new_n626_));
AND2X2 AND2X2_2236 ( .A(u0_csc_mask_3_), .B(\wb_addr_i[24] ), .Y(u0_u1__abc_72579_new_n627_));
AND2X2 AND2X2_2237 ( .A(u0_csc1_19_), .B(u0_csc_mask_3_), .Y(u0_u1__abc_72579_new_n629_));
AND2X2 AND2X2_2238 ( .A(u0_u1__abc_72579_new_n630_), .B(u0_u1__abc_72579_new_n632_), .Y(u0_u1__abc_72579_new_n633_));
AND2X2 AND2X2_2239 ( .A(u0_u1__abc_72579_new_n626_), .B(u0_u1__abc_72579_new_n633_), .Y(u0_u1__abc_72579_new_n634_));
AND2X2 AND2X2_224 ( .A(u0__abc_76628_new_n1389_), .B(u0__abc_76628_new_n1391_), .Y(u0__abc_76628_new_n1392_));
AND2X2 AND2X2_2240 ( .A(u0_u1__abc_72579_new_n619_), .B(u0_u1__abc_72579_new_n634_), .Y(u0_u1__abc_72579_new_n635_));
AND2X2 AND2X2_2241 ( .A(u0_u1__abc_72579_new_n635_), .B(u0_u1__abc_72579_new_n604_), .Y(u0_u1__abc_72579_new_n636_));
AND2X2 AND2X2_2242 ( .A(u0_u1__abc_72579_new_n636_), .B(u0_u1__abc_72579_new_n596_), .Y(u0_u1__abc_72579_new_n637_));
AND2X2 AND2X2_2243 ( .A(u0_u1__abc_72579_new_n637_), .B(u0_u1__abc_72579_new_n573_), .Y(u0_u1_wp_err));
AND2X2 AND2X2_2244 ( .A(u0_u1__abc_72579_new_n637_), .B(u0_u1__abc_72579_new_n639_), .Y(u0_cs1));
AND2X2 AND2X2_2245 ( .A(u0_u1__abc_72579_new_n642_), .B(u0_init_req1), .Y(u0_u1__abc_72579_new_n643_));
AND2X2 AND2X2_2246 ( .A(u0_u1__abc_72579_new_n644_), .B(u0_csc1_0_), .Y(u0_u1__abc_72579_new_n645_));
AND2X2 AND2X2_2247 ( .A(u0_u1__abc_72579_new_n645_), .B(u0_u1_init_req_we), .Y(u0_u1__abc_72579_new_n646_));
AND2X2 AND2X2_2248 ( .A(u0_u1__abc_72579_new_n203_), .B(u0_u1__abc_72579_new_n646_), .Y(u0_u1__abc_72579_new_n647_));
AND2X2 AND2X2_2249 ( .A(u1__abc_73140_new_n265_), .B(u1__abc_73140_new_n260_), .Y(u1__abc_73140_new_n266_));
AND2X2 AND2X2_225 ( .A(u0__abc_76628_new_n1170__bF_buf4), .B(sp_tms_9_), .Y(u0__abc_76628_new_n1394_));
AND2X2 AND2X2_2250 ( .A(u1__abc_73140_new_n267_), .B(csc_s_4_), .Y(u1__abc_73140_new_n268_));
AND2X2 AND2X2_2251 ( .A(u1__abc_73140_new_n263_), .B(csc_s_7_), .Y(u1__abc_73140_new_n269_));
AND2X2 AND2X2_2252 ( .A(u1__abc_73140_new_n268__bF_buf4), .B(u1__abc_73140_new_n269_), .Y(u1__abc_73140_new_n270_));
AND2X2 AND2X2_2253 ( .A(u1__abc_73140_new_n266_), .B(u1__abc_73140_new_n271_), .Y(u1__abc_73140_new_n272_));
AND2X2 AND2X2_2254 ( .A(u1__abc_73140_new_n273_), .B(u1__abc_73140_new_n268__bF_buf3), .Y(u1__abc_73140_new_n274_));
AND2X2 AND2X2_2255 ( .A(u1__abc_73140_new_n261_), .B(csc_s_5_), .Y(u1__abc_73140_new_n275_));
AND2X2 AND2X2_2256 ( .A(csc_s_7_), .B(csc_s_6_), .Y(u1__abc_73140_new_n276_));
AND2X2 AND2X2_2257 ( .A(u1__abc_73140_new_n277_), .B(u1__abc_73140_new_n275__bF_buf4), .Y(u1__abc_73140_new_n278_));
AND2X2 AND2X2_2258 ( .A(u1__abc_73140_new_n272_), .B(u1__abc_73140_new_n280_), .Y(page_size_10_));
AND2X2 AND2X2_2259 ( .A(u1__abc_73140_new_n282_), .B(bank_adr_0_), .Y(u1__abc_73140_new_n283_));
AND2X2 AND2X2_226 ( .A(spec_req_cs_5_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1395_));
AND2X2 AND2X2_2260 ( .A(page_size_10_), .B(\wb_addr_i[12] ), .Y(u1__abc_73140_new_n284_));
AND2X2 AND2X2_2261 ( .A(page_size_8_), .B(\wb_addr_i[10] ), .Y(u1__abc_73140_new_n285_));
AND2X2 AND2X2_2262 ( .A(page_size_9_), .B(\wb_addr_i[11] ), .Y(u1__abc_73140_new_n287_));
AND2X2 AND2X2_2263 ( .A(u1__abc_73140_new_n269_), .B(u1__abc_73140_new_n275__bF_buf3), .Y(u1__abc_73140_new_n292_));
AND2X2 AND2X2_2264 ( .A(u1__abc_73140_new_n296_), .B(u1__abc_73140_new_n271_), .Y(u1__abc_73140_new_n297_));
AND2X2 AND2X2_2265 ( .A(u1__abc_73140_new_n298_), .B(csc_s_6_), .Y(u1__abc_73140_new_n299_));
AND2X2 AND2X2_2266 ( .A(u1__abc_73140_new_n299_), .B(u1__abc_73140_new_n275__bF_buf1), .Y(u1__abc_73140_new_n300_));
AND2X2 AND2X2_2267 ( .A(u1__abc_73140_new_n303_), .B(u1__abc_73140_new_n299_), .Y(u1__abc_73140_new_n304_));
AND2X2 AND2X2_2268 ( .A(u1__abc_73140_new_n302_), .B(u1__abc_73140_new_n305_), .Y(u1__abc_73140_new_n306_));
AND2X2 AND2X2_2269 ( .A(u1__abc_73140_new_n306_), .B(u1__abc_73140_new_n297_), .Y(u1__abc_73140_new_n307_));
AND2X2 AND2X2_227 ( .A(u0__abc_76628_new_n1397_), .B(u0__abc_76628_new_n1179__bF_buf2), .Y(u0__abc_76628_new_n1398_));
AND2X2 AND2X2_2270 ( .A(u1__abc_73140_new_n307_), .B(u1__abc_73140_new_n294_), .Y(u1__abc_73140_new_n308_));
AND2X2 AND2X2_2271 ( .A(u1__abc_73140_new_n308_), .B(\wb_addr_i[25] ), .Y(u1__abc_73140_new_n309_));
AND2X2 AND2X2_2272 ( .A(u1__abc_73140_new_n293_), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n310_));
AND2X2 AND2X2_2273 ( .A(u1__abc_73140_new_n311_), .B(\wb_addr_i[24] ), .Y(u1__abc_73140_new_n312_));
AND2X2 AND2X2_2274 ( .A(u1__abc_73140_new_n301_), .B(\wb_addr_i[22] ), .Y(u1__abc_73140_new_n313_));
AND2X2 AND2X2_2275 ( .A(u1__abc_73140_new_n275__bF_buf0), .B(\wb_addr_i[21] ), .Y(u1__abc_73140_new_n315_));
AND2X2 AND2X2_2276 ( .A(u1__abc_73140_new_n315_), .B(u1__abc_73140_new_n273_), .Y(u1__abc_73140_new_n316_));
AND2X2 AND2X2_2277 ( .A(u1__abc_73140_new_n321_), .B(cs_le_bF_buf3), .Y(u1__abc_73140_new_n322_));
AND2X2 AND2X2_2278 ( .A(u1__abc_73140_new_n322_), .B(u1__abc_73140_new_n290_), .Y(u1__abc_73140_new_n323_));
AND2X2 AND2X2_2279 ( .A(u1__abc_73140_new_n282_), .B(bank_adr_1_), .Y(u1__abc_73140_new_n325_));
AND2X2 AND2X2_228 ( .A(u0__abc_76628_new_n1398_), .B(u0__abc_76628_new_n1396_), .Y(u0__abc_76628_new_n1399_));
AND2X2 AND2X2_2280 ( .A(page_size_10_), .B(\wb_addr_i[13] ), .Y(u1__abc_73140_new_n326_));
AND2X2 AND2X2_2281 ( .A(page_size_8_), .B(\wb_addr_i[11] ), .Y(u1__abc_73140_new_n327_));
AND2X2 AND2X2_2282 ( .A(page_size_9_), .B(\wb_addr_i[12] ), .Y(u1__abc_73140_new_n328_));
AND2X2 AND2X2_2283 ( .A(u1__abc_73140_new_n308_), .B(\wb_addr_i[26] ), .Y(u1__abc_73140_new_n332_));
AND2X2 AND2X2_2284 ( .A(u1__abc_73140_new_n293_), .B(\wb_addr_i[24] ), .Y(u1__abc_73140_new_n333_));
AND2X2 AND2X2_2285 ( .A(u1__abc_73140_new_n301_), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n334_));
AND2X2 AND2X2_2286 ( .A(u1__abc_73140_new_n311_), .B(\wb_addr_i[25] ), .Y(u1__abc_73140_new_n335_));
AND2X2 AND2X2_2287 ( .A(u1__abc_73140_new_n275__bF_buf4), .B(\wb_addr_i[22] ), .Y(u1__abc_73140_new_n336_));
AND2X2 AND2X2_2288 ( .A(u1__abc_73140_new_n336_), .B(u1__abc_73140_new_n273_), .Y(u1__abc_73140_new_n337_));
AND2X2 AND2X2_2289 ( .A(u1__abc_73140_new_n342_), .B(cs_le_bF_buf2), .Y(u1__abc_73140_new_n343_));
AND2X2 AND2X2_229 ( .A(u0__abc_76628_new_n1400_), .B(u0__abc_76628_new_n1175__bF_buf2), .Y(u0__abc_76628_new_n1401_));
AND2X2 AND2X2_2290 ( .A(u1__abc_73140_new_n343_), .B(u1__abc_73140_new_n331_), .Y(u1__abc_73140_new_n344_));
AND2X2 AND2X2_2291 ( .A(u1__abc_73140_new_n282_), .B(row_adr_0_bF_buf3_), .Y(u1__abc_73140_new_n346_));
AND2X2 AND2X2_2292 ( .A(page_size_10_), .B(\wb_addr_i[14] ), .Y(u1__abc_73140_new_n347_));
AND2X2 AND2X2_2293 ( .A(page_size_8_), .B(\wb_addr_i[12] ), .Y(u1__abc_73140_new_n348_));
AND2X2 AND2X2_2294 ( .A(page_size_9_), .B(\wb_addr_i[13] ), .Y(u1__abc_73140_new_n349_));
AND2X2 AND2X2_2295 ( .A(u1__abc_73140_new_n353_), .B(cs_le_bF_buf1), .Y(u1__abc_73140_new_n354_));
AND2X2 AND2X2_2296 ( .A(u1__abc_73140_new_n354_), .B(u1__abc_73140_new_n352_), .Y(u1__abc_73140_new_n355_));
AND2X2 AND2X2_2297 ( .A(u1__abc_73140_new_n282_), .B(row_adr_1_bF_buf3_), .Y(u1__abc_73140_new_n357_));
AND2X2 AND2X2_2298 ( .A(u1__abc_73140_new_n303_), .B(u1__abc_73140_new_n269_), .Y(u1__abc_73140_new_n360_));
AND2X2 AND2X2_2299 ( .A(u1__abc_73140_new_n266_), .B(u1__abc_73140_new_n361_), .Y(u1__abc_73140_new_n362_));
AND2X2 AND2X2_23 ( .A(_abc_85006_new_n305_), .B(_abc_85006_new_n306_), .Y(tms_s_5_));
AND2X2 AND2X2_230 ( .A(spec_req_cs_4_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1402_));
AND2X2 AND2X2_2300 ( .A(u1__abc_73140_new_n362_), .B(u1__abc_73140_new_n297_), .Y(u1__abc_73140_new_n363_));
AND2X2 AND2X2_2301 ( .A(u1__abc_73140_new_n363_), .B(u1__abc_73140_new_n359_), .Y(u1__abc_73140_new_n364_));
AND2X2 AND2X2_2302 ( .A(u1__abc_73140_new_n364_), .B(\wb_addr_i[15] ), .Y(u1__abc_73140_new_n365_));
AND2X2 AND2X2_2303 ( .A(page_size_9_), .B(\wb_addr_i[14] ), .Y(u1__abc_73140_new_n366_));
AND2X2 AND2X2_2304 ( .A(u1__abc_73140_new_n360_), .B(\wb_addr_i[15] ), .Y(u1__abc_73140_new_n367_));
AND2X2 AND2X2_2305 ( .A(page_size_8_), .B(\wb_addr_i[13] ), .Y(u1__abc_73140_new_n368_));
AND2X2 AND2X2_2306 ( .A(u1__abc_73140_new_n373_), .B(cs_le_bF_buf0), .Y(u1__abc_73140_new_n374_));
AND2X2 AND2X2_2307 ( .A(u1__abc_73140_new_n374_), .B(u1__abc_73140_new_n372_), .Y(u1__abc_73140_new_n375_));
AND2X2 AND2X2_2308 ( .A(u1__abc_73140_new_n282_), .B(row_adr_2_bF_buf3_), .Y(u1__abc_73140_new_n377_));
AND2X2 AND2X2_2309 ( .A(u1__abc_73140_new_n364_), .B(\wb_addr_i[16] ), .Y(u1__abc_73140_new_n379_));
AND2X2 AND2X2_231 ( .A(u0__abc_76628_new_n1403_), .B(u0__abc_76628_new_n1174__bF_buf2), .Y(u0__abc_76628_new_n1404_));
AND2X2 AND2X2_2310 ( .A(page_size_9_), .B(\wb_addr_i[15] ), .Y(u1__abc_73140_new_n380_));
AND2X2 AND2X2_2311 ( .A(u1__abc_73140_new_n360_), .B(\wb_addr_i[16] ), .Y(u1__abc_73140_new_n381_));
AND2X2 AND2X2_2312 ( .A(page_size_8_), .B(\wb_addr_i[14] ), .Y(u1__abc_73140_new_n382_));
AND2X2 AND2X2_2313 ( .A(u1__abc_73140_new_n386_), .B(cs_le_bF_buf4), .Y(u1__abc_73140_new_n387_));
AND2X2 AND2X2_2314 ( .A(u1__abc_73140_new_n387_), .B(u1__abc_73140_new_n378_), .Y(u1__abc_73140_new_n388_));
AND2X2 AND2X2_2315 ( .A(u1__abc_73140_new_n282_), .B(row_adr_3_bF_buf3_), .Y(u1__abc_73140_new_n390_));
AND2X2 AND2X2_2316 ( .A(u1__abc_73140_new_n364_), .B(\wb_addr_i[17] ), .Y(u1__abc_73140_new_n392_));
AND2X2 AND2X2_2317 ( .A(page_size_9_), .B(\wb_addr_i[16] ), .Y(u1__abc_73140_new_n393_));
AND2X2 AND2X2_2318 ( .A(u1__abc_73140_new_n360_), .B(\wb_addr_i[17] ), .Y(u1__abc_73140_new_n394_));
AND2X2 AND2X2_2319 ( .A(page_size_8_), .B(\wb_addr_i[15] ), .Y(u1__abc_73140_new_n395_));
AND2X2 AND2X2_232 ( .A(spec_req_cs_3_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1405_));
AND2X2 AND2X2_2320 ( .A(u1__abc_73140_new_n399_), .B(cs_le_bF_buf3), .Y(u1__abc_73140_new_n400_));
AND2X2 AND2X2_2321 ( .A(u1__abc_73140_new_n400_), .B(u1__abc_73140_new_n391_), .Y(u1__abc_73140_new_n401_));
AND2X2 AND2X2_2322 ( .A(u1__abc_73140_new_n282_), .B(row_adr_4_bF_buf3_), .Y(u1__abc_73140_new_n403_));
AND2X2 AND2X2_2323 ( .A(u1__abc_73140_new_n364_), .B(\wb_addr_i[18] ), .Y(u1__abc_73140_new_n404_));
AND2X2 AND2X2_2324 ( .A(page_size_9_), .B(\wb_addr_i[17] ), .Y(u1__abc_73140_new_n405_));
AND2X2 AND2X2_2325 ( .A(u1__abc_73140_new_n360_), .B(\wb_addr_i[18] ), .Y(u1__abc_73140_new_n406_));
AND2X2 AND2X2_2326 ( .A(page_size_8_), .B(\wb_addr_i[16] ), .Y(u1__abc_73140_new_n407_));
AND2X2 AND2X2_2327 ( .A(u1__abc_73140_new_n412_), .B(cs_le_bF_buf2), .Y(u1__abc_73140_new_n413_));
AND2X2 AND2X2_2328 ( .A(u1__abc_73140_new_n413_), .B(u1__abc_73140_new_n411_), .Y(u1__abc_73140_new_n414_));
AND2X2 AND2X2_2329 ( .A(u1__abc_73140_new_n282_), .B(row_adr_5_bF_buf3_), .Y(u1__abc_73140_new_n416_));
AND2X2 AND2X2_233 ( .A(u0__abc_76628_new_n1406_), .B(u0__abc_76628_new_n1173__bF_buf2), .Y(u0__abc_76628_new_n1407_));
AND2X2 AND2X2_2330 ( .A(u1__abc_73140_new_n364_), .B(\wb_addr_i[19] ), .Y(u1__abc_73140_new_n418_));
AND2X2 AND2X2_2331 ( .A(page_size_9_), .B(\wb_addr_i[18] ), .Y(u1__abc_73140_new_n419_));
AND2X2 AND2X2_2332 ( .A(u1__abc_73140_new_n360_), .B(\wb_addr_i[19] ), .Y(u1__abc_73140_new_n420_));
AND2X2 AND2X2_2333 ( .A(page_size_8_), .B(\wb_addr_i[17] ), .Y(u1__abc_73140_new_n421_));
AND2X2 AND2X2_2334 ( .A(u1__abc_73140_new_n425_), .B(cs_le_bF_buf1), .Y(u1__abc_73140_new_n426_));
AND2X2 AND2X2_2335 ( .A(u1__abc_73140_new_n426_), .B(u1__abc_73140_new_n417_), .Y(u1__abc_73140_new_n427_));
AND2X2 AND2X2_2336 ( .A(u1__abc_73140_new_n282_), .B(row_adr_6_bF_buf3_), .Y(u1__abc_73140_new_n429_));
AND2X2 AND2X2_2337 ( .A(u1__abc_73140_new_n364_), .B(\wb_addr_i[20] ), .Y(u1__abc_73140_new_n431_));
AND2X2 AND2X2_2338 ( .A(page_size_9_), .B(\wb_addr_i[19] ), .Y(u1__abc_73140_new_n432_));
AND2X2 AND2X2_2339 ( .A(u1__abc_73140_new_n360_), .B(\wb_addr_i[20] ), .Y(u1__abc_73140_new_n433_));
AND2X2 AND2X2_234 ( .A(spec_req_cs_2_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1408_));
AND2X2 AND2X2_2340 ( .A(page_size_8_), .B(\wb_addr_i[18] ), .Y(u1__abc_73140_new_n434_));
AND2X2 AND2X2_2341 ( .A(u1__abc_73140_new_n438_), .B(cs_le_bF_buf0), .Y(u1__abc_73140_new_n439_));
AND2X2 AND2X2_2342 ( .A(u1__abc_73140_new_n439_), .B(u1__abc_73140_new_n430_), .Y(u1__abc_73140_new_n440_));
AND2X2 AND2X2_2343 ( .A(u1__abc_73140_new_n282_), .B(row_adr_7_bF_buf3_), .Y(u1__abc_73140_new_n442_));
AND2X2 AND2X2_2344 ( .A(page_size_10_), .B(\wb_addr_i[21] ), .Y(u1__abc_73140_new_n444_));
AND2X2 AND2X2_2345 ( .A(page_size_9_), .B(\wb_addr_i[20] ), .Y(u1__abc_73140_new_n445_));
AND2X2 AND2X2_2346 ( .A(page_size_8_), .B(\wb_addr_i[19] ), .Y(u1__abc_73140_new_n446_));
AND2X2 AND2X2_2347 ( .A(u1__abc_73140_new_n449_), .B(cs_le_bF_buf4), .Y(u1__abc_73140_new_n450_));
AND2X2 AND2X2_2348 ( .A(u1__abc_73140_new_n450_), .B(u1__abc_73140_new_n443_), .Y(u1__abc_73140_new_n451_));
AND2X2 AND2X2_2349 ( .A(u1__abc_73140_new_n282_), .B(row_adr_8_bF_buf3_), .Y(u1__abc_73140_new_n453_));
AND2X2 AND2X2_235 ( .A(u0__abc_76628_new_n1409_), .B(u0__abc_76628_new_n1172__bF_buf2), .Y(u0__abc_76628_new_n1410_));
AND2X2 AND2X2_2350 ( .A(page_size_10_), .B(\wb_addr_i[22] ), .Y(u1__abc_73140_new_n455_));
AND2X2 AND2X2_2351 ( .A(page_size_9_), .B(\wb_addr_i[21] ), .Y(u1__abc_73140_new_n456_));
AND2X2 AND2X2_2352 ( .A(page_size_8_), .B(\wb_addr_i[20] ), .Y(u1__abc_73140_new_n457_));
AND2X2 AND2X2_2353 ( .A(u1__abc_73140_new_n460_), .B(cs_le_bF_buf3), .Y(u1__abc_73140_new_n461_));
AND2X2 AND2X2_2354 ( .A(u1__abc_73140_new_n461_), .B(u1__abc_73140_new_n454_), .Y(u1__abc_73140_new_n462_));
AND2X2 AND2X2_2355 ( .A(u1__abc_73140_new_n282_), .B(row_adr_9_bF_buf3_), .Y(u1__abc_73140_new_n464_));
AND2X2 AND2X2_2356 ( .A(u1__abc_73140_new_n364_), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n466_));
AND2X2 AND2X2_2357 ( .A(u1__abc_73140_new_n358_), .B(\wb_addr_i[21] ), .Y(u1__abc_73140_new_n467_));
AND2X2 AND2X2_2358 ( .A(u1__abc_73140_new_n270_), .B(\wb_addr_i[22] ), .Y(u1__abc_73140_new_n468_));
AND2X2 AND2X2_2359 ( .A(u1__abc_73140_new_n360_), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n470_));
AND2X2 AND2X2_236 ( .A(spec_req_cs_1_bF_buf5_), .B(u0_tms1_9_), .Y(u0__abc_76628_new_n1411_));
AND2X2 AND2X2_2360 ( .A(u1__abc_73140_new_n291_), .B(\wb_addr_i[22] ), .Y(u1__abc_73140_new_n471_));
AND2X2 AND2X2_2361 ( .A(u1__abc_73140_new_n476_), .B(cs_le_bF_buf2), .Y(u1__abc_73140_new_n477_));
AND2X2 AND2X2_2362 ( .A(u1__abc_73140_new_n477_), .B(u1__abc_73140_new_n465_), .Y(u1__abc_73140_new_n478_));
AND2X2 AND2X2_2363 ( .A(u1__abc_73140_new_n282_), .B(row_adr_10_bF_buf3_), .Y(u1__abc_73140_new_n480_));
AND2X2 AND2X2_2364 ( .A(u1__abc_73140_new_n364_), .B(\wb_addr_i[24] ), .Y(u1__abc_73140_new_n482_));
AND2X2 AND2X2_2365 ( .A(u1__abc_73140_new_n336_), .B(u1__abc_73140_new_n269_), .Y(u1__abc_73140_new_n483_));
AND2X2 AND2X2_2366 ( .A(u1__abc_73140_new_n360_), .B(\wb_addr_i[24] ), .Y(u1__abc_73140_new_n486_));
AND2X2 AND2X2_2367 ( .A(u1__abc_73140_new_n268__bF_buf2), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n487_));
AND2X2 AND2X2_2368 ( .A(u1__abc_73140_new_n487_), .B(u1__abc_73140_new_n269_), .Y(u1__abc_73140_new_n488_));
AND2X2 AND2X2_2369 ( .A(u1__abc_73140_new_n291_), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n490_));
AND2X2 AND2X2_237 ( .A(u0__abc_76628_new_n1169__bF_buf3), .B(u0__abc_76628_new_n1414_), .Y(u0__abc_76628_new_n1415_));
AND2X2 AND2X2_2370 ( .A(u1__abc_73140_new_n494_), .B(cs_le_bF_buf1), .Y(u1__abc_73140_new_n495_));
AND2X2 AND2X2_2371 ( .A(u1__abc_73140_new_n495_), .B(u1__abc_73140_new_n481_), .Y(u1__abc_73140_new_n496_));
AND2X2 AND2X2_2372 ( .A(u1__abc_73140_new_n282_), .B(row_adr_11_bF_buf3_), .Y(u1__abc_73140_new_n498_));
AND2X2 AND2X2_2373 ( .A(page_size_10_), .B(\wb_addr_i[25] ), .Y(u1__abc_73140_new_n502_));
AND2X2 AND2X2_2374 ( .A(page_size_9_), .B(\wb_addr_i[24] ), .Y(u1__abc_73140_new_n503_));
AND2X2 AND2X2_2375 ( .A(u1__abc_73140_new_n358_), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n504_));
AND2X2 AND2X2_2376 ( .A(u1__abc_73140_new_n507_), .B(cs_le_bF_buf0), .Y(u1__abc_73140_new_n508_));
AND2X2 AND2X2_2377 ( .A(u1__abc_73140_new_n508_), .B(u1__abc_73140_new_n501_), .Y(u1__abc_73140_new_n509_));
AND2X2 AND2X2_2378 ( .A(u1__abc_73140_new_n270_), .B(\wb_addr_i[25] ), .Y(u1__abc_73140_new_n511_));
AND2X2 AND2X2_2379 ( .A(u1__abc_73140_new_n360_), .B(\wb_addr_i[26] ), .Y(u1__abc_73140_new_n513_));
AND2X2 AND2X2_238 ( .A(u0__abc_76628_new_n1413_), .B(u0__abc_76628_new_n1415_), .Y(u0__abc_76628_new_n1416_));
AND2X2 AND2X2_2380 ( .A(u1__abc_73140_new_n275__bF_buf3), .B(\wb_addr_i[24] ), .Y(u1__abc_73140_new_n514_));
AND2X2 AND2X2_2381 ( .A(u1__abc_73140_new_n514_), .B(u1__abc_73140_new_n269_), .Y(u1__abc_73140_new_n515_));
AND2X2 AND2X2_2382 ( .A(u1__abc_73140_new_n517_), .B(u1__abc_73140_new_n519_), .Y(u1__abc_73140_new_n520_));
AND2X2 AND2X2_2383 ( .A(u1__abc_73140_new_n521_), .B(u1__abc_73140_new_n522_), .Y(u1__0row_adr_12_0__12_));
AND2X2 AND2X2_2384 ( .A(u1__abc_73140_new_n524_), .B(wb_stb_i_bF_buf3), .Y(u1__abc_73140_new_n525_));
AND2X2 AND2X2_2385 ( .A(mem_ack_r), .B(u1_wr_cycle), .Y(u1__abc_73140_new_n526_));
AND2X2 AND2X2_2386 ( .A(u1__abc_73140_new_n529_), .B(u1__abc_73140_new_n530_), .Y(u1__0col_adr_9_0__0_));
AND2X2 AND2X2_2387 ( .A(u1__abc_73140_new_n532_), .B(u1__abc_73140_new_n533_), .Y(u1__0col_adr_9_0__1_));
AND2X2 AND2X2_2388 ( .A(u1__abc_73140_new_n535_), .B(u1__abc_73140_new_n536_), .Y(u1__0col_adr_9_0__2_));
AND2X2 AND2X2_2389 ( .A(u1__abc_73140_new_n538_), .B(u1__abc_73140_new_n539_), .Y(u1__0col_adr_9_0__3_));
AND2X2 AND2X2_239 ( .A(u0__abc_76628_new_n1170__bF_buf3), .B(sp_tms_10_), .Y(u0__abc_76628_new_n1418_));
AND2X2 AND2X2_2390 ( .A(u1__abc_73140_new_n541_), .B(u1__abc_73140_new_n542_), .Y(u1__0col_adr_9_0__4_));
AND2X2 AND2X2_2391 ( .A(u1__abc_73140_new_n544_), .B(u1__abc_73140_new_n545_), .Y(u1__0col_adr_9_0__5_));
AND2X2 AND2X2_2392 ( .A(u1__abc_73140_new_n547_), .B(u1__abc_73140_new_n548_), .Y(u1__0col_adr_9_0__6_));
AND2X2 AND2X2_2393 ( .A(u1__abc_73140_new_n550_), .B(u1__abc_73140_new_n551_), .Y(u1__0col_adr_9_0__7_));
AND2X2 AND2X2_2394 ( .A(u1__abc_73140_new_n528_), .B(u1_col_adr_8_), .Y(u1__abc_73140_new_n553_));
AND2X2 AND2X2_2395 ( .A(u1__abc_73140_new_n527_), .B(\wb_addr_i[10] ), .Y(u1__abc_73140_new_n554_));
AND2X2 AND2X2_2396 ( .A(u1__abc_73140_new_n280_), .B(u1__abc_73140_new_n554_), .Y(u1__abc_73140_new_n555_));
AND2X2 AND2X2_2397 ( .A(u1__abc_73140_new_n528_), .B(u1_col_adr_9_), .Y(u1__abc_73140_new_n557_));
AND2X2 AND2X2_2398 ( .A(u1__abc_73140_new_n527_), .B(\wb_addr_i[11] ), .Y(u1__abc_73140_new_n558_));
AND2X2 AND2X2_2399 ( .A(page_size_10_), .B(u1__abc_73140_new_n558_), .Y(u1__abc_73140_new_n559_));
AND2X2 AND2X2_24 ( .A(_abc_85006_new_n308_), .B(_abc_85006_new_n309_), .Y(tms_s_6_));
AND2X2 AND2X2_240 ( .A(spec_req_cs_5_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1419_));
AND2X2 AND2X2_2400 ( .A(u1__abc_73140_new_n564_), .B(u1__abc_73140_new_n562_), .Y(u1__abc_73140_new_n565_));
AND2X2 AND2X2_2401 ( .A(u1__abc_73140_new_n295_), .B(u1__abc_73140_new_n262_), .Y(u1__abc_73140_new_n567_));
AND2X2 AND2X2_2402 ( .A(u1__abc_73140_new_n567__bF_buf3), .B(\wb_addr_i[0] ), .Y(u1__abc_73140_new_n568_));
AND2X2 AND2X2_2403 ( .A(u1__abc_73140_new_n275__bF_buf2), .B(\wb_addr_i[2] ), .Y(u1__abc_73140_new_n569_));
AND2X2 AND2X2_2404 ( .A(u1__abc_73140_new_n268__bF_buf1), .B(\wb_addr_i[1] ), .Y(u1__abc_73140_new_n571_));
AND2X2 AND2X2_2405 ( .A(u1__abc_73140_new_n574_), .B(u1__abc_73140_new_n566_), .Y(u1__0acs_addr_23_0__0_));
AND2X2 AND2X2_2406 ( .A(u1__abc_73140_new_n577_), .B(u1__abc_73140_new_n576_), .Y(u1__abc_73140_new_n578_));
AND2X2 AND2X2_2407 ( .A(u1__abc_73140_new_n567__bF_buf2), .B(\wb_addr_i[1] ), .Y(u1__abc_73140_new_n580_));
AND2X2 AND2X2_2408 ( .A(u1__abc_73140_new_n268__bF_buf0), .B(\wb_addr_i[2] ), .Y(u1__abc_73140_new_n581_));
AND2X2 AND2X2_2409 ( .A(u1__abc_73140_new_n275__bF_buf1), .B(\wb_addr_i[3] ), .Y(u1__abc_73140_new_n582_));
AND2X2 AND2X2_241 ( .A(u0__abc_76628_new_n1421_), .B(u0__abc_76628_new_n1179__bF_buf1), .Y(u0__abc_76628_new_n1422_));
AND2X2 AND2X2_2410 ( .A(u1__abc_73140_new_n585_), .B(u1__abc_73140_new_n579_), .Y(u1__0acs_addr_23_0__1_));
AND2X2 AND2X2_2411 ( .A(u1__abc_73140_new_n588_), .B(u1__abc_73140_new_n587_), .Y(u1__abc_73140_new_n589_));
AND2X2 AND2X2_2412 ( .A(u1__abc_73140_new_n567__bF_buf1), .B(\wb_addr_i[2] ), .Y(u1__abc_73140_new_n591_));
AND2X2 AND2X2_2413 ( .A(u1__abc_73140_new_n275__bF_buf0), .B(\wb_addr_i[4] ), .Y(u1__abc_73140_new_n592_));
AND2X2 AND2X2_2414 ( .A(u1__abc_73140_new_n268__bF_buf4), .B(\wb_addr_i[3] ), .Y(u1__abc_73140_new_n593_));
AND2X2 AND2X2_2415 ( .A(u1__abc_73140_new_n596_), .B(u1__abc_73140_new_n590_), .Y(u1__0acs_addr_23_0__2_));
AND2X2 AND2X2_2416 ( .A(u1__abc_73140_new_n599_), .B(u1__abc_73140_new_n598_), .Y(u1__abc_73140_new_n600_));
AND2X2 AND2X2_2417 ( .A(u1__abc_73140_new_n567__bF_buf0), .B(\wb_addr_i[3] ), .Y(u1__abc_73140_new_n602_));
AND2X2 AND2X2_2418 ( .A(u1__abc_73140_new_n275__bF_buf4), .B(\wb_addr_i[5] ), .Y(u1__abc_73140_new_n603_));
AND2X2 AND2X2_2419 ( .A(u1__abc_73140_new_n268__bF_buf3), .B(\wb_addr_i[4] ), .Y(u1__abc_73140_new_n604_));
AND2X2 AND2X2_242 ( .A(u0__abc_76628_new_n1422_), .B(u0__abc_76628_new_n1420_), .Y(u0__abc_76628_new_n1423_));
AND2X2 AND2X2_2420 ( .A(u1__abc_73140_new_n607_), .B(u1__abc_73140_new_n601_), .Y(u1__0acs_addr_23_0__3_));
AND2X2 AND2X2_2421 ( .A(u1__abc_73140_new_n610_), .B(u1__abc_73140_new_n609_), .Y(u1__abc_73140_new_n611_));
AND2X2 AND2X2_2422 ( .A(u1__abc_73140_new_n567__bF_buf3), .B(\wb_addr_i[4] ), .Y(u1__abc_73140_new_n613_));
AND2X2 AND2X2_2423 ( .A(u1__abc_73140_new_n275__bF_buf3), .B(\wb_addr_i[6] ), .Y(u1__abc_73140_new_n614_));
AND2X2 AND2X2_2424 ( .A(u1__abc_73140_new_n268__bF_buf2), .B(\wb_addr_i[5] ), .Y(u1__abc_73140_new_n615_));
AND2X2 AND2X2_2425 ( .A(u1__abc_73140_new_n618_), .B(u1__abc_73140_new_n612_), .Y(u1__0acs_addr_23_0__4_));
AND2X2 AND2X2_2426 ( .A(u1__abc_73140_new_n621_), .B(u1__abc_73140_new_n620_), .Y(u1__abc_73140_new_n622_));
AND2X2 AND2X2_2427 ( .A(u1__abc_73140_new_n567__bF_buf2), .B(\wb_addr_i[5] ), .Y(u1__abc_73140_new_n624_));
AND2X2 AND2X2_2428 ( .A(u1__abc_73140_new_n275__bF_buf2), .B(\wb_addr_i[7] ), .Y(u1__abc_73140_new_n625_));
AND2X2 AND2X2_2429 ( .A(u1__abc_73140_new_n268__bF_buf1), .B(\wb_addr_i[6] ), .Y(u1__abc_73140_new_n626_));
AND2X2 AND2X2_243 ( .A(u0__abc_76628_new_n1424_), .B(u0__abc_76628_new_n1175__bF_buf1), .Y(u0__abc_76628_new_n1425_));
AND2X2 AND2X2_2430 ( .A(u1__abc_73140_new_n629_), .B(u1__abc_73140_new_n623_), .Y(u1__0acs_addr_23_0__5_));
AND2X2 AND2X2_2431 ( .A(u1__abc_73140_new_n632_), .B(u1__abc_73140_new_n631_), .Y(u1__abc_73140_new_n633_));
AND2X2 AND2X2_2432 ( .A(u1__abc_73140_new_n567__bF_buf1), .B(\wb_addr_i[6] ), .Y(u1__abc_73140_new_n635_));
AND2X2 AND2X2_2433 ( .A(u1__abc_73140_new_n268__bF_buf0), .B(\wb_addr_i[7] ), .Y(u1__abc_73140_new_n636_));
AND2X2 AND2X2_2434 ( .A(u1__abc_73140_new_n275__bF_buf1), .B(\wb_addr_i[8] ), .Y(u1__abc_73140_new_n637_));
AND2X2 AND2X2_2435 ( .A(u1__abc_73140_new_n640_), .B(u1__abc_73140_new_n634_), .Y(u1__0acs_addr_23_0__6_));
AND2X2 AND2X2_2436 ( .A(u1__abc_73140_new_n643_), .B(u1__abc_73140_new_n642_), .Y(u1__abc_73140_new_n644_));
AND2X2 AND2X2_2437 ( .A(u1__abc_73140_new_n567__bF_buf0), .B(\wb_addr_i[7] ), .Y(u1__abc_73140_new_n646_));
AND2X2 AND2X2_2438 ( .A(u1__abc_73140_new_n275__bF_buf0), .B(\wb_addr_i[9] ), .Y(u1__abc_73140_new_n647_));
AND2X2 AND2X2_2439 ( .A(u1__abc_73140_new_n268__bF_buf4), .B(\wb_addr_i[8] ), .Y(u1__abc_73140_new_n648_));
AND2X2 AND2X2_244 ( .A(spec_req_cs_4_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1426_));
AND2X2 AND2X2_2440 ( .A(u1__abc_73140_new_n651_), .B(u1__abc_73140_new_n645_), .Y(u1__0acs_addr_23_0__7_));
AND2X2 AND2X2_2441 ( .A(u1__abc_73140_new_n654_), .B(u1__abc_73140_new_n653_), .Y(u1__abc_73140_new_n655_));
AND2X2 AND2X2_2442 ( .A(u1__abc_73140_new_n567__bF_buf3), .B(\wb_addr_i[8] ), .Y(u1__abc_73140_new_n657_));
AND2X2 AND2X2_2443 ( .A(u1__abc_73140_new_n275__bF_buf4), .B(\wb_addr_i[10] ), .Y(u1__abc_73140_new_n658_));
AND2X2 AND2X2_2444 ( .A(u1__abc_73140_new_n268__bF_buf3), .B(\wb_addr_i[9] ), .Y(u1__abc_73140_new_n659_));
AND2X2 AND2X2_2445 ( .A(u1__abc_73140_new_n662_), .B(u1__abc_73140_new_n656_), .Y(u1__0acs_addr_23_0__8_));
AND2X2 AND2X2_2446 ( .A(u1__abc_73140_new_n665_), .B(u1__abc_73140_new_n664_), .Y(u1__abc_73140_new_n666_));
AND2X2 AND2X2_2447 ( .A(u1__abc_73140_new_n567__bF_buf2), .B(\wb_addr_i[9] ), .Y(u1__abc_73140_new_n668_));
AND2X2 AND2X2_2448 ( .A(u1__abc_73140_new_n268__bF_buf2), .B(\wb_addr_i[10] ), .Y(u1__abc_73140_new_n669_));
AND2X2 AND2X2_2449 ( .A(u1__abc_73140_new_n275__bF_buf3), .B(\wb_addr_i[11] ), .Y(u1__abc_73140_new_n670_));
AND2X2 AND2X2_245 ( .A(u0__abc_76628_new_n1427_), .B(u0__abc_76628_new_n1174__bF_buf1), .Y(u0__abc_76628_new_n1428_));
AND2X2 AND2X2_2450 ( .A(u1__abc_73140_new_n673_), .B(u1__abc_73140_new_n667_), .Y(u1__0acs_addr_23_0__9_));
AND2X2 AND2X2_2451 ( .A(u1__abc_73140_new_n676_), .B(u1__abc_73140_new_n675_), .Y(u1__abc_73140_new_n677_));
AND2X2 AND2X2_2452 ( .A(u1__abc_73140_new_n567__bF_buf1), .B(\wb_addr_i[10] ), .Y(u1__abc_73140_new_n679_));
AND2X2 AND2X2_2453 ( .A(u1__abc_73140_new_n275__bF_buf2), .B(\wb_addr_i[12] ), .Y(u1__abc_73140_new_n680_));
AND2X2 AND2X2_2454 ( .A(u1__abc_73140_new_n268__bF_buf1), .B(\wb_addr_i[11] ), .Y(u1__abc_73140_new_n681_));
AND2X2 AND2X2_2455 ( .A(u1__abc_73140_new_n684_), .B(u1__abc_73140_new_n678_), .Y(u1__0acs_addr_23_0__10_));
AND2X2 AND2X2_2456 ( .A(u1__abc_73140_new_n687_), .B(u1__abc_73140_new_n686_), .Y(u1__abc_73140_new_n688_));
AND2X2 AND2X2_2457 ( .A(u1__abc_73140_new_n567__bF_buf0), .B(\wb_addr_i[11] ), .Y(u1__abc_73140_new_n690_));
AND2X2 AND2X2_2458 ( .A(u1__abc_73140_new_n275__bF_buf1), .B(\wb_addr_i[13] ), .Y(u1__abc_73140_new_n691_));
AND2X2 AND2X2_2459 ( .A(u1__abc_73140_new_n268__bF_buf0), .B(\wb_addr_i[12] ), .Y(u1__abc_73140_new_n692_));
AND2X2 AND2X2_246 ( .A(spec_req_cs_3_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1429_));
AND2X2 AND2X2_2460 ( .A(u1__abc_73140_new_n695_), .B(u1__abc_73140_new_n689_), .Y(u1__0acs_addr_23_0__11_));
AND2X2 AND2X2_2461 ( .A(u1__abc_73140_new_n698_), .B(u1__abc_73140_new_n697_), .Y(u1__abc_73140_new_n699_));
AND2X2 AND2X2_2462 ( .A(u1__abc_73140_new_n567__bF_buf3), .B(\wb_addr_i[12] ), .Y(u1__abc_73140_new_n701_));
AND2X2 AND2X2_2463 ( .A(u1__abc_73140_new_n275__bF_buf0), .B(\wb_addr_i[14] ), .Y(u1__abc_73140_new_n702_));
AND2X2 AND2X2_2464 ( .A(u1__abc_73140_new_n268__bF_buf4), .B(\wb_addr_i[13] ), .Y(u1__abc_73140_new_n703_));
AND2X2 AND2X2_2465 ( .A(u1__abc_73140_new_n706_), .B(u1__abc_73140_new_n700_), .Y(u1__0acs_addr_23_0__12_));
AND2X2 AND2X2_2466 ( .A(u1__abc_73140_new_n709_), .B(u1__abc_73140_new_n708_), .Y(u1__abc_73140_new_n710_));
AND2X2 AND2X2_2467 ( .A(u1__abc_73140_new_n567__bF_buf2), .B(\wb_addr_i[13] ), .Y(u1__abc_73140_new_n712_));
AND2X2 AND2X2_2468 ( .A(u1__abc_73140_new_n275__bF_buf4), .B(\wb_addr_i[15] ), .Y(u1__abc_73140_new_n713_));
AND2X2 AND2X2_2469 ( .A(u1__abc_73140_new_n268__bF_buf3), .B(\wb_addr_i[14] ), .Y(u1__abc_73140_new_n714_));
AND2X2 AND2X2_247 ( .A(u0__abc_76628_new_n1430_), .B(u0__abc_76628_new_n1173__bF_buf1), .Y(u0__abc_76628_new_n1431_));
AND2X2 AND2X2_2470 ( .A(u1__abc_73140_new_n717_), .B(u1__abc_73140_new_n711_), .Y(u1__0acs_addr_23_0__13_));
AND2X2 AND2X2_2471 ( .A(u1__abc_73140_new_n720_), .B(u1__abc_73140_new_n719_), .Y(u1__abc_73140_new_n721_));
AND2X2 AND2X2_2472 ( .A(u1__abc_73140_new_n567__bF_buf1), .B(\wb_addr_i[14] ), .Y(u1__abc_73140_new_n723_));
AND2X2 AND2X2_2473 ( .A(u1__abc_73140_new_n268__bF_buf2), .B(\wb_addr_i[15] ), .Y(u1__abc_73140_new_n724_));
AND2X2 AND2X2_2474 ( .A(u1__abc_73140_new_n275__bF_buf3), .B(\wb_addr_i[16] ), .Y(u1__abc_73140_new_n725_));
AND2X2 AND2X2_2475 ( .A(u1__abc_73140_new_n728_), .B(u1__abc_73140_new_n722_), .Y(u1__0acs_addr_23_0__14_));
AND2X2 AND2X2_2476 ( .A(u1__abc_73140_new_n731_), .B(u1__abc_73140_new_n730_), .Y(u1__abc_73140_new_n732_));
AND2X2 AND2X2_2477 ( .A(u1__abc_73140_new_n567__bF_buf0), .B(\wb_addr_i[15] ), .Y(u1__abc_73140_new_n734_));
AND2X2 AND2X2_2478 ( .A(u1__abc_73140_new_n275__bF_buf2), .B(\wb_addr_i[17] ), .Y(u1__abc_73140_new_n735_));
AND2X2 AND2X2_2479 ( .A(u1__abc_73140_new_n268__bF_buf1), .B(\wb_addr_i[16] ), .Y(u1__abc_73140_new_n736_));
AND2X2 AND2X2_248 ( .A(spec_req_cs_2_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1432_));
AND2X2 AND2X2_2480 ( .A(u1__abc_73140_new_n739_), .B(u1__abc_73140_new_n733_), .Y(u1__0acs_addr_23_0__15_));
AND2X2 AND2X2_2481 ( .A(u1__abc_73140_new_n742_), .B(u1__abc_73140_new_n741_), .Y(u1__abc_73140_new_n743_));
AND2X2 AND2X2_2482 ( .A(u1__abc_73140_new_n567__bF_buf3), .B(\wb_addr_i[16] ), .Y(u1__abc_73140_new_n745_));
AND2X2 AND2X2_2483 ( .A(u1__abc_73140_new_n275__bF_buf1), .B(\wb_addr_i[18] ), .Y(u1__abc_73140_new_n746_));
AND2X2 AND2X2_2484 ( .A(u1__abc_73140_new_n268__bF_buf0), .B(\wb_addr_i[17] ), .Y(u1__abc_73140_new_n747_));
AND2X2 AND2X2_2485 ( .A(u1__abc_73140_new_n750_), .B(u1__abc_73140_new_n744_), .Y(u1__0acs_addr_23_0__16_));
AND2X2 AND2X2_2486 ( .A(u1__abc_73140_new_n753_), .B(u1__abc_73140_new_n752_), .Y(u1__abc_73140_new_n754_));
AND2X2 AND2X2_2487 ( .A(u1__abc_73140_new_n567__bF_buf2), .B(\wb_addr_i[17] ), .Y(u1__abc_73140_new_n756_));
AND2X2 AND2X2_2488 ( .A(u1__abc_73140_new_n268__bF_buf4), .B(\wb_addr_i[18] ), .Y(u1__abc_73140_new_n757_));
AND2X2 AND2X2_2489 ( .A(u1__abc_73140_new_n275__bF_buf0), .B(\wb_addr_i[19] ), .Y(u1__abc_73140_new_n758_));
AND2X2 AND2X2_249 ( .A(u0__abc_76628_new_n1433_), .B(u0__abc_76628_new_n1172__bF_buf1), .Y(u0__abc_76628_new_n1434_));
AND2X2 AND2X2_2490 ( .A(u1__abc_73140_new_n761_), .B(u1__abc_73140_new_n755_), .Y(u1__0acs_addr_23_0__17_));
AND2X2 AND2X2_2491 ( .A(u1__abc_73140_new_n764_), .B(u1__abc_73140_new_n763_), .Y(u1__abc_73140_new_n765_));
AND2X2 AND2X2_2492 ( .A(u1__abc_73140_new_n567__bF_buf1), .B(\wb_addr_i[18] ), .Y(u1__abc_73140_new_n767_));
AND2X2 AND2X2_2493 ( .A(u1__abc_73140_new_n275__bF_buf4), .B(\wb_addr_i[20] ), .Y(u1__abc_73140_new_n768_));
AND2X2 AND2X2_2494 ( .A(u1__abc_73140_new_n268__bF_buf3), .B(\wb_addr_i[19] ), .Y(u1__abc_73140_new_n769_));
AND2X2 AND2X2_2495 ( .A(u1__abc_73140_new_n772_), .B(u1__abc_73140_new_n766_), .Y(u1__0acs_addr_23_0__18_));
AND2X2 AND2X2_2496 ( .A(u1__abc_73140_new_n775_), .B(u1__abc_73140_new_n774_), .Y(u1__abc_73140_new_n776_));
AND2X2 AND2X2_2497 ( .A(u1__abc_73140_new_n567__bF_buf0), .B(\wb_addr_i[19] ), .Y(u1__abc_73140_new_n778_));
AND2X2 AND2X2_2498 ( .A(u1__abc_73140_new_n268__bF_buf2), .B(\wb_addr_i[20] ), .Y(u1__abc_73140_new_n779_));
AND2X2 AND2X2_2499 ( .A(u1__abc_73140_new_n782_), .B(u1__abc_73140_new_n777_), .Y(u1__0acs_addr_23_0__19_));
AND2X2 AND2X2_25 ( .A(_abc_85006_new_n311_), .B(_abc_85006_new_n312_), .Y(tms_s_7_));
AND2X2 AND2X2_250 ( .A(spec_req_cs_1_bF_buf4_), .B(u0_tms1_10_), .Y(u0__abc_76628_new_n1435_));
AND2X2 AND2X2_2500 ( .A(u1__abc_73140_new_n785_), .B(u1__abc_73140_new_n784_), .Y(u1__abc_73140_new_n786_));
AND2X2 AND2X2_2501 ( .A(u1__abc_73140_new_n567__bF_buf3), .B(\wb_addr_i[20] ), .Y(u1__abc_73140_new_n788_));
AND2X2 AND2X2_2502 ( .A(u1__abc_73140_new_n268__bF_buf1), .B(\wb_addr_i[21] ), .Y(u1__abc_73140_new_n789_));
AND2X2 AND2X2_2503 ( .A(u1__abc_73140_new_n792_), .B(u1__abc_73140_new_n787_), .Y(u1__0acs_addr_23_0__20_));
AND2X2 AND2X2_2504 ( .A(u1__abc_73140_new_n795_), .B(u1__abc_73140_new_n794_), .Y(u1__abc_73140_new_n796_));
AND2X2 AND2X2_2505 ( .A(u1__abc_73140_new_n567__bF_buf2), .B(\wb_addr_i[21] ), .Y(u1__abc_73140_new_n798_));
AND2X2 AND2X2_2506 ( .A(u1__abc_73140_new_n275__bF_buf3), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n799_));
AND2X2 AND2X2_2507 ( .A(u1__abc_73140_new_n268__bF_buf0), .B(\wb_addr_i[22] ), .Y(u1__abc_73140_new_n800_));
AND2X2 AND2X2_2508 ( .A(u1__abc_73140_new_n803_), .B(u1__abc_73140_new_n797_), .Y(u1__0acs_addr_23_0__21_));
AND2X2 AND2X2_2509 ( .A(u1__abc_73140_new_n806_), .B(u1__abc_73140_new_n805_), .Y(u1__abc_73140_new_n807_));
AND2X2 AND2X2_251 ( .A(u0__abc_76628_new_n1169__bF_buf2), .B(u0__abc_76628_new_n1438_), .Y(u0__abc_76628_new_n1439_));
AND2X2 AND2X2_2510 ( .A(u1__abc_73140_new_n567__bF_buf1), .B(\wb_addr_i[22] ), .Y(u1__abc_73140_new_n809_));
AND2X2 AND2X2_2511 ( .A(u1__abc_73140_new_n812_), .B(u1__abc_73140_new_n808_), .Y(u1__0acs_addr_23_0__22_));
AND2X2 AND2X2_2512 ( .A(u1__abc_73140_new_n815_), .B(u1__abc_73140_new_n814_), .Y(u1__abc_73140_new_n816_));
AND2X2 AND2X2_2513 ( .A(u1__abc_73140_new_n567__bF_buf0), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n818_));
AND2X2 AND2X2_2514 ( .A(u1__abc_73140_new_n268__bF_buf4), .B(\wb_addr_i[24] ), .Y(u1__abc_73140_new_n819_));
AND2X2 AND2X2_2515 ( .A(u1__abc_73140_new_n275__bF_buf2), .B(\wb_addr_i[25] ), .Y(u1__abc_73140_new_n820_));
AND2X2 AND2X2_2516 ( .A(u1__abc_73140_new_n823_), .B(u1__abc_73140_new_n817_), .Y(u1__0acs_addr_23_0__23_));
AND2X2 AND2X2_2517 ( .A(u1__abc_73140_new_n827_), .B(u1__abc_73140_new_n825_), .Y(u1__0sram_addr_23_0__0_));
AND2X2 AND2X2_2518 ( .A(u1__abc_73140_new_n830_), .B(u1__abc_73140_new_n829_), .Y(u1__0sram_addr_23_0__1_));
AND2X2 AND2X2_2519 ( .A(u1__abc_73140_new_n833_), .B(u1__abc_73140_new_n832_), .Y(u1__0sram_addr_23_0__2_));
AND2X2 AND2X2_252 ( .A(u0__abc_76628_new_n1437_), .B(u0__abc_76628_new_n1439_), .Y(u0__abc_76628_new_n1440_));
AND2X2 AND2X2_2520 ( .A(u1__abc_73140_new_n836_), .B(u1__abc_73140_new_n835_), .Y(u1__0sram_addr_23_0__3_));
AND2X2 AND2X2_2521 ( .A(u1__abc_73140_new_n839_), .B(u1__abc_73140_new_n838_), .Y(u1__0sram_addr_23_0__4_));
AND2X2 AND2X2_2522 ( .A(u1__abc_73140_new_n842_), .B(u1__abc_73140_new_n841_), .Y(u1__0sram_addr_23_0__5_));
AND2X2 AND2X2_2523 ( .A(u1__abc_73140_new_n845_), .B(u1__abc_73140_new_n844_), .Y(u1__0sram_addr_23_0__6_));
AND2X2 AND2X2_2524 ( .A(u1__abc_73140_new_n848_), .B(u1__abc_73140_new_n847_), .Y(u1__0sram_addr_23_0__7_));
AND2X2 AND2X2_2525 ( .A(u1__abc_73140_new_n851_), .B(u1__abc_73140_new_n850_), .Y(u1__0sram_addr_23_0__8_));
AND2X2 AND2X2_2526 ( .A(u1__abc_73140_new_n854_), .B(u1__abc_73140_new_n853_), .Y(u1__0sram_addr_23_0__9_));
AND2X2 AND2X2_2527 ( .A(u1__abc_73140_new_n857_), .B(u1__abc_73140_new_n856_), .Y(u1__0sram_addr_23_0__10_));
AND2X2 AND2X2_2528 ( .A(u1__abc_73140_new_n860_), .B(u1__abc_73140_new_n859_), .Y(u1__0sram_addr_23_0__11_));
AND2X2 AND2X2_2529 ( .A(u1__abc_73140_new_n863_), .B(u1__abc_73140_new_n862_), .Y(u1__0sram_addr_23_0__12_));
AND2X2 AND2X2_253 ( .A(u0__abc_76628_new_n1170__bF_buf2), .B(sp_tms_11_), .Y(u0__abc_76628_new_n1442_));
AND2X2 AND2X2_2530 ( .A(u1__abc_73140_new_n866_), .B(u1__abc_73140_new_n865_), .Y(u1__0sram_addr_23_0__13_));
AND2X2 AND2X2_2531 ( .A(u1__abc_73140_new_n869_), .B(u1__abc_73140_new_n868_), .Y(u1__0sram_addr_23_0__14_));
AND2X2 AND2X2_2532 ( .A(u1__abc_73140_new_n872_), .B(u1__abc_73140_new_n871_), .Y(u1__0sram_addr_23_0__15_));
AND2X2 AND2X2_2533 ( .A(u1__abc_73140_new_n875_), .B(u1__abc_73140_new_n874_), .Y(u1__0sram_addr_23_0__16_));
AND2X2 AND2X2_2534 ( .A(u1__abc_73140_new_n878_), .B(u1__abc_73140_new_n877_), .Y(u1__0sram_addr_23_0__17_));
AND2X2 AND2X2_2535 ( .A(u1__abc_73140_new_n881_), .B(u1__abc_73140_new_n880_), .Y(u1__0sram_addr_23_0__18_));
AND2X2 AND2X2_2536 ( .A(u1__abc_73140_new_n884_), .B(u1__abc_73140_new_n883_), .Y(u1__0sram_addr_23_0__19_));
AND2X2 AND2X2_2537 ( .A(u1__abc_73140_new_n887_), .B(u1__abc_73140_new_n886_), .Y(u1__0sram_addr_23_0__20_));
AND2X2 AND2X2_2538 ( .A(u1__abc_73140_new_n890_), .B(u1__abc_73140_new_n889_), .Y(u1__0sram_addr_23_0__21_));
AND2X2 AND2X2_2539 ( .A(u1__abc_73140_new_n893_), .B(u1__abc_73140_new_n892_), .Y(u1__0sram_addr_23_0__22_));
AND2X2 AND2X2_254 ( .A(spec_req_cs_5_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1443_));
AND2X2 AND2X2_2540 ( .A(u1__abc_73140_new_n896_), .B(u1__abc_73140_new_n895_), .Y(u1__0sram_addr_23_0__23_));
AND2X2 AND2X2_2541 ( .A(u1__abc_73140_new_n899_), .B(csc_s_2_), .Y(u1__abc_73140_new_n900_));
AND2X2 AND2X2_2542 ( .A(csc_s_1_), .B(u1_wr_hold), .Y(u1__abc_73140_new_n903_));
AND2X2 AND2X2_2543 ( .A(u1__abc_73140_new_n902_), .B(u1__abc_73140_new_n903_), .Y(u1__abc_73140_new_n904_));
AND2X2 AND2X2_2544 ( .A(u1__abc_73140_new_n907_), .B(u1__abc_73140_new_n905_), .Y(u1__abc_73140_new_n908_));
AND2X2 AND2X2_2545 ( .A(u1__abc_73140_new_n899_), .B(u1__abc_73140_new_n910_), .Y(u1__abc_73140_new_n911_));
AND2X2 AND2X2_2546 ( .A(u1__abc_73140_new_n914_), .B(u1__abc_73140_new_n912__bF_buf3), .Y(u1__abc_73140_new_n915_));
AND2X2 AND2X2_2547 ( .A(u1__abc_73140_new_n909_), .B(u1__abc_73140_new_n915_), .Y(u1__abc_73140_new_n916_));
AND2X2 AND2X2_2548 ( .A(u1__abc_73140_new_n917_), .B(lmr_sel_bF_buf3), .Y(u1__abc_73140_new_n918_));
AND2X2 AND2X2_2549 ( .A(u1__abc_73140_new_n922_), .B(u1__abc_73140_new_n923_), .Y(u1__abc_73140_new_n924_));
AND2X2 AND2X2_255 ( .A(u0__abc_76628_new_n1445_), .B(u0__abc_76628_new_n1179__bF_buf0), .Y(u0__abc_76628_new_n1446_));
AND2X2 AND2X2_2550 ( .A(u1__abc_73140_new_n925_), .B(u1__abc_73140_new_n920_), .Y(u1__abc_73140_new_n926_));
AND2X2 AND2X2_2551 ( .A(u1__abc_73140_new_n926_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n927_));
AND2X2 AND2X2_2552 ( .A(u1__abc_73140_new_n930_), .B(u1__abc_73140_new_n929_), .Y(u1__abc_73140_new_n931_));
AND2X2 AND2X2_2553 ( .A(u1__abc_73140_new_n933_), .B(u1__abc_73140_new_n912__bF_buf2), .Y(u1__abc_73140_new_n934_));
AND2X2 AND2X2_2554 ( .A(u1__abc_73140_new_n932_), .B(u1__abc_73140_new_n934_), .Y(u1__abc_73140_new_n935_));
AND2X2 AND2X2_2555 ( .A(u1__abc_73140_new_n937_), .B(u1__abc_73140_new_n938_), .Y(u1__abc_73140_new_n939_));
AND2X2 AND2X2_2556 ( .A(u1__abc_73140_new_n940_), .B(u1__abc_73140_new_n936_), .Y(u1__abc_73140_new_n941_));
AND2X2 AND2X2_2557 ( .A(u1__abc_73140_new_n941_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n942_));
AND2X2 AND2X2_2558 ( .A(u1__abc_73140_new_n945_), .B(u1__abc_73140_new_n944_), .Y(u1__abc_73140_new_n946_));
AND2X2 AND2X2_2559 ( .A(u1__abc_73140_new_n948_), .B(u1__abc_73140_new_n912__bF_buf1), .Y(u1__abc_73140_new_n949_));
AND2X2 AND2X2_256 ( .A(u0__abc_76628_new_n1446_), .B(u0__abc_76628_new_n1444_), .Y(u0__abc_76628_new_n1447_));
AND2X2 AND2X2_2560 ( .A(u1__abc_73140_new_n947_), .B(u1__abc_73140_new_n949_), .Y(u1__abc_73140_new_n950_));
AND2X2 AND2X2_2561 ( .A(u1__abc_73140_new_n952_), .B(u1__abc_73140_new_n953_), .Y(u1__abc_73140_new_n954_));
AND2X2 AND2X2_2562 ( .A(u1__abc_73140_new_n955_), .B(u1__abc_73140_new_n951_), .Y(u1__abc_73140_new_n956_));
AND2X2 AND2X2_2563 ( .A(u1__abc_73140_new_n956_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n957_));
AND2X2 AND2X2_2564 ( .A(u1__abc_73140_new_n960_), .B(u1__abc_73140_new_n959_), .Y(u1__abc_73140_new_n961_));
AND2X2 AND2X2_2565 ( .A(u1__abc_73140_new_n963_), .B(u1__abc_73140_new_n912__bF_buf0), .Y(u1__abc_73140_new_n964_));
AND2X2 AND2X2_2566 ( .A(u1__abc_73140_new_n962_), .B(u1__abc_73140_new_n964_), .Y(u1__abc_73140_new_n965_));
AND2X2 AND2X2_2567 ( .A(u1__abc_73140_new_n967_), .B(u1__abc_73140_new_n968_), .Y(u1__abc_73140_new_n969_));
AND2X2 AND2X2_2568 ( .A(u1__abc_73140_new_n970_), .B(u1__abc_73140_new_n966_), .Y(u1__abc_73140_new_n971_));
AND2X2 AND2X2_2569 ( .A(u1__abc_73140_new_n971_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n972_));
AND2X2 AND2X2_257 ( .A(u0__abc_76628_new_n1448_), .B(u0__abc_76628_new_n1175__bF_buf0), .Y(u0__abc_76628_new_n1449_));
AND2X2 AND2X2_2570 ( .A(u1__abc_73140_new_n975_), .B(u1__abc_73140_new_n974_), .Y(u1__abc_73140_new_n976_));
AND2X2 AND2X2_2571 ( .A(u1__abc_73140_new_n978_), .B(u1__abc_73140_new_n912__bF_buf3), .Y(u1__abc_73140_new_n979_));
AND2X2 AND2X2_2572 ( .A(u1__abc_73140_new_n977_), .B(u1__abc_73140_new_n979_), .Y(u1__abc_73140_new_n980_));
AND2X2 AND2X2_2573 ( .A(u1__abc_73140_new_n982_), .B(u1__abc_73140_new_n983_), .Y(u1__abc_73140_new_n984_));
AND2X2 AND2X2_2574 ( .A(u1__abc_73140_new_n985_), .B(u1__abc_73140_new_n981_), .Y(u1__abc_73140_new_n986_));
AND2X2 AND2X2_2575 ( .A(u1__abc_73140_new_n986_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n987_));
AND2X2 AND2X2_2576 ( .A(u1__abc_73140_new_n990_), .B(u1__abc_73140_new_n989_), .Y(u1__abc_73140_new_n991_));
AND2X2 AND2X2_2577 ( .A(u1__abc_73140_new_n993_), .B(u1__abc_73140_new_n912__bF_buf2), .Y(u1__abc_73140_new_n994_));
AND2X2 AND2X2_2578 ( .A(u1__abc_73140_new_n992_), .B(u1__abc_73140_new_n994_), .Y(u1__abc_73140_new_n995_));
AND2X2 AND2X2_2579 ( .A(u1__abc_73140_new_n997_), .B(u1__abc_73140_new_n998_), .Y(u1__abc_73140_new_n999_));
AND2X2 AND2X2_258 ( .A(spec_req_cs_4_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1450_));
AND2X2 AND2X2_2580 ( .A(u1__abc_73140_new_n1000_), .B(u1__abc_73140_new_n996_), .Y(u1__abc_73140_new_n1001_));
AND2X2 AND2X2_2581 ( .A(u1__abc_73140_new_n1001_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n1002_));
AND2X2 AND2X2_2582 ( .A(u1__abc_73140_new_n1005_), .B(u1__abc_73140_new_n1004_), .Y(u1__abc_73140_new_n1006_));
AND2X2 AND2X2_2583 ( .A(u1__abc_73140_new_n1008_), .B(u1__abc_73140_new_n912__bF_buf1), .Y(u1__abc_73140_new_n1009_));
AND2X2 AND2X2_2584 ( .A(u1__abc_73140_new_n1007_), .B(u1__abc_73140_new_n1009_), .Y(u1__abc_73140_new_n1010_));
AND2X2 AND2X2_2585 ( .A(u1__abc_73140_new_n1012_), .B(u1__abc_73140_new_n1013_), .Y(u1__abc_73140_new_n1014_));
AND2X2 AND2X2_2586 ( .A(u1__abc_73140_new_n1015_), .B(u1__abc_73140_new_n1011_), .Y(u1__abc_73140_new_n1016_));
AND2X2 AND2X2_2587 ( .A(u1__abc_73140_new_n1016_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n1017_));
AND2X2 AND2X2_2588 ( .A(u1__abc_73140_new_n1020_), .B(u1__abc_73140_new_n1019_), .Y(u1__abc_73140_new_n1021_));
AND2X2 AND2X2_2589 ( .A(u1__abc_73140_new_n1023_), .B(u1__abc_73140_new_n912__bF_buf0), .Y(u1__abc_73140_new_n1024_));
AND2X2 AND2X2_259 ( .A(u0__abc_76628_new_n1451_), .B(u0__abc_76628_new_n1174__bF_buf0), .Y(u0__abc_76628_new_n1452_));
AND2X2 AND2X2_2590 ( .A(u1__abc_73140_new_n1022_), .B(u1__abc_73140_new_n1024_), .Y(u1__abc_73140_new_n1025_));
AND2X2 AND2X2_2591 ( .A(u1__abc_73140_new_n1027_), .B(u1__abc_73140_new_n1028_), .Y(u1__abc_73140_new_n1029_));
AND2X2 AND2X2_2592 ( .A(u1__abc_73140_new_n1030_), .B(u1__abc_73140_new_n1026_), .Y(u1__abc_73140_new_n1031_));
AND2X2 AND2X2_2593 ( .A(u1__abc_73140_new_n1031_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n1032_));
AND2X2 AND2X2_2594 ( .A(u1__abc_73140_new_n1035_), .B(u1__abc_73140_new_n1034_), .Y(u1__abc_73140_new_n1036_));
AND2X2 AND2X2_2595 ( .A(u1__abc_73140_new_n1038_), .B(u1__abc_73140_new_n912__bF_buf3), .Y(u1__abc_73140_new_n1039_));
AND2X2 AND2X2_2596 ( .A(u1__abc_73140_new_n1037_), .B(u1__abc_73140_new_n1039_), .Y(u1__abc_73140_new_n1040_));
AND2X2 AND2X2_2597 ( .A(u1__abc_73140_new_n1042_), .B(u1__abc_73140_new_n1043_), .Y(u1__abc_73140_new_n1044_));
AND2X2 AND2X2_2598 ( .A(u1__abc_73140_new_n1045_), .B(u1__abc_73140_new_n1041_), .Y(u1__abc_73140_new_n1046_));
AND2X2 AND2X2_2599 ( .A(u1__abc_73140_new_n1046_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n1047_));
AND2X2 AND2X2_26 ( .A(_abc_85006_new_n314_), .B(_abc_85006_new_n315_), .Y(tms_s_8_));
AND2X2 AND2X2_260 ( .A(spec_req_cs_3_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1453_));
AND2X2 AND2X2_2600 ( .A(u1__abc_73140_new_n1050_), .B(u1__abc_73140_new_n1049_), .Y(u1__abc_73140_new_n1051_));
AND2X2 AND2X2_2601 ( .A(u1__abc_73140_new_n1053_), .B(u1__abc_73140_new_n912__bF_buf2), .Y(u1__abc_73140_new_n1054_));
AND2X2 AND2X2_2602 ( .A(u1__abc_73140_new_n1052_), .B(u1__abc_73140_new_n1054_), .Y(u1__abc_73140_new_n1055_));
AND2X2 AND2X2_2603 ( .A(u1__abc_73140_new_n1057_), .B(u1__abc_73140_new_n1058_), .Y(u1__abc_73140_new_n1059_));
AND2X2 AND2X2_2604 ( .A(u1__abc_73140_new_n1060_), .B(u1__abc_73140_new_n1056_), .Y(u1__abc_73140_new_n1061_));
AND2X2 AND2X2_2605 ( .A(u1__abc_73140_new_n1061_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n1062_));
AND2X2 AND2X2_2606 ( .A(u1__abc_73140_new_n1065_), .B(u1__abc_73140_new_n1064_), .Y(u1__abc_73140_new_n1066_));
AND2X2 AND2X2_2607 ( .A(u1__abc_73140_new_n1068_), .B(u1__abc_73140_new_n912__bF_buf1), .Y(u1__abc_73140_new_n1069_));
AND2X2 AND2X2_2608 ( .A(u1__abc_73140_new_n1067_), .B(u1__abc_73140_new_n1069_), .Y(u1__abc_73140_new_n1070_));
AND2X2 AND2X2_2609 ( .A(row_adr_11_bF_buf2_), .B(row_sel), .Y(u1__abc_73140_new_n1072_));
AND2X2 AND2X2_261 ( .A(u0__abc_76628_new_n1454_), .B(u0__abc_76628_new_n1173__bF_buf0), .Y(u0__abc_76628_new_n1455_));
AND2X2 AND2X2_2610 ( .A(u1__abc_73140_new_n911_), .B(u1__abc_73140_new_n1073_), .Y(u1__abc_73140_new_n1074_));
AND2X2 AND2X2_2611 ( .A(u1__abc_73140_new_n1074_), .B(u1__abc_73140_new_n1071_), .Y(u1__abc_73140_new_n1075_));
AND2X2 AND2X2_2612 ( .A(u1__abc_73140_new_n1078_), .B(u1__abc_73140_new_n1077_), .Y(u1__abc_73140_new_n1079_));
AND2X2 AND2X2_2613 ( .A(u1__abc_73140_new_n1081_), .B(u1__abc_73140_new_n912__bF_buf0), .Y(u1__abc_73140_new_n1082_));
AND2X2 AND2X2_2614 ( .A(u1__abc_73140_new_n1080_), .B(u1__abc_73140_new_n1082_), .Y(u1__abc_73140_new_n1083_));
AND2X2 AND2X2_2615 ( .A(row_adr_12_bF_buf2_), .B(row_sel), .Y(u1__abc_73140_new_n1085_));
AND2X2 AND2X2_2616 ( .A(u1__abc_73140_new_n911_), .B(u1__abc_73140_new_n1086_), .Y(u1__abc_73140_new_n1087_));
AND2X2 AND2X2_2617 ( .A(u1__abc_73140_new_n1087_), .B(u1__abc_73140_new_n1084_), .Y(u1__abc_73140_new_n1088_));
AND2X2 AND2X2_2618 ( .A(u1__abc_73140_new_n1091_), .B(u1__abc_73140_new_n1090_), .Y(u1__abc_73140_new_n1092_));
AND2X2 AND2X2_2619 ( .A(u1__abc_73140_new_n1094_), .B(u1__abc_73140_new_n912__bF_buf3), .Y(u1__abc_73140_new_n1095_));
AND2X2 AND2X2_262 ( .A(spec_req_cs_2_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1456_));
AND2X2 AND2X2_2620 ( .A(u1__abc_73140_new_n1093_), .B(u1__abc_73140_new_n1095_), .Y(u1__abc_73140_new_n1096_));
AND2X2 AND2X2_2621 ( .A(u1__abc_73140_new_n911_), .B(bank_adr_0_), .Y(u1__abc_73140_new_n1097_));
AND2X2 AND2X2_2622 ( .A(u1__abc_73140_new_n1100_), .B(u1__abc_73140_new_n1099_), .Y(u1__abc_73140_new_n1101_));
AND2X2 AND2X2_2623 ( .A(u1__abc_73140_new_n1103_), .B(u1__abc_73140_new_n912__bF_buf2), .Y(u1__abc_73140_new_n1104_));
AND2X2 AND2X2_2624 ( .A(u1__abc_73140_new_n1102_), .B(u1__abc_73140_new_n1104_), .Y(u1__abc_73140_new_n1105_));
AND2X2 AND2X2_2625 ( .A(u1__abc_73140_new_n911_), .B(bank_adr_1_), .Y(u1__abc_73140_new_n1106_));
AND2X2 AND2X2_2626 ( .A(u1__abc_73140_new_n906__bF_buf1), .B(\wb_addr_i[17] ), .Y(u1__abc_73140_new_n1108_));
AND2X2 AND2X2_2627 ( .A(u1__abc_73140_new_n904__bF_buf4), .B(u1_sram_addr_15_), .Y(u1__abc_73140_new_n1109_));
AND2X2 AND2X2_2628 ( .A(u1__abc_73140_new_n912__bF_buf1), .B(u1__abc_73140_new_n1112_), .Y(u1__abc_73140_new_n1113_));
AND2X2 AND2X2_2629 ( .A(u1__abc_73140_new_n1111_), .B(u1__abc_73140_new_n1113_), .Y(mc_addr_d_15_));
AND2X2 AND2X2_263 ( .A(u0__abc_76628_new_n1457_), .B(u0__abc_76628_new_n1172__bF_buf0), .Y(u0__abc_76628_new_n1458_));
AND2X2 AND2X2_2630 ( .A(u1__abc_73140_new_n906__bF_buf0), .B(\wb_addr_i[18] ), .Y(u1__abc_73140_new_n1115_));
AND2X2 AND2X2_2631 ( .A(u1__abc_73140_new_n904__bF_buf3), .B(u1_sram_addr_16_), .Y(u1__abc_73140_new_n1116_));
AND2X2 AND2X2_2632 ( .A(u1__abc_73140_new_n912__bF_buf0), .B(u1__abc_73140_new_n1119_), .Y(u1__abc_73140_new_n1120_));
AND2X2 AND2X2_2633 ( .A(u1__abc_73140_new_n1118_), .B(u1__abc_73140_new_n1120_), .Y(mc_addr_d_16_));
AND2X2 AND2X2_2634 ( .A(u1__abc_73140_new_n906__bF_buf3), .B(\wb_addr_i[19] ), .Y(u1__abc_73140_new_n1122_));
AND2X2 AND2X2_2635 ( .A(u1__abc_73140_new_n904__bF_buf2), .B(u1_sram_addr_17_), .Y(u1__abc_73140_new_n1123_));
AND2X2 AND2X2_2636 ( .A(u1__abc_73140_new_n912__bF_buf3), .B(u1__abc_73140_new_n1126_), .Y(u1__abc_73140_new_n1127_));
AND2X2 AND2X2_2637 ( .A(u1__abc_73140_new_n1125_), .B(u1__abc_73140_new_n1127_), .Y(mc_addr_d_17_));
AND2X2 AND2X2_2638 ( .A(u1__abc_73140_new_n906__bF_buf2), .B(\wb_addr_i[20] ), .Y(u1__abc_73140_new_n1129_));
AND2X2 AND2X2_2639 ( .A(u1__abc_73140_new_n904__bF_buf1), .B(u1_sram_addr_18_), .Y(u1__abc_73140_new_n1130_));
AND2X2 AND2X2_264 ( .A(spec_req_cs_1_bF_buf3_), .B(u0_tms1_11_), .Y(u0__abc_76628_new_n1459_));
AND2X2 AND2X2_2640 ( .A(u1__abc_73140_new_n912__bF_buf2), .B(u1__abc_73140_new_n1133_), .Y(u1__abc_73140_new_n1134_));
AND2X2 AND2X2_2641 ( .A(u1__abc_73140_new_n1132_), .B(u1__abc_73140_new_n1134_), .Y(mc_addr_d_18_));
AND2X2 AND2X2_2642 ( .A(u1__abc_73140_new_n906__bF_buf1), .B(\wb_addr_i[21] ), .Y(u1__abc_73140_new_n1136_));
AND2X2 AND2X2_2643 ( .A(u1__abc_73140_new_n904__bF_buf0), .B(u1_sram_addr_19_), .Y(u1__abc_73140_new_n1137_));
AND2X2 AND2X2_2644 ( .A(u1__abc_73140_new_n912__bF_buf1), .B(u1__abc_73140_new_n1140_), .Y(u1__abc_73140_new_n1141_));
AND2X2 AND2X2_2645 ( .A(u1__abc_73140_new_n1139_), .B(u1__abc_73140_new_n1141_), .Y(mc_addr_d_19_));
AND2X2 AND2X2_2646 ( .A(u1__abc_73140_new_n906__bF_buf0), .B(\wb_addr_i[22] ), .Y(u1__abc_73140_new_n1143_));
AND2X2 AND2X2_2647 ( .A(u1__abc_73140_new_n904__bF_buf4), .B(u1_sram_addr_20_), .Y(u1__abc_73140_new_n1144_));
AND2X2 AND2X2_2648 ( .A(u1__abc_73140_new_n912__bF_buf0), .B(u1__abc_73140_new_n1147_), .Y(u1__abc_73140_new_n1148_));
AND2X2 AND2X2_2649 ( .A(u1__abc_73140_new_n1146_), .B(u1__abc_73140_new_n1148_), .Y(mc_addr_d_20_));
AND2X2 AND2X2_265 ( .A(u0__abc_76628_new_n1169__bF_buf1), .B(u0__abc_76628_new_n1462_), .Y(u0__abc_76628_new_n1463_));
AND2X2 AND2X2_2650 ( .A(u1__abc_73140_new_n906__bF_buf3), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n1150_));
AND2X2 AND2X2_2651 ( .A(u1__abc_73140_new_n904__bF_buf3), .B(u1_sram_addr_21_), .Y(u1__abc_73140_new_n1151_));
AND2X2 AND2X2_2652 ( .A(u1__abc_73140_new_n912__bF_buf3), .B(u1__abc_73140_new_n1154_), .Y(u1__abc_73140_new_n1155_));
AND2X2 AND2X2_2653 ( .A(u1__abc_73140_new_n1153_), .B(u1__abc_73140_new_n1155_), .Y(mc_addr_d_21_));
AND2X2 AND2X2_2654 ( .A(u1__abc_73140_new_n906__bF_buf2), .B(\wb_addr_i[24] ), .Y(u1__abc_73140_new_n1157_));
AND2X2 AND2X2_2655 ( .A(u1__abc_73140_new_n904__bF_buf2), .B(u1_sram_addr_22_), .Y(u1__abc_73140_new_n1158_));
AND2X2 AND2X2_2656 ( .A(u1__abc_73140_new_n912__bF_buf2), .B(u1__abc_73140_new_n1161_), .Y(u1__abc_73140_new_n1162_));
AND2X2 AND2X2_2657 ( .A(u1__abc_73140_new_n1160_), .B(u1__abc_73140_new_n1162_), .Y(mc_addr_d_22_));
AND2X2 AND2X2_2658 ( .A(u1__abc_73140_new_n904__bF_buf1), .B(u1_sram_addr_23_), .Y(u1__abc_73140_new_n1164_));
AND2X2 AND2X2_2659 ( .A(u1__abc_73140_new_n906__bF_buf1), .B(\wb_addr_i[25] ), .Y(u1__abc_73140_new_n1165_));
AND2X2 AND2X2_266 ( .A(u0__abc_76628_new_n1461_), .B(u0__abc_76628_new_n1463_), .Y(u0__abc_76628_new_n1464_));
AND2X2 AND2X2_2660 ( .A(u1__abc_73140_new_n912__bF_buf1), .B(u1__abc_73140_new_n1168_), .Y(u1__abc_73140_new_n1169_));
AND2X2 AND2X2_2661 ( .A(u1__abc_73140_new_n1167_), .B(u1__abc_73140_new_n1169_), .Y(mc_addr_d_23_));
AND2X2 AND2X2_2662 ( .A(u1__abc_73140_new_n1171_), .B(u1__abc_73140_new_n1172_), .Y(u1__abc_73140_new_n1173_));
AND2X2 AND2X2_2663 ( .A(u1__abc_73140_new_n912__bF_buf0), .B(u1__abc_73140_new_n1175_), .Y(u1__abc_73140_new_n1176_));
AND2X2 AND2X2_2664 ( .A(u1__abc_73140_new_n1174_), .B(u1__abc_73140_new_n1176_), .Y(u1__abc_73140_new_n1177_));
AND2X2 AND2X2_2665 ( .A(u1__abc_73140_new_n1178_), .B(u1__abc_73140_new_n1179_), .Y(u1__abc_73140_new_n1180_));
AND2X2 AND2X2_2666 ( .A(u1__abc_73140_new_n1182_), .B(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n1183_));
AND2X2 AND2X2_2667 ( .A(u1__abc_73140_new_n1183_), .B(u1__abc_73140_new_n1181_), .Y(u1__abc_73140_new_n1184_));
AND2X2 AND2X2_2668 ( .A(u1_acs_addr_0_), .B(u1_acs_addr_1_), .Y(u1_u0__abc_73035_new_n51_));
AND2X2 AND2X2_2669 ( .A(u1_u0__abc_73035_new_n52_), .B(u1_u0__abc_73035_new_n53_), .Y(u1_u0__0out_r_12_0__1_));
AND2X2 AND2X2_267 ( .A(u0__abc_76628_new_n1170__bF_buf1), .B(sp_tms_12_), .Y(u0__abc_76628_new_n1466_));
AND2X2 AND2X2_2670 ( .A(u1_u0__abc_73035_new_n51_), .B(u1_acs_addr_2_), .Y(u1_u0__abc_73035_new_n55_));
AND2X2 AND2X2_2671 ( .A(u1_u0__abc_73035_new_n56_), .B(u1_u0__abc_73035_new_n57_), .Y(u1_u0__0out_r_12_0__2_));
AND2X2 AND2X2_2672 ( .A(u1_u0__abc_73035_new_n55_), .B(u1_acs_addr_3_), .Y(u1_u0__abc_73035_new_n59_));
AND2X2 AND2X2_2673 ( .A(u1_u0__abc_73035_new_n60_), .B(u1_u0__abc_73035_new_n61_), .Y(u1_u0__0out_r_12_0__3_));
AND2X2 AND2X2_2674 ( .A(u1_u0__abc_73035_new_n59_), .B(u1_acs_addr_4_), .Y(u1_u0__abc_73035_new_n63_));
AND2X2 AND2X2_2675 ( .A(u1_u0__abc_73035_new_n64_), .B(u1_u0__abc_73035_new_n65_), .Y(u1_u0__0out_r_12_0__4_));
AND2X2 AND2X2_2676 ( .A(u1_acs_addr_4_), .B(u1_acs_addr_5_), .Y(u1_u0__abc_73035_new_n68_));
AND2X2 AND2X2_2677 ( .A(u1_u0__abc_73035_new_n59_), .B(u1_u0__abc_73035_new_n68_), .Y(u1_u0__abc_73035_new_n69_));
AND2X2 AND2X2_2678 ( .A(u1_u0__abc_73035_new_n67_), .B(u1_u0__abc_73035_new_n70_), .Y(u1_u0__0out_r_12_0__5_));
AND2X2 AND2X2_2679 ( .A(u1_u0__abc_73035_new_n69_), .B(u1_acs_addr_6_), .Y(u1_u0__abc_73035_new_n72_));
AND2X2 AND2X2_268 ( .A(spec_req_cs_5_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1467_));
AND2X2 AND2X2_2680 ( .A(u1_u0__abc_73035_new_n73_), .B(u1_u0__abc_73035_new_n74_), .Y(u1_u0__0out_r_12_0__6_));
AND2X2 AND2X2_2681 ( .A(u1_acs_addr_6_), .B(u1_acs_addr_7_), .Y(u1_u0__abc_73035_new_n77_));
AND2X2 AND2X2_2682 ( .A(u1_u0__abc_73035_new_n68_), .B(u1_u0__abc_73035_new_n77_), .Y(u1_u0__abc_73035_new_n78_));
AND2X2 AND2X2_2683 ( .A(u1_u0__abc_73035_new_n59_), .B(u1_u0__abc_73035_new_n78_), .Y(u1_u0__abc_73035_new_n79_));
AND2X2 AND2X2_2684 ( .A(u1_u0__abc_73035_new_n76_), .B(u1_u0__abc_73035_new_n80_), .Y(u1_u0__0out_r_12_0__7_));
AND2X2 AND2X2_2685 ( .A(u1_u0__abc_73035_new_n79_), .B(u1_acs_addr_8_), .Y(u1_u0__abc_73035_new_n82_));
AND2X2 AND2X2_2686 ( .A(u1_u0__abc_73035_new_n83_), .B(u1_u0__abc_73035_new_n84_), .Y(u1_u0__0out_r_12_0__8_));
AND2X2 AND2X2_2687 ( .A(u1_acs_addr_8_), .B(u1_acs_addr_9_), .Y(u1_u0__abc_73035_new_n87_));
AND2X2 AND2X2_2688 ( .A(u1_u0__abc_73035_new_n79_), .B(u1_u0__abc_73035_new_n87_), .Y(u1_u0__abc_73035_new_n88_));
AND2X2 AND2X2_2689 ( .A(u1_u0__abc_73035_new_n86_), .B(u1_u0__abc_73035_new_n89_), .Y(u1_u0__0out_r_12_0__9_));
AND2X2 AND2X2_269 ( .A(u0__abc_76628_new_n1469_), .B(u0__abc_76628_new_n1179__bF_buf5), .Y(u0__abc_76628_new_n1470_));
AND2X2 AND2X2_2690 ( .A(u1_u0__abc_73035_new_n88_), .B(u1_acs_addr_10_), .Y(u1_u0__abc_73035_new_n91_));
AND2X2 AND2X2_2691 ( .A(u1_u0__abc_73035_new_n92_), .B(u1_u0__abc_73035_new_n93_), .Y(u1_u0__0out_r_12_0__10_));
AND2X2 AND2X2_2692 ( .A(u1_acs_addr_10_), .B(u1_acs_addr_11_), .Y(u1_u0__abc_73035_new_n95_));
AND2X2 AND2X2_2693 ( .A(u1_u0__abc_73035_new_n87_), .B(u1_u0__abc_73035_new_n95_), .Y(u1_u0__abc_73035_new_n96_));
AND2X2 AND2X2_2694 ( .A(u1_u0__abc_73035_new_n79_), .B(u1_u0__abc_73035_new_n96_), .Y(u1_u0__0out_r_12_0__12_));
AND2X2 AND2X2_2695 ( .A(u1_u0__abc_73035_new_n99_), .B(u1_u0__abc_73035_new_n98_), .Y(u1_u0__0out_r_12_0__11_));
AND2X2 AND2X2_2696 ( .A(u1_u0_inc_next), .B(u1_acs_addr_12_), .Y(u1_u0__abc_73035_new_n102_));
AND2X2 AND2X2_2697 ( .A(u1_u0__abc_73035_new_n102_), .B(u1_acs_addr_13_), .Y(u1_u0__abc_73035_new_n103_));
AND2X2 AND2X2_2698 ( .A(u1_u0__abc_73035_new_n104_), .B(u1_u0__abc_73035_new_n105_), .Y(u1_acs_addr_pl1_13_));
AND2X2 AND2X2_2699 ( .A(u1_u0__abc_73035_new_n103_), .B(u1_acs_addr_14_), .Y(u1_u0__abc_73035_new_n107_));
AND2X2 AND2X2_27 ( .A(_abc_85006_new_n317_), .B(_abc_85006_new_n318_), .Y(tms_s_9_));
AND2X2 AND2X2_270 ( .A(u0__abc_76628_new_n1470_), .B(u0__abc_76628_new_n1468_), .Y(u0__abc_76628_new_n1471_));
AND2X2 AND2X2_2700 ( .A(u1_u0__abc_73035_new_n108_), .B(u1_u0__abc_73035_new_n109_), .Y(u1_acs_addr_pl1_14_));
AND2X2 AND2X2_2701 ( .A(u1_acs_addr_14_), .B(u1_acs_addr_15_), .Y(u1_u0__abc_73035_new_n112_));
AND2X2 AND2X2_2702 ( .A(u1_u0__abc_73035_new_n103_), .B(u1_u0__abc_73035_new_n112_), .Y(u1_u0__abc_73035_new_n113_));
AND2X2 AND2X2_2703 ( .A(u1_u0__abc_73035_new_n111_), .B(u1_u0__abc_73035_new_n114_), .Y(u1_acs_addr_pl1_15_));
AND2X2 AND2X2_2704 ( .A(u1_u0__abc_73035_new_n113_), .B(u1_acs_addr_16_), .Y(u1_u0__abc_73035_new_n116_));
AND2X2 AND2X2_2705 ( .A(u1_u0__abc_73035_new_n117_), .B(u1_u0__abc_73035_new_n118_), .Y(u1_acs_addr_pl1_16_));
AND2X2 AND2X2_2706 ( .A(u1_acs_addr_16_), .B(u1_acs_addr_17_), .Y(u1_u0__abc_73035_new_n121_));
AND2X2 AND2X2_2707 ( .A(u1_u0__abc_73035_new_n113_), .B(u1_u0__abc_73035_new_n121_), .Y(u1_u0__abc_73035_new_n122_));
AND2X2 AND2X2_2708 ( .A(u1_u0__abc_73035_new_n120_), .B(u1_u0__abc_73035_new_n123_), .Y(u1_acs_addr_pl1_17_));
AND2X2 AND2X2_2709 ( .A(u1_u0__abc_73035_new_n122_), .B(u1_acs_addr_18_), .Y(u1_u0__abc_73035_new_n125_));
AND2X2 AND2X2_271 ( .A(u0__abc_76628_new_n1472_), .B(u0__abc_76628_new_n1175__bF_buf5), .Y(u0__abc_76628_new_n1473_));
AND2X2 AND2X2_2710 ( .A(u1_u0__abc_73035_new_n126_), .B(u1_u0__abc_73035_new_n127_), .Y(u1_acs_addr_pl1_18_));
AND2X2 AND2X2_2711 ( .A(u1_acs_addr_18_), .B(u1_acs_addr_19_), .Y(u1_u0__abc_73035_new_n130_));
AND2X2 AND2X2_2712 ( .A(u1_u0__abc_73035_new_n121_), .B(u1_u0__abc_73035_new_n130_), .Y(u1_u0__abc_73035_new_n131_));
AND2X2 AND2X2_2713 ( .A(u1_u0__abc_73035_new_n113_), .B(u1_u0__abc_73035_new_n131_), .Y(u1_u0__abc_73035_new_n132_));
AND2X2 AND2X2_2714 ( .A(u1_u0__abc_73035_new_n129_), .B(u1_u0__abc_73035_new_n133_), .Y(u1_acs_addr_pl1_19_));
AND2X2 AND2X2_2715 ( .A(u1_u0__abc_73035_new_n132_), .B(u1_acs_addr_20_), .Y(u1_u0__abc_73035_new_n135_));
AND2X2 AND2X2_2716 ( .A(u1_u0__abc_73035_new_n136_), .B(u1_u0__abc_73035_new_n137_), .Y(u1_acs_addr_pl1_20_));
AND2X2 AND2X2_2717 ( .A(u1_acs_addr_20_), .B(u1_acs_addr_21_), .Y(u1_u0__abc_73035_new_n140_));
AND2X2 AND2X2_2718 ( .A(u1_u0__abc_73035_new_n132_), .B(u1_u0__abc_73035_new_n140_), .Y(u1_u0__abc_73035_new_n141_));
AND2X2 AND2X2_2719 ( .A(u1_u0__abc_73035_new_n139_), .B(u1_u0__abc_73035_new_n142_), .Y(u1_acs_addr_pl1_21_));
AND2X2 AND2X2_272 ( .A(spec_req_cs_4_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1474_));
AND2X2 AND2X2_2720 ( .A(u1_u0__abc_73035_new_n141_), .B(u1_acs_addr_22_), .Y(u1_u0__abc_73035_new_n144_));
AND2X2 AND2X2_2721 ( .A(u1_u0__abc_73035_new_n145_), .B(u1_u0__abc_73035_new_n146_), .Y(u1_acs_addr_pl1_22_));
AND2X2 AND2X2_2722 ( .A(u1_u0__abc_73035_new_n144_), .B(u1_acs_addr_23_), .Y(u1_u0__abc_73035_new_n149_));
AND2X2 AND2X2_2723 ( .A(u1_u0__abc_73035_new_n150_), .B(u1_u0__abc_73035_new_n148_), .Y(u1_acs_addr_pl1_23_));
AND2X2 AND2X2_2724 ( .A(u1_u0__abc_73035_new_n152_), .B(u1_u0__abc_73035_new_n153_), .Y(u1_acs_addr_pl1_12_));
AND2X2 AND2X2_2725 ( .A(bank_set), .B(obct_cs_0_), .Y(u2_bank_set_0));
AND2X2 AND2X2_2726 ( .A(bank_set), .B(obct_cs_1_), .Y(u2_bank_set_1));
AND2X2 AND2X2_2727 ( .A(obct_cs_0_), .B(bank_clr), .Y(u2_bank_clr_0));
AND2X2 AND2X2_2728 ( .A(obct_cs_1_), .B(bank_clr), .Y(u2_bank_clr_1));
AND2X2 AND2X2_2729 ( .A(obct_cs_0_), .B(bank_clr_all), .Y(u2__abc_75448_new_n80_));
AND2X2 AND2X2_273 ( .A(u0__abc_76628_new_n1475_), .B(u0__abc_76628_new_n1174__bF_buf5), .Y(u0__abc_76628_new_n1476_));
AND2X2 AND2X2_2730 ( .A(obct_cs_1_), .B(bank_clr_all), .Y(u2__abc_75448_new_n82_));
AND2X2 AND2X2_2731 ( .A(obct_cs_4_), .B(1'h0), .Y(u2__abc_75448_new_n96_));
AND2X2 AND2X2_2732 ( .A(obct_cs_2_), .B(1'h0), .Y(u2__abc_75448_new_n97_));
AND2X2 AND2X2_2733 ( .A(obct_cs_5_), .B(1'h0), .Y(u2__abc_75448_new_n99_));
AND2X2 AND2X2_2734 ( .A(obct_cs_3_), .B(1'h0), .Y(u2__abc_75448_new_n100_));
AND2X2 AND2X2_2735 ( .A(obct_cs_1_), .B(u2_bank_open_1), .Y(u2__abc_75448_new_n103_));
AND2X2 AND2X2_2736 ( .A(obct_cs_0_), .B(u2_bank_open_0), .Y(u2__abc_75448_new_n104_));
AND2X2 AND2X2_2737 ( .A(obct_cs_7_), .B(1'h0), .Y(u2__abc_75448_new_n106_));
AND2X2 AND2X2_2738 ( .A(obct_cs_6_), .B(1'h0), .Y(u2__abc_75448_new_n107_));
AND2X2 AND2X2_2739 ( .A(obct_cs_4_), .B(1'h0), .Y(u2__abc_75448_new_n111_));
AND2X2 AND2X2_274 ( .A(spec_req_cs_3_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1477_));
AND2X2 AND2X2_2740 ( .A(obct_cs_2_), .B(1'h0), .Y(u2__abc_75448_new_n112_));
AND2X2 AND2X2_2741 ( .A(obct_cs_5_), .B(1'h0), .Y(u2__abc_75448_new_n114_));
AND2X2 AND2X2_2742 ( .A(obct_cs_3_), .B(1'h0), .Y(u2__abc_75448_new_n115_));
AND2X2 AND2X2_2743 ( .A(obct_cs_1_), .B(u2_row_same_1), .Y(u2__abc_75448_new_n118_));
AND2X2 AND2X2_2744 ( .A(obct_cs_0_), .B(u2_row_same_0), .Y(u2__abc_75448_new_n119_));
AND2X2 AND2X2_2745 ( .A(obct_cs_7_), .B(1'h0), .Y(u2__abc_75448_new_n121_));
AND2X2 AND2X2_2746 ( .A(obct_cs_6_), .B(1'h0), .Y(u2__abc_75448_new_n122_));
AND2X2 AND2X2_2747 ( .A(bank_adr_0_), .B(bank_adr_1_), .Y(u2_u0__abc_74955_new_n136_));
AND2X2 AND2X2_2748 ( .A(u2_u0__abc_74955_new_n136_), .B(u2_bank_set_0), .Y(u2_u0__abc_74955_new_n137_));
AND2X2 AND2X2_2749 ( .A(u2_u0__abc_74955_new_n137__bF_buf3), .B(u2_u0__abc_74955_new_n139_), .Y(u2_u0__abc_74955_new_n140_));
AND2X2 AND2X2_275 ( .A(u0__abc_76628_new_n1478_), .B(u0__abc_76628_new_n1173__bF_buf5), .Y(u0__abc_76628_new_n1479_));
AND2X2 AND2X2_2750 ( .A(u2_u0__abc_74955_new_n141_), .B(u2_u0__abc_74955_new_n138_), .Y(u2_u0__0b3_last_row_12_0__0_));
AND2X2 AND2X2_2751 ( .A(u2_u0__abc_74955_new_n137__bF_buf1), .B(u2_u0__abc_74955_new_n144_), .Y(u2_u0__abc_74955_new_n145_));
AND2X2 AND2X2_2752 ( .A(u2_u0__abc_74955_new_n146_), .B(u2_u0__abc_74955_new_n143_), .Y(u2_u0__0b3_last_row_12_0__1_));
AND2X2 AND2X2_2753 ( .A(u2_u0__abc_74955_new_n137__bF_buf4), .B(u2_u0__abc_74955_new_n149_), .Y(u2_u0__abc_74955_new_n150_));
AND2X2 AND2X2_2754 ( .A(u2_u0__abc_74955_new_n151_), .B(u2_u0__abc_74955_new_n148_), .Y(u2_u0__0b3_last_row_12_0__2_));
AND2X2 AND2X2_2755 ( .A(u2_u0__abc_74955_new_n137__bF_buf2), .B(u2_u0__abc_74955_new_n154_), .Y(u2_u0__abc_74955_new_n155_));
AND2X2 AND2X2_2756 ( .A(u2_u0__abc_74955_new_n156_), .B(u2_u0__abc_74955_new_n153_), .Y(u2_u0__0b3_last_row_12_0__3_));
AND2X2 AND2X2_2757 ( .A(u2_u0__abc_74955_new_n137__bF_buf0), .B(u2_u0__abc_74955_new_n159_), .Y(u2_u0__abc_74955_new_n160_));
AND2X2 AND2X2_2758 ( .A(u2_u0__abc_74955_new_n161_), .B(u2_u0__abc_74955_new_n158_), .Y(u2_u0__0b3_last_row_12_0__4_));
AND2X2 AND2X2_2759 ( .A(u2_u0__abc_74955_new_n137__bF_buf3), .B(u2_u0__abc_74955_new_n164_), .Y(u2_u0__abc_74955_new_n165_));
AND2X2 AND2X2_276 ( .A(spec_req_cs_2_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1480_));
AND2X2 AND2X2_2760 ( .A(u2_u0__abc_74955_new_n166_), .B(u2_u0__abc_74955_new_n163_), .Y(u2_u0__0b3_last_row_12_0__5_));
AND2X2 AND2X2_2761 ( .A(u2_u0__abc_74955_new_n137__bF_buf1), .B(u2_u0__abc_74955_new_n169_), .Y(u2_u0__abc_74955_new_n170_));
AND2X2 AND2X2_2762 ( .A(u2_u0__abc_74955_new_n171_), .B(u2_u0__abc_74955_new_n168_), .Y(u2_u0__0b3_last_row_12_0__6_));
AND2X2 AND2X2_2763 ( .A(u2_u0__abc_74955_new_n137__bF_buf4), .B(u2_u0__abc_74955_new_n174_), .Y(u2_u0__abc_74955_new_n175_));
AND2X2 AND2X2_2764 ( .A(u2_u0__abc_74955_new_n176_), .B(u2_u0__abc_74955_new_n173_), .Y(u2_u0__0b3_last_row_12_0__7_));
AND2X2 AND2X2_2765 ( .A(u2_u0__abc_74955_new_n137__bF_buf2), .B(u2_u0__abc_74955_new_n179_), .Y(u2_u0__abc_74955_new_n180_));
AND2X2 AND2X2_2766 ( .A(u2_u0__abc_74955_new_n181_), .B(u2_u0__abc_74955_new_n178_), .Y(u2_u0__0b3_last_row_12_0__8_));
AND2X2 AND2X2_2767 ( .A(u2_u0__abc_74955_new_n137__bF_buf0), .B(u2_u0__abc_74955_new_n184_), .Y(u2_u0__abc_74955_new_n185_));
AND2X2 AND2X2_2768 ( .A(u2_u0__abc_74955_new_n186_), .B(u2_u0__abc_74955_new_n183_), .Y(u2_u0__0b3_last_row_12_0__9_));
AND2X2 AND2X2_2769 ( .A(u2_u0__abc_74955_new_n137__bF_buf3), .B(u2_u0__abc_74955_new_n189_), .Y(u2_u0__abc_74955_new_n190_));
AND2X2 AND2X2_277 ( .A(u0__abc_76628_new_n1481_), .B(u0__abc_76628_new_n1172__bF_buf5), .Y(u0__abc_76628_new_n1482_));
AND2X2 AND2X2_2770 ( .A(u2_u0__abc_74955_new_n191_), .B(u2_u0__abc_74955_new_n188_), .Y(u2_u0__0b3_last_row_12_0__10_));
AND2X2 AND2X2_2771 ( .A(u2_u0__abc_74955_new_n137__bF_buf1), .B(u2_u0__abc_74955_new_n194_), .Y(u2_u0__abc_74955_new_n195_));
AND2X2 AND2X2_2772 ( .A(u2_u0__abc_74955_new_n196_), .B(u2_u0__abc_74955_new_n193_), .Y(u2_u0__0b3_last_row_12_0__11_));
AND2X2 AND2X2_2773 ( .A(u2_u0__abc_74955_new_n137__bF_buf4), .B(u2_u0__abc_74955_new_n199_), .Y(u2_u0__abc_74955_new_n200_));
AND2X2 AND2X2_2774 ( .A(u2_u0__abc_74955_new_n201_), .B(u2_u0__abc_74955_new_n198_), .Y(u2_u0__0b3_last_row_12_0__12_));
AND2X2 AND2X2_2775 ( .A(u2_u0__abc_74955_new_n203_), .B(u2_u0__abc_74955_new_n204_), .Y(u2_u0__abc_74955_new_n205_));
AND2X2 AND2X2_2776 ( .A(u2_u0__abc_74955_new_n205_), .B(u2_bank_set_0), .Y(u2_u0__abc_74955_new_n206_));
AND2X2 AND2X2_2777 ( .A(u2_u0__abc_74955_new_n209_), .B(u2_u0__abc_74955_new_n207_), .Y(u2_u0__0b0_last_row_12_0__0_));
AND2X2 AND2X2_2778 ( .A(u2_u0__abc_74955_new_n212_), .B(u2_u0__abc_74955_new_n211_), .Y(u2_u0__0b0_last_row_12_0__1_));
AND2X2 AND2X2_2779 ( .A(u2_u0__abc_74955_new_n215_), .B(u2_u0__abc_74955_new_n214_), .Y(u2_u0__0b0_last_row_12_0__2_));
AND2X2 AND2X2_278 ( .A(spec_req_cs_1_bF_buf2_), .B(u0_tms1_12_), .Y(u0__abc_76628_new_n1483_));
AND2X2 AND2X2_2780 ( .A(u2_u0__abc_74955_new_n218_), .B(u2_u0__abc_74955_new_n217_), .Y(u2_u0__0b0_last_row_12_0__3_));
AND2X2 AND2X2_2781 ( .A(u2_u0__abc_74955_new_n221_), .B(u2_u0__abc_74955_new_n220_), .Y(u2_u0__0b0_last_row_12_0__4_));
AND2X2 AND2X2_2782 ( .A(u2_u0__abc_74955_new_n224_), .B(u2_u0__abc_74955_new_n223_), .Y(u2_u0__0b0_last_row_12_0__5_));
AND2X2 AND2X2_2783 ( .A(u2_u0__abc_74955_new_n227_), .B(u2_u0__abc_74955_new_n226_), .Y(u2_u0__0b0_last_row_12_0__6_));
AND2X2 AND2X2_2784 ( .A(u2_u0__abc_74955_new_n230_), .B(u2_u0__abc_74955_new_n229_), .Y(u2_u0__0b0_last_row_12_0__7_));
AND2X2 AND2X2_2785 ( .A(u2_u0__abc_74955_new_n233_), .B(u2_u0__abc_74955_new_n232_), .Y(u2_u0__0b0_last_row_12_0__8_));
AND2X2 AND2X2_2786 ( .A(u2_u0__abc_74955_new_n236_), .B(u2_u0__abc_74955_new_n235_), .Y(u2_u0__0b0_last_row_12_0__9_));
AND2X2 AND2X2_2787 ( .A(u2_u0__abc_74955_new_n239_), .B(u2_u0__abc_74955_new_n238_), .Y(u2_u0__0b0_last_row_12_0__10_));
AND2X2 AND2X2_2788 ( .A(u2_u0__abc_74955_new_n242_), .B(u2_u0__abc_74955_new_n241_), .Y(u2_u0__0b0_last_row_12_0__11_));
AND2X2 AND2X2_2789 ( .A(u2_u0__abc_74955_new_n245_), .B(u2_u0__abc_74955_new_n244_), .Y(u2_u0__0b0_last_row_12_0__12_));
AND2X2 AND2X2_279 ( .A(u0__abc_76628_new_n1169__bF_buf0), .B(u0__abc_76628_new_n1486_), .Y(u0__abc_76628_new_n1487_));
AND2X2 AND2X2_2790 ( .A(u2_u0__abc_74955_new_n204_), .B(bank_adr_0_), .Y(u2_u0__abc_74955_new_n247_));
AND2X2 AND2X2_2791 ( .A(u2_u0__abc_74955_new_n247_), .B(u2_bank_set_0), .Y(u2_u0__abc_74955_new_n248_));
AND2X2 AND2X2_2792 ( .A(u2_u0__abc_74955_new_n251_), .B(u2_u0__abc_74955_new_n249_), .Y(u2_u0__0b1_last_row_12_0__0_));
AND2X2 AND2X2_2793 ( .A(u2_u0__abc_74955_new_n254_), .B(u2_u0__abc_74955_new_n253_), .Y(u2_u0__0b1_last_row_12_0__1_));
AND2X2 AND2X2_2794 ( .A(u2_u0__abc_74955_new_n257_), .B(u2_u0__abc_74955_new_n256_), .Y(u2_u0__0b1_last_row_12_0__2_));
AND2X2 AND2X2_2795 ( .A(u2_u0__abc_74955_new_n260_), .B(u2_u0__abc_74955_new_n259_), .Y(u2_u0__0b1_last_row_12_0__3_));
AND2X2 AND2X2_2796 ( .A(u2_u0__abc_74955_new_n263_), .B(u2_u0__abc_74955_new_n262_), .Y(u2_u0__0b1_last_row_12_0__4_));
AND2X2 AND2X2_2797 ( .A(u2_u0__abc_74955_new_n266_), .B(u2_u0__abc_74955_new_n265_), .Y(u2_u0__0b1_last_row_12_0__5_));
AND2X2 AND2X2_2798 ( .A(u2_u0__abc_74955_new_n269_), .B(u2_u0__abc_74955_new_n268_), .Y(u2_u0__0b1_last_row_12_0__6_));
AND2X2 AND2X2_2799 ( .A(u2_u0__abc_74955_new_n272_), .B(u2_u0__abc_74955_new_n271_), .Y(u2_u0__0b1_last_row_12_0__7_));
AND2X2 AND2X2_28 ( .A(_abc_85006_new_n320_), .B(_abc_85006_new_n321_), .Y(tms_s_10_));
AND2X2 AND2X2_280 ( .A(u0__abc_76628_new_n1485_), .B(u0__abc_76628_new_n1487_), .Y(u0__abc_76628_new_n1488_));
AND2X2 AND2X2_2800 ( .A(u2_u0__abc_74955_new_n275_), .B(u2_u0__abc_74955_new_n274_), .Y(u2_u0__0b1_last_row_12_0__8_));
AND2X2 AND2X2_2801 ( .A(u2_u0__abc_74955_new_n278_), .B(u2_u0__abc_74955_new_n277_), .Y(u2_u0__0b1_last_row_12_0__9_));
AND2X2 AND2X2_2802 ( .A(u2_u0__abc_74955_new_n281_), .B(u2_u0__abc_74955_new_n280_), .Y(u2_u0__0b1_last_row_12_0__10_));
AND2X2 AND2X2_2803 ( .A(u2_u0__abc_74955_new_n284_), .B(u2_u0__abc_74955_new_n283_), .Y(u2_u0__0b1_last_row_12_0__11_));
AND2X2 AND2X2_2804 ( .A(u2_u0__abc_74955_new_n287_), .B(u2_u0__abc_74955_new_n286_), .Y(u2_u0__0b1_last_row_12_0__12_));
AND2X2 AND2X2_2805 ( .A(u2_u0__abc_74955_new_n203_), .B(bank_adr_1_), .Y(u2_u0__abc_74955_new_n289_));
AND2X2 AND2X2_2806 ( .A(u2_u0__abc_74955_new_n289_), .B(u2_bank_set_0), .Y(u2_u0__abc_74955_new_n290_));
AND2X2 AND2X2_2807 ( .A(u2_u0__abc_74955_new_n293_), .B(u2_u0__abc_74955_new_n291_), .Y(u2_u0__0b2_last_row_12_0__0_));
AND2X2 AND2X2_2808 ( .A(u2_u0__abc_74955_new_n296_), .B(u2_u0__abc_74955_new_n295_), .Y(u2_u0__0b2_last_row_12_0__1_));
AND2X2 AND2X2_2809 ( .A(u2_u0__abc_74955_new_n299_), .B(u2_u0__abc_74955_new_n298_), .Y(u2_u0__0b2_last_row_12_0__2_));
AND2X2 AND2X2_281 ( .A(u0__abc_76628_new_n1170__bF_buf0), .B(sp_tms_13_), .Y(u0__abc_76628_new_n1490_));
AND2X2 AND2X2_2810 ( .A(u2_u0__abc_74955_new_n302_), .B(u2_u0__abc_74955_new_n301_), .Y(u2_u0__0b2_last_row_12_0__3_));
AND2X2 AND2X2_2811 ( .A(u2_u0__abc_74955_new_n305_), .B(u2_u0__abc_74955_new_n304_), .Y(u2_u0__0b2_last_row_12_0__4_));
AND2X2 AND2X2_2812 ( .A(u2_u0__abc_74955_new_n308_), .B(u2_u0__abc_74955_new_n307_), .Y(u2_u0__0b2_last_row_12_0__5_));
AND2X2 AND2X2_2813 ( .A(u2_u0__abc_74955_new_n311_), .B(u2_u0__abc_74955_new_n310_), .Y(u2_u0__0b2_last_row_12_0__6_));
AND2X2 AND2X2_2814 ( .A(u2_u0__abc_74955_new_n314_), .B(u2_u0__abc_74955_new_n313_), .Y(u2_u0__0b2_last_row_12_0__7_));
AND2X2 AND2X2_2815 ( .A(u2_u0__abc_74955_new_n317_), .B(u2_u0__abc_74955_new_n316_), .Y(u2_u0__0b2_last_row_12_0__8_));
AND2X2 AND2X2_2816 ( .A(u2_u0__abc_74955_new_n320_), .B(u2_u0__abc_74955_new_n319_), .Y(u2_u0__0b2_last_row_12_0__9_));
AND2X2 AND2X2_2817 ( .A(u2_u0__abc_74955_new_n323_), .B(u2_u0__abc_74955_new_n322_), .Y(u2_u0__0b2_last_row_12_0__10_));
AND2X2 AND2X2_2818 ( .A(u2_u0__abc_74955_new_n326_), .B(u2_u0__abc_74955_new_n325_), .Y(u2_u0__0b2_last_row_12_0__11_));
AND2X2 AND2X2_2819 ( .A(u2_u0__abc_74955_new_n329_), .B(u2_u0__abc_74955_new_n328_), .Y(u2_u0__0b2_last_row_12_0__12_));
AND2X2 AND2X2_282 ( .A(spec_req_cs_5_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1491_));
AND2X2 AND2X2_2820 ( .A(u2_u0__abc_74955_new_n333_), .B(u2_u0__abc_74955_new_n335_), .Y(u2_u0__abc_74955_new_n336_));
AND2X2 AND2X2_2821 ( .A(u2_u0__abc_74955_new_n336_), .B(u2_u0__abc_74955_new_n331_), .Y(u2_u0__abc_74955_new_n337_));
AND2X2 AND2X2_2822 ( .A(u2_u0__abc_74955_new_n338_), .B(u2_u0__abc_74955_new_n340_), .Y(u2_u0__abc_74955_new_n341_));
AND2X2 AND2X2_2823 ( .A(u2_u0__abc_74955_new_n343_), .B(u2_u0__abc_74955_new_n344_), .Y(u2_u0__abc_74955_new_n345_));
AND2X2 AND2X2_2824 ( .A(u2_u0__abc_74955_new_n341_), .B(u2_u0__abc_74955_new_n345_), .Y(u2_u0__abc_74955_new_n346_));
AND2X2 AND2X2_2825 ( .A(u2_u0__abc_74955_new_n346_), .B(u2_u0__abc_74955_new_n337_), .Y(u2_u0__abc_74955_new_n347_));
AND2X2 AND2X2_2826 ( .A(u2_u0__abc_74955_new_n348_), .B(u2_u0__abc_74955_new_n139_), .Y(u2_u0__abc_74955_new_n349_));
AND2X2 AND2X2_2827 ( .A(u2_u0_b3_last_row_0_), .B(row_adr_0_bF_buf1_), .Y(u2_u0__abc_74955_new_n350_));
AND2X2 AND2X2_2828 ( .A(u2_u0__abc_74955_new_n352_), .B(u2_u0__abc_74955_new_n136_), .Y(u2_u0__abc_74955_new_n353_));
AND2X2 AND2X2_2829 ( .A(u2_u0__abc_74955_new_n351_), .B(u2_u0__abc_74955_new_n353_), .Y(u2_u0__abc_74955_new_n354_));
AND2X2 AND2X2_283 ( .A(u0__abc_76628_new_n1493_), .B(u0__abc_76628_new_n1179__bF_buf4), .Y(u0__abc_76628_new_n1494_));
AND2X2 AND2X2_2830 ( .A(u2_u0__abc_74955_new_n356_), .B(u2_u0__abc_74955_new_n357_), .Y(u2_u0__abc_74955_new_n358_));
AND2X2 AND2X2_2831 ( .A(u2_u0__abc_74955_new_n360_), .B(u2_u0__abc_74955_new_n361_), .Y(u2_u0__abc_74955_new_n362_));
AND2X2 AND2X2_2832 ( .A(u2_u0__abc_74955_new_n358_), .B(u2_u0__abc_74955_new_n362_), .Y(u2_u0__abc_74955_new_n363_));
AND2X2 AND2X2_2833 ( .A(u2_u0__abc_74955_new_n363_), .B(u2_u0__abc_74955_new_n354_), .Y(u2_u0__abc_74955_new_n364_));
AND2X2 AND2X2_2834 ( .A(u2_u0__abc_74955_new_n347_), .B(u2_u0__abc_74955_new_n364_), .Y(u2_u0__abc_74955_new_n365_));
AND2X2 AND2X2_2835 ( .A(u2_u0__abc_74955_new_n366_), .B(u2_u0__abc_74955_new_n368_), .Y(u2_u0__abc_74955_new_n369_));
AND2X2 AND2X2_2836 ( .A(u2_u0__abc_74955_new_n370_), .B(u2_u0__abc_74955_new_n372_), .Y(u2_u0__abc_74955_new_n373_));
AND2X2 AND2X2_2837 ( .A(u2_u0__abc_74955_new_n369_), .B(u2_u0__abc_74955_new_n373_), .Y(u2_u0__abc_74955_new_n374_));
AND2X2 AND2X2_2838 ( .A(u2_u0__abc_74955_new_n376_), .B(u2_u0__abc_74955_new_n377_), .Y(u2_u0__abc_74955_new_n378_));
AND2X2 AND2X2_2839 ( .A(u2_u0__abc_74955_new_n380_), .B(u2_u0__abc_74955_new_n381_), .Y(u2_u0__abc_74955_new_n382_));
AND2X2 AND2X2_284 ( .A(u0__abc_76628_new_n1494_), .B(u0__abc_76628_new_n1492_), .Y(u0__abc_76628_new_n1495_));
AND2X2 AND2X2_2840 ( .A(u2_u0__abc_74955_new_n378_), .B(u2_u0__abc_74955_new_n382_), .Y(u2_u0__abc_74955_new_n383_));
AND2X2 AND2X2_2841 ( .A(u2_u0__abc_74955_new_n384_), .B(u2_u0__abc_74955_new_n386_), .Y(u2_u0__abc_74955_new_n387_));
AND2X2 AND2X2_2842 ( .A(u2_u0__abc_74955_new_n389_), .B(u2_u0__abc_74955_new_n390_), .Y(u2_u0__abc_74955_new_n391_));
AND2X2 AND2X2_2843 ( .A(u2_u0__abc_74955_new_n387_), .B(u2_u0__abc_74955_new_n391_), .Y(u2_u0__abc_74955_new_n392_));
AND2X2 AND2X2_2844 ( .A(u2_u0__abc_74955_new_n383_), .B(u2_u0__abc_74955_new_n392_), .Y(u2_u0__abc_74955_new_n393_));
AND2X2 AND2X2_2845 ( .A(u2_u0__abc_74955_new_n393_), .B(u2_u0__abc_74955_new_n374_), .Y(u2_u0__abc_74955_new_n394_));
AND2X2 AND2X2_2846 ( .A(u2_u0__abc_74955_new_n365_), .B(u2_u0__abc_74955_new_n394_), .Y(u2_u0__abc_74955_new_n395_));
AND2X2 AND2X2_2847 ( .A(u2_u0__abc_74955_new_n396_), .B(u2_u0__abc_74955_new_n397_), .Y(u2_u0__abc_74955_new_n398_));
AND2X2 AND2X2_2848 ( .A(u2_u0__abc_74955_new_n398_), .B(u2_u0__abc_74955_new_n400_), .Y(u2_u0__abc_74955_new_n401_));
AND2X2 AND2X2_2849 ( .A(u2_u0__abc_74955_new_n402_), .B(u2_u0__abc_74955_new_n404_), .Y(u2_u0__abc_74955_new_n405_));
AND2X2 AND2X2_285 ( .A(u0__abc_76628_new_n1496_), .B(u0__abc_76628_new_n1175__bF_buf4), .Y(u0__abc_76628_new_n1497_));
AND2X2 AND2X2_2850 ( .A(u2_u0__abc_74955_new_n406_), .B(u2_u0__abc_74955_new_n408_), .Y(u2_u0__abc_74955_new_n409_));
AND2X2 AND2X2_2851 ( .A(u2_u0__abc_74955_new_n405_), .B(u2_u0__abc_74955_new_n409_), .Y(u2_u0__abc_74955_new_n410_));
AND2X2 AND2X2_2852 ( .A(u2_u0__abc_74955_new_n410_), .B(u2_u0__abc_74955_new_n401_), .Y(u2_u0__abc_74955_new_n411_));
AND2X2 AND2X2_2853 ( .A(u2_u0__abc_74955_new_n412_), .B(u2_u0__abc_74955_new_n414_), .Y(u2_u0__abc_74955_new_n415_));
AND2X2 AND2X2_2854 ( .A(u2_u0__abc_74955_new_n416_), .B(u2_u0__abc_74955_new_n418_), .Y(u2_u0__abc_74955_new_n419_));
AND2X2 AND2X2_2855 ( .A(u2_u0__abc_74955_new_n415_), .B(u2_u0__abc_74955_new_n419_), .Y(u2_u0__abc_74955_new_n420_));
AND2X2 AND2X2_2856 ( .A(u2_u0__abc_74955_new_n421_), .B(u2_u0__abc_74955_new_n423_), .Y(u2_u0__abc_74955_new_n424_));
AND2X2 AND2X2_2857 ( .A(u2_u0__abc_74955_new_n426_), .B(u2_u0__abc_74955_new_n247_), .Y(u2_u0__abc_74955_new_n427_));
AND2X2 AND2X2_2858 ( .A(u2_u0__abc_74955_new_n424_), .B(u2_u0__abc_74955_new_n427_), .Y(u2_u0__abc_74955_new_n428_));
AND2X2 AND2X2_2859 ( .A(u2_u0__abc_74955_new_n420_), .B(u2_u0__abc_74955_new_n428_), .Y(u2_u0__abc_74955_new_n429_));
AND2X2 AND2X2_286 ( .A(spec_req_cs_4_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1498_));
AND2X2 AND2X2_2860 ( .A(u2_u0__abc_74955_new_n411_), .B(u2_u0__abc_74955_new_n429_), .Y(u2_u0__abc_74955_new_n430_));
AND2X2 AND2X2_2861 ( .A(u2_u0__abc_74955_new_n432_), .B(u2_u0__abc_74955_new_n433_), .Y(u2_u0__abc_74955_new_n434_));
AND2X2 AND2X2_2862 ( .A(u2_u0__abc_74955_new_n436_), .B(u2_u0__abc_74955_new_n437_), .Y(u2_u0__abc_74955_new_n438_));
AND2X2 AND2X2_2863 ( .A(u2_u0__abc_74955_new_n434_), .B(u2_u0__abc_74955_new_n438_), .Y(u2_u0__abc_74955_new_n439_));
AND2X2 AND2X2_2864 ( .A(u2_u0__abc_74955_new_n441_), .B(u2_u0__abc_74955_new_n442_), .Y(u2_u0__abc_74955_new_n443_));
AND2X2 AND2X2_2865 ( .A(u2_u0__abc_74955_new_n445_), .B(u2_u0__abc_74955_new_n446_), .Y(u2_u0__abc_74955_new_n447_));
AND2X2 AND2X2_2866 ( .A(u2_u0__abc_74955_new_n443_), .B(u2_u0__abc_74955_new_n447_), .Y(u2_u0__abc_74955_new_n448_));
AND2X2 AND2X2_2867 ( .A(u2_u0__abc_74955_new_n449_), .B(u2_u0__abc_74955_new_n451_), .Y(u2_u0__abc_74955_new_n452_));
AND2X2 AND2X2_2868 ( .A(u2_u0__abc_74955_new_n453_), .B(u2_u0__abc_74955_new_n455_), .Y(u2_u0__abc_74955_new_n456_));
AND2X2 AND2X2_2869 ( .A(u2_u0__abc_74955_new_n452_), .B(u2_u0__abc_74955_new_n456_), .Y(u2_u0__abc_74955_new_n457_));
AND2X2 AND2X2_287 ( .A(u0__abc_76628_new_n1499_), .B(u0__abc_76628_new_n1174__bF_buf4), .Y(u0__abc_76628_new_n1500_));
AND2X2 AND2X2_2870 ( .A(u2_u0__abc_74955_new_n448_), .B(u2_u0__abc_74955_new_n457_), .Y(u2_u0__abc_74955_new_n458_));
AND2X2 AND2X2_2871 ( .A(u2_u0__abc_74955_new_n458_), .B(u2_u0__abc_74955_new_n439_), .Y(u2_u0__abc_74955_new_n459_));
AND2X2 AND2X2_2872 ( .A(u2_u0__abc_74955_new_n430_), .B(u2_u0__abc_74955_new_n459_), .Y(u2_u0__abc_74955_new_n460_));
AND2X2 AND2X2_2873 ( .A(u2_u0__abc_74955_new_n464_), .B(u2_u0__abc_74955_new_n465_), .Y(u2_u0__abc_74955_new_n466_));
AND2X2 AND2X2_2874 ( .A(u2_u0__abc_74955_new_n466_), .B(u2_u0__abc_74955_new_n463_), .Y(u2_u0__abc_74955_new_n467_));
AND2X2 AND2X2_2875 ( .A(u2_u0__abc_74955_new_n468_), .B(u2_u0__abc_74955_new_n470_), .Y(u2_u0__abc_74955_new_n471_));
AND2X2 AND2X2_2876 ( .A(u2_u0__abc_74955_new_n473_), .B(u2_u0__abc_74955_new_n474_), .Y(u2_u0__abc_74955_new_n475_));
AND2X2 AND2X2_2877 ( .A(u2_u0__abc_74955_new_n471_), .B(u2_u0__abc_74955_new_n475_), .Y(u2_u0__abc_74955_new_n476_));
AND2X2 AND2X2_2878 ( .A(u2_u0__abc_74955_new_n478_), .B(u2_u0__abc_74955_new_n480_), .Y(u2_u0__abc_74955_new_n481_));
AND2X2 AND2X2_2879 ( .A(u2_u0__abc_74955_new_n482_), .B(u2_u0__abc_74955_new_n483_), .Y(u2_u0__abc_74955_new_n484_));
AND2X2 AND2X2_288 ( .A(spec_req_cs_3_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1501_));
AND2X2 AND2X2_2880 ( .A(u2_u0__abc_74955_new_n481_), .B(u2_u0__abc_74955_new_n484_), .Y(u2_u0__abc_74955_new_n485_));
AND2X2 AND2X2_2881 ( .A(u2_u0__abc_74955_new_n476_), .B(u2_u0__abc_74955_new_n485_), .Y(u2_u0__abc_74955_new_n486_));
AND2X2 AND2X2_2882 ( .A(u2_u0__abc_74955_new_n486_), .B(u2_u0__abc_74955_new_n467_), .Y(u2_u0__abc_74955_new_n487_));
AND2X2 AND2X2_2883 ( .A(u2_u0__abc_74955_new_n139_), .B(u2_u0__abc_74955_new_n488_), .Y(u2_u0__abc_74955_new_n489_));
AND2X2 AND2X2_2884 ( .A(row_adr_0_bF_buf3_), .B(u2_u0_b0_last_row_0_), .Y(u2_u0__abc_74955_new_n490_));
AND2X2 AND2X2_2885 ( .A(u2_u0__abc_74955_new_n493_), .B(u2_u0__abc_74955_new_n494_), .Y(u2_u0__abc_74955_new_n495_));
AND2X2 AND2X2_2886 ( .A(u2_u0__abc_74955_new_n491_), .B(u2_u0__abc_74955_new_n495_), .Y(u2_u0__abc_74955_new_n496_));
AND2X2 AND2X2_2887 ( .A(u2_u0__abc_74955_new_n497_), .B(u2_u0__abc_74955_new_n499_), .Y(u2_u0__abc_74955_new_n500_));
AND2X2 AND2X2_2888 ( .A(u2_u0__abc_74955_new_n502_), .B(u2_u0__abc_74955_new_n205_), .Y(u2_u0__abc_74955_new_n503_));
AND2X2 AND2X2_2889 ( .A(u2_u0__abc_74955_new_n500_), .B(u2_u0__abc_74955_new_n503_), .Y(u2_u0__abc_74955_new_n504_));
AND2X2 AND2X2_289 ( .A(u0__abc_76628_new_n1502_), .B(u0__abc_76628_new_n1173__bF_buf4), .Y(u0__abc_76628_new_n1503_));
AND2X2 AND2X2_2890 ( .A(u2_u0__abc_74955_new_n496_), .B(u2_u0__abc_74955_new_n504_), .Y(u2_u0__abc_74955_new_n505_));
AND2X2 AND2X2_2891 ( .A(u2_u0__abc_74955_new_n507_), .B(u2_u0__abc_74955_new_n509_), .Y(u2_u0__abc_74955_new_n510_));
AND2X2 AND2X2_2892 ( .A(u2_u0__abc_74955_new_n511_), .B(u2_u0__abc_74955_new_n512_), .Y(u2_u0__abc_74955_new_n513_));
AND2X2 AND2X2_2893 ( .A(u2_u0__abc_74955_new_n510_), .B(u2_u0__abc_74955_new_n513_), .Y(u2_u0__abc_74955_new_n514_));
AND2X2 AND2X2_2894 ( .A(u2_u0__abc_74955_new_n515_), .B(u2_u0__abc_74955_new_n517_), .Y(u2_u0__abc_74955_new_n518_));
AND2X2 AND2X2_2895 ( .A(u2_u0__abc_74955_new_n519_), .B(u2_u0__abc_74955_new_n521_), .Y(u2_u0__abc_74955_new_n522_));
AND2X2 AND2X2_2896 ( .A(u2_u0__abc_74955_new_n518_), .B(u2_u0__abc_74955_new_n522_), .Y(u2_u0__abc_74955_new_n523_));
AND2X2 AND2X2_2897 ( .A(u2_u0__abc_74955_new_n514_), .B(u2_u0__abc_74955_new_n523_), .Y(u2_u0__abc_74955_new_n524_));
AND2X2 AND2X2_2898 ( .A(u2_u0__abc_74955_new_n524_), .B(u2_u0__abc_74955_new_n505_), .Y(u2_u0__abc_74955_new_n525_));
AND2X2 AND2X2_2899 ( .A(u2_u0__abc_74955_new_n487_), .B(u2_u0__abc_74955_new_n525_), .Y(u2_u0__abc_74955_new_n526_));
AND2X2 AND2X2_29 ( .A(_abc_85006_new_n323_), .B(_abc_85006_new_n324_), .Y(tms_s_11_));
AND2X2 AND2X2_290 ( .A(spec_req_cs_2_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1504_));
AND2X2 AND2X2_2900 ( .A(u2_u0__abc_74955_new_n529_), .B(u2_u0__abc_74955_new_n530_), .Y(u2_u0__abc_74955_new_n531_));
AND2X2 AND2X2_2901 ( .A(u2_u0__abc_74955_new_n531_), .B(u2_u0__abc_74955_new_n528_), .Y(u2_u0__abc_74955_new_n532_));
AND2X2 AND2X2_2902 ( .A(u2_u0__abc_74955_new_n534_), .B(u2_u0__abc_74955_new_n535_), .Y(u2_u0__abc_74955_new_n536_));
AND2X2 AND2X2_2903 ( .A(u2_u0__abc_74955_new_n538_), .B(u2_u0__abc_74955_new_n539_), .Y(u2_u0__abc_74955_new_n540_));
AND2X2 AND2X2_2904 ( .A(u2_u0__abc_74955_new_n536_), .B(u2_u0__abc_74955_new_n540_), .Y(u2_u0__abc_74955_new_n541_));
AND2X2 AND2X2_2905 ( .A(u2_u0__abc_74955_new_n541_), .B(u2_u0__abc_74955_new_n532_), .Y(u2_u0__abc_74955_new_n542_));
AND2X2 AND2X2_2906 ( .A(u2_u0__abc_74955_new_n543_), .B(u2_u0__abc_74955_new_n545_), .Y(u2_u0__abc_74955_new_n546_));
AND2X2 AND2X2_2907 ( .A(u2_u0__abc_74955_new_n547_), .B(u2_u0__abc_74955_new_n549_), .Y(u2_u0__abc_74955_new_n550_));
AND2X2 AND2X2_2908 ( .A(u2_u0__abc_74955_new_n546_), .B(u2_u0__abc_74955_new_n550_), .Y(u2_u0__abc_74955_new_n551_));
AND2X2 AND2X2_2909 ( .A(u2_u0__abc_74955_new_n552_), .B(u2_u0__abc_74955_new_n554_), .Y(u2_u0__abc_74955_new_n555_));
AND2X2 AND2X2_291 ( .A(u0__abc_76628_new_n1505_), .B(u0__abc_76628_new_n1172__bF_buf4), .Y(u0__abc_76628_new_n1506_));
AND2X2 AND2X2_2910 ( .A(u2_u0__abc_74955_new_n556_), .B(u2_u0__abc_74955_new_n558_), .Y(u2_u0__abc_74955_new_n559_));
AND2X2 AND2X2_2911 ( .A(u2_u0__abc_74955_new_n555_), .B(u2_u0__abc_74955_new_n559_), .Y(u2_u0__abc_74955_new_n560_));
AND2X2 AND2X2_2912 ( .A(u2_u0__abc_74955_new_n551_), .B(u2_u0__abc_74955_new_n560_), .Y(u2_u0__abc_74955_new_n561_));
AND2X2 AND2X2_2913 ( .A(u2_u0__abc_74955_new_n561_), .B(u2_u0__abc_74955_new_n542_), .Y(u2_u0__abc_74955_new_n562_));
AND2X2 AND2X2_2914 ( .A(u2_u0__abc_74955_new_n564_), .B(u2_u0__abc_74955_new_n565_), .Y(u2_u0__abc_74955_new_n566_));
AND2X2 AND2X2_2915 ( .A(u2_u0__abc_74955_new_n568_), .B(u2_u0__abc_74955_new_n569_), .Y(u2_u0__abc_74955_new_n570_));
AND2X2 AND2X2_2916 ( .A(u2_u0__abc_74955_new_n566_), .B(u2_u0__abc_74955_new_n570_), .Y(u2_u0__abc_74955_new_n571_));
AND2X2 AND2X2_2917 ( .A(u2_u0__abc_74955_new_n572_), .B(u2_u0__abc_74955_new_n574_), .Y(u2_u0__abc_74955_new_n575_));
AND2X2 AND2X2_2918 ( .A(u2_u0__abc_74955_new_n576_), .B(u2_u0__abc_74955_new_n578_), .Y(u2_u0__abc_74955_new_n579_));
AND2X2 AND2X2_2919 ( .A(u2_u0__abc_74955_new_n575_), .B(u2_u0__abc_74955_new_n579_), .Y(u2_u0__abc_74955_new_n580_));
AND2X2 AND2X2_292 ( .A(spec_req_cs_1_bF_buf1_), .B(u0_tms1_13_), .Y(u0__abc_76628_new_n1507_));
AND2X2 AND2X2_2920 ( .A(u2_u0__abc_74955_new_n581_), .B(u2_u0__abc_74955_new_n583_), .Y(u2_u0__abc_74955_new_n584_));
AND2X2 AND2X2_2921 ( .A(u2_u0__abc_74955_new_n586_), .B(u2_u0__abc_74955_new_n289_), .Y(u2_u0__abc_74955_new_n587_));
AND2X2 AND2X2_2922 ( .A(u2_u0__abc_74955_new_n584_), .B(u2_u0__abc_74955_new_n587_), .Y(u2_u0__abc_74955_new_n588_));
AND2X2 AND2X2_2923 ( .A(u2_u0__abc_74955_new_n580_), .B(u2_u0__abc_74955_new_n588_), .Y(u2_u0__abc_74955_new_n589_));
AND2X2 AND2X2_2924 ( .A(u2_u0__abc_74955_new_n589_), .B(u2_u0__abc_74955_new_n571_), .Y(u2_u0__abc_74955_new_n590_));
AND2X2 AND2X2_2925 ( .A(u2_u0__abc_74955_new_n562_), .B(u2_u0__abc_74955_new_n590_), .Y(u2_u0__abc_74955_new_n591_));
AND2X2 AND2X2_2926 ( .A(u2_u0__abc_74955_new_n289_), .B(u2_u0_bank2_open), .Y(u2_u0__abc_74955_new_n594_));
AND2X2 AND2X2_2927 ( .A(u2_u0__abc_74955_new_n136_), .B(u2_u0_bank3_open), .Y(u2_u0__abc_74955_new_n595_));
AND2X2 AND2X2_2928 ( .A(u2_u0__abc_74955_new_n205_), .B(u2_u0_bank0_open), .Y(u2_u0__abc_74955_new_n597_));
AND2X2 AND2X2_2929 ( .A(u2_u0__abc_74955_new_n247_), .B(u2_u0_bank1_open), .Y(u2_u0__abc_74955_new_n598_));
AND2X2 AND2X2_293 ( .A(u0__abc_76628_new_n1169__bF_buf6), .B(u0__abc_76628_new_n1510_), .Y(u0__abc_76628_new_n1511_));
AND2X2 AND2X2_2930 ( .A(u2_u0__abc_74955_new_n604_), .B(u2_u0_bank2_open), .Y(u2_u0__abc_74955_new_n605_));
AND2X2 AND2X2_2931 ( .A(u2_u0__abc_74955_new_n603_), .B(u2_u0__abc_74955_new_n605_), .Y(u2_u0__abc_74955_new_n606_));
AND2X2 AND2X2_2932 ( .A(u2_u0__abc_74955_new_n136_), .B(u2_bank_clr_0), .Y(u2_u0__abc_74955_new_n608_));
AND2X2 AND2X2_2933 ( .A(u2_u0__abc_74955_new_n604_), .B(u2_u0_bank3_open), .Y(u2_u0__abc_74955_new_n610_));
AND2X2 AND2X2_2934 ( .A(u2_u0__abc_74955_new_n609_), .B(u2_u0__abc_74955_new_n610_), .Y(u2_u0__abc_74955_new_n611_));
AND2X2 AND2X2_2935 ( .A(u2_u0__abc_74955_new_n604_), .B(u2_u0_bank1_open), .Y(u2_u0__abc_74955_new_n618_));
AND2X2 AND2X2_2936 ( .A(u2_u0__abc_74955_new_n617_), .B(u2_u0__abc_74955_new_n618_), .Y(u2_u0__abc_74955_new_n619_));
AND2X2 AND2X2_2937 ( .A(u2_u0__abc_74955_new_n604_), .B(u2_u0_bank0_open), .Y(u2_u0__abc_74955_new_n623_));
AND2X2 AND2X2_2938 ( .A(u2_u0__abc_74955_new_n622_), .B(u2_u0__abc_74955_new_n623_), .Y(u2_u0__abc_74955_new_n624_));
AND2X2 AND2X2_2939 ( .A(bank_adr_0_), .B(bank_adr_1_), .Y(u2_u1__abc_74955_new_n136_));
AND2X2 AND2X2_294 ( .A(u0__abc_76628_new_n1509_), .B(u0__abc_76628_new_n1511_), .Y(u0__abc_76628_new_n1512_));
AND2X2 AND2X2_2940 ( .A(u2_u1__abc_74955_new_n136_), .B(u2_bank_set_1), .Y(u2_u1__abc_74955_new_n137_));
AND2X2 AND2X2_2941 ( .A(u2_u1__abc_74955_new_n137__bF_buf3), .B(u2_u1__abc_74955_new_n139_), .Y(u2_u1__abc_74955_new_n140_));
AND2X2 AND2X2_2942 ( .A(u2_u1__abc_74955_new_n141_), .B(u2_u1__abc_74955_new_n138_), .Y(u2_u1__0b3_last_row_12_0__0_));
AND2X2 AND2X2_2943 ( .A(u2_u1__abc_74955_new_n137__bF_buf1), .B(u2_u1__abc_74955_new_n144_), .Y(u2_u1__abc_74955_new_n145_));
AND2X2 AND2X2_2944 ( .A(u2_u1__abc_74955_new_n146_), .B(u2_u1__abc_74955_new_n143_), .Y(u2_u1__0b3_last_row_12_0__1_));
AND2X2 AND2X2_2945 ( .A(u2_u1__abc_74955_new_n137__bF_buf4), .B(u2_u1__abc_74955_new_n149_), .Y(u2_u1__abc_74955_new_n150_));
AND2X2 AND2X2_2946 ( .A(u2_u1__abc_74955_new_n151_), .B(u2_u1__abc_74955_new_n148_), .Y(u2_u1__0b3_last_row_12_0__2_));
AND2X2 AND2X2_2947 ( .A(u2_u1__abc_74955_new_n137__bF_buf2), .B(u2_u1__abc_74955_new_n154_), .Y(u2_u1__abc_74955_new_n155_));
AND2X2 AND2X2_2948 ( .A(u2_u1__abc_74955_new_n156_), .B(u2_u1__abc_74955_new_n153_), .Y(u2_u1__0b3_last_row_12_0__3_));
AND2X2 AND2X2_2949 ( .A(u2_u1__abc_74955_new_n137__bF_buf0), .B(u2_u1__abc_74955_new_n159_), .Y(u2_u1__abc_74955_new_n160_));
AND2X2 AND2X2_295 ( .A(u0__abc_76628_new_n1170__bF_buf6), .B(sp_tms_14_), .Y(u0__abc_76628_new_n1514_));
AND2X2 AND2X2_2950 ( .A(u2_u1__abc_74955_new_n161_), .B(u2_u1__abc_74955_new_n158_), .Y(u2_u1__0b3_last_row_12_0__4_));
AND2X2 AND2X2_2951 ( .A(u2_u1__abc_74955_new_n137__bF_buf3), .B(u2_u1__abc_74955_new_n164_), .Y(u2_u1__abc_74955_new_n165_));
AND2X2 AND2X2_2952 ( .A(u2_u1__abc_74955_new_n166_), .B(u2_u1__abc_74955_new_n163_), .Y(u2_u1__0b3_last_row_12_0__5_));
AND2X2 AND2X2_2953 ( .A(u2_u1__abc_74955_new_n137__bF_buf1), .B(u2_u1__abc_74955_new_n169_), .Y(u2_u1__abc_74955_new_n170_));
AND2X2 AND2X2_2954 ( .A(u2_u1__abc_74955_new_n171_), .B(u2_u1__abc_74955_new_n168_), .Y(u2_u1__0b3_last_row_12_0__6_));
AND2X2 AND2X2_2955 ( .A(u2_u1__abc_74955_new_n137__bF_buf4), .B(u2_u1__abc_74955_new_n174_), .Y(u2_u1__abc_74955_new_n175_));
AND2X2 AND2X2_2956 ( .A(u2_u1__abc_74955_new_n176_), .B(u2_u1__abc_74955_new_n173_), .Y(u2_u1__0b3_last_row_12_0__7_));
AND2X2 AND2X2_2957 ( .A(u2_u1__abc_74955_new_n137__bF_buf2), .B(u2_u1__abc_74955_new_n179_), .Y(u2_u1__abc_74955_new_n180_));
AND2X2 AND2X2_2958 ( .A(u2_u1__abc_74955_new_n181_), .B(u2_u1__abc_74955_new_n178_), .Y(u2_u1__0b3_last_row_12_0__8_));
AND2X2 AND2X2_2959 ( .A(u2_u1__abc_74955_new_n137__bF_buf0), .B(u2_u1__abc_74955_new_n184_), .Y(u2_u1__abc_74955_new_n185_));
AND2X2 AND2X2_296 ( .A(spec_req_cs_5_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1515_));
AND2X2 AND2X2_2960 ( .A(u2_u1__abc_74955_new_n186_), .B(u2_u1__abc_74955_new_n183_), .Y(u2_u1__0b3_last_row_12_0__9_));
AND2X2 AND2X2_2961 ( .A(u2_u1__abc_74955_new_n137__bF_buf3), .B(u2_u1__abc_74955_new_n189_), .Y(u2_u1__abc_74955_new_n190_));
AND2X2 AND2X2_2962 ( .A(u2_u1__abc_74955_new_n191_), .B(u2_u1__abc_74955_new_n188_), .Y(u2_u1__0b3_last_row_12_0__10_));
AND2X2 AND2X2_2963 ( .A(u2_u1__abc_74955_new_n137__bF_buf1), .B(u2_u1__abc_74955_new_n194_), .Y(u2_u1__abc_74955_new_n195_));
AND2X2 AND2X2_2964 ( .A(u2_u1__abc_74955_new_n196_), .B(u2_u1__abc_74955_new_n193_), .Y(u2_u1__0b3_last_row_12_0__11_));
AND2X2 AND2X2_2965 ( .A(u2_u1__abc_74955_new_n137__bF_buf4), .B(u2_u1__abc_74955_new_n199_), .Y(u2_u1__abc_74955_new_n200_));
AND2X2 AND2X2_2966 ( .A(u2_u1__abc_74955_new_n201_), .B(u2_u1__abc_74955_new_n198_), .Y(u2_u1__0b3_last_row_12_0__12_));
AND2X2 AND2X2_2967 ( .A(u2_u1__abc_74955_new_n203_), .B(u2_u1__abc_74955_new_n204_), .Y(u2_u1__abc_74955_new_n205_));
AND2X2 AND2X2_2968 ( .A(u2_u1__abc_74955_new_n205_), .B(u2_bank_set_1), .Y(u2_u1__abc_74955_new_n206_));
AND2X2 AND2X2_2969 ( .A(u2_u1__abc_74955_new_n209_), .B(u2_u1__abc_74955_new_n207_), .Y(u2_u1__0b0_last_row_12_0__0_));
AND2X2 AND2X2_297 ( .A(u0__abc_76628_new_n1517_), .B(u0__abc_76628_new_n1179__bF_buf3), .Y(u0__abc_76628_new_n1518_));
AND2X2 AND2X2_2970 ( .A(u2_u1__abc_74955_new_n212_), .B(u2_u1__abc_74955_new_n211_), .Y(u2_u1__0b0_last_row_12_0__1_));
AND2X2 AND2X2_2971 ( .A(u2_u1__abc_74955_new_n215_), .B(u2_u1__abc_74955_new_n214_), .Y(u2_u1__0b0_last_row_12_0__2_));
AND2X2 AND2X2_2972 ( .A(u2_u1__abc_74955_new_n218_), .B(u2_u1__abc_74955_new_n217_), .Y(u2_u1__0b0_last_row_12_0__3_));
AND2X2 AND2X2_2973 ( .A(u2_u1__abc_74955_new_n221_), .B(u2_u1__abc_74955_new_n220_), .Y(u2_u1__0b0_last_row_12_0__4_));
AND2X2 AND2X2_2974 ( .A(u2_u1__abc_74955_new_n224_), .B(u2_u1__abc_74955_new_n223_), .Y(u2_u1__0b0_last_row_12_0__5_));
AND2X2 AND2X2_2975 ( .A(u2_u1__abc_74955_new_n227_), .B(u2_u1__abc_74955_new_n226_), .Y(u2_u1__0b0_last_row_12_0__6_));
AND2X2 AND2X2_2976 ( .A(u2_u1__abc_74955_new_n230_), .B(u2_u1__abc_74955_new_n229_), .Y(u2_u1__0b0_last_row_12_0__7_));
AND2X2 AND2X2_2977 ( .A(u2_u1__abc_74955_new_n233_), .B(u2_u1__abc_74955_new_n232_), .Y(u2_u1__0b0_last_row_12_0__8_));
AND2X2 AND2X2_2978 ( .A(u2_u1__abc_74955_new_n236_), .B(u2_u1__abc_74955_new_n235_), .Y(u2_u1__0b0_last_row_12_0__9_));
AND2X2 AND2X2_2979 ( .A(u2_u1__abc_74955_new_n239_), .B(u2_u1__abc_74955_new_n238_), .Y(u2_u1__0b0_last_row_12_0__10_));
AND2X2 AND2X2_298 ( .A(u0__abc_76628_new_n1518_), .B(u0__abc_76628_new_n1516_), .Y(u0__abc_76628_new_n1519_));
AND2X2 AND2X2_2980 ( .A(u2_u1__abc_74955_new_n242_), .B(u2_u1__abc_74955_new_n241_), .Y(u2_u1__0b0_last_row_12_0__11_));
AND2X2 AND2X2_2981 ( .A(u2_u1__abc_74955_new_n245_), .B(u2_u1__abc_74955_new_n244_), .Y(u2_u1__0b0_last_row_12_0__12_));
AND2X2 AND2X2_2982 ( .A(u2_u1__abc_74955_new_n204_), .B(bank_adr_0_), .Y(u2_u1__abc_74955_new_n247_));
AND2X2 AND2X2_2983 ( .A(u2_u1__abc_74955_new_n247_), .B(u2_bank_set_1), .Y(u2_u1__abc_74955_new_n248_));
AND2X2 AND2X2_2984 ( .A(u2_u1__abc_74955_new_n251_), .B(u2_u1__abc_74955_new_n249_), .Y(u2_u1__0b1_last_row_12_0__0_));
AND2X2 AND2X2_2985 ( .A(u2_u1__abc_74955_new_n254_), .B(u2_u1__abc_74955_new_n253_), .Y(u2_u1__0b1_last_row_12_0__1_));
AND2X2 AND2X2_2986 ( .A(u2_u1__abc_74955_new_n257_), .B(u2_u1__abc_74955_new_n256_), .Y(u2_u1__0b1_last_row_12_0__2_));
AND2X2 AND2X2_2987 ( .A(u2_u1__abc_74955_new_n260_), .B(u2_u1__abc_74955_new_n259_), .Y(u2_u1__0b1_last_row_12_0__3_));
AND2X2 AND2X2_2988 ( .A(u2_u1__abc_74955_new_n263_), .B(u2_u1__abc_74955_new_n262_), .Y(u2_u1__0b1_last_row_12_0__4_));
AND2X2 AND2X2_2989 ( .A(u2_u1__abc_74955_new_n266_), .B(u2_u1__abc_74955_new_n265_), .Y(u2_u1__0b1_last_row_12_0__5_));
AND2X2 AND2X2_299 ( .A(u0__abc_76628_new_n1520_), .B(u0__abc_76628_new_n1175__bF_buf3), .Y(u0__abc_76628_new_n1521_));
AND2X2 AND2X2_2990 ( .A(u2_u1__abc_74955_new_n269_), .B(u2_u1__abc_74955_new_n268_), .Y(u2_u1__0b1_last_row_12_0__6_));
AND2X2 AND2X2_2991 ( .A(u2_u1__abc_74955_new_n272_), .B(u2_u1__abc_74955_new_n271_), .Y(u2_u1__0b1_last_row_12_0__7_));
AND2X2 AND2X2_2992 ( .A(u2_u1__abc_74955_new_n275_), .B(u2_u1__abc_74955_new_n274_), .Y(u2_u1__0b1_last_row_12_0__8_));
AND2X2 AND2X2_2993 ( .A(u2_u1__abc_74955_new_n278_), .B(u2_u1__abc_74955_new_n277_), .Y(u2_u1__0b1_last_row_12_0__9_));
AND2X2 AND2X2_2994 ( .A(u2_u1__abc_74955_new_n281_), .B(u2_u1__abc_74955_new_n280_), .Y(u2_u1__0b1_last_row_12_0__10_));
AND2X2 AND2X2_2995 ( .A(u2_u1__abc_74955_new_n284_), .B(u2_u1__abc_74955_new_n283_), .Y(u2_u1__0b1_last_row_12_0__11_));
AND2X2 AND2X2_2996 ( .A(u2_u1__abc_74955_new_n287_), .B(u2_u1__abc_74955_new_n286_), .Y(u2_u1__0b1_last_row_12_0__12_));
AND2X2 AND2X2_2997 ( .A(u2_u1__abc_74955_new_n203_), .B(bank_adr_1_), .Y(u2_u1__abc_74955_new_n289_));
AND2X2 AND2X2_2998 ( .A(u2_u1__abc_74955_new_n289_), .B(u2_bank_set_1), .Y(u2_u1__abc_74955_new_n290_));
AND2X2 AND2X2_2999 ( .A(u2_u1__abc_74955_new_n293_), .B(u2_u1__abc_74955_new_n291_), .Y(u2_u1__0b2_last_row_12_0__0_));
AND2X2 AND2X2_3 ( .A(_abc_85006_new_n244_), .B(_abc_85006_new_n246_), .Y(obct_cs_0_));
AND2X2 AND2X2_30 ( .A(_abc_85006_new_n326_), .B(_abc_85006_new_n327_), .Y(tms_s_12_));
AND2X2 AND2X2_300 ( .A(spec_req_cs_4_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1522_));
AND2X2 AND2X2_3000 ( .A(u2_u1__abc_74955_new_n296_), .B(u2_u1__abc_74955_new_n295_), .Y(u2_u1__0b2_last_row_12_0__1_));
AND2X2 AND2X2_3001 ( .A(u2_u1__abc_74955_new_n299_), .B(u2_u1__abc_74955_new_n298_), .Y(u2_u1__0b2_last_row_12_0__2_));
AND2X2 AND2X2_3002 ( .A(u2_u1__abc_74955_new_n302_), .B(u2_u1__abc_74955_new_n301_), .Y(u2_u1__0b2_last_row_12_0__3_));
AND2X2 AND2X2_3003 ( .A(u2_u1__abc_74955_new_n305_), .B(u2_u1__abc_74955_new_n304_), .Y(u2_u1__0b2_last_row_12_0__4_));
AND2X2 AND2X2_3004 ( .A(u2_u1__abc_74955_new_n308_), .B(u2_u1__abc_74955_new_n307_), .Y(u2_u1__0b2_last_row_12_0__5_));
AND2X2 AND2X2_3005 ( .A(u2_u1__abc_74955_new_n311_), .B(u2_u1__abc_74955_new_n310_), .Y(u2_u1__0b2_last_row_12_0__6_));
AND2X2 AND2X2_3006 ( .A(u2_u1__abc_74955_new_n314_), .B(u2_u1__abc_74955_new_n313_), .Y(u2_u1__0b2_last_row_12_0__7_));
AND2X2 AND2X2_3007 ( .A(u2_u1__abc_74955_new_n317_), .B(u2_u1__abc_74955_new_n316_), .Y(u2_u1__0b2_last_row_12_0__8_));
AND2X2 AND2X2_3008 ( .A(u2_u1__abc_74955_new_n320_), .B(u2_u1__abc_74955_new_n319_), .Y(u2_u1__0b2_last_row_12_0__9_));
AND2X2 AND2X2_3009 ( .A(u2_u1__abc_74955_new_n323_), .B(u2_u1__abc_74955_new_n322_), .Y(u2_u1__0b2_last_row_12_0__10_));
AND2X2 AND2X2_301 ( .A(u0__abc_76628_new_n1523_), .B(u0__abc_76628_new_n1174__bF_buf3), .Y(u0__abc_76628_new_n1524_));
AND2X2 AND2X2_3010 ( .A(u2_u1__abc_74955_new_n326_), .B(u2_u1__abc_74955_new_n325_), .Y(u2_u1__0b2_last_row_12_0__11_));
AND2X2 AND2X2_3011 ( .A(u2_u1__abc_74955_new_n329_), .B(u2_u1__abc_74955_new_n328_), .Y(u2_u1__0b2_last_row_12_0__12_));
AND2X2 AND2X2_3012 ( .A(u2_u1__abc_74955_new_n333_), .B(u2_u1__abc_74955_new_n335_), .Y(u2_u1__abc_74955_new_n336_));
AND2X2 AND2X2_3013 ( .A(u2_u1__abc_74955_new_n336_), .B(u2_u1__abc_74955_new_n331_), .Y(u2_u1__abc_74955_new_n337_));
AND2X2 AND2X2_3014 ( .A(u2_u1__abc_74955_new_n338_), .B(u2_u1__abc_74955_new_n340_), .Y(u2_u1__abc_74955_new_n341_));
AND2X2 AND2X2_3015 ( .A(u2_u1__abc_74955_new_n343_), .B(u2_u1__abc_74955_new_n344_), .Y(u2_u1__abc_74955_new_n345_));
AND2X2 AND2X2_3016 ( .A(u2_u1__abc_74955_new_n341_), .B(u2_u1__abc_74955_new_n345_), .Y(u2_u1__abc_74955_new_n346_));
AND2X2 AND2X2_3017 ( .A(u2_u1__abc_74955_new_n346_), .B(u2_u1__abc_74955_new_n337_), .Y(u2_u1__abc_74955_new_n347_));
AND2X2 AND2X2_3018 ( .A(u2_u1__abc_74955_new_n348_), .B(u2_u1__abc_74955_new_n139_), .Y(u2_u1__abc_74955_new_n349_));
AND2X2 AND2X2_3019 ( .A(u2_u1_b3_last_row_0_), .B(row_adr_0_bF_buf1_), .Y(u2_u1__abc_74955_new_n350_));
AND2X2 AND2X2_302 ( .A(spec_req_cs_3_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1525_));
AND2X2 AND2X2_3020 ( .A(u2_u1__abc_74955_new_n352_), .B(u2_u1__abc_74955_new_n136_), .Y(u2_u1__abc_74955_new_n353_));
AND2X2 AND2X2_3021 ( .A(u2_u1__abc_74955_new_n351_), .B(u2_u1__abc_74955_new_n353_), .Y(u2_u1__abc_74955_new_n354_));
AND2X2 AND2X2_3022 ( .A(u2_u1__abc_74955_new_n356_), .B(u2_u1__abc_74955_new_n357_), .Y(u2_u1__abc_74955_new_n358_));
AND2X2 AND2X2_3023 ( .A(u2_u1__abc_74955_new_n360_), .B(u2_u1__abc_74955_new_n361_), .Y(u2_u1__abc_74955_new_n362_));
AND2X2 AND2X2_3024 ( .A(u2_u1__abc_74955_new_n358_), .B(u2_u1__abc_74955_new_n362_), .Y(u2_u1__abc_74955_new_n363_));
AND2X2 AND2X2_3025 ( .A(u2_u1__abc_74955_new_n363_), .B(u2_u1__abc_74955_new_n354_), .Y(u2_u1__abc_74955_new_n364_));
AND2X2 AND2X2_3026 ( .A(u2_u1__abc_74955_new_n347_), .B(u2_u1__abc_74955_new_n364_), .Y(u2_u1__abc_74955_new_n365_));
AND2X2 AND2X2_3027 ( .A(u2_u1__abc_74955_new_n366_), .B(u2_u1__abc_74955_new_n368_), .Y(u2_u1__abc_74955_new_n369_));
AND2X2 AND2X2_3028 ( .A(u2_u1__abc_74955_new_n370_), .B(u2_u1__abc_74955_new_n372_), .Y(u2_u1__abc_74955_new_n373_));
AND2X2 AND2X2_3029 ( .A(u2_u1__abc_74955_new_n369_), .B(u2_u1__abc_74955_new_n373_), .Y(u2_u1__abc_74955_new_n374_));
AND2X2 AND2X2_303 ( .A(u0__abc_76628_new_n1526_), .B(u0__abc_76628_new_n1173__bF_buf3), .Y(u0__abc_76628_new_n1527_));
AND2X2 AND2X2_3030 ( .A(u2_u1__abc_74955_new_n376_), .B(u2_u1__abc_74955_new_n377_), .Y(u2_u1__abc_74955_new_n378_));
AND2X2 AND2X2_3031 ( .A(u2_u1__abc_74955_new_n380_), .B(u2_u1__abc_74955_new_n381_), .Y(u2_u1__abc_74955_new_n382_));
AND2X2 AND2X2_3032 ( .A(u2_u1__abc_74955_new_n378_), .B(u2_u1__abc_74955_new_n382_), .Y(u2_u1__abc_74955_new_n383_));
AND2X2 AND2X2_3033 ( .A(u2_u1__abc_74955_new_n384_), .B(u2_u1__abc_74955_new_n386_), .Y(u2_u1__abc_74955_new_n387_));
AND2X2 AND2X2_3034 ( .A(u2_u1__abc_74955_new_n389_), .B(u2_u1__abc_74955_new_n390_), .Y(u2_u1__abc_74955_new_n391_));
AND2X2 AND2X2_3035 ( .A(u2_u1__abc_74955_new_n387_), .B(u2_u1__abc_74955_new_n391_), .Y(u2_u1__abc_74955_new_n392_));
AND2X2 AND2X2_3036 ( .A(u2_u1__abc_74955_new_n383_), .B(u2_u1__abc_74955_new_n392_), .Y(u2_u1__abc_74955_new_n393_));
AND2X2 AND2X2_3037 ( .A(u2_u1__abc_74955_new_n393_), .B(u2_u1__abc_74955_new_n374_), .Y(u2_u1__abc_74955_new_n394_));
AND2X2 AND2X2_3038 ( .A(u2_u1__abc_74955_new_n365_), .B(u2_u1__abc_74955_new_n394_), .Y(u2_u1__abc_74955_new_n395_));
AND2X2 AND2X2_3039 ( .A(u2_u1__abc_74955_new_n396_), .B(u2_u1__abc_74955_new_n397_), .Y(u2_u1__abc_74955_new_n398_));
AND2X2 AND2X2_304 ( .A(spec_req_cs_2_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1528_));
AND2X2 AND2X2_3040 ( .A(u2_u1__abc_74955_new_n398_), .B(u2_u1__abc_74955_new_n400_), .Y(u2_u1__abc_74955_new_n401_));
AND2X2 AND2X2_3041 ( .A(u2_u1__abc_74955_new_n402_), .B(u2_u1__abc_74955_new_n404_), .Y(u2_u1__abc_74955_new_n405_));
AND2X2 AND2X2_3042 ( .A(u2_u1__abc_74955_new_n406_), .B(u2_u1__abc_74955_new_n408_), .Y(u2_u1__abc_74955_new_n409_));
AND2X2 AND2X2_3043 ( .A(u2_u1__abc_74955_new_n405_), .B(u2_u1__abc_74955_new_n409_), .Y(u2_u1__abc_74955_new_n410_));
AND2X2 AND2X2_3044 ( .A(u2_u1__abc_74955_new_n410_), .B(u2_u1__abc_74955_new_n401_), .Y(u2_u1__abc_74955_new_n411_));
AND2X2 AND2X2_3045 ( .A(u2_u1__abc_74955_new_n412_), .B(u2_u1__abc_74955_new_n414_), .Y(u2_u1__abc_74955_new_n415_));
AND2X2 AND2X2_3046 ( .A(u2_u1__abc_74955_new_n416_), .B(u2_u1__abc_74955_new_n418_), .Y(u2_u1__abc_74955_new_n419_));
AND2X2 AND2X2_3047 ( .A(u2_u1__abc_74955_new_n415_), .B(u2_u1__abc_74955_new_n419_), .Y(u2_u1__abc_74955_new_n420_));
AND2X2 AND2X2_3048 ( .A(u2_u1__abc_74955_new_n421_), .B(u2_u1__abc_74955_new_n423_), .Y(u2_u1__abc_74955_new_n424_));
AND2X2 AND2X2_3049 ( .A(u2_u1__abc_74955_new_n426_), .B(u2_u1__abc_74955_new_n247_), .Y(u2_u1__abc_74955_new_n427_));
AND2X2 AND2X2_305 ( .A(u0__abc_76628_new_n1529_), .B(u0__abc_76628_new_n1172__bF_buf3), .Y(u0__abc_76628_new_n1530_));
AND2X2 AND2X2_3050 ( .A(u2_u1__abc_74955_new_n424_), .B(u2_u1__abc_74955_new_n427_), .Y(u2_u1__abc_74955_new_n428_));
AND2X2 AND2X2_3051 ( .A(u2_u1__abc_74955_new_n420_), .B(u2_u1__abc_74955_new_n428_), .Y(u2_u1__abc_74955_new_n429_));
AND2X2 AND2X2_3052 ( .A(u2_u1__abc_74955_new_n411_), .B(u2_u1__abc_74955_new_n429_), .Y(u2_u1__abc_74955_new_n430_));
AND2X2 AND2X2_3053 ( .A(u2_u1__abc_74955_new_n432_), .B(u2_u1__abc_74955_new_n433_), .Y(u2_u1__abc_74955_new_n434_));
AND2X2 AND2X2_3054 ( .A(u2_u1__abc_74955_new_n436_), .B(u2_u1__abc_74955_new_n437_), .Y(u2_u1__abc_74955_new_n438_));
AND2X2 AND2X2_3055 ( .A(u2_u1__abc_74955_new_n434_), .B(u2_u1__abc_74955_new_n438_), .Y(u2_u1__abc_74955_new_n439_));
AND2X2 AND2X2_3056 ( .A(u2_u1__abc_74955_new_n441_), .B(u2_u1__abc_74955_new_n442_), .Y(u2_u1__abc_74955_new_n443_));
AND2X2 AND2X2_3057 ( .A(u2_u1__abc_74955_new_n445_), .B(u2_u1__abc_74955_new_n446_), .Y(u2_u1__abc_74955_new_n447_));
AND2X2 AND2X2_3058 ( .A(u2_u1__abc_74955_new_n443_), .B(u2_u1__abc_74955_new_n447_), .Y(u2_u1__abc_74955_new_n448_));
AND2X2 AND2X2_3059 ( .A(u2_u1__abc_74955_new_n449_), .B(u2_u1__abc_74955_new_n451_), .Y(u2_u1__abc_74955_new_n452_));
AND2X2 AND2X2_306 ( .A(spec_req_cs_1_bF_buf0_), .B(u0_tms1_14_), .Y(u0__abc_76628_new_n1531_));
AND2X2 AND2X2_3060 ( .A(u2_u1__abc_74955_new_n453_), .B(u2_u1__abc_74955_new_n455_), .Y(u2_u1__abc_74955_new_n456_));
AND2X2 AND2X2_3061 ( .A(u2_u1__abc_74955_new_n452_), .B(u2_u1__abc_74955_new_n456_), .Y(u2_u1__abc_74955_new_n457_));
AND2X2 AND2X2_3062 ( .A(u2_u1__abc_74955_new_n448_), .B(u2_u1__abc_74955_new_n457_), .Y(u2_u1__abc_74955_new_n458_));
AND2X2 AND2X2_3063 ( .A(u2_u1__abc_74955_new_n458_), .B(u2_u1__abc_74955_new_n439_), .Y(u2_u1__abc_74955_new_n459_));
AND2X2 AND2X2_3064 ( .A(u2_u1__abc_74955_new_n430_), .B(u2_u1__abc_74955_new_n459_), .Y(u2_u1__abc_74955_new_n460_));
AND2X2 AND2X2_3065 ( .A(u2_u1__abc_74955_new_n464_), .B(u2_u1__abc_74955_new_n465_), .Y(u2_u1__abc_74955_new_n466_));
AND2X2 AND2X2_3066 ( .A(u2_u1__abc_74955_new_n466_), .B(u2_u1__abc_74955_new_n463_), .Y(u2_u1__abc_74955_new_n467_));
AND2X2 AND2X2_3067 ( .A(u2_u1__abc_74955_new_n468_), .B(u2_u1__abc_74955_new_n470_), .Y(u2_u1__abc_74955_new_n471_));
AND2X2 AND2X2_3068 ( .A(u2_u1__abc_74955_new_n473_), .B(u2_u1__abc_74955_new_n474_), .Y(u2_u1__abc_74955_new_n475_));
AND2X2 AND2X2_3069 ( .A(u2_u1__abc_74955_new_n471_), .B(u2_u1__abc_74955_new_n475_), .Y(u2_u1__abc_74955_new_n476_));
AND2X2 AND2X2_307 ( .A(u0__abc_76628_new_n1169__bF_buf5), .B(u0__abc_76628_new_n1534_), .Y(u0__abc_76628_new_n1535_));
AND2X2 AND2X2_3070 ( .A(u2_u1__abc_74955_new_n478_), .B(u2_u1__abc_74955_new_n480_), .Y(u2_u1__abc_74955_new_n481_));
AND2X2 AND2X2_3071 ( .A(u2_u1__abc_74955_new_n482_), .B(u2_u1__abc_74955_new_n483_), .Y(u2_u1__abc_74955_new_n484_));
AND2X2 AND2X2_3072 ( .A(u2_u1__abc_74955_new_n481_), .B(u2_u1__abc_74955_new_n484_), .Y(u2_u1__abc_74955_new_n485_));
AND2X2 AND2X2_3073 ( .A(u2_u1__abc_74955_new_n476_), .B(u2_u1__abc_74955_new_n485_), .Y(u2_u1__abc_74955_new_n486_));
AND2X2 AND2X2_3074 ( .A(u2_u1__abc_74955_new_n486_), .B(u2_u1__abc_74955_new_n467_), .Y(u2_u1__abc_74955_new_n487_));
AND2X2 AND2X2_3075 ( .A(u2_u1__abc_74955_new_n139_), .B(u2_u1__abc_74955_new_n488_), .Y(u2_u1__abc_74955_new_n489_));
AND2X2 AND2X2_3076 ( .A(row_adr_0_bF_buf3_), .B(u2_u1_b0_last_row_0_), .Y(u2_u1__abc_74955_new_n490_));
AND2X2 AND2X2_3077 ( .A(u2_u1__abc_74955_new_n493_), .B(u2_u1__abc_74955_new_n494_), .Y(u2_u1__abc_74955_new_n495_));
AND2X2 AND2X2_3078 ( .A(u2_u1__abc_74955_new_n491_), .B(u2_u1__abc_74955_new_n495_), .Y(u2_u1__abc_74955_new_n496_));
AND2X2 AND2X2_3079 ( .A(u2_u1__abc_74955_new_n497_), .B(u2_u1__abc_74955_new_n499_), .Y(u2_u1__abc_74955_new_n500_));
AND2X2 AND2X2_308 ( .A(u0__abc_76628_new_n1533_), .B(u0__abc_76628_new_n1535_), .Y(u0__abc_76628_new_n1536_));
AND2X2 AND2X2_3080 ( .A(u2_u1__abc_74955_new_n502_), .B(u2_u1__abc_74955_new_n205_), .Y(u2_u1__abc_74955_new_n503_));
AND2X2 AND2X2_3081 ( .A(u2_u1__abc_74955_new_n500_), .B(u2_u1__abc_74955_new_n503_), .Y(u2_u1__abc_74955_new_n504_));
AND2X2 AND2X2_3082 ( .A(u2_u1__abc_74955_new_n496_), .B(u2_u1__abc_74955_new_n504_), .Y(u2_u1__abc_74955_new_n505_));
AND2X2 AND2X2_3083 ( .A(u2_u1__abc_74955_new_n507_), .B(u2_u1__abc_74955_new_n509_), .Y(u2_u1__abc_74955_new_n510_));
AND2X2 AND2X2_3084 ( .A(u2_u1__abc_74955_new_n511_), .B(u2_u1__abc_74955_new_n512_), .Y(u2_u1__abc_74955_new_n513_));
AND2X2 AND2X2_3085 ( .A(u2_u1__abc_74955_new_n510_), .B(u2_u1__abc_74955_new_n513_), .Y(u2_u1__abc_74955_new_n514_));
AND2X2 AND2X2_3086 ( .A(u2_u1__abc_74955_new_n515_), .B(u2_u1__abc_74955_new_n517_), .Y(u2_u1__abc_74955_new_n518_));
AND2X2 AND2X2_3087 ( .A(u2_u1__abc_74955_new_n519_), .B(u2_u1__abc_74955_new_n521_), .Y(u2_u1__abc_74955_new_n522_));
AND2X2 AND2X2_3088 ( .A(u2_u1__abc_74955_new_n518_), .B(u2_u1__abc_74955_new_n522_), .Y(u2_u1__abc_74955_new_n523_));
AND2X2 AND2X2_3089 ( .A(u2_u1__abc_74955_new_n514_), .B(u2_u1__abc_74955_new_n523_), .Y(u2_u1__abc_74955_new_n524_));
AND2X2 AND2X2_309 ( .A(u0__abc_76628_new_n1170__bF_buf5), .B(sp_tms_15_), .Y(u0__abc_76628_new_n1538_));
AND2X2 AND2X2_3090 ( .A(u2_u1__abc_74955_new_n524_), .B(u2_u1__abc_74955_new_n505_), .Y(u2_u1__abc_74955_new_n525_));
AND2X2 AND2X2_3091 ( .A(u2_u1__abc_74955_new_n487_), .B(u2_u1__abc_74955_new_n525_), .Y(u2_u1__abc_74955_new_n526_));
AND2X2 AND2X2_3092 ( .A(u2_u1__abc_74955_new_n529_), .B(u2_u1__abc_74955_new_n530_), .Y(u2_u1__abc_74955_new_n531_));
AND2X2 AND2X2_3093 ( .A(u2_u1__abc_74955_new_n531_), .B(u2_u1__abc_74955_new_n528_), .Y(u2_u1__abc_74955_new_n532_));
AND2X2 AND2X2_3094 ( .A(u2_u1__abc_74955_new_n534_), .B(u2_u1__abc_74955_new_n535_), .Y(u2_u1__abc_74955_new_n536_));
AND2X2 AND2X2_3095 ( .A(u2_u1__abc_74955_new_n538_), .B(u2_u1__abc_74955_new_n539_), .Y(u2_u1__abc_74955_new_n540_));
AND2X2 AND2X2_3096 ( .A(u2_u1__abc_74955_new_n536_), .B(u2_u1__abc_74955_new_n540_), .Y(u2_u1__abc_74955_new_n541_));
AND2X2 AND2X2_3097 ( .A(u2_u1__abc_74955_new_n541_), .B(u2_u1__abc_74955_new_n532_), .Y(u2_u1__abc_74955_new_n542_));
AND2X2 AND2X2_3098 ( .A(u2_u1__abc_74955_new_n543_), .B(u2_u1__abc_74955_new_n545_), .Y(u2_u1__abc_74955_new_n546_));
AND2X2 AND2X2_3099 ( .A(u2_u1__abc_74955_new_n547_), .B(u2_u1__abc_74955_new_n549_), .Y(u2_u1__abc_74955_new_n550_));
AND2X2 AND2X2_31 ( .A(_abc_85006_new_n329_), .B(_abc_85006_new_n330_), .Y(tms_s_13_));
AND2X2 AND2X2_310 ( .A(spec_req_cs_5_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1539_));
AND2X2 AND2X2_3100 ( .A(u2_u1__abc_74955_new_n546_), .B(u2_u1__abc_74955_new_n550_), .Y(u2_u1__abc_74955_new_n551_));
AND2X2 AND2X2_3101 ( .A(u2_u1__abc_74955_new_n552_), .B(u2_u1__abc_74955_new_n554_), .Y(u2_u1__abc_74955_new_n555_));
AND2X2 AND2X2_3102 ( .A(u2_u1__abc_74955_new_n556_), .B(u2_u1__abc_74955_new_n558_), .Y(u2_u1__abc_74955_new_n559_));
AND2X2 AND2X2_3103 ( .A(u2_u1__abc_74955_new_n555_), .B(u2_u1__abc_74955_new_n559_), .Y(u2_u1__abc_74955_new_n560_));
AND2X2 AND2X2_3104 ( .A(u2_u1__abc_74955_new_n551_), .B(u2_u1__abc_74955_new_n560_), .Y(u2_u1__abc_74955_new_n561_));
AND2X2 AND2X2_3105 ( .A(u2_u1__abc_74955_new_n561_), .B(u2_u1__abc_74955_new_n542_), .Y(u2_u1__abc_74955_new_n562_));
AND2X2 AND2X2_3106 ( .A(u2_u1__abc_74955_new_n564_), .B(u2_u1__abc_74955_new_n565_), .Y(u2_u1__abc_74955_new_n566_));
AND2X2 AND2X2_3107 ( .A(u2_u1__abc_74955_new_n568_), .B(u2_u1__abc_74955_new_n569_), .Y(u2_u1__abc_74955_new_n570_));
AND2X2 AND2X2_3108 ( .A(u2_u1__abc_74955_new_n566_), .B(u2_u1__abc_74955_new_n570_), .Y(u2_u1__abc_74955_new_n571_));
AND2X2 AND2X2_3109 ( .A(u2_u1__abc_74955_new_n572_), .B(u2_u1__abc_74955_new_n574_), .Y(u2_u1__abc_74955_new_n575_));
AND2X2 AND2X2_311 ( .A(u0__abc_76628_new_n1541_), .B(u0__abc_76628_new_n1179__bF_buf2), .Y(u0__abc_76628_new_n1542_));
AND2X2 AND2X2_3110 ( .A(u2_u1__abc_74955_new_n576_), .B(u2_u1__abc_74955_new_n578_), .Y(u2_u1__abc_74955_new_n579_));
AND2X2 AND2X2_3111 ( .A(u2_u1__abc_74955_new_n575_), .B(u2_u1__abc_74955_new_n579_), .Y(u2_u1__abc_74955_new_n580_));
AND2X2 AND2X2_3112 ( .A(u2_u1__abc_74955_new_n581_), .B(u2_u1__abc_74955_new_n583_), .Y(u2_u1__abc_74955_new_n584_));
AND2X2 AND2X2_3113 ( .A(u2_u1__abc_74955_new_n586_), .B(u2_u1__abc_74955_new_n289_), .Y(u2_u1__abc_74955_new_n587_));
AND2X2 AND2X2_3114 ( .A(u2_u1__abc_74955_new_n584_), .B(u2_u1__abc_74955_new_n587_), .Y(u2_u1__abc_74955_new_n588_));
AND2X2 AND2X2_3115 ( .A(u2_u1__abc_74955_new_n580_), .B(u2_u1__abc_74955_new_n588_), .Y(u2_u1__abc_74955_new_n589_));
AND2X2 AND2X2_3116 ( .A(u2_u1__abc_74955_new_n589_), .B(u2_u1__abc_74955_new_n571_), .Y(u2_u1__abc_74955_new_n590_));
AND2X2 AND2X2_3117 ( .A(u2_u1__abc_74955_new_n562_), .B(u2_u1__abc_74955_new_n590_), .Y(u2_u1__abc_74955_new_n591_));
AND2X2 AND2X2_3118 ( .A(u2_u1__abc_74955_new_n289_), .B(u2_u1_bank2_open), .Y(u2_u1__abc_74955_new_n594_));
AND2X2 AND2X2_3119 ( .A(u2_u1__abc_74955_new_n136_), .B(u2_u1_bank3_open), .Y(u2_u1__abc_74955_new_n595_));
AND2X2 AND2X2_312 ( .A(u0__abc_76628_new_n1542_), .B(u0__abc_76628_new_n1540_), .Y(u0__abc_76628_new_n1543_));
AND2X2 AND2X2_3120 ( .A(u2_u1__abc_74955_new_n205_), .B(u2_u1_bank0_open), .Y(u2_u1__abc_74955_new_n597_));
AND2X2 AND2X2_3121 ( .A(u2_u1__abc_74955_new_n247_), .B(u2_u1_bank1_open), .Y(u2_u1__abc_74955_new_n598_));
AND2X2 AND2X2_3122 ( .A(u2_u1__abc_74955_new_n604_), .B(u2_u1_bank2_open), .Y(u2_u1__abc_74955_new_n605_));
AND2X2 AND2X2_3123 ( .A(u2_u1__abc_74955_new_n603_), .B(u2_u1__abc_74955_new_n605_), .Y(u2_u1__abc_74955_new_n606_));
AND2X2 AND2X2_3124 ( .A(u2_u1__abc_74955_new_n136_), .B(u2_bank_clr_1), .Y(u2_u1__abc_74955_new_n608_));
AND2X2 AND2X2_3125 ( .A(u2_u1__abc_74955_new_n604_), .B(u2_u1_bank3_open), .Y(u2_u1__abc_74955_new_n610_));
AND2X2 AND2X2_3126 ( .A(u2_u1__abc_74955_new_n609_), .B(u2_u1__abc_74955_new_n610_), .Y(u2_u1__abc_74955_new_n611_));
AND2X2 AND2X2_3127 ( .A(u2_u1__abc_74955_new_n604_), .B(u2_u1_bank1_open), .Y(u2_u1__abc_74955_new_n618_));
AND2X2 AND2X2_3128 ( .A(u2_u1__abc_74955_new_n617_), .B(u2_u1__abc_74955_new_n618_), .Y(u2_u1__abc_74955_new_n619_));
AND2X2 AND2X2_3129 ( .A(u2_u1__abc_74955_new_n604_), .B(u2_u1_bank0_open), .Y(u2_u1__abc_74955_new_n623_));
AND2X2 AND2X2_313 ( .A(u0__abc_76628_new_n1544_), .B(u0__abc_76628_new_n1175__bF_buf2), .Y(u0__abc_76628_new_n1545_));
AND2X2 AND2X2_3130 ( .A(u2_u1__abc_74955_new_n622_), .B(u2_u1__abc_74955_new_n623_), .Y(u2_u1__abc_74955_new_n624_));
AND2X2 AND2X2_3131 ( .A(\wb_data_i[3] ), .B(\wb_data_i[2] ), .Y(u3__abc_74070_new_n281_));
AND2X2 AND2X2_3132 ( .A(u3__abc_74070_new_n282_), .B(u3__abc_74070_new_n280_), .Y(u3__abc_74070_new_n283_));
AND2X2 AND2X2_3133 ( .A(u3__abc_74070_new_n286_), .B(u3__abc_74070_new_n288_), .Y(u3__abc_74070_new_n289_));
AND2X2 AND2X2_3134 ( .A(u3__abc_74070_new_n284_), .B(u3__abc_74070_new_n289_), .Y(u3__abc_74070_new_n290_));
AND2X2 AND2X2_3135 ( .A(u3__abc_74070_new_n291_), .B(u3__abc_74070_new_n292_), .Y(u3__abc_74070_new_n293_));
AND2X2 AND2X2_3136 ( .A(\wb_data_i[7] ), .B(\wb_data_i[6] ), .Y(u3__abc_74070_new_n296_));
AND2X2 AND2X2_3137 ( .A(u3__abc_74070_new_n297_), .B(u3__abc_74070_new_n295_), .Y(u3__abc_74070_new_n298_));
AND2X2 AND2X2_3138 ( .A(u3__abc_74070_new_n301_), .B(u3__abc_74070_new_n303_), .Y(u3__abc_74070_new_n304_));
AND2X2 AND2X2_3139 ( .A(u3__abc_74070_new_n305_), .B(u3__abc_74070_new_n299_), .Y(u3__abc_74070_new_n306_));
AND2X2 AND2X2_314 ( .A(spec_req_cs_4_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1546_));
AND2X2 AND2X2_3140 ( .A(u3__abc_74070_new_n304_), .B(u3__abc_74070_new_n298_), .Y(u3__abc_74070_new_n307_));
AND2X2 AND2X2_3141 ( .A(u3__abc_74070_new_n310_), .B(u3__abc_74070_new_n311_), .Y(u3__abc_74070_new_n312_));
AND2X2 AND2X2_3142 ( .A(u3__abc_74070_new_n313_), .B(u3__abc_74070_new_n278_), .Y(u3__0mc_dp_o_3_0__0_));
AND2X2 AND2X2_3143 ( .A(\wb_data_i[11] ), .B(\wb_data_i[10] ), .Y(u3__abc_74070_new_n317_));
AND2X2 AND2X2_3144 ( .A(u3__abc_74070_new_n318_), .B(u3__abc_74070_new_n316_), .Y(u3__abc_74070_new_n319_));
AND2X2 AND2X2_3145 ( .A(u3__abc_74070_new_n321_), .B(u3__abc_74070_new_n323_), .Y(u3__abc_74070_new_n324_));
AND2X2 AND2X2_3146 ( .A(u3__abc_74070_new_n325_), .B(u3__abc_74070_new_n319_), .Y(u3__abc_74070_new_n326_));
AND2X2 AND2X2_3147 ( .A(u3__abc_74070_new_n327_), .B(u3__abc_74070_new_n328_), .Y(u3__abc_74070_new_n329_));
AND2X2 AND2X2_3148 ( .A(\wb_data_i[15] ), .B(\wb_data_i[14] ), .Y(u3__abc_74070_new_n332_));
AND2X2 AND2X2_3149 ( .A(u3__abc_74070_new_n333_), .B(u3__abc_74070_new_n331_), .Y(u3__abc_74070_new_n334_));
AND2X2 AND2X2_315 ( .A(u0__abc_76628_new_n1547_), .B(u0__abc_76628_new_n1174__bF_buf2), .Y(u0__abc_76628_new_n1548_));
AND2X2 AND2X2_3150 ( .A(u3__abc_74070_new_n337_), .B(u3__abc_74070_new_n339_), .Y(u3__abc_74070_new_n340_));
AND2X2 AND2X2_3151 ( .A(u3__abc_74070_new_n341_), .B(u3__abc_74070_new_n335_), .Y(u3__abc_74070_new_n342_));
AND2X2 AND2X2_3152 ( .A(u3__abc_74070_new_n340_), .B(u3__abc_74070_new_n334_), .Y(u3__abc_74070_new_n343_));
AND2X2 AND2X2_3153 ( .A(u3__abc_74070_new_n346_), .B(u3__abc_74070_new_n347_), .Y(u3__abc_74070_new_n348_));
AND2X2 AND2X2_3154 ( .A(u3__abc_74070_new_n349_), .B(u3__abc_74070_new_n315_), .Y(u3__0mc_dp_o_3_0__1_));
AND2X2 AND2X2_3155 ( .A(\wb_data_i[19] ), .B(\wb_data_i[18] ), .Y(u3__abc_74070_new_n352_));
AND2X2 AND2X2_3156 ( .A(u3__abc_74070_new_n353_), .B(u3__abc_74070_new_n351_), .Y(u3__abc_74070_new_n354_));
AND2X2 AND2X2_3157 ( .A(u3__abc_74070_new_n356_), .B(u3__abc_74070_new_n358_), .Y(u3__abc_74070_new_n359_));
AND2X2 AND2X2_3158 ( .A(u3__abc_74070_new_n360_), .B(u3__abc_74070_new_n354_), .Y(u3__abc_74070_new_n361_));
AND2X2 AND2X2_3159 ( .A(u3__abc_74070_new_n362_), .B(u3__abc_74070_new_n363_), .Y(u3__abc_74070_new_n364_));
AND2X2 AND2X2_316 ( .A(spec_req_cs_3_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1549_));
AND2X2 AND2X2_3160 ( .A(\wb_data_i[23] ), .B(\wb_data_i[22] ), .Y(u3__abc_74070_new_n366_));
AND2X2 AND2X2_3161 ( .A(u3__abc_74070_new_n367_), .B(u3__abc_74070_new_n365_), .Y(u3__abc_74070_new_n368_));
AND2X2 AND2X2_3162 ( .A(u3__abc_74070_new_n371_), .B(u3__abc_74070_new_n373_), .Y(u3__abc_74070_new_n374_));
AND2X2 AND2X2_3163 ( .A(u3__abc_74070_new_n375_), .B(u3__abc_74070_new_n369_), .Y(u3__abc_74070_new_n376_));
AND2X2 AND2X2_3164 ( .A(u3__abc_74070_new_n374_), .B(u3__abc_74070_new_n368_), .Y(u3__abc_74070_new_n377_));
AND2X2 AND2X2_3165 ( .A(u3__abc_74070_new_n379_), .B(u3__abc_74070_new_n364_), .Y(u3__abc_74070_new_n380_));
AND2X2 AND2X2_3166 ( .A(u3__abc_74070_new_n381_), .B(u3__abc_74070_new_n378_), .Y(u3__abc_74070_new_n382_));
AND2X2 AND2X2_3167 ( .A(u3__abc_74070_new_n383_), .B(u3__abc_74070_new_n277__bF_buf2), .Y(u3__abc_74070_new_n384_));
AND2X2 AND2X2_3168 ( .A(u3__abc_74070_new_n279__bF_buf3), .B(mc_dp_od_2_), .Y(u3__abc_74070_new_n385_));
AND2X2 AND2X2_3169 ( .A(\wb_data_i[27] ), .B(\wb_data_i[26] ), .Y(u3__abc_74070_new_n388_));
AND2X2 AND2X2_317 ( .A(u0__abc_76628_new_n1550_), .B(u0__abc_76628_new_n1173__bF_buf2), .Y(u0__abc_76628_new_n1551_));
AND2X2 AND2X2_3170 ( .A(u3__abc_74070_new_n389_), .B(u3__abc_74070_new_n387_), .Y(u3__abc_74070_new_n390_));
AND2X2 AND2X2_3171 ( .A(u3__abc_74070_new_n392_), .B(u3__abc_74070_new_n394_), .Y(u3__abc_74070_new_n395_));
AND2X2 AND2X2_3172 ( .A(u3__abc_74070_new_n396_), .B(u3__abc_74070_new_n390_), .Y(u3__abc_74070_new_n397_));
AND2X2 AND2X2_3173 ( .A(u3__abc_74070_new_n398_), .B(u3__abc_74070_new_n399_), .Y(u3__abc_74070_new_n400_));
AND2X2 AND2X2_3174 ( .A(\wb_data_i[31] ), .B(\wb_data_i[30] ), .Y(u3__abc_74070_new_n402_));
AND2X2 AND2X2_3175 ( .A(u3__abc_74070_new_n403_), .B(u3__abc_74070_new_n401_), .Y(u3__abc_74070_new_n404_));
AND2X2 AND2X2_3176 ( .A(u3__abc_74070_new_n407_), .B(u3__abc_74070_new_n409_), .Y(u3__abc_74070_new_n410_));
AND2X2 AND2X2_3177 ( .A(u3__abc_74070_new_n411_), .B(u3__abc_74070_new_n405_), .Y(u3__abc_74070_new_n412_));
AND2X2 AND2X2_3178 ( .A(u3__abc_74070_new_n410_), .B(u3__abc_74070_new_n404_), .Y(u3__abc_74070_new_n413_));
AND2X2 AND2X2_3179 ( .A(u3__abc_74070_new_n415_), .B(u3__abc_74070_new_n400_), .Y(u3__abc_74070_new_n416_));
AND2X2 AND2X2_318 ( .A(spec_req_cs_2_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1552_));
AND2X2 AND2X2_3180 ( .A(u3__abc_74070_new_n417_), .B(u3__abc_74070_new_n414_), .Y(u3__abc_74070_new_n418_));
AND2X2 AND2X2_3181 ( .A(u3__abc_74070_new_n419_), .B(u3__abc_74070_new_n277__bF_buf1), .Y(u3__abc_74070_new_n420_));
AND2X2 AND2X2_3182 ( .A(u3__abc_74070_new_n279__bF_buf2), .B(mc_dp_od_3_), .Y(u3__abc_74070_new_n421_));
AND2X2 AND2X2_3183 ( .A(u3__abc_74070_new_n425_), .B(u3__abc_74070_new_n423_), .Y(u3__0byte2_7_0__0_));
AND2X2 AND2X2_3184 ( .A(u3__abc_74070_new_n428_), .B(u3__abc_74070_new_n427_), .Y(u3__0byte2_7_0__1_));
AND2X2 AND2X2_3185 ( .A(u3__abc_74070_new_n431_), .B(u3__abc_74070_new_n430_), .Y(u3__0byte2_7_0__2_));
AND2X2 AND2X2_3186 ( .A(u3__abc_74070_new_n434_), .B(u3__abc_74070_new_n433_), .Y(u3__0byte2_7_0__3_));
AND2X2 AND2X2_3187 ( .A(u3__abc_74070_new_n437_), .B(u3__abc_74070_new_n436_), .Y(u3__0byte2_7_0__4_));
AND2X2 AND2X2_3188 ( .A(u3__abc_74070_new_n440_), .B(u3__abc_74070_new_n439_), .Y(u3__0byte2_7_0__5_));
AND2X2 AND2X2_3189 ( .A(u3__abc_74070_new_n443_), .B(u3__abc_74070_new_n442_), .Y(u3__0byte2_7_0__6_));
AND2X2 AND2X2_319 ( .A(u0__abc_76628_new_n1553_), .B(u0__abc_76628_new_n1172__bF_buf2), .Y(u0__abc_76628_new_n1554_));
AND2X2 AND2X2_3190 ( .A(u3__abc_74070_new_n446_), .B(u3__abc_74070_new_n445_), .Y(u3__0byte2_7_0__7_));
AND2X2 AND2X2_3191 ( .A(u3__abc_74070_new_n448_), .B(u3__abc_74070_new_n449__bF_buf3), .Y(u3__abc_74070_new_n450_));
AND2X2 AND2X2_3192 ( .A(u3__abc_74070_new_n450__bF_buf3), .B(pack_le1), .Y(u3__abc_74070_new_n451_));
AND2X2 AND2X2_3193 ( .A(u3__abc_74070_new_n449__bF_buf2), .B(csc_4_), .Y(u3__abc_74070_new_n452_));
AND2X2 AND2X2_3194 ( .A(u3__abc_74070_new_n452__bF_buf3), .B(pack_le0), .Y(u3__abc_74070_new_n453_));
AND2X2 AND2X2_3195 ( .A(u3__abc_74070_new_n455_), .B(u3__abc_74070_new_n456_), .Y(u3__abc_74070_new_n457_));
AND2X2 AND2X2_3196 ( .A(u3__abc_74070_new_n458_), .B(u3__abc_74070_new_n460_), .Y(u3__0byte1_7_0__0_));
AND2X2 AND2X2_3197 ( .A(u3__abc_74070_new_n462_), .B(u3__abc_74070_new_n463_), .Y(u3__abc_74070_new_n464_));
AND2X2 AND2X2_3198 ( .A(u3__abc_74070_new_n465_), .B(u3__abc_74070_new_n466_), .Y(u3__0byte1_7_0__1_));
AND2X2 AND2X2_3199 ( .A(u3__abc_74070_new_n468_), .B(u3__abc_74070_new_n469_), .Y(u3__abc_74070_new_n470_));
AND2X2 AND2X2_32 ( .A(_abc_85006_new_n332_), .B(_abc_85006_new_n333_), .Y(tms_s_14_));
AND2X2 AND2X2_320 ( .A(spec_req_cs_1_bF_buf5_), .B(u0_tms1_15_), .Y(u0__abc_76628_new_n1555_));
AND2X2 AND2X2_3200 ( .A(u3__abc_74070_new_n471_), .B(u3__abc_74070_new_n472_), .Y(u3__0byte1_7_0__2_));
AND2X2 AND2X2_3201 ( .A(u3__abc_74070_new_n474_), .B(u3__abc_74070_new_n475_), .Y(u3__abc_74070_new_n476_));
AND2X2 AND2X2_3202 ( .A(u3__abc_74070_new_n477_), .B(u3__abc_74070_new_n478_), .Y(u3__0byte1_7_0__3_));
AND2X2 AND2X2_3203 ( .A(u3__abc_74070_new_n480_), .B(u3__abc_74070_new_n481_), .Y(u3__abc_74070_new_n482_));
AND2X2 AND2X2_3204 ( .A(u3__abc_74070_new_n483_), .B(u3__abc_74070_new_n484_), .Y(u3__0byte1_7_0__4_));
AND2X2 AND2X2_3205 ( .A(u3__abc_74070_new_n486_), .B(u3__abc_74070_new_n487_), .Y(u3__abc_74070_new_n488_));
AND2X2 AND2X2_3206 ( .A(u3__abc_74070_new_n489_), .B(u3__abc_74070_new_n490_), .Y(u3__0byte1_7_0__5_));
AND2X2 AND2X2_3207 ( .A(u3__abc_74070_new_n492_), .B(u3__abc_74070_new_n493_), .Y(u3__abc_74070_new_n494_));
AND2X2 AND2X2_3208 ( .A(u3__abc_74070_new_n495_), .B(u3__abc_74070_new_n496_), .Y(u3__0byte1_7_0__6_));
AND2X2 AND2X2_3209 ( .A(u3__abc_74070_new_n498_), .B(u3__abc_74070_new_n499_), .Y(u3__abc_74070_new_n500_));
AND2X2 AND2X2_321 ( .A(u0__abc_76628_new_n1169__bF_buf4), .B(u0__abc_76628_new_n1558_), .Y(u0__abc_76628_new_n1559_));
AND2X2 AND2X2_3210 ( .A(u3__abc_74070_new_n501_), .B(u3__abc_74070_new_n502_), .Y(u3__0byte1_7_0__7_));
AND2X2 AND2X2_3211 ( .A(u3__abc_74070_new_n506_), .B(u3__abc_74070_new_n504_), .Y(u3__0byte0_7_0__0_));
AND2X2 AND2X2_3212 ( .A(u3__abc_74070_new_n509_), .B(u3__abc_74070_new_n508_), .Y(u3__0byte0_7_0__1_));
AND2X2 AND2X2_3213 ( .A(u3__abc_74070_new_n512_), .B(u3__abc_74070_new_n511_), .Y(u3__0byte0_7_0__2_));
AND2X2 AND2X2_3214 ( .A(u3__abc_74070_new_n515_), .B(u3__abc_74070_new_n514_), .Y(u3__0byte0_7_0__3_));
AND2X2 AND2X2_3215 ( .A(u3__abc_74070_new_n518_), .B(u3__abc_74070_new_n517_), .Y(u3__0byte0_7_0__4_));
AND2X2 AND2X2_3216 ( .A(u3__abc_74070_new_n521_), .B(u3__abc_74070_new_n520_), .Y(u3__0byte0_7_0__5_));
AND2X2 AND2X2_3217 ( .A(u3__abc_74070_new_n524_), .B(u3__abc_74070_new_n523_), .Y(u3__0byte0_7_0__6_));
AND2X2 AND2X2_3218 ( .A(u3__abc_74070_new_n527_), .B(u3__abc_74070_new_n526_), .Y(u3__0byte0_7_0__7_));
AND2X2 AND2X2_3219 ( .A(u3__abc_74070_new_n529_), .B(u3__abc_74070_new_n530_), .Y(u3__0mc_data_o_31_0__0_));
AND2X2 AND2X2_322 ( .A(u0__abc_76628_new_n1557_), .B(u0__abc_76628_new_n1559_), .Y(u0__abc_76628_new_n1560_));
AND2X2 AND2X2_3220 ( .A(u3__abc_74070_new_n532_), .B(u3__abc_74070_new_n533_), .Y(u3__0mc_data_o_31_0__1_));
AND2X2 AND2X2_3221 ( .A(u3__abc_74070_new_n535_), .B(u3__abc_74070_new_n536_), .Y(u3__0mc_data_o_31_0__2_));
AND2X2 AND2X2_3222 ( .A(u3__abc_74070_new_n538_), .B(u3__abc_74070_new_n539_), .Y(u3__0mc_data_o_31_0__3_));
AND2X2 AND2X2_3223 ( .A(u3__abc_74070_new_n541_), .B(u3__abc_74070_new_n542_), .Y(u3__0mc_data_o_31_0__4_));
AND2X2 AND2X2_3224 ( .A(u3__abc_74070_new_n544_), .B(u3__abc_74070_new_n545_), .Y(u3__0mc_data_o_31_0__5_));
AND2X2 AND2X2_3225 ( .A(u3__abc_74070_new_n547_), .B(u3__abc_74070_new_n548_), .Y(u3__0mc_data_o_31_0__6_));
AND2X2 AND2X2_3226 ( .A(u3__abc_74070_new_n550_), .B(u3__abc_74070_new_n551_), .Y(u3__0mc_data_o_31_0__7_));
AND2X2 AND2X2_3227 ( .A(u3__abc_74070_new_n553_), .B(u3__abc_74070_new_n554_), .Y(u3__0mc_data_o_31_0__8_));
AND2X2 AND2X2_3228 ( .A(u3__abc_74070_new_n556_), .B(u3__abc_74070_new_n557_), .Y(u3__0mc_data_o_31_0__9_));
AND2X2 AND2X2_3229 ( .A(u3__abc_74070_new_n559_), .B(u3__abc_74070_new_n560_), .Y(u3__0mc_data_o_31_0__10_));
AND2X2 AND2X2_323 ( .A(u0__abc_76628_new_n1170__bF_buf4), .B(sp_tms_16_), .Y(u0__abc_76628_new_n1562_));
AND2X2 AND2X2_3230 ( .A(u3__abc_74070_new_n562_), .B(u3__abc_74070_new_n563_), .Y(u3__0mc_data_o_31_0__11_));
AND2X2 AND2X2_3231 ( .A(u3__abc_74070_new_n565_), .B(u3__abc_74070_new_n566_), .Y(u3__0mc_data_o_31_0__12_));
AND2X2 AND2X2_3232 ( .A(u3__abc_74070_new_n568_), .B(u3__abc_74070_new_n569_), .Y(u3__0mc_data_o_31_0__13_));
AND2X2 AND2X2_3233 ( .A(u3__abc_74070_new_n571_), .B(u3__abc_74070_new_n572_), .Y(u3__0mc_data_o_31_0__14_));
AND2X2 AND2X2_3234 ( .A(u3__abc_74070_new_n574_), .B(u3__abc_74070_new_n575_), .Y(u3__0mc_data_o_31_0__15_));
AND2X2 AND2X2_3235 ( .A(u3__abc_74070_new_n577_), .B(u3__abc_74070_new_n578_), .Y(u3__0mc_data_o_31_0__16_));
AND2X2 AND2X2_3236 ( .A(u3__abc_74070_new_n580_), .B(u3__abc_74070_new_n581_), .Y(u3__0mc_data_o_31_0__17_));
AND2X2 AND2X2_3237 ( .A(u3__abc_74070_new_n583_), .B(u3__abc_74070_new_n584_), .Y(u3__0mc_data_o_31_0__18_));
AND2X2 AND2X2_3238 ( .A(u3__abc_74070_new_n586_), .B(u3__abc_74070_new_n587_), .Y(u3__0mc_data_o_31_0__19_));
AND2X2 AND2X2_3239 ( .A(u3__abc_74070_new_n589_), .B(u3__abc_74070_new_n590_), .Y(u3__0mc_data_o_31_0__20_));
AND2X2 AND2X2_324 ( .A(spec_req_cs_5_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1563_));
AND2X2 AND2X2_3240 ( .A(u3__abc_74070_new_n592_), .B(u3__abc_74070_new_n593_), .Y(u3__0mc_data_o_31_0__21_));
AND2X2 AND2X2_3241 ( .A(u3__abc_74070_new_n595_), .B(u3__abc_74070_new_n596_), .Y(u3__0mc_data_o_31_0__22_));
AND2X2 AND2X2_3242 ( .A(u3__abc_74070_new_n598_), .B(u3__abc_74070_new_n599_), .Y(u3__0mc_data_o_31_0__23_));
AND2X2 AND2X2_3243 ( .A(u3__abc_74070_new_n601_), .B(u3__abc_74070_new_n602_), .Y(u3__0mc_data_o_31_0__24_));
AND2X2 AND2X2_3244 ( .A(u3__abc_74070_new_n604_), .B(u3__abc_74070_new_n605_), .Y(u3__0mc_data_o_31_0__25_));
AND2X2 AND2X2_3245 ( .A(u3__abc_74070_new_n607_), .B(u3__abc_74070_new_n608_), .Y(u3__0mc_data_o_31_0__26_));
AND2X2 AND2X2_3246 ( .A(u3__abc_74070_new_n610_), .B(u3__abc_74070_new_n611_), .Y(u3__0mc_data_o_31_0__27_));
AND2X2 AND2X2_3247 ( .A(u3__abc_74070_new_n613_), .B(u3__abc_74070_new_n614_), .Y(u3__0mc_data_o_31_0__28_));
AND2X2 AND2X2_3248 ( .A(u3__abc_74070_new_n616_), .B(u3__abc_74070_new_n617_), .Y(u3__0mc_data_o_31_0__29_));
AND2X2 AND2X2_3249 ( .A(u3__abc_74070_new_n619_), .B(u3__abc_74070_new_n620_), .Y(u3__0mc_data_o_31_0__30_));
AND2X2 AND2X2_325 ( .A(u0__abc_76628_new_n1565_), .B(u0__abc_76628_new_n1179__bF_buf1), .Y(u0__abc_76628_new_n1566_));
AND2X2 AND2X2_3250 ( .A(u3__abc_74070_new_n622_), .B(u3__abc_74070_new_n623_), .Y(u3__0mc_data_o_31_0__31_));
AND2X2 AND2X2_3251 ( .A(u3__abc_74070_new_n627_), .B(u3__abc_74070_new_n626_), .Y(u3__abc_74070_new_n628_));
AND2X2 AND2X2_3252 ( .A(u3__abc_74070_new_n629_), .B(u3__abc_74070_new_n630_), .Y(mem_dout_0_));
AND2X2 AND2X2_3253 ( .A(u3__abc_74070_new_n633_), .B(u3__abc_74070_new_n632_), .Y(u3__abc_74070_new_n634_));
AND2X2 AND2X2_3254 ( .A(u3__abc_74070_new_n635_), .B(u3__abc_74070_new_n636_), .Y(mem_dout_1_));
AND2X2 AND2X2_3255 ( .A(u3__abc_74070_new_n639_), .B(u3__abc_74070_new_n638_), .Y(u3__abc_74070_new_n640_));
AND2X2 AND2X2_3256 ( .A(u3__abc_74070_new_n641_), .B(u3__abc_74070_new_n642_), .Y(mem_dout_2_));
AND2X2 AND2X2_3257 ( .A(u3__abc_74070_new_n645_), .B(u3__abc_74070_new_n644_), .Y(u3__abc_74070_new_n646_));
AND2X2 AND2X2_3258 ( .A(u3__abc_74070_new_n647_), .B(u3__abc_74070_new_n648_), .Y(mem_dout_3_));
AND2X2 AND2X2_3259 ( .A(u3__abc_74070_new_n651_), .B(u3__abc_74070_new_n650_), .Y(u3__abc_74070_new_n652_));
AND2X2 AND2X2_326 ( .A(u0__abc_76628_new_n1566_), .B(u0__abc_76628_new_n1564_), .Y(u0__abc_76628_new_n1567_));
AND2X2 AND2X2_3260 ( .A(u3__abc_74070_new_n653_), .B(u3__abc_74070_new_n654_), .Y(mem_dout_4_));
AND2X2 AND2X2_3261 ( .A(u3__abc_74070_new_n657_), .B(u3__abc_74070_new_n656_), .Y(u3__abc_74070_new_n658_));
AND2X2 AND2X2_3262 ( .A(u3__abc_74070_new_n659_), .B(u3__abc_74070_new_n660_), .Y(mem_dout_5_));
AND2X2 AND2X2_3263 ( .A(u3__abc_74070_new_n663_), .B(u3__abc_74070_new_n662_), .Y(u3__abc_74070_new_n664_));
AND2X2 AND2X2_3264 ( .A(u3__abc_74070_new_n665_), .B(u3__abc_74070_new_n666_), .Y(mem_dout_6_));
AND2X2 AND2X2_3265 ( .A(u3__abc_74070_new_n669_), .B(u3__abc_74070_new_n668_), .Y(u3__abc_74070_new_n670_));
AND2X2 AND2X2_3266 ( .A(u3__abc_74070_new_n671_), .B(u3__abc_74070_new_n672_), .Y(mem_dout_7_));
AND2X2 AND2X2_3267 ( .A(u3__abc_74070_new_n675_), .B(u3__abc_74070_new_n674_), .Y(u3__abc_74070_new_n676_));
AND2X2 AND2X2_3268 ( .A(u3__abc_74070_new_n677_), .B(u3__abc_74070_new_n678_), .Y(mem_dout_8_));
AND2X2 AND2X2_3269 ( .A(u3__abc_74070_new_n681_), .B(u3__abc_74070_new_n680_), .Y(u3__abc_74070_new_n682_));
AND2X2 AND2X2_327 ( .A(u0__abc_76628_new_n1568_), .B(u0__abc_76628_new_n1175__bF_buf1), .Y(u0__abc_76628_new_n1569_));
AND2X2 AND2X2_3270 ( .A(u3__abc_74070_new_n683_), .B(u3__abc_74070_new_n684_), .Y(mem_dout_9_));
AND2X2 AND2X2_3271 ( .A(u3__abc_74070_new_n687_), .B(u3__abc_74070_new_n686_), .Y(u3__abc_74070_new_n688_));
AND2X2 AND2X2_3272 ( .A(u3__abc_74070_new_n689_), .B(u3__abc_74070_new_n690_), .Y(mem_dout_10_));
AND2X2 AND2X2_3273 ( .A(u3__abc_74070_new_n693_), .B(u3__abc_74070_new_n692_), .Y(u3__abc_74070_new_n694_));
AND2X2 AND2X2_3274 ( .A(u3__abc_74070_new_n695_), .B(u3__abc_74070_new_n696_), .Y(mem_dout_11_));
AND2X2 AND2X2_3275 ( .A(u3__abc_74070_new_n699_), .B(u3__abc_74070_new_n698_), .Y(u3__abc_74070_new_n700_));
AND2X2 AND2X2_3276 ( .A(u3__abc_74070_new_n701_), .B(u3__abc_74070_new_n702_), .Y(mem_dout_12_));
AND2X2 AND2X2_3277 ( .A(u3__abc_74070_new_n705_), .B(u3__abc_74070_new_n704_), .Y(u3__abc_74070_new_n706_));
AND2X2 AND2X2_3278 ( .A(u3__abc_74070_new_n707_), .B(u3__abc_74070_new_n708_), .Y(mem_dout_13_));
AND2X2 AND2X2_3279 ( .A(u3__abc_74070_new_n711_), .B(u3__abc_74070_new_n710_), .Y(u3__abc_74070_new_n712_));
AND2X2 AND2X2_328 ( .A(spec_req_cs_4_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1570_));
AND2X2 AND2X2_3280 ( .A(u3__abc_74070_new_n713_), .B(u3__abc_74070_new_n714_), .Y(mem_dout_14_));
AND2X2 AND2X2_3281 ( .A(u3__abc_74070_new_n717_), .B(u3__abc_74070_new_n716_), .Y(u3__abc_74070_new_n718_));
AND2X2 AND2X2_3282 ( .A(u3__abc_74070_new_n719_), .B(u3__abc_74070_new_n720_), .Y(mem_dout_15_));
AND2X2 AND2X2_3283 ( .A(u3__abc_74070_new_n452__bF_buf2), .B(mc_data_ir_0_), .Y(u3__abc_74070_new_n722_));
AND2X2 AND2X2_3284 ( .A(csc_5_bF_buf0_), .B(mc_data_ir_16_), .Y(u3__abc_74070_new_n723_));
AND2X2 AND2X2_3285 ( .A(u3__abc_74070_new_n450__bF_buf2), .B(u3_byte2_0_), .Y(u3__abc_74070_new_n725_));
AND2X2 AND2X2_3286 ( .A(u3__abc_74070_new_n727_), .B(u3__abc_74070_new_n728_), .Y(mem_dout_16_));
AND2X2 AND2X2_3287 ( .A(u3__abc_74070_new_n452__bF_buf1), .B(mc_data_ir_1_), .Y(u3__abc_74070_new_n730_));
AND2X2 AND2X2_3288 ( .A(csc_5_bF_buf4_), .B(mc_data_ir_17_), .Y(u3__abc_74070_new_n731_));
AND2X2 AND2X2_3289 ( .A(u3__abc_74070_new_n450__bF_buf1), .B(u3_byte2_1_), .Y(u3__abc_74070_new_n733_));
AND2X2 AND2X2_329 ( .A(u0__abc_76628_new_n1571_), .B(u0__abc_76628_new_n1174__bF_buf1), .Y(u0__abc_76628_new_n1572_));
AND2X2 AND2X2_3290 ( .A(u3__abc_74070_new_n735_), .B(u3__abc_74070_new_n736_), .Y(mem_dout_17_));
AND2X2 AND2X2_3291 ( .A(u3__abc_74070_new_n452__bF_buf0), .B(mc_data_ir_2_), .Y(u3__abc_74070_new_n738_));
AND2X2 AND2X2_3292 ( .A(csc_5_bF_buf3_), .B(mc_data_ir_18_), .Y(u3__abc_74070_new_n739_));
AND2X2 AND2X2_3293 ( .A(u3__abc_74070_new_n450__bF_buf0), .B(u3_byte2_2_), .Y(u3__abc_74070_new_n741_));
AND2X2 AND2X2_3294 ( .A(u3__abc_74070_new_n743_), .B(u3__abc_74070_new_n744_), .Y(mem_dout_18_));
AND2X2 AND2X2_3295 ( .A(u3__abc_74070_new_n452__bF_buf3), .B(mc_data_ir_3_), .Y(u3__abc_74070_new_n746_));
AND2X2 AND2X2_3296 ( .A(csc_5_bF_buf2_), .B(mc_data_ir_19_), .Y(u3__abc_74070_new_n747_));
AND2X2 AND2X2_3297 ( .A(u3__abc_74070_new_n450__bF_buf3), .B(u3_byte2_3_), .Y(u3__abc_74070_new_n749_));
AND2X2 AND2X2_3298 ( .A(u3__abc_74070_new_n751_), .B(u3__abc_74070_new_n752_), .Y(mem_dout_19_));
AND2X2 AND2X2_3299 ( .A(u3__abc_74070_new_n452__bF_buf2), .B(mc_data_ir_4_), .Y(u3__abc_74070_new_n754_));
AND2X2 AND2X2_33 ( .A(_abc_85006_new_n335_), .B(_abc_85006_new_n336_), .Y(tms_s_15_));
AND2X2 AND2X2_330 ( .A(spec_req_cs_3_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1573_));
AND2X2 AND2X2_3300 ( .A(csc_5_bF_buf1_), .B(mc_data_ir_20_), .Y(u3__abc_74070_new_n755_));
AND2X2 AND2X2_3301 ( .A(u3__abc_74070_new_n450__bF_buf2), .B(u3_byte2_4_), .Y(u3__abc_74070_new_n757_));
AND2X2 AND2X2_3302 ( .A(u3__abc_74070_new_n759_), .B(u3__abc_74070_new_n760_), .Y(mem_dout_20_));
AND2X2 AND2X2_3303 ( .A(u3__abc_74070_new_n452__bF_buf1), .B(mc_data_ir_5_), .Y(u3__abc_74070_new_n762_));
AND2X2 AND2X2_3304 ( .A(csc_5_bF_buf0_), .B(mc_data_ir_21_), .Y(u3__abc_74070_new_n763_));
AND2X2 AND2X2_3305 ( .A(u3__abc_74070_new_n450__bF_buf1), .B(u3_byte2_5_), .Y(u3__abc_74070_new_n765_));
AND2X2 AND2X2_3306 ( .A(u3__abc_74070_new_n767_), .B(u3__abc_74070_new_n768_), .Y(mem_dout_21_));
AND2X2 AND2X2_3307 ( .A(u3__abc_74070_new_n452__bF_buf0), .B(mc_data_ir_6_), .Y(u3__abc_74070_new_n770_));
AND2X2 AND2X2_3308 ( .A(csc_5_bF_buf4_), .B(mc_data_ir_22_), .Y(u3__abc_74070_new_n771_));
AND2X2 AND2X2_3309 ( .A(u3__abc_74070_new_n450__bF_buf0), .B(u3_byte2_6_), .Y(u3__abc_74070_new_n773_));
AND2X2 AND2X2_331 ( .A(u0__abc_76628_new_n1574_), .B(u0__abc_76628_new_n1173__bF_buf1), .Y(u0__abc_76628_new_n1575_));
AND2X2 AND2X2_3310 ( .A(u3__abc_74070_new_n775_), .B(u3__abc_74070_new_n776_), .Y(mem_dout_22_));
AND2X2 AND2X2_3311 ( .A(u3__abc_74070_new_n452__bF_buf3), .B(mc_data_ir_7_), .Y(u3__abc_74070_new_n778_));
AND2X2 AND2X2_3312 ( .A(csc_5_bF_buf3_), .B(mc_data_ir_23_), .Y(u3__abc_74070_new_n779_));
AND2X2 AND2X2_3313 ( .A(u3__abc_74070_new_n450__bF_buf3), .B(u3_byte2_7_), .Y(u3__abc_74070_new_n781_));
AND2X2 AND2X2_3314 ( .A(u3__abc_74070_new_n783_), .B(u3__abc_74070_new_n784_), .Y(mem_dout_23_));
AND2X2 AND2X2_3315 ( .A(u3__abc_74070_new_n452__bF_buf2), .B(mc_data_ir_8_), .Y(u3__abc_74070_new_n786_));
AND2X2 AND2X2_3316 ( .A(csc_5_bF_buf2_), .B(mc_data_ir_24_), .Y(u3__abc_74070_new_n787_));
AND2X2 AND2X2_3317 ( .A(u3__abc_74070_new_n450__bF_buf2), .B(mc_data_ir_0_), .Y(u3__abc_74070_new_n789_));
AND2X2 AND2X2_3318 ( .A(u3__abc_74070_new_n791_), .B(u3__abc_74070_new_n792_), .Y(mem_dout_24_));
AND2X2 AND2X2_3319 ( .A(u3__abc_74070_new_n452__bF_buf1), .B(mc_data_ir_9_), .Y(u3__abc_74070_new_n794_));
AND2X2 AND2X2_332 ( .A(spec_req_cs_2_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1576_));
AND2X2 AND2X2_3320 ( .A(csc_5_bF_buf1_), .B(mc_data_ir_25_), .Y(u3__abc_74070_new_n795_));
AND2X2 AND2X2_3321 ( .A(u3__abc_74070_new_n450__bF_buf1), .B(mc_data_ir_1_), .Y(u3__abc_74070_new_n797_));
AND2X2 AND2X2_3322 ( .A(u3__abc_74070_new_n799_), .B(u3__abc_74070_new_n800_), .Y(mem_dout_25_));
AND2X2 AND2X2_3323 ( .A(u3__abc_74070_new_n452__bF_buf0), .B(mc_data_ir_10_), .Y(u3__abc_74070_new_n802_));
AND2X2 AND2X2_3324 ( .A(csc_5_bF_buf0_), .B(mc_data_ir_26_), .Y(u3__abc_74070_new_n803_));
AND2X2 AND2X2_3325 ( .A(u3__abc_74070_new_n450__bF_buf0), .B(mc_data_ir_2_), .Y(u3__abc_74070_new_n805_));
AND2X2 AND2X2_3326 ( .A(u3__abc_74070_new_n807_), .B(u3__abc_74070_new_n808_), .Y(mem_dout_26_));
AND2X2 AND2X2_3327 ( .A(u3__abc_74070_new_n452__bF_buf3), .B(mc_data_ir_11_), .Y(u3__abc_74070_new_n810_));
AND2X2 AND2X2_3328 ( .A(csc_5_bF_buf4_), .B(mc_data_ir_27_), .Y(u3__abc_74070_new_n811_));
AND2X2 AND2X2_3329 ( .A(u3__abc_74070_new_n450__bF_buf3), .B(mc_data_ir_3_), .Y(u3__abc_74070_new_n813_));
AND2X2 AND2X2_333 ( .A(u0__abc_76628_new_n1577_), .B(u0__abc_76628_new_n1172__bF_buf1), .Y(u0__abc_76628_new_n1578_));
AND2X2 AND2X2_3330 ( .A(u3__abc_74070_new_n815_), .B(u3__abc_74070_new_n816_), .Y(mem_dout_27_));
AND2X2 AND2X2_3331 ( .A(u3__abc_74070_new_n452__bF_buf2), .B(mc_data_ir_12_), .Y(u3__abc_74070_new_n818_));
AND2X2 AND2X2_3332 ( .A(csc_5_bF_buf3_), .B(mc_data_ir_28_), .Y(u3__abc_74070_new_n819_));
AND2X2 AND2X2_3333 ( .A(u3__abc_74070_new_n450__bF_buf2), .B(mc_data_ir_4_), .Y(u3__abc_74070_new_n821_));
AND2X2 AND2X2_3334 ( .A(u3__abc_74070_new_n823_), .B(u3__abc_74070_new_n824_), .Y(mem_dout_28_));
AND2X2 AND2X2_3335 ( .A(u3__abc_74070_new_n452__bF_buf1), .B(mc_data_ir_13_), .Y(u3__abc_74070_new_n826_));
AND2X2 AND2X2_3336 ( .A(csc_5_bF_buf2_), .B(mc_data_ir_29_), .Y(u3__abc_74070_new_n827_));
AND2X2 AND2X2_3337 ( .A(u3__abc_74070_new_n450__bF_buf1), .B(mc_data_ir_5_), .Y(u3__abc_74070_new_n829_));
AND2X2 AND2X2_3338 ( .A(u3__abc_74070_new_n831_), .B(u3__abc_74070_new_n832_), .Y(mem_dout_29_));
AND2X2 AND2X2_3339 ( .A(u3__abc_74070_new_n452__bF_buf0), .B(mc_data_ir_14_), .Y(u3__abc_74070_new_n834_));
AND2X2 AND2X2_334 ( .A(spec_req_cs_1_bF_buf4_), .B(u0_tms1_16_), .Y(u0__abc_76628_new_n1579_));
AND2X2 AND2X2_3340 ( .A(csc_5_bF_buf1_), .B(mc_data_ir_30_), .Y(u3__abc_74070_new_n835_));
AND2X2 AND2X2_3341 ( .A(u3__abc_74070_new_n450__bF_buf0), .B(mc_data_ir_6_), .Y(u3__abc_74070_new_n837_));
AND2X2 AND2X2_3342 ( .A(u3__abc_74070_new_n839_), .B(u3__abc_74070_new_n840_), .Y(mem_dout_30_));
AND2X2 AND2X2_3343 ( .A(u3__abc_74070_new_n452__bF_buf3), .B(mc_data_ir_15_), .Y(u3__abc_74070_new_n842_));
AND2X2 AND2X2_3344 ( .A(csc_5_bF_buf0_), .B(mc_data_ir_31_), .Y(u3__abc_74070_new_n843_));
AND2X2 AND2X2_3345 ( .A(u3__abc_74070_new_n450__bF_buf3), .B(mc_data_ir_7_), .Y(u3__abc_74070_new_n845_));
AND2X2 AND2X2_3346 ( .A(u3__abc_74070_new_n847_), .B(u3__abc_74070_new_n848_), .Y(mem_dout_31_));
AND2X2 AND2X2_3347 ( .A(wb_stb_i_bF_buf1), .B(wb_we_i), .Y(u3__abc_74070_new_n851_));
AND2X2 AND2X2_3348 ( .A(mem_ack_r), .B(u3_wb_read_go), .Y(u3_re));
AND2X2 AND2X2_3349 ( .A(u3_rd_fifo_out_22_), .B(u3_rd_fifo_out_23_), .Y(u3__abc_74070_new_n855_));
AND2X2 AND2X2_335 ( .A(u0__abc_76628_new_n1169__bF_buf3), .B(u0__abc_76628_new_n1582_), .Y(u0__abc_76628_new_n1583_));
AND2X2 AND2X2_3350 ( .A(u3__abc_74070_new_n856_), .B(u3__abc_74070_new_n854_), .Y(u3__abc_74070_new_n857_));
AND2X2 AND2X2_3351 ( .A(u3__abc_74070_new_n859_), .B(u3__abc_74070_new_n861_), .Y(u3__abc_74070_new_n862_));
AND2X2 AND2X2_3352 ( .A(u3__abc_74070_new_n862_), .B(u3_rd_fifo_out_34_), .Y(u3__abc_74070_new_n863_));
AND2X2 AND2X2_3353 ( .A(u3__abc_74070_new_n860_), .B(u3_rd_fifo_out_16_), .Y(u3__abc_74070_new_n865_));
AND2X2 AND2X2_3354 ( .A(u3__abc_74070_new_n858_), .B(u3_rd_fifo_out_17_), .Y(u3__abc_74070_new_n866_));
AND2X2 AND2X2_3355 ( .A(u3__abc_74070_new_n867_), .B(u3__abc_74070_new_n864_), .Y(u3__abc_74070_new_n868_));
AND2X2 AND2X2_3356 ( .A(u3__abc_74070_new_n869_), .B(u3__abc_74070_new_n857_), .Y(u3__abc_74070_new_n870_));
AND2X2 AND2X2_3357 ( .A(u3__abc_74070_new_n872_), .B(u3__abc_74070_new_n873_), .Y(u3__abc_74070_new_n874_));
AND2X2 AND2X2_3358 ( .A(u3__abc_74070_new_n874_), .B(u3__abc_74070_new_n871_), .Y(u3__abc_74070_new_n875_));
AND2X2 AND2X2_3359 ( .A(u3_rd_fifo_out_20_), .B(u3_rd_fifo_out_21_), .Y(u3__abc_74070_new_n879_));
AND2X2 AND2X2_336 ( .A(u0__abc_76628_new_n1581_), .B(u0__abc_76628_new_n1583_), .Y(u0__abc_76628_new_n1584_));
AND2X2 AND2X2_3360 ( .A(u3__abc_74070_new_n880_), .B(u3__abc_74070_new_n878_), .Y(u3__abc_74070_new_n881_));
AND2X2 AND2X2_3361 ( .A(u3__abc_74070_new_n882_), .B(u3_rd_fifo_out_18_), .Y(u3__abc_74070_new_n883_));
AND2X2 AND2X2_3362 ( .A(u3__abc_74070_new_n884_), .B(u3__abc_74070_new_n885_), .Y(u3__abc_74070_new_n886_));
AND2X2 AND2X2_3363 ( .A(u3__abc_74070_new_n890_), .B(u3__abc_74070_new_n887_), .Y(u3__abc_74070_new_n891_));
AND2X2 AND2X2_3364 ( .A(u3__abc_74070_new_n894_), .B(\wb_sel_i[2] ), .Y(u3__abc_74070_new_n895_));
AND2X2 AND2X2_3365 ( .A(u3__abc_74070_new_n895_), .B(u3__abc_74070_new_n893_), .Y(u3__abc_74070_new_n896_));
AND2X2 AND2X2_3366 ( .A(u3_rd_fifo_out_30_), .B(u3_rd_fifo_out_31_), .Y(u3__abc_74070_new_n898_));
AND2X2 AND2X2_3367 ( .A(u3__abc_74070_new_n899_), .B(u3__abc_74070_new_n897_), .Y(u3__abc_74070_new_n900_));
AND2X2 AND2X2_3368 ( .A(u3__abc_74070_new_n901_), .B(u3__abc_74070_new_n902_), .Y(u3__abc_74070_new_n903_));
AND2X2 AND2X2_3369 ( .A(u3_rd_fifo_out_24_), .B(u3_rd_fifo_out_25_), .Y(u3__abc_74070_new_n904_));
AND2X2 AND2X2_337 ( .A(u0__abc_76628_new_n1170__bF_buf3), .B(sp_tms_17_), .Y(u0__abc_76628_new_n1586_));
AND2X2 AND2X2_3370 ( .A(u3__abc_74070_new_n905_), .B(u3_rd_fifo_out_35_), .Y(u3__abc_74070_new_n906_));
AND2X2 AND2X2_3371 ( .A(u3__abc_74070_new_n909_), .B(u3__abc_74070_new_n908_), .Y(u3__abc_74070_new_n910_));
AND2X2 AND2X2_3372 ( .A(u3__abc_74070_new_n910_), .B(u3__abc_74070_new_n907_), .Y(u3__abc_74070_new_n911_));
AND2X2 AND2X2_3373 ( .A(u3__abc_74070_new_n912_), .B(u3__abc_74070_new_n900_), .Y(u3__abc_74070_new_n913_));
AND2X2 AND2X2_3374 ( .A(u3__abc_74070_new_n916_), .B(u3__abc_74070_new_n915_), .Y(u3__abc_74070_new_n917_));
AND2X2 AND2X2_3375 ( .A(u3__abc_74070_new_n917_), .B(u3__abc_74070_new_n914_), .Y(u3__abc_74070_new_n918_));
AND2X2 AND2X2_3376 ( .A(u3_rd_fifo_out_28_), .B(u3_rd_fifo_out_29_), .Y(u3__abc_74070_new_n922_));
AND2X2 AND2X2_3377 ( .A(u3__abc_74070_new_n923_), .B(u3__abc_74070_new_n921_), .Y(u3__abc_74070_new_n924_));
AND2X2 AND2X2_3378 ( .A(u3__abc_74070_new_n925_), .B(u3_rd_fifo_out_26_), .Y(u3__abc_74070_new_n926_));
AND2X2 AND2X2_3379 ( .A(u3__abc_74070_new_n927_), .B(u3__abc_74070_new_n928_), .Y(u3__abc_74070_new_n929_));
AND2X2 AND2X2_338 ( .A(spec_req_cs_5_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1587_));
AND2X2 AND2X2_3380 ( .A(u3__abc_74070_new_n933_), .B(u3__abc_74070_new_n930_), .Y(u3__abc_74070_new_n934_));
AND2X2 AND2X2_3381 ( .A(u3__abc_74070_new_n937_), .B(\wb_sel_i[3] ), .Y(u3__abc_74070_new_n938_));
AND2X2 AND2X2_3382 ( .A(u3__abc_74070_new_n938_), .B(u3__abc_74070_new_n936_), .Y(u3__abc_74070_new_n939_));
AND2X2 AND2X2_3383 ( .A(u3_rd_fifo_out_14_), .B(u3_rd_fifo_out_15_), .Y(u3__abc_74070_new_n942_));
AND2X2 AND2X2_3384 ( .A(u3__abc_74070_new_n943_), .B(u3__abc_74070_new_n941_), .Y(u3__abc_74070_new_n944_));
AND2X2 AND2X2_3385 ( .A(u3_rd_fifo_out_8_), .B(u3_rd_fifo_out_9_), .Y(u3__abc_74070_new_n948_));
AND2X2 AND2X2_3386 ( .A(u3__abc_74070_new_n949_), .B(u3__abc_74070_new_n947_), .Y(u3__abc_74070_new_n950_));
AND2X2 AND2X2_3387 ( .A(u3__abc_74070_new_n952_), .B(u3__abc_74070_new_n953_), .Y(u3__abc_74070_new_n954_));
AND2X2 AND2X2_3388 ( .A(u3__abc_74070_new_n956_), .B(u3__abc_74070_new_n951_), .Y(u3__abc_74070_new_n957_));
AND2X2 AND2X2_3389 ( .A(u3__abc_74070_new_n955_), .B(u3_rd_fifo_out_33_), .Y(u3__abc_74070_new_n959_));
AND2X2 AND2X2_339 ( .A(u0__abc_76628_new_n1589_), .B(u0__abc_76628_new_n1179__bF_buf0), .Y(u0__abc_76628_new_n1590_));
AND2X2 AND2X2_3390 ( .A(u3__abc_74070_new_n950_), .B(u3__abc_74070_new_n946_), .Y(u3__abc_74070_new_n960_));
AND2X2 AND2X2_3391 ( .A(u3__abc_74070_new_n958_), .B(u3__abc_74070_new_n962_), .Y(u3__abc_74070_new_n963_));
AND2X2 AND2X2_3392 ( .A(u3_rd_fifo_out_12_), .B(u3_rd_fifo_out_13_), .Y(u3__abc_74070_new_n966_));
AND2X2 AND2X2_3393 ( .A(u3__abc_74070_new_n967_), .B(u3__abc_74070_new_n965_), .Y(u3__abc_74070_new_n968_));
AND2X2 AND2X2_3394 ( .A(u3__abc_74070_new_n970_), .B(u3_rd_fifo_out_10_), .Y(u3__abc_74070_new_n971_));
AND2X2 AND2X2_3395 ( .A(u3__abc_74070_new_n972_), .B(u3__abc_74070_new_n973_), .Y(u3__abc_74070_new_n974_));
AND2X2 AND2X2_3396 ( .A(u3__abc_74070_new_n975_), .B(u3__abc_74070_new_n969_), .Y(u3__abc_74070_new_n976_));
AND2X2 AND2X2_3397 ( .A(u3__abc_74070_new_n974_), .B(u3__abc_74070_new_n968_), .Y(u3__abc_74070_new_n977_));
AND2X2 AND2X2_3398 ( .A(u3__abc_74070_new_n981_), .B(\wb_sel_i[1] ), .Y(u3__abc_74070_new_n982_));
AND2X2 AND2X2_3399 ( .A(u3__abc_74070_new_n982_), .B(u3__abc_74070_new_n980_), .Y(u3__abc_74070_new_n983_));
AND2X2 AND2X2_34 ( .A(_abc_85006_new_n338_), .B(_abc_85006_new_n339_), .Y(tms_s_16_));
AND2X2 AND2X2_340 ( .A(u0__abc_76628_new_n1590_), .B(u0__abc_76628_new_n1588_), .Y(u0__abc_76628_new_n1591_));
AND2X2 AND2X2_3400 ( .A(u3_rd_fifo_out_6_), .B(u3_rd_fifo_out_7_), .Y(u3__abc_74070_new_n985_));
AND2X2 AND2X2_3401 ( .A(u3__abc_74070_new_n986_), .B(u3__abc_74070_new_n984_), .Y(u3__abc_74070_new_n987_));
AND2X2 AND2X2_3402 ( .A(u3_rd_fifo_out_0_), .B(u3_rd_fifo_out_1_), .Y(u3__abc_74070_new_n991_));
AND2X2 AND2X2_3403 ( .A(u3__abc_74070_new_n992_), .B(u3__abc_74070_new_n990_), .Y(u3__abc_74070_new_n993_));
AND2X2 AND2X2_3404 ( .A(u3__abc_74070_new_n996_), .B(u3__abc_74070_new_n998_), .Y(u3__abc_74070_new_n999_));
AND2X2 AND2X2_3405 ( .A(u3__abc_74070_new_n1000_), .B(u3__abc_74070_new_n994_), .Y(u3__abc_74070_new_n1001_));
AND2X2 AND2X2_3406 ( .A(u3__abc_74070_new_n999_), .B(u3_rd_fifo_out_32_), .Y(u3__abc_74070_new_n1003_));
AND2X2 AND2X2_3407 ( .A(u3__abc_74070_new_n993_), .B(u3__abc_74070_new_n989_), .Y(u3__abc_74070_new_n1004_));
AND2X2 AND2X2_3408 ( .A(u3__abc_74070_new_n1002_), .B(u3__abc_74070_new_n1006_), .Y(u3__abc_74070_new_n1007_));
AND2X2 AND2X2_3409 ( .A(u3_rd_fifo_out_4_), .B(u3_rd_fifo_out_5_), .Y(u3__abc_74070_new_n1010_));
AND2X2 AND2X2_341 ( .A(u0__abc_76628_new_n1592_), .B(u0__abc_76628_new_n1175__bF_buf0), .Y(u0__abc_76628_new_n1593_));
AND2X2 AND2X2_3410 ( .A(u3__abc_74070_new_n1011_), .B(u3__abc_74070_new_n1009_), .Y(u3__abc_74070_new_n1012_));
AND2X2 AND2X2_3411 ( .A(u3__abc_74070_new_n1014_), .B(u3_rd_fifo_out_2_), .Y(u3__abc_74070_new_n1015_));
AND2X2 AND2X2_3412 ( .A(u3__abc_74070_new_n1016_), .B(u3__abc_74070_new_n1017_), .Y(u3__abc_74070_new_n1018_));
AND2X2 AND2X2_3413 ( .A(u3__abc_74070_new_n1019_), .B(u3__abc_74070_new_n1013_), .Y(u3__abc_74070_new_n1020_));
AND2X2 AND2X2_3414 ( .A(u3__abc_74070_new_n1018_), .B(u3__abc_74070_new_n1012_), .Y(u3__abc_74070_new_n1021_));
AND2X2 AND2X2_3415 ( .A(u3__abc_74070_new_n1025_), .B(\wb_sel_i[0] ), .Y(u3__abc_74070_new_n1026_));
AND2X2 AND2X2_3416 ( .A(u3__abc_74070_new_n1026_), .B(u3__abc_74070_new_n1024_), .Y(u3__abc_74070_new_n1027_));
AND2X2 AND2X2_3417 ( .A(u3__abc_74070_new_n1030_), .B(mem_ack), .Y(u3__abc_74070_new_n1031_));
AND2X2 AND2X2_3418 ( .A(u3__abc_74070_new_n1031_), .B(u3_pen), .Y(u3__abc_74070_new_n1032_));
AND2X2 AND2X2_3419 ( .A(u3__abc_74070_new_n1029_), .B(u3__abc_74070_new_n1032_), .Y(par_err));
AND2X2 AND2X2_342 ( .A(spec_req_cs_4_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1594_));
AND2X2 AND2X2_3420 ( .A(u3_u0_wr_adr_1_), .B(dv), .Y(u3_u0__abc_75526_new_n382_));
AND2X2 AND2X2_3421 ( .A(u3_u0__abc_75526_new_n382__bF_buf6), .B(u3_u0__abc_75526_new_n384_), .Y(u3_u0__abc_75526_new_n385_));
AND2X2 AND2X2_3422 ( .A(u3_u0__abc_75526_new_n386_), .B(u3_u0__abc_75526_new_n383_), .Y(u3_u0__0r1_35_0__0_));
AND2X2 AND2X2_3423 ( .A(u3_u0__abc_75526_new_n382__bF_buf4), .B(u3_u0__abc_75526_new_n389_), .Y(u3_u0__abc_75526_new_n390_));
AND2X2 AND2X2_3424 ( .A(u3_u0__abc_75526_new_n391_), .B(u3_u0__abc_75526_new_n388_), .Y(u3_u0__0r1_35_0__1_));
AND2X2 AND2X2_3425 ( .A(u3_u0__abc_75526_new_n382__bF_buf2), .B(u3_u0__abc_75526_new_n394_), .Y(u3_u0__abc_75526_new_n395_));
AND2X2 AND2X2_3426 ( .A(u3_u0__abc_75526_new_n396_), .B(u3_u0__abc_75526_new_n393_), .Y(u3_u0__0r1_35_0__2_));
AND2X2 AND2X2_3427 ( .A(u3_u0__abc_75526_new_n382__bF_buf0), .B(u3_u0__abc_75526_new_n399_), .Y(u3_u0__abc_75526_new_n400_));
AND2X2 AND2X2_3428 ( .A(u3_u0__abc_75526_new_n401_), .B(u3_u0__abc_75526_new_n398_), .Y(u3_u0__0r1_35_0__3_));
AND2X2 AND2X2_3429 ( .A(u3_u0__abc_75526_new_n382__bF_buf6), .B(u3_u0__abc_75526_new_n404_), .Y(u3_u0__abc_75526_new_n405_));
AND2X2 AND2X2_343 ( .A(u0__abc_76628_new_n1595_), .B(u0__abc_76628_new_n1174__bF_buf0), .Y(u0__abc_76628_new_n1596_));
AND2X2 AND2X2_3430 ( .A(u3_u0__abc_75526_new_n406_), .B(u3_u0__abc_75526_new_n403_), .Y(u3_u0__0r1_35_0__4_));
AND2X2 AND2X2_3431 ( .A(u3_u0__abc_75526_new_n382__bF_buf4), .B(u3_u0__abc_75526_new_n409_), .Y(u3_u0__abc_75526_new_n410_));
AND2X2 AND2X2_3432 ( .A(u3_u0__abc_75526_new_n411_), .B(u3_u0__abc_75526_new_n408_), .Y(u3_u0__0r1_35_0__5_));
AND2X2 AND2X2_3433 ( .A(u3_u0__abc_75526_new_n382__bF_buf2), .B(u3_u0__abc_75526_new_n414_), .Y(u3_u0__abc_75526_new_n415_));
AND2X2 AND2X2_3434 ( .A(u3_u0__abc_75526_new_n416_), .B(u3_u0__abc_75526_new_n413_), .Y(u3_u0__0r1_35_0__6_));
AND2X2 AND2X2_3435 ( .A(u3_u0__abc_75526_new_n382__bF_buf0), .B(u3_u0__abc_75526_new_n419_), .Y(u3_u0__abc_75526_new_n420_));
AND2X2 AND2X2_3436 ( .A(u3_u0__abc_75526_new_n421_), .B(u3_u0__abc_75526_new_n418_), .Y(u3_u0__0r1_35_0__7_));
AND2X2 AND2X2_3437 ( .A(u3_u0__abc_75526_new_n382__bF_buf6), .B(u3_u0__abc_75526_new_n424_), .Y(u3_u0__abc_75526_new_n425_));
AND2X2 AND2X2_3438 ( .A(u3_u0__abc_75526_new_n426_), .B(u3_u0__abc_75526_new_n423_), .Y(u3_u0__0r1_35_0__8_));
AND2X2 AND2X2_3439 ( .A(u3_u0__abc_75526_new_n382__bF_buf4), .B(u3_u0__abc_75526_new_n429_), .Y(u3_u0__abc_75526_new_n430_));
AND2X2 AND2X2_344 ( .A(spec_req_cs_3_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1597_));
AND2X2 AND2X2_3440 ( .A(u3_u0__abc_75526_new_n431_), .B(u3_u0__abc_75526_new_n428_), .Y(u3_u0__0r1_35_0__9_));
AND2X2 AND2X2_3441 ( .A(u3_u0__abc_75526_new_n382__bF_buf2), .B(u3_u0__abc_75526_new_n434_), .Y(u3_u0__abc_75526_new_n435_));
AND2X2 AND2X2_3442 ( .A(u3_u0__abc_75526_new_n436_), .B(u3_u0__abc_75526_new_n433_), .Y(u3_u0__0r1_35_0__10_));
AND2X2 AND2X2_3443 ( .A(u3_u0__abc_75526_new_n382__bF_buf0), .B(u3_u0__abc_75526_new_n439_), .Y(u3_u0__abc_75526_new_n440_));
AND2X2 AND2X2_3444 ( .A(u3_u0__abc_75526_new_n441_), .B(u3_u0__abc_75526_new_n438_), .Y(u3_u0__0r1_35_0__11_));
AND2X2 AND2X2_3445 ( .A(u3_u0__abc_75526_new_n382__bF_buf6), .B(u3_u0__abc_75526_new_n444_), .Y(u3_u0__abc_75526_new_n445_));
AND2X2 AND2X2_3446 ( .A(u3_u0__abc_75526_new_n446_), .B(u3_u0__abc_75526_new_n443_), .Y(u3_u0__0r1_35_0__12_));
AND2X2 AND2X2_3447 ( .A(u3_u0__abc_75526_new_n382__bF_buf4), .B(u3_u0__abc_75526_new_n449_), .Y(u3_u0__abc_75526_new_n450_));
AND2X2 AND2X2_3448 ( .A(u3_u0__abc_75526_new_n451_), .B(u3_u0__abc_75526_new_n448_), .Y(u3_u0__0r1_35_0__13_));
AND2X2 AND2X2_3449 ( .A(u3_u0__abc_75526_new_n382__bF_buf2), .B(u3_u0__abc_75526_new_n454_), .Y(u3_u0__abc_75526_new_n455_));
AND2X2 AND2X2_345 ( .A(u0__abc_76628_new_n1598_), .B(u0__abc_76628_new_n1173__bF_buf0), .Y(u0__abc_76628_new_n1599_));
AND2X2 AND2X2_3450 ( .A(u3_u0__abc_75526_new_n456_), .B(u3_u0__abc_75526_new_n453_), .Y(u3_u0__0r1_35_0__14_));
AND2X2 AND2X2_3451 ( .A(u3_u0__abc_75526_new_n382__bF_buf0), .B(u3_u0__abc_75526_new_n459_), .Y(u3_u0__abc_75526_new_n460_));
AND2X2 AND2X2_3452 ( .A(u3_u0__abc_75526_new_n461_), .B(u3_u0__abc_75526_new_n458_), .Y(u3_u0__0r1_35_0__15_));
AND2X2 AND2X2_3453 ( .A(u3_u0__abc_75526_new_n382__bF_buf6), .B(u3_u0__abc_75526_new_n464_), .Y(u3_u0__abc_75526_new_n465_));
AND2X2 AND2X2_3454 ( .A(u3_u0__abc_75526_new_n466_), .B(u3_u0__abc_75526_new_n463_), .Y(u3_u0__0r1_35_0__16_));
AND2X2 AND2X2_3455 ( .A(u3_u0__abc_75526_new_n382__bF_buf4), .B(u3_u0__abc_75526_new_n469_), .Y(u3_u0__abc_75526_new_n470_));
AND2X2 AND2X2_3456 ( .A(u3_u0__abc_75526_new_n471_), .B(u3_u0__abc_75526_new_n468_), .Y(u3_u0__0r1_35_0__17_));
AND2X2 AND2X2_3457 ( .A(u3_u0__abc_75526_new_n382__bF_buf2), .B(u3_u0__abc_75526_new_n474_), .Y(u3_u0__abc_75526_new_n475_));
AND2X2 AND2X2_3458 ( .A(u3_u0__abc_75526_new_n476_), .B(u3_u0__abc_75526_new_n473_), .Y(u3_u0__0r1_35_0__18_));
AND2X2 AND2X2_3459 ( .A(u3_u0__abc_75526_new_n382__bF_buf0), .B(u3_u0__abc_75526_new_n479_), .Y(u3_u0__abc_75526_new_n480_));
AND2X2 AND2X2_346 ( .A(spec_req_cs_2_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1600_));
AND2X2 AND2X2_3460 ( .A(u3_u0__abc_75526_new_n481_), .B(u3_u0__abc_75526_new_n478_), .Y(u3_u0__0r1_35_0__19_));
AND2X2 AND2X2_3461 ( .A(u3_u0__abc_75526_new_n382__bF_buf6), .B(u3_u0__abc_75526_new_n484_), .Y(u3_u0__abc_75526_new_n485_));
AND2X2 AND2X2_3462 ( .A(u3_u0__abc_75526_new_n486_), .B(u3_u0__abc_75526_new_n483_), .Y(u3_u0__0r1_35_0__20_));
AND2X2 AND2X2_3463 ( .A(u3_u0__abc_75526_new_n382__bF_buf4), .B(u3_u0__abc_75526_new_n489_), .Y(u3_u0__abc_75526_new_n490_));
AND2X2 AND2X2_3464 ( .A(u3_u0__abc_75526_new_n491_), .B(u3_u0__abc_75526_new_n488_), .Y(u3_u0__0r1_35_0__21_));
AND2X2 AND2X2_3465 ( .A(u3_u0__abc_75526_new_n382__bF_buf2), .B(u3_u0__abc_75526_new_n494_), .Y(u3_u0__abc_75526_new_n495_));
AND2X2 AND2X2_3466 ( .A(u3_u0__abc_75526_new_n496_), .B(u3_u0__abc_75526_new_n493_), .Y(u3_u0__0r1_35_0__22_));
AND2X2 AND2X2_3467 ( .A(u3_u0__abc_75526_new_n382__bF_buf0), .B(u3_u0__abc_75526_new_n499_), .Y(u3_u0__abc_75526_new_n500_));
AND2X2 AND2X2_3468 ( .A(u3_u0__abc_75526_new_n501_), .B(u3_u0__abc_75526_new_n498_), .Y(u3_u0__0r1_35_0__23_));
AND2X2 AND2X2_3469 ( .A(u3_u0__abc_75526_new_n382__bF_buf6), .B(u3_u0__abc_75526_new_n504_), .Y(u3_u0__abc_75526_new_n505_));
AND2X2 AND2X2_347 ( .A(u0__abc_76628_new_n1601_), .B(u0__abc_76628_new_n1172__bF_buf0), .Y(u0__abc_76628_new_n1602_));
AND2X2 AND2X2_3470 ( .A(u3_u0__abc_75526_new_n506_), .B(u3_u0__abc_75526_new_n503_), .Y(u3_u0__0r1_35_0__24_));
AND2X2 AND2X2_3471 ( .A(u3_u0__abc_75526_new_n382__bF_buf4), .B(u3_u0__abc_75526_new_n509_), .Y(u3_u0__abc_75526_new_n510_));
AND2X2 AND2X2_3472 ( .A(u3_u0__abc_75526_new_n511_), .B(u3_u0__abc_75526_new_n508_), .Y(u3_u0__0r1_35_0__25_));
AND2X2 AND2X2_3473 ( .A(u3_u0__abc_75526_new_n382__bF_buf2), .B(u3_u0__abc_75526_new_n514_), .Y(u3_u0__abc_75526_new_n515_));
AND2X2 AND2X2_3474 ( .A(u3_u0__abc_75526_new_n516_), .B(u3_u0__abc_75526_new_n513_), .Y(u3_u0__0r1_35_0__26_));
AND2X2 AND2X2_3475 ( .A(u3_u0__abc_75526_new_n382__bF_buf0), .B(u3_u0__abc_75526_new_n519_), .Y(u3_u0__abc_75526_new_n520_));
AND2X2 AND2X2_3476 ( .A(u3_u0__abc_75526_new_n521_), .B(u3_u0__abc_75526_new_n518_), .Y(u3_u0__0r1_35_0__27_));
AND2X2 AND2X2_3477 ( .A(u3_u0__abc_75526_new_n382__bF_buf6), .B(u3_u0__abc_75526_new_n524_), .Y(u3_u0__abc_75526_new_n525_));
AND2X2 AND2X2_3478 ( .A(u3_u0__abc_75526_new_n526_), .B(u3_u0__abc_75526_new_n523_), .Y(u3_u0__0r1_35_0__28_));
AND2X2 AND2X2_3479 ( .A(u3_u0__abc_75526_new_n382__bF_buf4), .B(u3_u0__abc_75526_new_n529_), .Y(u3_u0__abc_75526_new_n530_));
AND2X2 AND2X2_348 ( .A(spec_req_cs_1_bF_buf3_), .B(u0_tms1_17_), .Y(u0__abc_76628_new_n1603_));
AND2X2 AND2X2_3480 ( .A(u3_u0__abc_75526_new_n531_), .B(u3_u0__abc_75526_new_n528_), .Y(u3_u0__0r1_35_0__29_));
AND2X2 AND2X2_3481 ( .A(u3_u0__abc_75526_new_n382__bF_buf2), .B(u3_u0__abc_75526_new_n534_), .Y(u3_u0__abc_75526_new_n535_));
AND2X2 AND2X2_3482 ( .A(u3_u0__abc_75526_new_n536_), .B(u3_u0__abc_75526_new_n533_), .Y(u3_u0__0r1_35_0__30_));
AND2X2 AND2X2_3483 ( .A(u3_u0__abc_75526_new_n382__bF_buf0), .B(u3_u0__abc_75526_new_n539_), .Y(u3_u0__abc_75526_new_n540_));
AND2X2 AND2X2_3484 ( .A(u3_u0__abc_75526_new_n541_), .B(u3_u0__abc_75526_new_n538_), .Y(u3_u0__0r1_35_0__31_));
AND2X2 AND2X2_3485 ( .A(u3_u0__abc_75526_new_n382__bF_buf6), .B(u3_u0__abc_75526_new_n544_), .Y(u3_u0__abc_75526_new_n545_));
AND2X2 AND2X2_3486 ( .A(u3_u0__abc_75526_new_n546_), .B(u3_u0__abc_75526_new_n543_), .Y(u3_u0__0r1_35_0__32_));
AND2X2 AND2X2_3487 ( .A(u3_u0__abc_75526_new_n382__bF_buf4), .B(u3_u0__abc_75526_new_n549_), .Y(u3_u0__abc_75526_new_n550_));
AND2X2 AND2X2_3488 ( .A(u3_u0__abc_75526_new_n551_), .B(u3_u0__abc_75526_new_n548_), .Y(u3_u0__0r1_35_0__33_));
AND2X2 AND2X2_3489 ( .A(u3_u0__abc_75526_new_n382__bF_buf2), .B(u3_u0__abc_75526_new_n554_), .Y(u3_u0__abc_75526_new_n555_));
AND2X2 AND2X2_349 ( .A(u0__abc_76628_new_n1169__bF_buf2), .B(u0__abc_76628_new_n1606_), .Y(u0__abc_76628_new_n1607_));
AND2X2 AND2X2_3490 ( .A(u3_u0__abc_75526_new_n556_), .B(u3_u0__abc_75526_new_n553_), .Y(u3_u0__0r1_35_0__34_));
AND2X2 AND2X2_3491 ( .A(u3_u0__abc_75526_new_n382__bF_buf0), .B(u3_u0__abc_75526_new_n559_), .Y(u3_u0__abc_75526_new_n560_));
AND2X2 AND2X2_3492 ( .A(u3_u0__abc_75526_new_n561_), .B(u3_u0__abc_75526_new_n558_), .Y(u3_u0__0r1_35_0__35_));
AND2X2 AND2X2_3493 ( .A(dv), .B(u3_u0_wr_adr_3_), .Y(u3_u0__abc_75526_new_n563_));
AND2X2 AND2X2_3494 ( .A(u3_u0__abc_75526_new_n563__bF_buf6), .B(u3_u0__abc_75526_new_n384_), .Y(u3_u0__abc_75526_new_n565_));
AND2X2 AND2X2_3495 ( .A(u3_u0__abc_75526_new_n566_), .B(u3_u0__abc_75526_new_n564_), .Y(u3_u0__0r3_35_0__0_));
AND2X2 AND2X2_3496 ( .A(u3_u0__abc_75526_new_n563__bF_buf4), .B(u3_u0__abc_75526_new_n389_), .Y(u3_u0__abc_75526_new_n569_));
AND2X2 AND2X2_3497 ( .A(u3_u0__abc_75526_new_n570_), .B(u3_u0__abc_75526_new_n568_), .Y(u3_u0__0r3_35_0__1_));
AND2X2 AND2X2_3498 ( .A(u3_u0__abc_75526_new_n563__bF_buf2), .B(u3_u0__abc_75526_new_n394_), .Y(u3_u0__abc_75526_new_n573_));
AND2X2 AND2X2_3499 ( .A(u3_u0__abc_75526_new_n574_), .B(u3_u0__abc_75526_new_n572_), .Y(u3_u0__0r3_35_0__2_));
AND2X2 AND2X2_35 ( .A(_abc_85006_new_n341_), .B(_abc_85006_new_n342_), .Y(tms_s_17_));
AND2X2 AND2X2_350 ( .A(u0__abc_76628_new_n1605_), .B(u0__abc_76628_new_n1607_), .Y(u0__abc_76628_new_n1608_));
AND2X2 AND2X2_3500 ( .A(u3_u0__abc_75526_new_n563__bF_buf0), .B(u3_u0__abc_75526_new_n399_), .Y(u3_u0__abc_75526_new_n577_));
AND2X2 AND2X2_3501 ( .A(u3_u0__abc_75526_new_n578_), .B(u3_u0__abc_75526_new_n576_), .Y(u3_u0__0r3_35_0__3_));
AND2X2 AND2X2_3502 ( .A(u3_u0__abc_75526_new_n563__bF_buf6), .B(u3_u0__abc_75526_new_n404_), .Y(u3_u0__abc_75526_new_n581_));
AND2X2 AND2X2_3503 ( .A(u3_u0__abc_75526_new_n582_), .B(u3_u0__abc_75526_new_n580_), .Y(u3_u0__0r3_35_0__4_));
AND2X2 AND2X2_3504 ( .A(u3_u0__abc_75526_new_n563__bF_buf4), .B(u3_u0__abc_75526_new_n409_), .Y(u3_u0__abc_75526_new_n585_));
AND2X2 AND2X2_3505 ( .A(u3_u0__abc_75526_new_n586_), .B(u3_u0__abc_75526_new_n584_), .Y(u3_u0__0r3_35_0__5_));
AND2X2 AND2X2_3506 ( .A(u3_u0__abc_75526_new_n563__bF_buf2), .B(u3_u0__abc_75526_new_n414_), .Y(u3_u0__abc_75526_new_n589_));
AND2X2 AND2X2_3507 ( .A(u3_u0__abc_75526_new_n590_), .B(u3_u0__abc_75526_new_n588_), .Y(u3_u0__0r3_35_0__6_));
AND2X2 AND2X2_3508 ( .A(u3_u0__abc_75526_new_n563__bF_buf0), .B(u3_u0__abc_75526_new_n419_), .Y(u3_u0__abc_75526_new_n593_));
AND2X2 AND2X2_3509 ( .A(u3_u0__abc_75526_new_n594_), .B(u3_u0__abc_75526_new_n592_), .Y(u3_u0__0r3_35_0__7_));
AND2X2 AND2X2_351 ( .A(u0__abc_76628_new_n1170__bF_buf2), .B(sp_tms_18_), .Y(u0__abc_76628_new_n1610_));
AND2X2 AND2X2_3510 ( .A(u3_u0__abc_75526_new_n563__bF_buf6), .B(u3_u0__abc_75526_new_n424_), .Y(u3_u0__abc_75526_new_n597_));
AND2X2 AND2X2_3511 ( .A(u3_u0__abc_75526_new_n598_), .B(u3_u0__abc_75526_new_n596_), .Y(u3_u0__0r3_35_0__8_));
AND2X2 AND2X2_3512 ( .A(u3_u0__abc_75526_new_n563__bF_buf4), .B(u3_u0__abc_75526_new_n429_), .Y(u3_u0__abc_75526_new_n601_));
AND2X2 AND2X2_3513 ( .A(u3_u0__abc_75526_new_n602_), .B(u3_u0__abc_75526_new_n600_), .Y(u3_u0__0r3_35_0__9_));
AND2X2 AND2X2_3514 ( .A(u3_u0__abc_75526_new_n563__bF_buf2), .B(u3_u0__abc_75526_new_n434_), .Y(u3_u0__abc_75526_new_n605_));
AND2X2 AND2X2_3515 ( .A(u3_u0__abc_75526_new_n606_), .B(u3_u0__abc_75526_new_n604_), .Y(u3_u0__0r3_35_0__10_));
AND2X2 AND2X2_3516 ( .A(u3_u0__abc_75526_new_n563__bF_buf0), .B(u3_u0__abc_75526_new_n439_), .Y(u3_u0__abc_75526_new_n609_));
AND2X2 AND2X2_3517 ( .A(u3_u0__abc_75526_new_n610_), .B(u3_u0__abc_75526_new_n608_), .Y(u3_u0__0r3_35_0__11_));
AND2X2 AND2X2_3518 ( .A(u3_u0__abc_75526_new_n563__bF_buf6), .B(u3_u0__abc_75526_new_n444_), .Y(u3_u0__abc_75526_new_n613_));
AND2X2 AND2X2_3519 ( .A(u3_u0__abc_75526_new_n614_), .B(u3_u0__abc_75526_new_n612_), .Y(u3_u0__0r3_35_0__12_));
AND2X2 AND2X2_352 ( .A(spec_req_cs_5_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1611_));
AND2X2 AND2X2_3520 ( .A(u3_u0__abc_75526_new_n563__bF_buf4), .B(u3_u0__abc_75526_new_n449_), .Y(u3_u0__abc_75526_new_n617_));
AND2X2 AND2X2_3521 ( .A(u3_u0__abc_75526_new_n618_), .B(u3_u0__abc_75526_new_n616_), .Y(u3_u0__0r3_35_0__13_));
AND2X2 AND2X2_3522 ( .A(u3_u0__abc_75526_new_n563__bF_buf2), .B(u3_u0__abc_75526_new_n454_), .Y(u3_u0__abc_75526_new_n621_));
AND2X2 AND2X2_3523 ( .A(u3_u0__abc_75526_new_n622_), .B(u3_u0__abc_75526_new_n620_), .Y(u3_u0__0r3_35_0__14_));
AND2X2 AND2X2_3524 ( .A(u3_u0__abc_75526_new_n563__bF_buf0), .B(u3_u0__abc_75526_new_n459_), .Y(u3_u0__abc_75526_new_n625_));
AND2X2 AND2X2_3525 ( .A(u3_u0__abc_75526_new_n626_), .B(u3_u0__abc_75526_new_n624_), .Y(u3_u0__0r3_35_0__15_));
AND2X2 AND2X2_3526 ( .A(u3_u0__abc_75526_new_n563__bF_buf6), .B(u3_u0__abc_75526_new_n464_), .Y(u3_u0__abc_75526_new_n629_));
AND2X2 AND2X2_3527 ( .A(u3_u0__abc_75526_new_n630_), .B(u3_u0__abc_75526_new_n628_), .Y(u3_u0__0r3_35_0__16_));
AND2X2 AND2X2_3528 ( .A(u3_u0__abc_75526_new_n563__bF_buf4), .B(u3_u0__abc_75526_new_n469_), .Y(u3_u0__abc_75526_new_n633_));
AND2X2 AND2X2_3529 ( .A(u3_u0__abc_75526_new_n634_), .B(u3_u0__abc_75526_new_n632_), .Y(u3_u0__0r3_35_0__17_));
AND2X2 AND2X2_353 ( .A(u0__abc_76628_new_n1613_), .B(u0__abc_76628_new_n1179__bF_buf5), .Y(u0__abc_76628_new_n1614_));
AND2X2 AND2X2_3530 ( .A(u3_u0__abc_75526_new_n563__bF_buf2), .B(u3_u0__abc_75526_new_n474_), .Y(u3_u0__abc_75526_new_n637_));
AND2X2 AND2X2_3531 ( .A(u3_u0__abc_75526_new_n638_), .B(u3_u0__abc_75526_new_n636_), .Y(u3_u0__0r3_35_0__18_));
AND2X2 AND2X2_3532 ( .A(u3_u0__abc_75526_new_n563__bF_buf0), .B(u3_u0__abc_75526_new_n479_), .Y(u3_u0__abc_75526_new_n641_));
AND2X2 AND2X2_3533 ( .A(u3_u0__abc_75526_new_n642_), .B(u3_u0__abc_75526_new_n640_), .Y(u3_u0__0r3_35_0__19_));
AND2X2 AND2X2_3534 ( .A(u3_u0__abc_75526_new_n563__bF_buf6), .B(u3_u0__abc_75526_new_n484_), .Y(u3_u0__abc_75526_new_n645_));
AND2X2 AND2X2_3535 ( .A(u3_u0__abc_75526_new_n646_), .B(u3_u0__abc_75526_new_n644_), .Y(u3_u0__0r3_35_0__20_));
AND2X2 AND2X2_3536 ( .A(u3_u0__abc_75526_new_n563__bF_buf4), .B(u3_u0__abc_75526_new_n489_), .Y(u3_u0__abc_75526_new_n649_));
AND2X2 AND2X2_3537 ( .A(u3_u0__abc_75526_new_n650_), .B(u3_u0__abc_75526_new_n648_), .Y(u3_u0__0r3_35_0__21_));
AND2X2 AND2X2_3538 ( .A(u3_u0__abc_75526_new_n563__bF_buf2), .B(u3_u0__abc_75526_new_n494_), .Y(u3_u0__abc_75526_new_n653_));
AND2X2 AND2X2_3539 ( .A(u3_u0__abc_75526_new_n654_), .B(u3_u0__abc_75526_new_n652_), .Y(u3_u0__0r3_35_0__22_));
AND2X2 AND2X2_354 ( .A(u0__abc_76628_new_n1614_), .B(u0__abc_76628_new_n1612_), .Y(u0__abc_76628_new_n1615_));
AND2X2 AND2X2_3540 ( .A(u3_u0__abc_75526_new_n563__bF_buf0), .B(u3_u0__abc_75526_new_n499_), .Y(u3_u0__abc_75526_new_n657_));
AND2X2 AND2X2_3541 ( .A(u3_u0__abc_75526_new_n658_), .B(u3_u0__abc_75526_new_n656_), .Y(u3_u0__0r3_35_0__23_));
AND2X2 AND2X2_3542 ( .A(u3_u0__abc_75526_new_n563__bF_buf6), .B(u3_u0__abc_75526_new_n504_), .Y(u3_u0__abc_75526_new_n661_));
AND2X2 AND2X2_3543 ( .A(u3_u0__abc_75526_new_n662_), .B(u3_u0__abc_75526_new_n660_), .Y(u3_u0__0r3_35_0__24_));
AND2X2 AND2X2_3544 ( .A(u3_u0__abc_75526_new_n563__bF_buf4), .B(u3_u0__abc_75526_new_n509_), .Y(u3_u0__abc_75526_new_n665_));
AND2X2 AND2X2_3545 ( .A(u3_u0__abc_75526_new_n666_), .B(u3_u0__abc_75526_new_n664_), .Y(u3_u0__0r3_35_0__25_));
AND2X2 AND2X2_3546 ( .A(u3_u0__abc_75526_new_n563__bF_buf2), .B(u3_u0__abc_75526_new_n514_), .Y(u3_u0__abc_75526_new_n669_));
AND2X2 AND2X2_3547 ( .A(u3_u0__abc_75526_new_n670_), .B(u3_u0__abc_75526_new_n668_), .Y(u3_u0__0r3_35_0__26_));
AND2X2 AND2X2_3548 ( .A(u3_u0__abc_75526_new_n563__bF_buf0), .B(u3_u0__abc_75526_new_n519_), .Y(u3_u0__abc_75526_new_n673_));
AND2X2 AND2X2_3549 ( .A(u3_u0__abc_75526_new_n674_), .B(u3_u0__abc_75526_new_n672_), .Y(u3_u0__0r3_35_0__27_));
AND2X2 AND2X2_355 ( .A(u0__abc_76628_new_n1616_), .B(u0__abc_76628_new_n1175__bF_buf5), .Y(u0__abc_76628_new_n1617_));
AND2X2 AND2X2_3550 ( .A(u3_u0__abc_75526_new_n563__bF_buf6), .B(u3_u0__abc_75526_new_n524_), .Y(u3_u0__abc_75526_new_n677_));
AND2X2 AND2X2_3551 ( .A(u3_u0__abc_75526_new_n678_), .B(u3_u0__abc_75526_new_n676_), .Y(u3_u0__0r3_35_0__28_));
AND2X2 AND2X2_3552 ( .A(u3_u0__abc_75526_new_n563__bF_buf4), .B(u3_u0__abc_75526_new_n529_), .Y(u3_u0__abc_75526_new_n681_));
AND2X2 AND2X2_3553 ( .A(u3_u0__abc_75526_new_n682_), .B(u3_u0__abc_75526_new_n680_), .Y(u3_u0__0r3_35_0__29_));
AND2X2 AND2X2_3554 ( .A(u3_u0__abc_75526_new_n563__bF_buf2), .B(u3_u0__abc_75526_new_n534_), .Y(u3_u0__abc_75526_new_n685_));
AND2X2 AND2X2_3555 ( .A(u3_u0__abc_75526_new_n686_), .B(u3_u0__abc_75526_new_n684_), .Y(u3_u0__0r3_35_0__30_));
AND2X2 AND2X2_3556 ( .A(u3_u0__abc_75526_new_n563__bF_buf0), .B(u3_u0__abc_75526_new_n539_), .Y(u3_u0__abc_75526_new_n689_));
AND2X2 AND2X2_3557 ( .A(u3_u0__abc_75526_new_n690_), .B(u3_u0__abc_75526_new_n688_), .Y(u3_u0__0r3_35_0__31_));
AND2X2 AND2X2_3558 ( .A(u3_u0__abc_75526_new_n563__bF_buf6), .B(u3_u0__abc_75526_new_n544_), .Y(u3_u0__abc_75526_new_n693_));
AND2X2 AND2X2_3559 ( .A(u3_u0__abc_75526_new_n694_), .B(u3_u0__abc_75526_new_n692_), .Y(u3_u0__0r3_35_0__32_));
AND2X2 AND2X2_356 ( .A(spec_req_cs_4_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1618_));
AND2X2 AND2X2_3560 ( .A(u3_u0__abc_75526_new_n563__bF_buf4), .B(u3_u0__abc_75526_new_n549_), .Y(u3_u0__abc_75526_new_n697_));
AND2X2 AND2X2_3561 ( .A(u3_u0__abc_75526_new_n698_), .B(u3_u0__abc_75526_new_n696_), .Y(u3_u0__0r3_35_0__33_));
AND2X2 AND2X2_3562 ( .A(u3_u0__abc_75526_new_n563__bF_buf2), .B(u3_u0__abc_75526_new_n554_), .Y(u3_u0__abc_75526_new_n701_));
AND2X2 AND2X2_3563 ( .A(u3_u0__abc_75526_new_n702_), .B(u3_u0__abc_75526_new_n700_), .Y(u3_u0__0r3_35_0__34_));
AND2X2 AND2X2_3564 ( .A(u3_u0__abc_75526_new_n563__bF_buf0), .B(u3_u0__abc_75526_new_n559_), .Y(u3_u0__abc_75526_new_n705_));
AND2X2 AND2X2_3565 ( .A(u3_u0__abc_75526_new_n706_), .B(u3_u0__abc_75526_new_n704_), .Y(u3_u0__0r3_35_0__35_));
AND2X2 AND2X2_3566 ( .A(dv), .B(u3_u0_wr_adr_2_), .Y(u3_u0__abc_75526_new_n708_));
AND2X2 AND2X2_3567 ( .A(u3_u0__abc_75526_new_n708__bF_buf6), .B(u3_u0__abc_75526_new_n384_), .Y(u3_u0__abc_75526_new_n710_));
AND2X2 AND2X2_3568 ( .A(u3_u0__abc_75526_new_n711_), .B(u3_u0__abc_75526_new_n709_), .Y(u3_u0__0r2_35_0__0_));
AND2X2 AND2X2_3569 ( .A(u3_u0__abc_75526_new_n708__bF_buf4), .B(u3_u0__abc_75526_new_n389_), .Y(u3_u0__abc_75526_new_n714_));
AND2X2 AND2X2_357 ( .A(u0__abc_76628_new_n1619_), .B(u0__abc_76628_new_n1174__bF_buf5), .Y(u0__abc_76628_new_n1620_));
AND2X2 AND2X2_3570 ( .A(u3_u0__abc_75526_new_n715_), .B(u3_u0__abc_75526_new_n713_), .Y(u3_u0__0r2_35_0__1_));
AND2X2 AND2X2_3571 ( .A(u3_u0__abc_75526_new_n708__bF_buf2), .B(u3_u0__abc_75526_new_n394_), .Y(u3_u0__abc_75526_new_n718_));
AND2X2 AND2X2_3572 ( .A(u3_u0__abc_75526_new_n719_), .B(u3_u0__abc_75526_new_n717_), .Y(u3_u0__0r2_35_0__2_));
AND2X2 AND2X2_3573 ( .A(u3_u0__abc_75526_new_n708__bF_buf0), .B(u3_u0__abc_75526_new_n399_), .Y(u3_u0__abc_75526_new_n722_));
AND2X2 AND2X2_3574 ( .A(u3_u0__abc_75526_new_n723_), .B(u3_u0__abc_75526_new_n721_), .Y(u3_u0__0r2_35_0__3_));
AND2X2 AND2X2_3575 ( .A(u3_u0__abc_75526_new_n708__bF_buf6), .B(u3_u0__abc_75526_new_n404_), .Y(u3_u0__abc_75526_new_n726_));
AND2X2 AND2X2_3576 ( .A(u3_u0__abc_75526_new_n727_), .B(u3_u0__abc_75526_new_n725_), .Y(u3_u0__0r2_35_0__4_));
AND2X2 AND2X2_3577 ( .A(u3_u0__abc_75526_new_n708__bF_buf4), .B(u3_u0__abc_75526_new_n409_), .Y(u3_u0__abc_75526_new_n730_));
AND2X2 AND2X2_3578 ( .A(u3_u0__abc_75526_new_n731_), .B(u3_u0__abc_75526_new_n729_), .Y(u3_u0__0r2_35_0__5_));
AND2X2 AND2X2_3579 ( .A(u3_u0__abc_75526_new_n708__bF_buf2), .B(u3_u0__abc_75526_new_n414_), .Y(u3_u0__abc_75526_new_n734_));
AND2X2 AND2X2_358 ( .A(spec_req_cs_3_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1621_));
AND2X2 AND2X2_3580 ( .A(u3_u0__abc_75526_new_n735_), .B(u3_u0__abc_75526_new_n733_), .Y(u3_u0__0r2_35_0__6_));
AND2X2 AND2X2_3581 ( .A(u3_u0__abc_75526_new_n708__bF_buf0), .B(u3_u0__abc_75526_new_n419_), .Y(u3_u0__abc_75526_new_n738_));
AND2X2 AND2X2_3582 ( .A(u3_u0__abc_75526_new_n739_), .B(u3_u0__abc_75526_new_n737_), .Y(u3_u0__0r2_35_0__7_));
AND2X2 AND2X2_3583 ( .A(u3_u0__abc_75526_new_n708__bF_buf6), .B(u3_u0__abc_75526_new_n424_), .Y(u3_u0__abc_75526_new_n742_));
AND2X2 AND2X2_3584 ( .A(u3_u0__abc_75526_new_n743_), .B(u3_u0__abc_75526_new_n741_), .Y(u3_u0__0r2_35_0__8_));
AND2X2 AND2X2_3585 ( .A(u3_u0__abc_75526_new_n708__bF_buf4), .B(u3_u0__abc_75526_new_n429_), .Y(u3_u0__abc_75526_new_n746_));
AND2X2 AND2X2_3586 ( .A(u3_u0__abc_75526_new_n747_), .B(u3_u0__abc_75526_new_n745_), .Y(u3_u0__0r2_35_0__9_));
AND2X2 AND2X2_3587 ( .A(u3_u0__abc_75526_new_n708__bF_buf2), .B(u3_u0__abc_75526_new_n434_), .Y(u3_u0__abc_75526_new_n750_));
AND2X2 AND2X2_3588 ( .A(u3_u0__abc_75526_new_n751_), .B(u3_u0__abc_75526_new_n749_), .Y(u3_u0__0r2_35_0__10_));
AND2X2 AND2X2_3589 ( .A(u3_u0__abc_75526_new_n708__bF_buf0), .B(u3_u0__abc_75526_new_n439_), .Y(u3_u0__abc_75526_new_n754_));
AND2X2 AND2X2_359 ( .A(u0__abc_76628_new_n1622_), .B(u0__abc_76628_new_n1173__bF_buf5), .Y(u0__abc_76628_new_n1623_));
AND2X2 AND2X2_3590 ( .A(u3_u0__abc_75526_new_n755_), .B(u3_u0__abc_75526_new_n753_), .Y(u3_u0__0r2_35_0__11_));
AND2X2 AND2X2_3591 ( .A(u3_u0__abc_75526_new_n708__bF_buf6), .B(u3_u0__abc_75526_new_n444_), .Y(u3_u0__abc_75526_new_n758_));
AND2X2 AND2X2_3592 ( .A(u3_u0__abc_75526_new_n759_), .B(u3_u0__abc_75526_new_n757_), .Y(u3_u0__0r2_35_0__12_));
AND2X2 AND2X2_3593 ( .A(u3_u0__abc_75526_new_n708__bF_buf4), .B(u3_u0__abc_75526_new_n449_), .Y(u3_u0__abc_75526_new_n762_));
AND2X2 AND2X2_3594 ( .A(u3_u0__abc_75526_new_n763_), .B(u3_u0__abc_75526_new_n761_), .Y(u3_u0__0r2_35_0__13_));
AND2X2 AND2X2_3595 ( .A(u3_u0__abc_75526_new_n708__bF_buf2), .B(u3_u0__abc_75526_new_n454_), .Y(u3_u0__abc_75526_new_n766_));
AND2X2 AND2X2_3596 ( .A(u3_u0__abc_75526_new_n767_), .B(u3_u0__abc_75526_new_n765_), .Y(u3_u0__0r2_35_0__14_));
AND2X2 AND2X2_3597 ( .A(u3_u0__abc_75526_new_n708__bF_buf0), .B(u3_u0__abc_75526_new_n459_), .Y(u3_u0__abc_75526_new_n770_));
AND2X2 AND2X2_3598 ( .A(u3_u0__abc_75526_new_n771_), .B(u3_u0__abc_75526_new_n769_), .Y(u3_u0__0r2_35_0__15_));
AND2X2 AND2X2_3599 ( .A(u3_u0__abc_75526_new_n708__bF_buf6), .B(u3_u0__abc_75526_new_n464_), .Y(u3_u0__abc_75526_new_n774_));
AND2X2 AND2X2_36 ( .A(_abc_85006_new_n344_), .B(_abc_85006_new_n345_), .Y(tms_s_18_));
AND2X2 AND2X2_360 ( .A(spec_req_cs_2_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1624_));
AND2X2 AND2X2_3600 ( .A(u3_u0__abc_75526_new_n775_), .B(u3_u0__abc_75526_new_n773_), .Y(u3_u0__0r2_35_0__16_));
AND2X2 AND2X2_3601 ( .A(u3_u0__abc_75526_new_n708__bF_buf4), .B(u3_u0__abc_75526_new_n469_), .Y(u3_u0__abc_75526_new_n778_));
AND2X2 AND2X2_3602 ( .A(u3_u0__abc_75526_new_n779_), .B(u3_u0__abc_75526_new_n777_), .Y(u3_u0__0r2_35_0__17_));
AND2X2 AND2X2_3603 ( .A(u3_u0__abc_75526_new_n708__bF_buf2), .B(u3_u0__abc_75526_new_n474_), .Y(u3_u0__abc_75526_new_n782_));
AND2X2 AND2X2_3604 ( .A(u3_u0__abc_75526_new_n783_), .B(u3_u0__abc_75526_new_n781_), .Y(u3_u0__0r2_35_0__18_));
AND2X2 AND2X2_3605 ( .A(u3_u0__abc_75526_new_n708__bF_buf0), .B(u3_u0__abc_75526_new_n479_), .Y(u3_u0__abc_75526_new_n786_));
AND2X2 AND2X2_3606 ( .A(u3_u0__abc_75526_new_n787_), .B(u3_u0__abc_75526_new_n785_), .Y(u3_u0__0r2_35_0__19_));
AND2X2 AND2X2_3607 ( .A(u3_u0__abc_75526_new_n708__bF_buf6), .B(u3_u0__abc_75526_new_n484_), .Y(u3_u0__abc_75526_new_n790_));
AND2X2 AND2X2_3608 ( .A(u3_u0__abc_75526_new_n791_), .B(u3_u0__abc_75526_new_n789_), .Y(u3_u0__0r2_35_0__20_));
AND2X2 AND2X2_3609 ( .A(u3_u0__abc_75526_new_n708__bF_buf4), .B(u3_u0__abc_75526_new_n489_), .Y(u3_u0__abc_75526_new_n794_));
AND2X2 AND2X2_361 ( .A(u0__abc_76628_new_n1625_), .B(u0__abc_76628_new_n1172__bF_buf5), .Y(u0__abc_76628_new_n1626_));
AND2X2 AND2X2_3610 ( .A(u3_u0__abc_75526_new_n795_), .B(u3_u0__abc_75526_new_n793_), .Y(u3_u0__0r2_35_0__21_));
AND2X2 AND2X2_3611 ( .A(u3_u0__abc_75526_new_n708__bF_buf2), .B(u3_u0__abc_75526_new_n494_), .Y(u3_u0__abc_75526_new_n798_));
AND2X2 AND2X2_3612 ( .A(u3_u0__abc_75526_new_n799_), .B(u3_u0__abc_75526_new_n797_), .Y(u3_u0__0r2_35_0__22_));
AND2X2 AND2X2_3613 ( .A(u3_u0__abc_75526_new_n708__bF_buf0), .B(u3_u0__abc_75526_new_n499_), .Y(u3_u0__abc_75526_new_n802_));
AND2X2 AND2X2_3614 ( .A(u3_u0__abc_75526_new_n803_), .B(u3_u0__abc_75526_new_n801_), .Y(u3_u0__0r2_35_0__23_));
AND2X2 AND2X2_3615 ( .A(u3_u0__abc_75526_new_n708__bF_buf6), .B(u3_u0__abc_75526_new_n504_), .Y(u3_u0__abc_75526_new_n806_));
AND2X2 AND2X2_3616 ( .A(u3_u0__abc_75526_new_n807_), .B(u3_u0__abc_75526_new_n805_), .Y(u3_u0__0r2_35_0__24_));
AND2X2 AND2X2_3617 ( .A(u3_u0__abc_75526_new_n708__bF_buf4), .B(u3_u0__abc_75526_new_n509_), .Y(u3_u0__abc_75526_new_n810_));
AND2X2 AND2X2_3618 ( .A(u3_u0__abc_75526_new_n811_), .B(u3_u0__abc_75526_new_n809_), .Y(u3_u0__0r2_35_0__25_));
AND2X2 AND2X2_3619 ( .A(u3_u0__abc_75526_new_n708__bF_buf2), .B(u3_u0__abc_75526_new_n514_), .Y(u3_u0__abc_75526_new_n814_));
AND2X2 AND2X2_362 ( .A(spec_req_cs_1_bF_buf2_), .B(u0_tms1_18_), .Y(u0__abc_76628_new_n1627_));
AND2X2 AND2X2_3620 ( .A(u3_u0__abc_75526_new_n815_), .B(u3_u0__abc_75526_new_n813_), .Y(u3_u0__0r2_35_0__26_));
AND2X2 AND2X2_3621 ( .A(u3_u0__abc_75526_new_n708__bF_buf0), .B(u3_u0__abc_75526_new_n519_), .Y(u3_u0__abc_75526_new_n818_));
AND2X2 AND2X2_3622 ( .A(u3_u0__abc_75526_new_n819_), .B(u3_u0__abc_75526_new_n817_), .Y(u3_u0__0r2_35_0__27_));
AND2X2 AND2X2_3623 ( .A(u3_u0__abc_75526_new_n708__bF_buf6), .B(u3_u0__abc_75526_new_n524_), .Y(u3_u0__abc_75526_new_n822_));
AND2X2 AND2X2_3624 ( .A(u3_u0__abc_75526_new_n823_), .B(u3_u0__abc_75526_new_n821_), .Y(u3_u0__0r2_35_0__28_));
AND2X2 AND2X2_3625 ( .A(u3_u0__abc_75526_new_n708__bF_buf4), .B(u3_u0__abc_75526_new_n529_), .Y(u3_u0__abc_75526_new_n826_));
AND2X2 AND2X2_3626 ( .A(u3_u0__abc_75526_new_n827_), .B(u3_u0__abc_75526_new_n825_), .Y(u3_u0__0r2_35_0__29_));
AND2X2 AND2X2_3627 ( .A(u3_u0__abc_75526_new_n708__bF_buf2), .B(u3_u0__abc_75526_new_n534_), .Y(u3_u0__abc_75526_new_n830_));
AND2X2 AND2X2_3628 ( .A(u3_u0__abc_75526_new_n831_), .B(u3_u0__abc_75526_new_n829_), .Y(u3_u0__0r2_35_0__30_));
AND2X2 AND2X2_3629 ( .A(u3_u0__abc_75526_new_n708__bF_buf0), .B(u3_u0__abc_75526_new_n539_), .Y(u3_u0__abc_75526_new_n834_));
AND2X2 AND2X2_363 ( .A(u0__abc_76628_new_n1169__bF_buf1), .B(u0__abc_76628_new_n1630_), .Y(u0__abc_76628_new_n1631_));
AND2X2 AND2X2_3630 ( .A(u3_u0__abc_75526_new_n835_), .B(u3_u0__abc_75526_new_n833_), .Y(u3_u0__0r2_35_0__31_));
AND2X2 AND2X2_3631 ( .A(u3_u0__abc_75526_new_n708__bF_buf6), .B(u3_u0__abc_75526_new_n544_), .Y(u3_u0__abc_75526_new_n838_));
AND2X2 AND2X2_3632 ( .A(u3_u0__abc_75526_new_n839_), .B(u3_u0__abc_75526_new_n837_), .Y(u3_u0__0r2_35_0__32_));
AND2X2 AND2X2_3633 ( .A(u3_u0__abc_75526_new_n708__bF_buf4), .B(u3_u0__abc_75526_new_n549_), .Y(u3_u0__abc_75526_new_n842_));
AND2X2 AND2X2_3634 ( .A(u3_u0__abc_75526_new_n843_), .B(u3_u0__abc_75526_new_n841_), .Y(u3_u0__0r2_35_0__33_));
AND2X2 AND2X2_3635 ( .A(u3_u0__abc_75526_new_n708__bF_buf2), .B(u3_u0__abc_75526_new_n554_), .Y(u3_u0__abc_75526_new_n846_));
AND2X2 AND2X2_3636 ( .A(u3_u0__abc_75526_new_n847_), .B(u3_u0__abc_75526_new_n845_), .Y(u3_u0__0r2_35_0__34_));
AND2X2 AND2X2_3637 ( .A(u3_u0__abc_75526_new_n708__bF_buf0), .B(u3_u0__abc_75526_new_n559_), .Y(u3_u0__abc_75526_new_n850_));
AND2X2 AND2X2_3638 ( .A(u3_u0__abc_75526_new_n851_), .B(u3_u0__abc_75526_new_n849_), .Y(u3_u0__0r2_35_0__35_));
AND2X2 AND2X2_3639 ( .A(u3_u0__abc_75526_new_n853_), .B(u3_u0_rd_adr_0_), .Y(u3_u0__abc_75526_new_n854_));
AND2X2 AND2X2_364 ( .A(u0__abc_76628_new_n1629_), .B(u0__abc_76628_new_n1631_), .Y(u0__abc_76628_new_n1632_));
AND2X2 AND2X2_3640 ( .A(u3_u0_rd_adr_3_), .B(u3_re), .Y(u3_u0__abc_75526_new_n855_));
AND2X2 AND2X2_3641 ( .A(u3_u0_rd_adr_0_), .B(u3_re), .Y(u3_u0__abc_75526_new_n859_));
AND2X2 AND2X2_3642 ( .A(u3_u0__abc_75526_new_n853_), .B(u3_u0_rd_adr_1_), .Y(u3_u0__abc_75526_new_n860_));
AND2X2 AND2X2_3643 ( .A(u3_u0__abc_75526_new_n861_), .B(u3_u0__abc_75526_new_n858_), .Y(u3_u0__0rd_adr_3_0__1_));
AND2X2 AND2X2_3644 ( .A(u3_re), .B(u3_u0_rd_adr_1_), .Y(u3_u0__abc_75526_new_n863_));
AND2X2 AND2X2_3645 ( .A(u3_u0__abc_75526_new_n853_), .B(u3_u0_rd_adr_2_), .Y(u3_u0__abc_75526_new_n864_));
AND2X2 AND2X2_3646 ( .A(u3_u0__abc_75526_new_n865_), .B(u3_u0__abc_75526_new_n858_), .Y(u3_u0__0rd_adr_3_0__2_));
AND2X2 AND2X2_3647 ( .A(u3_re), .B(u3_u0_rd_adr_2_), .Y(u3_u0__abc_75526_new_n867_));
AND2X2 AND2X2_3648 ( .A(u3_u0__abc_75526_new_n853_), .B(u3_u0_rd_adr_3_), .Y(u3_u0__abc_75526_new_n868_));
AND2X2 AND2X2_3649 ( .A(u3_u0__abc_75526_new_n869_), .B(u3_u0__abc_75526_new_n858_), .Y(u3_u0__0rd_adr_3_0__3_));
AND2X2 AND2X2_365 ( .A(u0__abc_76628_new_n1170__bF_buf1), .B(sp_tms_19_), .Y(u0__abc_76628_new_n1634_));
AND2X2 AND2X2_3650 ( .A(u3_u0__abc_75526_new_n871_), .B(u3_u0_wr_adr_0_), .Y(u3_u0__abc_75526_new_n872_));
AND2X2 AND2X2_3651 ( .A(u3_u0__abc_75526_new_n871_), .B(u3_u0_wr_adr_1_), .Y(u3_u0__abc_75526_new_n875_));
AND2X2 AND2X2_3652 ( .A(dv), .B(u3_u0_wr_adr_0_), .Y(u3_u0__abc_75526_new_n876_));
AND2X2 AND2X2_3653 ( .A(u3_u0__abc_75526_new_n877_), .B(u3_u0__abc_75526_new_n858_), .Y(u3_u0__0wr_adr_3_0__1_));
AND2X2 AND2X2_3654 ( .A(u3_u0__abc_75526_new_n871_), .B(u3_u0_wr_adr_2_), .Y(u3_u0__abc_75526_new_n879_));
AND2X2 AND2X2_3655 ( .A(u3_u0__abc_75526_new_n880_), .B(u3_u0__abc_75526_new_n858_), .Y(u3_u0__0wr_adr_3_0__2_));
AND2X2 AND2X2_3656 ( .A(u3_u0__abc_75526_new_n871_), .B(u3_u0_wr_adr_3_), .Y(u3_u0__abc_75526_new_n882_));
AND2X2 AND2X2_3657 ( .A(u3_u0__abc_75526_new_n883_), .B(u3_u0__abc_75526_new_n858_), .Y(u3_u0__0wr_adr_3_0__3_));
AND2X2 AND2X2_3658 ( .A(u3_u0__abc_75526_new_n876__bF_buf5), .B(u3_u0__abc_75526_new_n384_), .Y(u3_u0__abc_75526_new_n886_));
AND2X2 AND2X2_3659 ( .A(u3_u0__abc_75526_new_n887_), .B(u3_u0__abc_75526_new_n885_), .Y(u3_u0__0r0_35_0__0_));
AND2X2 AND2X2_366 ( .A(spec_req_cs_5_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1635_));
AND2X2 AND2X2_3660 ( .A(u3_u0__abc_75526_new_n876__bF_buf3), .B(u3_u0__abc_75526_new_n389_), .Y(u3_u0__abc_75526_new_n890_));
AND2X2 AND2X2_3661 ( .A(u3_u0__abc_75526_new_n891_), .B(u3_u0__abc_75526_new_n889_), .Y(u3_u0__0r0_35_0__1_));
AND2X2 AND2X2_3662 ( .A(u3_u0__abc_75526_new_n876__bF_buf1), .B(u3_u0__abc_75526_new_n394_), .Y(u3_u0__abc_75526_new_n894_));
AND2X2 AND2X2_3663 ( .A(u3_u0__abc_75526_new_n895_), .B(u3_u0__abc_75526_new_n893_), .Y(u3_u0__0r0_35_0__2_));
AND2X2 AND2X2_3664 ( .A(u3_u0__abc_75526_new_n876__bF_buf7), .B(u3_u0__abc_75526_new_n399_), .Y(u3_u0__abc_75526_new_n898_));
AND2X2 AND2X2_3665 ( .A(u3_u0__abc_75526_new_n899_), .B(u3_u0__abc_75526_new_n897_), .Y(u3_u0__0r0_35_0__3_));
AND2X2 AND2X2_3666 ( .A(u3_u0__abc_75526_new_n876__bF_buf5), .B(u3_u0__abc_75526_new_n404_), .Y(u3_u0__abc_75526_new_n902_));
AND2X2 AND2X2_3667 ( .A(u3_u0__abc_75526_new_n903_), .B(u3_u0__abc_75526_new_n901_), .Y(u3_u0__0r0_35_0__4_));
AND2X2 AND2X2_3668 ( .A(u3_u0__abc_75526_new_n876__bF_buf3), .B(u3_u0__abc_75526_new_n409_), .Y(u3_u0__abc_75526_new_n906_));
AND2X2 AND2X2_3669 ( .A(u3_u0__abc_75526_new_n907_), .B(u3_u0__abc_75526_new_n905_), .Y(u3_u0__0r0_35_0__5_));
AND2X2 AND2X2_367 ( .A(u0__abc_76628_new_n1637_), .B(u0__abc_76628_new_n1179__bF_buf4), .Y(u0__abc_76628_new_n1638_));
AND2X2 AND2X2_3670 ( .A(u3_u0__abc_75526_new_n876__bF_buf1), .B(u3_u0__abc_75526_new_n414_), .Y(u3_u0__abc_75526_new_n910_));
AND2X2 AND2X2_3671 ( .A(u3_u0__abc_75526_new_n911_), .B(u3_u0__abc_75526_new_n909_), .Y(u3_u0__0r0_35_0__6_));
AND2X2 AND2X2_3672 ( .A(u3_u0__abc_75526_new_n876__bF_buf7), .B(u3_u0__abc_75526_new_n419_), .Y(u3_u0__abc_75526_new_n914_));
AND2X2 AND2X2_3673 ( .A(u3_u0__abc_75526_new_n915_), .B(u3_u0__abc_75526_new_n913_), .Y(u3_u0__0r0_35_0__7_));
AND2X2 AND2X2_3674 ( .A(u3_u0__abc_75526_new_n876__bF_buf5), .B(u3_u0__abc_75526_new_n424_), .Y(u3_u0__abc_75526_new_n918_));
AND2X2 AND2X2_3675 ( .A(u3_u0__abc_75526_new_n919_), .B(u3_u0__abc_75526_new_n917_), .Y(u3_u0__0r0_35_0__8_));
AND2X2 AND2X2_3676 ( .A(u3_u0__abc_75526_new_n876__bF_buf3), .B(u3_u0__abc_75526_new_n429_), .Y(u3_u0__abc_75526_new_n922_));
AND2X2 AND2X2_3677 ( .A(u3_u0__abc_75526_new_n923_), .B(u3_u0__abc_75526_new_n921_), .Y(u3_u0__0r0_35_0__9_));
AND2X2 AND2X2_3678 ( .A(u3_u0__abc_75526_new_n876__bF_buf1), .B(u3_u0__abc_75526_new_n434_), .Y(u3_u0__abc_75526_new_n926_));
AND2X2 AND2X2_3679 ( .A(u3_u0__abc_75526_new_n927_), .B(u3_u0__abc_75526_new_n925_), .Y(u3_u0__0r0_35_0__10_));
AND2X2 AND2X2_368 ( .A(u0__abc_76628_new_n1638_), .B(u0__abc_76628_new_n1636_), .Y(u0__abc_76628_new_n1639_));
AND2X2 AND2X2_3680 ( .A(u3_u0__abc_75526_new_n876__bF_buf7), .B(u3_u0__abc_75526_new_n439_), .Y(u3_u0__abc_75526_new_n930_));
AND2X2 AND2X2_3681 ( .A(u3_u0__abc_75526_new_n931_), .B(u3_u0__abc_75526_new_n929_), .Y(u3_u0__0r0_35_0__11_));
AND2X2 AND2X2_3682 ( .A(u3_u0__abc_75526_new_n876__bF_buf5), .B(u3_u0__abc_75526_new_n444_), .Y(u3_u0__abc_75526_new_n934_));
AND2X2 AND2X2_3683 ( .A(u3_u0__abc_75526_new_n935_), .B(u3_u0__abc_75526_new_n933_), .Y(u3_u0__0r0_35_0__12_));
AND2X2 AND2X2_3684 ( .A(u3_u0__abc_75526_new_n876__bF_buf3), .B(u3_u0__abc_75526_new_n449_), .Y(u3_u0__abc_75526_new_n938_));
AND2X2 AND2X2_3685 ( .A(u3_u0__abc_75526_new_n939_), .B(u3_u0__abc_75526_new_n937_), .Y(u3_u0__0r0_35_0__13_));
AND2X2 AND2X2_3686 ( .A(u3_u0__abc_75526_new_n876__bF_buf1), .B(u3_u0__abc_75526_new_n454_), .Y(u3_u0__abc_75526_new_n942_));
AND2X2 AND2X2_3687 ( .A(u3_u0__abc_75526_new_n943_), .B(u3_u0__abc_75526_new_n941_), .Y(u3_u0__0r0_35_0__14_));
AND2X2 AND2X2_3688 ( .A(u3_u0__abc_75526_new_n876__bF_buf7), .B(u3_u0__abc_75526_new_n459_), .Y(u3_u0__abc_75526_new_n946_));
AND2X2 AND2X2_3689 ( .A(u3_u0__abc_75526_new_n947_), .B(u3_u0__abc_75526_new_n945_), .Y(u3_u0__0r0_35_0__15_));
AND2X2 AND2X2_369 ( .A(u0__abc_76628_new_n1640_), .B(u0__abc_76628_new_n1175__bF_buf4), .Y(u0__abc_76628_new_n1641_));
AND2X2 AND2X2_3690 ( .A(u3_u0__abc_75526_new_n876__bF_buf5), .B(u3_u0__abc_75526_new_n464_), .Y(u3_u0__abc_75526_new_n950_));
AND2X2 AND2X2_3691 ( .A(u3_u0__abc_75526_new_n951_), .B(u3_u0__abc_75526_new_n949_), .Y(u3_u0__0r0_35_0__16_));
AND2X2 AND2X2_3692 ( .A(u3_u0__abc_75526_new_n876__bF_buf3), .B(u3_u0__abc_75526_new_n469_), .Y(u3_u0__abc_75526_new_n954_));
AND2X2 AND2X2_3693 ( .A(u3_u0__abc_75526_new_n955_), .B(u3_u0__abc_75526_new_n953_), .Y(u3_u0__0r0_35_0__17_));
AND2X2 AND2X2_3694 ( .A(u3_u0__abc_75526_new_n876__bF_buf1), .B(u3_u0__abc_75526_new_n474_), .Y(u3_u0__abc_75526_new_n958_));
AND2X2 AND2X2_3695 ( .A(u3_u0__abc_75526_new_n959_), .B(u3_u0__abc_75526_new_n957_), .Y(u3_u0__0r0_35_0__18_));
AND2X2 AND2X2_3696 ( .A(u3_u0__abc_75526_new_n876__bF_buf7), .B(u3_u0__abc_75526_new_n479_), .Y(u3_u0__abc_75526_new_n962_));
AND2X2 AND2X2_3697 ( .A(u3_u0__abc_75526_new_n963_), .B(u3_u0__abc_75526_new_n961_), .Y(u3_u0__0r0_35_0__19_));
AND2X2 AND2X2_3698 ( .A(u3_u0__abc_75526_new_n876__bF_buf5), .B(u3_u0__abc_75526_new_n484_), .Y(u3_u0__abc_75526_new_n966_));
AND2X2 AND2X2_3699 ( .A(u3_u0__abc_75526_new_n967_), .B(u3_u0__abc_75526_new_n965_), .Y(u3_u0__0r0_35_0__20_));
AND2X2 AND2X2_37 ( .A(_abc_85006_new_n347_), .B(_abc_85006_new_n348_), .Y(tms_s_19_));
AND2X2 AND2X2_370 ( .A(spec_req_cs_4_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1642_));
AND2X2 AND2X2_3700 ( .A(u3_u0__abc_75526_new_n876__bF_buf3), .B(u3_u0__abc_75526_new_n489_), .Y(u3_u0__abc_75526_new_n970_));
AND2X2 AND2X2_3701 ( .A(u3_u0__abc_75526_new_n971_), .B(u3_u0__abc_75526_new_n969_), .Y(u3_u0__0r0_35_0__21_));
AND2X2 AND2X2_3702 ( .A(u3_u0__abc_75526_new_n876__bF_buf1), .B(u3_u0__abc_75526_new_n494_), .Y(u3_u0__abc_75526_new_n974_));
AND2X2 AND2X2_3703 ( .A(u3_u0__abc_75526_new_n975_), .B(u3_u0__abc_75526_new_n973_), .Y(u3_u0__0r0_35_0__22_));
AND2X2 AND2X2_3704 ( .A(u3_u0__abc_75526_new_n876__bF_buf7), .B(u3_u0__abc_75526_new_n499_), .Y(u3_u0__abc_75526_new_n978_));
AND2X2 AND2X2_3705 ( .A(u3_u0__abc_75526_new_n979_), .B(u3_u0__abc_75526_new_n977_), .Y(u3_u0__0r0_35_0__23_));
AND2X2 AND2X2_3706 ( .A(u3_u0__abc_75526_new_n876__bF_buf5), .B(u3_u0__abc_75526_new_n504_), .Y(u3_u0__abc_75526_new_n982_));
AND2X2 AND2X2_3707 ( .A(u3_u0__abc_75526_new_n983_), .B(u3_u0__abc_75526_new_n981_), .Y(u3_u0__0r0_35_0__24_));
AND2X2 AND2X2_3708 ( .A(u3_u0__abc_75526_new_n876__bF_buf3), .B(u3_u0__abc_75526_new_n509_), .Y(u3_u0__abc_75526_new_n986_));
AND2X2 AND2X2_3709 ( .A(u3_u0__abc_75526_new_n987_), .B(u3_u0__abc_75526_new_n985_), .Y(u3_u0__0r0_35_0__25_));
AND2X2 AND2X2_371 ( .A(u0__abc_76628_new_n1643_), .B(u0__abc_76628_new_n1174__bF_buf4), .Y(u0__abc_76628_new_n1644_));
AND2X2 AND2X2_3710 ( .A(u3_u0__abc_75526_new_n876__bF_buf1), .B(u3_u0__abc_75526_new_n514_), .Y(u3_u0__abc_75526_new_n990_));
AND2X2 AND2X2_3711 ( .A(u3_u0__abc_75526_new_n991_), .B(u3_u0__abc_75526_new_n989_), .Y(u3_u0__0r0_35_0__26_));
AND2X2 AND2X2_3712 ( .A(u3_u0__abc_75526_new_n876__bF_buf7), .B(u3_u0__abc_75526_new_n519_), .Y(u3_u0__abc_75526_new_n994_));
AND2X2 AND2X2_3713 ( .A(u3_u0__abc_75526_new_n995_), .B(u3_u0__abc_75526_new_n993_), .Y(u3_u0__0r0_35_0__27_));
AND2X2 AND2X2_3714 ( .A(u3_u0__abc_75526_new_n876__bF_buf5), .B(u3_u0__abc_75526_new_n524_), .Y(u3_u0__abc_75526_new_n998_));
AND2X2 AND2X2_3715 ( .A(u3_u0__abc_75526_new_n999_), .B(u3_u0__abc_75526_new_n997_), .Y(u3_u0__0r0_35_0__28_));
AND2X2 AND2X2_3716 ( .A(u3_u0__abc_75526_new_n876__bF_buf3), .B(u3_u0__abc_75526_new_n529_), .Y(u3_u0__abc_75526_new_n1002_));
AND2X2 AND2X2_3717 ( .A(u3_u0__abc_75526_new_n1003_), .B(u3_u0__abc_75526_new_n1001_), .Y(u3_u0__0r0_35_0__29_));
AND2X2 AND2X2_3718 ( .A(u3_u0__abc_75526_new_n876__bF_buf1), .B(u3_u0__abc_75526_new_n534_), .Y(u3_u0__abc_75526_new_n1006_));
AND2X2 AND2X2_3719 ( .A(u3_u0__abc_75526_new_n1007_), .B(u3_u0__abc_75526_new_n1005_), .Y(u3_u0__0r0_35_0__30_));
AND2X2 AND2X2_372 ( .A(spec_req_cs_3_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1645_));
AND2X2 AND2X2_3720 ( .A(u3_u0__abc_75526_new_n876__bF_buf7), .B(u3_u0__abc_75526_new_n539_), .Y(u3_u0__abc_75526_new_n1010_));
AND2X2 AND2X2_3721 ( .A(u3_u0__abc_75526_new_n1011_), .B(u3_u0__abc_75526_new_n1009_), .Y(u3_u0__0r0_35_0__31_));
AND2X2 AND2X2_3722 ( .A(u3_u0__abc_75526_new_n876__bF_buf5), .B(u3_u0__abc_75526_new_n544_), .Y(u3_u0__abc_75526_new_n1014_));
AND2X2 AND2X2_3723 ( .A(u3_u0__abc_75526_new_n1015_), .B(u3_u0__abc_75526_new_n1013_), .Y(u3_u0__0r0_35_0__32_));
AND2X2 AND2X2_3724 ( .A(u3_u0__abc_75526_new_n876__bF_buf3), .B(u3_u0__abc_75526_new_n549_), .Y(u3_u0__abc_75526_new_n1018_));
AND2X2 AND2X2_3725 ( .A(u3_u0__abc_75526_new_n1019_), .B(u3_u0__abc_75526_new_n1017_), .Y(u3_u0__0r0_35_0__33_));
AND2X2 AND2X2_3726 ( .A(u3_u0__abc_75526_new_n876__bF_buf1), .B(u3_u0__abc_75526_new_n554_), .Y(u3_u0__abc_75526_new_n1022_));
AND2X2 AND2X2_3727 ( .A(u3_u0__abc_75526_new_n1023_), .B(u3_u0__abc_75526_new_n1021_), .Y(u3_u0__0r0_35_0__34_));
AND2X2 AND2X2_3728 ( .A(u3_u0__abc_75526_new_n876__bF_buf7), .B(u3_u0__abc_75526_new_n559_), .Y(u3_u0__abc_75526_new_n1026_));
AND2X2 AND2X2_3729 ( .A(u3_u0__abc_75526_new_n1027_), .B(u3_u0__abc_75526_new_n1025_), .Y(u3_u0__0r0_35_0__35_));
AND2X2 AND2X2_373 ( .A(u0__abc_76628_new_n1646_), .B(u0__abc_76628_new_n1173__bF_buf4), .Y(u0__abc_76628_new_n1647_));
AND2X2 AND2X2_3730 ( .A(u3_u0__abc_75526_new_n1029_), .B(u3_u0__abc_75526_new_n1030_), .Y(u3_u0__abc_75526_new_n1031_));
AND2X2 AND2X2_3731 ( .A(u3_u0__abc_75526_new_n1032_), .B(u3_u0_rd_adr_3_), .Y(u3_u0__abc_75526_new_n1033_));
AND2X2 AND2X2_3732 ( .A(u3_u0__abc_75526_new_n1031_), .B(u3_u0__abc_75526_new_n1033_), .Y(u3_u0__abc_75526_new_n1034_));
AND2X2 AND2X2_3733 ( .A(u3_u0__abc_75526_new_n1038_), .B(u3_u0__abc_75526_new_n1041_), .Y(u3_u0__abc_75526_new_n1042_));
AND2X2 AND2X2_3734 ( .A(u3_u0__abc_75526_new_n1042_), .B(u3_u0__abc_75526_new_n1035_), .Y(u3_u0__abc_75526_new_n1043_));
AND2X2 AND2X2_3735 ( .A(u3_u0__abc_75526_new_n1043__bF_buf5), .B(u3_u0_r0_0_), .Y(u3_u0__abc_75526_new_n1044_));
AND2X2 AND2X2_3736 ( .A(u3_u0__abc_75526_new_n1034__bF_buf4), .B(u3_u0_r3_0_), .Y(u3_u0__abc_75526_new_n1045_));
AND2X2 AND2X2_3737 ( .A(u3_u0__abc_75526_new_n1029_), .B(u3_u0__abc_75526_new_n1046_), .Y(u3_u0__abc_75526_new_n1047_));
AND2X2 AND2X2_3738 ( .A(u3_u0__abc_75526_new_n1032_), .B(u3_u0_rd_adr_1_), .Y(u3_u0__abc_75526_new_n1048_));
AND2X2 AND2X2_3739 ( .A(u3_u0__abc_75526_new_n1047_), .B(u3_u0__abc_75526_new_n1048_), .Y(u3_u0__abc_75526_new_n1049_));
AND2X2 AND2X2_374 ( .A(spec_req_cs_2_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1648_));
AND2X2 AND2X2_3740 ( .A(u3_u0__abc_75526_new_n1049__bF_buf5), .B(u3_u0_r1_0_), .Y(u3_u0__abc_75526_new_n1050_));
AND2X2 AND2X2_3741 ( .A(u3_u0__abc_75526_new_n1046_), .B(u3_u0_rd_adr_2_), .Y(u3_u0__abc_75526_new_n1051_));
AND2X2 AND2X2_3742 ( .A(u3_u0__abc_75526_new_n1031_), .B(u3_u0__abc_75526_new_n1051_), .Y(u3_u0__abc_75526_new_n1052_));
AND2X2 AND2X2_3743 ( .A(u3_u0__abc_75526_new_n1052__bF_buf5), .B(u3_u0_r2_0_), .Y(u3_u0__abc_75526_new_n1053_));
AND2X2 AND2X2_3744 ( .A(u3_u0__abc_75526_new_n1043__bF_buf4), .B(u3_u0_r0_1_), .Y(u3_u0__abc_75526_new_n1057_));
AND2X2 AND2X2_3745 ( .A(u3_u0__abc_75526_new_n1034__bF_buf3), .B(u3_u0_r3_1_), .Y(u3_u0__abc_75526_new_n1058_));
AND2X2 AND2X2_3746 ( .A(u3_u0__abc_75526_new_n1049__bF_buf4), .B(u3_u0_r1_1_), .Y(u3_u0__abc_75526_new_n1059_));
AND2X2 AND2X2_3747 ( .A(u3_u0__abc_75526_new_n1052__bF_buf4), .B(u3_u0_r2_1_), .Y(u3_u0__abc_75526_new_n1060_));
AND2X2 AND2X2_3748 ( .A(u3_u0__abc_75526_new_n1043__bF_buf3), .B(u3_u0_r0_2_), .Y(u3_u0__abc_75526_new_n1064_));
AND2X2 AND2X2_3749 ( .A(u3_u0__abc_75526_new_n1034__bF_buf2), .B(u3_u0_r3_2_), .Y(u3_u0__abc_75526_new_n1065_));
AND2X2 AND2X2_375 ( .A(u0__abc_76628_new_n1649_), .B(u0__abc_76628_new_n1172__bF_buf4), .Y(u0__abc_76628_new_n1650_));
AND2X2 AND2X2_3750 ( .A(u3_u0__abc_75526_new_n1049__bF_buf3), .B(u3_u0_r1_2_), .Y(u3_u0__abc_75526_new_n1066_));
AND2X2 AND2X2_3751 ( .A(u3_u0__abc_75526_new_n1052__bF_buf3), .B(u3_u0_r2_2_), .Y(u3_u0__abc_75526_new_n1067_));
AND2X2 AND2X2_3752 ( .A(u3_u0__abc_75526_new_n1043__bF_buf2), .B(u3_u0_r0_3_), .Y(u3_u0__abc_75526_new_n1071_));
AND2X2 AND2X2_3753 ( .A(u3_u0__abc_75526_new_n1034__bF_buf1), .B(u3_u0_r3_3_), .Y(u3_u0__abc_75526_new_n1072_));
AND2X2 AND2X2_3754 ( .A(u3_u0__abc_75526_new_n1049__bF_buf2), .B(u3_u0_r1_3_), .Y(u3_u0__abc_75526_new_n1073_));
AND2X2 AND2X2_3755 ( .A(u3_u0__abc_75526_new_n1052__bF_buf2), .B(u3_u0_r2_3_), .Y(u3_u0__abc_75526_new_n1074_));
AND2X2 AND2X2_3756 ( .A(u3_u0__abc_75526_new_n1043__bF_buf1), .B(u3_u0_r0_4_), .Y(u3_u0__abc_75526_new_n1078_));
AND2X2 AND2X2_3757 ( .A(u3_u0__abc_75526_new_n1034__bF_buf0), .B(u3_u0_r3_4_), .Y(u3_u0__abc_75526_new_n1079_));
AND2X2 AND2X2_3758 ( .A(u3_u0__abc_75526_new_n1049__bF_buf1), .B(u3_u0_r1_4_), .Y(u3_u0__abc_75526_new_n1080_));
AND2X2 AND2X2_3759 ( .A(u3_u0__abc_75526_new_n1052__bF_buf1), .B(u3_u0_r2_4_), .Y(u3_u0__abc_75526_new_n1081_));
AND2X2 AND2X2_376 ( .A(spec_req_cs_1_bF_buf1_), .B(u0_tms1_19_), .Y(u0__abc_76628_new_n1651_));
AND2X2 AND2X2_3760 ( .A(u3_u0__abc_75526_new_n1043__bF_buf0), .B(u3_u0_r0_5_), .Y(u3_u0__abc_75526_new_n1085_));
AND2X2 AND2X2_3761 ( .A(u3_u0__abc_75526_new_n1034__bF_buf5), .B(u3_u0_r3_5_), .Y(u3_u0__abc_75526_new_n1086_));
AND2X2 AND2X2_3762 ( .A(u3_u0__abc_75526_new_n1049__bF_buf0), .B(u3_u0_r1_5_), .Y(u3_u0__abc_75526_new_n1087_));
AND2X2 AND2X2_3763 ( .A(u3_u0__abc_75526_new_n1052__bF_buf0), .B(u3_u0_r2_5_), .Y(u3_u0__abc_75526_new_n1088_));
AND2X2 AND2X2_3764 ( .A(u3_u0__abc_75526_new_n1043__bF_buf5), .B(u3_u0_r0_6_), .Y(u3_u0__abc_75526_new_n1092_));
AND2X2 AND2X2_3765 ( .A(u3_u0__abc_75526_new_n1034__bF_buf4), .B(u3_u0_r3_6_), .Y(u3_u0__abc_75526_new_n1093_));
AND2X2 AND2X2_3766 ( .A(u3_u0__abc_75526_new_n1049__bF_buf5), .B(u3_u0_r1_6_), .Y(u3_u0__abc_75526_new_n1094_));
AND2X2 AND2X2_3767 ( .A(u3_u0__abc_75526_new_n1052__bF_buf5), .B(u3_u0_r2_6_), .Y(u3_u0__abc_75526_new_n1095_));
AND2X2 AND2X2_3768 ( .A(u3_u0__abc_75526_new_n1043__bF_buf4), .B(u3_u0_r0_7_), .Y(u3_u0__abc_75526_new_n1099_));
AND2X2 AND2X2_3769 ( .A(u3_u0__abc_75526_new_n1034__bF_buf3), .B(u3_u0_r3_7_), .Y(u3_u0__abc_75526_new_n1100_));
AND2X2 AND2X2_377 ( .A(u0__abc_76628_new_n1169__bF_buf0), .B(u0__abc_76628_new_n1654_), .Y(u0__abc_76628_new_n1655_));
AND2X2 AND2X2_3770 ( .A(u3_u0__abc_75526_new_n1049__bF_buf4), .B(u3_u0_r1_7_), .Y(u3_u0__abc_75526_new_n1101_));
AND2X2 AND2X2_3771 ( .A(u3_u0__abc_75526_new_n1052__bF_buf4), .B(u3_u0_r2_7_), .Y(u3_u0__abc_75526_new_n1102_));
AND2X2 AND2X2_3772 ( .A(u3_u0__abc_75526_new_n1043__bF_buf3), .B(u3_u0_r0_8_), .Y(u3_u0__abc_75526_new_n1106_));
AND2X2 AND2X2_3773 ( .A(u3_u0__abc_75526_new_n1034__bF_buf2), .B(u3_u0_r3_8_), .Y(u3_u0__abc_75526_new_n1107_));
AND2X2 AND2X2_3774 ( .A(u3_u0__abc_75526_new_n1049__bF_buf3), .B(u3_u0_r1_8_), .Y(u3_u0__abc_75526_new_n1108_));
AND2X2 AND2X2_3775 ( .A(u3_u0__abc_75526_new_n1052__bF_buf3), .B(u3_u0_r2_8_), .Y(u3_u0__abc_75526_new_n1109_));
AND2X2 AND2X2_3776 ( .A(u3_u0__abc_75526_new_n1043__bF_buf2), .B(u3_u0_r0_9_), .Y(u3_u0__abc_75526_new_n1113_));
AND2X2 AND2X2_3777 ( .A(u3_u0__abc_75526_new_n1034__bF_buf1), .B(u3_u0_r3_9_), .Y(u3_u0__abc_75526_new_n1114_));
AND2X2 AND2X2_3778 ( .A(u3_u0__abc_75526_new_n1049__bF_buf2), .B(u3_u0_r1_9_), .Y(u3_u0__abc_75526_new_n1115_));
AND2X2 AND2X2_3779 ( .A(u3_u0__abc_75526_new_n1052__bF_buf2), .B(u3_u0_r2_9_), .Y(u3_u0__abc_75526_new_n1116_));
AND2X2 AND2X2_378 ( .A(u0__abc_76628_new_n1653_), .B(u0__abc_76628_new_n1655_), .Y(u0__abc_76628_new_n1656_));
AND2X2 AND2X2_3780 ( .A(u3_u0__abc_75526_new_n1043__bF_buf1), .B(u3_u0_r0_10_), .Y(u3_u0__abc_75526_new_n1120_));
AND2X2 AND2X2_3781 ( .A(u3_u0__abc_75526_new_n1034__bF_buf0), .B(u3_u0_r3_10_), .Y(u3_u0__abc_75526_new_n1121_));
AND2X2 AND2X2_3782 ( .A(u3_u0__abc_75526_new_n1049__bF_buf1), .B(u3_u0_r1_10_), .Y(u3_u0__abc_75526_new_n1122_));
AND2X2 AND2X2_3783 ( .A(u3_u0__abc_75526_new_n1052__bF_buf1), .B(u3_u0_r2_10_), .Y(u3_u0__abc_75526_new_n1123_));
AND2X2 AND2X2_3784 ( .A(u3_u0__abc_75526_new_n1043__bF_buf0), .B(u3_u0_r0_11_), .Y(u3_u0__abc_75526_new_n1127_));
AND2X2 AND2X2_3785 ( .A(u3_u0__abc_75526_new_n1034__bF_buf5), .B(u3_u0_r3_11_), .Y(u3_u0__abc_75526_new_n1128_));
AND2X2 AND2X2_3786 ( .A(u3_u0__abc_75526_new_n1049__bF_buf0), .B(u3_u0_r1_11_), .Y(u3_u0__abc_75526_new_n1129_));
AND2X2 AND2X2_3787 ( .A(u3_u0__abc_75526_new_n1052__bF_buf0), .B(u3_u0_r2_11_), .Y(u3_u0__abc_75526_new_n1130_));
AND2X2 AND2X2_3788 ( .A(u3_u0__abc_75526_new_n1043__bF_buf5), .B(u3_u0_r0_12_), .Y(u3_u0__abc_75526_new_n1134_));
AND2X2 AND2X2_3789 ( .A(u3_u0__abc_75526_new_n1034__bF_buf4), .B(u3_u0_r3_12_), .Y(u3_u0__abc_75526_new_n1135_));
AND2X2 AND2X2_379 ( .A(u0__abc_76628_new_n1170__bF_buf0), .B(sp_tms_20_), .Y(u0__abc_76628_new_n1658_));
AND2X2 AND2X2_3790 ( .A(u3_u0__abc_75526_new_n1049__bF_buf5), .B(u3_u0_r1_12_), .Y(u3_u0__abc_75526_new_n1136_));
AND2X2 AND2X2_3791 ( .A(u3_u0__abc_75526_new_n1052__bF_buf5), .B(u3_u0_r2_12_), .Y(u3_u0__abc_75526_new_n1137_));
AND2X2 AND2X2_3792 ( .A(u3_u0__abc_75526_new_n1043__bF_buf4), .B(u3_u0_r0_13_), .Y(u3_u0__abc_75526_new_n1141_));
AND2X2 AND2X2_3793 ( .A(u3_u0__abc_75526_new_n1034__bF_buf3), .B(u3_u0_r3_13_), .Y(u3_u0__abc_75526_new_n1142_));
AND2X2 AND2X2_3794 ( .A(u3_u0__abc_75526_new_n1049__bF_buf4), .B(u3_u0_r1_13_), .Y(u3_u0__abc_75526_new_n1143_));
AND2X2 AND2X2_3795 ( .A(u3_u0__abc_75526_new_n1052__bF_buf4), .B(u3_u0_r2_13_), .Y(u3_u0__abc_75526_new_n1144_));
AND2X2 AND2X2_3796 ( .A(u3_u0__abc_75526_new_n1043__bF_buf3), .B(u3_u0_r0_14_), .Y(u3_u0__abc_75526_new_n1148_));
AND2X2 AND2X2_3797 ( .A(u3_u0__abc_75526_new_n1034__bF_buf2), .B(u3_u0_r3_14_), .Y(u3_u0__abc_75526_new_n1149_));
AND2X2 AND2X2_3798 ( .A(u3_u0__abc_75526_new_n1049__bF_buf3), .B(u3_u0_r1_14_), .Y(u3_u0__abc_75526_new_n1150_));
AND2X2 AND2X2_3799 ( .A(u3_u0__abc_75526_new_n1052__bF_buf3), .B(u3_u0_r2_14_), .Y(u3_u0__abc_75526_new_n1151_));
AND2X2 AND2X2_38 ( .A(_abc_85006_new_n350_), .B(_abc_85006_new_n351_), .Y(tms_s_20_));
AND2X2 AND2X2_380 ( .A(spec_req_cs_5_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1659_));
AND2X2 AND2X2_3800 ( .A(u3_u0__abc_75526_new_n1043__bF_buf2), .B(u3_u0_r0_15_), .Y(u3_u0__abc_75526_new_n1155_));
AND2X2 AND2X2_3801 ( .A(u3_u0__abc_75526_new_n1034__bF_buf1), .B(u3_u0_r3_15_), .Y(u3_u0__abc_75526_new_n1156_));
AND2X2 AND2X2_3802 ( .A(u3_u0__abc_75526_new_n1049__bF_buf2), .B(u3_u0_r1_15_), .Y(u3_u0__abc_75526_new_n1157_));
AND2X2 AND2X2_3803 ( .A(u3_u0__abc_75526_new_n1052__bF_buf2), .B(u3_u0_r2_15_), .Y(u3_u0__abc_75526_new_n1158_));
AND2X2 AND2X2_3804 ( .A(u3_u0__abc_75526_new_n1043__bF_buf1), .B(u3_u0_r0_16_), .Y(u3_u0__abc_75526_new_n1162_));
AND2X2 AND2X2_3805 ( .A(u3_u0__abc_75526_new_n1034__bF_buf0), .B(u3_u0_r3_16_), .Y(u3_u0__abc_75526_new_n1163_));
AND2X2 AND2X2_3806 ( .A(u3_u0__abc_75526_new_n1049__bF_buf1), .B(u3_u0_r1_16_), .Y(u3_u0__abc_75526_new_n1164_));
AND2X2 AND2X2_3807 ( .A(u3_u0__abc_75526_new_n1052__bF_buf1), .B(u3_u0_r2_16_), .Y(u3_u0__abc_75526_new_n1165_));
AND2X2 AND2X2_3808 ( .A(u3_u0__abc_75526_new_n1043__bF_buf0), .B(u3_u0_r0_17_), .Y(u3_u0__abc_75526_new_n1169_));
AND2X2 AND2X2_3809 ( .A(u3_u0__abc_75526_new_n1034__bF_buf5), .B(u3_u0_r3_17_), .Y(u3_u0__abc_75526_new_n1170_));
AND2X2 AND2X2_381 ( .A(u0__abc_76628_new_n1661_), .B(u0__abc_76628_new_n1179__bF_buf3), .Y(u0__abc_76628_new_n1662_));
AND2X2 AND2X2_3810 ( .A(u3_u0__abc_75526_new_n1049__bF_buf0), .B(u3_u0_r1_17_), .Y(u3_u0__abc_75526_new_n1171_));
AND2X2 AND2X2_3811 ( .A(u3_u0__abc_75526_new_n1052__bF_buf0), .B(u3_u0_r2_17_), .Y(u3_u0__abc_75526_new_n1172_));
AND2X2 AND2X2_3812 ( .A(u3_u0__abc_75526_new_n1043__bF_buf5), .B(u3_u0_r0_18_), .Y(u3_u0__abc_75526_new_n1176_));
AND2X2 AND2X2_3813 ( .A(u3_u0__abc_75526_new_n1034__bF_buf4), .B(u3_u0_r3_18_), .Y(u3_u0__abc_75526_new_n1177_));
AND2X2 AND2X2_3814 ( .A(u3_u0__abc_75526_new_n1049__bF_buf5), .B(u3_u0_r1_18_), .Y(u3_u0__abc_75526_new_n1178_));
AND2X2 AND2X2_3815 ( .A(u3_u0__abc_75526_new_n1052__bF_buf5), .B(u3_u0_r2_18_), .Y(u3_u0__abc_75526_new_n1179_));
AND2X2 AND2X2_3816 ( .A(u3_u0__abc_75526_new_n1043__bF_buf4), .B(u3_u0_r0_19_), .Y(u3_u0__abc_75526_new_n1183_));
AND2X2 AND2X2_3817 ( .A(u3_u0__abc_75526_new_n1034__bF_buf3), .B(u3_u0_r3_19_), .Y(u3_u0__abc_75526_new_n1184_));
AND2X2 AND2X2_3818 ( .A(u3_u0__abc_75526_new_n1049__bF_buf4), .B(u3_u0_r1_19_), .Y(u3_u0__abc_75526_new_n1185_));
AND2X2 AND2X2_3819 ( .A(u3_u0__abc_75526_new_n1052__bF_buf4), .B(u3_u0_r2_19_), .Y(u3_u0__abc_75526_new_n1186_));
AND2X2 AND2X2_382 ( .A(u0__abc_76628_new_n1662_), .B(u0__abc_76628_new_n1660_), .Y(u0__abc_76628_new_n1663_));
AND2X2 AND2X2_3820 ( .A(u3_u0__abc_75526_new_n1043__bF_buf3), .B(u3_u0_r0_20_), .Y(u3_u0__abc_75526_new_n1190_));
AND2X2 AND2X2_3821 ( .A(u3_u0__abc_75526_new_n1034__bF_buf2), .B(u3_u0_r3_20_), .Y(u3_u0__abc_75526_new_n1191_));
AND2X2 AND2X2_3822 ( .A(u3_u0__abc_75526_new_n1049__bF_buf3), .B(u3_u0_r1_20_), .Y(u3_u0__abc_75526_new_n1192_));
AND2X2 AND2X2_3823 ( .A(u3_u0__abc_75526_new_n1052__bF_buf3), .B(u3_u0_r2_20_), .Y(u3_u0__abc_75526_new_n1193_));
AND2X2 AND2X2_3824 ( .A(u3_u0__abc_75526_new_n1043__bF_buf2), .B(u3_u0_r0_21_), .Y(u3_u0__abc_75526_new_n1197_));
AND2X2 AND2X2_3825 ( .A(u3_u0__abc_75526_new_n1034__bF_buf1), .B(u3_u0_r3_21_), .Y(u3_u0__abc_75526_new_n1198_));
AND2X2 AND2X2_3826 ( .A(u3_u0__abc_75526_new_n1049__bF_buf2), .B(u3_u0_r1_21_), .Y(u3_u0__abc_75526_new_n1199_));
AND2X2 AND2X2_3827 ( .A(u3_u0__abc_75526_new_n1052__bF_buf2), .B(u3_u0_r2_21_), .Y(u3_u0__abc_75526_new_n1200_));
AND2X2 AND2X2_3828 ( .A(u3_u0__abc_75526_new_n1043__bF_buf1), .B(u3_u0_r0_22_), .Y(u3_u0__abc_75526_new_n1204_));
AND2X2 AND2X2_3829 ( .A(u3_u0__abc_75526_new_n1034__bF_buf0), .B(u3_u0_r3_22_), .Y(u3_u0__abc_75526_new_n1205_));
AND2X2 AND2X2_383 ( .A(u0__abc_76628_new_n1664_), .B(u0__abc_76628_new_n1175__bF_buf3), .Y(u0__abc_76628_new_n1665_));
AND2X2 AND2X2_3830 ( .A(u3_u0__abc_75526_new_n1049__bF_buf1), .B(u3_u0_r1_22_), .Y(u3_u0__abc_75526_new_n1206_));
AND2X2 AND2X2_3831 ( .A(u3_u0__abc_75526_new_n1052__bF_buf1), .B(u3_u0_r2_22_), .Y(u3_u0__abc_75526_new_n1207_));
AND2X2 AND2X2_3832 ( .A(u3_u0__abc_75526_new_n1043__bF_buf0), .B(u3_u0_r0_23_), .Y(u3_u0__abc_75526_new_n1211_));
AND2X2 AND2X2_3833 ( .A(u3_u0__abc_75526_new_n1034__bF_buf5), .B(u3_u0_r3_23_), .Y(u3_u0__abc_75526_new_n1212_));
AND2X2 AND2X2_3834 ( .A(u3_u0__abc_75526_new_n1049__bF_buf0), .B(u3_u0_r1_23_), .Y(u3_u0__abc_75526_new_n1213_));
AND2X2 AND2X2_3835 ( .A(u3_u0__abc_75526_new_n1052__bF_buf0), .B(u3_u0_r2_23_), .Y(u3_u0__abc_75526_new_n1214_));
AND2X2 AND2X2_3836 ( .A(u3_u0__abc_75526_new_n1043__bF_buf5), .B(u3_u0_r0_24_), .Y(u3_u0__abc_75526_new_n1218_));
AND2X2 AND2X2_3837 ( .A(u3_u0__abc_75526_new_n1034__bF_buf4), .B(u3_u0_r3_24_), .Y(u3_u0__abc_75526_new_n1219_));
AND2X2 AND2X2_3838 ( .A(u3_u0__abc_75526_new_n1049__bF_buf5), .B(u3_u0_r1_24_), .Y(u3_u0__abc_75526_new_n1220_));
AND2X2 AND2X2_3839 ( .A(u3_u0__abc_75526_new_n1052__bF_buf5), .B(u3_u0_r2_24_), .Y(u3_u0__abc_75526_new_n1221_));
AND2X2 AND2X2_384 ( .A(spec_req_cs_4_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1666_));
AND2X2 AND2X2_3840 ( .A(u3_u0__abc_75526_new_n1043__bF_buf4), .B(u3_u0_r0_25_), .Y(u3_u0__abc_75526_new_n1225_));
AND2X2 AND2X2_3841 ( .A(u3_u0__abc_75526_new_n1034__bF_buf3), .B(u3_u0_r3_25_), .Y(u3_u0__abc_75526_new_n1226_));
AND2X2 AND2X2_3842 ( .A(u3_u0__abc_75526_new_n1049__bF_buf4), .B(u3_u0_r1_25_), .Y(u3_u0__abc_75526_new_n1227_));
AND2X2 AND2X2_3843 ( .A(u3_u0__abc_75526_new_n1052__bF_buf4), .B(u3_u0_r2_25_), .Y(u3_u0__abc_75526_new_n1228_));
AND2X2 AND2X2_3844 ( .A(u3_u0__abc_75526_new_n1043__bF_buf3), .B(u3_u0_r0_26_), .Y(u3_u0__abc_75526_new_n1232_));
AND2X2 AND2X2_3845 ( .A(u3_u0__abc_75526_new_n1034__bF_buf2), .B(u3_u0_r3_26_), .Y(u3_u0__abc_75526_new_n1233_));
AND2X2 AND2X2_3846 ( .A(u3_u0__abc_75526_new_n1049__bF_buf3), .B(u3_u0_r1_26_), .Y(u3_u0__abc_75526_new_n1234_));
AND2X2 AND2X2_3847 ( .A(u3_u0__abc_75526_new_n1052__bF_buf3), .B(u3_u0_r2_26_), .Y(u3_u0__abc_75526_new_n1235_));
AND2X2 AND2X2_3848 ( .A(u3_u0__abc_75526_new_n1043__bF_buf2), .B(u3_u0_r0_27_), .Y(u3_u0__abc_75526_new_n1239_));
AND2X2 AND2X2_3849 ( .A(u3_u0__abc_75526_new_n1034__bF_buf1), .B(u3_u0_r3_27_), .Y(u3_u0__abc_75526_new_n1240_));
AND2X2 AND2X2_385 ( .A(u0__abc_76628_new_n1667_), .B(u0__abc_76628_new_n1174__bF_buf3), .Y(u0__abc_76628_new_n1668_));
AND2X2 AND2X2_3850 ( .A(u3_u0__abc_75526_new_n1049__bF_buf2), .B(u3_u0_r1_27_), .Y(u3_u0__abc_75526_new_n1241_));
AND2X2 AND2X2_3851 ( .A(u3_u0__abc_75526_new_n1052__bF_buf2), .B(u3_u0_r2_27_), .Y(u3_u0__abc_75526_new_n1242_));
AND2X2 AND2X2_3852 ( .A(u3_u0__abc_75526_new_n1043__bF_buf1), .B(u3_u0_r0_28_), .Y(u3_u0__abc_75526_new_n1246_));
AND2X2 AND2X2_3853 ( .A(u3_u0__abc_75526_new_n1034__bF_buf0), .B(u3_u0_r3_28_), .Y(u3_u0__abc_75526_new_n1247_));
AND2X2 AND2X2_3854 ( .A(u3_u0__abc_75526_new_n1049__bF_buf1), .B(u3_u0_r1_28_), .Y(u3_u0__abc_75526_new_n1248_));
AND2X2 AND2X2_3855 ( .A(u3_u0__abc_75526_new_n1052__bF_buf1), .B(u3_u0_r2_28_), .Y(u3_u0__abc_75526_new_n1249_));
AND2X2 AND2X2_3856 ( .A(u3_u0__abc_75526_new_n1043__bF_buf0), .B(u3_u0_r0_29_), .Y(u3_u0__abc_75526_new_n1253_));
AND2X2 AND2X2_3857 ( .A(u3_u0__abc_75526_new_n1034__bF_buf5), .B(u3_u0_r3_29_), .Y(u3_u0__abc_75526_new_n1254_));
AND2X2 AND2X2_3858 ( .A(u3_u0__abc_75526_new_n1049__bF_buf0), .B(u3_u0_r1_29_), .Y(u3_u0__abc_75526_new_n1255_));
AND2X2 AND2X2_3859 ( .A(u3_u0__abc_75526_new_n1052__bF_buf0), .B(u3_u0_r2_29_), .Y(u3_u0__abc_75526_new_n1256_));
AND2X2 AND2X2_386 ( .A(spec_req_cs_3_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1669_));
AND2X2 AND2X2_3860 ( .A(u3_u0__abc_75526_new_n1043__bF_buf5), .B(u3_u0_r0_30_), .Y(u3_u0__abc_75526_new_n1260_));
AND2X2 AND2X2_3861 ( .A(u3_u0__abc_75526_new_n1034__bF_buf4), .B(u3_u0_r3_30_), .Y(u3_u0__abc_75526_new_n1261_));
AND2X2 AND2X2_3862 ( .A(u3_u0__abc_75526_new_n1049__bF_buf5), .B(u3_u0_r1_30_), .Y(u3_u0__abc_75526_new_n1262_));
AND2X2 AND2X2_3863 ( .A(u3_u0__abc_75526_new_n1052__bF_buf5), .B(u3_u0_r2_30_), .Y(u3_u0__abc_75526_new_n1263_));
AND2X2 AND2X2_3864 ( .A(u3_u0__abc_75526_new_n1043__bF_buf4), .B(u3_u0_r0_31_), .Y(u3_u0__abc_75526_new_n1267_));
AND2X2 AND2X2_3865 ( .A(u3_u0__abc_75526_new_n1034__bF_buf3), .B(u3_u0_r3_31_), .Y(u3_u0__abc_75526_new_n1268_));
AND2X2 AND2X2_3866 ( .A(u3_u0__abc_75526_new_n1049__bF_buf4), .B(u3_u0_r1_31_), .Y(u3_u0__abc_75526_new_n1269_));
AND2X2 AND2X2_3867 ( .A(u3_u0__abc_75526_new_n1052__bF_buf4), .B(u3_u0_r2_31_), .Y(u3_u0__abc_75526_new_n1270_));
AND2X2 AND2X2_3868 ( .A(u3_u0__abc_75526_new_n1043__bF_buf3), .B(u3_u0_r0_32_), .Y(u3_u0__abc_75526_new_n1274_));
AND2X2 AND2X2_3869 ( .A(u3_u0__abc_75526_new_n1034__bF_buf2), .B(u3_u0_r3_32_), .Y(u3_u0__abc_75526_new_n1275_));
AND2X2 AND2X2_387 ( .A(u0__abc_76628_new_n1670_), .B(u0__abc_76628_new_n1173__bF_buf3), .Y(u0__abc_76628_new_n1671_));
AND2X2 AND2X2_3870 ( .A(u3_u0__abc_75526_new_n1049__bF_buf3), .B(u3_u0_r1_32_), .Y(u3_u0__abc_75526_new_n1276_));
AND2X2 AND2X2_3871 ( .A(u3_u0__abc_75526_new_n1052__bF_buf3), .B(u3_u0_r2_32_), .Y(u3_u0__abc_75526_new_n1277_));
AND2X2 AND2X2_3872 ( .A(u3_u0__abc_75526_new_n1043__bF_buf2), .B(u3_u0_r0_33_), .Y(u3_u0__abc_75526_new_n1281_));
AND2X2 AND2X2_3873 ( .A(u3_u0__abc_75526_new_n1034__bF_buf1), .B(u3_u0_r3_33_), .Y(u3_u0__abc_75526_new_n1282_));
AND2X2 AND2X2_3874 ( .A(u3_u0__abc_75526_new_n1049__bF_buf2), .B(u3_u0_r1_33_), .Y(u3_u0__abc_75526_new_n1283_));
AND2X2 AND2X2_3875 ( .A(u3_u0__abc_75526_new_n1052__bF_buf2), .B(u3_u0_r2_33_), .Y(u3_u0__abc_75526_new_n1284_));
AND2X2 AND2X2_3876 ( .A(u3_u0__abc_75526_new_n1043__bF_buf1), .B(u3_u0_r0_34_), .Y(u3_u0__abc_75526_new_n1288_));
AND2X2 AND2X2_3877 ( .A(u3_u0__abc_75526_new_n1034__bF_buf0), .B(u3_u0_r3_34_), .Y(u3_u0__abc_75526_new_n1289_));
AND2X2 AND2X2_3878 ( .A(u3_u0__abc_75526_new_n1049__bF_buf1), .B(u3_u0_r1_34_), .Y(u3_u0__abc_75526_new_n1290_));
AND2X2 AND2X2_3879 ( .A(u3_u0__abc_75526_new_n1052__bF_buf1), .B(u3_u0_r2_34_), .Y(u3_u0__abc_75526_new_n1291_));
AND2X2 AND2X2_388 ( .A(spec_req_cs_2_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1672_));
AND2X2 AND2X2_3880 ( .A(u3_u0__abc_75526_new_n1043__bF_buf0), .B(u3_u0_r0_35_), .Y(u3_u0__abc_75526_new_n1295_));
AND2X2 AND2X2_3881 ( .A(u3_u0__abc_75526_new_n1034__bF_buf5), .B(u3_u0_r3_35_), .Y(u3_u0__abc_75526_new_n1296_));
AND2X2 AND2X2_3882 ( .A(u3_u0__abc_75526_new_n1049__bF_buf0), .B(u3_u0_r1_35_), .Y(u3_u0__abc_75526_new_n1297_));
AND2X2 AND2X2_3883 ( .A(u3_u0__abc_75526_new_n1052__bF_buf0), .B(u3_u0_r2_35_), .Y(u3_u0__abc_75526_new_n1298_));
AND2X2 AND2X2_3884 ( .A(u4_ps_cnt_3_), .B(rfr_ps_val_3_), .Y(u4__abc_76448_new_n73_));
AND2X2 AND2X2_3885 ( .A(u4__abc_76448_new_n74_), .B(u4__abc_76448_new_n72_), .Y(u4__abc_76448_new_n75_));
AND2X2 AND2X2_3886 ( .A(u4_ps_cnt_2_), .B(rfr_ps_val_2_), .Y(u4__abc_76448_new_n77_));
AND2X2 AND2X2_3887 ( .A(u4__abc_76448_new_n78_), .B(u4__abc_76448_new_n76_), .Y(u4__abc_76448_new_n79_));
AND2X2 AND2X2_3888 ( .A(u4_ps_cnt_7_), .B(rfr_ps_val_7_), .Y(u4__abc_76448_new_n82_));
AND2X2 AND2X2_3889 ( .A(u4__abc_76448_new_n83_), .B(u4__abc_76448_new_n81_), .Y(u4__abc_76448_new_n84_));
AND2X2 AND2X2_389 ( .A(u0__abc_76628_new_n1673_), .B(u0__abc_76628_new_n1172__bF_buf3), .Y(u0__abc_76628_new_n1674_));
AND2X2 AND2X2_3890 ( .A(u4_ps_cnt_6_), .B(rfr_ps_val_6_), .Y(u4__abc_76448_new_n86_));
AND2X2 AND2X2_3891 ( .A(u4__abc_76448_new_n87_), .B(u4__abc_76448_new_n85_), .Y(u4__abc_76448_new_n88_));
AND2X2 AND2X2_3892 ( .A(u4__abc_76448_new_n91_), .B(u4_ps_cnt_0_), .Y(u4__abc_76448_new_n92_));
AND2X2 AND2X2_3893 ( .A(u4__abc_76448_new_n93_), .B(rfr_ps_val_0_), .Y(u4__abc_76448_new_n94_));
AND2X2 AND2X2_3894 ( .A(u4__abc_76448_new_n96_), .B(u4_ps_cnt_1_), .Y(u4__abc_76448_new_n97_));
AND2X2 AND2X2_3895 ( .A(u4__abc_76448_new_n98_), .B(rfr_ps_val_1_), .Y(u4__abc_76448_new_n99_));
AND2X2 AND2X2_3896 ( .A(u4__abc_76448_new_n102_), .B(u4_ps_cnt_4_), .Y(u4__abc_76448_new_n103_));
AND2X2 AND2X2_3897 ( .A(u4__abc_76448_new_n104_), .B(rfr_ps_val_4_), .Y(u4__abc_76448_new_n105_));
AND2X2 AND2X2_3898 ( .A(u4__abc_76448_new_n107_), .B(rfr_ps_val_5_), .Y(u4__abc_76448_new_n108_));
AND2X2 AND2X2_3899 ( .A(u4__abc_76448_new_n109_), .B(u4_ps_cnt_5_), .Y(u4__abc_76448_new_n110_));
AND2X2 AND2X2_39 ( .A(_abc_85006_new_n353_), .B(_abc_85006_new_n354_), .Y(tms_s_21_));
AND2X2 AND2X2_390 ( .A(spec_req_cs_1_bF_buf0_), .B(u0_tms1_20_), .Y(u0__abc_76628_new_n1675_));
AND2X2 AND2X2_3900 ( .A(u4__abc_76448_new_n117_), .B(u4__abc_76448_new_n116_), .Y(u4__0rfr_req_0_0_));
AND2X2 AND2X2_3901 ( .A(u4_rfr_ce), .B(u4_rfr_cnt_0_), .Y(u4__abc_76448_new_n119_));
AND2X2 AND2X2_3902 ( .A(u4__abc_76448_new_n121_), .B(u4__abc_76448_new_n116_), .Y(u4__abc_76448_new_n122_));
AND2X2 AND2X2_3903 ( .A(u4__abc_76448_new_n122_), .B(u4__abc_76448_new_n120_), .Y(u4__0rfr_cnt_7_0__0_));
AND2X2 AND2X2_3904 ( .A(u4__abc_76448_new_n119_), .B(u4_rfr_cnt_1_), .Y(u4__abc_76448_new_n124_));
AND2X2 AND2X2_3905 ( .A(u4__abc_76448_new_n126_), .B(u4__abc_76448_new_n116_), .Y(u4__abc_76448_new_n127_));
AND2X2 AND2X2_3906 ( .A(u4__abc_76448_new_n127_), .B(u4__abc_76448_new_n125_), .Y(u4__0rfr_cnt_7_0__1_));
AND2X2 AND2X2_3907 ( .A(u4_rfr_cnt_0_), .B(u4_rfr_cnt_1_), .Y(u4__abc_76448_new_n129_));
AND2X2 AND2X2_3908 ( .A(u4__abc_76448_new_n129_), .B(u4_rfr_cnt_2_), .Y(u4__abc_76448_new_n130_));
AND2X2 AND2X2_3909 ( .A(u4__abc_76448_new_n130_), .B(u4_rfr_ce), .Y(u4__abc_76448_new_n131_));
AND2X2 AND2X2_391 ( .A(u0__abc_76628_new_n1169__bF_buf6), .B(u0__abc_76628_new_n1678_), .Y(u0__abc_76628_new_n1679_));
AND2X2 AND2X2_3910 ( .A(u4__abc_76448_new_n133_), .B(u4__abc_76448_new_n116_), .Y(u4__abc_76448_new_n134_));
AND2X2 AND2X2_3911 ( .A(u4__abc_76448_new_n134_), .B(u4__abc_76448_new_n132_), .Y(u4__0rfr_cnt_7_0__2_));
AND2X2 AND2X2_3912 ( .A(u4__abc_76448_new_n130_), .B(u4_rfr_cnt_3_), .Y(u4__abc_76448_new_n136_));
AND2X2 AND2X2_3913 ( .A(u4__abc_76448_new_n136_), .B(u4_rfr_ce), .Y(u4__abc_76448_new_n137_));
AND2X2 AND2X2_3914 ( .A(u4__abc_76448_new_n139_), .B(u4__abc_76448_new_n116_), .Y(u4__abc_76448_new_n140_));
AND2X2 AND2X2_3915 ( .A(u4__abc_76448_new_n140_), .B(u4__abc_76448_new_n138_), .Y(u4__0rfr_cnt_7_0__3_));
AND2X2 AND2X2_3916 ( .A(u4_rfr_cnt_3_), .B(u4_rfr_cnt_4_), .Y(u4__abc_76448_new_n143_));
AND2X2 AND2X2_3917 ( .A(u4__abc_76448_new_n130_), .B(u4__abc_76448_new_n143_), .Y(u4__abc_76448_new_n144_));
AND2X2 AND2X2_3918 ( .A(u4__abc_76448_new_n144_), .B(u4_rfr_ce), .Y(u4__abc_76448_new_n145_));
AND2X2 AND2X2_3919 ( .A(u4__abc_76448_new_n146_), .B(u4__abc_76448_new_n116_), .Y(u4__abc_76448_new_n147_));
AND2X2 AND2X2_392 ( .A(u0__abc_76628_new_n1677_), .B(u0__abc_76628_new_n1679_), .Y(u0__abc_76628_new_n1680_));
AND2X2 AND2X2_3920 ( .A(u4__abc_76448_new_n147_), .B(u4__abc_76448_new_n142_), .Y(u4__0rfr_cnt_7_0__4_));
AND2X2 AND2X2_3921 ( .A(u4__abc_76448_new_n144_), .B(u4_rfr_cnt_5_), .Y(u4__abc_76448_new_n149_));
AND2X2 AND2X2_3922 ( .A(u4__abc_76448_new_n149_), .B(u4_rfr_ce), .Y(u4__abc_76448_new_n150_));
AND2X2 AND2X2_3923 ( .A(u4__abc_76448_new_n152_), .B(u4__abc_76448_new_n116_), .Y(u4__abc_76448_new_n153_));
AND2X2 AND2X2_3924 ( .A(u4__abc_76448_new_n153_), .B(u4__abc_76448_new_n151_), .Y(u4__0rfr_cnt_7_0__5_));
AND2X2 AND2X2_3925 ( .A(u4_rfr_cnt_5_), .B(u4_rfr_cnt_6_), .Y(u4__abc_76448_new_n156_));
AND2X2 AND2X2_3926 ( .A(u4__abc_76448_new_n145_), .B(u4__abc_76448_new_n156_), .Y(u4__abc_76448_new_n157_));
AND2X2 AND2X2_3927 ( .A(u4__abc_76448_new_n158_), .B(u4__abc_76448_new_n116_), .Y(u4__abc_76448_new_n159_));
AND2X2 AND2X2_3928 ( .A(u4__abc_76448_new_n159_), .B(u4__abc_76448_new_n155_), .Y(u4__0rfr_cnt_7_0__6_));
AND2X2 AND2X2_3929 ( .A(u4__abc_76448_new_n157_), .B(u4_rfr_cnt_7_), .Y(u4__abc_76448_new_n161_));
AND2X2 AND2X2_393 ( .A(u0__abc_76628_new_n1170__bF_buf6), .B(sp_tms_21_), .Y(u0__abc_76628_new_n1682_));
AND2X2 AND2X2_3930 ( .A(u4__abc_76448_new_n163_), .B(u4__abc_76448_new_n116_), .Y(u4__abc_76448_new_n164_));
AND2X2 AND2X2_3931 ( .A(u4__abc_76448_new_n164_), .B(u4__abc_76448_new_n162_), .Y(u4__0rfr_cnt_7_0__7_));
AND2X2 AND2X2_3932 ( .A(u4__abc_76448_new_n102_), .B(u4__abc_76448_new_n109_), .Y(u4__abc_76448_new_n166_));
AND2X2 AND2X2_3933 ( .A(u4__abc_76448_new_n167_), .B(u4__abc_76448_new_n168_), .Y(u4__abc_76448_new_n169_));
AND2X2 AND2X2_3934 ( .A(u4__abc_76448_new_n166_), .B(u4__abc_76448_new_n169_), .Y(u4__abc_76448_new_n170_));
AND2X2 AND2X2_3935 ( .A(u4__abc_76448_new_n91_), .B(u4__abc_76448_new_n96_), .Y(u4__abc_76448_new_n171_));
AND2X2 AND2X2_3936 ( .A(u4__abc_76448_new_n172_), .B(u4__abc_76448_new_n173_), .Y(u4__abc_76448_new_n174_));
AND2X2 AND2X2_3937 ( .A(u4__abc_76448_new_n171_), .B(u4__abc_76448_new_n174_), .Y(u4__abc_76448_new_n175_));
AND2X2 AND2X2_3938 ( .A(u4__abc_76448_new_n170_), .B(u4__abc_76448_new_n175_), .Y(u4__abc_76448_new_n176_));
AND2X2 AND2X2_3939 ( .A(u4_ps_cnt_0_), .B(u4_rfr_en), .Y(u4__abc_76448_new_n179_));
AND2X2 AND2X2_394 ( .A(spec_req_cs_5_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1683_));
AND2X2 AND2X2_3940 ( .A(u4__abc_76448_new_n180_), .B(u4__abc_76448_new_n181_), .Y(u4__abc_76448_new_n182_));
AND2X2 AND2X2_3941 ( .A(u4__abc_76448_new_n177_), .B(u4__abc_76448_new_n182_), .Y(u4__0ps_cnt_7_0__0_));
AND2X2 AND2X2_3942 ( .A(u4__abc_76448_new_n179_), .B(u4_ps_cnt_1_), .Y(u4__abc_76448_new_n184_));
AND2X2 AND2X2_3943 ( .A(u4__abc_76448_new_n185_), .B(u4__abc_76448_new_n186_), .Y(u4__abc_76448_new_n187_));
AND2X2 AND2X2_3944 ( .A(u4__abc_76448_new_n177_), .B(u4__abc_76448_new_n187_), .Y(u4__0ps_cnt_7_0__1_));
AND2X2 AND2X2_3945 ( .A(u4__abc_76448_new_n184_), .B(u4_ps_cnt_2_), .Y(u4__abc_76448_new_n190_));
AND2X2 AND2X2_3946 ( .A(u4__abc_76448_new_n191_), .B(u4__abc_76448_new_n189_), .Y(u4__abc_76448_new_n192_));
AND2X2 AND2X2_3947 ( .A(u4__abc_76448_new_n177_), .B(u4__abc_76448_new_n192_), .Y(u4__0ps_cnt_7_0__2_));
AND2X2 AND2X2_3948 ( .A(u4__abc_76448_new_n190_), .B(u4_ps_cnt_3_), .Y(u4__abc_76448_new_n195_));
AND2X2 AND2X2_3949 ( .A(u4__abc_76448_new_n196_), .B(u4__abc_76448_new_n194_), .Y(u4__abc_76448_new_n197_));
AND2X2 AND2X2_395 ( .A(u0__abc_76628_new_n1685_), .B(u0__abc_76628_new_n1179__bF_buf2), .Y(u0__abc_76628_new_n1686_));
AND2X2 AND2X2_3950 ( .A(u4__abc_76448_new_n177_), .B(u4__abc_76448_new_n197_), .Y(u4__0ps_cnt_7_0__3_));
AND2X2 AND2X2_3951 ( .A(u4__abc_76448_new_n195_), .B(u4_ps_cnt_4_), .Y(u4__abc_76448_new_n200_));
AND2X2 AND2X2_3952 ( .A(u4__abc_76448_new_n201_), .B(u4__abc_76448_new_n199_), .Y(u4__abc_76448_new_n202_));
AND2X2 AND2X2_3953 ( .A(u4__abc_76448_new_n177_), .B(u4__abc_76448_new_n202_), .Y(u4__0ps_cnt_7_0__4_));
AND2X2 AND2X2_3954 ( .A(u4_ps_cnt_3_), .B(u4_ps_cnt_4_), .Y(u4__abc_76448_new_n204_));
AND2X2 AND2X2_3955 ( .A(u4__abc_76448_new_n204_), .B(u4_ps_cnt_5_), .Y(u4__abc_76448_new_n205_));
AND2X2 AND2X2_3956 ( .A(u4__abc_76448_new_n190_), .B(u4__abc_76448_new_n205_), .Y(u4__abc_76448_new_n206_));
AND2X2 AND2X2_3957 ( .A(u4__abc_76448_new_n208_), .B(u4__abc_76448_new_n207_), .Y(u4__abc_76448_new_n209_));
AND2X2 AND2X2_3958 ( .A(u4__abc_76448_new_n177_), .B(u4__abc_76448_new_n209_), .Y(u4__0ps_cnt_7_0__5_));
AND2X2 AND2X2_3959 ( .A(u4__abc_76448_new_n206_), .B(u4__abc_76448_new_n211_), .Y(u4__abc_76448_new_n212_));
AND2X2 AND2X2_396 ( .A(u0__abc_76628_new_n1686_), .B(u0__abc_76628_new_n1684_), .Y(u0__abc_76628_new_n1687_));
AND2X2 AND2X2_3960 ( .A(u4__abc_76448_new_n207_), .B(u4_ps_cnt_6_), .Y(u4__abc_76448_new_n213_));
AND2X2 AND2X2_3961 ( .A(u4__abc_76448_new_n177_), .B(u4__abc_76448_new_n214_), .Y(u4__0ps_cnt_7_0__6_));
AND2X2 AND2X2_3962 ( .A(u4__abc_76448_new_n206_), .B(u4_ps_cnt_6_), .Y(u4__abc_76448_new_n216_));
AND2X2 AND2X2_3963 ( .A(u4__abc_76448_new_n216_), .B(u4_ps_cnt_7_), .Y(u4__abc_76448_new_n217_));
AND2X2 AND2X2_3964 ( .A(u4__abc_76448_new_n218_), .B(u4__abc_76448_new_n219_), .Y(u4__abc_76448_new_n220_));
AND2X2 AND2X2_3965 ( .A(u4__abc_76448_new_n220_), .B(u4__abc_76448_new_n177_), .Y(u4__0ps_cnt_7_0__7_));
AND2X2 AND2X2_3966 ( .A(u4__abc_76448_new_n224_), .B(ref_int_1_), .Y(u4__abc_76448_new_n225_));
AND2X2 AND2X2_3967 ( .A(u4__abc_76448_new_n225_), .B(u4__abc_76448_new_n130_), .Y(u4__abc_76448_new_n226_));
AND2X2 AND2X2_3968 ( .A(u4__abc_76448_new_n228_), .B(u4_rfr_cnt_0_), .Y(u4__abc_76448_new_n229_));
AND2X2 AND2X2_3969 ( .A(u4__abc_76448_new_n227_), .B(u4__abc_76448_new_n229_), .Y(u4__abc_76448_new_n230_));
AND2X2 AND2X2_397 ( .A(u0__abc_76628_new_n1688_), .B(u0__abc_76628_new_n1175__bF_buf2), .Y(u0__abc_76628_new_n1689_));
AND2X2 AND2X2_3970 ( .A(u4__abc_76448_new_n231_), .B(u4__abc_76448_new_n222_), .Y(u4__abc_76448_new_n232_));
AND2X2 AND2X2_3971 ( .A(u4__abc_76448_new_n233_), .B(u4__abc_76448_new_n228_), .Y(u4__abc_76448_new_n234_));
AND2X2 AND2X2_3972 ( .A(u4_rfr_cnt_7_), .B(ref_int_1_), .Y(u4__abc_76448_new_n235_));
AND2X2 AND2X2_3973 ( .A(u4__abc_76448_new_n236_), .B(u4__abc_76448_new_n156_), .Y(u4__abc_76448_new_n237_));
AND2X2 AND2X2_3974 ( .A(u4__abc_76448_new_n144_), .B(ref_int_2_), .Y(u4__abc_76448_new_n239_));
AND2X2 AND2X2_3975 ( .A(u4__abc_76448_new_n238_), .B(u4__abc_76448_new_n239_), .Y(u4__abc_76448_new_n240_));
AND2X2 AND2X2_3976 ( .A(u4__abc_76448_new_n241_), .B(u4_rfr_early), .Y(u4__0rfr_clr_0_0_));
AND2X2 AND2X2_3977 ( .A(u5__abc_81276_new_n368_), .B(u5__abc_81276_new_n369_), .Y(u5__abc_81276_new_n370_));
AND2X2 AND2X2_3978 ( .A(u5__abc_81276_new_n370_), .B(u5__abc_81276_new_n367_), .Y(u5__abc_81276_new_n371_));
AND2X2 AND2X2_3979 ( .A(u5__abc_81276_new_n371_), .B(u5__abc_81276_new_n366_), .Y(u5__abc_81276_new_n372_));
AND2X2 AND2X2_398 ( .A(spec_req_cs_4_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1690_));
AND2X2 AND2X2_3980 ( .A(u5__abc_81276_new_n373_), .B(u5__abc_81276_new_n374_), .Y(u5__abc_81276_new_n375_));
AND2X2 AND2X2_3981 ( .A(u5__abc_81276_new_n376_), .B(u5__abc_81276_new_n377_), .Y(u5__abc_81276_new_n378_));
AND2X2 AND2X2_3982 ( .A(u5__abc_81276_new_n375_), .B(u5__abc_81276_new_n378_), .Y(u5__abc_81276_new_n379_));
AND2X2 AND2X2_3983 ( .A(u5__abc_81276_new_n382_), .B(u5__abc_81276_new_n380_), .Y(u5__abc_81276_new_n383_));
AND2X2 AND2X2_3984 ( .A(u5__abc_81276_new_n383_), .B(u5__abc_81276_new_n379_), .Y(u5__abc_81276_new_n384_));
AND2X2 AND2X2_3985 ( .A(u5__abc_81276_new_n384_), .B(u5__abc_81276_new_n372_), .Y(u5__abc_81276_new_n385_));
AND2X2 AND2X2_3986 ( .A(u5__abc_81276_new_n387_), .B(u5__abc_81276_new_n388_), .Y(u5__abc_81276_new_n389_));
AND2X2 AND2X2_3987 ( .A(u5__abc_81276_new_n390_), .B(u5__abc_81276_new_n391_), .Y(u5__abc_81276_new_n392_));
AND2X2 AND2X2_3988 ( .A(u5__abc_81276_new_n389_), .B(u5__abc_81276_new_n392_), .Y(u5__abc_81276_new_n393_));
AND2X2 AND2X2_3989 ( .A(u5__abc_81276_new_n394_), .B(u5__abc_81276_new_n395_), .Y(u5__abc_81276_new_n396_));
AND2X2 AND2X2_399 ( .A(u0__abc_76628_new_n1691_), .B(u0__abc_76628_new_n1174__bF_buf2), .Y(u0__abc_76628_new_n1692_));
AND2X2 AND2X2_3990 ( .A(u5__abc_81276_new_n397_), .B(u5__abc_81276_new_n398_), .Y(u5__abc_81276_new_n399_));
AND2X2 AND2X2_3991 ( .A(u5__abc_81276_new_n396_), .B(u5__abc_81276_new_n399_), .Y(u5__abc_81276_new_n400_));
AND2X2 AND2X2_3992 ( .A(u5__abc_81276_new_n393_), .B(u5__abc_81276_new_n400_), .Y(u5__abc_81276_new_n401_));
AND2X2 AND2X2_3993 ( .A(u5__abc_81276_new_n402_), .B(u5__abc_81276_new_n403_), .Y(u5__abc_81276_new_n404_));
AND2X2 AND2X2_3994 ( .A(u5__abc_81276_new_n405_), .B(u5__abc_81276_new_n406_), .Y(u5__abc_81276_new_n407_));
AND2X2 AND2X2_3995 ( .A(u5__abc_81276_new_n404_), .B(u5__abc_81276_new_n407_), .Y(u5__abc_81276_new_n408_));
AND2X2 AND2X2_3996 ( .A(u5__abc_81276_new_n409_), .B(u5__abc_81276_new_n410_), .Y(u5__abc_81276_new_n411_));
AND2X2 AND2X2_3997 ( .A(u5__abc_81276_new_n412_), .B(u5__abc_81276_new_n413_), .Y(u5__abc_81276_new_n414_));
AND2X2 AND2X2_3998 ( .A(u5__abc_81276_new_n411_), .B(u5__abc_81276_new_n414_), .Y(u5__abc_81276_new_n415_));
AND2X2 AND2X2_3999 ( .A(u5__abc_81276_new_n408_), .B(u5__abc_81276_new_n415_), .Y(u5__abc_81276_new_n416_));
AND2X2 AND2X2_4 ( .A(_abc_85006_new_n248_), .B(_abc_85006_new_n249_), .Y(_abc_85006_new_n250_));
AND2X2 AND2X2_40 ( .A(_abc_85006_new_n356_), .B(_abc_85006_new_n357_), .Y(tms_s_22_));
AND2X2 AND2X2_400 ( .A(spec_req_cs_3_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1693_));
AND2X2 AND2X2_4000 ( .A(u5__abc_81276_new_n401__bF_buf3), .B(u5__abc_81276_new_n416__bF_buf3), .Y(u5__abc_81276_new_n417_));
AND2X2 AND2X2_4001 ( .A(u5__abc_81276_new_n418_), .B(u5__abc_81276_new_n419_), .Y(u5__abc_81276_new_n420_));
AND2X2 AND2X2_4002 ( .A(u5__abc_81276_new_n421_), .B(u5__abc_81276_new_n422_), .Y(u5__abc_81276_new_n423_));
AND2X2 AND2X2_4003 ( .A(u5__abc_81276_new_n420_), .B(u5__abc_81276_new_n423_), .Y(u5__abc_81276_new_n424_));
AND2X2 AND2X2_4004 ( .A(u5__abc_81276_new_n425_), .B(u5__abc_81276_new_n426_), .Y(u5__abc_81276_new_n427_));
AND2X2 AND2X2_4005 ( .A(u5__abc_81276_new_n428_), .B(u5__abc_81276_new_n429_), .Y(u5__abc_81276_new_n430_));
AND2X2 AND2X2_4006 ( .A(u5__abc_81276_new_n427_), .B(u5__abc_81276_new_n430_), .Y(u5__abc_81276_new_n431_));
AND2X2 AND2X2_4007 ( .A(u5__abc_81276_new_n424_), .B(u5__abc_81276_new_n431_), .Y(u5__abc_81276_new_n432_));
AND2X2 AND2X2_4008 ( .A(u5__abc_81276_new_n433_), .B(u5__abc_81276_new_n434_), .Y(u5__abc_81276_new_n435_));
AND2X2 AND2X2_4009 ( .A(u5__abc_81276_new_n436_), .B(u5__abc_81276_new_n437_), .Y(u5__abc_81276_new_n438_));
AND2X2 AND2X2_401 ( .A(u0__abc_76628_new_n1694_), .B(u0__abc_76628_new_n1173__bF_buf2), .Y(u0__abc_76628_new_n1695_));
AND2X2 AND2X2_4010 ( .A(u5__abc_81276_new_n435_), .B(u5__abc_81276_new_n438_), .Y(u5__abc_81276_new_n439_));
AND2X2 AND2X2_4011 ( .A(u5__abc_81276_new_n440_), .B(u5__abc_81276_new_n441_), .Y(u5__abc_81276_new_n442_));
AND2X2 AND2X2_4012 ( .A(u5__abc_81276_new_n443_), .B(u5__abc_81276_new_n444_), .Y(u5__abc_81276_new_n445_));
AND2X2 AND2X2_4013 ( .A(u5__abc_81276_new_n442_), .B(u5__abc_81276_new_n445_), .Y(u5__abc_81276_new_n446_));
AND2X2 AND2X2_4014 ( .A(u5__abc_81276_new_n439_), .B(u5__abc_81276_new_n446_), .Y(u5__abc_81276_new_n447_));
AND2X2 AND2X2_4015 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n447_), .Y(u5__abc_81276_new_n448_));
AND2X2 AND2X2_4016 ( .A(u5__abc_81276_new_n417__bF_buf3), .B(u5__abc_81276_new_n448__bF_buf5), .Y(u5__abc_81276_new_n449_));
AND2X2 AND2X2_4017 ( .A(u5__abc_81276_new_n450_), .B(u5__abc_81276_new_n451_), .Y(u5__abc_81276_new_n452_));
AND2X2 AND2X2_4018 ( .A(u5__abc_81276_new_n453_), .B(u5__abc_81276_new_n454_), .Y(u5__abc_81276_new_n455_));
AND2X2 AND2X2_4019 ( .A(u5__abc_81276_new_n452_), .B(u5__abc_81276_new_n455_), .Y(u5__abc_81276_new_n456_));
AND2X2 AND2X2_402 ( .A(spec_req_cs_2_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1696_));
AND2X2 AND2X2_4020 ( .A(u5__abc_81276_new_n457_), .B(u5__abc_81276_new_n458_), .Y(u5__abc_81276_new_n459_));
AND2X2 AND2X2_4021 ( .A(u5__abc_81276_new_n460_), .B(u5__abc_81276_new_n461_), .Y(u5__abc_81276_new_n462_));
AND2X2 AND2X2_4022 ( .A(u5__abc_81276_new_n459_), .B(u5__abc_81276_new_n462_), .Y(u5__abc_81276_new_n463_));
AND2X2 AND2X2_4023 ( .A(u5__abc_81276_new_n456_), .B(u5__abc_81276_new_n463_), .Y(u5__abc_81276_new_n464_));
AND2X2 AND2X2_4024 ( .A(u5__abc_81276_new_n465_), .B(u5__abc_81276_new_n466_), .Y(u5__abc_81276_new_n467_));
AND2X2 AND2X2_4025 ( .A(u5__abc_81276_new_n468_), .B(u5__abc_81276_new_n469_), .Y(u5__abc_81276_new_n470_));
AND2X2 AND2X2_4026 ( .A(u5__abc_81276_new_n467_), .B(u5__abc_81276_new_n470_), .Y(u5__abc_81276_new_n471_));
AND2X2 AND2X2_4027 ( .A(u5__abc_81276_new_n472_), .B(u5__abc_81276_new_n473_), .Y(u5__abc_81276_new_n474_));
AND2X2 AND2X2_4028 ( .A(u5__abc_81276_new_n475_), .B(u5__abc_81276_new_n476_), .Y(u5__abc_81276_new_n477_));
AND2X2 AND2X2_4029 ( .A(u5__abc_81276_new_n474_), .B(u5__abc_81276_new_n477_), .Y(u5__abc_81276_new_n478_));
AND2X2 AND2X2_403 ( .A(u0__abc_76628_new_n1697_), .B(u0__abc_76628_new_n1172__bF_buf2), .Y(u0__abc_76628_new_n1698_));
AND2X2 AND2X2_4030 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n478_), .Y(u5__abc_81276_new_n479_));
AND2X2 AND2X2_4031 ( .A(u5__abc_81276_new_n464__bF_buf3), .B(u5__abc_81276_new_n479__bF_buf3), .Y(u5__abc_81276_new_n480_));
AND2X2 AND2X2_4032 ( .A(u5__abc_81276_new_n481_), .B(u5__abc_81276_new_n482_), .Y(u5__abc_81276_new_n483_));
AND2X2 AND2X2_4033 ( .A(u5__abc_81276_new_n484_), .B(u5__abc_81276_new_n485_), .Y(u5__abc_81276_new_n486_));
AND2X2 AND2X2_4034 ( .A(u5__abc_81276_new_n483_), .B(u5__abc_81276_new_n486_), .Y(u5__abc_81276_new_n487_));
AND2X2 AND2X2_4035 ( .A(u5__abc_81276_new_n488_), .B(u5__abc_81276_new_n489_), .Y(u5__abc_81276_new_n490_));
AND2X2 AND2X2_4036 ( .A(u5__abc_81276_new_n491_), .B(u5__abc_81276_new_n492_), .Y(u5__abc_81276_new_n493_));
AND2X2 AND2X2_4037 ( .A(u5__abc_81276_new_n494_), .B(u5__abc_81276_new_n495_), .Y(u5__abc_81276_new_n496_));
AND2X2 AND2X2_4038 ( .A(u5__abc_81276_new_n493_), .B(u5__abc_81276_new_n496_), .Y(u5__abc_81276_new_n497_));
AND2X2 AND2X2_4039 ( .A(u5__abc_81276_new_n497_), .B(u5__abc_81276_new_n490__bF_buf10), .Y(u5__abc_81276_new_n498_));
AND2X2 AND2X2_404 ( .A(spec_req_cs_1_bF_buf5_), .B(u0_tms1_21_), .Y(u0__abc_76628_new_n1699_));
AND2X2 AND2X2_4040 ( .A(u5__abc_81276_new_n498_), .B(u5__abc_81276_new_n487_), .Y(u5__abc_81276_new_n499_));
AND2X2 AND2X2_4041 ( .A(u5__abc_81276_new_n480__bF_buf4), .B(u5__abc_81276_new_n499_), .Y(u5__abc_81276_new_n500_));
AND2X2 AND2X2_4042 ( .A(u5__abc_81276_new_n449__bF_buf7), .B(u5__abc_81276_new_n500_), .Y(u5__abc_81276_new_n501_));
AND2X2 AND2X2_4043 ( .A(u5__abc_81276_new_n502_), .B(u5__abc_81276_new_n503_), .Y(u5__abc_81276_new_n504_));
AND2X2 AND2X2_4044 ( .A(u5__abc_81276_new_n505_), .B(u5__abc_81276_new_n506_), .Y(u5__abc_81276_new_n507_));
AND2X2 AND2X2_4045 ( .A(u5__abc_81276_new_n504_), .B(u5__abc_81276_new_n507_), .Y(u5__abc_81276_new_n508_));
AND2X2 AND2X2_4046 ( .A(u5__abc_81276_new_n509_), .B(u5__abc_81276_new_n510_), .Y(u5__abc_81276_new_n511_));
AND2X2 AND2X2_4047 ( .A(u5__abc_81276_new_n512_), .B(u5_state_30_), .Y(u5__abc_81276_new_n513_));
AND2X2 AND2X2_4048 ( .A(u5__abc_81276_new_n511_), .B(u5__abc_81276_new_n513_), .Y(u5__abc_81276_new_n514_));
AND2X2 AND2X2_4049 ( .A(u5__abc_81276_new_n508_), .B(u5__abc_81276_new_n514_), .Y(u5__abc_81276_new_n515_));
AND2X2 AND2X2_405 ( .A(u0__abc_76628_new_n1169__bF_buf5), .B(u0__abc_76628_new_n1702_), .Y(u0__abc_76628_new_n1703_));
AND2X2 AND2X2_4050 ( .A(u5__abc_81276_new_n501_), .B(u5__abc_81276_new_n515_), .Y(u5__abc_81276_new_n516_));
AND2X2 AND2X2_4051 ( .A(u5__abc_81276_new_n487_), .B(u5__abc_81276_new_n497_), .Y(u5__abc_81276_new_n517_));
AND2X2 AND2X2_4052 ( .A(u5__abc_81276_new_n518_), .B(u5__abc_81276_new_n512_), .Y(u5__abc_81276_new_n519_));
AND2X2 AND2X2_4053 ( .A(u5__abc_81276_new_n511_), .B(u5__abc_81276_new_n519_), .Y(u5__abc_81276_new_n520_));
AND2X2 AND2X2_4054 ( .A(u5__abc_81276_new_n508_), .B(u5__abc_81276_new_n520_), .Y(u5__abc_81276_new_n521_));
AND2X2 AND2X2_4055 ( .A(u5__abc_81276_new_n517_), .B(u5__abc_81276_new_n521__bF_buf3), .Y(u5__abc_81276_new_n522_));
AND2X2 AND2X2_4056 ( .A(u5__abc_81276_new_n480__bF_buf3), .B(u5__abc_81276_new_n522__bF_buf4), .Y(u5__abc_81276_new_n523_));
AND2X2 AND2X2_4057 ( .A(u5__abc_81276_new_n444_), .B(u5_state_32_), .Y(u5__abc_81276_new_n524_));
AND2X2 AND2X2_4058 ( .A(u5__abc_81276_new_n490__bF_buf9), .B(u5__abc_81276_new_n524_), .Y(u5__abc_81276_new_n525_));
AND2X2 AND2X2_4059 ( .A(u5__abc_81276_new_n525_), .B(u5__abc_81276_new_n442_), .Y(u5__abc_81276_new_n526_));
AND2X2 AND2X2_406 ( .A(u0__abc_76628_new_n1701_), .B(u0__abc_76628_new_n1703_), .Y(u0__abc_76628_new_n1704_));
AND2X2 AND2X2_4060 ( .A(u5__abc_81276_new_n526_), .B(u5__abc_81276_new_n439_), .Y(u5__abc_81276_new_n527_));
AND2X2 AND2X2_4061 ( .A(u5__abc_81276_new_n527_), .B(u5__abc_81276_new_n432_), .Y(u5__abc_81276_new_n528_));
AND2X2 AND2X2_4062 ( .A(u5__abc_81276_new_n528_), .B(u5__abc_81276_new_n417__bF_buf2), .Y(u5__abc_81276_new_n529_));
AND2X2 AND2X2_4063 ( .A(u5__abc_81276_new_n529_), .B(u5__abc_81276_new_n523__bF_buf7), .Y(u5__abc_81276_new_n530_));
AND2X2 AND2X2_4064 ( .A(u5__abc_81276_new_n480__bF_buf2), .B(u5__abc_81276_new_n498_), .Y(u5__abc_81276_new_n531_));
AND2X2 AND2X2_4065 ( .A(u5__abc_81276_new_n449__bF_buf6), .B(u5__abc_81276_new_n531_), .Y(u5__abc_81276_new_n532_));
AND2X2 AND2X2_4066 ( .A(u5__abc_81276_new_n518_), .B(u5_state_31_), .Y(u5__abc_81276_new_n533_));
AND2X2 AND2X2_4067 ( .A(u5__abc_81276_new_n511_), .B(u5__abc_81276_new_n533_), .Y(u5__abc_81276_new_n534_));
AND2X2 AND2X2_4068 ( .A(u5__abc_81276_new_n487_), .B(u5__abc_81276_new_n534_), .Y(u5__abc_81276_new_n535_));
AND2X2 AND2X2_4069 ( .A(u5__abc_81276_new_n535_), .B(u5__abc_81276_new_n508_), .Y(u5__abc_81276_new_n536_));
AND2X2 AND2X2_407 ( .A(u0__abc_76628_new_n1170__bF_buf5), .B(sp_tms_22_), .Y(u0__abc_76628_new_n1706_));
AND2X2 AND2X2_4070 ( .A(u5__abc_81276_new_n532_), .B(u5__abc_81276_new_n536_), .Y(u5__abc_81276_new_n537_));
AND2X2 AND2X2_4071 ( .A(u5__abc_81276_new_n506_), .B(u5_state_25_), .Y(u5__abc_81276_new_n540_));
AND2X2 AND2X2_4072 ( .A(u5__abc_81276_new_n490__bF_buf8), .B(u5__abc_81276_new_n540_), .Y(u5__abc_81276_new_n541_));
AND2X2 AND2X2_4073 ( .A(u5__abc_81276_new_n541_), .B(u5__abc_81276_new_n504_), .Y(u5__abc_81276_new_n542_));
AND2X2 AND2X2_4074 ( .A(u5__abc_81276_new_n517_), .B(u5__abc_81276_new_n542_), .Y(u5__abc_81276_new_n543_));
AND2X2 AND2X2_4075 ( .A(u5__abc_81276_new_n480__bF_buf1), .B(u5__abc_81276_new_n543_), .Y(u5__abc_81276_new_n544_));
AND2X2 AND2X2_4076 ( .A(u5__abc_81276_new_n449__bF_buf5), .B(u5__abc_81276_new_n544_), .Y(u5__abc_81276_new_n545_));
AND2X2 AND2X2_4077 ( .A(u5__abc_81276_new_n545_), .B(u5__abc_81276_new_n520_), .Y(u5__abc_81276_new_n546_));
AND2X2 AND2X2_4078 ( .A(u5__abc_81276_new_n502_), .B(u5_state_26_), .Y(u5__abc_81276_new_n548_));
AND2X2 AND2X2_4079 ( .A(u5__abc_81276_new_n490__bF_buf7), .B(u5__abc_81276_new_n548_), .Y(u5__abc_81276_new_n549_));
AND2X2 AND2X2_408 ( .A(spec_req_cs_5_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1707_));
AND2X2 AND2X2_4080 ( .A(u5__abc_81276_new_n549_), .B(u5__abc_81276_new_n507_), .Y(u5__abc_81276_new_n550_));
AND2X2 AND2X2_4081 ( .A(u5__abc_81276_new_n517_), .B(u5__abc_81276_new_n550_), .Y(u5__abc_81276_new_n551_));
AND2X2 AND2X2_4082 ( .A(u5__abc_81276_new_n480__bF_buf0), .B(u5__abc_81276_new_n551_), .Y(u5__abc_81276_new_n552_));
AND2X2 AND2X2_4083 ( .A(u5__abc_81276_new_n449__bF_buf4), .B(u5__abc_81276_new_n552_), .Y(u5__abc_81276_new_n553_));
AND2X2 AND2X2_4084 ( .A(u5__abc_81276_new_n553_), .B(u5__abc_81276_new_n520_), .Y(u5__abc_81276_new_n554_));
AND2X2 AND2X2_4085 ( .A(u5__abc_81276_new_n547_), .B(u5__abc_81276_new_n555_), .Y(u5__abc_81276_new_n556_));
AND2X2 AND2X2_4086 ( .A(u5__abc_81276_new_n417__bF_buf1), .B(u5__abc_81276_new_n432_), .Y(u5__abc_81276_new_n557_));
AND2X2 AND2X2_4087 ( .A(u5__abc_81276_new_n490__bF_buf6), .B(u5_state_35_), .Y(u5__abc_81276_new_n558_));
AND2X2 AND2X2_4088 ( .A(u5__abc_81276_new_n445_), .B(u5__abc_81276_new_n441_), .Y(u5__abc_81276_new_n559_));
AND2X2 AND2X2_4089 ( .A(u5__abc_81276_new_n439_), .B(u5__abc_81276_new_n559_), .Y(u5__abc_81276_new_n560_));
AND2X2 AND2X2_409 ( .A(u0__abc_76628_new_n1709_), .B(u0__abc_76628_new_n1179__bF_buf1), .Y(u0__abc_76628_new_n1710_));
AND2X2 AND2X2_4090 ( .A(u5__abc_81276_new_n560_), .B(u5__abc_81276_new_n558_), .Y(u5__abc_81276_new_n561_));
AND2X2 AND2X2_4091 ( .A(u5__abc_81276_new_n557_), .B(u5__abc_81276_new_n561_), .Y(u5__abc_81276_new_n562_));
AND2X2 AND2X2_4092 ( .A(u5__abc_81276_new_n562_), .B(u5__abc_81276_new_n523__bF_buf6), .Y(u5__abc_81276_new_n563_));
AND2X2 AND2X2_4093 ( .A(u5__abc_81276_new_n511_), .B(u5__abc_81276_new_n512_), .Y(u5__abc_81276_new_n565_));
AND2X2 AND2X2_4094 ( .A(u5__abc_81276_new_n490__bF_buf5), .B(u5_state_30_), .Y(u5__abc_81276_new_n566_));
AND2X2 AND2X2_4095 ( .A(u5__abc_81276_new_n565_), .B(u5__abc_81276_new_n566_), .Y(u5__abc_81276_new_n567_));
AND2X2 AND2X2_4096 ( .A(u5__abc_81276_new_n567_), .B(u5__abc_81276_new_n508_), .Y(u5__abc_81276_new_n568_));
AND2X2 AND2X2_4097 ( .A(u5__abc_81276_new_n480__bF_buf4), .B(u5__abc_81276_new_n568_), .Y(u5__abc_81276_new_n569_));
AND2X2 AND2X2_4098 ( .A(u5__abc_81276_new_n449__bF_buf3), .B(u5__abc_81276_new_n569_), .Y(u5__abc_81276_new_n570_));
AND2X2 AND2X2_4099 ( .A(u5__abc_81276_new_n570_), .B(u5__abc_81276_new_n517_), .Y(u5__abc_81276_new_n571_));
AND2X2 AND2X2_41 ( .A(_abc_85006_new_n359_), .B(_abc_85006_new_n360_), .Y(tms_s_23_));
AND2X2 AND2X2_410 ( .A(u0__abc_76628_new_n1710_), .B(u0__abc_76628_new_n1708_), .Y(u0__abc_76628_new_n1711_));
AND2X2 AND2X2_4100 ( .A(u5__abc_81276_new_n490__bF_buf4), .B(u5_state_32_), .Y(u5__abc_81276_new_n573_));
AND2X2 AND2X2_4101 ( .A(u5__abc_81276_new_n442_), .B(u5__abc_81276_new_n444_), .Y(u5__abc_81276_new_n574_));
AND2X2 AND2X2_4102 ( .A(u5__abc_81276_new_n439_), .B(u5__abc_81276_new_n574_), .Y(u5__abc_81276_new_n575_));
AND2X2 AND2X2_4103 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n575_), .Y(u5__abc_81276_new_n576_));
AND2X2 AND2X2_4104 ( .A(u5__abc_81276_new_n576_), .B(u5__abc_81276_new_n573_), .Y(u5__abc_81276_new_n577_));
AND2X2 AND2X2_4105 ( .A(u5__abc_81276_new_n577_), .B(u5__abc_81276_new_n417__bF_buf0), .Y(u5__abc_81276_new_n578_));
AND2X2 AND2X2_4106 ( .A(u5__abc_81276_new_n578_), .B(u5__abc_81276_new_n523__bF_buf5), .Y(u5__abc_81276_new_n579_));
AND2X2 AND2X2_4107 ( .A(u5__abc_81276_new_n572_), .B(u5__abc_81276_new_n580_), .Y(u5__abc_81276_new_n581_));
AND2X2 AND2X2_4108 ( .A(u5__abc_81276_new_n519_), .B(u5__abc_81276_new_n509_), .Y(u5__abc_81276_new_n582_));
AND2X2 AND2X2_4109 ( .A(u5__abc_81276_new_n508_), .B(u5__abc_81276_new_n582_), .Y(u5__abc_81276_new_n583_));
AND2X2 AND2X2_411 ( .A(u0__abc_76628_new_n1712_), .B(u0__abc_76628_new_n1175__bF_buf1), .Y(u0__abc_76628_new_n1713_));
AND2X2 AND2X2_4110 ( .A(u5__abc_81276_new_n499_), .B(u5__abc_81276_new_n583_), .Y(u5__abc_81276_new_n584_));
AND2X2 AND2X2_4111 ( .A(u5__abc_81276_new_n584_), .B(u5__abc_81276_new_n480__bF_buf3), .Y(u5__abc_81276_new_n585_));
AND2X2 AND2X2_4112 ( .A(u5__abc_81276_new_n449__bF_buf2), .B(u5_state_28_), .Y(u5__abc_81276_new_n586_));
AND2X2 AND2X2_4113 ( .A(u5__abc_81276_new_n586_), .B(u5__abc_81276_new_n585_), .Y(u5__abc_81276_new_n587_));
AND2X2 AND2X2_4114 ( .A(u5__abc_81276_new_n581_), .B(u5__abc_81276_new_n588_), .Y(u5__abc_81276_new_n589_));
AND2X2 AND2X2_4115 ( .A(u5__abc_81276_new_n510_), .B(u5_state_29_), .Y(u5__abc_81276_new_n590_));
AND2X2 AND2X2_4116 ( .A(u5__abc_81276_new_n508_), .B(u5__abc_81276_new_n519_), .Y(u5__abc_81276_new_n591_));
AND2X2 AND2X2_4117 ( .A(u5__abc_81276_new_n591_), .B(u5__abc_81276_new_n590_), .Y(u5__abc_81276_new_n592_));
AND2X2 AND2X2_4118 ( .A(u5__abc_81276_new_n499_), .B(u5__abc_81276_new_n592_), .Y(u5__abc_81276_new_n593_));
AND2X2 AND2X2_4119 ( .A(u5__abc_81276_new_n593_), .B(u5__abc_81276_new_n480__bF_buf2), .Y(u5__abc_81276_new_n594_));
AND2X2 AND2X2_412 ( .A(spec_req_cs_4_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1714_));
AND2X2 AND2X2_4120 ( .A(u5__abc_81276_new_n594_), .B(u5__abc_81276_new_n449__bF_buf1), .Y(u5__abc_81276_new_n595_));
AND2X2 AND2X2_4121 ( .A(u5__abc_81276_new_n507_), .B(u5__abc_81276_new_n503_), .Y(u5__abc_81276_new_n597_));
AND2X2 AND2X2_4122 ( .A(u5__abc_81276_new_n520_), .B(u5__abc_81276_new_n597_), .Y(u5__abc_81276_new_n598_));
AND2X2 AND2X2_4123 ( .A(u5__abc_81276_new_n499_), .B(u5__abc_81276_new_n598_), .Y(u5__abc_81276_new_n599_));
AND2X2 AND2X2_4124 ( .A(u5__abc_81276_new_n599_), .B(u5__abc_81276_new_n480__bF_buf1), .Y(u5__abc_81276_new_n600_));
AND2X2 AND2X2_4125 ( .A(u5__abc_81276_new_n449__bF_buf0), .B(u5_state_27_), .Y(u5__abc_81276_new_n601_));
AND2X2 AND2X2_4126 ( .A(u5__abc_81276_new_n601_), .B(u5__abc_81276_new_n600_), .Y(u5__abc_81276_new_n602_));
AND2X2 AND2X2_4127 ( .A(u5__abc_81276_new_n603_), .B(u5__abc_81276_new_n596_), .Y(u5__abc_81276_new_n604_));
AND2X2 AND2X2_4128 ( .A(u5__abc_81276_new_n589_), .B(u5__abc_81276_new_n604_), .Y(u5__abc_81276_new_n605_));
AND2X2 AND2X2_4129 ( .A(u5__abc_81276_new_n605_), .B(u5__abc_81276_new_n564_), .Y(u5__abc_81276_new_n606_));
AND2X2 AND2X2_413 ( .A(u0__abc_76628_new_n1715_), .B(u0__abc_76628_new_n1174__bF_buf1), .Y(u0__abc_76628_new_n1716_));
AND2X2 AND2X2_4130 ( .A(u5__abc_81276_new_n606_), .B(u5__abc_81276_new_n556_), .Y(u5__abc_81276_new_n607_));
AND2X2 AND2X2_4131 ( .A(u5__abc_81276_new_n482_), .B(u5_state_19_), .Y(u5__abc_81276_new_n608_));
AND2X2 AND2X2_4132 ( .A(u5__abc_81276_new_n486_), .B(u5__abc_81276_new_n608_), .Y(u5__abc_81276_new_n609_));
AND2X2 AND2X2_4133 ( .A(u5__abc_81276_new_n521__bF_buf2), .B(u5__abc_81276_new_n609_), .Y(u5__abc_81276_new_n610_));
AND2X2 AND2X2_4134 ( .A(u5__abc_81276_new_n532_), .B(u5__abc_81276_new_n610_), .Y(u5__abc_81276_new_n611_));
AND2X2 AND2X2_4135 ( .A(u5__abc_81276_new_n485_), .B(u5_state_17_), .Y(u5__abc_81276_new_n613_));
AND2X2 AND2X2_4136 ( .A(u5__abc_81276_new_n483_), .B(u5__abc_81276_new_n613_), .Y(u5__abc_81276_new_n614_));
AND2X2 AND2X2_4137 ( .A(u5__abc_81276_new_n498_), .B(u5__abc_81276_new_n614_), .Y(u5__abc_81276_new_n615_));
AND2X2 AND2X2_4138 ( .A(u5__abc_81276_new_n480__bF_buf0), .B(u5__abc_81276_new_n615_), .Y(u5__abc_81276_new_n616_));
AND2X2 AND2X2_4139 ( .A(u5__abc_81276_new_n449__bF_buf7), .B(u5__abc_81276_new_n616_), .Y(u5__abc_81276_new_n617_));
AND2X2 AND2X2_414 ( .A(spec_req_cs_3_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1717_));
AND2X2 AND2X2_4140 ( .A(u5__abc_81276_new_n617_), .B(u5__abc_81276_new_n521__bF_buf1), .Y(u5__abc_81276_new_n618_));
AND2X2 AND2X2_4141 ( .A(u5__abc_81276_new_n612_), .B(u5__abc_81276_new_n619_), .Y(u5__abc_81276_new_n620_));
AND2X2 AND2X2_4142 ( .A(u5__abc_81276_new_n484_), .B(u5_state_16_), .Y(u5__abc_81276_new_n621_));
AND2X2 AND2X2_4143 ( .A(u5__abc_81276_new_n483_), .B(u5__abc_81276_new_n621_), .Y(u5__abc_81276_new_n622_));
AND2X2 AND2X2_4144 ( .A(u5__abc_81276_new_n521__bF_buf0), .B(u5__abc_81276_new_n622_), .Y(u5__abc_81276_new_n623_));
AND2X2 AND2X2_4145 ( .A(u5__abc_81276_new_n532_), .B(u5__abc_81276_new_n623_), .Y(u5__abc_81276_new_n624_));
AND2X2 AND2X2_4146 ( .A(u5__abc_81276_new_n481_), .B(u5_state_18_), .Y(u5__abc_81276_new_n626_));
AND2X2 AND2X2_4147 ( .A(u5__abc_81276_new_n486_), .B(u5__abc_81276_new_n626_), .Y(u5__abc_81276_new_n627_));
AND2X2 AND2X2_4148 ( .A(u5__abc_81276_new_n521__bF_buf3), .B(u5__abc_81276_new_n627_), .Y(u5__abc_81276_new_n628_));
AND2X2 AND2X2_4149 ( .A(u5__abc_81276_new_n532_), .B(u5__abc_81276_new_n628_), .Y(u5__abc_81276_new_n629_));
AND2X2 AND2X2_415 ( .A(u0__abc_76628_new_n1718_), .B(u0__abc_76628_new_n1173__bF_buf1), .Y(u0__abc_76628_new_n1719_));
AND2X2 AND2X2_4150 ( .A(u5__abc_81276_new_n625_), .B(u5__abc_81276_new_n630_), .Y(u5__abc_81276_new_n631_));
AND2X2 AND2X2_4151 ( .A(u5__abc_81276_new_n505_), .B(u5_state_24_), .Y(u5__abc_81276_new_n632_));
AND2X2 AND2X2_4152 ( .A(u5__abc_81276_new_n490__bF_buf3), .B(u5__abc_81276_new_n632_), .Y(u5__abc_81276_new_n633_));
AND2X2 AND2X2_4153 ( .A(u5__abc_81276_new_n633_), .B(u5__abc_81276_new_n504_), .Y(u5__abc_81276_new_n634_));
AND2X2 AND2X2_4154 ( .A(u5__abc_81276_new_n517_), .B(u5__abc_81276_new_n634_), .Y(u5__abc_81276_new_n635_));
AND2X2 AND2X2_4155 ( .A(u5__abc_81276_new_n480__bF_buf4), .B(u5__abc_81276_new_n635_), .Y(u5__abc_81276_new_n636_));
AND2X2 AND2X2_4156 ( .A(u5__abc_81276_new_n449__bF_buf6), .B(u5__abc_81276_new_n636_), .Y(u5__abc_81276_new_n637_));
AND2X2 AND2X2_4157 ( .A(u5__abc_81276_new_n637_), .B(u5__abc_81276_new_n520_), .Y(u5__abc_81276_new_n638_));
AND2X2 AND2X2_4158 ( .A(u5__abc_81276_new_n493_), .B(u5__abc_81276_new_n490__bF_buf2), .Y(u5__abc_81276_new_n640_));
AND2X2 AND2X2_4159 ( .A(u5__abc_81276_new_n495_), .B(u5_state_23_), .Y(u5__abc_81276_new_n641_));
AND2X2 AND2X2_416 ( .A(spec_req_cs_2_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1720_));
AND2X2 AND2X2_4160 ( .A(u5__abc_81276_new_n487_), .B(u5__abc_81276_new_n641_), .Y(u5__abc_81276_new_n642_));
AND2X2 AND2X2_4161 ( .A(u5__abc_81276_new_n642_), .B(u5__abc_81276_new_n640_), .Y(u5__abc_81276_new_n643_));
AND2X2 AND2X2_4162 ( .A(u5__abc_81276_new_n480__bF_buf3), .B(u5__abc_81276_new_n643_), .Y(u5__abc_81276_new_n644_));
AND2X2 AND2X2_4163 ( .A(u5__abc_81276_new_n449__bF_buf5), .B(u5__abc_81276_new_n644_), .Y(u5__abc_81276_new_n645_));
AND2X2 AND2X2_4164 ( .A(u5__abc_81276_new_n645_), .B(u5__abc_81276_new_n521__bF_buf2), .Y(u5__abc_81276_new_n646_));
AND2X2 AND2X2_4165 ( .A(u5__abc_81276_new_n639_), .B(u5__abc_81276_new_n647_), .Y(u5__abc_81276_new_n648_));
AND2X2 AND2X2_4166 ( .A(u5__abc_81276_new_n494_), .B(u5_state_22_), .Y(u5__abc_81276_new_n649_));
AND2X2 AND2X2_4167 ( .A(u5__abc_81276_new_n487_), .B(u5__abc_81276_new_n649_), .Y(u5__abc_81276_new_n650_));
AND2X2 AND2X2_4168 ( .A(u5__abc_81276_new_n650_), .B(u5__abc_81276_new_n640_), .Y(u5__abc_81276_new_n651_));
AND2X2 AND2X2_4169 ( .A(u5__abc_81276_new_n480__bF_buf2), .B(u5__abc_81276_new_n651_), .Y(u5__abc_81276_new_n652_));
AND2X2 AND2X2_417 ( .A(u0__abc_76628_new_n1721_), .B(u0__abc_76628_new_n1172__bF_buf1), .Y(u0__abc_76628_new_n1722_));
AND2X2 AND2X2_4170 ( .A(u5__abc_81276_new_n449__bF_buf4), .B(u5__abc_81276_new_n652_), .Y(u5__abc_81276_new_n653_));
AND2X2 AND2X2_4171 ( .A(u5__abc_81276_new_n653_), .B(u5__abc_81276_new_n521__bF_buf1), .Y(u5__abc_81276_new_n654_));
AND2X2 AND2X2_4172 ( .A(u5__abc_81276_new_n492_), .B(u5_state_20_), .Y(u5__abc_81276_new_n660_));
AND2X2 AND2X2_4173 ( .A(u5__abc_81276_new_n487_), .B(u5__abc_81276_new_n660_), .Y(u5__abc_81276_new_n661_));
AND2X2 AND2X2_4174 ( .A(u5__abc_81276_new_n659_), .B(u5__abc_81276_new_n661_), .Y(u5__abc_81276_new_n662_));
AND2X2 AND2X2_4175 ( .A(u5__abc_81276_new_n662_), .B(u5__abc_81276_new_n480__bF_buf1), .Y(u5__abc_81276_new_n663_));
AND2X2 AND2X2_4176 ( .A(u5__abc_81276_new_n663_), .B(u5__abc_81276_new_n449__bF_buf3), .Y(u5__abc_81276_new_n664_));
AND2X2 AND2X2_4177 ( .A(u5__abc_81276_new_n664_), .B(u5__abc_81276_new_n521__bF_buf0), .Y(u5__abc_81276_new_n665_));
AND2X2 AND2X2_4178 ( .A(u5__abc_81276_new_n666_), .B(u5__abc_81276_new_n655_), .Y(u5__abc_81276_new_n667_));
AND2X2 AND2X2_4179 ( .A(u5__abc_81276_new_n667_), .B(u5__abc_81276_new_n648_), .Y(u5__abc_81276_new_n668_));
AND2X2 AND2X2_418 ( .A(spec_req_cs_1_bF_buf4_), .B(u0_tms1_22_), .Y(u0__abc_76628_new_n1723_));
AND2X2 AND2X2_4180 ( .A(u5__abc_81276_new_n668_), .B(u5__abc_81276_new_n631_), .Y(u5__abc_81276_new_n669_));
AND2X2 AND2X2_4181 ( .A(u5__abc_81276_new_n669_), .B(u5__abc_81276_new_n620_), .Y(u5__abc_81276_new_n670_));
AND2X2 AND2X2_4182 ( .A(u5__abc_81276_new_n607_), .B(u5__abc_81276_new_n670_), .Y(u5__abc_81276_new_n671_));
AND2X2 AND2X2_4183 ( .A(u5__abc_81276_new_n410_), .B(u5_state_51_), .Y(u5__abc_81276_new_n672_));
AND2X2 AND2X2_4184 ( .A(u5__abc_81276_new_n490__bF_buf0), .B(u5__abc_81276_new_n672_), .Y(u5__abc_81276_new_n673_));
AND2X2 AND2X2_4185 ( .A(u5__abc_81276_new_n673_), .B(u5__abc_81276_new_n414_), .Y(u5__abc_81276_new_n674_));
AND2X2 AND2X2_4186 ( .A(u5__abc_81276_new_n674_), .B(u5__abc_81276_new_n408_), .Y(u5__abc_81276_new_n675_));
AND2X2 AND2X2_4187 ( .A(u5__abc_81276_new_n675_), .B(u5__abc_81276_new_n401__bF_buf2), .Y(u5__abc_81276_new_n676_));
AND2X2 AND2X2_4188 ( .A(u5__abc_81276_new_n676_), .B(u5__abc_81276_new_n448__bF_buf4), .Y(u5__abc_81276_new_n677_));
AND2X2 AND2X2_4189 ( .A(u5__abc_81276_new_n677_), .B(u5__abc_81276_new_n523__bF_buf4), .Y(u5__abc_81276_new_n678_));
AND2X2 AND2X2_419 ( .A(u0__abc_76628_new_n1169__bF_buf4), .B(u0__abc_76628_new_n1726_), .Y(u0__abc_76628_new_n1727_));
AND2X2 AND2X2_4190 ( .A(u5__abc_81276_new_n409_), .B(u5_state_50_), .Y(u5__abc_81276_new_n679_));
AND2X2 AND2X2_4191 ( .A(u5__abc_81276_new_n490__bF_buf10), .B(u5__abc_81276_new_n679_), .Y(u5__abc_81276_new_n680_));
AND2X2 AND2X2_4192 ( .A(u5__abc_81276_new_n680_), .B(u5__abc_81276_new_n414_), .Y(u5__abc_81276_new_n681_));
AND2X2 AND2X2_4193 ( .A(u5__abc_81276_new_n681_), .B(u5__abc_81276_new_n408_), .Y(u5__abc_81276_new_n682_));
AND2X2 AND2X2_4194 ( .A(u5__abc_81276_new_n682_), .B(u5__abc_81276_new_n401__bF_buf1), .Y(u5__abc_81276_new_n683_));
AND2X2 AND2X2_4195 ( .A(u5__abc_81276_new_n683_), .B(u5__abc_81276_new_n448__bF_buf3), .Y(u5__abc_81276_new_n684_));
AND2X2 AND2X2_4196 ( .A(u5__abc_81276_new_n684_), .B(u5__abc_81276_new_n523__bF_buf3), .Y(u5__abc_81276_new_n685_));
AND2X2 AND2X2_4197 ( .A(u5__abc_81276_new_n468_), .B(u5_state_4_), .Y(u5__abc_81276_new_n688_));
AND2X2 AND2X2_4198 ( .A(u5__abc_81276_new_n467_), .B(u5__abc_81276_new_n490__bF_buf9), .Y(u5__abc_81276_new_n689_));
AND2X2 AND2X2_4199 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n689_), .Y(u5__abc_81276_new_n690_));
AND2X2 AND2X2_42 ( .A(_abc_85006_new_n362_), .B(_abc_85006_new_n363_), .Y(tms_s_24_));
AND2X2 AND2X2_420 ( .A(u0__abc_76628_new_n1725_), .B(u0__abc_76628_new_n1727_), .Y(u0__abc_76628_new_n1728_));
AND2X2 AND2X2_4200 ( .A(u5__abc_81276_new_n690_), .B(u5__abc_81276_new_n688_), .Y(u5__abc_81276_new_n691_));
AND2X2 AND2X2_4201 ( .A(u5__abc_81276_new_n691_), .B(u5__abc_81276_new_n464__bF_buf2), .Y(u5__abc_81276_new_n692_));
AND2X2 AND2X2_4202 ( .A(u5__abc_81276_new_n449__bF_buf2), .B(u5__abc_81276_new_n692_), .Y(u5__abc_81276_new_n693_));
AND2X2 AND2X2_4203 ( .A(u5__abc_81276_new_n693_), .B(u5__abc_81276_new_n522__bF_buf3), .Y(u5__abc_81276_new_n694_));
AND2X2 AND2X2_4204 ( .A(u5__abc_81276_new_n490__bF_buf8), .B(u5_state_49_), .Y(u5__abc_81276_new_n696_));
AND2X2 AND2X2_4205 ( .A(u5__abc_81276_new_n411_), .B(u5__abc_81276_new_n413_), .Y(u5__abc_81276_new_n697_));
AND2X2 AND2X2_4206 ( .A(u5__abc_81276_new_n408_), .B(u5__abc_81276_new_n697_), .Y(u5__abc_81276_new_n698_));
AND2X2 AND2X2_4207 ( .A(u5__abc_81276_new_n401__bF_buf0), .B(u5__abc_81276_new_n698_), .Y(u5__abc_81276_new_n699_));
AND2X2 AND2X2_4208 ( .A(u5__abc_81276_new_n699_), .B(u5__abc_81276_new_n696_), .Y(u5__abc_81276_new_n700_));
AND2X2 AND2X2_4209 ( .A(u5__abc_81276_new_n700_), .B(u5__abc_81276_new_n448__bF_buf2), .Y(u5__abc_81276_new_n701_));
AND2X2 AND2X2_421 ( .A(u0__abc_76628_new_n1170__bF_buf4), .B(sp_tms_23_), .Y(u0__abc_76628_new_n1730_));
AND2X2 AND2X2_4210 ( .A(u5__abc_81276_new_n701_), .B(u5__abc_81276_new_n523__bF_buf2), .Y(u5__abc_81276_new_n702_));
AND2X2 AND2X2_4211 ( .A(u5__abc_81276_new_n695_), .B(u5__abc_81276_new_n703_), .Y(u5__abc_81276_new_n704_));
AND2X2 AND2X2_4212 ( .A(u5__abc_81276_new_n687_), .B(u5__abc_81276_new_n704_), .Y(u5__abc_81276_new_n705_));
AND2X2 AND2X2_4213 ( .A(u5__abc_81276_new_n417__bF_buf3), .B(u5__abc_81276_new_n447_), .Y(u5__abc_81276_new_n706_));
AND2X2 AND2X2_4214 ( .A(u5__abc_81276_new_n490__bF_buf7), .B(u5_state_40_), .Y(u5__abc_81276_new_n707_));
AND2X2 AND2X2_4215 ( .A(u5__abc_81276_new_n427_), .B(u5__abc_81276_new_n429_), .Y(u5__abc_81276_new_n708_));
AND2X2 AND2X2_4216 ( .A(u5__abc_81276_new_n707_), .B(u5__abc_81276_new_n708_), .Y(u5__abc_81276_new_n709_));
AND2X2 AND2X2_4217 ( .A(u5__abc_81276_new_n709_), .B(u5__abc_81276_new_n424_), .Y(u5__abc_81276_new_n710_));
AND2X2 AND2X2_4218 ( .A(u5__abc_81276_new_n523__bF_buf1), .B(u5__abc_81276_new_n710_), .Y(u5__abc_81276_new_n711_));
AND2X2 AND2X2_4219 ( .A(u5__abc_81276_new_n711_), .B(u5__abc_81276_new_n706_), .Y(u5__abc_81276_new_n712_));
AND2X2 AND2X2_422 ( .A(spec_req_cs_5_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1731_));
AND2X2 AND2X2_4220 ( .A(u5__abc_81276_new_n490__bF_buf6), .B(u5_state_48_), .Y(u5__abc_81276_new_n714_));
AND2X2 AND2X2_4221 ( .A(u5__abc_81276_new_n411_), .B(u5__abc_81276_new_n412_), .Y(u5__abc_81276_new_n715_));
AND2X2 AND2X2_4222 ( .A(u5__abc_81276_new_n408_), .B(u5__abc_81276_new_n715_), .Y(u5__abc_81276_new_n716_));
AND2X2 AND2X2_4223 ( .A(u5__abc_81276_new_n401__bF_buf3), .B(u5__abc_81276_new_n716_), .Y(u5__abc_81276_new_n717_));
AND2X2 AND2X2_4224 ( .A(u5__abc_81276_new_n717_), .B(u5__abc_81276_new_n714_), .Y(u5__abc_81276_new_n718_));
AND2X2 AND2X2_4225 ( .A(u5__abc_81276_new_n718_), .B(u5__abc_81276_new_n448__bF_buf1), .Y(u5__abc_81276_new_n719_));
AND2X2 AND2X2_4226 ( .A(u5__abc_81276_new_n719_), .B(u5__abc_81276_new_n523__bF_buf0), .Y(u5__abc_81276_new_n720_));
AND2X2 AND2X2_4227 ( .A(u5__abc_81276_new_n431_), .B(u5__abc_81276_new_n419_), .Y(u5__abc_81276_new_n722_));
AND2X2 AND2X2_4228 ( .A(u5__abc_81276_new_n490__bF_buf5), .B(u5_state_47_), .Y(u5__abc_81276_new_n723_));
AND2X2 AND2X2_4229 ( .A(u5__abc_81276_new_n723_), .B(u5__abc_81276_new_n423_), .Y(u5__abc_81276_new_n724_));
AND2X2 AND2X2_423 ( .A(u0__abc_76628_new_n1733_), .B(u0__abc_76628_new_n1179__bF_buf0), .Y(u0__abc_76628_new_n1734_));
AND2X2 AND2X2_4230 ( .A(u5__abc_81276_new_n722_), .B(u5__abc_81276_new_n724_), .Y(u5__abc_81276_new_n725_));
AND2X2 AND2X2_4231 ( .A(u5__abc_81276_new_n706_), .B(u5__abc_81276_new_n725_), .Y(u5__abc_81276_new_n726_));
AND2X2 AND2X2_4232 ( .A(u5__abc_81276_new_n726_), .B(u5__abc_81276_new_n523__bF_buf7), .Y(u5__abc_81276_new_n727_));
AND2X2 AND2X2_4233 ( .A(u5__abc_81276_new_n728_), .B(u5__abc_81276_new_n721_), .Y(u5__abc_81276_new_n729_));
AND2X2 AND2X2_4234 ( .A(u5__abc_81276_new_n446_), .B(u5__abc_81276_new_n434_), .Y(u5__abc_81276_new_n730_));
AND2X2 AND2X2_4235 ( .A(u5__abc_81276_new_n490__bF_buf4), .B(u5_state_39_), .Y(u5__abc_81276_new_n731_));
AND2X2 AND2X2_4236 ( .A(u5__abc_81276_new_n731_), .B(u5__abc_81276_new_n438_), .Y(u5__abc_81276_new_n732_));
AND2X2 AND2X2_4237 ( .A(u5__abc_81276_new_n730_), .B(u5__abc_81276_new_n732_), .Y(u5__abc_81276_new_n733_));
AND2X2 AND2X2_4238 ( .A(u5__abc_81276_new_n523__bF_buf6), .B(u5__abc_81276_new_n733_), .Y(u5__abc_81276_new_n734_));
AND2X2 AND2X2_4239 ( .A(u5__abc_81276_new_n734_), .B(u5__abc_81276_new_n557_), .Y(u5__abc_81276_new_n735_));
AND2X2 AND2X2_424 ( .A(u0__abc_76628_new_n1734_), .B(u0__abc_76628_new_n1732_), .Y(u0__abc_76628_new_n1735_));
AND2X2 AND2X2_4240 ( .A(u5__abc_81276_new_n729_), .B(u5__abc_81276_new_n736_), .Y(u5__abc_81276_new_n737_));
AND2X2 AND2X2_4241 ( .A(u5__abc_81276_new_n737_), .B(u5__abc_81276_new_n713_), .Y(u5__abc_81276_new_n738_));
AND2X2 AND2X2_4242 ( .A(u5__abc_81276_new_n738_), .B(u5__abc_81276_new_n705_), .Y(u5__abc_81276_new_n739_));
AND2X2 AND2X2_4243 ( .A(u5__abc_81276_new_n490__bF_buf3), .B(u5_state_42_), .Y(u5__abc_81276_new_n740_));
AND2X2 AND2X2_4244 ( .A(u5__abc_81276_new_n430_), .B(u5__abc_81276_new_n425_), .Y(u5__abc_81276_new_n741_));
AND2X2 AND2X2_4245 ( .A(u5__abc_81276_new_n740_), .B(u5__abc_81276_new_n741_), .Y(u5__abc_81276_new_n742_));
AND2X2 AND2X2_4246 ( .A(u5__abc_81276_new_n742_), .B(u5__abc_81276_new_n424_), .Y(u5__abc_81276_new_n743_));
AND2X2 AND2X2_4247 ( .A(u5__abc_81276_new_n523__bF_buf5), .B(u5__abc_81276_new_n743_), .Y(u5__abc_81276_new_n744_));
AND2X2 AND2X2_4248 ( .A(u5__abc_81276_new_n744_), .B(u5__abc_81276_new_n706_), .Y(u5__abc_81276_new_n745_));
AND2X2 AND2X2_4249 ( .A(u5__abc_81276_new_n446_), .B(u5__abc_81276_new_n437_), .Y(u5__abc_81276_new_n747_));
AND2X2 AND2X2_425 ( .A(u0__abc_76628_new_n1736_), .B(u0__abc_76628_new_n1175__bF_buf0), .Y(u0__abc_76628_new_n1737_));
AND2X2 AND2X2_4250 ( .A(u5__abc_81276_new_n490__bF_buf2), .B(u5_state_37_), .Y(u5__abc_81276_new_n748_));
AND2X2 AND2X2_4251 ( .A(u5__abc_81276_new_n748_), .B(u5__abc_81276_new_n435_), .Y(u5__abc_81276_new_n749_));
AND2X2 AND2X2_4252 ( .A(u5__abc_81276_new_n747_), .B(u5__abc_81276_new_n749_), .Y(u5__abc_81276_new_n750_));
AND2X2 AND2X2_4253 ( .A(u5__abc_81276_new_n523__bF_buf4), .B(u5__abc_81276_new_n750_), .Y(u5__abc_81276_new_n751_));
AND2X2 AND2X2_4254 ( .A(u5__abc_81276_new_n751_), .B(u5__abc_81276_new_n557_), .Y(u5__abc_81276_new_n752_));
AND2X2 AND2X2_4255 ( .A(u5__abc_81276_new_n746_), .B(u5__abc_81276_new_n753_), .Y(u5__abc_81276_new_n754_));
AND2X2 AND2X2_4256 ( .A(u5__abc_81276_new_n431_), .B(u5__abc_81276_new_n418_), .Y(u5__abc_81276_new_n755_));
AND2X2 AND2X2_4257 ( .A(u5__abc_81276_new_n490__bF_buf1), .B(u5_state_46_), .Y(u5__abc_81276_new_n756_));
AND2X2 AND2X2_4258 ( .A(u5__abc_81276_new_n756_), .B(u5__abc_81276_new_n423_), .Y(u5__abc_81276_new_n757_));
AND2X2 AND2X2_4259 ( .A(u5__abc_81276_new_n447_), .B(u5__abc_81276_new_n757_), .Y(u5__abc_81276_new_n758_));
AND2X2 AND2X2_426 ( .A(spec_req_cs_4_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1738_));
AND2X2 AND2X2_4260 ( .A(u5__abc_81276_new_n758_), .B(u5__abc_81276_new_n755_), .Y(u5__abc_81276_new_n759_));
AND2X2 AND2X2_4261 ( .A(u5__abc_81276_new_n759_), .B(u5__abc_81276_new_n417__bF_buf2), .Y(u5__abc_81276_new_n760_));
AND2X2 AND2X2_4262 ( .A(u5__abc_81276_new_n760_), .B(u5__abc_81276_new_n523__bF_buf3), .Y(u5__abc_81276_new_n761_));
AND2X2 AND2X2_4263 ( .A(u5__abc_81276_new_n431_), .B(u5__abc_81276_new_n422_), .Y(u5__abc_81276_new_n762_));
AND2X2 AND2X2_4264 ( .A(u5__abc_81276_new_n490__bF_buf0), .B(u5_state_45_), .Y(u5__abc_81276_new_n763_));
AND2X2 AND2X2_4265 ( .A(u5__abc_81276_new_n763_), .B(u5__abc_81276_new_n420_), .Y(u5__abc_81276_new_n764_));
AND2X2 AND2X2_4266 ( .A(u5__abc_81276_new_n762_), .B(u5__abc_81276_new_n764_), .Y(u5__abc_81276_new_n765_));
AND2X2 AND2X2_4267 ( .A(u5__abc_81276_new_n523__bF_buf2), .B(u5__abc_81276_new_n765_), .Y(u5__abc_81276_new_n766_));
AND2X2 AND2X2_4268 ( .A(u5__abc_81276_new_n766_), .B(u5__abc_81276_new_n706_), .Y(u5__abc_81276_new_n767_));
AND2X2 AND2X2_4269 ( .A(u5__abc_81276_new_n446_), .B(u5__abc_81276_new_n433_), .Y(u5__abc_81276_new_n770_));
AND2X2 AND2X2_427 ( .A(u0__abc_76628_new_n1739_), .B(u0__abc_76628_new_n1174__bF_buf0), .Y(u0__abc_76628_new_n1740_));
AND2X2 AND2X2_4270 ( .A(u5__abc_81276_new_n490__bF_buf10), .B(u5_state_38_), .Y(u5__abc_81276_new_n771_));
AND2X2 AND2X2_4271 ( .A(u5__abc_81276_new_n771_), .B(u5__abc_81276_new_n438_), .Y(u5__abc_81276_new_n772_));
AND2X2 AND2X2_4272 ( .A(u5__abc_81276_new_n770_), .B(u5__abc_81276_new_n772_), .Y(u5__abc_81276_new_n773_));
AND2X2 AND2X2_4273 ( .A(u5__abc_81276_new_n523__bF_buf1), .B(u5__abc_81276_new_n773_), .Y(u5__abc_81276_new_n774_));
AND2X2 AND2X2_4274 ( .A(u5__abc_81276_new_n774_), .B(u5__abc_81276_new_n557_), .Y(u5__abc_81276_new_n775_));
AND2X2 AND2X2_4275 ( .A(u5__abc_81276_new_n431_), .B(u5__abc_81276_new_n421_), .Y(u5__abc_81276_new_n777_));
AND2X2 AND2X2_4276 ( .A(u5__abc_81276_new_n490__bF_buf9), .B(u5_state_44_), .Y(u5__abc_81276_new_n778_));
AND2X2 AND2X2_4277 ( .A(u5__abc_81276_new_n778_), .B(u5__abc_81276_new_n420_), .Y(u5__abc_81276_new_n779_));
AND2X2 AND2X2_4278 ( .A(u5__abc_81276_new_n777_), .B(u5__abc_81276_new_n779_), .Y(u5__abc_81276_new_n780_));
AND2X2 AND2X2_4279 ( .A(u5__abc_81276_new_n523__bF_buf0), .B(u5__abc_81276_new_n780_), .Y(u5__abc_81276_new_n781_));
AND2X2 AND2X2_428 ( .A(spec_req_cs_3_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1741_));
AND2X2 AND2X2_4280 ( .A(u5__abc_81276_new_n781_), .B(u5__abc_81276_new_n706_), .Y(u5__abc_81276_new_n782_));
AND2X2 AND2X2_4281 ( .A(u5__abc_81276_new_n776_), .B(u5__abc_81276_new_n783_), .Y(u5__abc_81276_new_n784_));
AND2X2 AND2X2_4282 ( .A(u5__abc_81276_new_n769_), .B(u5__abc_81276_new_n784_), .Y(u5__abc_81276_new_n785_));
AND2X2 AND2X2_4283 ( .A(u5__abc_81276_new_n490__bF_buf8), .B(u5_state_43_), .Y(u5__abc_81276_new_n786_));
AND2X2 AND2X2_4284 ( .A(u5__abc_81276_new_n430_), .B(u5__abc_81276_new_n426_), .Y(u5__abc_81276_new_n787_));
AND2X2 AND2X2_4285 ( .A(u5__abc_81276_new_n424_), .B(u5__abc_81276_new_n787_), .Y(u5__abc_81276_new_n788_));
AND2X2 AND2X2_4286 ( .A(u5__abc_81276_new_n788_), .B(u5__abc_81276_new_n786_), .Y(u5__abc_81276_new_n789_));
AND2X2 AND2X2_4287 ( .A(u5__abc_81276_new_n523__bF_buf7), .B(u5__abc_81276_new_n789_), .Y(u5__abc_81276_new_n790_));
AND2X2 AND2X2_4288 ( .A(u5__abc_81276_new_n790_), .B(u5__abc_81276_new_n706_), .Y(u5__abc_81276_new_n791_));
AND2X2 AND2X2_4289 ( .A(u5__abc_81276_new_n490__bF_buf7), .B(u5_state_41_), .Y(u5__abc_81276_new_n793_));
AND2X2 AND2X2_429 ( .A(u0__abc_76628_new_n1742_), .B(u0__abc_76628_new_n1173__bF_buf0), .Y(u0__abc_76628_new_n1743_));
AND2X2 AND2X2_4290 ( .A(u5__abc_81276_new_n427_), .B(u5__abc_81276_new_n428_), .Y(u5__abc_81276_new_n794_));
AND2X2 AND2X2_4291 ( .A(u5__abc_81276_new_n424_), .B(u5__abc_81276_new_n794_), .Y(u5__abc_81276_new_n795_));
AND2X2 AND2X2_4292 ( .A(u5__abc_81276_new_n447_), .B(u5__abc_81276_new_n795_), .Y(u5__abc_81276_new_n796_));
AND2X2 AND2X2_4293 ( .A(u5__abc_81276_new_n796_), .B(u5__abc_81276_new_n793_), .Y(u5__abc_81276_new_n797_));
AND2X2 AND2X2_4294 ( .A(u5__abc_81276_new_n797_), .B(u5__abc_81276_new_n417__bF_buf1), .Y(u5__abc_81276_new_n798_));
AND2X2 AND2X2_4295 ( .A(u5__abc_81276_new_n798_), .B(u5__abc_81276_new_n523__bF_buf6), .Y(u5__abc_81276_new_n799_));
AND2X2 AND2X2_4296 ( .A(u5__abc_81276_new_n792_), .B(u5__abc_81276_new_n800_), .Y(u5__abc_81276_new_n801_));
AND2X2 AND2X2_4297 ( .A(u5__abc_81276_new_n785_), .B(u5__abc_81276_new_n801_), .Y(u5__abc_81276_new_n802_));
AND2X2 AND2X2_4298 ( .A(u5__abc_81276_new_n802_), .B(u5__abc_81276_new_n754_), .Y(u5__abc_81276_new_n803_));
AND2X2 AND2X2_4299 ( .A(u5__abc_81276_new_n803_), .B(u5__abc_81276_new_n739_), .Y(u5__abc_81276_new_n804_));
AND2X2 AND2X2_43 ( .A(_abc_85006_new_n365_), .B(_abc_85006_new_n366_), .Y(tms_s_25_));
AND2X2 AND2X2_430 ( .A(spec_req_cs_2_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1744_));
AND2X2 AND2X2_4300 ( .A(u5__abc_81276_new_n490__bF_buf6), .B(u5_state_8_), .Y(u5__abc_81276_new_n805_));
AND2X2 AND2X2_4301 ( .A(u5__abc_81276_new_n459_), .B(u5__abc_81276_new_n460_), .Y(u5__abc_81276_new_n806_));
AND2X2 AND2X2_4302 ( .A(u5__abc_81276_new_n456_), .B(u5__abc_81276_new_n806_), .Y(u5__abc_81276_new_n807_));
AND2X2 AND2X2_4303 ( .A(u5__abc_81276_new_n807_), .B(u5__abc_81276_new_n805_), .Y(u5__abc_81276_new_n808_));
AND2X2 AND2X2_4304 ( .A(u5__abc_81276_new_n808_), .B(u5__abc_81276_new_n479__bF_buf2), .Y(u5__abc_81276_new_n809_));
AND2X2 AND2X2_4305 ( .A(u5__abc_81276_new_n449__bF_buf1), .B(u5__abc_81276_new_n809_), .Y(u5__abc_81276_new_n810_));
AND2X2 AND2X2_4306 ( .A(u5__abc_81276_new_n810_), .B(u5__abc_81276_new_n522__bF_buf2), .Y(u5__abc_81276_new_n811_));
AND2X2 AND2X2_4307 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n466_), .Y(u5__abc_81276_new_n813_));
AND2X2 AND2X2_4308 ( .A(u5__abc_81276_new_n490__bF_buf5), .B(u5_state_7_), .Y(u5__abc_81276_new_n814_));
AND2X2 AND2X2_4309 ( .A(u5__abc_81276_new_n814_), .B(u5__abc_81276_new_n470_), .Y(u5__abc_81276_new_n815_));
AND2X2 AND2X2_431 ( .A(u0__abc_76628_new_n1745_), .B(u0__abc_76628_new_n1172__bF_buf0), .Y(u0__abc_76628_new_n1746_));
AND2X2 AND2X2_4310 ( .A(u5__abc_81276_new_n813_), .B(u5__abc_81276_new_n815_), .Y(u5__abc_81276_new_n816_));
AND2X2 AND2X2_4311 ( .A(u5__abc_81276_new_n816_), .B(u5__abc_81276_new_n464__bF_buf1), .Y(u5__abc_81276_new_n817_));
AND2X2 AND2X2_4312 ( .A(u5__abc_81276_new_n449__bF_buf0), .B(u5__abc_81276_new_n817_), .Y(u5__abc_81276_new_n818_));
AND2X2 AND2X2_4313 ( .A(u5__abc_81276_new_n818_), .B(u5__abc_81276_new_n522__bF_buf1), .Y(u5__abc_81276_new_n819_));
AND2X2 AND2X2_4314 ( .A(u5__abc_81276_new_n812_), .B(u5__abc_81276_new_n820_), .Y(u5__abc_81276_new_n821_));
AND2X2 AND2X2_4315 ( .A(u5__abc_81276_new_n490__bF_buf4), .B(u5_state_9_), .Y(u5__abc_81276_new_n822_));
AND2X2 AND2X2_4316 ( .A(u5__abc_81276_new_n459_), .B(u5__abc_81276_new_n461_), .Y(u5__abc_81276_new_n823_));
AND2X2 AND2X2_4317 ( .A(u5__abc_81276_new_n456_), .B(u5__abc_81276_new_n823_), .Y(u5__abc_81276_new_n824_));
AND2X2 AND2X2_4318 ( .A(u5__abc_81276_new_n824_), .B(u5__abc_81276_new_n822_), .Y(u5__abc_81276_new_n825_));
AND2X2 AND2X2_4319 ( .A(u5__abc_81276_new_n825_), .B(u5__abc_81276_new_n479__bF_buf1), .Y(u5__abc_81276_new_n826_));
AND2X2 AND2X2_432 ( .A(spec_req_cs_1_bF_buf3_), .B(u0_tms1_23_), .Y(u0__abc_76628_new_n1747_));
AND2X2 AND2X2_4320 ( .A(u5__abc_81276_new_n449__bF_buf7), .B(u5__abc_81276_new_n826_), .Y(u5__abc_81276_new_n827_));
AND2X2 AND2X2_4321 ( .A(u5__abc_81276_new_n827_), .B(u5__abc_81276_new_n522__bF_buf0), .Y(u5__abc_81276_new_n828_));
AND2X2 AND2X2_4322 ( .A(u5__abc_81276_new_n490__bF_buf3), .B(u5_state_13_), .Y(u5__abc_81276_new_n830_));
AND2X2 AND2X2_4323 ( .A(u5__abc_81276_new_n463_), .B(u5__abc_81276_new_n453_), .Y(u5__abc_81276_new_n831_));
AND2X2 AND2X2_4324 ( .A(u5__abc_81276_new_n831_), .B(u5__abc_81276_new_n830_), .Y(u5__abc_81276_new_n832_));
AND2X2 AND2X2_4325 ( .A(u5__abc_81276_new_n479__bF_buf0), .B(u5__abc_81276_new_n452_), .Y(u5__abc_81276_new_n833_));
AND2X2 AND2X2_4326 ( .A(u5__abc_81276_new_n833_), .B(u5__abc_81276_new_n832_), .Y(u5__abc_81276_new_n834_));
AND2X2 AND2X2_4327 ( .A(u5__abc_81276_new_n834_), .B(u5__abc_81276_new_n522__bF_buf4), .Y(u5__abc_81276_new_n835_));
AND2X2 AND2X2_4328 ( .A(u5__abc_81276_new_n835_), .B(u5__abc_81276_new_n449__bF_buf6), .Y(u5__abc_81276_new_n836_));
AND2X2 AND2X2_4329 ( .A(u5__abc_81276_new_n829_), .B(u5__abc_81276_new_n837_), .Y(u5__abc_81276_new_n838_));
AND2X2 AND2X2_433 ( .A(u0__abc_76628_new_n1169__bF_buf3), .B(u0__abc_76628_new_n1750_), .Y(u0__abc_76628_new_n1751_));
AND2X2 AND2X2_4330 ( .A(u5__abc_81276_new_n462_), .B(u5__abc_81276_new_n457_), .Y(u5__abc_81276_new_n839_));
AND2X2 AND2X2_4331 ( .A(u5__abc_81276_new_n456_), .B(u5__abc_81276_new_n839_), .Y(u5__abc_81276_new_n840_));
AND2X2 AND2X2_4332 ( .A(u5__abc_81276_new_n479__bF_buf3), .B(u5__abc_81276_new_n840_), .Y(u5__abc_81276_new_n841_));
AND2X2 AND2X2_4333 ( .A(u5__abc_81276_new_n522__bF_buf3), .B(u5__abc_81276_new_n841_), .Y(u5__abc_81276_new_n842_));
AND2X2 AND2X2_4334 ( .A(u5__abc_81276_new_n490__bF_buf2), .B(u5_state_10_), .Y(u5__abc_81276_new_n843_));
AND2X2 AND2X2_4335 ( .A(u5__abc_81276_new_n449__bF_buf5), .B(u5__abc_81276_new_n843_), .Y(u5__abc_81276_new_n844_));
AND2X2 AND2X2_4336 ( .A(u5__abc_81276_new_n844_), .B(u5__abc_81276_new_n842_), .Y(u5__abc_81276_new_n845_));
AND2X2 AND2X2_4337 ( .A(u5__abc_81276_new_n490__bF_buf1), .B(u5_state_14_), .Y(u5__abc_81276_new_n847_));
AND2X2 AND2X2_4338 ( .A(u5__abc_81276_new_n847_), .B(u5__abc_81276_new_n455_), .Y(u5__abc_81276_new_n848_));
AND2X2 AND2X2_4339 ( .A(u5__abc_81276_new_n479__bF_buf2), .B(u5__abc_81276_new_n848_), .Y(u5__abc_81276_new_n849_));
AND2X2 AND2X2_434 ( .A(u0__abc_76628_new_n1749_), .B(u0__abc_76628_new_n1751_), .Y(u0__abc_76628_new_n1752_));
AND2X2 AND2X2_4340 ( .A(u5__abc_81276_new_n522__bF_buf2), .B(u5__abc_81276_new_n849_), .Y(u5__abc_81276_new_n850_));
AND2X2 AND2X2_4341 ( .A(u5__abc_81276_new_n463_), .B(u5__abc_81276_new_n450_), .Y(u5__abc_81276_new_n851_));
AND2X2 AND2X2_4342 ( .A(u5__abc_81276_new_n449__bF_buf4), .B(u5__abc_81276_new_n851_), .Y(u5__abc_81276_new_n852_));
AND2X2 AND2X2_4343 ( .A(u5__abc_81276_new_n852_), .B(u5__abc_81276_new_n850_), .Y(u5__abc_81276_new_n853_));
AND2X2 AND2X2_4344 ( .A(u5__abc_81276_new_n846_), .B(u5__abc_81276_new_n854_), .Y(u5__abc_81276_new_n855_));
AND2X2 AND2X2_4345 ( .A(u5__abc_81276_new_n855_), .B(u5__abc_81276_new_n838_), .Y(u5__abc_81276_new_n856_));
AND2X2 AND2X2_4346 ( .A(u5__abc_81276_new_n469_), .B(u5_state_5_), .Y(u5__abc_81276_new_n857_));
AND2X2 AND2X2_4347 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n857_), .Y(u5__abc_81276_new_n858_));
AND2X2 AND2X2_4348 ( .A(u5__abc_81276_new_n464__bF_buf0), .B(u5__abc_81276_new_n858_), .Y(u5__abc_81276_new_n859_));
AND2X2 AND2X2_4349 ( .A(u5__abc_81276_new_n859_), .B(u5__abc_81276_new_n689_), .Y(u5__abc_81276_new_n860_));
AND2X2 AND2X2_435 ( .A(u0__abc_76628_new_n1170__bF_buf3), .B(sp_tms_24_), .Y(u0__abc_76628_new_n1754_));
AND2X2 AND2X2_4350 ( .A(u5__abc_81276_new_n449__bF_buf3), .B(u5__abc_81276_new_n860_), .Y(u5__abc_81276_new_n861_));
AND2X2 AND2X2_4351 ( .A(u5__abc_81276_new_n861_), .B(u5__abc_81276_new_n522__bF_buf1), .Y(u5__abc_81276_new_n862_));
AND2X2 AND2X2_4352 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n465_), .Y(u5__abc_81276_new_n864_));
AND2X2 AND2X2_4353 ( .A(u5__abc_81276_new_n490__bF_buf0), .B(u5_state_6_), .Y(u5__abc_81276_new_n865_));
AND2X2 AND2X2_4354 ( .A(u5__abc_81276_new_n865_), .B(u5__abc_81276_new_n470_), .Y(u5__abc_81276_new_n866_));
AND2X2 AND2X2_4355 ( .A(u5__abc_81276_new_n464__bF_buf3), .B(u5__abc_81276_new_n866_), .Y(u5__abc_81276_new_n867_));
AND2X2 AND2X2_4356 ( .A(u5__abc_81276_new_n867_), .B(u5__abc_81276_new_n864_), .Y(u5__abc_81276_new_n868_));
AND2X2 AND2X2_4357 ( .A(u5__abc_81276_new_n868_), .B(u5__abc_81276_new_n522__bF_buf0), .Y(u5__abc_81276_new_n869_));
AND2X2 AND2X2_4358 ( .A(u5__abc_81276_new_n869_), .B(u5__abc_81276_new_n449__bF_buf2), .Y(u5__abc_81276_new_n870_));
AND2X2 AND2X2_4359 ( .A(u5__abc_81276_new_n863_), .B(u5__abc_81276_new_n871_), .Y(u5__abc_81276_new_n872_));
AND2X2 AND2X2_436 ( .A(spec_req_cs_5_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1755_));
AND2X2 AND2X2_4360 ( .A(u5__abc_81276_new_n856_), .B(u5__abc_81276_new_n872_), .Y(u5__abc_81276_new_n873_));
AND2X2 AND2X2_4361 ( .A(u5__abc_81276_new_n873_), .B(u5__abc_81276_new_n821_), .Y(u5__abc_81276_new_n874_));
AND2X2 AND2X2_4362 ( .A(u5__abc_81276_new_n490__bF_buf10), .B(u5_state_1_), .Y(u5__abc_81276_new_n875_));
AND2X2 AND2X2_4363 ( .A(u5__abc_81276_new_n474_), .B(u5__abc_81276_new_n476_), .Y(u5__abc_81276_new_n876_));
AND2X2 AND2X2_4364 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n876_), .Y(u5__abc_81276_new_n877_));
AND2X2 AND2X2_4365 ( .A(u5__abc_81276_new_n464__bF_buf2), .B(u5__abc_81276_new_n877_), .Y(u5__abc_81276_new_n878_));
AND2X2 AND2X2_4366 ( .A(u5__abc_81276_new_n878_), .B(u5__abc_81276_new_n875_), .Y(u5__abc_81276_new_n879_));
AND2X2 AND2X2_4367 ( .A(u5__abc_81276_new_n879_), .B(u5__abc_81276_new_n522__bF_buf4), .Y(u5__abc_81276_new_n880_));
AND2X2 AND2X2_4368 ( .A(u5__abc_81276_new_n880_), .B(u5__abc_81276_new_n449__bF_buf1), .Y(u5__abc_81276_new_n881_));
AND2X2 AND2X2_4369 ( .A(u5__abc_81276_new_n490__bF_buf9), .B(u5_state_0_), .Y(u5__abc_81276_new_n883_));
AND2X2 AND2X2_437 ( .A(u0__abc_76628_new_n1757_), .B(u0__abc_76628_new_n1179__bF_buf5), .Y(u0__abc_76628_new_n1758_));
AND2X2 AND2X2_4370 ( .A(u5__abc_81276_new_n474_), .B(u5__abc_81276_new_n475_), .Y(u5__abc_81276_new_n884_));
AND2X2 AND2X2_4371 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n884_), .Y(u5__abc_81276_new_n885_));
AND2X2 AND2X2_4372 ( .A(u5__abc_81276_new_n464__bF_buf1), .B(u5__abc_81276_new_n885_), .Y(u5__abc_81276_new_n886_));
AND2X2 AND2X2_4373 ( .A(u5__abc_81276_new_n886_), .B(u5__abc_81276_new_n883_), .Y(u5__abc_81276_new_n887_));
AND2X2 AND2X2_4374 ( .A(u5__abc_81276_new_n887_), .B(u5__abc_81276_new_n522__bF_buf3), .Y(u5__abc_81276_new_n888_));
AND2X2 AND2X2_4375 ( .A(u5__abc_81276_new_n888_), .B(u5__abc_81276_new_n449__bF_buf0), .Y(u5__abc_81276_new_n889_));
AND2X2 AND2X2_4376 ( .A(u5__abc_81276_new_n882_), .B(u5__abc_81276_new_n890_), .Y(u5__abc_81276_new_n891_));
AND2X2 AND2X2_4377 ( .A(u5__abc_81276_new_n511_), .B(u5__abc_81276_new_n518_), .Y(u5__abc_81276_new_n892_));
AND2X2 AND2X2_4378 ( .A(u5__abc_81276_new_n508_), .B(u5__abc_81276_new_n892_), .Y(u5__abc_81276_new_n893_));
AND2X2 AND2X2_4379 ( .A(u5__abc_81276_new_n490__bF_buf8), .B(u5_state_31_), .Y(u5__abc_81276_new_n894_));
AND2X2 AND2X2_438 ( .A(u0__abc_76628_new_n1758_), .B(u0__abc_76628_new_n1756_), .Y(u0__abc_76628_new_n1759_));
AND2X2 AND2X2_4380 ( .A(u5__abc_81276_new_n893_), .B(u5__abc_81276_new_n894_), .Y(u5__abc_81276_new_n895_));
AND2X2 AND2X2_4381 ( .A(u5__abc_81276_new_n895_), .B(u5__abc_81276_new_n517_), .Y(u5__abc_81276_new_n896_));
AND2X2 AND2X2_4382 ( .A(u5__abc_81276_new_n449__bF_buf7), .B(u5__abc_81276_new_n896_), .Y(u5__abc_81276_new_n897_));
AND2X2 AND2X2_4383 ( .A(u5__abc_81276_new_n897_), .B(u5__abc_81276_new_n480__bF_buf0), .Y(u5__abc_81276_new_n898_));
AND2X2 AND2X2_4384 ( .A(u5__abc_81276_new_n490__bF_buf7), .B(u5_state_34_), .Y(u5__abc_81276_new_n900_));
AND2X2 AND2X2_4385 ( .A(u5__abc_81276_new_n445_), .B(u5__abc_81276_new_n440_), .Y(u5__abc_81276_new_n901_));
AND2X2 AND2X2_4386 ( .A(u5__abc_81276_new_n439_), .B(u5__abc_81276_new_n901_), .Y(u5__abc_81276_new_n902_));
AND2X2 AND2X2_4387 ( .A(u5__abc_81276_new_n902_), .B(u5__abc_81276_new_n900_), .Y(u5__abc_81276_new_n903_));
AND2X2 AND2X2_4388 ( .A(u5__abc_81276_new_n523__bF_buf5), .B(u5__abc_81276_new_n903_), .Y(u5__abc_81276_new_n904_));
AND2X2 AND2X2_4389 ( .A(u5__abc_81276_new_n904_), .B(u5__abc_81276_new_n557_), .Y(u5__abc_81276_new_n905_));
AND2X2 AND2X2_439 ( .A(u0__abc_76628_new_n1760_), .B(u0__abc_76628_new_n1175__bF_buf5), .Y(u0__abc_76628_new_n1761_));
AND2X2 AND2X2_4390 ( .A(u5__abc_81276_new_n899_), .B(u5__abc_81276_new_n906_), .Y(u5__abc_81276_new_n907_));
AND2X2 AND2X2_4391 ( .A(u5__abc_81276_new_n907_), .B(u5__abc_81276_new_n891_), .Y(u5__abc_81276_new_n908_));
AND2X2 AND2X2_4392 ( .A(u5__abc_81276_new_n490__bF_buf6), .B(u5_state_33_), .Y(u5__abc_81276_new_n909_));
AND2X2 AND2X2_4393 ( .A(u5__abc_81276_new_n442_), .B(u5__abc_81276_new_n443_), .Y(u5__abc_81276_new_n910_));
AND2X2 AND2X2_4394 ( .A(u5__abc_81276_new_n439_), .B(u5__abc_81276_new_n910_), .Y(u5__abc_81276_new_n911_));
AND2X2 AND2X2_4395 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n911_), .Y(u5__abc_81276_new_n912_));
AND2X2 AND2X2_4396 ( .A(u5__abc_81276_new_n912_), .B(u5__abc_81276_new_n909_), .Y(u5__abc_81276_new_n913_));
AND2X2 AND2X2_4397 ( .A(u5__abc_81276_new_n913_), .B(u5__abc_81276_new_n417__bF_buf0), .Y(u5__abc_81276_new_n914_));
AND2X2 AND2X2_4398 ( .A(u5__abc_81276_new_n914_), .B(u5__abc_81276_new_n523__bF_buf4), .Y(u5__abc_81276_new_n915_));
AND2X2 AND2X2_4399 ( .A(u5__abc_81276_new_n922_), .B(u5__abc_81276_new_n521__bF_buf3), .Y(u5__abc_81276_new_n923_));
AND2X2 AND2X2_44 ( .A(_abc_85006_new_n368_), .B(_abc_85006_new_n369_), .Y(tms_s_26_));
AND2X2 AND2X2_440 ( .A(spec_req_cs_4_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1762_));
AND2X2 AND2X2_4400 ( .A(u5__abc_81276_new_n480__bF_buf4), .B(u5__abc_81276_new_n659_), .Y(u5__abc_81276_new_n924_));
AND2X2 AND2X2_4401 ( .A(u5__abc_81276_new_n449__bF_buf6), .B(u5__abc_81276_new_n924_), .Y(u5__abc_81276_new_n925_));
AND2X2 AND2X2_4402 ( .A(u5__abc_81276_new_n925_), .B(u5__abc_81276_new_n923_), .Y(u5__abc_81276_new_n926_));
AND2X2 AND2X2_4403 ( .A(u5__abc_81276_new_n927_), .B(u5__abc_81276_new_n916_), .Y(u5__abc_81276_new_n928_));
AND2X2 AND2X2_4404 ( .A(u5__abc_81276_new_n463_), .B(u5__abc_81276_new_n454_), .Y(u5__abc_81276_new_n929_));
AND2X2 AND2X2_4405 ( .A(u5__abc_81276_new_n490__bF_buf5), .B(u5_state_12_), .Y(u5__abc_81276_new_n930_));
AND2X2 AND2X2_4406 ( .A(u5__abc_81276_new_n930_), .B(u5__abc_81276_new_n452_), .Y(u5__abc_81276_new_n931_));
AND2X2 AND2X2_4407 ( .A(u5__abc_81276_new_n929_), .B(u5__abc_81276_new_n931_), .Y(u5__abc_81276_new_n932_));
AND2X2 AND2X2_4408 ( .A(u5__abc_81276_new_n932_), .B(u5__abc_81276_new_n479__bF_buf1), .Y(u5__abc_81276_new_n933_));
AND2X2 AND2X2_4409 ( .A(u5__abc_81276_new_n449__bF_buf5), .B(u5__abc_81276_new_n933_), .Y(u5__abc_81276_new_n934_));
AND2X2 AND2X2_441 ( .A(u0__abc_76628_new_n1763_), .B(u0__abc_76628_new_n1174__bF_buf5), .Y(u0__abc_76628_new_n1764_));
AND2X2 AND2X2_4410 ( .A(u5__abc_81276_new_n934_), .B(u5__abc_81276_new_n522__bF_buf2), .Y(u5__abc_81276_new_n935_));
AND2X2 AND2X2_4411 ( .A(u5__abc_81276_new_n463_), .B(u5__abc_81276_new_n451_), .Y(u5__abc_81276_new_n937_));
AND2X2 AND2X2_4412 ( .A(u5__abc_81276_new_n490__bF_buf4), .B(u5_state_15_), .Y(u5__abc_81276_new_n938_));
AND2X2 AND2X2_4413 ( .A(u5__abc_81276_new_n938_), .B(u5__abc_81276_new_n455_), .Y(u5__abc_81276_new_n939_));
AND2X2 AND2X2_4414 ( .A(u5__abc_81276_new_n937_), .B(u5__abc_81276_new_n939_), .Y(u5__abc_81276_new_n940_));
AND2X2 AND2X2_4415 ( .A(u5__abc_81276_new_n940_), .B(u5__abc_81276_new_n479__bF_buf0), .Y(u5__abc_81276_new_n941_));
AND2X2 AND2X2_4416 ( .A(u5__abc_81276_new_n449__bF_buf4), .B(u5__abc_81276_new_n941_), .Y(u5__abc_81276_new_n942_));
AND2X2 AND2X2_4417 ( .A(u5__abc_81276_new_n942_), .B(u5__abc_81276_new_n522__bF_buf1), .Y(u5__abc_81276_new_n943_));
AND2X2 AND2X2_4418 ( .A(u5__abc_81276_new_n936_), .B(u5__abc_81276_new_n944_), .Y(u5__abc_81276_new_n945_));
AND2X2 AND2X2_4419 ( .A(u5__abc_81276_new_n945_), .B(u5__abc_81276_new_n928_), .Y(u5__abc_81276_new_n946_));
AND2X2 AND2X2_442 ( .A(spec_req_cs_3_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1765_));
AND2X2 AND2X2_4420 ( .A(u5__abc_81276_new_n908_), .B(u5__abc_81276_new_n946_), .Y(u5__abc_81276_new_n947_));
AND2X2 AND2X2_4421 ( .A(u5__abc_81276_new_n449__bF_buf3), .B(u5__abc_81276_new_n523__bF_buf3), .Y(u5__abc_81276_new_n948_));
AND2X2 AND2X2_4422 ( .A(u5__abc_81276_new_n489_), .B(u5_state_65_), .Y(u5__abc_81276_new_n949_));
AND2X2 AND2X2_4423 ( .A(u5__abc_81276_new_n948_), .B(u5__abc_81276_new_n949_), .Y(u5__abc_81276_new_n950_));
AND2X2 AND2X2_4424 ( .A(u5__abc_81276_new_n400_), .B(u5__abc_81276_new_n387_), .Y(u5__abc_81276_new_n952_));
AND2X2 AND2X2_4425 ( .A(u5__abc_81276_new_n490__bF_buf3), .B(u5_state_62_), .Y(u5__abc_81276_new_n953_));
AND2X2 AND2X2_4426 ( .A(u5__abc_81276_new_n953_), .B(u5__abc_81276_new_n392_), .Y(u5__abc_81276_new_n954_));
AND2X2 AND2X2_4427 ( .A(u5__abc_81276_new_n416__bF_buf2), .B(u5__abc_81276_new_n954_), .Y(u5__abc_81276_new_n955_));
AND2X2 AND2X2_4428 ( .A(u5__abc_81276_new_n955_), .B(u5__abc_81276_new_n952_), .Y(u5__abc_81276_new_n956_));
AND2X2 AND2X2_4429 ( .A(u5__abc_81276_new_n956_), .B(u5__abc_81276_new_n448__bF_buf0), .Y(u5__abc_81276_new_n957_));
AND2X2 AND2X2_443 ( .A(u0__abc_76628_new_n1766_), .B(u0__abc_76628_new_n1173__bF_buf5), .Y(u0__abc_76628_new_n1767_));
AND2X2 AND2X2_4430 ( .A(u5__abc_81276_new_n957_), .B(u5__abc_81276_new_n523__bF_buf2), .Y(u5__abc_81276_new_n958_));
AND2X2 AND2X2_4431 ( .A(u5__abc_81276_new_n951_), .B(u5__abc_81276_new_n959_), .Y(u5__abc_81276_new_n960_));
AND2X2 AND2X2_4432 ( .A(u5__abc_81276_new_n400_), .B(u5__abc_81276_new_n391_), .Y(u5__abc_81276_new_n961_));
AND2X2 AND2X2_4433 ( .A(u5__abc_81276_new_n490__bF_buf2), .B(u5_state_61_), .Y(u5__abc_81276_new_n962_));
AND2X2 AND2X2_4434 ( .A(u5__abc_81276_new_n962_), .B(u5__abc_81276_new_n389_), .Y(u5__abc_81276_new_n963_));
AND2X2 AND2X2_4435 ( .A(u5__abc_81276_new_n416__bF_buf1), .B(u5__abc_81276_new_n963_), .Y(u5__abc_81276_new_n964_));
AND2X2 AND2X2_4436 ( .A(u5__abc_81276_new_n964_), .B(u5__abc_81276_new_n961_), .Y(u5__abc_81276_new_n965_));
AND2X2 AND2X2_4437 ( .A(u5__abc_81276_new_n965_), .B(u5__abc_81276_new_n448__bF_buf5), .Y(u5__abc_81276_new_n966_));
AND2X2 AND2X2_4438 ( .A(u5__abc_81276_new_n966_), .B(u5__abc_81276_new_n523__bF_buf1), .Y(u5__abc_81276_new_n967_));
AND2X2 AND2X2_4439 ( .A(u5__abc_81276_new_n400_), .B(u5__abc_81276_new_n390_), .Y(u5__abc_81276_new_n968_));
AND2X2 AND2X2_444 ( .A(spec_req_cs_2_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1768_));
AND2X2 AND2X2_4440 ( .A(u5__abc_81276_new_n490__bF_buf1), .B(u5_state_60_), .Y(u5__abc_81276_new_n969_));
AND2X2 AND2X2_4441 ( .A(u5__abc_81276_new_n969_), .B(u5__abc_81276_new_n389_), .Y(u5__abc_81276_new_n970_));
AND2X2 AND2X2_4442 ( .A(u5__abc_81276_new_n416__bF_buf0), .B(u5__abc_81276_new_n970_), .Y(u5__abc_81276_new_n971_));
AND2X2 AND2X2_4443 ( .A(u5__abc_81276_new_n971_), .B(u5__abc_81276_new_n968_), .Y(u5__abc_81276_new_n972_));
AND2X2 AND2X2_4444 ( .A(u5__abc_81276_new_n972_), .B(u5__abc_81276_new_n448__bF_buf4), .Y(u5__abc_81276_new_n973_));
AND2X2 AND2X2_4445 ( .A(u5__abc_81276_new_n973_), .B(u5__abc_81276_new_n523__bF_buf0), .Y(u5__abc_81276_new_n974_));
AND2X2 AND2X2_4446 ( .A(u5__abc_81276_new_n490__bF_buf0), .B(u5_state_2_), .Y(u5__abc_81276_new_n976_));
AND2X2 AND2X2_4447 ( .A(u5__abc_81276_new_n477_), .B(u5__abc_81276_new_n472_), .Y(u5__abc_81276_new_n977_));
AND2X2 AND2X2_4448 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n977_), .Y(u5__abc_81276_new_n978_));
AND2X2 AND2X2_4449 ( .A(u5__abc_81276_new_n978_), .B(u5__abc_81276_new_n976_), .Y(u5__abc_81276_new_n979_));
AND2X2 AND2X2_445 ( .A(u0__abc_76628_new_n1769_), .B(u0__abc_76628_new_n1172__bF_buf5), .Y(u0__abc_76628_new_n1770_));
AND2X2 AND2X2_4450 ( .A(u5__abc_81276_new_n979_), .B(u5__abc_81276_new_n464__bF_buf0), .Y(u5__abc_81276_new_n980_));
AND2X2 AND2X2_4451 ( .A(u5__abc_81276_new_n449__bF_buf2), .B(u5__abc_81276_new_n980_), .Y(u5__abc_81276_new_n981_));
AND2X2 AND2X2_4452 ( .A(u5__abc_81276_new_n981_), .B(u5__abc_81276_new_n522__bF_buf0), .Y(u5__abc_81276_new_n982_));
AND2X2 AND2X2_4453 ( .A(u5__abc_81276_new_n490__bF_buf10), .B(u5_state_3_), .Y(u5__abc_81276_new_n983_));
AND2X2 AND2X2_4454 ( .A(u5__abc_81276_new_n477_), .B(u5__abc_81276_new_n473_), .Y(u5__abc_81276_new_n984_));
AND2X2 AND2X2_4455 ( .A(u5__abc_81276_new_n983_), .B(u5__abc_81276_new_n984_), .Y(u5__abc_81276_new_n985_));
AND2X2 AND2X2_4456 ( .A(u5__abc_81276_new_n464__bF_buf3), .B(u5__abc_81276_new_n471_), .Y(u5__abc_81276_new_n986_));
AND2X2 AND2X2_4457 ( .A(u5__abc_81276_new_n986_), .B(u5__abc_81276_new_n985_), .Y(u5__abc_81276_new_n987_));
AND2X2 AND2X2_4458 ( .A(u5__abc_81276_new_n449__bF_buf1), .B(u5__abc_81276_new_n987_), .Y(u5__abc_81276_new_n988_));
AND2X2 AND2X2_4459 ( .A(u5__abc_81276_new_n988_), .B(u5__abc_81276_new_n522__bF_buf4), .Y(u5__abc_81276_new_n989_));
AND2X2 AND2X2_446 ( .A(spec_req_cs_1_bF_buf2_), .B(u0_tms1_24_), .Y(u0__abc_76628_new_n1771_));
AND2X2 AND2X2_4460 ( .A(u5__abc_81276_new_n488_), .B(u5_state_64_), .Y(u5__abc_81276_new_n993_));
AND2X2 AND2X2_4461 ( .A(u5__abc_81276_new_n948_), .B(u5__abc_81276_new_n993_), .Y(u5__abc_81276_new_n994_));
AND2X2 AND2X2_4462 ( .A(u5__abc_81276_new_n490__bF_buf9), .B(u5_state_63_), .Y(u5__abc_81276_new_n996_));
AND2X2 AND2X2_4463 ( .A(u5__abc_81276_new_n400_), .B(u5__abc_81276_new_n388_), .Y(u5__abc_81276_new_n997_));
AND2X2 AND2X2_4464 ( .A(u5__abc_81276_new_n997_), .B(u5__abc_81276_new_n996_), .Y(u5__abc_81276_new_n998_));
AND2X2 AND2X2_4465 ( .A(u5__abc_81276_new_n416__bF_buf3), .B(u5__abc_81276_new_n392_), .Y(u5__abc_81276_new_n999_));
AND2X2 AND2X2_4466 ( .A(u5__abc_81276_new_n999_), .B(u5__abc_81276_new_n998_), .Y(u5__abc_81276_new_n1000_));
AND2X2 AND2X2_4467 ( .A(u5__abc_81276_new_n1000_), .B(u5__abc_81276_new_n448__bF_buf3), .Y(u5__abc_81276_new_n1001_));
AND2X2 AND2X2_4468 ( .A(u5__abc_81276_new_n1001_), .B(u5__abc_81276_new_n523__bF_buf7), .Y(u5__abc_81276_new_n1002_));
AND2X2 AND2X2_4469 ( .A(u5__abc_81276_new_n995_), .B(u5__abc_81276_new_n1003_), .Y(u5__abc_81276_new_n1004_));
AND2X2 AND2X2_447 ( .A(u0__abc_76628_new_n1169__bF_buf2), .B(u0__abc_76628_new_n1774_), .Y(u0__abc_76628_new_n1775_));
AND2X2 AND2X2_4470 ( .A(u5__abc_81276_new_n992_), .B(u5__abc_81276_new_n1004_), .Y(u5__abc_81276_new_n1005_));
AND2X2 AND2X2_4471 ( .A(u5__abc_81276_new_n1005_), .B(u5__abc_81276_new_n960_), .Y(u5__abc_81276_new_n1006_));
AND2X2 AND2X2_4472 ( .A(u5__abc_81276_new_n1006_), .B(u5__abc_81276_new_n947_), .Y(u5__abc_81276_new_n1007_));
AND2X2 AND2X2_4473 ( .A(u5__abc_81276_new_n1007_), .B(u5__abc_81276_new_n874_), .Y(u5__abc_81276_new_n1008_));
AND2X2 AND2X2_4474 ( .A(u5__abc_81276_new_n1009_), .B(u5_mc_adv_r), .Y(u5__abc_81276_new_n1010_));
AND2X2 AND2X2_4475 ( .A(u5__abc_81276_new_n490__bF_buf8), .B(u5_state_11_), .Y(u5__abc_81276_new_n1011_));
AND2X2 AND2X2_4476 ( .A(u5__abc_81276_new_n462_), .B(u5__abc_81276_new_n458_), .Y(u5__abc_81276_new_n1012_));
AND2X2 AND2X2_4477 ( .A(u5__abc_81276_new_n456_), .B(u5__abc_81276_new_n1012_), .Y(u5__abc_81276_new_n1013_));
AND2X2 AND2X2_4478 ( .A(u5__abc_81276_new_n1013_), .B(u5__abc_81276_new_n1011_), .Y(u5__abc_81276_new_n1014_));
AND2X2 AND2X2_4479 ( .A(u5__abc_81276_new_n1014_), .B(u5__abc_81276_new_n479__bF_buf3), .Y(u5__abc_81276_new_n1015_));
AND2X2 AND2X2_448 ( .A(u0__abc_76628_new_n1773_), .B(u0__abc_76628_new_n1775_), .Y(u0__abc_76628_new_n1776_));
AND2X2 AND2X2_4480 ( .A(u5__abc_81276_new_n449__bF_buf0), .B(u5__abc_81276_new_n1015_), .Y(u5__abc_81276_new_n1016_));
AND2X2 AND2X2_4481 ( .A(u5__abc_81276_new_n1016_), .B(u5__abc_81276_new_n522__bF_buf3), .Y(u5__abc_81276_new_n1017_));
AND2X2 AND2X2_4482 ( .A(u5__abc_81276_new_n490__bF_buf7), .B(u5_state_36_), .Y(u5__abc_81276_new_n1019_));
AND2X2 AND2X2_4483 ( .A(u5__abc_81276_new_n1019_), .B(u5__abc_81276_new_n435_), .Y(u5__abc_81276_new_n1020_));
AND2X2 AND2X2_4484 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n1020_), .Y(u5__abc_81276_new_n1021_));
AND2X2 AND2X2_4485 ( .A(u5__abc_81276_new_n446_), .B(u5__abc_81276_new_n436_), .Y(u5__abc_81276_new_n1022_));
AND2X2 AND2X2_4486 ( .A(u5__abc_81276_new_n417__bF_buf3), .B(u5__abc_81276_new_n1022_), .Y(u5__abc_81276_new_n1023_));
AND2X2 AND2X2_4487 ( .A(u5__abc_81276_new_n523__bF_buf6), .B(u5__abc_81276_new_n1023_), .Y(u5__abc_81276_new_n1024_));
AND2X2 AND2X2_4488 ( .A(u5__abc_81276_new_n1024_), .B(u5__abc_81276_new_n1021_), .Y(u5__abc_81276_new_n1025_));
AND2X2 AND2X2_4489 ( .A(u5__abc_81276_new_n490__bF_buf6), .B(u5_state_59_), .Y(u5__abc_81276_new_n1027_));
AND2X2 AND2X2_449 ( .A(u0__abc_76628_new_n1170__bF_buf2), .B(sp_tms_25_), .Y(u0__abc_76628_new_n1778_));
AND2X2 AND2X2_4490 ( .A(u5__abc_81276_new_n399_), .B(u5__abc_81276_new_n395_), .Y(u5__abc_81276_new_n1028_));
AND2X2 AND2X2_4491 ( .A(u5__abc_81276_new_n393_), .B(u5__abc_81276_new_n1028_), .Y(u5__abc_81276_new_n1029_));
AND2X2 AND2X2_4492 ( .A(u5__abc_81276_new_n416__bF_buf2), .B(u5__abc_81276_new_n1029_), .Y(u5__abc_81276_new_n1030_));
AND2X2 AND2X2_4493 ( .A(u5__abc_81276_new_n1030_), .B(u5__abc_81276_new_n1027_), .Y(u5__abc_81276_new_n1031_));
AND2X2 AND2X2_4494 ( .A(u5__abc_81276_new_n1031_), .B(u5__abc_81276_new_n448__bF_buf2), .Y(u5__abc_81276_new_n1032_));
AND2X2 AND2X2_4495 ( .A(u5__abc_81276_new_n1032_), .B(u5__abc_81276_new_n523__bF_buf5), .Y(u5__abc_81276_new_n1033_));
AND2X2 AND2X2_4496 ( .A(u5__abc_81276_new_n490__bF_buf5), .B(u5_state_57_), .Y(u5__abc_81276_new_n1035_));
AND2X2 AND2X2_4497 ( .A(u5__abc_81276_new_n396_), .B(u5__abc_81276_new_n398_), .Y(u5__abc_81276_new_n1036_));
AND2X2 AND2X2_4498 ( .A(u5__abc_81276_new_n393_), .B(u5__abc_81276_new_n1036_), .Y(u5__abc_81276_new_n1037_));
AND2X2 AND2X2_4499 ( .A(u5__abc_81276_new_n416__bF_buf1), .B(u5__abc_81276_new_n1037_), .Y(u5__abc_81276_new_n1038_));
AND2X2 AND2X2_45 ( .A(_abc_85006_new_n371_), .B(_abc_85006_new_n372_), .Y(tms_s_27_));
AND2X2 AND2X2_450 ( .A(spec_req_cs_5_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1779_));
AND2X2 AND2X2_4500 ( .A(u5__abc_81276_new_n1038_), .B(u5__abc_81276_new_n1035_), .Y(u5__abc_81276_new_n1039_));
AND2X2 AND2X2_4501 ( .A(u5__abc_81276_new_n1039_), .B(u5__abc_81276_new_n448__bF_buf1), .Y(u5__abc_81276_new_n1040_));
AND2X2 AND2X2_4502 ( .A(u5__abc_81276_new_n1040_), .B(u5__abc_81276_new_n523__bF_buf4), .Y(u5__abc_81276_new_n1041_));
AND2X2 AND2X2_4503 ( .A(u5__abc_81276_new_n1034_), .B(u5__abc_81276_new_n1042_), .Y(u5__abc_81276_new_n1043_));
AND2X2 AND2X2_4504 ( .A(u5__abc_81276_new_n490__bF_buf4), .B(u5_state_58_), .Y(u5__abc_81276_new_n1044_));
AND2X2 AND2X2_4505 ( .A(u5__abc_81276_new_n399_), .B(u5__abc_81276_new_n394_), .Y(u5__abc_81276_new_n1045_));
AND2X2 AND2X2_4506 ( .A(u5__abc_81276_new_n393_), .B(u5__abc_81276_new_n1045_), .Y(u5__abc_81276_new_n1046_));
AND2X2 AND2X2_4507 ( .A(u5__abc_81276_new_n416__bF_buf0), .B(u5__abc_81276_new_n1046_), .Y(u5__abc_81276_new_n1047_));
AND2X2 AND2X2_4508 ( .A(u5__abc_81276_new_n1047_), .B(u5__abc_81276_new_n1044_), .Y(u5__abc_81276_new_n1048_));
AND2X2 AND2X2_4509 ( .A(u5__abc_81276_new_n1048_), .B(u5__abc_81276_new_n448__bF_buf0), .Y(u5__abc_81276_new_n1049_));
AND2X2 AND2X2_451 ( .A(u0__abc_76628_new_n1781_), .B(u0__abc_76628_new_n1179__bF_buf4), .Y(u0__abc_76628_new_n1782_));
AND2X2 AND2X2_4510 ( .A(u5__abc_81276_new_n1049_), .B(u5__abc_81276_new_n523__bF_buf3), .Y(u5__abc_81276_new_n1050_));
AND2X2 AND2X2_4511 ( .A(u5__abc_81276_new_n1043_), .B(u5__abc_81276_new_n1051_), .Y(u5__abc_81276_new_n1052_));
AND2X2 AND2X2_4512 ( .A(u5__abc_81276_new_n1052_), .B(u5__abc_81276_new_n1026_), .Y(u5__abc_81276_new_n1053_));
AND2X2 AND2X2_4513 ( .A(u5__abc_81276_new_n490__bF_buf3), .B(u5_state_56_), .Y(u5__abc_81276_new_n1054_));
AND2X2 AND2X2_4514 ( .A(u5__abc_81276_new_n396_), .B(u5__abc_81276_new_n397_), .Y(u5__abc_81276_new_n1055_));
AND2X2 AND2X2_4515 ( .A(u5__abc_81276_new_n393_), .B(u5__abc_81276_new_n1055_), .Y(u5__abc_81276_new_n1056_));
AND2X2 AND2X2_4516 ( .A(u5__abc_81276_new_n416__bF_buf3), .B(u5__abc_81276_new_n1056_), .Y(u5__abc_81276_new_n1057_));
AND2X2 AND2X2_4517 ( .A(u5__abc_81276_new_n1057_), .B(u5__abc_81276_new_n1054_), .Y(u5__abc_81276_new_n1058_));
AND2X2 AND2X2_4518 ( .A(u5__abc_81276_new_n1058_), .B(u5__abc_81276_new_n448__bF_buf5), .Y(u5__abc_81276_new_n1059_));
AND2X2 AND2X2_4519 ( .A(u5__abc_81276_new_n1059_), .B(u5__abc_81276_new_n523__bF_buf2), .Y(u5__abc_81276_new_n1060_));
AND2X2 AND2X2_452 ( .A(u0__abc_76628_new_n1782_), .B(u0__abc_76628_new_n1780_), .Y(u0__abc_76628_new_n1783_));
AND2X2 AND2X2_4520 ( .A(u5__abc_81276_new_n415_), .B(u5__abc_81276_new_n403_), .Y(u5__abc_81276_new_n1061_));
AND2X2 AND2X2_4521 ( .A(u5__abc_81276_new_n490__bF_buf2), .B(u5_state_55_), .Y(u5__abc_81276_new_n1062_));
AND2X2 AND2X2_4522 ( .A(u5__abc_81276_new_n1062_), .B(u5__abc_81276_new_n407_), .Y(u5__abc_81276_new_n1063_));
AND2X2 AND2X2_4523 ( .A(u5__abc_81276_new_n401__bF_buf2), .B(u5__abc_81276_new_n1063_), .Y(u5__abc_81276_new_n1064_));
AND2X2 AND2X2_4524 ( .A(u5__abc_81276_new_n1064_), .B(u5__abc_81276_new_n1061_), .Y(u5__abc_81276_new_n1065_));
AND2X2 AND2X2_4525 ( .A(u5__abc_81276_new_n1065_), .B(u5__abc_81276_new_n448__bF_buf4), .Y(u5__abc_81276_new_n1066_));
AND2X2 AND2X2_4526 ( .A(u5__abc_81276_new_n1066_), .B(u5__abc_81276_new_n523__bF_buf1), .Y(u5__abc_81276_new_n1067_));
AND2X2 AND2X2_4527 ( .A(u5__abc_81276_new_n415_), .B(u5__abc_81276_new_n405_), .Y(u5__abc_81276_new_n1070_));
AND2X2 AND2X2_4528 ( .A(u5__abc_81276_new_n490__bF_buf1), .B(u5_state_52_), .Y(u5__abc_81276_new_n1071_));
AND2X2 AND2X2_4529 ( .A(u5__abc_81276_new_n1071_), .B(u5__abc_81276_new_n404_), .Y(u5__abc_81276_new_n1072_));
AND2X2 AND2X2_453 ( .A(u0__abc_76628_new_n1784_), .B(u0__abc_76628_new_n1175__bF_buf4), .Y(u0__abc_76628_new_n1785_));
AND2X2 AND2X2_4530 ( .A(u5__abc_81276_new_n401__bF_buf1), .B(u5__abc_81276_new_n1072_), .Y(u5__abc_81276_new_n1073_));
AND2X2 AND2X2_4531 ( .A(u5__abc_81276_new_n1073_), .B(u5__abc_81276_new_n1070_), .Y(u5__abc_81276_new_n1074_));
AND2X2 AND2X2_4532 ( .A(u5__abc_81276_new_n1074_), .B(u5__abc_81276_new_n448__bF_buf3), .Y(u5__abc_81276_new_n1075_));
AND2X2 AND2X2_4533 ( .A(u5__abc_81276_new_n1075_), .B(u5__abc_81276_new_n523__bF_buf0), .Y(u5__abc_81276_new_n1076_));
AND2X2 AND2X2_4534 ( .A(u5__abc_81276_new_n415_), .B(u5__abc_81276_new_n406_), .Y(u5__abc_81276_new_n1078_));
AND2X2 AND2X2_4535 ( .A(u5__abc_81276_new_n490__bF_buf0), .B(u5_state_53_), .Y(u5__abc_81276_new_n1079_));
AND2X2 AND2X2_4536 ( .A(u5__abc_81276_new_n1079_), .B(u5__abc_81276_new_n404_), .Y(u5__abc_81276_new_n1080_));
AND2X2 AND2X2_4537 ( .A(u5__abc_81276_new_n401__bF_buf0), .B(u5__abc_81276_new_n1080_), .Y(u5__abc_81276_new_n1081_));
AND2X2 AND2X2_4538 ( .A(u5__abc_81276_new_n1081_), .B(u5__abc_81276_new_n1078_), .Y(u5__abc_81276_new_n1082_));
AND2X2 AND2X2_4539 ( .A(u5__abc_81276_new_n1082_), .B(u5__abc_81276_new_n448__bF_buf2), .Y(u5__abc_81276_new_n1083_));
AND2X2 AND2X2_454 ( .A(spec_req_cs_4_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1786_));
AND2X2 AND2X2_4540 ( .A(u5__abc_81276_new_n1083_), .B(u5__abc_81276_new_n523__bF_buf7), .Y(u5__abc_81276_new_n1084_));
AND2X2 AND2X2_4541 ( .A(u5__abc_81276_new_n1077_), .B(u5__abc_81276_new_n1085_), .Y(u5__abc_81276_new_n1086_));
AND2X2 AND2X2_4542 ( .A(u5__abc_81276_new_n1069_), .B(u5__abc_81276_new_n1086_), .Y(u5__abc_81276_new_n1087_));
AND2X2 AND2X2_4543 ( .A(u5__abc_81276_new_n1053_), .B(u5__abc_81276_new_n1087_), .Y(u5__abc_81276_new_n1088_));
AND2X2 AND2X2_4544 ( .A(u5__abc_81276_new_n1088_), .B(u5__abc_81276_new_n1018_), .Y(u5__abc_81276_new_n1089_));
AND2X2 AND2X2_4545 ( .A(u5__abc_81276_new_n1089_), .B(u5__abc_81276_new_n1010_), .Y(u5__abc_81276_new_n1090_));
AND2X2 AND2X2_4546 ( .A(u5__abc_81276_new_n1008_), .B(u5__abc_81276_new_n1090_), .Y(u5__abc_81276_new_n1091_));
AND2X2 AND2X2_4547 ( .A(u5__abc_81276_new_n1091_), .B(u5__abc_81276_new_n804_), .Y(u5__abc_81276_new_n1092_));
AND2X2 AND2X2_4548 ( .A(u5__abc_81276_new_n1092_), .B(u5__abc_81276_new_n671_), .Y(u5__abc_81276_new_n1093_));
AND2X2 AND2X2_4549 ( .A(u5__abc_81276_new_n1094_), .B(u5_wb_cycle), .Y(u5__abc_81276_new_n1095_));
AND2X2 AND2X2_455 ( .A(u0__abc_76628_new_n1787_), .B(u0__abc_76628_new_n1174__bF_buf4), .Y(u0__abc_76628_new_n1788_));
AND2X2 AND2X2_4550 ( .A(u5_burst_act_rd), .B(u5_cke_o_del), .Y(u5__abc_81276_new_n1096_));
AND2X2 AND2X2_4551 ( .A(u5__abc_81276_new_n1095_), .B(u5__abc_81276_new_n1096_), .Y(u5__abc_81276_new_n1097_));
AND2X2 AND2X2_4552 ( .A(u5__abc_81276_new_n1017_), .B(u5__abc_81276_new_n1097_), .Y(u5__abc_81276_new_n1098_));
AND2X2 AND2X2_4553 ( .A(u5__abc_81276_new_n1101_), .B(u5__abc_81276_new_n1102_), .Y(u5__abc_81276_new_n1103_));
AND2X2 AND2X2_4554 ( .A(u5__abc_81276_new_n1104_), .B(u5__abc_81276_new_n1105_), .Y(u5__abc_81276_new_n1106_));
AND2X2 AND2X2_4555 ( .A(u5__abc_81276_new_n1103_), .B(u5__abc_81276_new_n1106_), .Y(u5__abc_81276_new_n1107_));
AND2X2 AND2X2_4556 ( .A(u5__abc_81276_new_n1108_), .B(u5__abc_81276_new_n1109_), .Y(u5__abc_81276_new_n1110_));
AND2X2 AND2X2_4557 ( .A(u5__abc_81276_new_n1111_), .B(u5__abc_81276_new_n1112_), .Y(u5__abc_81276_new_n1113_));
AND2X2 AND2X2_4558 ( .A(u5__abc_81276_new_n1110_), .B(u5__abc_81276_new_n1113_), .Y(u5__abc_81276_new_n1114_));
AND2X2 AND2X2_4559 ( .A(u5__abc_81276_new_n1107_), .B(u5__abc_81276_new_n1114_), .Y(u5_timer_is_zero));
AND2X2 AND2X2_456 ( .A(spec_req_cs_3_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1789_));
AND2X2 AND2X2_4560 ( .A(u5__abc_81276_new_n1116_), .B(u5__abc_81276_new_n1117_), .Y(u5__abc_81276_new_n1118_));
AND2X2 AND2X2_4561 ( .A(u5__abc_81276_new_n1119_), .B(u5__abc_81276_new_n1120_), .Y(u5__abc_81276_new_n1121_));
AND2X2 AND2X2_4562 ( .A(u5__abc_81276_new_n1118_), .B(u5__abc_81276_new_n1121_), .Y(u5__0ir_cnt_done_0_0_));
AND2X2 AND2X2_4563 ( .A(u5__abc_81276_new_n1123_), .B(u5__abc_81276_new_n1124_), .Y(u5__0no_wb_cycle_0_0_));
AND2X2 AND2X2_4564 ( .A(u5__abc_81276_new_n523__bF_buf6), .B(u5__abc_81276_new_n490__bF_buf10), .Y(u5__abc_81276_new_n1126_));
AND2X2 AND2X2_4565 ( .A(u5__abc_81276_new_n387_), .B(u5_state_62_), .Y(u5__abc_81276_new_n1127_));
AND2X2 AND2X2_4566 ( .A(u5__abc_81276_new_n392_), .B(u5__abc_81276_new_n1127_), .Y(u5__abc_81276_new_n1128_));
AND2X2 AND2X2_4567 ( .A(u5__abc_81276_new_n400_), .B(u5__abc_81276_new_n1128_), .Y(u5__abc_81276_new_n1129_));
AND2X2 AND2X2_4568 ( .A(u5__abc_81276_new_n416__bF_buf2), .B(u5__abc_81276_new_n1129_), .Y(u5__abc_81276_new_n1130_));
AND2X2 AND2X2_4569 ( .A(u5__abc_81276_new_n448__bF_buf1), .B(u5__abc_81276_new_n1130_), .Y(u5__abc_81276_new_n1131_));
AND2X2 AND2X2_457 ( .A(u0__abc_76628_new_n1790_), .B(u0__abc_76628_new_n1173__bF_buf4), .Y(u0__abc_76628_new_n1791_));
AND2X2 AND2X2_4570 ( .A(u5__abc_81276_new_n1126__bF_buf3), .B(u5__abc_81276_new_n1131_), .Y(u5__abc_81276_new_n1132_));
AND2X2 AND2X2_4571 ( .A(u5__abc_81276_new_n951_), .B(u5__abc_81276_new_n1133_), .Y(u5__abc_81276_new_n1134_));
AND2X2 AND2X2_4572 ( .A(u5__abc_81276_new_n416__bF_buf1), .B(u5__abc_81276_new_n389_), .Y(u5__abc_81276_new_n1135_));
AND2X2 AND2X2_4573 ( .A(u5__abc_81276_new_n448__bF_buf0), .B(u5__abc_81276_new_n1135_), .Y(u5__abc_81276_new_n1136_));
AND2X2 AND2X2_4574 ( .A(u5__abc_81276_new_n523__bF_buf5), .B(u5__abc_81276_new_n1136_), .Y(u5__abc_81276_new_n1137_));
AND2X2 AND2X2_4575 ( .A(u5__abc_81276_new_n391_), .B(u5_state_61_), .Y(u5__abc_81276_new_n1138_));
AND2X2 AND2X2_4576 ( .A(u5__abc_81276_new_n490__bF_buf9), .B(u5__abc_81276_new_n1138_), .Y(u5__abc_81276_new_n1139_));
AND2X2 AND2X2_4577 ( .A(u5__abc_81276_new_n400_), .B(u5__abc_81276_new_n1139_), .Y(u5__abc_81276_new_n1140_));
AND2X2 AND2X2_4578 ( .A(u5__abc_81276_new_n1137_), .B(u5__abc_81276_new_n1140_), .Y(u5__abc_81276_new_n1141_));
AND2X2 AND2X2_4579 ( .A(u5__abc_81276_new_n390_), .B(u5_state_60_), .Y(u5__abc_81276_new_n1143_));
AND2X2 AND2X2_458 ( .A(spec_req_cs_2_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1792_));
AND2X2 AND2X2_4580 ( .A(u5__abc_81276_new_n490__bF_buf8), .B(u5__abc_81276_new_n1143_), .Y(u5__abc_81276_new_n1144_));
AND2X2 AND2X2_4581 ( .A(u5__abc_81276_new_n400_), .B(u5__abc_81276_new_n1144_), .Y(u5__abc_81276_new_n1145_));
AND2X2 AND2X2_4582 ( .A(u5__abc_81276_new_n1137_), .B(u5__abc_81276_new_n1145_), .Y(u5__abc_81276_new_n1146_));
AND2X2 AND2X2_4583 ( .A(u5__abc_81276_new_n1142_), .B(u5__abc_81276_new_n1147_), .Y(u5__abc_81276_new_n1148_));
AND2X2 AND2X2_4584 ( .A(u5__abc_81276_new_n449__bF_buf7), .B(u5__abc_81276_new_n522__bF_buf2), .Y(u5__abc_81276_new_n1149_));
AND2X2 AND2X2_4585 ( .A(u5__abc_81276_new_n477_), .B(u5__abc_81276_new_n490__bF_buf7), .Y(u5__abc_81276_new_n1150_));
AND2X2 AND2X2_4586 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n1150_), .Y(u5__abc_81276_new_n1151_));
AND2X2 AND2X2_4587 ( .A(u5__abc_81276_new_n472_), .B(u5_state_2_), .Y(u5__abc_81276_new_n1152_));
AND2X2 AND2X2_4588 ( .A(u5__abc_81276_new_n464__bF_buf2), .B(u5__abc_81276_new_n1152_), .Y(u5__abc_81276_new_n1153_));
AND2X2 AND2X2_4589 ( .A(u5__abc_81276_new_n1153_), .B(u5__abc_81276_new_n1151_), .Y(u5__abc_81276_new_n1154_));
AND2X2 AND2X2_459 ( .A(u0__abc_76628_new_n1793_), .B(u0__abc_76628_new_n1172__bF_buf4), .Y(u0__abc_76628_new_n1794_));
AND2X2 AND2X2_4590 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1154_), .Y(u5__abc_81276_new_n1155_));
AND2X2 AND2X2_4591 ( .A(u5__abc_81276_new_n473_), .B(u5_state_3_), .Y(u5__abc_81276_new_n1157_));
AND2X2 AND2X2_4592 ( .A(u5__abc_81276_new_n464__bF_buf1), .B(u5__abc_81276_new_n1157_), .Y(u5__abc_81276_new_n1158_));
AND2X2 AND2X2_4593 ( .A(u5__abc_81276_new_n1158_), .B(u5__abc_81276_new_n1151_), .Y(u5__abc_81276_new_n1159_));
AND2X2 AND2X2_4594 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1159_), .Y(u5__abc_81276_new_n1160_));
AND2X2 AND2X2_4595 ( .A(u5__abc_81276_new_n1156_), .B(u5__abc_81276_new_n1161_), .Y(u5__abc_81276_new_n1162_));
AND2X2 AND2X2_4596 ( .A(u5__abc_81276_new_n1148_), .B(u5__abc_81276_new_n1162_), .Y(u5__abc_81276_new_n1163_));
AND2X2 AND2X2_4597 ( .A(u5__abc_81276_new_n388_), .B(u5_state_63_), .Y(u5__abc_81276_new_n1164_));
AND2X2 AND2X2_4598 ( .A(u5__abc_81276_new_n490__bF_buf6), .B(u5__abc_81276_new_n1164_), .Y(u5__abc_81276_new_n1165_));
AND2X2 AND2X2_4599 ( .A(u5__abc_81276_new_n1165_), .B(u5__abc_81276_new_n392_), .Y(u5__abc_81276_new_n1166_));
AND2X2 AND2X2_46 ( .A(_abc_85006_new_n389_), .B(_abc_85006_new_n390_), .Y(csc_s_1_));
AND2X2 AND2X2_460 ( .A(spec_req_cs_1_bF_buf1_), .B(u0_tms1_25_), .Y(u0__abc_76628_new_n1795_));
AND2X2 AND2X2_4600 ( .A(u5__abc_81276_new_n1166_), .B(u5__abc_81276_new_n400_), .Y(u5__abc_81276_new_n1167_));
AND2X2 AND2X2_4601 ( .A(u5__abc_81276_new_n1167_), .B(u5__abc_81276_new_n416__bF_buf0), .Y(u5__abc_81276_new_n1168_));
AND2X2 AND2X2_4602 ( .A(u5__abc_81276_new_n1168_), .B(u5__abc_81276_new_n448__bF_buf5), .Y(u5__abc_81276_new_n1169_));
AND2X2 AND2X2_4603 ( .A(u5__abc_81276_new_n1169_), .B(u5__abc_81276_new_n523__bF_buf4), .Y(u5__abc_81276_new_n1170_));
AND2X2 AND2X2_4604 ( .A(u5__abc_81276_new_n995_), .B(u5__abc_81276_new_n1171_), .Y(u5__abc_81276_new_n1172_));
AND2X2 AND2X2_4605 ( .A(u5__abc_81276_new_n1163_), .B(u5__abc_81276_new_n1172_), .Y(u5__abc_81276_new_n1173_));
AND2X2 AND2X2_4606 ( .A(u5__abc_81276_new_n1173_), .B(u5__abc_81276_new_n1134_), .Y(u5__abc_81276_new_n1174_));
AND2X2 AND2X2_4607 ( .A(u5__abc_81276_new_n448__bF_buf4), .B(u5__abc_81276_new_n393_), .Y(u5__abc_81276_new_n1175_));
AND2X2 AND2X2_4608 ( .A(u5__abc_81276_new_n523__bF_buf3), .B(u5__abc_81276_new_n1175_), .Y(u5__abc_81276_new_n1176_));
AND2X2 AND2X2_4609 ( .A(u5__abc_81276_new_n397_), .B(u5_state_56_), .Y(u5__abc_81276_new_n1177_));
AND2X2 AND2X2_461 ( .A(u0__abc_76628_new_n1169__bF_buf1), .B(u0__abc_76628_new_n1798_), .Y(u0__abc_76628_new_n1799_));
AND2X2 AND2X2_4610 ( .A(u5__abc_81276_new_n490__bF_buf5), .B(u5__abc_81276_new_n1177_), .Y(u5__abc_81276_new_n1178_));
AND2X2 AND2X2_4611 ( .A(u5__abc_81276_new_n1178_), .B(u5__abc_81276_new_n396_), .Y(u5__abc_81276_new_n1179_));
AND2X2 AND2X2_4612 ( .A(u5__abc_81276_new_n416__bF_buf3), .B(u5__abc_81276_new_n1179_), .Y(u5__abc_81276_new_n1180_));
AND2X2 AND2X2_4613 ( .A(u5__abc_81276_new_n1176_), .B(u5__abc_81276_new_n1180_), .Y(u5__abc_81276_new_n1181_));
AND2X2 AND2X2_4614 ( .A(u5__abc_81276_new_n448__bF_buf3), .B(u5__abc_81276_new_n401__bF_buf3), .Y(u5__abc_81276_new_n1184_));
AND2X2 AND2X2_4615 ( .A(u5__abc_81276_new_n1193_), .B(u5__abc_81276_new_n1182_), .Y(u5__abc_81276_new_n1194_));
AND2X2 AND2X2_4616 ( .A(u5__abc_81276_new_n523__bF_buf1), .B(u5__abc_81276_new_n1184_), .Y(u5__abc_81276_new_n1195_));
AND2X2 AND2X2_4617 ( .A(u5__abc_81276_new_n405_), .B(u5_state_52_), .Y(u5__abc_81276_new_n1196_));
AND2X2 AND2X2_4618 ( .A(u5__abc_81276_new_n490__bF_buf4), .B(u5__abc_81276_new_n1196_), .Y(u5__abc_81276_new_n1197_));
AND2X2 AND2X2_4619 ( .A(u5__abc_81276_new_n1197_), .B(u5__abc_81276_new_n404_), .Y(u5__abc_81276_new_n1198_));
AND2X2 AND2X2_462 ( .A(u0__abc_76628_new_n1797_), .B(u0__abc_76628_new_n1799_), .Y(u0__abc_76628_new_n1800_));
AND2X2 AND2X2_4620 ( .A(u5__abc_81276_new_n1198_), .B(u5__abc_81276_new_n415_), .Y(u5__abc_81276_new_n1199_));
AND2X2 AND2X2_4621 ( .A(u5__abc_81276_new_n1195_), .B(u5__abc_81276_new_n1199_), .Y(u5__abc_81276_new_n1200_));
AND2X2 AND2X2_4622 ( .A(u5__abc_81276_new_n406_), .B(u5_state_53_), .Y(u5__abc_81276_new_n1202_));
AND2X2 AND2X2_4623 ( .A(u5__abc_81276_new_n490__bF_buf3), .B(u5__abc_81276_new_n1202_), .Y(u5__abc_81276_new_n1203_));
AND2X2 AND2X2_4624 ( .A(u5__abc_81276_new_n1203_), .B(u5__abc_81276_new_n404_), .Y(u5__abc_81276_new_n1204_));
AND2X2 AND2X2_4625 ( .A(u5__abc_81276_new_n1204_), .B(u5__abc_81276_new_n415_), .Y(u5__abc_81276_new_n1205_));
AND2X2 AND2X2_4626 ( .A(u5__abc_81276_new_n1195_), .B(u5__abc_81276_new_n1205_), .Y(u5__abc_81276_new_n1206_));
AND2X2 AND2X2_4627 ( .A(u5__abc_81276_new_n1201_), .B(u5__abc_81276_new_n1207_), .Y(u5__abc_81276_new_n1208_));
AND2X2 AND2X2_4628 ( .A(u5__abc_81276_new_n1194_), .B(u5__abc_81276_new_n1208_), .Y(u5__abc_81276_new_n1209_));
AND2X2 AND2X2_4629 ( .A(u5__abc_81276_new_n416__bF_buf2), .B(u5__abc_81276_new_n393_), .Y(u5__abc_81276_new_n1210_));
AND2X2 AND2X2_463 ( .A(u0__abc_76628_new_n1170__bF_buf1), .B(sp_tms_26_), .Y(u0__abc_76628_new_n1802_));
AND2X2 AND2X2_4630 ( .A(u5__abc_81276_new_n395_), .B(u5_state_59_), .Y(u5__abc_81276_new_n1211_));
AND2X2 AND2X2_4631 ( .A(u5__abc_81276_new_n399_), .B(u5__abc_81276_new_n1211_), .Y(u5__abc_81276_new_n1212_));
AND2X2 AND2X2_4632 ( .A(u5__abc_81276_new_n448__bF_buf2), .B(u5__abc_81276_new_n1212_), .Y(u5__abc_81276_new_n1213_));
AND2X2 AND2X2_4633 ( .A(u5__abc_81276_new_n1213_), .B(u5__abc_81276_new_n1210_), .Y(u5__abc_81276_new_n1214_));
AND2X2 AND2X2_4634 ( .A(u5__abc_81276_new_n1126__bF_buf2), .B(u5__abc_81276_new_n1214_), .Y(u5__abc_81276_new_n1215_));
AND2X2 AND2X2_4635 ( .A(u5__abc_81276_new_n1225_), .B(u5__abc_81276_new_n1216_), .Y(u5__abc_81276_new_n1226_));
AND2X2 AND2X2_4636 ( .A(u5__abc_81276_new_n398_), .B(u5_state_57_), .Y(u5__abc_81276_new_n1227_));
AND2X2 AND2X2_4637 ( .A(u5__abc_81276_new_n490__bF_buf2), .B(u5__abc_81276_new_n1227_), .Y(u5__abc_81276_new_n1228_));
AND2X2 AND2X2_4638 ( .A(u5__abc_81276_new_n1228_), .B(u5__abc_81276_new_n396_), .Y(u5__abc_81276_new_n1229_));
AND2X2 AND2X2_4639 ( .A(u5__abc_81276_new_n416__bF_buf1), .B(u5__abc_81276_new_n1229_), .Y(u5__abc_81276_new_n1230_));
AND2X2 AND2X2_464 ( .A(spec_req_cs_5_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1803_));
AND2X2 AND2X2_4640 ( .A(u5__abc_81276_new_n1176_), .B(u5__abc_81276_new_n1230_), .Y(u5__abc_81276_new_n1231_));
AND2X2 AND2X2_4641 ( .A(u5__abc_81276_new_n402_), .B(u5_state_54_), .Y(u5__abc_81276_new_n1233_));
AND2X2 AND2X2_4642 ( .A(u5__abc_81276_new_n490__bF_buf1), .B(u5__abc_81276_new_n1233_), .Y(u5__abc_81276_new_n1234_));
AND2X2 AND2X2_4643 ( .A(u5__abc_81276_new_n1234_), .B(u5__abc_81276_new_n407_), .Y(u5__abc_81276_new_n1235_));
AND2X2 AND2X2_4644 ( .A(u5__abc_81276_new_n1235_), .B(u5__abc_81276_new_n415_), .Y(u5__abc_81276_new_n1236_));
AND2X2 AND2X2_4645 ( .A(u5__abc_81276_new_n1195_), .B(u5__abc_81276_new_n1236_), .Y(u5__abc_81276_new_n1237_));
AND2X2 AND2X2_4646 ( .A(u5__abc_81276_new_n1232_), .B(u5__abc_81276_new_n1238_), .Y(u5__abc_81276_new_n1239_));
AND2X2 AND2X2_4647 ( .A(u5__abc_81276_new_n1226_), .B(u5__abc_81276_new_n1239_), .Y(u5__abc_81276_new_n1240_));
AND2X2 AND2X2_4648 ( .A(u5__abc_81276_new_n1240_), .B(u5__abc_81276_new_n1209_), .Y(u5__abc_81276_new_n1241_));
AND2X2 AND2X2_4649 ( .A(u5__abc_81276_new_n1174_), .B(u5__abc_81276_new_n1241_), .Y(u5__abc_81276_new_n1242_));
AND2X2 AND2X2_465 ( .A(u0__abc_76628_new_n1805_), .B(u0__abc_76628_new_n1179__bF_buf3), .Y(u0__abc_76628_new_n1806_));
AND2X2 AND2X2_4650 ( .A(u5__abc_81276_new_n434_), .B(u5_state_39_), .Y(u5__abc_81276_new_n1243_));
AND2X2 AND2X2_4651 ( .A(u5__abc_81276_new_n438_), .B(u5__abc_81276_new_n1243_), .Y(u5__abc_81276_new_n1244_));
AND2X2 AND2X2_4652 ( .A(u5__abc_81276_new_n446_), .B(u5__abc_81276_new_n1244_), .Y(u5__abc_81276_new_n1245_));
AND2X2 AND2X2_4653 ( .A(u5__abc_81276_new_n557_), .B(u5__abc_81276_new_n1245_), .Y(u5__abc_81276_new_n1246_));
AND2X2 AND2X2_4654 ( .A(u5__abc_81276_new_n1126__bF_buf1), .B(u5__abc_81276_new_n1246_), .Y(u5__abc_81276_new_n1247_));
AND2X2 AND2X2_4655 ( .A(u5__abc_81276_new_n433_), .B(u5_state_38_), .Y(u5__abc_81276_new_n1249_));
AND2X2 AND2X2_4656 ( .A(u5__abc_81276_new_n438_), .B(u5__abc_81276_new_n1249_), .Y(u5__abc_81276_new_n1250_));
AND2X2 AND2X2_4657 ( .A(u5__abc_81276_new_n446_), .B(u5__abc_81276_new_n1250_), .Y(u5__abc_81276_new_n1251_));
AND2X2 AND2X2_4658 ( .A(u5__abc_81276_new_n557_), .B(u5__abc_81276_new_n1251_), .Y(u5__abc_81276_new_n1252_));
AND2X2 AND2X2_4659 ( .A(u5__abc_81276_new_n1126__bF_buf0), .B(u5__abc_81276_new_n1252_), .Y(u5__abc_81276_new_n1253_));
AND2X2 AND2X2_466 ( .A(u0__abc_76628_new_n1806_), .B(u0__abc_76628_new_n1804_), .Y(u0__abc_76628_new_n1807_));
AND2X2 AND2X2_4660 ( .A(u5__abc_81276_new_n1248_), .B(u5__abc_81276_new_n1254_), .Y(u5__abc_81276_new_n1255_));
AND2X2 AND2X2_4661 ( .A(u5__abc_81276_new_n429_), .B(u5_state_40_), .Y(u5__abc_81276_new_n1256_));
AND2X2 AND2X2_4662 ( .A(u5__abc_81276_new_n427_), .B(u5__abc_81276_new_n1256_), .Y(u5__abc_81276_new_n1257_));
AND2X2 AND2X2_4663 ( .A(u5__abc_81276_new_n424_), .B(u5__abc_81276_new_n1257_), .Y(u5__abc_81276_new_n1258_));
AND2X2 AND2X2_4664 ( .A(u5__abc_81276_new_n706_), .B(u5__abc_81276_new_n1258_), .Y(u5__abc_81276_new_n1259_));
AND2X2 AND2X2_4665 ( .A(u5__abc_81276_new_n1126__bF_buf3), .B(u5__abc_81276_new_n1259_), .Y(u5__abc_81276_new_n1260_));
AND2X2 AND2X2_4666 ( .A(u5__abc_81276_new_n419_), .B(u5_state_47_), .Y(u5__abc_81276_new_n1262_));
AND2X2 AND2X2_4667 ( .A(u5__abc_81276_new_n423_), .B(u5__abc_81276_new_n1262_), .Y(u5__abc_81276_new_n1263_));
AND2X2 AND2X2_4668 ( .A(u5__abc_81276_new_n431_), .B(u5__abc_81276_new_n1263_), .Y(u5__abc_81276_new_n1264_));
AND2X2 AND2X2_4669 ( .A(u5__abc_81276_new_n706_), .B(u5__abc_81276_new_n1264_), .Y(u5__abc_81276_new_n1265_));
AND2X2 AND2X2_467 ( .A(u0__abc_76628_new_n1808_), .B(u0__abc_76628_new_n1175__bF_buf3), .Y(u0__abc_76628_new_n1809_));
AND2X2 AND2X2_4670 ( .A(u5__abc_81276_new_n1126__bF_buf2), .B(u5__abc_81276_new_n1265_), .Y(u5__abc_81276_new_n1266_));
AND2X2 AND2X2_4671 ( .A(u5__abc_81276_new_n1261_), .B(u5__abc_81276_new_n1267_), .Y(u5__abc_81276_new_n1268_));
AND2X2 AND2X2_4672 ( .A(u5__abc_81276_new_n1255_), .B(u5__abc_81276_new_n1268_), .Y(u5__abc_81276_new_n1269_));
AND2X2 AND2X2_4673 ( .A(u5__abc_81276_new_n1195_), .B(u5__abc_81276_new_n682_), .Y(u5__abc_81276_new_n1270_));
AND2X2 AND2X2_4674 ( .A(u5__abc_81276_new_n1195_), .B(u5__abc_81276_new_n675_), .Y(u5__abc_81276_new_n1272_));
AND2X2 AND2X2_4675 ( .A(u5__abc_81276_new_n1271_), .B(u5__abc_81276_new_n1273_), .Y(u5__abc_81276_new_n1274_));
AND2X2 AND2X2_4676 ( .A(u5__abc_81276_new_n448__bF_buf0), .B(u5__abc_81276_new_n408_), .Y(u5__abc_81276_new_n1275_));
AND2X2 AND2X2_4677 ( .A(u5__abc_81276_new_n523__bF_buf0), .B(u5__abc_81276_new_n1275_), .Y(u5__abc_81276_new_n1276_));
AND2X2 AND2X2_4678 ( .A(u5__abc_81276_new_n413_), .B(u5_state_49_), .Y(u5__abc_81276_new_n1277_));
AND2X2 AND2X2_4679 ( .A(u5__abc_81276_new_n490__bF_buf0), .B(u5__abc_81276_new_n1277_), .Y(u5__abc_81276_new_n1278_));
AND2X2 AND2X2_468 ( .A(spec_req_cs_4_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1810_));
AND2X2 AND2X2_4680 ( .A(u5__abc_81276_new_n1278_), .B(u5__abc_81276_new_n411_), .Y(u5__abc_81276_new_n1279_));
AND2X2 AND2X2_4681 ( .A(u5__abc_81276_new_n401__bF_buf2), .B(u5__abc_81276_new_n1279_), .Y(u5__abc_81276_new_n1280_));
AND2X2 AND2X2_4682 ( .A(u5__abc_81276_new_n1276_), .B(u5__abc_81276_new_n1280_), .Y(u5__abc_81276_new_n1281_));
AND2X2 AND2X2_4683 ( .A(u5__abc_81276_new_n412_), .B(u5_state_48_), .Y(u5__abc_81276_new_n1283_));
AND2X2 AND2X2_4684 ( .A(u5__abc_81276_new_n490__bF_buf10), .B(u5__abc_81276_new_n1283_), .Y(u5__abc_81276_new_n1284_));
AND2X2 AND2X2_4685 ( .A(u5__abc_81276_new_n1284_), .B(u5__abc_81276_new_n411_), .Y(u5__abc_81276_new_n1285_));
AND2X2 AND2X2_4686 ( .A(u5__abc_81276_new_n401__bF_buf1), .B(u5__abc_81276_new_n1285_), .Y(u5__abc_81276_new_n1286_));
AND2X2 AND2X2_4687 ( .A(u5__abc_81276_new_n1276_), .B(u5__abc_81276_new_n1286_), .Y(u5__abc_81276_new_n1287_));
AND2X2 AND2X2_4688 ( .A(u5__abc_81276_new_n1282_), .B(u5__abc_81276_new_n1288_), .Y(u5__abc_81276_new_n1289_));
AND2X2 AND2X2_4689 ( .A(u5__abc_81276_new_n1274_), .B(u5__abc_81276_new_n1289_), .Y(u5__abc_81276_new_n1290_));
AND2X2 AND2X2_469 ( .A(u0__abc_76628_new_n1811_), .B(u0__abc_76628_new_n1174__bF_buf3), .Y(u0__abc_76628_new_n1812_));
AND2X2 AND2X2_4690 ( .A(u5__abc_81276_new_n1269_), .B(u5__abc_81276_new_n1290_), .Y(u5__abc_81276_new_n1291_));
AND2X2 AND2X2_4691 ( .A(u5__abc_81276_new_n421_), .B(u5_state_44_), .Y(u5__abc_81276_new_n1292_));
AND2X2 AND2X2_4692 ( .A(u5__abc_81276_new_n420_), .B(u5__abc_81276_new_n1292_), .Y(u5__abc_81276_new_n1293_));
AND2X2 AND2X2_4693 ( .A(u5__abc_81276_new_n431_), .B(u5__abc_81276_new_n1293_), .Y(u5__abc_81276_new_n1294_));
AND2X2 AND2X2_4694 ( .A(u5__abc_81276_new_n706_), .B(u5__abc_81276_new_n1294_), .Y(u5__abc_81276_new_n1295_));
AND2X2 AND2X2_4695 ( .A(u5__abc_81276_new_n1126__bF_buf1), .B(u5__abc_81276_new_n1295_), .Y(u5__abc_81276_new_n1296_));
AND2X2 AND2X2_4696 ( .A(u5__abc_81276_new_n426_), .B(u5_state_43_), .Y(u5__abc_81276_new_n1298_));
AND2X2 AND2X2_4697 ( .A(u5__abc_81276_new_n430_), .B(u5__abc_81276_new_n1298_), .Y(u5__abc_81276_new_n1299_));
AND2X2 AND2X2_4698 ( .A(u5__abc_81276_new_n424_), .B(u5__abc_81276_new_n1299_), .Y(u5__abc_81276_new_n1300_));
AND2X2 AND2X2_4699 ( .A(u5__abc_81276_new_n706_), .B(u5__abc_81276_new_n1300_), .Y(u5__abc_81276_new_n1301_));
AND2X2 AND2X2_47 ( .A(_abc_85006_new_n392_), .B(_abc_85006_new_n393_), .Y(csc_s_2_));
AND2X2 AND2X2_470 ( .A(spec_req_cs_3_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1813_));
AND2X2 AND2X2_4700 ( .A(u5__abc_81276_new_n1126__bF_buf0), .B(u5__abc_81276_new_n1301_), .Y(u5__abc_81276_new_n1302_));
AND2X2 AND2X2_4701 ( .A(u5__abc_81276_new_n1297_), .B(u5__abc_81276_new_n1303_), .Y(u5__abc_81276_new_n1304_));
AND2X2 AND2X2_4702 ( .A(u5__abc_81276_new_n418_), .B(u5_state_46_), .Y(u5__abc_81276_new_n1305_));
AND2X2 AND2X2_4703 ( .A(u5__abc_81276_new_n423_), .B(u5__abc_81276_new_n1305_), .Y(u5__abc_81276_new_n1306_));
AND2X2 AND2X2_4704 ( .A(u5__abc_81276_new_n431_), .B(u5__abc_81276_new_n1306_), .Y(u5__abc_81276_new_n1307_));
AND2X2 AND2X2_4705 ( .A(u5__abc_81276_new_n706_), .B(u5__abc_81276_new_n1307_), .Y(u5__abc_81276_new_n1308_));
AND2X2 AND2X2_4706 ( .A(u5__abc_81276_new_n1126__bF_buf3), .B(u5__abc_81276_new_n1308_), .Y(u5__abc_81276_new_n1309_));
AND2X2 AND2X2_4707 ( .A(u5__abc_81276_new_n422_), .B(u5_state_45_), .Y(u5__abc_81276_new_n1311_));
AND2X2 AND2X2_4708 ( .A(u5__abc_81276_new_n420_), .B(u5__abc_81276_new_n1311_), .Y(u5__abc_81276_new_n1312_));
AND2X2 AND2X2_4709 ( .A(u5__abc_81276_new_n431_), .B(u5__abc_81276_new_n1312_), .Y(u5__abc_81276_new_n1313_));
AND2X2 AND2X2_471 ( .A(u0__abc_76628_new_n1814_), .B(u0__abc_76628_new_n1173__bF_buf3), .Y(u0__abc_76628_new_n1815_));
AND2X2 AND2X2_4710 ( .A(u5__abc_81276_new_n706_), .B(u5__abc_81276_new_n1313_), .Y(u5__abc_81276_new_n1314_));
AND2X2 AND2X2_4711 ( .A(u5__abc_81276_new_n1126__bF_buf2), .B(u5__abc_81276_new_n1314_), .Y(u5__abc_81276_new_n1315_));
AND2X2 AND2X2_4712 ( .A(u5__abc_81276_new_n1310_), .B(u5__abc_81276_new_n1316_), .Y(u5__abc_81276_new_n1317_));
AND2X2 AND2X2_4713 ( .A(u5__abc_81276_new_n1304_), .B(u5__abc_81276_new_n1317_), .Y(u5__abc_81276_new_n1318_));
AND2X2 AND2X2_4714 ( .A(u5__abc_81276_new_n425_), .B(u5_state_42_), .Y(u5__abc_81276_new_n1319_));
AND2X2 AND2X2_4715 ( .A(u5__abc_81276_new_n430_), .B(u5__abc_81276_new_n1319_), .Y(u5__abc_81276_new_n1320_));
AND2X2 AND2X2_4716 ( .A(u5__abc_81276_new_n424_), .B(u5__abc_81276_new_n1320_), .Y(u5__abc_81276_new_n1321_));
AND2X2 AND2X2_4717 ( .A(u5__abc_81276_new_n706_), .B(u5__abc_81276_new_n1321_), .Y(u5__abc_81276_new_n1322_));
AND2X2 AND2X2_4718 ( .A(u5__abc_81276_new_n1126__bF_buf1), .B(u5__abc_81276_new_n1322_), .Y(u5__abc_81276_new_n1323_));
AND2X2 AND2X2_4719 ( .A(u5__abc_81276_new_n428_), .B(u5_state_41_), .Y(u5__abc_81276_new_n1325_));
AND2X2 AND2X2_472 ( .A(spec_req_cs_2_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1816_));
AND2X2 AND2X2_4720 ( .A(u5__abc_81276_new_n427_), .B(u5__abc_81276_new_n1325_), .Y(u5__abc_81276_new_n1326_));
AND2X2 AND2X2_4721 ( .A(u5__abc_81276_new_n424_), .B(u5__abc_81276_new_n1326_), .Y(u5__abc_81276_new_n1327_));
AND2X2 AND2X2_4722 ( .A(u5__abc_81276_new_n706_), .B(u5__abc_81276_new_n1327_), .Y(u5__abc_81276_new_n1328_));
AND2X2 AND2X2_4723 ( .A(u5__abc_81276_new_n1126__bF_buf0), .B(u5__abc_81276_new_n1328_), .Y(u5__abc_81276_new_n1329_));
AND2X2 AND2X2_4724 ( .A(u5__abc_81276_new_n1324_), .B(u5__abc_81276_new_n1330_), .Y(u5__abc_81276_new_n1331_));
AND2X2 AND2X2_4725 ( .A(u5__abc_81276_new_n437_), .B(u5_state_37_), .Y(u5__abc_81276_new_n1332_));
AND2X2 AND2X2_4726 ( .A(u5__abc_81276_new_n435_), .B(u5__abc_81276_new_n1332_), .Y(u5__abc_81276_new_n1333_));
AND2X2 AND2X2_4727 ( .A(u5__abc_81276_new_n446_), .B(u5__abc_81276_new_n1333_), .Y(u5__abc_81276_new_n1334_));
AND2X2 AND2X2_4728 ( .A(u5__abc_81276_new_n557_), .B(u5__abc_81276_new_n1334_), .Y(u5__abc_81276_new_n1335_));
AND2X2 AND2X2_4729 ( .A(u5__abc_81276_new_n1126__bF_buf3), .B(u5__abc_81276_new_n1335_), .Y(u5__abc_81276_new_n1336_));
AND2X2 AND2X2_473 ( .A(u0__abc_76628_new_n1817_), .B(u0__abc_76628_new_n1172__bF_buf3), .Y(u0__abc_76628_new_n1818_));
AND2X2 AND2X2_4730 ( .A(u5__abc_81276_new_n436_), .B(u5_state_36_), .Y(u5__abc_81276_new_n1338_));
AND2X2 AND2X2_4731 ( .A(u5__abc_81276_new_n435_), .B(u5__abc_81276_new_n1338_), .Y(u5__abc_81276_new_n1339_));
AND2X2 AND2X2_4732 ( .A(u5__abc_81276_new_n446_), .B(u5__abc_81276_new_n1339_), .Y(u5__abc_81276_new_n1340_));
AND2X2 AND2X2_4733 ( .A(u5__abc_81276_new_n557_), .B(u5__abc_81276_new_n1340_), .Y(u5__abc_81276_new_n1341_));
AND2X2 AND2X2_4734 ( .A(u5__abc_81276_new_n1126__bF_buf2), .B(u5__abc_81276_new_n1341_), .Y(u5__abc_81276_new_n1342_));
AND2X2 AND2X2_4735 ( .A(u5__abc_81276_new_n1337_), .B(u5__abc_81276_new_n1343_), .Y(u5__abc_81276_new_n1344_));
AND2X2 AND2X2_4736 ( .A(u5__abc_81276_new_n1331_), .B(u5__abc_81276_new_n1344_), .Y(u5__abc_81276_new_n1345_));
AND2X2 AND2X2_4737 ( .A(u5__abc_81276_new_n1318_), .B(u5__abc_81276_new_n1345_), .Y(u5__abc_81276_new_n1346_));
AND2X2 AND2X2_4738 ( .A(u5__abc_81276_new_n1291_), .B(u5__abc_81276_new_n1346_), .Y(u5__abc_81276_new_n1347_));
AND2X2 AND2X2_4739 ( .A(u5__abc_81276_new_n1242_), .B(u5__abc_81276_new_n1347_), .Y(u5__abc_81276_new_n1348_));
AND2X2 AND2X2_474 ( .A(spec_req_cs_1_bF_buf0_), .B(u0_tms1_26_), .Y(u0__abc_76628_new_n1819_));
AND2X2 AND2X2_4740 ( .A(u5__abc_81276_new_n449__bF_buf6), .B(u5__abc_81276_new_n480__bF_buf3), .Y(u5__abc_81276_new_n1349_));
AND2X2 AND2X2_4741 ( .A(u5__abc_81276_new_n662_), .B(u5__abc_81276_new_n521__bF_buf2), .Y(u5__abc_81276_new_n1350_));
AND2X2 AND2X2_4742 ( .A(u5__abc_81276_new_n1349_), .B(u5__abc_81276_new_n1350_), .Y(u5__abc_81276_new_n1351_));
AND2X2 AND2X2_4743 ( .A(u5__abc_81276_new_n630_), .B(u5__abc_81276_new_n612_), .Y(u5__abc_81276_new_n1353_));
AND2X2 AND2X2_4744 ( .A(u5__abc_81276_new_n1353_), .B(u5__abc_81276_new_n1352_), .Y(u5__abc_81276_new_n1354_));
AND2X2 AND2X2_4745 ( .A(u5__abc_81276_new_n651_), .B(u5__abc_81276_new_n521__bF_buf1), .Y(u5__abc_81276_new_n1355_));
AND2X2 AND2X2_4746 ( .A(u5__abc_81276_new_n1349_), .B(u5__abc_81276_new_n1355_), .Y(u5__abc_81276_new_n1356_));
AND2X2 AND2X2_4747 ( .A(u5__abc_81276_new_n504_), .B(u5__abc_81276_new_n540_), .Y(u5__abc_81276_new_n1358_));
AND2X2 AND2X2_4748 ( .A(u5__abc_81276_new_n520_), .B(u5__abc_81276_new_n1358_), .Y(u5__abc_81276_new_n1359_));
AND2X2 AND2X2_4749 ( .A(u5__abc_81276_new_n501_), .B(u5__abc_81276_new_n1359_), .Y(u5__abc_81276_new_n1360_));
AND2X2 AND2X2_475 ( .A(u0__abc_76628_new_n1169__bF_buf0), .B(u0__abc_76628_new_n1822_), .Y(u0__abc_76628_new_n1823_));
AND2X2 AND2X2_4750 ( .A(u5__abc_81276_new_n643_), .B(u5__abc_81276_new_n521__bF_buf0), .Y(u5__abc_81276_new_n1362_));
AND2X2 AND2X2_4751 ( .A(u5__abc_81276_new_n1349_), .B(u5__abc_81276_new_n1362_), .Y(u5__abc_81276_new_n1363_));
AND2X2 AND2X2_4752 ( .A(u5__abc_81276_new_n1361_), .B(u5__abc_81276_new_n1364_), .Y(u5__abc_81276_new_n1365_));
AND2X2 AND2X2_4753 ( .A(u5__abc_81276_new_n507_), .B(u5__abc_81276_new_n548_), .Y(u5__abc_81276_new_n1366_));
AND2X2 AND2X2_4754 ( .A(u5__abc_81276_new_n520_), .B(u5__abc_81276_new_n1366_), .Y(u5__abc_81276_new_n1367_));
AND2X2 AND2X2_4755 ( .A(u5__abc_81276_new_n501_), .B(u5__abc_81276_new_n1367_), .Y(u5__abc_81276_new_n1368_));
AND2X2 AND2X2_4756 ( .A(u5__abc_81276_new_n634_), .B(u5__abc_81276_new_n520_), .Y(u5__abc_81276_new_n1370_));
AND2X2 AND2X2_4757 ( .A(u5__abc_81276_new_n1370_), .B(u5__abc_81276_new_n517_), .Y(u5__abc_81276_new_n1371_));
AND2X2 AND2X2_4758 ( .A(u5__abc_81276_new_n1349_), .B(u5__abc_81276_new_n1371_), .Y(u5__abc_81276_new_n1372_));
AND2X2 AND2X2_4759 ( .A(u5__abc_81276_new_n1369_), .B(u5__abc_81276_new_n1373_), .Y(u5__abc_81276_new_n1374_));
AND2X2 AND2X2_476 ( .A(u0__abc_76628_new_n1821_), .B(u0__abc_76628_new_n1823_), .Y(u0__abc_76628_new_n1824_));
AND2X2 AND2X2_4760 ( .A(u5__abc_81276_new_n1365_), .B(u5__abc_81276_new_n1374_), .Y(u5__abc_81276_new_n1375_));
AND2X2 AND2X2_4761 ( .A(u5__abc_81276_new_n1375_), .B(u5__abc_81276_new_n1357_), .Y(u5__abc_81276_new_n1376_));
AND2X2 AND2X2_4762 ( .A(u5__abc_81276_new_n1376_), .B(u5__abc_81276_new_n1354_), .Y(u5__abc_81276_new_n1377_));
AND2X2 AND2X2_4763 ( .A(u5__abc_81276_new_n509_), .B(u5_state_28_), .Y(u5__abc_81276_new_n1380_));
AND2X2 AND2X2_4764 ( .A(u5__abc_81276_new_n591_), .B(u5__abc_81276_new_n1380_), .Y(u5__abc_81276_new_n1381_));
AND2X2 AND2X2_4765 ( .A(u5__abc_81276_new_n501_), .B(u5__abc_81276_new_n1381_), .Y(u5__abc_81276_new_n1382_));
AND2X2 AND2X2_4766 ( .A(u5__abc_81276_new_n1379_), .B(u5__abc_81276_new_n1383_), .Y(u5__abc_81276_new_n1384_));
AND2X2 AND2X2_4767 ( .A(u5__abc_81276_new_n1384_), .B(u5__abc_81276_new_n1378_), .Y(u5__abc_81276_new_n1385_));
AND2X2 AND2X2_4768 ( .A(u5__abc_81276_new_n443_), .B(u5_state_33_), .Y(u5__abc_81276_new_n1386_));
AND2X2 AND2X2_4769 ( .A(u5__abc_81276_new_n442_), .B(u5__abc_81276_new_n1386_), .Y(u5__abc_81276_new_n1387_));
AND2X2 AND2X2_477 ( .A(u0__abc_76628_new_n1170__bF_buf0), .B(sp_tms_27_), .Y(u0__abc_76628_new_n1826_));
AND2X2 AND2X2_4770 ( .A(u5__abc_81276_new_n439_), .B(u5__abc_81276_new_n1387_), .Y(u5__abc_81276_new_n1388_));
AND2X2 AND2X2_4771 ( .A(u5__abc_81276_new_n557_), .B(u5__abc_81276_new_n1388_), .Y(u5__abc_81276_new_n1389_));
AND2X2 AND2X2_4772 ( .A(u5__abc_81276_new_n1126__bF_buf1), .B(u5__abc_81276_new_n1389_), .Y(u5__abc_81276_new_n1390_));
AND2X2 AND2X2_4773 ( .A(u5__abc_81276_new_n1391_), .B(u5__abc_81276_new_n1398_), .Y(u5__abc_81276_new_n1399_));
AND2X2 AND2X2_4774 ( .A(u5__abc_81276_new_n463_), .B(u5__abc_81276_new_n452_), .Y(u5__abc_81276_new_n1400_));
AND2X2 AND2X2_4775 ( .A(u5__abc_81276_new_n454_), .B(u5_state_12_), .Y(u5__abc_81276_new_n1401_));
AND2X2 AND2X2_4776 ( .A(u5__abc_81276_new_n490__bF_buf9), .B(u5__abc_81276_new_n1401_), .Y(u5__abc_81276_new_n1402_));
AND2X2 AND2X2_4777 ( .A(u5__abc_81276_new_n479__bF_buf2), .B(u5__abc_81276_new_n1402_), .Y(u5__abc_81276_new_n1403_));
AND2X2 AND2X2_4778 ( .A(u5__abc_81276_new_n1403_), .B(u5__abc_81276_new_n1400_), .Y(u5__abc_81276_new_n1404_));
AND2X2 AND2X2_4779 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1404_), .Y(u5__abc_81276_new_n1405_));
AND2X2 AND2X2_478 ( .A(spec_req_cs_5_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1827_));
AND2X2 AND2X2_4780 ( .A(u5__abc_81276_new_n451_), .B(u5_state_15_), .Y(u5__abc_81276_new_n1407_));
AND2X2 AND2X2_4781 ( .A(u5__abc_81276_new_n490__bF_buf8), .B(u5__abc_81276_new_n1407_), .Y(u5__abc_81276_new_n1408_));
AND2X2 AND2X2_4782 ( .A(u5__abc_81276_new_n1408_), .B(u5__abc_81276_new_n455_), .Y(u5__abc_81276_new_n1409_));
AND2X2 AND2X2_4783 ( .A(u5__abc_81276_new_n1409_), .B(u5__abc_81276_new_n463_), .Y(u5__abc_81276_new_n1410_));
AND2X2 AND2X2_4784 ( .A(u5__abc_81276_new_n1410_), .B(u5__abc_81276_new_n479__bF_buf1), .Y(u5__abc_81276_new_n1411_));
AND2X2 AND2X2_4785 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1411_), .Y(u5__abc_81276_new_n1412_));
AND2X2 AND2X2_4786 ( .A(u5__abc_81276_new_n1406_), .B(u5__abc_81276_new_n1413_), .Y(u5__abc_81276_new_n1414_));
AND2X2 AND2X2_4787 ( .A(u5__abc_81276_new_n1414_), .B(u5__abc_81276_new_n1399_), .Y(u5__abc_81276_new_n1415_));
AND2X2 AND2X2_4788 ( .A(u5__abc_81276_new_n440_), .B(u5_state_34_), .Y(u5__abc_81276_new_n1417_));
AND2X2 AND2X2_4789 ( .A(u5__abc_81276_new_n445_), .B(u5__abc_81276_new_n1417_), .Y(u5__abc_81276_new_n1418_));
AND2X2 AND2X2_479 ( .A(u0__abc_76628_new_n1829_), .B(u0__abc_76628_new_n1179__bF_buf2), .Y(u0__abc_76628_new_n1830_));
AND2X2 AND2X2_4790 ( .A(u5__abc_81276_new_n439_), .B(u5__abc_81276_new_n1418_), .Y(u5__abc_81276_new_n1419_));
AND2X2 AND2X2_4791 ( .A(u5__abc_81276_new_n557_), .B(u5__abc_81276_new_n1419_), .Y(u5__abc_81276_new_n1420_));
AND2X2 AND2X2_4792 ( .A(u5__abc_81276_new_n1126__bF_buf0), .B(u5__abc_81276_new_n1420_), .Y(u5__abc_81276_new_n1421_));
AND2X2 AND2X2_4793 ( .A(u5__abc_81276_new_n1416_), .B(u5__abc_81276_new_n1422_), .Y(u5__abc_81276_new_n1423_));
AND2X2 AND2X2_4794 ( .A(u5__abc_81276_new_n441_), .B(u5_state_35_), .Y(u5__abc_81276_new_n1424_));
AND2X2 AND2X2_4795 ( .A(u5__abc_81276_new_n445_), .B(u5__abc_81276_new_n1424_), .Y(u5__abc_81276_new_n1425_));
AND2X2 AND2X2_4796 ( .A(u5__abc_81276_new_n439_), .B(u5__abc_81276_new_n1425_), .Y(u5__abc_81276_new_n1426_));
AND2X2 AND2X2_4797 ( .A(u5__abc_81276_new_n557_), .B(u5__abc_81276_new_n1426_), .Y(u5__abc_81276_new_n1427_));
AND2X2 AND2X2_4798 ( .A(u5__abc_81276_new_n1126__bF_buf3), .B(u5__abc_81276_new_n1427_), .Y(u5__abc_81276_new_n1428_));
AND2X2 AND2X2_4799 ( .A(u5__abc_81276_new_n503_), .B(u5_state_27_), .Y(u5__abc_81276_new_n1430_));
AND2X2 AND2X2_48 ( .A(_abc_85006_new_n395_), .B(_abc_85006_new_n396_), .Y(csc_s_3_));
AND2X2 AND2X2_480 ( .A(u0__abc_76628_new_n1830_), .B(u0__abc_76628_new_n1828_), .Y(u0__abc_76628_new_n1831_));
AND2X2 AND2X2_4800 ( .A(u5__abc_81276_new_n507_), .B(u5__abc_81276_new_n1430_), .Y(u5__abc_81276_new_n1431_));
AND2X2 AND2X2_4801 ( .A(u5__abc_81276_new_n520_), .B(u5__abc_81276_new_n1431_), .Y(u5__abc_81276_new_n1432_));
AND2X2 AND2X2_4802 ( .A(u5__abc_81276_new_n501_), .B(u5__abc_81276_new_n1432_), .Y(u5__abc_81276_new_n1433_));
AND2X2 AND2X2_4803 ( .A(u5__abc_81276_new_n1429_), .B(u5__abc_81276_new_n1434_), .Y(u5__abc_81276_new_n1435_));
AND2X2 AND2X2_4804 ( .A(u5__abc_81276_new_n1423_), .B(u5__abc_81276_new_n1435_), .Y(u5__abc_81276_new_n1436_));
AND2X2 AND2X2_4805 ( .A(u5__abc_81276_new_n1436_), .B(u5__abc_81276_new_n1415_), .Y(u5__abc_81276_new_n1437_));
AND2X2 AND2X2_4806 ( .A(u5__abc_81276_new_n1437_), .B(u5__abc_81276_new_n1385_), .Y(u5__abc_81276_new_n1438_));
AND2X2 AND2X2_4807 ( .A(u5__abc_81276_new_n453_), .B(u5_state_13_), .Y(u5__abc_81276_new_n1439_));
AND2X2 AND2X2_4808 ( .A(u5__abc_81276_new_n490__bF_buf7), .B(u5__abc_81276_new_n1439_), .Y(u5__abc_81276_new_n1440_));
AND2X2 AND2X2_4809 ( .A(u5__abc_81276_new_n479__bF_buf0), .B(u5__abc_81276_new_n1440_), .Y(u5__abc_81276_new_n1441_));
AND2X2 AND2X2_481 ( .A(u0__abc_76628_new_n1832_), .B(u0__abc_76628_new_n1175__bF_buf2), .Y(u0__abc_76628_new_n1833_));
AND2X2 AND2X2_4810 ( .A(u5__abc_81276_new_n1441_), .B(u5__abc_81276_new_n1400_), .Y(u5__abc_81276_new_n1442_));
AND2X2 AND2X2_4811 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1442_), .Y(u5__abc_81276_new_n1443_));
AND2X2 AND2X2_4812 ( .A(u5__abc_81276_new_n479__bF_buf3), .B(u5__abc_81276_new_n456_), .Y(u5__abc_81276_new_n1445_));
AND2X2 AND2X2_4813 ( .A(u5__abc_81276_new_n460_), .B(u5_state_8_), .Y(u5__abc_81276_new_n1446_));
AND2X2 AND2X2_4814 ( .A(u5__abc_81276_new_n490__bF_buf6), .B(u5__abc_81276_new_n1446_), .Y(u5__abc_81276_new_n1447_));
AND2X2 AND2X2_4815 ( .A(u5__abc_81276_new_n1447_), .B(u5__abc_81276_new_n459_), .Y(u5__abc_81276_new_n1448_));
AND2X2 AND2X2_4816 ( .A(u5__abc_81276_new_n1445_), .B(u5__abc_81276_new_n1448_), .Y(u5__abc_81276_new_n1449_));
AND2X2 AND2X2_4817 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1449_), .Y(u5__abc_81276_new_n1450_));
AND2X2 AND2X2_4818 ( .A(u5__abc_81276_new_n1444_), .B(u5__abc_81276_new_n1451_), .Y(u5__abc_81276_new_n1452_));
AND2X2 AND2X2_4819 ( .A(u5__abc_81276_new_n461_), .B(u5_state_9_), .Y(u5__abc_81276_new_n1453_));
AND2X2 AND2X2_482 ( .A(spec_req_cs_4_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1834_));
AND2X2 AND2X2_4820 ( .A(u5__abc_81276_new_n490__bF_buf5), .B(u5__abc_81276_new_n1453_), .Y(u5__abc_81276_new_n1454_));
AND2X2 AND2X2_4821 ( .A(u5__abc_81276_new_n1454_), .B(u5__abc_81276_new_n459_), .Y(u5__abc_81276_new_n1455_));
AND2X2 AND2X2_4822 ( .A(u5__abc_81276_new_n1445_), .B(u5__abc_81276_new_n1455_), .Y(u5__abc_81276_new_n1456_));
AND2X2 AND2X2_4823 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1456_), .Y(u5__abc_81276_new_n1457_));
AND2X2 AND2X2_4824 ( .A(u5__abc_81276_new_n450_), .B(u5_state_14_), .Y(u5__abc_81276_new_n1459_));
AND2X2 AND2X2_4825 ( .A(u5__abc_81276_new_n490__bF_buf4), .B(u5__abc_81276_new_n1459_), .Y(u5__abc_81276_new_n1460_));
AND2X2 AND2X2_4826 ( .A(u5__abc_81276_new_n1460_), .B(u5__abc_81276_new_n455_), .Y(u5__abc_81276_new_n1461_));
AND2X2 AND2X2_4827 ( .A(u5__abc_81276_new_n1461_), .B(u5__abc_81276_new_n463_), .Y(u5__abc_81276_new_n1462_));
AND2X2 AND2X2_4828 ( .A(u5__abc_81276_new_n1462_), .B(u5__abc_81276_new_n479__bF_buf2), .Y(u5__abc_81276_new_n1463_));
AND2X2 AND2X2_4829 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1463_), .Y(u5__abc_81276_new_n1464_));
AND2X2 AND2X2_483 ( .A(u0__abc_76628_new_n1835_), .B(u0__abc_76628_new_n1174__bF_buf2), .Y(u0__abc_76628_new_n1836_));
AND2X2 AND2X2_4830 ( .A(u5__abc_81276_new_n1458_), .B(u5__abc_81276_new_n1465_), .Y(u5__abc_81276_new_n1466_));
AND2X2 AND2X2_4831 ( .A(u5__abc_81276_new_n1452_), .B(u5__abc_81276_new_n1466_), .Y(u5__abc_81276_new_n1467_));
AND2X2 AND2X2_4832 ( .A(u5__abc_81276_new_n458_), .B(u5_state_11_), .Y(u5__abc_81276_new_n1468_));
AND2X2 AND2X2_4833 ( .A(u5__abc_81276_new_n490__bF_buf3), .B(u5__abc_81276_new_n1468_), .Y(u5__abc_81276_new_n1469_));
AND2X2 AND2X2_4834 ( .A(u5__abc_81276_new_n1469_), .B(u5__abc_81276_new_n462_), .Y(u5__abc_81276_new_n1470_));
AND2X2 AND2X2_4835 ( .A(u5__abc_81276_new_n1445_), .B(u5__abc_81276_new_n1470_), .Y(u5__abc_81276_new_n1471_));
AND2X2 AND2X2_4836 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1471_), .Y(u5__abc_81276_new_n1472_));
AND2X2 AND2X2_4837 ( .A(u5__abc_81276_new_n457_), .B(u5_state_10_), .Y(u5__abc_81276_new_n1474_));
AND2X2 AND2X2_4838 ( .A(u5__abc_81276_new_n490__bF_buf2), .B(u5__abc_81276_new_n1474_), .Y(u5__abc_81276_new_n1475_));
AND2X2 AND2X2_4839 ( .A(u5__abc_81276_new_n1475_), .B(u5__abc_81276_new_n462_), .Y(u5__abc_81276_new_n1476_));
AND2X2 AND2X2_484 ( .A(spec_req_cs_3_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1837_));
AND2X2 AND2X2_4840 ( .A(u5__abc_81276_new_n1445_), .B(u5__abc_81276_new_n1476_), .Y(u5__abc_81276_new_n1477_));
AND2X2 AND2X2_4841 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1477_), .Y(u5__abc_81276_new_n1478_));
AND2X2 AND2X2_4842 ( .A(u5__abc_81276_new_n1473_), .B(u5__abc_81276_new_n1479_), .Y(u5__abc_81276_new_n1480_));
AND2X2 AND2X2_4843 ( .A(u5__abc_81276_new_n464__bF_buf0), .B(u5__abc_81276_new_n470_), .Y(u5__abc_81276_new_n1481_));
AND2X2 AND2X2_4844 ( .A(u5__abc_81276_new_n465_), .B(u5_state_6_), .Y(u5__abc_81276_new_n1482_));
AND2X2 AND2X2_4845 ( .A(u5__abc_81276_new_n490__bF_buf1), .B(u5__abc_81276_new_n1482_), .Y(u5__abc_81276_new_n1483_));
AND2X2 AND2X2_4846 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n1483_), .Y(u5__abc_81276_new_n1484_));
AND2X2 AND2X2_4847 ( .A(u5__abc_81276_new_n1481_), .B(u5__abc_81276_new_n1484_), .Y(u5__abc_81276_new_n1485_));
AND2X2 AND2X2_4848 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1485_), .Y(u5__abc_81276_new_n1486_));
AND2X2 AND2X2_4849 ( .A(u5__abc_81276_new_n466_), .B(u5_state_7_), .Y(u5__abc_81276_new_n1488_));
AND2X2 AND2X2_485 ( .A(u0__abc_76628_new_n1838_), .B(u0__abc_76628_new_n1173__bF_buf2), .Y(u0__abc_76628_new_n1839_));
AND2X2 AND2X2_4850 ( .A(u5__abc_81276_new_n490__bF_buf0), .B(u5__abc_81276_new_n1488_), .Y(u5__abc_81276_new_n1489_));
AND2X2 AND2X2_4851 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n1489_), .Y(u5__abc_81276_new_n1490_));
AND2X2 AND2X2_4852 ( .A(u5__abc_81276_new_n1481_), .B(u5__abc_81276_new_n1490_), .Y(u5__abc_81276_new_n1491_));
AND2X2 AND2X2_4853 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1491_), .Y(u5__abc_81276_new_n1492_));
AND2X2 AND2X2_4854 ( .A(u5__abc_81276_new_n1487_), .B(u5__abc_81276_new_n1493_), .Y(u5__abc_81276_new_n1494_));
AND2X2 AND2X2_4855 ( .A(u5__abc_81276_new_n1480_), .B(u5__abc_81276_new_n1494_), .Y(u5__abc_81276_new_n1495_));
AND2X2 AND2X2_4856 ( .A(u5__abc_81276_new_n1467_), .B(u5__abc_81276_new_n1495_), .Y(u5__abc_81276_new_n1496_));
AND2X2 AND2X2_4857 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n688_), .Y(u5__abc_81276_new_n1497_));
AND2X2 AND2X2_4858 ( .A(u5__abc_81276_new_n1497_), .B(u5__abc_81276_new_n689_), .Y(u5__abc_81276_new_n1498_));
AND2X2 AND2X2_4859 ( .A(u5__abc_81276_new_n1498_), .B(u5__abc_81276_new_n464__bF_buf3), .Y(u5__abc_81276_new_n1499_));
AND2X2 AND2X2_486 ( .A(spec_req_cs_2_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1840_));
AND2X2 AND2X2_4860 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1499_), .Y(u5__abc_81276_new_n1500_));
AND2X2 AND2X2_4861 ( .A(u5__abc_81276_new_n858_), .B(u5__abc_81276_new_n689_), .Y(u5__abc_81276_new_n1502_));
AND2X2 AND2X2_4862 ( .A(u5__abc_81276_new_n1502_), .B(u5__abc_81276_new_n464__bF_buf2), .Y(u5__abc_81276_new_n1503_));
AND2X2 AND2X2_4863 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1503_), .Y(u5__abc_81276_new_n1504_));
AND2X2 AND2X2_4864 ( .A(u5__abc_81276_new_n1501_), .B(u5__abc_81276_new_n1505_), .Y(u5__abc_81276_new_n1506_));
AND2X2 AND2X2_4865 ( .A(u5__abc_81276_new_n501_), .B(u5__abc_81276_new_n592_), .Y(u5__abc_81276_new_n1507_));
AND2X2 AND2X2_4866 ( .A(u5__abc_81276_new_n521__bF_buf2), .B(u5__abc_81276_new_n614_), .Y(u5__abc_81276_new_n1509_));
AND2X2 AND2X2_4867 ( .A(u5__abc_81276_new_n532_), .B(u5__abc_81276_new_n1509_), .Y(u5__abc_81276_new_n1510_));
AND2X2 AND2X2_4868 ( .A(u5__abc_81276_new_n1508_), .B(u5__abc_81276_new_n1511_), .Y(u5__abc_81276_new_n1512_));
AND2X2 AND2X2_4869 ( .A(u5__abc_81276_new_n464__bF_buf1), .B(u5__abc_81276_new_n474_), .Y(u5__abc_81276_new_n1513_));
AND2X2 AND2X2_487 ( .A(u0__abc_76628_new_n1841_), .B(u0__abc_76628_new_n1172__bF_buf2), .Y(u0__abc_76628_new_n1842_));
AND2X2 AND2X2_4870 ( .A(u5__abc_81276_new_n475_), .B(u5_state_0_), .Y(u5__abc_81276_new_n1514_));
AND2X2 AND2X2_4871 ( .A(u5__abc_81276_new_n490__bF_buf10), .B(u5__abc_81276_new_n1514_), .Y(u5__abc_81276_new_n1515_));
AND2X2 AND2X2_4872 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n1515_), .Y(u5__abc_81276_new_n1516_));
AND2X2 AND2X2_4873 ( .A(u5__abc_81276_new_n1513_), .B(u5__abc_81276_new_n1516_), .Y(u5__abc_81276_new_n1517_));
AND2X2 AND2X2_4874 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1517_), .Y(u5__abc_81276_new_n1518_));
AND2X2 AND2X2_4875 ( .A(u5__abc_81276_new_n625_), .B(u5__abc_81276_new_n1519_), .Y(u5__abc_81276_new_n1520_));
AND2X2 AND2X2_4876 ( .A(u5__abc_81276_new_n1512_), .B(u5__abc_81276_new_n1520_), .Y(u5__abc_81276_new_n1521_));
AND2X2 AND2X2_4877 ( .A(u5__abc_81276_new_n1521_), .B(u5__abc_81276_new_n1506_), .Y(u5__abc_81276_new_n1522_));
AND2X2 AND2X2_4878 ( .A(u5__abc_81276_new_n1496_), .B(u5__abc_81276_new_n1522_), .Y(u5__abc_81276_new_n1523_));
AND2X2 AND2X2_4879 ( .A(u5__abc_81276_new_n1523_), .B(u5__abc_81276_new_n1438_), .Y(u5__abc_81276_new_n1524_));
AND2X2 AND2X2_488 ( .A(spec_req_cs_1_bF_buf5_), .B(u0_tms1_27_), .Y(u0__abc_76628_new_n1843_));
AND2X2 AND2X2_4880 ( .A(u5__abc_81276_new_n1524_), .B(u5__abc_81276_new_n1377_), .Y(u5__abc_81276_new_n1525_));
AND2X2 AND2X2_4881 ( .A(u5__abc_81276_new_n1525_), .B(u5__abc_81276_new_n1348_), .Y(u5__abc_81276_new_n1526_));
AND2X2 AND2X2_4882 ( .A(u5__abc_81276_new_n1526__bF_buf3), .B(rfr_req), .Y(u5__abc_81276_new_n1527_));
AND2X2 AND2X2_4883 ( .A(u5__abc_81276_new_n1529_), .B(rfr_ack), .Y(u5__abc_81276_new_n1530_));
AND2X2 AND2X2_4884 ( .A(csc_s_2_), .B(csc_s_1_), .Y(u5__abc_81276_new_n1534_));
AND2X2 AND2X2_4885 ( .A(u5__abc_81276_new_n1534_), .B(u5__abc_81276_new_n1533_), .Y(u5__abc_81276_new_n1535_));
AND2X2 AND2X2_4886 ( .A(u5__abc_81276_new_n1536_), .B(u1_wb_write_go), .Y(u5__abc_81276_new_n1537_));
AND2X2 AND2X2_4887 ( .A(u5__abc_81276_new_n1535_), .B(u5__abc_81276_new_n1537_), .Y(u5__abc_81276_new_n1538_));
AND2X2 AND2X2_4888 ( .A(u5__abc_81276_new_n1547_), .B(u5_lookup_ready2), .Y(u5__abc_81276_new_n1548_));
AND2X2 AND2X2_4889 ( .A(u5__abc_81276_new_n1546_), .B(u5__abc_81276_new_n1548_), .Y(u5__abc_81276_new_n1549_));
AND2X2 AND2X2_489 ( .A(u0__abc_76628_new_n1169__bF_buf6), .B(u0__abc_76628_new_n1846_), .Y(u0__abc_76628_new_n1847_));
AND2X2 AND2X2_4890 ( .A(u5_lookup_ready2), .B(lmr_req), .Y(u5__abc_81276_new_n1550_));
AND2X2 AND2X2_4891 ( .A(u5__abc_81276_new_n1552_), .B(u5_susp_req_r), .Y(u5__abc_81276_new_n1553_));
AND2X2 AND2X2_4892 ( .A(u5__abc_81276_new_n1554_), .B(u5__abc_81276_new_n1551_), .Y(u5__abc_81276_new_n1555_));
AND2X2 AND2X2_4893 ( .A(u5__abc_81276_new_n1556_), .B(u5__abc_81276_new_n1557_), .Y(u5__abc_81276_new_n1558_));
AND2X2 AND2X2_4894 ( .A(u5__abc_81276_new_n1555_), .B(u5__abc_81276_new_n1558_), .Y(u5__abc_81276_new_n1559_));
AND2X2 AND2X2_4895 ( .A(u5__abc_81276_new_n1549_), .B(u5__abc_81276_new_n1559_), .Y(u5__abc_81276_new_n1560_));
AND2X2 AND2X2_4896 ( .A(u5__abc_81276_new_n1526__bF_buf2), .B(u5__abc_81276_new_n1562_), .Y(u5__abc_81276_new_n1563_));
AND2X2 AND2X2_4897 ( .A(u5__abc_81276_new_n1207_), .B(u5__abc_81276_new_n1238_), .Y(u5__abc_81276_new_n1564_));
AND2X2 AND2X2_4898 ( .A(u5__abc_81276_new_n1194_), .B(u5__abc_81276_new_n1564_), .Y(u5__abc_81276_new_n1565_));
AND2X2 AND2X2_4899 ( .A(u5__abc_81276_new_n1473_), .B(u5__abc_81276_new_n1406_), .Y(u5__abc_81276_new_n1566_));
AND2X2 AND2X2_49 ( .A(_abc_85006_new_n398_), .B(_abc_85006_new_n399_), .Y(csc_s_4_));
AND2X2 AND2X2_490 ( .A(u0__abc_76628_new_n1845_), .B(u0__abc_76628_new_n1847_), .Y(u0__abc_76628_new_n1848_));
AND2X2 AND2X2_4900 ( .A(u5__abc_81276_new_n1566_), .B(u5__abc_81276_new_n1399_), .Y(u5__abc_81276_new_n1567_));
AND2X2 AND2X2_4901 ( .A(u5__abc_81276_new_n1385_), .B(u5__abc_81276_new_n1567_), .Y(u5__abc_81276_new_n1568_));
AND2X2 AND2X2_4902 ( .A(u5__abc_81276_new_n1568_), .B(u5__abc_81276_new_n1565_), .Y(u5__abc_81276_new_n1569_));
AND2X2 AND2X2_4903 ( .A(u5__abc_81276_new_n1273_), .B(u5__abc_81276_new_n1261_), .Y(u5__abc_81276_new_n1570_));
AND2X2 AND2X2_4904 ( .A(u5__abc_81276_new_n1451_), .B(u5__abc_81276_new_n1493_), .Y(u5__abc_81276_new_n1571_));
AND2X2 AND2X2_4905 ( .A(u5__abc_81276_new_n1571_), .B(u5__abc_81276_new_n1365_), .Y(u5__abc_81276_new_n1572_));
AND2X2 AND2X2_4906 ( .A(u5__abc_81276_new_n1572_), .B(u5__abc_81276_new_n1570_), .Y(u5__abc_81276_new_n1573_));
AND2X2 AND2X2_4907 ( .A(u5__abc_81276_new_n1429_), .B(u5__abc_81276_new_n1519_), .Y(u5__abc_81276_new_n1574_));
AND2X2 AND2X2_4908 ( .A(u5__abc_81276_new_n612_), .B(u5__abc_81276_new_n1505_), .Y(u5__abc_81276_new_n1575_));
AND2X2 AND2X2_4909 ( .A(u5__abc_81276_new_n1574_), .B(u5__abc_81276_new_n1575_), .Y(u5__abc_81276_new_n1576_));
AND2X2 AND2X2_491 ( .A(u0__abc_76628_new_n1168_), .B(cs_le_d), .Y(u0__abc_76628_new_n1946_));
AND2X2 AND2X2_4910 ( .A(u5__abc_81276_new_n1162_), .B(u5__abc_81276_new_n1423_), .Y(u5__abc_81276_new_n1577_));
AND2X2 AND2X2_4911 ( .A(u5__abc_81276_new_n1576_), .B(u5__abc_81276_new_n1577_), .Y(u5__abc_81276_new_n1578_));
AND2X2 AND2X2_4912 ( .A(u5__abc_81276_new_n1232_), .B(u5__abc_81276_new_n1479_), .Y(u5__abc_81276_new_n1579_));
AND2X2 AND2X2_4913 ( .A(u5__abc_81276_new_n1579_), .B(u5__abc_81276_new_n1216_), .Y(u5__abc_81276_new_n1580_));
AND2X2 AND2X2_4914 ( .A(u5__abc_81276_new_n1580_), .B(u5__abc_81276_new_n1134_), .Y(u5__abc_81276_new_n1581_));
AND2X2 AND2X2_4915 ( .A(u5__abc_81276_new_n1578_), .B(u5__abc_81276_new_n1581_), .Y(u5__abc_81276_new_n1582_));
AND2X2 AND2X2_4916 ( .A(u5__abc_81276_new_n1582_), .B(u5__abc_81276_new_n1573_), .Y(u5__abc_81276_new_n1583_));
AND2X2 AND2X2_4917 ( .A(u5__abc_81276_new_n1583_), .B(u5__abc_81276_new_n1569_), .Y(u5__abc_81276_new_n1584_));
AND2X2 AND2X2_4918 ( .A(u5__abc_81276_new_n1585_), .B(u5_tmr_done_bF_buf3), .Y(u5__abc_81276_new_n1586_));
AND2X2 AND2X2_4919 ( .A(u5__abc_81276_new_n624_), .B(u5__abc_81276_new_n1587_), .Y(u5__abc_81276_new_n1588_));
AND2X2 AND2X2_492 ( .A(u0__abc_76628_new_n1947__bF_buf3), .B(sp_csc_1_), .Y(u0__abc_76628_new_n1972_));
AND2X2 AND2X2_4920 ( .A(u5__abc_81276_new_n1589_), .B(u5__abc_81276_new_n1458_), .Y(u5__abc_81276_new_n1590_));
AND2X2 AND2X2_4921 ( .A(u5__abc_81276_new_n1584_), .B(u5__abc_81276_new_n1590_), .Y(u5__abc_81276_new_n1591_));
AND2X2 AND2X2_4922 ( .A(u5__abc_81276_new_n1324_), .B(u5__abc_81276_new_n1337_), .Y(u5__abc_81276_new_n1592_));
AND2X2 AND2X2_4923 ( .A(u5__abc_81276_new_n1310_), .B(u5__abc_81276_new_n1297_), .Y(u5__abc_81276_new_n1593_));
AND2X2 AND2X2_4924 ( .A(u5__abc_81276_new_n1592_), .B(u5__abc_81276_new_n1593_), .Y(u5__abc_81276_new_n1594_));
AND2X2 AND2X2_4925 ( .A(u5__abc_81276_new_n1316_), .B(u5__abc_81276_new_n1254_), .Y(u5__abc_81276_new_n1595_));
AND2X2 AND2X2_4926 ( .A(u5__abc_81276_new_n1303_), .B(u5__abc_81276_new_n1330_), .Y(u5__abc_81276_new_n1596_));
AND2X2 AND2X2_4927 ( .A(u5__abc_81276_new_n1595_), .B(u5__abc_81276_new_n1596_), .Y(u5__abc_81276_new_n1597_));
AND2X2 AND2X2_4928 ( .A(u5__abc_81276_new_n1594_), .B(u5__abc_81276_new_n1597_), .Y(u5__abc_81276_new_n1598_));
AND2X2 AND2X2_4929 ( .A(u5__abc_81276_new_n1248_), .B(u5__abc_81276_new_n1201_), .Y(u5__abc_81276_new_n1599_));
AND2X2 AND2X2_493 ( .A(spec_req_cs_5_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1973_));
AND2X2 AND2X2_4930 ( .A(u5__abc_81276_new_n1599_), .B(u5__abc_81276_new_n1343_), .Y(u5__abc_81276_new_n1600_));
AND2X2 AND2X2_4931 ( .A(u5__abc_81276_new_n1600_), .B(u5__abc_81276_new_n1148_), .Y(u5__abc_81276_new_n1601_));
AND2X2 AND2X2_4932 ( .A(u5__abc_81276_new_n1598_), .B(u5__abc_81276_new_n1601_), .Y(u5__abc_81276_new_n1602_));
AND2X2 AND2X2_4933 ( .A(u5__abc_81276_new_n1271_), .B(u5__abc_81276_new_n1282_), .Y(u5__abc_81276_new_n1603_));
AND2X2 AND2X2_4934 ( .A(u5__abc_81276_new_n1603_), .B(u5__abc_81276_new_n1487_), .Y(u5__abc_81276_new_n1604_));
AND2X2 AND2X2_4935 ( .A(u5__abc_81276_new_n1606_), .B(u5__abc_81276_new_n1607_), .Y(u5__abc_81276_new_n1608_));
AND2X2 AND2X2_4936 ( .A(u5__abc_81276_new_n1608_), .B(u5__abc_81276_new_n1605_), .Y(u5__abc_81276_new_n1609_));
AND2X2 AND2X2_4937 ( .A(u5__abc_81276_new_n1610_), .B(u5_wb_cycle), .Y(u5__abc_81276_new_n1611_));
AND2X2 AND2X2_4938 ( .A(u5__0burst_act_rd_0_0_), .B(u5__abc_81276_new_n1613_), .Y(u5__abc_81276_new_n1614_));
AND2X2 AND2X2_4939 ( .A(u5__abc_81276_new_n1614_), .B(u5__abc_81276_new_n1612_), .Y(u5__abc_81276_new_n1615_));
AND2X2 AND2X2_494 ( .A(u0__abc_76628_new_n1975_), .B(u0__abc_76628_new_n1179__bF_buf1), .Y(u0__abc_76628_new_n1976_));
AND2X2 AND2X2_4940 ( .A(u5__abc_81276_new_n1613_), .B(u5__abc_81276_new_n1094_), .Y(u5__abc_81276_new_n1616_));
AND2X2 AND2X2_4941 ( .A(u5__abc_81276_new_n1616_), .B(u5_wb_wait), .Y(u5__abc_81276_new_n1617_));
AND2X2 AND2X2_4942 ( .A(u5__abc_81276_new_n1618_), .B(u5__abc_81276_new_n1619_), .Y(u5__abc_81276_new_n1620_));
AND2X2 AND2X2_4943 ( .A(u5__abc_81276_new_n1620_), .B(u5__abc_81276_new_n1615_), .Y(u5__abc_81276_new_n1621_));
AND2X2 AND2X2_4944 ( .A(u5__abc_81276_new_n1622_), .B(u5__abc_81276_new_n1464_), .Y(u5__abc_81276_new_n1623_));
AND2X2 AND2X2_4945 ( .A(u5__abc_81276_new_n1625_), .B(u5__abc_81276_new_n1604_), .Y(u5__abc_81276_new_n1626_));
AND2X2 AND2X2_4946 ( .A(u5__abc_81276_new_n994_), .B(u5_tmr_done_bF_buf2), .Y(u5__abc_81276_new_n1627_));
AND2X2 AND2X2_4947 ( .A(u5__abc_81276_new_n1512_), .B(u5__abc_81276_new_n1373_), .Y(u5__abc_81276_new_n1629_));
AND2X2 AND2X2_4948 ( .A(u5__abc_81276_new_n1629_), .B(u5__abc_81276_new_n1628_), .Y(u5__abc_81276_new_n1630_));
AND2X2 AND2X2_4949 ( .A(u5__abc_81276_new_n1626_), .B(u5__abc_81276_new_n1630_), .Y(u5__abc_81276_new_n1631_));
AND2X2 AND2X2_495 ( .A(u0__abc_76628_new_n1976_), .B(u0__abc_76628_new_n1974_), .Y(u0__abc_76628_new_n1977_));
AND2X2 AND2X2_4950 ( .A(u5__abc_81276_new_n1631_), .B(u5__abc_81276_new_n1602_), .Y(u5__abc_81276_new_n1632_));
AND2X2 AND2X2_4951 ( .A(u5__abc_81276_new_n1591_), .B(u5__abc_81276_new_n1632_), .Y(u5__abc_81276_new_n1633_));
AND2X2 AND2X2_4952 ( .A(u5_cmd_del_0_), .B(u1_wr_cycle), .Y(u5__abc_81276_new_n1636_));
AND2X2 AND2X2_4953 ( .A(u5_cmd_0_), .B(u5__abc_81276_new_n1637_), .Y(u5__abc_81276_new_n1638_));
AND2X2 AND2X2_4954 ( .A(u5__abc_81276_new_n1434_), .B(u5__abc_81276_new_n1357_), .Y(u5__abc_81276_new_n1644_));
AND2X2 AND2X2_4955 ( .A(u5__abc_81276_new_n1644_), .B(u5__abc_81276_new_n630_), .Y(u5__abc_81276_new_n1645_));
AND2X2 AND2X2_4956 ( .A(u5__abc_81276_new_n1501_), .B(u5__abc_81276_new_n1413_), .Y(u5__abc_81276_new_n1646_));
AND2X2 AND2X2_4957 ( .A(u5__abc_81276_new_n1645_), .B(u5__abc_81276_new_n1646_), .Y(u5__abc_81276_new_n1647_));
AND2X2 AND2X2_4958 ( .A(u5__abc_81276_new_n1288_), .B(u5__abc_81276_new_n1267_), .Y(u5__abc_81276_new_n1649_));
AND2X2 AND2X2_4959 ( .A(u5__abc_81276_new_n1225_), .B(u5__abc_81276_new_n1171_), .Y(u5__abc_81276_new_n1650_));
AND2X2 AND2X2_496 ( .A(u0__abc_76628_new_n1978_), .B(u0__abc_76628_new_n1175__bF_buf1), .Y(u0__abc_76628_new_n1979_));
AND2X2 AND2X2_4960 ( .A(u5__abc_81276_new_n1650_), .B(u5__abc_81276_new_n1649_), .Y(u5__abc_81276_new_n1651_));
AND2X2 AND2X2_4961 ( .A(u5__abc_81276_new_n1464_), .B(u5__abc_81276_new_n1655_), .Y(u5__abc_81276_new_n1656_));
AND2X2 AND2X2_4962 ( .A(u1_wr_cycle), .B(u5_cmd_del_1_), .Y(u5__abc_81276_new_n1662_));
AND2X2 AND2X2_4963 ( .A(u5_cmd_1_), .B(u5__abc_81276_new_n1637_), .Y(u5__abc_81276_new_n1663_));
AND2X2 AND2X2_4964 ( .A(u5__abc_81276_new_n1603_), .B(u5__abc_81276_new_n1413_), .Y(u5__abc_81276_new_n1665_));
AND2X2 AND2X2_4965 ( .A(u5__abc_81276_new_n1486_), .B(u5_wb_wait_r), .Y(u5__abc_81276_new_n1666_));
AND2X2 AND2X2_4966 ( .A(u5__abc_81276_new_n1444_), .B(u5__abc_81276_new_n1465_), .Y(u5__abc_81276_new_n1668_));
AND2X2 AND2X2_4967 ( .A(u5__abc_81276_new_n1668_), .B(u5__abc_81276_new_n1667_), .Y(u5__abc_81276_new_n1669_));
AND2X2 AND2X2_4968 ( .A(u5__abc_81276_new_n1665_), .B(u5__abc_81276_new_n1669_), .Y(u5__abc_81276_new_n1670_));
AND2X2 AND2X2_4969 ( .A(u5__abc_81276_new_n1670_), .B(u5__abc_81276_new_n1651_), .Y(u5__abc_81276_new_n1671_));
AND2X2 AND2X2_497 ( .A(spec_req_cs_4_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1980_));
AND2X2 AND2X2_4970 ( .A(u5__abc_81276_new_n1591_), .B(u5__abc_81276_new_n1671_), .Y(u5__abc_81276_new_n1672_));
AND2X2 AND2X2_4971 ( .A(u1_wr_cycle), .B(u5_cmd_del_2_), .Y(u5__abc_81276_new_n1675_));
AND2X2 AND2X2_4972 ( .A(u5_cmd_2_), .B(u5__abc_81276_new_n1637_), .Y(u5__abc_81276_new_n1676_));
AND2X2 AND2X2_4973 ( .A(u5__abc_81276_new_n1679_), .B(mc_c_oe_d), .Y(u5__abc_81276_new_n1680_));
AND2X2 AND2X2_4974 ( .A(u5__abc_81276_new_n1686_), .B(u5__abc_81276_new_n1281_), .Y(u5__abc_81276_new_n1687_));
AND2X2 AND2X2_4975 ( .A(u5__abc_81276_new_n1526__bF_buf0), .B(u5__abc_81276_new_n1560_), .Y(u5__abc_81276_new_n1689_));
AND2X2 AND2X2_4976 ( .A(u5__abc_81276_new_n1123_), .B(u5__abc_81276_new_n1536_), .Y(u5__abc_81276_new_n1693_));
AND2X2 AND2X2_4977 ( .A(u5__abc_81276_new_n1692_), .B(u5__abc_81276_new_n1693_), .Y(u5__abc_81276_new_n1694_));
AND2X2 AND2X2_4978 ( .A(u5__abc_81276_new_n1689_), .B(u5__abc_81276_new_n1694_), .Y(u5__abc_81276_new_n1695_));
AND2X2 AND2X2_4979 ( .A(u5__abc_81276_new_n1695_), .B(u5__abc_81276_new_n1688_), .Y(u5__abc_81276_new_n1696_));
AND2X2 AND2X2_498 ( .A(u0__abc_76628_new_n1981_), .B(u0__abc_76628_new_n1174__bF_buf1), .Y(u0__abc_76628_new_n1982_));
AND2X2 AND2X2_4980 ( .A(u5__abc_81276_new_n1535_), .B(u5__abc_81276_new_n1536_), .Y(u5__abc_81276_new_n1697_));
AND2X2 AND2X2_4981 ( .A(u5__abc_81276_new_n1689_), .B(u5__abc_81276_new_n1697_), .Y(u5__abc_81276_new_n1698_));
AND2X2 AND2X2_4982 ( .A(u5__abc_81276_new_n1486_), .B(u5__abc_81276_new_n1699_), .Y(u5__abc_81276_new_n1700_));
AND2X2 AND2X2_4983 ( .A(u5__abc_81276_new_n624_), .B(u5__abc_81276_new_n1586_), .Y(u5__abc_81276_new_n1702_));
AND2X2 AND2X2_4984 ( .A(u5__abc_81276_new_n1458_), .B(u5__abc_81276_new_n1444_), .Y(u5__abc_81276_new_n1706_));
AND2X2 AND2X2_4985 ( .A(u5__abc_81276_new_n1270_), .B(u5__abc_81276_new_n1708_), .Y(u5__abc_81276_new_n1709_));
AND2X2 AND2X2_4986 ( .A(u5__abc_81276_new_n994_), .B(u5__abc_81276_new_n1712_), .Y(u5__abc_81276_new_n1713_));
AND2X2 AND2X2_4987 ( .A(u5__abc_81276_new_n1714_), .B(u5__abc_81276_new_n1464_), .Y(u5__abc_81276_new_n1715_));
AND2X2 AND2X2_4988 ( .A(u1_wr_cycle), .B(u5_cmd_del_3_), .Y(u5__abc_81276_new_n1724_));
AND2X2 AND2X2_4989 ( .A(u5_cmd_3_), .B(u5__abc_81276_new_n1637_), .Y(u5__abc_81276_new_n1725_));
AND2X2 AND2X2_499 ( .A(spec_req_cs_3_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1983_));
AND2X2 AND2X2_4990 ( .A(u5__abc_81276_new_n1533_), .B(csc_s_2_), .Y(u5__abc_81276_new_n1727_));
AND2X2 AND2X2_4991 ( .A(u5__abc_81276_new_n1728_), .B(u5__abc_81276_new_n1537_), .Y(u5__abc_81276_new_n1729_));
AND2X2 AND2X2_4992 ( .A(u5__abc_81276_new_n1689_), .B(u5__abc_81276_new_n1729_), .Y(u5__abc_81276_new_n1730_));
AND2X2 AND2X2_4993 ( .A(u5__abc_81276_new_n1450_), .B(u5__abc_81276_new_n1537_), .Y(u5__abc_81276_new_n1733_));
AND2X2 AND2X2_4994 ( .A(u5__abc_81276_new_n1215_), .B(u5__abc_81276_new_n1537_), .Y(u5__abc_81276_new_n1734_));
AND2X2 AND2X2_4995 ( .A(u1_wr_cycle), .B(u5_data_oe_r2), .Y(u5__abc_81276_new_n1740_));
AND2X2 AND2X2_4996 ( .A(u5_data_oe_d), .B(u5__abc_81276_new_n1637_), .Y(u5__abc_81276_new_n1741_));
AND2X2 AND2X2_4997 ( .A(u5__abc_81276_new_n1501_), .B(u5__abc_81276_new_n1273_), .Y(u5__abc_81276_new_n1743_));
AND2X2 AND2X2_4998 ( .A(u5__abc_81276_new_n1603_), .B(u5__abc_81276_new_n1743_), .Y(u5__abc_81276_new_n1744_));
AND2X2 AND2X2_4999 ( .A(u5__abc_81276_new_n1649_), .B(u5__abc_81276_new_n1248_), .Y(u5__abc_81276_new_n1745_));
AND2X2 AND2X2_5 ( .A(_abc_85006_new_n251_), .B(_abc_85006_new_n252_), .Y(obct_cs_1_));
AND2X2 AND2X2_50 ( .A(_abc_85006_new_n401_), .B(_abc_85006_new_n402_), .Y(csc_s_5_));
AND2X2 AND2X2_500 ( .A(u0__abc_76628_new_n1984_), .B(u0__abc_76628_new_n1173__bF_buf1), .Y(u0__abc_76628_new_n1985_));
AND2X2 AND2X2_5000 ( .A(u5__abc_81276_new_n1745_), .B(u5__abc_81276_new_n1261_), .Y(u5__abc_81276_new_n1746_));
AND2X2 AND2X2_5001 ( .A(u5__abc_81276_new_n1746_), .B(u5__abc_81276_new_n1744_), .Y(u5__abc_81276_new_n1747_));
AND2X2 AND2X2_5002 ( .A(u5__abc_81276_new_n1174_), .B(u5__abc_81276_new_n1747_), .Y(u5__abc_81276_new_n1748_));
AND2X2 AND2X2_5003 ( .A(u5__abc_81276_new_n1749_), .B(u5__abc_81276_new_n1750_), .Y(u5__abc_81276_new_n1751_));
AND2X2 AND2X2_5004 ( .A(u5__abc_81276_new_n1304_), .B(u5__abc_81276_new_n1751_), .Y(u5__abc_81276_new_n1752_));
AND2X2 AND2X2_5005 ( .A(u5__abc_81276_new_n1310_), .B(u5__abc_81276_new_n1254_), .Y(u5__abc_81276_new_n1753_));
AND2X2 AND2X2_5006 ( .A(u5__abc_81276_new_n1752_), .B(u5__abc_81276_new_n1753_), .Y(u5__abc_81276_new_n1754_));
AND2X2 AND2X2_5007 ( .A(u5__abc_81276_new_n1754_), .B(u5__abc_81276_new_n1345_), .Y(u5__abc_81276_new_n1755_));
AND2X2 AND2X2_5008 ( .A(u5__abc_81276_new_n1755_), .B(u5__abc_81276_new_n1241_), .Y(u5__abc_81276_new_n1756_));
AND2X2 AND2X2_5009 ( .A(u5__abc_81276_new_n1748_), .B(u5__abc_81276_new_n1756_), .Y(u5__abc_81276_new_n1757_));
AND2X2 AND2X2_501 ( .A(spec_req_cs_2_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1986_));
AND2X2 AND2X2_5010 ( .A(u5__abc_81276_new_n1434_), .B(u5__abc_81276_new_n1508_), .Y(u5__abc_81276_new_n1758_));
AND2X2 AND2X2_5011 ( .A(u5__abc_81276_new_n1758_), .B(u5__abc_81276_new_n1384_), .Y(u5__abc_81276_new_n1759_));
AND2X2 AND2X2_5012 ( .A(u5__abc_81276_new_n1429_), .B(u5__abc_81276_new_n1369_), .Y(u5__abc_81276_new_n1760_));
AND2X2 AND2X2_5013 ( .A(u5__abc_81276_new_n1361_), .B(u5__abc_81276_new_n1373_), .Y(u5__abc_81276_new_n1761_));
AND2X2 AND2X2_5014 ( .A(u5__abc_81276_new_n1760_), .B(u5__abc_81276_new_n1761_), .Y(u5__abc_81276_new_n1762_));
AND2X2 AND2X2_5015 ( .A(u5__abc_81276_new_n1759_), .B(u5__abc_81276_new_n1762_), .Y(u5__abc_81276_new_n1763_));
AND2X2 AND2X2_5016 ( .A(u5__abc_81276_new_n476_), .B(u5_state_1_), .Y(u5__abc_81276_new_n1764_));
AND2X2 AND2X2_5017 ( .A(u5__abc_81276_new_n490__bF_buf9), .B(u5__abc_81276_new_n1764_), .Y(u5__abc_81276_new_n1765_));
AND2X2 AND2X2_5018 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n1765_), .Y(u5__abc_81276_new_n1766_));
AND2X2 AND2X2_5019 ( .A(u5__abc_81276_new_n1513_), .B(u5__abc_81276_new_n1766_), .Y(u5__abc_81276_new_n1767_));
AND2X2 AND2X2_502 ( .A(u0__abc_76628_new_n1987_), .B(u0__abc_76628_new_n1172__bF_buf1), .Y(u0__abc_76628_new_n1988_));
AND2X2 AND2X2_5020 ( .A(u5__abc_81276_new_n1149_), .B(u5__abc_81276_new_n1767_), .Y(u5__abc_81276_new_n1768_));
AND2X2 AND2X2_5021 ( .A(u5__abc_81276_new_n625_), .B(u5__abc_81276_new_n1769_), .Y(u5__abc_81276_new_n1770_));
AND2X2 AND2X2_5022 ( .A(u5__abc_81276_new_n1364_), .B(u5__abc_81276_new_n1352_), .Y(u5__abc_81276_new_n1771_));
AND2X2 AND2X2_5023 ( .A(u5__abc_81276_new_n612_), .B(u5__abc_81276_new_n1357_), .Y(u5__abc_81276_new_n1772_));
AND2X2 AND2X2_5024 ( .A(u5__abc_81276_new_n1771_), .B(u5__abc_81276_new_n1772_), .Y(u5__abc_81276_new_n1773_));
AND2X2 AND2X2_5025 ( .A(u5__abc_81276_new_n630_), .B(u5__abc_81276_new_n1511_), .Y(u5__abc_81276_new_n1774_));
AND2X2 AND2X2_5026 ( .A(u5__abc_81276_new_n1773_), .B(u5__abc_81276_new_n1774_), .Y(u5__abc_81276_new_n1775_));
AND2X2 AND2X2_5027 ( .A(u5__abc_81276_new_n1775_), .B(u5__abc_81276_new_n1770_), .Y(u5__abc_81276_new_n1776_));
AND2X2 AND2X2_5028 ( .A(u5__abc_81276_new_n1776_), .B(u5__abc_81276_new_n1763_), .Y(u5__abc_81276_new_n1777_));
AND2X2 AND2X2_5029 ( .A(u5__abc_81276_new_n1479_), .B(u5__abc_81276_new_n1465_), .Y(u5__abc_81276_new_n1778_));
AND2X2 AND2X2_503 ( .A(spec_req_cs_1_bF_buf4_), .B(u0_csc1_1_), .Y(u0__abc_76628_new_n1989_));
AND2X2 AND2X2_5030 ( .A(u5__abc_81276_new_n1706_), .B(u5__abc_81276_new_n1778_), .Y(u5__abc_81276_new_n1779_));
AND2X2 AND2X2_5031 ( .A(u5__abc_81276_new_n1505_), .B(u5__abc_81276_new_n1487_), .Y(u5__abc_81276_new_n1780_));
AND2X2 AND2X2_5032 ( .A(u5__abc_81276_new_n1780_), .B(u5__abc_81276_new_n1571_), .Y(u5__abc_81276_new_n1781_));
AND2X2 AND2X2_5033 ( .A(u5__abc_81276_new_n1779_), .B(u5__abc_81276_new_n1781_), .Y(u5__abc_81276_new_n1782_));
AND2X2 AND2X2_5034 ( .A(u5__abc_81276_new_n1519_), .B(u5__abc_81276_new_n1422_), .Y(u5__abc_81276_new_n1783_));
AND2X2 AND2X2_5035 ( .A(u5__abc_81276_new_n1416_), .B(u5__abc_81276_new_n1391_), .Y(u5__abc_81276_new_n1784_));
AND2X2 AND2X2_5036 ( .A(u5__abc_81276_new_n1413_), .B(u5__abc_81276_new_n1398_), .Y(u5__abc_81276_new_n1785_));
AND2X2 AND2X2_5037 ( .A(u5__abc_81276_new_n1784_), .B(u5__abc_81276_new_n1785_), .Y(u5__abc_81276_new_n1786_));
AND2X2 AND2X2_5038 ( .A(u5__abc_81276_new_n1786_), .B(u5__abc_81276_new_n1783_), .Y(u5__abc_81276_new_n1787_));
AND2X2 AND2X2_5039 ( .A(u5__abc_81276_new_n1787_), .B(u5__abc_81276_new_n1566_), .Y(u5__abc_81276_new_n1788_));
AND2X2 AND2X2_504 ( .A(u0__abc_76628_new_n1946__bF_buf2), .B(u0__abc_76628_new_n1992_), .Y(u0__abc_76628_new_n1993_));
AND2X2 AND2X2_5040 ( .A(u5__abc_81276_new_n1788_), .B(u5__abc_81276_new_n1782_), .Y(u5__abc_81276_new_n1789_));
AND2X2 AND2X2_5041 ( .A(u5__abc_81276_new_n1777_), .B(u5__abc_81276_new_n1789_), .Y(u5__abc_81276_new_n1790_));
AND2X2 AND2X2_5042 ( .A(u5__abc_81276_new_n1790_), .B(u5__abc_81276_new_n1378_), .Y(u5__abc_81276_new_n1791_));
AND2X2 AND2X2_5043 ( .A(u5__abc_81276_new_n1791_), .B(u5__abc_81276_new_n1757_), .Y(u5_pack_le2_d));
AND2X2 AND2X2_5044 ( .A(u5__abc_81276_new_n1494_), .B(u5__abc_81276_new_n1506_), .Y(u5__abc_81276_new_n1793_));
AND2X2 AND2X2_5045 ( .A(u5__abc_81276_new_n1458_), .B(u5__abc_81276_new_n1451_), .Y(u5__abc_81276_new_n1794_));
AND2X2 AND2X2_5046 ( .A(u5__abc_81276_new_n1793_), .B(u5__abc_81276_new_n1794_), .Y(u5__abc_81276_new_n1795_));
AND2X2 AND2X2_5047 ( .A(u5__abc_81276_new_n1406_), .B(u5__abc_81276_new_n1479_), .Y(u5__abc_81276_new_n1796_));
AND2X2 AND2X2_5048 ( .A(u5__abc_81276_new_n1796_), .B(u5__abc_81276_new_n1094_), .Y(u5__abc_81276_new_n1797_));
AND2X2 AND2X2_5049 ( .A(u5__abc_81276_new_n1795_), .B(u5__abc_81276_new_n1797_), .Y(u5__abc_81276_new_n1798_));
AND2X2 AND2X2_505 ( .A(u0__abc_76628_new_n1991_), .B(u0__abc_76628_new_n1993_), .Y(u0__abc_76628_new_n1994_));
AND2X2 AND2X2_5050 ( .A(u5__abc_81276_new_n1348_), .B(u5__abc_81276_new_n1798_), .Y(u5__abc_81276_new_n1799_));
AND2X2 AND2X2_5051 ( .A(u5__abc_81276_new_n1775_), .B(u5__abc_81276_new_n1761_), .Y(u5__abc_81276_new_n1800_));
AND2X2 AND2X2_5052 ( .A(u5__abc_81276_new_n1759_), .B(u5__abc_81276_new_n1378_), .Y(u5__abc_81276_new_n1801_));
AND2X2 AND2X2_5053 ( .A(u5__abc_81276_new_n1760_), .B(u5__abc_81276_new_n1770_), .Y(u5__abc_81276_new_n1802_));
AND2X2 AND2X2_5054 ( .A(u5__abc_81276_new_n1801_), .B(u5__abc_81276_new_n1802_), .Y(u5__abc_81276_new_n1803_));
AND2X2 AND2X2_5055 ( .A(u5__abc_81276_new_n1803_), .B(u5__abc_81276_new_n1787_), .Y(u5__abc_81276_new_n1804_));
AND2X2 AND2X2_5056 ( .A(u5__abc_81276_new_n1804_), .B(u5__abc_81276_new_n1800_), .Y(u5__abc_81276_new_n1805_));
AND2X2 AND2X2_5057 ( .A(u5__abc_81276_new_n1799_), .B(u5__abc_81276_new_n1805_), .Y(u5_cnt_next));
AND2X2 AND2X2_5058 ( .A(u5__abc_81276_new_n1378_), .B(u5_kro), .Y(u5__abc_81276_new_n1807_));
AND2X2 AND2X2_5059 ( .A(u5__abc_81276_new_n1487_), .B(u5__abc_81276_new_n1451_), .Y(u5__abc_81276_new_n1808_));
AND2X2 AND2X2_506 ( .A(u0__abc_76628_new_n1947__bF_buf2), .B(sp_csc_2_), .Y(u0__abc_76628_new_n1996_));
AND2X2 AND2X2_5060 ( .A(u5__abc_81276_new_n1808_), .B(u5__abc_81276_new_n1807_), .Y(u5__abc_81276_new_n1809_));
AND2X2 AND2X2_5061 ( .A(u5__abc_81276_new_n1809_), .B(u5__abc_81276_new_n1506_), .Y(u5__abc_81276_new_n1810_));
AND2X2 AND2X2_5062 ( .A(u5__abc_81276_new_n1810_), .B(u5__abc_81276_new_n1779_), .Y(u5__abc_81276_new_n1811_));
AND2X2 AND2X2_5063 ( .A(u5__abc_81276_new_n1788_), .B(u5__abc_81276_new_n1811_), .Y(u5__abc_81276_new_n1812_));
AND2X2 AND2X2_5064 ( .A(u5__abc_81276_new_n1777_), .B(u5__abc_81276_new_n1812_), .Y(u5__abc_81276_new_n1813_));
AND2X2 AND2X2_5065 ( .A(u5__abc_81276_new_n1813_), .B(u5__abc_81276_new_n1348_), .Y(bank_set));
AND2X2 AND2X2_5066 ( .A(u5__abc_81276_new_n1818_), .B(u5__abc_81276_new_n1816_), .Y(u5__abc_81276_new_n1819_));
AND2X2 AND2X2_5067 ( .A(u5__abc_81276_new_n1819_), .B(u5__abc_81276_new_n1815_), .Y(u5__abc_81276_new_n1820_));
AND2X2 AND2X2_5068 ( .A(wb_we_i), .B(wb_stb_i_bF_buf0), .Y(u5__abc_81276_new_n1822_));
AND2X2 AND2X2_5069 ( .A(u5__abc_81276_new_n1536_), .B(u5__abc_81276_new_n1824_), .Y(u5__abc_81276_new_n1825_));
AND2X2 AND2X2_507 ( .A(spec_req_cs_5_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1997_));
AND2X2 AND2X2_5070 ( .A(u5__abc_81276_new_n1825_), .B(u3_wb_read_go), .Y(u5__abc_81276_new_n1826_));
AND2X2 AND2X2_5071 ( .A(u5__abc_81276_new_n1826_), .B(u5__abc_81276_new_n1823_), .Y(u5__abc_81276_new_n1827_));
AND2X2 AND2X2_5072 ( .A(u5__abc_81276_new_n1821_), .B(u5__abc_81276_new_n1827_), .Y(u5__abc_81276_new_n1828_));
AND2X2 AND2X2_5073 ( .A(u5__abc_81276_new_n1688_), .B(csc_s_1_), .Y(u5__abc_81276_new_n1830_));
AND2X2 AND2X2_5074 ( .A(u5__abc_81276_new_n1830_), .B(u5__abc_81276_new_n1533_), .Y(u5__abc_81276_new_n1831_));
AND2X2 AND2X2_5075 ( .A(u5__abc_81276_new_n1831_), .B(u5__abc_81276_new_n1537_), .Y(u5__abc_81276_new_n1832_));
AND2X2 AND2X2_5076 ( .A(u5__abc_81276_new_n1689_), .B(u5__abc_81276_new_n1832_), .Y(u5__abc_81276_new_n1833_));
AND2X2 AND2X2_5077 ( .A(u5__abc_81276_new_n1835_), .B(u5__0burst_act_rd_0_0_), .Y(u5__abc_81276_new_n1836_));
AND2X2 AND2X2_5078 ( .A(u5__abc_81276_new_n1537_), .B(u5__abc_81276_new_n1824_), .Y(u5__abc_81276_new_n1837_));
AND2X2 AND2X2_5079 ( .A(u5__abc_81276_new_n1837_), .B(u1_wr_cycle), .Y(u5__abc_81276_new_n1838_));
AND2X2 AND2X2_508 ( .A(u0__abc_76628_new_n1999_), .B(u0__abc_76628_new_n1179__bF_buf0), .Y(u0__abc_76628_new_n2000_));
AND2X2 AND2X2_5080 ( .A(u5__abc_81276_new_n1464_), .B(u5__abc_81276_new_n1838_), .Y(u5__abc_81276_new_n1839_));
AND2X2 AND2X2_5081 ( .A(u5__abc_81276_new_n1837_), .B(u5_cmd_asserted_bF_buf3), .Y(u5__abc_81276_new_n1840_));
AND2X2 AND2X2_5082 ( .A(u5__abc_81276_new_n1840_), .B(u5_wb_cycle), .Y(u5__abc_81276_new_n1841_));
AND2X2 AND2X2_5083 ( .A(u5__abc_81276_new_n1443_), .B(u5__abc_81276_new_n1841_), .Y(u5__abc_81276_new_n1842_));
AND2X2 AND2X2_5084 ( .A(u5__abc_81276_new_n1836_), .B(u5__abc_81276_new_n1843_), .Y(u5__abc_81276_new_n1844_));
AND2X2 AND2X2_5085 ( .A(u5__abc_81276_new_n995_), .B(u5__abc_81276_new_n1142_), .Y(u5__abc_81276_new_n1845_));
AND2X2 AND2X2_5086 ( .A(u5__abc_81276_new_n1570_), .B(u5__abc_81276_new_n951_), .Y(u5__abc_81276_new_n1847_));
AND2X2 AND2X2_5087 ( .A(u5__abc_81276_new_n1849_), .B(u5__abc_81276_new_n1840_), .Y(u5__abc_81276_new_n1850_));
AND2X2 AND2X2_5088 ( .A(u1_wb_write_go), .B(u5_tmr_done_bF_buf0), .Y(u5__abc_81276_new_n1851_));
AND2X2 AND2X2_5089 ( .A(u5__abc_81276_new_n1851_), .B(u5__abc_81276_new_n1824_), .Y(u5__abc_81276_new_n1852_));
AND2X2 AND2X2_509 ( .A(u0__abc_76628_new_n2000_), .B(u0__abc_76628_new_n1998_), .Y(u0__abc_76628_new_n2001_));
AND2X2 AND2X2_5090 ( .A(u5__abc_81276_new_n1492_), .B(u5__abc_81276_new_n1852_), .Y(u5__abc_81276_new_n1853_));
AND2X2 AND2X2_5091 ( .A(u5__abc_81276_new_n1450_), .B(u5__abc_81276_new_n1837_), .Y(u5__abc_81276_new_n1854_));
AND2X2 AND2X2_5092 ( .A(u5__abc_81276_new_n1858_), .B(u5__abc_81276_new_n1846_), .Y(u5__abc_81276_new_n1859_));
AND2X2 AND2X2_5093 ( .A(u5__abc_81276_new_n1863_), .B(u5__abc_81276_new_n1829_), .Y(u5__abc_81276_new_n1864_));
AND2X2 AND2X2_5094 ( .A(wb_stb_i_bF_buf5), .B(u5_wb_first), .Y(u5__abc_81276_new_n1867_));
AND2X2 AND2X2_5095 ( .A(u5__abc_81276_new_n1865_), .B(u5__abc_81276_new_n1868_), .Y(u5__0wb_stb_first_0_0_));
AND2X2 AND2X2_5096 ( .A(u5__abc_81276_new_n1034_), .B(u5__abc_81276_new_n1051_), .Y(u5__abc_81276_new_n1871_));
AND2X2 AND2X2_5097 ( .A(u5__abc_81276_new_n415_), .B(u5__abc_81276_new_n402_), .Y(u5__abc_81276_new_n1872_));
AND2X2 AND2X2_5098 ( .A(u5__abc_81276_new_n490__bF_buf8), .B(u5_state_54_), .Y(u5__abc_81276_new_n1873_));
AND2X2 AND2X2_5099 ( .A(u5__abc_81276_new_n1873_), .B(u5__abc_81276_new_n407_), .Y(u5__abc_81276_new_n1874_));
AND2X2 AND2X2_51 ( .A(_abc_85006_new_n404_), .B(_abc_85006_new_n405_), .Y(csc_s_6_));
AND2X2 AND2X2_510 ( .A(u0__abc_76628_new_n2002_), .B(u0__abc_76628_new_n1175__bF_buf0), .Y(u0__abc_76628_new_n2003_));
AND2X2 AND2X2_5100 ( .A(u5__abc_81276_new_n401__bF_buf0), .B(u5__abc_81276_new_n1874_), .Y(u5__abc_81276_new_n1875_));
AND2X2 AND2X2_5101 ( .A(u5__abc_81276_new_n1875_), .B(u5__abc_81276_new_n1872_), .Y(u5__abc_81276_new_n1876_));
AND2X2 AND2X2_5102 ( .A(u5__abc_81276_new_n1876_), .B(u5__abc_81276_new_n448__bF_buf5), .Y(u5__abc_81276_new_n1877_));
AND2X2 AND2X2_5103 ( .A(u5__abc_81276_new_n1877_), .B(u5__abc_81276_new_n523__bF_buf7), .Y(u5__abc_81276_new_n1878_));
AND2X2 AND2X2_5104 ( .A(u5__abc_81276_new_n1042_), .B(u5__abc_81276_new_n1879_), .Y(u5__abc_81276_new_n1880_));
AND2X2 AND2X2_5105 ( .A(u5__abc_81276_new_n1871_), .B(u5__abc_81276_new_n1880_), .Y(u5__abc_81276_new_n1881_));
AND2X2 AND2X2_5106 ( .A(u5__abc_81276_new_n1087_), .B(u5__abc_81276_new_n1881_), .Y(u5__abc_81276_new_n1882_));
AND2X2 AND2X2_5107 ( .A(u5__abc_81276_new_n1006_), .B(u5__abc_81276_new_n1882_), .Y(u5__abc_81276_new_n1883_));
AND2X2 AND2X2_5108 ( .A(u5__abc_81276_new_n703_), .B(u5__abc_81276_new_n721_), .Y(u5__abc_81276_new_n1884_));
AND2X2 AND2X2_5109 ( .A(u5__abc_81276_new_n1884_), .B(u5__abc_81276_new_n713_), .Y(u5__abc_81276_new_n1885_));
AND2X2 AND2X2_511 ( .A(spec_req_cs_4_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n2004_));
AND2X2 AND2X2_5110 ( .A(u5__abc_81276_new_n1885_), .B(u5__abc_81276_new_n728_), .Y(u5__abc_81276_new_n1886_));
AND2X2 AND2X2_5111 ( .A(u5__abc_81276_new_n736_), .B(u5__abc_81276_new_n776_), .Y(u5__abc_81276_new_n1887_));
AND2X2 AND2X2_5112 ( .A(u5__abc_81276_new_n687_), .B(u5__abc_81276_new_n1887_), .Y(u5__abc_81276_new_n1888_));
AND2X2 AND2X2_5113 ( .A(u5__abc_81276_new_n1886_), .B(u5__abc_81276_new_n1888_), .Y(u5__abc_81276_new_n1889_));
AND2X2 AND2X2_5114 ( .A(u5__abc_81276_new_n783_), .B(u5__abc_81276_new_n792_), .Y(u5__abc_81276_new_n1890_));
AND2X2 AND2X2_5115 ( .A(u5__abc_81276_new_n769_), .B(u5__abc_81276_new_n1890_), .Y(u5__abc_81276_new_n1891_));
AND2X2 AND2X2_5116 ( .A(u5__abc_81276_new_n746_), .B(u5__abc_81276_new_n800_), .Y(u5__abc_81276_new_n1892_));
AND2X2 AND2X2_5117 ( .A(u5__abc_81276_new_n753_), .B(u5__abc_81276_new_n1026_), .Y(u5__abc_81276_new_n1893_));
AND2X2 AND2X2_5118 ( .A(u5__abc_81276_new_n1893_), .B(u5__abc_81276_new_n1892_), .Y(u5__abc_81276_new_n1894_));
AND2X2 AND2X2_5119 ( .A(u5__abc_81276_new_n1891_), .B(u5__abc_81276_new_n1894_), .Y(u5__abc_81276_new_n1895_));
AND2X2 AND2X2_512 ( .A(u0__abc_76628_new_n2005_), .B(u0__abc_76628_new_n1174__bF_buf0), .Y(u0__abc_76628_new_n2006_));
AND2X2 AND2X2_5120 ( .A(u5__abc_81276_new_n1889_), .B(u5__abc_81276_new_n1895_), .Y(u5__abc_81276_new_n1896_));
AND2X2 AND2X2_5121 ( .A(u5__abc_81276_new_n1883_), .B(u5__abc_81276_new_n1896_), .Y(u5__abc_81276_new_n1897_));
AND2X2 AND2X2_5122 ( .A(u5__abc_81276_new_n603_), .B(u5__abc_81276_new_n564_), .Y(u5__abc_81276_new_n1898_));
AND2X2 AND2X2_5123 ( .A(u5__abc_81276_new_n946_), .B(u5__abc_81276_new_n1898_), .Y(u5__abc_81276_new_n1899_));
AND2X2 AND2X2_5124 ( .A(u5__abc_81276_new_n589_), .B(u5__abc_81276_new_n907_), .Y(u5__abc_81276_new_n1900_));
AND2X2 AND2X2_5125 ( .A(u5__abc_81276_new_n1899_), .B(u5__abc_81276_new_n1900_), .Y(u5__abc_81276_new_n1901_));
AND2X2 AND2X2_5126 ( .A(u5__abc_81276_new_n854_), .B(u5__abc_81276_new_n837_), .Y(u5__abc_81276_new_n1902_));
AND2X2 AND2X2_5127 ( .A(u5__abc_81276_new_n812_), .B(u5__abc_81276_new_n829_), .Y(u5__abc_81276_new_n1903_));
AND2X2 AND2X2_5128 ( .A(u5__abc_81276_new_n1903_), .B(u5__abc_81276_new_n1902_), .Y(u5__abc_81276_new_n1904_));
AND2X2 AND2X2_5129 ( .A(u5__abc_81276_new_n846_), .B(u5__abc_81276_new_n1018_), .Y(u5__abc_81276_new_n1905_));
AND2X2 AND2X2_513 ( .A(spec_req_cs_3_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n2007_));
AND2X2 AND2X2_5130 ( .A(u5__abc_81276_new_n820_), .B(u5__abc_81276_new_n871_), .Y(u5__abc_81276_new_n1906_));
AND2X2 AND2X2_5131 ( .A(u5__abc_81276_new_n1905_), .B(u5__abc_81276_new_n1906_), .Y(u5__abc_81276_new_n1907_));
AND2X2 AND2X2_5132 ( .A(u5__abc_81276_new_n1904_), .B(u5__abc_81276_new_n1907_), .Y(u5__abc_81276_new_n1908_));
AND2X2 AND2X2_5133 ( .A(u5__abc_81276_new_n695_), .B(u5__abc_81276_new_n863_), .Y(u5__abc_81276_new_n1909_));
AND2X2 AND2X2_5134 ( .A(u5__abc_81276_new_n619_), .B(u5__abc_81276_new_n596_), .Y(u5__abc_81276_new_n1910_));
AND2X2 AND2X2_5135 ( .A(u5__abc_81276_new_n1909_), .B(u5__abc_81276_new_n1910_), .Y(u5__abc_81276_new_n1911_));
AND2X2 AND2X2_5136 ( .A(u5__abc_81276_new_n1908_), .B(u5__abc_81276_new_n1911_), .Y(u5__abc_81276_new_n1912_));
AND2X2 AND2X2_5137 ( .A(u5__abc_81276_new_n556_), .B(u5__abc_81276_new_n648_), .Y(u5__abc_81276_new_n1913_));
AND2X2 AND2X2_5138 ( .A(u5__abc_81276_new_n667_), .B(u5__abc_81276_new_n1353_), .Y(u5__abc_81276_new_n1914_));
AND2X2 AND2X2_5139 ( .A(u5__abc_81276_new_n1914_), .B(u5__abc_81276_new_n1913_), .Y(u5__abc_81276_new_n1915_));
AND2X2 AND2X2_514 ( .A(u0__abc_76628_new_n2008_), .B(u0__abc_76628_new_n1173__bF_buf0), .Y(u0__abc_76628_new_n2009_));
AND2X2 AND2X2_5140 ( .A(u5__abc_81276_new_n625_), .B(u5__abc_81276_new_n890_), .Y(u5__abc_81276_new_n1916_));
AND2X2 AND2X2_5141 ( .A(u5__abc_81276_new_n1915_), .B(u5__abc_81276_new_n1916_), .Y(u5__abc_81276_new_n1917_));
AND2X2 AND2X2_5142 ( .A(u5__abc_81276_new_n1917_), .B(u5__abc_81276_new_n1912_), .Y(u5__abc_81276_new_n1918_));
AND2X2 AND2X2_5143 ( .A(u5__abc_81276_new_n1918_), .B(u5__abc_81276_new_n1901_), .Y(u5__abc_81276_new_n1919_));
AND2X2 AND2X2_5144 ( .A(u5__abc_81276_new_n1897_), .B(u5__abc_81276_new_n1919_), .Y(u5__abc_81276_new_n1920_));
AND2X2 AND2X2_5145 ( .A(u5__abc_81276_new_n1920_), .B(u5__abc_81276_new_n1585_), .Y(u5__abc_81276_new_n1921_));
AND2X2 AND2X2_5146 ( .A(u5__abc_81276_new_n1870_), .B(u5__abc_81276_new_n1921_), .Y(u5__abc_81276_new_n1922_));
AND2X2 AND2X2_5147 ( .A(u5__abc_81276_new_n467_), .B(u5__abc_81276_new_n857_), .Y(u5__abc_81276_new_n1923_));
AND2X2 AND2X2_5148 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n1923_), .Y(u5__abc_81276_new_n1924_));
AND2X2 AND2X2_5149 ( .A(u5__abc_81276_new_n464__bF_buf0), .B(u5__abc_81276_new_n1924_), .Y(u5__abc_81276_new_n1925_));
AND2X2 AND2X2_515 ( .A(spec_req_cs_2_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n2010_));
AND2X2 AND2X2_5150 ( .A(u5__abc_81276_new_n522__bF_buf1), .B(u5__abc_81276_new_n1925_), .Y(u5__abc_81276_new_n1926_));
AND2X2 AND2X2_5151 ( .A(u5__abc_81276_new_n449__bF_buf4), .B(u5__abc_81276_new_n1926_), .Y(u5__abc_81276_new_n1927_));
AND2X2 AND2X2_5152 ( .A(u5__abc_81276_new_n1927_), .B(u5__abc_81276_new_n490__bF_buf7), .Y(u5__abc_81276_new_n1928_));
AND2X2 AND2X2_5153 ( .A(u5__abc_81276_new_n467_), .B(u5__abc_81276_new_n688_), .Y(u5__abc_81276_new_n1930_));
AND2X2 AND2X2_5154 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n1930_), .Y(u5__abc_81276_new_n1931_));
AND2X2 AND2X2_5155 ( .A(u5__abc_81276_new_n464__bF_buf3), .B(u5__abc_81276_new_n1931_), .Y(u5__abc_81276_new_n1932_));
AND2X2 AND2X2_5156 ( .A(u5__abc_81276_new_n522__bF_buf0), .B(u5__abc_81276_new_n1932_), .Y(u5__abc_81276_new_n1933_));
AND2X2 AND2X2_5157 ( .A(u5__abc_81276_new_n449__bF_buf3), .B(u5__abc_81276_new_n1933_), .Y(u5__abc_81276_new_n1934_));
AND2X2 AND2X2_5158 ( .A(u5__abc_81276_new_n1934_), .B(u5__abc_81276_new_n490__bF_buf6), .Y(u5__abc_81276_new_n1935_));
AND2X2 AND2X2_5159 ( .A(u5__abc_81276_new_n1929_), .B(u5__abc_81276_new_n1936_), .Y(u5__abc_81276_new_n1937_));
AND2X2 AND2X2_516 ( .A(u0__abc_76628_new_n2011_), .B(u0__abc_76628_new_n1172__bF_buf0), .Y(u0__abc_76628_new_n2012_));
AND2X2 AND2X2_5160 ( .A(u5__abc_81276_new_n592_), .B(u5__abc_81276_new_n517_), .Y(u5__abc_81276_new_n1938_));
AND2X2 AND2X2_5161 ( .A(u5__abc_81276_new_n1938_), .B(u5__abc_81276_new_n480__bF_buf1), .Y(u5__abc_81276_new_n1939_));
AND2X2 AND2X2_5162 ( .A(u5__abc_81276_new_n1939_), .B(u5__abc_81276_new_n449__bF_buf2), .Y(u5__abc_81276_new_n1940_));
AND2X2 AND2X2_5163 ( .A(u5__abc_81276_new_n1940_), .B(u5__abc_81276_new_n490__bF_buf5), .Y(u5__abc_81276_new_n1941_));
AND2X2 AND2X2_5164 ( .A(u5__abc_81276_new_n497_), .B(u5__abc_81276_new_n614_), .Y(u5__abc_81276_new_n1943_));
AND2X2 AND2X2_5165 ( .A(u5__abc_81276_new_n521__bF_buf1), .B(u5__abc_81276_new_n1943_), .Y(u5__abc_81276_new_n1944_));
AND2X2 AND2X2_5166 ( .A(u5__abc_81276_new_n480__bF_buf0), .B(u5__abc_81276_new_n1944_), .Y(u5__abc_81276_new_n1945_));
AND2X2 AND2X2_5167 ( .A(u5__abc_81276_new_n449__bF_buf1), .B(u5__abc_81276_new_n1945_), .Y(u5__abc_81276_new_n1946_));
AND2X2 AND2X2_5168 ( .A(u5__abc_81276_new_n1946_), .B(u5__abc_81276_new_n490__bF_buf4), .Y(u5__abc_81276_new_n1947_));
AND2X2 AND2X2_5169 ( .A(u5__abc_81276_new_n1942_), .B(u5__abc_81276_new_n1948_), .Y(u5__abc_81276_new_n1949_));
AND2X2 AND2X2_517 ( .A(spec_req_cs_1_bF_buf3_), .B(u0_csc1_2_), .Y(u0__abc_76628_new_n2013_));
AND2X2 AND2X2_5170 ( .A(u5__abc_81276_new_n442_), .B(u5__abc_81276_new_n524_), .Y(u5__abc_81276_new_n1950_));
AND2X2 AND2X2_5171 ( .A(u5__abc_81276_new_n439_), .B(u5__abc_81276_new_n1950_), .Y(u5__abc_81276_new_n1951_));
AND2X2 AND2X2_5172 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n1951_), .Y(u5__abc_81276_new_n1952_));
AND2X2 AND2X2_5173 ( .A(u5__abc_81276_new_n417__bF_buf2), .B(u5__abc_81276_new_n1952_), .Y(u5__abc_81276_new_n1953_));
AND2X2 AND2X2_5174 ( .A(u5__abc_81276_new_n523__bF_buf6), .B(u5__abc_81276_new_n1953_), .Y(u5__abc_81276_new_n1954_));
AND2X2 AND2X2_5175 ( .A(u5__abc_81276_new_n1954_), .B(u5__abc_81276_new_n490__bF_buf3), .Y(u5__abc_81276_new_n1955_));
AND2X2 AND2X2_5176 ( .A(u5__abc_81276_new_n517_), .B(u5__abc_81276_new_n515_), .Y(u5__abc_81276_new_n1957_));
AND2X2 AND2X2_5177 ( .A(u5__abc_81276_new_n480__bF_buf4), .B(u5__abc_81276_new_n1957_), .Y(u5__abc_81276_new_n1958_));
AND2X2 AND2X2_5178 ( .A(u5__abc_81276_new_n449__bF_buf0), .B(u5__abc_81276_new_n1958_), .Y(u5__abc_81276_new_n1959_));
AND2X2 AND2X2_5179 ( .A(u5__abc_81276_new_n1381_), .B(u5__abc_81276_new_n517_), .Y(u5__abc_81276_new_n1961_));
AND2X2 AND2X2_518 ( .A(u0__abc_76628_new_n1946__bF_buf1), .B(u0__abc_76628_new_n2016_), .Y(u0__abc_76628_new_n2017_));
AND2X2 AND2X2_5180 ( .A(u5__abc_81276_new_n1961_), .B(u5__abc_81276_new_n480__bF_buf3), .Y(u5__abc_81276_new_n1962_));
AND2X2 AND2X2_5181 ( .A(u5__abc_81276_new_n1962_), .B(u5__abc_81276_new_n449__bF_buf7), .Y(u5__abc_81276_new_n1963_));
AND2X2 AND2X2_5182 ( .A(u5__abc_81276_new_n1964_), .B(u5__abc_81276_new_n1960_), .Y(u5__abc_81276_new_n1965_));
AND2X2 AND2X2_5183 ( .A(u5__abc_81276_new_n1966_), .B(u5__abc_81276_new_n1435_), .Y(u5__abc_81276_new_n1967_));
AND2X2 AND2X2_5184 ( .A(u5__abc_81276_new_n1967_), .B(u5__abc_81276_new_n1956_), .Y(u5__abc_81276_new_n1968_));
AND2X2 AND2X2_5185 ( .A(u5__abc_81276_new_n517_), .B(u5__abc_81276_new_n1367_), .Y(u5__abc_81276_new_n1969_));
AND2X2 AND2X2_5186 ( .A(u5__abc_81276_new_n480__bF_buf2), .B(u5__abc_81276_new_n1969_), .Y(u5__abc_81276_new_n1970_));
AND2X2 AND2X2_5187 ( .A(u5__abc_81276_new_n449__bF_buf6), .B(u5__abc_81276_new_n1970_), .Y(u5__abc_81276_new_n1971_));
AND2X2 AND2X2_5188 ( .A(u5__abc_81276_new_n517_), .B(u5__abc_81276_new_n1359_), .Y(u5__abc_81276_new_n1972_));
AND2X2 AND2X2_5189 ( .A(u5__abc_81276_new_n480__bF_buf1), .B(u5__abc_81276_new_n1972_), .Y(u5__abc_81276_new_n1973_));
AND2X2 AND2X2_519 ( .A(u0__abc_76628_new_n2015_), .B(u0__abc_76628_new_n2017_), .Y(u0__abc_76628_new_n2018_));
AND2X2 AND2X2_5190 ( .A(u5__abc_81276_new_n449__bF_buf5), .B(u5__abc_81276_new_n1973_), .Y(u5__abc_81276_new_n1974_));
AND2X2 AND2X2_5191 ( .A(u5__abc_81276_new_n1975_), .B(u5__abc_81276_new_n490__bF_buf2), .Y(u5__abc_81276_new_n1976_));
AND2X2 AND2X2_5192 ( .A(u5__abc_81276_new_n504_), .B(u5__abc_81276_new_n632_), .Y(u5__abc_81276_new_n1978_));
AND2X2 AND2X2_5193 ( .A(u5__abc_81276_new_n520_), .B(u5__abc_81276_new_n1978_), .Y(u5__abc_81276_new_n1979_));
AND2X2 AND2X2_5194 ( .A(u5__abc_81276_new_n517_), .B(u5__abc_81276_new_n1979_), .Y(u5__abc_81276_new_n1980_));
AND2X2 AND2X2_5195 ( .A(u5__abc_81276_new_n480__bF_buf0), .B(u5__abc_81276_new_n1980_), .Y(u5__abc_81276_new_n1981_));
AND2X2 AND2X2_5196 ( .A(u5__abc_81276_new_n449__bF_buf4), .B(u5__abc_81276_new_n1981_), .Y(u5__abc_81276_new_n1982_));
AND2X2 AND2X2_5197 ( .A(u5__abc_81276_new_n493_), .B(u5__abc_81276_new_n641_), .Y(u5__abc_81276_new_n1983_));
AND2X2 AND2X2_5198 ( .A(u5__abc_81276_new_n487_), .B(u5__abc_81276_new_n1983_), .Y(u5__abc_81276_new_n1984_));
AND2X2 AND2X2_5199 ( .A(u5__abc_81276_new_n521__bF_buf0), .B(u5__abc_81276_new_n1984_), .Y(u5__abc_81276_new_n1985_));
AND2X2 AND2X2_52 ( .A(_abc_85006_new_n407_), .B(_abc_85006_new_n408_), .Y(csc_s_7_));
AND2X2 AND2X2_520 ( .A(u0__abc_76628_new_n1947__bF_buf1), .B(sp_csc_3_), .Y(u0__abc_76628_new_n2020_));
AND2X2 AND2X2_5200 ( .A(u5__abc_81276_new_n480__bF_buf4), .B(u5__abc_81276_new_n1985_), .Y(u5__abc_81276_new_n1986_));
AND2X2 AND2X2_5201 ( .A(u5__abc_81276_new_n449__bF_buf3), .B(u5__abc_81276_new_n1986_), .Y(u5__abc_81276_new_n1987_));
AND2X2 AND2X2_5202 ( .A(u5__abc_81276_new_n1988_), .B(u5__abc_81276_new_n490__bF_buf1), .Y(u5__abc_81276_new_n1989_));
AND2X2 AND2X2_5203 ( .A(u5__abc_81276_new_n1977_), .B(u5__abc_81276_new_n1990_), .Y(u5__abc_81276_new_n1991_));
AND2X2 AND2X2_5204 ( .A(u5__abc_81276_new_n493_), .B(u5__abc_81276_new_n649_), .Y(u5__abc_81276_new_n1992_));
AND2X2 AND2X2_5205 ( .A(u5__abc_81276_new_n487_), .B(u5__abc_81276_new_n1992_), .Y(u5__abc_81276_new_n1993_));
AND2X2 AND2X2_5206 ( .A(u5__abc_81276_new_n521__bF_buf3), .B(u5__abc_81276_new_n1993_), .Y(u5__abc_81276_new_n1994_));
AND2X2 AND2X2_5207 ( .A(u5__abc_81276_new_n480__bF_buf3), .B(u5__abc_81276_new_n1994_), .Y(u5__abc_81276_new_n1995_));
AND2X2 AND2X2_5208 ( .A(u5__abc_81276_new_n449__bF_buf2), .B(u5__abc_81276_new_n1995_), .Y(u5__abc_81276_new_n1996_));
AND2X2 AND2X2_5209 ( .A(u5__abc_81276_new_n496_), .B(u5__abc_81276_new_n660_), .Y(u5__abc_81276_new_n1997_));
AND2X2 AND2X2_521 ( .A(spec_req_cs_5_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n2021_));
AND2X2 AND2X2_5210 ( .A(u5__abc_81276_new_n487_), .B(u5__abc_81276_new_n1997_), .Y(u5__abc_81276_new_n1998_));
AND2X2 AND2X2_5211 ( .A(u5__abc_81276_new_n521__bF_buf2), .B(u5__abc_81276_new_n1998_), .Y(u5__abc_81276_new_n1999_));
AND2X2 AND2X2_5212 ( .A(u5__abc_81276_new_n480__bF_buf2), .B(u5__abc_81276_new_n1999_), .Y(u5__abc_81276_new_n2000_));
AND2X2 AND2X2_5213 ( .A(u5__abc_81276_new_n449__bF_buf1), .B(u5__abc_81276_new_n2000_), .Y(u5__abc_81276_new_n2001_));
AND2X2 AND2X2_5214 ( .A(u5__abc_81276_new_n2002_), .B(u5__abc_81276_new_n490__bF_buf0), .Y(u5__abc_81276_new_n2003_));
AND2X2 AND2X2_5215 ( .A(u5__abc_81276_new_n497_), .B(u5__abc_81276_new_n609_), .Y(u5__abc_81276_new_n2005_));
AND2X2 AND2X2_5216 ( .A(u5__abc_81276_new_n521__bF_buf1), .B(u5__abc_81276_new_n2005_), .Y(u5__abc_81276_new_n2006_));
AND2X2 AND2X2_5217 ( .A(u5__abc_81276_new_n480__bF_buf1), .B(u5__abc_81276_new_n2006_), .Y(u5__abc_81276_new_n2007_));
AND2X2 AND2X2_5218 ( .A(u5__abc_81276_new_n449__bF_buf0), .B(u5__abc_81276_new_n2007_), .Y(u5__abc_81276_new_n2008_));
AND2X2 AND2X2_5219 ( .A(u5__abc_81276_new_n497_), .B(u5__abc_81276_new_n627_), .Y(u5__abc_81276_new_n2009_));
AND2X2 AND2X2_522 ( .A(u0__abc_76628_new_n2023_), .B(u0__abc_76628_new_n1179__bF_buf5), .Y(u0__abc_76628_new_n2024_));
AND2X2 AND2X2_5220 ( .A(u5__abc_81276_new_n521__bF_buf0), .B(u5__abc_81276_new_n2009_), .Y(u5__abc_81276_new_n2010_));
AND2X2 AND2X2_5221 ( .A(u5__abc_81276_new_n480__bF_buf0), .B(u5__abc_81276_new_n2010_), .Y(u5__abc_81276_new_n2011_));
AND2X2 AND2X2_5222 ( .A(u5__abc_81276_new_n449__bF_buf7), .B(u5__abc_81276_new_n2011_), .Y(u5__abc_81276_new_n2012_));
AND2X2 AND2X2_5223 ( .A(u5__abc_81276_new_n2013_), .B(u5__abc_81276_new_n490__bF_buf10), .Y(u5__abc_81276_new_n2014_));
AND2X2 AND2X2_5224 ( .A(u5__abc_81276_new_n2004_), .B(u5__abc_81276_new_n2015_), .Y(u5__abc_81276_new_n2016_));
AND2X2 AND2X2_5225 ( .A(u5__abc_81276_new_n1991_), .B(u5__abc_81276_new_n2016_), .Y(u5__abc_81276_new_n2017_));
AND2X2 AND2X2_5226 ( .A(u5__abc_81276_new_n1968_), .B(u5__abc_81276_new_n2017_), .Y(u5__abc_81276_new_n2018_));
AND2X2 AND2X2_5227 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n1388_), .Y(u5__abc_81276_new_n2019_));
AND2X2 AND2X2_5228 ( .A(u5__abc_81276_new_n417__bF_buf1), .B(u5__abc_81276_new_n2019_), .Y(u5__abc_81276_new_n2020_));
AND2X2 AND2X2_5229 ( .A(u5__abc_81276_new_n523__bF_buf5), .B(u5__abc_81276_new_n2020_), .Y(u5__abc_81276_new_n2021_));
AND2X2 AND2X2_523 ( .A(u0__abc_76628_new_n2024_), .B(u0__abc_76628_new_n2022_), .Y(u0__abc_76628_new_n2025_));
AND2X2 AND2X2_5230 ( .A(u5__abc_81276_new_n2022_), .B(u5__abc_81276_new_n496_), .Y(u5__abc_81276_new_n2023_));
AND2X2 AND2X2_5231 ( .A(u5__abc_81276_new_n2023_), .B(u5__abc_81276_new_n487_), .Y(u5__abc_81276_new_n2024_));
AND2X2 AND2X2_5232 ( .A(u5__abc_81276_new_n2024_), .B(u5__abc_81276_new_n521__bF_buf3), .Y(u5__abc_81276_new_n2025_));
AND2X2 AND2X2_5233 ( .A(u5__abc_81276_new_n2025_), .B(u5__abc_81276_new_n480__bF_buf4), .Y(u5__abc_81276_new_n2026_));
AND2X2 AND2X2_5234 ( .A(u5__abc_81276_new_n2026_), .B(u5__abc_81276_new_n449__bF_buf6), .Y(u5__abc_81276_new_n2027_));
AND2X2 AND2X2_5235 ( .A(u5__abc_81276_new_n2028_), .B(u5__abc_81276_new_n490__bF_buf9), .Y(u5__abc_81276_new_n2029_));
AND2X2 AND2X2_5236 ( .A(u5__abc_81276_new_n452_), .B(u5__abc_81276_new_n1401_), .Y(u5__abc_81276_new_n2031_));
AND2X2 AND2X2_5237 ( .A(u5__abc_81276_new_n463_), .B(u5__abc_81276_new_n2031_), .Y(u5__abc_81276_new_n2032_));
AND2X2 AND2X2_5238 ( .A(u5__abc_81276_new_n479__bF_buf1), .B(u5__abc_81276_new_n2032_), .Y(u5__abc_81276_new_n2033_));
AND2X2 AND2X2_5239 ( .A(u5__abc_81276_new_n522__bF_buf4), .B(u5__abc_81276_new_n2033_), .Y(u5__abc_81276_new_n2034_));
AND2X2 AND2X2_524 ( .A(u0__abc_76628_new_n2026_), .B(u0__abc_76628_new_n1175__bF_buf5), .Y(u0__abc_76628_new_n2027_));
AND2X2 AND2X2_5240 ( .A(u5__abc_81276_new_n449__bF_buf5), .B(u5__abc_81276_new_n2034_), .Y(u5__abc_81276_new_n2035_));
AND2X2 AND2X2_5241 ( .A(u5__abc_81276_new_n455_), .B(u5__abc_81276_new_n1407_), .Y(u5__abc_81276_new_n2036_));
AND2X2 AND2X2_5242 ( .A(u5__abc_81276_new_n463_), .B(u5__abc_81276_new_n2036_), .Y(u5__abc_81276_new_n2037_));
AND2X2 AND2X2_5243 ( .A(u5__abc_81276_new_n479__bF_buf0), .B(u5__abc_81276_new_n2037_), .Y(u5__abc_81276_new_n2038_));
AND2X2 AND2X2_5244 ( .A(u5__abc_81276_new_n522__bF_buf3), .B(u5__abc_81276_new_n2038_), .Y(u5__abc_81276_new_n2039_));
AND2X2 AND2X2_5245 ( .A(u5__abc_81276_new_n449__bF_buf4), .B(u5__abc_81276_new_n2039_), .Y(u5__abc_81276_new_n2040_));
AND2X2 AND2X2_5246 ( .A(u5__abc_81276_new_n2041_), .B(u5__abc_81276_new_n490__bF_buf8), .Y(u5__abc_81276_new_n2042_));
AND2X2 AND2X2_5247 ( .A(u5__abc_81276_new_n2030_), .B(u5__abc_81276_new_n2043_), .Y(u5__abc_81276_new_n2044_));
AND2X2 AND2X2_5248 ( .A(u5__abc_81276_new_n508_), .B(u5__abc_81276_new_n534_), .Y(u5__abc_81276_new_n2045_));
AND2X2 AND2X2_5249 ( .A(u5__abc_81276_new_n517_), .B(u5__abc_81276_new_n2045_), .Y(u5__abc_81276_new_n2046_));
AND2X2 AND2X2_525 ( .A(spec_req_cs_4_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n2028_));
AND2X2 AND2X2_5250 ( .A(u5__abc_81276_new_n480__bF_buf3), .B(u5__abc_81276_new_n2046_), .Y(u5__abc_81276_new_n2047_));
AND2X2 AND2X2_5251 ( .A(u5__abc_81276_new_n449__bF_buf3), .B(u5__abc_81276_new_n2047_), .Y(u5__abc_81276_new_n2048_));
AND2X2 AND2X2_5252 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n1419_), .Y(u5__abc_81276_new_n2049_));
AND2X2 AND2X2_5253 ( .A(u5__abc_81276_new_n417__bF_buf0), .B(u5__abc_81276_new_n2049_), .Y(u5__abc_81276_new_n2050_));
AND2X2 AND2X2_5254 ( .A(u5__abc_81276_new_n523__bF_buf4), .B(u5__abc_81276_new_n2050_), .Y(u5__abc_81276_new_n2051_));
AND2X2 AND2X2_5255 ( .A(u5__abc_81276_new_n2052_), .B(u5__abc_81276_new_n490__bF_buf7), .Y(u5__abc_81276_new_n2053_));
AND2X2 AND2X2_5256 ( .A(u5__abc_81276_new_n497_), .B(u5__abc_81276_new_n622_), .Y(u5__abc_81276_new_n2055_));
AND2X2 AND2X2_5257 ( .A(u5__abc_81276_new_n521__bF_buf2), .B(u5__abc_81276_new_n2055_), .Y(u5__abc_81276_new_n2056_));
AND2X2 AND2X2_5258 ( .A(u5__abc_81276_new_n480__bF_buf2), .B(u5__abc_81276_new_n2056_), .Y(u5__abc_81276_new_n2057_));
AND2X2 AND2X2_5259 ( .A(u5__abc_81276_new_n449__bF_buf2), .B(u5__abc_81276_new_n2057_), .Y(u5__abc_81276_new_n2058_));
AND2X2 AND2X2_526 ( .A(u0__abc_76628_new_n2029_), .B(u0__abc_76628_new_n1174__bF_buf5), .Y(u0__abc_76628_new_n2030_));
AND2X2 AND2X2_5260 ( .A(u5__abc_81276_new_n474_), .B(u5__abc_81276_new_n1514_), .Y(u5__abc_81276_new_n2060_));
AND2X2 AND2X2_5261 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n2060_), .Y(u5__abc_81276_new_n2061_));
AND2X2 AND2X2_5262 ( .A(u5__abc_81276_new_n464__bF_buf2), .B(u5__abc_81276_new_n2061_), .Y(u5__abc_81276_new_n2062_));
AND2X2 AND2X2_5263 ( .A(u5__abc_81276_new_n522__bF_buf2), .B(u5__abc_81276_new_n2062_), .Y(u5__abc_81276_new_n2063_));
AND2X2 AND2X2_5264 ( .A(u5__abc_81276_new_n449__bF_buf1), .B(u5__abc_81276_new_n2063_), .Y(u5__abc_81276_new_n2064_));
AND2X2 AND2X2_5265 ( .A(u5__abc_81276_new_n2059_), .B(u5__abc_81276_new_n2065_), .Y(u5__abc_81276_new_n2066_));
AND2X2 AND2X2_5266 ( .A(u5__abc_81276_new_n2054_), .B(u5__abc_81276_new_n2067_), .Y(u5__abc_81276_new_n2068_));
AND2X2 AND2X2_5267 ( .A(u5__abc_81276_new_n2044_), .B(u5__abc_81276_new_n2068_), .Y(u5__abc_81276_new_n2069_));
AND2X2 AND2X2_5268 ( .A(u5__abc_81276_new_n462_), .B(u5__abc_81276_new_n1468_), .Y(u5__abc_81276_new_n2070_));
AND2X2 AND2X2_5269 ( .A(u5__abc_81276_new_n456_), .B(u5__abc_81276_new_n2070_), .Y(u5__abc_81276_new_n2071_));
AND2X2 AND2X2_527 ( .A(spec_req_cs_3_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n2031_));
AND2X2 AND2X2_5270 ( .A(u5__abc_81276_new_n479__bF_buf3), .B(u5__abc_81276_new_n2071_), .Y(u5__abc_81276_new_n2072_));
AND2X2 AND2X2_5271 ( .A(u5__abc_81276_new_n522__bF_buf1), .B(u5__abc_81276_new_n2072_), .Y(u5__abc_81276_new_n2073_));
AND2X2 AND2X2_5272 ( .A(u5__abc_81276_new_n449__bF_buf0), .B(u5__abc_81276_new_n2073_), .Y(u5__abc_81276_new_n2074_));
AND2X2 AND2X2_5273 ( .A(u5__abc_81276_new_n462_), .B(u5__abc_81276_new_n1474_), .Y(u5__abc_81276_new_n2075_));
AND2X2 AND2X2_5274 ( .A(u5__abc_81276_new_n456_), .B(u5__abc_81276_new_n2075_), .Y(u5__abc_81276_new_n2076_));
AND2X2 AND2X2_5275 ( .A(u5__abc_81276_new_n479__bF_buf2), .B(u5__abc_81276_new_n2076_), .Y(u5__abc_81276_new_n2077_));
AND2X2 AND2X2_5276 ( .A(u5__abc_81276_new_n522__bF_buf0), .B(u5__abc_81276_new_n2077_), .Y(u5__abc_81276_new_n2078_));
AND2X2 AND2X2_5277 ( .A(u5__abc_81276_new_n449__bF_buf7), .B(u5__abc_81276_new_n2078_), .Y(u5__abc_81276_new_n2079_));
AND2X2 AND2X2_5278 ( .A(u5__abc_81276_new_n2080_), .B(u5__abc_81276_new_n490__bF_buf6), .Y(u5__abc_81276_new_n2081_));
AND2X2 AND2X2_5279 ( .A(u5__abc_81276_new_n459_), .B(u5__abc_81276_new_n1453_), .Y(u5__abc_81276_new_n2083_));
AND2X2 AND2X2_528 ( .A(u0__abc_76628_new_n2032_), .B(u0__abc_76628_new_n1173__bF_buf5), .Y(u0__abc_76628_new_n2033_));
AND2X2 AND2X2_5280 ( .A(u5__abc_81276_new_n456_), .B(u5__abc_81276_new_n2083_), .Y(u5__abc_81276_new_n2084_));
AND2X2 AND2X2_5281 ( .A(u5__abc_81276_new_n479__bF_buf1), .B(u5__abc_81276_new_n2084_), .Y(u5__abc_81276_new_n2085_));
AND2X2 AND2X2_5282 ( .A(u5__abc_81276_new_n522__bF_buf4), .B(u5__abc_81276_new_n2085_), .Y(u5__abc_81276_new_n2086_));
AND2X2 AND2X2_5283 ( .A(u5__abc_81276_new_n449__bF_buf6), .B(u5__abc_81276_new_n2086_), .Y(u5__abc_81276_new_n2087_));
AND2X2 AND2X2_5284 ( .A(u5__abc_81276_new_n455_), .B(u5__abc_81276_new_n1459_), .Y(u5__abc_81276_new_n2088_));
AND2X2 AND2X2_5285 ( .A(u5__abc_81276_new_n463_), .B(u5__abc_81276_new_n2088_), .Y(u5__abc_81276_new_n2089_));
AND2X2 AND2X2_5286 ( .A(u5__abc_81276_new_n479__bF_buf0), .B(u5__abc_81276_new_n2089_), .Y(u5__abc_81276_new_n2090_));
AND2X2 AND2X2_5287 ( .A(u5__abc_81276_new_n522__bF_buf3), .B(u5__abc_81276_new_n2090_), .Y(u5__abc_81276_new_n2091_));
AND2X2 AND2X2_5288 ( .A(u5__abc_81276_new_n449__bF_buf5), .B(u5__abc_81276_new_n2091_), .Y(u5__abc_81276_new_n2092_));
AND2X2 AND2X2_5289 ( .A(u5__abc_81276_new_n2093_), .B(u5__abc_81276_new_n490__bF_buf5), .Y(u5__abc_81276_new_n2094_));
AND2X2 AND2X2_529 ( .A(spec_req_cs_2_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n2034_));
AND2X2 AND2X2_5290 ( .A(u5__abc_81276_new_n2082_), .B(u5__abc_81276_new_n2095_), .Y(u5__abc_81276_new_n2096_));
AND2X2 AND2X2_5291 ( .A(u5__abc_81276_new_n452_), .B(u5__abc_81276_new_n1439_), .Y(u5__abc_81276_new_n2097_));
AND2X2 AND2X2_5292 ( .A(u5__abc_81276_new_n463_), .B(u5__abc_81276_new_n2097_), .Y(u5__abc_81276_new_n2098_));
AND2X2 AND2X2_5293 ( .A(u5__abc_81276_new_n479__bF_buf3), .B(u5__abc_81276_new_n2098_), .Y(u5__abc_81276_new_n2099_));
AND2X2 AND2X2_5294 ( .A(u5__abc_81276_new_n522__bF_buf2), .B(u5__abc_81276_new_n2099_), .Y(u5__abc_81276_new_n2100_));
AND2X2 AND2X2_5295 ( .A(u5__abc_81276_new_n449__bF_buf4), .B(u5__abc_81276_new_n2100_), .Y(u5__abc_81276_new_n2101_));
AND2X2 AND2X2_5296 ( .A(u5__abc_81276_new_n459_), .B(u5__abc_81276_new_n1446_), .Y(u5__abc_81276_new_n2102_));
AND2X2 AND2X2_5297 ( .A(u5__abc_81276_new_n456_), .B(u5__abc_81276_new_n2102_), .Y(u5__abc_81276_new_n2103_));
AND2X2 AND2X2_5298 ( .A(u5__abc_81276_new_n479__bF_buf2), .B(u5__abc_81276_new_n2103_), .Y(u5__abc_81276_new_n2104_));
AND2X2 AND2X2_5299 ( .A(u5__abc_81276_new_n522__bF_buf1), .B(u5__abc_81276_new_n2104_), .Y(u5__abc_81276_new_n2105_));
AND2X2 AND2X2_53 ( .A(_abc_85006_new_n413_), .B(_abc_85006_new_n414_), .Y(u1_bas));
AND2X2 AND2X2_530 ( .A(u0__abc_76628_new_n2035_), .B(u0__abc_76628_new_n1172__bF_buf5), .Y(u0__abc_76628_new_n2036_));
AND2X2 AND2X2_5300 ( .A(u5__abc_81276_new_n449__bF_buf3), .B(u5__abc_81276_new_n2105_), .Y(u5__abc_81276_new_n2106_));
AND2X2 AND2X2_5301 ( .A(u5__abc_81276_new_n2107_), .B(u5__abc_81276_new_n490__bF_buf4), .Y(u5__abc_81276_new_n2108_));
AND2X2 AND2X2_5302 ( .A(u5__abc_81276_new_n470_), .B(u5__abc_81276_new_n1488_), .Y(u5__abc_81276_new_n2110_));
AND2X2 AND2X2_5303 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n2110_), .Y(u5__abc_81276_new_n2111_));
AND2X2 AND2X2_5304 ( .A(u5__abc_81276_new_n464__bF_buf1), .B(u5__abc_81276_new_n2111_), .Y(u5__abc_81276_new_n2112_));
AND2X2 AND2X2_5305 ( .A(u5__abc_81276_new_n522__bF_buf0), .B(u5__abc_81276_new_n2112_), .Y(u5__abc_81276_new_n2113_));
AND2X2 AND2X2_5306 ( .A(u5__abc_81276_new_n449__bF_buf2), .B(u5__abc_81276_new_n2113_), .Y(u5__abc_81276_new_n2114_));
AND2X2 AND2X2_5307 ( .A(u5__abc_81276_new_n470_), .B(u5__abc_81276_new_n1482_), .Y(u5__abc_81276_new_n2115_));
AND2X2 AND2X2_5308 ( .A(u5__abc_81276_new_n478_), .B(u5__abc_81276_new_n2115_), .Y(u5__abc_81276_new_n2116_));
AND2X2 AND2X2_5309 ( .A(u5__abc_81276_new_n464__bF_buf0), .B(u5__abc_81276_new_n2116_), .Y(u5__abc_81276_new_n2117_));
AND2X2 AND2X2_531 ( .A(spec_req_cs_1_bF_buf2_), .B(u0_csc1_3_), .Y(u0__abc_76628_new_n2037_));
AND2X2 AND2X2_5310 ( .A(u5__abc_81276_new_n522__bF_buf4), .B(u5__abc_81276_new_n2117_), .Y(u5__abc_81276_new_n2118_));
AND2X2 AND2X2_5311 ( .A(u5__abc_81276_new_n449__bF_buf1), .B(u5__abc_81276_new_n2118_), .Y(u5__abc_81276_new_n2119_));
AND2X2 AND2X2_5312 ( .A(u5__abc_81276_new_n2120_), .B(u5__abc_81276_new_n490__bF_buf3), .Y(u5__abc_81276_new_n2121_));
AND2X2 AND2X2_5313 ( .A(u5__abc_81276_new_n2109_), .B(u5__abc_81276_new_n2122_), .Y(u5__abc_81276_new_n2123_));
AND2X2 AND2X2_5314 ( .A(u5__abc_81276_new_n2096_), .B(u5__abc_81276_new_n2123_), .Y(u5__abc_81276_new_n2124_));
AND2X2 AND2X2_5315 ( .A(u5__abc_81276_new_n2069_), .B(u5__abc_81276_new_n2124_), .Y(u5__abc_81276_new_n2125_));
AND2X2 AND2X2_5316 ( .A(u5__abc_81276_new_n2018_), .B(u5__abc_81276_new_n2125_), .Y(u5__abc_81276_new_n2126_));
AND2X2 AND2X2_5317 ( .A(u5__abc_81276_new_n414_), .B(u5__abc_81276_new_n672_), .Y(u5__abc_81276_new_n2127_));
AND2X2 AND2X2_5318 ( .A(u5__abc_81276_new_n408_), .B(u5__abc_81276_new_n2127_), .Y(u5__abc_81276_new_n2128_));
AND2X2 AND2X2_5319 ( .A(u5__abc_81276_new_n401__bF_buf3), .B(u5__abc_81276_new_n2128_), .Y(u5__abc_81276_new_n2129_));
AND2X2 AND2X2_532 ( .A(u0__abc_76628_new_n1946__bF_buf0), .B(u0__abc_76628_new_n2040_), .Y(u0__abc_76628_new_n2041_));
AND2X2 AND2X2_5320 ( .A(u5__abc_81276_new_n448__bF_buf4), .B(u5__abc_81276_new_n2129_), .Y(u5__abc_81276_new_n2130_));
AND2X2 AND2X2_5321 ( .A(u5__abc_81276_new_n523__bF_buf3), .B(u5__abc_81276_new_n2130_), .Y(u5__abc_81276_new_n2131_));
AND2X2 AND2X2_5322 ( .A(u5__abc_81276_new_n414_), .B(u5__abc_81276_new_n679_), .Y(u5__abc_81276_new_n2132_));
AND2X2 AND2X2_5323 ( .A(u5__abc_81276_new_n408_), .B(u5__abc_81276_new_n2132_), .Y(u5__abc_81276_new_n2133_));
AND2X2 AND2X2_5324 ( .A(u5__abc_81276_new_n401__bF_buf2), .B(u5__abc_81276_new_n2133_), .Y(u5__abc_81276_new_n2134_));
AND2X2 AND2X2_5325 ( .A(u5__abc_81276_new_n448__bF_buf3), .B(u5__abc_81276_new_n2134_), .Y(u5__abc_81276_new_n2135_));
AND2X2 AND2X2_5326 ( .A(u5__abc_81276_new_n523__bF_buf2), .B(u5__abc_81276_new_n2135_), .Y(u5__abc_81276_new_n2136_));
AND2X2 AND2X2_5327 ( .A(u5__abc_81276_new_n2137_), .B(u5__abc_81276_new_n490__bF_buf2), .Y(u5__abc_81276_new_n2138_));
AND2X2 AND2X2_5328 ( .A(u5__abc_81276_new_n411_), .B(u5__abc_81276_new_n1277_), .Y(u5__abc_81276_new_n2139_));
AND2X2 AND2X2_5329 ( .A(u5__abc_81276_new_n408_), .B(u5__abc_81276_new_n2139_), .Y(u5__abc_81276_new_n2140_));
AND2X2 AND2X2_533 ( .A(u0__abc_76628_new_n2039_), .B(u0__abc_76628_new_n2041_), .Y(u0__abc_76628_new_n2042_));
AND2X2 AND2X2_5330 ( .A(u5__abc_81276_new_n401__bF_buf1), .B(u5__abc_81276_new_n2140_), .Y(u5__abc_81276_new_n2141_));
AND2X2 AND2X2_5331 ( .A(u5__abc_81276_new_n448__bF_buf2), .B(u5__abc_81276_new_n2141_), .Y(u5__abc_81276_new_n2142_));
AND2X2 AND2X2_5332 ( .A(u5__abc_81276_new_n523__bF_buf1), .B(u5__abc_81276_new_n2142_), .Y(u5__abc_81276_new_n2143_));
AND2X2 AND2X2_5333 ( .A(u5__abc_81276_new_n411_), .B(u5__abc_81276_new_n1283_), .Y(u5__abc_81276_new_n2144_));
AND2X2 AND2X2_5334 ( .A(u5__abc_81276_new_n408_), .B(u5__abc_81276_new_n2144_), .Y(u5__abc_81276_new_n2145_));
AND2X2 AND2X2_5335 ( .A(u5__abc_81276_new_n401__bF_buf0), .B(u5__abc_81276_new_n2145_), .Y(u5__abc_81276_new_n2146_));
AND2X2 AND2X2_5336 ( .A(u5__abc_81276_new_n448__bF_buf1), .B(u5__abc_81276_new_n2146_), .Y(u5__abc_81276_new_n2147_));
AND2X2 AND2X2_5337 ( .A(u5__abc_81276_new_n523__bF_buf0), .B(u5__abc_81276_new_n2147_), .Y(u5__abc_81276_new_n2148_));
AND2X2 AND2X2_5338 ( .A(u5__abc_81276_new_n2149_), .B(u5__abc_81276_new_n490__bF_buf1), .Y(u5__abc_81276_new_n2150_));
AND2X2 AND2X2_5339 ( .A(u5__abc_81276_new_n447_), .B(u5__abc_81276_new_n1264_), .Y(u5__abc_81276_new_n2152_));
AND2X2 AND2X2_534 ( .A(u0__abc_76628_new_n1947__bF_buf0), .B(sp_csc_4_), .Y(u0__abc_76628_new_n2044_));
AND2X2 AND2X2_5340 ( .A(u5__abc_81276_new_n417__bF_buf3), .B(u5__abc_81276_new_n2152_), .Y(u5__abc_81276_new_n2153_));
AND2X2 AND2X2_5341 ( .A(u5__abc_81276_new_n523__bF_buf7), .B(u5__abc_81276_new_n2153_), .Y(u5__abc_81276_new_n2154_));
AND2X2 AND2X2_5342 ( .A(u5__abc_81276_new_n447_), .B(u5__abc_81276_new_n1258_), .Y(u5__abc_81276_new_n2155_));
AND2X2 AND2X2_5343 ( .A(u5__abc_81276_new_n417__bF_buf2), .B(u5__abc_81276_new_n2155_), .Y(u5__abc_81276_new_n2156_));
AND2X2 AND2X2_5344 ( .A(u5__abc_81276_new_n523__bF_buf6), .B(u5__abc_81276_new_n2156_), .Y(u5__abc_81276_new_n2157_));
AND2X2 AND2X2_5345 ( .A(u5__abc_81276_new_n2158_), .B(u5__abc_81276_new_n490__bF_buf0), .Y(u5__abc_81276_new_n2159_));
AND2X2 AND2X2_5346 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n1245_), .Y(u5__abc_81276_new_n2160_));
AND2X2 AND2X2_5347 ( .A(u5__abc_81276_new_n417__bF_buf1), .B(u5__abc_81276_new_n2160_), .Y(u5__abc_81276_new_n2161_));
AND2X2 AND2X2_5348 ( .A(u5__abc_81276_new_n523__bF_buf5), .B(u5__abc_81276_new_n2161_), .Y(u5__abc_81276_new_n2162_));
AND2X2 AND2X2_5349 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n1251_), .Y(u5__abc_81276_new_n2163_));
AND2X2 AND2X2_535 ( .A(spec_req_cs_5_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n2045_));
AND2X2 AND2X2_5350 ( .A(u5__abc_81276_new_n417__bF_buf0), .B(u5__abc_81276_new_n2163_), .Y(u5__abc_81276_new_n2164_));
AND2X2 AND2X2_5351 ( .A(u5__abc_81276_new_n523__bF_buf4), .B(u5__abc_81276_new_n2164_), .Y(u5__abc_81276_new_n2165_));
AND2X2 AND2X2_5352 ( .A(u5__abc_81276_new_n2166_), .B(u5__abc_81276_new_n490__bF_buf10), .Y(u5__abc_81276_new_n2167_));
AND2X2 AND2X2_5353 ( .A(u5__abc_81276_new_n1308_), .B(u5__abc_81276_new_n523__bF_buf3), .Y(u5__abc_81276_new_n2170_));
AND2X2 AND2X2_5354 ( .A(u5__abc_81276_new_n447_), .B(u5__abc_81276_new_n1313_), .Y(u5__abc_81276_new_n2171_));
AND2X2 AND2X2_5355 ( .A(u5__abc_81276_new_n417__bF_buf3), .B(u5__abc_81276_new_n2171_), .Y(u5__abc_81276_new_n2172_));
AND2X2 AND2X2_5356 ( .A(u5__abc_81276_new_n523__bF_buf2), .B(u5__abc_81276_new_n2172_), .Y(u5__abc_81276_new_n2173_));
AND2X2 AND2X2_5357 ( .A(u5__abc_81276_new_n2174_), .B(u5__abc_81276_new_n490__bF_buf9), .Y(u5__abc_81276_new_n2175_));
AND2X2 AND2X2_5358 ( .A(u5__abc_81276_new_n447_), .B(u5__abc_81276_new_n1294_), .Y(u5__abc_81276_new_n2176_));
AND2X2 AND2X2_5359 ( .A(u5__abc_81276_new_n417__bF_buf2), .B(u5__abc_81276_new_n2176_), .Y(u5__abc_81276_new_n2177_));
AND2X2 AND2X2_536 ( .A(u0__abc_76628_new_n2047_), .B(u0__abc_76628_new_n1179__bF_buf4), .Y(u0__abc_76628_new_n2048_));
AND2X2 AND2X2_5360 ( .A(u5__abc_81276_new_n523__bF_buf1), .B(u5__abc_81276_new_n2177_), .Y(u5__abc_81276_new_n2178_));
AND2X2 AND2X2_5361 ( .A(u5__abc_81276_new_n447_), .B(u5__abc_81276_new_n1300_), .Y(u5__abc_81276_new_n2179_));
AND2X2 AND2X2_5362 ( .A(u5__abc_81276_new_n417__bF_buf1), .B(u5__abc_81276_new_n2179_), .Y(u5__abc_81276_new_n2180_));
AND2X2 AND2X2_5363 ( .A(u5__abc_81276_new_n523__bF_buf0), .B(u5__abc_81276_new_n2180_), .Y(u5__abc_81276_new_n2181_));
AND2X2 AND2X2_5364 ( .A(u5__abc_81276_new_n2182_), .B(u5__abc_81276_new_n490__bF_buf8), .Y(u5__abc_81276_new_n2183_));
AND2X2 AND2X2_5365 ( .A(u5__abc_81276_new_n447_), .B(u5__abc_81276_new_n1321_), .Y(u5__abc_81276_new_n2185_));
AND2X2 AND2X2_5366 ( .A(u5__abc_81276_new_n417__bF_buf0), .B(u5__abc_81276_new_n2185_), .Y(u5__abc_81276_new_n2186_));
AND2X2 AND2X2_5367 ( .A(u5__abc_81276_new_n523__bF_buf7), .B(u5__abc_81276_new_n2186_), .Y(u5__abc_81276_new_n2187_));
AND2X2 AND2X2_5368 ( .A(u5__abc_81276_new_n447_), .B(u5__abc_81276_new_n1327_), .Y(u5__abc_81276_new_n2188_));
AND2X2 AND2X2_5369 ( .A(u5__abc_81276_new_n417__bF_buf3), .B(u5__abc_81276_new_n2188_), .Y(u5__abc_81276_new_n2189_));
AND2X2 AND2X2_537 ( .A(u0__abc_76628_new_n2048_), .B(u0__abc_76628_new_n2046_), .Y(u0__abc_76628_new_n2049_));
AND2X2 AND2X2_5370 ( .A(u5__abc_81276_new_n523__bF_buf6), .B(u5__abc_81276_new_n2189_), .Y(u5__abc_81276_new_n2190_));
AND2X2 AND2X2_5371 ( .A(u5__abc_81276_new_n2191_), .B(u5__abc_81276_new_n490__bF_buf7), .Y(u5__abc_81276_new_n2192_));
AND2X2 AND2X2_5372 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n1334_), .Y(u5__abc_81276_new_n2193_));
AND2X2 AND2X2_5373 ( .A(u5__abc_81276_new_n417__bF_buf2), .B(u5__abc_81276_new_n2193_), .Y(u5__abc_81276_new_n2194_));
AND2X2 AND2X2_5374 ( .A(u5__abc_81276_new_n523__bF_buf5), .B(u5__abc_81276_new_n2194_), .Y(u5__abc_81276_new_n2195_));
AND2X2 AND2X2_5375 ( .A(u5__abc_81276_new_n432_), .B(u5__abc_81276_new_n1340_), .Y(u5__abc_81276_new_n2196_));
AND2X2 AND2X2_5376 ( .A(u5__abc_81276_new_n417__bF_buf1), .B(u5__abc_81276_new_n2196_), .Y(u5__abc_81276_new_n2197_));
AND2X2 AND2X2_5377 ( .A(u5__abc_81276_new_n523__bF_buf4), .B(u5__abc_81276_new_n2197_), .Y(u5__abc_81276_new_n2198_));
AND2X2 AND2X2_5378 ( .A(u5__abc_81276_new_n2199_), .B(u5__abc_81276_new_n490__bF_buf6), .Y(u5__abc_81276_new_n2200_));
AND2X2 AND2X2_5379 ( .A(u5__abc_81276_new_n948_), .B(u5__abc_81276_new_n2204_), .Y(u5__abc_81276_new_n2205_));
AND2X2 AND2X2_538 ( .A(u0__abc_76628_new_n2050_), .B(u0__abc_76628_new_n1175__bF_buf4), .Y(u0__abc_76628_new_n2051_));
AND2X2 AND2X2_5380 ( .A(u5__abc_81276_new_n523__bF_buf3), .B(u5__abc_81276_new_n1131_), .Y(u5__abc_81276_new_n2206_));
AND2X2 AND2X2_5381 ( .A(u5__abc_81276_new_n392_), .B(u5__abc_81276_new_n1164_), .Y(u5__abc_81276_new_n2207_));
AND2X2 AND2X2_5382 ( .A(u5__abc_81276_new_n400_), .B(u5__abc_81276_new_n2207_), .Y(u5__abc_81276_new_n2208_));
AND2X2 AND2X2_5383 ( .A(u5__abc_81276_new_n416__bF_buf0), .B(u5__abc_81276_new_n2208_), .Y(u5__abc_81276_new_n2209_));
AND2X2 AND2X2_5384 ( .A(u5__abc_81276_new_n448__bF_buf0), .B(u5__abc_81276_new_n2209_), .Y(u5__abc_81276_new_n2210_));
AND2X2 AND2X2_5385 ( .A(u5__abc_81276_new_n523__bF_buf2), .B(u5__abc_81276_new_n2210_), .Y(u5__abc_81276_new_n2211_));
AND2X2 AND2X2_5386 ( .A(u5__abc_81276_new_n2212_), .B(u5__abc_81276_new_n490__bF_buf5), .Y(u5__abc_81276_new_n2213_));
AND2X2 AND2X2_5387 ( .A(u5__abc_81276_new_n389_), .B(u5__abc_81276_new_n1143_), .Y(u5__abc_81276_new_n2215_));
AND2X2 AND2X2_5388 ( .A(u5__abc_81276_new_n400_), .B(u5__abc_81276_new_n2215_), .Y(u5__abc_81276_new_n2216_));
AND2X2 AND2X2_5389 ( .A(u5__abc_81276_new_n416__bF_buf3), .B(u5__abc_81276_new_n2216_), .Y(u5__abc_81276_new_n2217_));
AND2X2 AND2X2_539 ( .A(spec_req_cs_4_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n2052_));
AND2X2 AND2X2_5390 ( .A(u5__abc_81276_new_n448__bF_buf5), .B(u5__abc_81276_new_n2217_), .Y(u5__abc_81276_new_n2218_));
AND2X2 AND2X2_5391 ( .A(u5__abc_81276_new_n523__bF_buf1), .B(u5__abc_81276_new_n2218_), .Y(u5__abc_81276_new_n2219_));
AND2X2 AND2X2_5392 ( .A(u5__abc_81276_new_n389_), .B(u5__abc_81276_new_n1138_), .Y(u5__abc_81276_new_n2220_));
AND2X2 AND2X2_5393 ( .A(u5__abc_81276_new_n400_), .B(u5__abc_81276_new_n2220_), .Y(u5__abc_81276_new_n2221_));
AND2X2 AND2X2_5394 ( .A(u5__abc_81276_new_n416__bF_buf2), .B(u5__abc_81276_new_n2221_), .Y(u5__abc_81276_new_n2222_));
AND2X2 AND2X2_5395 ( .A(u5__abc_81276_new_n448__bF_buf4), .B(u5__abc_81276_new_n2222_), .Y(u5__abc_81276_new_n2223_));
AND2X2 AND2X2_5396 ( .A(u5__abc_81276_new_n523__bF_buf0), .B(u5__abc_81276_new_n2223_), .Y(u5__abc_81276_new_n2224_));
AND2X2 AND2X2_5397 ( .A(u5__abc_81276_new_n2225_), .B(u5__abc_81276_new_n490__bF_buf4), .Y(u5__abc_81276_new_n2226_));
AND2X2 AND2X2_5398 ( .A(u5__abc_81276_new_n477_), .B(u5__abc_81276_new_n1157_), .Y(u5__abc_81276_new_n2227_));
AND2X2 AND2X2_5399 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n2227_), .Y(u5__abc_81276_new_n2228_));
AND2X2 AND2X2_54 ( .A(_abc_85006_new_n416_), .B(_abc_85006_new_n417_), .Y(u5_kro));
AND2X2 AND2X2_540 ( .A(u0__abc_76628_new_n2053_), .B(u0__abc_76628_new_n1174__bF_buf4), .Y(u0__abc_76628_new_n2054_));
AND2X2 AND2X2_5400 ( .A(u5__abc_81276_new_n464__bF_buf3), .B(u5__abc_81276_new_n2228_), .Y(u5__abc_81276_new_n2229_));
AND2X2 AND2X2_5401 ( .A(u5__abc_81276_new_n522__bF_buf3), .B(u5__abc_81276_new_n2229_), .Y(u5__abc_81276_new_n2230_));
AND2X2 AND2X2_5402 ( .A(u5__abc_81276_new_n449__bF_buf0), .B(u5__abc_81276_new_n2230_), .Y(u5__abc_81276_new_n2231_));
AND2X2 AND2X2_5403 ( .A(u5__abc_81276_new_n477_), .B(u5__abc_81276_new_n1152_), .Y(u5__abc_81276_new_n2232_));
AND2X2 AND2X2_5404 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n2232_), .Y(u5__abc_81276_new_n2233_));
AND2X2 AND2X2_5405 ( .A(u5__abc_81276_new_n464__bF_buf2), .B(u5__abc_81276_new_n2233_), .Y(u5__abc_81276_new_n2234_));
AND2X2 AND2X2_5406 ( .A(u5__abc_81276_new_n522__bF_buf2), .B(u5__abc_81276_new_n2234_), .Y(u5__abc_81276_new_n2235_));
AND2X2 AND2X2_5407 ( .A(u5__abc_81276_new_n449__bF_buf7), .B(u5__abc_81276_new_n2235_), .Y(u5__abc_81276_new_n2236_));
AND2X2 AND2X2_5408 ( .A(u5__abc_81276_new_n2237_), .B(u5__abc_81276_new_n490__bF_buf3), .Y(u5__abc_81276_new_n2238_));
AND2X2 AND2X2_5409 ( .A(u5__abc_81276_new_n393_), .B(u5__abc_81276_new_n1212_), .Y(u5__abc_81276_new_n2241_));
AND2X2 AND2X2_541 ( .A(spec_req_cs_3_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n2055_));
AND2X2 AND2X2_5410 ( .A(u5__abc_81276_new_n416__bF_buf1), .B(u5__abc_81276_new_n2241_), .Y(u5__abc_81276_new_n2242_));
AND2X2 AND2X2_5411 ( .A(u5__abc_81276_new_n448__bF_buf3), .B(u5__abc_81276_new_n2242_), .Y(u5__abc_81276_new_n2243_));
AND2X2 AND2X2_5412 ( .A(u5__abc_81276_new_n523__bF_buf7), .B(u5__abc_81276_new_n2243_), .Y(u5__abc_81276_new_n2244_));
AND2X2 AND2X2_5413 ( .A(u5__abc_81276_new_n2245_), .B(u5__abc_81276_new_n399_), .Y(u5__abc_81276_new_n2246_));
AND2X2 AND2X2_5414 ( .A(u5__abc_81276_new_n2246_), .B(u5__abc_81276_new_n393_), .Y(u5__abc_81276_new_n2247_));
AND2X2 AND2X2_5415 ( .A(u5__abc_81276_new_n2247_), .B(u5__abc_81276_new_n416__bF_buf0), .Y(u5__abc_81276_new_n2248_));
AND2X2 AND2X2_5416 ( .A(u5__abc_81276_new_n2248_), .B(u5__abc_81276_new_n448__bF_buf2), .Y(u5__abc_81276_new_n2249_));
AND2X2 AND2X2_5417 ( .A(u5__abc_81276_new_n2249_), .B(u5__abc_81276_new_n523__bF_buf6), .Y(u5__abc_81276_new_n2250_));
AND2X2 AND2X2_5418 ( .A(u5__abc_81276_new_n2251_), .B(u5__abc_81276_new_n490__bF_buf2), .Y(u5__abc_81276_new_n2252_));
AND2X2 AND2X2_5419 ( .A(u5__abc_81276_new_n396_), .B(u5__abc_81276_new_n1227_), .Y(u5__abc_81276_new_n2253_));
AND2X2 AND2X2_542 ( .A(u0__abc_76628_new_n2056_), .B(u0__abc_76628_new_n1173__bF_buf4), .Y(u0__abc_76628_new_n2057_));
AND2X2 AND2X2_5420 ( .A(u5__abc_81276_new_n393_), .B(u5__abc_81276_new_n2253_), .Y(u5__abc_81276_new_n2254_));
AND2X2 AND2X2_5421 ( .A(u5__abc_81276_new_n416__bF_buf3), .B(u5__abc_81276_new_n2254_), .Y(u5__abc_81276_new_n2255_));
AND2X2 AND2X2_5422 ( .A(u5__abc_81276_new_n448__bF_buf1), .B(u5__abc_81276_new_n2255_), .Y(u5__abc_81276_new_n2256_));
AND2X2 AND2X2_5423 ( .A(u5__abc_81276_new_n523__bF_buf5), .B(u5__abc_81276_new_n2256_), .Y(u5__abc_81276_new_n2257_));
AND2X2 AND2X2_5424 ( .A(u5__abc_81276_new_n396_), .B(u5__abc_81276_new_n1177_), .Y(u5__abc_81276_new_n2258_));
AND2X2 AND2X2_5425 ( .A(u5__abc_81276_new_n393_), .B(u5__abc_81276_new_n2258_), .Y(u5__abc_81276_new_n2259_));
AND2X2 AND2X2_5426 ( .A(u5__abc_81276_new_n416__bF_buf2), .B(u5__abc_81276_new_n2259_), .Y(u5__abc_81276_new_n2260_));
AND2X2 AND2X2_5427 ( .A(u5__abc_81276_new_n448__bF_buf0), .B(u5__abc_81276_new_n2260_), .Y(u5__abc_81276_new_n2261_));
AND2X2 AND2X2_5428 ( .A(u5__abc_81276_new_n523__bF_buf4), .B(u5__abc_81276_new_n2261_), .Y(u5__abc_81276_new_n2262_));
AND2X2 AND2X2_5429 ( .A(u5__abc_81276_new_n2263_), .B(u5__abc_81276_new_n490__bF_buf1), .Y(u5__abc_81276_new_n2264_));
AND2X2 AND2X2_543 ( .A(spec_req_cs_2_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n2058_));
AND2X2 AND2X2_5430 ( .A(u5__abc_81276_new_n404_), .B(u5__abc_81276_new_n1202_), .Y(u5__abc_81276_new_n2266_));
AND2X2 AND2X2_5431 ( .A(u5__abc_81276_new_n415_), .B(u5__abc_81276_new_n2266_), .Y(u5__abc_81276_new_n2267_));
AND2X2 AND2X2_5432 ( .A(u5__abc_81276_new_n401__bF_buf3), .B(u5__abc_81276_new_n2267_), .Y(u5__abc_81276_new_n2268_));
AND2X2 AND2X2_5433 ( .A(u5__abc_81276_new_n448__bF_buf5), .B(u5__abc_81276_new_n2268_), .Y(u5__abc_81276_new_n2269_));
AND2X2 AND2X2_5434 ( .A(u5__abc_81276_new_n523__bF_buf3), .B(u5__abc_81276_new_n2269_), .Y(u5__abc_81276_new_n2270_));
AND2X2 AND2X2_5435 ( .A(u5__abc_81276_new_n404_), .B(u5__abc_81276_new_n1196_), .Y(u5__abc_81276_new_n2271_));
AND2X2 AND2X2_5436 ( .A(u5__abc_81276_new_n415_), .B(u5__abc_81276_new_n2271_), .Y(u5__abc_81276_new_n2272_));
AND2X2 AND2X2_5437 ( .A(u5__abc_81276_new_n401__bF_buf2), .B(u5__abc_81276_new_n2272_), .Y(u5__abc_81276_new_n2273_));
AND2X2 AND2X2_5438 ( .A(u5__abc_81276_new_n448__bF_buf4), .B(u5__abc_81276_new_n2273_), .Y(u5__abc_81276_new_n2274_));
AND2X2 AND2X2_5439 ( .A(u5__abc_81276_new_n523__bF_buf2), .B(u5__abc_81276_new_n2274_), .Y(u5__abc_81276_new_n2275_));
AND2X2 AND2X2_544 ( .A(u0__abc_76628_new_n2059_), .B(u0__abc_76628_new_n1172__bF_buf4), .Y(u0__abc_76628_new_n2060_));
AND2X2 AND2X2_5440 ( .A(u5__abc_81276_new_n2276_), .B(u5__abc_81276_new_n490__bF_buf0), .Y(u5__abc_81276_new_n2277_));
AND2X2 AND2X2_5441 ( .A(u5__abc_81276_new_n2278_), .B(u5__abc_81276_new_n407_), .Y(u5__abc_81276_new_n2279_));
AND2X2 AND2X2_5442 ( .A(u5__abc_81276_new_n2279_), .B(u5__abc_81276_new_n415_), .Y(u5__abc_81276_new_n2280_));
AND2X2 AND2X2_5443 ( .A(u5__abc_81276_new_n2280_), .B(u5__abc_81276_new_n401__bF_buf1), .Y(u5__abc_81276_new_n2281_));
AND2X2 AND2X2_5444 ( .A(u5__abc_81276_new_n2281_), .B(u5__abc_81276_new_n448__bF_buf3), .Y(u5__abc_81276_new_n2282_));
AND2X2 AND2X2_5445 ( .A(u5__abc_81276_new_n2282_), .B(u5__abc_81276_new_n523__bF_buf1), .Y(u5__abc_81276_new_n2283_));
AND2X2 AND2X2_5446 ( .A(u5__abc_81276_new_n407_), .B(u5__abc_81276_new_n1233_), .Y(u5__abc_81276_new_n2284_));
AND2X2 AND2X2_5447 ( .A(u5__abc_81276_new_n415_), .B(u5__abc_81276_new_n2284_), .Y(u5__abc_81276_new_n2285_));
AND2X2 AND2X2_5448 ( .A(u5__abc_81276_new_n401__bF_buf0), .B(u5__abc_81276_new_n2285_), .Y(u5__abc_81276_new_n2286_));
AND2X2 AND2X2_5449 ( .A(u5__abc_81276_new_n448__bF_buf2), .B(u5__abc_81276_new_n2286_), .Y(u5__abc_81276_new_n2287_));
AND2X2 AND2X2_545 ( .A(spec_req_cs_1_bF_buf1_), .B(u0_csc1_4_), .Y(u0__abc_76628_new_n2061_));
AND2X2 AND2X2_5450 ( .A(u5__abc_81276_new_n523__bF_buf0), .B(u5__abc_81276_new_n2287_), .Y(u5__abc_81276_new_n2288_));
AND2X2 AND2X2_5451 ( .A(u5__abc_81276_new_n2289_), .B(u5__abc_81276_new_n490__bF_buf10), .Y(u5__abc_81276_new_n2290_));
AND2X2 AND2X2_5452 ( .A(u5__abc_81276_new_n2295_), .B(u5__abc_81276_new_n2126_), .Y(u5__abc_81276_new_n2296_));
AND2X2 AND2X2_5453 ( .A(u5__abc_81276_new_n2296_), .B(u5__abc_81276_new_n1949_), .Y(u5__abc_81276_new_n2297_));
AND2X2 AND2X2_5454 ( .A(u5__abc_81276_new_n2297_), .B(u5__abc_81276_new_n1937_), .Y(u5__abc_81276_new_n2298_));
AND2X2 AND2X2_5455 ( .A(u5__abc_81276_new_n2299_), .B(u5_ap_en), .Y(u5__abc_81276_new_n2300_));
AND2X2 AND2X2_5456 ( .A(u5__abc_81276_new_n1232_), .B(u5__abc_81276_new_n1343_), .Y(u5__abc_81276_new_n2302_));
AND2X2 AND2X2_5457 ( .A(u5__abc_81276_new_n1226_), .B(u5__abc_81276_new_n2302_), .Y(u5__abc_81276_new_n2303_));
AND2X2 AND2X2_5458 ( .A(u5__abc_81276_new_n2303_), .B(u5__abc_81276_new_n1565_), .Y(u5__abc_81276_new_n2304_));
AND2X2 AND2X2_5459 ( .A(u5__abc_81276_new_n2304_), .B(u5__abc_81276_new_n1598_), .Y(u5__abc_81276_new_n2305_));
AND2X2 AND2X2_546 ( .A(u0__abc_76628_new_n1946__bF_buf3), .B(u0__abc_76628_new_n2064_), .Y(u0__abc_76628_new_n2065_));
AND2X2 AND2X2_5460 ( .A(u5__abc_81276_new_n1748_), .B(u5__abc_81276_new_n2305_), .Y(u5__abc_81276_new_n2306_));
AND2X2 AND2X2_5461 ( .A(u5__abc_81276_new_n1791_), .B(u5__abc_81276_new_n2306_), .Y(u5__abc_81276_new_n2307_));
AND2X2 AND2X2_5462 ( .A(u5__abc_81276_new_n2309_), .B(u5__abc_81276_new_n1607_), .Y(u5__abc_81276_new_n2310_));
AND2X2 AND2X2_5463 ( .A(u5__abc_81276_new_n2309_), .B(u5__abc_81276_new_n1606_), .Y(u5__abc_81276_new_n2312_));
AND2X2 AND2X2_5464 ( .A(u5__abc_81276_new_n2309_), .B(u5__abc_81276_new_n1605_), .Y(u5__abc_81276_new_n2314_));
AND2X2 AND2X2_5465 ( .A(u5__abc_81276_new_n2313_), .B(u5__abc_81276_new_n2315_), .Y(u5__abc_81276_new_n2316_));
AND2X2 AND2X2_5466 ( .A(u5__abc_81276_new_n2316_), .B(u5__abc_81276_new_n2311_), .Y(u5__abc_81276_new_n2317_));
AND2X2 AND2X2_5467 ( .A(u5__abc_81276_new_n2317_), .B(u5__abc_81276_new_n1526__bF_buf3), .Y(u5__abc_81276_new_n2318_));
AND2X2 AND2X2_5468 ( .A(u5__abc_81276_new_n2318_), .B(1'h0), .Y(u5__abc_81276_new_n2319_));
AND2X2 AND2X2_5469 ( .A(u5__abc_81276_new_n1607_), .B(tms_s_0_), .Y(u5__abc_81276_new_n2321_));
AND2X2 AND2X2_547 ( .A(u0__abc_76628_new_n2063_), .B(u0__abc_76628_new_n2065_), .Y(u0__abc_76628_new_n2066_));
AND2X2 AND2X2_5470 ( .A(u5__abc_81276_new_n2314_), .B(u5__abc_81276_new_n2321_), .Y(u5__abc_81276_new_n2322_));
AND2X2 AND2X2_5471 ( .A(u5__abc_81276_new_n1608_), .B(tms_s_1_), .Y(u5__abc_81276_new_n2326_));
AND2X2 AND2X2_5472 ( .A(u5__abc_81276_new_n2309_), .B(u5__abc_81276_new_n2326_), .Y(u5__abc_81276_new_n2327_));
AND2X2 AND2X2_5473 ( .A(u5__abc_81276_new_n2325_), .B(u5__abc_81276_new_n2328_), .Y(u5__abc_81276_new_n2329_));
AND2X2 AND2X2_5474 ( .A(u5__abc_81276_new_n2329_), .B(u5__abc_81276_new_n2324_), .Y(u5__abc_81276_new_n2330_));
AND2X2 AND2X2_5475 ( .A(dv), .B(u5__abc_81276_new_n1637_), .Y(u5__abc_81276_new_n2332_));
AND2X2 AND2X2_5476 ( .A(u5__abc_81276_new_n1862_), .B(u1_wr_cycle), .Y(u5__abc_81276_new_n2333_));
AND2X2 AND2X2_5477 ( .A(u5__abc_81276_new_n2334_), .B(u5__abc_81276_new_n369_), .Y(u5__abc_81276_new_n2335_));
AND2X2 AND2X2_5478 ( .A(u5__abc_81276_new_n2336_), .B(u5_burst_cnt_0_), .Y(u5__abc_81276_new_n2337_));
AND2X2 AND2X2_5479 ( .A(u5__abc_81276_new_n2338_), .B(u5__abc_81276_new_n2299_), .Y(u5__abc_81276_new_n2339_));
AND2X2 AND2X2_548 ( .A(u0__abc_76628_new_n1947__bF_buf3), .B(sp_csc_5_), .Y(u0__abc_76628_new_n2068_));
AND2X2 AND2X2_5480 ( .A(u5__abc_81276_new_n2340_), .B(u5__abc_81276_new_n2308_), .Y(u5__0burst_cnt_10_0__0_));
AND2X2 AND2X2_5481 ( .A(u5__abc_81276_new_n2342_), .B(u5_burst_cnt_1_), .Y(u5__abc_81276_new_n2343_));
AND2X2 AND2X2_5482 ( .A(u5__abc_81276_new_n2334_), .B(u5__abc_81276_new_n370_), .Y(u5__abc_81276_new_n2344_));
AND2X2 AND2X2_5483 ( .A(u5__abc_81276_new_n2317_), .B(1'h0), .Y(u5__abc_81276_new_n2347_));
AND2X2 AND2X2_5484 ( .A(u5__abc_81276_new_n2348_), .B(u5__abc_81276_new_n2308_), .Y(u5__abc_81276_new_n2349_));
AND2X2 AND2X2_5485 ( .A(u5__abc_81276_new_n2346_), .B(u5__abc_81276_new_n2349_), .Y(u5__0burst_cnt_10_0__1_));
AND2X2 AND2X2_5486 ( .A(u5__abc_81276_new_n2334_), .B(u5__abc_81276_new_n371_), .Y(u5__abc_81276_new_n2351_));
AND2X2 AND2X2_5487 ( .A(u5__abc_81276_new_n2352_), .B(u5_burst_cnt_2_), .Y(u5__abc_81276_new_n2353_));
AND2X2 AND2X2_5488 ( .A(u5__abc_81276_new_n2354_), .B(u5__abc_81276_new_n2320_), .Y(u5__abc_81276_new_n2355_));
AND2X2 AND2X2_5489 ( .A(u5__abc_81276_new_n2318_), .B(1'h0), .Y(u5__abc_81276_new_n2356_));
AND2X2 AND2X2_549 ( .A(spec_req_cs_5_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n2069_));
AND2X2 AND2X2_5490 ( .A(u5__abc_81276_new_n2327_), .B(u5__abc_81276_new_n1526__bF_buf0), .Y(u5__abc_81276_new_n2357_));
AND2X2 AND2X2_5491 ( .A(u5__abc_81276_new_n2361_), .B(u5_burst_cnt_3_), .Y(u5__abc_81276_new_n2362_));
AND2X2 AND2X2_5492 ( .A(u5__abc_81276_new_n2334_), .B(u5__abc_81276_new_n372_), .Y(u5__abc_81276_new_n2363_));
AND2X2 AND2X2_5493 ( .A(u5__abc_81276_new_n2316_), .B(u5__abc_81276_new_n2366_), .Y(u5__abc_81276_new_n2367_));
AND2X2 AND2X2_5494 ( .A(u5__abc_81276_new_n2368_), .B(u5__abc_81276_new_n2308_), .Y(u5__abc_81276_new_n2369_));
AND2X2 AND2X2_5495 ( .A(u5__abc_81276_new_n2365_), .B(u5__abc_81276_new_n2369_), .Y(u5__0burst_cnt_10_0__3_));
AND2X2 AND2X2_5496 ( .A(u5__abc_81276_new_n2317_), .B(1'h0), .Y(u5__abc_81276_new_n2371_));
AND2X2 AND2X2_5497 ( .A(u5__abc_81276_new_n2373_), .B(u5_burst_cnt_4_), .Y(u5__abc_81276_new_n2374_));
AND2X2 AND2X2_5498 ( .A(u5__abc_81276_new_n2363_), .B(u5__abc_81276_new_n374_), .Y(u5__abc_81276_new_n2375_));
AND2X2 AND2X2_5499 ( .A(u5__abc_81276_new_n2377_), .B(u5__abc_81276_new_n2372_), .Y(u5__abc_81276_new_n2378_));
AND2X2 AND2X2_55 ( .A(wb_stb_i_bF_buf5), .B(wb_cyc_i), .Y(_abc_85006_new_n484_));
AND2X2 AND2X2_550 ( .A(u0__abc_76628_new_n2071_), .B(u0__abc_76628_new_n1179__bF_buf3), .Y(u0__abc_76628_new_n2072_));
AND2X2 AND2X2_5500 ( .A(u5__abc_81276_new_n2378_), .B(u5__abc_81276_new_n2308_), .Y(u5__0burst_cnt_10_0__4_));
AND2X2 AND2X2_5501 ( .A(u5__abc_81276_new_n2375_), .B(u5__abc_81276_new_n373_), .Y(u5__abc_81276_new_n2380_));
AND2X2 AND2X2_5502 ( .A(u5__abc_81276_new_n2381_), .B(u5_burst_cnt_5_), .Y(u5__abc_81276_new_n2382_));
AND2X2 AND2X2_5503 ( .A(u5__abc_81276_new_n2317_), .B(1'h0), .Y(u5__abc_81276_new_n2385_));
AND2X2 AND2X2_5504 ( .A(u5__abc_81276_new_n2386_), .B(u5__abc_81276_new_n2308_), .Y(u5__abc_81276_new_n2387_));
AND2X2 AND2X2_5505 ( .A(u5__abc_81276_new_n2384_), .B(u5__abc_81276_new_n2387_), .Y(u5__0burst_cnt_10_0__5_));
AND2X2 AND2X2_5506 ( .A(u5__abc_81276_new_n2389_), .B(u5_burst_cnt_6_), .Y(u5__abc_81276_new_n2390_));
AND2X2 AND2X2_5507 ( .A(u5__abc_81276_new_n2380_), .B(u5__abc_81276_new_n377_), .Y(u5__abc_81276_new_n2391_));
AND2X2 AND2X2_5508 ( .A(u5__abc_81276_new_n2317_), .B(1'h0), .Y(u5__abc_81276_new_n2394_));
AND2X2 AND2X2_5509 ( .A(u5__abc_81276_new_n2395_), .B(u5__abc_81276_new_n2308_), .Y(u5__abc_81276_new_n2396_));
AND2X2 AND2X2_551 ( .A(u0__abc_76628_new_n2072_), .B(u0__abc_76628_new_n2070_), .Y(u0__abc_76628_new_n2073_));
AND2X2 AND2X2_5510 ( .A(u5__abc_81276_new_n2393_), .B(u5__abc_81276_new_n2396_), .Y(u5__0burst_cnt_10_0__6_));
AND2X2 AND2X2_5511 ( .A(u5__abc_81276_new_n372_), .B(u5__abc_81276_new_n375_), .Y(u5__abc_81276_new_n2398_));
AND2X2 AND2X2_5512 ( .A(u5__abc_81276_new_n2398_), .B(u5__abc_81276_new_n377_), .Y(u5__abc_81276_new_n2399_));
AND2X2 AND2X2_5513 ( .A(u5__abc_81276_new_n2402_), .B(u5__abc_81276_new_n2400_), .Y(u5__abc_81276_new_n2403_));
AND2X2 AND2X2_5514 ( .A(u5__abc_81276_new_n2404_), .B(u5__abc_81276_new_n2405_), .Y(u5__abc_81276_new_n2406_));
AND2X2 AND2X2_5515 ( .A(u5__abc_81276_new_n2317_), .B(1'h0), .Y(u5__abc_81276_new_n2408_));
AND2X2 AND2X2_5516 ( .A(u5__abc_81276_new_n2409_), .B(u5__abc_81276_new_n2308_), .Y(u5__abc_81276_new_n2410_));
AND2X2 AND2X2_5517 ( .A(u5__abc_81276_new_n2407_), .B(u5__abc_81276_new_n2410_), .Y(u5__0burst_cnt_10_0__7_));
AND2X2 AND2X2_5518 ( .A(u5__abc_81276_new_n2363_), .B(u5__abc_81276_new_n379_), .Y(u5__abc_81276_new_n2412_));
AND2X2 AND2X2_5519 ( .A(u5__abc_81276_new_n2413_), .B(u5_burst_cnt_8_), .Y(u5__abc_81276_new_n2414_));
AND2X2 AND2X2_552 ( .A(u0__abc_76628_new_n2074_), .B(u0__abc_76628_new_n1175__bF_buf3), .Y(u0__abc_76628_new_n2075_));
AND2X2 AND2X2_5520 ( .A(u5__abc_81276_new_n2412_), .B(u5__abc_81276_new_n2415_), .Y(u5__abc_81276_new_n2416_));
AND2X2 AND2X2_5521 ( .A(u5__abc_81276_new_n2317_), .B(page_size_8_), .Y(u5__abc_81276_new_n2419_));
AND2X2 AND2X2_5522 ( .A(u5__abc_81276_new_n2420_), .B(u5__abc_81276_new_n2308_), .Y(u5__abc_81276_new_n2421_));
AND2X2 AND2X2_5523 ( .A(u5__abc_81276_new_n2418_), .B(u5__abc_81276_new_n2421_), .Y(u5__0burst_cnt_10_0__8_));
AND2X2 AND2X2_5524 ( .A(u5__abc_81276_new_n2423_), .B(u5_burst_cnt_9_), .Y(u5__abc_81276_new_n2424_));
AND2X2 AND2X2_5525 ( .A(u5__abc_81276_new_n2412_), .B(u5__abc_81276_new_n382_), .Y(u5__abc_81276_new_n2425_));
AND2X2 AND2X2_5526 ( .A(u5__abc_81276_new_n2317_), .B(page_size_9_), .Y(u5__abc_81276_new_n2428_));
AND2X2 AND2X2_5527 ( .A(u5__abc_81276_new_n2429_), .B(u5__abc_81276_new_n2308_), .Y(u5__abc_81276_new_n2430_));
AND2X2 AND2X2_5528 ( .A(u5__abc_81276_new_n2427_), .B(u5__abc_81276_new_n2430_), .Y(u5__0burst_cnt_10_0__9_));
AND2X2 AND2X2_5529 ( .A(u5__abc_81276_new_n372_), .B(u5__abc_81276_new_n379_), .Y(u5__abc_81276_new_n2432_));
AND2X2 AND2X2_553 ( .A(spec_req_cs_4_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n2076_));
AND2X2 AND2X2_5530 ( .A(u5__abc_81276_new_n2432_), .B(u5__abc_81276_new_n382_), .Y(u5__abc_81276_new_n2433_));
AND2X2 AND2X2_5531 ( .A(u5__abc_81276_new_n2436_), .B(u5__abc_81276_new_n2434_), .Y(u5__abc_81276_new_n2437_));
AND2X2 AND2X2_5532 ( .A(u5__abc_81276_new_n2438_), .B(u5__abc_81276_new_n2439_), .Y(u5__abc_81276_new_n2440_));
AND2X2 AND2X2_5533 ( .A(u5__abc_81276_new_n2317_), .B(page_size_10_), .Y(u5__abc_81276_new_n2442_));
AND2X2 AND2X2_5534 ( .A(u5__abc_81276_new_n2443_), .B(u5__abc_81276_new_n2308_), .Y(u5__abc_81276_new_n2444_));
AND2X2 AND2X2_5535 ( .A(u5__abc_81276_new_n2441_), .B(u5__abc_81276_new_n2444_), .Y(u5__0burst_cnt_10_0__10_));
AND2X2 AND2X2_5536 ( .A(u5__abc_81276_new_n1769_), .B(u5__abc_81276_new_n1519_), .Y(u5__abc_81276_new_n2446_));
AND2X2 AND2X2_5537 ( .A(u5__abc_81276_new_n625_), .B(u5__abc_81276_new_n1511_), .Y(u5__abc_81276_new_n2447_));
AND2X2 AND2X2_5538 ( .A(u5__abc_81276_new_n2446_), .B(u5__abc_81276_new_n2447_), .Y(u5__abc_81276_new_n2448_));
AND2X2 AND2X2_5539 ( .A(u5__abc_81276_new_n2448_), .B(u5__abc_81276_new_n1354_), .Y(u5__abc_81276_new_n2449_));
AND2X2 AND2X2_554 ( .A(u0__abc_76628_new_n2077_), .B(u0__abc_76628_new_n1174__bF_buf3), .Y(u0__abc_76628_new_n2078_));
AND2X2 AND2X2_5540 ( .A(u5__abc_81276_new_n2449_), .B(u5__abc_81276_new_n1357_), .Y(u5__abc_81276_new_n2450_));
AND2X2 AND2X2_5541 ( .A(u5__abc_81276_new_n1760_), .B(u5__abc_81276_new_n1361_), .Y(u5__abc_81276_new_n2451_));
AND2X2 AND2X2_5542 ( .A(u5__abc_81276_new_n1378_), .B(u5_cmd_asserted_bF_buf2), .Y(u5__abc_81276_new_n2452_));
AND2X2 AND2X2_5543 ( .A(u5__abc_81276_new_n2452_), .B(u5__abc_81276_new_n1364_), .Y(u5__abc_81276_new_n2453_));
AND2X2 AND2X2_5544 ( .A(u5__abc_81276_new_n2451_), .B(u5__abc_81276_new_n2453_), .Y(u5__abc_81276_new_n2454_));
AND2X2 AND2X2_5545 ( .A(u5__abc_81276_new_n2454_), .B(u5__abc_81276_new_n1759_), .Y(u5__abc_81276_new_n2455_));
AND2X2 AND2X2_5546 ( .A(u5__abc_81276_new_n2450_), .B(u5__abc_81276_new_n2455_), .Y(u5__abc_81276_new_n2456_));
AND2X2 AND2X2_5547 ( .A(u5__abc_81276_new_n1423_), .B(u5__abc_81276_new_n1480_), .Y(u5__abc_81276_new_n2457_));
AND2X2 AND2X2_5548 ( .A(u5__abc_81276_new_n2457_), .B(u5__abc_81276_new_n1415_), .Y(u5__abc_81276_new_n2458_));
AND2X2 AND2X2_5549 ( .A(u5__abc_81276_new_n1467_), .B(u5__abc_81276_new_n1793_), .Y(u5__abc_81276_new_n2459_));
AND2X2 AND2X2_555 ( .A(spec_req_cs_3_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n2079_));
AND2X2 AND2X2_5550 ( .A(u5__abc_81276_new_n2459_), .B(u5__abc_81276_new_n2458_), .Y(u5__abc_81276_new_n2460_));
AND2X2 AND2X2_5551 ( .A(u5__abc_81276_new_n2456_), .B(u5__abc_81276_new_n2460_), .Y(u5__abc_81276_new_n2461_));
AND2X2 AND2X2_5552 ( .A(u5__abc_81276_new_n1348_), .B(u5__abc_81276_new_n2461_), .Y(u5__abc_81276_new_n2462_));
AND2X2 AND2X2_5553 ( .A(u5__abc_81276_new_n2462_), .B(u5__abc_81276_new_n1117_), .Y(u5__abc_81276_new_n2463_));
AND2X2 AND2X2_5554 ( .A(u5__abc_81276_new_n2464_), .B(u5_ir_cnt_0_), .Y(u5__abc_81276_new_n2465_));
AND2X2 AND2X2_5555 ( .A(u5__abc_81276_new_n1348_), .B(u5__abc_81276_new_n1763_), .Y(u5__abc_81276_new_n2467_));
AND2X2 AND2X2_5556 ( .A(u5__abc_81276_new_n1353_), .B(u5__abc_81276_new_n1378_), .Y(u5__abc_81276_new_n2468_));
AND2X2 AND2X2_5557 ( .A(u5__abc_81276_new_n2468_), .B(u5__abc_81276_new_n1771_), .Y(u5__abc_81276_new_n2469_));
AND2X2 AND2X2_5558 ( .A(u5__abc_81276_new_n2469_), .B(u5__abc_81276_new_n2448_), .Y(u5__abc_81276_new_n2470_));
AND2X2 AND2X2_5559 ( .A(u5__abc_81276_new_n2460_), .B(u5__abc_81276_new_n2470_), .Y(u5__abc_81276_new_n2471_));
AND2X2 AND2X2_556 ( .A(u0__abc_76628_new_n2080_), .B(u0__abc_76628_new_n1173__bF_buf3), .Y(u0__abc_76628_new_n2081_));
AND2X2 AND2X2_5560 ( .A(u5__abc_81276_new_n2467_), .B(u5__abc_81276_new_n2471_), .Y(u5__abc_81276_new_n2472_));
AND2X2 AND2X2_5561 ( .A(u5__abc_81276_new_n2466_), .B(u5__abc_81276_new_n2473_), .Y(u5__0ir_cnt_3_0__0_));
AND2X2 AND2X2_5562 ( .A(u5__abc_81276_new_n2463_), .B(u5__abc_81276_new_n1116_), .Y(u5__abc_81276_new_n2475_));
AND2X2 AND2X2_5563 ( .A(u5__abc_81276_new_n2477_), .B(u5__abc_81276_new_n2473_), .Y(u5__abc_81276_new_n2478_));
AND2X2 AND2X2_5564 ( .A(u5__abc_81276_new_n2478_), .B(u5__abc_81276_new_n2476_), .Y(u5__abc_81276_new_n2479_));
AND2X2 AND2X2_5565 ( .A(u5__abc_81276_new_n2476_), .B(u5_ir_cnt_2_), .Y(u5__abc_81276_new_n2481_));
AND2X2 AND2X2_5566 ( .A(u5__abc_81276_new_n2475_), .B(u5__abc_81276_new_n1120_), .Y(u5__abc_81276_new_n2482_));
AND2X2 AND2X2_5567 ( .A(u5__abc_81276_new_n2483_), .B(u5__abc_81276_new_n2473_), .Y(u5__0ir_cnt_3_0__2_));
AND2X2 AND2X2_5568 ( .A(u5__abc_81276_new_n2482_), .B(u5_ir_cnt_3_), .Y(u5__abc_81276_new_n2485_));
AND2X2 AND2X2_5569 ( .A(u5__abc_81276_new_n2486_), .B(u5__abc_81276_new_n2487_), .Y(u5__abc_81276_new_n2488_));
AND2X2 AND2X2_557 ( .A(spec_req_cs_2_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n2082_));
AND2X2 AND2X2_5570 ( .A(u5__abc_81276_new_n2488_), .B(u5__abc_81276_new_n2473_), .Y(u5__0ir_cnt_3_0__3_));
AND2X2 AND2X2_5571 ( .A(u5__abc_81276_new_n1385_), .B(u5__abc_81276_new_n1508_), .Y(u5__abc_81276_new_n2490_));
AND2X2 AND2X2_5572 ( .A(u5__abc_81276_new_n612_), .B(u5__abc_81276_new_n1511_), .Y(u5__abc_81276_new_n2491_));
AND2X2 AND2X2_5573 ( .A(u5__abc_81276_new_n2491_), .B(u5__abc_81276_new_n1771_), .Y(u5__abc_81276_new_n2492_));
AND2X2 AND2X2_5574 ( .A(u5__abc_81276_new_n1762_), .B(u5__abc_81276_new_n2492_), .Y(u5__abc_81276_new_n2493_));
AND2X2 AND2X2_5575 ( .A(u5__abc_81276_new_n2493_), .B(u5__abc_81276_new_n2490_), .Y(u5__abc_81276_new_n2494_));
AND2X2 AND2X2_5576 ( .A(u5__abc_81276_new_n2446_), .B(u5__abc_81276_new_n1423_), .Y(u5__abc_81276_new_n2495_));
AND2X2 AND2X2_5577 ( .A(u5__abc_81276_new_n2495_), .B(u5__abc_81276_new_n1586_), .Y(u5__abc_81276_new_n2496_));
AND2X2 AND2X2_5578 ( .A(u5__abc_81276_new_n2496_), .B(u5__abc_81276_new_n1567_), .Y(u5__abc_81276_new_n2497_));
AND2X2 AND2X2_5579 ( .A(u5__abc_81276_new_n2497_), .B(u5__abc_81276_new_n1782_), .Y(u5__abc_81276_new_n2498_));
AND2X2 AND2X2_558 ( .A(u0__abc_76628_new_n2083_), .B(u0__abc_76628_new_n1172__bF_buf3), .Y(u0__abc_76628_new_n2084_));
AND2X2 AND2X2_5580 ( .A(u5__abc_81276_new_n2498_), .B(u5__abc_81276_new_n2494_), .Y(u5__abc_81276_new_n2499_));
AND2X2 AND2X2_5581 ( .A(u5__abc_81276_new_n1348_), .B(u5__abc_81276_new_n2499_), .Y(u5__abc_81276_new_n2500_));
AND2X2 AND2X2_5582 ( .A(u5__abc_81276_new_n1506_), .B(u5__abc_81276_new_n1699_), .Y(u5__abc_81276_new_n2502_));
AND2X2 AND2X2_5583 ( .A(u5__abc_81276_new_n1571_), .B(u5__abc_81276_new_n1378_), .Y(u5__abc_81276_new_n2503_));
AND2X2 AND2X2_5584 ( .A(u5__abc_81276_new_n1779_), .B(u5__abc_81276_new_n2503_), .Y(u5__abc_81276_new_n2504_));
AND2X2 AND2X2_5585 ( .A(u5__abc_81276_new_n2504_), .B(u5__abc_81276_new_n2502_), .Y(u5__abc_81276_new_n2505_));
AND2X2 AND2X2_5586 ( .A(u5__abc_81276_new_n2505_), .B(u5__abc_81276_new_n1788_), .Y(u5__abc_81276_new_n2506_));
AND2X2 AND2X2_5587 ( .A(u5__abc_81276_new_n1777_), .B(u5__abc_81276_new_n2506_), .Y(u5__abc_81276_new_n2507_));
AND2X2 AND2X2_5588 ( .A(u5__abc_81276_new_n2507_), .B(u5__abc_81276_new_n1348_), .Y(u5__abc_81276_new_n2508_));
AND2X2 AND2X2_5589 ( .A(u5__abc_81276_new_n1778_), .B(u5__abc_81276_new_n1378_), .Y(u5__abc_81276_new_n2510_));
AND2X2 AND2X2_559 ( .A(spec_req_cs_1_bF_buf0_), .B(u0_csc1_5_), .Y(u0__abc_76628_new_n2085_));
AND2X2 AND2X2_5590 ( .A(u5__abc_81276_new_n2510_), .B(u5__abc_81276_new_n1452_), .Y(u5__abc_81276_new_n2511_));
AND2X2 AND2X2_5591 ( .A(u5__abc_81276_new_n2511_), .B(u5__abc_81276_new_n1793_), .Y(u5__abc_81276_new_n2512_));
AND2X2 AND2X2_5592 ( .A(u5__abc_81276_new_n1788_), .B(u5__abc_81276_new_n2512_), .Y(u5__abc_81276_new_n2513_));
AND2X2 AND2X2_5593 ( .A(u5__abc_81276_new_n1777_), .B(u5__abc_81276_new_n2513_), .Y(u5__abc_81276_new_n2514_));
AND2X2 AND2X2_5594 ( .A(u5__abc_81276_new_n2514_), .B(u5__abc_81276_new_n1348_), .Y(u5__abc_81276_new_n2515_));
AND2X2 AND2X2_5595 ( .A(u5__abc_81276_new_n1801_), .B(u5__abc_81276_new_n1429_), .Y(u5__abc_81276_new_n2519_));
AND2X2 AND2X2_5596 ( .A(u5__abc_81276_new_n2519_), .B(u5__abc_81276_new_n2458_), .Y(u5__abc_81276_new_n2520_));
AND2X2 AND2X2_5597 ( .A(u5__abc_81276_new_n1242_), .B(u5__abc_81276_new_n2520_), .Y(u5__abc_81276_new_n2521_));
AND2X2 AND2X2_5598 ( .A(u5__abc_81276_new_n631_), .B(u5__abc_81276_new_n2446_), .Y(u5__abc_81276_new_n2522_));
AND2X2 AND2X2_5599 ( .A(u5__abc_81276_new_n1365_), .B(u5__abc_81276_new_n1772_), .Y(u5__abc_81276_new_n2523_));
AND2X2 AND2X2_56 ( .A(_abc_85006_new_n483_), .B(_abc_85006_new_n484_), .Y(not_mem_cyc));
AND2X2 AND2X2_560 ( .A(u0__abc_76628_new_n1946__bF_buf2), .B(u0__abc_76628_new_n2088_), .Y(u0__abc_76628_new_n2089_));
AND2X2 AND2X2_5600 ( .A(u5__abc_81276_new_n2522_), .B(u5__abc_81276_new_n2523_), .Y(u5__abc_81276_new_n2524_));
AND2X2 AND2X2_5601 ( .A(u5__abc_81276_new_n2459_), .B(u5__abc_81276_new_n2524_), .Y(u5__abc_81276_new_n2525_));
AND2X2 AND2X2_5602 ( .A(u5__abc_81276_new_n1347_), .B(u5__abc_81276_new_n2525_), .Y(u5__abc_81276_new_n2526_));
AND2X2 AND2X2_5603 ( .A(u5__abc_81276_new_n2521_), .B(u5__abc_81276_new_n2526_), .Y(u5__abc_81276_new_n2527_));
AND2X2 AND2X2_5604 ( .A(u5__abc_81276_new_n1383_), .B(u5__abc_81276_new_n1378_), .Y(u5__abc_81276_new_n2530_));
AND2X2 AND2X2_5605 ( .A(u5__abc_81276_new_n1758_), .B(u5__abc_81276_new_n2530_), .Y(u5__abc_81276_new_n2531_));
AND2X2 AND2X2_5606 ( .A(u5__abc_81276_new_n1762_), .B(u5__abc_81276_new_n2531_), .Y(u5__abc_81276_new_n2532_));
AND2X2 AND2X2_5607 ( .A(u5__abc_81276_new_n1776_), .B(u5__abc_81276_new_n2532_), .Y(u5__abc_81276_new_n2533_));
AND2X2 AND2X2_5608 ( .A(u5__abc_81276_new_n1480_), .B(u5__abc_81276_new_n1783_), .Y(u5__abc_81276_new_n2534_));
AND2X2 AND2X2_5609 ( .A(u5__abc_81276_new_n2534_), .B(u5__abc_81276_new_n1415_), .Y(u5__abc_81276_new_n2535_));
AND2X2 AND2X2_561 ( .A(u0__abc_76628_new_n2087_), .B(u0__abc_76628_new_n2089_), .Y(u0__abc_76628_new_n2090_));
AND2X2 AND2X2_5610 ( .A(u5__abc_81276_new_n2459_), .B(u5__abc_81276_new_n2535_), .Y(u5__abc_81276_new_n2536_));
AND2X2 AND2X2_5611 ( .A(u5__abc_81276_new_n2533_), .B(u5__abc_81276_new_n2536_), .Y(u5__abc_81276_new_n2537_));
AND2X2 AND2X2_5612 ( .A(u5__abc_81276_new_n1348_), .B(u5__abc_81276_new_n2537_), .Y(u5__abc_81276_new_n2538_));
AND2X2 AND2X2_5613 ( .A(u5__abc_81276_new_n2540_), .B(u5__abc_81276_new_n1102_), .Y(u5__abc_81276_new_n2541_));
AND2X2 AND2X2_5614 ( .A(u5_mc_le), .B(u5_timer_0_), .Y(u5__abc_81276_new_n2542_));
AND2X2 AND2X2_5615 ( .A(u5__abc_81276_new_n1801_), .B(u5__abc_81276_new_n1375_), .Y(u5__abc_81276_new_n2545_));
AND2X2 AND2X2_5616 ( .A(u5__abc_81276_new_n2450_), .B(u5__abc_81276_new_n2545_), .Y(u5__abc_81276_new_n2546_));
AND2X2 AND2X2_5617 ( .A(u5__abc_81276_new_n2546_), .B(u5__abc_81276_new_n2460_), .Y(u5__abc_81276_new_n2547_));
AND2X2 AND2X2_5618 ( .A(u5__abc_81276_new_n2547_), .B(u5__abc_81276_new_n1348_), .Y(u5__abc_81276_new_n2548_));
AND2X2 AND2X2_5619 ( .A(u5__abc_81276_new_n2528_), .B(u5__abc_81276_new_n2549_), .Y(u5__abc_81276_new_n2550_));
AND2X2 AND2X2_562 ( .A(u0__abc_76628_new_n1947__bF_buf2), .B(sp_csc_6_), .Y(u0__abc_76628_new_n2092_));
AND2X2 AND2X2_5620 ( .A(u5__abc_81276_new_n2529_), .B(u5__abc_81276_new_n2552_), .Y(u5__abc_81276_new_n2553_));
AND2X2 AND2X2_5621 ( .A(u5__abc_81276_new_n2554_), .B(u5__abc_81276_new_n2517_), .Y(u5__abc_81276_new_n2555_));
AND2X2 AND2X2_5622 ( .A(u5__abc_81276_new_n2556_), .B(u5__abc_81276_new_n2559_), .Y(u5__abc_81276_new_n2560_));
AND2X2 AND2X2_5623 ( .A(u5__abc_81276_new_n1907_), .B(u5__abc_81276_new_n1903_), .Y(u5__abc_81276_new_n2565_));
AND2X2 AND2X2_5624 ( .A(u5__abc_81276_new_n2565_), .B(u5__abc_81276_new_n1909_), .Y(u5__abc_81276_new_n2566_));
AND2X2 AND2X2_5625 ( .A(u5__abc_81276_new_n2566_), .B(u5__abc_81276_new_n947_), .Y(u5__abc_81276_new_n2567_));
AND2X2 AND2X2_5626 ( .A(u5__abc_81276_new_n1897_), .B(u5__abc_81276_new_n671_), .Y(u5__abc_81276_new_n2568_));
AND2X2 AND2X2_5627 ( .A(u5__abc_81276_new_n2568_), .B(u5__abc_81276_new_n2567_), .Y(u5__abc_81276_new_n2569_));
AND2X2 AND2X2_5628 ( .A(u5__abc_81276_new_n2564_), .B(u5__abc_81276_new_n2570_), .Y(u5__abc_81276_new_n2571_));
AND2X2 AND2X2_5629 ( .A(u5__abc_81276_new_n2561_), .B(u5__abc_81276_new_n2571_), .Y(u5__abc_81276_new_n2572_));
AND2X2 AND2X2_563 ( .A(spec_req_cs_5_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n2093_));
AND2X2 AND2X2_5630 ( .A(u5__abc_81276_new_n2562_), .B(u5__abc_81276_new_n2574_), .Y(u5__abc_81276_new_n2575_));
AND2X2 AND2X2_5631 ( .A(u5__abc_81276_new_n2576_), .B(u5__abc_81276_new_n2569_), .Y(u5__abc_81276_new_n2577_));
AND2X2 AND2X2_5632 ( .A(u5__abc_81276_new_n2577_), .B(u5__abc_81276_new_n2573_), .Y(u5__abc_81276_new_n2578_));
AND2X2 AND2X2_5633 ( .A(u5__abc_81276_new_n2580_), .B(u5__abc_81276_new_n1533_), .Y(u5__abc_81276_new_n2581_));
AND2X2 AND2X2_5634 ( .A(u5__abc_81276_new_n1920_), .B(u5__abc_81276_new_n2583_), .Y(u5__abc_81276_new_n2584_));
AND2X2 AND2X2_5635 ( .A(u5__abc_81276_new_n927_), .B(u5__abc_81276_new_n944_), .Y(u5__abc_81276_new_n2586_));
AND2X2 AND2X2_5636 ( .A(u5__abc_81276_new_n936_), .B(u5__abc_81276_new_n1018_), .Y(u5__abc_81276_new_n2587_));
AND2X2 AND2X2_5637 ( .A(u5__abc_81276_new_n906_), .B(u5__abc_81276_new_n890_), .Y(u5__abc_81276_new_n2588_));
AND2X2 AND2X2_5638 ( .A(u5__abc_81276_new_n899_), .B(u5__abc_81276_new_n916_), .Y(u5__abc_81276_new_n2589_));
AND2X2 AND2X2_5639 ( .A(u5__abc_81276_new_n2588_), .B(u5__abc_81276_new_n2589_), .Y(u5__abc_81276_new_n2590_));
AND2X2 AND2X2_564 ( .A(u0__abc_76628_new_n2095_), .B(u0__abc_76628_new_n1179__bF_buf2), .Y(u0__abc_76628_new_n2096_));
AND2X2 AND2X2_5640 ( .A(u5__abc_81276_new_n2590_), .B(u5__abc_81276_new_n2587_), .Y(u5__abc_81276_new_n2591_));
AND2X2 AND2X2_5641 ( .A(u5__abc_81276_new_n2591_), .B(u5__abc_81276_new_n2586_), .Y(u5__abc_81276_new_n2592_));
AND2X2 AND2X2_5642 ( .A(u5__abc_81276_new_n874_), .B(u5__abc_81276_new_n2592_), .Y(u5__abc_81276_new_n2593_));
AND2X2 AND2X2_5643 ( .A(u5__abc_81276_new_n671_), .B(u5__abc_81276_new_n2593_), .Y(u5__abc_81276_new_n2594_));
AND2X2 AND2X2_5644 ( .A(u5__abc_81276_new_n959_), .B(u5__abc_81276_new_n2596_), .Y(u5__abc_81276_new_n2597_));
AND2X2 AND2X2_5645 ( .A(u5__abc_81276_new_n2595_), .B(u5__abc_81276_new_n2597_), .Y(u5__abc_81276_new_n2598_));
AND2X2 AND2X2_5646 ( .A(u5__abc_81276_new_n1069_), .B(u5__abc_81276_new_n1879_), .Y(u5__abc_81276_new_n2599_));
AND2X2 AND2X2_5647 ( .A(u5__abc_81276_new_n2599_), .B(u5__abc_81276_new_n1085_), .Y(u5__abc_81276_new_n2600_));
AND2X2 AND2X2_5648 ( .A(u5__abc_81276_new_n2600_), .B(u5__abc_81276_new_n1053_), .Y(u5__abc_81276_new_n2601_));
AND2X2 AND2X2_5649 ( .A(u5__abc_81276_new_n995_), .B(u5__abc_81276_new_n1077_), .Y(u5__abc_81276_new_n2602_));
AND2X2 AND2X2_565 ( .A(u0__abc_76628_new_n2096_), .B(u0__abc_76628_new_n2094_), .Y(u0__abc_76628_new_n2097_));
AND2X2 AND2X2_5650 ( .A(u5__abc_81276_new_n951_), .B(u5__abc_81276_new_n1003_), .Y(u5__abc_81276_new_n2603_));
AND2X2 AND2X2_5651 ( .A(u5__abc_81276_new_n2602_), .B(u5__abc_81276_new_n2603_), .Y(u5__abc_81276_new_n2604_));
AND2X2 AND2X2_5652 ( .A(u5__abc_81276_new_n2601_), .B(u5__abc_81276_new_n2604_), .Y(u5__abc_81276_new_n2605_));
AND2X2 AND2X2_5653 ( .A(u5__abc_81276_new_n2605_), .B(u5__abc_81276_new_n2598_), .Y(u5__abc_81276_new_n2606_));
AND2X2 AND2X2_5654 ( .A(u5__abc_81276_new_n2606_), .B(u5__abc_81276_new_n804_), .Y(u5__abc_81276_new_n2607_));
AND2X2 AND2X2_5655 ( .A(u5__abc_81276_new_n2607_), .B(u5__abc_81276_new_n2594_), .Y(u5__abc_81276_new_n2608_));
AND2X2 AND2X2_5656 ( .A(u5__abc_81276_new_n2585_), .B(u5__abc_81276_new_n2608_), .Y(u5__abc_81276_new_n2609_));
AND2X2 AND2X2_5657 ( .A(u5__abc_81276_new_n2206_), .B(u5__abc_81276_new_n490__bF_buf9), .Y(u5__abc_81276_new_n2612_));
AND2X2 AND2X2_5658 ( .A(u5__abc_81276_new_n1268_), .B(u5__abc_81276_new_n1506_), .Y(u5__abc_81276_new_n2613_));
AND2X2 AND2X2_5659 ( .A(u5__abc_81276_new_n1290_), .B(u5__abc_81276_new_n2613_), .Y(u5__abc_81276_new_n2614_));
AND2X2 AND2X2_566 ( .A(u0__abc_76628_new_n2098_), .B(u0__abc_76628_new_n1175__bF_buf2), .Y(u0__abc_76628_new_n2099_));
AND2X2 AND2X2_5660 ( .A(u5__abc_81276_new_n1255_), .B(u5__abc_81276_new_n1331_), .Y(u5__abc_81276_new_n2615_));
AND2X2 AND2X2_5661 ( .A(u5__abc_81276_new_n1318_), .B(u5__abc_81276_new_n2615_), .Y(u5__abc_81276_new_n2616_));
AND2X2 AND2X2_5662 ( .A(u5__abc_81276_new_n2614_), .B(u5__abc_81276_new_n2616_), .Y(u5__abc_81276_new_n2617_));
AND2X2 AND2X2_5663 ( .A(u5__abc_81276_new_n951_), .B(u5__abc_81276_new_n995_), .Y(u5__abc_81276_new_n2618_));
AND2X2 AND2X2_5664 ( .A(u5__abc_81276_new_n1147_), .B(u5__abc_81276_new_n1171_), .Y(u5__abc_81276_new_n2619_));
AND2X2 AND2X2_5665 ( .A(u5__abc_81276_new_n1239_), .B(u5__abc_81276_new_n2619_), .Y(u5__abc_81276_new_n2620_));
AND2X2 AND2X2_5666 ( .A(u5__abc_81276_new_n2620_), .B(u5__abc_81276_new_n2618_), .Y(u5__abc_81276_new_n2621_));
AND2X2 AND2X2_5667 ( .A(u5__abc_81276_new_n1226_), .B(u5__abc_81276_new_n1344_), .Y(u5__abc_81276_new_n2622_));
AND2X2 AND2X2_5668 ( .A(u5__abc_81276_new_n1162_), .B(u5_tmr_done_bF_buf3), .Y(u5__abc_81276_new_n2623_));
AND2X2 AND2X2_5669 ( .A(u5__abc_81276_new_n1209_), .B(u5__abc_81276_new_n2623_), .Y(u5__abc_81276_new_n2624_));
AND2X2 AND2X2_567 ( .A(spec_req_cs_4_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n2100_));
AND2X2 AND2X2_5670 ( .A(u5__abc_81276_new_n2624_), .B(u5__abc_81276_new_n2622_), .Y(u5__abc_81276_new_n2625_));
AND2X2 AND2X2_5671 ( .A(u5__abc_81276_new_n2625_), .B(u5__abc_81276_new_n2621_), .Y(u5__abc_81276_new_n2626_));
AND2X2 AND2X2_5672 ( .A(u5__abc_81276_new_n2626_), .B(u5__abc_81276_new_n2617_), .Y(u5__abc_81276_new_n2627_));
AND2X2 AND2X2_5673 ( .A(u5__abc_81276_new_n1373_), .B(u5__abc_81276_new_n1364_), .Y(u5__abc_81276_new_n2628_));
AND2X2 AND2X2_5674 ( .A(u5__abc_81276_new_n2491_), .B(u5__abc_81276_new_n2628_), .Y(u5__abc_81276_new_n2629_));
AND2X2 AND2X2_5675 ( .A(u5__abc_81276_new_n1357_), .B(u5__abc_81276_new_n1352_), .Y(u5__abc_81276_new_n2630_));
AND2X2 AND2X2_5676 ( .A(u5__abc_81276_new_n2629_), .B(u5__abc_81276_new_n2630_), .Y(u5__abc_81276_new_n2631_));
AND2X2 AND2X2_5677 ( .A(u5__abc_81276_new_n2631_), .B(u5__abc_81276_new_n631_), .Y(u5__abc_81276_new_n2632_));
AND2X2 AND2X2_5678 ( .A(u5__abc_81276_new_n2632_), .B(u5__abc_81276_new_n1801_), .Y(u5__abc_81276_new_n2633_));
AND2X2 AND2X2_5679 ( .A(u5__abc_81276_new_n2633_), .B(u5__abc_81276_new_n2451_), .Y(u5__abc_81276_new_n2634_));
AND2X2 AND2X2_568 ( .A(u0__abc_76628_new_n2101_), .B(u0__abc_76628_new_n1174__bF_buf2), .Y(u0__abc_76628_new_n2102_));
AND2X2 AND2X2_5680 ( .A(u5__abc_81276_new_n2495_), .B(u5__abc_81276_new_n1415_), .Y(u5__abc_81276_new_n2635_));
AND2X2 AND2X2_5681 ( .A(u5__abc_81276_new_n1496_), .B(u5__abc_81276_new_n2635_), .Y(u5__abc_81276_new_n2636_));
AND2X2 AND2X2_5682 ( .A(u5__abc_81276_new_n2634_), .B(u5__abc_81276_new_n2636_), .Y(u5__abc_81276_new_n2637_));
AND2X2 AND2X2_5683 ( .A(u5__abc_81276_new_n2637_), .B(u5__abc_81276_new_n2627_), .Y(u5__abc_81276_new_n2638_));
AND2X2 AND2X2_5684 ( .A(u5__abc_81276_new_n1526__bF_buf1), .B(u5__abc_81276_new_n2583_), .Y(u5__abc_81276_new_n2641_));
AND2X2 AND2X2_5685 ( .A(u5__abc_81276_new_n2634_), .B(u5__abc_81276_new_n1789_), .Y(u5__abc_81276_new_n2643_));
AND2X2 AND2X2_5686 ( .A(u5__abc_81276_new_n1747_), .B(u5__abc_81276_new_n1598_), .Y(u5__abc_81276_new_n2644_));
AND2X2 AND2X2_5687 ( .A(u5__abc_81276_new_n951_), .B(u5__abc_81276_new_n1201_), .Y(u5__abc_81276_new_n2645_));
AND2X2 AND2X2_5688 ( .A(u5__abc_81276_new_n1172_), .B(u5__abc_81276_new_n2645_), .Y(u5__abc_81276_new_n2646_));
AND2X2 AND2X2_5689 ( .A(u5__abc_81276_new_n1133_), .B(u5__abc_81276_new_n1142_), .Y(u5__abc_81276_new_n2647_));
AND2X2 AND2X2_569 ( .A(spec_req_cs_3_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n2103_));
AND2X2 AND2X2_5690 ( .A(u5__abc_81276_new_n1162_), .B(u5__abc_81276_new_n2647_), .Y(u5__abc_81276_new_n2648_));
AND2X2 AND2X2_5691 ( .A(u5__abc_81276_new_n2304_), .B(u5__abc_81276_new_n2648_), .Y(u5__abc_81276_new_n2649_));
AND2X2 AND2X2_5692 ( .A(u5__abc_81276_new_n2649_), .B(u5__abc_81276_new_n2646_), .Y(u5__abc_81276_new_n2650_));
AND2X2 AND2X2_5693 ( .A(u5__abc_81276_new_n2650_), .B(u5__abc_81276_new_n2644_), .Y(u5__abc_81276_new_n2651_));
AND2X2 AND2X2_5694 ( .A(u5__abc_81276_new_n2643_), .B(u5__abc_81276_new_n2651_), .Y(u5__abc_81276_new_n2652_));
AND2X2 AND2X2_5695 ( .A(u5__abc_81276_new_n2642_), .B(u5__abc_81276_new_n2652_), .Y(u5__abc_81276_new_n2653_));
AND2X2 AND2X2_5696 ( .A(u5__abc_81276_new_n2655_), .B(u5__abc_81276_new_n2640_), .Y(u5__abc_81276_new_n2656_));
AND2X2 AND2X2_5697 ( .A(u5__abc_81276_new_n2611_), .B(u5__abc_81276_new_n2656_), .Y(u5__abc_81276_new_n2657_));
AND2X2 AND2X2_5698 ( .A(u5__abc_81276_new_n1526__bF_buf0), .B(u5__abc_81276_new_n2659_), .Y(u5__abc_81276_new_n2660_));
AND2X2 AND2X2_5699 ( .A(u5__abc_81276_new_n995_), .B(u5__abc_81276_new_n1201_), .Y(u5__abc_81276_new_n2662_));
AND2X2 AND2X2_57 ( .A(u0__abc_76628_new_n1100_), .B(u0_lmr_req0), .Y(u0__abc_76628_new_n1101_));
AND2X2 AND2X2_570 ( .A(u0__abc_76628_new_n2104_), .B(u0__abc_76628_new_n1173__bF_buf2), .Y(u0__abc_76628_new_n2105_));
AND2X2 AND2X2_5700 ( .A(u5__abc_81276_new_n1163_), .B(u5__abc_81276_new_n2662_), .Y(u5__abc_81276_new_n2663_));
AND2X2 AND2X2_5701 ( .A(u5__abc_81276_new_n2304_), .B(u5__abc_81276_new_n2663_), .Y(u5__abc_81276_new_n2664_));
AND2X2 AND2X2_5702 ( .A(u5__abc_81276_new_n2644_), .B(u5__abc_81276_new_n2664_), .Y(u5__abc_81276_new_n2665_));
AND2X2 AND2X2_5703 ( .A(u5__abc_81276_new_n2665_), .B(u5__abc_81276_new_n1134_), .Y(u5__abc_81276_new_n2666_));
AND2X2 AND2X2_5704 ( .A(u5__abc_81276_new_n2643_), .B(u5__abc_81276_new_n2666_), .Y(u5__abc_81276_new_n2667_));
AND2X2 AND2X2_5705 ( .A(u5__abc_81276_new_n2661_), .B(u5__abc_81276_new_n2667_), .Y(u5__abc_81276_new_n2668_));
AND2X2 AND2X2_5706 ( .A(u5__abc_81276_new_n2669_), .B(u5__abc_81276_new_n2639_), .Y(u5__abc_81276_new_n2670_));
AND2X2 AND2X2_5707 ( .A(u5__abc_81276_new_n2672_), .B(u5__abc_81276_new_n2675_), .Y(u5__0timer_7_0__0_));
AND2X2 AND2X2_5708 ( .A(u5__abc_81276_new_n2685_), .B(u5_timer_1_), .Y(u5__abc_81276_new_n2686_));
AND2X2 AND2X2_5709 ( .A(u5__abc_81276_new_n2541_), .B(u5__abc_81276_new_n1101_), .Y(u5__abc_81276_new_n2687_));
AND2X2 AND2X2_571 ( .A(spec_req_cs_2_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n2106_));
AND2X2 AND2X2_5710 ( .A(u5__abc_81276_new_n2550_), .B(u5__abc_81276_new_n2689_), .Y(u5__abc_81276_new_n2690_));
AND2X2 AND2X2_5711 ( .A(u5__abc_81276_new_n2684_), .B(u5__abc_81276_new_n2692_), .Y(u5__abc_81276_new_n2693_));
AND2X2 AND2X2_5712 ( .A(u5__abc_81276_new_n2694_), .B(u5__abc_81276_new_n2682_), .Y(u5__abc_81276_new_n2695_));
AND2X2 AND2X2_5713 ( .A(u5__abc_81276_new_n2696_), .B(u5__abc_81276_new_n2680_), .Y(u5__abc_81276_new_n2697_));
AND2X2 AND2X2_5714 ( .A(u5__abc_81276_new_n2700_), .B(u5__abc_81276_new_n2570_), .Y(u5__abc_81276_new_n2701_));
AND2X2 AND2X2_5715 ( .A(u5__abc_81276_new_n2698_), .B(u5__abc_81276_new_n2701_), .Y(u5__abc_81276_new_n2702_));
AND2X2 AND2X2_5716 ( .A(u5__abc_81276_new_n2703_), .B(u5__abc_81276_new_n2699_), .Y(u5__abc_81276_new_n2704_));
AND2X2 AND2X2_5717 ( .A(u5__abc_81276_new_n2705_), .B(u5__abc_81276_new_n2706_), .Y(u5__abc_81276_new_n2707_));
AND2X2 AND2X2_5718 ( .A(u5__abc_81276_new_n2711_), .B(u5__abc_81276_new_n2569_), .Y(u5__abc_81276_new_n2712_));
AND2X2 AND2X2_5719 ( .A(u5__abc_81276_new_n2712_), .B(u5__abc_81276_new_n2708_), .Y(u5__abc_81276_new_n2713_));
AND2X2 AND2X2_572 ( .A(u0__abc_76628_new_n2107_), .B(u0__abc_76628_new_n1172__bF_buf2), .Y(u0__abc_76628_new_n2108_));
AND2X2 AND2X2_5720 ( .A(u5__abc_81276_new_n2716_), .B(u5__abc_81276_new_n2640_), .Y(u5__abc_81276_new_n2717_));
AND2X2 AND2X2_5721 ( .A(u5__abc_81276_new_n2715_), .B(u5__abc_81276_new_n2717_), .Y(u5__abc_81276_new_n2718_));
AND2X2 AND2X2_5722 ( .A(u5__abc_81276_new_n2719_), .B(u5__abc_81276_new_n2639_), .Y(u5__abc_81276_new_n2720_));
AND2X2 AND2X2_5723 ( .A(u5__abc_81276_new_n2722_), .B(u5__abc_81276_new_n2678_), .Y(u5__0timer_7_0__1_));
AND2X2 AND2X2_5724 ( .A(u5__abc_81276_new_n2707_), .B(u5__abc_81276_new_n2575_), .Y(u5__abc_81276_new_n2726_));
AND2X2 AND2X2_5725 ( .A(u5__abc_81276_new_n2711_), .B(u5__abc_81276_new_n2705_), .Y(u5__abc_81276_new_n2730_));
AND2X2 AND2X2_5726 ( .A(u5__abc_81276_new_n2731_), .B(u5__abc_81276_new_n2569_), .Y(u5__abc_81276_new_n2732_));
AND2X2 AND2X2_5727 ( .A(u5__abc_81276_new_n2732_), .B(u5__abc_81276_new_n2728_), .Y(u5__abc_81276_new_n2733_));
AND2X2 AND2X2_5728 ( .A(u5__abc_81276_new_n1683_), .B(u5__abc_81276_new_n2508_), .Y(u5__abc_81276_new_n2734_));
AND2X2 AND2X2_5729 ( .A(u5__abc_81276_new_n2030_), .B(u5__abc_81276_new_n2054_), .Y(u5__abc_81276_new_n2736_));
AND2X2 AND2X2_573 ( .A(spec_req_cs_1_bF_buf5_), .B(u0_csc1_6_), .Y(u0__abc_76628_new_n2109_));
AND2X2 AND2X2_5730 ( .A(u5__abc_81276_new_n2043_), .B(u5__abc_81276_new_n2082_), .Y(u5__abc_81276_new_n2737_));
AND2X2 AND2X2_5731 ( .A(u5__abc_81276_new_n2736_), .B(u5__abc_81276_new_n2737_), .Y(u5__abc_81276_new_n2738_));
AND2X2 AND2X2_5732 ( .A(u5__abc_81276_new_n2122_), .B(u5__abc_81276_new_n1937_), .Y(u5__abc_81276_new_n2739_));
AND2X2 AND2X2_5733 ( .A(u5__abc_81276_new_n2095_), .B(u5__abc_81276_new_n2109_), .Y(u5__abc_81276_new_n2740_));
AND2X2 AND2X2_5734 ( .A(u5__abc_81276_new_n2740_), .B(u5__abc_81276_new_n2739_), .Y(u5__abc_81276_new_n2741_));
AND2X2 AND2X2_5735 ( .A(u5__abc_81276_new_n2738_), .B(u5__abc_81276_new_n2741_), .Y(u5__abc_81276_new_n2742_));
AND2X2 AND2X2_5736 ( .A(u5__abc_81276_new_n1959_), .B(u5__abc_81276_new_n490__bF_buf8), .Y(u5__abc_81276_new_n2743_));
AND2X2 AND2X2_5737 ( .A(u5__abc_81276_new_n1963_), .B(u5__abc_81276_new_n490__bF_buf7), .Y(u5__abc_81276_new_n2746_));
AND2X2 AND2X2_5738 ( .A(u5__abc_81276_new_n2748_), .B(u5__abc_81276_new_n1435_), .Y(u5__abc_81276_new_n2749_));
AND2X2 AND2X2_5739 ( .A(u5__abc_81276_new_n2749_), .B(u5__abc_81276_new_n2745_), .Y(u5__abc_81276_new_n2750_));
AND2X2 AND2X2_574 ( .A(u0__abc_76628_new_n1946__bF_buf1), .B(u0__abc_76628_new_n2112_), .Y(u0__abc_76628_new_n2113_));
AND2X2 AND2X2_5740 ( .A(u5__abc_81276_new_n1974_), .B(u5__abc_81276_new_n490__bF_buf6), .Y(u5__abc_81276_new_n2751_));
AND2X2 AND2X2_5741 ( .A(u5__abc_81276_new_n1987_), .B(u5__abc_81276_new_n490__bF_buf5), .Y(u5__abc_81276_new_n2753_));
AND2X2 AND2X2_5742 ( .A(u5__abc_81276_new_n2752_), .B(u5__abc_81276_new_n2754_), .Y(u5__abc_81276_new_n2755_));
AND2X2 AND2X2_5743 ( .A(u5__abc_81276_new_n2008_), .B(u5__abc_81276_new_n490__bF_buf4), .Y(u5__abc_81276_new_n2756_));
AND2X2 AND2X2_5744 ( .A(u5__abc_81276_new_n1996_), .B(u5__abc_81276_new_n490__bF_buf3), .Y(u5__abc_81276_new_n2758_));
AND2X2 AND2X2_5745 ( .A(u5__abc_81276_new_n2757_), .B(u5__abc_81276_new_n2759_), .Y(u5__abc_81276_new_n2760_));
AND2X2 AND2X2_5746 ( .A(u5__abc_81276_new_n2755_), .B(u5__abc_81276_new_n2760_), .Y(u5__abc_81276_new_n2761_));
AND2X2 AND2X2_5747 ( .A(u5__abc_81276_new_n474_), .B(u5__abc_81276_new_n1764_), .Y(u5__abc_81276_new_n2762_));
AND2X2 AND2X2_5748 ( .A(u5__abc_81276_new_n471_), .B(u5__abc_81276_new_n2762_), .Y(u5__abc_81276_new_n2763_));
AND2X2 AND2X2_5749 ( .A(u5__abc_81276_new_n464__bF_buf1), .B(u5__abc_81276_new_n2763_), .Y(u5__abc_81276_new_n2764_));
AND2X2 AND2X2_575 ( .A(u0__abc_76628_new_n2111_), .B(u0__abc_76628_new_n2113_), .Y(u0__abc_76628_new_n2114_));
AND2X2 AND2X2_5750 ( .A(u5__abc_81276_new_n522__bF_buf1), .B(u5__abc_81276_new_n2764_), .Y(u5__abc_81276_new_n2765_));
AND2X2 AND2X2_5751 ( .A(u5__abc_81276_new_n449__bF_buf6), .B(u5__abc_81276_new_n2765_), .Y(u5__abc_81276_new_n2766_));
AND2X2 AND2X2_5752 ( .A(u5__abc_81276_new_n2766_), .B(u5__abc_81276_new_n490__bF_buf2), .Y(u5__abc_81276_new_n2767_));
AND2X2 AND2X2_5753 ( .A(u5__abc_81276_new_n2064_), .B(u5__abc_81276_new_n490__bF_buf1), .Y(u5__abc_81276_new_n2768_));
AND2X2 AND2X2_5754 ( .A(u5__abc_81276_new_n2058_), .B(u5__abc_81276_new_n490__bF_buf0), .Y(u5__abc_81276_new_n2771_));
AND2X2 AND2X2_5755 ( .A(u5__abc_81276_new_n2012_), .B(u5__abc_81276_new_n490__bF_buf10), .Y(u5__abc_81276_new_n2773_));
AND2X2 AND2X2_5756 ( .A(u5__abc_81276_new_n2772_), .B(u5__abc_81276_new_n2774_), .Y(u5__abc_81276_new_n2775_));
AND2X2 AND2X2_5757 ( .A(u5__abc_81276_new_n2770_), .B(u5__abc_81276_new_n2775_), .Y(u5__abc_81276_new_n2776_));
AND2X2 AND2X2_5758 ( .A(u5__abc_81276_new_n2776_), .B(u5__abc_81276_new_n2761_), .Y(u5__abc_81276_new_n2777_));
AND2X2 AND2X2_5759 ( .A(u5__abc_81276_new_n2750_), .B(u5__abc_81276_new_n2777_), .Y(u5__abc_81276_new_n2778_));
AND2X2 AND2X2_576 ( .A(u0__abc_76628_new_n1947__bF_buf1), .B(sp_csc_7_), .Y(u0__abc_76628_new_n2116_));
AND2X2 AND2X2_5760 ( .A(u5__abc_81276_new_n2778_), .B(u5__abc_81276_new_n2742_), .Y(u5__abc_81276_new_n2779_));
AND2X2 AND2X2_5761 ( .A(u5__abc_81276_new_n2295_), .B(u5__abc_81276_new_n2779_), .Y(u5__abc_81276_new_n2780_));
AND2X2 AND2X2_5762 ( .A(u5__abc_81276_new_n2781_), .B(u5__abc_81276_new_n2780_), .Y(u5__abc_81276_new_n2782_));
AND2X2 AND2X2_5763 ( .A(u5__abc_81276_new_n2783_), .B(u5_timer_2_), .Y(u5__abc_81276_new_n2784_));
AND2X2 AND2X2_5764 ( .A(u5__abc_81276_new_n2687_), .B(u5__abc_81276_new_n1105_), .Y(u5__abc_81276_new_n2785_));
AND2X2 AND2X2_5765 ( .A(u5__abc_81276_new_n2550_), .B(u5__abc_81276_new_n2787_), .Y(u5__abc_81276_new_n2788_));
AND2X2 AND2X2_5766 ( .A(u5__abc_81276_new_n2558_), .B(u5__abc_81276_new_n2516_), .Y(u5__abc_81276_new_n2790_));
AND2X2 AND2X2_5767 ( .A(u5__abc_81276_new_n2789_), .B(u5__abc_81276_new_n2790_), .Y(u5__abc_81276_new_n2791_));
AND2X2 AND2X2_5768 ( .A(u5__abc_81276_new_n2793_), .B(u5__abc_81276_new_n2570_), .Y(u5__abc_81276_new_n2794_));
AND2X2 AND2X2_5769 ( .A(u5__abc_81276_new_n2792_), .B(u5__abc_81276_new_n2794_), .Y(u5__abc_81276_new_n2795_));
AND2X2 AND2X2_577 ( .A(spec_req_cs_5_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n2117_));
AND2X2 AND2X2_5770 ( .A(u5__abc_81276_new_n2797_), .B(u5__abc_81276_new_n2724_), .Y(u5__abc_81276_new_n2798_));
AND2X2 AND2X2_5771 ( .A(u5__abc_81276_new_n2798_), .B(u5__abc_81276_new_n2640_), .Y(u5__abc_81276_new_n2799_));
AND2X2 AND2X2_5772 ( .A(u5__abc_81276_new_n2800_), .B(u5__abc_81276_new_n2639_), .Y(u5__abc_81276_new_n2801_));
AND2X2 AND2X2_5773 ( .A(u5__abc_81276_new_n2803_), .B(u5__abc_81276_new_n2805_), .Y(u5__0timer_7_0__2_));
AND2X2 AND2X2_5774 ( .A(u5__abc_81276_new_n2727_), .B(u5__abc_81276_new_n2725_), .Y(u5__abc_81276_new_n2811_));
AND2X2 AND2X2_5775 ( .A(u5__abc_81276_new_n2810_), .B(u5__abc_81276_new_n2812_), .Y(u5__abc_81276_new_n2813_));
AND2X2 AND2X2_5776 ( .A(u5__abc_81276_new_n2813_), .B(u5__abc_81276_new_n2569_), .Y(u5__abc_81276_new_n2814_));
AND2X2 AND2X2_5777 ( .A(u5__abc_81276_new_n2808_), .B(u5__abc_81276_new_n2501_), .Y(u5__abc_81276_new_n2815_));
AND2X2 AND2X2_5778 ( .A(u5__abc_81276_new_n2816_), .B(u5__abc_81276_new_n2780_), .Y(u5__abc_81276_new_n2817_));
AND2X2 AND2X2_5779 ( .A(u5__abc_81276_new_n2540_), .B(u5__abc_81276_new_n1107_), .Y(u5__abc_81276_new_n2818_));
AND2X2 AND2X2_578 ( .A(u0__abc_76628_new_n2119_), .B(u0__abc_76628_new_n1179__bF_buf1), .Y(u0__abc_76628_new_n2120_));
AND2X2 AND2X2_5780 ( .A(u5__abc_81276_new_n2819_), .B(u5_timer_3_), .Y(u5__abc_81276_new_n2820_));
AND2X2 AND2X2_5781 ( .A(u5__abc_81276_new_n2690_), .B(u5__abc_81276_new_n2821_), .Y(u5__abc_81276_new_n2822_));
AND2X2 AND2X2_5782 ( .A(u5__abc_81276_new_n572_), .B(u5__abc_81276_new_n588_), .Y(u5__abc_81276_new_n2824_));
AND2X2 AND2X2_5783 ( .A(u5__abc_81276_new_n2824_), .B(u5__abc_81276_new_n604_), .Y(u5__abc_81276_new_n2825_));
AND2X2 AND2X2_5784 ( .A(u5__abc_81276_new_n555_), .B(u5__abc_81276_new_n564_), .Y(u5__abc_81276_new_n2826_));
AND2X2 AND2X2_5785 ( .A(u5__abc_81276_new_n2826_), .B(u5__abc_81276_new_n547_), .Y(u5__abc_81276_new_n2827_));
AND2X2 AND2X2_5786 ( .A(u5__abc_81276_new_n2827_), .B(u5__abc_81276_new_n639_), .Y(u5__abc_81276_new_n2828_));
AND2X2 AND2X2_5787 ( .A(u5__abc_81276_new_n2828_), .B(u5__abc_81276_new_n2825_), .Y(u5__abc_81276_new_n2829_));
AND2X2 AND2X2_5788 ( .A(u5__abc_81276_new_n625_), .B(u5__abc_81276_new_n882_), .Y(u5__abc_81276_new_n2830_));
AND2X2 AND2X2_5789 ( .A(u5__abc_81276_new_n666_), .B(u5__abc_81276_new_n647_), .Y(u5__abc_81276_new_n2831_));
AND2X2 AND2X2_579 ( .A(u0__abc_76628_new_n2120_), .B(u0__abc_76628_new_n2118_), .Y(u0__abc_76628_new_n2121_));
AND2X2 AND2X2_5790 ( .A(u5__abc_81276_new_n612_), .B(u5__abc_81276_new_n655_), .Y(u5__abc_81276_new_n2832_));
AND2X2 AND2X2_5791 ( .A(u5__abc_81276_new_n2831_), .B(u5__abc_81276_new_n2832_), .Y(u5__abc_81276_new_n2833_));
AND2X2 AND2X2_5792 ( .A(u5__abc_81276_new_n630_), .B(u5__abc_81276_new_n619_), .Y(u5__abc_81276_new_n2834_));
AND2X2 AND2X2_5793 ( .A(u5__abc_81276_new_n2833_), .B(u5__abc_81276_new_n2834_), .Y(u5__abc_81276_new_n2835_));
AND2X2 AND2X2_5794 ( .A(u5__abc_81276_new_n2835_), .B(u5__abc_81276_new_n2830_), .Y(u5__abc_81276_new_n2836_));
AND2X2 AND2X2_5795 ( .A(u5__abc_81276_new_n2836_), .B(u5__abc_81276_new_n2829_), .Y(u5__abc_81276_new_n2837_));
AND2X2 AND2X2_5796 ( .A(u5__abc_81276_new_n812_), .B(u5__abc_81276_new_n837_), .Y(u5__abc_81276_new_n2838_));
AND2X2 AND2X2_5797 ( .A(u5__abc_81276_new_n1909_), .B(u5__abc_81276_new_n1906_), .Y(u5__abc_81276_new_n2839_));
AND2X2 AND2X2_5798 ( .A(u5__abc_81276_new_n2839_), .B(u5__abc_81276_new_n580_), .Y(u5__abc_81276_new_n2840_));
AND2X2 AND2X2_5799 ( .A(u5__abc_81276_new_n2840_), .B(u5__abc_81276_new_n855_), .Y(u5__abc_81276_new_n2841_));
AND2X2 AND2X2_58 ( .A(u0_init_req0), .B(init_req), .Y(u0__abc_76628_new_n1102_));
AND2X2 AND2X2_580 ( .A(u0__abc_76628_new_n2122_), .B(u0__abc_76628_new_n1175__bF_buf1), .Y(u0__abc_76628_new_n2123_));
AND2X2 AND2X2_5800 ( .A(u5__abc_81276_new_n2841_), .B(u5__abc_81276_new_n2838_), .Y(u5__abc_81276_new_n2842_));
AND2X2 AND2X2_5801 ( .A(u5__abc_81276_new_n2837_), .B(u5__abc_81276_new_n2842_), .Y(u5__abc_81276_new_n2843_));
AND2X2 AND2X2_5802 ( .A(u5__abc_81276_new_n1897_), .B(u5__abc_81276_new_n2843_), .Y(u5__abc_81276_new_n2844_));
AND2X2 AND2X2_5803 ( .A(u5__abc_81276_new_n2844_), .B(u5__abc_81276_new_n2592_), .Y(u5__abc_81276_new_n2845_));
AND2X2 AND2X2_5804 ( .A(u5__abc_81276_new_n2846_), .B(u5__abc_81276_new_n2558_), .Y(u5__abc_81276_new_n2847_));
AND2X2 AND2X2_5805 ( .A(u5__abc_81276_new_n2847_), .B(u5__abc_81276_new_n2563_), .Y(u5__abc_81276_new_n2848_));
AND2X2 AND2X2_5806 ( .A(u5__abc_81276_new_n2823_), .B(u5__abc_81276_new_n2848_), .Y(u5__abc_81276_new_n2849_));
AND2X2 AND2X2_5807 ( .A(u5__abc_81276_new_n2850_), .B(u5__abc_81276_new_n2570_), .Y(u5__abc_81276_new_n2851_));
AND2X2 AND2X2_5808 ( .A(u5__abc_81276_new_n2855_), .B(u5__abc_81276_new_n2640_), .Y(u5__abc_81276_new_n2856_));
AND2X2 AND2X2_5809 ( .A(u5__abc_81276_new_n2853_), .B(u5__abc_81276_new_n2856_), .Y(u5__abc_81276_new_n2857_));
AND2X2 AND2X2_581 ( .A(spec_req_cs_4_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n2124_));
AND2X2 AND2X2_5810 ( .A(u5__abc_81276_new_n2858_), .B(u5__abc_81276_new_n2639_), .Y(u5__abc_81276_new_n2859_));
AND2X2 AND2X2_5811 ( .A(u5__abc_81276_new_n2861_), .B(u5__abc_81276_new_n2807_), .Y(u5__0timer_7_0__3_));
AND2X2 AND2X2_5812 ( .A(u5__abc_81276_new_n2673_), .B(u5__abc_81276_new_n2640_), .Y(u5__abc_81276_new_n2863_));
AND2X2 AND2X2_5813 ( .A(u5__abc_81276_new_n2635_), .B(u5__abc_81276_new_n1480_), .Y(u5__abc_81276_new_n2864_));
AND2X2 AND2X2_5814 ( .A(u5__abc_81276_new_n2864_), .B(u5__abc_81276_new_n1795_), .Y(u5__abc_81276_new_n2865_));
AND2X2 AND2X2_5815 ( .A(u5__abc_81276_new_n2634_), .B(u5__abc_81276_new_n1348_), .Y(u5__abc_81276_new_n2866_));
AND2X2 AND2X2_5816 ( .A(u5__abc_81276_new_n2866_), .B(u5__abc_81276_new_n2865_), .Y(u5__abc_81276_new_n2867_));
AND2X2 AND2X2_5817 ( .A(u5__abc_81276_new_n2528_), .B(u5__abc_81276_new_n2689_), .Y(u5__abc_81276_new_n2869_));
AND2X2 AND2X2_5818 ( .A(u5__abc_81276_new_n2869_), .B(u5__abc_81276_new_n2868_), .Y(u5__abc_81276_new_n2870_));
AND2X2 AND2X2_5819 ( .A(u5__abc_81276_new_n2870_), .B(u5__abc_81276_new_n2563_), .Y(u5__abc_81276_new_n2871_));
AND2X2 AND2X2_582 ( .A(u0__abc_76628_new_n2125_), .B(u0__abc_76628_new_n1174__bF_buf1), .Y(u0__abc_76628_new_n2126_));
AND2X2 AND2X2_5820 ( .A(u5__abc_81276_new_n2790_), .B(u5__abc_81276_new_n2549_), .Y(u5__abc_81276_new_n2872_));
AND2X2 AND2X2_5821 ( .A(u5__abc_81276_new_n2818_), .B(u5__abc_81276_new_n1109_), .Y(u5__abc_81276_new_n2873_));
AND2X2 AND2X2_5822 ( .A(u5__abc_81276_new_n2874_), .B(u5_timer_4_), .Y(u5__abc_81276_new_n2875_));
AND2X2 AND2X2_5823 ( .A(u5__abc_81276_new_n2654_), .B(u5__abc_81276_new_n2876_), .Y(u5__abc_81276_new_n2877_));
AND2X2 AND2X2_5824 ( .A(u5__abc_81276_new_n2877_), .B(u5__abc_81276_new_n2872_), .Y(u5__abc_81276_new_n2878_));
AND2X2 AND2X2_5825 ( .A(u5__abc_81276_new_n2878_), .B(u5__abc_81276_new_n2871_), .Y(u5__abc_81276_new_n2879_));
AND2X2 AND2X2_5826 ( .A(u5__abc_81276_new_n2509_), .B(u5__abc_81276_new_n2653_), .Y(u5__abc_81276_new_n2880_));
AND2X2 AND2X2_5827 ( .A(u5__abc_81276_new_n2881_), .B(u5__abc_81276_new_n2863_), .Y(u5__0timer_7_0__4_));
AND2X2 AND2X2_5828 ( .A(u5__abc_81276_new_n2873_), .B(u5__abc_81276_new_n1108_), .Y(u5__abc_81276_new_n2883_));
AND2X2 AND2X2_5829 ( .A(u5__abc_81276_new_n2884_), .B(u5_timer_5_), .Y(u5__abc_81276_new_n2885_));
AND2X2 AND2X2_583 ( .A(spec_req_cs_3_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n2127_));
AND2X2 AND2X2_5830 ( .A(u5__abc_81276_new_n2871_), .B(u5__abc_81276_new_n2872_), .Y(u5__abc_81276_new_n2887_));
AND2X2 AND2X2_5831 ( .A(u5__abc_81276_new_n2887_), .B(u5__abc_81276_new_n2886_), .Y(u5__abc_81276_new_n2888_));
AND2X2 AND2X2_5832 ( .A(u5__abc_81276_new_n2890_), .B(u5__abc_81276_new_n2863_), .Y(u5__abc_81276_new_n2891_));
AND2X2 AND2X2_5833 ( .A(u5__abc_81276_new_n2889_), .B(u5__abc_81276_new_n2891_), .Y(u5__0timer_7_0__5_));
AND2X2 AND2X2_5834 ( .A(u5__abc_81276_new_n2893_), .B(u5_timer_6_), .Y(u5__abc_81276_new_n2894_));
AND2X2 AND2X2_5835 ( .A(u5__abc_81276_new_n1108_), .B(u5__abc_81276_new_n1112_), .Y(u5__abc_81276_new_n2895_));
AND2X2 AND2X2_5836 ( .A(u5__abc_81276_new_n2873_), .B(u5__abc_81276_new_n2895_), .Y(u5__abc_81276_new_n2896_));
AND2X2 AND2X2_5837 ( .A(u5__abc_81276_new_n2887_), .B(u5__abc_81276_new_n2897_), .Y(u5__abc_81276_new_n2898_));
AND2X2 AND2X2_5838 ( .A(u5__abc_81276_new_n2901_), .B(u5__abc_81276_new_n2863_), .Y(u5__abc_81276_new_n2902_));
AND2X2 AND2X2_5839 ( .A(u5__abc_81276_new_n2899_), .B(u5__abc_81276_new_n2902_), .Y(u5__0timer_7_0__6_));
AND2X2 AND2X2_584 ( .A(u0__abc_76628_new_n2128_), .B(u0__abc_76628_new_n1173__bF_buf1), .Y(u0__abc_76628_new_n2129_));
AND2X2 AND2X2_5840 ( .A(u5__abc_81276_new_n2904_), .B(u5_timer_7_), .Y(u5__abc_81276_new_n2905_));
AND2X2 AND2X2_5841 ( .A(u5__abc_81276_new_n2887_), .B(u5__abc_81276_new_n2905_), .Y(u5__abc_81276_new_n2906_));
AND2X2 AND2X2_5842 ( .A(u5__abc_81276_new_n2909_), .B(u5__abc_81276_new_n2863_), .Y(u5__abc_81276_new_n2910_));
AND2X2 AND2X2_5843 ( .A(u5__abc_81276_new_n2907_), .B(u5__abc_81276_new_n2910_), .Y(u5__0timer_7_0__7_));
AND2X2 AND2X2_5844 ( .A(u5__abc_81276_new_n1526__bF_buf3), .B(u5__abc_81276_new_n1535_), .Y(u5__abc_81276_new_n2912_));
AND2X2 AND2X2_5845 ( .A(u5__abc_81276_new_n2703_), .B(u5__abc_81276_new_n2912_), .Y(u5__abc_81276_new_n2913_));
AND2X2 AND2X2_5846 ( .A(u5__abc_81276_new_n1242_), .B(u5__abc_81276_new_n1346_), .Y(u5__abc_81276_new_n2914_));
AND2X2 AND2X2_5847 ( .A(u5__abc_81276_new_n1271_), .B(u5__abc_81276_new_n1501_), .Y(u5__abc_81276_new_n2915_));
AND2X2 AND2X2_5848 ( .A(u5__abc_81276_new_n1289_), .B(u5__abc_81276_new_n2915_), .Y(u5__abc_81276_new_n2916_));
AND2X2 AND2X2_5849 ( .A(u5__abc_81276_new_n1269_), .B(u5__abc_81276_new_n2916_), .Y(u5__abc_81276_new_n2917_));
AND2X2 AND2X2_585 ( .A(spec_req_cs_2_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n2130_));
AND2X2 AND2X2_5850 ( .A(u5__abc_81276_new_n2914_), .B(u5__abc_81276_new_n2917_), .Y(u5__abc_81276_new_n2918_));
AND2X2 AND2X2_5851 ( .A(u5__abc_81276_new_n1791_), .B(u5__abc_81276_new_n2918_), .Y(u5__abc_81276_new_n2919_));
AND2X2 AND2X2_5852 ( .A(u5__abc_81276_new_n1744_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n2922_));
AND2X2 AND2X2_5853 ( .A(u5__abc_81276_new_n2922_), .B(u5__abc_81276_new_n1269_), .Y(u5__abc_81276_new_n2923_));
AND2X2 AND2X2_5854 ( .A(u5__abc_81276_new_n2914_), .B(u5__abc_81276_new_n2923_), .Y(u5__abc_81276_new_n2924_));
AND2X2 AND2X2_5855 ( .A(u5__abc_81276_new_n1791_), .B(u5__abc_81276_new_n2924_), .Y(u5__abc_81276_new_n2925_));
AND2X2 AND2X2_5856 ( .A(u5__abc_81276_new_n1744_), .B(u5__abc_81276_new_n1254_), .Y(u5__abc_81276_new_n2927_));
AND2X2 AND2X2_5857 ( .A(u5__abc_81276_new_n2927_), .B(u5__abc_81276_new_n1745_), .Y(u5__abc_81276_new_n2928_));
AND2X2 AND2X2_5858 ( .A(u5__abc_81276_new_n2914_), .B(u5__abc_81276_new_n2928_), .Y(u5__abc_81276_new_n2929_));
AND2X2 AND2X2_5859 ( .A(u5__abc_81276_new_n1791_), .B(u5__abc_81276_new_n2929_), .Y(u5__abc_81276_new_n2930_));
AND2X2 AND2X2_586 ( .A(u0__abc_76628_new_n2131_), .B(u0__abc_76628_new_n1172__bF_buf1), .Y(u0__abc_76628_new_n2132_));
AND2X2 AND2X2_5860 ( .A(u5__abc_81276_new_n2920_), .B(u5__abc_81276_new_n2931_), .Y(u5__abc_81276_new_n2932_));
AND2X2 AND2X2_5861 ( .A(u5__abc_81276_new_n2942_), .B(u5__abc_81276_new_n2934_), .Y(u5__abc_81276_new_n2943_));
AND2X2 AND2X2_5862 ( .A(u5__abc_81276_new_n1594_), .B(u5__abc_81276_new_n2448_), .Y(u5__abc_81276_new_n2944_));
AND2X2 AND2X2_5863 ( .A(u5__abc_81276_new_n1291_), .B(u5__abc_81276_new_n2944_), .Y(u5__abc_81276_new_n2945_));
AND2X2 AND2X2_5864 ( .A(u5__abc_81276_new_n2945_), .B(u5__abc_81276_new_n2459_), .Y(u5__abc_81276_new_n2946_));
AND2X2 AND2X2_5865 ( .A(u5__abc_81276_new_n2946_), .B(u5__abc_81276_new_n1377_), .Y(u5__abc_81276_new_n2947_));
AND2X2 AND2X2_5866 ( .A(u5__abc_81276_new_n2947_), .B(u5__abc_81276_new_n2521_), .Y(u5__abc_81276_new_n2948_));
AND2X2 AND2X2_5867 ( .A(u5__abc_81276_new_n2950_), .B(u5__abc_81276_new_n2926_), .Y(u5__abc_81276_new_n2951_));
AND2X2 AND2X2_5868 ( .A(u5__abc_81276_new_n2921_), .B(u5__abc_81276_new_n2951_), .Y(u5__abc_81276_new_n2952_));
AND2X2 AND2X2_5869 ( .A(u5__abc_81276_new_n1287_), .B(u5__abc_81276_new_n2953__bF_buf3), .Y(u5__abc_81276_new_n2954_));
AND2X2 AND2X2_587 ( .A(spec_req_cs_1_bF_buf4_), .B(u0_csc1_7_), .Y(u0__abc_76628_new_n2133_));
AND2X2 AND2X2_5870 ( .A(u5__abc_81276_new_n1255_), .B(u5__abc_81276_new_n1261_), .Y(u5__abc_81276_new_n2955_));
AND2X2 AND2X2_5871 ( .A(u5__abc_81276_new_n1290_), .B(u5__abc_81276_new_n1506_), .Y(u5__abc_81276_new_n2956_));
AND2X2 AND2X2_5872 ( .A(u5__abc_81276_new_n2956_), .B(u5__abc_81276_new_n2955_), .Y(u5__abc_81276_new_n2957_));
AND2X2 AND2X2_5873 ( .A(u5__abc_81276_new_n2957_), .B(u5__abc_81276_new_n1346_), .Y(u5__abc_81276_new_n2958_));
AND2X2 AND2X2_5874 ( .A(u5__abc_81276_new_n1242_), .B(u5__abc_81276_new_n2958_), .Y(u5__abc_81276_new_n2959_));
AND2X2 AND2X2_5875 ( .A(u5__abc_81276_new_n2637_), .B(u5__abc_81276_new_n2959_), .Y(u5__abc_81276_new_n2960_));
AND2X2 AND2X2_5876 ( .A(u5__abc_81276_new_n1526__bF_buf2), .B(u5__abc_81276_new_n2963_), .Y(u5__abc_81276_new_n2964_));
AND2X2 AND2X2_5877 ( .A(u5__abc_81276_new_n2643_), .B(u5__abc_81276_new_n2306_), .Y(u5__abc_81276_new_n2966_));
AND2X2 AND2X2_5878 ( .A(u5__abc_81276_new_n2965_), .B(u5__abc_81276_new_n2966_), .Y(u5__abc_81276_new_n2967_));
AND2X2 AND2X2_5879 ( .A(u5__abc_81276_new_n2971_), .B(u5__abc_81276_new_n2969_), .Y(u5__abc_81276_new_n2972_));
AND2X2 AND2X2_588 ( .A(u0__abc_76628_new_n1946__bF_buf0), .B(u0__abc_76628_new_n2136_), .Y(u0__abc_76628_new_n2137_));
AND2X2 AND2X2_5880 ( .A(u5__abc_81276_new_n2962_), .B(u5__abc_81276_new_n2972_), .Y(u5__abc_81276_new_n2973_));
AND2X2 AND2X2_5881 ( .A(u5__abc_81276_new_n2557_), .B(u5__abc_81276_new_n2912_), .Y(u5__abc_81276_new_n2975_));
AND2X2 AND2X2_5882 ( .A(u5__abc_81276_new_n1883_), .B(u5__abc_81276_new_n1895_), .Y(u5__abc_81276_new_n2976_));
AND2X2 AND2X2_5883 ( .A(u5__abc_81276_new_n2837_), .B(u5__abc_81276_new_n2593_), .Y(u5__abc_81276_new_n2977_));
AND2X2 AND2X2_5884 ( .A(u5__abc_81276_new_n713_), .B(u5__abc_81276_new_n728_), .Y(u5__abc_81276_new_n2978_));
AND2X2 AND2X2_5885 ( .A(u5__abc_81276_new_n1887_), .B(u5__abc_81276_new_n2978_), .Y(u5__abc_81276_new_n2979_));
AND2X2 AND2X2_5886 ( .A(u5__abc_81276_new_n580_), .B(u5__abc_81276_new_n2980_), .Y(u5__abc_81276_new_n2981_));
AND2X2 AND2X2_5887 ( .A(u5__abc_81276_new_n1884_), .B(u5__abc_81276_new_n2981_), .Y(u5__abc_81276_new_n2982_));
AND2X2 AND2X2_5888 ( .A(u5__abc_81276_new_n2982_), .B(u5__abc_81276_new_n695_), .Y(u5__abc_81276_new_n2983_));
AND2X2 AND2X2_5889 ( .A(u5__abc_81276_new_n2983_), .B(u5__abc_81276_new_n2979_), .Y(u5__abc_81276_new_n2984_));
AND2X2 AND2X2_589 ( .A(u0__abc_76628_new_n2135_), .B(u0__abc_76628_new_n2137_), .Y(u0__abc_76628_new_n2138_));
AND2X2 AND2X2_5890 ( .A(u5__abc_81276_new_n2977_), .B(u5__abc_81276_new_n2984_), .Y(u5__abc_81276_new_n2985_));
AND2X2 AND2X2_5891 ( .A(u5__abc_81276_new_n2985_), .B(u5__abc_81276_new_n2976_), .Y(u5__abc_81276_new_n2986_));
AND2X2 AND2X2_5892 ( .A(u5__abc_81276_new_n2313_), .B(u5__abc_81276_new_n2948_), .Y(u5__abc_81276_new_n2987_));
AND2X2 AND2X2_5893 ( .A(u5__abc_81276_new_n776_), .B(u5__abc_81276_new_n580_), .Y(u5__abc_81276_new_n2988_));
AND2X2 AND2X2_5894 ( .A(u5__abc_81276_new_n705_), .B(u5__abc_81276_new_n2988_), .Y(u5__abc_81276_new_n2989_));
AND2X2 AND2X2_5895 ( .A(u5__abc_81276_new_n2976_), .B(u5__abc_81276_new_n2989_), .Y(u5__abc_81276_new_n2990_));
AND2X2 AND2X2_5896 ( .A(u5__abc_81276_new_n2990_), .B(u5__abc_81276_new_n737_), .Y(u5__abc_81276_new_n2991_));
AND2X2 AND2X2_5897 ( .A(u5__abc_81276_new_n2991_), .B(u5__abc_81276_new_n2977_), .Y(u5__abc_81276_new_n2992_));
AND2X2 AND2X2_5898 ( .A(u5__abc_81276_new_n2839_), .B(u5__abc_81276_new_n754_), .Y(u5__abc_81276_new_n2993_));
AND2X2 AND2X2_5899 ( .A(u5__abc_81276_new_n619_), .B(u5__abc_81276_new_n890_), .Y(u5__abc_81276_new_n2994_));
AND2X2 AND2X2_59 ( .A(u0__abc_76628_new_n1104_), .B(u0_sreq_cs_le), .Y(u0__abc_76628_new_n1105_));
AND2X2 AND2X2_590 ( .A(u0__abc_76628_new_n1947__bF_buf0), .B(sp_csc_9_), .Y(u0__abc_76628_new_n2164_));
AND2X2 AND2X2_5900 ( .A(u5__abc_81276_new_n2830_), .B(u5__abc_81276_new_n2994_), .Y(u5__abc_81276_new_n2995_));
AND2X2 AND2X2_5901 ( .A(u5__abc_81276_new_n2995_), .B(u5__abc_81276_new_n2997_), .Y(u5__abc_81276_new_n2998_));
AND2X2 AND2X2_5902 ( .A(u5__abc_81276_new_n2993_), .B(u5__abc_81276_new_n2998_), .Y(u5__abc_81276_new_n2999_));
AND2X2 AND2X2_5903 ( .A(u5__abc_81276_new_n2999_), .B(u5__abc_81276_new_n1904_), .Y(u5__abc_81276_new_n3000_));
AND2X2 AND2X2_5904 ( .A(u5__abc_81276_new_n1883_), .B(u5__abc_81276_new_n3000_), .Y(u5__abc_81276_new_n3001_));
AND2X2 AND2X2_5905 ( .A(u5__abc_81276_new_n945_), .B(u5__abc_81276_new_n1905_), .Y(u5__abc_81276_new_n3002_));
AND2X2 AND2X2_5906 ( .A(u5__abc_81276_new_n906_), .B(u5__abc_81276_new_n927_), .Y(u5__abc_81276_new_n3003_));
AND2X2 AND2X2_5907 ( .A(u5__abc_81276_new_n3002_), .B(u5__abc_81276_new_n3003_), .Y(u5__abc_81276_new_n3004_));
AND2X2 AND2X2_5908 ( .A(u5__abc_81276_new_n3004_), .B(u5__abc_81276_new_n2589_), .Y(u5__abc_81276_new_n3005_));
AND2X2 AND2X2_5909 ( .A(u5__abc_81276_new_n3005_), .B(u5__abc_81276_new_n606_), .Y(u5__abc_81276_new_n3006_));
AND2X2 AND2X2_591 ( .A(spec_req_cs_5_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n2165_));
AND2X2 AND2X2_5910 ( .A(u5__abc_81276_new_n1889_), .B(u5__abc_81276_new_n1915_), .Y(u5__abc_81276_new_n3007_));
AND2X2 AND2X2_5911 ( .A(u5__abc_81276_new_n3006_), .B(u5__abc_81276_new_n3007_), .Y(u5__abc_81276_new_n3008_));
AND2X2 AND2X2_5912 ( .A(u5__abc_81276_new_n3001_), .B(u5__abc_81276_new_n3008_), .Y(u5__abc_81276_new_n3009_));
AND2X2 AND2X2_5913 ( .A(u5_timer2_1_), .B(u5_timer2_0_), .Y(u5__abc_81276_new_n3012_));
AND2X2 AND2X2_5914 ( .A(u5__abc_81276_new_n3010_), .B(u5__abc_81276_new_n3013_), .Y(u5__abc_81276_new_n3014_));
AND2X2 AND2X2_5915 ( .A(u5__abc_81276_new_n3014_), .B(u5__abc_81276_new_n2942_), .Y(u5__abc_81276_new_n3015_));
AND2X2 AND2X2_5916 ( .A(u5__abc_81276_new_n3017_), .B(u5__abc_81276_new_n3019_), .Y(u5__abc_81276_new_n3020_));
AND2X2 AND2X2_5917 ( .A(u5__abc_81276_new_n3023_), .B(u5__abc_81276_new_n2926_), .Y(u5__abc_81276_new_n3024_));
AND2X2 AND2X2_5918 ( .A(u5__abc_81276_new_n3021_), .B(u5__abc_81276_new_n3024_), .Y(u5__abc_81276_new_n3025_));
AND2X2 AND2X2_5919 ( .A(u5__abc_81276_new_n2703_), .B(u5__abc_81276_new_n2925_), .Y(u5__abc_81276_new_n3026_));
AND2X2 AND2X2_592 ( .A(u0__abc_76628_new_n2167_), .B(u0__abc_76628_new_n1179__bF_buf0), .Y(u0__abc_76628_new_n2168_));
AND2X2 AND2X2_5920 ( .A(u5__abc_81276_new_n2969_), .B(u5__abc_81276_new_n2970_), .Y(u5__abc_81276_new_n3029_));
AND2X2 AND2X2_5921 ( .A(u5__abc_81276_new_n2677_), .B(u5__abc_81276_new_n2969_), .Y(u5__abc_81276_new_n3030_));
AND2X2 AND2X2_5922 ( .A(u5__abc_81276_new_n3028_), .B(u5__abc_81276_new_n3031_), .Y(u5__abc_81276_new_n3032_));
AND2X2 AND2X2_5923 ( .A(u5__abc_81276_new_n2315_), .B(u5__abc_81276_new_n3009_), .Y(u5__abc_81276_new_n3038_));
AND2X2 AND2X2_5924 ( .A(u5__abc_81276_new_n2935_), .B(u5_timer2_2_), .Y(u5__abc_81276_new_n3040_));
AND2X2 AND2X2_5925 ( .A(u5__abc_81276_new_n3010_), .B(u5__abc_81276_new_n3041_), .Y(u5__abc_81276_new_n3042_));
AND2X2 AND2X2_5926 ( .A(u5__abc_81276_new_n3042_), .B(u5__abc_81276_new_n2942_), .Y(u5__abc_81276_new_n3043_));
AND2X2 AND2X2_5927 ( .A(u5__abc_81276_new_n3045_), .B(u5__abc_81276_new_n3037_), .Y(u5__abc_81276_new_n3046_));
AND2X2 AND2X2_5928 ( .A(u5__abc_81276_new_n3047_), .B(u5__abc_81276_new_n3036_), .Y(u5__abc_81276_new_n3048_));
AND2X2 AND2X2_5929 ( .A(u5__abc_81276_new_n3050_), .B(u5__abc_81276_new_n2970_), .Y(u5__abc_81276_new_n3051_));
AND2X2 AND2X2_593 ( .A(u0__abc_76628_new_n2168_), .B(u0__abc_76628_new_n2166_), .Y(u0__abc_76628_new_n2169_));
AND2X2 AND2X2_5930 ( .A(u5__abc_81276_new_n3049_), .B(u5__abc_81276_new_n3051_), .Y(u5__abc_81276_new_n3052_));
AND2X2 AND2X2_5931 ( .A(u5__abc_81276_new_n3053_), .B(u5__abc_81276_new_n3054_), .Y(u5__abc_81276_new_n3055_));
AND2X2 AND2X2_5932 ( .A(u5__abc_81276_new_n3056_), .B(u5__abc_81276_new_n3035_), .Y(u5__0timer2_8_0__2_));
AND2X2 AND2X2_5933 ( .A(u5__abc_81276_new_n1683_), .B(u5__abc_81276_new_n2912_), .Y(u5__abc_81276_new_n3058_));
AND2X2 AND2X2_5934 ( .A(u5__abc_81276_new_n2574_), .B(u5__abc_81276_new_n2969_), .Y(u5__abc_81276_new_n3059_));
AND2X2 AND2X2_5935 ( .A(u5__abc_81276_new_n2311_), .B(u5__abc_81276_new_n2948_), .Y(u5__abc_81276_new_n3061_));
AND2X2 AND2X2_5936 ( .A(u5__abc_81276_new_n2936_), .B(u5_timer2_3_), .Y(u5__abc_81276_new_n3063_));
AND2X2 AND2X2_5937 ( .A(u5__abc_81276_new_n3010_), .B(u5__abc_81276_new_n3064_), .Y(u5__abc_81276_new_n3065_));
AND2X2 AND2X2_5938 ( .A(u5__abc_81276_new_n3065_), .B(u5__abc_81276_new_n2942_), .Y(u5__abc_81276_new_n3066_));
AND2X2 AND2X2_5939 ( .A(u5__abc_81276_new_n3068_), .B(u5__abc_81276_new_n3069_), .Y(u5__abc_81276_new_n3070_));
AND2X2 AND2X2_594 ( .A(u0__abc_76628_new_n2170_), .B(u0__abc_76628_new_n1175__bF_buf0), .Y(u0__abc_76628_new_n2171_));
AND2X2 AND2X2_5940 ( .A(u5__abc_81276_new_n3072_), .B(u5__abc_81276_new_n2926_), .Y(u5__abc_81276_new_n3073_));
AND2X2 AND2X2_5941 ( .A(u5__abc_81276_new_n3071_), .B(u5__abc_81276_new_n3073_), .Y(u5__abc_81276_new_n3074_));
AND2X2 AND2X2_5942 ( .A(u5__abc_81276_new_n2679_), .B(u5__abc_81276_new_n2925_), .Y(u5__abc_81276_new_n3075_));
AND2X2 AND2X2_5943 ( .A(u5__abc_81276_new_n3077_), .B(u5__abc_81276_new_n3060_), .Y(u5__abc_81276_new_n3078_));
AND2X2 AND2X2_5944 ( .A(u5__abc_81276_new_n2562_), .B(u5__abc_81276_new_n2912_), .Y(u5__abc_81276_new_n3080_));
AND2X2 AND2X2_5945 ( .A(u5__abc_81276_new_n2854_), .B(u5__abc_81276_new_n3009_), .Y(u5__abc_81276_new_n3081_));
AND2X2 AND2X2_5946 ( .A(u5__abc_81276_new_n2937_), .B(u5_timer2_4_), .Y(u5__abc_81276_new_n3083_));
AND2X2 AND2X2_5947 ( .A(u5__abc_81276_new_n3010_), .B(u5__abc_81276_new_n3084_), .Y(u5__abc_81276_new_n3085_));
AND2X2 AND2X2_5948 ( .A(u5__abc_81276_new_n3085_), .B(u5__abc_81276_new_n2942_), .Y(u5__abc_81276_new_n3086_));
AND2X2 AND2X2_5949 ( .A(u5__abc_81276_new_n3088_), .B(u5__abc_81276_new_n3089_), .Y(u5__abc_81276_new_n3090_));
AND2X2 AND2X2_595 ( .A(spec_req_cs_4_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n2172_));
AND2X2 AND2X2_5950 ( .A(u5__abc_81276_new_n3092_), .B(u5__abc_81276_new_n2926_), .Y(u5__abc_81276_new_n3093_));
AND2X2 AND2X2_5951 ( .A(u5__abc_81276_new_n3091_), .B(u5__abc_81276_new_n3093_), .Y(u5__abc_81276_new_n3094_));
AND2X2 AND2X2_5952 ( .A(u5__abc_81276_new_n1683_), .B(u5__abc_81276_new_n2925_), .Y(u5__abc_81276_new_n3095_));
AND2X2 AND2X2_5953 ( .A(u5__abc_81276_new_n3096_), .B(u5__abc_81276_new_n3029_), .Y(u5__abc_81276_new_n3097_));
AND2X2 AND2X2_5954 ( .A(u5__abc_81276_new_n2699_), .B(u5__abc_81276_new_n2912_), .Y(u5__abc_81276_new_n3099_));
AND2X2 AND2X2_5955 ( .A(u5__abc_81276_new_n2938_), .B(u5_timer2_5_), .Y(u5__abc_81276_new_n3103_));
AND2X2 AND2X2_5956 ( .A(u5__abc_81276_new_n2942_), .B(u5__abc_81276_new_n3104_), .Y(u5__abc_81276_new_n3105_));
AND2X2 AND2X2_5957 ( .A(u5__abc_81276_new_n2931_), .B(u5__abc_81276_new_n3106_), .Y(u5__abc_81276_new_n3107_));
AND2X2 AND2X2_5958 ( .A(u5__abc_81276_new_n3101_), .B(u5__abc_81276_new_n3107_), .Y(u5__abc_81276_new_n3108_));
AND2X2 AND2X2_5959 ( .A(u5__abc_81276_new_n3029_), .B(u5__abc_81276_new_n2926_), .Y(u5__abc_81276_new_n3111_));
AND2X2 AND2X2_596 ( .A(u0__abc_76628_new_n2173_), .B(u0__abc_76628_new_n1174__bF_buf0), .Y(u0__abc_76628_new_n2174_));
AND2X2 AND2X2_5960 ( .A(u5__abc_81276_new_n3111_), .B(u5__abc_81276_new_n3110_), .Y(u5__abc_81276_new_n3112_));
AND2X2 AND2X2_5961 ( .A(u5__abc_81276_new_n3109_), .B(u5__abc_81276_new_n3112_), .Y(u5__abc_81276_new_n3113_));
AND2X2 AND2X2_5962 ( .A(u5__abc_81276_new_n2725_), .B(u5__abc_81276_new_n2912_), .Y(u5__abc_81276_new_n3115_));
AND2X2 AND2X2_5963 ( .A(u5__abc_81276_new_n2681_), .B(u5__abc_81276_new_n3009_), .Y(u5__abc_81276_new_n3116_));
AND2X2 AND2X2_5964 ( .A(u5__abc_81276_new_n2939_), .B(u5_timer2_6_), .Y(u5__abc_81276_new_n3118_));
AND2X2 AND2X2_5965 ( .A(u5__abc_81276_new_n2942_), .B(u5__abc_81276_new_n3119_), .Y(u5__abc_81276_new_n3120_));
AND2X2 AND2X2_5966 ( .A(u5__abc_81276_new_n3010_), .B(u5__abc_81276_new_n3120_), .Y(u5__abc_81276_new_n3121_));
AND2X2 AND2X2_5967 ( .A(u5__abc_81276_new_n3111_), .B(u5__abc_81276_new_n2932_), .Y(u5__abc_81276_new_n3123_));
AND2X2 AND2X2_5968 ( .A(u5__abc_81276_new_n3123_), .B(u5__abc_81276_new_n3122_), .Y(u5__abc_81276_new_n3124_));
AND2X2 AND2X2_5969 ( .A(u5__abc_81276_new_n2808_), .B(u5__abc_81276_new_n2912_), .Y(u5__abc_81276_new_n3126_));
AND2X2 AND2X2_597 ( .A(spec_req_cs_3_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n2175_));
AND2X2 AND2X2_5970 ( .A(u5__abc_81276_new_n2900_), .B(u5__abc_81276_new_n3009_), .Y(u5__abc_81276_new_n3127_));
AND2X2 AND2X2_5971 ( .A(u5__abc_81276_new_n3128_), .B(u5_timer2_8_), .Y(u5__abc_81276_new_n3129_));
AND2X2 AND2X2_5972 ( .A(u5__abc_81276_new_n2940_), .B(u5_timer2_7_), .Y(u5__abc_81276_new_n3130_));
AND2X2 AND2X2_5973 ( .A(u5__abc_81276_new_n3010_), .B(u5__abc_81276_new_n3131_), .Y(u5__abc_81276_new_n3132_));
AND2X2 AND2X2_5974 ( .A(u5__abc_81276_new_n3123_), .B(u5__abc_81276_new_n3133_), .Y(u5__abc_81276_new_n3134_));
AND2X2 AND2X2_5975 ( .A(u5__abc_81276_new_n2518_), .B(u5__abc_81276_new_n2912_), .Y(u5__abc_81276_new_n3136_));
AND2X2 AND2X2_5976 ( .A(u5__abc_81276_new_n2908_), .B(u5__abc_81276_new_n3009_), .Y(u5__abc_81276_new_n3137_));
AND2X2 AND2X2_5977 ( .A(u5__abc_81276_new_n2941_), .B(u5_timer2_8_), .Y(u5__abc_81276_new_n3138_));
AND2X2 AND2X2_5978 ( .A(u5__abc_81276_new_n3010_), .B(u5__abc_81276_new_n3138_), .Y(u5__abc_81276_new_n3139_));
AND2X2 AND2X2_5979 ( .A(u5__abc_81276_new_n3123_), .B(u5__abc_81276_new_n3140_), .Y(u5__abc_81276_new_n3141_));
AND2X2 AND2X2_598 ( .A(u0__abc_76628_new_n2176_), .B(u0__abc_76628_new_n1173__bF_buf0), .Y(u0__abc_76628_new_n2177_));
AND2X2 AND2X2_5980 ( .A(dv), .B(u5__abc_81276_new_n1829_), .Y(u5__abc_81276_new_n3144_));
AND2X2 AND2X2_5981 ( .A(u5__abc_81276_new_n3151_), .B(u5__abc_81276_new_n3150_), .Y(u5__abc_81276_new_n3152_));
AND2X2 AND2X2_5982 ( .A(u5__abc_81276_new_n3152_), .B(u5__abc_81276_new_n3149_), .Y(u5__0ack_cnt_3_0__0_));
AND2X2 AND2X2_5983 ( .A(u5_ack_cnt_1_), .B(u5_ack_cnt_0_), .Y(u5__abc_81276_new_n3155_));
AND2X2 AND2X2_5984 ( .A(u5__abc_81276_new_n3154_), .B(u5__abc_81276_new_n3157_), .Y(u5__abc_81276_new_n3158_));
AND2X2 AND2X2_5985 ( .A(u5__abc_81276_new_n3144_), .B(u5__abc_81276_new_n3156_), .Y(u5__abc_81276_new_n3160_));
AND2X2 AND2X2_5986 ( .A(u5__abc_81276_new_n3161_), .B(u5__abc_81276_new_n3150_), .Y(u5__abc_81276_new_n3162_));
AND2X2 AND2X2_5987 ( .A(u5__abc_81276_new_n3159_), .B(u5__abc_81276_new_n3162_), .Y(u5__0ack_cnt_3_0__1_));
AND2X2 AND2X2_5988 ( .A(u5__abc_81276_new_n3146_), .B(u5__abc_81276_new_n1818_), .Y(u5__abc_81276_new_n3164_));
AND2X2 AND2X2_5989 ( .A(u5__abc_81276_new_n3144_), .B(u5__abc_81276_new_n3155_), .Y(u5__abc_81276_new_n3165_));
AND2X2 AND2X2_599 ( .A(spec_req_cs_2_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n2178_));
AND2X2 AND2X2_5990 ( .A(u5__abc_81276_new_n3169_), .B(u5__abc_81276_new_n3150_), .Y(u5__abc_81276_new_n3170_));
AND2X2 AND2X2_5991 ( .A(u5__abc_81276_new_n3170_), .B(u5__abc_81276_new_n3168_), .Y(u5__0ack_cnt_3_0__2_));
AND2X2 AND2X2_5992 ( .A(u5__abc_81276_new_n3173_), .B(u5_ack_cnt_3_), .Y(u5__abc_81276_new_n3174_));
AND2X2 AND2X2_5993 ( .A(u5__abc_81276_new_n3155_), .B(u5_ack_cnt_2_), .Y(u5__abc_81276_new_n3176_));
AND2X2 AND2X2_5994 ( .A(u5__abc_81276_new_n3176_), .B(u5__abc_81276_new_n1815_), .Y(u5__abc_81276_new_n3177_));
AND2X2 AND2X2_5995 ( .A(u5__abc_81276_new_n3178_), .B(u5__abc_81276_new_n3179_), .Y(u5__abc_81276_new_n3180_));
AND2X2 AND2X2_5996 ( .A(u5__abc_81276_new_n3144_), .B(u5__abc_81276_new_n3180_), .Y(u5__abc_81276_new_n3181_));
AND2X2 AND2X2_5997 ( .A(u5__abc_81276_new_n3182_), .B(u5__abc_81276_new_n3150_), .Y(u5__abc_81276_new_n3183_));
AND2X2 AND2X2_5998 ( .A(u5__abc_81276_new_n3175_), .B(u5__abc_81276_new_n3183_), .Y(u5__0ack_cnt_3_0__3_));
AND2X2 AND2X2_5999 ( .A(u5__abc_81276_new_n3186_), .B(u5__abc_81276_new_n3185_), .Y(u5__0cmd_asserted2_0_0_));
AND2X2 AND2X2_6 ( .A(_abc_85006_new_n254_), .B(_abc_85006_new_n255_), .Y(_abc_85006_new_n256_));
AND2X2 AND2X2_60 ( .A(u0__abc_76628_new_n1106_), .B(u0__abc_76628_new_n1107_), .Y(u0__0spec_req_cs_7_0__0_));
AND2X2 AND2X2_600 ( .A(u0__abc_76628_new_n2179_), .B(u0__abc_76628_new_n1172__bF_buf0), .Y(u0__abc_76628_new_n2180_));
AND2X2 AND2X2_6000 ( .A(u5_mc_le), .B(u5_cmd_asserted_bF_buf3), .Y(u5__abc_81276_new_n3188_));
AND2X2 AND2X2_6001 ( .A(u5_cmd_3_), .B(u5__0mc_le_0_0_), .Y(u5__abc_81276_new_n3189_));
AND2X2 AND2X2_6002 ( .A(u5__abc_81276_new_n3192_), .B(u5__abc_81276_new_n3191_), .Y(u5__0mc_adv_r_0_0_));
AND2X2 AND2X2_6003 ( .A(u5__abc_81276_new_n1879_), .B(u5__abc_81276_new_n1708_), .Y(u5__abc_81276_new_n3194_));
AND2X2 AND2X2_6004 ( .A(u5__abc_81276_new_n1232_), .B(u5__abc_81276_new_n1201_), .Y(u5__abc_81276_new_n3196_));
AND2X2 AND2X2_6005 ( .A(u5__abc_81276_new_n1194_), .B(u5__abc_81276_new_n3196_), .Y(u5__abc_81276_new_n3197_));
AND2X2 AND2X2_6006 ( .A(u5__abc_81276_new_n2622_), .B(u5__abc_81276_new_n3197_), .Y(u5__abc_81276_new_n3198_));
AND2X2 AND2X2_6007 ( .A(u5__abc_81276_new_n1174_), .B(u5__abc_81276_new_n3198_), .Y(u5__abc_81276_new_n3199_));
AND2X2 AND2X2_6008 ( .A(u5__abc_81276_new_n3199_), .B(u5__abc_81276_new_n2617_), .Y(u5__abc_81276_new_n3200_));
AND2X2 AND2X2_6009 ( .A(u5__abc_81276_new_n2637_), .B(u5__abc_81276_new_n3200_), .Y(u5__abc_81276_new_n3201_));
AND2X2 AND2X2_601 ( .A(spec_req_cs_1_bF_buf3_), .B(u0_csc1_9_), .Y(u0__abc_76628_new_n2181_));
AND2X2 AND2X2_6010 ( .A(u5__abc_81276_new_n3201_), .B(u5__abc_81276_new_n3195_), .Y(mc_adv_d));
AND2X2 AND2X2_6011 ( .A(u5_mc_le), .B(u5_mc_adv_r1), .Y(u5__abc_81276_new_n3203_));
AND2X2 AND2X2_6012 ( .A(mc_adv_d), .B(u5__0mc_le_0_0_), .Y(u5__abc_81276_new_n3204_));
AND2X2 AND2X2_6013 ( .A(u5__abc_81276_new_n3206_), .B(u5__abc_81276_new_n1712_), .Y(u5__abc_81276_new_n3207_));
AND2X2 AND2X2_6014 ( .A(u5__abc_81276_new_n3212_), .B(u5__abc_81276_new_n3210_), .Y(u5__abc_81276_new_n3213_));
AND2X2 AND2X2_6015 ( .A(u5__abc_81276_new_n3213_), .B(u5__abc_81276_new_n1559_), .Y(u5__abc_81276_new_n3214_));
AND2X2 AND2X2_6016 ( .A(u5__abc_81276_new_n1526__bF_buf1), .B(u5__abc_81276_new_n3214_), .Y(u5__abc_81276_new_n3215_));
AND2X2 AND2X2_6017 ( .A(u5__abc_81276_new_n3216_), .B(u5_state_0_), .Y(u5_next_state_0_));
AND2X2 AND2X2_6018 ( .A(u5__abc_81276_new_n3214_), .B(u5_state_1_), .Y(u5__abc_81276_new_n3218_));
AND2X2 AND2X2_6019 ( .A(u5_wb_cycle), .B(u5_wb_wait), .Y(u5__abc_81276_new_n3220_));
AND2X2 AND2X2_602 ( .A(u0__abc_76628_new_n1946__bF_buf3), .B(u0__abc_76628_new_n2184_), .Y(u0__abc_76628_new_n2185_));
AND2X2 AND2X2_6020 ( .A(u5__abc_81276_new_n3222_), .B(u5__abc_81276_new_n3219_), .Y(u5__abc_81276_new_n3223_));
AND2X2 AND2X2_6021 ( .A(u5__abc_81276_new_n989_), .B(u5__abc_81276_new_n3224_), .Y(u5__abc_81276_new_n3225_));
AND2X2 AND2X2_6022 ( .A(u5__abc_81276_new_n3206_), .B(u5__abc_81276_new_n3227_), .Y(u5__abc_81276_new_n3228_));
AND2X2 AND2X2_6023 ( .A(u5_kro), .B(u5_tmr_done_bF_buf1), .Y(u5__abc_81276_new_n3229_));
AND2X2 AND2X2_6024 ( .A(u5__abc_81276_new_n1586_), .B(u5_cmd_asserted_bF_buf2), .Y(u5__abc_81276_new_n3230_));
AND2X2 AND2X2_6025 ( .A(u5__abc_81276_new_n3231_), .B(u5_state_1_), .Y(u5__abc_81276_new_n3232_));
AND2X2 AND2X2_6026 ( .A(u5__abc_81276_new_n624_), .B(u5__abc_81276_new_n3233_), .Y(u5__abc_81276_new_n3234_));
AND2X2 AND2X2_6027 ( .A(u5__abc_81276_new_n3239_), .B(u5__abc_81276_new_n3238_), .Y(u5__abc_81276_new_n3240_));
AND2X2 AND2X2_6028 ( .A(u5__abc_81276_new_n1612_), .B(u3_wb_read_go), .Y(u5__abc_81276_new_n3243_));
AND2X2 AND2X2_6029 ( .A(u5__abc_81276_new_n3245_), .B(u5__abc_81276_new_n3242_), .Y(u5__abc_81276_new_n3246_));
AND2X2 AND2X2_603 ( .A(u0__abc_76628_new_n2183_), .B(u0__abc_76628_new_n2185_), .Y(u0__abc_76628_new_n2186_));
AND2X2 AND2X2_6030 ( .A(u5__abc_81276_new_n3246_), .B(u5__abc_81276_new_n3241_), .Y(u5__abc_81276_new_n3247_));
AND2X2 AND2X2_6031 ( .A(u5__abc_81276_new_n1610_), .B(u5__abc_81276_new_n1552_), .Y(u5__abc_81276_new_n3249_));
AND2X2 AND2X2_6032 ( .A(u5__abc_81276_new_n3252_), .B(u5__abc_81276_new_n1464_), .Y(u5__abc_81276_new_n3253_));
AND2X2 AND2X2_6033 ( .A(u5__abc_81276_new_n3251_), .B(u5__abc_81276_new_n3253_), .Y(u5__abc_81276_new_n3254_));
AND2X2 AND2X2_6034 ( .A(u5__abc_81276_new_n1412_), .B(u5__abc_81276_new_n2953__bF_buf2), .Y(u5__abc_81276_new_n3255_));
AND2X2 AND2X2_6035 ( .A(u5__abc_81276_new_n3256_), .B(u5_state_2_), .Y(u5__abc_81276_new_n3257_));
AND2X2 AND2X2_6036 ( .A(u5__abc_81276_new_n3259_), .B(u5__abc_81276_new_n3258_), .Y(u5__abc_81276_new_n3260_));
AND2X2 AND2X2_6037 ( .A(u5__abc_81276_new_n1428_), .B(u5__abc_81276_new_n3261_), .Y(u5__abc_81276_new_n3262_));
AND2X2 AND2X2_6038 ( .A(u5__abc_81276_new_n1821_), .B(u5__abc_81276_new_n1123_), .Y(u5__abc_81276_new_n3265_));
AND2X2 AND2X2_6039 ( .A(u5__abc_81276_new_n3266_), .B(u5__abc_81276_new_n1825_), .Y(u5__abc_81276_new_n3267_));
AND2X2 AND2X2_604 ( .A(u0__abc_76628_new_n1947__bF_buf3), .B(sp_csc_10_), .Y(u0__abc_76628_new_n2188_));
AND2X2 AND2X2_6040 ( .A(u5__abc_81276_new_n1585_), .B(u5__abc_81276_new_n3238_), .Y(u5__abc_81276_new_n3269_));
AND2X2 AND2X2_6041 ( .A(u5__abc_81276_new_n3266_), .B(u5__abc_81276_new_n3269_), .Y(u5__abc_81276_new_n3270_));
AND2X2 AND2X2_6042 ( .A(u5__abc_81276_new_n1405_), .B(u5__abc_81276_new_n3271_), .Y(u5__abc_81276_new_n3272_));
AND2X2 AND2X2_6043 ( .A(u5__abc_81276_new_n3272_), .B(u5__abc_81276_new_n3268_), .Y(u5__abc_81276_new_n3273_));
AND2X2 AND2X2_6044 ( .A(u5__abc_81276_new_n624_), .B(u5__abc_81276_new_n3275_), .Y(u5__abc_81276_new_n3276_));
AND2X2 AND2X2_6045 ( .A(u5__abc_81276_new_n3276_), .B(u5__abc_81276_new_n3274_), .Y(u5__abc_81276_new_n3277_));
AND2X2 AND2X2_6046 ( .A(u5__abc_81276_new_n3239_), .B(u5_wb_cycle), .Y(u5__abc_81276_new_n3282_));
AND2X2 AND2X2_6047 ( .A(u5__abc_81276_new_n1123_), .B(u5_ap_en), .Y(u5__abc_81276_new_n3284_));
AND2X2 AND2X2_6048 ( .A(u5__abc_81276_new_n3283_), .B(u5__abc_81276_new_n3284_), .Y(u5__abc_81276_new_n3285_));
AND2X2 AND2X2_6049 ( .A(u5__abc_81276_new_n1443_), .B(u5__abc_81276_new_n3258_), .Y(u5__abc_81276_new_n3288_));
AND2X2 AND2X2_605 ( .A(spec_req_cs_5_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n2189_));
AND2X2 AND2X2_6050 ( .A(u5__abc_81276_new_n3287_), .B(u5__abc_81276_new_n3288_), .Y(u5__abc_81276_new_n3289_));
AND2X2 AND2X2_6051 ( .A(u5__abc_81276_new_n3214_), .B(u5_state_3_), .Y(u5__abc_81276_new_n3292_));
AND2X2 AND2X2_6052 ( .A(u5__abc_81276_new_n1526__bF_buf0), .B(u5__abc_81276_new_n3292_), .Y(u5__abc_81276_new_n3293_));
AND2X2 AND2X2_6053 ( .A(u5__abc_81276_new_n3294_), .B(u5_state_3_), .Y(u5__abc_81276_new_n3295_));
AND2X2 AND2X2_6054 ( .A(u5__abc_81276_new_n1160_), .B(u5__abc_81276_new_n3295_), .Y(u5__abc_81276_new_n3296_));
AND2X2 AND2X2_6055 ( .A(u5__abc_81276_new_n1555_), .B(u5__abc_81276_new_n1556_), .Y(u5__abc_81276_new_n3299_));
AND2X2 AND2X2_6056 ( .A(u5__abc_81276_new_n3209_), .B(u5_state_4_), .Y(u5__abc_81276_new_n3300_));
AND2X2 AND2X2_6057 ( .A(u5__abc_81276_new_n3301_), .B(u5__abc_81276_new_n3299_), .Y(u5__abc_81276_new_n3302_));
AND2X2 AND2X2_6058 ( .A(u5__abc_81276_new_n1536_), .B(u5_lookup_ready2), .Y(u5__abc_81276_new_n3305_));
AND2X2 AND2X2_6059 ( .A(u5_kro), .B(bank_open), .Y(u5__abc_81276_new_n3306_));
AND2X2 AND2X2_606 ( .A(u0__abc_76628_new_n2191_), .B(u0__abc_76628_new_n1179__bF_buf5), .Y(u0__abc_76628_new_n2192_));
AND2X2 AND2X2_6060 ( .A(u5__abc_81276_new_n3305_), .B(u5__abc_81276_new_n3306_), .Y(u5__abc_81276_new_n3307_));
AND2X2 AND2X2_6061 ( .A(u5__abc_81276_new_n3307_), .B(u5__abc_81276_new_n3304_), .Y(u5__abc_81276_new_n3308_));
AND2X2 AND2X2_6062 ( .A(u5__abc_81276_new_n3303_), .B(u5__abc_81276_new_n3308_), .Y(u5__abc_81276_new_n3309_));
AND2X2 AND2X2_6063 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_4_), .Y(u5__abc_81276_new_n3310_));
AND2X2 AND2X2_6064 ( .A(u5__abc_81276_new_n3311_), .B(u5__abc_81276_new_n3302_), .Y(u5__abc_81276_new_n3312_));
AND2X2 AND2X2_6065 ( .A(u5__abc_81276_new_n1526__bF_buf3), .B(u5__abc_81276_new_n3313_), .Y(u5__abc_81276_new_n3314_));
AND2X2 AND2X2_6066 ( .A(u5__abc_81276_new_n694_), .B(u5__abc_81276_new_n2953__bF_buf0), .Y(u5__abc_81276_new_n3315_));
AND2X2 AND2X2_6067 ( .A(u5__abc_81276_new_n1504_), .B(u5__abc_81276_new_n1712_), .Y(u5__abc_81276_new_n3317_));
AND2X2 AND2X2_6068 ( .A(u5__abc_81276_new_n3318_), .B(u5_state_5_), .Y(u5__abc_81276_new_n3319_));
AND2X2 AND2X2_6069 ( .A(u5__abc_81276_new_n1500_), .B(u5__abc_81276_new_n3320_), .Y(u5__abc_81276_new_n3321_));
AND2X2 AND2X2_607 ( .A(u0__abc_76628_new_n2192_), .B(u0__abc_76628_new_n2190_), .Y(u0__abc_76628_new_n2193_));
AND2X2 AND2X2_6070 ( .A(u5__abc_81276_new_n1920_), .B(u5__abc_81276_new_n1558_), .Y(u5__abc_81276_new_n3323_));
AND2X2 AND2X2_6071 ( .A(u5__abc_81276_new_n3210_), .B(u5__abc_81276_new_n1555_), .Y(u5__abc_81276_new_n3324_));
AND2X2 AND2X2_6072 ( .A(u5__abc_81276_new_n1728_), .B(u5__abc_81276_new_n1536_), .Y(u5__abc_81276_new_n3325_));
AND2X2 AND2X2_6073 ( .A(u5__abc_81276_new_n3326_), .B(u5__abc_81276_new_n3327_), .Y(u5__abc_81276_new_n3328_));
AND2X2 AND2X2_6074 ( .A(u5__abc_81276_new_n3303_), .B(u5__abc_81276_new_n3305_), .Y(u5__abc_81276_new_n3330_));
AND2X2 AND2X2_6075 ( .A(u5__abc_81276_new_n3330_), .B(u5__abc_81276_new_n1549_), .Y(u5__abc_81276_new_n3331_));
AND2X2 AND2X2_6076 ( .A(u5__abc_81276_new_n3332_), .B(u5__abc_81276_new_n3329_), .Y(u5__abc_81276_new_n3333_));
AND2X2 AND2X2_6077 ( .A(u5__abc_81276_new_n3333_), .B(u5__abc_81276_new_n3324_), .Y(u5__abc_81276_new_n3334_));
AND2X2 AND2X2_6078 ( .A(u5__abc_81276_new_n3323__bF_buf3), .B(u5__abc_81276_new_n3334_), .Y(u5__abc_81276_new_n3335_));
AND2X2 AND2X2_6079 ( .A(u5_tmr_done_bF_buf0), .B(rfr_ack), .Y(u5__abc_81276_new_n3336_));
AND2X2 AND2X2_608 ( .A(u0__abc_76628_new_n2194_), .B(u0__abc_76628_new_n1175__bF_buf5), .Y(u0__abc_76628_new_n2195_));
AND2X2 AND2X2_6080 ( .A(u5__abc_81276_new_n3337_), .B(u5__abc_81276_new_n3338_), .Y(u5__abc_81276_new_n3339_));
AND2X2 AND2X2_6081 ( .A(u5__abc_81276_new_n1928_), .B(u5__abc_81276_new_n3339_), .Y(u5__abc_81276_new_n3340_));
AND2X2 AND2X2_6082 ( .A(u5__abc_81276_new_n2119_), .B(u5__abc_81276_new_n490__bF_buf9), .Y(u5__abc_81276_new_n3341_));
AND2X2 AND2X2_6083 ( .A(u5__abc_81276_new_n2953__bF_buf3), .B(u5_state_6_), .Y(u5__abc_81276_new_n3342_));
AND2X2 AND2X2_6084 ( .A(u5__abc_81276_new_n3341_), .B(u5__abc_81276_new_n3342_), .Y(u5__abc_81276_new_n3343_));
AND2X2 AND2X2_6085 ( .A(u5__abc_81276_new_n3212_), .B(u5__abc_81276_new_n1555_), .Y(u5__abc_81276_new_n3346_));
AND2X2 AND2X2_6086 ( .A(u5__abc_81276_new_n3346_), .B(u5__abc_81276_new_n3210_), .Y(u5__abc_81276_new_n3347_));
AND2X2 AND2X2_6087 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_7_), .Y(u5__abc_81276_new_n3348_));
AND2X2 AND2X2_6088 ( .A(u5__abc_81276_new_n3323__bF_buf2), .B(u5__abc_81276_new_n3348_), .Y(u5__abc_81276_new_n3349_));
AND2X2 AND2X2_6089 ( .A(u5__abc_81276_new_n3341_), .B(u5__abc_81276_new_n3350_), .Y(u5__abc_81276_new_n3351_));
AND2X2 AND2X2_609 ( .A(spec_req_cs_4_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n2196_));
AND2X2 AND2X2_6090 ( .A(u5__abc_81276_new_n2114_), .B(u5__abc_81276_new_n490__bF_buf8), .Y(u5__abc_81276_new_n3352_));
AND2X2 AND2X2_6091 ( .A(u5__abc_81276_new_n1699_), .B(u5_tmr_done_bF_buf2), .Y(u5__abc_81276_new_n3354_));
AND2X2 AND2X2_6092 ( .A(u5__abc_81276_new_n3355_), .B(u5__abc_81276_new_n3353_), .Y(u5__abc_81276_new_n3356_));
AND2X2 AND2X2_6093 ( .A(u5__abc_81276_new_n3356_), .B(u5_state_7_), .Y(u5__abc_81276_new_n3357_));
AND2X2 AND2X2_6094 ( .A(u5__abc_81276_new_n3352_), .B(u5__abc_81276_new_n3357_), .Y(u5__abc_81276_new_n3358_));
AND2X2 AND2X2_6095 ( .A(u5__abc_81276_new_n3323__bF_buf1), .B(u5__abc_81276_new_n3324_), .Y(u5__abc_81276_new_n3361_));
AND2X2 AND2X2_6096 ( .A(u5__abc_81276_new_n3362_), .B(u5_state_8_), .Y(u5__abc_81276_new_n3363_));
AND2X2 AND2X2_6097 ( .A(u5__abc_81276_new_n3307_), .B(row_same), .Y(u5__abc_81276_new_n3364_));
AND2X2 AND2X2_6098 ( .A(u5__abc_81276_new_n3365_), .B(u5__abc_81276_new_n3303_), .Y(u5__abc_81276_new_n3366_));
AND2X2 AND2X2_6099 ( .A(u5_state_8_), .B(u5_wb_wait), .Y(u5__abc_81276_new_n3367_));
AND2X2 AND2X2_61 ( .A(u0__abc_76628_new_n1109_), .B(spec_req_cs_1_bF_buf4_), .Y(u0__abc_76628_new_n1110_));
AND2X2 AND2X2_610 ( .A(u0__abc_76628_new_n2197_), .B(u0__abc_76628_new_n1174__bF_buf5), .Y(u0__abc_76628_new_n2198_));
AND2X2 AND2X2_6100 ( .A(u5__abc_81276_new_n1728_), .B(u5__abc_81276_new_n3367_), .Y(u5__abc_81276_new_n3368_));
AND2X2 AND2X2_6101 ( .A(u5__abc_81276_new_n3370_), .B(u5__abc_81276_new_n3371_), .Y(u5__abc_81276_new_n3372_));
AND2X2 AND2X2_6102 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3372_), .Y(u5__abc_81276_new_n3373_));
AND2X2 AND2X2_6103 ( .A(u5__abc_81276_new_n1536_), .B(u5_kro), .Y(u5__abc_81276_new_n3374_));
AND2X2 AND2X2_6104 ( .A(u5_state_8_), .B(u5_wb_wait_r), .Y(u5__abc_81276_new_n3375_));
AND2X2 AND2X2_6105 ( .A(u5__abc_81276_new_n3374_), .B(u5__abc_81276_new_n3375_), .Y(u5__abc_81276_new_n3376_));
AND2X2 AND2X2_6106 ( .A(u5__abc_81276_new_n3376_), .B(u5__abc_81276_new_n2658_), .Y(u5__abc_81276_new_n3377_));
AND2X2 AND2X2_6107 ( .A(u5__abc_81276_new_n1450_), .B(u5__abc_81276_new_n3378_), .Y(u5__abc_81276_new_n3379_));
AND2X2 AND2X2_6108 ( .A(u5__abc_81276_new_n1549_), .B(u5__abc_81276_new_n1728_), .Y(u5__abc_81276_new_n3381_));
AND2X2 AND2X2_6109 ( .A(u5_state_9_), .B(u5_wb_wait), .Y(u5__abc_81276_new_n3383_));
AND2X2 AND2X2_611 ( .A(spec_req_cs_3_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n2199_));
AND2X2 AND2X2_6110 ( .A(u5__abc_81276_new_n3303_), .B(u5__abc_81276_new_n3362_), .Y(u5__abc_81276_new_n3384_));
AND2X2 AND2X2_6111 ( .A(u5__abc_81276_new_n3386_), .B(u5__abc_81276_new_n3382_), .Y(u5__abc_81276_new_n3387_));
AND2X2 AND2X2_6112 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3387_), .Y(u5__abc_81276_new_n3388_));
AND2X2 AND2X2_6113 ( .A(u5_kro), .B(u5_wb_wait_r), .Y(u5__abc_81276_new_n3389_));
AND2X2 AND2X2_6114 ( .A(u5__abc_81276_new_n3389_), .B(u5__abc_81276_new_n460_), .Y(u5__abc_81276_new_n3390_));
AND2X2 AND2X2_6115 ( .A(u5__abc_81276_new_n1457_), .B(u5__abc_81276_new_n2953__bF_buf2), .Y(u5__abc_81276_new_n3392_));
AND2X2 AND2X2_6116 ( .A(u5__abc_81276_new_n3393_), .B(u5__abc_81276_new_n3353_), .Y(u5__abc_81276_new_n3394_));
AND2X2 AND2X2_6117 ( .A(u5__abc_81276_new_n1492_), .B(u5__abc_81276_new_n3394_), .Y(u5__abc_81276_new_n3395_));
AND2X2 AND2X2_6118 ( .A(u5__abc_81276_new_n1450_), .B(u5__abc_81276_new_n3396_), .Y(u5__abc_81276_new_n3397_));
AND2X2 AND2X2_6119 ( .A(u5__abc_81276_new_n3399_), .B(u5__abc_81276_new_n3391_), .Y(u5__abc_81276_new_n3400_));
AND2X2 AND2X2_612 ( .A(u0__abc_76628_new_n2200_), .B(u0__abc_76628_new_n1173__bF_buf5), .Y(u0__abc_76628_new_n2201_));
AND2X2 AND2X2_6120 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_10_), .Y(u5__abc_81276_new_n3402_));
AND2X2 AND2X2_6121 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3402_), .Y(u5__abc_81276_new_n3403_));
AND2X2 AND2X2_6122 ( .A(u5__abc_81276_new_n1457_), .B(u5_cmd_asserted_bF_buf2), .Y(u5__abc_81276_new_n3404_));
AND2X2 AND2X2_6123 ( .A(u5__abc_81276_new_n1478_), .B(u5__abc_81276_new_n1712_), .Y(u5__abc_81276_new_n3405_));
AND2X2 AND2X2_6124 ( .A(u5__abc_81276_new_n1836_), .B(u5_state_11_), .Y(u5__abc_81276_new_n3408_));
AND2X2 AND2X2_6125 ( .A(u5_wb_cycle), .B(u1_wb_write_go), .Y(u5__abc_81276_new_n3410_));
AND2X2 AND2X2_6126 ( .A(u5__abc_81276_new_n1472_), .B(u5__abc_81276_new_n3411_), .Y(u5__abc_81276_new_n3412_));
AND2X2 AND2X2_6127 ( .A(u5__abc_81276_new_n3409_), .B(u5__abc_81276_new_n3412_), .Y(u5__abc_81276_new_n3413_));
AND2X2 AND2X2_6128 ( .A(u5__abc_81276_new_n3413_), .B(u5__abc_81276_new_n3408_), .Y(u5__abc_81276_new_n3414_));
AND2X2 AND2X2_6129 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_11_), .Y(u5__abc_81276_new_n3415_));
AND2X2 AND2X2_613 ( .A(spec_req_cs_2_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n2202_));
AND2X2 AND2X2_6130 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3415_), .Y(u5__abc_81276_new_n3416_));
AND2X2 AND2X2_6131 ( .A(u5__abc_81276_new_n1478_), .B(u5__abc_81276_new_n3417_), .Y(u5__abc_81276_new_n3418_));
AND2X2 AND2X2_6132 ( .A(u5__abc_81276_new_n3413_), .B(u5__abc_81276_new_n3421_), .Y(u5__abc_81276_new_n3422_));
AND2X2 AND2X2_6133 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_12_), .Y(u5__abc_81276_new_n3423_));
AND2X2 AND2X2_6134 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3423_), .Y(u5__abc_81276_new_n3424_));
AND2X2 AND2X2_6135 ( .A(u5__abc_81276_new_n3425_), .B(u5_state_12_), .Y(u5__abc_81276_new_n3426_));
AND2X2 AND2X2_6136 ( .A(u5__abc_81276_new_n3272_), .B(u5__abc_81276_new_n3426_), .Y(u5__abc_81276_new_n3427_));
AND2X2 AND2X2_6137 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_13_), .Y(u5__abc_81276_new_n3430_));
AND2X2 AND2X2_6138 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3430_), .Y(u5__abc_81276_new_n3431_));
AND2X2 AND2X2_6139 ( .A(u5__abc_81276_new_n1443_), .B(u5__abc_81276_new_n2953__bF_buf1), .Y(u5__abc_81276_new_n3432_));
AND2X2 AND2X2_614 ( .A(u0__abc_76628_new_n2203_), .B(u0__abc_76628_new_n1172__bF_buf5), .Y(u0__abc_76628_new_n2204_));
AND2X2 AND2X2_6140 ( .A(u5__abc_81276_new_n1492_), .B(u5__abc_81276_new_n1851_), .Y(u5__abc_81276_new_n3433_));
AND2X2 AND2X2_6141 ( .A(u5__abc_81276_new_n1123_), .B(u5_cmd_asserted_bF_buf0), .Y(u5__abc_81276_new_n3440_));
AND2X2 AND2X2_6142 ( .A(u5__abc_81276_new_n3441_), .B(u5__abc_81276_new_n3439_), .Y(u5__abc_81276_new_n3442_));
AND2X2 AND2X2_6143 ( .A(u5__abc_81276_new_n1443_), .B(u5__abc_81276_new_n3442_), .Y(u5__abc_81276_new_n3443_));
AND2X2 AND2X2_6144 ( .A(u5__abc_81276_new_n3438_), .B(u5__abc_81276_new_n3443_), .Y(u5__abc_81276_new_n3444_));
AND2X2 AND2X2_6145 ( .A(u5__abc_81276_new_n3215__bF_buf2), .B(u5_state_14_), .Y(u5__abc_81276_new_n3445_));
AND2X2 AND2X2_6146 ( .A(u5__abc_81276_new_n3447_), .B(u5__abc_81276_new_n3446_), .Y(u5__abc_81276_new_n3448_));
AND2X2 AND2X2_6147 ( .A(u5__abc_81276_new_n1836_), .B(u5__abc_81276_new_n3448_), .Y(u5__abc_81276_new_n3449_));
AND2X2 AND2X2_6148 ( .A(u5__abc_81276_new_n3450_), .B(u5__abc_81276_new_n1623_), .Y(u5__abc_81276_new_n3451_));
AND2X2 AND2X2_6149 ( .A(u5__abc_81276_new_n943_), .B(u5__abc_81276_new_n2953__bF_buf3), .Y(u5__abc_81276_new_n3454_));
AND2X2 AND2X2_615 ( .A(spec_req_cs_1_bF_buf2_), .B(u0_csc1_10_), .Y(u0__abc_76628_new_n2205_));
AND2X2 AND2X2_6150 ( .A(u5_state_15_), .B(u5_wb_wait), .Y(u5__abc_81276_new_n3456_));
AND2X2 AND2X2_6151 ( .A(u5__abc_81276_new_n3457_), .B(u5__abc_81276_new_n3455_), .Y(u5__abc_81276_new_n3458_));
AND2X2 AND2X2_6152 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3458_), .Y(u5__abc_81276_new_n3459_));
AND2X2 AND2X2_6153 ( .A(u5__abc_81276_new_n2953__bF_buf2), .B(u5_state_15_), .Y(u5__abc_81276_new_n3460_));
AND2X2 AND2X2_6154 ( .A(u5__abc_81276_new_n1614_), .B(u5__abc_81276_new_n3440_), .Y(u5__abc_81276_new_n3461_));
AND2X2 AND2X2_6155 ( .A(u5__abc_81276_new_n3462_), .B(u5__abc_81276_new_n836_), .Y(u5__abc_81276_new_n3463_));
AND2X2 AND2X2_6156 ( .A(u5__abc_81276_new_n1836_), .B(u5__abc_81276_new_n3466_), .Y(u5__abc_81276_new_n3467_));
AND2X2 AND2X2_6157 ( .A(u5__abc_81276_new_n3468_), .B(u5__abc_81276_new_n1472_), .Y(u5__abc_81276_new_n3469_));
AND2X2 AND2X2_6158 ( .A(u5__abc_81276_new_n3446_), .B(u5_state_15_), .Y(u5__abc_81276_new_n3471_));
AND2X2 AND2X2_6159 ( .A(u5__abc_81276_new_n1836_), .B(u5__abc_81276_new_n3471_), .Y(u5__abc_81276_new_n3472_));
AND2X2 AND2X2_616 ( .A(u0__abc_76628_new_n1946__bF_buf2), .B(u0__abc_76628_new_n2208_), .Y(u0__abc_76628_new_n2209_));
AND2X2 AND2X2_6160 ( .A(u5__abc_81276_new_n3473_), .B(u5__abc_81276_new_n3447_), .Y(u5__abc_81276_new_n3474_));
AND2X2 AND2X2_6161 ( .A(u5__abc_81276_new_n3475_), .B(u5__abc_81276_new_n3253_), .Y(u5__abc_81276_new_n3476_));
AND2X2 AND2X2_6162 ( .A(u5__abc_81276_new_n1123_), .B(u5__abc_81276_new_n3238_), .Y(u5__abc_81276_new_n3478_));
AND2X2 AND2X2_6163 ( .A(u5__abc_81276_new_n3283_), .B(u5__abc_81276_new_n3478_), .Y(u5__abc_81276_new_n3479_));
AND2X2 AND2X2_6164 ( .A(u5__abc_81276_new_n3480_), .B(u5__abc_81276_new_n3288_), .Y(u5__abc_81276_new_n3481_));
AND2X2 AND2X2_6165 ( .A(u5__abc_81276_new_n3438_), .B(u5__abc_81276_new_n3481_), .Y(u5__abc_81276_new_n3482_));
AND2X2 AND2X2_6166 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_16_), .Y(u5__abc_81276_new_n3483_));
AND2X2 AND2X2_6167 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3483_), .Y(u5__abc_81276_new_n3484_));
AND2X2 AND2X2_6168 ( .A(u5__abc_81276_new_n3231_), .B(u5_state_16_), .Y(u5__abc_81276_new_n3485_));
AND2X2 AND2X2_6169 ( .A(u5__abc_81276_new_n3276_), .B(u5__abc_81276_new_n3485_), .Y(u5__abc_81276_new_n3486_));
AND2X2 AND2X2_617 ( .A(u0__abc_76628_new_n2207_), .B(u0__abc_76628_new_n2209_), .Y(u0__abc_76628_new_n2210_));
AND2X2 AND2X2_6170 ( .A(u5__abc_81276_new_n3425_), .B(u5_state_16_), .Y(u5__abc_81276_new_n3487_));
AND2X2 AND2X2_6171 ( .A(u5__abc_81276_new_n3488_), .B(u5__abc_81276_new_n1405_), .Y(u5__abc_81276_new_n3489_));
AND2X2 AND2X2_6172 ( .A(u5__abc_81276_new_n1412_), .B(u5__abc_81276_new_n3490_), .Y(u5__abc_81276_new_n3491_));
AND2X2 AND2X2_6173 ( .A(u5__abc_81276_new_n3446_), .B(u5_state_16_), .Y(u5__abc_81276_new_n3496_));
AND2X2 AND2X2_6174 ( .A(u5__abc_81276_new_n1836_), .B(u5__abc_81276_new_n3496_), .Y(u5__abc_81276_new_n3497_));
AND2X2 AND2X2_6175 ( .A(u5__abc_81276_new_n3242_), .B(u5__abc_81276_new_n3447_), .Y(u5__abc_81276_new_n3499_));
AND2X2 AND2X2_6176 ( .A(u5__abc_81276_new_n3498_), .B(u5__abc_81276_new_n3499_), .Y(u5__abc_81276_new_n3500_));
AND2X2 AND2X2_6177 ( .A(u5__abc_81276_new_n3501_), .B(u5__abc_81276_new_n3253_), .Y(u5__abc_81276_new_n3502_));
AND2X2 AND2X2_6178 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_17_), .Y(u5__abc_81276_new_n3504_));
AND2X2 AND2X2_6179 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3504_), .Y(u5__abc_81276_new_n3505_));
AND2X2 AND2X2_618 ( .A(u0__abc_76628_new_n1170__bF_buf6), .B(tms_0_), .Y(u0__abc_76628_new_n2716_));
AND2X2 AND2X2_6180 ( .A(u5__abc_81276_new_n2953__bF_buf0), .B(u5_state_17_), .Y(u5__abc_81276_new_n3506_));
AND2X2 AND2X2_6181 ( .A(u5__abc_81276_new_n3508_), .B(u5__abc_81276_new_n3506_), .Y(u5__abc_81276_new_n3509_));
AND2X2 AND2X2_6182 ( .A(u5__abc_81276_new_n1382_), .B(u5__abc_81276_new_n1712_), .Y(u5__abc_81276_new_n3511_));
AND2X2 AND2X2_6183 ( .A(u5__abc_81276_new_n3512_), .B(u5__abc_81276_new_n3510_), .Y(u5__abc_81276_new_n3513_));
AND2X2 AND2X2_6184 ( .A(u5__abc_81276_new_n1712_), .B(u5_state_17_), .Y(u5__abc_81276_new_n3514_));
AND2X2 AND2X2_6185 ( .A(u5__abc_81276_new_n1504_), .B(u5__abc_81276_new_n3515_), .Y(u5__abc_81276_new_n3516_));
AND2X2 AND2X2_6186 ( .A(u5__abc_81276_new_n1554_), .B(u5_state_18_), .Y(u5__abc_81276_new_n3520_));
AND2X2 AND2X2_6187 ( .A(u5__abc_81276_new_n3213_), .B(u5__abc_81276_new_n3520_), .Y(u5__abc_81276_new_n3521_));
AND2X2 AND2X2_6188 ( .A(u5__abc_81276_new_n3323__bF_buf0), .B(u5__abc_81276_new_n3522_), .Y(u5__abc_81276_new_n3523_));
AND2X2 AND2X2_6189 ( .A(u5__abc_81276_new_n629_), .B(u5__abc_81276_new_n2953__bF_buf3), .Y(u5__abc_81276_new_n3524_));
AND2X2 AND2X2_619 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2721_));
AND2X2 AND2X2_6190 ( .A(u5__abc_81276_new_n1555_), .B(u5_state_19_), .Y(u5__abc_81276_new_n3526_));
AND2X2 AND2X2_6191 ( .A(u5__abc_81276_new_n3213_), .B(u5__abc_81276_new_n3526_), .Y(u5__abc_81276_new_n3527_));
AND2X2 AND2X2_6192 ( .A(u5__abc_81276_new_n3323__bF_buf3), .B(u5__abc_81276_new_n3527_), .Y(u5__abc_81276_new_n3528_));
AND2X2 AND2X2_6193 ( .A(u5__abc_81276_new_n1712_), .B(u5_state_19_), .Y(u5__abc_81276_new_n3529_));
AND2X2 AND2X2_6194 ( .A(u5__abc_81276_new_n611_), .B(u5__abc_81276_new_n3529_), .Y(u5__abc_81276_new_n3530_));
AND2X2 AND2X2_6195 ( .A(u5__abc_81276_new_n629_), .B(u5__abc_81276_new_n3531_), .Y(u5__abc_81276_new_n3532_));
AND2X2 AND2X2_6196 ( .A(u5__abc_81276_new_n1526__bF_buf2), .B(u5__abc_81276_new_n1557_), .Y(u5__abc_81276_new_n3535_));
AND2X2 AND2X2_6197 ( .A(u5__abc_81276_new_n3299_), .B(u5_state_20_), .Y(u5__abc_81276_new_n3536_));
AND2X2 AND2X2_6198 ( .A(u5__abc_81276_new_n3213_), .B(u5__abc_81276_new_n3536_), .Y(u5__abc_81276_new_n3537_));
AND2X2 AND2X2_6199 ( .A(u5__abc_81276_new_n3535_), .B(u5__abc_81276_new_n3537_), .Y(u5__abc_81276_new_n3538_));
AND2X2 AND2X2_62 ( .A(u0__abc_76628_new_n1100_), .B(u0_lmr_req1), .Y(u0__abc_76628_new_n1111_));
AND2X2 AND2X2_620 ( .A(u0__abc_76628_new_n2725_), .B(u0__abc_76628_new_n2724__bF_buf5), .Y(u0__abc_76628_new_n2726_));
AND2X2 AND2X2_6200 ( .A(u5__abc_81276_new_n611_), .B(u5__abc_81276_new_n3539_), .Y(u5__abc_81276_new_n3540_));
AND2X2 AND2X2_6201 ( .A(u5__abc_81276_new_n2953__bF_buf2), .B(u5_state_20_), .Y(u5__abc_81276_new_n3541_));
AND2X2 AND2X2_6202 ( .A(u5__abc_81276_new_n3259_), .B(u5__abc_81276_new_n3541_), .Y(u5__abc_81276_new_n3542_));
AND2X2 AND2X2_6203 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_21_), .Y(u5__abc_81276_new_n3545_));
AND2X2 AND2X2_6204 ( .A(u5__abc_81276_new_n3535_), .B(u5__abc_81276_new_n3546_), .Y(u5_next_state_21_));
AND2X2 AND2X2_6205 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_22_), .Y(u5__abc_81276_new_n3548_));
AND2X2 AND2X2_6206 ( .A(u5__abc_81276_new_n3323__bF_buf2), .B(u5__abc_81276_new_n3548_), .Y(u5__abc_81276_new_n3549_));
AND2X2 AND2X2_6207 ( .A(u5__abc_81276_new_n2953__bF_buf1), .B(u5_state_22_), .Y(u5__abc_81276_new_n3551_));
AND2X2 AND2X2_6208 ( .A(u5__abc_81276_new_n1356_), .B(u5__abc_81276_new_n3551_), .Y(u5__abc_81276_new_n3552_));
AND2X2 AND2X2_6209 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_23_), .Y(u5__abc_81276_new_n3555_));
AND2X2 AND2X2_621 ( .A(u0__abc_76628_new_n2726_), .B(u0__abc_76628_new_n2723_), .Y(u0__abc_76628_new_n2727_));
AND2X2 AND2X2_6210 ( .A(u5__abc_81276_new_n3323__bF_buf1), .B(u5__abc_81276_new_n3555_), .Y(u5__abc_81276_new_n3556_));
AND2X2 AND2X2_6211 ( .A(u5__abc_81276_new_n1356_), .B(u5__abc_81276_new_n3557_), .Y(u5__abc_81276_new_n3558_));
AND2X2 AND2X2_6212 ( .A(u5__abc_81276_new_n1712_), .B(u5_state_23_), .Y(u5__abc_81276_new_n3559_));
AND2X2 AND2X2_6213 ( .A(u5__abc_81276_new_n1363_), .B(u5__abc_81276_new_n3559_), .Y(u5__abc_81276_new_n3560_));
AND2X2 AND2X2_6214 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_24_), .Y(u5__abc_81276_new_n3563_));
AND2X2 AND2X2_6215 ( .A(u5__abc_81276_new_n3323__bF_buf0), .B(u5__abc_81276_new_n3563_), .Y(u5__abc_81276_new_n3564_));
AND2X2 AND2X2_6216 ( .A(u5_tmr_done_bF_buf2), .B(u5_ir_cnt_done), .Y(u5__abc_81276_new_n3565_));
AND2X2 AND2X2_6217 ( .A(u5__abc_81276_new_n3568_), .B(u5__abc_81276_new_n3569_), .Y(u5__abc_81276_new_n3570_));
AND2X2 AND2X2_6218 ( .A(u5__abc_81276_new_n3570_), .B(u5__abc_81276_new_n3567_), .Y(u5__abc_81276_new_n3571_));
AND2X2 AND2X2_6219 ( .A(u5__abc_81276_new_n638_), .B(u5__abc_81276_new_n2953__bF_buf0), .Y(u5__abc_81276_new_n3572_));
AND2X2 AND2X2_622 ( .A(u0__abc_76628_new_n2728_), .B(u0__abc_76628_new_n2720__bF_buf5), .Y(u0__abc_76628_new_n2729_));
AND2X2 AND2X2_6220 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_25_), .Y(u5__abc_81276_new_n3575_));
AND2X2 AND2X2_6221 ( .A(u5__abc_81276_new_n3323__bF_buf3), .B(u5__abc_81276_new_n3575_), .Y(u5__abc_81276_new_n3576_));
AND2X2 AND2X2_6222 ( .A(u5__abc_81276_new_n1372_), .B(u5__abc_81276_new_n3577_), .Y(u5__abc_81276_new_n3578_));
AND2X2 AND2X2_6223 ( .A(u5__abc_81276_new_n1712_), .B(u5_state_25_), .Y(u5__abc_81276_new_n3579_));
AND2X2 AND2X2_6224 ( .A(u5__abc_81276_new_n1360_), .B(u5__abc_81276_new_n3579_), .Y(u5__abc_81276_new_n3580_));
AND2X2 AND2X2_6225 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_26_), .Y(u5__abc_81276_new_n3583_));
AND2X2 AND2X2_6226 ( .A(u5__abc_81276_new_n3323__bF_buf2), .B(u5__abc_81276_new_n3583_), .Y(u5__abc_81276_new_n3584_));
AND2X2 AND2X2_6227 ( .A(u5__abc_81276_new_n1712_), .B(u5_state_26_), .Y(u5__abc_81276_new_n3585_));
AND2X2 AND2X2_6228 ( .A(u5__abc_81276_new_n1360_), .B(u5__abc_81276_new_n3586_), .Y(u5__abc_81276_new_n3587_));
AND2X2 AND2X2_6229 ( .A(u5__abc_81276_new_n2953__bF_buf3), .B(u5_state_26_), .Y(u5__abc_81276_new_n3588_));
AND2X2 AND2X2_623 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2730_));
AND2X2 AND2X2_6230 ( .A(u5__abc_81276_new_n3259_), .B(u5__abc_81276_new_n3588_), .Y(u5__abc_81276_new_n3589_));
AND2X2 AND2X2_6231 ( .A(u5__abc_81276_new_n3323__bF_buf1), .B(u5__abc_81276_new_n1551_), .Y(u5__abc_81276_new_n3592_));
AND2X2 AND2X2_6232 ( .A(u5__abc_81276_new_n3213_), .B(u5_state_27_), .Y(u5__abc_81276_new_n3593_));
AND2X2 AND2X2_6233 ( .A(u5__abc_81276_new_n3592_), .B(u5__abc_81276_new_n3594_), .Y(u5__abc_81276_new_n3595_));
AND2X2 AND2X2_6234 ( .A(u5__abc_81276_new_n602_), .B(u5__abc_81276_new_n2953__bF_buf2), .Y(u5__abc_81276_new_n3596_));
AND2X2 AND2X2_6235 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_28_), .Y(u5__abc_81276_new_n3598_));
AND2X2 AND2X2_6236 ( .A(u5__abc_81276_new_n3323__bF_buf0), .B(u5__abc_81276_new_n3598_), .Y(u5__abc_81276_new_n3599_));
AND2X2 AND2X2_6237 ( .A(u5__abc_81276_new_n1433_), .B(u5__abc_81276_new_n3600_), .Y(u5__abc_81276_new_n3601_));
AND2X2 AND2X2_6238 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_29_), .Y(u5__abc_81276_new_n3604_));
AND2X2 AND2X2_6239 ( .A(u5__abc_81276_new_n3323__bF_buf3), .B(u5__abc_81276_new_n3604_), .Y(u5__abc_81276_new_n3605_));
AND2X2 AND2X2_624 ( .A(u0__abc_76628_new_n2731_), .B(u0__abc_76628_new_n2719__bF_buf5), .Y(u0__abc_76628_new_n2732_));
AND2X2 AND2X2_6240 ( .A(u5__abc_81276_new_n2746_), .B(u5__abc_81276_new_n3606_), .Y(u5__abc_81276_new_n3607_));
AND2X2 AND2X2_6241 ( .A(u5__abc_81276_new_n2953__bF_buf1), .B(u5_state_29_), .Y(u5__abc_81276_new_n3608_));
AND2X2 AND2X2_6242 ( .A(u5__abc_81276_new_n1941_), .B(u5__abc_81276_new_n3608_), .Y(u5__abc_81276_new_n3609_));
AND2X2 AND2X2_6243 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_30_), .Y(u5__abc_81276_new_n3612_));
AND2X2 AND2X2_6244 ( .A(u5__abc_81276_new_n3323__bF_buf2), .B(u5__abc_81276_new_n3612_), .Y(u5__abc_81276_new_n3613_));
AND2X2 AND2X2_6245 ( .A(u5__abc_81276_new_n1941_), .B(u5__abc_81276_new_n3614_), .Y(u5__abc_81276_new_n3615_));
AND2X2 AND2X2_6246 ( .A(u5__abc_81276_new_n3616_), .B(u5_state_30_), .Y(u5__abc_81276_new_n3617_));
AND2X2 AND2X2_6247 ( .A(u5__abc_81276_new_n2743_), .B(u5__abc_81276_new_n3617_), .Y(u5__abc_81276_new_n3618_));
AND2X2 AND2X2_6248 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_31_), .Y(u5__abc_81276_new_n3621_));
AND2X2 AND2X2_6249 ( .A(u5__abc_81276_new_n3323__bF_buf1), .B(u5__abc_81276_new_n3621_), .Y(u5__abc_81276_new_n3622_));
AND2X2 AND2X2_625 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2733_));
AND2X2 AND2X2_6250 ( .A(u5__abc_81276_new_n516_), .B(u5__abc_81276_new_n3623_), .Y(u5__abc_81276_new_n3624_));
AND2X2 AND2X2_6251 ( .A(u5__abc_81276_new_n3347_), .B(u5_state_32_), .Y(u5__abc_81276_new_n3626_));
AND2X2 AND2X2_6252 ( .A(u5__abc_81276_new_n3323__bF_buf0), .B(u5__abc_81276_new_n3626_), .Y(u5__abc_81276_new_n3627_));
AND2X2 AND2X2_6253 ( .A(u5__abc_81276_new_n1712_), .B(u5_state_32_), .Y(u5__abc_81276_new_n3628_));
AND2X2 AND2X2_6254 ( .A(u5__abc_81276_new_n530_), .B(u5__abc_81276_new_n3628_), .Y(u5__abc_81276_new_n3629_));
AND2X2 AND2X2_6255 ( .A(u5__abc_81276_new_n3633_), .B(u5__abc_81276_new_n3346_), .Y(u5__abc_81276_new_n3634_));
AND2X2 AND2X2_6256 ( .A(u5__abc_81276_new_n3323__bF_buf3), .B(u5__abc_81276_new_n3634_), .Y(u5_next_state_33_));
AND2X2 AND2X2_6257 ( .A(u5__abc_81276_new_n3215__bF_buf1), .B(u5_state_34_), .Y(u5__abc_81276_new_n3636_));
AND2X2 AND2X2_6258 ( .A(u5__abc_81276_new_n3215__bF_buf0), .B(u5_state_35_), .Y(u5__abc_81276_new_n3638_));
AND2X2 AND2X2_6259 ( .A(u5__abc_81276_new_n1428_), .B(mc_br_r), .Y(u5__abc_81276_new_n3639_));
AND2X2 AND2X2_626 ( .A(u0__abc_76628_new_n2734_), .B(u0__abc_76628_new_n2718__bF_buf5), .Y(u0__abc_76628_new_n2735_));
AND2X2 AND2X2_6260 ( .A(u5__abc_81276_new_n3326_), .B(u5__abc_81276_new_n3362_), .Y(u5__abc_81276_new_n3642_));
AND2X2 AND2X2_6261 ( .A(u5__abc_81276_new_n3642_), .B(u5_state_36_), .Y(u5__abc_81276_new_n3643_));
AND2X2 AND2X2_6262 ( .A(u5__abc_81276_new_n1727_), .B(u5__abc_81276_new_n1690_), .Y(u5__abc_81276_new_n3644_));
AND2X2 AND2X2_6263 ( .A(u5__abc_81276_new_n3644_), .B(u5__abc_81276_new_n1693_), .Y(u5__abc_81276_new_n3645_));
AND2X2 AND2X2_6264 ( .A(u5__abc_81276_new_n3324_), .B(u5__abc_81276_new_n3648_), .Y(u5__abc_81276_new_n3649_));
AND2X2 AND2X2_6265 ( .A(u5__abc_81276_new_n3647_), .B(u5__abc_81276_new_n3649_), .Y(u5__abc_81276_new_n3650_));
AND2X2 AND2X2_6266 ( .A(u5__abc_81276_new_n3323__bF_buf2), .B(u5__abc_81276_new_n3650_), .Y(u5_next_state_36_));
AND2X2 AND2X2_6267 ( .A(u5__abc_81276_new_n3215__bF_buf4), .B(u5_state_37_), .Y(u5__abc_81276_new_n3652_));
AND2X2 AND2X2_6268 ( .A(u5__abc_81276_new_n1708_), .B(u5_state_37_), .Y(u5__abc_81276_new_n3654_));
AND2X2 AND2X2_6269 ( .A(u5__abc_81276_new_n3653_), .B(u5__abc_81276_new_n3654_), .Y(u5__abc_81276_new_n3655_));
AND2X2 AND2X2_627 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2736_));
AND2X2 AND2X2_6270 ( .A(u5__abc_81276_new_n3215__bF_buf3), .B(u5_state_38_), .Y(u5__abc_81276_new_n3658_));
AND2X2 AND2X2_6271 ( .A(u5__abc_81276_new_n2195_), .B(u5__abc_81276_new_n490__bF_buf7), .Y(u5__abc_81276_new_n3659_));
AND2X2 AND2X2_6272 ( .A(u5__abc_81276_new_n1750_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3661_));
AND2X2 AND2X2_6273 ( .A(u5__abc_81276_new_n3662_), .B(u5__abc_81276_new_n3660_), .Y(u5__abc_81276_new_n3663_));
AND2X2 AND2X2_6274 ( .A(u5__abc_81276_new_n3659_), .B(u5__abc_81276_new_n3663_), .Y(u5__abc_81276_new_n3664_));
AND2X2 AND2X2_6275 ( .A(u5__abc_81276_new_n3215__bF_buf2), .B(u5_state_39_), .Y(u5__abc_81276_new_n3666_));
AND2X2 AND2X2_6276 ( .A(u5__abc_81276_new_n761_), .B(u5__abc_81276_new_n3667_), .Y(u5__abc_81276_new_n3668_));
AND2X2 AND2X2_6277 ( .A(u5__abc_81276_new_n3215__bF_buf1), .B(u5_state_40_), .Y(u5__abc_81276_new_n3671_));
AND2X2 AND2X2_6278 ( .A(u5__abc_81276_new_n3215__bF_buf0), .B(u5_state_41_), .Y(u5__abc_81276_new_n3673_));
AND2X2 AND2X2_6279 ( .A(u5__abc_81276_new_n3674_), .B(u5__abc_81276_new_n3675_), .Y(u5__abc_81276_new_n3676_));
AND2X2 AND2X2_628 ( .A(u0__abc_76628_new_n2737_), .B(u0__abc_76628_new_n2717__bF_buf5), .Y(u0__abc_76628_new_n2738_));
AND2X2 AND2X2_6280 ( .A(u5__abc_81276_new_n3659_), .B(u5__abc_81276_new_n3676_), .Y(u5__abc_81276_new_n3677_));
AND2X2 AND2X2_6281 ( .A(u5__abc_81276_new_n3215__bF_buf4), .B(u5_state_42_), .Y(u5__abc_81276_new_n3679_));
AND2X2 AND2X2_6282 ( .A(u5__abc_81276_new_n1708_), .B(u5_state_42_), .Y(u5__abc_81276_new_n3680_));
AND2X2 AND2X2_6283 ( .A(u5__abc_81276_new_n1323_), .B(u5__abc_81276_new_n3680_), .Y(u5__abc_81276_new_n3681_));
AND2X2 AND2X2_6284 ( .A(u5__abc_81276_new_n1323_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3684_));
AND2X2 AND2X2_6285 ( .A(u5__abc_81276_new_n3686_), .B(u5__abc_81276_new_n3685_), .Y(u5_next_state_43_));
AND2X2 AND2X2_6286 ( .A(u5__abc_81276_new_n3215__bF_buf2), .B(u5_state_44_), .Y(u5__abc_81276_new_n3688_));
AND2X2 AND2X2_6287 ( .A(u5__abc_81276_new_n1708_), .B(u5_state_44_), .Y(u5__abc_81276_new_n3689_));
AND2X2 AND2X2_6288 ( .A(u5__abc_81276_new_n2996_), .B(u5__abc_81276_new_n3689_), .Y(u5__abc_81276_new_n3690_));
AND2X2 AND2X2_6289 ( .A(u5__abc_81276_new_n3215__bF_buf1), .B(u5_state_45_), .Y(u5__abc_81276_new_n3693_));
AND2X2 AND2X2_629 ( .A(u0_tms1_0_), .B(u0_cs1_bF_buf4), .Y(u0__abc_76628_new_n2739_));
AND2X2 AND2X2_6290 ( .A(u5__abc_81276_new_n1750_), .B(csc_s_4_), .Y(u5__abc_81276_new_n3695_));
AND2X2 AND2X2_6291 ( .A(u5__abc_81276_new_n1336_), .B(u5__abc_81276_new_n3696_), .Y(u5__abc_81276_new_n3697_));
AND2X2 AND2X2_6292 ( .A(u5__abc_81276_new_n3698_), .B(u5__abc_81276_new_n3694_), .Y(u5__abc_81276_new_n3699_));
AND2X2 AND2X2_6293 ( .A(u5__abc_81276_new_n3215__bF_buf0), .B(u5_state_46_), .Y(u5__abc_81276_new_n3701_));
AND2X2 AND2X2_6294 ( .A(u5__abc_81276_new_n1708_), .B(u5_state_46_), .Y(u5__abc_81276_new_n3702_));
AND2X2 AND2X2_6295 ( .A(u5__abc_81276_new_n1309_), .B(u5__abc_81276_new_n3702_), .Y(u5__abc_81276_new_n3703_));
AND2X2 AND2X2_6296 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_47_), .Y(u5__abc_81276_new_n3706_));
AND2X2 AND2X2_6297 ( .A(u5__abc_81276_new_n3644_), .B(u5__abc_81276_new_n1537_), .Y(u5__abc_81276_new_n3707_));
AND2X2 AND2X2_6298 ( .A(u5__abc_81276_new_n1549_), .B(u5__abc_81276_new_n3707_), .Y(u5__abc_81276_new_n3708_));
AND2X2 AND2X2_6299 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3709_), .Y(u5_next_state_47_));
AND2X2 AND2X2_63 ( .A(init_req), .B(u0_init_req1), .Y(u0__abc_76628_new_n1112_));
AND2X2 AND2X2_630 ( .A(u0__abc_76628_new_n1169__bF_buf5), .B(u0__abc_76628_new_n2743_), .Y(u0__abc_76628_new_n2744_));
AND2X2 AND2X2_6300 ( .A(u5__abc_81276_new_n1708_), .B(u5_state_48_), .Y(u5__abc_81276_new_n3711_));
AND2X2 AND2X2_6301 ( .A(u5__abc_81276_new_n720_), .B(u5__abc_81276_new_n3711_), .Y(u5__abc_81276_new_n3712_));
AND2X2 AND2X2_6302 ( .A(u5__abc_81276_new_n3215__bF_buf4), .B(u5_state_48_), .Y(u5__abc_81276_new_n3713_));
AND2X2 AND2X2_6303 ( .A(u5__abc_81276_new_n1287_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3716_));
AND2X2 AND2X2_6304 ( .A(u5__abc_81276_new_n3718_), .B(u5__abc_81276_new_n3717_), .Y(u5_next_state_49_));
AND2X2 AND2X2_6305 ( .A(u5__abc_81276_new_n3215__bF_buf2), .B(u5_state_50_), .Y(u5__abc_81276_new_n3720_));
AND2X2 AND2X2_6306 ( .A(u5__abc_81276_new_n1270_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3723_));
AND2X2 AND2X2_6307 ( .A(u5__abc_81276_new_n3725_), .B(u5__abc_81276_new_n3724_), .Y(u5_next_state_51_));
AND2X2 AND2X2_6308 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_52_), .Y(u5__abc_81276_new_n3727_));
AND2X2 AND2X2_6309 ( .A(u5__abc_81276_new_n1831_), .B(u5__abc_81276_new_n1693_), .Y(u5__abc_81276_new_n3728_));
AND2X2 AND2X2_631 ( .A(u0__abc_76628_new_n2741_), .B(u0__abc_76628_new_n2744_), .Y(u0__abc_76628_new_n2745_));
AND2X2 AND2X2_6310 ( .A(u5__abc_81276_new_n1549_), .B(u5__abc_81276_new_n3728_), .Y(u5__abc_81276_new_n3729_));
AND2X2 AND2X2_6311 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3730_), .Y(u5__abc_81276_new_n3731_));
AND2X2 AND2X2_6312 ( .A(u5__abc_81276_new_n1181_), .B(u3_wb_read_go), .Y(u5__abc_81276_new_n3733_));
AND2X2 AND2X2_6313 ( .A(u5__abc_81276_new_n3733_), .B(u5__abc_81276_new_n3732_), .Y(u5__abc_81276_new_n3734_));
AND2X2 AND2X2_6314 ( .A(u5__abc_81276_new_n2953__bF_buf0), .B(u5_state_52_), .Y(u5__abc_81276_new_n3735_));
AND2X2 AND2X2_6315 ( .A(u5__abc_81276_new_n1200_), .B(u5__abc_81276_new_n3735_), .Y(u5__abc_81276_new_n3736_));
AND2X2 AND2X2_6316 ( .A(u5__abc_81276_new_n3215__bF_buf0), .B(u5_state_53_), .Y(u5__abc_81276_new_n3739_));
AND2X2 AND2X2_6317 ( .A(u5__abc_81276_new_n1206_), .B(u5__abc_81276_new_n1708_), .Y(u5__abc_81276_new_n3740_));
AND2X2 AND2X2_6318 ( .A(u5__abc_81276_new_n1200_), .B(u5__abc_81276_new_n3741_), .Y(u5__abc_81276_new_n3742_));
AND2X2 AND2X2_6319 ( .A(u5__abc_81276_new_n1836_), .B(u3_wb_read_go), .Y(u5__abc_81276_new_n3745_));
AND2X2 AND2X2_632 ( .A(u0__abc_76628_new_n1170__bF_buf5), .B(tms_1_), .Y(u0__abc_76628_new_n2747_));
AND2X2 AND2X2_6320 ( .A(u5__abc_81276_new_n3745_), .B(u5__abc_81276_new_n1237_), .Y(u5__abc_81276_new_n3746_));
AND2X2 AND2X2_6321 ( .A(u5__abc_81276_new_n1206_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3747_));
AND2X2 AND2X2_6322 ( .A(u5__abc_81276_new_n3749_), .B(u5__abc_81276_new_n3748_), .Y(u5__abc_81276_new_n3750_));
AND2X2 AND2X2_6323 ( .A(u5__abc_81276_new_n3753_), .B(u5__abc_81276_new_n1237_), .Y(u5__abc_81276_new_n3754_));
AND2X2 AND2X2_6324 ( .A(u5_state_55_), .B(u5_wb_wait), .Y(u5__abc_81276_new_n3756_));
AND2X2 AND2X2_6325 ( .A(u5__abc_81276_new_n3757_), .B(u5__abc_81276_new_n3755_), .Y(u5__abc_81276_new_n3758_));
AND2X2 AND2X2_6326 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3758_), .Y(u5__abc_81276_new_n3759_));
AND2X2 AND2X2_6327 ( .A(u5__abc_81276_new_n3760_), .B(u5__abc_81276_new_n1821_), .Y(u5__abc_81276_new_n3761_));
AND2X2 AND2X2_6328 ( .A(u5__abc_81276_new_n3761_), .B(u3_wb_read_go), .Y(u5__abc_81276_new_n3762_));
AND2X2 AND2X2_6329 ( .A(u5_state_56_), .B(u5_wb_wait), .Y(u5__abc_81276_new_n3766_));
AND2X2 AND2X2_633 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2748_));
AND2X2 AND2X2_6330 ( .A(u5__abc_81276_new_n3767_), .B(u5__abc_81276_new_n3765_), .Y(u5__abc_81276_new_n3768_));
AND2X2 AND2X2_6331 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3768_), .Y(u5__abc_81276_new_n3769_));
AND2X2 AND2X2_6332 ( .A(u5__abc_81276_new_n3733_), .B(u5__abc_81276_new_n3766_), .Y(u5__abc_81276_new_n3770_));
AND2X2 AND2X2_6333 ( .A(u5__abc_81276_new_n3771_), .B(u3_wb_read_go), .Y(u5__abc_81276_new_n3772_));
AND2X2 AND2X2_6334 ( .A(u5__abc_81276_new_n3760_), .B(u5__abc_81276_new_n3772_), .Y(u5__abc_81276_new_n3773_));
AND2X2 AND2X2_6335 ( .A(u5__abc_81276_new_n3215__bF_buf3), .B(u5_state_57_), .Y(u5__abc_81276_new_n3776_));
AND2X2 AND2X2_6336 ( .A(u5__abc_81276_new_n3777_), .B(u5__abc_81276_new_n1124_), .Y(u5__abc_81276_new_n3778_));
AND2X2 AND2X2_6337 ( .A(u5_wb_wait), .B(u5_cmd_asserted_bF_buf0), .Y(u5__abc_81276_new_n3779_));
AND2X2 AND2X2_6338 ( .A(u5__abc_81276_new_n3781_), .B(u5__abc_81276_new_n3780_), .Y(u5__abc_81276_new_n3782_));
AND2X2 AND2X2_6339 ( .A(u5__abc_81276_new_n1849_), .B(u5__abc_81276_new_n3782_), .Y(u5__abc_81276_new_n3783_));
AND2X2 AND2X2_634 ( .A(u0__abc_76628_new_n2750_), .B(u0__abc_76628_new_n2724__bF_buf4), .Y(u0__abc_76628_new_n2751_));
AND2X2 AND2X2_6340 ( .A(u5__abc_81276_new_n1215_), .B(u5__abc_81276_new_n1693_), .Y(u5__abc_81276_new_n3784_));
AND2X2 AND2X2_6341 ( .A(u5__abc_81276_new_n1549_), .B(u5__abc_81276_new_n1832_), .Y(u5__abc_81276_new_n3788_));
AND2X2 AND2X2_6342 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_58_), .Y(u5__abc_81276_new_n3789_));
AND2X2 AND2X2_6343 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3790_), .Y(u5__abc_81276_new_n3791_));
AND2X2 AND2X2_6344 ( .A(u5__abc_81276_new_n3780_), .B(u5_state_58_), .Y(u5__abc_81276_new_n3792_));
AND2X2 AND2X2_6345 ( .A(u5__abc_81276_new_n3792_), .B(u5__abc_81276_new_n3441_), .Y(u5__abc_81276_new_n3793_));
AND2X2 AND2X2_6346 ( .A(u5__abc_81276_new_n1849_), .B(u5__abc_81276_new_n3793_), .Y(u5__abc_81276_new_n3794_));
AND2X2 AND2X2_6347 ( .A(u5__abc_81276_new_n3215__bF_buf2), .B(u5_state_59_), .Y(u5__abc_81276_new_n3797_));
AND2X2 AND2X2_6348 ( .A(u5__abc_81276_new_n3441_), .B(u5_state_59_), .Y(u5__abc_81276_new_n3798_));
AND2X2 AND2X2_6349 ( .A(u5__abc_81276_new_n1849_), .B(u5__abc_81276_new_n3799_), .Y(u5__abc_81276_new_n3800_));
AND2X2 AND2X2_635 ( .A(u0__abc_76628_new_n2751_), .B(u0__abc_76628_new_n2749_), .Y(u0__abc_76628_new_n2752_));
AND2X2 AND2X2_6350 ( .A(u5__abc_81276_new_n1215_), .B(u5_wb_wait), .Y(u5__abc_81276_new_n3801_));
AND2X2 AND2X2_6351 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_60_), .Y(u5__abc_81276_new_n3804_));
AND2X2 AND2X2_6352 ( .A(u5__abc_81276_new_n1697_), .B(u5__abc_81276_new_n1123_), .Y(u5__abc_81276_new_n3805_));
AND2X2 AND2X2_6353 ( .A(u5__abc_81276_new_n1549_), .B(u5__abc_81276_new_n3805_), .Y(u5__abc_81276_new_n3806_));
AND2X2 AND2X2_6354 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3807_), .Y(u5__abc_81276_new_n3808_));
AND2X2 AND2X2_6355 ( .A(u5__abc_81276_new_n1708_), .B(u5__abc_81276_new_n3809_), .Y(u5__abc_81276_new_n3810_));
AND2X2 AND2X2_6356 ( .A(u5__abc_81276_new_n3810_), .B(u5_state_60_), .Y(u5__abc_81276_new_n3811_));
AND2X2 AND2X2_6357 ( .A(u5__abc_81276_new_n1146_), .B(u5__abc_81276_new_n3811_), .Y(u5__abc_81276_new_n3812_));
AND2X2 AND2X2_6358 ( .A(u5__abc_81276_new_n3215__bF_buf1), .B(u5_state_61_), .Y(u5__abc_81276_new_n3814_));
AND2X2 AND2X2_6359 ( .A(u5__abc_81276_new_n1712_), .B(u5_state_61_), .Y(u5__abc_81276_new_n3815_));
AND2X2 AND2X2_636 ( .A(u0__abc_76628_new_n2753_), .B(u0__abc_76628_new_n2720__bF_buf4), .Y(u0__abc_76628_new_n2754_));
AND2X2 AND2X2_6360 ( .A(u5__abc_81276_new_n1141_), .B(u5__abc_81276_new_n3815_), .Y(u5__abc_81276_new_n3816_));
AND2X2 AND2X2_6361 ( .A(u5__abc_81276_new_n1708_), .B(u5_state_61_), .Y(u5__abc_81276_new_n3817_));
AND2X2 AND2X2_6362 ( .A(u5__abc_81276_new_n1146_), .B(u5__abc_81276_new_n3818_), .Y(u5__abc_81276_new_n3819_));
AND2X2 AND2X2_6363 ( .A(u5__abc_81276_new_n1141_), .B(u5_tmr_done_bF_buf3), .Y(u5__abc_81276_new_n3822_));
AND2X2 AND2X2_6364 ( .A(u5__abc_81276_new_n3824_), .B(u5__abc_81276_new_n3823_), .Y(u5_next_state_62_));
AND2X2 AND2X2_6365 ( .A(u5__abc_81276_new_n1549_), .B(u5__abc_81276_new_n1538_), .Y(u5__abc_81276_new_n3826_));
AND2X2 AND2X2_6366 ( .A(u5__abc_81276_new_n3212_), .B(u5_state_63_), .Y(u5__abc_81276_new_n3827_));
AND2X2 AND2X2_6367 ( .A(u5__abc_81276_new_n3361_), .B(u5__abc_81276_new_n3828_), .Y(u5__abc_81276_new_n3829_));
AND2X2 AND2X2_6368 ( .A(u5__abc_81276_new_n1002_), .B(u5__abc_81276_new_n3810_), .Y(u5__abc_81276_new_n3830_));
AND2X2 AND2X2_6369 ( .A(u5__abc_81276_new_n3215__bF_buf4), .B(u5_state_64_), .Y(u5__abc_81276_new_n3832_));
AND2X2 AND2X2_637 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2755_));
AND2X2 AND2X2_6370 ( .A(u5__abc_81276_new_n1708_), .B(u5_state_64_), .Y(u5__abc_81276_new_n3833_));
AND2X2 AND2X2_6371 ( .A(u5__abc_81276_new_n1170_), .B(u5__abc_81276_new_n3834_), .Y(u5__abc_81276_new_n3835_));
AND2X2 AND2X2_6372 ( .A(u5__abc_81276_new_n3215__bF_buf3), .B(u5_state_65_), .Y(u5__abc_81276_new_n3839_));
AND2X2 AND2X2_6373 ( .A(u5__abc_81276_new_n3840_), .B(u5__abc_81276_new_n3809_), .Y(u5__abc_81276_new_n3841_));
AND2X2 AND2X2_6374 ( .A(u5__abc_81276_new_n3842_), .B(u5__abc_81276_new_n3838_), .Y(u5_next_state_65_));
AND2X2 AND2X2_6375 ( .A(u5__abc_81276_new_n1315_), .B(u5__abc_81276_new_n3844_), .Y(u5__abc_81276_new_n3845_));
AND2X2 AND2X2_6376 ( .A(u5__abc_81276_new_n1324_), .B(u5__abc_81276_new_n1303_), .Y(u5__abc_81276_new_n3847_));
AND2X2 AND2X2_6377 ( .A(u5__abc_81276_new_n1593_), .B(u5__abc_81276_new_n3847_), .Y(u5__abc_81276_new_n3848_));
AND2X2 AND2X2_6378 ( .A(u5__abc_81276_new_n1255_), .B(u5__abc_81276_new_n1344_), .Y(u5__abc_81276_new_n3849_));
AND2X2 AND2X2_6379 ( .A(u5__abc_81276_new_n3848_), .B(u5__abc_81276_new_n3849_), .Y(u5__abc_81276_new_n3850_));
AND2X2 AND2X2_638 ( .A(u0__abc_76628_new_n2756_), .B(u0__abc_76628_new_n2719__bF_buf4), .Y(u0__abc_76628_new_n2757_));
AND2X2 AND2X2_6380 ( .A(u5__abc_81276_new_n2614_), .B(u5__abc_81276_new_n3850_), .Y(u5__abc_81276_new_n3851_));
AND2X2 AND2X2_6381 ( .A(u5__abc_81276_new_n1242_), .B(u5__abc_81276_new_n3851_), .Y(u5__abc_81276_new_n3852_));
AND2X2 AND2X2_6382 ( .A(u5__abc_81276_new_n2637_), .B(u5__abc_81276_new_n3852_), .Y(u5__abc_81276_new_n3853_));
AND2X2 AND2X2_6383 ( .A(u5__abc_81276_new_n3853_), .B(u5__abc_81276_new_n3846_), .Y(u5_pack_le0_d));
AND2X2 AND2X2_6384 ( .A(u5__abc_81276_new_n1836_), .B(u5__abc_81276_new_n1095_), .Y(u5__abc_81276_new_n3855_));
AND2X2 AND2X2_6385 ( .A(u5__abc_81276_new_n2569_), .B(u5__abc_81276_new_n854_), .Y(u5__abc_81276_new_n3859_));
AND2X2 AND2X2_6386 ( .A(u5__abc_81276_new_n3858_), .B(u5__abc_81276_new_n3859_), .Y(u5__abc_81276_new_n3860_));
AND2X2 AND2X2_6387 ( .A(u5__abc_81276_new_n3860_), .B(u5__abc_81276_new_n3857_), .Y(u5__abc_81276_new_n3861_));
AND2X2 AND2X2_6388 ( .A(u5__abc_81276_new_n3862_), .B(u5__abc_81276_new_n3863_), .Y(u5__abc_81276_new_n3864_));
AND2X2 AND2X2_6389 ( .A(u5__abc_81276_new_n853_), .B(u5__abc_81276_new_n3864_), .Y(u5__abc_81276_new_n3865_));
AND2X2 AND2X2_639 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2758_));
AND2X2 AND2X2_6390 ( .A(u5__abc_81276_new_n3866_), .B(u5__abc_81276_new_n603_), .Y(u5__abc_81276_new_n3867_));
AND2X2 AND2X2_6391 ( .A(u5__abc_81276_new_n589_), .B(u5__abc_81276_new_n3867_), .Y(u5__abc_81276_new_n3868_));
AND2X2 AND2X2_6392 ( .A(u5__abc_81276_new_n670_), .B(u5__abc_81276_new_n3868_), .Y(u5__abc_81276_new_n3869_));
AND2X2 AND2X2_6393 ( .A(u5__abc_81276_new_n3869_), .B(u5__abc_81276_new_n2567_), .Y(u5__abc_81276_new_n3870_));
AND2X2 AND2X2_6394 ( .A(u5__abc_81276_new_n3870_), .B(u5__abc_81276_new_n2827_), .Y(u5__abc_81276_new_n3871_));
AND2X2 AND2X2_6395 ( .A(u5__abc_81276_new_n3871_), .B(u5__abc_81276_new_n1897_), .Y(u5__abc_81276_new_n3872_));
AND2X2 AND2X2_6396 ( .A(u5__abc_81276_new_n1558_), .B(u5__abc_81276_new_n1550_), .Y(u5__abc_81276_new_n3876_));
AND2X2 AND2X2_6397 ( .A(u5__abc_81276_new_n1511_), .B(u5__abc_81276_new_n3876_), .Y(u5__abc_81276_new_n3877_));
AND2X2 AND2X2_6398 ( .A(u5__abc_81276_new_n3877_), .B(u5__abc_81276_new_n1357_), .Y(u5__abc_81276_new_n3878_));
AND2X2 AND2X2_6399 ( .A(u5__abc_81276_new_n3878_), .B(u5__abc_81276_new_n1520_), .Y(u5__abc_81276_new_n3879_));
AND2X2 AND2X2_64 ( .A(u0__abc_76628_new_n1105_), .B(u0__abc_76628_new_n1113_), .Y(u0__abc_76628_new_n1114_));
AND2X2 AND2X2_640 ( .A(u0__abc_76628_new_n2759_), .B(u0__abc_76628_new_n2718__bF_buf4), .Y(u0__abc_76628_new_n2760_));
AND2X2 AND2X2_6400 ( .A(u5__abc_81276_new_n3879_), .B(u5__abc_81276_new_n1913_), .Y(u5__abc_81276_new_n3880_));
AND2X2 AND2X2_6401 ( .A(u5__abc_81276_new_n3880_), .B(u5__abc_81276_new_n2459_), .Y(u5__abc_81276_new_n3881_));
AND2X2 AND2X2_6402 ( .A(u5__abc_81276_new_n2520_), .B(u5__abc_81276_new_n3881_), .Y(u5__abc_81276_new_n3882_));
AND2X2 AND2X2_6403 ( .A(u5__abc_81276_new_n1348_), .B(u5__abc_81276_new_n3882_), .Y(u5__abc_81276_new_n3883_));
AND2X2 AND2X2_6404 ( .A(u5__abc_81276_new_n3890_), .B(u5__abc_81276_new_n3891_), .Y(u5__abc_81276_new_n3892_));
AND2X2 AND2X2_6405 ( .A(u5__0no_wb_cycle_0_0_), .B(u5__abc_81276_new_n3892_), .Y(u5__abc_81276_new_n3893_));
AND2X2 AND2X2_6406 ( .A(u5__abc_81276_new_n3893_), .B(u5__abc_81276_new_n1558_), .Y(u5__abc_81276_new_n3894_));
AND2X2 AND2X2_6407 ( .A(u5__abc_81276_new_n1428_), .B(u5__abc_81276_new_n3894_), .Y(u5__abc_81276_new_n3895_));
AND2X2 AND2X2_6408 ( .A(u5__abc_81276_new_n1414_), .B(u5__abc_81276_new_n1480_), .Y(u5__abc_81276_new_n3896_));
AND2X2 AND2X2_6409 ( .A(u5__abc_81276_new_n1416_), .B(u5__abc_81276_new_n1398_), .Y(u5__abc_81276_new_n3897_));
AND2X2 AND2X2_641 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2761_));
AND2X2 AND2X2_6410 ( .A(u5__abc_81276_new_n2446_), .B(u5__abc_81276_new_n3897_), .Y(u5__abc_81276_new_n3898_));
AND2X2 AND2X2_6411 ( .A(u5__abc_81276_new_n2451_), .B(u5__abc_81276_new_n3898_), .Y(u5__abc_81276_new_n3899_));
AND2X2 AND2X2_6412 ( .A(u5__abc_81276_new_n3899_), .B(u5__abc_81276_new_n3896_), .Y(u5__abc_81276_new_n3900_));
AND2X2 AND2X2_6413 ( .A(u5__abc_81276_new_n3900_), .B(u5__abc_81276_new_n2459_), .Y(u5__abc_81276_new_n3901_));
AND2X2 AND2X2_6414 ( .A(u5__abc_81276_new_n2633_), .B(u5__abc_81276_new_n3901_), .Y(u5__abc_81276_new_n3902_));
AND2X2 AND2X2_6415 ( .A(u5__abc_81276_new_n3902_), .B(u5__abc_81276_new_n1348_), .Y(u5__abc_81276_new_n3903_));
AND2X2 AND2X2_6416 ( .A(u5__abc_81276_new_n1549_), .B(u5__abc_81276_new_n3325_), .Y(u5__abc_81276_new_n3906_));
AND2X2 AND2X2_6417 ( .A(u5__abc_81276_new_n3535_), .B(u5__abc_81276_new_n3907_), .Y(u5__abc_81276_new_n3908_));
AND2X2 AND2X2_6418 ( .A(u5__abc_81276_new_n1526__bF_buf1), .B(u5_wb_stb_first), .Y(u5__abc_81276_new_n3909_));
AND2X2 AND2X2_6419 ( .A(u5__abc_81276_new_n1536_), .B(u5_tmr_done_bF_buf2), .Y(u5__abc_81276_new_n3910_));
AND2X2 AND2X2_642 ( .A(u0__abc_76628_new_n2762_), .B(u0__abc_76628_new_n2717__bF_buf4), .Y(u0__abc_76628_new_n2763_));
AND2X2 AND2X2_6420 ( .A(u5__abc_81276_new_n1155_), .B(u5__abc_81276_new_n3910_), .Y(u5__abc_81276_new_n3911_));
AND2X2 AND2X2_6421 ( .A(u5__abc_81276_new_n1160_), .B(u5__abc_81276_new_n3222_), .Y(u5__abc_81276_new_n3912_));
AND2X2 AND2X2_6422 ( .A(u5__abc_81276_new_n3914_), .B(u5_wb_cycle), .Y(u5__abc_81276_new_n3915_));
AND2X2 AND2X2_6423 ( .A(u5__abc_81276_new_n1547_), .B(u5__abc_81276_new_n3229_), .Y(u5__abc_81276_new_n3916_));
AND2X2 AND2X2_6424 ( .A(u5__abc_81276_new_n3916_), .B(u5__abc_81276_new_n3374_), .Y(u5__abc_81276_new_n3917_));
AND2X2 AND2X2_6425 ( .A(u5__abc_81276_new_n624_), .B(u5__abc_81276_new_n3917_), .Y(u5__abc_81276_new_n3918_));
AND2X2 AND2X2_6426 ( .A(u5__abc_81276_new_n1526__bF_buf0), .B(u5__abc_81276_new_n3928_), .Y(u5__abc_81276_new_n3929_));
AND2X2 AND2X2_6427 ( .A(u5__abc_81276_new_n1361_), .B(rfr_ack), .Y(u5__abc_81276_new_n3947_));
AND2X2 AND2X2_6428 ( .A(u5__abc_81276_new_n3947_), .B(u5__abc_81276_new_n1429_), .Y(u5__abc_81276_new_n3948_));
AND2X2 AND2X2_6429 ( .A(u5__abc_81276_new_n3948_), .B(u5__abc_81276_new_n1770_), .Y(u5__abc_81276_new_n3949_));
AND2X2 AND2X2_643 ( .A(u0_tms1_1_), .B(u0_cs1_bF_buf3), .Y(u0__abc_76628_new_n2764_));
AND2X2 AND2X2_6430 ( .A(u5__abc_81276_new_n3949_), .B(u5__abc_81276_new_n2629_), .Y(u5__abc_81276_new_n3950_));
AND2X2 AND2X2_6431 ( .A(u5__abc_81276_new_n3950_), .B(u5__abc_81276_new_n2490_), .Y(u5__abc_81276_new_n3951_));
AND2X2 AND2X2_6432 ( .A(u5__abc_81276_new_n1348_), .B(u5__abc_81276_new_n1789_), .Y(u5__abc_81276_new_n3952_));
AND2X2 AND2X2_6433 ( .A(u5__abc_81276_new_n3952_), .B(u5__abc_81276_new_n3951_), .Y(u5__abc_81276_new_n3953_));
AND2X2 AND2X2_6434 ( .A(u5__abc_81276_new_n630_), .B(u5__abc_81276_new_n3957_), .Y(u5__abc_81276_new_n3958_));
AND2X2 AND2X2_6435 ( .A(u5__abc_81276_new_n1770_), .B(u5__abc_81276_new_n3958_), .Y(u5__abc_81276_new_n3959_));
AND2X2 AND2X2_6436 ( .A(u5__abc_81276_new_n2451_), .B(u5__abc_81276_new_n3959_), .Y(u5__abc_81276_new_n3960_));
AND2X2 AND2X2_6437 ( .A(u5__abc_81276_new_n1801_), .B(u5__abc_81276_new_n3960_), .Y(u5__abc_81276_new_n3961_));
AND2X2 AND2X2_6438 ( .A(u5__abc_81276_new_n3961_), .B(u5__abc_81276_new_n2631_), .Y(u5__abc_81276_new_n3962_));
AND2X2 AND2X2_6439 ( .A(u5__abc_81276_new_n3952_), .B(u5__abc_81276_new_n3962_), .Y(u5__abc_81276_new_n3963_));
AND2X2 AND2X2_644 ( .A(u0__abc_76628_new_n1169__bF_buf4), .B(u0__abc_76628_new_n2767_), .Y(u0__abc_76628_new_n2768_));
AND2X2 AND2X2_6440 ( .A(u5__abc_81276_new_n1316_), .B(u5__abc_81276_new_n3661_), .Y(u5__abc_81276_new_n3965_));
AND2X2 AND2X2_6441 ( .A(u5__abc_81276_new_n3965_), .B(u5__abc_81276_new_n1343_), .Y(u5__abc_81276_new_n3966_));
AND2X2 AND2X2_6442 ( .A(u5__abc_81276_new_n1596_), .B(u5__abc_81276_new_n1780_), .Y(u5__abc_81276_new_n3967_));
AND2X2 AND2X2_6443 ( .A(u5__abc_81276_new_n3967_), .B(u5__abc_81276_new_n3966_), .Y(u5__abc_81276_new_n3968_));
AND2X2 AND2X2_6444 ( .A(u5__abc_81276_new_n3968_), .B(u5__abc_81276_new_n1779_), .Y(u5__abc_81276_new_n3969_));
AND2X2 AND2X2_6445 ( .A(u5__abc_81276_new_n1571_), .B(u5__abc_81276_new_n1566_), .Y(u5__abc_81276_new_n3970_));
AND2X2 AND2X2_6446 ( .A(u5__abc_81276_new_n3970_), .B(u5__abc_81276_new_n1753_), .Y(u5__abc_81276_new_n3971_));
AND2X2 AND2X2_6447 ( .A(u5__abc_81276_new_n1241_), .B(u5__abc_81276_new_n3971_), .Y(u5__abc_81276_new_n3972_));
AND2X2 AND2X2_6448 ( .A(u5__abc_81276_new_n3972_), .B(u5__abc_81276_new_n3969_), .Y(u5__abc_81276_new_n3973_));
AND2X2 AND2X2_6449 ( .A(u5__abc_81276_new_n3973_), .B(u5__abc_81276_new_n1748_), .Y(u5__abc_81276_new_n3974_));
AND2X2 AND2X2_645 ( .A(u0__abc_76628_new_n2766_), .B(u0__abc_76628_new_n2768_), .Y(u0__abc_76628_new_n2769_));
AND2X2 AND2X2_6450 ( .A(u5__abc_81276_new_n3974_), .B(u5__abc_81276_new_n1805_), .Y(u5__abc_81276_new_n3975_));
AND2X2 AND2X2_6451 ( .A(u5__abc_81276_new_n3976_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3977_));
AND2X2 AND2X2_6452 ( .A(u5__abc_81276_new_n1467_), .B(u5__abc_81276_new_n1480_), .Y(u5__abc_81276_new_n3979_));
AND2X2 AND2X2_6453 ( .A(u5__abc_81276_new_n3979_), .B(u5__abc_81276_new_n2502_), .Y(u5__abc_81276_new_n3980_));
AND2X2 AND2X2_6454 ( .A(u5__abc_81276_new_n3980_), .B(u5__abc_81276_new_n2635_), .Y(u5__abc_81276_new_n3981_));
AND2X2 AND2X2_6455 ( .A(u5__abc_81276_new_n2866_), .B(u5__abc_81276_new_n3981_), .Y(u5__abc_81276_new_n3982_));
AND2X2 AND2X2_6456 ( .A(u5__abc_81276_new_n2635_), .B(u5__abc_81276_new_n1746_), .Y(u5__abc_81276_new_n3984_));
AND2X2 AND2X2_6457 ( .A(u5__abc_81276_new_n3984_), .B(u5__abc_81276_new_n2646_), .Y(u5__abc_81276_new_n3985_));
AND2X2 AND2X2_6458 ( .A(u5__abc_81276_new_n1273_), .B(u5__abc_81276_new_n1147_), .Y(u5__abc_81276_new_n3986_));
AND2X2 AND2X2_6459 ( .A(u5__abc_81276_new_n1161_), .B(u5__abc_81276_new_n1458_), .Y(u5__abc_81276_new_n3987_));
AND2X2 AND2X2_646 ( .A(u0__abc_76628_new_n1170__bF_buf4), .B(tms_2_), .Y(u0__abc_76628_new_n2771_));
AND2X2 AND2X2_6460 ( .A(u5__abc_81276_new_n3986_), .B(u5__abc_81276_new_n3987_), .Y(u5__abc_81276_new_n3988_));
AND2X2 AND2X2_6461 ( .A(u5__abc_81276_new_n1603_), .B(u5__abc_81276_new_n1780_), .Y(u5__abc_81276_new_n3989_));
AND2X2 AND2X2_6462 ( .A(u5__abc_81276_new_n1480_), .B(u5__abc_81276_new_n2647_), .Y(u5__abc_81276_new_n3990_));
AND2X2 AND2X2_6463 ( .A(u5__abc_81276_new_n3989_), .B(u5__abc_81276_new_n3990_), .Y(u5__abc_81276_new_n3991_));
AND2X2 AND2X2_6464 ( .A(u5__abc_81276_new_n3991_), .B(u5__abc_81276_new_n3988_), .Y(u5__abc_81276_new_n3992_));
AND2X2 AND2X2_6465 ( .A(u5__abc_81276_new_n2305_), .B(u5__abc_81276_new_n3992_), .Y(u5__abc_81276_new_n3993_));
AND2X2 AND2X2_6466 ( .A(u5__abc_81276_new_n3993_), .B(u5__abc_81276_new_n2494_), .Y(u5__abc_81276_new_n3994_));
AND2X2 AND2X2_6467 ( .A(u5__abc_81276_new_n3994_), .B(u5__abc_81276_new_n3985_), .Y(u5__abc_81276_new_n3995_));
AND2X2 AND2X2_6468 ( .A(u5__abc_81276_new_n1501_), .B(u5_cmd_a10_r), .Y(u5__abc_81276_new_n3996_));
AND2X2 AND2X2_6469 ( .A(u5__abc_81276_new_n3996_), .B(u5__abc_81276_new_n625_), .Y(u5__abc_81276_new_n3997_));
AND2X2 AND2X2_647 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2772_));
AND2X2 AND2X2_6470 ( .A(u5__abc_81276_new_n1571_), .B(u5__abc_81276_new_n1668_), .Y(u5__abc_81276_new_n3998_));
AND2X2 AND2X2_6471 ( .A(u5__abc_81276_new_n3998_), .B(u5__abc_81276_new_n3997_), .Y(u5__abc_81276_new_n3999_));
AND2X2 AND2X2_6472 ( .A(u5__abc_81276_new_n3999_), .B(u5__abc_81276_new_n1645_), .Y(u5__abc_81276_new_n4000_));
AND2X2 AND2X2_6473 ( .A(u5__abc_81276_new_n3995_), .B(u5__abc_81276_new_n4000_), .Y(u5__abc_81276_new_n4001_));
AND2X2 AND2X2_6474 ( .A(u5__abc_81276_new_n1668_), .B(u5__abc_81276_new_n3353_), .Y(u5__abc_81276_new_n4006_));
AND2X2 AND2X2_6475 ( .A(u5__abc_81276_new_n4006_), .B(u5__abc_81276_new_n4005_), .Y(u5__abc_81276_new_n4007_));
AND2X2 AND2X2_6476 ( .A(u5__abc_81276_new_n4008_), .B(u5__abc_81276_new_n3238_), .Y(u5__abc_81276_new_n4009_));
AND2X2 AND2X2_6477 ( .A(u5__abc_81276_new_n1450_), .B(u5__abc_81276_new_n4010_), .Y(u5__abc_81276_new_n4011_));
AND2X2 AND2X2_6478 ( .A(u5__abc_81276_new_n1668_), .B(u5__abc_81276_new_n1493_), .Y(u5__abc_81276_new_n4013_));
AND2X2 AND2X2_6479 ( .A(u5__abc_81276_new_n4013_), .B(u5__abc_81276_new_n4012_), .Y(u5__abc_81276_new_n4014_));
AND2X2 AND2X2_648 ( .A(u0__abc_76628_new_n2774_), .B(u0__abc_76628_new_n2724__bF_buf3), .Y(u0__abc_76628_new_n2775_));
AND2X2 AND2X2_6480 ( .A(u5__abc_81276_new_n1588_), .B(u5_cmd_a10_r), .Y(u5__abc_81276_new_n4016_));
AND2X2 AND2X2_6481 ( .A(u5__abc_81276_new_n1500_), .B(rfr_ack), .Y(u5__abc_81276_new_n4018_));
AND2X2 AND2X2_6482 ( .A(u5__abc_81276_new_n1645_), .B(u5__abc_81276_new_n4019_), .Y(u5__abc_81276_new_n4020_));
AND2X2 AND2X2_6483 ( .A(u5__abc_81276_new_n4020_), .B(u5__abc_81276_new_n4017_), .Y(u5__abc_81276_new_n4021_));
AND2X2 AND2X2_6484 ( .A(u5__abc_81276_new_n4015_), .B(u5__abc_81276_new_n4021_), .Y(u5__abc_81276_new_n4022_));
AND2X2 AND2X2_6485 ( .A(u5__abc_81276_new_n4003_), .B(u5__abc_81276_new_n4022_), .Y(u5__abc_81276_new_n4023_));
AND2X2 AND2X2_6486 ( .A(u5__abc_81276_new_n4023_), .B(u5__abc_81276_new_n4002_), .Y(u5__abc_81276_new_n4024_));
AND2X2 AND2X2_6487 ( .A(u5__abc_81276_new_n1148_), .B(u5__abc_81276_new_n1254_), .Y(u5__abc_81276_new_n4028_));
AND2X2 AND2X2_6488 ( .A(u5__abc_81276_new_n4028_), .B(u5__abc_81276_new_n1208_), .Y(u5__abc_81276_new_n4029_));
AND2X2 AND2X2_6489 ( .A(u5__abc_81276_new_n1346_), .B(u5__abc_81276_new_n4029_), .Y(u5__abc_81276_new_n4030_));
AND2X2 AND2X2_649 ( .A(u0__abc_76628_new_n2775_), .B(u0__abc_76628_new_n2773_), .Y(u0__abc_76628_new_n2776_));
AND2X2 AND2X2_6490 ( .A(u5__abc_81276_new_n4027_), .B(u5__abc_81276_new_n4030_), .Y(u5__abc_81276_new_n4031_));
AND2X2 AND2X2_6491 ( .A(u5__abc_81276_new_n4031_), .B(u5__abc_81276_new_n4026_), .Y(u5__0oe__0_0_));
AND2X2 AND2X2_6492 ( .A(u5__abc_81276_new_n1595_), .B(u5__abc_81276_new_n1378_), .Y(u5__abc_81276_new_n4033_));
AND2X2 AND2X2_6493 ( .A(u5__abc_81276_new_n4033_), .B(u5__abc_81276_new_n1593_), .Y(u5__abc_81276_new_n4034_));
AND2X2 AND2X2_6494 ( .A(u5__abc_81276_new_n4034_), .B(u5__abc_81276_new_n1345_), .Y(u5__abc_81276_new_n4035_));
AND2X2 AND2X2_6495 ( .A(u5__abc_81276_new_n4035_), .B(u5__abc_81276_new_n1241_), .Y(u5__abc_81276_new_n4036_));
AND2X2 AND2X2_6496 ( .A(u5__abc_81276_new_n1748_), .B(u5__abc_81276_new_n4036_), .Y(u5__abc_81276_new_n4037_));
AND2X2 AND2X2_6497 ( .A(u5__abc_81276_new_n1790_), .B(u5__abc_81276_new_n4037_), .Y(u5_pack_le1_d));
AND2X2 AND2X2_6498 ( .A(u5__abc_81276_new_n1133_), .B(u5__abc_81276_new_n1171_), .Y(u5__abc_81276_new_n4039_));
AND2X2 AND2X2_6499 ( .A(u5__abc_81276_new_n2665_), .B(u5__abc_81276_new_n4039_), .Y(u5__abc_81276_new_n4040_));
AND2X2 AND2X2_65 ( .A(u0__abc_76628_new_n1109_), .B(spec_req_cs_2_bF_buf4_), .Y(u0__abc_76628_new_n1116_));
AND2X2 AND2X2_650 ( .A(u0__abc_76628_new_n2777_), .B(u0__abc_76628_new_n2720__bF_buf3), .Y(u0__abc_76628_new_n2778_));
AND2X2 AND2X2_6500 ( .A(u5__abc_81276_new_n1791_), .B(u5__abc_81276_new_n4040_), .Y(err));
AND2X2 AND2X2_6501 ( .A(u5__abc_81276_new_n2459_), .B(u5__abc_81276_new_n2449_), .Y(u5__abc_81276_new_n4042_));
AND2X2 AND2X2_6502 ( .A(u5__abc_81276_new_n2520_), .B(u5__abc_81276_new_n4042_), .Y(u5__abc_81276_new_n4043_));
AND2X2 AND2X2_6503 ( .A(u5__abc_81276_new_n1348_), .B(u5__abc_81276_new_n4043_), .Y(init_ack));
AND2X2 AND2X2_6504 ( .A(u5_wb_cycle), .B(u5_cnt), .Y(u5__abc_81276_new_n4045_));
AND2X2 AND2X2_6505 ( .A(u5__abc_81276_new_n1836_), .B(u5__abc_81276_new_n4045_), .Y(u5__abc_81276_new_n4046_));
AND2X2 AND2X2_6506 ( .A(u5__abc_81276_new_n4049_), .B(u5__abc_81276_new_n572_), .Y(u5__abc_81276_new_n4050_));
AND2X2 AND2X2_6507 ( .A(u5__abc_81276_new_n4050_), .B(u5__abc_81276_new_n4048_), .Y(u5__abc_81276_new_n4051_));
AND2X2 AND2X2_6508 ( .A(u5__abc_81276_new_n4059_), .B(u5_cke_r), .Y(u5__0cke__0_0_));
AND2X2 AND2X2_6509 ( .A(wb_stb_i_bF_buf4), .B(wb_cyc_i), .Y(u5__abc_81276_new_n4061_));
AND2X2 AND2X2_651 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2779_));
AND2X2 AND2X2_6510 ( .A(u5__abc_81276_new_n4061_), .B(cs_le_bF_buf2), .Y(u5__0lookup_ready1_0_0_));
AND2X2 AND2X2_6511 ( .A(u5__abc_81276_new_n4061_), .B(u5_lookup_ready1), .Y(u5__0lookup_ready2_0_0_));
AND2X2 AND2X2_6512 ( .A(u5__abc_81276_new_n3100_), .B(u5__abc_81276_new_n4064_), .Y(u5__abc_81276_new_n4065_));
AND2X2 AND2X2_6513 ( .A(u5__abc_81276_new_n4065_), .B(u5__abc_81276_new_n3034_), .Y(u5__abc_81276_new_n4066_));
AND2X2 AND2X2_6514 ( .A(u5__abc_81276_new_n4066_), .B(u5__abc_81276_new_n2926_), .Y(u5__abc_81276_new_n4067_));
AND2X2 AND2X2_6515 ( .A(u5__abc_81276_new_n2970_), .B(u5__abc_81276_new_n2932_), .Y(u5__abc_81276_new_n4068_));
AND2X2 AND2X2_6516 ( .A(u5__abc_81276_new_n4068_), .B(u5__abc_81276_new_n4067_), .Y(u5__0tmr2_done_0_0_));
AND2X2 AND2X2_6517 ( .A(u5__abc_81276_new_n3592_), .B(u5__abc_81276_new_n1553_), .Y(u5__abc_81276_new_n4070_));
AND2X2 AND2X2_6518 ( .A(u5__abc_81276_new_n4079_), .B(susp_sel), .Y(u5__abc_81276_new_n4080_));
AND2X2 AND2X2_6519 ( .A(u5_wb_cycle), .B(wb_cyc_i), .Y(u5__abc_81276_new_n4083_));
AND2X2 AND2X2_652 ( .A(u0__abc_76628_new_n2780_), .B(u0__abc_76628_new_n2719__bF_buf3), .Y(u0__abc_76628_new_n2781_));
AND2X2 AND2X2_6520 ( .A(u5__abc_81276_new_n4083_), .B(u5__abc_81276_new_n4082_), .Y(u5__abc_81276_new_n4084_));
AND2X2 AND2X2_6521 ( .A(u5__abc_81276_new_n1689_), .B(u5__abc_81276_new_n3330_), .Y(u5__abc_81276_new_n4088_));
AND2X2 AND2X2_6522 ( .A(u5__abc_81276_new_n4089_), .B(u5__abc_81276_new_n4086_), .Y(u5__abc_81276_new_n4090_));
AND2X2 AND2X2_6523 ( .A(u5__abc_81276_new_n2320_), .B(u1_wr_cycle), .Y(u5__abc_81276_new_n4091_));
AND2X2 AND2X2_6524 ( .A(wb_cyc_i), .B(wb_stb_i_bF_buf3), .Y(u6__abc_85257_new_n133_));
AND2X2 AND2X2_6525 ( .A(u6__abc_85257_new_n136_), .B(u6__abc_85257_new_n137_), .Y(u6__abc_85257_new_n138_));
AND2X2 AND2X2_6526 ( .A(u6__abc_85257_new_n138_), .B(u6__abc_85257_new_n135_), .Y(u6__abc_85257_new_n139_));
AND2X2 AND2X2_6527 ( .A(u6__abc_85257_new_n142_), .B(u6__abc_85257_new_n143_), .Y(u6__abc_85257_new_n144_));
AND2X2 AND2X2_6528 ( .A(u6__abc_85257_new_n144_), .B(u6__abc_85257_new_n141_), .Y(u6__abc_85257_new_n145_));
AND2X2 AND2X2_6529 ( .A(u6__abc_85257_new_n145__bF_buf5), .B(mem_ack), .Y(u6__abc_85257_new_n146_));
AND2X2 AND2X2_653 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2782_));
AND2X2 AND2X2_6530 ( .A(u6__abc_85257_new_n140_), .B(u6__abc_85257_new_n146_), .Y(u6__abc_85257_new_n147_));
AND2X2 AND2X2_6531 ( .A(u6__abc_85257_new_n141_), .B(\wb_addr_i[29] ), .Y(u6__abc_85257_new_n148_));
AND2X2 AND2X2_6532 ( .A(u6__abc_85257_new_n149_), .B(\wb_addr_i[30] ), .Y(u6__abc_85257_new_n150_));
AND2X2 AND2X2_6533 ( .A(u6__abc_85257_new_n150_), .B(u6__abc_85257_new_n133_), .Y(u6__abc_85257_new_n151_));
AND2X2 AND2X2_6534 ( .A(u6__abc_85257_new_n151_), .B(u6__abc_85257_new_n148_), .Y(u6__abc_85257_new_n152_));
AND2X2 AND2X2_6535 ( .A(u6__abc_85257_new_n156_), .B(u6__abc_85257_new_n154_), .Y(u6__0wb_data_o_31_0__0_));
AND2X2 AND2X2_6536 ( .A(u6__abc_85257_new_n159_), .B(u6__abc_85257_new_n158_), .Y(u6__0wb_data_o_31_0__1_));
AND2X2 AND2X2_6537 ( .A(u6__abc_85257_new_n162_), .B(u6__abc_85257_new_n161_), .Y(u6__0wb_data_o_31_0__2_));
AND2X2 AND2X2_6538 ( .A(u6__abc_85257_new_n165_), .B(u6__abc_85257_new_n164_), .Y(u6__0wb_data_o_31_0__3_));
AND2X2 AND2X2_6539 ( .A(u6__abc_85257_new_n168_), .B(u6__abc_85257_new_n167_), .Y(u6__0wb_data_o_31_0__4_));
AND2X2 AND2X2_654 ( .A(u0__abc_76628_new_n2783_), .B(u0__abc_76628_new_n2718__bF_buf3), .Y(u0__abc_76628_new_n2784_));
AND2X2 AND2X2_6540 ( .A(u6__abc_85257_new_n171_), .B(u6__abc_85257_new_n170_), .Y(u6__0wb_data_o_31_0__5_));
AND2X2 AND2X2_6541 ( .A(u6__abc_85257_new_n174_), .B(u6__abc_85257_new_n173_), .Y(u6__0wb_data_o_31_0__6_));
AND2X2 AND2X2_6542 ( .A(u6__abc_85257_new_n177_), .B(u6__abc_85257_new_n176_), .Y(u6__0wb_data_o_31_0__7_));
AND2X2 AND2X2_6543 ( .A(u6__abc_85257_new_n180_), .B(u6__abc_85257_new_n179_), .Y(u6__0wb_data_o_31_0__8_));
AND2X2 AND2X2_6544 ( .A(u6__abc_85257_new_n183_), .B(u6__abc_85257_new_n182_), .Y(u6__0wb_data_o_31_0__9_));
AND2X2 AND2X2_6545 ( .A(u6__abc_85257_new_n186_), .B(u6__abc_85257_new_n185_), .Y(u6__0wb_data_o_31_0__10_));
AND2X2 AND2X2_6546 ( .A(u6__abc_85257_new_n189_), .B(u6__abc_85257_new_n188_), .Y(u6__0wb_data_o_31_0__11_));
AND2X2 AND2X2_6547 ( .A(u6__abc_85257_new_n192_), .B(u6__abc_85257_new_n191_), .Y(u6__0wb_data_o_31_0__12_));
AND2X2 AND2X2_6548 ( .A(u6__abc_85257_new_n195_), .B(u6__abc_85257_new_n194_), .Y(u6__0wb_data_o_31_0__13_));
AND2X2 AND2X2_6549 ( .A(u6__abc_85257_new_n198_), .B(u6__abc_85257_new_n197_), .Y(u6__0wb_data_o_31_0__14_));
AND2X2 AND2X2_655 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2785_));
AND2X2 AND2X2_6550 ( .A(u6__abc_85257_new_n201_), .B(u6__abc_85257_new_n200_), .Y(u6__0wb_data_o_31_0__15_));
AND2X2 AND2X2_6551 ( .A(u6__abc_85257_new_n204_), .B(u6__abc_85257_new_n203_), .Y(u6__0wb_data_o_31_0__16_));
AND2X2 AND2X2_6552 ( .A(u6__abc_85257_new_n207_), .B(u6__abc_85257_new_n206_), .Y(u6__0wb_data_o_31_0__17_));
AND2X2 AND2X2_6553 ( .A(u6__abc_85257_new_n210_), .B(u6__abc_85257_new_n209_), .Y(u6__0wb_data_o_31_0__18_));
AND2X2 AND2X2_6554 ( .A(u6__abc_85257_new_n213_), .B(u6__abc_85257_new_n212_), .Y(u6__0wb_data_o_31_0__19_));
AND2X2 AND2X2_6555 ( .A(u6__abc_85257_new_n216_), .B(u6__abc_85257_new_n215_), .Y(u6__0wb_data_o_31_0__20_));
AND2X2 AND2X2_6556 ( .A(u6__abc_85257_new_n219_), .B(u6__abc_85257_new_n218_), .Y(u6__0wb_data_o_31_0__21_));
AND2X2 AND2X2_6557 ( .A(u6__abc_85257_new_n222_), .B(u6__abc_85257_new_n221_), .Y(u6__0wb_data_o_31_0__22_));
AND2X2 AND2X2_6558 ( .A(u6__abc_85257_new_n225_), .B(u6__abc_85257_new_n224_), .Y(u6__0wb_data_o_31_0__23_));
AND2X2 AND2X2_6559 ( .A(u6__abc_85257_new_n228_), .B(u6__abc_85257_new_n227_), .Y(u6__0wb_data_o_31_0__24_));
AND2X2 AND2X2_656 ( .A(u0__abc_76628_new_n2786_), .B(u0__abc_76628_new_n2717__bF_buf3), .Y(u0__abc_76628_new_n2787_));
AND2X2 AND2X2_6560 ( .A(u6__abc_85257_new_n231_), .B(u6__abc_85257_new_n230_), .Y(u6__0wb_data_o_31_0__25_));
AND2X2 AND2X2_6561 ( .A(u6__abc_85257_new_n234_), .B(u6__abc_85257_new_n233_), .Y(u6__0wb_data_o_31_0__26_));
AND2X2 AND2X2_6562 ( .A(u6__abc_85257_new_n237_), .B(u6__abc_85257_new_n236_), .Y(u6__0wb_data_o_31_0__27_));
AND2X2 AND2X2_6563 ( .A(u6__abc_85257_new_n240_), .B(u6__abc_85257_new_n239_), .Y(u6__0wb_data_o_31_0__28_));
AND2X2 AND2X2_6564 ( .A(u6__abc_85257_new_n243_), .B(u6__abc_85257_new_n242_), .Y(u6__0wb_data_o_31_0__29_));
AND2X2 AND2X2_6565 ( .A(u6__abc_85257_new_n246_), .B(u6__abc_85257_new_n245_), .Y(u6__0wb_data_o_31_0__30_));
AND2X2 AND2X2_6566 ( .A(u6__abc_85257_new_n249_), .B(u6__abc_85257_new_n248_), .Y(u6__0wb_data_o_31_0__31_));
AND2X2 AND2X2_6567 ( .A(u6__abc_85257_new_n133_), .B(wb_we_i), .Y(u6__abc_85257_new_n251_));
AND2X2 AND2X2_6568 ( .A(u6__abc_85257_new_n134_), .B(u1_wr_hold), .Y(u6__abc_85257_new_n252_));
AND2X2 AND2X2_6569 ( .A(u6__abc_85257_new_n254_), .B(u6_rmw_en), .Y(u6__abc_85257_new_n255_));
AND2X2 AND2X2_657 ( .A(u0_tms1_2_), .B(u0_cs1_bF_buf2), .Y(u0__abc_76628_new_n2788_));
AND2X2 AND2X2_6570 ( .A(u6__abc_85257_new_n251_), .B(u6__abc_85257_new_n255_), .Y(u6__0rmw_r_0_0_));
AND2X2 AND2X2_6571 ( .A(u6__abc_85257_new_n145__bF_buf1), .B(wb_stb_i_bF_buf2), .Y(u6__abc_85257_new_n258_));
AND2X2 AND2X2_6572 ( .A(u6__abc_85257_new_n258_), .B(u6__abc_85257_new_n257_), .Y(u6__abc_85257_new_n259_));
AND2X2 AND2X2_6573 ( .A(u6__abc_85257_new_n262_), .B(u6__abc_85257_new_n261_), .Y(u6__abc_85257_new_n263_));
AND2X2 AND2X2_6574 ( .A(u6__abc_85257_new_n263_), .B(wb_cyc_i), .Y(u6__abc_85257_new_n264_));
AND2X2 AND2X2_6575 ( .A(u6__abc_85257_new_n260_), .B(u6__abc_85257_new_n264_), .Y(u6__0read_go_r1_0_0_));
AND2X2 AND2X2_6576 ( .A(wb_cyc_i), .B(u6_read_go_r1), .Y(u6__0read_go_r_0_0_));
AND2X2 AND2X2_6577 ( .A(u6__abc_85257_new_n263_), .B(u6__0read_go_r_0_0_), .Y(u3_wb_read_go));
AND2X2 AND2X2_6578 ( .A(u6__abc_85257_new_n258_), .B(wb_we_i), .Y(u6__abc_85257_new_n268_));
AND2X2 AND2X2_6579 ( .A(u6__abc_85257_new_n269_), .B(wb_cyc_i), .Y(u6__0write_go_r1_0_0_));
AND2X2 AND2X2_658 ( .A(u0__abc_76628_new_n1169__bF_buf3), .B(u0__abc_76628_new_n2791_), .Y(u0__abc_76628_new_n2792_));
AND2X2 AND2X2_6580 ( .A(wb_cyc_i), .B(u6_write_go_r1), .Y(u6__abc_85257_new_n273_));
AND2X2 AND2X2_6581 ( .A(u6__abc_85257_new_n272_), .B(u6__abc_85257_new_n273_), .Y(u6__0write_go_r_0_0_));
AND2X2 AND2X2_6582 ( .A(u6__abc_85257_new_n263_), .B(u6__0write_go_r_0_0_), .Y(u1_wb_write_go));
AND2X2 AND2X2_6583 ( .A(u6__abc_85257_new_n276_), .B(u6__abc_85257_new_n277_), .Y(u6__abc_85257_new_n278_));
AND2X2 AND2X2_6584 ( .A(u6__abc_85257_new_n278_), .B(u6__abc_85257_new_n133_), .Y(u6__abc_85257_new_n279_));
AND2X2 AND2X2_6585 ( .A(u6__abc_85257_new_n145__bF_buf0), .B(u6__abc_85257_new_n279_), .Y(u6__abc_85257_new_n280_));
AND2X2 AND2X2_6586 ( .A(u6__abc_85257_new_n149_), .B(u6_wb_first_r), .Y(u6__abc_85257_new_n282_));
AND2X2 AND2X2_6587 ( .A(u6__abc_85257_new_n282_), .B(u6__abc_85257_new_n281_), .Y(u6__abc_85257_new_n283_));
AND2X2 AND2X2_6588 ( .A(u6__abc_85257_new_n145__bF_buf5), .B(u6__abc_85257_new_n281_), .Y(u6__abc_85257_new_n286_));
AND2X2 AND2X2_6589 ( .A(u6__abc_85257_new_n285_), .B(u6__abc_85257_new_n286_), .Y(u6__0wb_err_0_0_));
AND2X2 AND2X2_659 ( .A(u0__abc_76628_new_n2790_), .B(u0__abc_76628_new_n2792_), .Y(u0__abc_76628_new_n2793_));
AND2X2 AND2X2_6590 ( .A(u6__abc_85257_new_n271_), .B(wb_cyc_i), .Y(u6__abc_85257_new_n289_));
AND2X2 AND2X2_6591 ( .A(u6__abc_85257_new_n288_), .B(u6__abc_85257_new_n289_), .Y(u5_wb_wait));
AND2X2 AND2X2_6592 ( .A(wb_cyc_i), .B(u6_rmw_en), .Y(u6__abc_85257_new_n291_));
AND2X2 AND2X2_6593 ( .A(u7__abc_74830_new_n75_), .B(data_oe), .Y(u7__abc_74830_new_n76_));
AND2X2 AND2X2_6594 ( .A(u7__abc_74830_new_n79_), .B(u7__abc_74830_new_n77_), .Y(u7__abc_74830_new_n80_));
AND2X2 AND2X2_6595 ( .A(u7__abc_74830_new_n83_), .B(data_oe), .Y(u7__abc_74830_new_n84_));
AND2X2 AND2X2_6596 ( .A(u7__abc_74830_new_n86_), .B(data_oe), .Y(u7__abc_74830_new_n87_));
AND2X2 AND2X2_6597 ( .A(u7__abc_74830_new_n89_), .B(data_oe), .Y(u7__abc_74830_new_n90_));
AND2X2 AND2X2_6598 ( .A(wb_stb_i_bF_buf0), .B(wb_cyc_i), .Y(u7__abc_74830_new_n92_));
AND2X2 AND2X2_6599 ( .A(u7__abc_74830_new_n92_), .B(\wb_sel_i[0] ), .Y(u7__abc_74830_new_n93_));
AND2X2 AND2X2_66 ( .A(u0__abc_76628_new_n1100_), .B(1'h0), .Y(u0__abc_76628_new_n1117_));
AND2X2 AND2X2_660 ( .A(u0__abc_76628_new_n1170__bF_buf3), .B(tms_3_), .Y(u0__abc_76628_new_n2795_));
AND2X2 AND2X2_6600 ( .A(u7__abc_74830_new_n94_), .B(u7_mc_dqm_r_0_), .Y(u7__abc_74830_new_n95_));
AND2X2 AND2X2_6601 ( .A(u7__abc_74830_new_n92_), .B(\wb_sel_i[1] ), .Y(u7__abc_74830_new_n97_));
AND2X2 AND2X2_6602 ( .A(u7__abc_74830_new_n94_), .B(u7_mc_dqm_r_1_), .Y(u7__abc_74830_new_n98_));
AND2X2 AND2X2_6603 ( .A(u7__abc_74830_new_n92_), .B(\wb_sel_i[2] ), .Y(u7__abc_74830_new_n100_));
AND2X2 AND2X2_6604 ( .A(u7__abc_74830_new_n94_), .B(u7_mc_dqm_r_2_), .Y(u7__abc_74830_new_n101_));
AND2X2 AND2X2_6605 ( .A(u7__abc_74830_new_n92_), .B(\wb_sel_i[3] ), .Y(u7__abc_74830_new_n103_));
AND2X2 AND2X2_6606 ( .A(u7__abc_74830_new_n94_), .B(u7_mc_dqm_r_3_), .Y(u7__abc_74830_new_n104_));
AND2X2 AND2X2_6607 ( .A(spec_req_cs_0_bF_buf5_), .B(lmr_sel_bF_buf1), .Y(u7__abc_74830_new_n110_));
AND2X2 AND2X2_6608 ( .A(u7__abc_74830_new_n109_), .B(u7__abc_74830_new_n111_), .Y(u7__abc_74830_new_n112_));
AND2X2 AND2X2_6609 ( .A(u7__abc_74830_new_n112_), .B(u7__abc_74830_new_n107_), .Y(u7__abc_74830_new_n113_));
AND2X2 AND2X2_661 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2796_));
AND2X2 AND2X2_6610 ( .A(u7__abc_74830_new_n106_), .B(u7__abc_74830_new_n115_), .Y(u7__abc_74830_new_n116_));
AND2X2 AND2X2_6611 ( .A(lmr_sel_bF_buf6), .B(spec_req_cs_1_bF_buf5_), .Y(u7__abc_74830_new_n121_));
AND2X2 AND2X2_6612 ( .A(u7__abc_74830_new_n120_), .B(u7__abc_74830_new_n122_), .Y(u7__abc_74830_new_n123_));
AND2X2 AND2X2_6613 ( .A(u7__abc_74830_new_n123_), .B(u7__abc_74830_new_n107_), .Y(u7__abc_74830_new_n124_));
AND2X2 AND2X2_6614 ( .A(u7__abc_74830_new_n106_), .B(u7__abc_74830_new_n125_), .Y(u7__abc_74830_new_n126_));
AND2X2 AND2X2_6615 ( .A(lmr_sel_bF_buf4), .B(spec_req_cs_2_bF_buf1_), .Y(u7__abc_74830_new_n131_));
AND2X2 AND2X2_6616 ( .A(u7__abc_74830_new_n130_), .B(u7__abc_74830_new_n132_), .Y(u7__abc_74830_new_n133_));
AND2X2 AND2X2_6617 ( .A(u7__abc_74830_new_n133_), .B(u7__abc_74830_new_n107_), .Y(u7__abc_74830_new_n134_));
AND2X2 AND2X2_6618 ( .A(u7__abc_74830_new_n106_), .B(u7__abc_74830_new_n135_), .Y(u7__abc_74830_new_n136_));
AND2X2 AND2X2_6619 ( .A(lmr_sel_bF_buf2), .B(spec_req_cs_3_bF_buf1_), .Y(u7__abc_74830_new_n141_));
AND2X2 AND2X2_662 ( .A(u0__abc_76628_new_n2798_), .B(u0__abc_76628_new_n2724__bF_buf2), .Y(u0__abc_76628_new_n2799_));
AND2X2 AND2X2_6620 ( .A(u7__abc_74830_new_n140_), .B(u7__abc_74830_new_n142_), .Y(u7__abc_74830_new_n143_));
AND2X2 AND2X2_6621 ( .A(u7__abc_74830_new_n143_), .B(u7__abc_74830_new_n107_), .Y(u7__abc_74830_new_n144_));
AND2X2 AND2X2_6622 ( .A(u7__abc_74830_new_n106_), .B(u7__abc_74830_new_n145_), .Y(u7__abc_74830_new_n146_));
AND2X2 AND2X2_6623 ( .A(lmr_sel_bF_buf0), .B(spec_req_cs_4_bF_buf1_), .Y(u7__abc_74830_new_n151_));
AND2X2 AND2X2_6624 ( .A(u7__abc_74830_new_n150_), .B(u7__abc_74830_new_n152_), .Y(u7__abc_74830_new_n153_));
AND2X2 AND2X2_6625 ( .A(u7__abc_74830_new_n153_), .B(u7__abc_74830_new_n107_), .Y(u7__abc_74830_new_n154_));
AND2X2 AND2X2_6626 ( .A(u7__abc_74830_new_n106_), .B(u7__abc_74830_new_n155_), .Y(u7__abc_74830_new_n156_));
AND2X2 AND2X2_6627 ( .A(lmr_sel_bF_buf5), .B(spec_req_cs_5_bF_buf1_), .Y(u7__abc_74830_new_n161_));
AND2X2 AND2X2_6628 ( .A(u7__abc_74830_new_n160_), .B(u7__abc_74830_new_n162_), .Y(u7__abc_74830_new_n163_));
AND2X2 AND2X2_6629 ( .A(u7__abc_74830_new_n163_), .B(u7__abc_74830_new_n107_), .Y(u7__abc_74830_new_n164_));
AND2X2 AND2X2_663 ( .A(u0__abc_76628_new_n2799_), .B(u0__abc_76628_new_n2797_), .Y(u0__abc_76628_new_n2800_));
AND2X2 AND2X2_6630 ( .A(u7__abc_74830_new_n106_), .B(u7__abc_74830_new_n165_), .Y(u7__abc_74830_new_n166_));
AND2X2 AND2X2_6631 ( .A(lmr_sel_bF_buf3), .B(spec_req_cs_6_bF_buf1_), .Y(u7__abc_74830_new_n171_));
AND2X2 AND2X2_6632 ( .A(u7__abc_74830_new_n170_), .B(u7__abc_74830_new_n172_), .Y(u7__abc_74830_new_n173_));
AND2X2 AND2X2_6633 ( .A(u7__abc_74830_new_n173_), .B(u7__abc_74830_new_n107_), .Y(u7__abc_74830_new_n174_));
AND2X2 AND2X2_6634 ( .A(u7__abc_74830_new_n106_), .B(u7__abc_74830_new_n175_), .Y(u7__abc_74830_new_n176_));
AND2X2 AND2X2_6635 ( .A(lmr_sel_bF_buf1), .B(spec_req_cs_7_), .Y(u7__abc_74830_new_n181_));
AND2X2 AND2X2_6636 ( .A(u7__abc_74830_new_n180_), .B(u7__abc_74830_new_n182_), .Y(u7__abc_74830_new_n183_));
AND2X2 AND2X2_6637 ( .A(u7__abc_74830_new_n183_), .B(u7__abc_74830_new_n107_), .Y(u7__abc_74830_new_n184_));
AND2X2 AND2X2_6638 ( .A(u7__abc_74830_new_n106_), .B(u7__abc_74830_new_n185_), .Y(u7__abc_74830_new_n186_));
AND2X2 AND2X2_6639 ( .A(u7__abc_74830_new_n191_), .B(u7__abc_74830_new_n192_), .Y(u7__0mc_rp_0_0_));
AND2X2 AND2X2_664 ( .A(u0__abc_76628_new_n2801_), .B(u0__abc_76628_new_n2720__bF_buf2), .Y(u0__abc_76628_new_n2802_));
AND2X2 AND2X2_6640 ( .A(data_oe), .B(mc_c_oe_d), .Y(u7__abc_74830_new_n195_));
AND2X2 AND2X2_6641 ( .A(u7__abc_74830_new_n195_), .B(u7__abc_74830_new_n194_), .Y(u7__0mc_data_oe_0_0_));
AND2X2 AND2X2_665 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2803_));
AND2X2 AND2X2_666 ( .A(u0__abc_76628_new_n2804_), .B(u0__abc_76628_new_n2719__bF_buf2), .Y(u0__abc_76628_new_n2805_));
AND2X2 AND2X2_667 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2806_));
AND2X2 AND2X2_668 ( .A(u0__abc_76628_new_n2807_), .B(u0__abc_76628_new_n2718__bF_buf2), .Y(u0__abc_76628_new_n2808_));
AND2X2 AND2X2_669 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2809_));
AND2X2 AND2X2_67 ( .A(init_req), .B(1'h0), .Y(u0__abc_76628_new_n1118_));
AND2X2 AND2X2_670 ( .A(u0__abc_76628_new_n2810_), .B(u0__abc_76628_new_n2717__bF_buf2), .Y(u0__abc_76628_new_n2811_));
AND2X2 AND2X2_671 ( .A(u0_tms1_3_), .B(u0_cs1_bF_buf1), .Y(u0__abc_76628_new_n2812_));
AND2X2 AND2X2_672 ( .A(u0__abc_76628_new_n1169__bF_buf2), .B(u0__abc_76628_new_n2815_), .Y(u0__abc_76628_new_n2816_));
AND2X2 AND2X2_673 ( .A(u0__abc_76628_new_n2814_), .B(u0__abc_76628_new_n2816_), .Y(u0__abc_76628_new_n2817_));
AND2X2 AND2X2_674 ( .A(u0__abc_76628_new_n1170__bF_buf2), .B(tms_4_), .Y(u0__abc_76628_new_n2819_));
AND2X2 AND2X2_675 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2820_));
AND2X2 AND2X2_676 ( .A(u0__abc_76628_new_n2822_), .B(u0__abc_76628_new_n2724__bF_buf1), .Y(u0__abc_76628_new_n2823_));
AND2X2 AND2X2_677 ( .A(u0__abc_76628_new_n2823_), .B(u0__abc_76628_new_n2821_), .Y(u0__abc_76628_new_n2824_));
AND2X2 AND2X2_678 ( .A(u0__abc_76628_new_n2825_), .B(u0__abc_76628_new_n2720__bF_buf1), .Y(u0__abc_76628_new_n2826_));
AND2X2 AND2X2_679 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2827_));
AND2X2 AND2X2_68 ( .A(u0__abc_76628_new_n1105_), .B(u0__abc_76628_new_n1120_), .Y(u0__abc_76628_new_n1121_));
AND2X2 AND2X2_680 ( .A(u0__abc_76628_new_n2828_), .B(u0__abc_76628_new_n2719__bF_buf1), .Y(u0__abc_76628_new_n2829_));
AND2X2 AND2X2_681 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2830_));
AND2X2 AND2X2_682 ( .A(u0__abc_76628_new_n2831_), .B(u0__abc_76628_new_n2718__bF_buf1), .Y(u0__abc_76628_new_n2832_));
AND2X2 AND2X2_683 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2833_));
AND2X2 AND2X2_684 ( .A(u0__abc_76628_new_n2834_), .B(u0__abc_76628_new_n2717__bF_buf1), .Y(u0__abc_76628_new_n2835_));
AND2X2 AND2X2_685 ( .A(u0_tms1_4_), .B(u0_cs1_bF_buf0), .Y(u0__abc_76628_new_n2836_));
AND2X2 AND2X2_686 ( .A(u0__abc_76628_new_n1169__bF_buf1), .B(u0__abc_76628_new_n2839_), .Y(u0__abc_76628_new_n2840_));
AND2X2 AND2X2_687 ( .A(u0__abc_76628_new_n2838_), .B(u0__abc_76628_new_n2840_), .Y(u0__abc_76628_new_n2841_));
AND2X2 AND2X2_688 ( .A(u0__abc_76628_new_n1170__bF_buf1), .B(tms_5_), .Y(u0__abc_76628_new_n2843_));
AND2X2 AND2X2_689 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2844_));
AND2X2 AND2X2_69 ( .A(u0__abc_76628_new_n1121_), .B(u0__abc_76628_new_n1119_), .Y(u0__abc_76628_new_n1122_));
AND2X2 AND2X2_690 ( .A(u0__abc_76628_new_n2846_), .B(u0__abc_76628_new_n2724__bF_buf0), .Y(u0__abc_76628_new_n2847_));
AND2X2 AND2X2_691 ( .A(u0__abc_76628_new_n2847_), .B(u0__abc_76628_new_n2845_), .Y(u0__abc_76628_new_n2848_));
AND2X2 AND2X2_692 ( .A(u0__abc_76628_new_n2849_), .B(u0__abc_76628_new_n2720__bF_buf0), .Y(u0__abc_76628_new_n2850_));
AND2X2 AND2X2_693 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2851_));
AND2X2 AND2X2_694 ( .A(u0__abc_76628_new_n2852_), .B(u0__abc_76628_new_n2719__bF_buf0), .Y(u0__abc_76628_new_n2853_));
AND2X2 AND2X2_695 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2854_));
AND2X2 AND2X2_696 ( .A(u0__abc_76628_new_n2855_), .B(u0__abc_76628_new_n2718__bF_buf0), .Y(u0__abc_76628_new_n2856_));
AND2X2 AND2X2_697 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2857_));
AND2X2 AND2X2_698 ( .A(u0__abc_76628_new_n2858_), .B(u0__abc_76628_new_n2717__bF_buf0), .Y(u0__abc_76628_new_n2859_));
AND2X2 AND2X2_699 ( .A(u0_tms1_5_), .B(u0_cs1_bF_buf5), .Y(u0__abc_76628_new_n2860_));
AND2X2 AND2X2_7 ( .A(_abc_85006_new_n257_), .B(_abc_85006_new_n258_), .Y(obct_cs_2_));
AND2X2 AND2X2_70 ( .A(u0__abc_76628_new_n1109_), .B(spec_req_cs_3_bF_buf4_), .Y(u0__abc_76628_new_n1124_));
AND2X2 AND2X2_700 ( .A(u0__abc_76628_new_n1169__bF_buf0), .B(u0__abc_76628_new_n2863_), .Y(u0__abc_76628_new_n2864_));
AND2X2 AND2X2_701 ( .A(u0__abc_76628_new_n2862_), .B(u0__abc_76628_new_n2864_), .Y(u0__abc_76628_new_n2865_));
AND2X2 AND2X2_702 ( .A(u0__abc_76628_new_n1170__bF_buf0), .B(tms_6_), .Y(u0__abc_76628_new_n2867_));
AND2X2 AND2X2_703 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2868_));
AND2X2 AND2X2_704 ( .A(u0__abc_76628_new_n2870_), .B(u0__abc_76628_new_n2724__bF_buf5), .Y(u0__abc_76628_new_n2871_));
AND2X2 AND2X2_705 ( .A(u0__abc_76628_new_n2871_), .B(u0__abc_76628_new_n2869_), .Y(u0__abc_76628_new_n2872_));
AND2X2 AND2X2_706 ( .A(u0__abc_76628_new_n2873_), .B(u0__abc_76628_new_n2720__bF_buf5), .Y(u0__abc_76628_new_n2874_));
AND2X2 AND2X2_707 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2875_));
AND2X2 AND2X2_708 ( .A(u0__abc_76628_new_n2876_), .B(u0__abc_76628_new_n2719__bF_buf5), .Y(u0__abc_76628_new_n2877_));
AND2X2 AND2X2_709 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2878_));
AND2X2 AND2X2_71 ( .A(u0__abc_76628_new_n1100_), .B(1'h0), .Y(u0__abc_76628_new_n1126_));
AND2X2 AND2X2_710 ( .A(u0__abc_76628_new_n2879_), .B(u0__abc_76628_new_n2718__bF_buf5), .Y(u0__abc_76628_new_n2880_));
AND2X2 AND2X2_711 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2881_));
AND2X2 AND2X2_712 ( .A(u0__abc_76628_new_n2882_), .B(u0__abc_76628_new_n2717__bF_buf5), .Y(u0__abc_76628_new_n2883_));
AND2X2 AND2X2_713 ( .A(u0_tms1_6_), .B(u0_cs1_bF_buf4), .Y(u0__abc_76628_new_n2884_));
AND2X2 AND2X2_714 ( .A(u0__abc_76628_new_n1169__bF_buf6), .B(u0__abc_76628_new_n2887_), .Y(u0__abc_76628_new_n2888_));
AND2X2 AND2X2_715 ( .A(u0__abc_76628_new_n2886_), .B(u0__abc_76628_new_n2888_), .Y(u0__abc_76628_new_n2889_));
AND2X2 AND2X2_716 ( .A(u0__abc_76628_new_n1170__bF_buf6), .B(tms_7_), .Y(u0__abc_76628_new_n2891_));
AND2X2 AND2X2_717 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2892_));
AND2X2 AND2X2_718 ( .A(u0__abc_76628_new_n2894_), .B(u0__abc_76628_new_n2724__bF_buf4), .Y(u0__abc_76628_new_n2895_));
AND2X2 AND2X2_719 ( .A(u0__abc_76628_new_n2895_), .B(u0__abc_76628_new_n2893_), .Y(u0__abc_76628_new_n2896_));
AND2X2 AND2X2_72 ( .A(init_req), .B(1'h0), .Y(u0__abc_76628_new_n1127_));
AND2X2 AND2X2_720 ( .A(u0__abc_76628_new_n2897_), .B(u0__abc_76628_new_n2720__bF_buf4), .Y(u0__abc_76628_new_n2898_));
AND2X2 AND2X2_721 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2899_));
AND2X2 AND2X2_722 ( .A(u0__abc_76628_new_n2900_), .B(u0__abc_76628_new_n2719__bF_buf4), .Y(u0__abc_76628_new_n2901_));
AND2X2 AND2X2_723 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2902_));
AND2X2 AND2X2_724 ( .A(u0__abc_76628_new_n2903_), .B(u0__abc_76628_new_n2718__bF_buf4), .Y(u0__abc_76628_new_n2904_));
AND2X2 AND2X2_725 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2905_));
AND2X2 AND2X2_726 ( .A(u0__abc_76628_new_n2906_), .B(u0__abc_76628_new_n2717__bF_buf4), .Y(u0__abc_76628_new_n2907_));
AND2X2 AND2X2_727 ( .A(u0_tms1_7_), .B(u0_cs1_bF_buf3), .Y(u0__abc_76628_new_n2908_));
AND2X2 AND2X2_728 ( .A(u0__abc_76628_new_n1169__bF_buf5), .B(u0__abc_76628_new_n2911_), .Y(u0__abc_76628_new_n2912_));
AND2X2 AND2X2_729 ( .A(u0__abc_76628_new_n2910_), .B(u0__abc_76628_new_n2912_), .Y(u0__abc_76628_new_n2913_));
AND2X2 AND2X2_73 ( .A(u0__abc_76628_new_n1125_), .B(u0__abc_76628_new_n1128_), .Y(u0__abc_76628_new_n1129_));
AND2X2 AND2X2_730 ( .A(u0__abc_76628_new_n1170__bF_buf5), .B(tms_8_), .Y(u0__abc_76628_new_n2915_));
AND2X2 AND2X2_731 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2916_));
AND2X2 AND2X2_732 ( .A(u0__abc_76628_new_n2918_), .B(u0__abc_76628_new_n2724__bF_buf3), .Y(u0__abc_76628_new_n2919_));
AND2X2 AND2X2_733 ( .A(u0__abc_76628_new_n2919_), .B(u0__abc_76628_new_n2917_), .Y(u0__abc_76628_new_n2920_));
AND2X2 AND2X2_734 ( .A(u0__abc_76628_new_n2921_), .B(u0__abc_76628_new_n2720__bF_buf3), .Y(u0__abc_76628_new_n2922_));
AND2X2 AND2X2_735 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2923_));
AND2X2 AND2X2_736 ( .A(u0__abc_76628_new_n2924_), .B(u0__abc_76628_new_n2719__bF_buf3), .Y(u0__abc_76628_new_n2925_));
AND2X2 AND2X2_737 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2926_));
AND2X2 AND2X2_738 ( .A(u0__abc_76628_new_n2927_), .B(u0__abc_76628_new_n2718__bF_buf3), .Y(u0__abc_76628_new_n2928_));
AND2X2 AND2X2_739 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2929_));
AND2X2 AND2X2_74 ( .A(u0__abc_76628_new_n1121_), .B(u0__abc_76628_new_n1129_), .Y(u0__abc_76628_new_n1130_));
AND2X2 AND2X2_740 ( .A(u0__abc_76628_new_n2930_), .B(u0__abc_76628_new_n2717__bF_buf3), .Y(u0__abc_76628_new_n2931_));
AND2X2 AND2X2_741 ( .A(u0_tms1_8_), .B(u0_cs1_bF_buf2), .Y(u0__abc_76628_new_n2932_));
AND2X2 AND2X2_742 ( .A(u0__abc_76628_new_n1169__bF_buf4), .B(u0__abc_76628_new_n2935_), .Y(u0__abc_76628_new_n2936_));
AND2X2 AND2X2_743 ( .A(u0__abc_76628_new_n2934_), .B(u0__abc_76628_new_n2936_), .Y(u0__abc_76628_new_n2937_));
AND2X2 AND2X2_744 ( .A(u0__abc_76628_new_n1170__bF_buf4), .B(tms_9_), .Y(u0__abc_76628_new_n2939_));
AND2X2 AND2X2_745 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2940_));
AND2X2 AND2X2_746 ( .A(u0__abc_76628_new_n2942_), .B(u0__abc_76628_new_n2724__bF_buf2), .Y(u0__abc_76628_new_n2943_));
AND2X2 AND2X2_747 ( .A(u0__abc_76628_new_n2943_), .B(u0__abc_76628_new_n2941_), .Y(u0__abc_76628_new_n2944_));
AND2X2 AND2X2_748 ( .A(u0__abc_76628_new_n2945_), .B(u0__abc_76628_new_n2720__bF_buf2), .Y(u0__abc_76628_new_n2946_));
AND2X2 AND2X2_749 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2947_));
AND2X2 AND2X2_75 ( .A(u0__abc_76628_new_n1109_), .B(spec_req_cs_4_bF_buf4_), .Y(u0__abc_76628_new_n1132_));
AND2X2 AND2X2_750 ( .A(u0__abc_76628_new_n2948_), .B(u0__abc_76628_new_n2719__bF_buf2), .Y(u0__abc_76628_new_n2949_));
AND2X2 AND2X2_751 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2950_));
AND2X2 AND2X2_752 ( .A(u0__abc_76628_new_n2951_), .B(u0__abc_76628_new_n2718__bF_buf2), .Y(u0__abc_76628_new_n2952_));
AND2X2 AND2X2_753 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2953_));
AND2X2 AND2X2_754 ( .A(u0__abc_76628_new_n2954_), .B(u0__abc_76628_new_n2717__bF_buf2), .Y(u0__abc_76628_new_n2955_));
AND2X2 AND2X2_755 ( .A(u0_tms1_9_), .B(u0_cs1_bF_buf1), .Y(u0__abc_76628_new_n2956_));
AND2X2 AND2X2_756 ( .A(u0__abc_76628_new_n1169__bF_buf3), .B(u0__abc_76628_new_n2959_), .Y(u0__abc_76628_new_n2960_));
AND2X2 AND2X2_757 ( .A(u0__abc_76628_new_n2958_), .B(u0__abc_76628_new_n2960_), .Y(u0__abc_76628_new_n2961_));
AND2X2 AND2X2_758 ( .A(u0__abc_76628_new_n1170__bF_buf3), .B(tms_10_), .Y(u0__abc_76628_new_n2963_));
AND2X2 AND2X2_759 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2964_));
AND2X2 AND2X2_76 ( .A(u0__abc_76628_new_n1100_), .B(1'h0), .Y(u0__abc_76628_new_n1133_));
AND2X2 AND2X2_760 ( .A(u0__abc_76628_new_n2966_), .B(u0__abc_76628_new_n2724__bF_buf1), .Y(u0__abc_76628_new_n2967_));
AND2X2 AND2X2_761 ( .A(u0__abc_76628_new_n2967_), .B(u0__abc_76628_new_n2965_), .Y(u0__abc_76628_new_n2968_));
AND2X2 AND2X2_762 ( .A(u0__abc_76628_new_n2969_), .B(u0__abc_76628_new_n2720__bF_buf1), .Y(u0__abc_76628_new_n2970_));
AND2X2 AND2X2_763 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2971_));
AND2X2 AND2X2_764 ( .A(u0__abc_76628_new_n2972_), .B(u0__abc_76628_new_n2719__bF_buf1), .Y(u0__abc_76628_new_n2973_));
AND2X2 AND2X2_765 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2974_));
AND2X2 AND2X2_766 ( .A(u0__abc_76628_new_n2975_), .B(u0__abc_76628_new_n2718__bF_buf1), .Y(u0__abc_76628_new_n2976_));
AND2X2 AND2X2_767 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2977_));
AND2X2 AND2X2_768 ( .A(u0__abc_76628_new_n2978_), .B(u0__abc_76628_new_n2717__bF_buf1), .Y(u0__abc_76628_new_n2979_));
AND2X2 AND2X2_769 ( .A(u0_tms1_10_), .B(u0_cs1_bF_buf0), .Y(u0__abc_76628_new_n2980_));
AND2X2 AND2X2_77 ( .A(init_req), .B(1'h0), .Y(u0__abc_76628_new_n1134_));
AND2X2 AND2X2_770 ( .A(u0__abc_76628_new_n1169__bF_buf2), .B(u0__abc_76628_new_n2983_), .Y(u0__abc_76628_new_n2984_));
AND2X2 AND2X2_771 ( .A(u0__abc_76628_new_n2982_), .B(u0__abc_76628_new_n2984_), .Y(u0__abc_76628_new_n2985_));
AND2X2 AND2X2_772 ( .A(u0__abc_76628_new_n1170__bF_buf2), .B(tms_11_), .Y(u0__abc_76628_new_n2987_));
AND2X2 AND2X2_773 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2988_));
AND2X2 AND2X2_774 ( .A(u0__abc_76628_new_n2990_), .B(u0__abc_76628_new_n2724__bF_buf0), .Y(u0__abc_76628_new_n2991_));
AND2X2 AND2X2_775 ( .A(u0__abc_76628_new_n2991_), .B(u0__abc_76628_new_n2989_), .Y(u0__abc_76628_new_n2992_));
AND2X2 AND2X2_776 ( .A(u0__abc_76628_new_n2993_), .B(u0__abc_76628_new_n2720__bF_buf0), .Y(u0__abc_76628_new_n2994_));
AND2X2 AND2X2_777 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2995_));
AND2X2 AND2X2_778 ( .A(u0__abc_76628_new_n2996_), .B(u0__abc_76628_new_n2719__bF_buf0), .Y(u0__abc_76628_new_n2997_));
AND2X2 AND2X2_779 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2998_));
AND2X2 AND2X2_78 ( .A(u0__abc_76628_new_n1125_), .B(u0__abc_76628_new_n1136_), .Y(u0__abc_76628_new_n1137_));
AND2X2 AND2X2_780 ( .A(u0__abc_76628_new_n2999_), .B(u0__abc_76628_new_n2718__bF_buf0), .Y(u0__abc_76628_new_n3000_));
AND2X2 AND2X2_781 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3001_));
AND2X2 AND2X2_782 ( .A(u0__abc_76628_new_n3002_), .B(u0__abc_76628_new_n2717__bF_buf0), .Y(u0__abc_76628_new_n3003_));
AND2X2 AND2X2_783 ( .A(u0_tms1_11_), .B(u0_cs1_bF_buf5), .Y(u0__abc_76628_new_n3004_));
AND2X2 AND2X2_784 ( .A(u0__abc_76628_new_n1169__bF_buf1), .B(u0__abc_76628_new_n3007_), .Y(u0__abc_76628_new_n3008_));
AND2X2 AND2X2_785 ( .A(u0__abc_76628_new_n3006_), .B(u0__abc_76628_new_n3008_), .Y(u0__abc_76628_new_n3009_));
AND2X2 AND2X2_786 ( .A(u0__abc_76628_new_n1170__bF_buf1), .B(tms_12_), .Y(u0__abc_76628_new_n3011_));
AND2X2 AND2X2_787 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3012_));
AND2X2 AND2X2_788 ( .A(u0__abc_76628_new_n3014_), .B(u0__abc_76628_new_n2724__bF_buf5), .Y(u0__abc_76628_new_n3015_));
AND2X2 AND2X2_789 ( .A(u0__abc_76628_new_n3015_), .B(u0__abc_76628_new_n3013_), .Y(u0__abc_76628_new_n3016_));
AND2X2 AND2X2_79 ( .A(u0__abc_76628_new_n1121_), .B(u0__abc_76628_new_n1137_), .Y(u0__abc_76628_new_n1138_));
AND2X2 AND2X2_790 ( .A(u0__abc_76628_new_n3017_), .B(u0__abc_76628_new_n2720__bF_buf5), .Y(u0__abc_76628_new_n3018_));
AND2X2 AND2X2_791 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3019_));
AND2X2 AND2X2_792 ( .A(u0__abc_76628_new_n3020_), .B(u0__abc_76628_new_n2719__bF_buf5), .Y(u0__abc_76628_new_n3021_));
AND2X2 AND2X2_793 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3022_));
AND2X2 AND2X2_794 ( .A(u0__abc_76628_new_n3023_), .B(u0__abc_76628_new_n2718__bF_buf5), .Y(u0__abc_76628_new_n3024_));
AND2X2 AND2X2_795 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3025_));
AND2X2 AND2X2_796 ( .A(u0__abc_76628_new_n3026_), .B(u0__abc_76628_new_n2717__bF_buf5), .Y(u0__abc_76628_new_n3027_));
AND2X2 AND2X2_797 ( .A(u0_tms1_12_), .B(u0_cs1_bF_buf4), .Y(u0__abc_76628_new_n3028_));
AND2X2 AND2X2_798 ( .A(u0__abc_76628_new_n1169__bF_buf0), .B(u0__abc_76628_new_n3031_), .Y(u0__abc_76628_new_n3032_));
AND2X2 AND2X2_799 ( .A(u0__abc_76628_new_n3030_), .B(u0__abc_76628_new_n3032_), .Y(u0__abc_76628_new_n3033_));
AND2X2 AND2X2_8 ( .A(_abc_85006_new_n260_), .B(_abc_85006_new_n261_), .Y(_abc_85006_new_n262_));
AND2X2 AND2X2_80 ( .A(u0__abc_76628_new_n1138_), .B(u0__abc_76628_new_n1135_), .Y(u0__abc_76628_new_n1139_));
AND2X2 AND2X2_800 ( .A(u0__abc_76628_new_n1170__bF_buf0), .B(tms_13_), .Y(u0__abc_76628_new_n3035_));
AND2X2 AND2X2_801 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3036_));
AND2X2 AND2X2_802 ( .A(u0__abc_76628_new_n3038_), .B(u0__abc_76628_new_n2724__bF_buf4), .Y(u0__abc_76628_new_n3039_));
AND2X2 AND2X2_803 ( .A(u0__abc_76628_new_n3039_), .B(u0__abc_76628_new_n3037_), .Y(u0__abc_76628_new_n3040_));
AND2X2 AND2X2_804 ( .A(u0__abc_76628_new_n3041_), .B(u0__abc_76628_new_n2720__bF_buf4), .Y(u0__abc_76628_new_n3042_));
AND2X2 AND2X2_805 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3043_));
AND2X2 AND2X2_806 ( .A(u0__abc_76628_new_n3044_), .B(u0__abc_76628_new_n2719__bF_buf4), .Y(u0__abc_76628_new_n3045_));
AND2X2 AND2X2_807 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3046_));
AND2X2 AND2X2_808 ( .A(u0__abc_76628_new_n3047_), .B(u0__abc_76628_new_n2718__bF_buf4), .Y(u0__abc_76628_new_n3048_));
AND2X2 AND2X2_809 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3049_));
AND2X2 AND2X2_81 ( .A(u0__abc_76628_new_n1109_), .B(spec_req_cs_5_bF_buf4_), .Y(u0__abc_76628_new_n1141_));
AND2X2 AND2X2_810 ( .A(u0__abc_76628_new_n3050_), .B(u0__abc_76628_new_n2717__bF_buf4), .Y(u0__abc_76628_new_n3051_));
AND2X2 AND2X2_811 ( .A(u0_tms1_13_), .B(u0_cs1_bF_buf3), .Y(u0__abc_76628_new_n3052_));
AND2X2 AND2X2_812 ( .A(u0__abc_76628_new_n1169__bF_buf6), .B(u0__abc_76628_new_n3055_), .Y(u0__abc_76628_new_n3056_));
AND2X2 AND2X2_813 ( .A(u0__abc_76628_new_n3054_), .B(u0__abc_76628_new_n3056_), .Y(u0__abc_76628_new_n3057_));
AND2X2 AND2X2_814 ( .A(u0__abc_76628_new_n1170__bF_buf6), .B(tms_14_), .Y(u0__abc_76628_new_n3059_));
AND2X2 AND2X2_815 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3060_));
AND2X2 AND2X2_816 ( .A(u0__abc_76628_new_n3062_), .B(u0__abc_76628_new_n2724__bF_buf3), .Y(u0__abc_76628_new_n3063_));
AND2X2 AND2X2_817 ( .A(u0__abc_76628_new_n3063_), .B(u0__abc_76628_new_n3061_), .Y(u0__abc_76628_new_n3064_));
AND2X2 AND2X2_818 ( .A(u0__abc_76628_new_n3065_), .B(u0__abc_76628_new_n2720__bF_buf3), .Y(u0__abc_76628_new_n3066_));
AND2X2 AND2X2_819 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3067_));
AND2X2 AND2X2_82 ( .A(u0__abc_76628_new_n1100_), .B(1'h0), .Y(u0__abc_76628_new_n1143_));
AND2X2 AND2X2_820 ( .A(u0__abc_76628_new_n3068_), .B(u0__abc_76628_new_n2719__bF_buf3), .Y(u0__abc_76628_new_n3069_));
AND2X2 AND2X2_821 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3070_));
AND2X2 AND2X2_822 ( .A(u0__abc_76628_new_n3071_), .B(u0__abc_76628_new_n2718__bF_buf3), .Y(u0__abc_76628_new_n3072_));
AND2X2 AND2X2_823 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3073_));
AND2X2 AND2X2_824 ( .A(u0__abc_76628_new_n3074_), .B(u0__abc_76628_new_n2717__bF_buf3), .Y(u0__abc_76628_new_n3075_));
AND2X2 AND2X2_825 ( .A(u0_tms1_14_), .B(u0_cs1_bF_buf2), .Y(u0__abc_76628_new_n3076_));
AND2X2 AND2X2_826 ( .A(u0__abc_76628_new_n1169__bF_buf5), .B(u0__abc_76628_new_n3079_), .Y(u0__abc_76628_new_n3080_));
AND2X2 AND2X2_827 ( .A(u0__abc_76628_new_n3078_), .B(u0__abc_76628_new_n3080_), .Y(u0__abc_76628_new_n3081_));
AND2X2 AND2X2_828 ( .A(u0__abc_76628_new_n1170__bF_buf5), .B(tms_15_), .Y(u0__abc_76628_new_n3083_));
AND2X2 AND2X2_829 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3084_));
AND2X2 AND2X2_83 ( .A(init_req), .B(1'h0), .Y(u0__abc_76628_new_n1144_));
AND2X2 AND2X2_830 ( .A(u0__abc_76628_new_n3086_), .B(u0__abc_76628_new_n2724__bF_buf2), .Y(u0__abc_76628_new_n3087_));
AND2X2 AND2X2_831 ( .A(u0__abc_76628_new_n3087_), .B(u0__abc_76628_new_n3085_), .Y(u0__abc_76628_new_n3088_));
AND2X2 AND2X2_832 ( .A(u0__abc_76628_new_n3089_), .B(u0__abc_76628_new_n2720__bF_buf2), .Y(u0__abc_76628_new_n3090_));
AND2X2 AND2X2_833 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3091_));
AND2X2 AND2X2_834 ( .A(u0__abc_76628_new_n3092_), .B(u0__abc_76628_new_n2719__bF_buf2), .Y(u0__abc_76628_new_n3093_));
AND2X2 AND2X2_835 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3094_));
AND2X2 AND2X2_836 ( .A(u0__abc_76628_new_n3095_), .B(u0__abc_76628_new_n2718__bF_buf2), .Y(u0__abc_76628_new_n3096_));
AND2X2 AND2X2_837 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3097_));
AND2X2 AND2X2_838 ( .A(u0__abc_76628_new_n3098_), .B(u0__abc_76628_new_n2717__bF_buf2), .Y(u0__abc_76628_new_n3099_));
AND2X2 AND2X2_839 ( .A(u0_tms1_15_), .B(u0_cs1_bF_buf1), .Y(u0__abc_76628_new_n3100_));
AND2X2 AND2X2_84 ( .A(u0__abc_76628_new_n1142_), .B(u0__abc_76628_new_n1145_), .Y(u0__abc_76628_new_n1146_));
AND2X2 AND2X2_840 ( .A(u0__abc_76628_new_n1169__bF_buf4), .B(u0__abc_76628_new_n3103_), .Y(u0__abc_76628_new_n3104_));
AND2X2 AND2X2_841 ( .A(u0__abc_76628_new_n3102_), .B(u0__abc_76628_new_n3104_), .Y(u0__abc_76628_new_n3105_));
AND2X2 AND2X2_842 ( .A(u0__abc_76628_new_n1170__bF_buf4), .B(tms_16_), .Y(u0__abc_76628_new_n3107_));
AND2X2 AND2X2_843 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3108_));
AND2X2 AND2X2_844 ( .A(u0__abc_76628_new_n3110_), .B(u0__abc_76628_new_n2724__bF_buf1), .Y(u0__abc_76628_new_n3111_));
AND2X2 AND2X2_845 ( .A(u0__abc_76628_new_n3111_), .B(u0__abc_76628_new_n3109_), .Y(u0__abc_76628_new_n3112_));
AND2X2 AND2X2_846 ( .A(u0__abc_76628_new_n3113_), .B(u0__abc_76628_new_n2720__bF_buf1), .Y(u0__abc_76628_new_n3114_));
AND2X2 AND2X2_847 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3115_));
AND2X2 AND2X2_848 ( .A(u0__abc_76628_new_n3116_), .B(u0__abc_76628_new_n2719__bF_buf1), .Y(u0__abc_76628_new_n3117_));
AND2X2 AND2X2_849 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3118_));
AND2X2 AND2X2_85 ( .A(u0__abc_76628_new_n1138_), .B(u0__abc_76628_new_n1146_), .Y(u0__abc_76628_new_n1147_));
AND2X2 AND2X2_850 ( .A(u0__abc_76628_new_n3119_), .B(u0__abc_76628_new_n2718__bF_buf1), .Y(u0__abc_76628_new_n3120_));
AND2X2 AND2X2_851 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3121_));
AND2X2 AND2X2_852 ( .A(u0__abc_76628_new_n3122_), .B(u0__abc_76628_new_n2717__bF_buf1), .Y(u0__abc_76628_new_n3123_));
AND2X2 AND2X2_853 ( .A(u0_tms1_16_), .B(u0_cs1_bF_buf0), .Y(u0__abc_76628_new_n3124_));
AND2X2 AND2X2_854 ( .A(u0__abc_76628_new_n1169__bF_buf3), .B(u0__abc_76628_new_n3127_), .Y(u0__abc_76628_new_n3128_));
AND2X2 AND2X2_855 ( .A(u0__abc_76628_new_n3126_), .B(u0__abc_76628_new_n3128_), .Y(u0__abc_76628_new_n3129_));
AND2X2 AND2X2_856 ( .A(u0__abc_76628_new_n1170__bF_buf3), .B(tms_17_), .Y(u0__abc_76628_new_n3131_));
AND2X2 AND2X2_857 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3132_));
AND2X2 AND2X2_858 ( .A(u0__abc_76628_new_n3134_), .B(u0__abc_76628_new_n2724__bF_buf0), .Y(u0__abc_76628_new_n3135_));
AND2X2 AND2X2_859 ( .A(u0__abc_76628_new_n3135_), .B(u0__abc_76628_new_n3133_), .Y(u0__abc_76628_new_n3136_));
AND2X2 AND2X2_86 ( .A(u0__abc_76628_new_n1109_), .B(spec_req_cs_6_bF_buf4_), .Y(u0__abc_76628_new_n1149_));
AND2X2 AND2X2_860 ( .A(u0__abc_76628_new_n3137_), .B(u0__abc_76628_new_n2720__bF_buf0), .Y(u0__abc_76628_new_n3138_));
AND2X2 AND2X2_861 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3139_));
AND2X2 AND2X2_862 ( .A(u0__abc_76628_new_n3140_), .B(u0__abc_76628_new_n2719__bF_buf0), .Y(u0__abc_76628_new_n3141_));
AND2X2 AND2X2_863 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3142_));
AND2X2 AND2X2_864 ( .A(u0__abc_76628_new_n3143_), .B(u0__abc_76628_new_n2718__bF_buf0), .Y(u0__abc_76628_new_n3144_));
AND2X2 AND2X2_865 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3145_));
AND2X2 AND2X2_866 ( .A(u0__abc_76628_new_n3146_), .B(u0__abc_76628_new_n2717__bF_buf0), .Y(u0__abc_76628_new_n3147_));
AND2X2 AND2X2_867 ( .A(u0_tms1_17_), .B(u0_cs1_bF_buf5), .Y(u0__abc_76628_new_n3148_));
AND2X2 AND2X2_868 ( .A(u0__abc_76628_new_n1169__bF_buf2), .B(u0__abc_76628_new_n3151_), .Y(u0__abc_76628_new_n3152_));
AND2X2 AND2X2_869 ( .A(u0__abc_76628_new_n3150_), .B(u0__abc_76628_new_n3152_), .Y(u0__abc_76628_new_n3153_));
AND2X2 AND2X2_87 ( .A(u0__abc_76628_new_n1100_), .B(1'h0), .Y(u0__abc_76628_new_n1150_));
AND2X2 AND2X2_870 ( .A(u0__abc_76628_new_n1170__bF_buf2), .B(tms_18_), .Y(u0__abc_76628_new_n3155_));
AND2X2 AND2X2_871 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3156_));
AND2X2 AND2X2_872 ( .A(u0__abc_76628_new_n3158_), .B(u0__abc_76628_new_n2724__bF_buf5), .Y(u0__abc_76628_new_n3159_));
AND2X2 AND2X2_873 ( .A(u0__abc_76628_new_n3159_), .B(u0__abc_76628_new_n3157_), .Y(u0__abc_76628_new_n3160_));
AND2X2 AND2X2_874 ( .A(u0__abc_76628_new_n3161_), .B(u0__abc_76628_new_n2720__bF_buf5), .Y(u0__abc_76628_new_n3162_));
AND2X2 AND2X2_875 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3163_));
AND2X2 AND2X2_876 ( .A(u0__abc_76628_new_n3164_), .B(u0__abc_76628_new_n2719__bF_buf5), .Y(u0__abc_76628_new_n3165_));
AND2X2 AND2X2_877 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3166_));
AND2X2 AND2X2_878 ( .A(u0__abc_76628_new_n3167_), .B(u0__abc_76628_new_n2718__bF_buf5), .Y(u0__abc_76628_new_n3168_));
AND2X2 AND2X2_879 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3169_));
AND2X2 AND2X2_88 ( .A(init_req), .B(1'h0), .Y(u0__abc_76628_new_n1151_));
AND2X2 AND2X2_880 ( .A(u0__abc_76628_new_n3170_), .B(u0__abc_76628_new_n2717__bF_buf5), .Y(u0__abc_76628_new_n3171_));
AND2X2 AND2X2_881 ( .A(u0_tms1_18_), .B(u0_cs1_bF_buf4), .Y(u0__abc_76628_new_n3172_));
AND2X2 AND2X2_882 ( .A(u0__abc_76628_new_n1169__bF_buf1), .B(u0__abc_76628_new_n3175_), .Y(u0__abc_76628_new_n3176_));
AND2X2 AND2X2_883 ( .A(u0__abc_76628_new_n3174_), .B(u0__abc_76628_new_n3176_), .Y(u0__abc_76628_new_n3177_));
AND2X2 AND2X2_884 ( .A(u0__abc_76628_new_n1170__bF_buf1), .B(tms_19_), .Y(u0__abc_76628_new_n3179_));
AND2X2 AND2X2_885 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3180_));
AND2X2 AND2X2_886 ( .A(u0__abc_76628_new_n3182_), .B(u0__abc_76628_new_n2724__bF_buf4), .Y(u0__abc_76628_new_n3183_));
AND2X2 AND2X2_887 ( .A(u0__abc_76628_new_n3183_), .B(u0__abc_76628_new_n3181_), .Y(u0__abc_76628_new_n3184_));
AND2X2 AND2X2_888 ( .A(u0__abc_76628_new_n3185_), .B(u0__abc_76628_new_n2720__bF_buf4), .Y(u0__abc_76628_new_n3186_));
AND2X2 AND2X2_889 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3187_));
AND2X2 AND2X2_89 ( .A(u0__abc_76628_new_n1142_), .B(u0__abc_76628_new_n1153_), .Y(u0__abc_76628_new_n1154_));
AND2X2 AND2X2_890 ( .A(u0__abc_76628_new_n3188_), .B(u0__abc_76628_new_n2719__bF_buf4), .Y(u0__abc_76628_new_n3189_));
AND2X2 AND2X2_891 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3190_));
AND2X2 AND2X2_892 ( .A(u0__abc_76628_new_n3191_), .B(u0__abc_76628_new_n2718__bF_buf4), .Y(u0__abc_76628_new_n3192_));
AND2X2 AND2X2_893 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3193_));
AND2X2 AND2X2_894 ( .A(u0__abc_76628_new_n3194_), .B(u0__abc_76628_new_n2717__bF_buf4), .Y(u0__abc_76628_new_n3195_));
AND2X2 AND2X2_895 ( .A(u0_tms1_19_), .B(u0_cs1_bF_buf3), .Y(u0__abc_76628_new_n3196_));
AND2X2 AND2X2_896 ( .A(u0__abc_76628_new_n1169__bF_buf0), .B(u0__abc_76628_new_n3199_), .Y(u0__abc_76628_new_n3200_));
AND2X2 AND2X2_897 ( .A(u0__abc_76628_new_n3198_), .B(u0__abc_76628_new_n3200_), .Y(u0__abc_76628_new_n3201_));
AND2X2 AND2X2_898 ( .A(u0__abc_76628_new_n1170__bF_buf0), .B(tms_20_), .Y(u0__abc_76628_new_n3203_));
AND2X2 AND2X2_899 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3204_));
AND2X2 AND2X2_9 ( .A(_abc_85006_new_n263_), .B(_abc_85006_new_n264_), .Y(obct_cs_3_));
AND2X2 AND2X2_90 ( .A(u0__abc_76628_new_n1154_), .B(u0__abc_76628_new_n1152_), .Y(u0__abc_76628_new_n1155_));
AND2X2 AND2X2_900 ( .A(u0__abc_76628_new_n3206_), .B(u0__abc_76628_new_n2724__bF_buf3), .Y(u0__abc_76628_new_n3207_));
AND2X2 AND2X2_901 ( .A(u0__abc_76628_new_n3207_), .B(u0__abc_76628_new_n3205_), .Y(u0__abc_76628_new_n3208_));
AND2X2 AND2X2_902 ( .A(u0__abc_76628_new_n3209_), .B(u0__abc_76628_new_n2720__bF_buf3), .Y(u0__abc_76628_new_n3210_));
AND2X2 AND2X2_903 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3211_));
AND2X2 AND2X2_904 ( .A(u0__abc_76628_new_n3212_), .B(u0__abc_76628_new_n2719__bF_buf3), .Y(u0__abc_76628_new_n3213_));
AND2X2 AND2X2_905 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3214_));
AND2X2 AND2X2_906 ( .A(u0__abc_76628_new_n3215_), .B(u0__abc_76628_new_n2718__bF_buf3), .Y(u0__abc_76628_new_n3216_));
AND2X2 AND2X2_907 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3217_));
AND2X2 AND2X2_908 ( .A(u0__abc_76628_new_n3218_), .B(u0__abc_76628_new_n2717__bF_buf3), .Y(u0__abc_76628_new_n3219_));
AND2X2 AND2X2_909 ( .A(u0_tms1_20_), .B(u0_cs1_bF_buf2), .Y(u0__abc_76628_new_n3220_));
AND2X2 AND2X2_91 ( .A(u0__abc_76628_new_n1138_), .B(u0__abc_76628_new_n1155_), .Y(u0__abc_76628_new_n1156_));
AND2X2 AND2X2_910 ( .A(u0__abc_76628_new_n1169__bF_buf6), .B(u0__abc_76628_new_n3223_), .Y(u0__abc_76628_new_n3224_));
AND2X2 AND2X2_911 ( .A(u0__abc_76628_new_n3222_), .B(u0__abc_76628_new_n3224_), .Y(u0__abc_76628_new_n3225_));
AND2X2 AND2X2_912 ( .A(u0__abc_76628_new_n1170__bF_buf6), .B(tms_21_), .Y(u0__abc_76628_new_n3227_));
AND2X2 AND2X2_913 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3228_));
AND2X2 AND2X2_914 ( .A(u0__abc_76628_new_n3230_), .B(u0__abc_76628_new_n2724__bF_buf2), .Y(u0__abc_76628_new_n3231_));
AND2X2 AND2X2_915 ( .A(u0__abc_76628_new_n3231_), .B(u0__abc_76628_new_n3229_), .Y(u0__abc_76628_new_n3232_));
AND2X2 AND2X2_916 ( .A(u0__abc_76628_new_n3233_), .B(u0__abc_76628_new_n2720__bF_buf2), .Y(u0__abc_76628_new_n3234_));
AND2X2 AND2X2_917 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3235_));
AND2X2 AND2X2_918 ( .A(u0__abc_76628_new_n3236_), .B(u0__abc_76628_new_n2719__bF_buf2), .Y(u0__abc_76628_new_n3237_));
AND2X2 AND2X2_919 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3238_));
AND2X2 AND2X2_92 ( .A(u0__abc_76628_new_n1109_), .B(spec_req_cs_7_), .Y(u0__abc_76628_new_n1158_));
AND2X2 AND2X2_920 ( .A(u0__abc_76628_new_n3239_), .B(u0__abc_76628_new_n2718__bF_buf2), .Y(u0__abc_76628_new_n3240_));
AND2X2 AND2X2_921 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3241_));
AND2X2 AND2X2_922 ( .A(u0__abc_76628_new_n3242_), .B(u0__abc_76628_new_n2717__bF_buf2), .Y(u0__abc_76628_new_n3243_));
AND2X2 AND2X2_923 ( .A(u0_tms1_21_), .B(u0_cs1_bF_buf1), .Y(u0__abc_76628_new_n3244_));
AND2X2 AND2X2_924 ( .A(u0__abc_76628_new_n1169__bF_buf5), .B(u0__abc_76628_new_n3247_), .Y(u0__abc_76628_new_n3248_));
AND2X2 AND2X2_925 ( .A(u0__abc_76628_new_n3246_), .B(u0__abc_76628_new_n3248_), .Y(u0__abc_76628_new_n3249_));
AND2X2 AND2X2_926 ( .A(u0__abc_76628_new_n1170__bF_buf5), .B(tms_22_), .Y(u0__abc_76628_new_n3251_));
AND2X2 AND2X2_927 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3252_));
AND2X2 AND2X2_928 ( .A(u0__abc_76628_new_n3254_), .B(u0__abc_76628_new_n2724__bF_buf1), .Y(u0__abc_76628_new_n3255_));
AND2X2 AND2X2_929 ( .A(u0__abc_76628_new_n3255_), .B(u0__abc_76628_new_n3253_), .Y(u0__abc_76628_new_n3256_));
AND2X2 AND2X2_93 ( .A(u0__abc_76628_new_n1161_), .B(u0__abc_76628_new_n1160_), .Y(u0__abc_76628_new_n1162_));
AND2X2 AND2X2_930 ( .A(u0__abc_76628_new_n3257_), .B(u0__abc_76628_new_n2720__bF_buf1), .Y(u0__abc_76628_new_n3258_));
AND2X2 AND2X2_931 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3259_));
AND2X2 AND2X2_932 ( .A(u0__abc_76628_new_n3260_), .B(u0__abc_76628_new_n2719__bF_buf1), .Y(u0__abc_76628_new_n3261_));
AND2X2 AND2X2_933 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3262_));
AND2X2 AND2X2_934 ( .A(u0__abc_76628_new_n3263_), .B(u0__abc_76628_new_n2718__bF_buf1), .Y(u0__abc_76628_new_n3264_));
AND2X2 AND2X2_935 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3265_));
AND2X2 AND2X2_936 ( .A(u0__abc_76628_new_n3266_), .B(u0__abc_76628_new_n2717__bF_buf1), .Y(u0__abc_76628_new_n3267_));
AND2X2 AND2X2_937 ( .A(u0_tms1_22_), .B(u0_cs1_bF_buf0), .Y(u0__abc_76628_new_n3268_));
AND2X2 AND2X2_938 ( .A(u0__abc_76628_new_n1169__bF_buf4), .B(u0__abc_76628_new_n3271_), .Y(u0__abc_76628_new_n3272_));
AND2X2 AND2X2_939 ( .A(u0__abc_76628_new_n3270_), .B(u0__abc_76628_new_n3272_), .Y(u0__abc_76628_new_n3273_));
AND2X2 AND2X2_94 ( .A(u0__abc_76628_new_n1159_), .B(u0__abc_76628_new_n1162_), .Y(u0__abc_76628_new_n1163_));
AND2X2 AND2X2_940 ( .A(u0__abc_76628_new_n1170__bF_buf4), .B(tms_23_), .Y(u0__abc_76628_new_n3275_));
AND2X2 AND2X2_941 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3276_));
AND2X2 AND2X2_942 ( .A(u0__abc_76628_new_n3278_), .B(u0__abc_76628_new_n2724__bF_buf0), .Y(u0__abc_76628_new_n3279_));
AND2X2 AND2X2_943 ( .A(u0__abc_76628_new_n3279_), .B(u0__abc_76628_new_n3277_), .Y(u0__abc_76628_new_n3280_));
AND2X2 AND2X2_944 ( .A(u0__abc_76628_new_n3281_), .B(u0__abc_76628_new_n2720__bF_buf0), .Y(u0__abc_76628_new_n3282_));
AND2X2 AND2X2_945 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3283_));
AND2X2 AND2X2_946 ( .A(u0__abc_76628_new_n3284_), .B(u0__abc_76628_new_n2719__bF_buf0), .Y(u0__abc_76628_new_n3285_));
AND2X2 AND2X2_947 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3286_));
AND2X2 AND2X2_948 ( .A(u0__abc_76628_new_n3287_), .B(u0__abc_76628_new_n2718__bF_buf0), .Y(u0__abc_76628_new_n3288_));
AND2X2 AND2X2_949 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3289_));
AND2X2 AND2X2_95 ( .A(u0__abc_76628_new_n1154_), .B(u0__abc_76628_new_n1163_), .Y(u0__abc_76628_new_n1164_));
AND2X2 AND2X2_950 ( .A(u0__abc_76628_new_n3290_), .B(u0__abc_76628_new_n2717__bF_buf0), .Y(u0__abc_76628_new_n3291_));
AND2X2 AND2X2_951 ( .A(u0_tms1_23_), .B(u0_cs1_bF_buf5), .Y(u0__abc_76628_new_n3292_));
AND2X2 AND2X2_952 ( .A(u0__abc_76628_new_n1169__bF_buf3), .B(u0__abc_76628_new_n3295_), .Y(u0__abc_76628_new_n3296_));
AND2X2 AND2X2_953 ( .A(u0__abc_76628_new_n3294_), .B(u0__abc_76628_new_n3296_), .Y(u0__abc_76628_new_n3297_));
AND2X2 AND2X2_954 ( .A(u0__abc_76628_new_n1170__bF_buf3), .B(tms_24_), .Y(u0__abc_76628_new_n3299_));
AND2X2 AND2X2_955 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3300_));
AND2X2 AND2X2_956 ( .A(u0__abc_76628_new_n3302_), .B(u0__abc_76628_new_n2724__bF_buf5), .Y(u0__abc_76628_new_n3303_));
AND2X2 AND2X2_957 ( .A(u0__abc_76628_new_n3303_), .B(u0__abc_76628_new_n3301_), .Y(u0__abc_76628_new_n3304_));
AND2X2 AND2X2_958 ( .A(u0__abc_76628_new_n3305_), .B(u0__abc_76628_new_n2720__bF_buf5), .Y(u0__abc_76628_new_n3306_));
AND2X2 AND2X2_959 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3307_));
AND2X2 AND2X2_96 ( .A(u0__abc_76628_new_n1138_), .B(u0__abc_76628_new_n1164_), .Y(u0__abc_76628_new_n1165_));
AND2X2 AND2X2_960 ( .A(u0__abc_76628_new_n3308_), .B(u0__abc_76628_new_n2719__bF_buf5), .Y(u0__abc_76628_new_n3309_));
AND2X2 AND2X2_961 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3310_));
AND2X2 AND2X2_962 ( .A(u0__abc_76628_new_n3311_), .B(u0__abc_76628_new_n2718__bF_buf5), .Y(u0__abc_76628_new_n3312_));
AND2X2 AND2X2_963 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3313_));
AND2X2 AND2X2_964 ( .A(u0__abc_76628_new_n3314_), .B(u0__abc_76628_new_n2717__bF_buf5), .Y(u0__abc_76628_new_n3315_));
AND2X2 AND2X2_965 ( .A(u0_tms1_24_), .B(u0_cs1_bF_buf4), .Y(u0__abc_76628_new_n3316_));
AND2X2 AND2X2_966 ( .A(u0__abc_76628_new_n1169__bF_buf2), .B(u0__abc_76628_new_n3319_), .Y(u0__abc_76628_new_n3320_));
AND2X2 AND2X2_967 ( .A(u0__abc_76628_new_n3318_), .B(u0__abc_76628_new_n3320_), .Y(u0__abc_76628_new_n3321_));
AND2X2 AND2X2_968 ( .A(u0__abc_76628_new_n1170__bF_buf2), .B(tms_25_), .Y(u0__abc_76628_new_n3323_));
AND2X2 AND2X2_969 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3324_));
AND2X2 AND2X2_97 ( .A(wb_stb_i_bF_buf4), .B(wb_cyc_i), .Y(u0__abc_76628_new_n1168_));
AND2X2 AND2X2_970 ( .A(u0__abc_76628_new_n3326_), .B(u0__abc_76628_new_n2724__bF_buf4), .Y(u0__abc_76628_new_n3327_));
AND2X2 AND2X2_971 ( .A(u0__abc_76628_new_n3327_), .B(u0__abc_76628_new_n3325_), .Y(u0__abc_76628_new_n3328_));
AND2X2 AND2X2_972 ( .A(u0__abc_76628_new_n3329_), .B(u0__abc_76628_new_n2720__bF_buf4), .Y(u0__abc_76628_new_n3330_));
AND2X2 AND2X2_973 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3331_));
AND2X2 AND2X2_974 ( .A(u0__abc_76628_new_n3332_), .B(u0__abc_76628_new_n2719__bF_buf4), .Y(u0__abc_76628_new_n3333_));
AND2X2 AND2X2_975 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3334_));
AND2X2 AND2X2_976 ( .A(u0__abc_76628_new_n3335_), .B(u0__abc_76628_new_n2718__bF_buf4), .Y(u0__abc_76628_new_n3336_));
AND2X2 AND2X2_977 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3337_));
AND2X2 AND2X2_978 ( .A(u0__abc_76628_new_n3338_), .B(u0__abc_76628_new_n2717__bF_buf4), .Y(u0__abc_76628_new_n3339_));
AND2X2 AND2X2_979 ( .A(u0_tms1_25_), .B(u0_cs1_bF_buf3), .Y(u0__abc_76628_new_n3340_));
AND2X2 AND2X2_98 ( .A(u0__abc_76628_new_n1167_), .B(u0__abc_76628_new_n1168_), .Y(u0__abc_76628_new_n1169_));
AND2X2 AND2X2_980 ( .A(u0__abc_76628_new_n1169__bF_buf1), .B(u0__abc_76628_new_n3343_), .Y(u0__abc_76628_new_n3344_));
AND2X2 AND2X2_981 ( .A(u0__abc_76628_new_n3342_), .B(u0__abc_76628_new_n3344_), .Y(u0__abc_76628_new_n3345_));
AND2X2 AND2X2_982 ( .A(u0__abc_76628_new_n1170__bF_buf1), .B(tms_26_), .Y(u0__abc_76628_new_n3347_));
AND2X2 AND2X2_983 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3348_));
AND2X2 AND2X2_984 ( .A(u0__abc_76628_new_n3350_), .B(u0__abc_76628_new_n2724__bF_buf3), .Y(u0__abc_76628_new_n3351_));
AND2X2 AND2X2_985 ( .A(u0__abc_76628_new_n3351_), .B(u0__abc_76628_new_n3349_), .Y(u0__abc_76628_new_n3352_));
AND2X2 AND2X2_986 ( .A(u0__abc_76628_new_n3353_), .B(u0__abc_76628_new_n2720__bF_buf3), .Y(u0__abc_76628_new_n3354_));
AND2X2 AND2X2_987 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3355_));
AND2X2 AND2X2_988 ( .A(u0__abc_76628_new_n3356_), .B(u0__abc_76628_new_n2719__bF_buf3), .Y(u0__abc_76628_new_n3357_));
AND2X2 AND2X2_989 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3358_));
AND2X2 AND2X2_99 ( .A(u0__abc_76628_new_n1170__bF_buf6), .B(sp_tms_0_), .Y(u0__abc_76628_new_n1171_));
AND2X2 AND2X2_990 ( .A(u0__abc_76628_new_n3359_), .B(u0__abc_76628_new_n2718__bF_buf3), .Y(u0__abc_76628_new_n3360_));
AND2X2 AND2X2_991 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3361_));
AND2X2 AND2X2_992 ( .A(u0__abc_76628_new_n3362_), .B(u0__abc_76628_new_n2717__bF_buf3), .Y(u0__abc_76628_new_n3363_));
AND2X2 AND2X2_993 ( .A(u0_tms1_26_), .B(u0_cs1_bF_buf2), .Y(u0__abc_76628_new_n3364_));
AND2X2 AND2X2_994 ( .A(u0__abc_76628_new_n1169__bF_buf0), .B(u0__abc_76628_new_n3367_), .Y(u0__abc_76628_new_n3368_));
AND2X2 AND2X2_995 ( .A(u0__abc_76628_new_n3366_), .B(u0__abc_76628_new_n3368_), .Y(u0__abc_76628_new_n3369_));
AND2X2 AND2X2_996 ( .A(u0__abc_76628_new_n1170__bF_buf0), .B(tms_27_), .Y(u0__abc_76628_new_n3371_));
AND2X2 AND2X2_997 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3372_));
AND2X2 AND2X2_998 ( .A(u0__abc_76628_new_n3374_), .B(u0__abc_76628_new_n2724__bF_buf2), .Y(u0__abc_76628_new_n3375_));
AND2X2 AND2X2_999 ( .A(u0__abc_76628_new_n3375_), .B(u0__abc_76628_new_n3373_), .Y(u0__abc_76628_new_n3376_));
BUFX2 BUFX2_1 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf1_));
BUFX2 BUFX2_10 ( .A(u5__abc_81276_new_n479_), .Y(u5__abc_81276_new_n479__bF_buf1));
BUFX2 BUFX2_100 ( .A(_auto_iopadmap_cc_368_execute_85420_6_), .Y(\mc_addr_pad_o[6] ));
BUFX2 BUFX2_101 ( .A(_auto_iopadmap_cc_368_execute_85420_7_), .Y(\mc_addr_pad_o[7] ));
BUFX2 BUFX2_102 ( .A(_auto_iopadmap_cc_368_execute_85420_8_), .Y(\mc_addr_pad_o[8] ));
BUFX2 BUFX2_103 ( .A(_auto_iopadmap_cc_368_execute_85420_9_), .Y(\mc_addr_pad_o[9] ));
BUFX2 BUFX2_104 ( .A(_auto_iopadmap_cc_368_execute_85420_10_), .Y(\mc_addr_pad_o[10] ));
BUFX2 BUFX2_105 ( .A(_auto_iopadmap_cc_368_execute_85420_11_), .Y(\mc_addr_pad_o[11] ));
BUFX2 BUFX2_106 ( .A(_auto_iopadmap_cc_368_execute_85420_12_), .Y(\mc_addr_pad_o[12] ));
BUFX2 BUFX2_107 ( .A(_auto_iopadmap_cc_368_execute_85420_13_), .Y(\mc_addr_pad_o[13] ));
BUFX2 BUFX2_108 ( .A(_auto_iopadmap_cc_368_execute_85420_14_), .Y(\mc_addr_pad_o[14] ));
BUFX2 BUFX2_109 ( .A(_auto_iopadmap_cc_368_execute_85420_15_), .Y(\mc_addr_pad_o[15] ));
BUFX2 BUFX2_11 ( .A(u5__abc_81276_new_n479_), .Y(u5__abc_81276_new_n479__bF_buf0));
BUFX2 BUFX2_110 ( .A(_auto_iopadmap_cc_368_execute_85420_16_), .Y(\mc_addr_pad_o[16] ));
BUFX2 BUFX2_111 ( .A(_auto_iopadmap_cc_368_execute_85420_17_), .Y(\mc_addr_pad_o[17] ));
BUFX2 BUFX2_112 ( .A(_auto_iopadmap_cc_368_execute_85420_18_), .Y(\mc_addr_pad_o[18] ));
BUFX2 BUFX2_113 ( .A(_auto_iopadmap_cc_368_execute_85420_19_), .Y(\mc_addr_pad_o[19] ));
BUFX2 BUFX2_114 ( .A(_auto_iopadmap_cc_368_execute_85420_20_), .Y(\mc_addr_pad_o[20] ));
BUFX2 BUFX2_115 ( .A(_auto_iopadmap_cc_368_execute_85420_21_), .Y(\mc_addr_pad_o[21] ));
BUFX2 BUFX2_116 ( .A(_auto_iopadmap_cc_368_execute_85420_22_), .Y(\mc_addr_pad_o[22] ));
BUFX2 BUFX2_117 ( .A(_auto_iopadmap_cc_368_execute_85420_23_), .Y(\mc_addr_pad_o[23] ));
BUFX2 BUFX2_118 ( .A(_auto_iopadmap_cc_368_execute_85445), .Y(mc_adsc_pad_o_));
BUFX2 BUFX2_119 ( .A(_auto_iopadmap_cc_368_execute_85447), .Y(mc_adv_pad_o_));
BUFX2 BUFX2_12 ( .A(u0__abc_76628_new_n4541_), .Y(u0__abc_76628_new_n4541__bF_buf3));
BUFX2 BUFX2_120 ( .A(_auto_iopadmap_cc_368_execute_85449), .Y(mc_bg_pad_o));
BUFX2 BUFX2_121 ( .A(_auto_iopadmap_cc_368_execute_85451), .Y(mc_cas_pad_o_));
BUFX2 BUFX2_122 ( .A(_auto_iopadmap_cc_368_execute_85453), .Y(mc_cke_pad_o_));
BUFX2 BUFX2_123 ( .A(_auto_iopadmap_cc_368_execute_85455), .Y(mc_coe_pad_coe_o));
BUFX2 BUFX2_124 ( .A(_auto_iopadmap_cc_368_execute_85457_0_), .Y(\mc_cs_pad_o_[0] ));
BUFX2 BUFX2_125 ( .A(_auto_iopadmap_cc_368_execute_85457_1_), .Y(\mc_cs_pad_o_[1] ));
BUFX2 BUFX2_126 ( .A(_auto_iopadmap_cc_368_execute_85457_2_), .Y(\mc_cs_pad_o_[2] ));
BUFX2 BUFX2_127 ( .A(_auto_iopadmap_cc_368_execute_85457_3_), .Y(\mc_cs_pad_o_[3] ));
BUFX2 BUFX2_128 ( .A(_auto_iopadmap_cc_368_execute_85457_4_), .Y(\mc_cs_pad_o_[4] ));
BUFX2 BUFX2_129 ( .A(_auto_iopadmap_cc_368_execute_85457_5_), .Y(\mc_cs_pad_o_[5] ));
BUFX2 BUFX2_13 ( .A(u0__abc_76628_new_n4541_), .Y(u0__abc_76628_new_n4541__bF_buf2));
BUFX2 BUFX2_130 ( .A(_auto_iopadmap_cc_368_execute_85457_6_), .Y(\mc_cs_pad_o_[6] ));
BUFX2 BUFX2_131 ( .A(_auto_iopadmap_cc_368_execute_85457_7_), .Y(\mc_cs_pad_o_[7] ));
BUFX2 BUFX2_132 ( .A(_auto_iopadmap_cc_368_execute_85466_0_), .Y(\mc_data_pad_o[0] ));
BUFX2 BUFX2_133 ( .A(_auto_iopadmap_cc_368_execute_85466_1_), .Y(\mc_data_pad_o[1] ));
BUFX2 BUFX2_134 ( .A(_auto_iopadmap_cc_368_execute_85466_2_), .Y(\mc_data_pad_o[2] ));
BUFX2 BUFX2_135 ( .A(_auto_iopadmap_cc_368_execute_85466_3_), .Y(\mc_data_pad_o[3] ));
BUFX2 BUFX2_136 ( .A(_auto_iopadmap_cc_368_execute_85466_4_), .Y(\mc_data_pad_o[4] ));
BUFX2 BUFX2_137 ( .A(_auto_iopadmap_cc_368_execute_85466_5_), .Y(\mc_data_pad_o[5] ));
BUFX2 BUFX2_138 ( .A(_auto_iopadmap_cc_368_execute_85466_6_), .Y(\mc_data_pad_o[6] ));
BUFX2 BUFX2_139 ( .A(_auto_iopadmap_cc_368_execute_85466_7_), .Y(\mc_data_pad_o[7] ));
BUFX2 BUFX2_14 ( .A(u0__abc_76628_new_n4541_), .Y(u0__abc_76628_new_n4541__bF_buf1));
BUFX2 BUFX2_140 ( .A(_auto_iopadmap_cc_368_execute_85466_8_), .Y(\mc_data_pad_o[8] ));
BUFX2 BUFX2_141 ( .A(_auto_iopadmap_cc_368_execute_85466_9_), .Y(\mc_data_pad_o[9] ));
BUFX2 BUFX2_142 ( .A(_auto_iopadmap_cc_368_execute_85466_10_), .Y(\mc_data_pad_o[10] ));
BUFX2 BUFX2_143 ( .A(_auto_iopadmap_cc_368_execute_85466_11_), .Y(\mc_data_pad_o[11] ));
BUFX2 BUFX2_144 ( .A(_auto_iopadmap_cc_368_execute_85466_12_), .Y(\mc_data_pad_o[12] ));
BUFX2 BUFX2_145 ( .A(_auto_iopadmap_cc_368_execute_85466_13_), .Y(\mc_data_pad_o[13] ));
BUFX2 BUFX2_146 ( .A(_auto_iopadmap_cc_368_execute_85466_14_), .Y(\mc_data_pad_o[14] ));
BUFX2 BUFX2_147 ( .A(_auto_iopadmap_cc_368_execute_85466_15_), .Y(\mc_data_pad_o[15] ));
BUFX2 BUFX2_148 ( .A(_auto_iopadmap_cc_368_execute_85466_16_), .Y(\mc_data_pad_o[16] ));
BUFX2 BUFX2_149 ( .A(_auto_iopadmap_cc_368_execute_85466_17_), .Y(\mc_data_pad_o[17] ));
BUFX2 BUFX2_15 ( .A(u0__abc_76628_new_n4541_), .Y(u0__abc_76628_new_n4541__bF_buf0));
BUFX2 BUFX2_150 ( .A(_auto_iopadmap_cc_368_execute_85466_18_), .Y(\mc_data_pad_o[18] ));
BUFX2 BUFX2_151 ( .A(_auto_iopadmap_cc_368_execute_85466_19_), .Y(\mc_data_pad_o[19] ));
BUFX2 BUFX2_152 ( .A(_auto_iopadmap_cc_368_execute_85466_20_), .Y(\mc_data_pad_o[20] ));
BUFX2 BUFX2_153 ( .A(_auto_iopadmap_cc_368_execute_85466_21_), .Y(\mc_data_pad_o[21] ));
BUFX2 BUFX2_154 ( .A(_auto_iopadmap_cc_368_execute_85466_22_), .Y(\mc_data_pad_o[22] ));
BUFX2 BUFX2_155 ( .A(_auto_iopadmap_cc_368_execute_85466_23_), .Y(\mc_data_pad_o[23] ));
BUFX2 BUFX2_156 ( .A(_auto_iopadmap_cc_368_execute_85466_24_), .Y(\mc_data_pad_o[24] ));
BUFX2 BUFX2_157 ( .A(_auto_iopadmap_cc_368_execute_85466_25_), .Y(\mc_data_pad_o[25] ));
BUFX2 BUFX2_158 ( .A(_auto_iopadmap_cc_368_execute_85466_26_), .Y(\mc_data_pad_o[26] ));
BUFX2 BUFX2_159 ( .A(_auto_iopadmap_cc_368_execute_85466_27_), .Y(\mc_data_pad_o[27] ));
BUFX2 BUFX2_16 ( .A(u5__abc_81276_new_n2953_), .Y(u5__abc_81276_new_n2953__bF_buf3));
BUFX2 BUFX2_160 ( .A(_auto_iopadmap_cc_368_execute_85466_28_), .Y(\mc_data_pad_o[28] ));
BUFX2 BUFX2_161 ( .A(_auto_iopadmap_cc_368_execute_85466_29_), .Y(\mc_data_pad_o[29] ));
BUFX2 BUFX2_162 ( .A(_auto_iopadmap_cc_368_execute_85466_30_), .Y(\mc_data_pad_o[30] ));
BUFX2 BUFX2_163 ( .A(_auto_iopadmap_cc_368_execute_85466_31_), .Y(\mc_data_pad_o[31] ));
BUFX2 BUFX2_164 ( .A(_auto_iopadmap_cc_368_execute_85499), .Y(mc_doe_pad_doe_o));
BUFX2 BUFX2_165 ( .A(_auto_iopadmap_cc_368_execute_85501_0_), .Y(\mc_dp_pad_o[0] ));
BUFX2 BUFX2_166 ( .A(_auto_iopadmap_cc_368_execute_85501_1_), .Y(\mc_dp_pad_o[1] ));
BUFX2 BUFX2_167 ( .A(_auto_iopadmap_cc_368_execute_85501_2_), .Y(\mc_dp_pad_o[2] ));
BUFX2 BUFX2_168 ( .A(_auto_iopadmap_cc_368_execute_85501_3_), .Y(\mc_dp_pad_o[3] ));
BUFX2 BUFX2_169 ( .A(_auto_iopadmap_cc_368_execute_85506_0_), .Y(\mc_dqm_pad_o[0] ));
BUFX2 BUFX2_17 ( .A(u5__abc_81276_new_n2953_), .Y(u5__abc_81276_new_n2953__bF_buf2));
BUFX2 BUFX2_170 ( .A(_auto_iopadmap_cc_368_execute_85506_1_), .Y(\mc_dqm_pad_o[1] ));
BUFX2 BUFX2_171 ( .A(_auto_iopadmap_cc_368_execute_85506_2_), .Y(\mc_dqm_pad_o[2] ));
BUFX2 BUFX2_172 ( .A(_auto_iopadmap_cc_368_execute_85506_3_), .Y(\mc_dqm_pad_o[3] ));
BUFX2 BUFX2_173 ( .A(_auto_iopadmap_cc_368_execute_85511), .Y(mc_oe_pad_o_));
BUFX2 BUFX2_174 ( .A(_auto_iopadmap_cc_368_execute_85513), .Y(mc_ras_pad_o_));
BUFX2 BUFX2_175 ( .A(_auto_iopadmap_cc_368_execute_85515), .Y(mc_rp_pad_o_));
BUFX2 BUFX2_176 ( .A(u0_csr_1_), .Y(mc_vpen_pad_o));
BUFX2 BUFX2_177 ( .A(_auto_iopadmap_cc_368_execute_85519), .Y(mc_we_pad_o_));
BUFX2 BUFX2_178 ( .A(_auto_iopadmap_cc_368_execute_85521), .Y(mc_zz_pad_o));
BUFX2 BUFX2_179 ( .A(_auto_iopadmap_cc_368_execute_85523_0_), .Y(\poc_o[0] ));
BUFX2 BUFX2_18 ( .A(u5__abc_81276_new_n2953_), .Y(u5__abc_81276_new_n2953__bF_buf1));
BUFX2 BUFX2_180 ( .A(_auto_iopadmap_cc_368_execute_85523_1_), .Y(\poc_o[1] ));
BUFX2 BUFX2_181 ( .A(_auto_iopadmap_cc_368_execute_85523_2_), .Y(\poc_o[2] ));
BUFX2 BUFX2_182 ( .A(_auto_iopadmap_cc_368_execute_85523_3_), .Y(\poc_o[3] ));
BUFX2 BUFX2_183 ( .A(_auto_iopadmap_cc_368_execute_85523_4_), .Y(\poc_o[4] ));
BUFX2 BUFX2_184 ( .A(_auto_iopadmap_cc_368_execute_85523_5_), .Y(\poc_o[5] ));
BUFX2 BUFX2_185 ( .A(_auto_iopadmap_cc_368_execute_85523_6_), .Y(\poc_o[6] ));
BUFX2 BUFX2_186 ( .A(_auto_iopadmap_cc_368_execute_85523_7_), .Y(\poc_o[7] ));
BUFX2 BUFX2_187 ( .A(_auto_iopadmap_cc_368_execute_85523_8_), .Y(\poc_o[8] ));
BUFX2 BUFX2_188 ( .A(_auto_iopadmap_cc_368_execute_85523_9_), .Y(\poc_o[9] ));
BUFX2 BUFX2_189 ( .A(_auto_iopadmap_cc_368_execute_85523_10_), .Y(\poc_o[10] ));
BUFX2 BUFX2_19 ( .A(u5__abc_81276_new_n2953_), .Y(u5__abc_81276_new_n2953__bF_buf0));
BUFX2 BUFX2_190 ( .A(_auto_iopadmap_cc_368_execute_85523_11_), .Y(\poc_o[11] ));
BUFX2 BUFX2_191 ( .A(_auto_iopadmap_cc_368_execute_85523_12_), .Y(\poc_o[12] ));
BUFX2 BUFX2_192 ( .A(_auto_iopadmap_cc_368_execute_85523_13_), .Y(\poc_o[13] ));
BUFX2 BUFX2_193 ( .A(_auto_iopadmap_cc_368_execute_85523_14_), .Y(\poc_o[14] ));
BUFX2 BUFX2_194 ( .A(_auto_iopadmap_cc_368_execute_85523_15_), .Y(\poc_o[15] ));
BUFX2 BUFX2_195 ( .A(_auto_iopadmap_cc_368_execute_85523_16_), .Y(\poc_o[16] ));
BUFX2 BUFX2_196 ( .A(_auto_iopadmap_cc_368_execute_85523_17_), .Y(\poc_o[17] ));
BUFX2 BUFX2_197 ( .A(_auto_iopadmap_cc_368_execute_85523_18_), .Y(\poc_o[18] ));
BUFX2 BUFX2_198 ( .A(_auto_iopadmap_cc_368_execute_85523_19_), .Y(\poc_o[19] ));
BUFX2 BUFX2_199 ( .A(_auto_iopadmap_cc_368_execute_85523_20_), .Y(\poc_o[20] ));
BUFX2 BUFX2_2 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf0_));
BUFX2 BUFX2_20 ( .A(u0__abc_76628_new_n4438_), .Y(u0__abc_76628_new_n4438__bF_buf1));
BUFX2 BUFX2_200 ( .A(_auto_iopadmap_cc_368_execute_85523_21_), .Y(\poc_o[21] ));
BUFX2 BUFX2_201 ( .A(_auto_iopadmap_cc_368_execute_85523_22_), .Y(\poc_o[22] ));
BUFX2 BUFX2_202 ( .A(_auto_iopadmap_cc_368_execute_85523_23_), .Y(\poc_o[23] ));
BUFX2 BUFX2_203 ( .A(_auto_iopadmap_cc_368_execute_85523_24_), .Y(\poc_o[24] ));
BUFX2 BUFX2_204 ( .A(_auto_iopadmap_cc_368_execute_85523_25_), .Y(\poc_o[25] ));
BUFX2 BUFX2_205 ( .A(_auto_iopadmap_cc_368_execute_85523_26_), .Y(\poc_o[26] ));
BUFX2 BUFX2_206 ( .A(_auto_iopadmap_cc_368_execute_85523_27_), .Y(\poc_o[27] ));
BUFX2 BUFX2_207 ( .A(_auto_iopadmap_cc_368_execute_85523_28_), .Y(\poc_o[28] ));
BUFX2 BUFX2_208 ( .A(_auto_iopadmap_cc_368_execute_85523_29_), .Y(\poc_o[29] ));
BUFX2 BUFX2_209 ( .A(_auto_iopadmap_cc_368_execute_85523_30_), .Y(\poc_o[30] ));
BUFX2 BUFX2_21 ( .A(u0__abc_76628_new_n4438_), .Y(u0__abc_76628_new_n4438__bF_buf0));
BUFX2 BUFX2_210 ( .A(_auto_iopadmap_cc_368_execute_85523_31_), .Y(\poc_o[31] ));
BUFX2 BUFX2_211 ( .A(_auto_iopadmap_cc_368_execute_85556), .Y(suspended_o));
BUFX2 BUFX2_212 ( .A(_auto_iopadmap_cc_368_execute_85558), .Y(wb_ack_o));
BUFX2 BUFX2_213 ( .A(_auto_iopadmap_cc_368_execute_85560_0_), .Y(\wb_data_o[0] ));
BUFX2 BUFX2_214 ( .A(_auto_iopadmap_cc_368_execute_85560_1_), .Y(\wb_data_o[1] ));
BUFX2 BUFX2_215 ( .A(_auto_iopadmap_cc_368_execute_85560_2_), .Y(\wb_data_o[2] ));
BUFX2 BUFX2_216 ( .A(_auto_iopadmap_cc_368_execute_85560_3_), .Y(\wb_data_o[3] ));
BUFX2 BUFX2_217 ( .A(_auto_iopadmap_cc_368_execute_85560_4_), .Y(\wb_data_o[4] ));
BUFX2 BUFX2_218 ( .A(_auto_iopadmap_cc_368_execute_85560_5_), .Y(\wb_data_o[5] ));
BUFX2 BUFX2_219 ( .A(_auto_iopadmap_cc_368_execute_85560_6_), .Y(\wb_data_o[6] ));
BUFX2 BUFX2_22 ( .A(u1__abc_73140_new_n275_), .Y(u1__abc_73140_new_n275__bF_buf1));
BUFX2 BUFX2_220 ( .A(_auto_iopadmap_cc_368_execute_85560_7_), .Y(\wb_data_o[7] ));
BUFX2 BUFX2_221 ( .A(_auto_iopadmap_cc_368_execute_85560_8_), .Y(\wb_data_o[8] ));
BUFX2 BUFX2_222 ( .A(_auto_iopadmap_cc_368_execute_85560_9_), .Y(\wb_data_o[9] ));
BUFX2 BUFX2_223 ( .A(_auto_iopadmap_cc_368_execute_85560_10_), .Y(\wb_data_o[10] ));
BUFX2 BUFX2_224 ( .A(_auto_iopadmap_cc_368_execute_85560_11_), .Y(\wb_data_o[11] ));
BUFX2 BUFX2_225 ( .A(_auto_iopadmap_cc_368_execute_85560_12_), .Y(\wb_data_o[12] ));
BUFX2 BUFX2_226 ( .A(_auto_iopadmap_cc_368_execute_85560_13_), .Y(\wb_data_o[13] ));
BUFX2 BUFX2_227 ( .A(_auto_iopadmap_cc_368_execute_85560_14_), .Y(\wb_data_o[14] ));
BUFX2 BUFX2_228 ( .A(_auto_iopadmap_cc_368_execute_85560_15_), .Y(\wb_data_o[15] ));
BUFX2 BUFX2_229 ( .A(_auto_iopadmap_cc_368_execute_85560_16_), .Y(\wb_data_o[16] ));
BUFX2 BUFX2_23 ( .A(u1__abc_73140_new_n275_), .Y(u1__abc_73140_new_n275__bF_buf0));
BUFX2 BUFX2_230 ( .A(_auto_iopadmap_cc_368_execute_85560_17_), .Y(\wb_data_o[17] ));
BUFX2 BUFX2_231 ( .A(_auto_iopadmap_cc_368_execute_85560_18_), .Y(\wb_data_o[18] ));
BUFX2 BUFX2_232 ( .A(_auto_iopadmap_cc_368_execute_85560_19_), .Y(\wb_data_o[19] ));
BUFX2 BUFX2_233 ( .A(_auto_iopadmap_cc_368_execute_85560_20_), .Y(\wb_data_o[20] ));
BUFX2 BUFX2_234 ( .A(_auto_iopadmap_cc_368_execute_85560_21_), .Y(\wb_data_o[21] ));
BUFX2 BUFX2_235 ( .A(_auto_iopadmap_cc_368_execute_85560_22_), .Y(\wb_data_o[22] ));
BUFX2 BUFX2_236 ( .A(_auto_iopadmap_cc_368_execute_85560_23_), .Y(\wb_data_o[23] ));
BUFX2 BUFX2_237 ( .A(_auto_iopadmap_cc_368_execute_85560_24_), .Y(\wb_data_o[24] ));
BUFX2 BUFX2_238 ( .A(_auto_iopadmap_cc_368_execute_85560_25_), .Y(\wb_data_o[25] ));
BUFX2 BUFX2_239 ( .A(_auto_iopadmap_cc_368_execute_85560_26_), .Y(\wb_data_o[26] ));
BUFX2 BUFX2_24 ( .A(u5__abc_81276_new_n3215_), .Y(u5__abc_81276_new_n3215__bF_buf2));
BUFX2 BUFX2_240 ( .A(_auto_iopadmap_cc_368_execute_85560_27_), .Y(\wb_data_o[27] ));
BUFX2 BUFX2_241 ( .A(_auto_iopadmap_cc_368_execute_85560_28_), .Y(\wb_data_o[28] ));
BUFX2 BUFX2_242 ( .A(_auto_iopadmap_cc_368_execute_85560_29_), .Y(\wb_data_o[29] ));
BUFX2 BUFX2_243 ( .A(_auto_iopadmap_cc_368_execute_85560_30_), .Y(\wb_data_o[30] ));
BUFX2 BUFX2_244 ( .A(_auto_iopadmap_cc_368_execute_85560_31_), .Y(\wb_data_o[31] ));
BUFX2 BUFX2_245 ( .A(_auto_iopadmap_cc_368_execute_85593), .Y(wb_err_o));
BUFX2 BUFX2_25 ( .A(u5__abc_81276_new_n3215_), .Y(u5__abc_81276_new_n3215__bF_buf1));
BUFX2 BUFX2_26 ( .A(u5__abc_81276_new_n3215_), .Y(u5__abc_81276_new_n3215__bF_buf0));
BUFX2 BUFX2_27 ( .A(u5__abc_81276_new_n464_), .Y(u5__abc_81276_new_n464__bF_buf0));
BUFX2 BUFX2_28 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf1_));
BUFX2 BUFX2_29 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf0_));
BUFX2 BUFX2_3 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf1_));
BUFX2 BUFX2_30 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf1_));
BUFX2 BUFX2_31 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf0_));
BUFX2 BUFX2_32 ( .A(u3__abc_74070_new_n450_), .Y(u3__abc_74070_new_n450__bF_buf3));
BUFX2 BUFX2_33 ( .A(u3__abc_74070_new_n450_), .Y(u3__abc_74070_new_n450__bF_buf2));
BUFX2 BUFX2_34 ( .A(u3__abc_74070_new_n450_), .Y(u3__abc_74070_new_n450__bF_buf1));
BUFX2 BUFX2_35 ( .A(u3__abc_74070_new_n450_), .Y(u3__abc_74070_new_n450__bF_buf0));
BUFX2 BUFX2_36 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf1_));
BUFX2 BUFX2_37 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf0_));
BUFX2 BUFX2_38 ( .A(u5__abc_81276_new_n417_), .Y(u5__abc_81276_new_n417__bF_buf0));
BUFX2 BUFX2_39 ( .A(u2_u1__abc_74955_new_n137_), .Y(u2_u1__abc_74955_new_n137__bF_buf1));
BUFX2 BUFX2_4 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf0_));
BUFX2 BUFX2_40 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf1_));
BUFX2 BUFX2_41 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf0_));
BUFX2 BUFX2_42 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf3_));
BUFX2 BUFX2_43 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf1_));
BUFX2 BUFX2_44 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf0_));
BUFX2 BUFX2_45 ( .A(cs_le), .Y(cs_le_bF_buf0));
BUFX2 BUFX2_46 ( .A(u5__abc_81276_new_n3323_), .Y(u5__abc_81276_new_n3323__bF_buf3));
BUFX2 BUFX2_47 ( .A(u5__abc_81276_new_n3323_), .Y(u5__abc_81276_new_n3323__bF_buf2));
BUFX2 BUFX2_48 ( .A(u5__abc_81276_new_n3323_), .Y(u5__abc_81276_new_n3323__bF_buf1));
BUFX2 BUFX2_49 ( .A(u5__abc_81276_new_n3323_), .Y(u5__abc_81276_new_n3323__bF_buf0));
BUFX2 BUFX2_5 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf1_));
BUFX2 BUFX2_50 ( .A(u5_tmr_done), .Y(u5_tmr_done_bF_buf3));
BUFX2 BUFX2_51 ( .A(u5_tmr_done), .Y(u5_tmr_done_bF_buf2));
BUFX2 BUFX2_52 ( .A(u5_tmr_done), .Y(u5_tmr_done_bF_buf0));
BUFX2 BUFX2_53 ( .A(u0__abc_76628_new_n1947_), .Y(u0__abc_76628_new_n1947__bF_buf3));
BUFX2 BUFX2_54 ( .A(u0__abc_76628_new_n1947_), .Y(u0__abc_76628_new_n1947__bF_buf2));
BUFX2 BUFX2_55 ( .A(u0__abc_76628_new_n1947_), .Y(u0__abc_76628_new_n1947__bF_buf1));
BUFX2 BUFX2_56 ( .A(u0__abc_76628_new_n1947_), .Y(u0__abc_76628_new_n1947__bF_buf0));
BUFX2 BUFX2_57 ( .A(u0__abc_76628_new_n4437_), .Y(u0__abc_76628_new_n4437__bF_buf0));
BUFX2 BUFX2_58 ( .A(u3__abc_74070_new_n452_), .Y(u3__abc_74070_new_n452__bF_buf3));
BUFX2 BUFX2_59 ( .A(u3__abc_74070_new_n452_), .Y(u3__abc_74070_new_n452__bF_buf2));
BUFX2 BUFX2_6 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf0_));
BUFX2 BUFX2_60 ( .A(u3__abc_74070_new_n452_), .Y(u3__abc_74070_new_n452__bF_buf1));
BUFX2 BUFX2_61 ( .A(u3__abc_74070_new_n452_), .Y(u3__abc_74070_new_n452__bF_buf0));
BUFX2 BUFX2_62 ( .A(u5_cmd_asserted), .Y(u5_cmd_asserted_bF_buf2));
BUFX2 BUFX2_63 ( .A(u3__abc_74070_new_n449_), .Y(u3__abc_74070_new_n449__bF_buf1));
BUFX2 BUFX2_64 ( .A(u3__abc_74070_new_n449_), .Y(u3__abc_74070_new_n449__bF_buf0));
BUFX2 BUFX2_65 ( .A(u1__abc_73140_new_n268_), .Y(u1__abc_73140_new_n268__bF_buf3));
BUFX2 BUFX2_66 ( .A(u1__abc_73140_new_n268_), .Y(u1__abc_73140_new_n268__bF_buf2));
BUFX2 BUFX2_67 ( .A(u1__abc_73140_new_n268_), .Y(u1__abc_73140_new_n268__bF_buf1));
BUFX2 BUFX2_68 ( .A(u1__abc_73140_new_n268_), .Y(u1__abc_73140_new_n268__bF_buf0));
BUFX2 BUFX2_69 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf1_));
BUFX2 BUFX2_7 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf1_));
BUFX2 BUFX2_70 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf0_));
BUFX2 BUFX2_71 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf1_));
BUFX2 BUFX2_72 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf0_));
BUFX2 BUFX2_73 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf1_));
BUFX2 BUFX2_74 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf0_));
BUFX2 BUFX2_75 ( .A(u5__abc_81276_new_n416_), .Y(u5__abc_81276_new_n416__bF_buf1));
BUFX2 BUFX2_76 ( .A(u5__abc_81276_new_n416_), .Y(u5__abc_81276_new_n416__bF_buf0));
BUFX2 BUFX2_77 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf1_));
BUFX2 BUFX2_78 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf0_));
BUFX2 BUFX2_79 ( .A(u5__abc_81276_new_n401_), .Y(u5__abc_81276_new_n401__bF_buf3));
BUFX2 BUFX2_8 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf0_));
BUFX2 BUFX2_80 ( .A(u5__abc_81276_new_n401_), .Y(u5__abc_81276_new_n401__bF_buf2));
BUFX2 BUFX2_81 ( .A(u5__abc_81276_new_n401_), .Y(u5__abc_81276_new_n401__bF_buf1));
BUFX2 BUFX2_82 ( .A(u5__abc_81276_new_n401_), .Y(u5__abc_81276_new_n401__bF_buf0));
BUFX2 BUFX2_83 ( .A(u0__abc_76628_new_n1946_), .Y(u0__abc_76628_new_n1946__bF_buf2));
BUFX2 BUFX2_84 ( .A(u0__abc_76628_new_n1946_), .Y(u0__abc_76628_new_n1946__bF_buf1));
BUFX2 BUFX2_85 ( .A(u0__abc_76628_new_n1946_), .Y(u0__abc_76628_new_n1946__bF_buf0));
BUFX2 BUFX2_86 ( .A(u1_bas), .Y(u1_bas_bF_buf1));
BUFX2 BUFX2_87 ( .A(u1_bas), .Y(u1_bas_bF_buf0));
BUFX2 BUFX2_88 ( .A(u5__abc_81276_new_n1126_), .Y(u5__abc_81276_new_n1126__bF_buf3));
BUFX2 BUFX2_89 ( .A(u5__abc_81276_new_n1126_), .Y(u5__abc_81276_new_n1126__bF_buf2));
BUFX2 BUFX2_9 ( .A(u2_u0__abc_74955_new_n137_), .Y(u2_u0__abc_74955_new_n137__bF_buf1));
BUFX2 BUFX2_90 ( .A(u5__abc_81276_new_n1126_), .Y(u5__abc_81276_new_n1126__bF_buf1));
BUFX2 BUFX2_91 ( .A(u5__abc_81276_new_n1126_), .Y(u5__abc_81276_new_n1126__bF_buf0));
BUFX2 BUFX2_92 ( .A(u5__abc_81276_new_n521_), .Y(u5__abc_81276_new_n521__bF_buf1));
BUFX2 BUFX2_93 ( .A(u5__abc_81276_new_n521_), .Y(u5__abc_81276_new_n521__bF_buf0));
BUFX2 BUFX2_94 ( .A(_auto_iopadmap_cc_368_execute_85420_0_), .Y(\mc_addr_pad_o[0] ));
BUFX2 BUFX2_95 ( .A(_auto_iopadmap_cc_368_execute_85420_1_), .Y(\mc_addr_pad_o[1] ));
BUFX2 BUFX2_96 ( .A(_auto_iopadmap_cc_368_execute_85420_2_), .Y(\mc_addr_pad_o[2] ));
BUFX2 BUFX2_97 ( .A(_auto_iopadmap_cc_368_execute_85420_3_), .Y(\mc_addr_pad_o[3] ));
BUFX2 BUFX2_98 ( .A(_auto_iopadmap_cc_368_execute_85420_4_), .Y(\mc_addr_pad_o[4] ));
BUFX2 BUFX2_99 ( .A(_auto_iopadmap_cc_368_execute_85420_5_), .Y(\mc_addr_pad_o[5] ));
BUFX4 BUFX4_1 ( .A(clk_i), .Y(clk_i_hier0_bF_buf8));
BUFX4 BUFX4_10 ( .A(u0_u0__abc_72207_new_n354_), .Y(u0_u0__abc_72207_new_n354__bF_buf4));
BUFX4 BUFX4_100 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf72));
BUFX4 BUFX4_101 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf71));
BUFX4 BUFX4_102 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf70));
BUFX4 BUFX4_103 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf69));
BUFX4 BUFX4_104 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf68));
BUFX4 BUFX4_105 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf67));
BUFX4 BUFX4_106 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf66));
BUFX4 BUFX4_107 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf65));
BUFX4 BUFX4_108 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf64));
BUFX4 BUFX4_109 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf63));
BUFX4 BUFX4_11 ( .A(u0_u0__abc_72207_new_n354_), .Y(u0_u0__abc_72207_new_n354__bF_buf3));
BUFX4 BUFX4_110 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf62));
BUFX4 BUFX4_111 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf61));
BUFX4 BUFX4_112 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf60));
BUFX4 BUFX4_113 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf59));
BUFX4 BUFX4_114 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf58));
BUFX4 BUFX4_115 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf57));
BUFX4 BUFX4_116 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf56));
BUFX4 BUFX4_117 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf55));
BUFX4 BUFX4_118 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf54));
BUFX4 BUFX4_119 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf53));
BUFX4 BUFX4_12 ( .A(u0_u0__abc_72207_new_n354_), .Y(u0_u0__abc_72207_new_n354__bF_buf2));
BUFX4 BUFX4_120 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf52));
BUFX4 BUFX4_121 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf51));
BUFX4 BUFX4_122 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf50));
BUFX4 BUFX4_123 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf49));
BUFX4 BUFX4_124 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf48));
BUFX4 BUFX4_125 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf47));
BUFX4 BUFX4_126 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf46));
BUFX4 BUFX4_127 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf45));
BUFX4 BUFX4_128 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf44));
BUFX4 BUFX4_129 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf43));
BUFX4 BUFX4_13 ( .A(u0_u0__abc_72207_new_n354_), .Y(u0_u0__abc_72207_new_n354__bF_buf1));
BUFX4 BUFX4_130 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf42));
BUFX4 BUFX4_131 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf41));
BUFX4 BUFX4_132 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf40));
BUFX4 BUFX4_133 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf39));
BUFX4 BUFX4_134 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf38));
BUFX4 BUFX4_135 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf37));
BUFX4 BUFX4_136 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf36));
BUFX4 BUFX4_137 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf35));
BUFX4 BUFX4_138 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf34));
BUFX4 BUFX4_139 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf33));
BUFX4 BUFX4_14 ( .A(u0_u0__abc_72207_new_n354_), .Y(u0_u0__abc_72207_new_n354__bF_buf0));
BUFX4 BUFX4_140 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf32));
BUFX4 BUFX4_141 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf31));
BUFX4 BUFX4_142 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf30));
BUFX4 BUFX4_143 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf29));
BUFX4 BUFX4_144 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf28));
BUFX4 BUFX4_145 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf27));
BUFX4 BUFX4_146 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf26));
BUFX4 BUFX4_147 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf25));
BUFX4 BUFX4_148 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf24));
BUFX4 BUFX4_149 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf23));
BUFX4 BUFX4_15 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf3_));
BUFX4 BUFX4_150 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf22));
BUFX4 BUFX4_151 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf21));
BUFX4 BUFX4_152 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf20));
BUFX4 BUFX4_153 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf19));
BUFX4 BUFX4_154 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf18));
BUFX4 BUFX4_155 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf17));
BUFX4 BUFX4_156 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf16));
BUFX4 BUFX4_157 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf15));
BUFX4 BUFX4_158 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf14));
BUFX4 BUFX4_159 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf13));
BUFX4 BUFX4_16 ( .A(row_adr_7_), .Y(row_adr_7_bF_buf2_));
BUFX4 BUFX4_160 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf12));
BUFX4 BUFX4_161 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf11));
BUFX4 BUFX4_162 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf10));
BUFX4 BUFX4_163 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf9));
BUFX4 BUFX4_164 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf8));
BUFX4 BUFX4_165 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf7));
BUFX4 BUFX4_166 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf6));
BUFX4 BUFX4_167 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf5));
BUFX4 BUFX4_168 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf4));
BUFX4 BUFX4_169 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf3));
BUFX4 BUFX4_17 ( .A(u3_u0__abc_75526_new_n876_), .Y(u3_u0__abc_75526_new_n876__bF_buf7));
BUFX4 BUFX4_170 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf2));
BUFX4 BUFX4_171 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf1));
BUFX4 BUFX4_172 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf0));
BUFX4 BUFX4_173 ( .A(u2_u0__abc_74955_new_n137_), .Y(u2_u0__abc_74955_new_n137__bF_buf4));
BUFX4 BUFX4_174 ( .A(u2_u0__abc_74955_new_n137_), .Y(u2_u0__abc_74955_new_n137__bF_buf3));
BUFX4 BUFX4_175 ( .A(u2_u0__abc_74955_new_n137_), .Y(u2_u0__abc_74955_new_n137__bF_buf2));
BUFX4 BUFX4_176 ( .A(u2_u0__abc_74955_new_n137_), .Y(u2_u0__abc_74955_new_n137__bF_buf0));
BUFX4 BUFX4_177 ( .A(u0__abc_76628_new_n4547_), .Y(u0__abc_76628_new_n4547__bF_buf4));
BUFX4 BUFX4_178 ( .A(u0__abc_76628_new_n4547_), .Y(u0__abc_76628_new_n4547__bF_buf3));
BUFX4 BUFX4_179 ( .A(u0__abc_76628_new_n4547_), .Y(u0__abc_76628_new_n4547__bF_buf2));
BUFX4 BUFX4_18 ( .A(u3_u0__abc_75526_new_n876_), .Y(u3_u0__abc_75526_new_n876__bF_buf6));
BUFX4 BUFX4_180 ( .A(u0__abc_76628_new_n4547_), .Y(u0__abc_76628_new_n4547__bF_buf1));
BUFX4 BUFX4_181 ( .A(u0__abc_76628_new_n4547_), .Y(u0__abc_76628_new_n4547__bF_buf0));
BUFX4 BUFX4_182 ( .A(u5__abc_81276_new_n479_), .Y(u5__abc_81276_new_n479__bF_buf3));
BUFX4 BUFX4_183 ( .A(u5__abc_81276_new_n479_), .Y(u5__abc_81276_new_n479__bF_buf2));
BUFX4 BUFX4_184 ( .A(u3_u0__abc_75526_new_n382_), .Y(u3_u0__abc_75526_new_n382__bF_buf7));
BUFX4 BUFX4_185 ( .A(u3_u0__abc_75526_new_n382_), .Y(u3_u0__abc_75526_new_n382__bF_buf6));
BUFX4 BUFX4_186 ( .A(u3_u0__abc_75526_new_n382_), .Y(u3_u0__abc_75526_new_n382__bF_buf5));
BUFX4 BUFX4_187 ( .A(u3_u0__abc_75526_new_n382_), .Y(u3_u0__abc_75526_new_n382__bF_buf4));
BUFX4 BUFX4_188 ( .A(u3_u0__abc_75526_new_n382_), .Y(u3_u0__abc_75526_new_n382__bF_buf3));
BUFX4 BUFX4_189 ( .A(u3_u0__abc_75526_new_n382_), .Y(u3_u0__abc_75526_new_n382__bF_buf2));
BUFX4 BUFX4_19 ( .A(u3_u0__abc_75526_new_n876_), .Y(u3_u0__abc_75526_new_n876__bF_buf5));
BUFX4 BUFX4_190 ( .A(u3_u0__abc_75526_new_n382_), .Y(u3_u0__abc_75526_new_n382__bF_buf1));
BUFX4 BUFX4_191 ( .A(u3_u0__abc_75526_new_n382_), .Y(u3_u0__abc_75526_new_n382__bF_buf0));
BUFX4 BUFX4_192 ( .A(u3__abc_74070_new_n277_), .Y(u3__abc_74070_new_n277__bF_buf5));
BUFX4 BUFX4_193 ( .A(u3__abc_74070_new_n277_), .Y(u3__abc_74070_new_n277__bF_buf4));
BUFX4 BUFX4_194 ( .A(u3__abc_74070_new_n277_), .Y(u3__abc_74070_new_n277__bF_buf3));
BUFX4 BUFX4_195 ( .A(u3__abc_74070_new_n277_), .Y(u3__abc_74070_new_n277__bF_buf2));
BUFX4 BUFX4_196 ( .A(u3__abc_74070_new_n277_), .Y(u3__abc_74070_new_n277__bF_buf1));
BUFX4 BUFX4_197 ( .A(u3__abc_74070_new_n277_), .Y(u3__abc_74070_new_n277__bF_buf0));
BUFX4 BUFX4_198 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf5_));
BUFX4 BUFX4_199 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf4_));
BUFX4 BUFX4_2 ( .A(clk_i), .Y(clk_i_hier0_bF_buf7));
BUFX4 BUFX4_20 ( .A(u3_u0__abc_75526_new_n876_), .Y(u3_u0__abc_75526_new_n876__bF_buf4));
BUFX4 BUFX4_200 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf3_));
BUFX4 BUFX4_201 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf2_));
BUFX4 BUFX4_202 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf1_));
BUFX4 BUFX4_203 ( .A(spec_req_cs_5_), .Y(spec_req_cs_5_bF_buf0_));
BUFX4 BUFX4_204 ( .A(u0__abc_76628_new_n2742_), .Y(u0__abc_76628_new_n2742__bF_buf5));
BUFX4 BUFX4_205 ( .A(u0__abc_76628_new_n2742_), .Y(u0__abc_76628_new_n2742__bF_buf4));
BUFX4 BUFX4_206 ( .A(u0__abc_76628_new_n2742_), .Y(u0__abc_76628_new_n2742__bF_buf3));
BUFX4 BUFX4_207 ( .A(u0__abc_76628_new_n2742_), .Y(u0__abc_76628_new_n2742__bF_buf2));
BUFX4 BUFX4_208 ( .A(u0__abc_76628_new_n2742_), .Y(u0__abc_76628_new_n2742__bF_buf1));
BUFX4 BUFX4_209 ( .A(u0__abc_76628_new_n2742_), .Y(u0__abc_76628_new_n2742__bF_buf0));
BUFX4 BUFX4_21 ( .A(u3_u0__abc_75526_new_n876_), .Y(u3_u0__abc_75526_new_n876__bF_buf3));
BUFX4 BUFX4_210 ( .A(u0__abc_76628_new_n4503_), .Y(u0__abc_76628_new_n4503__bF_buf4));
BUFX4 BUFX4_211 ( .A(u0__abc_76628_new_n4503_), .Y(u0__abc_76628_new_n4503__bF_buf3));
BUFX4 BUFX4_212 ( .A(u0__abc_76628_new_n4503_), .Y(u0__abc_76628_new_n4503__bF_buf2));
BUFX4 BUFX4_213 ( .A(u0__abc_76628_new_n4503_), .Y(u0__abc_76628_new_n4503__bF_buf1));
BUFX4 BUFX4_214 ( .A(u0__abc_76628_new_n4503_), .Y(u0__abc_76628_new_n4503__bF_buf0));
BUFX4 BUFX4_215 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf5_));
BUFX4 BUFX4_216 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf4_));
BUFX4 BUFX4_217 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf3_));
BUFX4 BUFX4_218 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf2_));
BUFX4 BUFX4_219 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf1_));
BUFX4 BUFX4_22 ( .A(u3_u0__abc_75526_new_n876_), .Y(u3_u0__abc_75526_new_n876__bF_buf2));
BUFX4 BUFX4_220 ( .A(spec_req_cs_2_), .Y(spec_req_cs_2_bF_buf0_));
BUFX4 BUFX4_221 ( .A(csc_5_), .Y(csc_5_bF_buf4_));
BUFX4 BUFX4_222 ( .A(csc_5_), .Y(csc_5_bF_buf3_));
BUFX4 BUFX4_223 ( .A(csc_5_), .Y(csc_5_bF_buf2_));
BUFX4 BUFX4_224 ( .A(csc_5_), .Y(csc_5_bF_buf1_));
BUFX4 BUFX4_225 ( .A(csc_5_), .Y(csc_5_bF_buf0_));
BUFX4 BUFX4_226 ( .A(u0__abc_76628_new_n4500_), .Y(u0__abc_76628_new_n4500__bF_buf4));
BUFX4 BUFX4_227 ( .A(u0__abc_76628_new_n4500_), .Y(u0__abc_76628_new_n4500__bF_buf3));
BUFX4 BUFX4_228 ( .A(u0__abc_76628_new_n4500_), .Y(u0__abc_76628_new_n4500__bF_buf2));
BUFX4 BUFX4_229 ( .A(u0__abc_76628_new_n4500_), .Y(u0__abc_76628_new_n4500__bF_buf1));
BUFX4 BUFX4_23 ( .A(u3_u0__abc_75526_new_n876_), .Y(u3_u0__abc_75526_new_n876__bF_buf1));
BUFX4 BUFX4_230 ( .A(u0__abc_76628_new_n4500_), .Y(u0__abc_76628_new_n4500__bF_buf0));
BUFX4 BUFX4_231 ( .A(u0__abc_76628_new_n4438_), .Y(u0__abc_76628_new_n4438__bF_buf3));
BUFX4 BUFX4_232 ( .A(u0__abc_76628_new_n4438_), .Y(u0__abc_76628_new_n4438__bF_buf2));
BUFX4 BUFX4_233 ( .A(u1__abc_73140_new_n563_), .Y(u1__abc_73140_new_n563__bF_buf3));
BUFX4 BUFX4_234 ( .A(u1__abc_73140_new_n563_), .Y(u1__abc_73140_new_n563__bF_buf2));
BUFX4 BUFX4_235 ( .A(u1__abc_73140_new_n563_), .Y(u1__abc_73140_new_n563__bF_buf1));
BUFX4 BUFX4_236 ( .A(u1__abc_73140_new_n563_), .Y(u1__abc_73140_new_n563__bF_buf0));
BUFX4 BUFX4_237 ( .A(u0_u1__0lmr_req_we_0_0_), .Y(u0_u1__0lmr_req_we_0_0_bF_buf7_));
BUFX4 BUFX4_238 ( .A(u0_u1__0lmr_req_we_0_0_), .Y(u0_u1__0lmr_req_we_0_0_bF_buf6_));
BUFX4 BUFX4_239 ( .A(u0_u1__0lmr_req_we_0_0_), .Y(u0_u1__0lmr_req_we_0_0_bF_buf5_));
BUFX4 BUFX4_24 ( .A(u3_u0__abc_75526_new_n876_), .Y(u3_u0__abc_75526_new_n876__bF_buf0));
BUFX4 BUFX4_240 ( .A(u0_u1__0lmr_req_we_0_0_), .Y(u0_u1__0lmr_req_we_0_0_bF_buf4_));
BUFX4 BUFX4_241 ( .A(u0_u1__0lmr_req_we_0_0_), .Y(u0_u1__0lmr_req_we_0_0_bF_buf3_));
BUFX4 BUFX4_242 ( .A(u0_u1__0lmr_req_we_0_0_), .Y(u0_u1__0lmr_req_we_0_0_bF_buf2_));
BUFX4 BUFX4_243 ( .A(u0_u1__0lmr_req_we_0_0_), .Y(u0_u1__0lmr_req_we_0_0_bF_buf1_));
BUFX4 BUFX4_244 ( .A(u0_u1__0lmr_req_we_0_0_), .Y(u0_u1__0lmr_req_we_0_0_bF_buf0_));
BUFX4 BUFX4_245 ( .A(u1__abc_73140_new_n275_), .Y(u1__abc_73140_new_n275__bF_buf4));
BUFX4 BUFX4_246 ( .A(u1__abc_73140_new_n275_), .Y(u1__abc_73140_new_n275__bF_buf3));
BUFX4 BUFX4_247 ( .A(u1__abc_73140_new_n275_), .Y(u1__abc_73140_new_n275__bF_buf2));
BUFX4 BUFX4_248 ( .A(u1__abc_73140_new_n904_), .Y(u1__abc_73140_new_n904__bF_buf4));
BUFX4 BUFX4_249 ( .A(u1__abc_73140_new_n904_), .Y(u1__abc_73140_new_n904__bF_buf3));
BUFX4 BUFX4_25 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf3_));
BUFX4 BUFX4_250 ( .A(u1__abc_73140_new_n904_), .Y(u1__abc_73140_new_n904__bF_buf2));
BUFX4 BUFX4_251 ( .A(u1__abc_73140_new_n904_), .Y(u1__abc_73140_new_n904__bF_buf1));
BUFX4 BUFX4_252 ( .A(u1__abc_73140_new_n904_), .Y(u1__abc_73140_new_n904__bF_buf0));
BUFX4 BUFX4_253 ( .A(u5__abc_81276_new_n523_), .Y(u5__abc_81276_new_n523__bF_buf7));
BUFX4 BUFX4_254 ( .A(u5__abc_81276_new_n523_), .Y(u5__abc_81276_new_n523__bF_buf6));
BUFX4 BUFX4_255 ( .A(u5__abc_81276_new_n523_), .Y(u5__abc_81276_new_n523__bF_buf5));
BUFX4 BUFX4_256 ( .A(u5__abc_81276_new_n523_), .Y(u5__abc_81276_new_n523__bF_buf4));
BUFX4 BUFX4_257 ( .A(u5__abc_81276_new_n523_), .Y(u5__abc_81276_new_n523__bF_buf3));
BUFX4 BUFX4_258 ( .A(u5__abc_81276_new_n523_), .Y(u5__abc_81276_new_n523__bF_buf2));
BUFX4 BUFX4_259 ( .A(u5__abc_81276_new_n523_), .Y(u5__abc_81276_new_n523__bF_buf1));
BUFX4 BUFX4_26 ( .A(row_adr_10_), .Y(row_adr_10_bF_buf2_));
BUFX4 BUFX4_260 ( .A(u5__abc_81276_new_n523_), .Y(u5__abc_81276_new_n523__bF_buf0));
BUFX4 BUFX4_261 ( .A(u5__abc_81276_new_n3215_), .Y(u5__abc_81276_new_n3215__bF_buf4));
BUFX4 BUFX4_262 ( .A(u5__abc_81276_new_n3215_), .Y(u5__abc_81276_new_n3215__bF_buf3));
BUFX4 BUFX4_263 ( .A(u5__abc_81276_new_n464_), .Y(u5__abc_81276_new_n464__bF_buf3));
BUFX4 BUFX4_264 ( .A(u5__abc_81276_new_n464_), .Y(u5__abc_81276_new_n464__bF_buf2));
BUFX4 BUFX4_265 ( .A(u5__abc_81276_new_n464_), .Y(u5__abc_81276_new_n464__bF_buf1));
BUFX4 BUFX4_266 ( .A(u0_u0__abc_72207_new_n224_), .Y(u0_u0__abc_72207_new_n224__bF_buf4));
BUFX4 BUFX4_267 ( .A(u0_u0__abc_72207_new_n224_), .Y(u0_u0__abc_72207_new_n224__bF_buf3));
BUFX4 BUFX4_268 ( .A(u0_u0__abc_72207_new_n224_), .Y(u0_u0__abc_72207_new_n224__bF_buf2));
BUFX4 BUFX4_269 ( .A(u0_u0__abc_72207_new_n224_), .Y(u0_u0__abc_72207_new_n224__bF_buf1));
BUFX4 BUFX4_27 ( .A(u0__abc_76628_new_n1173_), .Y(u0__abc_76628_new_n1173__bF_buf5));
BUFX4 BUFX4_270 ( .A(u0_u0__abc_72207_new_n224_), .Y(u0_u0__abc_72207_new_n224__bF_buf0));
BUFX4 BUFX4_271 ( .A(u3_u0__abc_75526_new_n708_), .Y(u3_u0__abc_75526_new_n708__bF_buf7));
BUFX4 BUFX4_272 ( .A(u3_u0__abc_75526_new_n708_), .Y(u3_u0__abc_75526_new_n708__bF_buf6));
BUFX4 BUFX4_273 ( .A(u3_u0__abc_75526_new_n708_), .Y(u3_u0__abc_75526_new_n708__bF_buf5));
BUFX4 BUFX4_274 ( .A(u3_u0__abc_75526_new_n708_), .Y(u3_u0__abc_75526_new_n708__bF_buf4));
BUFX4 BUFX4_275 ( .A(u3_u0__abc_75526_new_n708_), .Y(u3_u0__abc_75526_new_n708__bF_buf3));
BUFX4 BUFX4_276 ( .A(u3_u0__abc_75526_new_n708_), .Y(u3_u0__abc_75526_new_n708__bF_buf2));
BUFX4 BUFX4_277 ( .A(u3_u0__abc_75526_new_n708_), .Y(u3_u0__abc_75526_new_n708__bF_buf1));
BUFX4 BUFX4_278 ( .A(u3_u0__abc_75526_new_n708_), .Y(u3_u0__abc_75526_new_n708__bF_buf0));
BUFX4 BUFX4_279 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf3_));
BUFX4 BUFX4_28 ( .A(u0__abc_76628_new_n1173_), .Y(u0__abc_76628_new_n1173__bF_buf4));
BUFX4 BUFX4_280 ( .A(row_adr_9_), .Y(row_adr_9_bF_buf2_));
BUFX4 BUFX4_281 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf3_));
BUFX4 BUFX4_282 ( .A(row_adr_12_), .Y(row_adr_12_bF_buf2_));
BUFX4 BUFX4_283 ( .A(u0__abc_76628_new_n1175_), .Y(u0__abc_76628_new_n1175__bF_buf5));
BUFX4 BUFX4_284 ( .A(u0__abc_76628_new_n1175_), .Y(u0__abc_76628_new_n1175__bF_buf4));
BUFX4 BUFX4_285 ( .A(u0__abc_76628_new_n1175_), .Y(u0__abc_76628_new_n1175__bF_buf3));
BUFX4 BUFX4_286 ( .A(u0__abc_76628_new_n1175_), .Y(u0__abc_76628_new_n1175__bF_buf2));
BUFX4 BUFX4_287 ( .A(u0__abc_76628_new_n1175_), .Y(u0__abc_76628_new_n1175__bF_buf1));
BUFX4 BUFX4_288 ( .A(u0__abc_76628_new_n1175_), .Y(u0__abc_76628_new_n1175__bF_buf0));
BUFX4 BUFX4_289 ( .A(u0__abc_76628_new_n2724_), .Y(u0__abc_76628_new_n2724__bF_buf5));
BUFX4 BUFX4_29 ( .A(u0__abc_76628_new_n1173_), .Y(u0__abc_76628_new_n1173__bF_buf3));
BUFX4 BUFX4_290 ( .A(u0__abc_76628_new_n2724_), .Y(u0__abc_76628_new_n2724__bF_buf4));
BUFX4 BUFX4_291 ( .A(u0__abc_76628_new_n2724_), .Y(u0__abc_76628_new_n2724__bF_buf3));
BUFX4 BUFX4_292 ( .A(u0__abc_76628_new_n2724_), .Y(u0__abc_76628_new_n2724__bF_buf2));
BUFX4 BUFX4_293 ( .A(u0__abc_76628_new_n2724_), .Y(u0__abc_76628_new_n2724__bF_buf1));
BUFX4 BUFX4_294 ( .A(u0__abc_76628_new_n2724_), .Y(u0__abc_76628_new_n2724__bF_buf0));
BUFX4 BUFX4_295 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf3_));
BUFX4 BUFX4_296 ( .A(row_adr_6_), .Y(row_adr_6_bF_buf2_));
BUFX4 BUFX4_297 ( .A(u0__abc_76628_new_n1172_), .Y(u0__abc_76628_new_n1172__bF_buf5));
BUFX4 BUFX4_298 ( .A(u0__abc_76628_new_n1172_), .Y(u0__abc_76628_new_n1172__bF_buf4));
BUFX4 BUFX4_299 ( .A(u0__abc_76628_new_n1172_), .Y(u0__abc_76628_new_n1172__bF_buf3));
BUFX4 BUFX4_3 ( .A(clk_i), .Y(clk_i_hier0_bF_buf6));
BUFX4 BUFX4_30 ( .A(u0__abc_76628_new_n1173_), .Y(u0__abc_76628_new_n1173__bF_buf2));
BUFX4 BUFX4_300 ( .A(u0__abc_76628_new_n1172_), .Y(u0__abc_76628_new_n1172__bF_buf2));
BUFX4 BUFX4_301 ( .A(u0__abc_76628_new_n1172_), .Y(u0__abc_76628_new_n1172__bF_buf1));
BUFX4 BUFX4_302 ( .A(u0__abc_76628_new_n1172_), .Y(u0__abc_76628_new_n1172__bF_buf0));
BUFX4 BUFX4_303 ( .A(u0__abc_76628_new_n4523_), .Y(u0__abc_76628_new_n4523__bF_buf4));
BUFX4 BUFX4_304 ( .A(u0__abc_76628_new_n4523_), .Y(u0__abc_76628_new_n4523__bF_buf3));
BUFX4 BUFX4_305 ( .A(u0__abc_76628_new_n4523_), .Y(u0__abc_76628_new_n4523__bF_buf2));
BUFX4 BUFX4_306 ( .A(u0__abc_76628_new_n4523_), .Y(u0__abc_76628_new_n4523__bF_buf1));
BUFX4 BUFX4_307 ( .A(u0__abc_76628_new_n4523_), .Y(u0__abc_76628_new_n4523__bF_buf0));
BUFX4 BUFX4_308 ( .A(lmr_sel), .Y(lmr_sel_bF_buf6));
BUFX4 BUFX4_309 ( .A(lmr_sel), .Y(lmr_sel_bF_buf5));
BUFX4 BUFX4_31 ( .A(u0__abc_76628_new_n1173_), .Y(u0__abc_76628_new_n1173__bF_buf1));
BUFX4 BUFX4_310 ( .A(lmr_sel), .Y(lmr_sel_bF_buf4));
BUFX4 BUFX4_311 ( .A(lmr_sel), .Y(lmr_sel_bF_buf3));
BUFX4 BUFX4_312 ( .A(lmr_sel), .Y(lmr_sel_bF_buf2));
BUFX4 BUFX4_313 ( .A(lmr_sel), .Y(lmr_sel_bF_buf1));
BUFX4 BUFX4_314 ( .A(lmr_sel), .Y(lmr_sel_bF_buf0));
BUFX4 BUFX4_315 ( .A(u0__abc_76628_new_n1169_), .Y(u0__abc_76628_new_n1169__bF_buf6));
BUFX4 BUFX4_316 ( .A(u0__abc_76628_new_n1169_), .Y(u0__abc_76628_new_n1169__bF_buf5));
BUFX4 BUFX4_317 ( .A(u0__abc_76628_new_n1169_), .Y(u0__abc_76628_new_n1169__bF_buf4));
BUFX4 BUFX4_318 ( .A(u0__abc_76628_new_n1169_), .Y(u0__abc_76628_new_n1169__bF_buf3));
BUFX4 BUFX4_319 ( .A(u0__abc_76628_new_n1169_), .Y(u0__abc_76628_new_n1169__bF_buf2));
BUFX4 BUFX4_32 ( .A(u0__abc_76628_new_n1173_), .Y(u0__abc_76628_new_n1173__bF_buf0));
BUFX4 BUFX4_320 ( .A(u0__abc_76628_new_n1169_), .Y(u0__abc_76628_new_n1169__bF_buf1));
BUFX4 BUFX4_321 ( .A(u0__abc_76628_new_n1169_), .Y(u0__abc_76628_new_n1169__bF_buf0));
BUFX4 BUFX4_322 ( .A(u0__abc_76628_new_n4558_), .Y(u0__abc_76628_new_n4558__bF_buf4));
BUFX4 BUFX4_323 ( .A(u0__abc_76628_new_n4558_), .Y(u0__abc_76628_new_n4558__bF_buf3));
BUFX4 BUFX4_324 ( .A(u0__abc_76628_new_n4558_), .Y(u0__abc_76628_new_n4558__bF_buf2));
BUFX4 BUFX4_325 ( .A(u0__abc_76628_new_n4558_), .Y(u0__abc_76628_new_n4558__bF_buf1));
BUFX4 BUFX4_326 ( .A(u0__abc_76628_new_n4558_), .Y(u0__abc_76628_new_n4558__bF_buf0));
BUFX4 BUFX4_327 ( .A(u5__abc_81276_new_n417_), .Y(u5__abc_81276_new_n417__bF_buf3));
BUFX4 BUFX4_328 ( .A(u5__abc_81276_new_n417_), .Y(u5__abc_81276_new_n417__bF_buf2));
BUFX4 BUFX4_329 ( .A(u5__abc_81276_new_n417_), .Y(u5__abc_81276_new_n417__bF_buf1));
BUFX4 BUFX4_33 ( .A(u0__abc_76628_new_n4562_), .Y(u0__abc_76628_new_n4562__bF_buf4));
BUFX4 BUFX4_330 ( .A(u2_u1__abc_74955_new_n137_), .Y(u2_u1__abc_74955_new_n137__bF_buf4));
BUFX4 BUFX4_331 ( .A(u2_u1__abc_74955_new_n137_), .Y(u2_u1__abc_74955_new_n137__bF_buf3));
BUFX4 BUFX4_332 ( .A(u2_u1__abc_74955_new_n137_), .Y(u2_u1__abc_74955_new_n137__bF_buf2));
BUFX4 BUFX4_333 ( .A(u2_u1__abc_74955_new_n137_), .Y(u2_u1__abc_74955_new_n137__bF_buf0));
BUFX4 BUFX4_334 ( .A(u0__abc_76628_new_n2718_), .Y(u0__abc_76628_new_n2718__bF_buf5));
BUFX4 BUFX4_335 ( .A(u0__abc_76628_new_n2718_), .Y(u0__abc_76628_new_n2718__bF_buf4));
BUFX4 BUFX4_336 ( .A(u0__abc_76628_new_n2718_), .Y(u0__abc_76628_new_n2718__bF_buf3));
BUFX4 BUFX4_337 ( .A(u0__abc_76628_new_n2718_), .Y(u0__abc_76628_new_n2718__bF_buf2));
BUFX4 BUFX4_338 ( .A(u0__abc_76628_new_n2718_), .Y(u0__abc_76628_new_n2718__bF_buf1));
BUFX4 BUFX4_339 ( .A(u0__abc_76628_new_n2718_), .Y(u0__abc_76628_new_n2718__bF_buf0));
BUFX4 BUFX4_34 ( .A(u0__abc_76628_new_n4562_), .Y(u0__abc_76628_new_n4562__bF_buf3));
BUFX4 BUFX4_340 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf3_));
BUFX4 BUFX4_341 ( .A(row_adr_3_), .Y(row_adr_3_bF_buf2_));
BUFX4 BUFX4_342 ( .A(u0__abc_76628_new_n4520_), .Y(u0__abc_76628_new_n4520__bF_buf4));
BUFX4 BUFX4_343 ( .A(u0__abc_76628_new_n4520_), .Y(u0__abc_76628_new_n4520__bF_buf3));
BUFX4 BUFX4_344 ( .A(u0__abc_76628_new_n4520_), .Y(u0__abc_76628_new_n4520__bF_buf2));
BUFX4 BUFX4_345 ( .A(u0__abc_76628_new_n4520_), .Y(u0__abc_76628_new_n4520__bF_buf1));
BUFX4 BUFX4_346 ( .A(u0__abc_76628_new_n4520_), .Y(u0__abc_76628_new_n4520__bF_buf0));
BUFX4 BUFX4_347 ( .A(u0__abc_76628_new_n4517_), .Y(u0__abc_76628_new_n4517__bF_buf4));
BUFX4 BUFX4_348 ( .A(u0__abc_76628_new_n4517_), .Y(u0__abc_76628_new_n4517__bF_buf3));
BUFX4 BUFX4_349 ( .A(u0__abc_76628_new_n4517_), .Y(u0__abc_76628_new_n4517__bF_buf2));
BUFX4 BUFX4_35 ( .A(u0__abc_76628_new_n4562_), .Y(u0__abc_76628_new_n4562__bF_buf2));
BUFX4 BUFX4_350 ( .A(u0__abc_76628_new_n4517_), .Y(u0__abc_76628_new_n4517__bF_buf1));
BUFX4 BUFX4_351 ( .A(u0__abc_76628_new_n4517_), .Y(u0__abc_76628_new_n4517__bF_buf0));
BUFX4 BUFX4_352 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf10));
BUFX4 BUFX4_353 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf9));
BUFX4 BUFX4_354 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf8));
BUFX4 BUFX4_355 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf7));
BUFX4 BUFX4_356 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf6));
BUFX4 BUFX4_357 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf5));
BUFX4 BUFX4_358 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf4));
BUFX4 BUFX4_359 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf3));
BUFX4 BUFX4_36 ( .A(u0__abc_76628_new_n4562_), .Y(u0__abc_76628_new_n4562__bF_buf1));
BUFX4 BUFX4_360 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf2));
BUFX4 BUFX4_361 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf1));
BUFX4 BUFX4_362 ( .A(u5__abc_81276_new_n490_), .Y(u5__abc_81276_new_n490__bF_buf0));
BUFX4 BUFX4_363 ( .A(row_adr_0_), .Y(row_adr_0_bF_buf2_));
BUFX4 BUFX4_364 ( .A(u5__abc_81276_new_n449_), .Y(u5__abc_81276_new_n449__bF_buf7));
BUFX4 BUFX4_365 ( .A(u5__abc_81276_new_n449_), .Y(u5__abc_81276_new_n449__bF_buf6));
BUFX4 BUFX4_366 ( .A(u5__abc_81276_new_n449_), .Y(u5__abc_81276_new_n449__bF_buf5));
BUFX4 BUFX4_367 ( .A(u5__abc_81276_new_n449_), .Y(u5__abc_81276_new_n449__bF_buf4));
BUFX4 BUFX4_368 ( .A(u5__abc_81276_new_n449_), .Y(u5__abc_81276_new_n449__bF_buf3));
BUFX4 BUFX4_369 ( .A(u5__abc_81276_new_n449_), .Y(u5__abc_81276_new_n449__bF_buf2));
BUFX4 BUFX4_37 ( .A(u0__abc_76628_new_n4562_), .Y(u0__abc_76628_new_n4562__bF_buf0));
BUFX4 BUFX4_370 ( .A(u5__abc_81276_new_n449_), .Y(u5__abc_81276_new_n449__bF_buf1));
BUFX4 BUFX4_371 ( .A(u5__abc_81276_new_n449_), .Y(u5__abc_81276_new_n449__bF_buf0));
BUFX4 BUFX4_372 ( .A(cs_le), .Y(cs_le_bF_buf4));
BUFX4 BUFX4_373 ( .A(cs_le), .Y(cs_le_bF_buf3));
BUFX4 BUFX4_374 ( .A(cs_le), .Y(cs_le_bF_buf2));
BUFX4 BUFX4_375 ( .A(cs_le), .Y(cs_le_bF_buf1));
BUFX4 BUFX4_376 ( .A(u0__abc_76628_new_n4549_), .Y(u0__abc_76628_new_n4549__bF_buf4));
BUFX4 BUFX4_377 ( .A(u0__abc_76628_new_n4549_), .Y(u0__abc_76628_new_n4549__bF_buf3));
BUFX4 BUFX4_378 ( .A(u0__abc_76628_new_n4549_), .Y(u0__abc_76628_new_n4549__bF_buf2));
BUFX4 BUFX4_379 ( .A(u0__abc_76628_new_n4549_), .Y(u0__abc_76628_new_n4549__bF_buf1));
BUFX4 BUFX4_38 ( .A(u0__abc_76628_new_n2722_), .Y(u0__abc_76628_new_n2722__bF_buf5));
BUFX4 BUFX4_380 ( .A(u0__abc_76628_new_n4549_), .Y(u0__abc_76628_new_n4549__bF_buf0));
BUFX4 BUFX4_381 ( .A(u3__abc_74070_new_n279_), .Y(u3__abc_74070_new_n279__bF_buf5));
BUFX4 BUFX4_382 ( .A(u3__abc_74070_new_n279_), .Y(u3__abc_74070_new_n279__bF_buf4));
BUFX4 BUFX4_383 ( .A(u3__abc_74070_new_n279_), .Y(u3__abc_74070_new_n279__bF_buf3));
BUFX4 BUFX4_384 ( .A(u3__abc_74070_new_n279_), .Y(u3__abc_74070_new_n279__bF_buf2));
BUFX4 BUFX4_385 ( .A(u3__abc_74070_new_n279_), .Y(u3__abc_74070_new_n279__bF_buf1));
BUFX4 BUFX4_386 ( .A(u3__abc_74070_new_n279_), .Y(u3__abc_74070_new_n279__bF_buf0));
BUFX4 BUFX4_387 ( .A(u0_u1__abc_72579_new_n219_), .Y(u0_u1__abc_72579_new_n219__bF_buf7));
BUFX4 BUFX4_388 ( .A(u0_u1__abc_72579_new_n219_), .Y(u0_u1__abc_72579_new_n219__bF_buf6));
BUFX4 BUFX4_389 ( .A(u0_u1__abc_72579_new_n219_), .Y(u0_u1__abc_72579_new_n219__bF_buf5));
BUFX4 BUFX4_39 ( .A(u0__abc_76628_new_n2722_), .Y(u0__abc_76628_new_n2722__bF_buf4));
BUFX4 BUFX4_390 ( .A(u0_u1__abc_72579_new_n219_), .Y(u0_u1__abc_72579_new_n219__bF_buf4));
BUFX4 BUFX4_391 ( .A(u0_u1__abc_72579_new_n219_), .Y(u0_u1__abc_72579_new_n219__bF_buf3));
BUFX4 BUFX4_392 ( .A(u0_u1__abc_72579_new_n219_), .Y(u0_u1__abc_72579_new_n219__bF_buf2));
BUFX4 BUFX4_393 ( .A(u0_u1__abc_72579_new_n219_), .Y(u0_u1__abc_72579_new_n219__bF_buf1));
BUFX4 BUFX4_394 ( .A(u0_u1__abc_72579_new_n219_), .Y(u0_u1__abc_72579_new_n219__bF_buf0));
BUFX4 BUFX4_395 ( .A(next_adr), .Y(next_adr_bF_buf4));
BUFX4 BUFX4_396 ( .A(next_adr), .Y(next_adr_bF_buf3));
BUFX4 BUFX4_397 ( .A(next_adr), .Y(next_adr_bF_buf2));
BUFX4 BUFX4_398 ( .A(next_adr), .Y(next_adr_bF_buf1));
BUFX4 BUFX4_399 ( .A(next_adr), .Y(next_adr_bF_buf0));
BUFX4 BUFX4_4 ( .A(clk_i), .Y(clk_i_hier0_bF_buf5));
BUFX4 BUFX4_40 ( .A(u0__abc_76628_new_n2722_), .Y(u0__abc_76628_new_n2722__bF_buf3));
BUFX4 BUFX4_400 ( .A(u6__abc_85257_new_n145_), .Y(u6__abc_85257_new_n145__bF_buf5));
BUFX4 BUFX4_401 ( .A(u6__abc_85257_new_n145_), .Y(u6__abc_85257_new_n145__bF_buf4));
BUFX4 BUFX4_402 ( .A(u6__abc_85257_new_n145_), .Y(u6__abc_85257_new_n145__bF_buf3));
BUFX4 BUFX4_403 ( .A(u6__abc_85257_new_n145_), .Y(u6__abc_85257_new_n145__bF_buf2));
BUFX4 BUFX4_404 ( .A(u6__abc_85257_new_n145_), .Y(u6__abc_85257_new_n145__bF_buf1));
BUFX4 BUFX4_405 ( .A(u6__abc_85257_new_n145_), .Y(u6__abc_85257_new_n145__bF_buf0));
BUFX4 BUFX4_406 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf5_));
BUFX4 BUFX4_407 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf4_));
BUFX4 BUFX4_408 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf3_));
BUFX4 BUFX4_409 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf2_));
BUFX4 BUFX4_41 ( .A(u0__abc_76628_new_n2722_), .Y(u0__abc_76628_new_n2722__bF_buf2));
BUFX4 BUFX4_410 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf1_));
BUFX4 BUFX4_411 ( .A(spec_req_cs_4_), .Y(spec_req_cs_4_bF_buf0_));
BUFX4 BUFX4_412 ( .A(u0_cs0), .Y(u0_cs0_bF_buf5));
BUFX4 BUFX4_413 ( .A(u0_cs0), .Y(u0_cs0_bF_buf4));
BUFX4 BUFX4_414 ( .A(u0_cs0), .Y(u0_cs0_bF_buf3));
BUFX4 BUFX4_415 ( .A(u0_cs0), .Y(u0_cs0_bF_buf2));
BUFX4 BUFX4_416 ( .A(u0_cs0), .Y(u0_cs0_bF_buf1));
BUFX4 BUFX4_417 ( .A(u0_cs0), .Y(u0_cs0_bF_buf0));
BUFX4 BUFX4_418 ( .A(u0_cs1), .Y(u0_cs1_bF_buf5));
BUFX4 BUFX4_419 ( .A(u0_cs1), .Y(u0_cs1_bF_buf4));
BUFX4 BUFX4_42 ( .A(u0__abc_76628_new_n2722_), .Y(u0__abc_76628_new_n2722__bF_buf1));
BUFX4 BUFX4_420 ( .A(u0_cs1), .Y(u0_cs1_bF_buf3));
BUFX4 BUFX4_421 ( .A(u0_cs1), .Y(u0_cs1_bF_buf2));
BUFX4 BUFX4_422 ( .A(u0_cs1), .Y(u0_cs1_bF_buf1));
BUFX4 BUFX4_423 ( .A(u0_cs1), .Y(u0_cs1_bF_buf0));
BUFX4 BUFX4_424 ( .A(u5_tmr_done), .Y(u5_tmr_done_bF_buf1));
BUFX4 BUFX4_425 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf5_));
BUFX4 BUFX4_426 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf4_));
BUFX4 BUFX4_427 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf3_));
BUFX4 BUFX4_428 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf2_));
BUFX4 BUFX4_429 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf1_));
BUFX4 BUFX4_43 ( .A(u0__abc_76628_new_n2722_), .Y(u0__abc_76628_new_n2722__bF_buf0));
BUFX4 BUFX4_430 ( .A(spec_req_cs_1_), .Y(spec_req_cs_1_bF_buf0_));
BUFX4 BUFX4_431 ( .A(u1__abc_73140_new_n912_), .Y(u1__abc_73140_new_n912__bF_buf3));
BUFX4 BUFX4_432 ( .A(u1__abc_73140_new_n912_), .Y(u1__abc_73140_new_n912__bF_buf2));
BUFX4 BUFX4_433 ( .A(u1__abc_73140_new_n912_), .Y(u1__abc_73140_new_n912__bF_buf1));
BUFX4 BUFX4_434 ( .A(u1__abc_73140_new_n912_), .Y(u1__abc_73140_new_n912__bF_buf0));
BUFX4 BUFX4_435 ( .A(u3_u0__abc_75526_new_n563_), .Y(u3_u0__abc_75526_new_n563__bF_buf7));
BUFX4 BUFX4_436 ( .A(u3_u0__abc_75526_new_n563_), .Y(u3_u0__abc_75526_new_n563__bF_buf6));
BUFX4 BUFX4_437 ( .A(u3_u0__abc_75526_new_n563_), .Y(u3_u0__abc_75526_new_n563__bF_buf5));
BUFX4 BUFX4_438 ( .A(u3_u0__abc_75526_new_n563_), .Y(u3_u0__abc_75526_new_n563__bF_buf4));
BUFX4 BUFX4_439 ( .A(u3_u0__abc_75526_new_n563_), .Y(u3_u0__abc_75526_new_n563__bF_buf3));
BUFX4 BUFX4_44 ( .A(u0__abc_76628_new_n2719_), .Y(u0__abc_76628_new_n2719__bF_buf5));
BUFX4 BUFX4_440 ( .A(u3_u0__abc_75526_new_n563_), .Y(u3_u0__abc_75526_new_n563__bF_buf2));
BUFX4 BUFX4_441 ( .A(u3_u0__abc_75526_new_n563_), .Y(u3_u0__abc_75526_new_n563__bF_buf1));
BUFX4 BUFX4_442 ( .A(u3_u0__abc_75526_new_n563_), .Y(u3_u0__abc_75526_new_n563__bF_buf0));
BUFX4 BUFX4_443 ( .A(u0__abc_76628_new_n4437_), .Y(u0__abc_76628_new_n4437__bF_buf3));
BUFX4 BUFX4_444 ( .A(u0__abc_76628_new_n4437_), .Y(u0__abc_76628_new_n4437__bF_buf2));
BUFX4 BUFX4_445 ( .A(u0__abc_76628_new_n4437_), .Y(u0__abc_76628_new_n4437__bF_buf1));
BUFX4 BUFX4_446 ( .A(u1__abc_73140_new_n906_), .Y(u1__abc_73140_new_n906__bF_buf3));
BUFX4 BUFX4_447 ( .A(u1__abc_73140_new_n906_), .Y(u1__abc_73140_new_n906__bF_buf2));
BUFX4 BUFX4_448 ( .A(u1__abc_73140_new_n906_), .Y(u1__abc_73140_new_n906__bF_buf1));
BUFX4 BUFX4_449 ( .A(u1__abc_73140_new_n906_), .Y(u1__abc_73140_new_n906__bF_buf0));
BUFX4 BUFX4_45 ( .A(u0__abc_76628_new_n2719_), .Y(u0__abc_76628_new_n2719__bF_buf4));
BUFX4 BUFX4_450 ( .A(u0_u0__abc_72207_new_n361_), .Y(u0_u0__abc_72207_new_n361__bF_buf4));
BUFX4 BUFX4_451 ( .A(u0_u0__abc_72207_new_n361_), .Y(u0_u0__abc_72207_new_n361__bF_buf3));
BUFX4 BUFX4_452 ( .A(u0_u0__abc_72207_new_n361_), .Y(u0_u0__abc_72207_new_n361__bF_buf2));
BUFX4 BUFX4_453 ( .A(u0_u0__abc_72207_new_n361_), .Y(u0_u0__abc_72207_new_n361__bF_buf1));
BUFX4 BUFX4_454 ( .A(u0_u0__abc_72207_new_n361_), .Y(u0_u0__abc_72207_new_n361__bF_buf0));
BUFX4 BUFX4_455 ( .A(u0__abc_76628_new_n4531_), .Y(u0__abc_76628_new_n4531__bF_buf4));
BUFX4 BUFX4_456 ( .A(u0__abc_76628_new_n4531_), .Y(u0__abc_76628_new_n4531__bF_buf3));
BUFX4 BUFX4_457 ( .A(u0__abc_76628_new_n4531_), .Y(u0__abc_76628_new_n4531__bF_buf2));
BUFX4 BUFX4_458 ( .A(u0__abc_76628_new_n4531_), .Y(u0__abc_76628_new_n4531__bF_buf1));
BUFX4 BUFX4_459 ( .A(u0__abc_76628_new_n4531_), .Y(u0__abc_76628_new_n4531__bF_buf0));
BUFX4 BUFX4_46 ( .A(u0__abc_76628_new_n2719_), .Y(u0__abc_76628_new_n2719__bF_buf3));
BUFX4 BUFX4_460 ( .A(u5__abc_81276_new_n1682_), .Y(u5__abc_81276_new_n1682__bF_buf4));
BUFX4 BUFX4_461 ( .A(u5__abc_81276_new_n1682_), .Y(u5__abc_81276_new_n1682__bF_buf3));
BUFX4 BUFX4_462 ( .A(u5__abc_81276_new_n1682_), .Y(u5__abc_81276_new_n1682__bF_buf2));
BUFX4 BUFX4_463 ( .A(u5__abc_81276_new_n1682_), .Y(u5__abc_81276_new_n1682__bF_buf1));
BUFX4 BUFX4_464 ( .A(u5__abc_81276_new_n1682_), .Y(u5__abc_81276_new_n1682__bF_buf0));
BUFX4 BUFX4_465 ( .A(u5__abc_81276_new_n522_), .Y(u5__abc_81276_new_n522__bF_buf4));
BUFX4 BUFX4_466 ( .A(u5__abc_81276_new_n522_), .Y(u5__abc_81276_new_n522__bF_buf3));
BUFX4 BUFX4_467 ( .A(u5__abc_81276_new_n522_), .Y(u5__abc_81276_new_n522__bF_buf2));
BUFX4 BUFX4_468 ( .A(u5__abc_81276_new_n522_), .Y(u5__abc_81276_new_n522__bF_buf1));
BUFX4 BUFX4_469 ( .A(u5__abc_81276_new_n522_), .Y(u5__abc_81276_new_n522__bF_buf0));
BUFX4 BUFX4_47 ( .A(u0__abc_76628_new_n2719_), .Y(u0__abc_76628_new_n2719__bF_buf2));
BUFX4 BUFX4_470 ( .A(u0__abc_76628_new_n1177_), .Y(u0__abc_76628_new_n1177__bF_buf5));
BUFX4 BUFX4_471 ( .A(u0__abc_76628_new_n1177_), .Y(u0__abc_76628_new_n1177__bF_buf4));
BUFX4 BUFX4_472 ( .A(u0__abc_76628_new_n1177_), .Y(u0__abc_76628_new_n1177__bF_buf3));
BUFX4 BUFX4_473 ( .A(u0__abc_76628_new_n1177_), .Y(u0__abc_76628_new_n1177__bF_buf2));
BUFX4 BUFX4_474 ( .A(u0__abc_76628_new_n1177_), .Y(u0__abc_76628_new_n1177__bF_buf1));
BUFX4 BUFX4_475 ( .A(u0__abc_76628_new_n1177_), .Y(u0__abc_76628_new_n1177__bF_buf0));
BUFX4 BUFX4_476 ( .A(u0__abc_76628_new_n4528_), .Y(u0__abc_76628_new_n4528__bF_buf4));
BUFX4 BUFX4_477 ( .A(u0__abc_76628_new_n4528_), .Y(u0__abc_76628_new_n4528__bF_buf3));
BUFX4 BUFX4_478 ( .A(u0__abc_76628_new_n4528_), .Y(u0__abc_76628_new_n4528__bF_buf2));
BUFX4 BUFX4_479 ( .A(u0__abc_76628_new_n4528_), .Y(u0__abc_76628_new_n4528__bF_buf1));
BUFX4 BUFX4_48 ( .A(u0__abc_76628_new_n2719_), .Y(u0__abc_76628_new_n2719__bF_buf1));
BUFX4 BUFX4_480 ( .A(u0__abc_76628_new_n4528_), .Y(u0__abc_76628_new_n4528__bF_buf0));
BUFX4 BUFX4_481 ( .A(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562), .Y(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf3));
BUFX4 BUFX4_482 ( .A(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562), .Y(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf2));
BUFX4 BUFX4_483 ( .A(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562), .Y(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf1));
BUFX4 BUFX4_484 ( .A(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562), .Y(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf0));
BUFX4 BUFX4_485 ( .A(u0__abc_76628_new_n4566_), .Y(u0__abc_76628_new_n4566__bF_buf4));
BUFX4 BUFX4_486 ( .A(u0__abc_76628_new_n4566_), .Y(u0__abc_76628_new_n4566__bF_buf3));
BUFX4 BUFX4_487 ( .A(u0__abc_76628_new_n4566_), .Y(u0__abc_76628_new_n4566__bF_buf2));
BUFX4 BUFX4_488 ( .A(u0__abc_76628_new_n4566_), .Y(u0__abc_76628_new_n4566__bF_buf1));
BUFX4 BUFX4_489 ( .A(u0__abc_76628_new_n4566_), .Y(u0__abc_76628_new_n4566__bF_buf0));
BUFX4 BUFX4_49 ( .A(u0__abc_76628_new_n2719_), .Y(u0__abc_76628_new_n2719__bF_buf0));
BUFX4 BUFX4_490 ( .A(u5_cmd_asserted), .Y(u5_cmd_asserted_bF_buf3));
BUFX4 BUFX4_491 ( .A(u5_cmd_asserted), .Y(u5_cmd_asserted_bF_buf1));
BUFX4 BUFX4_492 ( .A(u5_cmd_asserted), .Y(u5_cmd_asserted_bF_buf0));
BUFX4 BUFX4_493 ( .A(u3__abc_74070_new_n449_), .Y(u3__abc_74070_new_n449__bF_buf3));
BUFX4 BUFX4_494 ( .A(u3__abc_74070_new_n449_), .Y(u3__abc_74070_new_n449__bF_buf2));
BUFX4 BUFX4_495 ( .A(u1__abc_73140_new_n268_), .Y(u1__abc_73140_new_n268__bF_buf4));
BUFX4 BUFX4_496 ( .A(u1__abc_73140_new_n900_), .Y(u1__abc_73140_new_n900__bF_buf4));
BUFX4 BUFX4_497 ( .A(u1__abc_73140_new_n900_), .Y(u1__abc_73140_new_n900__bF_buf3));
BUFX4 BUFX4_498 ( .A(u1__abc_73140_new_n900_), .Y(u1__abc_73140_new_n900__bF_buf2));
BUFX4 BUFX4_499 ( .A(u1__abc_73140_new_n900_), .Y(u1__abc_73140_new_n900__bF_buf1));
BUFX4 BUFX4_5 ( .A(clk_i), .Y(clk_i_hier0_bF_buf4));
BUFX4 BUFX4_50 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf3_));
BUFX4 BUFX4_500 ( .A(u1__abc_73140_new_n900_), .Y(u1__abc_73140_new_n900__bF_buf0));
BUFX4 BUFX4_501 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf3_));
BUFX4 BUFX4_502 ( .A(row_adr_8_), .Y(row_adr_8_bF_buf2_));
BUFX4 BUFX4_503 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf3_));
BUFX4 BUFX4_504 ( .A(row_adr_11_), .Y(row_adr_11_bF_buf2_));
BUFX4 BUFX4_505 ( .A(u0__abc_76628_new_n1174_), .Y(u0__abc_76628_new_n1174__bF_buf5));
BUFX4 BUFX4_506 ( .A(u0__abc_76628_new_n1174_), .Y(u0__abc_76628_new_n1174__bF_buf4));
BUFX4 BUFX4_507 ( .A(u0__abc_76628_new_n1174_), .Y(u0__abc_76628_new_n1174__bF_buf3));
BUFX4 BUFX4_508 ( .A(u0__abc_76628_new_n1174_), .Y(u0__abc_76628_new_n1174__bF_buf2));
BUFX4 BUFX4_509 ( .A(u0__abc_76628_new_n1174_), .Y(u0__abc_76628_new_n1174__bF_buf1));
BUFX4 BUFX4_51 ( .A(row_adr_4_), .Y(row_adr_4_bF_buf2_));
BUFX4 BUFX4_510 ( .A(u0__abc_76628_new_n1174_), .Y(u0__abc_76628_new_n1174__bF_buf0));
BUFX4 BUFX4_511 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf3_));
BUFX4 BUFX4_512 ( .A(row_adr_5_), .Y(row_adr_5_bF_buf2_));
BUFX4 BUFX4_513 ( .A(u0_u0_rst_r2), .Y(u0_u0_rst_r2_bF_buf5));
BUFX4 BUFX4_514 ( .A(u0_u0_rst_r2), .Y(u0_u0_rst_r2_bF_buf4));
BUFX4 BUFX4_515 ( .A(u0_u0_rst_r2), .Y(u0_u0_rst_r2_bF_buf3));
BUFX4 BUFX4_516 ( .A(u0_u0_rst_r2), .Y(u0_u0_rst_r2_bF_buf2));
BUFX4 BUFX4_517 ( .A(u0_u0_rst_r2), .Y(u0_u0_rst_r2_bF_buf1));
BUFX4 BUFX4_518 ( .A(u0_u0_rst_r2), .Y(u0_u0_rst_r2_bF_buf0));
BUFX4 BUFX4_519 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf5));
BUFX4 BUFX4_52 ( .A(u0__abc_76628_new_n1170_), .Y(u0__abc_76628_new_n1170__bF_buf6));
BUFX4 BUFX4_520 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf4));
BUFX4 BUFX4_521 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf3));
BUFX4 BUFX4_522 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf2));
BUFX4 BUFX4_523 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf1));
BUFX4 BUFX4_524 ( .A(wb_stb_i), .Y(wb_stb_i_bF_buf0));
BUFX4 BUFX4_525 ( .A(u0__abc_76628_new_n2720_), .Y(u0__abc_76628_new_n2720__bF_buf5));
BUFX4 BUFX4_526 ( .A(u0__abc_76628_new_n2720_), .Y(u0__abc_76628_new_n2720__bF_buf4));
BUFX4 BUFX4_527 ( .A(u0__abc_76628_new_n2720_), .Y(u0__abc_76628_new_n2720__bF_buf3));
BUFX4 BUFX4_528 ( .A(u0__abc_76628_new_n2720_), .Y(u0__abc_76628_new_n2720__bF_buf2));
BUFX4 BUFX4_529 ( .A(u0__abc_76628_new_n2720_), .Y(u0__abc_76628_new_n2720__bF_buf1));
BUFX4 BUFX4_53 ( .A(u0__abc_76628_new_n1170_), .Y(u0__abc_76628_new_n1170__bF_buf5));
BUFX4 BUFX4_530 ( .A(u0__abc_76628_new_n2720_), .Y(u0__abc_76628_new_n2720__bF_buf0));
BUFX4 BUFX4_531 ( .A(u5__abc_81276_new_n416_), .Y(u5__abc_81276_new_n416__bF_buf3));
BUFX4 BUFX4_532 ( .A(u5__abc_81276_new_n416_), .Y(u5__abc_81276_new_n416__bF_buf2));
BUFX4 BUFX4_533 ( .A(u0__abc_76628_new_n2717_), .Y(u0__abc_76628_new_n2717__bF_buf5));
BUFX4 BUFX4_534 ( .A(u0__abc_76628_new_n2717_), .Y(u0__abc_76628_new_n2717__bF_buf4));
BUFX4 BUFX4_535 ( .A(u0__abc_76628_new_n2717_), .Y(u0__abc_76628_new_n2717__bF_buf3));
BUFX4 BUFX4_536 ( .A(u0__abc_76628_new_n2717_), .Y(u0__abc_76628_new_n2717__bF_buf2));
BUFX4 BUFX4_537 ( .A(u0__abc_76628_new_n2717_), .Y(u0__abc_76628_new_n2717__bF_buf1));
BUFX4 BUFX4_538 ( .A(u0__abc_76628_new_n2717_), .Y(u0__abc_76628_new_n2717__bF_buf0));
BUFX4 BUFX4_539 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf3_));
BUFX4 BUFX4_54 ( .A(u0__abc_76628_new_n1170_), .Y(u0__abc_76628_new_n1170__bF_buf4));
BUFX4 BUFX4_540 ( .A(row_adr_2_), .Y(row_adr_2_bF_buf2_));
BUFX4 BUFX4_541 ( .A(u0__abc_76628_new_n4554_), .Y(u0__abc_76628_new_n4554__bF_buf4));
BUFX4 BUFX4_542 ( .A(u0__abc_76628_new_n4554_), .Y(u0__abc_76628_new_n4554__bF_buf3));
BUFX4 BUFX4_543 ( .A(u0__abc_76628_new_n4554_), .Y(u0__abc_76628_new_n4554__bF_buf2));
BUFX4 BUFX4_544 ( .A(u0__abc_76628_new_n4554_), .Y(u0__abc_76628_new_n4554__bF_buf1));
BUFX4 BUFX4_545 ( .A(u0__abc_76628_new_n4554_), .Y(u0__abc_76628_new_n4554__bF_buf0));
BUFX4 BUFX4_546 ( .A(u5__abc_81276_new_n448_), .Y(u5__abc_81276_new_n448__bF_buf5));
BUFX4 BUFX4_547 ( .A(u5__abc_81276_new_n448_), .Y(u5__abc_81276_new_n448__bF_buf4));
BUFX4 BUFX4_548 ( .A(u5__abc_81276_new_n448_), .Y(u5__abc_81276_new_n448__bF_buf3));
BUFX4 BUFX4_549 ( .A(u5__abc_81276_new_n448_), .Y(u5__abc_81276_new_n448__bF_buf2));
BUFX4 BUFX4_55 ( .A(u0__abc_76628_new_n1170_), .Y(u0__abc_76628_new_n1170__bF_buf3));
BUFX4 BUFX4_550 ( .A(u5__abc_81276_new_n448_), .Y(u5__abc_81276_new_n448__bF_buf1));
BUFX4 BUFX4_551 ( .A(u5__abc_81276_new_n448_), .Y(u5__abc_81276_new_n448__bF_buf0));
BUFX4 BUFX4_552 ( .A(_abc_85006_new_n240_), .Y(_abc_85006_new_n240__bF_buf5));
BUFX4 BUFX4_553 ( .A(_abc_85006_new_n240_), .Y(_abc_85006_new_n240__bF_buf4));
BUFX4 BUFX4_554 ( .A(_abc_85006_new_n240_), .Y(_abc_85006_new_n240__bF_buf3));
BUFX4 BUFX4_555 ( .A(_abc_85006_new_n240_), .Y(_abc_85006_new_n240__bF_buf2));
BUFX4 BUFX4_556 ( .A(_abc_85006_new_n240_), .Y(_abc_85006_new_n240__bF_buf1));
BUFX4 BUFX4_557 ( .A(_abc_85006_new_n240_), .Y(_abc_85006_new_n240__bF_buf0));
BUFX4 BUFX4_558 ( .A(u0__abc_76628_new_n1197_), .Y(u0__abc_76628_new_n1197__bF_buf5));
BUFX4 BUFX4_559 ( .A(u0__abc_76628_new_n1197_), .Y(u0__abc_76628_new_n1197__bF_buf4));
BUFX4 BUFX4_56 ( .A(u0__abc_76628_new_n1170_), .Y(u0__abc_76628_new_n1170__bF_buf2));
BUFX4 BUFX4_560 ( .A(u0__abc_76628_new_n1197_), .Y(u0__abc_76628_new_n1197__bF_buf3));
BUFX4 BUFX4_561 ( .A(u0__abc_76628_new_n1197_), .Y(u0__abc_76628_new_n1197__bF_buf2));
BUFX4 BUFX4_562 ( .A(u0__abc_76628_new_n1197_), .Y(u0__abc_76628_new_n1197__bF_buf1));
BUFX4 BUFX4_563 ( .A(u0__abc_76628_new_n1197_), .Y(u0__abc_76628_new_n1197__bF_buf0));
BUFX4 BUFX4_564 ( .A(u1__abc_73140_new_n826_), .Y(u1__abc_73140_new_n826__bF_buf3));
BUFX4 BUFX4_565 ( .A(u1__abc_73140_new_n826_), .Y(u1__abc_73140_new_n826__bF_buf2));
BUFX4 BUFX4_566 ( .A(u1__abc_73140_new_n826_), .Y(u1__abc_73140_new_n826__bF_buf1));
BUFX4 BUFX4_567 ( .A(u1__abc_73140_new_n826_), .Y(u1__abc_73140_new_n826__bF_buf0));
BUFX4 BUFX4_568 ( .A(u3__abc_74070_new_n625_), .Y(u3__abc_74070_new_n625__bF_buf4));
BUFX4 BUFX4_569 ( .A(u3__abc_74070_new_n625_), .Y(u3__abc_74070_new_n625__bF_buf3));
BUFX4 BUFX4_57 ( .A(u0__abc_76628_new_n1170_), .Y(u0__abc_76628_new_n1170__bF_buf1));
BUFX4 BUFX4_570 ( .A(u3__abc_74070_new_n625_), .Y(u3__abc_74070_new_n625__bF_buf2));
BUFX4 BUFX4_571 ( .A(u3__abc_74070_new_n625_), .Y(u3__abc_74070_new_n625__bF_buf1));
BUFX4 BUFX4_572 ( .A(u3__abc_74070_new_n625_), .Y(u3__abc_74070_new_n625__bF_buf0));
BUFX4 BUFX4_573 ( .A(u0__abc_76628_new_n4298_), .Y(u0__abc_76628_new_n4298__bF_buf4));
BUFX4 BUFX4_574 ( .A(u0__abc_76628_new_n4298_), .Y(u0__abc_76628_new_n4298__bF_buf3));
BUFX4 BUFX4_575 ( .A(u0__abc_76628_new_n4298_), .Y(u0__abc_76628_new_n4298__bF_buf2));
BUFX4 BUFX4_576 ( .A(u0__abc_76628_new_n4298_), .Y(u0__abc_76628_new_n4298__bF_buf1));
BUFX4 BUFX4_577 ( .A(u0__abc_76628_new_n4298_), .Y(u0__abc_76628_new_n4298__bF_buf0));
BUFX4 BUFX4_578 ( .A(u0__abc_76628_new_n4510_), .Y(u0__abc_76628_new_n4510__bF_buf4));
BUFX4 BUFX4_579 ( .A(u0__abc_76628_new_n4510_), .Y(u0__abc_76628_new_n4510__bF_buf3));
BUFX4 BUFX4_58 ( .A(u0__abc_76628_new_n1170_), .Y(u0__abc_76628_new_n1170__bF_buf0));
BUFX4 BUFX4_580 ( .A(u0__abc_76628_new_n4510_), .Y(u0__abc_76628_new_n4510__bF_buf2));
BUFX4 BUFX4_581 ( .A(u0__abc_76628_new_n4510_), .Y(u0__abc_76628_new_n4510__bF_buf1));
BUFX4 BUFX4_582 ( .A(u0__abc_76628_new_n4510_), .Y(u0__abc_76628_new_n4510__bF_buf0));
BUFX4 BUFX4_583 ( .A(u5__abc_81276_new_n1526_), .Y(u5__abc_81276_new_n1526__bF_buf3));
BUFX4 BUFX4_584 ( .A(u5__abc_81276_new_n1526_), .Y(u5__abc_81276_new_n1526__bF_buf2));
BUFX4 BUFX4_585 ( .A(u5__abc_81276_new_n1526_), .Y(u5__abc_81276_new_n1526__bF_buf1));
BUFX4 BUFX4_586 ( .A(u5__abc_81276_new_n1526_), .Y(u5__abc_81276_new_n1526__bF_buf0));
BUFX4 BUFX4_587 ( .A(u0__abc_76628_new_n4507_), .Y(u0__abc_76628_new_n4507__bF_buf4));
BUFX4 BUFX4_588 ( .A(u0__abc_76628_new_n4507_), .Y(u0__abc_76628_new_n4507__bF_buf3));
BUFX4 BUFX4_589 ( .A(u0__abc_76628_new_n4507_), .Y(u0__abc_76628_new_n4507__bF_buf2));
BUFX4 BUFX4_59 ( .A(u6__abc_85257_new_n155_), .Y(u6__abc_85257_new_n155__bF_buf4));
BUFX4 BUFX4_590 ( .A(u0__abc_76628_new_n4507_), .Y(u0__abc_76628_new_n4507__bF_buf1));
BUFX4 BUFX4_591 ( .A(u0__abc_76628_new_n4507_), .Y(u0__abc_76628_new_n4507__bF_buf0));
BUFX4 BUFX4_592 ( .A(u3_u0__abc_75526_new_n1052_), .Y(u3_u0__abc_75526_new_n1052__bF_buf5));
BUFX4 BUFX4_593 ( .A(u3_u0__abc_75526_new_n1052_), .Y(u3_u0__abc_75526_new_n1052__bF_buf4));
BUFX4 BUFX4_594 ( .A(u3_u0__abc_75526_new_n1052_), .Y(u3_u0__abc_75526_new_n1052__bF_buf3));
BUFX4 BUFX4_595 ( .A(u3_u0__abc_75526_new_n1052_), .Y(u3_u0__abc_75526_new_n1052__bF_buf2));
BUFX4 BUFX4_596 ( .A(u3_u0__abc_75526_new_n1052_), .Y(u3_u0__abc_75526_new_n1052__bF_buf1));
BUFX4 BUFX4_597 ( .A(u3_u0__abc_75526_new_n1052_), .Y(u3_u0__abc_75526_new_n1052__bF_buf0));
BUFX4 BUFX4_598 ( .A(u0__abc_76628_new_n4545_), .Y(u0__abc_76628_new_n4545__bF_buf4));
BUFX4 BUFX4_599 ( .A(u0__abc_76628_new_n4545_), .Y(u0__abc_76628_new_n4545__bF_buf3));
BUFX4 BUFX4_6 ( .A(clk_i), .Y(clk_i_hier0_bF_buf3));
BUFX4 BUFX4_60 ( .A(u6__abc_85257_new_n155_), .Y(u6__abc_85257_new_n155__bF_buf3));
BUFX4 BUFX4_600 ( .A(u0__abc_76628_new_n4545_), .Y(u0__abc_76628_new_n4545__bF_buf2));
BUFX4 BUFX4_601 ( .A(u0__abc_76628_new_n4545_), .Y(u0__abc_76628_new_n4545__bF_buf1));
BUFX4 BUFX4_602 ( .A(u0__abc_76628_new_n4545_), .Y(u0__abc_76628_new_n4545__bF_buf0));
BUFX4 BUFX4_603 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf5_));
BUFX4 BUFX4_604 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf4_));
BUFX4 BUFX4_605 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf3_));
BUFX4 BUFX4_606 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf2_));
BUFX4 BUFX4_607 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf1_));
BUFX4 BUFX4_608 ( .A(spec_req_cs_6_), .Y(spec_req_cs_6_bF_buf0_));
BUFX4 BUFX4_609 ( .A(u5__abc_81276_new_n480_), .Y(u5__abc_81276_new_n480__bF_buf4));
BUFX4 BUFX4_61 ( .A(u6__abc_85257_new_n155_), .Y(u6__abc_85257_new_n155__bF_buf2));
BUFX4 BUFX4_610 ( .A(u5__abc_81276_new_n480_), .Y(u5__abc_81276_new_n480__bF_buf3));
BUFX4 BUFX4_611 ( .A(u5__abc_81276_new_n480_), .Y(u5__abc_81276_new_n480__bF_buf2));
BUFX4 BUFX4_612 ( .A(u5__abc_81276_new_n480_), .Y(u5__abc_81276_new_n480__bF_buf1));
BUFX4 BUFX4_613 ( .A(u5__abc_81276_new_n480_), .Y(u5__abc_81276_new_n480__bF_buf0));
BUFX4 BUFX4_614 ( .A(u3_u0__abc_75526_new_n1049_), .Y(u3_u0__abc_75526_new_n1049__bF_buf5));
BUFX4 BUFX4_615 ( .A(u3_u0__abc_75526_new_n1049_), .Y(u3_u0__abc_75526_new_n1049__bF_buf4));
BUFX4 BUFX4_616 ( .A(u3_u0__abc_75526_new_n1049_), .Y(u3_u0__abc_75526_new_n1049__bF_buf3));
BUFX4 BUFX4_617 ( .A(u3_u0__abc_75526_new_n1049_), .Y(u3_u0__abc_75526_new_n1049__bF_buf2));
BUFX4 BUFX4_618 ( .A(u3_u0__abc_75526_new_n1049_), .Y(u3_u0__abc_75526_new_n1049__bF_buf1));
BUFX4 BUFX4_619 ( .A(u3_u0__abc_75526_new_n1049_), .Y(u3_u0__abc_75526_new_n1049__bF_buf0));
BUFX4 BUFX4_62 ( .A(u6__abc_85257_new_n155_), .Y(u6__abc_85257_new_n155__bF_buf1));
BUFX4 BUFX4_620 ( .A(u3__abc_74070_new_n275_), .Y(u3__abc_74070_new_n275__bF_buf4));
BUFX4 BUFX4_621 ( .A(u3__abc_74070_new_n275_), .Y(u3__abc_74070_new_n275__bF_buf3));
BUFX4 BUFX4_622 ( .A(u3__abc_74070_new_n275_), .Y(u3__abc_74070_new_n275__bF_buf2));
BUFX4 BUFX4_623 ( .A(u3__abc_74070_new_n275_), .Y(u3__abc_74070_new_n275__bF_buf1));
BUFX4 BUFX4_624 ( .A(u3__abc_74070_new_n275_), .Y(u3__abc_74070_new_n275__bF_buf0));
BUFX4 BUFX4_625 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf5_));
BUFX4 BUFX4_626 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf4_));
BUFX4 BUFX4_627 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf3_));
BUFX4 BUFX4_628 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf2_));
BUFX4 BUFX4_629 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf1_));
BUFX4 BUFX4_63 ( .A(u6__abc_85257_new_n155_), .Y(u6__abc_85257_new_n155__bF_buf0));
BUFX4 BUFX4_630 ( .A(spec_req_cs_3_), .Y(spec_req_cs_3_bF_buf0_));
BUFX4 BUFX4_631 ( .A(u1__abc_73140_new_n570_), .Y(u1__abc_73140_new_n570__bF_buf3));
BUFX4 BUFX4_632 ( .A(u1__abc_73140_new_n570_), .Y(u1__abc_73140_new_n570__bF_buf2));
BUFX4 BUFX4_633 ( .A(u1__abc_73140_new_n570_), .Y(u1__abc_73140_new_n570__bF_buf1));
BUFX4 BUFX4_634 ( .A(u1__abc_73140_new_n570_), .Y(u1__abc_73140_new_n570__bF_buf0));
BUFX4 BUFX4_635 ( .A(u0_rst_r3), .Y(u0_rst_r3_bF_buf4));
BUFX4 BUFX4_636 ( .A(u0_rst_r3), .Y(u0_rst_r3_bF_buf3));
BUFX4 BUFX4_637 ( .A(u0_rst_r3), .Y(u0_rst_r3_bF_buf2));
BUFX4 BUFX4_638 ( .A(u0_rst_r3), .Y(u0_rst_r3_bF_buf1));
BUFX4 BUFX4_639 ( .A(u0_rst_r3), .Y(u0_rst_r3_bF_buf0));
BUFX4 BUFX4_64 ( .A(u0__abc_76628_new_n4556_), .Y(u0__abc_76628_new_n4556__bF_buf4));
BUFX4 BUFX4_640 ( .A(u1__abc_73140_new_n567_), .Y(u1__abc_73140_new_n567__bF_buf3));
BUFX4 BUFX4_641 ( .A(u1__abc_73140_new_n567_), .Y(u1__abc_73140_new_n567__bF_buf2));
BUFX4 BUFX4_642 ( .A(u1__abc_73140_new_n567_), .Y(u1__abc_73140_new_n567__bF_buf1));
BUFX4 BUFX4_643 ( .A(u1__abc_73140_new_n567_), .Y(u1__abc_73140_new_n567__bF_buf0));
BUFX4 BUFX4_644 ( .A(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9));
BUFX4 BUFX4_645 ( .A(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8));
BUFX4 BUFX4_646 ( .A(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7));
BUFX4 BUFX4_647 ( .A(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6));
BUFX4 BUFX4_648 ( .A(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5));
BUFX4 BUFX4_649 ( .A(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4));
BUFX4 BUFX4_65 ( .A(u0__abc_76628_new_n4556_), .Y(u0__abc_76628_new_n4556__bF_buf3));
BUFX4 BUFX4_650 ( .A(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3));
BUFX4 BUFX4_651 ( .A(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2));
BUFX4 BUFX4_652 ( .A(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1));
BUFX4 BUFX4_653 ( .A(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0));
BUFX4 BUFX4_654 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf5_));
BUFX4 BUFX4_655 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf4_));
BUFX4 BUFX4_656 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf3_));
BUFX4 BUFX4_657 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf2_));
BUFX4 BUFX4_658 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf1_));
BUFX4 BUFX4_659 ( .A(spec_req_cs_0_), .Y(spec_req_cs_0_bF_buf0_));
BUFX4 BUFX4_66 ( .A(u0__abc_76628_new_n4556_), .Y(u0__abc_76628_new_n4556__bF_buf2));
BUFX4 BUFX4_660 ( .A(u3_u0__abc_75526_new_n1043_), .Y(u3_u0__abc_75526_new_n1043__bF_buf5));
BUFX4 BUFX4_661 ( .A(u3_u0__abc_75526_new_n1043_), .Y(u3_u0__abc_75526_new_n1043__bF_buf4));
BUFX4 BUFX4_662 ( .A(u3_u0__abc_75526_new_n1043_), .Y(u3_u0__abc_75526_new_n1043__bF_buf3));
BUFX4 BUFX4_663 ( .A(u3_u0__abc_75526_new_n1043_), .Y(u3_u0__abc_75526_new_n1043__bF_buf2));
BUFX4 BUFX4_664 ( .A(u3_u0__abc_75526_new_n1043_), .Y(u3_u0__abc_75526_new_n1043__bF_buf1));
BUFX4 BUFX4_665 ( .A(u3_u0__abc_75526_new_n1043_), .Y(u3_u0__abc_75526_new_n1043__bF_buf0));
BUFX4 BUFX4_666 ( .A(u0_u0__0lmr_req_we_0_0_), .Y(u0_u0__0lmr_req_we_0_0_bF_buf4_));
BUFX4 BUFX4_667 ( .A(u0_u0__0lmr_req_we_0_0_), .Y(u0_u0__0lmr_req_we_0_0_bF_buf3_));
BUFX4 BUFX4_668 ( .A(u0_u0__0lmr_req_we_0_0_), .Y(u0_u0__0lmr_req_we_0_0_bF_buf2_));
BUFX4 BUFX4_669 ( .A(u0_u0__0lmr_req_we_0_0_), .Y(u0_u0__0lmr_req_we_0_0_bF_buf1_));
BUFX4 BUFX4_67 ( .A(u0__abc_76628_new_n4556_), .Y(u0__abc_76628_new_n4556__bF_buf1));
BUFX4 BUFX4_670 ( .A(u0_u0__0lmr_req_we_0_0_), .Y(u0_u0__0lmr_req_we_0_0_bF_buf0_));
BUFX4 BUFX4_671 ( .A(u0__abc_76628_new_n1946_), .Y(u0__abc_76628_new_n1946__bF_buf3));
BUFX4 BUFX4_672 ( .A(u0_u1__0init_req_we_0_0_), .Y(u0_u1__0init_req_we_0_0_bF_buf7_));
BUFX4 BUFX4_673 ( .A(u0_u1__0init_req_we_0_0_), .Y(u0_u1__0init_req_we_0_0_bF_buf6_));
BUFX4 BUFX4_674 ( .A(u0_u1__0init_req_we_0_0_), .Y(u0_u1__0init_req_we_0_0_bF_buf5_));
BUFX4 BUFX4_675 ( .A(u0_u1__0init_req_we_0_0_), .Y(u0_u1__0init_req_we_0_0_bF_buf4_));
BUFX4 BUFX4_676 ( .A(u0_u1__0init_req_we_0_0_), .Y(u0_u1__0init_req_we_0_0_bF_buf3_));
BUFX4 BUFX4_677 ( .A(u0_u1__0init_req_we_0_0_), .Y(u0_u1__0init_req_we_0_0_bF_buf2_));
BUFX4 BUFX4_678 ( .A(u0_u1__0init_req_we_0_0_), .Y(u0_u1__0init_req_we_0_0_bF_buf1_));
BUFX4 BUFX4_679 ( .A(u0_u1__0init_req_we_0_0_), .Y(u0_u1__0init_req_we_0_0_bF_buf0_));
BUFX4 BUFX4_68 ( .A(u0__abc_76628_new_n4556_), .Y(u0__abc_76628_new_n4556__bF_buf0));
BUFX4 BUFX4_680 ( .A(u1_bas), .Y(u1_bas_bF_buf3));
BUFX4 BUFX4_681 ( .A(u1_bas), .Y(u1_bas_bF_buf2));
BUFX4 BUFX4_682 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10));
BUFX4 BUFX4_683 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9));
BUFX4 BUFX4_684 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8));
BUFX4 BUFX4_685 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7));
BUFX4 BUFX4_686 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6));
BUFX4 BUFX4_687 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5));
BUFX4 BUFX4_688 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4));
BUFX4 BUFX4_689 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3));
BUFX4 BUFX4_69 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf3_));
BUFX4 BUFX4_690 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2));
BUFX4 BUFX4_691 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1));
BUFX4 BUFX4_692 ( .A(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0));
BUFX4 BUFX4_693 ( .A(u0__abc_76628_new_n1179_), .Y(u0__abc_76628_new_n1179__bF_buf5));
BUFX4 BUFX4_694 ( .A(u0__abc_76628_new_n1179_), .Y(u0__abc_76628_new_n1179__bF_buf4));
BUFX4 BUFX4_695 ( .A(u0__abc_76628_new_n1179_), .Y(u0__abc_76628_new_n1179__bF_buf3));
BUFX4 BUFX4_696 ( .A(u0__abc_76628_new_n1179_), .Y(u0__abc_76628_new_n1179__bF_buf2));
BUFX4 BUFX4_697 ( .A(u0__abc_76628_new_n1179_), .Y(u0__abc_76628_new_n1179__bF_buf1));
BUFX4 BUFX4_698 ( .A(u0__abc_76628_new_n1179_), .Y(u0__abc_76628_new_n1179__bF_buf0));
BUFX4 BUFX4_699 ( .A(u1__abc_73140_new_n561_), .Y(u1__abc_73140_new_n561__bF_buf4));
BUFX4 BUFX4_7 ( .A(clk_i), .Y(clk_i_hier0_bF_buf2));
BUFX4 BUFX4_70 ( .A(row_adr_1_), .Y(row_adr_1_bF_buf2_));
BUFX4 BUFX4_700 ( .A(u1__abc_73140_new_n561_), .Y(u1__abc_73140_new_n561__bF_buf3));
BUFX4 BUFX4_701 ( .A(u1__abc_73140_new_n561_), .Y(u1__abc_73140_new_n561__bF_buf2));
BUFX4 BUFX4_702 ( .A(u1__abc_73140_new_n561_), .Y(u1__abc_73140_new_n561__bF_buf1));
BUFX4 BUFX4_703 ( .A(u1__abc_73140_new_n561_), .Y(u1__abc_73140_new_n561__bF_buf0));
BUFX4 BUFX4_704 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf10));
BUFX4 BUFX4_705 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf9));
BUFX4 BUFX4_706 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf8));
BUFX4 BUFX4_707 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf7));
BUFX4 BUFX4_708 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf6));
BUFX4 BUFX4_709 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf5));
BUFX4 BUFX4_71 ( .A(u0_u0__0init_req_we_0_0_), .Y(u0_u0__0init_req_we_0_0_bF_buf4_));
BUFX4 BUFX4_710 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf4));
BUFX4 BUFX4_711 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf3));
BUFX4 BUFX4_712 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf2));
BUFX4 BUFX4_713 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf1));
BUFX4 BUFX4_714 ( .A(mc_clk_i), .Y(mc_clk_i_bF_buf0));
BUFX4 BUFX4_715 ( .A(u5__abc_81276_new_n521_), .Y(u5__abc_81276_new_n521__bF_buf3));
BUFX4 BUFX4_716 ( .A(u5__abc_81276_new_n521_), .Y(u5__abc_81276_new_n521__bF_buf2));
BUFX4 BUFX4_717 ( .A(u3_u0__abc_75526_new_n1034_), .Y(u3_u0__abc_75526_new_n1034__bF_buf5));
BUFX4 BUFX4_718 ( .A(u3_u0__abc_75526_new_n1034_), .Y(u3_u0__abc_75526_new_n1034__bF_buf4));
BUFX4 BUFX4_719 ( .A(u3_u0__abc_75526_new_n1034_), .Y(u3_u0__abc_75526_new_n1034__bF_buf3));
BUFX4 BUFX4_72 ( .A(u0_u0__0init_req_we_0_0_), .Y(u0_u0__0init_req_we_0_0_bF_buf3_));
BUFX4 BUFX4_720 ( .A(u3_u0__abc_75526_new_n1034_), .Y(u3_u0__abc_75526_new_n1034__bF_buf2));
BUFX4 BUFX4_721 ( .A(u3_u0__abc_75526_new_n1034_), .Y(u3_u0__abc_75526_new_n1034__bF_buf1));
BUFX4 BUFX4_722 ( .A(u3_u0__abc_75526_new_n1034_), .Y(u3_u0__abc_75526_new_n1034__bF_buf0));
BUFX4 BUFX4_73 ( .A(u0_u0__0init_req_we_0_0_), .Y(u0_u0__0init_req_we_0_0_bF_buf2_));
BUFX4 BUFX4_74 ( .A(u0_u0__0init_req_we_0_0_), .Y(u0_u0__0init_req_we_0_0_bF_buf1_));
BUFX4 BUFX4_75 ( .A(u0_u0__0init_req_we_0_0_), .Y(u0_u0__0init_req_we_0_0_bF_buf0_));
BUFX4 BUFX4_76 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf96));
BUFX4 BUFX4_77 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf95));
BUFX4 BUFX4_78 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf94));
BUFX4 BUFX4_79 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf93));
BUFX4 BUFX4_8 ( .A(clk_i), .Y(clk_i_hier0_bF_buf1));
BUFX4 BUFX4_80 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf92));
BUFX4 BUFX4_81 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf91));
BUFX4 BUFX4_82 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf90));
BUFX4 BUFX4_83 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf89));
BUFX4 BUFX4_84 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf88));
BUFX4 BUFX4_85 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf87));
BUFX4 BUFX4_86 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf86));
BUFX4 BUFX4_87 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf85));
BUFX4 BUFX4_88 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf84));
BUFX4 BUFX4_89 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf83));
BUFX4 BUFX4_9 ( .A(clk_i), .Y(clk_i_hier0_bF_buf0));
BUFX4 BUFX4_90 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf82));
BUFX4 BUFX4_91 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf81));
BUFX4 BUFX4_92 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf80));
BUFX4 BUFX4_93 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf79));
BUFX4 BUFX4_94 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf78));
BUFX4 BUFX4_95 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf77));
BUFX4 BUFX4_96 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf76));
BUFX4 BUFX4_97 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf75));
BUFX4 BUFX4_98 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf74));
BUFX4 BUFX4_99 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf73));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_i_bF_buf96), .D(mem_ack), .Q(mem_ack_r));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_i_bF_buf87), .D(u0__0poc_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_85523_6_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_i_bF_buf64), .D(u0_u0__0csc_31_0__26_), .Q(u0_csc0_26_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_i_bF_buf63), .D(u0_u0__0csc_31_0__27_), .Q(u0_csc0_27_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_i_bF_buf62), .D(u0_u0__0csc_31_0__28_), .Q(u0_csc0_28_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_i_bF_buf61), .D(u0_u0__0csc_31_0__29_), .Q(u0_csc0_29_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_i_bF_buf60), .D(u0_u0__0csc_31_0__30_), .Q(u0_csc0_30_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_i_bF_buf59), .D(u0_u0__0csc_31_0__31_), .Q(u0_csc0_31_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_i_bF_buf58), .D(\wb_addr_i[2] ), .Q(u0_u0_addr_r_2_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_i_bF_buf57), .D(\wb_addr_i[3] ), .Q(u0_u0_addr_r_3_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_i_bF_buf56), .D(\wb_addr_i[4] ), .Q(u0_u0_addr_r_4_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_i_bF_buf55), .D(\wb_addr_i[5] ), .Q(u0_u0_addr_r_5_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_i_bF_buf86), .D(u0__0poc_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_85523_7_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_i_bF_buf54), .D(\wb_addr_i[6] ), .Q(u0_u0_addr_r_6_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_i_bF_buf47), .D(u0_u1__0tms_31_0__0_), .Q(u0_tms1_0_));
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_i_bF_buf46), .D(u0_u1__0tms_31_0__1_), .Q(u0_tms1_1_));
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_i_bF_buf45), .D(u0_u1__0tms_31_0__2_), .Q(u0_tms1_2_));
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_i_bF_buf44), .D(u0_u1__0tms_31_0__3_), .Q(u0_tms1_3_));
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_i_bF_buf43), .D(u0_u1__0tms_31_0__4_), .Q(u0_tms1_4_));
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_i_bF_buf42), .D(u0_u1__0tms_31_0__5_), .Q(u0_tms1_5_));
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_i_bF_buf41), .D(u0_u1__0tms_31_0__6_), .Q(u0_tms1_6_));
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_i_bF_buf40), .D(u0_u1__0tms_31_0__7_), .Q(u0_tms1_7_));
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_i_bF_buf39), .D(u0_u1__0tms_31_0__8_), .Q(u0_tms1_8_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_i_bF_buf85), .D(u0__0poc_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_85523_8_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_i_bF_buf38), .D(u0_u1__0tms_31_0__9_), .Q(u0_tms1_9_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_i_bF_buf37), .D(u0_u1__0tms_31_0__10_), .Q(u0_tms1_10_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_i_bF_buf36), .D(u0_u1__0tms_31_0__11_), .Q(u0_tms1_11_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_i_bF_buf35), .D(u0_u1__0tms_31_0__12_), .Q(u0_tms1_12_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_i_bF_buf34), .D(u0_u1__0tms_31_0__13_), .Q(u0_tms1_13_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_i_bF_buf33), .D(u0_u1__0tms_31_0__14_), .Q(u0_tms1_14_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_i_bF_buf32), .D(u0_u1__0tms_31_0__15_), .Q(u0_tms1_15_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_i_bF_buf31), .D(u0_u1__0tms_31_0__16_), .Q(u0_tms1_16_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_i_bF_buf30), .D(u0_u1__0tms_31_0__17_), .Q(u0_tms1_17_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_i_bF_buf29), .D(u0_u1__0tms_31_0__18_), .Q(u0_tms1_18_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_i_bF_buf84), .D(u0__0poc_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_85523_9_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_i_bF_buf28), .D(u0_u1__0tms_31_0__19_), .Q(u0_tms1_19_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_i_bF_buf27), .D(u0_u1__0tms_31_0__20_), .Q(u0_tms1_20_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_i_bF_buf26), .D(u0_u1__0tms_31_0__21_), .Q(u0_tms1_21_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_i_bF_buf25), .D(u0_u1__0tms_31_0__22_), .Q(u0_tms1_22_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_i_bF_buf24), .D(u0_u1__0tms_31_0__23_), .Q(u0_tms1_23_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_i_bF_buf23), .D(u0_u1__0tms_31_0__24_), .Q(u0_tms1_24_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_i_bF_buf22), .D(u0_u1__0tms_31_0__25_), .Q(u0_tms1_25_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_i_bF_buf21), .D(u0_u1__0tms_31_0__26_), .Q(u0_tms1_26_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_i_bF_buf20), .D(u0_u1__0tms_31_0__27_), .Q(u0_tms1_27_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_i_bF_buf19), .D(u0_u1__0tms_31_0__28_), .Q(u0_tms1_28_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_i_bF_buf83), .D(u0__0poc_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_85523_10_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_i_bF_buf18), .D(u0_u1__0tms_31_0__29_), .Q(u0_tms1_29_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_i_bF_buf17), .D(u0_u1__0tms_31_0__30_), .Q(u0_tms1_30_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_i_bF_buf16), .D(u0_u1__0tms_31_0__31_), .Q(u0_tms1_31_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_i_bF_buf15), .D(u0_u1__0csc_31_0__0_), .Q(u0_csc1_0_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_i_bF_buf14), .D(u0_u1__0csc_31_0__1_), .Q(u0_csc1_1_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_i_bF_buf13), .D(u0_u1__0csc_31_0__2_), .Q(u0_csc1_2_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_i_bF_buf12), .D(u0_u1__0csc_31_0__3_), .Q(u0_csc1_3_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_i_bF_buf11), .D(u0_u1__0csc_31_0__4_), .Q(u0_csc1_4_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_i_bF_buf10), .D(u0_u1__0csc_31_0__5_), .Q(u0_csc1_5_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_i_bF_buf9), .D(u0_u1__0csc_31_0__6_), .Q(u0_csc1_6_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_i_bF_buf82), .D(u0__0poc_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_85523_11_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_i_bF_buf8), .D(u0_u1__0csc_31_0__7_), .Q(u0_csc1_7_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_i_bF_buf7), .D(u0_u1__0csc_31_0__8_), .Q(u0_csc1_8_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_i_bF_buf6), .D(u0_u1__0csc_31_0__9_), .Q(u0_csc1_9_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_i_bF_buf5), .D(u0_u1__0csc_31_0__10_), .Q(u0_csc1_10_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_i_bF_buf4), .D(u0_u1__0csc_31_0__11_), .Q(u0_csc1_11_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_i_bF_buf3), .D(u0_u1__0csc_31_0__12_), .Q(u0_csc1_12_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_i_bF_buf2), .D(u0_u1__0csc_31_0__13_), .Q(u0_csc1_13_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_i_bF_buf1), .D(u0_u1__0csc_31_0__14_), .Q(u0_csc1_14_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_i_bF_buf0), .D(u0_u1__0csc_31_0__15_), .Q(u0_csc1_15_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_i_bF_buf96), .D(u0_u1__0csc_31_0__16_), .Q(u0_csc1_16_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_i_bF_buf81), .D(u0__0poc_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_85523_12_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_i_bF_buf95), .D(u0_u1__0csc_31_0__17_), .Q(u0_csc1_17_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_i_bF_buf94), .D(u0_u1__0csc_31_0__18_), .Q(u0_csc1_18_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_i_bF_buf93), .D(u0_u1__0csc_31_0__19_), .Q(u0_csc1_19_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_i_bF_buf92), .D(u0_u1__0csc_31_0__20_), .Q(u0_csc1_20_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_i_bF_buf91), .D(u0_u1__0csc_31_0__21_), .Q(u0_csc1_21_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_i_bF_buf90), .D(u0_u1__0csc_31_0__22_), .Q(u0_csc1_22_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_i_bF_buf89), .D(u0_u1__0csc_31_0__23_), .Q(u0_csc1_23_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_i_bF_buf88), .D(u0_u1__0csc_31_0__24_), .Q(u0_csc1_24_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_i_bF_buf87), .D(u0_u1__0csc_31_0__25_), .Q(u0_csc1_25_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_i_bF_buf86), .D(u0_u1__0csc_31_0__26_), .Q(u0_csc1_26_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_i_bF_buf80), .D(u0__0poc_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_85523_13_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_i_bF_buf85), .D(u0_u1__0csc_31_0__27_), .Q(u0_csc1_27_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_i_bF_buf84), .D(u0_u1__0csc_31_0__28_), .Q(u0_csc1_28_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_i_bF_buf83), .D(u0_u1__0csc_31_0__29_), .Q(u0_csc1_29_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_i_bF_buf82), .D(u0_u1__0csc_31_0__30_), .Q(u0_csc1_30_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_i_bF_buf81), .D(u0_u1__0csc_31_0__31_), .Q(u0_csc1_31_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_i_bF_buf80), .D(\wb_addr_i[2] ), .Q(u0_u1_addr_r_2_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_i_bF_buf79), .D(\wb_addr_i[3] ), .Q(u0_u1_addr_r_3_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_i_bF_buf78), .D(\wb_addr_i[4] ), .Q(u0_u1_addr_r_4_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_i_bF_buf77), .D(\wb_addr_i[5] ), .Q(u0_u1_addr_r_5_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_i_bF_buf76), .D(\wb_addr_i[6] ), .Q(u0_u1_addr_r_6_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_i_bF_buf79), .D(u0__0poc_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_85523_14_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_i_bF_buf69), .D(u1__0bank_adr_1_0__0_), .Q(bank_adr_0_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_i_bF_buf68), .D(u1__0bank_adr_1_0__1_), .Q(bank_adr_1_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_i_bF_buf67), .D(u1__0row_adr_12_0__0_), .Q(row_adr_0_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_i_bF_buf66), .D(u1__0row_adr_12_0__1_), .Q(row_adr_1_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_i_bF_buf65), .D(u1__0row_adr_12_0__2_), .Q(row_adr_2_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_i_bF_buf64), .D(u1__0row_adr_12_0__3_), .Q(row_adr_3_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_i_bF_buf63), .D(u1__0row_adr_12_0__4_), .Q(row_adr_4_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_i_bF_buf62), .D(u1__0row_adr_12_0__5_), .Q(row_adr_5_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_i_bF_buf61), .D(u1__0row_adr_12_0__6_), .Q(row_adr_6_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_i_bF_buf60), .D(u1__0row_adr_12_0__7_), .Q(row_adr_7_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_i_bF_buf78), .D(u0__0poc_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_85523_15_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_i_bF_buf59), .D(u1__0row_adr_12_0__8_), .Q(row_adr_8_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_i_bF_buf58), .D(u1__0row_adr_12_0__9_), .Q(row_adr_9_));
DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_i_bF_buf57), .D(u1__0row_adr_12_0__10_), .Q(row_adr_10_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_i_bF_buf56), .D(u1__0row_adr_12_0__11_), .Q(row_adr_11_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_i_bF_buf55), .D(u1__0row_adr_12_0__12_), .Q(row_adr_12_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_i_bF_buf54), .D(u1__0col_adr_9_0__0_), .Q(u1_col_adr_0_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_i_bF_buf53), .D(u1__0col_adr_9_0__1_), .Q(u1_col_adr_1_));
DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_i_bF_buf52), .D(u1__0col_adr_9_0__2_), .Q(u1_col_adr_2_));
DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_i_bF_buf51), .D(u1__0col_adr_9_0__3_), .Q(u1_col_adr_3_));
DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_i_bF_buf50), .D(u1__0col_adr_9_0__4_), .Q(u1_col_adr_4_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_i_bF_buf95), .D(lmr_ack), .Q(u0_lmr_ack_r));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_i_bF_buf77), .D(u0__0poc_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_85523_16_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_i_bF_buf49), .D(u1__0col_adr_9_0__5_), .Q(u1_col_adr_5_));
DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_i_bF_buf48), .D(u1__0col_adr_9_0__6_), .Q(u1_col_adr_6_));
DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_i_bF_buf47), .D(u1__0col_adr_9_0__7_), .Q(u1_col_adr_7_));
DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_i_bF_buf46), .D(u1__0col_adr_9_0__8_), .Q(u1_col_adr_8_));
DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_i_bF_buf45), .D(u1__0col_adr_9_0__9_), .Q(u1_col_adr_9_));
DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_i_bF_buf44), .D(u1__0acs_addr_23_0__0_), .Q(u1_acs_addr_0_));
DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_i_bF_buf43), .D(u1__0acs_addr_23_0__1_), .Q(u1_acs_addr_1_));
DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_i_bF_buf42), .D(u1__0acs_addr_23_0__2_), .Q(u1_acs_addr_2_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_i_bF_buf41), .D(u1__0acs_addr_23_0__3_), .Q(u1_acs_addr_3_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_i_bF_buf40), .D(u1__0acs_addr_23_0__4_), .Q(u1_acs_addr_4_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_i_bF_buf76), .D(u0__0poc_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_85523_17_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_i_bF_buf39), .D(u1__0acs_addr_23_0__5_), .Q(u1_acs_addr_5_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_i_bF_buf38), .D(u1__0acs_addr_23_0__6_), .Q(u1_acs_addr_6_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_i_bF_buf37), .D(u1__0acs_addr_23_0__7_), .Q(u1_acs_addr_7_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_i_bF_buf36), .D(u1__0acs_addr_23_0__8_), .Q(u1_acs_addr_8_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_i_bF_buf35), .D(u1__0acs_addr_23_0__9_), .Q(u1_acs_addr_9_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_i_bF_buf34), .D(u1__0acs_addr_23_0__10_), .Q(u1_acs_addr_10_));
DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_i_bF_buf33), .D(u1__0acs_addr_23_0__11_), .Q(u1_acs_addr_11_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_i_bF_buf32), .D(u1__0acs_addr_23_0__12_), .Q(u1_acs_addr_12_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_i_bF_buf31), .D(u1__0acs_addr_23_0__13_), .Q(u1_acs_addr_13_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_i_bF_buf30), .D(u1__0acs_addr_23_0__14_), .Q(u1_acs_addr_14_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_i_bF_buf75), .D(u0__0poc_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_85523_18_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_i_bF_buf29), .D(u1__0acs_addr_23_0__15_), .Q(u1_acs_addr_15_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_i_bF_buf28), .D(u1__0acs_addr_23_0__16_), .Q(u1_acs_addr_16_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_i_bF_buf27), .D(u1__0acs_addr_23_0__17_), .Q(u1_acs_addr_17_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_i_bF_buf26), .D(u1__0acs_addr_23_0__18_), .Q(u1_acs_addr_18_));
DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_i_bF_buf25), .D(u1__0acs_addr_23_0__19_), .Q(u1_acs_addr_19_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_i_bF_buf24), .D(u1__0acs_addr_23_0__20_), .Q(u1_acs_addr_20_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_i_bF_buf23), .D(u1__0acs_addr_23_0__21_), .Q(u1_acs_addr_21_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_i_bF_buf22), .D(u1__0acs_addr_23_0__22_), .Q(u1_acs_addr_22_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_i_bF_buf21), .D(u1__0acs_addr_23_0__23_), .Q(u1_acs_addr_23_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_i_bF_buf20), .D(u1__0sram_addr_23_0__0_), .Q(u1_sram_addr_0_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_i_bF_buf74), .D(u0__0poc_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_85523_19_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_i_bF_buf19), .D(u1__0sram_addr_23_0__1_), .Q(u1_sram_addr_1_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_i_bF_buf18), .D(u1__0sram_addr_23_0__2_), .Q(u1_sram_addr_2_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_i_bF_buf17), .D(u1__0sram_addr_23_0__3_), .Q(u1_sram_addr_3_));
DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_i_bF_buf16), .D(u1__0sram_addr_23_0__4_), .Q(u1_sram_addr_4_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_i_bF_buf15), .D(u1__0sram_addr_23_0__5_), .Q(u1_sram_addr_5_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_i_bF_buf14), .D(u1__0sram_addr_23_0__6_), .Q(u1_sram_addr_6_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_i_bF_buf13), .D(u1__0sram_addr_23_0__7_), .Q(u1_sram_addr_7_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_i_bF_buf12), .D(u1__0sram_addr_23_0__8_), .Q(u1_sram_addr_8_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_i_bF_buf11), .D(u1__0sram_addr_23_0__9_), .Q(u1_sram_addr_9_));
DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_i_bF_buf10), .D(u1__0sram_addr_23_0__10_), .Q(u1_sram_addr_10_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_i_bF_buf73), .D(u0__0poc_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_85523_20_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_i_bF_buf9), .D(u1__0sram_addr_23_0__11_), .Q(u1_sram_addr_11_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_i_bF_buf8), .D(u1__0sram_addr_23_0__12_), .Q(u1_sram_addr_12_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_i_bF_buf7), .D(u1__0sram_addr_23_0__13_), .Q(u1_sram_addr_13_));
DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_i_bF_buf6), .D(u1__0sram_addr_23_0__14_), .Q(u1_sram_addr_14_));
DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_i_bF_buf5), .D(u1__0sram_addr_23_0__15_), .Q(u1_sram_addr_15_));
DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_i_bF_buf4), .D(u1__0sram_addr_23_0__16_), .Q(u1_sram_addr_16_));
DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_i_bF_buf3), .D(u1__0sram_addr_23_0__17_), .Q(u1_sram_addr_17_));
DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_i_bF_buf2), .D(u1__0sram_addr_23_0__18_), .Q(u1_sram_addr_18_));
DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_i_bF_buf1), .D(u1__0sram_addr_23_0__19_), .Q(u1_sram_addr_19_));
DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_i_bF_buf0), .D(u1__0sram_addr_23_0__20_), .Q(u1_sram_addr_20_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_i_bF_buf72), .D(u0__0poc_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_85523_21_));
DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_i_bF_buf96), .D(u1__0sram_addr_23_0__21_), .Q(u1_sram_addr_21_));
DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_i_bF_buf95), .D(u1__0sram_addr_23_0__22_), .Q(u1_sram_addr_22_));
DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_i_bF_buf94), .D(u1__0sram_addr_23_0__23_), .Q(u1_sram_addr_23_));
DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_i_bF_buf93), .D(u1_u0__0out_r_12_0__0_), .Q(u1_acs_addr_pl1_0_));
DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_i_bF_buf92), .D(u1_u0__0out_r_12_0__1_), .Q(u1_acs_addr_pl1_1_));
DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_i_bF_buf91), .D(u1_u0__0out_r_12_0__2_), .Q(u1_acs_addr_pl1_2_));
DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_i_bF_buf90), .D(u1_u0__0out_r_12_0__3_), .Q(u1_acs_addr_pl1_3_));
DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_i_bF_buf89), .D(u1_u0__0out_r_12_0__4_), .Q(u1_acs_addr_pl1_4_));
DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_i_bF_buf88), .D(u1_u0__0out_r_12_0__5_), .Q(u1_acs_addr_pl1_5_));
DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_i_bF_buf87), .D(u1_u0__0out_r_12_0__6_), .Q(u1_acs_addr_pl1_6_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_i_bF_buf71), .D(u0__0poc_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_85523_22_));
DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_i_bF_buf86), .D(u1_u0__0out_r_12_0__7_), .Q(u1_acs_addr_pl1_7_));
DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_i_bF_buf85), .D(u1_u0__0out_r_12_0__8_), .Q(u1_acs_addr_pl1_8_));
DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_i_bF_buf84), .D(u1_u0__0out_r_12_0__9_), .Q(u1_acs_addr_pl1_9_));
DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_i_bF_buf83), .D(u1_u0__0out_r_12_0__10_), .Q(u1_acs_addr_pl1_10_));
DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_i_bF_buf82), .D(u1_u0__0out_r_12_0__11_), .Q(u1_acs_addr_pl1_11_));
DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_i_bF_buf81), .D(u1_u0__0out_r_12_0__12_), .Q(u1_u0_inc_next));
DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_i_bF_buf80), .D(u2__0row_same_0_0_), .Q(row_same));
DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_i_bF_buf79), .D(u2__0bank_open_0_0_), .Q(bank_open));
DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_i_bF_buf78), .D(u2_u0__0b3_last_row_12_0__0_), .Q(u2_u0_b3_last_row_0_));
DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_i_bF_buf77), .D(u2_u0__0b3_last_row_12_0__1_), .Q(u2_u0_b3_last_row_1_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_i_bF_buf70), .D(u0__0poc_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_85523_23_));
DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_i_bF_buf76), .D(u2_u0__0b3_last_row_12_0__2_), .Q(u2_u0_b3_last_row_2_));
DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_i_bF_buf75), .D(u2_u0__0b3_last_row_12_0__3_), .Q(u2_u0_b3_last_row_3_));
DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_i_bF_buf74), .D(u2_u0__0b3_last_row_12_0__4_), .Q(u2_u0_b3_last_row_4_));
DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_i_bF_buf73), .D(u2_u0__0b3_last_row_12_0__5_), .Q(u2_u0_b3_last_row_5_));
DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_i_bF_buf72), .D(u2_u0__0b3_last_row_12_0__6_), .Q(u2_u0_b3_last_row_6_));
DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_i_bF_buf71), .D(u2_u0__0b3_last_row_12_0__7_), .Q(u2_u0_b3_last_row_7_));
DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_i_bF_buf70), .D(u2_u0__0b3_last_row_12_0__8_), .Q(u2_u0_b3_last_row_8_));
DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_i_bF_buf69), .D(u2_u0__0b3_last_row_12_0__9_), .Q(u2_u0_b3_last_row_9_));
DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_i_bF_buf68), .D(u2_u0__0b3_last_row_12_0__10_), .Q(u2_u0_b3_last_row_10_));
DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_i_bF_buf67), .D(u2_u0__0b3_last_row_12_0__11_), .Q(u2_u0_b3_last_row_11_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_i_bF_buf69), .D(u0__0poc_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_85523_24_));
DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_i_bF_buf66), .D(u2_u0__0b3_last_row_12_0__12_), .Q(u2_u0_b3_last_row_12_));
DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_i_bF_buf65), .D(u2_u0__0b2_last_row_12_0__0_), .Q(u2_u0_b2_last_row_0_));
DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_i_bF_buf64), .D(u2_u0__0b2_last_row_12_0__1_), .Q(u2_u0_b2_last_row_1_));
DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_i_bF_buf63), .D(u2_u0__0b2_last_row_12_0__2_), .Q(u2_u0_b2_last_row_2_));
DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_i_bF_buf62), .D(u2_u0__0b2_last_row_12_0__3_), .Q(u2_u0_b2_last_row_3_));
DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_i_bF_buf61), .D(u2_u0__0b2_last_row_12_0__4_), .Q(u2_u0_b2_last_row_4_));
DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_i_bF_buf60), .D(u2_u0__0b2_last_row_12_0__5_), .Q(u2_u0_b2_last_row_5_));
DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_i_bF_buf59), .D(u2_u0__0b2_last_row_12_0__6_), .Q(u2_u0_b2_last_row_6_));
DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_i_bF_buf58), .D(u2_u0__0b2_last_row_12_0__7_), .Q(u2_u0_b2_last_row_7_));
DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_i_bF_buf57), .D(u2_u0__0b2_last_row_12_0__8_), .Q(u2_u0_b2_last_row_8_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_i_bF_buf68), .D(u0__0poc_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_85523_25_));
DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_i_bF_buf56), .D(u2_u0__0b2_last_row_12_0__9_), .Q(u2_u0_b2_last_row_9_));
DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_i_bF_buf55), .D(u2_u0__0b2_last_row_12_0__10_), .Q(u2_u0_b2_last_row_10_));
DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_i_bF_buf54), .D(u2_u0__0b2_last_row_12_0__11_), .Q(u2_u0_b2_last_row_11_));
DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_i_bF_buf53), .D(u2_u0__0b2_last_row_12_0__12_), .Q(u2_u0_b2_last_row_12_));
DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_i_bF_buf52), .D(u2_u0__0b1_last_row_12_0__0_), .Q(u2_u0_b1_last_row_0_));
DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_i_bF_buf51), .D(u2_u0__0b1_last_row_12_0__1_), .Q(u2_u0_b1_last_row_1_));
DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_i_bF_buf50), .D(u2_u0__0b1_last_row_12_0__2_), .Q(u2_u0_b1_last_row_2_));
DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_i_bF_buf49), .D(u2_u0__0b1_last_row_12_0__3_), .Q(u2_u0_b1_last_row_3_));
DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_i_bF_buf48), .D(u2_u0__0b1_last_row_12_0__4_), .Q(u2_u0_b1_last_row_4_));
DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_i_bF_buf47), .D(u2_u0__0b1_last_row_12_0__5_), .Q(u2_u0_b1_last_row_5_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_i_bF_buf94), .D(init_ack), .Q(u0_init_ack_r));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_i_bF_buf67), .D(u0__0poc_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_85523_26_));
DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_i_bF_buf46), .D(u2_u0__0b1_last_row_12_0__6_), .Q(u2_u0_b1_last_row_6_));
DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_i_bF_buf45), .D(u2_u0__0b1_last_row_12_0__7_), .Q(u2_u0_b1_last_row_7_));
DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_i_bF_buf44), .D(u2_u0__0b1_last_row_12_0__8_), .Q(u2_u0_b1_last_row_8_));
DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_i_bF_buf43), .D(u2_u0__0b1_last_row_12_0__9_), .Q(u2_u0_b1_last_row_9_));
DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_i_bF_buf42), .D(u2_u0__0b1_last_row_12_0__10_), .Q(u2_u0_b1_last_row_10_));
DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_i_bF_buf41), .D(u2_u0__0b1_last_row_12_0__11_), .Q(u2_u0_b1_last_row_11_));
DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_i_bF_buf40), .D(u2_u0__0b1_last_row_12_0__12_), .Q(u2_u0_b1_last_row_12_));
DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_i_bF_buf39), .D(u2_u0__0b0_last_row_12_0__0_), .Q(u2_u0_b0_last_row_0_));
DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_i_bF_buf38), .D(u2_u0__0b0_last_row_12_0__1_), .Q(u2_u0_b0_last_row_1_));
DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_i_bF_buf37), .D(u2_u0__0b0_last_row_12_0__2_), .Q(u2_u0_b0_last_row_2_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_i_bF_buf66), .D(u0__0poc_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_85523_27_));
DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_i_bF_buf36), .D(u2_u0__0b0_last_row_12_0__3_), .Q(u2_u0_b0_last_row_3_));
DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_i_bF_buf35), .D(u2_u0__0b0_last_row_12_0__4_), .Q(u2_u0_b0_last_row_4_));
DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_i_bF_buf34), .D(u2_u0__0b0_last_row_12_0__5_), .Q(u2_u0_b0_last_row_5_));
DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_i_bF_buf33), .D(u2_u0__0b0_last_row_12_0__6_), .Q(u2_u0_b0_last_row_6_));
DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_i_bF_buf32), .D(u2_u0__0b0_last_row_12_0__7_), .Q(u2_u0_b0_last_row_7_));
DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_i_bF_buf31), .D(u2_u0__0b0_last_row_12_0__8_), .Q(u2_u0_b0_last_row_8_));
DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_i_bF_buf30), .D(u2_u0__0b0_last_row_12_0__9_), .Q(u2_u0_b0_last_row_9_));
DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_i_bF_buf29), .D(u2_u0__0b0_last_row_12_0__10_), .Q(u2_u0_b0_last_row_10_));
DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_i_bF_buf28), .D(u2_u0__0b0_last_row_12_0__11_), .Q(u2_u0_b0_last_row_11_));
DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_i_bF_buf27), .D(u2_u0__0b0_last_row_12_0__12_), .Q(u2_u0_b0_last_row_12_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_i_bF_buf65), .D(u0__0poc_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_85523_28_));
DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_i_bF_buf22), .D(u2_u1__0b3_last_row_12_0__0_), .Q(u2_u1_b3_last_row_0_));
DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_i_bF_buf21), .D(u2_u1__0b3_last_row_12_0__1_), .Q(u2_u1_b3_last_row_1_));
DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_i_bF_buf20), .D(u2_u1__0b3_last_row_12_0__2_), .Q(u2_u1_b3_last_row_2_));
DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_i_bF_buf19), .D(u2_u1__0b3_last_row_12_0__3_), .Q(u2_u1_b3_last_row_3_));
DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_i_bF_buf18), .D(u2_u1__0b3_last_row_12_0__4_), .Q(u2_u1_b3_last_row_4_));
DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_i_bF_buf17), .D(u2_u1__0b3_last_row_12_0__5_), .Q(u2_u1_b3_last_row_5_));
DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_i_bF_buf16), .D(u2_u1__0b3_last_row_12_0__6_), .Q(u2_u1_b3_last_row_6_));
DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_i_bF_buf15), .D(u2_u1__0b3_last_row_12_0__7_), .Q(u2_u1_b3_last_row_7_));
DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_i_bF_buf14), .D(u2_u1__0b3_last_row_12_0__8_), .Q(u2_u1_b3_last_row_8_));
DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_i_bF_buf13), .D(u2_u1__0b3_last_row_12_0__9_), .Q(u2_u1_b3_last_row_9_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_i_bF_buf64), .D(u0__0poc_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_85523_29_));
DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_i_bF_buf12), .D(u2_u1__0b3_last_row_12_0__10_), .Q(u2_u1_b3_last_row_10_));
DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_i_bF_buf11), .D(u2_u1__0b3_last_row_12_0__11_), .Q(u2_u1_b3_last_row_11_));
DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_i_bF_buf10), .D(u2_u1__0b3_last_row_12_0__12_), .Q(u2_u1_b3_last_row_12_));
DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_i_bF_buf9), .D(u2_u1__0b2_last_row_12_0__0_), .Q(u2_u1_b2_last_row_0_));
DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_i_bF_buf8), .D(u2_u1__0b2_last_row_12_0__1_), .Q(u2_u1_b2_last_row_1_));
DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_i_bF_buf7), .D(u2_u1__0b2_last_row_12_0__2_), .Q(u2_u1_b2_last_row_2_));
DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_i_bF_buf6), .D(u2_u1__0b2_last_row_12_0__3_), .Q(u2_u1_b2_last_row_3_));
DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_i_bF_buf5), .D(u2_u1__0b2_last_row_12_0__4_), .Q(u2_u1_b2_last_row_4_));
DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_i_bF_buf4), .D(u2_u1__0b2_last_row_12_0__5_), .Q(u2_u1_b2_last_row_5_));
DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_i_bF_buf3), .D(u2_u1__0b2_last_row_12_0__6_), .Q(u2_u1_b2_last_row_6_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_i_bF_buf63), .D(u0__0poc_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_85523_30_));
DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_i_bF_buf2), .D(u2_u1__0b2_last_row_12_0__7_), .Q(u2_u1_b2_last_row_7_));
DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_i_bF_buf1), .D(u2_u1__0b2_last_row_12_0__8_), .Q(u2_u1_b2_last_row_8_));
DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_i_bF_buf0), .D(u2_u1__0b2_last_row_12_0__9_), .Q(u2_u1_b2_last_row_9_));
DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_i_bF_buf96), .D(u2_u1__0b2_last_row_12_0__10_), .Q(u2_u1_b2_last_row_10_));
DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_i_bF_buf95), .D(u2_u1__0b2_last_row_12_0__11_), .Q(u2_u1_b2_last_row_11_));
DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_i_bF_buf94), .D(u2_u1__0b2_last_row_12_0__12_), .Q(u2_u1_b2_last_row_12_));
DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_i_bF_buf93), .D(u2_u1__0b1_last_row_12_0__0_), .Q(u2_u1_b1_last_row_0_));
DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_i_bF_buf92), .D(u2_u1__0b1_last_row_12_0__1_), .Q(u2_u1_b1_last_row_1_));
DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_i_bF_buf91), .D(u2_u1__0b1_last_row_12_0__2_), .Q(u2_u1_b1_last_row_2_));
DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_i_bF_buf90), .D(u2_u1__0b1_last_row_12_0__3_), .Q(u2_u1_b1_last_row_3_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_i_bF_buf62), .D(u0__0poc_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_85523_31_));
DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_i_bF_buf89), .D(u2_u1__0b1_last_row_12_0__4_), .Q(u2_u1_b1_last_row_4_));
DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_i_bF_buf88), .D(u2_u1__0b1_last_row_12_0__5_), .Q(u2_u1_b1_last_row_5_));
DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_i_bF_buf87), .D(u2_u1__0b1_last_row_12_0__6_), .Q(u2_u1_b1_last_row_6_));
DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_i_bF_buf86), .D(u2_u1__0b1_last_row_12_0__7_), .Q(u2_u1_b1_last_row_7_));
DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_i_bF_buf85), .D(u2_u1__0b1_last_row_12_0__8_), .Q(u2_u1_b1_last_row_8_));
DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_i_bF_buf84), .D(u2_u1__0b1_last_row_12_0__9_), .Q(u2_u1_b1_last_row_9_));
DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_i_bF_buf83), .D(u2_u1__0b1_last_row_12_0__10_), .Q(u2_u1_b1_last_row_10_));
DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_i_bF_buf82), .D(u2_u1__0b1_last_row_12_0__11_), .Q(u2_u1_b1_last_row_11_));
DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_i_bF_buf81), .D(u2_u1__0b1_last_row_12_0__12_), .Q(u2_u1_b1_last_row_12_));
DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_i_bF_buf80), .D(u2_u1__0b0_last_row_12_0__0_), .Q(u2_u1_b0_last_row_0_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_i_bF_buf61), .D(mc_sts_ir), .Q(u0_csr_0_));
DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_i_bF_buf79), .D(u2_u1__0b0_last_row_12_0__1_), .Q(u2_u1_b0_last_row_1_));
DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_i_bF_buf78), .D(u2_u1__0b0_last_row_12_0__2_), .Q(u2_u1_b0_last_row_2_));
DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_i_bF_buf77), .D(u2_u1__0b0_last_row_12_0__3_), .Q(u2_u1_b0_last_row_3_));
DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_i_bF_buf76), .D(u2_u1__0b0_last_row_12_0__4_), .Q(u2_u1_b0_last_row_4_));
DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_i_bF_buf75), .D(u2_u1__0b0_last_row_12_0__5_), .Q(u2_u1_b0_last_row_5_));
DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_i_bF_buf74), .D(u2_u1__0b0_last_row_12_0__6_), .Q(u2_u1_b0_last_row_6_));
DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_i_bF_buf73), .D(u2_u1__0b0_last_row_12_0__7_), .Q(u2_u1_b0_last_row_7_));
DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_i_bF_buf72), .D(u2_u1__0b0_last_row_12_0__8_), .Q(u2_u1_b0_last_row_8_));
DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_i_bF_buf71), .D(u2_u1__0b0_last_row_12_0__9_), .Q(u2_u1_b0_last_row_9_));
DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_i_bF_buf70), .D(u2_u1__0b0_last_row_12_0__10_), .Q(u2_u1_b0_last_row_10_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_i_bF_buf60), .D(\wb_addr_i[2] ), .Q(u0_wb_addr_r_2_));
DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_i_bF_buf69), .D(u2_u1__0b0_last_row_12_0__11_), .Q(u2_u1_b0_last_row_11_));
DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_i_bF_buf68), .D(u2_u1__0b0_last_row_12_0__12_), .Q(u2_u1_b0_last_row_12_));
DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_i_bF_buf63), .D(u3__0mc_dp_o_3_0__0_), .Q(mc_dp_od_0_));
DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_i_bF_buf62), .D(u3__0mc_dp_o_3_0__1_), .Q(mc_dp_od_1_));
DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_i_bF_buf61), .D(u3__0mc_dp_o_3_0__2_), .Q(mc_dp_od_2_));
DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_i_bF_buf60), .D(u3__0mc_dp_o_3_0__3_), .Q(mc_dp_od_3_));
DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_i_bF_buf59), .D(u3__0byte2_7_0__0_), .Q(u3_byte2_0_));
DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_i_bF_buf58), .D(u3__0byte2_7_0__1_), .Q(u3_byte2_1_));
DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_i_bF_buf57), .D(u3__0byte2_7_0__2_), .Q(u3_byte2_2_));
DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_i_bF_buf56), .D(u3__0byte2_7_0__3_), .Q(u3_byte2_3_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_i_bF_buf59), .D(\wb_addr_i[3] ), .Q(u0_wb_addr_r_3_));
DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_i_bF_buf55), .D(u3__0byte2_7_0__4_), .Q(u3_byte2_4_));
DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_i_bF_buf54), .D(u3__0byte2_7_0__5_), .Q(u3_byte2_5_));
DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_i_bF_buf53), .D(u3__0byte2_7_0__6_), .Q(u3_byte2_6_));
DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_i_bF_buf52), .D(u3__0byte2_7_0__7_), .Q(u3_byte2_7_));
DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_i_bF_buf51), .D(u3__0byte1_7_0__0_), .Q(u3_byte1_0_));
DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_i_bF_buf50), .D(u3__0byte1_7_0__1_), .Q(u3_byte1_1_));
DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_i_bF_buf49), .D(u3__0byte1_7_0__2_), .Q(u3_byte1_2_));
DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_i_bF_buf48), .D(u3__0byte1_7_0__3_), .Q(u3_byte1_3_));
DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_i_bF_buf47), .D(u3__0byte1_7_0__4_), .Q(u3_byte1_4_));
DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_i_bF_buf46), .D(u3__0byte1_7_0__5_), .Q(u3_byte1_5_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_i_bF_buf58), .D(\wb_addr_i[4] ), .Q(u0_wb_addr_r_4_));
DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_i_bF_buf45), .D(u3__0byte1_7_0__6_), .Q(u3_byte1_6_));
DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_i_bF_buf44), .D(u3__0byte1_7_0__7_), .Q(u3_byte1_7_));
DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_i_bF_buf43), .D(u3__0byte0_7_0__0_), .Q(u3_byte0_0_));
DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_i_bF_buf42), .D(u3__0byte0_7_0__1_), .Q(u3_byte0_1_));
DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_i_bF_buf41), .D(u3__0byte0_7_0__2_), .Q(u3_byte0_2_));
DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_i_bF_buf40), .D(u3__0byte0_7_0__3_), .Q(u3_byte0_3_));
DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_i_bF_buf39), .D(u3__0byte0_7_0__4_), .Q(u3_byte0_4_));
DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_i_bF_buf38), .D(u3__0byte0_7_0__5_), .Q(u3_byte0_5_));
DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_i_bF_buf37), .D(u3__0byte0_7_0__6_), .Q(u3_byte0_6_));
DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_i_bF_buf36), .D(u3__0byte0_7_0__7_), .Q(u3_byte0_7_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_i_bF_buf93), .D(u0__0poc_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_85523_0_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_i_bF_buf57), .D(\wb_addr_i[5] ), .Q(u0_wb_addr_r_5_));
DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_i_bF_buf35), .D(u3__0mc_data_o_31_0__0_), .Q(mc_data_od_0_));
DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_i_bF_buf34), .D(u3__0mc_data_o_31_0__1_), .Q(mc_data_od_1_));
DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_i_bF_buf33), .D(u3__0mc_data_o_31_0__2_), .Q(mc_data_od_2_));
DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_i_bF_buf32), .D(u3__0mc_data_o_31_0__3_), .Q(mc_data_od_3_));
DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_i_bF_buf31), .D(u3__0mc_data_o_31_0__4_), .Q(mc_data_od_4_));
DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_i_bF_buf30), .D(u3__0mc_data_o_31_0__5_), .Q(mc_data_od_5_));
DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_i_bF_buf29), .D(u3__0mc_data_o_31_0__6_), .Q(mc_data_od_6_));
DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_i_bF_buf28), .D(u3__0mc_data_o_31_0__7_), .Q(mc_data_od_7_));
DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_i_bF_buf27), .D(u3__0mc_data_o_31_0__8_), .Q(mc_data_od_8_));
DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_i_bF_buf26), .D(u3__0mc_data_o_31_0__9_), .Q(mc_data_od_9_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_i_bF_buf56), .D(\wb_addr_i[6] ), .Q(u0_wb_addr_r_6_));
DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_i_bF_buf25), .D(u3__0mc_data_o_31_0__10_), .Q(mc_data_od_10_));
DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_i_bF_buf24), .D(u3__0mc_data_o_31_0__11_), .Q(mc_data_od_11_));
DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_i_bF_buf23), .D(u3__0mc_data_o_31_0__12_), .Q(mc_data_od_12_));
DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_i_bF_buf22), .D(u3__0mc_data_o_31_0__13_), .Q(mc_data_od_13_));
DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_i_bF_buf21), .D(u3__0mc_data_o_31_0__14_), .Q(mc_data_od_14_));
DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_i_bF_buf20), .D(u3__0mc_data_o_31_0__15_), .Q(mc_data_od_15_));
DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_i_bF_buf19), .D(u3__0mc_data_o_31_0__16_), .Q(mc_data_od_16_));
DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_i_bF_buf18), .D(u3__0mc_data_o_31_0__17_), .Q(mc_data_od_17_));
DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_i_bF_buf17), .D(u3__0mc_data_o_31_0__18_), .Q(mc_data_od_18_));
DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_i_bF_buf16), .D(u3__0mc_data_o_31_0__19_), .Q(mc_data_od_19_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_i_bF_buf25), .D(u0_u0__0tms_31_0__0_), .Q(u0_tms0_0_));
DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_i_bF_buf15), .D(u3__0mc_data_o_31_0__20_), .Q(mc_data_od_20_));
DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_i_bF_buf14), .D(u3__0mc_data_o_31_0__21_), .Q(mc_data_od_21_));
DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_i_bF_buf13), .D(u3__0mc_data_o_31_0__22_), .Q(mc_data_od_22_));
DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_i_bF_buf12), .D(u3__0mc_data_o_31_0__23_), .Q(mc_data_od_23_));
DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_i_bF_buf11), .D(u3__0mc_data_o_31_0__24_), .Q(mc_data_od_24_));
DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_i_bF_buf10), .D(u3__0mc_data_o_31_0__25_), .Q(mc_data_od_25_));
DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_i_bF_buf9), .D(u3__0mc_data_o_31_0__26_), .Q(mc_data_od_26_));
DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_i_bF_buf8), .D(u3__0mc_data_o_31_0__27_), .Q(mc_data_od_27_));
DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_i_bF_buf7), .D(u3__0mc_data_o_31_0__28_), .Q(mc_data_od_28_));
DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_i_bF_buf6), .D(u3__0mc_data_o_31_0__29_), .Q(mc_data_od_29_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_i_bF_buf24), .D(u0_u0__0tms_31_0__1_), .Q(u0_tms0_1_));
DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_i_bF_buf5), .D(u3__0mc_data_o_31_0__30_), .Q(mc_data_od_30_));
DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_i_bF_buf4), .D(u3__0mc_data_o_31_0__31_), .Q(mc_data_od_31_));
DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_i_bF_buf3), .D(u3_u0__0r3_35_0__0_), .Q(u3_u0_r3_0_));
DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_i_bF_buf2), .D(u3_u0__0r3_35_0__1_), .Q(u3_u0_r3_1_));
DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_i_bF_buf1), .D(u3_u0__0r3_35_0__2_), .Q(u3_u0_r3_2_));
DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_i_bF_buf0), .D(u3_u0__0r3_35_0__3_), .Q(u3_u0_r3_3_));
DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_i_bF_buf96), .D(u3_u0__0r3_35_0__4_), .Q(u3_u0_r3_4_));
DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_i_bF_buf95), .D(u3_u0__0r3_35_0__5_), .Q(u3_u0_r3_5_));
DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_i_bF_buf94), .D(u3_u0__0r3_35_0__6_), .Q(u3_u0_r3_6_));
DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_i_bF_buf93), .D(u3_u0__0r3_35_0__7_), .Q(u3_u0_r3_7_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_i_bF_buf23), .D(u0_u0__0tms_31_0__2_), .Q(u0_tms0_2_));
DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_i_bF_buf92), .D(u3_u0__0r3_35_0__8_), .Q(u3_u0_r3_8_));
DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_i_bF_buf91), .D(u3_u0__0r3_35_0__9_), .Q(u3_u0_r3_9_));
DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_i_bF_buf90), .D(u3_u0__0r3_35_0__10_), .Q(u3_u0_r3_10_));
DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_i_bF_buf89), .D(u3_u0__0r3_35_0__11_), .Q(u3_u0_r3_11_));
DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_i_bF_buf88), .D(u3_u0__0r3_35_0__12_), .Q(u3_u0_r3_12_));
DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_i_bF_buf87), .D(u3_u0__0r3_35_0__13_), .Q(u3_u0_r3_13_));
DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_i_bF_buf86), .D(u3_u0__0r3_35_0__14_), .Q(u3_u0_r3_14_));
DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_i_bF_buf85), .D(u3_u0__0r3_35_0__15_), .Q(u3_u0_r3_15_));
DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_i_bF_buf84), .D(u3_u0__0r3_35_0__16_), .Q(u3_u0_r3_16_));
DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_i_bF_buf83), .D(u3_u0__0r3_35_0__17_), .Q(u3_u0_r3_17_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_i_bF_buf22), .D(u0_u0__0tms_31_0__3_), .Q(u0_tms0_3_));
DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_i_bF_buf82), .D(u3_u0__0r3_35_0__18_), .Q(u3_u0_r3_18_));
DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_i_bF_buf81), .D(u3_u0__0r3_35_0__19_), .Q(u3_u0_r3_19_));
DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_i_bF_buf80), .D(u3_u0__0r3_35_0__20_), .Q(u3_u0_r3_20_));
DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_i_bF_buf79), .D(u3_u0__0r3_35_0__21_), .Q(u3_u0_r3_21_));
DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_i_bF_buf78), .D(u3_u0__0r3_35_0__22_), .Q(u3_u0_r3_22_));
DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_i_bF_buf77), .D(u3_u0__0r3_35_0__23_), .Q(u3_u0_r3_23_));
DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_i_bF_buf76), .D(u3_u0__0r3_35_0__24_), .Q(u3_u0_r3_24_));
DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_i_bF_buf75), .D(u3_u0__0r3_35_0__25_), .Q(u3_u0_r3_25_));
DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_i_bF_buf74), .D(u3_u0__0r3_35_0__26_), .Q(u3_u0_r3_26_));
DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_i_bF_buf73), .D(u3_u0__0r3_35_0__27_), .Q(u3_u0_r3_27_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_i_bF_buf21), .D(u0_u0__0tms_31_0__4_), .Q(u0_tms0_4_));
DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_i_bF_buf72), .D(u3_u0__0r3_35_0__28_), .Q(u3_u0_r3_28_));
DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_i_bF_buf71), .D(u3_u0__0r3_35_0__29_), .Q(u3_u0_r3_29_));
DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_i_bF_buf70), .D(u3_u0__0r3_35_0__30_), .Q(u3_u0_r3_30_));
DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_i_bF_buf69), .D(u3_u0__0r3_35_0__31_), .Q(u3_u0_r3_31_));
DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_i_bF_buf68), .D(u3_u0__0r3_35_0__32_), .Q(u3_u0_r3_32_));
DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_i_bF_buf67), .D(u3_u0__0r3_35_0__33_), .Q(u3_u0_r3_33_));
DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_i_bF_buf66), .D(u3_u0__0r3_35_0__34_), .Q(u3_u0_r3_34_));
DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_i_bF_buf65), .D(u3_u0__0r3_35_0__35_), .Q(u3_u0_r3_35_));
DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_i_bF_buf64), .D(u3_u0__0r2_35_0__0_), .Q(u3_u0_r2_0_));
DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_i_bF_buf63), .D(u3_u0__0r2_35_0__1_), .Q(u3_u0_r2_1_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_i_bF_buf20), .D(u0_u0__0tms_31_0__5_), .Q(u0_tms0_5_));
DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_i_bF_buf62), .D(u3_u0__0r2_35_0__2_), .Q(u3_u0_r2_2_));
DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_i_bF_buf61), .D(u3_u0__0r2_35_0__3_), .Q(u3_u0_r2_3_));
DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_i_bF_buf60), .D(u3_u0__0r2_35_0__4_), .Q(u3_u0_r2_4_));
DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_i_bF_buf59), .D(u3_u0__0r2_35_0__5_), .Q(u3_u0_r2_5_));
DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_i_bF_buf58), .D(u3_u0__0r2_35_0__6_), .Q(u3_u0_r2_6_));
DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_i_bF_buf57), .D(u3_u0__0r2_35_0__7_), .Q(u3_u0_r2_7_));
DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_i_bF_buf56), .D(u3_u0__0r2_35_0__8_), .Q(u3_u0_r2_8_));
DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_i_bF_buf55), .D(u3_u0__0r2_35_0__9_), .Q(u3_u0_r2_9_));
DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_i_bF_buf54), .D(u3_u0__0r2_35_0__10_), .Q(u3_u0_r2_10_));
DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_i_bF_buf53), .D(u3_u0__0r2_35_0__11_), .Q(u3_u0_r2_11_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_i_bF_buf19), .D(u0_u0__0tms_31_0__6_), .Q(u0_tms0_6_));
DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_i_bF_buf52), .D(u3_u0__0r2_35_0__12_), .Q(u3_u0_r2_12_));
DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_i_bF_buf51), .D(u3_u0__0r2_35_0__13_), .Q(u3_u0_r2_13_));
DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_i_bF_buf50), .D(u3_u0__0r2_35_0__14_), .Q(u3_u0_r2_14_));
DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_i_bF_buf49), .D(u3_u0__0r2_35_0__15_), .Q(u3_u0_r2_15_));
DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_i_bF_buf48), .D(u3_u0__0r2_35_0__16_), .Q(u3_u0_r2_16_));
DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_i_bF_buf47), .D(u3_u0__0r2_35_0__17_), .Q(u3_u0_r2_17_));
DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_i_bF_buf46), .D(u3_u0__0r2_35_0__18_), .Q(u3_u0_r2_18_));
DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_i_bF_buf45), .D(u3_u0__0r2_35_0__19_), .Q(u3_u0_r2_19_));
DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_i_bF_buf44), .D(u3_u0__0r2_35_0__20_), .Q(u3_u0_r2_20_));
DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_i_bF_buf43), .D(u3_u0__0r2_35_0__21_), .Q(u3_u0_r2_21_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_i_bF_buf18), .D(u0_u0__0tms_31_0__7_), .Q(u0_tms0_7_));
DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_i_bF_buf42), .D(u3_u0__0r2_35_0__22_), .Q(u3_u0_r2_22_));
DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_i_bF_buf41), .D(u3_u0__0r2_35_0__23_), .Q(u3_u0_r2_23_));
DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_i_bF_buf40), .D(u3_u0__0r2_35_0__24_), .Q(u3_u0_r2_24_));
DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_i_bF_buf39), .D(u3_u0__0r2_35_0__25_), .Q(u3_u0_r2_25_));
DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_i_bF_buf38), .D(u3_u0__0r2_35_0__26_), .Q(u3_u0_r2_26_));
DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_i_bF_buf37), .D(u3_u0__0r2_35_0__27_), .Q(u3_u0_r2_27_));
DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_i_bF_buf36), .D(u3_u0__0r2_35_0__28_), .Q(u3_u0_r2_28_));
DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_i_bF_buf35), .D(u3_u0__0r2_35_0__29_), .Q(u3_u0_r2_29_));
DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_i_bF_buf34), .D(u3_u0__0r2_35_0__30_), .Q(u3_u0_r2_30_));
DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_i_bF_buf33), .D(u3_u0__0r2_35_0__31_), .Q(u3_u0_r2_31_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_i_bF_buf92), .D(u0__0poc_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_85523_1_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_i_bF_buf17), .D(u0_u0__0tms_31_0__8_), .Q(u0_tms0_8_));
DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_i_bF_buf32), .D(u3_u0__0r2_35_0__32_), .Q(u3_u0_r2_32_));
DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_i_bF_buf31), .D(u3_u0__0r2_35_0__33_), .Q(u3_u0_r2_33_));
DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_i_bF_buf30), .D(u3_u0__0r2_35_0__34_), .Q(u3_u0_r2_34_));
DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_i_bF_buf29), .D(u3_u0__0r2_35_0__35_), .Q(u3_u0_r2_35_));
DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_i_bF_buf28), .D(u3_u0__0r1_35_0__0_), .Q(u3_u0_r1_0_));
DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_i_bF_buf27), .D(u3_u0__0r1_35_0__1_), .Q(u3_u0_r1_1_));
DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_i_bF_buf26), .D(u3_u0__0r1_35_0__2_), .Q(u3_u0_r1_2_));
DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_i_bF_buf25), .D(u3_u0__0r1_35_0__3_), .Q(u3_u0_r1_3_));
DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_i_bF_buf24), .D(u3_u0__0r1_35_0__4_), .Q(u3_u0_r1_4_));
DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_i_bF_buf23), .D(u3_u0__0r1_35_0__5_), .Q(u3_u0_r1_5_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_i_bF_buf16), .D(u0_u0__0tms_31_0__9_), .Q(u0_tms0_9_));
DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_i_bF_buf22), .D(u3_u0__0r1_35_0__6_), .Q(u3_u0_r1_6_));
DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_i_bF_buf21), .D(u3_u0__0r1_35_0__7_), .Q(u3_u0_r1_7_));
DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_i_bF_buf20), .D(u3_u0__0r1_35_0__8_), .Q(u3_u0_r1_8_));
DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_i_bF_buf19), .D(u3_u0__0r1_35_0__9_), .Q(u3_u0_r1_9_));
DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_i_bF_buf18), .D(u3_u0__0r1_35_0__10_), .Q(u3_u0_r1_10_));
DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_i_bF_buf17), .D(u3_u0__0r1_35_0__11_), .Q(u3_u0_r1_11_));
DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_i_bF_buf16), .D(u3_u0__0r1_35_0__12_), .Q(u3_u0_r1_12_));
DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_i_bF_buf15), .D(u3_u0__0r1_35_0__13_), .Q(u3_u0_r1_13_));
DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_i_bF_buf14), .D(u3_u0__0r1_35_0__14_), .Q(u3_u0_r1_14_));
DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_i_bF_buf13), .D(u3_u0__0r1_35_0__15_), .Q(u3_u0_r1_15_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_i_bF_buf15), .D(u0_u0__0tms_31_0__10_), .Q(u0_tms0_10_));
DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_i_bF_buf12), .D(u3_u0__0r1_35_0__16_), .Q(u3_u0_r1_16_));
DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_i_bF_buf11), .D(u3_u0__0r1_35_0__17_), .Q(u3_u0_r1_17_));
DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_i_bF_buf10), .D(u3_u0__0r1_35_0__18_), .Q(u3_u0_r1_18_));
DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_i_bF_buf9), .D(u3_u0__0r1_35_0__19_), .Q(u3_u0_r1_19_));
DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_i_bF_buf8), .D(u3_u0__0r1_35_0__20_), .Q(u3_u0_r1_20_));
DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_i_bF_buf7), .D(u3_u0__0r1_35_0__21_), .Q(u3_u0_r1_21_));
DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_i_bF_buf6), .D(u3_u0__0r1_35_0__22_), .Q(u3_u0_r1_22_));
DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_i_bF_buf5), .D(u3_u0__0r1_35_0__23_), .Q(u3_u0_r1_23_));
DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_i_bF_buf4), .D(u3_u0__0r1_35_0__24_), .Q(u3_u0_r1_24_));
DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_i_bF_buf3), .D(u3_u0__0r1_35_0__25_), .Q(u3_u0_r1_25_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_i_bF_buf14), .D(u0_u0__0tms_31_0__11_), .Q(u0_tms0_11_));
DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_i_bF_buf2), .D(u3_u0__0r1_35_0__26_), .Q(u3_u0_r1_26_));
DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_i_bF_buf1), .D(u3_u0__0r1_35_0__27_), .Q(u3_u0_r1_27_));
DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_i_bF_buf0), .D(u3_u0__0r1_35_0__28_), .Q(u3_u0_r1_28_));
DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_i_bF_buf96), .D(u3_u0__0r1_35_0__29_), .Q(u3_u0_r1_29_));
DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_i_bF_buf95), .D(u3_u0__0r1_35_0__30_), .Q(u3_u0_r1_30_));
DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_i_bF_buf94), .D(u3_u0__0r1_35_0__31_), .Q(u3_u0_r1_31_));
DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_i_bF_buf93), .D(u3_u0__0r1_35_0__32_), .Q(u3_u0_r1_32_));
DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_i_bF_buf92), .D(u3_u0__0r1_35_0__33_), .Q(u3_u0_r1_33_));
DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_i_bF_buf91), .D(u3_u0__0r1_35_0__34_), .Q(u3_u0_r1_34_));
DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_i_bF_buf90), .D(u3_u0__0r1_35_0__35_), .Q(u3_u0_r1_35_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_i_bF_buf13), .D(u0_u0__0tms_31_0__12_), .Q(u0_tms0_12_));
DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_i_bF_buf89), .D(u3_u0__0r0_35_0__0_), .Q(u3_u0_r0_0_));
DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_i_bF_buf88), .D(u3_u0__0r0_35_0__1_), .Q(u3_u0_r0_1_));
DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_i_bF_buf87), .D(u3_u0__0r0_35_0__2_), .Q(u3_u0_r0_2_));
DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_i_bF_buf86), .D(u3_u0__0r0_35_0__3_), .Q(u3_u0_r0_3_));
DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_i_bF_buf85), .D(u3_u0__0r0_35_0__4_), .Q(u3_u0_r0_4_));
DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_i_bF_buf84), .D(u3_u0__0r0_35_0__5_), .Q(u3_u0_r0_5_));
DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_i_bF_buf83), .D(u3_u0__0r0_35_0__6_), .Q(u3_u0_r0_6_));
DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_i_bF_buf82), .D(u3_u0__0r0_35_0__7_), .Q(u3_u0_r0_7_));
DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_i_bF_buf81), .D(u3_u0__0r0_35_0__8_), .Q(u3_u0_r0_8_));
DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_i_bF_buf80), .D(u3_u0__0r0_35_0__9_), .Q(u3_u0_r0_9_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_i_bF_buf12), .D(u0_u0__0tms_31_0__13_), .Q(u0_tms0_13_));
DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_i_bF_buf79), .D(u3_u0__0r0_35_0__10_), .Q(u3_u0_r0_10_));
DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_i_bF_buf78), .D(u3_u0__0r0_35_0__11_), .Q(u3_u0_r0_11_));
DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_i_bF_buf77), .D(u3_u0__0r0_35_0__12_), .Q(u3_u0_r0_12_));
DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_i_bF_buf76), .D(u3_u0__0r0_35_0__13_), .Q(u3_u0_r0_13_));
DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_i_bF_buf75), .D(u3_u0__0r0_35_0__14_), .Q(u3_u0_r0_14_));
DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_i_bF_buf74), .D(u3_u0__0r0_35_0__15_), .Q(u3_u0_r0_15_));
DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_i_bF_buf73), .D(u3_u0__0r0_35_0__16_), .Q(u3_u0_r0_16_));
DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_i_bF_buf72), .D(u3_u0__0r0_35_0__17_), .Q(u3_u0_r0_17_));
DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_i_bF_buf71), .D(u3_u0__0r0_35_0__18_), .Q(u3_u0_r0_18_));
DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_i_bF_buf70), .D(u3_u0__0r0_35_0__19_), .Q(u3_u0_r0_19_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_i_bF_buf11), .D(u0_u0__0tms_31_0__14_), .Q(u0_tms0_14_));
DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_i_bF_buf69), .D(u3_u0__0r0_35_0__20_), .Q(u3_u0_r0_20_));
DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_i_bF_buf68), .D(u3_u0__0r0_35_0__21_), .Q(u3_u0_r0_21_));
DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_i_bF_buf67), .D(u3_u0__0r0_35_0__22_), .Q(u3_u0_r0_22_));
DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_i_bF_buf66), .D(u3_u0__0r0_35_0__23_), .Q(u3_u0_r0_23_));
DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_i_bF_buf65), .D(u3_u0__0r0_35_0__24_), .Q(u3_u0_r0_24_));
DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_i_bF_buf64), .D(u3_u0__0r0_35_0__25_), .Q(u3_u0_r0_25_));
DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_i_bF_buf63), .D(u3_u0__0r0_35_0__26_), .Q(u3_u0_r0_26_));
DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_i_bF_buf62), .D(u3_u0__0r0_35_0__27_), .Q(u3_u0_r0_27_));
DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_i_bF_buf61), .D(u3_u0__0r0_35_0__28_), .Q(u3_u0_r0_28_));
DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_i_bF_buf60), .D(u3_u0__0r0_35_0__29_), .Q(u3_u0_r0_29_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_i_bF_buf10), .D(u0_u0__0tms_31_0__15_), .Q(u0_tms0_15_));
DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_i_bF_buf59), .D(u3_u0__0r0_35_0__30_), .Q(u3_u0_r0_30_));
DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_i_bF_buf58), .D(u3_u0__0r0_35_0__31_), .Q(u3_u0_r0_31_));
DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_i_bF_buf57), .D(u3_u0__0r0_35_0__32_), .Q(u3_u0_r0_32_));
DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_i_bF_buf56), .D(u3_u0__0r0_35_0__33_), .Q(u3_u0_r0_33_));
DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_i_bF_buf55), .D(u3_u0__0r0_35_0__34_), .Q(u3_u0_r0_34_));
DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_i_bF_buf54), .D(u3_u0__0r0_35_0__35_), .Q(u3_u0_r0_35_));
DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_i_bF_buf45), .D(u4__0rfr_clr_0_0_), .Q(u4_rfr_clr));
DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_i_bF_buf24), .D(u1_wb_write_go), .Q(u5_wb_write_go_r));
DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_i_bF_buf23), .D(cmd_a10), .Q(u5_cmd_a10_r));
DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_i_bF_buf22), .D(u5__0burst_act_rd_0_0_), .Q(u5_burst_act_rd));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_i_bF_buf9), .D(u0_u0__0tms_31_0__16_), .Q(u0_tms0_16_));
DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_i_bF_buf21), .D(u5__0burst_cnt_10_0__0_), .Q(u5_burst_cnt_0_));
DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_i_bF_buf20), .D(u5__0burst_cnt_10_0__1_), .Q(u5_burst_cnt_1_));
DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_i_bF_buf19), .D(u5__0burst_cnt_10_0__2_), .Q(u5_burst_cnt_2_));
DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_i_bF_buf18), .D(u5__0burst_cnt_10_0__3_), .Q(u5_burst_cnt_3_));
DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_i_bF_buf17), .D(u5__0burst_cnt_10_0__4_), .Q(u5_burst_cnt_4_));
DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_i_bF_buf16), .D(u5__0burst_cnt_10_0__5_), .Q(u5_burst_cnt_5_));
DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_i_bF_buf15), .D(u5__0burst_cnt_10_0__6_), .Q(u5_burst_cnt_6_));
DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_i_bF_buf14), .D(u5__0burst_cnt_10_0__7_), .Q(u5_burst_cnt_7_));
DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_i_bF_buf13), .D(u5__0burst_cnt_10_0__8_), .Q(u5_burst_cnt_8_));
DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_i_bF_buf12), .D(u5__0burst_cnt_10_0__9_), .Q(u5_burst_cnt_9_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_i_bF_buf8), .D(u0_u0__0tms_31_0__17_), .Q(u0_tms0_17_));
DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_i_bF_buf11), .D(u5__0burst_cnt_10_0__10_), .Q(u5_burst_cnt_10_));
DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_i_bF_buf10), .D(u5__0ir_cnt_done_0_0_), .Q(u5_ir_cnt_done));
DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_i_bF_buf9), .D(u5__0ir_cnt_3_0__0_), .Q(u5_ir_cnt_0_));
DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_i_bF_buf8), .D(u5__0ir_cnt_3_0__1_), .Q(u5_ir_cnt_1_));
DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_i_bF_buf7), .D(u5__0ir_cnt_3_0__2_), .Q(u5_ir_cnt_2_));
DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_i_bF_buf6), .D(u5__0ir_cnt_3_0__3_), .Q(u5_ir_cnt_3_));
DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_i_bF_buf5), .D(u5__0timer2_8_0__0_), .Q(u5_timer2_0_));
DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_i_bF_buf4), .D(u5__0timer2_8_0__1_), .Q(u5_timer2_1_));
DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_i_bF_buf3), .D(u5__0timer2_8_0__2_), .Q(u5_timer2_2_));
DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_i_bF_buf2), .D(u5__0timer2_8_0__3_), .Q(u5_timer2_3_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_i_bF_buf91), .D(u0__0poc_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_85523_2_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_i_bF_buf7), .D(u0_u0__0tms_31_0__18_), .Q(u0_tms0_18_));
DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_i_bF_buf1), .D(u5__0timer2_8_0__4_), .Q(u5_timer2_4_));
DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_i_bF_buf0), .D(u5__0timer2_8_0__5_), .Q(u5_timer2_5_));
DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_i_bF_buf96), .D(u5__0timer2_8_0__6_), .Q(u5_timer2_6_));
DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_i_bF_buf95), .D(u5__0timer2_8_0__7_), .Q(u5_timer2_7_));
DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_i_bF_buf94), .D(u5__0timer2_8_0__8_), .Q(u5_timer2_8_));
DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_i_bF_buf93), .D(u5_cnt_next), .Q(u5_cnt));
DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_i_bF_buf92), .D(u5_wb_wait_r2), .Q(u5_wb_wait_r));
DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_i_bF_buf91), .D(u5_wb_wait), .Q(u5_wb_wait_r2));
DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_i_bF_buf90), .D(u5_cke_o_r2), .Q(u5_cke_o_del));
DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_i_bF_buf89), .D(u5_cke_o_r1), .Q(u5_cke_o_r2));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_i_bF_buf6), .D(u0_u0__0tms_31_0__19_), .Q(u0_tms0_19_));
DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_i_bF_buf88), .D(_auto_iopadmap_cc_368_execute_85453), .Q(u5_cke_o_r1));
DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_i_bF_buf87), .D(u5__0cke__0_0_), .Q(_auto_iopadmap_cc_368_execute_85453));
DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_i_bF_buf86), .D(u5_cke_d), .Q(u5_cke_r));
DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_i_bF_buf85), .D(u5_pack_le2_d), .Q(pack_le2));
DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_i_bF_buf84), .D(u5_pack_le1_d), .Q(pack_le1));
DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_i_bF_buf83), .D(u5_pack_le0_d), .Q(pack_le0));
DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_i_bF_buf82), .D(cs_le_d), .Q(cs_le));
DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_i_bF_buf81), .D(cs_le_bF_buf1), .Q(u5_cs_le_r1));
DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_i_bF_buf80), .D(u5_cs_le_r1), .Q(u5_cs_le_r));
DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_i_bF_buf79), .D(u5_lmr_ack_d), .Q(lmr_ack));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_i_bF_buf5), .D(u0_u0__0tms_31_0__20_), .Q(u0_tms0_20_));
DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_i_bF_buf62), .D(u6__0wb_data_o_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_85560_0_));
DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_i_bF_buf61), .D(u6__0wb_data_o_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_85560_1_));
DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_i_bF_buf60), .D(u6__0wb_data_o_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_85560_2_));
DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_i_bF_buf59), .D(u6__0wb_data_o_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_85560_3_));
DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_i_bF_buf58), .D(u6__0wb_data_o_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_85560_4_));
DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_i_bF_buf57), .D(u6__0wb_data_o_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_85560_5_));
DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_i_bF_buf56), .D(u6__0wb_data_o_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_85560_6_));
DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_i_bF_buf55), .D(u6__0wb_data_o_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_85560_7_));
DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_i_bF_buf54), .D(u6__0wb_data_o_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_85560_8_));
DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_i_bF_buf53), .D(u6__0wb_data_o_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_85560_9_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_i_bF_buf4), .D(u0_u0__0tms_31_0__21_), .Q(u0_tms0_21_));
DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_i_bF_buf52), .D(u6__0wb_data_o_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_85560_10_));
DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_i_bF_buf51), .D(u6__0wb_data_o_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_85560_11_));
DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_i_bF_buf50), .D(u6__0wb_data_o_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_85560_12_));
DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_i_bF_buf49), .D(u6__0wb_data_o_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_85560_13_));
DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_i_bF_buf48), .D(u6__0wb_data_o_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_85560_14_));
DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_i_bF_buf47), .D(u6__0wb_data_o_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_85560_15_));
DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_i_bF_buf46), .D(u6__0wb_data_o_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_85560_16_));
DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_i_bF_buf45), .D(u6__0wb_data_o_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_85560_17_));
DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_i_bF_buf44), .D(u6__0wb_data_o_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_85560_18_));
DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_i_bF_buf43), .D(u6__0wb_data_o_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_85560_19_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_i_bF_buf3), .D(u0_u0__0tms_31_0__22_), .Q(u0_tms0_22_));
DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_i_bF_buf42), .D(u6__0wb_data_o_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_85560_20_));
DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_i_bF_buf41), .D(u6__0wb_data_o_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_85560_21_));
DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_i_bF_buf40), .D(u6__0wb_data_o_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_85560_22_));
DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_i_bF_buf39), .D(u6__0wb_data_o_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_85560_23_));
DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_i_bF_buf38), .D(u6__0wb_data_o_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_85560_24_));
DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_i_bF_buf37), .D(u6__0wb_data_o_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_85560_25_));
DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_i_bF_buf36), .D(u6__0wb_data_o_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_85560_26_));
DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_i_bF_buf35), .D(u6__0wb_data_o_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_85560_27_));
DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_i_bF_buf34), .D(u6__0wb_data_o_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_85560_28_));
DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_i_bF_buf33), .D(u6__0wb_data_o_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_85560_29_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_i_bF_buf2), .D(u0_u0__0tms_31_0__23_), .Q(u0_tms0_23_));
DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_i_bF_buf32), .D(u6__0wb_data_o_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_85560_30_));
DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_i_bF_buf31), .D(u6__0wb_data_o_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_85560_31_));
DFFPOSX1 DFFPOSX1_652 ( .CLK(mc_clk_i_bF_buf10), .D(u7__0mc_adv__0_0_), .Q(_auto_iopadmap_cc_368_execute_85447));
DFFPOSX1 DFFPOSX1_653 ( .CLK(mc_clk_i_bF_buf9), .D(u7__0mc_adsc__0_0_), .Q(_auto_iopadmap_cc_368_execute_85445));
DFFPOSX1 DFFPOSX1_654 ( .CLK(mc_clk_i_bF_buf8), .D(ras_), .Q(_auto_iopadmap_cc_368_execute_85513));
DFFPOSX1 DFFPOSX1_655 ( .CLK(mc_clk_i_bF_buf7), .D(cas_), .Q(_auto_iopadmap_cc_368_execute_85451));
DFFPOSX1 DFFPOSX1_656 ( .CLK(mc_clk_i_bF_buf6), .D(u5_we_), .Q(_auto_iopadmap_cc_368_execute_85519));
DFFPOSX1 DFFPOSX1_657 ( .CLK(mc_clk_i_bF_buf5), .D(u7__0mc_dqm_3_0__0_), .Q(_auto_iopadmap_cc_368_execute_85506_0_));
DFFPOSX1 DFFPOSX1_658 ( .CLK(mc_clk_i_bF_buf4), .D(u7__0mc_dqm_3_0__1_), .Q(_auto_iopadmap_cc_368_execute_85506_1_));
DFFPOSX1 DFFPOSX1_659 ( .CLK(mc_clk_i_bF_buf3), .D(u7__0mc_dqm_3_0__2_), .Q(_auto_iopadmap_cc_368_execute_85506_2_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_i_bF_buf1), .D(u0_u0__0tms_31_0__24_), .Q(u0_tms0_24_));
DFFPOSX1 DFFPOSX1_660 ( .CLK(mc_clk_i_bF_buf2), .D(u7__0mc_dqm_3_0__3_), .Q(_auto_iopadmap_cc_368_execute_85506_3_));
DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_i_bF_buf20), .D(u7_mc_dqm_r_0_), .Q(u7_mc_dqm_r2_0_));
DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_i_bF_buf19), .D(u7_mc_dqm_r_1_), .Q(u7_mc_dqm_r2_1_));
DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_i_bF_buf18), .D(u7_mc_dqm_r_2_), .Q(u7_mc_dqm_r2_2_));
DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_i_bF_buf17), .D(u7_mc_dqm_r_3_), .Q(u7_mc_dqm_r2_3_));
DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_i_bF_buf16), .D(u7__0mc_dqm_r_3_0__0_), .Q(u7_mc_dqm_r_0_));
DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_i_bF_buf15), .D(u7__0mc_dqm_r_3_0__1_), .Q(u7_mc_dqm_r_1_));
DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_i_bF_buf14), .D(u7__0mc_dqm_r_3_0__2_), .Q(u7_mc_dqm_r_2_));
DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_i_bF_buf13), .D(u7__0mc_dqm_r_3_0__3_), .Q(u7_mc_dqm_r_3_));
DFFPOSX1 DFFPOSX1_669 ( .CLK(mc_clk_i_bF_buf1), .D(mc_addr_d_0_), .Q(_auto_iopadmap_cc_368_execute_85420_0_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_i_bF_buf0), .D(u0_u0__0tms_31_0__25_), .Q(u0_tms0_25_));
DFFPOSX1 DFFPOSX1_670 ( .CLK(mc_clk_i_bF_buf0), .D(mc_addr_d_1_), .Q(_auto_iopadmap_cc_368_execute_85420_1_));
DFFPOSX1 DFFPOSX1_671 ( .CLK(mc_clk_i_bF_buf10), .D(mc_addr_d_2_), .Q(_auto_iopadmap_cc_368_execute_85420_2_));
DFFPOSX1 DFFPOSX1_672 ( .CLK(mc_clk_i_bF_buf9), .D(mc_addr_d_3_), .Q(_auto_iopadmap_cc_368_execute_85420_3_));
DFFPOSX1 DFFPOSX1_673 ( .CLK(mc_clk_i_bF_buf8), .D(mc_addr_d_4_), .Q(_auto_iopadmap_cc_368_execute_85420_4_));
DFFPOSX1 DFFPOSX1_674 ( .CLK(mc_clk_i_bF_buf7), .D(mc_addr_d_5_), .Q(_auto_iopadmap_cc_368_execute_85420_5_));
DFFPOSX1 DFFPOSX1_675 ( .CLK(mc_clk_i_bF_buf6), .D(mc_addr_d_6_), .Q(_auto_iopadmap_cc_368_execute_85420_6_));
DFFPOSX1 DFFPOSX1_676 ( .CLK(mc_clk_i_bF_buf5), .D(mc_addr_d_7_), .Q(_auto_iopadmap_cc_368_execute_85420_7_));
DFFPOSX1 DFFPOSX1_677 ( .CLK(mc_clk_i_bF_buf4), .D(mc_addr_d_8_), .Q(_auto_iopadmap_cc_368_execute_85420_8_));
DFFPOSX1 DFFPOSX1_678 ( .CLK(mc_clk_i_bF_buf3), .D(mc_addr_d_9_), .Q(_auto_iopadmap_cc_368_execute_85420_9_));
DFFPOSX1 DFFPOSX1_679 ( .CLK(mc_clk_i_bF_buf2), .D(mc_addr_d_10_), .Q(_auto_iopadmap_cc_368_execute_85420_10_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_i_bF_buf96), .D(u0_u0__0tms_31_0__26_), .Q(u0_tms0_26_));
DFFPOSX1 DFFPOSX1_680 ( .CLK(mc_clk_i_bF_buf1), .D(mc_addr_d_11_), .Q(_auto_iopadmap_cc_368_execute_85420_11_));
DFFPOSX1 DFFPOSX1_681 ( .CLK(mc_clk_i_bF_buf0), .D(mc_addr_d_12_), .Q(_auto_iopadmap_cc_368_execute_85420_12_));
DFFPOSX1 DFFPOSX1_682 ( .CLK(mc_clk_i_bF_buf10), .D(mc_addr_d_13_), .Q(_auto_iopadmap_cc_368_execute_85420_13_));
DFFPOSX1 DFFPOSX1_683 ( .CLK(mc_clk_i_bF_buf9), .D(mc_addr_d_14_), .Q(_auto_iopadmap_cc_368_execute_85420_14_));
DFFPOSX1 DFFPOSX1_684 ( .CLK(mc_clk_i_bF_buf8), .D(mc_addr_d_15_), .Q(_auto_iopadmap_cc_368_execute_85420_15_));
DFFPOSX1 DFFPOSX1_685 ( .CLK(mc_clk_i_bF_buf7), .D(mc_addr_d_16_), .Q(_auto_iopadmap_cc_368_execute_85420_16_));
DFFPOSX1 DFFPOSX1_686 ( .CLK(mc_clk_i_bF_buf6), .D(mc_addr_d_17_), .Q(_auto_iopadmap_cc_368_execute_85420_17_));
DFFPOSX1 DFFPOSX1_687 ( .CLK(mc_clk_i_bF_buf5), .D(mc_addr_d_18_), .Q(_auto_iopadmap_cc_368_execute_85420_18_));
DFFPOSX1 DFFPOSX1_688 ( .CLK(mc_clk_i_bF_buf4), .D(mc_addr_d_19_), .Q(_auto_iopadmap_cc_368_execute_85420_19_));
DFFPOSX1 DFFPOSX1_689 ( .CLK(mc_clk_i_bF_buf3), .D(mc_addr_d_20_), .Q(_auto_iopadmap_cc_368_execute_85420_20_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_i_bF_buf95), .D(u0_u0__0tms_31_0__27_), .Q(u0_tms0_27_));
DFFPOSX1 DFFPOSX1_690 ( .CLK(mc_clk_i_bF_buf2), .D(mc_addr_d_21_), .Q(_auto_iopadmap_cc_368_execute_85420_21_));
DFFPOSX1 DFFPOSX1_691 ( .CLK(mc_clk_i_bF_buf1), .D(mc_addr_d_22_), .Q(_auto_iopadmap_cc_368_execute_85420_22_));
DFFPOSX1 DFFPOSX1_692 ( .CLK(mc_clk_i_bF_buf0), .D(mc_addr_d_23_), .Q(_auto_iopadmap_cc_368_execute_85420_23_));
DFFPOSX1 DFFPOSX1_693 ( .CLK(mc_clk_i_bF_buf10), .D(mc_dp_od_0_), .Q(_auto_iopadmap_cc_368_execute_85501_0_));
DFFPOSX1 DFFPOSX1_694 ( .CLK(mc_clk_i_bF_buf9), .D(mc_dp_od_1_), .Q(_auto_iopadmap_cc_368_execute_85501_1_));
DFFPOSX1 DFFPOSX1_695 ( .CLK(mc_clk_i_bF_buf8), .D(mc_dp_od_2_), .Q(_auto_iopadmap_cc_368_execute_85501_2_));
DFFPOSX1 DFFPOSX1_696 ( .CLK(mc_clk_i_bF_buf7), .D(mc_dp_od_3_), .Q(_auto_iopadmap_cc_368_execute_85501_3_));
DFFPOSX1 DFFPOSX1_697 ( .CLK(mc_clk_i_bF_buf6), .D(mc_data_od_0_), .Q(_auto_iopadmap_cc_368_execute_85466_0_));
DFFPOSX1 DFFPOSX1_698 ( .CLK(mc_clk_i_bF_buf5), .D(mc_data_od_1_), .Q(_auto_iopadmap_cc_368_execute_85466_1_));
DFFPOSX1 DFFPOSX1_699 ( .CLK(mc_clk_i_bF_buf4), .D(mc_data_od_2_), .Q(_auto_iopadmap_cc_368_execute_85466_2_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_i_bF_buf90), .D(u0__0poc_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_85523_3_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_i_bF_buf94), .D(u0_u0__0tms_31_0__28_), .Q(u0_tms0_28_));
DFFPOSX1 DFFPOSX1_700 ( .CLK(mc_clk_i_bF_buf3), .D(mc_data_od_3_), .Q(_auto_iopadmap_cc_368_execute_85466_3_));
DFFPOSX1 DFFPOSX1_701 ( .CLK(mc_clk_i_bF_buf2), .D(mc_data_od_4_), .Q(_auto_iopadmap_cc_368_execute_85466_4_));
DFFPOSX1 DFFPOSX1_702 ( .CLK(mc_clk_i_bF_buf1), .D(mc_data_od_5_), .Q(_auto_iopadmap_cc_368_execute_85466_5_));
DFFPOSX1 DFFPOSX1_703 ( .CLK(mc_clk_i_bF_buf0), .D(mc_data_od_6_), .Q(_auto_iopadmap_cc_368_execute_85466_6_));
DFFPOSX1 DFFPOSX1_704 ( .CLK(mc_clk_i_bF_buf10), .D(mc_data_od_7_), .Q(_auto_iopadmap_cc_368_execute_85466_7_));
DFFPOSX1 DFFPOSX1_705 ( .CLK(mc_clk_i_bF_buf9), .D(mc_data_od_8_), .Q(_auto_iopadmap_cc_368_execute_85466_8_));
DFFPOSX1 DFFPOSX1_706 ( .CLK(mc_clk_i_bF_buf8), .D(mc_data_od_9_), .Q(_auto_iopadmap_cc_368_execute_85466_9_));
DFFPOSX1 DFFPOSX1_707 ( .CLK(mc_clk_i_bF_buf7), .D(mc_data_od_10_), .Q(_auto_iopadmap_cc_368_execute_85466_10_));
DFFPOSX1 DFFPOSX1_708 ( .CLK(mc_clk_i_bF_buf6), .D(mc_data_od_11_), .Q(_auto_iopadmap_cc_368_execute_85466_11_));
DFFPOSX1 DFFPOSX1_709 ( .CLK(mc_clk_i_bF_buf5), .D(mc_data_od_12_), .Q(_auto_iopadmap_cc_368_execute_85466_12_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_i_bF_buf93), .D(u0_u0__0tms_31_0__29_), .Q(u0_tms0_29_));
DFFPOSX1 DFFPOSX1_710 ( .CLK(mc_clk_i_bF_buf4), .D(mc_data_od_13_), .Q(_auto_iopadmap_cc_368_execute_85466_13_));
DFFPOSX1 DFFPOSX1_711 ( .CLK(mc_clk_i_bF_buf3), .D(mc_data_od_14_), .Q(_auto_iopadmap_cc_368_execute_85466_14_));
DFFPOSX1 DFFPOSX1_712 ( .CLK(mc_clk_i_bF_buf2), .D(mc_data_od_15_), .Q(_auto_iopadmap_cc_368_execute_85466_15_));
DFFPOSX1 DFFPOSX1_713 ( .CLK(mc_clk_i_bF_buf1), .D(mc_data_od_16_), .Q(_auto_iopadmap_cc_368_execute_85466_16_));
DFFPOSX1 DFFPOSX1_714 ( .CLK(mc_clk_i_bF_buf0), .D(mc_data_od_17_), .Q(_auto_iopadmap_cc_368_execute_85466_17_));
DFFPOSX1 DFFPOSX1_715 ( .CLK(mc_clk_i_bF_buf10), .D(mc_data_od_18_), .Q(_auto_iopadmap_cc_368_execute_85466_18_));
DFFPOSX1 DFFPOSX1_716 ( .CLK(mc_clk_i_bF_buf9), .D(mc_data_od_19_), .Q(_auto_iopadmap_cc_368_execute_85466_19_));
DFFPOSX1 DFFPOSX1_717 ( .CLK(mc_clk_i_bF_buf8), .D(mc_data_od_20_), .Q(_auto_iopadmap_cc_368_execute_85466_20_));
DFFPOSX1 DFFPOSX1_718 ( .CLK(mc_clk_i_bF_buf7), .D(mc_data_od_21_), .Q(_auto_iopadmap_cc_368_execute_85466_21_));
DFFPOSX1 DFFPOSX1_719 ( .CLK(mc_clk_i_bF_buf6), .D(mc_data_od_22_), .Q(_auto_iopadmap_cc_368_execute_85466_22_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_i_bF_buf92), .D(u0_u0__0tms_31_0__30_), .Q(u0_tms0_30_));
DFFPOSX1 DFFPOSX1_720 ( .CLK(mc_clk_i_bF_buf5), .D(mc_data_od_23_), .Q(_auto_iopadmap_cc_368_execute_85466_23_));
DFFPOSX1 DFFPOSX1_721 ( .CLK(mc_clk_i_bF_buf4), .D(mc_data_od_24_), .Q(_auto_iopadmap_cc_368_execute_85466_24_));
DFFPOSX1 DFFPOSX1_722 ( .CLK(mc_clk_i_bF_buf3), .D(mc_data_od_25_), .Q(_auto_iopadmap_cc_368_execute_85466_25_));
DFFPOSX1 DFFPOSX1_723 ( .CLK(mc_clk_i_bF_buf2), .D(mc_data_od_26_), .Q(_auto_iopadmap_cc_368_execute_85466_26_));
DFFPOSX1 DFFPOSX1_724 ( .CLK(mc_clk_i_bF_buf1), .D(mc_data_od_27_), .Q(_auto_iopadmap_cc_368_execute_85466_27_));
DFFPOSX1 DFFPOSX1_725 ( .CLK(mc_clk_i_bF_buf0), .D(mc_data_od_28_), .Q(_auto_iopadmap_cc_368_execute_85466_28_));
DFFPOSX1 DFFPOSX1_726 ( .CLK(mc_clk_i_bF_buf10), .D(mc_data_od_29_), .Q(_auto_iopadmap_cc_368_execute_85466_29_));
DFFPOSX1 DFFPOSX1_727 ( .CLK(mc_clk_i_bF_buf9), .D(mc_data_od_30_), .Q(_auto_iopadmap_cc_368_execute_85466_30_));
DFFPOSX1 DFFPOSX1_728 ( .CLK(mc_clk_i_bF_buf8), .D(mc_data_od_31_), .Q(_auto_iopadmap_cc_368_execute_85466_31_));
DFFPOSX1 DFFPOSX1_729 ( .CLK(mc_clk_i_bF_buf7), .D(mc_bg_d), .Q(_auto_iopadmap_cc_368_execute_85449));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_i_bF_buf91), .D(u0_u0__0tms_31_0__31_), .Q(u0_tms0_31_));
DFFPOSX1 DFFPOSX1_730 ( .CLK(mc_clk_i_bF_buf6), .D(mc_ack_pad_i), .Q(mc_ack_r));
DFFPOSX1 DFFPOSX1_731 ( .CLK(mc_clk_i_bF_buf5), .D(mc_br_pad_i), .Q(mc_br_r));
DFFPOSX1 DFFPOSX1_732 ( .CLK(mc_clk_i_bF_buf4), .D(u7__0mc_rp_0_0_), .Q(_auto_iopadmap_cc_368_execute_85515));
DFFPOSX1 DFFPOSX1_733 ( .CLK(mc_clk_i_bF_buf3), .D(mc_c_oe_d), .Q(_auto_iopadmap_cc_368_execute_85455));
DFFPOSX1 DFFPOSX1_734 ( .CLK(mc_clk_i_bF_buf2), .D(\mc_data_pad_i[0] ), .Q(mc_data_ir_0_));
DFFPOSX1 DFFPOSX1_735 ( .CLK(mc_clk_i_bF_buf1), .D(\mc_data_pad_i[1] ), .Q(mc_data_ir_1_));
DFFPOSX1 DFFPOSX1_736 ( .CLK(mc_clk_i_bF_buf0), .D(\mc_data_pad_i[2] ), .Q(mc_data_ir_2_));
DFFPOSX1 DFFPOSX1_737 ( .CLK(mc_clk_i_bF_buf10), .D(\mc_data_pad_i[3] ), .Q(mc_data_ir_3_));
DFFPOSX1 DFFPOSX1_738 ( .CLK(mc_clk_i_bF_buf9), .D(\mc_data_pad_i[4] ), .Q(mc_data_ir_4_));
DFFPOSX1 DFFPOSX1_739 ( .CLK(mc_clk_i_bF_buf8), .D(\mc_data_pad_i[5] ), .Q(mc_data_ir_5_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_i_bF_buf90), .D(u0_u0__0csc_31_0__0_), .Q(u0_csc0_0_));
DFFPOSX1 DFFPOSX1_740 ( .CLK(mc_clk_i_bF_buf7), .D(\mc_data_pad_i[6] ), .Q(mc_data_ir_6_));
DFFPOSX1 DFFPOSX1_741 ( .CLK(mc_clk_i_bF_buf6), .D(\mc_data_pad_i[7] ), .Q(mc_data_ir_7_));
DFFPOSX1 DFFPOSX1_742 ( .CLK(mc_clk_i_bF_buf5), .D(\mc_data_pad_i[8] ), .Q(mc_data_ir_8_));
DFFPOSX1 DFFPOSX1_743 ( .CLK(mc_clk_i_bF_buf4), .D(\mc_data_pad_i[9] ), .Q(mc_data_ir_9_));
DFFPOSX1 DFFPOSX1_744 ( .CLK(mc_clk_i_bF_buf3), .D(\mc_data_pad_i[10] ), .Q(mc_data_ir_10_));
DFFPOSX1 DFFPOSX1_745 ( .CLK(mc_clk_i_bF_buf2), .D(\mc_data_pad_i[11] ), .Q(mc_data_ir_11_));
DFFPOSX1 DFFPOSX1_746 ( .CLK(mc_clk_i_bF_buf1), .D(\mc_data_pad_i[12] ), .Q(mc_data_ir_12_));
DFFPOSX1 DFFPOSX1_747 ( .CLK(mc_clk_i_bF_buf0), .D(\mc_data_pad_i[13] ), .Q(mc_data_ir_13_));
DFFPOSX1 DFFPOSX1_748 ( .CLK(mc_clk_i_bF_buf10), .D(\mc_data_pad_i[14] ), .Q(mc_data_ir_14_));
DFFPOSX1 DFFPOSX1_749 ( .CLK(mc_clk_i_bF_buf9), .D(\mc_data_pad_i[15] ), .Q(mc_data_ir_15_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_i_bF_buf89), .D(u0_u0__0csc_31_0__1_), .Q(u0_csc0_1_));
DFFPOSX1 DFFPOSX1_750 ( .CLK(mc_clk_i_bF_buf8), .D(\mc_data_pad_i[16] ), .Q(mc_data_ir_16_));
DFFPOSX1 DFFPOSX1_751 ( .CLK(mc_clk_i_bF_buf7), .D(\mc_data_pad_i[17] ), .Q(mc_data_ir_17_));
DFFPOSX1 DFFPOSX1_752 ( .CLK(mc_clk_i_bF_buf6), .D(\mc_data_pad_i[18] ), .Q(mc_data_ir_18_));
DFFPOSX1 DFFPOSX1_753 ( .CLK(mc_clk_i_bF_buf5), .D(\mc_data_pad_i[19] ), .Q(mc_data_ir_19_));
DFFPOSX1 DFFPOSX1_754 ( .CLK(mc_clk_i_bF_buf4), .D(\mc_data_pad_i[20] ), .Q(mc_data_ir_20_));
DFFPOSX1 DFFPOSX1_755 ( .CLK(mc_clk_i_bF_buf3), .D(\mc_data_pad_i[21] ), .Q(mc_data_ir_21_));
DFFPOSX1 DFFPOSX1_756 ( .CLK(mc_clk_i_bF_buf2), .D(\mc_data_pad_i[22] ), .Q(mc_data_ir_22_));
DFFPOSX1 DFFPOSX1_757 ( .CLK(mc_clk_i_bF_buf1), .D(\mc_data_pad_i[23] ), .Q(mc_data_ir_23_));
DFFPOSX1 DFFPOSX1_758 ( .CLK(mc_clk_i_bF_buf0), .D(\mc_data_pad_i[24] ), .Q(mc_data_ir_24_));
DFFPOSX1 DFFPOSX1_759 ( .CLK(mc_clk_i_bF_buf10), .D(\mc_data_pad_i[25] ), .Q(mc_data_ir_25_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_i_bF_buf88), .D(u0_u0__0csc_31_0__2_), .Q(u0_csc0_2_));
DFFPOSX1 DFFPOSX1_760 ( .CLK(mc_clk_i_bF_buf9), .D(\mc_data_pad_i[26] ), .Q(mc_data_ir_26_));
DFFPOSX1 DFFPOSX1_761 ( .CLK(mc_clk_i_bF_buf8), .D(\mc_data_pad_i[27] ), .Q(mc_data_ir_27_));
DFFPOSX1 DFFPOSX1_762 ( .CLK(mc_clk_i_bF_buf7), .D(\mc_data_pad_i[28] ), .Q(mc_data_ir_28_));
DFFPOSX1 DFFPOSX1_763 ( .CLK(mc_clk_i_bF_buf6), .D(\mc_data_pad_i[29] ), .Q(mc_data_ir_29_));
DFFPOSX1 DFFPOSX1_764 ( .CLK(mc_clk_i_bF_buf5), .D(\mc_data_pad_i[30] ), .Q(mc_data_ir_30_));
DFFPOSX1 DFFPOSX1_765 ( .CLK(mc_clk_i_bF_buf4), .D(\mc_data_pad_i[31] ), .Q(mc_data_ir_31_));
DFFPOSX1 DFFPOSX1_766 ( .CLK(mc_clk_i_bF_buf3), .D(\mc_dp_pad_i[0] ), .Q(mc_data_ir_32_));
DFFPOSX1 DFFPOSX1_767 ( .CLK(mc_clk_i_bF_buf2), .D(\mc_dp_pad_i[1] ), .Q(mc_data_ir_33_));
DFFPOSX1 DFFPOSX1_768 ( .CLK(mc_clk_i_bF_buf1), .D(\mc_dp_pad_i[2] ), .Q(mc_data_ir_34_));
DFFPOSX1 DFFPOSX1_769 ( .CLK(mc_clk_i_bF_buf0), .D(\mc_dp_pad_i[3] ), .Q(mc_data_ir_35_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_i_bF_buf87), .D(u0_u0__0csc_31_0__3_), .Q(u0_csc0_3_));
DFFPOSX1 DFFPOSX1_770 ( .CLK(mc_clk_i_bF_buf10), .D(mc_sts_pad_i), .Q(mc_sts_ir));
DFFPOSX1 DFFPOSX1_771 ( .CLK(mc_clk_i_bF_buf9), .D(_auto_iopadmap_cc_368_execute_85556), .Q(_auto_iopadmap_cc_368_execute_85521));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_i_bF_buf86), .D(u0_u0__0csc_31_0__4_), .Q(u0_csc0_4_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_i_bF_buf85), .D(u0_u0__0csc_31_0__5_), .Q(u0_csc0_5_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_i_bF_buf89), .D(u0__0poc_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_85523_4_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_i_bF_buf84), .D(u0_u0__0csc_31_0__6_), .Q(u0_csc0_6_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_i_bF_buf83), .D(u0_u0__0csc_31_0__7_), .Q(u0_csc0_7_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_i_bF_buf82), .D(u0_u0__0csc_31_0__8_), .Q(u0_csc0_8_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_i_bF_buf81), .D(u0_u0__0csc_31_0__9_), .Q(u0_csc0_9_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_i_bF_buf80), .D(u0_u0__0csc_31_0__10_), .Q(u0_csc0_10_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_i_bF_buf79), .D(u0_u0__0csc_31_0__11_), .Q(u0_csc0_11_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_i_bF_buf78), .D(u0_u0__0csc_31_0__12_), .Q(u0_csc0_12_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_i_bF_buf77), .D(u0_u0__0csc_31_0__13_), .Q(u0_csc0_13_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_i_bF_buf76), .D(u0_u0__0csc_31_0__14_), .Q(u0_csc0_14_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_i_bF_buf75), .D(u0_u0__0csc_31_0__15_), .Q(u0_csc0_15_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_i_bF_buf88), .D(u0__0poc_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_85523_5_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_i_bF_buf74), .D(u0_u0__0csc_31_0__16_), .Q(u0_csc0_16_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_i_bF_buf73), .D(u0_u0__0csc_31_0__17_), .Q(u0_csc0_17_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_i_bF_buf72), .D(u0_u0__0csc_31_0__18_), .Q(u0_csc0_18_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_i_bF_buf71), .D(u0_u0__0csc_31_0__19_), .Q(u0_csc0_19_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_i_bF_buf70), .D(u0_u0__0csc_31_0__20_), .Q(u0_csc0_20_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_i_bF_buf69), .D(u0_u0__0csc_31_0__21_), .Q(u0_csc0_21_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_i_bF_buf68), .D(u0_u0__0csc_31_0__22_), .Q(u0_csc0_22_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_i_bF_buf67), .D(u0_u0__0csc_31_0__23_), .Q(u0_csc0_23_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_i_bF_buf66), .D(u0_u0__0csc_31_0__24_), .Q(u0_csc0_24_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_i_bF_buf65), .D(u0_u0__0csc_31_0__25_), .Q(u0_csc0_25_));
DFFSR DFFSR_1 ( .CLK(clk_i_bF_buf55), .D(u0__0lmr_req_0_0_), .Q(lmr_req), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10), .S(1'h1));
DFFSR DFFSR_10 ( .CLK(clk_i_bF_buf46), .D(u0__0spec_req_cs_7_0__6_), .Q(spec_req_cs_6_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1), .S(1'h1));
DFFSR DFFSR_100 ( .CLK(clk_i_bF_buf53), .D(u0__0csc_mask_r_10_0__2_), .Q(u0_csc_mask_2_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10));
DFFSR DFFSR_101 ( .CLK(clk_i_bF_buf52), .D(u0__0csc_mask_r_10_0__3_), .Q(u0_csc_mask_3_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9));
DFFSR DFFSR_102 ( .CLK(clk_i_bF_buf51), .D(u0__0csc_mask_r_10_0__4_), .Q(u0_csc_mask_4_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8));
DFFSR DFFSR_103 ( .CLK(clk_i_bF_buf50), .D(u0__0csc_mask_r_10_0__5_), .Q(u0_csc_mask_5_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7));
DFFSR DFFSR_104 ( .CLK(clk_i_bF_buf49), .D(u0__0csc_mask_r_10_0__6_), .Q(u0_csc_mask_6_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6));
DFFSR DFFSR_105 ( .CLK(clk_i_bF_buf48), .D(u0__0csc_mask_r_10_0__7_), .Q(u0_csc_mask_7_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5));
DFFSR DFFSR_106 ( .CLK(clk_i_bF_buf47), .D(u0__0csc_mask_r_10_0__8_), .Q(u0_csc_mask_8_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4));
DFFSR DFFSR_107 ( .CLK(clk_i_bF_buf46), .D(u0__0csc_mask_r_10_0__9_), .Q(u0_csc_mask_9_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3));
DFFSR DFFSR_108 ( .CLK(clk_i_bF_buf45), .D(u0__0csc_mask_r_10_0__10_), .Q(u0_csc_mask_10_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2));
DFFSR DFFSR_109 ( .CLK(clk_i_bF_buf44), .D(u0__0csr_r_10_1__0_), .Q(u0_csr_1_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1), .S(1'h1));
DFFSR DFFSR_11 ( .CLK(clk_i_bF_buf45), .D(u0__0spec_req_cs_7_0__7_), .Q(spec_req_cs_7_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0), .S(1'h1));
DFFSR DFFSR_110 ( .CLK(clk_i_bF_buf43), .D(u0__0csr_r_10_1__1_), .Q(fs), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0), .S(1'h1));
DFFSR DFFSR_111 ( .CLK(clk_i_bF_buf42), .D(u0__0csr_r_10_1__2_), .Q(u0_csr_3_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10), .S(1'h1));
DFFSR DFFSR_112 ( .CLK(clk_i_bF_buf41), .D(u0__0csr_r_10_1__3_), .Q(u0_csr_4_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9), .S(1'h1));
DFFSR DFFSR_113 ( .CLK(clk_i_bF_buf40), .D(u0__0csr_r_10_1__4_), .Q(u0_csr_5_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8), .S(1'h1));
DFFSR DFFSR_114 ( .CLK(clk_i_bF_buf39), .D(u0__0csr_r_10_1__5_), .Q(u0_csr_6_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7), .S(1'h1));
DFFSR DFFSR_115 ( .CLK(clk_i_bF_buf38), .D(u0__0csr_r_10_1__6_), .Q(u0_csr_7_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6), .S(1'h1));
DFFSR DFFSR_116 ( .CLK(clk_i_bF_buf37), .D(u0__0csr_r_10_1__7_), .Q(ref_int_0_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5), .S(1'h1));
DFFSR DFFSR_117 ( .CLK(clk_i_bF_buf36), .D(u0__0csr_r_10_1__8_), .Q(ref_int_1_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4), .S(1'h1));
DFFSR DFFSR_118 ( .CLK(clk_i_bF_buf35), .D(u0__0csr_r_10_1__9_), .Q(ref_int_2_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3), .S(1'h1));
DFFSR DFFSR_119 ( .CLK(clk_i_bF_buf34), .D(u0__0csr_r2_7_0__0_), .Q(rfr_ps_val_0_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2), .S(1'h1));
DFFSR DFFSR_12 ( .CLK(clk_i_bF_buf44), .D(u0__0sp_tms_31_0__0_), .Q(sp_tms_0_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10));
DFFSR DFFSR_120 ( .CLK(clk_i_bF_buf33), .D(u0__0csr_r2_7_0__1_), .Q(rfr_ps_val_1_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1), .S(1'h1));
DFFSR DFFSR_121 ( .CLK(clk_i_bF_buf32), .D(u0__0csr_r2_7_0__2_), .Q(rfr_ps_val_2_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0), .S(1'h1));
DFFSR DFFSR_122 ( .CLK(clk_i_bF_buf31), .D(u0__0csr_r2_7_0__3_), .Q(rfr_ps_val_3_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10), .S(1'h1));
DFFSR DFFSR_123 ( .CLK(clk_i_bF_buf30), .D(u0__0csr_r2_7_0__4_), .Q(rfr_ps_val_4_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9), .S(1'h1));
DFFSR DFFSR_124 ( .CLK(clk_i_bF_buf29), .D(u0__0csr_r2_7_0__5_), .Q(rfr_ps_val_5_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8), .S(1'h1));
DFFSR DFFSR_125 ( .CLK(clk_i_bF_buf28), .D(u0__0csr_r2_7_0__6_), .Q(rfr_ps_val_6_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7), .S(1'h1));
DFFSR DFFSR_126 ( .CLK(clk_i_bF_buf27), .D(u0__0csr_r2_7_0__7_), .Q(rfr_ps_val_7_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6), .S(1'h1));
DFFSR DFFSR_127 ( .CLK(clk_i_bF_buf26), .D(u0__0rf_we_0_0_), .Q(u0_rf_we), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5), .S(1'h1));
DFFSR DFFSR_128 ( .CLK(clk_i_bF_buf53), .D(u0_u0__0inited_0_0_), .Q(u0_u0_inited), .R(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494), .S(1'h1));
DFFSR DFFSR_129 ( .CLK(clk_i_bF_buf52), .D(u0_u0__0init_req_0_0_), .Q(u0_init_req0), .R(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494), .S(1'h1));
DFFSR DFFSR_13 ( .CLK(clk_i_bF_buf43), .D(u0__0sp_tms_31_0__1_), .Q(sp_tms_1_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9));
DFFSR DFFSR_130 ( .CLK(clk_i_bF_buf51), .D(u0_u0__0init_req_we_0_0_bF_buf2_), .Q(u0_u0_init_req_we), .R(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494), .S(1'h1));
DFFSR DFFSR_131 ( .CLK(clk_i_bF_buf50), .D(u0_u0__0lmr_req_0_0_), .Q(u0_lmr_req0), .R(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494), .S(1'h1));
DFFSR DFFSR_132 ( .CLK(clk_i_bF_buf49), .D(u0_u0__0lmr_req_we_0_0_bF_buf1_), .Q(u0_u0_lmr_req_we), .R(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494), .S(1'h1));
DFFSR DFFSR_133 ( .CLK(clk_i_bF_buf48), .D(1'h0), .Q(u0_u0_rst_r2), .R(1'h1), .S(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494));
DFFSR DFFSR_134 ( .CLK(clk_i_bF_buf75), .D(u0_u1__0inited_0_0_), .Q(u0_u1_inited), .R(u0_u1__abc_72579_auto_rtlil_cc_1942_NotGate_71506), .S(1'h1));
DFFSR DFFSR_135 ( .CLK(clk_i_bF_buf74), .D(u0_u1__0init_req_0_0_), .Q(u0_init_req1), .R(u0_u1__abc_72579_auto_rtlil_cc_1942_NotGate_71506), .S(1'h1));
DFFSR DFFSR_136 ( .CLK(clk_i_bF_buf73), .D(u0_u1__0init_req_we_0_0_bF_buf7_), .Q(u0_u1_init_req_we), .R(u0_u1__abc_72579_auto_rtlil_cc_1942_NotGate_71506), .S(1'h1));
DFFSR DFFSR_137 ( .CLK(clk_i_bF_buf72), .D(u0_u1__0lmr_req_0_0_), .Q(u0_lmr_req1), .R(u0_u1__abc_72579_auto_rtlil_cc_1942_NotGate_71506), .S(1'h1));
DFFSR DFFSR_138 ( .CLK(clk_i_bF_buf71), .D(u0_u1__0lmr_req_we_0_0_bF_buf7_), .Q(u0_u1_lmr_req_we), .R(u0_u1__abc_72579_auto_rtlil_cc_1942_NotGate_71506), .S(1'h1));
DFFSR DFFSR_139 ( .CLK(clk_i_bF_buf70), .D(1'h0), .Q(u0_u1_rst_r2), .R(1'h1), .S(u0_u1__abc_72579_auto_rtlil_cc_1942_NotGate_71506));
DFFSR DFFSR_14 ( .CLK(clk_i_bF_buf42), .D(u0__0sp_tms_31_0__2_), .Q(sp_tms_2_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8));
DFFSR DFFSR_140 ( .CLK(clk_i_bF_buf26), .D(u2_u0__0bank3_open_0_0_), .Q(u2_u0_bank3_open), .R(u2_u0__abc_74955_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_141 ( .CLK(clk_i_bF_buf25), .D(u2_u0__0bank2_open_0_0_), .Q(u2_u0_bank2_open), .R(u2_u0__abc_74955_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_142 ( .CLK(clk_i_bF_buf24), .D(u2_u0__0bank1_open_0_0_), .Q(u2_u0_bank1_open), .R(u2_u0__abc_74955_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_143 ( .CLK(clk_i_bF_buf23), .D(u2_u0__0bank0_open_0_0_), .Q(u2_u0_bank0_open), .R(u2_u0__abc_74955_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_144 ( .CLK(clk_i_bF_buf67), .D(u2_u1__0bank3_open_0_0_), .Q(u2_u1_bank3_open), .R(u2_u1__abc_74955_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_145 ( .CLK(clk_i_bF_buf66), .D(u2_u1__0bank2_open_0_0_), .Q(u2_u1_bank2_open), .R(u2_u1__abc_74955_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_146 ( .CLK(clk_i_bF_buf65), .D(u2_u1__0bank1_open_0_0_), .Q(u2_u1_bank1_open), .R(u2_u1__abc_74955_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_147 ( .CLK(clk_i_bF_buf64), .D(u2_u1__0bank0_open_0_0_), .Q(u2_u1_bank0_open), .R(u2_u1__abc_74955_auto_rtlil_cc_1942_NotGate_71538), .S(1'h1));
DFFSR DFFSR_148 ( .CLK(clk_i_bF_buf53), .D(u3_u0__0wr_adr_3_0__0_), .Q(u3_u0_wr_adr_0_), .R(1'h1), .S(u3_u0__abc_75526_auto_rtlil_cc_1942_NotGate_71546));
DFFSR DFFSR_149 ( .CLK(clk_i_bF_buf52), .D(u3_u0__0wr_adr_3_0__1_), .Q(u3_u0_wr_adr_1_), .R(u3_u0__abc_75526_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_15 ( .CLK(clk_i_bF_buf41), .D(u0__0sp_tms_31_0__3_), .Q(sp_tms_3_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7));
DFFSR DFFSR_150 ( .CLK(clk_i_bF_buf51), .D(u3_u0__0wr_adr_3_0__2_), .Q(u3_u0_wr_adr_2_), .R(u3_u0__abc_75526_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_151 ( .CLK(clk_i_bF_buf50), .D(u3_u0__0wr_adr_3_0__3_), .Q(u3_u0_wr_adr_3_), .R(u3_u0__abc_75526_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_152 ( .CLK(clk_i_bF_buf49), .D(u3_u0__0rd_adr_3_0__0_), .Q(u3_u0_rd_adr_0_), .R(1'h1), .S(u3_u0__abc_75526_auto_rtlil_cc_1942_NotGate_71546));
DFFSR DFFSR_153 ( .CLK(clk_i_bF_buf48), .D(u3_u0__0rd_adr_3_0__1_), .Q(u3_u0_rd_adr_1_), .R(u3_u0__abc_75526_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_154 ( .CLK(clk_i_bF_buf47), .D(u3_u0__0rd_adr_3_0__2_), .Q(u3_u0_rd_adr_2_), .R(u3_u0__abc_75526_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_155 ( .CLK(clk_i_bF_buf46), .D(u3_u0__0rd_adr_3_0__3_), .Q(u3_u0_rd_adr_3_), .R(u3_u0__abc_75526_auto_rtlil_cc_1942_NotGate_71546), .S(1'h1));
DFFSR DFFSR_156 ( .CLK(clk_i_bF_buf44), .D(u4__0rfr_req_0_0_), .Q(rfr_req), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf3), .S(1'h1));
DFFSR DFFSR_157 ( .CLK(clk_i_bF_buf43), .D(u4__0rfr_cnt_7_0__0_), .Q(u4_rfr_cnt_0_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf2), .S(1'h1));
DFFSR DFFSR_158 ( .CLK(clk_i_bF_buf42), .D(u4__0rfr_cnt_7_0__1_), .Q(u4_rfr_cnt_1_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf1), .S(1'h1));
DFFSR DFFSR_159 ( .CLK(clk_i_bF_buf41), .D(u4__0rfr_cnt_7_0__2_), .Q(u4_rfr_cnt_2_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf0), .S(1'h1));
DFFSR DFFSR_16 ( .CLK(clk_i_bF_buf40), .D(u0__0sp_tms_31_0__4_), .Q(sp_tms_4_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6));
DFFSR DFFSR_160 ( .CLK(clk_i_bF_buf40), .D(u4__0rfr_cnt_7_0__3_), .Q(u4_rfr_cnt_3_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf3), .S(1'h1));
DFFSR DFFSR_161 ( .CLK(clk_i_bF_buf39), .D(u4__0rfr_cnt_7_0__4_), .Q(u4_rfr_cnt_4_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf2), .S(1'h1));
DFFSR DFFSR_162 ( .CLK(clk_i_bF_buf38), .D(u4__0rfr_cnt_7_0__5_), .Q(u4_rfr_cnt_5_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf1), .S(1'h1));
DFFSR DFFSR_163 ( .CLK(clk_i_bF_buf37), .D(u4__0rfr_cnt_7_0__6_), .Q(u4_rfr_cnt_6_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf0), .S(1'h1));
DFFSR DFFSR_164 ( .CLK(clk_i_bF_buf36), .D(u4__0rfr_cnt_7_0__7_), .Q(u4_rfr_cnt_7_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf3), .S(1'h1));
DFFSR DFFSR_165 ( .CLK(clk_i_bF_buf35), .D(u4_ps_cnt_clr), .Q(u4_rfr_ce), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf2), .S(1'h1));
DFFSR DFFSR_166 ( .CLK(clk_i_bF_buf34), .D(u4__0rfr_early_0_0_), .Q(u4_rfr_early), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf1), .S(1'h1));
DFFSR DFFSR_167 ( .CLK(clk_i_bF_buf33), .D(u4__0ps_cnt_7_0__0_), .Q(u4_ps_cnt_0_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf0), .S(1'h1));
DFFSR DFFSR_168 ( .CLK(clk_i_bF_buf32), .D(u4__0ps_cnt_7_0__1_), .Q(u4_ps_cnt_1_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf3), .S(1'h1));
DFFSR DFFSR_169 ( .CLK(clk_i_bF_buf31), .D(u4__0ps_cnt_7_0__2_), .Q(u4_ps_cnt_2_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf2), .S(1'h1));
DFFSR DFFSR_17 ( .CLK(clk_i_bF_buf39), .D(u0__0sp_tms_31_0__5_), .Q(sp_tms_5_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5));
DFFSR DFFSR_170 ( .CLK(clk_i_bF_buf30), .D(u4__0ps_cnt_7_0__3_), .Q(u4_ps_cnt_3_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf1), .S(1'h1));
DFFSR DFFSR_171 ( .CLK(clk_i_bF_buf29), .D(u4__0ps_cnt_7_0__4_), .Q(u4_ps_cnt_4_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf0), .S(1'h1));
DFFSR DFFSR_172 ( .CLK(clk_i_bF_buf28), .D(u4__0ps_cnt_7_0__5_), .Q(u4_ps_cnt_5_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf3), .S(1'h1));
DFFSR DFFSR_173 ( .CLK(clk_i_bF_buf27), .D(u4__0ps_cnt_7_0__6_), .Q(u4_ps_cnt_6_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf2), .S(1'h1));
DFFSR DFFSR_174 ( .CLK(clk_i_bF_buf26), .D(u4__0ps_cnt_7_0__7_), .Q(u4_ps_cnt_7_), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf1), .S(1'h1));
DFFSR DFFSR_175 ( .CLK(clk_i_bF_buf25), .D(u4__0rfr_en_0_0_), .Q(u4_rfr_en), .R(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562_bF_buf0), .S(1'h1));
DFFSR DFFSR_176 ( .CLK(clk_i_bF_buf78), .D(u5_next_state_0_), .Q(u5_state_0_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9));
DFFSR DFFSR_177 ( .CLK(clk_i_bF_buf77), .D(u5_next_state_1_), .Q(u5_state_1_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8), .S(1'h1));
DFFSR DFFSR_178 ( .CLK(clk_i_bF_buf76), .D(u5_next_state_2_), .Q(u5_state_2_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_179 ( .CLK(clk_i_bF_buf75), .D(u5_next_state_3_), .Q(u5_state_3_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6), .S(1'h1));
DFFSR DFFSR_18 ( .CLK(clk_i_bF_buf38), .D(u0__0sp_tms_31_0__6_), .Q(sp_tms_6_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4));
DFFSR DFFSR_180 ( .CLK(clk_i_bF_buf74), .D(u5_next_state_4_), .Q(u5_state_4_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5), .S(1'h1));
DFFSR DFFSR_181 ( .CLK(clk_i_bF_buf73), .D(u5_next_state_5_), .Q(u5_state_5_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4), .S(1'h1));
DFFSR DFFSR_182 ( .CLK(clk_i_bF_buf72), .D(u5_next_state_6_), .Q(u5_state_6_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3), .S(1'h1));
DFFSR DFFSR_183 ( .CLK(clk_i_bF_buf71), .D(u5_next_state_7_), .Q(u5_state_7_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2), .S(1'h1));
DFFSR DFFSR_184 ( .CLK(clk_i_bF_buf70), .D(u5_next_state_8_), .Q(u5_state_8_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_185 ( .CLK(clk_i_bF_buf69), .D(u5_next_state_9_), .Q(u5_state_9_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0), .S(1'h1));
DFFSR DFFSR_186 ( .CLK(clk_i_bF_buf68), .D(u5_next_state_10_), .Q(u5_state_10_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9), .S(1'h1));
DFFSR DFFSR_187 ( .CLK(clk_i_bF_buf67), .D(u5_next_state_11_), .Q(u5_state_11_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8), .S(1'h1));
DFFSR DFFSR_188 ( .CLK(clk_i_bF_buf66), .D(u5_next_state_12_), .Q(u5_state_12_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_189 ( .CLK(clk_i_bF_buf65), .D(u5_next_state_13_), .Q(u5_state_13_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6), .S(1'h1));
DFFSR DFFSR_19 ( .CLK(clk_i_bF_buf37), .D(u0__0sp_tms_31_0__7_), .Q(sp_tms_7_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3));
DFFSR DFFSR_190 ( .CLK(clk_i_bF_buf64), .D(u5_next_state_14_), .Q(u5_state_14_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5), .S(1'h1));
DFFSR DFFSR_191 ( .CLK(clk_i_bF_buf63), .D(u5_next_state_15_), .Q(u5_state_15_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4), .S(1'h1));
DFFSR DFFSR_192 ( .CLK(clk_i_bF_buf62), .D(u5_next_state_16_), .Q(u5_state_16_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3), .S(1'h1));
DFFSR DFFSR_193 ( .CLK(clk_i_bF_buf61), .D(u5_next_state_17_), .Q(u5_state_17_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2), .S(1'h1));
DFFSR DFFSR_194 ( .CLK(clk_i_bF_buf60), .D(u5_next_state_18_), .Q(u5_state_18_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_195 ( .CLK(clk_i_bF_buf59), .D(u5_next_state_19_), .Q(u5_state_19_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0), .S(1'h1));
DFFSR DFFSR_196 ( .CLK(clk_i_bF_buf58), .D(u5_next_state_20_), .Q(u5_state_20_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9), .S(1'h1));
DFFSR DFFSR_197 ( .CLK(clk_i_bF_buf57), .D(u5_next_state_21_), .Q(u5_state_21_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8), .S(1'h1));
DFFSR DFFSR_198 ( .CLK(clk_i_bF_buf56), .D(u5_next_state_22_), .Q(u5_state_22_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_199 ( .CLK(clk_i_bF_buf55), .D(u5_next_state_23_), .Q(u5_state_23_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6), .S(1'h1));
DFFSR DFFSR_2 ( .CLK(clk_i_bF_buf54), .D(u0__0init_req_0_0_), .Q(init_req), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9), .S(1'h1));
DFFSR DFFSR_20 ( .CLK(clk_i_bF_buf36), .D(u0__0sp_tms_31_0__8_), .Q(sp_tms_8_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2));
DFFSR DFFSR_200 ( .CLK(clk_i_bF_buf54), .D(u5_next_state_24_), .Q(u5_state_24_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5), .S(1'h1));
DFFSR DFFSR_201 ( .CLK(clk_i_bF_buf53), .D(u5_next_state_25_), .Q(u5_state_25_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4), .S(1'h1));
DFFSR DFFSR_202 ( .CLK(clk_i_bF_buf52), .D(u5_next_state_26_), .Q(u5_state_26_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3), .S(1'h1));
DFFSR DFFSR_203 ( .CLK(clk_i_bF_buf51), .D(u5_next_state_27_), .Q(u5_state_27_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2), .S(1'h1));
DFFSR DFFSR_204 ( .CLK(clk_i_bF_buf50), .D(u5_next_state_28_), .Q(u5_state_28_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_205 ( .CLK(clk_i_bF_buf49), .D(u5_next_state_29_), .Q(u5_state_29_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0), .S(1'h1));
DFFSR DFFSR_206 ( .CLK(clk_i_bF_buf48), .D(u5_next_state_30_), .Q(u5_state_30_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9), .S(1'h1));
DFFSR DFFSR_207 ( .CLK(clk_i_bF_buf47), .D(u5_next_state_31_), .Q(u5_state_31_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8), .S(1'h1));
DFFSR DFFSR_208 ( .CLK(clk_i_bF_buf46), .D(u5_next_state_32_), .Q(u5_state_32_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_209 ( .CLK(clk_i_bF_buf45), .D(u5_next_state_33_), .Q(u5_state_33_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6), .S(1'h1));
DFFSR DFFSR_21 ( .CLK(clk_i_bF_buf35), .D(u0__0sp_tms_31_0__9_), .Q(sp_tms_9_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1));
DFFSR DFFSR_210 ( .CLK(clk_i_bF_buf44), .D(u5_next_state_34_), .Q(u5_state_34_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5), .S(1'h1));
DFFSR DFFSR_211 ( .CLK(clk_i_bF_buf43), .D(u5_next_state_35_), .Q(u5_state_35_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4), .S(1'h1));
DFFSR DFFSR_212 ( .CLK(clk_i_bF_buf42), .D(u5_next_state_36_), .Q(u5_state_36_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3), .S(1'h1));
DFFSR DFFSR_213 ( .CLK(clk_i_bF_buf41), .D(u5_next_state_37_), .Q(u5_state_37_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2), .S(1'h1));
DFFSR DFFSR_214 ( .CLK(clk_i_bF_buf40), .D(u5_next_state_38_), .Q(u5_state_38_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_215 ( .CLK(clk_i_bF_buf39), .D(u5_next_state_39_), .Q(u5_state_39_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0), .S(1'h1));
DFFSR DFFSR_216 ( .CLK(clk_i_bF_buf38), .D(u5_next_state_40_), .Q(u5_state_40_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9), .S(1'h1));
DFFSR DFFSR_217 ( .CLK(clk_i_bF_buf37), .D(u5_next_state_41_), .Q(u5_state_41_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8), .S(1'h1));
DFFSR DFFSR_218 ( .CLK(clk_i_bF_buf36), .D(u5_next_state_42_), .Q(u5_state_42_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_219 ( .CLK(clk_i_bF_buf35), .D(u5_next_state_43_), .Q(u5_state_43_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6), .S(1'h1));
DFFSR DFFSR_22 ( .CLK(clk_i_bF_buf34), .D(u0__0sp_tms_31_0__10_), .Q(sp_tms_10_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0));
DFFSR DFFSR_220 ( .CLK(clk_i_bF_buf34), .D(u5_next_state_44_), .Q(u5_state_44_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5), .S(1'h1));
DFFSR DFFSR_221 ( .CLK(clk_i_bF_buf33), .D(u5_next_state_45_), .Q(u5_state_45_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4), .S(1'h1));
DFFSR DFFSR_222 ( .CLK(clk_i_bF_buf32), .D(u5_next_state_46_), .Q(u5_state_46_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3), .S(1'h1));
DFFSR DFFSR_223 ( .CLK(clk_i_bF_buf31), .D(u5_next_state_47_), .Q(u5_state_47_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2), .S(1'h1));
DFFSR DFFSR_224 ( .CLK(clk_i_bF_buf30), .D(u5_next_state_48_), .Q(u5_state_48_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_225 ( .CLK(clk_i_bF_buf29), .D(u5_next_state_49_), .Q(u5_state_49_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0), .S(1'h1));
DFFSR DFFSR_226 ( .CLK(clk_i_bF_buf28), .D(u5_next_state_50_), .Q(u5_state_50_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9), .S(1'h1));
DFFSR DFFSR_227 ( .CLK(clk_i_bF_buf27), .D(u5_next_state_51_), .Q(u5_state_51_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8), .S(1'h1));
DFFSR DFFSR_228 ( .CLK(clk_i_bF_buf26), .D(u5_next_state_52_), .Q(u5_state_52_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_229 ( .CLK(clk_i_bF_buf25), .D(u5_next_state_53_), .Q(u5_state_53_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6), .S(1'h1));
DFFSR DFFSR_23 ( .CLK(clk_i_bF_buf33), .D(u0__0sp_tms_31_0__11_), .Q(sp_tms_11_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10));
DFFSR DFFSR_230 ( .CLK(clk_i_bF_buf24), .D(u5_next_state_54_), .Q(u5_state_54_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5), .S(1'h1));
DFFSR DFFSR_231 ( .CLK(clk_i_bF_buf23), .D(u5_next_state_55_), .Q(u5_state_55_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4), .S(1'h1));
DFFSR DFFSR_232 ( .CLK(clk_i_bF_buf22), .D(u5_next_state_56_), .Q(u5_state_56_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3), .S(1'h1));
DFFSR DFFSR_233 ( .CLK(clk_i_bF_buf21), .D(u5_next_state_57_), .Q(u5_state_57_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2), .S(1'h1));
DFFSR DFFSR_234 ( .CLK(clk_i_bF_buf20), .D(u5_next_state_58_), .Q(u5_state_58_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_235 ( .CLK(clk_i_bF_buf19), .D(u5_next_state_59_), .Q(u5_state_59_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0), .S(1'h1));
DFFSR DFFSR_236 ( .CLK(clk_i_bF_buf18), .D(u5_next_state_60_), .Q(u5_state_60_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9), .S(1'h1));
DFFSR DFFSR_237 ( .CLK(clk_i_bF_buf17), .D(u5_next_state_61_), .Q(u5_state_61_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8), .S(1'h1));
DFFSR DFFSR_238 ( .CLK(clk_i_bF_buf16), .D(u5_next_state_62_), .Q(u5_state_62_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_239 ( .CLK(clk_i_bF_buf15), .D(u5_next_state_63_), .Q(u5_state_63_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6), .S(1'h1));
DFFSR DFFSR_24 ( .CLK(clk_i_bF_buf32), .D(u0__0sp_tms_31_0__12_), .Q(sp_tms_12_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9));
DFFSR DFFSR_240 ( .CLK(clk_i_bF_buf14), .D(u5_next_state_64_), .Q(u5_state_64_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5), .S(1'h1));
DFFSR DFFSR_241 ( .CLK(clk_i_bF_buf13), .D(u5_next_state_65_), .Q(u5_state_65_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4), .S(1'h1));
DFFSR DFFSR_242 ( .CLK(clk_i_bF_buf12), .D(u5__0wb_stb_first_0_0_), .Q(u5_wb_stb_first), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3), .S(1'h1));
DFFSR DFFSR_243 ( .CLK(clk_i_bF_buf11), .D(dv), .Q(u5_dv_r), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2), .S(1'h1));
DFFSR DFFSR_244 ( .CLK(clk_i_bF_buf10), .D(u5__0ap_en_0_0_), .Q(u5_ap_en), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_245 ( .CLK(clk_i_bF_buf9), .D(u5_timer_is_zero), .Q(u5_tmr_done), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0), .S(1'h1));
DFFSR DFFSR_246 ( .CLK(clk_i_bF_buf8), .D(u5__0timer_7_0__0_), .Q(u5_timer_0_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9), .S(1'h1));
DFFSR DFFSR_247 ( .CLK(clk_i_bF_buf7), .D(u5__0timer_7_0__1_), .Q(u5_timer_1_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8));
DFFSR DFFSR_248 ( .CLK(clk_i_bF_buf6), .D(u5__0timer_7_0__2_), .Q(u5_timer_2_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_249 ( .CLK(clk_i_bF_buf5), .D(u5__0timer_7_0__3_), .Q(u5_timer_3_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6));
DFFSR DFFSR_25 ( .CLK(clk_i_bF_buf31), .D(u0__0sp_tms_31_0__13_), .Q(sp_tms_13_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8));
DFFSR DFFSR_250 ( .CLK(clk_i_bF_buf4), .D(u5__0timer_7_0__4_), .Q(u5_timer_4_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5));
DFFSR DFFSR_251 ( .CLK(clk_i_bF_buf3), .D(u5__0timer_7_0__5_), .Q(u5_timer_5_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4));
DFFSR DFFSR_252 ( .CLK(clk_i_bF_buf2), .D(u5__0timer_7_0__6_), .Q(u5_timer_6_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3));
DFFSR DFFSR_253 ( .CLK(clk_i_bF_buf1), .D(u5__0timer_7_0__7_), .Q(u5_timer_7_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2));
DFFSR DFFSR_254 ( .CLK(clk_i_bF_buf0), .D(u5__0tmr2_done_0_0_), .Q(u5_tmr2_done), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_255 ( .CLK(clk_i_bF_buf96), .D(u5__0susp_sel_r_0_0_), .Q(susp_sel), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0), .S(1'h1));
DFFSR DFFSR_256 ( .CLK(clk_i_bF_buf95), .D(u5_rfr_ack_d), .Q(rfr_ack), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9), .S(1'h1));
DFFSR DFFSR_257 ( .CLK(clk_i_bF_buf94), .D(u5_suspended_d), .Q(_auto_iopadmap_cc_368_execute_85556), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8), .S(1'h1));
DFFSR DFFSR_258 ( .CLK(clk_i_bF_buf93), .D(resume_req_i), .Q(u5_resume_req_r), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_259 ( .CLK(clk_i_bF_buf92), .D(susp_req_i), .Q(u5_susp_req_r), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6), .S(1'h1));
DFFSR DFFSR_26 ( .CLK(clk_i_bF_buf30), .D(u0__0sp_tms_31_0__14_), .Q(sp_tms_14_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7));
DFFSR DFFSR_260 ( .CLK(clk_i_bF_buf91), .D(u5__0ack_cnt_3_0__0_), .Q(u5_ack_cnt_0_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5), .S(1'h1));
DFFSR DFFSR_261 ( .CLK(clk_i_bF_buf90), .D(u5__0ack_cnt_3_0__1_), .Q(u5_ack_cnt_1_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4), .S(1'h1));
DFFSR DFFSR_262 ( .CLK(clk_i_bF_buf89), .D(u5__0ack_cnt_3_0__2_), .Q(u5_ack_cnt_2_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3), .S(1'h1));
DFFSR DFFSR_263 ( .CLK(clk_i_bF_buf88), .D(u5__0ack_cnt_3_0__3_), .Q(u5_ack_cnt_3_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2), .S(1'h1));
DFFSR DFFSR_264 ( .CLK(clk_i_bF_buf87), .D(u5__0no_wb_cycle_0_0_), .Q(u5_no_wb_cycle), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_265 ( .CLK(clk_i_bF_buf86), .D(u5__0wb_cycle_0_0_), .Q(u5_wb_cycle), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0), .S(1'h1));
DFFSR DFFSR_266 ( .CLK(clk_i_bF_buf85), .D(u5__0wr_cycle_0_0_), .Q(u1_wr_cycle), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9), .S(1'h1));
DFFSR DFFSR_267 ( .CLK(clk_i_bF_buf84), .D(u5__0lookup_ready2_0_0_), .Q(u5_lookup_ready2), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8), .S(1'h1));
DFFSR DFFSR_268 ( .CLK(clk_i_bF_buf83), .D(u5__0lookup_ready1_0_0_), .Q(u5_lookup_ready1), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_269 ( .CLK(clk_i_bF_buf82), .D(u5__0data_oe_0_0_), .Q(data_oe), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6), .S(1'h1));
DFFSR DFFSR_27 ( .CLK(clk_i_bF_buf29), .D(u0__0sp_tms_31_0__15_), .Q(sp_tms_15_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6));
DFFSR DFFSR_270 ( .CLK(clk_i_bF_buf81), .D(u5_data_oe_r), .Q(u5_data_oe_r2), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5), .S(1'h1));
DFFSR DFFSR_271 ( .CLK(clk_i_bF_buf80), .D(u5_data_oe_d), .Q(u5_data_oe_r), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4), .S(1'h1));
DFFSR DFFSR_272 ( .CLK(clk_i_bF_buf79), .D(u5__0oe__0_0_), .Q(oe_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3));
DFFSR DFFSR_273 ( .CLK(clk_i_bF_buf78), .D(u5__0cmd_asserted2_0_0_), .Q(u5_cmd_asserted2), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2), .S(1'h1));
DFFSR DFFSR_274 ( .CLK(clk_i_bF_buf77), .D(u5__0cmd_asserted_0_0_), .Q(u5_cmd_asserted), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_275 ( .CLK(clk_i_bF_buf76), .D(u5_cmd_r_0_), .Q(u5_cmd_del_0_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0));
DFFSR DFFSR_276 ( .CLK(clk_i_bF_buf75), .D(u5_cmd_r_1_), .Q(u5_cmd_del_1_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9));
DFFSR DFFSR_277 ( .CLK(clk_i_bF_buf74), .D(u5_cmd_r_2_), .Q(u5_cmd_del_2_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8));
DFFSR DFFSR_278 ( .CLK(clk_i_bF_buf73), .D(u5_cmd_r_3_), .Q(u5_cmd_del_3_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf7), .S(1'h1));
DFFSR DFFSR_279 ( .CLK(clk_i_bF_buf72), .D(u5_cmd_0_), .Q(u5_cmd_r_0_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf6));
DFFSR DFFSR_28 ( .CLK(clk_i_bF_buf28), .D(u0__0sp_tms_31_0__16_), .Q(sp_tms_16_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5));
DFFSR DFFSR_280 ( .CLK(clk_i_bF_buf71), .D(u5_cmd_1_), .Q(u5_cmd_r_1_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf5));
DFFSR DFFSR_281 ( .CLK(clk_i_bF_buf70), .D(u5_cmd_2_), .Q(u5_cmd_r_2_), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf4));
DFFSR DFFSR_282 ( .CLK(clk_i_bF_buf69), .D(u5_cmd_3_), .Q(u5_cmd_r_3_), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf3), .S(1'h1));
DFFSR DFFSR_283 ( .CLK(clk_i_bF_buf68), .D(mem_ack), .Q(u5_mem_ack_r), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf2), .S(1'h1));
DFFSR DFFSR_284 ( .CLK(clk_i_bF_buf67), .D(u5__0mc_adv_r_0_0_), .Q(u5_mc_adv_r), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf1), .S(1'h1));
DFFSR DFFSR_285 ( .CLK(clk_i_bF_buf66), .D(u5__0mc_adv_r1_0_0_), .Q(u5_mc_adv_r1), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf0), .S(1'h1));
DFFSR DFFSR_286 ( .CLK(clk_i_bF_buf65), .D(u5__0mc_le_0_0_), .Q(u5_mc_le), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_72182), .S(1'h1));
DFFSR DFFSR_287 ( .CLK(clk_i_bF_buf64), .D(u5_mc_c_oe_d), .Q(mc_c_oe_d), .R(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf9), .S(1'h1));
DFFSR DFFSR_288 ( .CLK(clk_i_bF_buf63), .D(1'h0), .Q(u5_rsts), .R(1'h1), .S(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962_bF_buf8));
DFFSR DFFSR_289 ( .CLK(clk_i_bF_buf30), .D(u6__0wb_err_0_0_), .Q(_auto_iopadmap_cc_368_execute_85593), .R(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_29 ( .CLK(clk_i_bF_buf27), .D(u0__0sp_tms_31_0__17_), .Q(sp_tms_17_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4));
DFFSR DFFSR_290 ( .CLK(clk_i_bF_buf29), .D(u6__0wb_ack_o_0_0_), .Q(_auto_iopadmap_cc_368_execute_85558), .R(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_291 ( .CLK(clk_i_bF_buf28), .D(u6__0wr_hold_0_0_), .Q(u1_wr_hold), .R(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_292 ( .CLK(clk_i_bF_buf27), .D(u6__0wb_first_r_0_0_), .Q(u6_wb_first_r), .R(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_293 ( .CLK(clk_i_bF_buf26), .D(u6__0write_go_r_0_0_), .Q(u6_write_go_r), .R(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_294 ( .CLK(clk_i_bF_buf25), .D(u6__0write_go_r1_0_0_), .Q(u6_write_go_r1), .R(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_295 ( .CLK(clk_i_bF_buf24), .D(u6__0read_go_r_0_0_), .Q(u6_read_go_r), .R(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_296 ( .CLK(clk_i_bF_buf23), .D(u6__0read_go_r1_0_0_), .Q(u6_read_go_r1), .R(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_297 ( .CLK(clk_i_bF_buf22), .D(u6__0rmw_r_0_0_), .Q(u6_rmw_r), .R(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_298 ( .CLK(clk_i_bF_buf21), .D(u6__0rmw_en_0_0_), .Q(u6_rmw_en), .R(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188), .S(1'h1));
DFFSR DFFSR_299 ( .CLK(mc_clk_i_bF_buf8), .D(u7__0mc_cs__7_7_), .Q(_auto_iopadmap_cc_368_execute_85457_7_), .R(1'h1), .S(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_3 ( .CLK(clk_i_bF_buf53), .D(u0__0sreq_cs_le_0_0_), .Q(u0_sreq_cs_le), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8), .S(1'h1));
DFFSR DFFSR_30 ( .CLK(clk_i_bF_buf26), .D(u0__0sp_tms_31_0__18_), .Q(sp_tms_18_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3));
DFFSR DFFSR_300 ( .CLK(mc_clk_i_bF_buf7), .D(u7__0mc_cs__6_6_), .Q(_auto_iopadmap_cc_368_execute_85457_6_), .R(1'h1), .S(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_301 ( .CLK(mc_clk_i_bF_buf6), .D(u7__0mc_cs__5_5_), .Q(_auto_iopadmap_cc_368_execute_85457_5_), .R(1'h1), .S(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_302 ( .CLK(mc_clk_i_bF_buf5), .D(u7__0mc_cs__4_4_), .Q(_auto_iopadmap_cc_368_execute_85457_4_), .R(1'h1), .S(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_303 ( .CLK(mc_clk_i_bF_buf4), .D(u7__0mc_cs__3_3_), .Q(_auto_iopadmap_cc_368_execute_85457_3_), .R(1'h1), .S(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_304 ( .CLK(mc_clk_i_bF_buf3), .D(u7__0mc_cs__2_2_), .Q(_auto_iopadmap_cc_368_execute_85457_2_), .R(1'h1), .S(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_305 ( .CLK(mc_clk_i_bF_buf2), .D(u7__0mc_cs__1_1_), .Q(_auto_iopadmap_cc_368_execute_85457_1_), .R(1'h1), .S(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_306 ( .CLK(mc_clk_i_bF_buf1), .D(u7__0mc_cs__0_0_), .Q(_auto_iopadmap_cc_368_execute_85457_0_), .R(1'h1), .S(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_307 ( .CLK(mc_clk_i_bF_buf0), .D(u7__0mc_oe__0_0_), .Q(_auto_iopadmap_cc_368_execute_85511), .R(1'h1), .S(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518));
DFFSR DFFSR_308 ( .CLK(mc_clk_i_bF_buf10), .D(u7__0mc_data_oe_0_0_), .Q(_auto_iopadmap_cc_368_execute_85499), .R(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518), .S(1'h1));
DFFSR DFFSR_31 ( .CLK(clk_i_bF_buf25), .D(u0__0sp_tms_31_0__19_), .Q(sp_tms_19_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2));
DFFSR DFFSR_32 ( .CLK(clk_i_bF_buf24), .D(u0__0sp_tms_31_0__20_), .Q(sp_tms_20_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1));
DFFSR DFFSR_33 ( .CLK(clk_i_bF_buf23), .D(u0__0sp_tms_31_0__21_), .Q(sp_tms_21_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0));
DFFSR DFFSR_34 ( .CLK(clk_i_bF_buf22), .D(u0__0sp_tms_31_0__22_), .Q(sp_tms_22_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10));
DFFSR DFFSR_35 ( .CLK(clk_i_bF_buf21), .D(u0__0sp_tms_31_0__23_), .Q(sp_tms_23_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9));
DFFSR DFFSR_36 ( .CLK(clk_i_bF_buf20), .D(u0__0sp_tms_31_0__24_), .Q(sp_tms_24_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8));
DFFSR DFFSR_37 ( .CLK(clk_i_bF_buf19), .D(u0__0sp_tms_31_0__25_), .Q(sp_tms_25_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7));
DFFSR DFFSR_38 ( .CLK(clk_i_bF_buf18), .D(u0__0sp_tms_31_0__26_), .Q(sp_tms_26_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6));
DFFSR DFFSR_39 ( .CLK(clk_i_bF_buf17), .D(u0__0sp_tms_31_0__27_), .Q(sp_tms_27_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5));
DFFSR DFFSR_4 ( .CLK(clk_i_bF_buf52), .D(u0__0spec_req_cs_7_0__0_), .Q(spec_req_cs_0_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7), .S(1'h1));
DFFSR DFFSR_40 ( .CLK(clk_i_bF_buf16), .D(u0__0sp_csc_31_0__1_), .Q(sp_csc_1_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4), .S(1'h1));
DFFSR DFFSR_41 ( .CLK(clk_i_bF_buf15), .D(u0__0sp_csc_31_0__2_), .Q(sp_csc_2_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3), .S(1'h1));
DFFSR DFFSR_42 ( .CLK(clk_i_bF_buf14), .D(u0__0sp_csc_31_0__3_), .Q(sp_csc_3_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2), .S(1'h1));
DFFSR DFFSR_43 ( .CLK(clk_i_bF_buf13), .D(u0__0sp_csc_31_0__4_), .Q(sp_csc_4_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1), .S(1'h1));
DFFSR DFFSR_44 ( .CLK(clk_i_bF_buf12), .D(u0__0sp_csc_31_0__5_), .Q(sp_csc_5_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0), .S(1'h1));
DFFSR DFFSR_45 ( .CLK(clk_i_bF_buf11), .D(u0__0sp_csc_31_0__6_), .Q(sp_csc_6_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10), .S(1'h1));
DFFSR DFFSR_46 ( .CLK(clk_i_bF_buf10), .D(u0__0sp_csc_31_0__7_), .Q(sp_csc_7_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9), .S(1'h1));
DFFSR DFFSR_47 ( .CLK(clk_i_bF_buf9), .D(u0__0sp_csc_31_0__9_), .Q(sp_csc_9_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8), .S(1'h1));
DFFSR DFFSR_48 ( .CLK(clk_i_bF_buf8), .D(u0__0sp_csc_31_0__10_), .Q(sp_csc_10_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7), .S(1'h1));
DFFSR DFFSR_49 ( .CLK(clk_i_bF_buf7), .D(u0__0tms_31_0__0_), .Q(tms_0_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6));
DFFSR DFFSR_5 ( .CLK(clk_i_bF_buf51), .D(u0__0spec_req_cs_7_0__1_), .Q(spec_req_cs_1_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6), .S(1'h1));
DFFSR DFFSR_50 ( .CLK(clk_i_bF_buf6), .D(u0__0tms_31_0__1_), .Q(tms_1_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5));
DFFSR DFFSR_51 ( .CLK(clk_i_bF_buf5), .D(u0__0tms_31_0__2_), .Q(tms_2_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4));
DFFSR DFFSR_52 ( .CLK(clk_i_bF_buf4), .D(u0__0tms_31_0__3_), .Q(tms_3_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3));
DFFSR DFFSR_53 ( .CLK(clk_i_bF_buf3), .D(u0__0tms_31_0__4_), .Q(tms_4_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2));
DFFSR DFFSR_54 ( .CLK(clk_i_bF_buf2), .D(u0__0tms_31_0__5_), .Q(tms_5_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1));
DFFSR DFFSR_55 ( .CLK(clk_i_bF_buf1), .D(u0__0tms_31_0__6_), .Q(tms_6_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0));
DFFSR DFFSR_56 ( .CLK(clk_i_bF_buf0), .D(u0__0tms_31_0__7_), .Q(tms_7_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10));
DFFSR DFFSR_57 ( .CLK(clk_i_bF_buf96), .D(u0__0tms_31_0__8_), .Q(tms_8_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9));
DFFSR DFFSR_58 ( .CLK(clk_i_bF_buf95), .D(u0__0tms_31_0__9_), .Q(tms_9_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8));
DFFSR DFFSR_59 ( .CLK(clk_i_bF_buf94), .D(u0__0tms_31_0__10_), .Q(tms_10_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7));
DFFSR DFFSR_6 ( .CLK(clk_i_bF_buf50), .D(u0__0spec_req_cs_7_0__2_), .Q(spec_req_cs_2_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5), .S(1'h1));
DFFSR DFFSR_60 ( .CLK(clk_i_bF_buf93), .D(u0__0tms_31_0__11_), .Q(tms_11_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6));
DFFSR DFFSR_61 ( .CLK(clk_i_bF_buf92), .D(u0__0tms_31_0__12_), .Q(tms_12_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5));
DFFSR DFFSR_62 ( .CLK(clk_i_bF_buf91), .D(u0__0tms_31_0__13_), .Q(tms_13_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4));
DFFSR DFFSR_63 ( .CLK(clk_i_bF_buf90), .D(u0__0tms_31_0__14_), .Q(tms_14_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3));
DFFSR DFFSR_64 ( .CLK(clk_i_bF_buf89), .D(u0__0tms_31_0__15_), .Q(tms_15_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2));
DFFSR DFFSR_65 ( .CLK(clk_i_bF_buf88), .D(u0__0tms_31_0__16_), .Q(tms_16_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1));
DFFSR DFFSR_66 ( .CLK(clk_i_bF_buf87), .D(u0__0tms_31_0__17_), .Q(tms_17_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0));
DFFSR DFFSR_67 ( .CLK(clk_i_bF_buf86), .D(u0__0tms_31_0__18_), .Q(tms_18_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10));
DFFSR DFFSR_68 ( .CLK(clk_i_bF_buf85), .D(u0__0tms_31_0__19_), .Q(tms_19_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9));
DFFSR DFFSR_69 ( .CLK(clk_i_bF_buf84), .D(u0__0tms_31_0__20_), .Q(tms_20_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8));
DFFSR DFFSR_7 ( .CLK(clk_i_bF_buf49), .D(u0__0spec_req_cs_7_0__3_), .Q(spec_req_cs_3_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4), .S(1'h1));
DFFSR DFFSR_70 ( .CLK(clk_i_bF_buf83), .D(u0__0tms_31_0__21_), .Q(tms_21_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7));
DFFSR DFFSR_71 ( .CLK(clk_i_bF_buf82), .D(u0__0tms_31_0__22_), .Q(tms_22_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6));
DFFSR DFFSR_72 ( .CLK(clk_i_bF_buf81), .D(u0__0tms_31_0__23_), .Q(tms_23_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5));
DFFSR DFFSR_73 ( .CLK(clk_i_bF_buf80), .D(u0__0tms_31_0__24_), .Q(tms_24_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4));
DFFSR DFFSR_74 ( .CLK(clk_i_bF_buf79), .D(u0__0tms_31_0__25_), .Q(tms_25_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3));
DFFSR DFFSR_75 ( .CLK(clk_i_bF_buf78), .D(u0__0tms_31_0__26_), .Q(tms_26_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2));
DFFSR DFFSR_76 ( .CLK(clk_i_bF_buf77), .D(u0__0tms_31_0__27_), .Q(tms_27_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1));
DFFSR DFFSR_77 ( .CLK(clk_i_bF_buf76), .D(u0__0csc_31_0__1_), .Q(csc_1_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0), .S(1'h1));
DFFSR DFFSR_78 ( .CLK(clk_i_bF_buf75), .D(u0__0csc_31_0__2_), .Q(csc_2_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10), .S(1'h1));
DFFSR DFFSR_79 ( .CLK(clk_i_bF_buf74), .D(u0__0csc_31_0__3_), .Q(csc_3_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9), .S(1'h1));
DFFSR DFFSR_8 ( .CLK(clk_i_bF_buf48), .D(u0__0spec_req_cs_7_0__4_), .Q(spec_req_cs_4_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3), .S(1'h1));
DFFSR DFFSR_80 ( .CLK(clk_i_bF_buf73), .D(u0__0csc_31_0__4_), .Q(csc_4_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8), .S(1'h1));
DFFSR DFFSR_81 ( .CLK(clk_i_bF_buf72), .D(u0__0csc_31_0__5_), .Q(csc_5_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7), .S(1'h1));
DFFSR DFFSR_82 ( .CLK(clk_i_bF_buf71), .D(u0__0csc_31_0__6_), .Q(csc_6_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6), .S(1'h1));
DFFSR DFFSR_83 ( .CLK(clk_i_bF_buf70), .D(u0__0csc_31_0__7_), .Q(csc_7_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5), .S(1'h1));
DFFSR DFFSR_84 ( .CLK(clk_i_bF_buf69), .D(u0__0csc_31_0__9_), .Q(csc_9_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4), .S(1'h1));
DFFSR DFFSR_85 ( .CLK(clk_i_bF_buf68), .D(u0__0csc_31_0__10_), .Q(csc_10_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3), .S(1'h1));
DFFSR DFFSR_86 ( .CLK(clk_i_bF_buf67), .D(u0__0csc_31_0__11_), .Q(u3_pen), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2), .S(1'h1));
DFFSR DFFSR_87 ( .CLK(clk_i_bF_buf66), .D(u0__0wp_err_0_0_), .Q(u0_wp_err), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1), .S(1'h1));
DFFSR DFFSR_88 ( .CLK(clk_i_bF_buf65), .D(u0__0cs_7_0__0_), .Q(cs_0_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0), .S(1'h1));
DFFSR DFFSR_89 ( .CLK(clk_i_bF_buf64), .D(u0__0cs_7_0__1_), .Q(cs_1_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf10), .S(1'h1));
DFFSR DFFSR_9 ( .CLK(clk_i_bF_buf47), .D(u0__0spec_req_cs_7_0__5_), .Q(spec_req_cs_5_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2), .S(1'h1));
DFFSR DFFSR_90 ( .CLK(clk_i_bF_buf63), .D(u0__0cs_7_0__2_), .Q(cs_2_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf9), .S(1'h1));
DFFSR DFFSR_91 ( .CLK(clk_i_bF_buf62), .D(u0__0cs_7_0__3_), .Q(cs_3_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf8), .S(1'h1));
DFFSR DFFSR_92 ( .CLK(clk_i_bF_buf61), .D(u0__0cs_7_0__4_), .Q(cs_4_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf7), .S(1'h1));
DFFSR DFFSR_93 ( .CLK(clk_i_bF_buf60), .D(u0__0cs_7_0__5_), .Q(cs_5_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf6), .S(1'h1));
DFFSR DFFSR_94 ( .CLK(clk_i_bF_buf59), .D(u0__0cs_7_0__6_), .Q(cs_6_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf5), .S(1'h1));
DFFSR DFFSR_95 ( .CLK(clk_i_bF_buf58), .D(u0__0cs_7_0__7_), .Q(cs_7_), .R(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf4), .S(1'h1));
DFFSR DFFSR_96 ( .CLK(clk_i_bF_buf57), .D(u0_rst_r2), .Q(u0_rst_r3), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf3));
DFFSR DFFSR_97 ( .CLK(clk_i_bF_buf56), .D(1'h0), .Q(u0_rst_r2), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf2));
DFFSR DFFSR_98 ( .CLK(clk_i_bF_buf55), .D(u0__0csc_mask_r_10_0__0_), .Q(u0_csc_mask_0_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf1));
DFFSR DFFSR_99 ( .CLK(clk_i_bF_buf54), .D(u0__0csc_mask_r_10_0__1_), .Q(u0_csc_mask_1_), .R(1'h1), .S(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602_bF_buf0));
INVX1 INVX1_1 ( .A(init_ack), .Y(_abc_85006_new_n238_));
INVX1 INVX1_10 ( .A(u0__abc_76628_new_n1152_), .Y(u0__abc_76628_new_n1159_));
INVX1 INVX1_100 ( .A(\wb_data_i[7] ), .Y(u0_u1__abc_72579_new_n262_));
INVX1 INVX1_1000 ( .A(u5__abc_81276_new_n920_), .Y(u5__abc_81276_new_n2022_));
INVX1 INVX1_1001 ( .A(u5__abc_81276_new_n2029_), .Y(u5__abc_81276_new_n2030_));
INVX1 INVX1_1002 ( .A(u5__abc_81276_new_n2042_), .Y(u5__abc_81276_new_n2043_));
INVX1 INVX1_1003 ( .A(u5__abc_81276_new_n2053_), .Y(u5__abc_81276_new_n2054_));
INVX1 INVX1_1004 ( .A(u5__abc_81276_new_n2058_), .Y(u5__abc_81276_new_n2059_));
INVX1 INVX1_1005 ( .A(u5__abc_81276_new_n2064_), .Y(u5__abc_81276_new_n2065_));
INVX1 INVX1_1006 ( .A(u5__abc_81276_new_n2081_), .Y(u5__abc_81276_new_n2082_));
INVX1 INVX1_1007 ( .A(u5__abc_81276_new_n2094_), .Y(u5__abc_81276_new_n2095_));
INVX1 INVX1_1008 ( .A(u5__abc_81276_new_n2108_), .Y(u5__abc_81276_new_n2109_));
INVX1 INVX1_1009 ( .A(u5__abc_81276_new_n2121_), .Y(u5__abc_81276_new_n2122_));
INVX1 INVX1_101 ( .A(u0_u1__abc_72579_new_n263_), .Y(u0_u1__abc_72579_new_n264_));
INVX1 INVX1_1010 ( .A(u5__abc_81276_new_n1220_), .Y(u5__abc_81276_new_n2245_));
INVX1 INVX1_1011 ( .A(u5__abc_81276_new_n1188_), .Y(u5__abc_81276_new_n2278_));
INVX1 INVX1_1012 ( .A(u5__abc_81276_new_n2294_), .Y(u5__abc_81276_new_n2295_));
INVX1 INVX1_1013 ( .A(u5__abc_81276_new_n1682__bF_buf2), .Y(u5__abc_81276_new_n2309_));
INVX1 INVX1_1014 ( .A(u5__abc_81276_new_n2310_), .Y(u5__abc_81276_new_n2311_));
INVX1 INVX1_1015 ( .A(u5__abc_81276_new_n2312_), .Y(u5__abc_81276_new_n2313_));
INVX1 INVX1_1016 ( .A(u5__abc_81276_new_n2314_), .Y(u5__abc_81276_new_n2315_));
INVX1 INVX1_1017 ( .A(u5__abc_81276_new_n1526__bF_buf2), .Y(u5__abc_81276_new_n2320_));
INVX1 INVX1_1018 ( .A(u5__abc_81276_new_n2323_), .Y(u5__abc_81276_new_n2324_));
INVX1 INVX1_1019 ( .A(u5__abc_81276_new_n2316_), .Y(u5__abc_81276_new_n2325_));
INVX1 INVX1_102 ( .A(\wb_data_i[8] ), .Y(u0_u1__abc_72579_new_n268_));
INVX1 INVX1_1020 ( .A(u5__abc_81276_new_n2327_), .Y(u5__abc_81276_new_n2328_));
INVX1 INVX1_1021 ( .A(u5__abc_81276_new_n2334_), .Y(u5__abc_81276_new_n2336_));
INVX1 INVX1_1022 ( .A(u5__abc_81276_new_n2335_), .Y(u5__abc_81276_new_n2342_));
INVX1 INVX1_1023 ( .A(u5__abc_81276_new_n2344_), .Y(u5__abc_81276_new_n2352_));
INVX1 INVX1_1024 ( .A(u5__abc_81276_new_n2351_), .Y(u5__abc_81276_new_n2361_));
INVX1 INVX1_1025 ( .A(u5__abc_81276_new_n2363_), .Y(u5__abc_81276_new_n2373_));
INVX1 INVX1_1026 ( .A(u5__abc_81276_new_n2375_), .Y(u5__abc_81276_new_n2381_));
INVX1 INVX1_1027 ( .A(u5__abc_81276_new_n2399_), .Y(u5__abc_81276_new_n2401_));
INVX1 INVX1_1028 ( .A(u5__abc_81276_new_n2412_), .Y(u5__abc_81276_new_n2413_));
INVX1 INVX1_1029 ( .A(u5_burst_cnt_8_), .Y(u5__abc_81276_new_n2415_));
INVX1 INVX1_103 ( .A(u0_u1__abc_72579_new_n269_), .Y(u0_u1__abc_72579_new_n270_));
INVX1 INVX1_1030 ( .A(u5__abc_81276_new_n2416_), .Y(u5__abc_81276_new_n2423_));
INVX1 INVX1_1031 ( .A(u5__abc_81276_new_n2433_), .Y(u5__abc_81276_new_n2435_));
INVX1 INVX1_1032 ( .A(u5__abc_81276_new_n2462_), .Y(u5__abc_81276_new_n2464_));
INVX1 INVX1_1033 ( .A(u5__abc_81276_new_n2472_), .Y(u5__abc_81276_new_n2473_));
INVX1 INVX1_1034 ( .A(u5__abc_81276_new_n2475_), .Y(u5__abc_81276_new_n2476_));
INVX1 INVX1_1035 ( .A(u5__abc_81276_new_n2479_), .Y(u5__0ir_cnt_3_0__1_));
INVX1 INVX1_1036 ( .A(u5__abc_81276_new_n2485_), .Y(u5__abc_81276_new_n2486_));
INVX1 INVX1_1037 ( .A(u5__abc_81276_new_n2515_), .Y(u5__abc_81276_new_n2516_));
INVX1 INVX1_1038 ( .A(u5__abc_81276_new_n2527_), .Y(u5__abc_81276_new_n2528_));
INVX1 INVX1_1039 ( .A(u5__abc_81276_new_n2539_), .Y(u5__abc_81276_new_n2540_));
INVX1 INVX1_104 ( .A(\wb_data_i[9] ), .Y(u0_u1__abc_72579_new_n274_));
INVX1 INVX1_1040 ( .A(u5__abc_81276_new_n2548_), .Y(u5__abc_81276_new_n2549_));
INVX1 INVX1_1041 ( .A(u5__abc_81276_new_n2550_), .Y(u5__abc_81276_new_n2551_));
INVX1 INVX1_1042 ( .A(u5__abc_81276_new_n2508_), .Y(u5__abc_81276_new_n2558_));
INVX1 INVX1_1043 ( .A(u5__abc_81276_new_n2569_), .Y(u5__abc_81276_new_n2570_));
INVX1 INVX1_1044 ( .A(u5__abc_81276_new_n2575_), .Y(u5__abc_81276_new_n2576_));
INVX1 INVX1_1045 ( .A(u5__abc_81276_new_n1693_), .Y(u5__abc_81276_new_n2579_));
INVX1 INVX1_1046 ( .A(u5__abc_81276_new_n1534_), .Y(u5__abc_81276_new_n2580_));
INVX1 INVX1_1047 ( .A(u5__abc_81276_new_n2584_), .Y(u5__abc_81276_new_n2585_));
INVX1 INVX1_1048 ( .A(u5__abc_81276_new_n990_), .Y(u5__abc_81276_new_n2595_));
INVX1 INVX1_1049 ( .A(u5__abc_81276_new_n967_), .Y(u5__abc_81276_new_n2596_));
INVX1 INVX1_105 ( .A(u0_u1__abc_72579_new_n275_), .Y(u0_u1__abc_72579_new_n276_));
INVX1 INVX1_1050 ( .A(u5__abc_81276_new_n2641_), .Y(u5__abc_81276_new_n2642_));
INVX1 INVX1_1051 ( .A(u5__abc_81276_new_n1537_), .Y(u5__abc_81276_new_n2658_));
INVX1 INVX1_1052 ( .A(u5__abc_81276_new_n2660_), .Y(u5__abc_81276_new_n2661_));
INVX1 INVX1_1053 ( .A(u5__abc_81276_new_n2541_), .Y(u5__abc_81276_new_n2685_));
INVX1 INVX1_1054 ( .A(u5__abc_81276_new_n2538_), .Y(u5__abc_81276_new_n2689_));
INVX1 INVX1_1055 ( .A(u5__abc_81276_new_n2690_), .Y(u5__abc_81276_new_n2691_));
INVX1 INVX1_1056 ( .A(u5__abc_81276_new_n2704_), .Y(u5__abc_81276_new_n2705_));
INVX1 INVX1_1057 ( .A(u5__abc_81276_new_n2706_), .Y(u5__abc_81276_new_n2709_));
INVX1 INVX1_1058 ( .A(u5__abc_81276_new_n2725_), .Y(u5__abc_81276_new_n2729_));
INVX1 INVX1_1059 ( .A(u5__abc_81276_new_n2744_), .Y(u5__abc_81276_new_n2745_));
INVX1 INVX1_106 ( .A(\wb_data_i[10] ), .Y(u0_u1__abc_72579_new_n280_));
INVX1 INVX1_1060 ( .A(u5__abc_81276_new_n2747_), .Y(u5__abc_81276_new_n2748_));
INVX1 INVX1_1061 ( .A(u5__abc_81276_new_n2751_), .Y(u5__abc_81276_new_n2752_));
INVX1 INVX1_1062 ( .A(u5__abc_81276_new_n2753_), .Y(u5__abc_81276_new_n2754_));
INVX1 INVX1_1063 ( .A(u5__abc_81276_new_n2756_), .Y(u5__abc_81276_new_n2757_));
INVX1 INVX1_1064 ( .A(u5__abc_81276_new_n2758_), .Y(u5__abc_81276_new_n2759_));
INVX1 INVX1_1065 ( .A(u5__abc_81276_new_n2769_), .Y(u5__abc_81276_new_n2770_));
INVX1 INVX1_1066 ( .A(u5__abc_81276_new_n2771_), .Y(u5__abc_81276_new_n2772_));
INVX1 INVX1_1067 ( .A(u5__abc_81276_new_n2773_), .Y(u5__abc_81276_new_n2774_));
INVX1 INVX1_1068 ( .A(u5__abc_81276_new_n2687_), .Y(u5__abc_81276_new_n2783_));
INVX1 INVX1_1069 ( .A(u5__abc_81276_new_n2808_), .Y(u5__abc_81276_new_n2809_));
INVX1 INVX1_107 ( .A(u0_u1__abc_72579_new_n281_), .Y(u0_u1__abc_72579_new_n282_));
INVX1 INVX1_1070 ( .A(u5__abc_81276_new_n2785_), .Y(u5__abc_81276_new_n2819_));
INVX1 INVX1_1071 ( .A(u5__abc_81276_new_n2845_), .Y(u5__abc_81276_new_n2846_));
INVX1 INVX1_1072 ( .A(u5__abc_81276_new_n2867_), .Y(u5__abc_81276_new_n2868_));
INVX1 INVX1_1073 ( .A(u5__abc_81276_new_n2818_), .Y(u5__abc_81276_new_n2874_));
INVX1 INVX1_1074 ( .A(u5__abc_81276_new_n2873_), .Y(u5__abc_81276_new_n2884_));
INVX1 INVX1_1075 ( .A(u5__abc_81276_new_n2883_), .Y(u5__abc_81276_new_n2893_));
INVX1 INVX1_1076 ( .A(u5__abc_81276_new_n2896_), .Y(u5__abc_81276_new_n2904_));
INVX1 INVX1_1077 ( .A(u5__abc_81276_new_n2919_), .Y(u5__abc_81276_new_n2920_));
INVX1 INVX1_1078 ( .A(u5__abc_81276_new_n2930_), .Y(u5__abc_81276_new_n2931_));
INVX1 INVX1_1079 ( .A(u5__abc_81276_new_n2932_), .Y(u5__abc_81276_new_n2933_));
INVX1 INVX1_108 ( .A(\wb_data_i[11] ), .Y(u0_u1__abc_72579_new_n286_));
INVX1 INVX1_1080 ( .A(u5_timer2_0_), .Y(u5__abc_81276_new_n2934_));
INVX1 INVX1_1081 ( .A(u5__abc_81276_new_n1831_), .Y(u5__abc_81276_new_n2963_));
INVX1 INVX1_1082 ( .A(u5__abc_81276_new_n2964_), .Y(u5__abc_81276_new_n2965_));
INVX1 INVX1_1083 ( .A(u5__abc_81276_new_n2968_), .Y(u5__abc_81276_new_n2969_));
INVX1 INVX1_1084 ( .A(u5__abc_81276_new_n2961_), .Y(u5__abc_81276_new_n2970_));
INVX1 INVX1_1085 ( .A(u5__abc_81276_new_n685_), .Y(u5__abc_81276_new_n2980_));
INVX1 INVX1_1086 ( .A(u5__abc_81276_new_n2996_), .Y(u5__abc_81276_new_n2997_));
INVX1 INVX1_1087 ( .A(u5__abc_81276_new_n2935_), .Y(u5__abc_81276_new_n3011_));
INVX1 INVX1_1088 ( .A(u5__abc_81276_new_n2992_), .Y(u5__abc_81276_new_n3018_));
INVX1 INVX1_1089 ( .A(u5__abc_81276_new_n2986_), .Y(u5__abc_81276_new_n3022_));
INVX1 INVX1_109 ( .A(u0_u1__abc_72579_new_n287_), .Y(u0_u1__abc_72579_new_n288_));
INVX1 INVX1_1090 ( .A(u5__abc_81276_new_n2912_), .Y(u5__abc_81276_new_n3034_));
INVX1 INVX1_1091 ( .A(u5__abc_81276_new_n2936_), .Y(u5__abc_81276_new_n3039_));
INVX1 INVX1_1092 ( .A(u5__abc_81276_new_n3029_), .Y(u5__abc_81276_new_n3053_));
INVX1 INVX1_1093 ( .A(u5__abc_81276_new_n2937_), .Y(u5__abc_81276_new_n3062_));
INVX1 INVX1_1094 ( .A(u5__abc_81276_new_n2938_), .Y(u5__abc_81276_new_n3082_));
INVX1 INVX1_1095 ( .A(u5__abc_81276_new_n2948_), .Y(u5__abc_81276_new_n3100_));
INVX1 INVX1_1096 ( .A(u5__abc_81276_new_n2939_), .Y(u5__abc_81276_new_n3102_));
INVX1 INVX1_1097 ( .A(u5__abc_81276_new_n2940_), .Y(u5__abc_81276_new_n3117_));
INVX1 INVX1_1098 ( .A(u5__abc_81276_new_n2941_), .Y(u5__abc_81276_new_n3128_));
INVX1 INVX1_1099 ( .A(u5_ack_cnt_0_), .Y(u5__abc_81276_new_n3143_));
INVX1 INVX1_11 ( .A(u0__abc_76628_new_n4259_), .Y(u0__abc_76628_new_n4268_));
INVX1 INVX1_110 ( .A(\wb_data_i[12] ), .Y(u0_u1__abc_72579_new_n292_));
INVX1 INVX1_1100 ( .A(u5__abc_81276_new_n3145_), .Y(u5__abc_81276_new_n3146_));
INVX1 INVX1_1101 ( .A(u5__abc_81276_new_n3147_), .Y(u5__abc_81276_new_n3148_));
INVX1 INVX1_1102 ( .A(u5_no_wb_cycle), .Y(u5__abc_81276_new_n3150_));
INVX1 INVX1_1103 ( .A(u5__abc_81276_new_n3160_), .Y(u5__abc_81276_new_n3161_));
INVX1 INVX1_1104 ( .A(u5__abc_81276_new_n3166_), .Y(u5__abc_81276_new_n3167_));
INVX1 INVX1_1105 ( .A(u5__abc_81276_new_n1819_), .Y(u5__abc_81276_new_n3172_));
INVX1 INVX1_1106 ( .A(u5__abc_81276_new_n3177_), .Y(u5__abc_81276_new_n3178_));
INVX1 INVX1_1107 ( .A(u5__abc_81276_new_n3181_), .Y(u5__abc_81276_new_n3182_));
INVX1 INVX1_1108 ( .A(mc_br_r), .Y(u5__abc_81276_new_n3208_));
INVX1 INVX1_1109 ( .A(u5__abc_81276_new_n3221_), .Y(u5__abc_81276_new_n3222_));
INVX1 INVX1_111 ( .A(u0_u1__abc_72579_new_n293_), .Y(u0_u1__abc_72579_new_n294_));
INVX1 INVX1_1110 ( .A(u5__abc_81276_new_n3230_), .Y(u5__abc_81276_new_n3231_));
INVX1 INVX1_1111 ( .A(u5__abc_81276_new_n3240_), .Y(u5__abc_81276_new_n3241_));
INVX1 INVX1_1112 ( .A(u5__abc_81276_new_n1615_), .Y(u5__abc_81276_new_n3242_));
INVX1 INVX1_1113 ( .A(u5__abc_81276_new_n3265_), .Y(u5__abc_81276_new_n3266_));
INVX1 INVX1_1114 ( .A(u5__abc_81276_new_n3270_), .Y(u5__abc_81276_new_n3271_));
INVX1 INVX1_1115 ( .A(u5__abc_81276_new_n3229_), .Y(u5__abc_81276_new_n3275_));
INVX1 INVX1_1116 ( .A(u5__abc_81276_new_n1614_), .Y(u5__abc_81276_new_n3283_));
INVX1 INVX1_1117 ( .A(u5__abc_81276_new_n3223_), .Y(u5__abc_81276_new_n3294_));
INVX1 INVX1_1118 ( .A(u5__abc_81276_new_n1728_), .Y(u5__abc_81276_new_n3303_));
INVX1 INVX1_1119 ( .A(row_same), .Y(u5__abc_81276_new_n3304_));
INVX1 INVX1_112 ( .A(\wb_data_i[13] ), .Y(u0_u1__abc_72579_new_n298_));
INVX1 INVX1_1120 ( .A(u5__abc_81276_new_n3325_), .Y(u5__abc_81276_new_n3326_));
INVX1 INVX1_1121 ( .A(u5__abc_81276_new_n3307_), .Y(u5__abc_81276_new_n3327_));
INVX1 INVX1_1122 ( .A(u5__abc_81276_new_n3336_), .Y(u5__abc_81276_new_n3337_));
INVX1 INVX1_1123 ( .A(u5__abc_81276_new_n1851_), .Y(u5__abc_81276_new_n3353_));
INVX1 INVX1_1124 ( .A(u5__abc_81276_new_n3354_), .Y(u5__abc_81276_new_n3355_));
INVX1 INVX1_1125 ( .A(u5__abc_81276_new_n3305_), .Y(u5__abc_81276_new_n3362_));
INVX1 INVX1_1126 ( .A(u5__abc_81276_new_n3390_), .Y(u5__abc_81276_new_n3391_));
INVX1 INVX1_1127 ( .A(u5__abc_81276_new_n3410_), .Y(u5__abc_81276_new_n3411_));
INVX1 INVX1_1128 ( .A(u5__abc_81276_new_n3267_), .Y(u5__abc_81276_new_n3425_));
INVX1 INVX1_1129 ( .A(u5__abc_81276_new_n3282_), .Y(u5__abc_81276_new_n3437_));
INVX1 INVX1_113 ( .A(u0_u1__abc_72579_new_n299_), .Y(u0_u1__abc_72579_new_n300_));
INVX1 INVX1_1130 ( .A(u5__abc_81276_new_n3440_), .Y(u5__abc_81276_new_n3441_));
INVX1 INVX1_1131 ( .A(u5__abc_81276_new_n3243_), .Y(u5__abc_81276_new_n3446_));
INVX1 INVX1_1132 ( .A(u5__abc_81276_new_n3249_), .Y(u5__abc_81276_new_n3447_));
INVX1 INVX1_1133 ( .A(u5__abc_81276_new_n1758_), .Y(u5__abc_81276_new_n3507_));
INVX1 INVX1_1134 ( .A(u5__abc_81276_new_n1398_), .Y(u5__abc_81276_new_n3550_));
INVX1 INVX1_1135 ( .A(u5__abc_81276_new_n3565_), .Y(u5__abc_81276_new_n3566_));
INVX1 INVX1_1136 ( .A(u5_resume_req_r), .Y(u5__abc_81276_new_n3616_));
INVX1 INVX1_1137 ( .A(u5__abc_81276_new_n3210_), .Y(u5__abc_81276_new_n3632_));
INVX1 INVX1_1138 ( .A(u5__abc_81276_new_n1592_), .Y(u5__abc_81276_new_n3653_));
INVX1 INVX1_1139 ( .A(u5__abc_81276_new_n3661_), .Y(u5__abc_81276_new_n3662_));
INVX1 INVX1_114 ( .A(\wb_data_i[14] ), .Y(u0_u1__abc_72579_new_n304_));
INVX1 INVX1_1140 ( .A(u5__abc_81276_new_n3745_), .Y(u5__abc_81276_new_n3752_));
INVX1 INVX1_1141 ( .A(u5__abc_81276_new_n1193_), .Y(u5__abc_81276_new_n3760_));
INVX1 INVX1_1142 ( .A(u5__abc_81276_new_n1194_), .Y(u5__abc_81276_new_n3777_));
INVX1 INVX1_1143 ( .A(u5__abc_81276_new_n3779_), .Y(u5__abc_81276_new_n3780_));
INVX1 INVX1_1144 ( .A(mc_ack_r), .Y(u5__abc_81276_new_n3809_));
INVX1 INVX1_1145 ( .A(u5__abc_81276_new_n2619_), .Y(u5__abc_81276_new_n3840_));
INVX1 INVX1_1146 ( .A(u5__abc_81276_new_n3695_), .Y(u5__abc_81276_new_n3844_));
INVX1 INVX1_1147 ( .A(u5__abc_81276_new_n3845_), .Y(u5__abc_81276_new_n3846_));
INVX1 INVX1_1148 ( .A(u5__abc_81276_new_n3855_), .Y(u5__abc_81276_new_n3856_));
INVX1 INVX1_1149 ( .A(u5__abc_81276_new_n3865_), .Y(u5__abc_81276_new_n3866_));
INVX1 INVX1_115 ( .A(u0_u1__abc_72579_new_n305_), .Y(u0_u1__abc_72579_new_n306_));
INVX1 INVX1_1150 ( .A(u5__abc_81276_new_n3872_), .Y(u5__abc_81276_new_n3873_));
INVX1 INVX1_1151 ( .A(u5__abc_81276_new_n1354_), .Y(u5__abc_81276_new_n3875_));
INVX1 INVX1_1152 ( .A(u5__abc_81276_new_n3196_), .Y(u5__abc_81276_new_n3885_));
INVX1 INVX1_1153 ( .A(lmr_req), .Y(u5__abc_81276_new_n3890_));
INVX1 INVX1_1154 ( .A(u5_susp_req_r), .Y(u5__abc_81276_new_n3891_));
INVX1 INVX1_1155 ( .A(u5__abc_81276_new_n3299_), .Y(u5__abc_81276_new_n3905_));
INVX1 INVX1_1156 ( .A(u5__abc_81276_new_n1559_), .Y(u5__abc_81276_new_n3927_));
INVX1 INVX1_1157 ( .A(u5__abc_81276_new_n1348_), .Y(u5__abc_81276_new_n3930_));
INVX1 INVX1_1158 ( .A(u5__abc_81276_new_n1800_), .Y(u5__abc_81276_new_n3931_));
INVX1 INVX1_1159 ( .A(u5__abc_81276_new_n3897_), .Y(u5__abc_81276_new_n3932_));
INVX1 INVX1_116 ( .A(\wb_data_i[15] ), .Y(u0_u1__abc_72579_new_n310_));
INVX1 INVX1_1160 ( .A(u5__abc_81276_new_n1520_), .Y(u5__abc_81276_new_n3933_));
INVX1 INVX1_1161 ( .A(u5__abc_81276_new_n3896_), .Y(u5__abc_81276_new_n3937_));
INVX1 INVX1_1162 ( .A(u5__abc_81276_new_n2459_), .Y(u5__abc_81276_new_n3940_));
INVX1 INVX1_1163 ( .A(u5__abc_81276_new_n2490_), .Y(u5__abc_81276_new_n3941_));
INVX1 INVX1_1164 ( .A(u5__abc_81276_new_n1645_), .Y(u5__abc_81276_new_n3954_));
INVX1 INVX1_1165 ( .A(rfr_ack), .Y(u5__abc_81276_new_n3957_));
INVX1 INVX1_1166 ( .A(u5__abc_81276_new_n4001_), .Y(u5__abc_81276_new_n4002_));
INVX1 INVX1_1167 ( .A(u5__abc_81276_new_n1733_), .Y(u5__abc_81276_new_n4005_));
INVX1 INVX1_1168 ( .A(u5__abc_81276_new_n4011_), .Y(u5__abc_81276_new_n4012_));
INVX1 INVX1_1169 ( .A(u5__abc_81276_new_n4016_), .Y(u5__abc_81276_new_n4017_));
INVX1 INVX1_117 ( .A(u0_u1__abc_72579_new_n311_), .Y(u0_u1__abc_72579_new_n312_));
INVX1 INVX1_1170 ( .A(u5__abc_81276_new_n4018_), .Y(u5__abc_81276_new_n4019_));
INVX1 INVX1_1171 ( .A(u5__abc_81276_new_n4024_), .Y(cmd_a10));
INVX1 INVX1_1172 ( .A(u5__abc_81276_new_n1695_), .Y(u5__abc_81276_new_n4026_));
INVX1 INVX1_1173 ( .A(u5__abc_81276_new_n3746_), .Y(u5__abc_81276_new_n4027_));
INVX1 INVX1_1174 ( .A(u5__abc_81276_new_n4046_), .Y(u5__abc_81276_new_n4047_));
INVX1 INVX1_1175 ( .A(u5__abc_81276_new_n2533_), .Y(u5__abc_81276_new_n4052_));
INVX1 INVX1_1176 ( .A(u5__abc_81276_new_n1787_), .Y(u5__abc_81276_new_n4053_));
INVX1 INVX1_1177 ( .A(u5__abc_81276_new_n1796_), .Y(u5__abc_81276_new_n4054_));
INVX1 INVX1_1178 ( .A(u5__abc_81276_new_n2942_), .Y(u5__abc_81276_new_n4064_));
INVX1 INVX1_1179 ( .A(u5__abc_81276_new_n2467_), .Y(u5__abc_81276_new_n4071_));
INVX1 INVX1_118 ( .A(\wb_data_i[16] ), .Y(u0_u1__abc_72579_new_n316_));
INVX1 INVX1_1180 ( .A(u5__abc_81276_new_n2460_), .Y(u5__abc_81276_new_n4072_));
INVX1 INVX1_1181 ( .A(u5__abc_81276_new_n2522_), .Y(u5__abc_81276_new_n4073_));
INVX1 INVX1_1182 ( .A(u5__abc_81276_new_n1773_), .Y(u5__abc_81276_new_n4074_));
INVX1 INVX1_1183 ( .A(u5__abc_81276_new_n2452_), .Y(u5__abc_81276_new_n4075_));
INVX1 INVX1_1184 ( .A(not_mem_cyc), .Y(u5__abc_81276_new_n4082_));
INVX1 INVX1_1185 ( .A(u5__abc_81276_new_n1571_), .Y(u5__abc_81276_new_n4087_));
INVX1 INVX1_1186 ( .A(u5_rsts), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_72182));
INVX1 INVX1_1187 ( .A(u6__abc_85257_new_n133_), .Y(u6__abc_85257_new_n134_));
INVX1 INVX1_1188 ( .A(u0_wp_err), .Y(u6__abc_85257_new_n135_));
INVX1 INVX1_1189 ( .A(err), .Y(u6__abc_85257_new_n136_));
INVX1 INVX1_119 ( .A(u0_u1__abc_72579_new_n317_), .Y(u0_u1__abc_72579_new_n318_));
INVX1 INVX1_1190 ( .A(par_err), .Y(u6__abc_85257_new_n137_));
INVX1 INVX1_1191 ( .A(\wb_addr_i[31] ), .Y(u6__abc_85257_new_n141_));
INVX1 INVX1_1192 ( .A(\wb_addr_i[30] ), .Y(u6__abc_85257_new_n142_));
INVX1 INVX1_1193 ( .A(\wb_addr_i[29] ), .Y(u6__abc_85257_new_n143_));
INVX1 INVX1_1194 ( .A(_auto_iopadmap_cc_368_execute_85558), .Y(u6__abc_85257_new_n149_));
INVX1 INVX1_1195 ( .A(u1_wr_hold), .Y(u6__abc_85257_new_n254_));
INVX1 INVX1_1196 ( .A(wb_we_i), .Y(u6__abc_85257_new_n257_));
INVX1 INVX1_1197 ( .A(u6_rmw_r), .Y(u6__abc_85257_new_n261_));
INVX1 INVX1_1198 ( .A(u6__0rmw_r_0_0_), .Y(u6__abc_85257_new_n262_));
INVX1 INVX1_1199 ( .A(wb_stb_i_bF_buf1), .Y(u6__abc_85257_new_n271_));
INVX1 INVX1_12 ( .A(u0__abc_76628_new_n4395_), .Y(u0__abc_76628_new_n4396_));
INVX1 INVX1_120 ( .A(\wb_data_i[17] ), .Y(u0_u1__abc_72579_new_n322_));
INVX1 INVX1_1200 ( .A(u6_read_go_r), .Y(u6__abc_85257_new_n276_));
INVX1 INVX1_1201 ( .A(u6_write_go_r), .Y(u6__abc_85257_new_n277_));
INVX1 INVX1_1202 ( .A(_auto_iopadmap_cc_368_execute_85593), .Y(u6__abc_85257_new_n281_));
INVX1 INVX1_1203 ( .A(u6__abc_85257_new_n140_), .Y(u6__abc_85257_new_n285_));
INVX1 INVX1_1204 ( .A(u7_mc_dqm_r2_0_), .Y(u7__abc_74830_new_n75_));
INVX1 INVX1_1205 ( .A(data_oe), .Y(u7__abc_74830_new_n77_));
INVX1 INVX1_1206 ( .A(u5_wb_cycle), .Y(u7__abc_74830_new_n78_));
INVX1 INVX1_1207 ( .A(u7_mc_dqm_r2_1_), .Y(u7__abc_74830_new_n83_));
INVX1 INVX1_1208 ( .A(u7_mc_dqm_r2_2_), .Y(u7__abc_74830_new_n86_));
INVX1 INVX1_1209 ( .A(u7_mc_dqm_r2_3_), .Y(u7__abc_74830_new_n89_));
INVX1 INVX1_121 ( .A(u0_u1__abc_72579_new_n323_), .Y(u0_u1__abc_72579_new_n324_));
INVX1 INVX1_1210 ( .A(u7__abc_74830_new_n92_), .Y(u7__abc_74830_new_n94_));
INVX1 INVX1_1211 ( .A(cs_0_), .Y(u7__abc_74830_new_n108_));
INVX1 INVX1_1212 ( .A(u7__abc_74830_new_n110_), .Y(u7__abc_74830_new_n111_));
INVX1 INVX1_1213 ( .A(cs_need_rfr_0_), .Y(u7__abc_74830_new_n115_));
INVX1 INVX1_1214 ( .A(cs_1_), .Y(u7__abc_74830_new_n119_));
INVX1 INVX1_1215 ( .A(u7__abc_74830_new_n121_), .Y(u7__abc_74830_new_n122_));
INVX1 INVX1_1216 ( .A(cs_need_rfr_1_), .Y(u7__abc_74830_new_n125_));
INVX1 INVX1_1217 ( .A(cs_2_), .Y(u7__abc_74830_new_n129_));
INVX1 INVX1_1218 ( .A(u7__abc_74830_new_n131_), .Y(u7__abc_74830_new_n132_));
INVX1 INVX1_1219 ( .A(cs_need_rfr_2_), .Y(u7__abc_74830_new_n135_));
INVX1 INVX1_122 ( .A(\wb_data_i[18] ), .Y(u0_u1__abc_72579_new_n328_));
INVX1 INVX1_1220 ( .A(cs_3_), .Y(u7__abc_74830_new_n139_));
INVX1 INVX1_1221 ( .A(u7__abc_74830_new_n141_), .Y(u7__abc_74830_new_n142_));
INVX1 INVX1_1222 ( .A(cs_need_rfr_3_), .Y(u7__abc_74830_new_n145_));
INVX1 INVX1_1223 ( .A(cs_4_), .Y(u7__abc_74830_new_n149_));
INVX1 INVX1_1224 ( .A(u7__abc_74830_new_n151_), .Y(u7__abc_74830_new_n152_));
INVX1 INVX1_1225 ( .A(cs_need_rfr_4_), .Y(u7__abc_74830_new_n155_));
INVX1 INVX1_1226 ( .A(cs_5_), .Y(u7__abc_74830_new_n159_));
INVX1 INVX1_1227 ( .A(u7__abc_74830_new_n161_), .Y(u7__abc_74830_new_n162_));
INVX1 INVX1_1228 ( .A(cs_need_rfr_5_), .Y(u7__abc_74830_new_n165_));
INVX1 INVX1_1229 ( .A(cs_6_), .Y(u7__abc_74830_new_n169_));
INVX1 INVX1_123 ( .A(u0_u1__abc_72579_new_n329_), .Y(u0_u1__abc_72579_new_n330_));
INVX1 INVX1_1230 ( .A(u7__abc_74830_new_n171_), .Y(u7__abc_74830_new_n172_));
INVX1 INVX1_1231 ( .A(cs_need_rfr_6_), .Y(u7__abc_74830_new_n175_));
INVX1 INVX1_1232 ( .A(cs_7_), .Y(u7__abc_74830_new_n179_));
INVX1 INVX1_1233 ( .A(u7__abc_74830_new_n181_), .Y(u7__abc_74830_new_n182_));
INVX1 INVX1_1234 ( .A(cs_need_rfr_7_), .Y(u7__abc_74830_new_n185_));
INVX1 INVX1_1235 ( .A(mc_adsc_d), .Y(u7__0mc_adsc__0_0_));
INVX1 INVX1_1236 ( .A(mc_adv_d), .Y(u7__0mc_adv__0_0_));
INVX1 INVX1_1237 ( .A(fs), .Y(u7__abc_74830_new_n191_));
INVX1 INVX1_1238 ( .A(_auto_iopadmap_cc_368_execute_85556), .Y(u7__abc_74830_new_n192_));
INVX1 INVX1_1239 ( .A(susp_sel), .Y(u7__abc_74830_new_n194_));
INVX1 INVX1_124 ( .A(\wb_data_i[19] ), .Y(u0_u1__abc_72579_new_n334_));
INVX1 INVX1_125 ( .A(u0_u1__abc_72579_new_n335_), .Y(u0_u1__abc_72579_new_n336_));
INVX1 INVX1_126 ( .A(\wb_data_i[20] ), .Y(u0_u1__abc_72579_new_n340_));
INVX1 INVX1_127 ( .A(u0_u1__abc_72579_new_n341_), .Y(u0_u1__abc_72579_new_n342_));
INVX1 INVX1_128 ( .A(\wb_data_i[21] ), .Y(u0_u1__abc_72579_new_n346_));
INVX1 INVX1_129 ( .A(u0_u1__abc_72579_new_n347_), .Y(u0_u1__abc_72579_new_n348_));
INVX1 INVX1_13 ( .A(u0_rf_we), .Y(u0__abc_76628_new_n4397_));
INVX1 INVX1_130 ( .A(\wb_data_i[22] ), .Y(u0_u1__abc_72579_new_n352_));
INVX1 INVX1_131 ( .A(u0_u1__abc_72579_new_n353_), .Y(u0_u1__abc_72579_new_n354_));
INVX1 INVX1_132 ( .A(\wb_data_i[23] ), .Y(u0_u1__abc_72579_new_n358_));
INVX1 INVX1_133 ( .A(u0_u1__abc_72579_new_n359_), .Y(u0_u1__abc_72579_new_n360_));
INVX1 INVX1_134 ( .A(\wb_data_i[24] ), .Y(u0_u1__abc_72579_new_n364_));
INVX1 INVX1_135 ( .A(u0_u1__abc_72579_new_n365_), .Y(u0_u1__abc_72579_new_n366_));
INVX1 INVX1_136 ( .A(\wb_data_i[25] ), .Y(u0_u1__abc_72579_new_n370_));
INVX1 INVX1_137 ( .A(u0_u1__abc_72579_new_n371_), .Y(u0_u1__abc_72579_new_n372_));
INVX1 INVX1_138 ( .A(\wb_data_i[26] ), .Y(u0_u1__abc_72579_new_n376_));
INVX1 INVX1_139 ( .A(u0_u1__abc_72579_new_n377_), .Y(u0_u1__abc_72579_new_n378_));
INVX1 INVX1_14 ( .A(u0__abc_76628_new_n4398_), .Y(u0__abc_76628_new_n4399_));
INVX1 INVX1_140 ( .A(\wb_data_i[27] ), .Y(u0_u1__abc_72579_new_n382_));
INVX1 INVX1_141 ( .A(u0_u1__abc_72579_new_n383_), .Y(u0_u1__abc_72579_new_n384_));
INVX1 INVX1_142 ( .A(\wb_data_i[28] ), .Y(u0_u1__abc_72579_new_n388_));
INVX1 INVX1_143 ( .A(u0_u1__abc_72579_new_n389_), .Y(u0_u1__abc_72579_new_n390_));
INVX1 INVX1_144 ( .A(\wb_data_i[29] ), .Y(u0_u1__abc_72579_new_n394_));
INVX1 INVX1_145 ( .A(u0_u1__abc_72579_new_n395_), .Y(u0_u1__abc_72579_new_n396_));
INVX1 INVX1_146 ( .A(\wb_data_i[30] ), .Y(u0_u1__abc_72579_new_n400_));
INVX1 INVX1_147 ( .A(u0_u1__abc_72579_new_n401_), .Y(u0_u1__abc_72579_new_n402_));
INVX1 INVX1_148 ( .A(\wb_data_i[31] ), .Y(u0_u1__abc_72579_new_n406_));
INVX1 INVX1_149 ( .A(u0_u1__abc_72579_new_n407_), .Y(u0_u1__abc_72579_new_n408_));
INVX1 INVX1_15 ( .A(\wb_addr_i[5] ), .Y(u0__abc_76628_new_n4493_));
INVX1 INVX1_150 ( .A(u0_u1_addr_r_2_), .Y(u0_u1__abc_72579_new_n411_));
INVX1 INVX1_151 ( .A(u0_u1__abc_72579_new_n414_), .Y(u0_u1__abc_72579_new_n415_));
INVX1 INVX1_152 ( .A(u0_u1__abc_72579_new_n419_), .Y(u0_u1__abc_72579_new_n420_));
INVX1 INVX1_153 ( .A(u0_u1__abc_72579_new_n424_), .Y(u0_u1__abc_72579_new_n425_));
INVX1 INVX1_154 ( .A(u0_u1__abc_72579_new_n429_), .Y(u0_u1__abc_72579_new_n430_));
INVX1 INVX1_155 ( .A(u0_u1__abc_72579_new_n434_), .Y(u0_u1__abc_72579_new_n435_));
INVX1 INVX1_156 ( .A(u0_u1__abc_72579_new_n439_), .Y(u0_u1__abc_72579_new_n440_));
INVX1 INVX1_157 ( .A(u0_u1__abc_72579_new_n444_), .Y(u0_u1__abc_72579_new_n445_));
INVX1 INVX1_158 ( .A(u0_u1__abc_72579_new_n449_), .Y(u0_u1__abc_72579_new_n450_));
INVX1 INVX1_159 ( .A(u0_u1__abc_72579_new_n454_), .Y(u0_u1__abc_72579_new_n455_));
INVX1 INVX1_16 ( .A(\wb_addr_i[4] ), .Y(u0__abc_76628_new_n4494_));
INVX1 INVX1_160 ( .A(u0_u1__abc_72579_new_n459_), .Y(u0_u1__abc_72579_new_n460_));
INVX1 INVX1_161 ( .A(u0_u1__abc_72579_new_n464_), .Y(u0_u1__abc_72579_new_n465_));
INVX1 INVX1_162 ( .A(u0_u1__abc_72579_new_n469_), .Y(u0_u1__abc_72579_new_n470_));
INVX1 INVX1_163 ( .A(u0_u1__abc_72579_new_n474_), .Y(u0_u1__abc_72579_new_n475_));
INVX1 INVX1_164 ( .A(u0_u1__abc_72579_new_n479_), .Y(u0_u1__abc_72579_new_n480_));
INVX1 INVX1_165 ( .A(u0_u1__abc_72579_new_n484_), .Y(u0_u1__abc_72579_new_n485_));
INVX1 INVX1_166 ( .A(u0_u1__abc_72579_new_n489_), .Y(u0_u1__abc_72579_new_n490_));
INVX1 INVX1_167 ( .A(u0_u1__abc_72579_new_n494_), .Y(u0_u1__abc_72579_new_n495_));
INVX1 INVX1_168 ( .A(u0_u1__abc_72579_new_n499_), .Y(u0_u1__abc_72579_new_n500_));
INVX1 INVX1_169 ( .A(u0_u1__abc_72579_new_n504_), .Y(u0_u1__abc_72579_new_n505_));
INVX1 INVX1_17 ( .A(\wb_addr_i[3] ), .Y(u0__abc_76628_new_n4497_));
INVX1 INVX1_170 ( .A(u0_u1__abc_72579_new_n509_), .Y(u0_u1__abc_72579_new_n510_));
INVX1 INVX1_171 ( .A(u0_u1__abc_72579_new_n514_), .Y(u0_u1__abc_72579_new_n515_));
INVX1 INVX1_172 ( .A(u0_u1__abc_72579_new_n519_), .Y(u0_u1__abc_72579_new_n520_));
INVX1 INVX1_173 ( .A(u0_u1__abc_72579_new_n524_), .Y(u0_u1__abc_72579_new_n525_));
INVX1 INVX1_174 ( .A(u0_u1__abc_72579_new_n529_), .Y(u0_u1__abc_72579_new_n530_));
INVX1 INVX1_175 ( .A(u0_u1__abc_72579_new_n534_), .Y(u0_u1__abc_72579_new_n535_));
INVX1 INVX1_176 ( .A(u0_u1__abc_72579_new_n539_), .Y(u0_u1__abc_72579_new_n540_));
INVX1 INVX1_177 ( .A(u0_u1__abc_72579_new_n544_), .Y(u0_u1__abc_72579_new_n545_));
INVX1 INVX1_178 ( .A(u0_u1__abc_72579_new_n549_), .Y(u0_u1__abc_72579_new_n550_));
INVX1 INVX1_179 ( .A(u0_u1__abc_72579_new_n554_), .Y(u0_u1__abc_72579_new_n555_));
INVX1 INVX1_18 ( .A(\wb_addr_i[2] ), .Y(u0__abc_76628_new_n4498_));
INVX1 INVX1_180 ( .A(u0_u1__abc_72579_new_n559_), .Y(u0_u1__abc_72579_new_n560_));
INVX1 INVX1_181 ( .A(u0_u1__abc_72579_new_n564_), .Y(u0_u1__abc_72579_new_n565_));
INVX1 INVX1_182 ( .A(u0_u1__abc_72579_new_n569_), .Y(u0_u1__abc_72579_new_n570_));
INVX1 INVX1_183 ( .A(u0_csc1_23_), .Y(u0_u1__abc_72579_new_n574_));
INVX1 INVX1_184 ( .A(\wb_addr_i[28] ), .Y(u0_u1__abc_72579_new_n575_));
INVX1 INVX1_185 ( .A(u0_csc_mask_7_), .Y(u0_u1__abc_72579_new_n577_));
INVX1 INVX1_186 ( .A(u0_csc_mask_6_), .Y(u0_u1__abc_72579_new_n582_));
INVX1 INVX1_187 ( .A(u0_csc1_22_), .Y(u0_u1__abc_72579_new_n583_));
INVX1 INVX1_188 ( .A(\wb_addr_i[27] ), .Y(u0_u1__abc_72579_new_n584_));
INVX1 INVX1_189 ( .A(u0_csc_mask_5_), .Y(u0_u1__abc_72579_new_n590_));
INVX1 INVX1_19 ( .A(u0__abc_76628_new_n4495_), .Y(u0__abc_76628_new_n4536_));
INVX1 INVX1_190 ( .A(u0_csc1_21_), .Y(u0_u1__abc_72579_new_n591_));
INVX1 INVX1_191 ( .A(\wb_addr_i[26] ), .Y(u0_u1__abc_72579_new_n592_));
INVX1 INVX1_192 ( .A(u0_csc_mask_0_), .Y(u0_u1__abc_72579_new_n598_));
INVX1 INVX1_193 ( .A(u0_csc1_16_), .Y(u0_u1__abc_72579_new_n599_));
INVX1 INVX1_194 ( .A(\wb_addr_i[21] ), .Y(u0_u1__abc_72579_new_n600_));
INVX1 INVX1_195 ( .A(u0_u1__abc_72579_new_n605_), .Y(u0_u1__abc_72579_new_n606_));
INVX1 INVX1_196 ( .A(u0_u1__abc_72579_new_n607_), .Y(u0_u1__abc_72579_new_n609_));
INVX1 INVX1_197 ( .A(u0_u1__abc_72579_new_n612_), .Y(u0_u1__abc_72579_new_n613_));
INVX1 INVX1_198 ( .A(u0_u1__abc_72579_new_n614_), .Y(u0_u1__abc_72579_new_n616_));
INVX1 INVX1_199 ( .A(u0_u1__abc_72579_new_n620_), .Y(u0_u1__abc_72579_new_n621_));
INVX1 INVX1_2 ( .A(lmr_ack), .Y(_abc_85006_new_n239_));
INVX1 INVX1_20 ( .A(\wb_addr_i[31] ), .Y(u0__abc_76628_new_n5652_));
INVX1 INVX1_200 ( .A(u0_u1__abc_72579_new_n622_), .Y(u0_u1__abc_72579_new_n624_));
INVX1 INVX1_201 ( .A(u0_u1__abc_72579_new_n627_), .Y(u0_u1__abc_72579_new_n628_));
INVX1 INVX1_202 ( .A(u0_u1__abc_72579_new_n629_), .Y(u0_u1__abc_72579_new_n631_));
INVX1 INVX1_203 ( .A(u0_u1__abc_72579_new_n573_), .Y(u0_u1__abc_72579_new_n639_));
INVX1 INVX1_204 ( .A(u0_init_ack1), .Y(u0_u1__abc_72579_new_n642_));
INVX1 INVX1_205 ( .A(u0_u1_inited), .Y(u0_u1__abc_72579_new_n644_));
INVX1 INVX1_206 ( .A(csc_s_4_), .Y(u1__abc_73140_new_n261_));
INVX1 INVX1_207 ( .A(csc_s_6_), .Y(u1__abc_73140_new_n263_));
INVX1 INVX1_208 ( .A(csc_s_5_), .Y(u1__abc_73140_new_n267_));
INVX1 INVX1_209 ( .A(u1__abc_73140_new_n270_), .Y(u1__abc_73140_new_n271_));
INVX1 INVX1_21 ( .A(u0_csc0_1_), .Y(u0__abc_76628_new_n5660_));
INVX1 INVX1_210 ( .A(u1__abc_73140_new_n259_), .Y(u1__abc_73140_new_n273_));
INVX1 INVX1_211 ( .A(u1__abc_73140_new_n276_), .Y(u1__abc_73140_new_n277_));
INVX1 INVX1_212 ( .A(page_size_8_), .Y(u1__abc_73140_new_n280_));
INVX1 INVX1_213 ( .A(u1__abc_73140_new_n266_), .Y(u1__abc_73140_new_n291_));
INVX1 INVX1_214 ( .A(u1__abc_73140_new_n293_), .Y(u1__abc_73140_new_n294_));
INVX1 INVX1_215 ( .A(u1__abc_73140_new_n275__bF_buf2), .Y(u1__abc_73140_new_n295_));
INVX1 INVX1_216 ( .A(csc_s_7_), .Y(u1__abc_73140_new_n298_));
INVX1 INVX1_217 ( .A(u1__abc_73140_new_n301_), .Y(u1__abc_73140_new_n302_));
INVX1 INVX1_218 ( .A(u1__abc_73140_new_n258_), .Y(u1__abc_73140_new_n303_));
INVX1 INVX1_219 ( .A(u1__abc_73140_new_n304_), .Y(u1__abc_73140_new_n305_));
INVX1 INVX1_22 ( .A(u0_csc0_2_), .Y(u0__abc_76628_new_n5661_));
INVX1 INVX1_220 ( .A(u1__abc_73140_new_n358_), .Y(u1__abc_73140_new_n359_));
INVX1 INVX1_221 ( .A(u1__abc_73140_new_n360_), .Y(u1__abc_73140_new_n361_));
INVX1 INVX1_222 ( .A(u1_wr_cycle), .Y(u1__abc_73140_new_n524_));
INVX1 INVX1_223 ( .A(u1__abc_73140_new_n898_), .Y(u1__abc_73140_new_n899_));
INVX1 INVX1_224 ( .A(u1__abc_73140_new_n901_), .Y(u1__abc_73140_new_n902_));
INVX1 INVX1_225 ( .A(csc_s_2_), .Y(u1__abc_73140_new_n910_));
INVX1 INVX1_226 ( .A(cas_), .Y(u1__abc_73140_new_n917_));
INVX1 INVX1_227 ( .A(u1_u0__abc_73035_new_n51_), .Y(u1_u0__abc_73035_new_n52_));
INVX1 INVX1_228 ( .A(u1_u0__abc_73035_new_n55_), .Y(u1_u0__abc_73035_new_n56_));
INVX1 INVX1_229 ( .A(u1_u0__abc_73035_new_n59_), .Y(u1_u0__abc_73035_new_n60_));
INVX1 INVX1_23 ( .A(u0_csc0_3_), .Y(u0__abc_76628_new_n5663_));
INVX1 INVX1_230 ( .A(u1_u0__abc_73035_new_n63_), .Y(u1_u0__abc_73035_new_n64_));
INVX1 INVX1_231 ( .A(u1_u0__abc_73035_new_n69_), .Y(u1_u0__abc_73035_new_n70_));
INVX1 INVX1_232 ( .A(u1_u0__abc_73035_new_n72_), .Y(u1_u0__abc_73035_new_n73_));
INVX1 INVX1_233 ( .A(u1_u0__abc_73035_new_n79_), .Y(u1_u0__abc_73035_new_n80_));
INVX1 INVX1_234 ( .A(u1_u0__abc_73035_new_n82_), .Y(u1_u0__abc_73035_new_n83_));
INVX1 INVX1_235 ( .A(u1_u0__abc_73035_new_n88_), .Y(u1_u0__abc_73035_new_n89_));
INVX1 INVX1_236 ( .A(u1_u0__abc_73035_new_n91_), .Y(u1_u0__abc_73035_new_n92_));
INVX1 INVX1_237 ( .A(u1_u0__0out_r_12_0__12_), .Y(u1_u0__abc_73035_new_n98_));
INVX1 INVX1_238 ( .A(u1_acs_addr_0_), .Y(u1_u0__0out_r_12_0__0_));
INVX1 INVX1_239 ( .A(u1_u0__abc_73035_new_n103_), .Y(u1_u0__abc_73035_new_n104_));
INVX1 INVX1_24 ( .A(u0_csc1_1_), .Y(u0__abc_76628_new_n5666_));
INVX1 INVX1_240 ( .A(u1_u0__abc_73035_new_n107_), .Y(u1_u0__abc_73035_new_n108_));
INVX1 INVX1_241 ( .A(u1_u0__abc_73035_new_n113_), .Y(u1_u0__abc_73035_new_n114_));
INVX1 INVX1_242 ( .A(u1_u0__abc_73035_new_n116_), .Y(u1_u0__abc_73035_new_n117_));
INVX1 INVX1_243 ( .A(u1_u0__abc_73035_new_n122_), .Y(u1_u0__abc_73035_new_n123_));
INVX1 INVX1_244 ( .A(u1_u0__abc_73035_new_n125_), .Y(u1_u0__abc_73035_new_n126_));
INVX1 INVX1_245 ( .A(u1_u0__abc_73035_new_n132_), .Y(u1_u0__abc_73035_new_n133_));
INVX1 INVX1_246 ( .A(u1_u0__abc_73035_new_n135_), .Y(u1_u0__abc_73035_new_n136_));
INVX1 INVX1_247 ( .A(u1_u0__abc_73035_new_n141_), .Y(u1_u0__abc_73035_new_n142_));
INVX1 INVX1_248 ( .A(u1_u0__abc_73035_new_n144_), .Y(u1_u0__abc_73035_new_n145_));
INVX1 INVX1_249 ( .A(u1_u0__abc_73035_new_n149_), .Y(u1_u0__abc_73035_new_n150_));
INVX1 INVX1_25 ( .A(u0_csc1_2_), .Y(u0__abc_76628_new_n5667_));
INVX1 INVX1_250 ( .A(u1_u0__abc_73035_new_n102_), .Y(u1_u0__abc_73035_new_n152_));
INVX1 INVX1_251 ( .A(u2_u0__abc_74955_new_n140_), .Y(u2_u0__abc_74955_new_n141_));
INVX1 INVX1_252 ( .A(u2_u0__abc_74955_new_n145_), .Y(u2_u0__abc_74955_new_n146_));
INVX1 INVX1_253 ( .A(u2_u0__abc_74955_new_n150_), .Y(u2_u0__abc_74955_new_n151_));
INVX1 INVX1_254 ( .A(u2_u0__abc_74955_new_n155_), .Y(u2_u0__abc_74955_new_n156_));
INVX1 INVX1_255 ( .A(u2_u0__abc_74955_new_n160_), .Y(u2_u0__abc_74955_new_n161_));
INVX1 INVX1_256 ( .A(u2_u0__abc_74955_new_n165_), .Y(u2_u0__abc_74955_new_n166_));
INVX1 INVX1_257 ( .A(u2_u0__abc_74955_new_n170_), .Y(u2_u0__abc_74955_new_n171_));
INVX1 INVX1_258 ( .A(u2_u0__abc_74955_new_n175_), .Y(u2_u0__abc_74955_new_n176_));
INVX1 INVX1_259 ( .A(u2_u0__abc_74955_new_n180_), .Y(u2_u0__abc_74955_new_n181_));
INVX1 INVX1_26 ( .A(u0_csc1_3_), .Y(u0__abc_76628_new_n5669_));
INVX1 INVX1_260 ( .A(u2_u0__abc_74955_new_n185_), .Y(u2_u0__abc_74955_new_n186_));
INVX1 INVX1_261 ( .A(u2_u0__abc_74955_new_n190_), .Y(u2_u0__abc_74955_new_n191_));
INVX1 INVX1_262 ( .A(u2_u0__abc_74955_new_n195_), .Y(u2_u0__abc_74955_new_n196_));
INVX1 INVX1_263 ( .A(u2_u0__abc_74955_new_n200_), .Y(u2_u0__abc_74955_new_n201_));
INVX1 INVX1_264 ( .A(bank_adr_0_), .Y(u2_u0__abc_74955_new_n203_));
INVX1 INVX1_265 ( .A(bank_adr_1_), .Y(u2_u0__abc_74955_new_n204_));
INVX1 INVX1_266 ( .A(u2_u0_b3_last_row_9_), .Y(u2_u0__abc_74955_new_n332_));
INVX1 INVX1_267 ( .A(u2_u0_b3_last_row_8_), .Y(u2_u0__abc_74955_new_n334_));
INVX1 INVX1_268 ( .A(u2_u0_b3_last_row_11_), .Y(u2_u0__abc_74955_new_n339_));
INVX1 INVX1_269 ( .A(u2_u0_b3_last_row_4_), .Y(u2_u0__abc_74955_new_n342_));
INVX1 INVX1_27 ( .A(1'h0), .Y(u0__abc_76628_new_n5672_));
INVX1 INVX1_270 ( .A(u2_u0_b3_last_row_0_), .Y(u2_u0__abc_74955_new_n348_));
INVX1 INVX1_271 ( .A(u2_u0_b3_last_row_7_), .Y(u2_u0__abc_74955_new_n355_));
INVX1 INVX1_272 ( .A(u2_u0_b3_last_row_5_), .Y(u2_u0__abc_74955_new_n359_));
INVX1 INVX1_273 ( .A(u2_u0_b3_last_row_12_), .Y(u2_u0__abc_74955_new_n367_));
INVX1 INVX1_274 ( .A(u2_u0_b3_last_row_10_), .Y(u2_u0__abc_74955_new_n371_));
INVX1 INVX1_275 ( .A(u2_u0_b3_last_row_3_), .Y(u2_u0__abc_74955_new_n375_));
INVX1 INVX1_276 ( .A(u2_u0_b3_last_row_1_), .Y(u2_u0__abc_74955_new_n379_));
INVX1 INVX1_277 ( .A(u2_u0_b3_last_row_6_), .Y(u2_u0__abc_74955_new_n385_));
INVX1 INVX1_278 ( .A(u2_u0_b3_last_row_2_), .Y(u2_u0__abc_74955_new_n388_));
INVX1 INVX1_279 ( .A(u2_u0_b1_last_row_0_), .Y(u2_u0__abc_74955_new_n399_));
INVX1 INVX1_28 ( .A(1'h0), .Y(u0__abc_76628_new_n5673_));
INVX1 INVX1_280 ( .A(u2_u0_b1_last_row_4_), .Y(u2_u0__abc_74955_new_n403_));
INVX1 INVX1_281 ( .A(u2_u0_b1_last_row_3_), .Y(u2_u0__abc_74955_new_n407_));
INVX1 INVX1_282 ( .A(u2_u0_b1_last_row_8_), .Y(u2_u0__abc_74955_new_n413_));
INVX1 INVX1_283 ( .A(u2_u0_b1_last_row_6_), .Y(u2_u0__abc_74955_new_n417_));
INVX1 INVX1_284 ( .A(u2_u0_b1_last_row_12_), .Y(u2_u0__abc_74955_new_n422_));
INVX1 INVX1_285 ( .A(u2_u0_b1_last_row_11_), .Y(u2_u0__abc_74955_new_n425_));
INVX1 INVX1_286 ( .A(u2_u0_b1_last_row_2_), .Y(u2_u0__abc_74955_new_n431_));
INVX1 INVX1_287 ( .A(u2_u0_b1_last_row_1_), .Y(u2_u0__abc_74955_new_n435_));
INVX1 INVX1_288 ( .A(u2_u0_b1_last_row_10_), .Y(u2_u0__abc_74955_new_n440_));
INVX1 INVX1_289 ( .A(u2_u0_b1_last_row_9_), .Y(u2_u0__abc_74955_new_n444_));
INVX1 INVX1_29 ( .A(1'h0), .Y(u0__abc_76628_new_n5675_));
INVX1 INVX1_290 ( .A(u2_u0_b1_last_row_7_), .Y(u2_u0__abc_74955_new_n450_));
INVX1 INVX1_291 ( .A(u2_u0_b1_last_row_5_), .Y(u2_u0__abc_74955_new_n454_));
INVX1 INVX1_292 ( .A(u2_u0_b0_last_row_9_), .Y(u2_u0__abc_74955_new_n462_));
INVX1 INVX1_293 ( .A(u2_u0_b0_last_row_12_), .Y(u2_u0__abc_74955_new_n469_));
INVX1 INVX1_294 ( .A(u2_u0_b0_last_row_3_), .Y(u2_u0__abc_74955_new_n472_));
INVX1 INVX1_295 ( .A(u2_u0_b0_last_row_2_), .Y(u2_u0__abc_74955_new_n477_));
INVX1 INVX1_296 ( .A(u2_u0_b0_last_row_6_), .Y(u2_u0__abc_74955_new_n479_));
INVX1 INVX1_297 ( .A(u2_u0_b0_last_row_0_), .Y(u2_u0__abc_74955_new_n488_));
INVX1 INVX1_298 ( .A(u2_u0_b0_last_row_1_), .Y(u2_u0__abc_74955_new_n492_));
INVX1 INVX1_299 ( .A(u2_u0_b0_last_row_5_), .Y(u2_u0__abc_74955_new_n498_));
INVX1 INVX1_3 ( .A(u0__abc_76628_new_n1103_), .Y(u0__abc_76628_new_n1104_));
INVX1 INVX1_30 ( .A(1'h0), .Y(u0__abc_76628_new_n5678_));
INVX1 INVX1_300 ( .A(u2_u0_b0_last_row_8_), .Y(u2_u0__abc_74955_new_n501_));
INVX1 INVX1_301 ( .A(u2_u0_b0_last_row_4_), .Y(u2_u0__abc_74955_new_n506_));
INVX1 INVX1_302 ( .A(u2_u0_b0_last_row_11_), .Y(u2_u0__abc_74955_new_n508_));
INVX1 INVX1_303 ( .A(u2_u0_b0_last_row_7_), .Y(u2_u0__abc_74955_new_n516_));
INVX1 INVX1_304 ( .A(u2_u0_b0_last_row_10_), .Y(u2_u0__abc_74955_new_n520_));
INVX1 INVX1_305 ( .A(u2_u0_b2_last_row_8_), .Y(u2_u0__abc_74955_new_n527_));
INVX1 INVX1_306 ( .A(u2_u0_b2_last_row_9_), .Y(u2_u0__abc_74955_new_n533_));
INVX1 INVX1_307 ( .A(u2_u0_b2_last_row_11_), .Y(u2_u0__abc_74955_new_n537_));
INVX1 INVX1_308 ( .A(u2_u0_b2_last_row_7_), .Y(u2_u0__abc_74955_new_n544_));
INVX1 INVX1_309 ( .A(u2_u0_b2_last_row_6_), .Y(u2_u0__abc_74955_new_n548_));
INVX1 INVX1_31 ( .A(1'h0), .Y(u0__abc_76628_new_n5679_));
INVX1 INVX1_310 ( .A(u2_u0_b2_last_row_3_), .Y(u2_u0__abc_74955_new_n553_));
INVX1 INVX1_311 ( .A(u2_u0_b2_last_row_2_), .Y(u2_u0__abc_74955_new_n557_));
INVX1 INVX1_312 ( .A(u2_u0_b2_last_row_12_), .Y(u2_u0__abc_74955_new_n563_));
INVX1 INVX1_313 ( .A(u2_u0_b2_last_row_10_), .Y(u2_u0__abc_74955_new_n567_));
INVX1 INVX1_314 ( .A(u2_u0_b2_last_row_4_), .Y(u2_u0__abc_74955_new_n573_));
INVX1 INVX1_315 ( .A(u2_u0_b2_last_row_5_), .Y(u2_u0__abc_74955_new_n577_));
INVX1 INVX1_316 ( .A(u2_u0_b2_last_row_0_), .Y(u2_u0__abc_74955_new_n582_));
INVX1 INVX1_317 ( .A(u2_u0_b2_last_row_1_), .Y(u2_u0__abc_74955_new_n585_));
INVX1 INVX1_318 ( .A(u2_bank_clr_0), .Y(u2_u0__abc_74955_new_n601_));
INVX1 INVX1_319 ( .A(u2_u0__abc_74955_new_n289_), .Y(u2_u0__abc_74955_new_n602_));
INVX1 INVX1_32 ( .A(1'h0), .Y(u0__abc_76628_new_n5681_));
INVX1 INVX1_320 ( .A(u2_bank_clr_all_0), .Y(u2_u0__abc_74955_new_n604_));
INVX1 INVX1_321 ( .A(u2_u0__abc_74955_new_n608_), .Y(u2_u0__abc_74955_new_n609_));
INVX1 INVX1_322 ( .A(u2_u0__abc_74955_new_n247_), .Y(u2_u0__abc_74955_new_n616_));
INVX1 INVX1_323 ( .A(u2_u0__abc_74955_new_n205_), .Y(u2_u0__abc_74955_new_n621_));
INVX1 INVX1_324 ( .A(u2_u1__abc_74955_new_n140_), .Y(u2_u1__abc_74955_new_n141_));
INVX1 INVX1_325 ( .A(u2_u1__abc_74955_new_n145_), .Y(u2_u1__abc_74955_new_n146_));
INVX1 INVX1_326 ( .A(u2_u1__abc_74955_new_n150_), .Y(u2_u1__abc_74955_new_n151_));
INVX1 INVX1_327 ( .A(u2_u1__abc_74955_new_n155_), .Y(u2_u1__abc_74955_new_n156_));
INVX1 INVX1_328 ( .A(u2_u1__abc_74955_new_n160_), .Y(u2_u1__abc_74955_new_n161_));
INVX1 INVX1_329 ( .A(u2_u1__abc_74955_new_n165_), .Y(u2_u1__abc_74955_new_n166_));
INVX1 INVX1_33 ( .A(1'h0), .Y(u0__abc_76628_new_n5684_));
INVX1 INVX1_330 ( .A(u2_u1__abc_74955_new_n170_), .Y(u2_u1__abc_74955_new_n171_));
INVX1 INVX1_331 ( .A(u2_u1__abc_74955_new_n175_), .Y(u2_u1__abc_74955_new_n176_));
INVX1 INVX1_332 ( .A(u2_u1__abc_74955_new_n180_), .Y(u2_u1__abc_74955_new_n181_));
INVX1 INVX1_333 ( .A(u2_u1__abc_74955_new_n185_), .Y(u2_u1__abc_74955_new_n186_));
INVX1 INVX1_334 ( .A(u2_u1__abc_74955_new_n190_), .Y(u2_u1__abc_74955_new_n191_));
INVX1 INVX1_335 ( .A(u2_u1__abc_74955_new_n195_), .Y(u2_u1__abc_74955_new_n196_));
INVX1 INVX1_336 ( .A(u2_u1__abc_74955_new_n200_), .Y(u2_u1__abc_74955_new_n201_));
INVX1 INVX1_337 ( .A(bank_adr_0_), .Y(u2_u1__abc_74955_new_n203_));
INVX1 INVX1_338 ( .A(bank_adr_1_), .Y(u2_u1__abc_74955_new_n204_));
INVX1 INVX1_339 ( .A(u2_u1_b3_last_row_9_), .Y(u2_u1__abc_74955_new_n332_));
INVX1 INVX1_34 ( .A(1'h0), .Y(u0__abc_76628_new_n5685_));
INVX1 INVX1_340 ( .A(u2_u1_b3_last_row_8_), .Y(u2_u1__abc_74955_new_n334_));
INVX1 INVX1_341 ( .A(u2_u1_b3_last_row_11_), .Y(u2_u1__abc_74955_new_n339_));
INVX1 INVX1_342 ( .A(u2_u1_b3_last_row_4_), .Y(u2_u1__abc_74955_new_n342_));
INVX1 INVX1_343 ( .A(u2_u1_b3_last_row_0_), .Y(u2_u1__abc_74955_new_n348_));
INVX1 INVX1_344 ( .A(u2_u1_b3_last_row_7_), .Y(u2_u1__abc_74955_new_n355_));
INVX1 INVX1_345 ( .A(u2_u1_b3_last_row_5_), .Y(u2_u1__abc_74955_new_n359_));
INVX1 INVX1_346 ( .A(u2_u1_b3_last_row_12_), .Y(u2_u1__abc_74955_new_n367_));
INVX1 INVX1_347 ( .A(u2_u1_b3_last_row_10_), .Y(u2_u1__abc_74955_new_n371_));
INVX1 INVX1_348 ( .A(u2_u1_b3_last_row_3_), .Y(u2_u1__abc_74955_new_n375_));
INVX1 INVX1_349 ( .A(u2_u1_b3_last_row_1_), .Y(u2_u1__abc_74955_new_n379_));
INVX1 INVX1_35 ( .A(1'h0), .Y(u0__abc_76628_new_n5687_));
INVX1 INVX1_350 ( .A(u2_u1_b3_last_row_6_), .Y(u2_u1__abc_74955_new_n385_));
INVX1 INVX1_351 ( .A(u2_u1_b3_last_row_2_), .Y(u2_u1__abc_74955_new_n388_));
INVX1 INVX1_352 ( .A(u2_u1_b1_last_row_0_), .Y(u2_u1__abc_74955_new_n399_));
INVX1 INVX1_353 ( .A(u2_u1_b1_last_row_4_), .Y(u2_u1__abc_74955_new_n403_));
INVX1 INVX1_354 ( .A(u2_u1_b1_last_row_3_), .Y(u2_u1__abc_74955_new_n407_));
INVX1 INVX1_355 ( .A(u2_u1_b1_last_row_8_), .Y(u2_u1__abc_74955_new_n413_));
INVX1 INVX1_356 ( .A(u2_u1_b1_last_row_6_), .Y(u2_u1__abc_74955_new_n417_));
INVX1 INVX1_357 ( .A(u2_u1_b1_last_row_12_), .Y(u2_u1__abc_74955_new_n422_));
INVX1 INVX1_358 ( .A(u2_u1_b1_last_row_11_), .Y(u2_u1__abc_74955_new_n425_));
INVX1 INVX1_359 ( .A(u2_u1_b1_last_row_2_), .Y(u2_u1__abc_74955_new_n431_));
INVX1 INVX1_36 ( .A(1'h0), .Y(u0__abc_76628_new_n5690_));
INVX1 INVX1_360 ( .A(u2_u1_b1_last_row_1_), .Y(u2_u1__abc_74955_new_n435_));
INVX1 INVX1_361 ( .A(u2_u1_b1_last_row_10_), .Y(u2_u1__abc_74955_new_n440_));
INVX1 INVX1_362 ( .A(u2_u1_b1_last_row_9_), .Y(u2_u1__abc_74955_new_n444_));
INVX1 INVX1_363 ( .A(u2_u1_b1_last_row_7_), .Y(u2_u1__abc_74955_new_n450_));
INVX1 INVX1_364 ( .A(u2_u1_b1_last_row_5_), .Y(u2_u1__abc_74955_new_n454_));
INVX1 INVX1_365 ( .A(u2_u1_b0_last_row_9_), .Y(u2_u1__abc_74955_new_n462_));
INVX1 INVX1_366 ( .A(u2_u1_b0_last_row_12_), .Y(u2_u1__abc_74955_new_n469_));
INVX1 INVX1_367 ( .A(u2_u1_b0_last_row_3_), .Y(u2_u1__abc_74955_new_n472_));
INVX1 INVX1_368 ( .A(u2_u1_b0_last_row_2_), .Y(u2_u1__abc_74955_new_n477_));
INVX1 INVX1_369 ( .A(u2_u1_b0_last_row_6_), .Y(u2_u1__abc_74955_new_n479_));
INVX1 INVX1_37 ( .A(1'h0), .Y(u0__abc_76628_new_n5691_));
INVX1 INVX1_370 ( .A(u2_u1_b0_last_row_0_), .Y(u2_u1__abc_74955_new_n488_));
INVX1 INVX1_371 ( .A(u2_u1_b0_last_row_1_), .Y(u2_u1__abc_74955_new_n492_));
INVX1 INVX1_372 ( .A(u2_u1_b0_last_row_5_), .Y(u2_u1__abc_74955_new_n498_));
INVX1 INVX1_373 ( .A(u2_u1_b0_last_row_8_), .Y(u2_u1__abc_74955_new_n501_));
INVX1 INVX1_374 ( .A(u2_u1_b0_last_row_4_), .Y(u2_u1__abc_74955_new_n506_));
INVX1 INVX1_375 ( .A(u2_u1_b0_last_row_11_), .Y(u2_u1__abc_74955_new_n508_));
INVX1 INVX1_376 ( .A(u2_u1_b0_last_row_7_), .Y(u2_u1__abc_74955_new_n516_));
INVX1 INVX1_377 ( .A(u2_u1_b0_last_row_10_), .Y(u2_u1__abc_74955_new_n520_));
INVX1 INVX1_378 ( .A(u2_u1_b2_last_row_8_), .Y(u2_u1__abc_74955_new_n527_));
INVX1 INVX1_379 ( .A(u2_u1_b2_last_row_9_), .Y(u2_u1__abc_74955_new_n533_));
INVX1 INVX1_38 ( .A(1'h0), .Y(u0__abc_76628_new_n5693_));
INVX1 INVX1_380 ( .A(u2_u1_b2_last_row_11_), .Y(u2_u1__abc_74955_new_n537_));
INVX1 INVX1_381 ( .A(u2_u1_b2_last_row_7_), .Y(u2_u1__abc_74955_new_n544_));
INVX1 INVX1_382 ( .A(u2_u1_b2_last_row_6_), .Y(u2_u1__abc_74955_new_n548_));
INVX1 INVX1_383 ( .A(u2_u1_b2_last_row_3_), .Y(u2_u1__abc_74955_new_n553_));
INVX1 INVX1_384 ( .A(u2_u1_b2_last_row_2_), .Y(u2_u1__abc_74955_new_n557_));
INVX1 INVX1_385 ( .A(u2_u1_b2_last_row_12_), .Y(u2_u1__abc_74955_new_n563_));
INVX1 INVX1_386 ( .A(u2_u1_b2_last_row_10_), .Y(u2_u1__abc_74955_new_n567_));
INVX1 INVX1_387 ( .A(u2_u1_b2_last_row_4_), .Y(u2_u1__abc_74955_new_n573_));
INVX1 INVX1_388 ( .A(u2_u1_b2_last_row_5_), .Y(u2_u1__abc_74955_new_n577_));
INVX1 INVX1_389 ( .A(u2_u1_b2_last_row_0_), .Y(u2_u1__abc_74955_new_n582_));
INVX1 INVX1_39 ( .A(1'h0), .Y(u0__abc_76628_new_n5696_));
INVX1 INVX1_390 ( .A(u2_u1_b2_last_row_1_), .Y(u2_u1__abc_74955_new_n585_));
INVX1 INVX1_391 ( .A(u2_bank_clr_1), .Y(u2_u1__abc_74955_new_n601_));
INVX1 INVX1_392 ( .A(u2_u1__abc_74955_new_n289_), .Y(u2_u1__abc_74955_new_n602_));
INVX1 INVX1_393 ( .A(u2_bank_clr_all_1), .Y(u2_u1__abc_74955_new_n604_));
INVX1 INVX1_394 ( .A(u2_u1__abc_74955_new_n608_), .Y(u2_u1__abc_74955_new_n609_));
INVX1 INVX1_395 ( .A(u2_u1__abc_74955_new_n247_), .Y(u2_u1__abc_74955_new_n616_));
INVX1 INVX1_396 ( .A(u2_u1__abc_74955_new_n205_), .Y(u2_u1__abc_74955_new_n621_));
INVX1 INVX1_397 ( .A(u3__abc_74070_new_n281_), .Y(u3__abc_74070_new_n282_));
INVX1 INVX1_398 ( .A(u3__abc_74070_new_n283_), .Y(u3__abc_74070_new_n284_));
INVX1 INVX1_399 ( .A(\wb_data_i[1] ), .Y(u3__abc_74070_new_n285_));
INVX1 INVX1_4 ( .A(u0__abc_76628_new_n1105_), .Y(u0__abc_76628_new_n1106_));
INVX1 INVX1_40 ( .A(1'h0), .Y(u0__abc_76628_new_n5697_));
INVX1 INVX1_400 ( .A(\wb_data_i[0] ), .Y(u3__abc_74070_new_n287_));
INVX1 INVX1_401 ( .A(u3__abc_74070_new_n290_), .Y(u3__abc_74070_new_n291_));
INVX1 INVX1_402 ( .A(u3__abc_74070_new_n293_), .Y(u3__abc_74070_new_n294_));
INVX1 INVX1_403 ( .A(u3__abc_74070_new_n296_), .Y(u3__abc_74070_new_n297_));
INVX1 INVX1_404 ( .A(u3__abc_74070_new_n298_), .Y(u3__abc_74070_new_n299_));
INVX1 INVX1_405 ( .A(\wb_data_i[5] ), .Y(u3__abc_74070_new_n300_));
INVX1 INVX1_406 ( .A(\wb_data_i[4] ), .Y(u3__abc_74070_new_n302_));
INVX1 INVX1_407 ( .A(u3__abc_74070_new_n304_), .Y(u3__abc_74070_new_n305_));
INVX1 INVX1_408 ( .A(u3__abc_74070_new_n308_), .Y(u3__abc_74070_new_n309_));
INVX1 INVX1_409 ( .A(u3__abc_74070_new_n317_), .Y(u3__abc_74070_new_n318_));
INVX1 INVX1_41 ( .A(1'h0), .Y(u0__abc_76628_new_n5699_));
INVX1 INVX1_410 ( .A(\wb_data_i[9] ), .Y(u3__abc_74070_new_n320_));
INVX1 INVX1_411 ( .A(\wb_data_i[8] ), .Y(u3__abc_74070_new_n322_));
INVX1 INVX1_412 ( .A(u3__abc_74070_new_n324_), .Y(u3__abc_74070_new_n325_));
INVX1 INVX1_413 ( .A(u3__abc_74070_new_n326_), .Y(u3__abc_74070_new_n327_));
INVX1 INVX1_414 ( .A(u3__abc_74070_new_n329_), .Y(u3__abc_74070_new_n330_));
INVX1 INVX1_415 ( .A(u3__abc_74070_new_n332_), .Y(u3__abc_74070_new_n333_));
INVX1 INVX1_416 ( .A(u3__abc_74070_new_n334_), .Y(u3__abc_74070_new_n335_));
INVX1 INVX1_417 ( .A(\wb_data_i[13] ), .Y(u3__abc_74070_new_n336_));
INVX1 INVX1_418 ( .A(\wb_data_i[12] ), .Y(u3__abc_74070_new_n338_));
INVX1 INVX1_419 ( .A(u3__abc_74070_new_n340_), .Y(u3__abc_74070_new_n341_));
INVX1 INVX1_42 ( .A(1'h0), .Y(u0__abc_76628_new_n5702_));
INVX1 INVX1_420 ( .A(u3__abc_74070_new_n344_), .Y(u3__abc_74070_new_n345_));
INVX1 INVX1_421 ( .A(u3__abc_74070_new_n352_), .Y(u3__abc_74070_new_n353_));
INVX1 INVX1_422 ( .A(\wb_data_i[17] ), .Y(u3__abc_74070_new_n355_));
INVX1 INVX1_423 ( .A(\wb_data_i[16] ), .Y(u3__abc_74070_new_n357_));
INVX1 INVX1_424 ( .A(u3__abc_74070_new_n359_), .Y(u3__abc_74070_new_n360_));
INVX1 INVX1_425 ( .A(u3__abc_74070_new_n361_), .Y(u3__abc_74070_new_n362_));
INVX1 INVX1_426 ( .A(u3__abc_74070_new_n366_), .Y(u3__abc_74070_new_n367_));
INVX1 INVX1_427 ( .A(u3__abc_74070_new_n368_), .Y(u3__abc_74070_new_n369_));
INVX1 INVX1_428 ( .A(\wb_data_i[21] ), .Y(u3__abc_74070_new_n370_));
INVX1 INVX1_429 ( .A(\wb_data_i[20] ), .Y(u3__abc_74070_new_n372_));
INVX1 INVX1_43 ( .A(1'h0), .Y(u0__abc_76628_new_n5703_));
INVX1 INVX1_430 ( .A(u3__abc_74070_new_n374_), .Y(u3__abc_74070_new_n375_));
INVX1 INVX1_431 ( .A(u3__abc_74070_new_n378_), .Y(u3__abc_74070_new_n379_));
INVX1 INVX1_432 ( .A(u3__abc_74070_new_n364_), .Y(u3__abc_74070_new_n381_));
INVX1 INVX1_433 ( .A(u3__abc_74070_new_n388_), .Y(u3__abc_74070_new_n389_));
INVX1 INVX1_434 ( .A(\wb_data_i[25] ), .Y(u3__abc_74070_new_n391_));
INVX1 INVX1_435 ( .A(\wb_data_i[24] ), .Y(u3__abc_74070_new_n393_));
INVX1 INVX1_436 ( .A(u3__abc_74070_new_n395_), .Y(u3__abc_74070_new_n396_));
INVX1 INVX1_437 ( .A(u3__abc_74070_new_n397_), .Y(u3__abc_74070_new_n398_));
INVX1 INVX1_438 ( .A(u3__abc_74070_new_n402_), .Y(u3__abc_74070_new_n403_));
INVX1 INVX1_439 ( .A(u3__abc_74070_new_n404_), .Y(u3__abc_74070_new_n405_));
INVX1 INVX1_44 ( .A(1'h0), .Y(u0__abc_76628_new_n5705_));
INVX1 INVX1_440 ( .A(\wb_data_i[29] ), .Y(u3__abc_74070_new_n406_));
INVX1 INVX1_441 ( .A(\wb_data_i[28] ), .Y(u3__abc_74070_new_n408_));
INVX1 INVX1_442 ( .A(u3__abc_74070_new_n410_), .Y(u3__abc_74070_new_n411_));
INVX1 INVX1_443 ( .A(u3__abc_74070_new_n414_), .Y(u3__abc_74070_new_n415_));
INVX1 INVX1_444 ( .A(u3__abc_74070_new_n400_), .Y(u3__abc_74070_new_n417_));
INVX1 INVX1_445 ( .A(csc_4_), .Y(u3__abc_74070_new_n448_));
INVX1 INVX1_446 ( .A(wb_cyc_i), .Y(u3__abc_74070_new_n850_));
INVX1 INVX1_447 ( .A(u3__abc_74070_new_n855_), .Y(u3__abc_74070_new_n856_));
INVX1 INVX1_448 ( .A(u3_rd_fifo_out_16_), .Y(u3__abc_74070_new_n858_));
INVX1 INVX1_449 ( .A(u3_rd_fifo_out_17_), .Y(u3__abc_74070_new_n860_));
INVX1 INVX1_45 ( .A(lmr_ack), .Y(u0__abc_76628_new_n5708_));
INVX1 INVX1_450 ( .A(u3_rd_fifo_out_34_), .Y(u3__abc_74070_new_n864_));
INVX1 INVX1_451 ( .A(u3__abc_74070_new_n857_), .Y(u3__abc_74070_new_n871_));
INVX1 INVX1_452 ( .A(u3__abc_74070_new_n876_), .Y(u3__abc_74070_new_n877_));
INVX1 INVX1_453 ( .A(u3__abc_74070_new_n879_), .Y(u3__abc_74070_new_n880_));
INVX1 INVX1_454 ( .A(u3_rd_fifo_out_19_), .Y(u3__abc_74070_new_n882_));
INVX1 INVX1_455 ( .A(u3__abc_74070_new_n883_), .Y(u3__abc_74070_new_n884_));
INVX1 INVX1_456 ( .A(u3__abc_74070_new_n881_), .Y(u3__abc_74070_new_n888_));
INVX1 INVX1_457 ( .A(u3__abc_74070_new_n886_), .Y(u3__abc_74070_new_n889_));
INVX1 INVX1_458 ( .A(u3__abc_74070_new_n891_), .Y(u3__abc_74070_new_n892_));
INVX1 INVX1_459 ( .A(u3__abc_74070_new_n898_), .Y(u3__abc_74070_new_n899_));
INVX1 INVX1_46 ( .A(init_ack), .Y(u0__abc_76628_new_n5710_));
INVX1 INVX1_460 ( .A(u3_rd_fifo_out_24_), .Y(u3__abc_74070_new_n901_));
INVX1 INVX1_461 ( .A(u3_rd_fifo_out_25_), .Y(u3__abc_74070_new_n902_));
INVX1 INVX1_462 ( .A(u3_rd_fifo_out_35_), .Y(u3__abc_74070_new_n907_));
INVX1 INVX1_463 ( .A(u3__abc_74070_new_n904_), .Y(u3__abc_74070_new_n909_));
INVX1 INVX1_464 ( .A(u3__abc_74070_new_n900_), .Y(u3__abc_74070_new_n914_));
INVX1 INVX1_465 ( .A(u3__abc_74070_new_n919_), .Y(u3__abc_74070_new_n920_));
INVX1 INVX1_466 ( .A(u3__abc_74070_new_n922_), .Y(u3__abc_74070_new_n923_));
INVX1 INVX1_467 ( .A(u3_rd_fifo_out_27_), .Y(u3__abc_74070_new_n925_));
INVX1 INVX1_468 ( .A(u3__abc_74070_new_n926_), .Y(u3__abc_74070_new_n927_));
INVX1 INVX1_469 ( .A(u3__abc_74070_new_n924_), .Y(u3__abc_74070_new_n931_));
INVX1 INVX1_47 ( .A(lmr_req), .Y(u0__abc_76628_new_n5712_));
INVX1 INVX1_470 ( .A(u3__abc_74070_new_n929_), .Y(u3__abc_74070_new_n932_));
INVX1 INVX1_471 ( .A(u3__abc_74070_new_n934_), .Y(u3__abc_74070_new_n935_));
INVX1 INVX1_472 ( .A(u3__abc_74070_new_n942_), .Y(u3__abc_74070_new_n943_));
INVX1 INVX1_473 ( .A(u3__abc_74070_new_n944_), .Y(u3__abc_74070_new_n945_));
INVX1 INVX1_474 ( .A(u3_rd_fifo_out_33_), .Y(u3__abc_74070_new_n946_));
INVX1 INVX1_475 ( .A(u3__abc_74070_new_n948_), .Y(u3__abc_74070_new_n949_));
INVX1 INVX1_476 ( .A(u3_rd_fifo_out_8_), .Y(u3__abc_74070_new_n952_));
INVX1 INVX1_477 ( .A(u3_rd_fifo_out_9_), .Y(u3__abc_74070_new_n953_));
INVX1 INVX1_478 ( .A(u3__abc_74070_new_n963_), .Y(u3__abc_74070_new_n964_));
INVX1 INVX1_479 ( .A(u3__abc_74070_new_n966_), .Y(u3__abc_74070_new_n967_));
INVX1 INVX1_48 ( .A(u0_u0__abc_72207_new_n206_), .Y(u0_u0__abc_72207_new_n207_));
INVX1 INVX1_480 ( .A(u3__abc_74070_new_n968_), .Y(u3__abc_74070_new_n969_));
INVX1 INVX1_481 ( .A(u3_rd_fifo_out_11_), .Y(u3__abc_74070_new_n970_));
INVX1 INVX1_482 ( .A(u3__abc_74070_new_n971_), .Y(u3__abc_74070_new_n972_));
INVX1 INVX1_483 ( .A(u3__abc_74070_new_n974_), .Y(u3__abc_74070_new_n975_));
INVX1 INVX1_484 ( .A(u3__abc_74070_new_n978_), .Y(u3__abc_74070_new_n979_));
INVX1 INVX1_485 ( .A(u3__abc_74070_new_n985_), .Y(u3__abc_74070_new_n986_));
INVX1 INVX1_486 ( .A(u3__abc_74070_new_n987_), .Y(u3__abc_74070_new_n988_));
INVX1 INVX1_487 ( .A(u3_rd_fifo_out_32_), .Y(u3__abc_74070_new_n989_));
INVX1 INVX1_488 ( .A(u3__abc_74070_new_n991_), .Y(u3__abc_74070_new_n992_));
INVX1 INVX1_489 ( .A(u3_rd_fifo_out_0_), .Y(u3__abc_74070_new_n995_));
INVX1 INVX1_49 ( .A(u0_u0__abc_72207_new_n208_), .Y(u0_u0__abc_72207_new_n210_));
INVX1 INVX1_490 ( .A(u3_rd_fifo_out_1_), .Y(u3__abc_74070_new_n997_));
INVX1 INVX1_491 ( .A(u3__abc_74070_new_n1007_), .Y(u3__abc_74070_new_n1008_));
INVX1 INVX1_492 ( .A(u3__abc_74070_new_n1010_), .Y(u3__abc_74070_new_n1011_));
INVX1 INVX1_493 ( .A(u3__abc_74070_new_n1012_), .Y(u3__abc_74070_new_n1013_));
INVX1 INVX1_494 ( .A(u3_rd_fifo_out_3_), .Y(u3__abc_74070_new_n1014_));
INVX1 INVX1_495 ( .A(u3__abc_74070_new_n1015_), .Y(u3__abc_74070_new_n1016_));
INVX1 INVX1_496 ( .A(u3__abc_74070_new_n1018_), .Y(u3__abc_74070_new_n1019_));
INVX1 INVX1_497 ( .A(u3__abc_74070_new_n1022_), .Y(u3__abc_74070_new_n1023_));
INVX1 INVX1_498 ( .A(wb_we_i), .Y(u3__abc_74070_new_n1030_));
INVX1 INVX1_499 ( .A(mc_data_ir_0_), .Y(u3_u0__abc_75526_new_n384_));
INVX1 INVX1_5 ( .A(u0__abc_76628_new_n1113_), .Y(u0__abc_76628_new_n1120_));
INVX1 INVX1_50 ( .A(u0_lmr_ack0), .Y(u0_u0__abc_72207_new_n211_));
INVX1 INVX1_500 ( .A(u3_u0__abc_75526_new_n385_), .Y(u3_u0__abc_75526_new_n386_));
INVX1 INVX1_501 ( .A(mc_data_ir_1_), .Y(u3_u0__abc_75526_new_n389_));
INVX1 INVX1_502 ( .A(u3_u0__abc_75526_new_n390_), .Y(u3_u0__abc_75526_new_n391_));
INVX1 INVX1_503 ( .A(mc_data_ir_2_), .Y(u3_u0__abc_75526_new_n394_));
INVX1 INVX1_504 ( .A(u3_u0__abc_75526_new_n395_), .Y(u3_u0__abc_75526_new_n396_));
INVX1 INVX1_505 ( .A(mc_data_ir_3_), .Y(u3_u0__abc_75526_new_n399_));
INVX1 INVX1_506 ( .A(u3_u0__abc_75526_new_n400_), .Y(u3_u0__abc_75526_new_n401_));
INVX1 INVX1_507 ( .A(mc_data_ir_4_), .Y(u3_u0__abc_75526_new_n404_));
INVX1 INVX1_508 ( .A(u3_u0__abc_75526_new_n405_), .Y(u3_u0__abc_75526_new_n406_));
INVX1 INVX1_509 ( .A(mc_data_ir_5_), .Y(u3_u0__abc_75526_new_n409_));
INVX1 INVX1_51 ( .A(u0_u0_addr_r_5_), .Y(u0_u0__abc_72207_new_n215_));
INVX1 INVX1_510 ( .A(u3_u0__abc_75526_new_n410_), .Y(u3_u0__abc_75526_new_n411_));
INVX1 INVX1_511 ( .A(mc_data_ir_6_), .Y(u3_u0__abc_75526_new_n414_));
INVX1 INVX1_512 ( .A(u3_u0__abc_75526_new_n415_), .Y(u3_u0__abc_75526_new_n416_));
INVX1 INVX1_513 ( .A(mc_data_ir_7_), .Y(u3_u0__abc_75526_new_n419_));
INVX1 INVX1_514 ( .A(u3_u0__abc_75526_new_n420_), .Y(u3_u0__abc_75526_new_n421_));
INVX1 INVX1_515 ( .A(mc_data_ir_8_), .Y(u3_u0__abc_75526_new_n424_));
INVX1 INVX1_516 ( .A(u3_u0__abc_75526_new_n425_), .Y(u3_u0__abc_75526_new_n426_));
INVX1 INVX1_517 ( .A(mc_data_ir_9_), .Y(u3_u0__abc_75526_new_n429_));
INVX1 INVX1_518 ( .A(u3_u0__abc_75526_new_n430_), .Y(u3_u0__abc_75526_new_n431_));
INVX1 INVX1_519 ( .A(mc_data_ir_10_), .Y(u3_u0__abc_75526_new_n434_));
INVX1 INVX1_52 ( .A(u0_u0_addr_r_6_), .Y(u0_u0__abc_72207_new_n217_));
INVX1 INVX1_520 ( .A(u3_u0__abc_75526_new_n435_), .Y(u3_u0__abc_75526_new_n436_));
INVX1 INVX1_521 ( .A(mc_data_ir_11_), .Y(u3_u0__abc_75526_new_n439_));
INVX1 INVX1_522 ( .A(u3_u0__abc_75526_new_n440_), .Y(u3_u0__abc_75526_new_n441_));
INVX1 INVX1_523 ( .A(mc_data_ir_12_), .Y(u3_u0__abc_75526_new_n444_));
INVX1 INVX1_524 ( .A(u3_u0__abc_75526_new_n445_), .Y(u3_u0__abc_75526_new_n446_));
INVX1 INVX1_525 ( .A(mc_data_ir_13_), .Y(u3_u0__abc_75526_new_n449_));
INVX1 INVX1_526 ( .A(u3_u0__abc_75526_new_n450_), .Y(u3_u0__abc_75526_new_n451_));
INVX1 INVX1_527 ( .A(mc_data_ir_14_), .Y(u3_u0__abc_75526_new_n454_));
INVX1 INVX1_528 ( .A(u3_u0__abc_75526_new_n455_), .Y(u3_u0__abc_75526_new_n456_));
INVX1 INVX1_529 ( .A(mc_data_ir_15_), .Y(u3_u0__abc_75526_new_n459_));
INVX1 INVX1_53 ( .A(u0_u0_addr_r_3_), .Y(u0_u0__abc_72207_new_n218_));
INVX1 INVX1_530 ( .A(u3_u0__abc_75526_new_n460_), .Y(u3_u0__abc_75526_new_n461_));
INVX1 INVX1_531 ( .A(mc_data_ir_16_), .Y(u3_u0__abc_75526_new_n464_));
INVX1 INVX1_532 ( .A(u3_u0__abc_75526_new_n465_), .Y(u3_u0__abc_75526_new_n466_));
INVX1 INVX1_533 ( .A(mc_data_ir_17_), .Y(u3_u0__abc_75526_new_n469_));
INVX1 INVX1_534 ( .A(u3_u0__abc_75526_new_n470_), .Y(u3_u0__abc_75526_new_n471_));
INVX1 INVX1_535 ( .A(mc_data_ir_18_), .Y(u3_u0__abc_75526_new_n474_));
INVX1 INVX1_536 ( .A(u3_u0__abc_75526_new_n475_), .Y(u3_u0__abc_75526_new_n476_));
INVX1 INVX1_537 ( .A(mc_data_ir_19_), .Y(u3_u0__abc_75526_new_n479_));
INVX1 INVX1_538 ( .A(u3_u0__abc_75526_new_n480_), .Y(u3_u0__abc_75526_new_n481_));
INVX1 INVX1_539 ( .A(mc_data_ir_20_), .Y(u3_u0__abc_75526_new_n484_));
INVX1 INVX1_54 ( .A(u0_u0_addr_r_2_), .Y(u0_u0__abc_72207_new_n352_));
INVX1 INVX1_540 ( .A(u3_u0__abc_75526_new_n485_), .Y(u3_u0__abc_75526_new_n486_));
INVX1 INVX1_541 ( .A(mc_data_ir_21_), .Y(u3_u0__abc_75526_new_n489_));
INVX1 INVX1_542 ( .A(u3_u0__abc_75526_new_n490_), .Y(u3_u0__abc_75526_new_n491_));
INVX1 INVX1_543 ( .A(mc_data_ir_22_), .Y(u3_u0__abc_75526_new_n494_));
INVX1 INVX1_544 ( .A(u3_u0__abc_75526_new_n495_), .Y(u3_u0__abc_75526_new_n496_));
INVX1 INVX1_545 ( .A(mc_data_ir_23_), .Y(u3_u0__abc_75526_new_n499_));
INVX1 INVX1_546 ( .A(u3_u0__abc_75526_new_n500_), .Y(u3_u0__abc_75526_new_n501_));
INVX1 INVX1_547 ( .A(mc_data_ir_24_), .Y(u3_u0__abc_75526_new_n504_));
INVX1 INVX1_548 ( .A(u3_u0__abc_75526_new_n505_), .Y(u3_u0__abc_75526_new_n506_));
INVX1 INVX1_549 ( .A(mc_data_ir_25_), .Y(u3_u0__abc_75526_new_n509_));
INVX1 INVX1_55 ( .A(u0_u0__abc_72207_new_n219_), .Y(u0_u0__abc_72207_new_n356_));
INVX1 INVX1_550 ( .A(u3_u0__abc_75526_new_n510_), .Y(u3_u0__abc_75526_new_n511_));
INVX1 INVX1_551 ( .A(mc_data_ir_26_), .Y(u3_u0__abc_75526_new_n514_));
INVX1 INVX1_552 ( .A(u3_u0__abc_75526_new_n515_), .Y(u3_u0__abc_75526_new_n516_));
INVX1 INVX1_553 ( .A(mc_data_ir_27_), .Y(u3_u0__abc_75526_new_n519_));
INVX1 INVX1_554 ( .A(u3_u0__abc_75526_new_n520_), .Y(u3_u0__abc_75526_new_n521_));
INVX1 INVX1_555 ( .A(mc_data_ir_28_), .Y(u3_u0__abc_75526_new_n524_));
INVX1 INVX1_556 ( .A(u3_u0__abc_75526_new_n525_), .Y(u3_u0__abc_75526_new_n526_));
INVX1 INVX1_557 ( .A(mc_data_ir_29_), .Y(u3_u0__abc_75526_new_n529_));
INVX1 INVX1_558 ( .A(u3_u0__abc_75526_new_n530_), .Y(u3_u0__abc_75526_new_n531_));
INVX1 INVX1_559 ( .A(mc_data_ir_30_), .Y(u3_u0__abc_75526_new_n534_));
INVX1 INVX1_56 ( .A(u0_rf_we), .Y(u0_u0__abc_72207_new_n357_));
INVX1 INVX1_560 ( .A(u3_u0__abc_75526_new_n535_), .Y(u3_u0__abc_75526_new_n536_));
INVX1 INVX1_561 ( .A(mc_data_ir_31_), .Y(u3_u0__abc_75526_new_n539_));
INVX1 INVX1_562 ( .A(u3_u0__abc_75526_new_n540_), .Y(u3_u0__abc_75526_new_n541_));
INVX1 INVX1_563 ( .A(mc_data_ir_32_), .Y(u3_u0__abc_75526_new_n544_));
INVX1 INVX1_564 ( .A(u3_u0__abc_75526_new_n545_), .Y(u3_u0__abc_75526_new_n546_));
INVX1 INVX1_565 ( .A(mc_data_ir_33_), .Y(u3_u0__abc_75526_new_n549_));
INVX1 INVX1_566 ( .A(u3_u0__abc_75526_new_n550_), .Y(u3_u0__abc_75526_new_n551_));
INVX1 INVX1_567 ( .A(mc_data_ir_34_), .Y(u3_u0__abc_75526_new_n554_));
INVX1 INVX1_568 ( .A(u3_u0__abc_75526_new_n555_), .Y(u3_u0__abc_75526_new_n556_));
INVX1 INVX1_569 ( .A(mc_data_ir_35_), .Y(u3_u0__abc_75526_new_n559_));
INVX1 INVX1_57 ( .A(u0_csc0_23_), .Y(u0_u0__abc_72207_new_n500_));
INVX1 INVX1_570 ( .A(u3_u0__abc_75526_new_n560_), .Y(u3_u0__abc_75526_new_n561_));
INVX1 INVX1_571 ( .A(u3_u0__abc_75526_new_n565_), .Y(u3_u0__abc_75526_new_n566_));
INVX1 INVX1_572 ( .A(u3_u0__abc_75526_new_n569_), .Y(u3_u0__abc_75526_new_n570_));
INVX1 INVX1_573 ( .A(u3_u0__abc_75526_new_n573_), .Y(u3_u0__abc_75526_new_n574_));
INVX1 INVX1_574 ( .A(u3_u0__abc_75526_new_n577_), .Y(u3_u0__abc_75526_new_n578_));
INVX1 INVX1_575 ( .A(u3_u0__abc_75526_new_n581_), .Y(u3_u0__abc_75526_new_n582_));
INVX1 INVX1_576 ( .A(u3_u0__abc_75526_new_n585_), .Y(u3_u0__abc_75526_new_n586_));
INVX1 INVX1_577 ( .A(u3_u0__abc_75526_new_n589_), .Y(u3_u0__abc_75526_new_n590_));
INVX1 INVX1_578 ( .A(u3_u0__abc_75526_new_n593_), .Y(u3_u0__abc_75526_new_n594_));
INVX1 INVX1_579 ( .A(u3_u0__abc_75526_new_n597_), .Y(u3_u0__abc_75526_new_n598_));
INVX1 INVX1_58 ( .A(\wb_addr_i[28] ), .Y(u0_u0__abc_72207_new_n501_));
INVX1 INVX1_580 ( .A(u3_u0__abc_75526_new_n601_), .Y(u3_u0__abc_75526_new_n602_));
INVX1 INVX1_581 ( .A(u3_u0__abc_75526_new_n605_), .Y(u3_u0__abc_75526_new_n606_));
INVX1 INVX1_582 ( .A(u3_u0__abc_75526_new_n609_), .Y(u3_u0__abc_75526_new_n610_));
INVX1 INVX1_583 ( .A(u3_u0__abc_75526_new_n613_), .Y(u3_u0__abc_75526_new_n614_));
INVX1 INVX1_584 ( .A(u3_u0__abc_75526_new_n617_), .Y(u3_u0__abc_75526_new_n618_));
INVX1 INVX1_585 ( .A(u3_u0__abc_75526_new_n621_), .Y(u3_u0__abc_75526_new_n622_));
INVX1 INVX1_586 ( .A(u3_u0__abc_75526_new_n625_), .Y(u3_u0__abc_75526_new_n626_));
INVX1 INVX1_587 ( .A(u3_u0__abc_75526_new_n629_), .Y(u3_u0__abc_75526_new_n630_));
INVX1 INVX1_588 ( .A(u3_u0__abc_75526_new_n633_), .Y(u3_u0__abc_75526_new_n634_));
INVX1 INVX1_589 ( .A(u3_u0__abc_75526_new_n637_), .Y(u3_u0__abc_75526_new_n638_));
INVX1 INVX1_59 ( .A(u0_csc_mask_7_), .Y(u0_u0__abc_72207_new_n503_));
INVX1 INVX1_590 ( .A(u3_u0__abc_75526_new_n641_), .Y(u3_u0__abc_75526_new_n642_));
INVX1 INVX1_591 ( .A(u3_u0__abc_75526_new_n645_), .Y(u3_u0__abc_75526_new_n646_));
INVX1 INVX1_592 ( .A(u3_u0__abc_75526_new_n649_), .Y(u3_u0__abc_75526_new_n650_));
INVX1 INVX1_593 ( .A(u3_u0__abc_75526_new_n653_), .Y(u3_u0__abc_75526_new_n654_));
INVX1 INVX1_594 ( .A(u3_u0__abc_75526_new_n657_), .Y(u3_u0__abc_75526_new_n658_));
INVX1 INVX1_595 ( .A(u3_u0__abc_75526_new_n661_), .Y(u3_u0__abc_75526_new_n662_));
INVX1 INVX1_596 ( .A(u3_u0__abc_75526_new_n665_), .Y(u3_u0__abc_75526_new_n666_));
INVX1 INVX1_597 ( .A(u3_u0__abc_75526_new_n669_), .Y(u3_u0__abc_75526_new_n670_));
INVX1 INVX1_598 ( .A(u3_u0__abc_75526_new_n673_), .Y(u3_u0__abc_75526_new_n674_));
INVX1 INVX1_599 ( .A(u3_u0__abc_75526_new_n677_), .Y(u3_u0__abc_75526_new_n678_));
INVX1 INVX1_6 ( .A(u0__abc_76628_new_n1119_), .Y(u0__abc_76628_new_n1125_));
INVX1 INVX1_60 ( .A(u0_csc_mask_6_), .Y(u0_u0__abc_72207_new_n508_));
INVX1 INVX1_600 ( .A(u3_u0__abc_75526_new_n681_), .Y(u3_u0__abc_75526_new_n682_));
INVX1 INVX1_601 ( .A(u3_u0__abc_75526_new_n685_), .Y(u3_u0__abc_75526_new_n686_));
INVX1 INVX1_602 ( .A(u3_u0__abc_75526_new_n689_), .Y(u3_u0__abc_75526_new_n690_));
INVX1 INVX1_603 ( .A(u3_u0__abc_75526_new_n693_), .Y(u3_u0__abc_75526_new_n694_));
INVX1 INVX1_604 ( .A(u3_u0__abc_75526_new_n697_), .Y(u3_u0__abc_75526_new_n698_));
INVX1 INVX1_605 ( .A(u3_u0__abc_75526_new_n701_), .Y(u3_u0__abc_75526_new_n702_));
INVX1 INVX1_606 ( .A(u3_u0__abc_75526_new_n705_), .Y(u3_u0__abc_75526_new_n706_));
INVX1 INVX1_607 ( .A(u3_u0__abc_75526_new_n710_), .Y(u3_u0__abc_75526_new_n711_));
INVX1 INVX1_608 ( .A(u3_u0__abc_75526_new_n714_), .Y(u3_u0__abc_75526_new_n715_));
INVX1 INVX1_609 ( .A(u3_u0__abc_75526_new_n718_), .Y(u3_u0__abc_75526_new_n719_));
INVX1 INVX1_61 ( .A(u0_csc0_22_), .Y(u0_u0__abc_72207_new_n509_));
INVX1 INVX1_610 ( .A(u3_u0__abc_75526_new_n722_), .Y(u3_u0__abc_75526_new_n723_));
INVX1 INVX1_611 ( .A(u3_u0__abc_75526_new_n726_), .Y(u3_u0__abc_75526_new_n727_));
INVX1 INVX1_612 ( .A(u3_u0__abc_75526_new_n730_), .Y(u3_u0__abc_75526_new_n731_));
INVX1 INVX1_613 ( .A(u3_u0__abc_75526_new_n734_), .Y(u3_u0__abc_75526_new_n735_));
INVX1 INVX1_614 ( .A(u3_u0__abc_75526_new_n738_), .Y(u3_u0__abc_75526_new_n739_));
INVX1 INVX1_615 ( .A(u3_u0__abc_75526_new_n742_), .Y(u3_u0__abc_75526_new_n743_));
INVX1 INVX1_616 ( .A(u3_u0__abc_75526_new_n746_), .Y(u3_u0__abc_75526_new_n747_));
INVX1 INVX1_617 ( .A(u3_u0__abc_75526_new_n750_), .Y(u3_u0__abc_75526_new_n751_));
INVX1 INVX1_618 ( .A(u3_u0__abc_75526_new_n754_), .Y(u3_u0__abc_75526_new_n755_));
INVX1 INVX1_619 ( .A(u3_u0__abc_75526_new_n758_), .Y(u3_u0__abc_75526_new_n759_));
INVX1 INVX1_62 ( .A(\wb_addr_i[27] ), .Y(u0_u0__abc_72207_new_n510_));
INVX1 INVX1_620 ( .A(u3_u0__abc_75526_new_n762_), .Y(u3_u0__abc_75526_new_n763_));
INVX1 INVX1_621 ( .A(u3_u0__abc_75526_new_n766_), .Y(u3_u0__abc_75526_new_n767_));
INVX1 INVX1_622 ( .A(u3_u0__abc_75526_new_n770_), .Y(u3_u0__abc_75526_new_n771_));
INVX1 INVX1_623 ( .A(u3_u0__abc_75526_new_n774_), .Y(u3_u0__abc_75526_new_n775_));
INVX1 INVX1_624 ( .A(u3_u0__abc_75526_new_n778_), .Y(u3_u0__abc_75526_new_n779_));
INVX1 INVX1_625 ( .A(u3_u0__abc_75526_new_n782_), .Y(u3_u0__abc_75526_new_n783_));
INVX1 INVX1_626 ( .A(u3_u0__abc_75526_new_n786_), .Y(u3_u0__abc_75526_new_n787_));
INVX1 INVX1_627 ( .A(u3_u0__abc_75526_new_n790_), .Y(u3_u0__abc_75526_new_n791_));
INVX1 INVX1_628 ( .A(u3_u0__abc_75526_new_n794_), .Y(u3_u0__abc_75526_new_n795_));
INVX1 INVX1_629 ( .A(u3_u0__abc_75526_new_n798_), .Y(u3_u0__abc_75526_new_n799_));
INVX1 INVX1_63 ( .A(u0_csc_mask_5_), .Y(u0_u0__abc_72207_new_n516_));
INVX1 INVX1_630 ( .A(u3_u0__abc_75526_new_n802_), .Y(u3_u0__abc_75526_new_n803_));
INVX1 INVX1_631 ( .A(u3_u0__abc_75526_new_n806_), .Y(u3_u0__abc_75526_new_n807_));
INVX1 INVX1_632 ( .A(u3_u0__abc_75526_new_n810_), .Y(u3_u0__abc_75526_new_n811_));
INVX1 INVX1_633 ( .A(u3_u0__abc_75526_new_n814_), .Y(u3_u0__abc_75526_new_n815_));
INVX1 INVX1_634 ( .A(u3_u0__abc_75526_new_n818_), .Y(u3_u0__abc_75526_new_n819_));
INVX1 INVX1_635 ( .A(u3_u0__abc_75526_new_n822_), .Y(u3_u0__abc_75526_new_n823_));
INVX1 INVX1_636 ( .A(u3_u0__abc_75526_new_n826_), .Y(u3_u0__abc_75526_new_n827_));
INVX1 INVX1_637 ( .A(u3_u0__abc_75526_new_n830_), .Y(u3_u0__abc_75526_new_n831_));
INVX1 INVX1_638 ( .A(u3_u0__abc_75526_new_n834_), .Y(u3_u0__abc_75526_new_n835_));
INVX1 INVX1_639 ( .A(u3_u0__abc_75526_new_n838_), .Y(u3_u0__abc_75526_new_n839_));
INVX1 INVX1_64 ( .A(u0_csc0_21_), .Y(u0_u0__abc_72207_new_n517_));
INVX1 INVX1_640 ( .A(u3_u0__abc_75526_new_n842_), .Y(u3_u0__abc_75526_new_n843_));
INVX1 INVX1_641 ( .A(u3_u0__abc_75526_new_n846_), .Y(u3_u0__abc_75526_new_n847_));
INVX1 INVX1_642 ( .A(u3_u0__abc_75526_new_n850_), .Y(u3_u0__abc_75526_new_n851_));
INVX1 INVX1_643 ( .A(u3_re), .Y(u3_u0__abc_75526_new_n853_));
INVX1 INVX1_644 ( .A(dv), .Y(u3_u0__abc_75526_new_n871_));
INVX1 INVX1_645 ( .A(u3_u0__abc_75526_new_n886_), .Y(u3_u0__abc_75526_new_n887_));
INVX1 INVX1_646 ( .A(u3_u0__abc_75526_new_n890_), .Y(u3_u0__abc_75526_new_n891_));
INVX1 INVX1_647 ( .A(u3_u0__abc_75526_new_n894_), .Y(u3_u0__abc_75526_new_n895_));
INVX1 INVX1_648 ( .A(u3_u0__abc_75526_new_n898_), .Y(u3_u0__abc_75526_new_n899_));
INVX1 INVX1_649 ( .A(u3_u0__abc_75526_new_n902_), .Y(u3_u0__abc_75526_new_n903_));
INVX1 INVX1_65 ( .A(\wb_addr_i[26] ), .Y(u0_u0__abc_72207_new_n518_));
INVX1 INVX1_650 ( .A(u3_u0__abc_75526_new_n906_), .Y(u3_u0__abc_75526_new_n907_));
INVX1 INVX1_651 ( .A(u3_u0__abc_75526_new_n910_), .Y(u3_u0__abc_75526_new_n911_));
INVX1 INVX1_652 ( .A(u3_u0__abc_75526_new_n914_), .Y(u3_u0__abc_75526_new_n915_));
INVX1 INVX1_653 ( .A(u3_u0__abc_75526_new_n918_), .Y(u3_u0__abc_75526_new_n919_));
INVX1 INVX1_654 ( .A(u3_u0__abc_75526_new_n922_), .Y(u3_u0__abc_75526_new_n923_));
INVX1 INVX1_655 ( .A(u3_u0__abc_75526_new_n926_), .Y(u3_u0__abc_75526_new_n927_));
INVX1 INVX1_656 ( .A(u3_u0__abc_75526_new_n930_), .Y(u3_u0__abc_75526_new_n931_));
INVX1 INVX1_657 ( .A(u3_u0__abc_75526_new_n934_), .Y(u3_u0__abc_75526_new_n935_));
INVX1 INVX1_658 ( .A(u3_u0__abc_75526_new_n938_), .Y(u3_u0__abc_75526_new_n939_));
INVX1 INVX1_659 ( .A(u3_u0__abc_75526_new_n942_), .Y(u3_u0__abc_75526_new_n943_));
INVX1 INVX1_66 ( .A(u0_csc_mask_0_), .Y(u0_u0__abc_72207_new_n524_));
INVX1 INVX1_660 ( .A(u3_u0__abc_75526_new_n946_), .Y(u3_u0__abc_75526_new_n947_));
INVX1 INVX1_661 ( .A(u3_u0__abc_75526_new_n950_), .Y(u3_u0__abc_75526_new_n951_));
INVX1 INVX1_662 ( .A(u3_u0__abc_75526_new_n954_), .Y(u3_u0__abc_75526_new_n955_));
INVX1 INVX1_663 ( .A(u3_u0__abc_75526_new_n958_), .Y(u3_u0__abc_75526_new_n959_));
INVX1 INVX1_664 ( .A(u3_u0__abc_75526_new_n962_), .Y(u3_u0__abc_75526_new_n963_));
INVX1 INVX1_665 ( .A(u3_u0__abc_75526_new_n966_), .Y(u3_u0__abc_75526_new_n967_));
INVX1 INVX1_666 ( .A(u3_u0__abc_75526_new_n970_), .Y(u3_u0__abc_75526_new_n971_));
INVX1 INVX1_667 ( .A(u3_u0__abc_75526_new_n974_), .Y(u3_u0__abc_75526_new_n975_));
INVX1 INVX1_668 ( .A(u3_u0__abc_75526_new_n978_), .Y(u3_u0__abc_75526_new_n979_));
INVX1 INVX1_669 ( .A(u3_u0__abc_75526_new_n982_), .Y(u3_u0__abc_75526_new_n983_));
INVX1 INVX1_67 ( .A(u0_csc0_16_), .Y(u0_u0__abc_72207_new_n525_));
INVX1 INVX1_670 ( .A(u3_u0__abc_75526_new_n986_), .Y(u3_u0__abc_75526_new_n987_));
INVX1 INVX1_671 ( .A(u3_u0__abc_75526_new_n990_), .Y(u3_u0__abc_75526_new_n991_));
INVX1 INVX1_672 ( .A(u3_u0__abc_75526_new_n994_), .Y(u3_u0__abc_75526_new_n995_));
INVX1 INVX1_673 ( .A(u3_u0__abc_75526_new_n998_), .Y(u3_u0__abc_75526_new_n999_));
INVX1 INVX1_674 ( .A(u3_u0__abc_75526_new_n1002_), .Y(u3_u0__abc_75526_new_n1003_));
INVX1 INVX1_675 ( .A(u3_u0__abc_75526_new_n1006_), .Y(u3_u0__abc_75526_new_n1007_));
INVX1 INVX1_676 ( .A(u3_u0__abc_75526_new_n1010_), .Y(u3_u0__abc_75526_new_n1011_));
INVX1 INVX1_677 ( .A(u3_u0__abc_75526_new_n1014_), .Y(u3_u0__abc_75526_new_n1015_));
INVX1 INVX1_678 ( .A(u3_u0__abc_75526_new_n1018_), .Y(u3_u0__abc_75526_new_n1019_));
INVX1 INVX1_679 ( .A(u3_u0__abc_75526_new_n1022_), .Y(u3_u0__abc_75526_new_n1023_));
INVX1 INVX1_68 ( .A(\wb_addr_i[21] ), .Y(u0_u0__abc_72207_new_n526_));
INVX1 INVX1_680 ( .A(u3_u0__abc_75526_new_n1026_), .Y(u3_u0__abc_75526_new_n1027_));
INVX1 INVX1_681 ( .A(u3_u0_rd_adr_0_), .Y(u3_u0__abc_75526_new_n1029_));
INVX1 INVX1_682 ( .A(u3_u0_rd_adr_1_), .Y(u3_u0__abc_75526_new_n1030_));
INVX1 INVX1_683 ( .A(u3_u0_rd_adr_2_), .Y(u3_u0__abc_75526_new_n1032_));
INVX1 INVX1_684 ( .A(u3_u0__abc_75526_new_n1034__bF_buf5), .Y(u3_u0__abc_75526_new_n1035_));
INVX1 INVX1_685 ( .A(u3_u0_rd_adr_3_), .Y(u3_u0__abc_75526_new_n1046_));
INVX1 INVX1_686 ( .A(u4__abc_76448_new_n73_), .Y(u4__abc_76448_new_n74_));
INVX1 INVX1_687 ( .A(u4__abc_76448_new_n77_), .Y(u4__abc_76448_new_n78_));
INVX1 INVX1_688 ( .A(u4__abc_76448_new_n82_), .Y(u4__abc_76448_new_n83_));
INVX1 INVX1_689 ( .A(u4__abc_76448_new_n86_), .Y(u4__abc_76448_new_n87_));
INVX1 INVX1_69 ( .A(u0_csc_mask_2_), .Y(u0_u0__abc_72207_new_n532_));
INVX1 INVX1_690 ( .A(rfr_ps_val_0_), .Y(u4__abc_76448_new_n91_));
INVX1 INVX1_691 ( .A(u4_ps_cnt_0_), .Y(u4__abc_76448_new_n93_));
INVX1 INVX1_692 ( .A(rfr_ps_val_1_), .Y(u4__abc_76448_new_n96_));
INVX1 INVX1_693 ( .A(u4_ps_cnt_1_), .Y(u4__abc_76448_new_n98_));
INVX1 INVX1_694 ( .A(rfr_ps_val_4_), .Y(u4__abc_76448_new_n102_));
INVX1 INVX1_695 ( .A(u4_ps_cnt_4_), .Y(u4__abc_76448_new_n104_));
INVX1 INVX1_696 ( .A(u4_ps_cnt_5_), .Y(u4__abc_76448_new_n107_));
INVX1 INVX1_697 ( .A(rfr_ps_val_5_), .Y(u4__abc_76448_new_n109_));
INVX1 INVX1_698 ( .A(u4__abc_76448_new_n114_), .Y(u4__0rfr_early_0_0_));
INVX1 INVX1_699 ( .A(u4__abc_76448_new_n119_), .Y(u4__abc_76448_new_n120_));
INVX1 INVX1_7 ( .A(u0__abc_76628_new_n1128_), .Y(u0__abc_76628_new_n1136_));
INVX1 INVX1_70 ( .A(u0_csc0_18_), .Y(u0_u0__abc_72207_new_n533_));
INVX1 INVX1_700 ( .A(u4__abc_76448_new_n124_), .Y(u4__abc_76448_new_n125_));
INVX1 INVX1_701 ( .A(u4__abc_76448_new_n131_), .Y(u4__abc_76448_new_n132_));
INVX1 INVX1_702 ( .A(u4__abc_76448_new_n137_), .Y(u4__abc_76448_new_n138_));
INVX1 INVX1_703 ( .A(u4__abc_76448_new_n145_), .Y(u4__abc_76448_new_n146_));
INVX1 INVX1_704 ( .A(u4__abc_76448_new_n150_), .Y(u4__abc_76448_new_n151_));
INVX1 INVX1_705 ( .A(u4__abc_76448_new_n157_), .Y(u4__abc_76448_new_n158_));
INVX1 INVX1_706 ( .A(u4__abc_76448_new_n161_), .Y(u4__abc_76448_new_n162_));
INVX1 INVX1_707 ( .A(rfr_ps_val_6_), .Y(u4__abc_76448_new_n167_));
INVX1 INVX1_708 ( .A(rfr_ps_val_7_), .Y(u4__abc_76448_new_n168_));
INVX1 INVX1_709 ( .A(rfr_ps_val_2_), .Y(u4__abc_76448_new_n172_));
INVX1 INVX1_71 ( .A(\wb_addr_i[23] ), .Y(u0_u0__abc_72207_new_n534_));
INVX1 INVX1_710 ( .A(rfr_ps_val_3_), .Y(u4__abc_76448_new_n173_));
INVX1 INVX1_711 ( .A(u4__abc_76448_new_n177_), .Y(u4_ps_cnt_clr));
INVX1 INVX1_712 ( .A(u4__abc_76448_new_n179_), .Y(u4__abc_76448_new_n180_));
INVX1 INVX1_713 ( .A(u4__abc_76448_new_n184_), .Y(u4__abc_76448_new_n185_));
INVX1 INVX1_714 ( .A(u4__abc_76448_new_n190_), .Y(u4__abc_76448_new_n191_));
INVX1 INVX1_715 ( .A(u4__abc_76448_new_n195_), .Y(u4__abc_76448_new_n196_));
INVX1 INVX1_716 ( .A(u4__abc_76448_new_n200_), .Y(u4__abc_76448_new_n201_));
INVX1 INVX1_717 ( .A(u4__abc_76448_new_n206_), .Y(u4__abc_76448_new_n207_));
INVX1 INVX1_718 ( .A(u4_ps_cnt_6_), .Y(u4__abc_76448_new_n211_));
INVX1 INVX1_719 ( .A(u4__abc_76448_new_n217_), .Y(u4__abc_76448_new_n218_));
INVX1 INVX1_72 ( .A(u0_u0__abc_72207_new_n538_), .Y(u0_u0__abc_72207_new_n539_));
INVX1 INVX1_720 ( .A(ref_int_2_), .Y(u4__abc_76448_new_n222_));
INVX1 INVX1_721 ( .A(ref_int_1_), .Y(u4__abc_76448_new_n228_));
INVX1 INVX1_722 ( .A(u5_burst_cnt_3_), .Y(u5__abc_81276_new_n366_));
INVX1 INVX1_723 ( .A(u5_burst_cnt_2_), .Y(u5__abc_81276_new_n367_));
INVX1 INVX1_724 ( .A(u5_burst_cnt_1_), .Y(u5__abc_81276_new_n368_));
INVX1 INVX1_725 ( .A(u5_burst_cnt_0_), .Y(u5__abc_81276_new_n369_));
INVX1 INVX1_726 ( .A(u5_burst_cnt_5_), .Y(u5__abc_81276_new_n373_));
INVX1 INVX1_727 ( .A(u5_burst_cnt_4_), .Y(u5__abc_81276_new_n374_));
INVX1 INVX1_728 ( .A(u5_burst_cnt_7_), .Y(u5__abc_81276_new_n376_));
INVX1 INVX1_729 ( .A(u5_burst_cnt_6_), .Y(u5__abc_81276_new_n377_));
INVX1 INVX1_73 ( .A(u0_u0__abc_72207_new_n540_), .Y(u0_u0__abc_72207_new_n542_));
INVX1 INVX1_730 ( .A(u5_burst_cnt_10_), .Y(u5__abc_81276_new_n380_));
INVX1 INVX1_731 ( .A(u5__abc_81276_new_n381_), .Y(u5__abc_81276_new_n382_));
INVX1 INVX1_732 ( .A(u5__abc_81276_new_n385_), .Y(u5__0burst_act_rd_0_0_));
INVX1 INVX1_733 ( .A(u5_state_63_), .Y(u5__abc_81276_new_n387_));
INVX1 INVX1_734 ( .A(u5_state_62_), .Y(u5__abc_81276_new_n388_));
INVX1 INVX1_735 ( .A(u5_state_61_), .Y(u5__abc_81276_new_n390_));
INVX1 INVX1_736 ( .A(u5_state_60_), .Y(u5__abc_81276_new_n391_));
INVX1 INVX1_737 ( .A(u5_state_59_), .Y(u5__abc_81276_new_n394_));
INVX1 INVX1_738 ( .A(u5_state_58_), .Y(u5__abc_81276_new_n395_));
INVX1 INVX1_739 ( .A(u5_state_57_), .Y(u5__abc_81276_new_n397_));
INVX1 INVX1_74 ( .A(u0_u0__abc_72207_new_n546_), .Y(u0_u0__abc_72207_new_n547_));
INVX1 INVX1_740 ( .A(u5_state_56_), .Y(u5__abc_81276_new_n398_));
INVX1 INVX1_741 ( .A(u5_state_55_), .Y(u5__abc_81276_new_n402_));
INVX1 INVX1_742 ( .A(u5_state_54_), .Y(u5__abc_81276_new_n403_));
INVX1 INVX1_743 ( .A(u5_state_53_), .Y(u5__abc_81276_new_n405_));
INVX1 INVX1_744 ( .A(u5_state_52_), .Y(u5__abc_81276_new_n406_));
INVX1 INVX1_745 ( .A(u5_state_51_), .Y(u5__abc_81276_new_n409_));
INVX1 INVX1_746 ( .A(u5_state_50_), .Y(u5__abc_81276_new_n410_));
INVX1 INVX1_747 ( .A(u5_state_49_), .Y(u5__abc_81276_new_n412_));
INVX1 INVX1_748 ( .A(u5_state_48_), .Y(u5__abc_81276_new_n413_));
INVX1 INVX1_749 ( .A(u5_state_47_), .Y(u5__abc_81276_new_n418_));
INVX1 INVX1_75 ( .A(u0_u0__abc_72207_new_n548_), .Y(u0_u0__abc_72207_new_n550_));
INVX1 INVX1_750 ( .A(u5_state_46_), .Y(u5__abc_81276_new_n419_));
INVX1 INVX1_751 ( .A(u5_state_45_), .Y(u5__abc_81276_new_n421_));
INVX1 INVX1_752 ( .A(u5_state_44_), .Y(u5__abc_81276_new_n422_));
INVX1 INVX1_753 ( .A(u5_state_43_), .Y(u5__abc_81276_new_n425_));
INVX1 INVX1_754 ( .A(u5_state_42_), .Y(u5__abc_81276_new_n426_));
INVX1 INVX1_755 ( .A(u5_state_40_), .Y(u5__abc_81276_new_n428_));
INVX1 INVX1_756 ( .A(u5_state_41_), .Y(u5__abc_81276_new_n429_));
INVX1 INVX1_757 ( .A(u5_state_39_), .Y(u5__abc_81276_new_n433_));
INVX1 INVX1_758 ( .A(u5_state_38_), .Y(u5__abc_81276_new_n434_));
INVX1 INVX1_759 ( .A(u5_state_37_), .Y(u5__abc_81276_new_n436_));
INVX1 INVX1_76 ( .A(u0_u0__abc_72207_new_n553_), .Y(u0_u0__abc_72207_new_n554_));
INVX1 INVX1_760 ( .A(u5_state_36_), .Y(u5__abc_81276_new_n437_));
INVX1 INVX1_761 ( .A(u5_state_35_), .Y(u5__abc_81276_new_n440_));
INVX1 INVX1_762 ( .A(u5_state_34_), .Y(u5__abc_81276_new_n441_));
INVX1 INVX1_763 ( .A(u5_state_32_), .Y(u5__abc_81276_new_n443_));
INVX1 INVX1_764 ( .A(u5_state_33_), .Y(u5__abc_81276_new_n444_));
INVX1 INVX1_765 ( .A(u5_state_15_), .Y(u5__abc_81276_new_n450_));
INVX1 INVX1_766 ( .A(u5_state_14_), .Y(u5__abc_81276_new_n451_));
INVX1 INVX1_767 ( .A(u5_state_12_), .Y(u5__abc_81276_new_n453_));
INVX1 INVX1_768 ( .A(u5_state_13_), .Y(u5__abc_81276_new_n454_));
INVX1 INVX1_769 ( .A(u5_state_11_), .Y(u5__abc_81276_new_n457_));
INVX1 INVX1_77 ( .A(u0_u0__abc_72207_new_n555_), .Y(u0_u0__abc_72207_new_n557_));
INVX1 INVX1_770 ( .A(u5_state_10_), .Y(u5__abc_81276_new_n458_));
INVX1 INVX1_771 ( .A(u5_state_9_), .Y(u5__abc_81276_new_n460_));
INVX1 INVX1_772 ( .A(u5_state_8_), .Y(u5__abc_81276_new_n461_));
INVX1 INVX1_773 ( .A(u5_state_7_), .Y(u5__abc_81276_new_n465_));
INVX1 INVX1_774 ( .A(u5_state_6_), .Y(u5__abc_81276_new_n466_));
INVX1 INVX1_775 ( .A(u5_state_5_), .Y(u5__abc_81276_new_n468_));
INVX1 INVX1_776 ( .A(u5_state_4_), .Y(u5__abc_81276_new_n469_));
INVX1 INVX1_777 ( .A(u5_state_3_), .Y(u5__abc_81276_new_n472_));
INVX1 INVX1_778 ( .A(u5_state_2_), .Y(u5__abc_81276_new_n473_));
INVX1 INVX1_779 ( .A(u5_state_1_), .Y(u5__abc_81276_new_n475_));
INVX1 INVX1_78 ( .A(u0_u0__abc_72207_new_n499_), .Y(u0_u0__abc_72207_new_n565_));
INVX1 INVX1_780 ( .A(u5_state_0_), .Y(u5__abc_81276_new_n476_));
INVX1 INVX1_781 ( .A(u5_state_19_), .Y(u5__abc_81276_new_n481_));
INVX1 INVX1_782 ( .A(u5_state_18_), .Y(u5__abc_81276_new_n482_));
INVX1 INVX1_783 ( .A(u5_state_17_), .Y(u5__abc_81276_new_n484_));
INVX1 INVX1_784 ( .A(u5_state_16_), .Y(u5__abc_81276_new_n485_));
INVX1 INVX1_785 ( .A(u5_state_65_), .Y(u5__abc_81276_new_n488_));
INVX1 INVX1_786 ( .A(u5_state_64_), .Y(u5__abc_81276_new_n489_));
INVX1 INVX1_787 ( .A(u5_state_20_), .Y(u5__abc_81276_new_n491_));
INVX1 INVX1_788 ( .A(u5_state_21_), .Y(u5__abc_81276_new_n492_));
INVX1 INVX1_789 ( .A(u5_state_23_), .Y(u5__abc_81276_new_n494_));
INVX1 INVX1_79 ( .A(u0_init_ack0), .Y(u0_u0__abc_72207_new_n568_));
INVX1 INVX1_790 ( .A(u5_state_22_), .Y(u5__abc_81276_new_n495_));
INVX1 INVX1_791 ( .A(u5_state_27_), .Y(u5__abc_81276_new_n502_));
INVX1 INVX1_792 ( .A(u5_state_26_), .Y(u5__abc_81276_new_n503_));
INVX1 INVX1_793 ( .A(u5_state_25_), .Y(u5__abc_81276_new_n505_));
INVX1 INVX1_794 ( .A(u5_state_24_), .Y(u5__abc_81276_new_n506_));
INVX1 INVX1_795 ( .A(u5_state_29_), .Y(u5__abc_81276_new_n509_));
INVX1 INVX1_796 ( .A(u5_state_28_), .Y(u5__abc_81276_new_n510_));
INVX1 INVX1_797 ( .A(u5_state_31_), .Y(u5__abc_81276_new_n512_));
INVX1 INVX1_798 ( .A(u5_state_30_), .Y(u5__abc_81276_new_n518_));
INVX1 INVX1_799 ( .A(u5__abc_81276_new_n546_), .Y(u5__abc_81276_new_n547_));
INVX1 INVX1_8 ( .A(u0__abc_76628_new_n1135_), .Y(u0__abc_76628_new_n1142_));
INVX1 INVX1_80 ( .A(u0_u0_inited), .Y(u0_u0__abc_72207_new_n570_));
INVX1 INVX1_800 ( .A(u5__abc_81276_new_n554_), .Y(u5__abc_81276_new_n555_));
INVX1 INVX1_801 ( .A(u5__abc_81276_new_n563_), .Y(u5__abc_81276_new_n564_));
INVX1 INVX1_802 ( .A(u5__abc_81276_new_n571_), .Y(u5__abc_81276_new_n572_));
INVX1 INVX1_803 ( .A(u5__abc_81276_new_n579_), .Y(u5__abc_81276_new_n580_));
INVX1 INVX1_804 ( .A(u5__abc_81276_new_n587_), .Y(u5__abc_81276_new_n588_));
INVX1 INVX1_805 ( .A(u5__abc_81276_new_n595_), .Y(u5__abc_81276_new_n596_));
INVX1 INVX1_806 ( .A(u5__abc_81276_new_n602_), .Y(u5__abc_81276_new_n603_));
INVX1 INVX1_807 ( .A(u5__abc_81276_new_n618_), .Y(u5__abc_81276_new_n619_));
INVX1 INVX1_808 ( .A(u5__abc_81276_new_n638_), .Y(u5__abc_81276_new_n639_));
INVX1 INVX1_809 ( .A(u5__abc_81276_new_n646_), .Y(u5__abc_81276_new_n647_));
INVX1 INVX1_81 ( .A(u0_u1__abc_72579_new_n202_), .Y(u0_u1__abc_72579_new_n203_));
INVX1 INVX1_810 ( .A(u5__abc_81276_new_n654_), .Y(u5__abc_81276_new_n655_));
INVX1 INVX1_811 ( .A(u5__abc_81276_new_n496_), .Y(u5__abc_81276_new_n657_));
INVX1 INVX1_812 ( .A(u5__abc_81276_new_n658_), .Y(u5__abc_81276_new_n659_));
INVX1 INVX1_813 ( .A(u5__abc_81276_new_n665_), .Y(u5__abc_81276_new_n666_));
INVX1 INVX1_814 ( .A(u5__abc_81276_new_n686_), .Y(u5__abc_81276_new_n687_));
INVX1 INVX1_815 ( .A(u5__abc_81276_new_n694_), .Y(u5__abc_81276_new_n695_));
INVX1 INVX1_816 ( .A(u5__abc_81276_new_n702_), .Y(u5__abc_81276_new_n703_));
INVX1 INVX1_817 ( .A(u5__abc_81276_new_n712_), .Y(u5__abc_81276_new_n713_));
INVX1 INVX1_818 ( .A(u5__abc_81276_new_n720_), .Y(u5__abc_81276_new_n721_));
INVX1 INVX1_819 ( .A(u5__abc_81276_new_n727_), .Y(u5__abc_81276_new_n728_));
INVX1 INVX1_82 ( .A(u0_u1__abc_72579_new_n204_), .Y(u0_u1__abc_72579_new_n206_));
INVX1 INVX1_820 ( .A(u5__abc_81276_new_n735_), .Y(u5__abc_81276_new_n736_));
INVX1 INVX1_821 ( .A(u5__abc_81276_new_n745_), .Y(u5__abc_81276_new_n746_));
INVX1 INVX1_822 ( .A(u5__abc_81276_new_n752_), .Y(u5__abc_81276_new_n753_));
INVX1 INVX1_823 ( .A(u5__abc_81276_new_n768_), .Y(u5__abc_81276_new_n769_));
INVX1 INVX1_824 ( .A(u5__abc_81276_new_n775_), .Y(u5__abc_81276_new_n776_));
INVX1 INVX1_825 ( .A(u5__abc_81276_new_n782_), .Y(u5__abc_81276_new_n783_));
INVX1 INVX1_826 ( .A(u5__abc_81276_new_n791_), .Y(u5__abc_81276_new_n792_));
INVX1 INVX1_827 ( .A(u5__abc_81276_new_n799_), .Y(u5__abc_81276_new_n800_));
INVX1 INVX1_828 ( .A(u5__abc_81276_new_n811_), .Y(u5__abc_81276_new_n812_));
INVX1 INVX1_829 ( .A(u5__abc_81276_new_n819_), .Y(u5__abc_81276_new_n820_));
INVX1 INVX1_83 ( .A(u0_lmr_ack1), .Y(u0_u1__abc_72579_new_n207_));
INVX1 INVX1_830 ( .A(u5__abc_81276_new_n828_), .Y(u5__abc_81276_new_n829_));
INVX1 INVX1_831 ( .A(u5__abc_81276_new_n836_), .Y(u5__abc_81276_new_n837_));
INVX1 INVX1_832 ( .A(u5__abc_81276_new_n845_), .Y(u5__abc_81276_new_n846_));
INVX1 INVX1_833 ( .A(u5__abc_81276_new_n853_), .Y(u5__abc_81276_new_n854_));
INVX1 INVX1_834 ( .A(u5__abc_81276_new_n862_), .Y(u5__abc_81276_new_n863_));
INVX1 INVX1_835 ( .A(u5__abc_81276_new_n870_), .Y(u5__abc_81276_new_n871_));
INVX1 INVX1_836 ( .A(u5__abc_81276_new_n881_), .Y(u5__abc_81276_new_n882_));
INVX1 INVX1_837 ( .A(u5__abc_81276_new_n889_), .Y(u5__abc_81276_new_n890_));
INVX1 INVX1_838 ( .A(u5__abc_81276_new_n898_), .Y(u5__abc_81276_new_n899_));
INVX1 INVX1_839 ( .A(u5__abc_81276_new_n905_), .Y(u5__abc_81276_new_n906_));
INVX1 INVX1_84 ( .A(u0_u1_addr_r_5_), .Y(u0_u1__abc_72579_new_n211_));
INVX1 INVX1_840 ( .A(u5__abc_81276_new_n915_), .Y(u5__abc_81276_new_n916_));
INVX1 INVX1_841 ( .A(u5__abc_81276_new_n921_), .Y(u5__abc_81276_new_n922_));
INVX1 INVX1_842 ( .A(u5__abc_81276_new_n926_), .Y(u5__abc_81276_new_n927_));
INVX1 INVX1_843 ( .A(u5__abc_81276_new_n935_), .Y(u5__abc_81276_new_n936_));
INVX1 INVX1_844 ( .A(u5__abc_81276_new_n943_), .Y(u5__abc_81276_new_n944_));
INVX1 INVX1_845 ( .A(u5__abc_81276_new_n958_), .Y(u5__abc_81276_new_n959_));
INVX1 INVX1_846 ( .A(u5__abc_81276_new_n991_), .Y(u5__abc_81276_new_n992_));
INVX1 INVX1_847 ( .A(u5__abc_81276_new_n1002_), .Y(u5__abc_81276_new_n1003_));
INVX1 INVX1_848 ( .A(u5_dv_r), .Y(u5__abc_81276_new_n1009_));
INVX1 INVX1_849 ( .A(u5__abc_81276_new_n1017_), .Y(u5__abc_81276_new_n1018_));
INVX1 INVX1_85 ( .A(u0_u1_addr_r_6_), .Y(u0_u1__abc_72579_new_n213_));
INVX1 INVX1_850 ( .A(u5__abc_81276_new_n1025_), .Y(u5__abc_81276_new_n1026_));
INVX1 INVX1_851 ( .A(u5__abc_81276_new_n1033_), .Y(u5__abc_81276_new_n1034_));
INVX1 INVX1_852 ( .A(u5__abc_81276_new_n1041_), .Y(u5__abc_81276_new_n1042_));
INVX1 INVX1_853 ( .A(u5__abc_81276_new_n1050_), .Y(u5__abc_81276_new_n1051_));
INVX1 INVX1_854 ( .A(u5__abc_81276_new_n1068_), .Y(u5__abc_81276_new_n1069_));
INVX1 INVX1_855 ( .A(u5__abc_81276_new_n1076_), .Y(u5__abc_81276_new_n1077_));
INVX1 INVX1_856 ( .A(u5__abc_81276_new_n1084_), .Y(u5__abc_81276_new_n1085_));
INVX1 INVX1_857 ( .A(u5_cnt), .Y(u5__abc_81276_new_n1094_));
INVX1 INVX1_858 ( .A(u5_timer_1_), .Y(u5__abc_81276_new_n1101_));
INVX1 INVX1_859 ( .A(u5_timer_0_), .Y(u5__abc_81276_new_n1102_));
INVX1 INVX1_86 ( .A(\wb_data_i[0] ), .Y(u0_u1__abc_72579_new_n220_));
INVX1 INVX1_860 ( .A(u5_timer_3_), .Y(u5__abc_81276_new_n1104_));
INVX1 INVX1_861 ( .A(u5_timer_2_), .Y(u5__abc_81276_new_n1105_));
INVX1 INVX1_862 ( .A(u5_timer_5_), .Y(u5__abc_81276_new_n1108_));
INVX1 INVX1_863 ( .A(u5_timer_4_), .Y(u5__abc_81276_new_n1109_));
INVX1 INVX1_864 ( .A(u5_timer_7_), .Y(u5__abc_81276_new_n1111_));
INVX1 INVX1_865 ( .A(u5_timer_6_), .Y(u5__abc_81276_new_n1112_));
INVX1 INVX1_866 ( .A(u5_ir_cnt_1_), .Y(u5__abc_81276_new_n1116_));
INVX1 INVX1_867 ( .A(u5_ir_cnt_0_), .Y(u5__abc_81276_new_n1117_));
INVX1 INVX1_868 ( .A(u5_ir_cnt_3_), .Y(u5__abc_81276_new_n1119_));
INVX1 INVX1_869 ( .A(u5_ir_cnt_2_), .Y(u5__abc_81276_new_n1120_));
INVX1 INVX1_87 ( .A(u0_u1__abc_72579_new_n221_), .Y(u0_u1__abc_72579_new_n222_));
INVX1 INVX1_870 ( .A(u3_wb_read_go), .Y(u5__abc_81276_new_n1124_));
INVX1 INVX1_871 ( .A(u5__abc_81276_new_n1132_), .Y(u5__abc_81276_new_n1133_));
INVX1 INVX1_872 ( .A(u5__abc_81276_new_n1141_), .Y(u5__abc_81276_new_n1142_));
INVX1 INVX1_873 ( .A(u5__abc_81276_new_n1146_), .Y(u5__abc_81276_new_n1147_));
INVX1 INVX1_874 ( .A(u5__abc_81276_new_n1155_), .Y(u5__abc_81276_new_n1156_));
INVX1 INVX1_875 ( .A(u5__abc_81276_new_n1160_), .Y(u5__abc_81276_new_n1161_));
INVX1 INVX1_876 ( .A(u5__abc_81276_new_n1170_), .Y(u5__abc_81276_new_n1171_));
INVX1 INVX1_877 ( .A(u5__abc_81276_new_n1181_), .Y(u5__abc_81276_new_n1182_));
INVX1 INVX1_878 ( .A(u5__abc_81276_new_n523__bF_buf2), .Y(u5__abc_81276_new_n1183_));
INVX1 INVX1_879 ( .A(u5__abc_81276_new_n1184_), .Y(u5__abc_81276_new_n1185_));
INVX1 INVX1_88 ( .A(\wb_data_i[1] ), .Y(u0_u1__abc_72579_new_n226_));
INVX1 INVX1_880 ( .A(u5__abc_81276_new_n415_), .Y(u5__abc_81276_new_n1186_));
INVX1 INVX1_881 ( .A(u5__abc_81276_new_n407_), .Y(u5__abc_81276_new_n1187_));
INVX1 INVX1_882 ( .A(u5__abc_81276_new_n1206_), .Y(u5__abc_81276_new_n1207_));
INVX1 INVX1_883 ( .A(u5__abc_81276_new_n1215_), .Y(u5__abc_81276_new_n1216_));
INVX1 INVX1_884 ( .A(u5__abc_81276_new_n1210_), .Y(u5__abc_81276_new_n1217_));
INVX1 INVX1_885 ( .A(u5__abc_81276_new_n448__bF_buf1), .Y(u5__abc_81276_new_n1218_));
INVX1 INVX1_886 ( .A(u5__abc_81276_new_n399_), .Y(u5__abc_81276_new_n1219_));
INVX1 INVX1_887 ( .A(u5__abc_81276_new_n1231_), .Y(u5__abc_81276_new_n1232_));
INVX1 INVX1_888 ( .A(u5__abc_81276_new_n1237_), .Y(u5__abc_81276_new_n1238_));
INVX1 INVX1_889 ( .A(u5__abc_81276_new_n1247_), .Y(u5__abc_81276_new_n1248_));
INVX1 INVX1_89 ( .A(u0_u1__abc_72579_new_n227_), .Y(u0_u1__abc_72579_new_n228_));
INVX1 INVX1_890 ( .A(u5__abc_81276_new_n1260_), .Y(u5__abc_81276_new_n1261_));
INVX1 INVX1_891 ( .A(u5__abc_81276_new_n1266_), .Y(u5__abc_81276_new_n1267_));
INVX1 INVX1_892 ( .A(u5__abc_81276_new_n1270_), .Y(u5__abc_81276_new_n1271_));
INVX1 INVX1_893 ( .A(u5__abc_81276_new_n1272_), .Y(u5__abc_81276_new_n1273_));
INVX1 INVX1_894 ( .A(u5__abc_81276_new_n1281_), .Y(u5__abc_81276_new_n1282_));
INVX1 INVX1_895 ( .A(u5__abc_81276_new_n1287_), .Y(u5__abc_81276_new_n1288_));
INVX1 INVX1_896 ( .A(u5__abc_81276_new_n1296_), .Y(u5__abc_81276_new_n1297_));
INVX1 INVX1_897 ( .A(u5__abc_81276_new_n1302_), .Y(u5__abc_81276_new_n1303_));
INVX1 INVX1_898 ( .A(u5__abc_81276_new_n1309_), .Y(u5__abc_81276_new_n1310_));
INVX1 INVX1_899 ( .A(u5__abc_81276_new_n1315_), .Y(u5__abc_81276_new_n1316_));
INVX1 INVX1_9 ( .A(u0__abc_76628_new_n1145_), .Y(u0__abc_76628_new_n1153_));
INVX1 INVX1_90 ( .A(\wb_data_i[2] ), .Y(u0_u1__abc_72579_new_n232_));
INVX1 INVX1_900 ( .A(u5__abc_81276_new_n1323_), .Y(u5__abc_81276_new_n1324_));
INVX1 INVX1_901 ( .A(u5__abc_81276_new_n1329_), .Y(u5__abc_81276_new_n1330_));
INVX1 INVX1_902 ( .A(u5__abc_81276_new_n1336_), .Y(u5__abc_81276_new_n1337_));
INVX1 INVX1_903 ( .A(u5__abc_81276_new_n1342_), .Y(u5__abc_81276_new_n1343_));
INVX1 INVX1_904 ( .A(u5__abc_81276_new_n1351_), .Y(u5__abc_81276_new_n1352_));
INVX1 INVX1_905 ( .A(u5__abc_81276_new_n1360_), .Y(u5__abc_81276_new_n1361_));
INVX1 INVX1_906 ( .A(u5__abc_81276_new_n1363_), .Y(u5__abc_81276_new_n1364_));
INVX1 INVX1_907 ( .A(u5__abc_81276_new_n1368_), .Y(u5__abc_81276_new_n1369_));
INVX1 INVX1_908 ( .A(u5__abc_81276_new_n1372_), .Y(u5__abc_81276_new_n1373_));
INVX1 INVX1_909 ( .A(u5__abc_81276_new_n516_), .Y(u5__abc_81276_new_n1379_));
INVX1 INVX1_91 ( .A(u0_u1__abc_72579_new_n233_), .Y(u0_u1__abc_72579_new_n234_));
INVX1 INVX1_910 ( .A(u5__abc_81276_new_n1382_), .Y(u5__abc_81276_new_n1383_));
INVX1 INVX1_911 ( .A(u5__abc_81276_new_n1390_), .Y(u5__abc_81276_new_n1391_));
INVX1 INVX1_912 ( .A(u5__abc_81276_new_n449__bF_buf5), .Y(u5__abc_81276_new_n1392_));
INVX1 INVX1_913 ( .A(u5__abc_81276_new_n480__bF_buf2), .Y(u5__abc_81276_new_n1393_));
INVX1 INVX1_914 ( .A(u5__abc_81276_new_n521__bF_buf3), .Y(u5__abc_81276_new_n1394_));
INVX1 INVX1_915 ( .A(u5__abc_81276_new_n1405_), .Y(u5__abc_81276_new_n1406_));
INVX1 INVX1_916 ( .A(u5__abc_81276_new_n1412_), .Y(u5__abc_81276_new_n1413_));
INVX1 INVX1_917 ( .A(u5__abc_81276_new_n537_), .Y(u5__abc_81276_new_n1416_));
INVX1 INVX1_918 ( .A(u5__abc_81276_new_n1421_), .Y(u5__abc_81276_new_n1422_));
INVX1 INVX1_919 ( .A(u5__abc_81276_new_n1433_), .Y(u5__abc_81276_new_n1434_));
INVX1 INVX1_92 ( .A(\wb_data_i[3] ), .Y(u0_u1__abc_72579_new_n238_));
INVX1 INVX1_920 ( .A(u5__abc_81276_new_n1443_), .Y(u5__abc_81276_new_n1444_));
INVX1 INVX1_921 ( .A(u5__abc_81276_new_n1450_), .Y(u5__abc_81276_new_n1451_));
INVX1 INVX1_922 ( .A(u5__abc_81276_new_n1464_), .Y(u5__abc_81276_new_n1465_));
INVX1 INVX1_923 ( .A(u5__abc_81276_new_n1472_), .Y(u5__abc_81276_new_n1473_));
INVX1 INVX1_924 ( .A(u5__abc_81276_new_n1478_), .Y(u5__abc_81276_new_n1479_));
INVX1 INVX1_925 ( .A(u5__abc_81276_new_n1486_), .Y(u5__abc_81276_new_n1487_));
INVX1 INVX1_926 ( .A(u5__abc_81276_new_n1492_), .Y(u5__abc_81276_new_n1493_));
INVX1 INVX1_927 ( .A(u5__abc_81276_new_n1504_), .Y(u5__abc_81276_new_n1505_));
INVX1 INVX1_928 ( .A(u5__abc_81276_new_n1507_), .Y(u5__abc_81276_new_n1508_));
INVX1 INVX1_929 ( .A(u5__abc_81276_new_n1518_), .Y(u5__abc_81276_new_n1519_));
INVX1 INVX1_93 ( .A(u0_u1__abc_72579_new_n239_), .Y(u0_u1__abc_72579_new_n240_));
INVX1 INVX1_930 ( .A(u5__abc_81276_new_n1512_), .Y(u5__abc_81276_new_n1528_));
INVX1 INVX1_931 ( .A(u5__abc_81276_new_n1506_), .Y(u5__abc_81276_new_n1529_));
INVX1 INVX1_932 ( .A(csc_s_3_), .Y(u5__abc_81276_new_n1533_));
INVX1 INVX1_933 ( .A(u5__abc_81276_new_n1538_), .Y(u5__abc_81276_new_n1539_));
INVX1 INVX1_934 ( .A(u5__0no_wb_cycle_0_0_), .Y(u5__abc_81276_new_n1547_));
INVX1 INVX1_935 ( .A(u5__abc_81276_new_n1550_), .Y(u5__abc_81276_new_n1551_));
INVX1 INVX1_936 ( .A(u5_wb_cycle), .Y(u5__abc_81276_new_n1552_));
INVX1 INVX1_937 ( .A(u5__abc_81276_new_n1553_), .Y(u5__abc_81276_new_n1554_));
INVX1 INVX1_938 ( .A(init_req), .Y(u5__abc_81276_new_n1556_));
INVX1 INVX1_939 ( .A(rfr_req), .Y(u5__abc_81276_new_n1557_));
INVX1 INVX1_94 ( .A(\wb_data_i[4] ), .Y(u0_u1__abc_72579_new_n244_));
INVX1 INVX1_940 ( .A(u5__abc_81276_new_n1560_), .Y(u5__abc_81276_new_n1561_));
INVX1 INVX1_941 ( .A(u5_kro), .Y(u5__abc_81276_new_n1585_));
INVX1 INVX1_942 ( .A(u5__abc_81276_new_n1586_), .Y(u5__abc_81276_new_n1587_));
INVX1 INVX1_943 ( .A(u5__abc_81276_new_n1588_), .Y(u5__abc_81276_new_n1589_));
INVX1 INVX1_944 ( .A(tms_s_1_), .Y(u5__abc_81276_new_n1605_));
INVX1 INVX1_945 ( .A(tms_s_0_), .Y(u5__abc_81276_new_n1606_));
INVX1 INVX1_946 ( .A(tms_s_2_), .Y(u5__abc_81276_new_n1607_));
INVX1 INVX1_947 ( .A(u5_wb_write_go_r), .Y(u5__abc_81276_new_n1612_));
INVX1 INVX1_948 ( .A(u5__abc_81276_new_n1610_), .Y(u5__abc_81276_new_n1613_));
INVX1 INVX1_949 ( .A(u5__abc_81276_new_n1617_), .Y(u5__abc_81276_new_n1618_));
INVX1 INVX1_95 ( .A(u0_u1__abc_72579_new_n245_), .Y(u0_u1__abc_72579_new_n246_));
INVX1 INVX1_950 ( .A(u5__abc_81276_new_n1621_), .Y(u5__abc_81276_new_n1622_));
INVX1 INVX1_951 ( .A(u5__abc_81276_new_n1623_), .Y(u5__abc_81276_new_n1624_));
INVX1 INVX1_952 ( .A(u5__abc_81276_new_n1627_), .Y(u5__abc_81276_new_n1628_));
INVX1 INVX1_953 ( .A(u5__abc_81276_new_n1633_), .Y(u5__abc_81276_new_n1634_));
INVX1 INVX1_954 ( .A(u5__abc_81276_new_n1602_), .Y(u5__abc_81276_new_n1640_));
INVX1 INVX1_955 ( .A(u5__abc_81276_new_n1584_), .Y(u5__abc_81276_new_n1643_));
INVX1 INVX1_956 ( .A(u5__abc_81276_new_n1647_), .Y(u5__abc_81276_new_n1648_));
INVX1 INVX1_957 ( .A(u5__abc_81276_new_n1651_), .Y(u5__abc_81276_new_n1652_));
INVX1 INVX1_958 ( .A(u5__abc_81276_new_n1604_), .Y(u5__abc_81276_new_n1654_));
INVX1 INVX1_959 ( .A(u5__abc_81276_new_n1611_), .Y(u5__abc_81276_new_n1655_));
INVX1 INVX1_96 ( .A(\wb_data_i[5] ), .Y(u0_u1__abc_72579_new_n250_));
INVX1 INVX1_960 ( .A(u5__abc_81276_new_n1666_), .Y(u5__abc_81276_new_n1667_));
INVX1 INVX1_961 ( .A(u5__abc_81276_new_n1672_), .Y(u5__abc_81276_new_n1673_));
INVX1 INVX1_962 ( .A(u5__abc_81276_new_n1678_), .Y(u5__abc_81276_new_n1679_));
INVX1 INVX1_963 ( .A(u5__abc_81276_new_n1680_), .Y(u5__abc_81276_new_n1681_));
INVX1 INVX1_964 ( .A(csc_s_2_), .Y(u5__abc_81276_new_n1688_));
INVX1 INVX1_965 ( .A(csc_s_1_), .Y(u5__abc_81276_new_n1690_));
INVX1 INVX1_966 ( .A(u5__abc_81276_new_n1691_), .Y(u5__abc_81276_new_n1692_));
INVX1 INVX1_967 ( .A(u5_wb_wait_r), .Y(u5__abc_81276_new_n1699_));
INVX1 INVX1_968 ( .A(u5__abc_81276_new_n1629_), .Y(u5__abc_81276_new_n1705_));
INVX1 INVX1_969 ( .A(u5__abc_81276_new_n1706_), .Y(u5__abc_81276_new_n1707_));
INVX1 INVX1_97 ( .A(u0_u1__abc_72579_new_n251_), .Y(u0_u1__abc_72579_new_n252_));
INVX1 INVX1_970 ( .A(u5__abc_81276_new_n1668_), .Y(u5__abc_81276_new_n1731_));
INVX1 INVX1_971 ( .A(csc_s_4_), .Y(u5__abc_81276_new_n1749_));
INVX1 INVX1_972 ( .A(csc_s_5_), .Y(u5__abc_81276_new_n1750_));
INVX1 INVX1_973 ( .A(u5__abc_81276_new_n1768_), .Y(u5__abc_81276_new_n1769_));
INVX1 INVX1_974 ( .A(u5_ack_cnt_3_), .Y(u5__abc_81276_new_n1815_));
INVX1 INVX1_975 ( .A(u5_ack_cnt_2_), .Y(u5__abc_81276_new_n1816_));
INVX1 INVX1_976 ( .A(u5__abc_81276_new_n1817_), .Y(u5__abc_81276_new_n1818_));
INVX1 INVX1_977 ( .A(u5__abc_81276_new_n1820_), .Y(u5__abc_81276_new_n1821_));
INVX1 INVX1_978 ( .A(u5__abc_81276_new_n1822_), .Y(u5__abc_81276_new_n1823_));
INVX1 INVX1_979 ( .A(u5_mem_ack_r), .Y(u5__abc_81276_new_n1824_));
INVX1 INVX1_98 ( .A(\wb_data_i[6] ), .Y(u0_u1__abc_72579_new_n256_));
INVX1 INVX1_980 ( .A(u5__abc_81276_new_n1828_), .Y(u5__abc_81276_new_n1829_));
INVX1 INVX1_981 ( .A(u5__abc_81276_new_n1609_), .Y(u5__abc_81276_new_n1834_));
INVX1 INVX1_982 ( .A(u5__abc_81276_new_n1847_), .Y(u5__abc_81276_new_n1848_));
INVX1 INVX1_983 ( .A(u5__abc_81276_new_n1857_), .Y(u5__abc_81276_new_n1858_));
INVX1 INVX1_984 ( .A(u5__abc_81276_new_n1859_), .Y(u5__abc_81276_new_n1860_));
INVX1 INVX1_985 ( .A(u5__abc_81276_new_n1862_), .Y(u5__abc_81276_new_n1863_));
INVX1 INVX1_986 ( .A(u5__abc_81276_new_n1865_), .Y(mem_ack));
INVX1 INVX1_987 ( .A(u5__abc_81276_new_n1835_), .Y(u5__abc_81276_new_n1870_));
INVX1 INVX1_988 ( .A(u5__abc_81276_new_n1878_), .Y(u5__abc_81276_new_n1879_));
INVX1 INVX1_989 ( .A(u5__abc_81276_new_n1928_), .Y(u5__abc_81276_new_n1929_));
INVX1 INVX1_99 ( .A(u0_u1__abc_72579_new_n257_), .Y(u0_u1__abc_72579_new_n258_));
INVX1 INVX1_990 ( .A(u5__abc_81276_new_n1935_), .Y(u5__abc_81276_new_n1936_));
INVX1 INVX1_991 ( .A(u5__abc_81276_new_n1941_), .Y(u5__abc_81276_new_n1942_));
INVX1 INVX1_992 ( .A(u5__abc_81276_new_n1947_), .Y(u5__abc_81276_new_n1948_));
INVX1 INVX1_993 ( .A(u5__abc_81276_new_n1955_), .Y(u5__abc_81276_new_n1956_));
INVX1 INVX1_994 ( .A(u5__abc_81276_new_n1959_), .Y(u5__abc_81276_new_n1960_));
INVX1 INVX1_995 ( .A(u5__abc_81276_new_n1963_), .Y(u5__abc_81276_new_n1964_));
INVX1 INVX1_996 ( .A(u5__abc_81276_new_n1976_), .Y(u5__abc_81276_new_n1977_));
INVX1 INVX1_997 ( .A(u5__abc_81276_new_n1989_), .Y(u5__abc_81276_new_n1990_));
INVX1 INVX1_998 ( .A(u5__abc_81276_new_n2003_), .Y(u5__abc_81276_new_n2004_));
INVX1 INVX1_999 ( .A(u5__abc_81276_new_n2014_), .Y(u5__abc_81276_new_n2015_));
INVX2 INVX2_1 ( .A(init_req), .Y(u0__abc_76628_new_n1100_));
INVX2 INVX2_10 ( .A(row_adr_6_bF_buf1_), .Y(u2_u0__abc_74955_new_n169_));
INVX2 INVX2_11 ( .A(row_adr_7_bF_buf1_), .Y(u2_u0__abc_74955_new_n174_));
INVX2 INVX2_12 ( .A(row_adr_8_bF_buf1_), .Y(u2_u0__abc_74955_new_n179_));
INVX2 INVX2_13 ( .A(row_adr_9_bF_buf1_), .Y(u2_u0__abc_74955_new_n184_));
INVX2 INVX2_14 ( .A(row_adr_10_bF_buf1_), .Y(u2_u0__abc_74955_new_n189_));
INVX2 INVX2_15 ( .A(row_adr_11_bF_buf1_), .Y(u2_u0__abc_74955_new_n194_));
INVX2 INVX2_16 ( .A(row_adr_12_bF_buf1_), .Y(u2_u0__abc_74955_new_n199_));
INVX2 INVX2_17 ( .A(rst_i), .Y(u2_u0__abc_74955_auto_rtlil_cc_1942_NotGate_71538));
INVX2 INVX2_18 ( .A(row_adr_0_bF_buf1_), .Y(u2_u1__abc_74955_new_n139_));
INVX2 INVX2_19 ( .A(row_adr_1_bF_buf1_), .Y(u2_u1__abc_74955_new_n144_));
INVX2 INVX2_2 ( .A(u0_sreq_cs_le), .Y(u0__abc_76628_new_n1109_));
INVX2 INVX2_20 ( .A(row_adr_2_bF_buf1_), .Y(u2_u1__abc_74955_new_n149_));
INVX2 INVX2_21 ( .A(row_adr_3_bF_buf1_), .Y(u2_u1__abc_74955_new_n154_));
INVX2 INVX2_22 ( .A(row_adr_4_bF_buf1_), .Y(u2_u1__abc_74955_new_n159_));
INVX2 INVX2_23 ( .A(row_adr_5_bF_buf1_), .Y(u2_u1__abc_74955_new_n164_));
INVX2 INVX2_24 ( .A(row_adr_6_bF_buf1_), .Y(u2_u1__abc_74955_new_n169_));
INVX2 INVX2_25 ( .A(row_adr_7_bF_buf1_), .Y(u2_u1__abc_74955_new_n174_));
INVX2 INVX2_26 ( .A(row_adr_8_bF_buf1_), .Y(u2_u1__abc_74955_new_n179_));
INVX2 INVX2_27 ( .A(row_adr_9_bF_buf1_), .Y(u2_u1__abc_74955_new_n184_));
INVX2 INVX2_28 ( .A(row_adr_10_bF_buf1_), .Y(u2_u1__abc_74955_new_n189_));
INVX2 INVX2_29 ( .A(row_adr_11_bF_buf1_), .Y(u2_u1__abc_74955_new_n194_));
INVX2 INVX2_3 ( .A(\wb_addr_i[6] ), .Y(u0__abc_76628_new_n4515_));
INVX2 INVX2_30 ( .A(row_adr_12_bF_buf1_), .Y(u2_u1__abc_74955_new_n199_));
INVX2 INVX2_31 ( .A(rst_i), .Y(u2_u1__abc_74955_auto_rtlil_cc_1942_NotGate_71538));
INVX2 INVX2_32 ( .A(u3_rd_fifo_clr), .Y(u3_u0__abc_75526_new_n858_));
INVX2 INVX2_33 ( .A(rfr_ack), .Y(u4__abc_76448_new_n116_));
INVX2 INVX2_34 ( .A(ref_int_0_), .Y(u4__abc_76448_new_n223_));
INVX2 INVX2_35 ( .A(u5__abc_81276_new_n611_), .Y(u5__abc_81276_new_n612_));
INVX2 INVX2_36 ( .A(u5__abc_81276_new_n624_), .Y(u5__abc_81276_new_n625_));
INVX2 INVX2_37 ( .A(u5__abc_81276_new_n629_), .Y(u5__abc_81276_new_n630_));
INVX2 INVX2_38 ( .A(u5__abc_81276_new_n490__bF_buf1), .Y(u5__abc_81276_new_n656_));
INVX2 INVX2_39 ( .A(u5__abc_81276_new_n950_), .Y(u5__abc_81276_new_n951_));
INVX2 INVX2_4 ( .A(row_adr_0_bF_buf1_), .Y(u2_u0__abc_74955_new_n139_));
INVX2 INVX2_40 ( .A(u5__abc_81276_new_n994_), .Y(u5__abc_81276_new_n995_));
INVX2 INVX2_41 ( .A(u5_mc_le), .Y(u5__0mc_le_0_0_));
INVX2 INVX2_42 ( .A(u1_wb_write_go), .Y(u5__abc_81276_new_n1123_));
INVX2 INVX2_43 ( .A(u5__abc_81276_new_n1200_), .Y(u5__abc_81276_new_n1201_));
INVX2 INVX2_44 ( .A(u5__abc_81276_new_n1253_), .Y(u5__abc_81276_new_n1254_));
INVX2 INVX2_45 ( .A(u5__abc_81276_new_n1356_), .Y(u5__abc_81276_new_n1357_));
INVX2 INVX2_46 ( .A(u5__abc_81276_new_n530_), .Y(u5__abc_81276_new_n1378_));
INVX2 INVX2_47 ( .A(u5__abc_81276_new_n1428_), .Y(u5__abc_81276_new_n1429_));
INVX2 INVX2_48 ( .A(u5__abc_81276_new_n1457_), .Y(u5__abc_81276_new_n1458_));
INVX2 INVX2_49 ( .A(u5__abc_81276_new_n1500_), .Y(u5__abc_81276_new_n1501_));
INVX2 INVX2_5 ( .A(row_adr_1_bF_buf1_), .Y(u2_u0__abc_74955_new_n144_));
INVX2 INVX2_50 ( .A(u5__abc_81276_new_n1510_), .Y(u5__abc_81276_new_n1511_));
INVX2 INVX2_51 ( .A(u1_wr_cycle), .Y(u5__abc_81276_new_n1637_));
INVX2 INVX2_52 ( .A(u5__abc_81276_new_n1225_), .Y(u5__abc_81276_new_n1849_));
INVX2 INVX2_53 ( .A(u5__abc_81276_new_n2307_), .Y(u5__abc_81276_new_n2308_));
INVX2 INVX2_54 ( .A(u5__abc_81276_new_n2501_), .Y(u5__abc_81276_new_n2563_));
INVX2 INVX2_55 ( .A(u5__abc_81276_new_n2639_), .Y(u5__abc_81276_new_n2640_));
INVX2 INVX2_56 ( .A(u5__abc_81276_new_n2653_), .Y(u5__abc_81276_new_n2654_));
INVX2 INVX2_57 ( .A(u5__abc_81276_new_n2668_), .Y(u5__abc_81276_new_n2673_));
INVX2 INVX2_58 ( .A(u5__abc_81276_new_n2925_), .Y(u5__abc_81276_new_n2926_));
INVX2 INVX2_59 ( .A(u5__abc_81276_new_n3009_), .Y(u5__abc_81276_new_n3010_));
INVX2 INVX2_6 ( .A(row_adr_2_bF_buf1_), .Y(u2_u0__abc_74955_new_n149_));
INVX2 INVX2_60 ( .A(u5__abc_81276_new_n1549_), .Y(u5__abc_81276_new_n3211_));
INVX2 INVX2_61 ( .A(u5_ap_en), .Y(u5__abc_81276_new_n3238_));
INVX2 INVX2_62 ( .A(u5__abc_81276_new_n1836_), .Y(u5__abc_81276_new_n3239_));
INVX2 INVX2_63 ( .A(u5__abc_81276_new_n1620_), .Y(u5__abc_81276_new_n3248_));
INVX2 INVX2_64 ( .A(u7__abc_74830_new_n106_), .Y(u7__abc_74830_new_n107_));
INVX2 INVX2_65 ( .A(cs_en), .Y(u7__abc_74830_new_n114_));
INVX2 INVX2_7 ( .A(row_adr_3_bF_buf1_), .Y(u2_u0__abc_74955_new_n154_));
INVX2 INVX2_8 ( .A(row_adr_4_bF_buf1_), .Y(u2_u0__abc_74955_new_n159_));
INVX2 INVX2_9 ( .A(row_adr_5_bF_buf1_), .Y(u2_u0__abc_74955_new_n164_));
INVX4 INVX4_1 ( .A(_abc_85006_new_n237_), .Y(_abc_85006_new_n245_));
INVX4 INVX4_10 ( .A(u1__abc_73140_new_n527_), .Y(u1__abc_73140_new_n528_));
INVX4 INVX4_11 ( .A(u1__abc_73140_new_n900__bF_buf3), .Y(u1__abc_73140_new_n913_));
INVX4 INVX4_12 ( .A(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n919_));
INVX4 INVX4_13 ( .A(row_sel), .Y(u1__abc_73140_new_n921_));
INVX4 INVX4_14 ( .A(u2_u0__abc_74955_new_n206_), .Y(u2_u0__abc_74955_new_n208_));
INVX4 INVX4_15 ( .A(u2_u0__abc_74955_new_n248_), .Y(u2_u0__abc_74955_new_n250_));
INVX4 INVX4_16 ( .A(u2_u0__abc_74955_new_n290_), .Y(u2_u0__abc_74955_new_n292_));
INVX4 INVX4_17 ( .A(u2_u1__abc_74955_new_n206_), .Y(u2_u1__abc_74955_new_n208_));
INVX4 INVX4_18 ( .A(u2_u1__abc_74955_new_n248_), .Y(u2_u1__abc_74955_new_n250_));
INVX4 INVX4_19 ( .A(u2_u1__abc_74955_new_n290_), .Y(u2_u1__abc_74955_new_n292_));
INVX4 INVX4_2 ( .A(u0__abc_76628_new_n1946__bF_buf3), .Y(u0__abc_76628_new_n1947_));
INVX4 INVX4_20 ( .A(pack_le2), .Y(u3__abc_74070_new_n424_));
INVX4 INVX4_21 ( .A(u3__abc_74070_new_n453_), .Y(u3__abc_74070_new_n454_));
INVX4 INVX4_22 ( .A(u3__abc_74070_new_n451_), .Y(u3__abc_74070_new_n459_));
INVX4 INVX4_23 ( .A(pack_le0), .Y(u3__abc_74070_new_n505_));
INVX4 INVX4_24 ( .A(rst_i), .Y(u3_u0__abc_75526_auto_rtlil_cc_1942_NotGate_71546));
INVX4 INVX4_25 ( .A(u5_wb_wait), .Y(u5__abc_81276_new_n1536_));
INVX4 INVX4_26 ( .A(u5_tmr2_done), .Y(u5__abc_81276_new_n1708_));
INVX4 INVX4_27 ( .A(u5_tmr_done_bF_buf1), .Y(u5__abc_81276_new_n1712_));
INVX4 INVX4_28 ( .A(u5__abc_81276_new_n2298_), .Y(u5__abc_81276_new_n2299_));
INVX4 INVX4_29 ( .A(u5_cmd_asserted_bF_buf1), .Y(u5__abc_81276_new_n2953_));
INVX4 INVX4_3 ( .A(cs_le_bF_buf2), .Y(u0__abc_76628_new_n4273_));
INVX4 INVX4_30 ( .A(rst_i), .Y(u7__abc_74830_auto_rtlil_cc_1942_NotGate_71518));
INVX4 INVX4_4 ( .A(u0__abc_76628_new_n4401_), .Y(u0__abc_76628_new_n4403_));
INVX4 INVX4_5 ( .A(rst_i), .Y(u0_u0__abc_72207_auto_rtlil_cc_1942_NotGate_71494));
INVX4 INVX4_6 ( .A(rst_i), .Y(u0_u1__abc_72579_auto_rtlil_cc_1942_NotGate_71506));
INVX4 INVX4_7 ( .A(cs_le_bF_buf4), .Y(u1__abc_73140_new_n282_));
INVX4 INVX4_8 ( .A(u1__abc_73140_new_n272_), .Y(page_size_9_));
INVX4 INVX4_9 ( .A(u1_bas_bF_buf2), .Y(u1__abc_73140_new_n314_));
INVX8 INVX8_1 ( .A(u0__abc_76628_new_n1169__bF_buf6), .Y(u0__abc_76628_new_n1170_));
INVX8 INVX8_10 ( .A(1'h0), .Y(u0__abc_76628_new_n2718_));
INVX8 INVX8_11 ( .A(1'h0), .Y(u0__abc_76628_new_n2719_));
INVX8 INVX8_12 ( .A(1'h0), .Y(u0__abc_76628_new_n2720_));
INVX8 INVX8_13 ( .A(1'h0), .Y(u0__abc_76628_new_n2722_));
INVX8 INVX8_14 ( .A(1'h0), .Y(u0__abc_76628_new_n2724_));
INVX8 INVX8_15 ( .A(u0_cs0_bF_buf4), .Y(u0__abc_76628_new_n2742_));
INVX8 INVX8_16 ( .A(u0_rst_r3_bF_buf3), .Y(u0__abc_76628_new_n4298_));
INVX8 INVX8_17 ( .A(u0__abc_76628_new_n4437__bF_buf3), .Y(u0__abc_76628_new_n4438_));
INVX8 INVX8_18 ( .A(rst_i), .Y(u0__abc_76628_auto_rtlil_cc_1942_NotGate_71602));
INVX8 INVX8_19 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf3_), .Y(u0_u0__abc_72207_new_n224_));
INVX8 INVX8_2 ( .A(spec_req_cs_1_bF_buf3_), .Y(u0__abc_76628_new_n1172_));
INVX8 INVX8_20 ( .A(u0_u0_rst_r2_bF_buf3), .Y(u0_u0__abc_72207_new_n354_));
INVX8 INVX8_21 ( .A(u0_u1_rst_r2), .Y(u0_u1__abc_72579_new_n219_));
INVX8 INVX8_22 ( .A(next_adr_bF_buf3), .Y(u1__abc_73140_new_n563_));
INVX8 INVX8_23 ( .A(u1__abc_73140_new_n561__bF_buf3), .Y(u1__abc_73140_new_n570_));
INVX8 INVX8_24 ( .A(wb_stb_i_bF_buf1), .Y(u1__abc_73140_new_n826_));
INVX8 INVX8_25 ( .A(u1__abc_73140_new_n904__bF_buf3), .Y(u1__abc_73140_new_n906_));
INVX8 INVX8_26 ( .A(u1__abc_73140_new_n911_), .Y(u1__abc_73140_new_n912_));
INVX8 INVX8_27 ( .A(u3__abc_74070_new_n277__bF_buf4), .Y(u3__abc_74070_new_n279_));
INVX8 INVX8_28 ( .A(csc_5_bF_buf2_), .Y(u3__abc_74070_new_n449_));
INVX8 INVX8_29 ( .A(u3__abc_74070_new_n275__bF_buf3), .Y(u3__abc_74070_new_n625_));
INVX8 INVX8_3 ( .A(spec_req_cs_2_bF_buf3_), .Y(u0__abc_76628_new_n1173_));
INVX8 INVX8_30 ( .A(rst_i), .Y(u4__abc_76448_auto_rtlil_cc_1942_NotGate_71562));
INVX8 INVX8_31 ( .A(rst_i), .Y(u5__abc_81276_auto_rtlil_cc_1942_NotGate_71962));
INVX8 INVX8_32 ( .A(u6__abc_85257_new_n145__bF_buf3), .Y(u6__abc_85257_new_n155_));
INVX8 INVX8_33 ( .A(rst_i), .Y(u6__abc_85257_auto_rtlil_cc_1942_NotGate_72188));
INVX8 INVX8_4 ( .A(spec_req_cs_3_bF_buf3_), .Y(u0__abc_76628_new_n1174_));
INVX8 INVX8_5 ( .A(spec_req_cs_4_bF_buf3_), .Y(u0__abc_76628_new_n1175_));
INVX8 INVX8_6 ( .A(spec_req_cs_6_bF_buf3_), .Y(u0__abc_76628_new_n1177_));
INVX8 INVX8_7 ( .A(spec_req_cs_5_bF_buf2_), .Y(u0__abc_76628_new_n1179_));
INVX8 INVX8_8 ( .A(spec_req_cs_0_bF_buf2_), .Y(u0__abc_76628_new_n1197_));
INVX8 INVX8_9 ( .A(u0_cs1_bF_buf5), .Y(u0__abc_76628_new_n2717_));
OR2X2 OR2X2_1 ( .A(init_ack), .B(lmr_ack), .Y(lmr_sel));
OR2X2 OR2X2_10 ( .A(_abc_85006_new_n245_), .B(cs_need_rfr_1_), .Y(_abc_85006_new_n252_));
OR2X2 OR2X2_100 ( .A(lmr_sel_bF_buf1), .B(csc_5_bF_buf4_), .Y(_abc_85006_new_n402_));
OR2X2 OR2X2_1000 ( .A(u0__abc_76628_new_n4438__bF_buf0), .B(u0_csr_4_), .Y(u0__abc_76628_new_n4448_));
OR2X2 OR2X2_1001 ( .A(u0__abc_76628_new_n4437__bF_buf3), .B(\wb_data_i[4] ), .Y(u0__abc_76628_new_n4449_));
OR2X2 OR2X2_1002 ( .A(u0__abc_76628_new_n4438__bF_buf3), .B(u0_csr_5_), .Y(u0__abc_76628_new_n4451_));
OR2X2 OR2X2_1003 ( .A(u0__abc_76628_new_n4437__bF_buf2), .B(\wb_data_i[5] ), .Y(u0__abc_76628_new_n4452_));
OR2X2 OR2X2_1004 ( .A(u0__abc_76628_new_n4438__bF_buf2), .B(u0_csr_6_), .Y(u0__abc_76628_new_n4454_));
OR2X2 OR2X2_1005 ( .A(u0__abc_76628_new_n4437__bF_buf1), .B(\wb_data_i[6] ), .Y(u0__abc_76628_new_n4455_));
OR2X2 OR2X2_1006 ( .A(u0__abc_76628_new_n4438__bF_buf1), .B(u0_csr_7_), .Y(u0__abc_76628_new_n4457_));
OR2X2 OR2X2_1007 ( .A(u0__abc_76628_new_n4437__bF_buf0), .B(\wb_data_i[7] ), .Y(u0__abc_76628_new_n4458_));
OR2X2 OR2X2_1008 ( .A(u0__abc_76628_new_n4438__bF_buf0), .B(ref_int_0_), .Y(u0__abc_76628_new_n4460_));
OR2X2 OR2X2_1009 ( .A(u0__abc_76628_new_n4437__bF_buf3), .B(\wb_data_i[8] ), .Y(u0__abc_76628_new_n4461_));
OR2X2 OR2X2_101 ( .A(_abc_85006_new_n240__bF_buf0), .B(sp_csc_6_), .Y(_abc_85006_new_n404_));
OR2X2 OR2X2_1010 ( .A(u0__abc_76628_new_n4438__bF_buf3), .B(ref_int_1_), .Y(u0__abc_76628_new_n4463_));
OR2X2 OR2X2_1011 ( .A(u0__abc_76628_new_n4437__bF_buf2), .B(\wb_data_i[9] ), .Y(u0__abc_76628_new_n4464_));
OR2X2 OR2X2_1012 ( .A(u0__abc_76628_new_n4438__bF_buf2), .B(ref_int_2_), .Y(u0__abc_76628_new_n4466_));
OR2X2 OR2X2_1013 ( .A(u0__abc_76628_new_n4437__bF_buf1), .B(\wb_data_i[10] ), .Y(u0__abc_76628_new_n4467_));
OR2X2 OR2X2_1014 ( .A(u0__abc_76628_new_n4438__bF_buf1), .B(rfr_ps_val_0_), .Y(u0__abc_76628_new_n4469_));
OR2X2 OR2X2_1015 ( .A(u0__abc_76628_new_n4437__bF_buf0), .B(\wb_data_i[24] ), .Y(u0__abc_76628_new_n4470_));
OR2X2 OR2X2_1016 ( .A(u0__abc_76628_new_n4438__bF_buf0), .B(rfr_ps_val_1_), .Y(u0__abc_76628_new_n4472_));
OR2X2 OR2X2_1017 ( .A(u0__abc_76628_new_n4437__bF_buf3), .B(\wb_data_i[25] ), .Y(u0__abc_76628_new_n4473_));
OR2X2 OR2X2_1018 ( .A(u0__abc_76628_new_n4438__bF_buf3), .B(rfr_ps_val_2_), .Y(u0__abc_76628_new_n4475_));
OR2X2 OR2X2_1019 ( .A(u0__abc_76628_new_n4437__bF_buf2), .B(\wb_data_i[26] ), .Y(u0__abc_76628_new_n4476_));
OR2X2 OR2X2_102 ( .A(lmr_sel_bF_buf0), .B(csc_6_), .Y(_abc_85006_new_n405_));
OR2X2 OR2X2_1020 ( .A(u0__abc_76628_new_n4438__bF_buf2), .B(rfr_ps_val_3_), .Y(u0__abc_76628_new_n4478_));
OR2X2 OR2X2_1021 ( .A(u0__abc_76628_new_n4437__bF_buf1), .B(\wb_data_i[27] ), .Y(u0__abc_76628_new_n4479_));
OR2X2 OR2X2_1022 ( .A(u0__abc_76628_new_n4438__bF_buf1), .B(rfr_ps_val_4_), .Y(u0__abc_76628_new_n4481_));
OR2X2 OR2X2_1023 ( .A(u0__abc_76628_new_n4437__bF_buf0), .B(\wb_data_i[28] ), .Y(u0__abc_76628_new_n4482_));
OR2X2 OR2X2_1024 ( .A(u0__abc_76628_new_n4438__bF_buf0), .B(rfr_ps_val_5_), .Y(u0__abc_76628_new_n4484_));
OR2X2 OR2X2_1025 ( .A(u0__abc_76628_new_n4437__bF_buf3), .B(\wb_data_i[29] ), .Y(u0__abc_76628_new_n4485_));
OR2X2 OR2X2_1026 ( .A(u0__abc_76628_new_n4438__bF_buf3), .B(rfr_ps_val_6_), .Y(u0__abc_76628_new_n4487_));
OR2X2 OR2X2_1027 ( .A(u0__abc_76628_new_n4437__bF_buf2), .B(\wb_data_i[30] ), .Y(u0__abc_76628_new_n4488_));
OR2X2 OR2X2_1028 ( .A(u0__abc_76628_new_n4438__bF_buf2), .B(rfr_ps_val_7_), .Y(u0__abc_76628_new_n4490_));
OR2X2 OR2X2_1029 ( .A(u0__abc_76628_new_n4437__bF_buf1), .B(\wb_data_i[31] ), .Y(u0__abc_76628_new_n4491_));
OR2X2 OR2X2_103 ( .A(_abc_85006_new_n240__bF_buf5), .B(sp_csc_7_), .Y(_abc_85006_new_n407_));
OR2X2 OR2X2_1030 ( .A(u0__abc_76628_new_n4501_), .B(u0__abc_76628_new_n4504_), .Y(u0__abc_76628_new_n4505_));
OR2X2 OR2X2_1031 ( .A(u0__abc_76628_new_n4508_), .B(u0__abc_76628_new_n4511_), .Y(u0__abc_76628_new_n4512_));
OR2X2 OR2X2_1032 ( .A(u0__abc_76628_new_n4505_), .B(u0__abc_76628_new_n4512_), .Y(u0__abc_76628_new_n4513_));
OR2X2 OR2X2_1033 ( .A(u0__abc_76628_new_n4521_), .B(u0__abc_76628_new_n4524_), .Y(u0__abc_76628_new_n4525_));
OR2X2 OR2X2_1034 ( .A(u0__abc_76628_new_n4525_), .B(u0__abc_76628_new_n4518_), .Y(u0__abc_76628_new_n4526_));
OR2X2 OR2X2_1035 ( .A(u0__abc_76628_new_n4529_), .B(u0__abc_76628_new_n4532_), .Y(u0__abc_76628_new_n4533_));
OR2X2 OR2X2_1036 ( .A(u0__abc_76628_new_n4526_), .B(u0__abc_76628_new_n4533_), .Y(u0__abc_76628_new_n4534_));
OR2X2 OR2X2_1037 ( .A(u0__abc_76628_new_n4534_), .B(u0__abc_76628_new_n4513_), .Y(u0__abc_76628_new_n4535_));
OR2X2 OR2X2_1038 ( .A(u0__abc_76628_new_n4499_), .B(u0__abc_76628_new_n4506_), .Y(u0__abc_76628_new_n4539_));
OR2X2 OR2X2_1039 ( .A(u0__abc_76628_new_n4540_), .B(u0__abc_76628_new_n4537_), .Y(u0__abc_76628_new_n4541_));
OR2X2 OR2X2_104 ( .A(lmr_sel_bF_buf6), .B(csc_7_), .Y(_abc_85006_new_n408_));
OR2X2 OR2X2_1040 ( .A(u0__abc_76628_new_n4548_), .B(u0__abc_76628_new_n4550_), .Y(u0__abc_76628_new_n4551_));
OR2X2 OR2X2_1041 ( .A(u0__abc_76628_new_n4551_), .B(u0__abc_76628_new_n4546_), .Y(u0__abc_76628_new_n4552_));
OR2X2 OR2X2_1042 ( .A(u0__abc_76628_new_n4552_), .B(u0__abc_76628_new_n4542_), .Y(u0__abc_76628_new_n4553_));
OR2X2 OR2X2_1043 ( .A(u0__abc_76628_new_n4559_), .B(u0__abc_76628_new_n4557_), .Y(u0__abc_76628_new_n4560_));
OR2X2 OR2X2_1044 ( .A(u0__abc_76628_new_n4560_), .B(u0__abc_76628_new_n4555_), .Y(u0__abc_76628_new_n4561_));
OR2X2 OR2X2_1045 ( .A(u0__abc_76628_new_n4565_), .B(u0__abc_76628_new_n4567_), .Y(u0__abc_76628_new_n4568_));
OR2X2 OR2X2_1046 ( .A(u0__abc_76628_new_n4568_), .B(u0__abc_76628_new_n4563_), .Y(u0__abc_76628_new_n4569_));
OR2X2 OR2X2_1047 ( .A(u0__abc_76628_new_n4561_), .B(u0__abc_76628_new_n4569_), .Y(u0__abc_76628_new_n4570_));
OR2X2 OR2X2_1048 ( .A(u0__abc_76628_new_n4570_), .B(u0__abc_76628_new_n4553_), .Y(u0__abc_76628_new_n4571_));
OR2X2 OR2X2_1049 ( .A(u0__abc_76628_new_n4571_), .B(u0__abc_76628_new_n4535_), .Y(rf_dout_0_));
OR2X2 OR2X2_105 ( .A(_abc_85006_new_n240__bF_buf4), .B(sp_csc_9_), .Y(_abc_85006_new_n413_));
OR2X2 OR2X2_1050 ( .A(u0__abc_76628_new_n4573_), .B(u0__abc_76628_new_n4574_), .Y(u0__abc_76628_new_n4575_));
OR2X2 OR2X2_1051 ( .A(u0__abc_76628_new_n4576_), .B(u0__abc_76628_new_n4577_), .Y(u0__abc_76628_new_n4578_));
OR2X2 OR2X2_1052 ( .A(u0__abc_76628_new_n4579_), .B(u0__abc_76628_new_n4580_), .Y(u0__abc_76628_new_n4581_));
OR2X2 OR2X2_1053 ( .A(u0__abc_76628_new_n4578_), .B(u0__abc_76628_new_n4581_), .Y(u0__abc_76628_new_n4582_));
OR2X2 OR2X2_1054 ( .A(u0__abc_76628_new_n4582_), .B(u0__abc_76628_new_n4575_), .Y(u0__abc_76628_new_n4583_));
OR2X2 OR2X2_1055 ( .A(u0__abc_76628_new_n4584_), .B(u0__abc_76628_new_n4585_), .Y(u0__abc_76628_new_n4586_));
OR2X2 OR2X2_1056 ( .A(u0__abc_76628_new_n4588_), .B(u0__abc_76628_new_n4587_), .Y(u0__abc_76628_new_n4589_));
OR2X2 OR2X2_1057 ( .A(u0__abc_76628_new_n4586_), .B(u0__abc_76628_new_n4589_), .Y(u0__abc_76628_new_n4590_));
OR2X2 OR2X2_1058 ( .A(u0__abc_76628_new_n4591_), .B(u0__abc_76628_new_n4592_), .Y(u0__abc_76628_new_n4593_));
OR2X2 OR2X2_1059 ( .A(u0__abc_76628_new_n4594_), .B(u0__abc_76628_new_n4595_), .Y(u0__abc_76628_new_n4596_));
OR2X2 OR2X2_106 ( .A(lmr_sel_bF_buf5), .B(csc_9_), .Y(_abc_85006_new_n414_));
OR2X2 OR2X2_1060 ( .A(u0__abc_76628_new_n4596_), .B(u0__abc_76628_new_n4593_), .Y(u0__abc_76628_new_n4597_));
OR2X2 OR2X2_1061 ( .A(u0__abc_76628_new_n4590_), .B(u0__abc_76628_new_n4597_), .Y(u0__abc_76628_new_n4598_));
OR2X2 OR2X2_1062 ( .A(u0__abc_76628_new_n4600_), .B(u0__abc_76628_new_n4601_), .Y(u0__abc_76628_new_n4602_));
OR2X2 OR2X2_1063 ( .A(u0__abc_76628_new_n4603_), .B(u0__abc_76628_new_n4604_), .Y(u0__abc_76628_new_n4605_));
OR2X2 OR2X2_1064 ( .A(u0__abc_76628_new_n4602_), .B(u0__abc_76628_new_n4605_), .Y(u0__abc_76628_new_n4606_));
OR2X2 OR2X2_1065 ( .A(u0__abc_76628_new_n4606_), .B(u0__abc_76628_new_n4599_), .Y(u0__abc_76628_new_n4607_));
OR2X2 OR2X2_1066 ( .A(u0__abc_76628_new_n4598_), .B(u0__abc_76628_new_n4607_), .Y(u0__abc_76628_new_n4608_));
OR2X2 OR2X2_1067 ( .A(u0__abc_76628_new_n4608_), .B(u0__abc_76628_new_n4583_), .Y(rf_dout_1_));
OR2X2 OR2X2_1068 ( .A(u0__abc_76628_new_n4610_), .B(u0__abc_76628_new_n4611_), .Y(u0__abc_76628_new_n4612_));
OR2X2 OR2X2_1069 ( .A(u0__abc_76628_new_n4613_), .B(u0__abc_76628_new_n4614_), .Y(u0__abc_76628_new_n4615_));
OR2X2 OR2X2_107 ( .A(_abc_85006_new_n240__bF_buf3), .B(sp_csc_10_), .Y(_abc_85006_new_n416_));
OR2X2 OR2X2_1070 ( .A(u0__abc_76628_new_n4616_), .B(u0__abc_76628_new_n4617_), .Y(u0__abc_76628_new_n4618_));
OR2X2 OR2X2_1071 ( .A(u0__abc_76628_new_n4615_), .B(u0__abc_76628_new_n4618_), .Y(u0__abc_76628_new_n4619_));
OR2X2 OR2X2_1072 ( .A(u0__abc_76628_new_n4619_), .B(u0__abc_76628_new_n4612_), .Y(u0__abc_76628_new_n4620_));
OR2X2 OR2X2_1073 ( .A(u0__abc_76628_new_n4621_), .B(u0__abc_76628_new_n4622_), .Y(u0__abc_76628_new_n4623_));
OR2X2 OR2X2_1074 ( .A(u0__abc_76628_new_n4624_), .B(u0__abc_76628_new_n4625_), .Y(u0__abc_76628_new_n4626_));
OR2X2 OR2X2_1075 ( .A(u0__abc_76628_new_n4623_), .B(u0__abc_76628_new_n4626_), .Y(u0__abc_76628_new_n4627_));
OR2X2 OR2X2_1076 ( .A(u0__abc_76628_new_n4628_), .B(u0__abc_76628_new_n4629_), .Y(u0__abc_76628_new_n4630_));
OR2X2 OR2X2_1077 ( .A(u0__abc_76628_new_n4631_), .B(u0__abc_76628_new_n4632_), .Y(u0__abc_76628_new_n4633_));
OR2X2 OR2X2_1078 ( .A(u0__abc_76628_new_n4630_), .B(u0__abc_76628_new_n4633_), .Y(u0__abc_76628_new_n4634_));
OR2X2 OR2X2_1079 ( .A(u0__abc_76628_new_n4634_), .B(u0__abc_76628_new_n4627_), .Y(u0__abc_76628_new_n4635_));
OR2X2 OR2X2_108 ( .A(lmr_sel_bF_buf4), .B(csc_10_), .Y(_abc_85006_new_n417_));
OR2X2 OR2X2_1080 ( .A(u0__abc_76628_new_n4638_), .B(u0__abc_76628_new_n4637_), .Y(u0__abc_76628_new_n4639_));
OR2X2 OR2X2_1081 ( .A(u0__abc_76628_new_n4640_), .B(u0__abc_76628_new_n4641_), .Y(u0__abc_76628_new_n4642_));
OR2X2 OR2X2_1082 ( .A(u0__abc_76628_new_n4642_), .B(u0__abc_76628_new_n4639_), .Y(u0__abc_76628_new_n4643_));
OR2X2 OR2X2_1083 ( .A(u0__abc_76628_new_n4643_), .B(u0__abc_76628_new_n4636_), .Y(u0__abc_76628_new_n4644_));
OR2X2 OR2X2_1084 ( .A(u0__abc_76628_new_n4635_), .B(u0__abc_76628_new_n4644_), .Y(u0__abc_76628_new_n4645_));
OR2X2 OR2X2_1085 ( .A(u0__abc_76628_new_n4645_), .B(u0__abc_76628_new_n4620_), .Y(rf_dout_2_));
OR2X2 OR2X2_1086 ( .A(u0__abc_76628_new_n4647_), .B(u0__abc_76628_new_n4648_), .Y(u0__abc_76628_new_n4649_));
OR2X2 OR2X2_1087 ( .A(u0__abc_76628_new_n4650_), .B(u0__abc_76628_new_n4651_), .Y(u0__abc_76628_new_n4652_));
OR2X2 OR2X2_1088 ( .A(u0__abc_76628_new_n4649_), .B(u0__abc_76628_new_n4652_), .Y(u0__abc_76628_new_n4653_));
OR2X2 OR2X2_1089 ( .A(u0__abc_76628_new_n4656_), .B(u0__abc_76628_new_n4655_), .Y(u0__abc_76628_new_n4657_));
OR2X2 OR2X2_109 ( .A(\wb_addr_i[31] ), .B(\wb_addr_i[30] ), .Y(_abc_85006_new_n482_));
OR2X2 OR2X2_1090 ( .A(u0__abc_76628_new_n4657_), .B(u0__abc_76628_new_n4654_), .Y(u0__abc_76628_new_n4658_));
OR2X2 OR2X2_1091 ( .A(u0__abc_76628_new_n4659_), .B(u0__abc_76628_new_n4660_), .Y(u0__abc_76628_new_n4661_));
OR2X2 OR2X2_1092 ( .A(u0__abc_76628_new_n4658_), .B(u0__abc_76628_new_n4661_), .Y(u0__abc_76628_new_n4662_));
OR2X2 OR2X2_1093 ( .A(u0__abc_76628_new_n4662_), .B(u0__abc_76628_new_n4653_), .Y(u0__abc_76628_new_n4663_));
OR2X2 OR2X2_1094 ( .A(u0__abc_76628_new_n4665_), .B(u0__abc_76628_new_n4666_), .Y(u0__abc_76628_new_n4667_));
OR2X2 OR2X2_1095 ( .A(u0__abc_76628_new_n4667_), .B(u0__abc_76628_new_n4668_), .Y(u0__abc_76628_new_n4669_));
OR2X2 OR2X2_1096 ( .A(u0__abc_76628_new_n4669_), .B(u0__abc_76628_new_n4664_), .Y(u0__abc_76628_new_n4670_));
OR2X2 OR2X2_1097 ( .A(u0__abc_76628_new_n4673_), .B(u0__abc_76628_new_n4672_), .Y(u0__abc_76628_new_n4674_));
OR2X2 OR2X2_1098 ( .A(u0__abc_76628_new_n4674_), .B(u0__abc_76628_new_n4671_), .Y(u0__abc_76628_new_n4675_));
OR2X2 OR2X2_1099 ( .A(u0__abc_76628_new_n4677_), .B(u0__abc_76628_new_n4678_), .Y(u0__abc_76628_new_n4679_));
OR2X2 OR2X2_11 ( .A(_abc_85006_new_n240__bF_buf3), .B(spec_req_cs_2_bF_buf5_), .Y(_abc_85006_new_n254_));
OR2X2 OR2X2_110 ( .A(_abc_85006_new_n482_), .B(\wb_addr_i[29] ), .Y(_abc_85006_new_n483_));
OR2X2 OR2X2_1100 ( .A(u0__abc_76628_new_n4679_), .B(u0__abc_76628_new_n4676_), .Y(u0__abc_76628_new_n4680_));
OR2X2 OR2X2_1101 ( .A(u0__abc_76628_new_n4675_), .B(u0__abc_76628_new_n4680_), .Y(u0__abc_76628_new_n4681_));
OR2X2 OR2X2_1102 ( .A(u0__abc_76628_new_n4681_), .B(u0__abc_76628_new_n4670_), .Y(u0__abc_76628_new_n4682_));
OR2X2 OR2X2_1103 ( .A(u0__abc_76628_new_n4682_), .B(u0__abc_76628_new_n4663_), .Y(rf_dout_3_));
OR2X2 OR2X2_1104 ( .A(u0__abc_76628_new_n4684_), .B(u0__abc_76628_new_n4685_), .Y(u0__abc_76628_new_n4686_));
OR2X2 OR2X2_1105 ( .A(u0__abc_76628_new_n4687_), .B(u0__abc_76628_new_n4688_), .Y(u0__abc_76628_new_n4689_));
OR2X2 OR2X2_1106 ( .A(u0__abc_76628_new_n4690_), .B(u0__abc_76628_new_n4691_), .Y(u0__abc_76628_new_n4692_));
OR2X2 OR2X2_1107 ( .A(u0__abc_76628_new_n4689_), .B(u0__abc_76628_new_n4692_), .Y(u0__abc_76628_new_n4693_));
OR2X2 OR2X2_1108 ( .A(u0__abc_76628_new_n4693_), .B(u0__abc_76628_new_n4686_), .Y(u0__abc_76628_new_n4694_));
OR2X2 OR2X2_1109 ( .A(u0__abc_76628_new_n4695_), .B(u0__abc_76628_new_n4696_), .Y(u0__abc_76628_new_n4697_));
OR2X2 OR2X2_111 ( .A(u0__abc_76628_new_n1101_), .B(u0__abc_76628_new_n1102_), .Y(u0__abc_76628_new_n1103_));
OR2X2 OR2X2_1110 ( .A(u0__abc_76628_new_n4698_), .B(u0__abc_76628_new_n4699_), .Y(u0__abc_76628_new_n4700_));
OR2X2 OR2X2_1111 ( .A(u0__abc_76628_new_n4697_), .B(u0__abc_76628_new_n4700_), .Y(u0__abc_76628_new_n4701_));
OR2X2 OR2X2_1112 ( .A(u0__abc_76628_new_n4702_), .B(u0__abc_76628_new_n4703_), .Y(u0__abc_76628_new_n4704_));
OR2X2 OR2X2_1113 ( .A(u0__abc_76628_new_n4706_), .B(u0__abc_76628_new_n4705_), .Y(u0__abc_76628_new_n4707_));
OR2X2 OR2X2_1114 ( .A(u0__abc_76628_new_n4704_), .B(u0__abc_76628_new_n4707_), .Y(u0__abc_76628_new_n4708_));
OR2X2 OR2X2_1115 ( .A(u0__abc_76628_new_n4701_), .B(u0__abc_76628_new_n4708_), .Y(u0__abc_76628_new_n4709_));
OR2X2 OR2X2_1116 ( .A(u0__abc_76628_new_n4712_), .B(u0__abc_76628_new_n4711_), .Y(u0__abc_76628_new_n4713_));
OR2X2 OR2X2_1117 ( .A(u0__abc_76628_new_n4714_), .B(u0__abc_76628_new_n4715_), .Y(u0__abc_76628_new_n4716_));
OR2X2 OR2X2_1118 ( .A(u0__abc_76628_new_n4716_), .B(u0__abc_76628_new_n4713_), .Y(u0__abc_76628_new_n4717_));
OR2X2 OR2X2_1119 ( .A(u0__abc_76628_new_n4717_), .B(u0__abc_76628_new_n4710_), .Y(u0__abc_76628_new_n4718_));
OR2X2 OR2X2_112 ( .A(spec_req_cs_0_bF_buf4_), .B(u0_sreq_cs_le), .Y(u0__abc_76628_new_n1107_));
OR2X2 OR2X2_1120 ( .A(u0__abc_76628_new_n4709_), .B(u0__abc_76628_new_n4718_), .Y(u0__abc_76628_new_n4719_));
OR2X2 OR2X2_1121 ( .A(u0__abc_76628_new_n4719_), .B(u0__abc_76628_new_n4694_), .Y(rf_dout_4_));
OR2X2 OR2X2_1122 ( .A(u0__abc_76628_new_n4721_), .B(u0__abc_76628_new_n4722_), .Y(u0__abc_76628_new_n4723_));
OR2X2 OR2X2_1123 ( .A(u0__abc_76628_new_n4724_), .B(u0__abc_76628_new_n4725_), .Y(u0__abc_76628_new_n4726_));
OR2X2 OR2X2_1124 ( .A(u0__abc_76628_new_n4723_), .B(u0__abc_76628_new_n4726_), .Y(u0__abc_76628_new_n4727_));
OR2X2 OR2X2_1125 ( .A(u0__abc_76628_new_n4729_), .B(u0__abc_76628_new_n4730_), .Y(u0__abc_76628_new_n4731_));
OR2X2 OR2X2_1126 ( .A(u0__abc_76628_new_n4731_), .B(u0__abc_76628_new_n4728_), .Y(u0__abc_76628_new_n4732_));
OR2X2 OR2X2_1127 ( .A(u0__abc_76628_new_n4733_), .B(u0__abc_76628_new_n4734_), .Y(u0__abc_76628_new_n4735_));
OR2X2 OR2X2_1128 ( .A(u0__abc_76628_new_n4732_), .B(u0__abc_76628_new_n4735_), .Y(u0__abc_76628_new_n4736_));
OR2X2 OR2X2_1129 ( .A(u0__abc_76628_new_n4736_), .B(u0__abc_76628_new_n4727_), .Y(u0__abc_76628_new_n4737_));
OR2X2 OR2X2_113 ( .A(u0__abc_76628_new_n1111_), .B(u0__abc_76628_new_n1112_), .Y(u0__abc_76628_new_n1113_));
OR2X2 OR2X2_1130 ( .A(u0__abc_76628_new_n4740_), .B(u0__abc_76628_new_n4741_), .Y(u0__abc_76628_new_n4742_));
OR2X2 OR2X2_1131 ( .A(u0__abc_76628_new_n4742_), .B(u0__abc_76628_new_n4739_), .Y(u0__abc_76628_new_n4743_));
OR2X2 OR2X2_1132 ( .A(u0__abc_76628_new_n4743_), .B(u0__abc_76628_new_n4738_), .Y(u0__abc_76628_new_n4744_));
OR2X2 OR2X2_1133 ( .A(u0__abc_76628_new_n4746_), .B(u0__abc_76628_new_n4747_), .Y(u0__abc_76628_new_n4748_));
OR2X2 OR2X2_1134 ( .A(u0__abc_76628_new_n4748_), .B(u0__abc_76628_new_n4745_), .Y(u0__abc_76628_new_n4749_));
OR2X2 OR2X2_1135 ( .A(u0__abc_76628_new_n4751_), .B(u0__abc_76628_new_n4752_), .Y(u0__abc_76628_new_n4753_));
OR2X2 OR2X2_1136 ( .A(u0__abc_76628_new_n4753_), .B(u0__abc_76628_new_n4750_), .Y(u0__abc_76628_new_n4754_));
OR2X2 OR2X2_1137 ( .A(u0__abc_76628_new_n4749_), .B(u0__abc_76628_new_n4754_), .Y(u0__abc_76628_new_n4755_));
OR2X2 OR2X2_1138 ( .A(u0__abc_76628_new_n4755_), .B(u0__abc_76628_new_n4744_), .Y(u0__abc_76628_new_n4756_));
OR2X2 OR2X2_1139 ( .A(u0__abc_76628_new_n4756_), .B(u0__abc_76628_new_n4737_), .Y(rf_dout_5_));
OR2X2 OR2X2_114 ( .A(u0__abc_76628_new_n1114_), .B(u0__abc_76628_new_n1110_), .Y(u0__0spec_req_cs_7_0__1_));
OR2X2 OR2X2_1140 ( .A(u0__abc_76628_new_n4758_), .B(u0__abc_76628_new_n4759_), .Y(u0__abc_76628_new_n4760_));
OR2X2 OR2X2_1141 ( .A(u0__abc_76628_new_n4761_), .B(u0__abc_76628_new_n4762_), .Y(u0__abc_76628_new_n4763_));
OR2X2 OR2X2_1142 ( .A(u0__abc_76628_new_n4764_), .B(u0__abc_76628_new_n4765_), .Y(u0__abc_76628_new_n4766_));
OR2X2 OR2X2_1143 ( .A(u0__abc_76628_new_n4763_), .B(u0__abc_76628_new_n4766_), .Y(u0__abc_76628_new_n4767_));
OR2X2 OR2X2_1144 ( .A(u0__abc_76628_new_n4767_), .B(u0__abc_76628_new_n4760_), .Y(u0__abc_76628_new_n4768_));
OR2X2 OR2X2_1145 ( .A(u0__abc_76628_new_n4769_), .B(u0__abc_76628_new_n4770_), .Y(u0__abc_76628_new_n4771_));
OR2X2 OR2X2_1146 ( .A(u0__abc_76628_new_n4772_), .B(u0__abc_76628_new_n4773_), .Y(u0__abc_76628_new_n4774_));
OR2X2 OR2X2_1147 ( .A(u0__abc_76628_new_n4771_), .B(u0__abc_76628_new_n4774_), .Y(u0__abc_76628_new_n4775_));
OR2X2 OR2X2_1148 ( .A(u0__abc_76628_new_n4776_), .B(u0__abc_76628_new_n4777_), .Y(u0__abc_76628_new_n4778_));
OR2X2 OR2X2_1149 ( .A(u0__abc_76628_new_n4780_), .B(u0__abc_76628_new_n4779_), .Y(u0__abc_76628_new_n4781_));
OR2X2 OR2X2_115 ( .A(u0__abc_76628_new_n1117_), .B(u0__abc_76628_new_n1118_), .Y(u0__abc_76628_new_n1119_));
OR2X2 OR2X2_1150 ( .A(u0__abc_76628_new_n4778_), .B(u0__abc_76628_new_n4781_), .Y(u0__abc_76628_new_n4782_));
OR2X2 OR2X2_1151 ( .A(u0__abc_76628_new_n4775_), .B(u0__abc_76628_new_n4782_), .Y(u0__abc_76628_new_n4783_));
OR2X2 OR2X2_1152 ( .A(u0__abc_76628_new_n4786_), .B(u0__abc_76628_new_n4785_), .Y(u0__abc_76628_new_n4787_));
OR2X2 OR2X2_1153 ( .A(u0__abc_76628_new_n4788_), .B(u0__abc_76628_new_n4789_), .Y(u0__abc_76628_new_n4790_));
OR2X2 OR2X2_1154 ( .A(u0__abc_76628_new_n4790_), .B(u0__abc_76628_new_n4787_), .Y(u0__abc_76628_new_n4791_));
OR2X2 OR2X2_1155 ( .A(u0__abc_76628_new_n4791_), .B(u0__abc_76628_new_n4784_), .Y(u0__abc_76628_new_n4792_));
OR2X2 OR2X2_1156 ( .A(u0__abc_76628_new_n4783_), .B(u0__abc_76628_new_n4792_), .Y(u0__abc_76628_new_n4793_));
OR2X2 OR2X2_1157 ( .A(u0__abc_76628_new_n4793_), .B(u0__abc_76628_new_n4768_), .Y(rf_dout_6_));
OR2X2 OR2X2_1158 ( .A(u0__abc_76628_new_n4795_), .B(u0__abc_76628_new_n4796_), .Y(u0__abc_76628_new_n4797_));
OR2X2 OR2X2_1159 ( .A(u0__abc_76628_new_n4798_), .B(u0__abc_76628_new_n4799_), .Y(u0__abc_76628_new_n4800_));
OR2X2 OR2X2_116 ( .A(u0__abc_76628_new_n1122_), .B(u0__abc_76628_new_n1116_), .Y(u0__0spec_req_cs_7_0__2_));
OR2X2 OR2X2_1160 ( .A(u0__abc_76628_new_n4797_), .B(u0__abc_76628_new_n4800_), .Y(u0__abc_76628_new_n4801_));
OR2X2 OR2X2_1161 ( .A(u0__abc_76628_new_n4802_), .B(u0__abc_76628_new_n4803_), .Y(u0__abc_76628_new_n4804_));
OR2X2 OR2X2_1162 ( .A(u0__abc_76628_new_n4807_), .B(u0__abc_76628_new_n4806_), .Y(u0__abc_76628_new_n4808_));
OR2X2 OR2X2_1163 ( .A(u0__abc_76628_new_n4808_), .B(u0__abc_76628_new_n4805_), .Y(u0__abc_76628_new_n4809_));
OR2X2 OR2X2_1164 ( .A(u0__abc_76628_new_n4809_), .B(u0__abc_76628_new_n4804_), .Y(u0__abc_76628_new_n4810_));
OR2X2 OR2X2_1165 ( .A(u0__abc_76628_new_n4810_), .B(u0__abc_76628_new_n4801_), .Y(u0__abc_76628_new_n4811_));
OR2X2 OR2X2_1166 ( .A(u0__abc_76628_new_n4814_), .B(u0__abc_76628_new_n4815_), .Y(u0__abc_76628_new_n4816_));
OR2X2 OR2X2_1167 ( .A(u0__abc_76628_new_n4816_), .B(u0__abc_76628_new_n4813_), .Y(u0__abc_76628_new_n4817_));
OR2X2 OR2X2_1168 ( .A(u0__abc_76628_new_n4817_), .B(u0__abc_76628_new_n4812_), .Y(u0__abc_76628_new_n4818_));
OR2X2 OR2X2_1169 ( .A(u0__abc_76628_new_n4820_), .B(u0__abc_76628_new_n4821_), .Y(u0__abc_76628_new_n4822_));
OR2X2 OR2X2_117 ( .A(u0__abc_76628_new_n1126_), .B(u0__abc_76628_new_n1127_), .Y(u0__abc_76628_new_n1128_));
OR2X2 OR2X2_1170 ( .A(u0__abc_76628_new_n4822_), .B(u0__abc_76628_new_n4819_), .Y(u0__abc_76628_new_n4823_));
OR2X2 OR2X2_1171 ( .A(u0__abc_76628_new_n4825_), .B(u0__abc_76628_new_n4826_), .Y(u0__abc_76628_new_n4827_));
OR2X2 OR2X2_1172 ( .A(u0__abc_76628_new_n4827_), .B(u0__abc_76628_new_n4824_), .Y(u0__abc_76628_new_n4828_));
OR2X2 OR2X2_1173 ( .A(u0__abc_76628_new_n4823_), .B(u0__abc_76628_new_n4828_), .Y(u0__abc_76628_new_n4829_));
OR2X2 OR2X2_1174 ( .A(u0__abc_76628_new_n4829_), .B(u0__abc_76628_new_n4818_), .Y(u0__abc_76628_new_n4830_));
OR2X2 OR2X2_1175 ( .A(u0__abc_76628_new_n4830_), .B(u0__abc_76628_new_n4811_), .Y(rf_dout_7_));
OR2X2 OR2X2_1176 ( .A(u0__abc_76628_new_n4832_), .B(u0__abc_76628_new_n4833_), .Y(u0__abc_76628_new_n4834_));
OR2X2 OR2X2_1177 ( .A(u0__abc_76628_new_n4835_), .B(u0__abc_76628_new_n4836_), .Y(u0__abc_76628_new_n4837_));
OR2X2 OR2X2_1178 ( .A(u0__abc_76628_new_n4838_), .B(u0__abc_76628_new_n4839_), .Y(u0__abc_76628_new_n4840_));
OR2X2 OR2X2_1179 ( .A(u0__abc_76628_new_n4840_), .B(u0__abc_76628_new_n4837_), .Y(u0__abc_76628_new_n4841_));
OR2X2 OR2X2_118 ( .A(u0__abc_76628_new_n1130_), .B(u0__abc_76628_new_n1124_), .Y(u0__0spec_req_cs_7_0__3_));
OR2X2 OR2X2_1180 ( .A(u0__abc_76628_new_n4841_), .B(u0__abc_76628_new_n4834_), .Y(u0__abc_76628_new_n4842_));
OR2X2 OR2X2_1181 ( .A(u0__abc_76628_new_n4843_), .B(u0__abc_76628_new_n4844_), .Y(u0__abc_76628_new_n4845_));
OR2X2 OR2X2_1182 ( .A(u0__abc_76628_new_n4847_), .B(u0__abc_76628_new_n4846_), .Y(u0__abc_76628_new_n4848_));
OR2X2 OR2X2_1183 ( .A(u0__abc_76628_new_n4845_), .B(u0__abc_76628_new_n4848_), .Y(u0__abc_76628_new_n4849_));
OR2X2 OR2X2_1184 ( .A(u0__abc_76628_new_n4851_), .B(u0__abc_76628_new_n4850_), .Y(u0__abc_76628_new_n4852_));
OR2X2 OR2X2_1185 ( .A(u0__abc_76628_new_n4853_), .B(u0__abc_76628_new_n4854_), .Y(u0__abc_76628_new_n4855_));
OR2X2 OR2X2_1186 ( .A(u0__abc_76628_new_n4852_), .B(u0__abc_76628_new_n4855_), .Y(u0__abc_76628_new_n4856_));
OR2X2 OR2X2_1187 ( .A(u0__abc_76628_new_n4849_), .B(u0__abc_76628_new_n4856_), .Y(u0__abc_76628_new_n4857_));
OR2X2 OR2X2_1188 ( .A(u0__abc_76628_new_n4859_), .B(u0__abc_76628_new_n4860_), .Y(u0__abc_76628_new_n4861_));
OR2X2 OR2X2_1189 ( .A(u0__abc_76628_new_n4862_), .B(u0__abc_76628_new_n4863_), .Y(u0__abc_76628_new_n4864_));
OR2X2 OR2X2_119 ( .A(u0__abc_76628_new_n1133_), .B(u0__abc_76628_new_n1134_), .Y(u0__abc_76628_new_n1135_));
OR2X2 OR2X2_1190 ( .A(u0__abc_76628_new_n4861_), .B(u0__abc_76628_new_n4864_), .Y(u0__abc_76628_new_n4865_));
OR2X2 OR2X2_1191 ( .A(u0__abc_76628_new_n4865_), .B(u0__abc_76628_new_n4858_), .Y(u0__abc_76628_new_n4866_));
OR2X2 OR2X2_1192 ( .A(u0__abc_76628_new_n4857_), .B(u0__abc_76628_new_n4866_), .Y(u0__abc_76628_new_n4867_));
OR2X2 OR2X2_1193 ( .A(u0__abc_76628_new_n4867_), .B(u0__abc_76628_new_n4842_), .Y(rf_dout_8_));
OR2X2 OR2X2_1194 ( .A(u0__abc_76628_new_n4869_), .B(u0__abc_76628_new_n4870_), .Y(u0__abc_76628_new_n4871_));
OR2X2 OR2X2_1195 ( .A(u0__abc_76628_new_n4872_), .B(u0__abc_76628_new_n4873_), .Y(u0__abc_76628_new_n4874_));
OR2X2 OR2X2_1196 ( .A(u0__abc_76628_new_n4871_), .B(u0__abc_76628_new_n4874_), .Y(u0__abc_76628_new_n4875_));
OR2X2 OR2X2_1197 ( .A(u0__abc_76628_new_n4878_), .B(u0__abc_76628_new_n4877_), .Y(u0__abc_76628_new_n4879_));
OR2X2 OR2X2_1198 ( .A(u0__abc_76628_new_n4879_), .B(u0__abc_76628_new_n4876_), .Y(u0__abc_76628_new_n4880_));
OR2X2 OR2X2_1199 ( .A(u0__abc_76628_new_n4881_), .B(u0__abc_76628_new_n4882_), .Y(u0__abc_76628_new_n4883_));
OR2X2 OR2X2_12 ( .A(lmr_sel_bF_buf4), .B(cs_2_), .Y(_abc_85006_new_n255_));
OR2X2 OR2X2_120 ( .A(u0__abc_76628_new_n1139_), .B(u0__abc_76628_new_n1132_), .Y(u0__0spec_req_cs_7_0__4_));
OR2X2 OR2X2_1200 ( .A(u0__abc_76628_new_n4880_), .B(u0__abc_76628_new_n4883_), .Y(u0__abc_76628_new_n4884_));
OR2X2 OR2X2_1201 ( .A(u0__abc_76628_new_n4884_), .B(u0__abc_76628_new_n4875_), .Y(u0__abc_76628_new_n4885_));
OR2X2 OR2X2_1202 ( .A(u0__abc_76628_new_n4887_), .B(u0__abc_76628_new_n4888_), .Y(u0__abc_76628_new_n4889_));
OR2X2 OR2X2_1203 ( .A(u0__abc_76628_new_n4889_), .B(u0__abc_76628_new_n4890_), .Y(u0__abc_76628_new_n4891_));
OR2X2 OR2X2_1204 ( .A(u0__abc_76628_new_n4891_), .B(u0__abc_76628_new_n4886_), .Y(u0__abc_76628_new_n4892_));
OR2X2 OR2X2_1205 ( .A(u0__abc_76628_new_n4895_), .B(u0__abc_76628_new_n4894_), .Y(u0__abc_76628_new_n4896_));
OR2X2 OR2X2_1206 ( .A(u0__abc_76628_new_n4896_), .B(u0__abc_76628_new_n4893_), .Y(u0__abc_76628_new_n4897_));
OR2X2 OR2X2_1207 ( .A(u0__abc_76628_new_n4899_), .B(u0__abc_76628_new_n4900_), .Y(u0__abc_76628_new_n4901_));
OR2X2 OR2X2_1208 ( .A(u0__abc_76628_new_n4901_), .B(u0__abc_76628_new_n4898_), .Y(u0__abc_76628_new_n4902_));
OR2X2 OR2X2_1209 ( .A(u0__abc_76628_new_n4897_), .B(u0__abc_76628_new_n4902_), .Y(u0__abc_76628_new_n4903_));
OR2X2 OR2X2_121 ( .A(u0__abc_76628_new_n1143_), .B(u0__abc_76628_new_n1144_), .Y(u0__abc_76628_new_n1145_));
OR2X2 OR2X2_1210 ( .A(u0__abc_76628_new_n4903_), .B(u0__abc_76628_new_n4892_), .Y(u0__abc_76628_new_n4904_));
OR2X2 OR2X2_1211 ( .A(u0__abc_76628_new_n4904_), .B(u0__abc_76628_new_n4885_), .Y(rf_dout_9_));
OR2X2 OR2X2_1212 ( .A(u0__abc_76628_new_n4906_), .B(u0__abc_76628_new_n4907_), .Y(u0__abc_76628_new_n4908_));
OR2X2 OR2X2_1213 ( .A(u0__abc_76628_new_n4909_), .B(u0__abc_76628_new_n4910_), .Y(u0__abc_76628_new_n4911_));
OR2X2 OR2X2_1214 ( .A(u0__abc_76628_new_n4912_), .B(u0__abc_76628_new_n4913_), .Y(u0__abc_76628_new_n4914_));
OR2X2 OR2X2_1215 ( .A(u0__abc_76628_new_n4911_), .B(u0__abc_76628_new_n4914_), .Y(u0__abc_76628_new_n4915_));
OR2X2 OR2X2_1216 ( .A(u0__abc_76628_new_n4915_), .B(u0__abc_76628_new_n4908_), .Y(u0__abc_76628_new_n4916_));
OR2X2 OR2X2_1217 ( .A(u0__abc_76628_new_n4917_), .B(u0__abc_76628_new_n4918_), .Y(u0__abc_76628_new_n4919_));
OR2X2 OR2X2_1218 ( .A(u0__abc_76628_new_n4920_), .B(u0__abc_76628_new_n4921_), .Y(u0__abc_76628_new_n4922_));
OR2X2 OR2X2_1219 ( .A(u0__abc_76628_new_n4919_), .B(u0__abc_76628_new_n4922_), .Y(u0__abc_76628_new_n4923_));
OR2X2 OR2X2_122 ( .A(u0__abc_76628_new_n1147_), .B(u0__abc_76628_new_n1141_), .Y(u0__0spec_req_cs_7_0__5_));
OR2X2 OR2X2_1220 ( .A(u0__abc_76628_new_n4924_), .B(u0__abc_76628_new_n4925_), .Y(u0__abc_76628_new_n4926_));
OR2X2 OR2X2_1221 ( .A(u0__abc_76628_new_n4928_), .B(u0__abc_76628_new_n4927_), .Y(u0__abc_76628_new_n4929_));
OR2X2 OR2X2_1222 ( .A(u0__abc_76628_new_n4926_), .B(u0__abc_76628_new_n4929_), .Y(u0__abc_76628_new_n4930_));
OR2X2 OR2X2_1223 ( .A(u0__abc_76628_new_n4923_), .B(u0__abc_76628_new_n4930_), .Y(u0__abc_76628_new_n4931_));
OR2X2 OR2X2_1224 ( .A(u0__abc_76628_new_n4934_), .B(u0__abc_76628_new_n4933_), .Y(u0__abc_76628_new_n4935_));
OR2X2 OR2X2_1225 ( .A(u0__abc_76628_new_n4936_), .B(u0__abc_76628_new_n4937_), .Y(u0__abc_76628_new_n4938_));
OR2X2 OR2X2_1226 ( .A(u0__abc_76628_new_n4938_), .B(u0__abc_76628_new_n4935_), .Y(u0__abc_76628_new_n4939_));
OR2X2 OR2X2_1227 ( .A(u0__abc_76628_new_n4939_), .B(u0__abc_76628_new_n4932_), .Y(u0__abc_76628_new_n4940_));
OR2X2 OR2X2_1228 ( .A(u0__abc_76628_new_n4931_), .B(u0__abc_76628_new_n4940_), .Y(u0__abc_76628_new_n4941_));
OR2X2 OR2X2_1229 ( .A(u0__abc_76628_new_n4941_), .B(u0__abc_76628_new_n4916_), .Y(rf_dout_10_));
OR2X2 OR2X2_123 ( .A(u0__abc_76628_new_n1150_), .B(u0__abc_76628_new_n1151_), .Y(u0__abc_76628_new_n1152_));
OR2X2 OR2X2_1230 ( .A(u0__abc_76628_new_n4943_), .B(u0__abc_76628_new_n4944_), .Y(u0__abc_76628_new_n4945_));
OR2X2 OR2X2_1231 ( .A(u0__abc_76628_new_n4946_), .B(u0__abc_76628_new_n4947_), .Y(u0__abc_76628_new_n4948_));
OR2X2 OR2X2_1232 ( .A(u0__abc_76628_new_n4950_), .B(u0__abc_76628_new_n4949_), .Y(u0__abc_76628_new_n4951_));
OR2X2 OR2X2_1233 ( .A(u0__abc_76628_new_n4948_), .B(u0__abc_76628_new_n4951_), .Y(u0__abc_76628_new_n4952_));
OR2X2 OR2X2_1234 ( .A(u0__abc_76628_new_n4952_), .B(u0__abc_76628_new_n4945_), .Y(u0__abc_76628_new_n4953_));
OR2X2 OR2X2_1235 ( .A(u0__abc_76628_new_n4955_), .B(u0__abc_76628_new_n4956_), .Y(u0__abc_76628_new_n4957_));
OR2X2 OR2X2_1236 ( .A(u0__abc_76628_new_n4957_), .B(u0__abc_76628_new_n4954_), .Y(u0__abc_76628_new_n4958_));
OR2X2 OR2X2_1237 ( .A(u0__abc_76628_new_n4959_), .B(u0__abc_76628_new_n4960_), .Y(u0__abc_76628_new_n4961_));
OR2X2 OR2X2_1238 ( .A(u0__abc_76628_new_n4963_), .B(u0__abc_76628_new_n4962_), .Y(u0__abc_76628_new_n4964_));
OR2X2 OR2X2_1239 ( .A(u0__abc_76628_new_n4964_), .B(u0__abc_76628_new_n4961_), .Y(u0__abc_76628_new_n4965_));
OR2X2 OR2X2_124 ( .A(u0__abc_76628_new_n1156_), .B(u0__abc_76628_new_n1149_), .Y(u0__0spec_req_cs_7_0__6_));
OR2X2 OR2X2_1240 ( .A(u0__abc_76628_new_n4966_), .B(u0__abc_76628_new_n4967_), .Y(u0__abc_76628_new_n4968_));
OR2X2 OR2X2_1241 ( .A(u0__abc_76628_new_n4969_), .B(u0__abc_76628_new_n4970_), .Y(u0__abc_76628_new_n4971_));
OR2X2 OR2X2_1242 ( .A(u0__abc_76628_new_n4968_), .B(u0__abc_76628_new_n4971_), .Y(u0__abc_76628_new_n4972_));
OR2X2 OR2X2_1243 ( .A(u0__abc_76628_new_n4972_), .B(u0__abc_76628_new_n4965_), .Y(u0__abc_76628_new_n4973_));
OR2X2 OR2X2_1244 ( .A(u0__abc_76628_new_n4973_), .B(u0__abc_76628_new_n4958_), .Y(u0__abc_76628_new_n4974_));
OR2X2 OR2X2_1245 ( .A(u0__abc_76628_new_n4974_), .B(u0__abc_76628_new_n4953_), .Y(rf_dout_11_));
OR2X2 OR2X2_1246 ( .A(u0__abc_76628_new_n4976_), .B(u0__abc_76628_new_n4977_), .Y(u0__abc_76628_new_n4978_));
OR2X2 OR2X2_1247 ( .A(u0__abc_76628_new_n4979_), .B(u0__abc_76628_new_n4980_), .Y(u0__abc_76628_new_n4981_));
OR2X2 OR2X2_1248 ( .A(u0__abc_76628_new_n4983_), .B(u0__abc_76628_new_n4982_), .Y(u0__abc_76628_new_n4984_));
OR2X2 OR2X2_1249 ( .A(u0__abc_76628_new_n4981_), .B(u0__abc_76628_new_n4984_), .Y(u0__abc_76628_new_n4985_));
OR2X2 OR2X2_125 ( .A(init_req), .B(1'h0), .Y(u0__abc_76628_new_n1160_));
OR2X2 OR2X2_1250 ( .A(u0__abc_76628_new_n4985_), .B(u0__abc_76628_new_n4978_), .Y(u0__abc_76628_new_n4986_));
OR2X2 OR2X2_1251 ( .A(u0__abc_76628_new_n4988_), .B(u0__abc_76628_new_n4989_), .Y(u0__abc_76628_new_n4990_));
OR2X2 OR2X2_1252 ( .A(u0__abc_76628_new_n4990_), .B(u0__abc_76628_new_n4987_), .Y(u0__abc_76628_new_n4991_));
OR2X2 OR2X2_1253 ( .A(u0__abc_76628_new_n4992_), .B(u0__abc_76628_new_n4993_), .Y(u0__abc_76628_new_n4994_));
OR2X2 OR2X2_1254 ( .A(u0__abc_76628_new_n4996_), .B(u0__abc_76628_new_n4995_), .Y(u0__abc_76628_new_n4997_));
OR2X2 OR2X2_1255 ( .A(u0__abc_76628_new_n4997_), .B(u0__abc_76628_new_n4994_), .Y(u0__abc_76628_new_n4998_));
OR2X2 OR2X2_1256 ( .A(u0__abc_76628_new_n4999_), .B(u0__abc_76628_new_n5000_), .Y(u0__abc_76628_new_n5001_));
OR2X2 OR2X2_1257 ( .A(u0__abc_76628_new_n5002_), .B(u0__abc_76628_new_n5003_), .Y(u0__abc_76628_new_n5004_));
OR2X2 OR2X2_1258 ( .A(u0__abc_76628_new_n5001_), .B(u0__abc_76628_new_n5004_), .Y(u0__abc_76628_new_n5005_));
OR2X2 OR2X2_1259 ( .A(u0__abc_76628_new_n5005_), .B(u0__abc_76628_new_n4998_), .Y(u0__abc_76628_new_n5006_));
OR2X2 OR2X2_126 ( .A(u0__abc_76628_new_n1100_), .B(1'h0), .Y(u0__abc_76628_new_n1161_));
OR2X2 OR2X2_1260 ( .A(u0__abc_76628_new_n5006_), .B(u0__abc_76628_new_n4991_), .Y(u0__abc_76628_new_n5007_));
OR2X2 OR2X2_1261 ( .A(u0__abc_76628_new_n5007_), .B(u0__abc_76628_new_n4986_), .Y(rf_dout_12_));
OR2X2 OR2X2_1262 ( .A(u0__abc_76628_new_n5009_), .B(u0__abc_76628_new_n5010_), .Y(u0__abc_76628_new_n5011_));
OR2X2 OR2X2_1263 ( .A(u0__abc_76628_new_n5012_), .B(u0__abc_76628_new_n5013_), .Y(u0__abc_76628_new_n5014_));
OR2X2 OR2X2_1264 ( .A(u0__abc_76628_new_n5015_), .B(u0__abc_76628_new_n5016_), .Y(u0__abc_76628_new_n5017_));
OR2X2 OR2X2_1265 ( .A(u0__abc_76628_new_n5014_), .B(u0__abc_76628_new_n5017_), .Y(u0__abc_76628_new_n5018_));
OR2X2 OR2X2_1266 ( .A(u0__abc_76628_new_n5018_), .B(u0__abc_76628_new_n5011_), .Y(u0__abc_76628_new_n5019_));
OR2X2 OR2X2_1267 ( .A(u0__abc_76628_new_n5021_), .B(u0__abc_76628_new_n5022_), .Y(u0__abc_76628_new_n5023_));
OR2X2 OR2X2_1268 ( .A(u0__abc_76628_new_n5023_), .B(u0__abc_76628_new_n5020_), .Y(u0__abc_76628_new_n5024_));
OR2X2 OR2X2_1269 ( .A(u0__abc_76628_new_n5025_), .B(u0__abc_76628_new_n5026_), .Y(u0__abc_76628_new_n5027_));
OR2X2 OR2X2_127 ( .A(u0__abc_76628_new_n1165_), .B(u0__abc_76628_new_n1158_), .Y(u0__0spec_req_cs_7_0__7_));
OR2X2 OR2X2_1270 ( .A(u0__abc_76628_new_n5028_), .B(u0__abc_76628_new_n5029_), .Y(u0__abc_76628_new_n5030_));
OR2X2 OR2X2_1271 ( .A(u0__abc_76628_new_n5030_), .B(u0__abc_76628_new_n5027_), .Y(u0__abc_76628_new_n5031_));
OR2X2 OR2X2_1272 ( .A(u0__abc_76628_new_n5032_), .B(u0__abc_76628_new_n5033_), .Y(u0__abc_76628_new_n5034_));
OR2X2 OR2X2_1273 ( .A(u0__abc_76628_new_n5035_), .B(u0__abc_76628_new_n5036_), .Y(u0__abc_76628_new_n5037_));
OR2X2 OR2X2_1274 ( .A(u0__abc_76628_new_n5037_), .B(u0__abc_76628_new_n5034_), .Y(u0__abc_76628_new_n5038_));
OR2X2 OR2X2_1275 ( .A(u0__abc_76628_new_n5031_), .B(u0__abc_76628_new_n5038_), .Y(u0__abc_76628_new_n5039_));
OR2X2 OR2X2_1276 ( .A(u0__abc_76628_new_n5039_), .B(u0__abc_76628_new_n5024_), .Y(u0__abc_76628_new_n5040_));
OR2X2 OR2X2_1277 ( .A(u0__abc_76628_new_n5040_), .B(u0__abc_76628_new_n5019_), .Y(rf_dout_13_));
OR2X2 OR2X2_1278 ( .A(u0__abc_76628_new_n5042_), .B(u0__abc_76628_new_n5043_), .Y(u0__abc_76628_new_n5044_));
OR2X2 OR2X2_1279 ( .A(u0__abc_76628_new_n5045_), .B(u0__abc_76628_new_n5046_), .Y(u0__abc_76628_new_n5047_));
OR2X2 OR2X2_128 ( .A(cs_le_d), .B(u0_rf_we), .Y(u0__abc_76628_new_n1167_));
OR2X2 OR2X2_1280 ( .A(u0__abc_76628_new_n5048_), .B(u0__abc_76628_new_n5049_), .Y(u0__abc_76628_new_n5050_));
OR2X2 OR2X2_1281 ( .A(u0__abc_76628_new_n5047_), .B(u0__abc_76628_new_n5050_), .Y(u0__abc_76628_new_n5051_));
OR2X2 OR2X2_1282 ( .A(u0__abc_76628_new_n5051_), .B(u0__abc_76628_new_n5044_), .Y(u0__abc_76628_new_n5052_));
OR2X2 OR2X2_1283 ( .A(u0__abc_76628_new_n5054_), .B(u0__abc_76628_new_n5055_), .Y(u0__abc_76628_new_n5056_));
OR2X2 OR2X2_1284 ( .A(u0__abc_76628_new_n5056_), .B(u0__abc_76628_new_n5053_), .Y(u0__abc_76628_new_n5057_));
OR2X2 OR2X2_1285 ( .A(u0__abc_76628_new_n5058_), .B(u0__abc_76628_new_n5059_), .Y(u0__abc_76628_new_n5060_));
OR2X2 OR2X2_1286 ( .A(u0__abc_76628_new_n5061_), .B(u0__abc_76628_new_n5062_), .Y(u0__abc_76628_new_n5063_));
OR2X2 OR2X2_1287 ( .A(u0__abc_76628_new_n5063_), .B(u0__abc_76628_new_n5060_), .Y(u0__abc_76628_new_n5064_));
OR2X2 OR2X2_1288 ( .A(u0__abc_76628_new_n5065_), .B(u0__abc_76628_new_n5066_), .Y(u0__abc_76628_new_n5067_));
OR2X2 OR2X2_1289 ( .A(u0__abc_76628_new_n5068_), .B(u0__abc_76628_new_n5069_), .Y(u0__abc_76628_new_n5070_));
OR2X2 OR2X2_129 ( .A(u0__abc_76628_new_n1177__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n1178_));
OR2X2 OR2X2_1290 ( .A(u0__abc_76628_new_n5070_), .B(u0__abc_76628_new_n5067_), .Y(u0__abc_76628_new_n5071_));
OR2X2 OR2X2_1291 ( .A(u0__abc_76628_new_n5064_), .B(u0__abc_76628_new_n5071_), .Y(u0__abc_76628_new_n5072_));
OR2X2 OR2X2_1292 ( .A(u0__abc_76628_new_n5072_), .B(u0__abc_76628_new_n5057_), .Y(u0__abc_76628_new_n5073_));
OR2X2 OR2X2_1293 ( .A(u0__abc_76628_new_n5073_), .B(u0__abc_76628_new_n5052_), .Y(rf_dout_14_));
OR2X2 OR2X2_1294 ( .A(u0__abc_76628_new_n5077_), .B(u0__abc_76628_new_n5076_), .Y(u0__abc_76628_new_n5078_));
OR2X2 OR2X2_1295 ( .A(u0__abc_76628_new_n5078_), .B(u0__abc_76628_new_n5075_), .Y(u0__abc_76628_new_n5079_));
OR2X2 OR2X2_1296 ( .A(u0__abc_76628_new_n5080_), .B(u0__abc_76628_new_n5081_), .Y(u0__abc_76628_new_n5082_));
OR2X2 OR2X2_1297 ( .A(u0__abc_76628_new_n5083_), .B(u0__abc_76628_new_n5084_), .Y(u0__abc_76628_new_n5085_));
OR2X2 OR2X2_1298 ( .A(u0__abc_76628_new_n5082_), .B(u0__abc_76628_new_n5085_), .Y(u0__abc_76628_new_n5086_));
OR2X2 OR2X2_1299 ( .A(u0__abc_76628_new_n5086_), .B(u0__abc_76628_new_n5079_), .Y(u0__abc_76628_new_n5087_));
OR2X2 OR2X2_13 ( .A(_abc_85006_new_n256_), .B(_abc_85006_new_n237_), .Y(_abc_85006_new_n257_));
OR2X2 OR2X2_130 ( .A(spec_req_cs_6_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1180_));
OR2X2 OR2X2_1300 ( .A(u0__abc_76628_new_n5090_), .B(u0__abc_76628_new_n5091_), .Y(u0__abc_76628_new_n5092_));
OR2X2 OR2X2_1301 ( .A(u0__abc_76628_new_n5092_), .B(u0__abc_76628_new_n5089_), .Y(u0__abc_76628_new_n5093_));
OR2X2 OR2X2_1302 ( .A(u0__abc_76628_new_n5093_), .B(u0__abc_76628_new_n5088_), .Y(u0__abc_76628_new_n5094_));
OR2X2 OR2X2_1303 ( .A(u0__abc_76628_new_n5096_), .B(u0__abc_76628_new_n5097_), .Y(u0__abc_76628_new_n5098_));
OR2X2 OR2X2_1304 ( .A(u0__abc_76628_new_n5098_), .B(u0__abc_76628_new_n5095_), .Y(u0__abc_76628_new_n5099_));
OR2X2 OR2X2_1305 ( .A(u0__abc_76628_new_n5101_), .B(u0__abc_76628_new_n5102_), .Y(u0__abc_76628_new_n5103_));
OR2X2 OR2X2_1306 ( .A(u0__abc_76628_new_n5103_), .B(u0__abc_76628_new_n5100_), .Y(u0__abc_76628_new_n5104_));
OR2X2 OR2X2_1307 ( .A(u0__abc_76628_new_n5099_), .B(u0__abc_76628_new_n5104_), .Y(u0__abc_76628_new_n5105_));
OR2X2 OR2X2_1308 ( .A(u0__abc_76628_new_n5105_), .B(u0__abc_76628_new_n5094_), .Y(u0__abc_76628_new_n5106_));
OR2X2 OR2X2_1309 ( .A(u0__abc_76628_new_n5106_), .B(u0__abc_76628_new_n5087_), .Y(rf_dout_15_));
OR2X2 OR2X2_131 ( .A(u0__abc_76628_new_n1182_), .B(u0__abc_76628_new_n1176_), .Y(u0__abc_76628_new_n1183_));
OR2X2 OR2X2_1310 ( .A(u0__abc_76628_new_n5108_), .B(u0__abc_76628_new_n5109_), .Y(u0__abc_76628_new_n5110_));
OR2X2 OR2X2_1311 ( .A(u0__abc_76628_new_n5112_), .B(u0__abc_76628_new_n5111_), .Y(u0__abc_76628_new_n5113_));
OR2X2 OR2X2_1312 ( .A(u0__abc_76628_new_n5114_), .B(u0__abc_76628_new_n5115_), .Y(u0__abc_76628_new_n5116_));
OR2X2 OR2X2_1313 ( .A(u0__abc_76628_new_n5113_), .B(u0__abc_76628_new_n5116_), .Y(u0__abc_76628_new_n5117_));
OR2X2 OR2X2_1314 ( .A(u0__abc_76628_new_n5117_), .B(u0__abc_76628_new_n5110_), .Y(u0__abc_76628_new_n5118_));
OR2X2 OR2X2_1315 ( .A(u0__abc_76628_new_n5120_), .B(u0__abc_76628_new_n5121_), .Y(u0__abc_76628_new_n5122_));
OR2X2 OR2X2_1316 ( .A(u0__abc_76628_new_n5122_), .B(u0__abc_76628_new_n5119_), .Y(u0__abc_76628_new_n5123_));
OR2X2 OR2X2_1317 ( .A(u0__abc_76628_new_n5125_), .B(u0__abc_76628_new_n5124_), .Y(u0__abc_76628_new_n5126_));
OR2X2 OR2X2_1318 ( .A(u0__abc_76628_new_n5127_), .B(u0__abc_76628_new_n5128_), .Y(u0__abc_76628_new_n5129_));
OR2X2 OR2X2_1319 ( .A(u0__abc_76628_new_n5129_), .B(u0__abc_76628_new_n5126_), .Y(u0__abc_76628_new_n5130_));
OR2X2 OR2X2_132 ( .A(u0__abc_76628_new_n1184_), .B(u0__abc_76628_new_n1185_), .Y(u0__abc_76628_new_n1186_));
OR2X2 OR2X2_1320 ( .A(u0__abc_76628_new_n5131_), .B(u0__abc_76628_new_n5132_), .Y(u0__abc_76628_new_n5133_));
OR2X2 OR2X2_1321 ( .A(u0__abc_76628_new_n5135_), .B(u0__abc_76628_new_n5134_), .Y(u0__abc_76628_new_n5136_));
OR2X2 OR2X2_1322 ( .A(u0__abc_76628_new_n5133_), .B(u0__abc_76628_new_n5136_), .Y(u0__abc_76628_new_n5137_));
OR2X2 OR2X2_1323 ( .A(u0__abc_76628_new_n5137_), .B(u0__abc_76628_new_n5130_), .Y(u0__abc_76628_new_n5138_));
OR2X2 OR2X2_1324 ( .A(u0__abc_76628_new_n5138_), .B(u0__abc_76628_new_n5123_), .Y(u0__abc_76628_new_n5139_));
OR2X2 OR2X2_1325 ( .A(u0__abc_76628_new_n5139_), .B(u0__abc_76628_new_n5118_), .Y(rf_dout_16_));
OR2X2 OR2X2_1326 ( .A(u0__abc_76628_new_n5141_), .B(u0__abc_76628_new_n5142_), .Y(u0__abc_76628_new_n5143_));
OR2X2 OR2X2_1327 ( .A(u0__abc_76628_new_n5144_), .B(u0__abc_76628_new_n5145_), .Y(u0__abc_76628_new_n5146_));
OR2X2 OR2X2_1328 ( .A(u0__abc_76628_new_n5148_), .B(u0__abc_76628_new_n5147_), .Y(u0__abc_76628_new_n5149_));
OR2X2 OR2X2_1329 ( .A(u0__abc_76628_new_n5146_), .B(u0__abc_76628_new_n5149_), .Y(u0__abc_76628_new_n5150_));
OR2X2 OR2X2_133 ( .A(u0__abc_76628_new_n1187_), .B(u0__abc_76628_new_n1188_), .Y(u0__abc_76628_new_n1189_));
OR2X2 OR2X2_1330 ( .A(u0__abc_76628_new_n5150_), .B(u0__abc_76628_new_n5143_), .Y(u0__abc_76628_new_n5151_));
OR2X2 OR2X2_1331 ( .A(u0__abc_76628_new_n5154_), .B(u0__abc_76628_new_n5153_), .Y(u0__abc_76628_new_n5155_));
OR2X2 OR2X2_1332 ( .A(u0__abc_76628_new_n5155_), .B(u0__abc_76628_new_n5152_), .Y(u0__abc_76628_new_n5156_));
OR2X2 OR2X2_1333 ( .A(u0__abc_76628_new_n5157_), .B(u0__abc_76628_new_n5158_), .Y(u0__abc_76628_new_n5159_));
OR2X2 OR2X2_1334 ( .A(u0__abc_76628_new_n5161_), .B(u0__abc_76628_new_n5160_), .Y(u0__abc_76628_new_n5162_));
OR2X2 OR2X2_1335 ( .A(u0__abc_76628_new_n5162_), .B(u0__abc_76628_new_n5159_), .Y(u0__abc_76628_new_n5163_));
OR2X2 OR2X2_1336 ( .A(u0__abc_76628_new_n5164_), .B(u0__abc_76628_new_n5165_), .Y(u0__abc_76628_new_n5166_));
OR2X2 OR2X2_1337 ( .A(u0__abc_76628_new_n5167_), .B(u0__abc_76628_new_n5168_), .Y(u0__abc_76628_new_n5169_));
OR2X2 OR2X2_1338 ( .A(u0__abc_76628_new_n5166_), .B(u0__abc_76628_new_n5169_), .Y(u0__abc_76628_new_n5170_));
OR2X2 OR2X2_1339 ( .A(u0__abc_76628_new_n5170_), .B(u0__abc_76628_new_n5163_), .Y(u0__abc_76628_new_n5171_));
OR2X2 OR2X2_134 ( .A(u0__abc_76628_new_n1190_), .B(u0__abc_76628_new_n1191_), .Y(u0__abc_76628_new_n1192_));
OR2X2 OR2X2_1340 ( .A(u0__abc_76628_new_n5171_), .B(u0__abc_76628_new_n5156_), .Y(u0__abc_76628_new_n5172_));
OR2X2 OR2X2_1341 ( .A(u0__abc_76628_new_n5172_), .B(u0__abc_76628_new_n5151_), .Y(rf_dout_17_));
OR2X2 OR2X2_1342 ( .A(u0__abc_76628_new_n5176_), .B(u0__abc_76628_new_n5175_), .Y(u0__abc_76628_new_n5177_));
OR2X2 OR2X2_1343 ( .A(u0__abc_76628_new_n5177_), .B(u0__abc_76628_new_n5174_), .Y(u0__abc_76628_new_n5178_));
OR2X2 OR2X2_1344 ( .A(u0__abc_76628_new_n5179_), .B(u0__abc_76628_new_n5180_), .Y(u0__abc_76628_new_n5181_));
OR2X2 OR2X2_1345 ( .A(u0__abc_76628_new_n5182_), .B(u0__abc_76628_new_n5183_), .Y(u0__abc_76628_new_n5184_));
OR2X2 OR2X2_1346 ( .A(u0__abc_76628_new_n5181_), .B(u0__abc_76628_new_n5184_), .Y(u0__abc_76628_new_n5185_));
OR2X2 OR2X2_1347 ( .A(u0__abc_76628_new_n5185_), .B(u0__abc_76628_new_n5178_), .Y(u0__abc_76628_new_n5186_));
OR2X2 OR2X2_1348 ( .A(u0__abc_76628_new_n5189_), .B(u0__abc_76628_new_n5190_), .Y(u0__abc_76628_new_n5191_));
OR2X2 OR2X2_1349 ( .A(u0__abc_76628_new_n5191_), .B(u0__abc_76628_new_n5188_), .Y(u0__abc_76628_new_n5192_));
OR2X2 OR2X2_135 ( .A(u0__abc_76628_new_n1194_), .B(spec_req_cs_0_bF_buf3_), .Y(u0__abc_76628_new_n1195_));
OR2X2 OR2X2_1350 ( .A(u0__abc_76628_new_n5192_), .B(u0__abc_76628_new_n5187_), .Y(u0__abc_76628_new_n5193_));
OR2X2 OR2X2_1351 ( .A(u0__abc_76628_new_n5195_), .B(u0__abc_76628_new_n5196_), .Y(u0__abc_76628_new_n5197_));
OR2X2 OR2X2_1352 ( .A(u0__abc_76628_new_n5197_), .B(u0__abc_76628_new_n5194_), .Y(u0__abc_76628_new_n5198_));
OR2X2 OR2X2_1353 ( .A(u0__abc_76628_new_n5200_), .B(u0__abc_76628_new_n5201_), .Y(u0__abc_76628_new_n5202_));
OR2X2 OR2X2_1354 ( .A(u0__abc_76628_new_n5202_), .B(u0__abc_76628_new_n5199_), .Y(u0__abc_76628_new_n5203_));
OR2X2 OR2X2_1355 ( .A(u0__abc_76628_new_n5198_), .B(u0__abc_76628_new_n5203_), .Y(u0__abc_76628_new_n5204_));
OR2X2 OR2X2_1356 ( .A(u0__abc_76628_new_n5204_), .B(u0__abc_76628_new_n5193_), .Y(u0__abc_76628_new_n5205_));
OR2X2 OR2X2_1357 ( .A(u0__abc_76628_new_n5205_), .B(u0__abc_76628_new_n5186_), .Y(rf_dout_18_));
OR2X2 OR2X2_1358 ( .A(u0__abc_76628_new_n5208_), .B(u0__abc_76628_new_n5209_), .Y(u0__abc_76628_new_n5210_));
OR2X2 OR2X2_1359 ( .A(u0__abc_76628_new_n5210_), .B(u0__abc_76628_new_n5207_), .Y(u0__abc_76628_new_n5211_));
OR2X2 OR2X2_136 ( .A(u0__abc_76628_new_n1193_), .B(u0__abc_76628_new_n1195_), .Y(u0__abc_76628_new_n1196_));
OR2X2 OR2X2_1360 ( .A(u0__abc_76628_new_n5212_), .B(u0__abc_76628_new_n5213_), .Y(u0__abc_76628_new_n5214_));
OR2X2 OR2X2_1361 ( .A(u0__abc_76628_new_n5211_), .B(u0__abc_76628_new_n5214_), .Y(u0__abc_76628_new_n5215_));
OR2X2 OR2X2_1362 ( .A(u0__abc_76628_new_n5217_), .B(u0__abc_76628_new_n5218_), .Y(u0__abc_76628_new_n5219_));
OR2X2 OR2X2_1363 ( .A(u0__abc_76628_new_n5219_), .B(u0__abc_76628_new_n5216_), .Y(u0__abc_76628_new_n5220_));
OR2X2 OR2X2_1364 ( .A(u0__abc_76628_new_n5223_), .B(u0__abc_76628_new_n5222_), .Y(u0__abc_76628_new_n5224_));
OR2X2 OR2X2_1365 ( .A(u0__abc_76628_new_n5224_), .B(u0__abc_76628_new_n5221_), .Y(u0__abc_76628_new_n5225_));
OR2X2 OR2X2_1366 ( .A(u0__abc_76628_new_n5220_), .B(u0__abc_76628_new_n5225_), .Y(u0__abc_76628_new_n5226_));
OR2X2 OR2X2_1367 ( .A(u0__abc_76628_new_n5229_), .B(u0__abc_76628_new_n5228_), .Y(u0__abc_76628_new_n5230_));
OR2X2 OR2X2_1368 ( .A(u0__abc_76628_new_n5230_), .B(u0__abc_76628_new_n5227_), .Y(u0__abc_76628_new_n5231_));
OR2X2 OR2X2_1369 ( .A(u0__abc_76628_new_n5233_), .B(u0__abc_76628_new_n5234_), .Y(u0__abc_76628_new_n5235_));
OR2X2 OR2X2_137 ( .A(u0__abc_76628_new_n1197__bF_buf5), .B(u0_tms0_0_), .Y(u0__abc_76628_new_n1198_));
OR2X2 OR2X2_1370 ( .A(u0__abc_76628_new_n5235_), .B(u0__abc_76628_new_n5232_), .Y(u0__abc_76628_new_n5236_));
OR2X2 OR2X2_1371 ( .A(u0__abc_76628_new_n5236_), .B(u0__abc_76628_new_n5231_), .Y(u0__abc_76628_new_n5237_));
OR2X2 OR2X2_1372 ( .A(u0__abc_76628_new_n5226_), .B(u0__abc_76628_new_n5237_), .Y(u0__abc_76628_new_n5238_));
OR2X2 OR2X2_1373 ( .A(u0__abc_76628_new_n5238_), .B(u0__abc_76628_new_n5215_), .Y(rf_dout_19_));
OR2X2 OR2X2_1374 ( .A(u0__abc_76628_new_n5242_), .B(u0__abc_76628_new_n5241_), .Y(u0__abc_76628_new_n5243_));
OR2X2 OR2X2_1375 ( .A(u0__abc_76628_new_n5243_), .B(u0__abc_76628_new_n5240_), .Y(u0__abc_76628_new_n5244_));
OR2X2 OR2X2_1376 ( .A(u0__abc_76628_new_n5245_), .B(u0__abc_76628_new_n5246_), .Y(u0__abc_76628_new_n5247_));
OR2X2 OR2X2_1377 ( .A(u0__abc_76628_new_n5248_), .B(u0__abc_76628_new_n5249_), .Y(u0__abc_76628_new_n5250_));
OR2X2 OR2X2_1378 ( .A(u0__abc_76628_new_n5247_), .B(u0__abc_76628_new_n5250_), .Y(u0__abc_76628_new_n5251_));
OR2X2 OR2X2_1379 ( .A(u0__abc_76628_new_n5251_), .B(u0__abc_76628_new_n5244_), .Y(u0__abc_76628_new_n5252_));
OR2X2 OR2X2_138 ( .A(u0__abc_76628_new_n1200_), .B(u0__abc_76628_new_n1171_), .Y(u0__0sp_tms_31_0__0_));
OR2X2 OR2X2_1380 ( .A(u0__abc_76628_new_n5255_), .B(u0__abc_76628_new_n5256_), .Y(u0__abc_76628_new_n5257_));
OR2X2 OR2X2_1381 ( .A(u0__abc_76628_new_n5257_), .B(u0__abc_76628_new_n5254_), .Y(u0__abc_76628_new_n5258_));
OR2X2 OR2X2_1382 ( .A(u0__abc_76628_new_n5258_), .B(u0__abc_76628_new_n5253_), .Y(u0__abc_76628_new_n5259_));
OR2X2 OR2X2_1383 ( .A(u0__abc_76628_new_n5261_), .B(u0__abc_76628_new_n5262_), .Y(u0__abc_76628_new_n5263_));
OR2X2 OR2X2_1384 ( .A(u0__abc_76628_new_n5263_), .B(u0__abc_76628_new_n5260_), .Y(u0__abc_76628_new_n5264_));
OR2X2 OR2X2_1385 ( .A(u0__abc_76628_new_n5266_), .B(u0__abc_76628_new_n5267_), .Y(u0__abc_76628_new_n5268_));
OR2X2 OR2X2_1386 ( .A(u0__abc_76628_new_n5268_), .B(u0__abc_76628_new_n5265_), .Y(u0__abc_76628_new_n5269_));
OR2X2 OR2X2_1387 ( .A(u0__abc_76628_new_n5264_), .B(u0__abc_76628_new_n5269_), .Y(u0__abc_76628_new_n5270_));
OR2X2 OR2X2_1388 ( .A(u0__abc_76628_new_n5270_), .B(u0__abc_76628_new_n5259_), .Y(u0__abc_76628_new_n5271_));
OR2X2 OR2X2_1389 ( .A(u0__abc_76628_new_n5271_), .B(u0__abc_76628_new_n5252_), .Y(rf_dout_20_));
OR2X2 OR2X2_139 ( .A(u0__abc_76628_new_n1177__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n1204_));
OR2X2 OR2X2_1390 ( .A(u0__abc_76628_new_n5273_), .B(u0__abc_76628_new_n5274_), .Y(u0__abc_76628_new_n5275_));
OR2X2 OR2X2_1391 ( .A(u0__abc_76628_new_n5276_), .B(u0__abc_76628_new_n5277_), .Y(u0__abc_76628_new_n5278_));
OR2X2 OR2X2_1392 ( .A(u0__abc_76628_new_n5279_), .B(u0__abc_76628_new_n5280_), .Y(u0__abc_76628_new_n5281_));
OR2X2 OR2X2_1393 ( .A(u0__abc_76628_new_n5278_), .B(u0__abc_76628_new_n5281_), .Y(u0__abc_76628_new_n5282_));
OR2X2 OR2X2_1394 ( .A(u0__abc_76628_new_n5282_), .B(u0__abc_76628_new_n5275_), .Y(u0__abc_76628_new_n5283_));
OR2X2 OR2X2_1395 ( .A(u0__abc_76628_new_n5285_), .B(u0__abc_76628_new_n5286_), .Y(u0__abc_76628_new_n5287_));
OR2X2 OR2X2_1396 ( .A(u0__abc_76628_new_n5287_), .B(u0__abc_76628_new_n5284_), .Y(u0__abc_76628_new_n5288_));
OR2X2 OR2X2_1397 ( .A(u0__abc_76628_new_n5289_), .B(u0__abc_76628_new_n5290_), .Y(u0__abc_76628_new_n5291_));
OR2X2 OR2X2_1398 ( .A(u0__abc_76628_new_n5292_), .B(u0__abc_76628_new_n5293_), .Y(u0__abc_76628_new_n5294_));
OR2X2 OR2X2_1399 ( .A(u0__abc_76628_new_n5294_), .B(u0__abc_76628_new_n5291_), .Y(u0__abc_76628_new_n5295_));
OR2X2 OR2X2_14 ( .A(_abc_85006_new_n245_), .B(cs_need_rfr_2_), .Y(_abc_85006_new_n258_));
OR2X2 OR2X2_140 ( .A(spec_req_cs_6_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1205_));
OR2X2 OR2X2_1400 ( .A(u0__abc_76628_new_n5296_), .B(u0__abc_76628_new_n5297_), .Y(u0__abc_76628_new_n5298_));
OR2X2 OR2X2_1401 ( .A(u0__abc_76628_new_n5300_), .B(u0__abc_76628_new_n5299_), .Y(u0__abc_76628_new_n5301_));
OR2X2 OR2X2_1402 ( .A(u0__abc_76628_new_n5301_), .B(u0__abc_76628_new_n5298_), .Y(u0__abc_76628_new_n5302_));
OR2X2 OR2X2_1403 ( .A(u0__abc_76628_new_n5295_), .B(u0__abc_76628_new_n5302_), .Y(u0__abc_76628_new_n5303_));
OR2X2 OR2X2_1404 ( .A(u0__abc_76628_new_n5303_), .B(u0__abc_76628_new_n5288_), .Y(u0__abc_76628_new_n5304_));
OR2X2 OR2X2_1405 ( .A(u0__abc_76628_new_n5304_), .B(u0__abc_76628_new_n5283_), .Y(rf_dout_21_));
OR2X2 OR2X2_1406 ( .A(u0__abc_76628_new_n5306_), .B(u0__abc_76628_new_n5307_), .Y(u0__abc_76628_new_n5308_));
OR2X2 OR2X2_1407 ( .A(u0__abc_76628_new_n5309_), .B(u0__abc_76628_new_n5310_), .Y(u0__abc_76628_new_n5311_));
OR2X2 OR2X2_1408 ( .A(u0__abc_76628_new_n5313_), .B(u0__abc_76628_new_n5312_), .Y(u0__abc_76628_new_n5314_));
OR2X2 OR2X2_1409 ( .A(u0__abc_76628_new_n5311_), .B(u0__abc_76628_new_n5314_), .Y(u0__abc_76628_new_n5315_));
OR2X2 OR2X2_141 ( .A(u0__abc_76628_new_n1207_), .B(u0__abc_76628_new_n1203_), .Y(u0__abc_76628_new_n1208_));
OR2X2 OR2X2_1410 ( .A(u0__abc_76628_new_n5315_), .B(u0__abc_76628_new_n5308_), .Y(u0__abc_76628_new_n5316_));
OR2X2 OR2X2_1411 ( .A(u0__abc_76628_new_n5318_), .B(u0__abc_76628_new_n5319_), .Y(u0__abc_76628_new_n5320_));
OR2X2 OR2X2_1412 ( .A(u0__abc_76628_new_n5320_), .B(u0__abc_76628_new_n5317_), .Y(u0__abc_76628_new_n5321_));
OR2X2 OR2X2_1413 ( .A(u0__abc_76628_new_n5322_), .B(u0__abc_76628_new_n5323_), .Y(u0__abc_76628_new_n5324_));
OR2X2 OR2X2_1414 ( .A(u0__abc_76628_new_n5326_), .B(u0__abc_76628_new_n5325_), .Y(u0__abc_76628_new_n5327_));
OR2X2 OR2X2_1415 ( .A(u0__abc_76628_new_n5327_), .B(u0__abc_76628_new_n5324_), .Y(u0__abc_76628_new_n5328_));
OR2X2 OR2X2_1416 ( .A(u0__abc_76628_new_n5329_), .B(u0__abc_76628_new_n5330_), .Y(u0__abc_76628_new_n5331_));
OR2X2 OR2X2_1417 ( .A(u0__abc_76628_new_n5332_), .B(u0__abc_76628_new_n5333_), .Y(u0__abc_76628_new_n5334_));
OR2X2 OR2X2_1418 ( .A(u0__abc_76628_new_n5331_), .B(u0__abc_76628_new_n5334_), .Y(u0__abc_76628_new_n5335_));
OR2X2 OR2X2_1419 ( .A(u0__abc_76628_new_n5335_), .B(u0__abc_76628_new_n5328_), .Y(u0__abc_76628_new_n5336_));
OR2X2 OR2X2_142 ( .A(u0__abc_76628_new_n1209_), .B(u0__abc_76628_new_n1210_), .Y(u0__abc_76628_new_n1211_));
OR2X2 OR2X2_1420 ( .A(u0__abc_76628_new_n5336_), .B(u0__abc_76628_new_n5321_), .Y(u0__abc_76628_new_n5337_));
OR2X2 OR2X2_1421 ( .A(u0__abc_76628_new_n5337_), .B(u0__abc_76628_new_n5316_), .Y(rf_dout_22_));
OR2X2 OR2X2_1422 ( .A(u0__abc_76628_new_n5339_), .B(u0__abc_76628_new_n5340_), .Y(u0__abc_76628_new_n5341_));
OR2X2 OR2X2_1423 ( .A(u0__abc_76628_new_n5343_), .B(u0__abc_76628_new_n5342_), .Y(u0__abc_76628_new_n5344_));
OR2X2 OR2X2_1424 ( .A(u0__abc_76628_new_n5345_), .B(u0__abc_76628_new_n5346_), .Y(u0__abc_76628_new_n5347_));
OR2X2 OR2X2_1425 ( .A(u0__abc_76628_new_n5344_), .B(u0__abc_76628_new_n5347_), .Y(u0__abc_76628_new_n5348_));
OR2X2 OR2X2_1426 ( .A(u0__abc_76628_new_n5348_), .B(u0__abc_76628_new_n5341_), .Y(u0__abc_76628_new_n5349_));
OR2X2 OR2X2_1427 ( .A(u0__abc_76628_new_n5351_), .B(u0__abc_76628_new_n5352_), .Y(u0__abc_76628_new_n5353_));
OR2X2 OR2X2_1428 ( .A(u0__abc_76628_new_n5353_), .B(u0__abc_76628_new_n5350_), .Y(u0__abc_76628_new_n5354_));
OR2X2 OR2X2_1429 ( .A(u0__abc_76628_new_n5356_), .B(u0__abc_76628_new_n5355_), .Y(u0__abc_76628_new_n5357_));
OR2X2 OR2X2_143 ( .A(u0__abc_76628_new_n1212_), .B(u0__abc_76628_new_n1213_), .Y(u0__abc_76628_new_n1214_));
OR2X2 OR2X2_1430 ( .A(u0__abc_76628_new_n5358_), .B(u0__abc_76628_new_n5359_), .Y(u0__abc_76628_new_n5360_));
OR2X2 OR2X2_1431 ( .A(u0__abc_76628_new_n5360_), .B(u0__abc_76628_new_n5357_), .Y(u0__abc_76628_new_n5361_));
OR2X2 OR2X2_1432 ( .A(u0__abc_76628_new_n5362_), .B(u0__abc_76628_new_n5363_), .Y(u0__abc_76628_new_n5364_));
OR2X2 OR2X2_1433 ( .A(u0__abc_76628_new_n5366_), .B(u0__abc_76628_new_n5365_), .Y(u0__abc_76628_new_n5367_));
OR2X2 OR2X2_1434 ( .A(u0__abc_76628_new_n5364_), .B(u0__abc_76628_new_n5367_), .Y(u0__abc_76628_new_n5368_));
OR2X2 OR2X2_1435 ( .A(u0__abc_76628_new_n5368_), .B(u0__abc_76628_new_n5361_), .Y(u0__abc_76628_new_n5369_));
OR2X2 OR2X2_1436 ( .A(u0__abc_76628_new_n5369_), .B(u0__abc_76628_new_n5354_), .Y(u0__abc_76628_new_n5370_));
OR2X2 OR2X2_1437 ( .A(u0__abc_76628_new_n5370_), .B(u0__abc_76628_new_n5349_), .Y(rf_dout_23_));
OR2X2 OR2X2_1438 ( .A(u0__abc_76628_new_n5372_), .B(u0__abc_76628_new_n5373_), .Y(u0__abc_76628_new_n5374_));
OR2X2 OR2X2_1439 ( .A(u0__abc_76628_new_n5376_), .B(u0__abc_76628_new_n5375_), .Y(u0__abc_76628_new_n5377_));
OR2X2 OR2X2_144 ( .A(u0__abc_76628_new_n1215_), .B(u0__abc_76628_new_n1216_), .Y(u0__abc_76628_new_n1217_));
OR2X2 OR2X2_1440 ( .A(u0__abc_76628_new_n5379_), .B(u0__abc_76628_new_n5378_), .Y(u0__abc_76628_new_n5380_));
OR2X2 OR2X2_1441 ( .A(u0__abc_76628_new_n5377_), .B(u0__abc_76628_new_n5380_), .Y(u0__abc_76628_new_n5381_));
OR2X2 OR2X2_1442 ( .A(u0__abc_76628_new_n5381_), .B(u0__abc_76628_new_n5374_), .Y(u0__abc_76628_new_n5382_));
OR2X2 OR2X2_1443 ( .A(u0__abc_76628_new_n5383_), .B(u0__abc_76628_new_n5384_), .Y(u0__abc_76628_new_n5385_));
OR2X2 OR2X2_1444 ( .A(u0__abc_76628_new_n5386_), .B(u0__abc_76628_new_n5387_), .Y(u0__abc_76628_new_n5388_));
OR2X2 OR2X2_1445 ( .A(u0__abc_76628_new_n5385_), .B(u0__abc_76628_new_n5388_), .Y(u0__abc_76628_new_n5389_));
OR2X2 OR2X2_1446 ( .A(u0__abc_76628_new_n5390_), .B(u0__abc_76628_new_n5391_), .Y(u0__abc_76628_new_n5392_));
OR2X2 OR2X2_1447 ( .A(u0__abc_76628_new_n5393_), .B(u0__abc_76628_new_n5394_), .Y(u0__abc_76628_new_n5395_));
OR2X2 OR2X2_1448 ( .A(u0__abc_76628_new_n5395_), .B(u0__abc_76628_new_n5392_), .Y(u0__abc_76628_new_n5396_));
OR2X2 OR2X2_1449 ( .A(u0__abc_76628_new_n5389_), .B(u0__abc_76628_new_n5396_), .Y(u0__abc_76628_new_n5397_));
OR2X2 OR2X2_145 ( .A(u0__abc_76628_new_n1219_), .B(spec_req_cs_0_bF_buf1_), .Y(u0__abc_76628_new_n1220_));
OR2X2 OR2X2_1450 ( .A(u0__abc_76628_new_n5400_), .B(u0__abc_76628_new_n5401_), .Y(u0__abc_76628_new_n5402_));
OR2X2 OR2X2_1451 ( .A(u0__abc_76628_new_n5402_), .B(u0__abc_76628_new_n5399_), .Y(u0__abc_76628_new_n5403_));
OR2X2 OR2X2_1452 ( .A(u0__abc_76628_new_n5403_), .B(u0__abc_76628_new_n5398_), .Y(u0__abc_76628_new_n5404_));
OR2X2 OR2X2_1453 ( .A(u0__abc_76628_new_n5397_), .B(u0__abc_76628_new_n5404_), .Y(u0__abc_76628_new_n5405_));
OR2X2 OR2X2_1454 ( .A(u0__abc_76628_new_n5405_), .B(u0__abc_76628_new_n5382_), .Y(rf_dout_24_));
OR2X2 OR2X2_1455 ( .A(u0__abc_76628_new_n5408_), .B(u0__abc_76628_new_n5407_), .Y(u0__abc_76628_new_n5409_));
OR2X2 OR2X2_1456 ( .A(u0__abc_76628_new_n5410_), .B(u0__abc_76628_new_n5411_), .Y(u0__abc_76628_new_n5412_));
OR2X2 OR2X2_1457 ( .A(u0__abc_76628_new_n5413_), .B(u0__abc_76628_new_n5414_), .Y(u0__abc_76628_new_n5415_));
OR2X2 OR2X2_1458 ( .A(u0__abc_76628_new_n5412_), .B(u0__abc_76628_new_n5415_), .Y(u0__abc_76628_new_n5416_));
OR2X2 OR2X2_1459 ( .A(u0__abc_76628_new_n5416_), .B(u0__abc_76628_new_n5409_), .Y(u0__abc_76628_new_n5417_));
OR2X2 OR2X2_146 ( .A(u0__abc_76628_new_n1218_), .B(u0__abc_76628_new_n1220_), .Y(u0__abc_76628_new_n1221_));
OR2X2 OR2X2_1460 ( .A(u0__abc_76628_new_n5419_), .B(u0__abc_76628_new_n5418_), .Y(u0__abc_76628_new_n5420_));
OR2X2 OR2X2_1461 ( .A(u0__abc_76628_new_n5422_), .B(u0__abc_76628_new_n5421_), .Y(u0__abc_76628_new_n5423_));
OR2X2 OR2X2_1462 ( .A(u0__abc_76628_new_n5420_), .B(u0__abc_76628_new_n5423_), .Y(u0__abc_76628_new_n5424_));
OR2X2 OR2X2_1463 ( .A(u0__abc_76628_new_n5425_), .B(u0__abc_76628_new_n5426_), .Y(u0__abc_76628_new_n5427_));
OR2X2 OR2X2_1464 ( .A(u0__abc_76628_new_n5428_), .B(u0__abc_76628_new_n5429_), .Y(u0__abc_76628_new_n5430_));
OR2X2 OR2X2_1465 ( .A(u0__abc_76628_new_n5427_), .B(u0__abc_76628_new_n5430_), .Y(u0__abc_76628_new_n5431_));
OR2X2 OR2X2_1466 ( .A(u0__abc_76628_new_n5424_), .B(u0__abc_76628_new_n5431_), .Y(u0__abc_76628_new_n5432_));
OR2X2 OR2X2_1467 ( .A(u0__abc_76628_new_n5435_), .B(u0__abc_76628_new_n5436_), .Y(u0__abc_76628_new_n5437_));
OR2X2 OR2X2_1468 ( .A(u0__abc_76628_new_n5437_), .B(u0__abc_76628_new_n5434_), .Y(u0__abc_76628_new_n5438_));
OR2X2 OR2X2_1469 ( .A(u0__abc_76628_new_n5438_), .B(u0__abc_76628_new_n5433_), .Y(u0__abc_76628_new_n5439_));
OR2X2 OR2X2_147 ( .A(u0__abc_76628_new_n1197__bF_buf4), .B(u0_tms0_1_), .Y(u0__abc_76628_new_n1222_));
OR2X2 OR2X2_1470 ( .A(u0__abc_76628_new_n5432_), .B(u0__abc_76628_new_n5439_), .Y(u0__abc_76628_new_n5440_));
OR2X2 OR2X2_1471 ( .A(u0__abc_76628_new_n5440_), .B(u0__abc_76628_new_n5417_), .Y(rf_dout_25_));
OR2X2 OR2X2_1472 ( .A(u0__abc_76628_new_n5444_), .B(u0__abc_76628_new_n5443_), .Y(u0__abc_76628_new_n5445_));
OR2X2 OR2X2_1473 ( .A(u0__abc_76628_new_n5445_), .B(u0__abc_76628_new_n5442_), .Y(u0__abc_76628_new_n5446_));
OR2X2 OR2X2_1474 ( .A(u0__abc_76628_new_n5448_), .B(u0__abc_76628_new_n5449_), .Y(u0__abc_76628_new_n5450_));
OR2X2 OR2X2_1475 ( .A(u0__abc_76628_new_n5450_), .B(u0__abc_76628_new_n5447_), .Y(u0__abc_76628_new_n5451_));
OR2X2 OR2X2_1476 ( .A(u0__abc_76628_new_n5451_), .B(u0__abc_76628_new_n5446_), .Y(u0__abc_76628_new_n5452_));
OR2X2 OR2X2_1477 ( .A(u0__abc_76628_new_n5455_), .B(u0__abc_76628_new_n5456_), .Y(u0__abc_76628_new_n5457_));
OR2X2 OR2X2_1478 ( .A(u0__abc_76628_new_n5457_), .B(u0__abc_76628_new_n5454_), .Y(u0__abc_76628_new_n5458_));
OR2X2 OR2X2_1479 ( .A(u0__abc_76628_new_n5458_), .B(u0__abc_76628_new_n5453_), .Y(u0__abc_76628_new_n5459_));
OR2X2 OR2X2_148 ( .A(u0__abc_76628_new_n1224_), .B(u0__abc_76628_new_n1202_), .Y(u0__0sp_tms_31_0__1_));
OR2X2 OR2X2_1480 ( .A(u0__abc_76628_new_n5452_), .B(u0__abc_76628_new_n5459_), .Y(u0__abc_76628_new_n5460_));
OR2X2 OR2X2_1481 ( .A(u0__abc_76628_new_n5462_), .B(u0__abc_76628_new_n5463_), .Y(u0__abc_76628_new_n5464_));
OR2X2 OR2X2_1482 ( .A(u0__abc_76628_new_n5464_), .B(u0__abc_76628_new_n5461_), .Y(u0__abc_76628_new_n5465_));
OR2X2 OR2X2_1483 ( .A(u0__abc_76628_new_n5467_), .B(u0__abc_76628_new_n5468_), .Y(u0__abc_76628_new_n5469_));
OR2X2 OR2X2_1484 ( .A(u0__abc_76628_new_n5469_), .B(u0__abc_76628_new_n5466_), .Y(u0__abc_76628_new_n5470_));
OR2X2 OR2X2_1485 ( .A(u0__abc_76628_new_n5472_), .B(u0__abc_76628_new_n5471_), .Y(u0__abc_76628_new_n5473_));
OR2X2 OR2X2_1486 ( .A(u0__abc_76628_new_n5470_), .B(u0__abc_76628_new_n5473_), .Y(u0__abc_76628_new_n5474_));
OR2X2 OR2X2_1487 ( .A(u0__abc_76628_new_n5474_), .B(u0__abc_76628_new_n5465_), .Y(u0__abc_76628_new_n5475_));
OR2X2 OR2X2_1488 ( .A(u0__abc_76628_new_n5460_), .B(u0__abc_76628_new_n5475_), .Y(rf_dout_26_));
OR2X2 OR2X2_1489 ( .A(u0__abc_76628_new_n5477_), .B(u0__abc_76628_new_n5478_), .Y(u0__abc_76628_new_n5479_));
OR2X2 OR2X2_149 ( .A(u0__abc_76628_new_n1177__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n1228_));
OR2X2 OR2X2_1490 ( .A(u0__abc_76628_new_n5480_), .B(u0__abc_76628_new_n5481_), .Y(u0__abc_76628_new_n5482_));
OR2X2 OR2X2_1491 ( .A(u0__abc_76628_new_n5483_), .B(u0__abc_76628_new_n5484_), .Y(u0__abc_76628_new_n5485_));
OR2X2 OR2X2_1492 ( .A(u0__abc_76628_new_n5482_), .B(u0__abc_76628_new_n5485_), .Y(u0__abc_76628_new_n5486_));
OR2X2 OR2X2_1493 ( .A(u0__abc_76628_new_n5486_), .B(u0__abc_76628_new_n5479_), .Y(u0__abc_76628_new_n5487_));
OR2X2 OR2X2_1494 ( .A(u0__abc_76628_new_n5488_), .B(u0__abc_76628_new_n5489_), .Y(u0__abc_76628_new_n5490_));
OR2X2 OR2X2_1495 ( .A(u0__abc_76628_new_n5491_), .B(u0__abc_76628_new_n5492_), .Y(u0__abc_76628_new_n5493_));
OR2X2 OR2X2_1496 ( .A(u0__abc_76628_new_n5490_), .B(u0__abc_76628_new_n5493_), .Y(u0__abc_76628_new_n5494_));
OR2X2 OR2X2_1497 ( .A(u0__abc_76628_new_n5496_), .B(u0__abc_76628_new_n5495_), .Y(u0__abc_76628_new_n5497_));
OR2X2 OR2X2_1498 ( .A(u0__abc_76628_new_n5498_), .B(u0__abc_76628_new_n5499_), .Y(u0__abc_76628_new_n5500_));
OR2X2 OR2X2_1499 ( .A(u0__abc_76628_new_n5497_), .B(u0__abc_76628_new_n5500_), .Y(u0__abc_76628_new_n5501_));
OR2X2 OR2X2_15 ( .A(_abc_85006_new_n240__bF_buf2), .B(spec_req_cs_3_bF_buf5_), .Y(_abc_85006_new_n260_));
OR2X2 OR2X2_150 ( .A(spec_req_cs_6_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1229_));
OR2X2 OR2X2_1500 ( .A(u0__abc_76628_new_n5501_), .B(u0__abc_76628_new_n5494_), .Y(u0__abc_76628_new_n5502_));
OR2X2 OR2X2_1501 ( .A(u0__abc_76628_new_n5505_), .B(u0__abc_76628_new_n5506_), .Y(u0__abc_76628_new_n5507_));
OR2X2 OR2X2_1502 ( .A(u0__abc_76628_new_n5507_), .B(u0__abc_76628_new_n5504_), .Y(u0__abc_76628_new_n5508_));
OR2X2 OR2X2_1503 ( .A(u0__abc_76628_new_n5508_), .B(u0__abc_76628_new_n5503_), .Y(u0__abc_76628_new_n5509_));
OR2X2 OR2X2_1504 ( .A(u0__abc_76628_new_n5502_), .B(u0__abc_76628_new_n5509_), .Y(u0__abc_76628_new_n5510_));
OR2X2 OR2X2_1505 ( .A(u0__abc_76628_new_n5510_), .B(u0__abc_76628_new_n5487_), .Y(rf_dout_27_));
OR2X2 OR2X2_1506 ( .A(u0__abc_76628_new_n5514_), .B(u0__abc_76628_new_n5513_), .Y(u0__abc_76628_new_n5515_));
OR2X2 OR2X2_1507 ( .A(u0__abc_76628_new_n5515_), .B(u0__abc_76628_new_n5512_), .Y(u0__abc_76628_new_n5516_));
OR2X2 OR2X2_1508 ( .A(u0__abc_76628_new_n5518_), .B(u0__abc_76628_new_n5519_), .Y(u0__abc_76628_new_n5520_));
OR2X2 OR2X2_1509 ( .A(u0__abc_76628_new_n5520_), .B(u0__abc_76628_new_n5517_), .Y(u0__abc_76628_new_n5521_));
OR2X2 OR2X2_151 ( .A(u0__abc_76628_new_n1231_), .B(u0__abc_76628_new_n1227_), .Y(u0__abc_76628_new_n1232_));
OR2X2 OR2X2_1510 ( .A(u0__abc_76628_new_n5521_), .B(u0__abc_76628_new_n5516_), .Y(u0__abc_76628_new_n5522_));
OR2X2 OR2X2_1511 ( .A(u0__abc_76628_new_n5525_), .B(u0__abc_76628_new_n5526_), .Y(u0__abc_76628_new_n5527_));
OR2X2 OR2X2_1512 ( .A(u0__abc_76628_new_n5527_), .B(u0__abc_76628_new_n5524_), .Y(u0__abc_76628_new_n5528_));
OR2X2 OR2X2_1513 ( .A(u0__abc_76628_new_n5528_), .B(u0__abc_76628_new_n5523_), .Y(u0__abc_76628_new_n5529_));
OR2X2 OR2X2_1514 ( .A(u0__abc_76628_new_n5522_), .B(u0__abc_76628_new_n5529_), .Y(u0__abc_76628_new_n5530_));
OR2X2 OR2X2_1515 ( .A(u0__abc_76628_new_n5532_), .B(u0__abc_76628_new_n5533_), .Y(u0__abc_76628_new_n5534_));
OR2X2 OR2X2_1516 ( .A(u0__abc_76628_new_n5534_), .B(u0__abc_76628_new_n5531_), .Y(u0__abc_76628_new_n5535_));
OR2X2 OR2X2_1517 ( .A(u0__abc_76628_new_n5537_), .B(u0__abc_76628_new_n5538_), .Y(u0__abc_76628_new_n5539_));
OR2X2 OR2X2_1518 ( .A(u0__abc_76628_new_n5539_), .B(u0__abc_76628_new_n5536_), .Y(u0__abc_76628_new_n5540_));
OR2X2 OR2X2_1519 ( .A(u0__abc_76628_new_n5542_), .B(u0__abc_76628_new_n5541_), .Y(u0__abc_76628_new_n5543_));
OR2X2 OR2X2_152 ( .A(u0__abc_76628_new_n1233_), .B(u0__abc_76628_new_n1234_), .Y(u0__abc_76628_new_n1235_));
OR2X2 OR2X2_1520 ( .A(u0__abc_76628_new_n5540_), .B(u0__abc_76628_new_n5543_), .Y(u0__abc_76628_new_n5544_));
OR2X2 OR2X2_1521 ( .A(u0__abc_76628_new_n5544_), .B(u0__abc_76628_new_n5535_), .Y(u0__abc_76628_new_n5545_));
OR2X2 OR2X2_1522 ( .A(u0__abc_76628_new_n5530_), .B(u0__abc_76628_new_n5545_), .Y(rf_dout_28_));
OR2X2 OR2X2_1523 ( .A(u0__abc_76628_new_n5547_), .B(u0__abc_76628_new_n5548_), .Y(u0__abc_76628_new_n5549_));
OR2X2 OR2X2_1524 ( .A(u0__abc_76628_new_n5551_), .B(u0__abc_76628_new_n5550_), .Y(u0__abc_76628_new_n5552_));
OR2X2 OR2X2_1525 ( .A(u0__abc_76628_new_n5553_), .B(u0__abc_76628_new_n5554_), .Y(u0__abc_76628_new_n5555_));
OR2X2 OR2X2_1526 ( .A(u0__abc_76628_new_n5552_), .B(u0__abc_76628_new_n5555_), .Y(u0__abc_76628_new_n5556_));
OR2X2 OR2X2_1527 ( .A(u0__abc_76628_new_n5556_), .B(u0__abc_76628_new_n5549_), .Y(u0__abc_76628_new_n5557_));
OR2X2 OR2X2_1528 ( .A(u0__abc_76628_new_n5559_), .B(u0__abc_76628_new_n5558_), .Y(u0__abc_76628_new_n5560_));
OR2X2 OR2X2_1529 ( .A(u0__abc_76628_new_n5562_), .B(u0__abc_76628_new_n5561_), .Y(u0__abc_76628_new_n5563_));
OR2X2 OR2X2_153 ( .A(u0__abc_76628_new_n1236_), .B(u0__abc_76628_new_n1237_), .Y(u0__abc_76628_new_n1238_));
OR2X2 OR2X2_1530 ( .A(u0__abc_76628_new_n5560_), .B(u0__abc_76628_new_n5563_), .Y(u0__abc_76628_new_n5564_));
OR2X2 OR2X2_1531 ( .A(u0__abc_76628_new_n5565_), .B(u0__abc_76628_new_n5566_), .Y(u0__abc_76628_new_n5567_));
OR2X2 OR2X2_1532 ( .A(u0__abc_76628_new_n5568_), .B(u0__abc_76628_new_n5569_), .Y(u0__abc_76628_new_n5570_));
OR2X2 OR2X2_1533 ( .A(u0__abc_76628_new_n5567_), .B(u0__abc_76628_new_n5570_), .Y(u0__abc_76628_new_n5571_));
OR2X2 OR2X2_1534 ( .A(u0__abc_76628_new_n5564_), .B(u0__abc_76628_new_n5571_), .Y(u0__abc_76628_new_n5572_));
OR2X2 OR2X2_1535 ( .A(u0__abc_76628_new_n5575_), .B(u0__abc_76628_new_n5576_), .Y(u0__abc_76628_new_n5577_));
OR2X2 OR2X2_1536 ( .A(u0__abc_76628_new_n5577_), .B(u0__abc_76628_new_n5574_), .Y(u0__abc_76628_new_n5578_));
OR2X2 OR2X2_1537 ( .A(u0__abc_76628_new_n5578_), .B(u0__abc_76628_new_n5573_), .Y(u0__abc_76628_new_n5579_));
OR2X2 OR2X2_1538 ( .A(u0__abc_76628_new_n5572_), .B(u0__abc_76628_new_n5579_), .Y(u0__abc_76628_new_n5580_));
OR2X2 OR2X2_1539 ( .A(u0__abc_76628_new_n5580_), .B(u0__abc_76628_new_n5557_), .Y(rf_dout_29_));
OR2X2 OR2X2_154 ( .A(u0__abc_76628_new_n1239_), .B(u0__abc_76628_new_n1240_), .Y(u0__abc_76628_new_n1241_));
OR2X2 OR2X2_1540 ( .A(u0__abc_76628_new_n5582_), .B(u0__abc_76628_new_n5583_), .Y(u0__abc_76628_new_n5584_));
OR2X2 OR2X2_1541 ( .A(u0__abc_76628_new_n5586_), .B(u0__abc_76628_new_n5585_), .Y(u0__abc_76628_new_n5587_));
OR2X2 OR2X2_1542 ( .A(u0__abc_76628_new_n5588_), .B(u0__abc_76628_new_n5589_), .Y(u0__abc_76628_new_n5590_));
OR2X2 OR2X2_1543 ( .A(u0__abc_76628_new_n5587_), .B(u0__abc_76628_new_n5590_), .Y(u0__abc_76628_new_n5591_));
OR2X2 OR2X2_1544 ( .A(u0__abc_76628_new_n5591_), .B(u0__abc_76628_new_n5584_), .Y(u0__abc_76628_new_n5592_));
OR2X2 OR2X2_1545 ( .A(u0__abc_76628_new_n5594_), .B(u0__abc_76628_new_n5593_), .Y(u0__abc_76628_new_n5595_));
OR2X2 OR2X2_1546 ( .A(u0__abc_76628_new_n5597_), .B(u0__abc_76628_new_n5596_), .Y(u0__abc_76628_new_n5598_));
OR2X2 OR2X2_1547 ( .A(u0__abc_76628_new_n5595_), .B(u0__abc_76628_new_n5598_), .Y(u0__abc_76628_new_n5599_));
OR2X2 OR2X2_1548 ( .A(u0__abc_76628_new_n5600_), .B(u0__abc_76628_new_n5601_), .Y(u0__abc_76628_new_n5602_));
OR2X2 OR2X2_1549 ( .A(u0__abc_76628_new_n5603_), .B(u0__abc_76628_new_n5604_), .Y(u0__abc_76628_new_n5605_));
OR2X2 OR2X2_155 ( .A(u0__abc_76628_new_n1243_), .B(spec_req_cs_0_bF_buf0_), .Y(u0__abc_76628_new_n1244_));
OR2X2 OR2X2_1550 ( .A(u0__abc_76628_new_n5602_), .B(u0__abc_76628_new_n5605_), .Y(u0__abc_76628_new_n5606_));
OR2X2 OR2X2_1551 ( .A(u0__abc_76628_new_n5599_), .B(u0__abc_76628_new_n5606_), .Y(u0__abc_76628_new_n5607_));
OR2X2 OR2X2_1552 ( .A(u0__abc_76628_new_n5610_), .B(u0__abc_76628_new_n5611_), .Y(u0__abc_76628_new_n5612_));
OR2X2 OR2X2_1553 ( .A(u0__abc_76628_new_n5612_), .B(u0__abc_76628_new_n5609_), .Y(u0__abc_76628_new_n5613_));
OR2X2 OR2X2_1554 ( .A(u0__abc_76628_new_n5613_), .B(u0__abc_76628_new_n5608_), .Y(u0__abc_76628_new_n5614_));
OR2X2 OR2X2_1555 ( .A(u0__abc_76628_new_n5607_), .B(u0__abc_76628_new_n5614_), .Y(u0__abc_76628_new_n5615_));
OR2X2 OR2X2_1556 ( .A(u0__abc_76628_new_n5615_), .B(u0__abc_76628_new_n5592_), .Y(rf_dout_30_));
OR2X2 OR2X2_1557 ( .A(u0__abc_76628_new_n5617_), .B(u0__abc_76628_new_n5618_), .Y(u0__abc_76628_new_n5619_));
OR2X2 OR2X2_1558 ( .A(u0__abc_76628_new_n5620_), .B(u0__abc_76628_new_n5621_), .Y(u0__abc_76628_new_n5622_));
OR2X2 OR2X2_1559 ( .A(u0__abc_76628_new_n5623_), .B(u0__abc_76628_new_n5624_), .Y(u0__abc_76628_new_n5625_));
OR2X2 OR2X2_156 ( .A(u0__abc_76628_new_n1242_), .B(u0__abc_76628_new_n1244_), .Y(u0__abc_76628_new_n1245_));
OR2X2 OR2X2_1560 ( .A(u0__abc_76628_new_n5625_), .B(u0__abc_76628_new_n5622_), .Y(u0__abc_76628_new_n5626_));
OR2X2 OR2X2_1561 ( .A(u0__abc_76628_new_n5626_), .B(u0__abc_76628_new_n5619_), .Y(u0__abc_76628_new_n5627_));
OR2X2 OR2X2_1562 ( .A(u0__abc_76628_new_n5629_), .B(u0__abc_76628_new_n5628_), .Y(u0__abc_76628_new_n5630_));
OR2X2 OR2X2_1563 ( .A(u0__abc_76628_new_n5632_), .B(u0__abc_76628_new_n5631_), .Y(u0__abc_76628_new_n5633_));
OR2X2 OR2X2_1564 ( .A(u0__abc_76628_new_n5630_), .B(u0__abc_76628_new_n5633_), .Y(u0__abc_76628_new_n5634_));
OR2X2 OR2X2_1565 ( .A(u0__abc_76628_new_n5635_), .B(u0__abc_76628_new_n5636_), .Y(u0__abc_76628_new_n5637_));
OR2X2 OR2X2_1566 ( .A(u0__abc_76628_new_n5638_), .B(u0__abc_76628_new_n5639_), .Y(u0__abc_76628_new_n5640_));
OR2X2 OR2X2_1567 ( .A(u0__abc_76628_new_n5637_), .B(u0__abc_76628_new_n5640_), .Y(u0__abc_76628_new_n5641_));
OR2X2 OR2X2_1568 ( .A(u0__abc_76628_new_n5634_), .B(u0__abc_76628_new_n5641_), .Y(u0__abc_76628_new_n5642_));
OR2X2 OR2X2_1569 ( .A(u0__abc_76628_new_n5645_), .B(u0__abc_76628_new_n5646_), .Y(u0__abc_76628_new_n5647_));
OR2X2 OR2X2_157 ( .A(u0__abc_76628_new_n1197__bF_buf3), .B(u0_tms0_2_), .Y(u0__abc_76628_new_n1246_));
OR2X2 OR2X2_1570 ( .A(u0__abc_76628_new_n5647_), .B(u0__abc_76628_new_n5644_), .Y(u0__abc_76628_new_n5648_));
OR2X2 OR2X2_1571 ( .A(u0__abc_76628_new_n5648_), .B(u0__abc_76628_new_n5643_), .Y(u0__abc_76628_new_n5649_));
OR2X2 OR2X2_1572 ( .A(u0__abc_76628_new_n5642_), .B(u0__abc_76628_new_n5649_), .Y(u0__abc_76628_new_n5650_));
OR2X2 OR2X2_1573 ( .A(u0__abc_76628_new_n5650_), .B(u0__abc_76628_new_n5627_), .Y(rf_dout_31_));
OR2X2 OR2X2_1574 ( .A(u0__abc_76628_new_n5713_), .B(u0__abc_76628_new_n5711_), .Y(u0__abc_76628_new_n5714_));
OR2X2 OR2X2_1575 ( .A(u0__abc_76628_new_n5714_), .B(u0__abc_76628_new_n5709_), .Y(u0__0sreq_cs_le_0_0_));
OR2X2 OR2X2_1576 ( .A(u0_init_req0), .B(u0_init_req1), .Y(u0__abc_76628_new_n5716_));
OR2X2 OR2X2_1577 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n5717_));
OR2X2 OR2X2_1578 ( .A(u0__abc_76628_new_n5716_), .B(u0__abc_76628_new_n5717_), .Y(u0__abc_76628_new_n5718_));
OR2X2 OR2X2_1579 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n5719_));
OR2X2 OR2X2_158 ( .A(u0__abc_76628_new_n1248_), .B(u0__abc_76628_new_n1226_), .Y(u0__0sp_tms_31_0__2_));
OR2X2 OR2X2_1580 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n5720_));
OR2X2 OR2X2_1581 ( .A(u0__abc_76628_new_n5719_), .B(u0__abc_76628_new_n5720_), .Y(u0__abc_76628_new_n5721_));
OR2X2 OR2X2_1582 ( .A(u0__abc_76628_new_n5718_), .B(u0__abc_76628_new_n5721_), .Y(u0__0init_req_0_0_));
OR2X2 OR2X2_1583 ( .A(u0_lmr_req0), .B(u0_lmr_req1), .Y(u0__abc_76628_new_n5723_));
OR2X2 OR2X2_1584 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n5724_));
OR2X2 OR2X2_1585 ( .A(u0__abc_76628_new_n5723_), .B(u0__abc_76628_new_n5724_), .Y(u0__abc_76628_new_n5725_));
OR2X2 OR2X2_1586 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n5726_));
OR2X2 OR2X2_1587 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n5727_));
OR2X2 OR2X2_1588 ( .A(u0__abc_76628_new_n5726_), .B(u0__abc_76628_new_n5727_), .Y(u0__abc_76628_new_n5728_));
OR2X2 OR2X2_1589 ( .A(u0__abc_76628_new_n5725_), .B(u0__abc_76628_new_n5728_), .Y(u0__0lmr_req_0_0_));
OR2X2 OR2X2_159 ( .A(u0__abc_76628_new_n1177__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n1252_));
OR2X2 OR2X2_1590 ( .A(u0_csc0_2_), .B(u0_csc0_1_), .Y(u0_u0__abc_72207_new_n205_));
OR2X2 OR2X2_1591 ( .A(u0_u0__abc_72207_new_n205_), .B(u0_csc0_3_), .Y(u0_u0__abc_72207_new_n206_));
OR2X2 OR2X2_1592 ( .A(u0_u0__abc_72207_new_n213_), .B(u0_u0__abc_72207_new_n209_), .Y(u0_u0__0lmr_req_0_0_));
OR2X2 OR2X2_1593 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf4_), .B(u0_tms0_0_), .Y(u0_u0__abc_72207_new_n223_));
OR2X2 OR2X2_1594 ( .A(u0_u0__abc_72207_new_n224__bF_buf4), .B(\wb_data_i[0] ), .Y(u0_u0__abc_72207_new_n225_));
OR2X2 OR2X2_1595 ( .A(u0_u0__abc_72207_new_n226_), .B(u0_u0_rst_r2_bF_buf5), .Y(u0_u0__0tms_31_0__0_));
OR2X2 OR2X2_1596 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf2_), .B(u0_tms0_1_), .Y(u0_u0__abc_72207_new_n228_));
OR2X2 OR2X2_1597 ( .A(u0_u0__abc_72207_new_n224__bF_buf3), .B(\wb_data_i[1] ), .Y(u0_u0__abc_72207_new_n229_));
OR2X2 OR2X2_1598 ( .A(u0_u0__abc_72207_new_n230_), .B(u0_u0_rst_r2_bF_buf4), .Y(u0_u0__0tms_31_0__1_));
OR2X2 OR2X2_1599 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms0_2_), .Y(u0_u0__abc_72207_new_n232_));
OR2X2 OR2X2_16 ( .A(lmr_sel_bF_buf3), .B(cs_3_), .Y(_abc_85006_new_n261_));
OR2X2 OR2X2_160 ( .A(spec_req_cs_6_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1253_));
OR2X2 OR2X2_1600 ( .A(u0_u0__abc_72207_new_n224__bF_buf2), .B(\wb_data_i[2] ), .Y(u0_u0__abc_72207_new_n233_));
OR2X2 OR2X2_1601 ( .A(u0_u0__abc_72207_new_n234_), .B(u0_u0_rst_r2_bF_buf3), .Y(u0_u0__0tms_31_0__2_));
OR2X2 OR2X2_1602 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf0_), .B(u0_tms0_3_), .Y(u0_u0__abc_72207_new_n236_));
OR2X2 OR2X2_1603 ( .A(u0_u0__abc_72207_new_n224__bF_buf1), .B(\wb_data_i[3] ), .Y(u0_u0__abc_72207_new_n237_));
OR2X2 OR2X2_1604 ( .A(u0_u0__abc_72207_new_n238_), .B(u0_u0_rst_r2_bF_buf2), .Y(u0_u0__0tms_31_0__3_));
OR2X2 OR2X2_1605 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf4_), .B(u0_tms0_4_), .Y(u0_u0__abc_72207_new_n240_));
OR2X2 OR2X2_1606 ( .A(u0_u0__abc_72207_new_n224__bF_buf0), .B(\wb_data_i[4] ), .Y(u0_u0__abc_72207_new_n241_));
OR2X2 OR2X2_1607 ( .A(u0_u0__abc_72207_new_n242_), .B(u0_u0_rst_r2_bF_buf1), .Y(u0_u0__0tms_31_0__4_));
OR2X2 OR2X2_1608 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms0_5_), .Y(u0_u0__abc_72207_new_n244_));
OR2X2 OR2X2_1609 ( .A(u0_u0__abc_72207_new_n224__bF_buf4), .B(\wb_data_i[5] ), .Y(u0_u0__abc_72207_new_n245_));
OR2X2 OR2X2_161 ( .A(u0__abc_76628_new_n1255_), .B(u0__abc_76628_new_n1251_), .Y(u0__abc_76628_new_n1256_));
OR2X2 OR2X2_1610 ( .A(u0_u0__abc_72207_new_n246_), .B(u0_u0_rst_r2_bF_buf0), .Y(u0_u0__0tms_31_0__5_));
OR2X2 OR2X2_1611 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf2_), .B(u0_tms0_6_), .Y(u0_u0__abc_72207_new_n248_));
OR2X2 OR2X2_1612 ( .A(u0_u0__abc_72207_new_n224__bF_buf3), .B(\wb_data_i[6] ), .Y(u0_u0__abc_72207_new_n249_));
OR2X2 OR2X2_1613 ( .A(u0_u0__abc_72207_new_n250_), .B(u0_u0_rst_r2_bF_buf5), .Y(u0_u0__0tms_31_0__6_));
OR2X2 OR2X2_1614 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms0_7_), .Y(u0_u0__abc_72207_new_n252_));
OR2X2 OR2X2_1615 ( .A(u0_u0__abc_72207_new_n224__bF_buf2), .B(\wb_data_i[7] ), .Y(u0_u0__abc_72207_new_n253_));
OR2X2 OR2X2_1616 ( .A(u0_u0__abc_72207_new_n254_), .B(u0_u0_rst_r2_bF_buf4), .Y(u0_u0__0tms_31_0__7_));
OR2X2 OR2X2_1617 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf0_), .B(u0_tms0_8_), .Y(u0_u0__abc_72207_new_n256_));
OR2X2 OR2X2_1618 ( .A(u0_u0__abc_72207_new_n224__bF_buf1), .B(\wb_data_i[8] ), .Y(u0_u0__abc_72207_new_n257_));
OR2X2 OR2X2_1619 ( .A(u0_u0__abc_72207_new_n258_), .B(u0_u0_rst_r2_bF_buf3), .Y(u0_u0__0tms_31_0__8_));
OR2X2 OR2X2_162 ( .A(u0__abc_76628_new_n1257_), .B(u0__abc_76628_new_n1258_), .Y(u0__abc_76628_new_n1259_));
OR2X2 OR2X2_1620 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf4_), .B(u0_tms0_9_), .Y(u0_u0__abc_72207_new_n260_));
OR2X2 OR2X2_1621 ( .A(u0_u0__abc_72207_new_n224__bF_buf0), .B(\wb_data_i[9] ), .Y(u0_u0__abc_72207_new_n261_));
OR2X2 OR2X2_1622 ( .A(u0_u0__abc_72207_new_n262_), .B(u0_u0_rst_r2_bF_buf2), .Y(u0_u0__0tms_31_0__9_));
OR2X2 OR2X2_1623 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms0_10_), .Y(u0_u0__abc_72207_new_n264_));
OR2X2 OR2X2_1624 ( .A(u0_u0__abc_72207_new_n224__bF_buf4), .B(\wb_data_i[10] ), .Y(u0_u0__abc_72207_new_n265_));
OR2X2 OR2X2_1625 ( .A(u0_u0__abc_72207_new_n266_), .B(u0_u0_rst_r2_bF_buf1), .Y(u0_u0__0tms_31_0__10_));
OR2X2 OR2X2_1626 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf2_), .B(u0_tms0_11_), .Y(u0_u0__abc_72207_new_n268_));
OR2X2 OR2X2_1627 ( .A(u0_u0__abc_72207_new_n224__bF_buf3), .B(\wb_data_i[11] ), .Y(u0_u0__abc_72207_new_n269_));
OR2X2 OR2X2_1628 ( .A(u0_u0__abc_72207_new_n270_), .B(u0_u0_rst_r2_bF_buf0), .Y(u0_u0__0tms_31_0__11_));
OR2X2 OR2X2_1629 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms0_12_), .Y(u0_u0__abc_72207_new_n272_));
OR2X2 OR2X2_163 ( .A(u0__abc_76628_new_n1260_), .B(u0__abc_76628_new_n1261_), .Y(u0__abc_76628_new_n1262_));
OR2X2 OR2X2_1630 ( .A(u0_u0__abc_72207_new_n224__bF_buf2), .B(\wb_data_i[12] ), .Y(u0_u0__abc_72207_new_n273_));
OR2X2 OR2X2_1631 ( .A(u0_u0__abc_72207_new_n274_), .B(u0_u0_rst_r2_bF_buf5), .Y(u0_u0__0tms_31_0__12_));
OR2X2 OR2X2_1632 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf0_), .B(u0_tms0_13_), .Y(u0_u0__abc_72207_new_n276_));
OR2X2 OR2X2_1633 ( .A(u0_u0__abc_72207_new_n224__bF_buf1), .B(\wb_data_i[13] ), .Y(u0_u0__abc_72207_new_n277_));
OR2X2 OR2X2_1634 ( .A(u0_u0__abc_72207_new_n278_), .B(u0_u0_rst_r2_bF_buf4), .Y(u0_u0__0tms_31_0__13_));
OR2X2 OR2X2_1635 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf4_), .B(u0_tms0_14_), .Y(u0_u0__abc_72207_new_n280_));
OR2X2 OR2X2_1636 ( .A(u0_u0__abc_72207_new_n224__bF_buf0), .B(\wb_data_i[14] ), .Y(u0_u0__abc_72207_new_n281_));
OR2X2 OR2X2_1637 ( .A(u0_u0__abc_72207_new_n282_), .B(u0_u0_rst_r2_bF_buf3), .Y(u0_u0__0tms_31_0__14_));
OR2X2 OR2X2_1638 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms0_15_), .Y(u0_u0__abc_72207_new_n284_));
OR2X2 OR2X2_1639 ( .A(u0_u0__abc_72207_new_n224__bF_buf4), .B(\wb_data_i[15] ), .Y(u0_u0__abc_72207_new_n285_));
OR2X2 OR2X2_164 ( .A(u0__abc_76628_new_n1263_), .B(u0__abc_76628_new_n1264_), .Y(u0__abc_76628_new_n1265_));
OR2X2 OR2X2_1640 ( .A(u0_u0__abc_72207_new_n286_), .B(u0_u0_rst_r2_bF_buf2), .Y(u0_u0__0tms_31_0__15_));
OR2X2 OR2X2_1641 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf2_), .B(u0_tms0_16_), .Y(u0_u0__abc_72207_new_n288_));
OR2X2 OR2X2_1642 ( .A(u0_u0__abc_72207_new_n224__bF_buf3), .B(\wb_data_i[16] ), .Y(u0_u0__abc_72207_new_n289_));
OR2X2 OR2X2_1643 ( .A(u0_u0__abc_72207_new_n290_), .B(u0_u0_rst_r2_bF_buf1), .Y(u0_u0__0tms_31_0__16_));
OR2X2 OR2X2_1644 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms0_17_), .Y(u0_u0__abc_72207_new_n292_));
OR2X2 OR2X2_1645 ( .A(u0_u0__abc_72207_new_n224__bF_buf2), .B(\wb_data_i[17] ), .Y(u0_u0__abc_72207_new_n293_));
OR2X2 OR2X2_1646 ( .A(u0_u0__abc_72207_new_n294_), .B(u0_u0_rst_r2_bF_buf0), .Y(u0_u0__0tms_31_0__17_));
OR2X2 OR2X2_1647 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf0_), .B(u0_tms0_18_), .Y(u0_u0__abc_72207_new_n296_));
OR2X2 OR2X2_1648 ( .A(u0_u0__abc_72207_new_n224__bF_buf1), .B(\wb_data_i[18] ), .Y(u0_u0__abc_72207_new_n297_));
OR2X2 OR2X2_1649 ( .A(u0_u0__abc_72207_new_n298_), .B(u0_u0_rst_r2_bF_buf5), .Y(u0_u0__0tms_31_0__18_));
OR2X2 OR2X2_165 ( .A(u0__abc_76628_new_n1267_), .B(spec_req_cs_0_bF_buf5_), .Y(u0__abc_76628_new_n1268_));
OR2X2 OR2X2_1650 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf4_), .B(u0_tms0_19_), .Y(u0_u0__abc_72207_new_n300_));
OR2X2 OR2X2_1651 ( .A(u0_u0__abc_72207_new_n224__bF_buf0), .B(\wb_data_i[19] ), .Y(u0_u0__abc_72207_new_n301_));
OR2X2 OR2X2_1652 ( .A(u0_u0__abc_72207_new_n302_), .B(u0_u0_rst_r2_bF_buf4), .Y(u0_u0__0tms_31_0__19_));
OR2X2 OR2X2_1653 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms0_20_), .Y(u0_u0__abc_72207_new_n304_));
OR2X2 OR2X2_1654 ( .A(u0_u0__abc_72207_new_n224__bF_buf4), .B(\wb_data_i[20] ), .Y(u0_u0__abc_72207_new_n305_));
OR2X2 OR2X2_1655 ( .A(u0_u0__abc_72207_new_n306_), .B(u0_u0_rst_r2_bF_buf3), .Y(u0_u0__0tms_31_0__20_));
OR2X2 OR2X2_1656 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf2_), .B(u0_tms0_21_), .Y(u0_u0__abc_72207_new_n308_));
OR2X2 OR2X2_1657 ( .A(u0_u0__abc_72207_new_n224__bF_buf3), .B(\wb_data_i[21] ), .Y(u0_u0__abc_72207_new_n309_));
OR2X2 OR2X2_1658 ( .A(u0_u0__abc_72207_new_n310_), .B(u0_u0_rst_r2_bF_buf2), .Y(u0_u0__0tms_31_0__21_));
OR2X2 OR2X2_1659 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms0_22_), .Y(u0_u0__abc_72207_new_n312_));
OR2X2 OR2X2_166 ( .A(u0__abc_76628_new_n1266_), .B(u0__abc_76628_new_n1268_), .Y(u0__abc_76628_new_n1269_));
OR2X2 OR2X2_1660 ( .A(u0_u0__abc_72207_new_n224__bF_buf2), .B(\wb_data_i[22] ), .Y(u0_u0__abc_72207_new_n313_));
OR2X2 OR2X2_1661 ( .A(u0_u0__abc_72207_new_n314_), .B(u0_u0_rst_r2_bF_buf1), .Y(u0_u0__0tms_31_0__22_));
OR2X2 OR2X2_1662 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf0_), .B(u0_tms0_23_), .Y(u0_u0__abc_72207_new_n316_));
OR2X2 OR2X2_1663 ( .A(u0_u0__abc_72207_new_n224__bF_buf1), .B(\wb_data_i[23] ), .Y(u0_u0__abc_72207_new_n317_));
OR2X2 OR2X2_1664 ( .A(u0_u0__abc_72207_new_n318_), .B(u0_u0_rst_r2_bF_buf0), .Y(u0_u0__0tms_31_0__23_));
OR2X2 OR2X2_1665 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf4_), .B(u0_tms0_24_), .Y(u0_u0__abc_72207_new_n320_));
OR2X2 OR2X2_1666 ( .A(u0_u0__abc_72207_new_n224__bF_buf0), .B(\wb_data_i[24] ), .Y(u0_u0__abc_72207_new_n321_));
OR2X2 OR2X2_1667 ( .A(u0_u0__abc_72207_new_n322_), .B(u0_u0_rst_r2_bF_buf5), .Y(u0_u0__0tms_31_0__24_));
OR2X2 OR2X2_1668 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms0_25_), .Y(u0_u0__abc_72207_new_n324_));
OR2X2 OR2X2_1669 ( .A(u0_u0__abc_72207_new_n224__bF_buf4), .B(\wb_data_i[25] ), .Y(u0_u0__abc_72207_new_n325_));
OR2X2 OR2X2_167 ( .A(u0__abc_76628_new_n1197__bF_buf2), .B(u0_tms0_3_), .Y(u0__abc_76628_new_n1270_));
OR2X2 OR2X2_1670 ( .A(u0_u0__abc_72207_new_n326_), .B(u0_u0_rst_r2_bF_buf4), .Y(u0_u0__0tms_31_0__25_));
OR2X2 OR2X2_1671 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf2_), .B(u0_tms0_26_), .Y(u0_u0__abc_72207_new_n328_));
OR2X2 OR2X2_1672 ( .A(u0_u0__abc_72207_new_n224__bF_buf3), .B(\wb_data_i[26] ), .Y(u0_u0__abc_72207_new_n329_));
OR2X2 OR2X2_1673 ( .A(u0_u0__abc_72207_new_n330_), .B(u0_u0_rst_r2_bF_buf3), .Y(u0_u0__0tms_31_0__26_));
OR2X2 OR2X2_1674 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms0_27_), .Y(u0_u0__abc_72207_new_n332_));
OR2X2 OR2X2_1675 ( .A(u0_u0__abc_72207_new_n224__bF_buf2), .B(\wb_data_i[27] ), .Y(u0_u0__abc_72207_new_n333_));
OR2X2 OR2X2_1676 ( .A(u0_u0__abc_72207_new_n334_), .B(u0_u0_rst_r2_bF_buf2), .Y(u0_u0__0tms_31_0__27_));
OR2X2 OR2X2_1677 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf0_), .B(u0_tms0_28_), .Y(u0_u0__abc_72207_new_n336_));
OR2X2 OR2X2_1678 ( .A(u0_u0__abc_72207_new_n224__bF_buf1), .B(\wb_data_i[28] ), .Y(u0_u0__abc_72207_new_n337_));
OR2X2 OR2X2_1679 ( .A(u0_u0__abc_72207_new_n338_), .B(u0_u0_rst_r2_bF_buf1), .Y(u0_u0__0tms_31_0__28_));
OR2X2 OR2X2_168 ( .A(u0__abc_76628_new_n1272_), .B(u0__abc_76628_new_n1250_), .Y(u0__0sp_tms_31_0__3_));
OR2X2 OR2X2_1680 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf4_), .B(u0_tms0_29_), .Y(u0_u0__abc_72207_new_n340_));
OR2X2 OR2X2_1681 ( .A(u0_u0__abc_72207_new_n224__bF_buf0), .B(\wb_data_i[29] ), .Y(u0_u0__abc_72207_new_n341_));
OR2X2 OR2X2_1682 ( .A(u0_u0__abc_72207_new_n342_), .B(u0_u0_rst_r2_bF_buf0), .Y(u0_u0__0tms_31_0__29_));
OR2X2 OR2X2_1683 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms0_30_), .Y(u0_u0__abc_72207_new_n344_));
OR2X2 OR2X2_1684 ( .A(u0_u0__abc_72207_new_n224__bF_buf4), .B(\wb_data_i[30] ), .Y(u0_u0__abc_72207_new_n345_));
OR2X2 OR2X2_1685 ( .A(u0_u0__abc_72207_new_n346_), .B(u0_u0_rst_r2_bF_buf5), .Y(u0_u0__0tms_31_0__30_));
OR2X2 OR2X2_1686 ( .A(u0_u0__0lmr_req_we_0_0_bF_buf2_), .B(u0_tms0_31_), .Y(u0_u0__abc_72207_new_n348_));
OR2X2 OR2X2_1687 ( .A(u0_u0__abc_72207_new_n224__bF_buf3), .B(\wb_data_i[31] ), .Y(u0_u0__abc_72207_new_n349_));
OR2X2 OR2X2_1688 ( .A(u0_u0__abc_72207_new_n350_), .B(u0_u0_rst_r2_bF_buf4), .Y(u0_u0__0tms_31_0__31_));
OR2X2 OR2X2_1689 ( .A(u0_u0__0init_req_we_0_0_bF_buf4_), .B(u0_csc0_0_), .Y(u0_u0__abc_72207_new_n355_));
OR2X2 OR2X2_169 ( .A(u0__abc_76628_new_n1177__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n1276_));
OR2X2 OR2X2_1690 ( .A(u0_u0_addr_r_6_), .B(u0_u0_addr_r_5_), .Y(u0_u0__abc_72207_new_n358_));
OR2X2 OR2X2_1691 ( .A(u0_u0__abc_72207_new_n358_), .B(u0_u0__abc_72207_new_n357_), .Y(u0_u0__abc_72207_new_n359_));
OR2X2 OR2X2_1692 ( .A(u0_u0__abc_72207_new_n359_), .B(u0_u0__abc_72207_new_n356_), .Y(u0_u0__abc_72207_new_n360_));
OR2X2 OR2X2_1693 ( .A(u0_u0__abc_72207_new_n360_), .B(u0_u0_addr_r_2_), .Y(u0_u0__abc_72207_new_n361_));
OR2X2 OR2X2_1694 ( .A(u0_u0__abc_72207_new_n361__bF_buf4), .B(\wb_data_i[0] ), .Y(u0_u0__abc_72207_new_n362_));
OR2X2 OR2X2_1695 ( .A(u0_u0__abc_72207_new_n365_), .B(u0_u0__abc_72207_new_n366_), .Y(u0_u0__abc_72207_new_n367_));
OR2X2 OR2X2_1696 ( .A(u0_u0__abc_72207_new_n364_), .B(u0_u0__abc_72207_new_n367_), .Y(u0_u0__0csc_31_0__0_));
OR2X2 OR2X2_1697 ( .A(u0_u0__0init_req_we_0_0_bF_buf3_), .B(u0_csc0_1_), .Y(u0_u0__abc_72207_new_n369_));
OR2X2 OR2X2_1698 ( .A(u0_u0__abc_72207_new_n361__bF_buf3), .B(\wb_data_i[1] ), .Y(u0_u0__abc_72207_new_n370_));
OR2X2 OR2X2_1699 ( .A(u0_u0__abc_72207_new_n372_), .B(u0_u0__abc_72207_new_n365_), .Y(u0_u0__0csc_31_0__1_));
OR2X2 OR2X2_17 ( .A(_abc_85006_new_n262_), .B(_abc_85006_new_n237_), .Y(_abc_85006_new_n263_));
OR2X2 OR2X2_170 ( .A(spec_req_cs_6_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1277_));
OR2X2 OR2X2_1700 ( .A(u0_u0__0init_req_we_0_0_bF_buf2_), .B(u0_csc0_2_), .Y(u0_u0__abc_72207_new_n374_));
OR2X2 OR2X2_1701 ( .A(u0_u0__abc_72207_new_n361__bF_buf2), .B(\wb_data_i[2] ), .Y(u0_u0__abc_72207_new_n375_));
OR2X2 OR2X2_1702 ( .A(u0_u0__abc_72207_new_n377_), .B(u0_u0__abc_72207_new_n366_), .Y(u0_u0__0csc_31_0__2_));
OR2X2 OR2X2_1703 ( .A(u0_u0__0init_req_we_0_0_bF_buf1_), .B(u0_csc0_3_), .Y(u0_u0__abc_72207_new_n379_));
OR2X2 OR2X2_1704 ( .A(u0_u0__abc_72207_new_n361__bF_buf1), .B(\wb_data_i[3] ), .Y(u0_u0__abc_72207_new_n380_));
OR2X2 OR2X2_1705 ( .A(u0_u0__0init_req_we_0_0_bF_buf0_), .B(u0_csc0_4_), .Y(u0_u0__abc_72207_new_n383_));
OR2X2 OR2X2_1706 ( .A(u0_u0__abc_72207_new_n361__bF_buf0), .B(\wb_data_i[4] ), .Y(u0_u0__abc_72207_new_n384_));
OR2X2 OR2X2_1707 ( .A(u0_u0__abc_72207_new_n385_), .B(u0_u0_rst_r2_bF_buf0), .Y(u0_u0__abc_72207_new_n386_));
OR2X2 OR2X2_1708 ( .A(u0_u0__abc_72207_new_n354__bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_0_), .Y(u0_u0__abc_72207_new_n387_));
OR2X2 OR2X2_1709 ( .A(u0_u0__0init_req_we_0_0_bF_buf4_), .B(u0_csc0_5_), .Y(u0_u0__abc_72207_new_n389_));
OR2X2 OR2X2_171 ( .A(u0__abc_76628_new_n1279_), .B(u0__abc_76628_new_n1275_), .Y(u0__abc_76628_new_n1280_));
OR2X2 OR2X2_1710 ( .A(u0_u0__abc_72207_new_n361__bF_buf4), .B(\wb_data_i[5] ), .Y(u0_u0__abc_72207_new_n390_));
OR2X2 OR2X2_1711 ( .A(u0_u0__abc_72207_new_n391_), .B(u0_u0_rst_r2_bF_buf5), .Y(u0_u0__abc_72207_new_n392_));
OR2X2 OR2X2_1712 ( .A(u0_u0__abc_72207_new_n354__bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_1_), .Y(u0_u0__abc_72207_new_n393_));
OR2X2 OR2X2_1713 ( .A(u0_u0__0init_req_we_0_0_bF_buf3_), .B(u0_csc0_6_), .Y(u0_u0__abc_72207_new_n395_));
OR2X2 OR2X2_1714 ( .A(u0_u0__abc_72207_new_n361__bF_buf3), .B(\wb_data_i[6] ), .Y(u0_u0__abc_72207_new_n396_));
OR2X2 OR2X2_1715 ( .A(u0_u0__0init_req_we_0_0_bF_buf2_), .B(u0_csc0_7_), .Y(u0_u0__abc_72207_new_n399_));
OR2X2 OR2X2_1716 ( .A(u0_u0__abc_72207_new_n361__bF_buf2), .B(\wb_data_i[7] ), .Y(u0_u0__abc_72207_new_n400_));
OR2X2 OR2X2_1717 ( .A(u0_u0__0init_req_we_0_0_bF_buf1_), .B(u0_csc0_8_), .Y(u0_u0__abc_72207_new_n403_));
OR2X2 OR2X2_1718 ( .A(u0_u0__abc_72207_new_n361__bF_buf1), .B(\wb_data_i[8] ), .Y(u0_u0__abc_72207_new_n404_));
OR2X2 OR2X2_1719 ( .A(u0_u0__0init_req_we_0_0_bF_buf0_), .B(u0_csc0_9_), .Y(u0_u0__abc_72207_new_n407_));
OR2X2 OR2X2_172 ( .A(u0__abc_76628_new_n1281_), .B(u0__abc_76628_new_n1282_), .Y(u0__abc_76628_new_n1283_));
OR2X2 OR2X2_1720 ( .A(u0_u0__abc_72207_new_n361__bF_buf0), .B(\wb_data_i[9] ), .Y(u0_u0__abc_72207_new_n408_));
OR2X2 OR2X2_1721 ( .A(u0_u0__0init_req_we_0_0_bF_buf4_), .B(u0_csc0_10_), .Y(u0_u0__abc_72207_new_n411_));
OR2X2 OR2X2_1722 ( .A(u0_u0__abc_72207_new_n361__bF_buf4), .B(\wb_data_i[10] ), .Y(u0_u0__abc_72207_new_n412_));
OR2X2 OR2X2_1723 ( .A(u0_u0__0init_req_we_0_0_bF_buf3_), .B(u0_csc0_11_), .Y(u0_u0__abc_72207_new_n415_));
OR2X2 OR2X2_1724 ( .A(u0_u0__abc_72207_new_n361__bF_buf3), .B(\wb_data_i[11] ), .Y(u0_u0__abc_72207_new_n416_));
OR2X2 OR2X2_1725 ( .A(u0_u0__0init_req_we_0_0_bF_buf2_), .B(u0_csc0_12_), .Y(u0_u0__abc_72207_new_n419_));
OR2X2 OR2X2_1726 ( .A(u0_u0__abc_72207_new_n361__bF_buf2), .B(\wb_data_i[12] ), .Y(u0_u0__abc_72207_new_n420_));
OR2X2 OR2X2_1727 ( .A(u0_u0__0init_req_we_0_0_bF_buf1_), .B(u0_csc0_13_), .Y(u0_u0__abc_72207_new_n423_));
OR2X2 OR2X2_1728 ( .A(u0_u0__abc_72207_new_n361__bF_buf1), .B(\wb_data_i[13] ), .Y(u0_u0__abc_72207_new_n424_));
OR2X2 OR2X2_1729 ( .A(u0_u0__0init_req_we_0_0_bF_buf0_), .B(u0_csc0_14_), .Y(u0_u0__abc_72207_new_n427_));
OR2X2 OR2X2_173 ( .A(u0__abc_76628_new_n1284_), .B(u0__abc_76628_new_n1285_), .Y(u0__abc_76628_new_n1286_));
OR2X2 OR2X2_1730 ( .A(u0_u0__abc_72207_new_n361__bF_buf0), .B(\wb_data_i[14] ), .Y(u0_u0__abc_72207_new_n428_));
OR2X2 OR2X2_1731 ( .A(u0_u0__0init_req_we_0_0_bF_buf4_), .B(u0_csc0_15_), .Y(u0_u0__abc_72207_new_n431_));
OR2X2 OR2X2_1732 ( .A(u0_u0__abc_72207_new_n361__bF_buf4), .B(\wb_data_i[15] ), .Y(u0_u0__abc_72207_new_n432_));
OR2X2 OR2X2_1733 ( .A(u0_u0__0init_req_we_0_0_bF_buf3_), .B(u0_csc0_16_), .Y(u0_u0__abc_72207_new_n435_));
OR2X2 OR2X2_1734 ( .A(u0_u0__abc_72207_new_n361__bF_buf3), .B(\wb_data_i[16] ), .Y(u0_u0__abc_72207_new_n436_));
OR2X2 OR2X2_1735 ( .A(u0_u0__0init_req_we_0_0_bF_buf2_), .B(u0_csc0_17_), .Y(u0_u0__abc_72207_new_n439_));
OR2X2 OR2X2_1736 ( .A(u0_u0__abc_72207_new_n361__bF_buf2), .B(\wb_data_i[17] ), .Y(u0_u0__abc_72207_new_n440_));
OR2X2 OR2X2_1737 ( .A(u0_u0__0init_req_we_0_0_bF_buf1_), .B(u0_csc0_18_), .Y(u0_u0__abc_72207_new_n443_));
OR2X2 OR2X2_1738 ( .A(u0_u0__abc_72207_new_n361__bF_buf1), .B(\wb_data_i[18] ), .Y(u0_u0__abc_72207_new_n444_));
OR2X2 OR2X2_1739 ( .A(u0_u0__0init_req_we_0_0_bF_buf0_), .B(u0_csc0_19_), .Y(u0_u0__abc_72207_new_n447_));
OR2X2 OR2X2_174 ( .A(u0__abc_76628_new_n1287_), .B(u0__abc_76628_new_n1288_), .Y(u0__abc_76628_new_n1289_));
OR2X2 OR2X2_1740 ( .A(u0_u0__abc_72207_new_n361__bF_buf0), .B(\wb_data_i[19] ), .Y(u0_u0__abc_72207_new_n448_));
OR2X2 OR2X2_1741 ( .A(u0_u0__0init_req_we_0_0_bF_buf4_), .B(u0_csc0_20_), .Y(u0_u0__abc_72207_new_n451_));
OR2X2 OR2X2_1742 ( .A(u0_u0__abc_72207_new_n361__bF_buf4), .B(\wb_data_i[20] ), .Y(u0_u0__abc_72207_new_n452_));
OR2X2 OR2X2_1743 ( .A(u0_u0__0init_req_we_0_0_bF_buf3_), .B(u0_csc0_21_), .Y(u0_u0__abc_72207_new_n455_));
OR2X2 OR2X2_1744 ( .A(u0_u0__abc_72207_new_n361__bF_buf3), .B(\wb_data_i[21] ), .Y(u0_u0__abc_72207_new_n456_));
OR2X2 OR2X2_1745 ( .A(u0_u0__0init_req_we_0_0_bF_buf2_), .B(u0_csc0_22_), .Y(u0_u0__abc_72207_new_n459_));
OR2X2 OR2X2_1746 ( .A(u0_u0__abc_72207_new_n361__bF_buf2), .B(\wb_data_i[22] ), .Y(u0_u0__abc_72207_new_n460_));
OR2X2 OR2X2_1747 ( .A(u0_u0__0init_req_we_0_0_bF_buf1_), .B(u0_csc0_23_), .Y(u0_u0__abc_72207_new_n463_));
OR2X2 OR2X2_1748 ( .A(u0_u0__abc_72207_new_n361__bF_buf1), .B(\wb_data_i[23] ), .Y(u0_u0__abc_72207_new_n464_));
OR2X2 OR2X2_1749 ( .A(u0_u0__0init_req_we_0_0_bF_buf0_), .B(u0_csc0_24_), .Y(u0_u0__abc_72207_new_n467_));
OR2X2 OR2X2_175 ( .A(u0__abc_76628_new_n1291_), .B(spec_req_cs_0_bF_buf4_), .Y(u0__abc_76628_new_n1292_));
OR2X2 OR2X2_1750 ( .A(u0_u0__abc_72207_new_n361__bF_buf0), .B(\wb_data_i[24] ), .Y(u0_u0__abc_72207_new_n468_));
OR2X2 OR2X2_1751 ( .A(u0_u0__0init_req_we_0_0_bF_buf4_), .B(u0_csc0_25_), .Y(u0_u0__abc_72207_new_n471_));
OR2X2 OR2X2_1752 ( .A(u0_u0__abc_72207_new_n361__bF_buf4), .B(\wb_data_i[25] ), .Y(u0_u0__abc_72207_new_n472_));
OR2X2 OR2X2_1753 ( .A(u0_u0__0init_req_we_0_0_bF_buf3_), .B(u0_csc0_26_), .Y(u0_u0__abc_72207_new_n475_));
OR2X2 OR2X2_1754 ( .A(u0_u0__abc_72207_new_n361__bF_buf3), .B(\wb_data_i[26] ), .Y(u0_u0__abc_72207_new_n476_));
OR2X2 OR2X2_1755 ( .A(u0_u0__0init_req_we_0_0_bF_buf2_), .B(u0_csc0_27_), .Y(u0_u0__abc_72207_new_n479_));
OR2X2 OR2X2_1756 ( .A(u0_u0__abc_72207_new_n361__bF_buf2), .B(\wb_data_i[27] ), .Y(u0_u0__abc_72207_new_n480_));
OR2X2 OR2X2_1757 ( .A(u0_u0__0init_req_we_0_0_bF_buf1_), .B(u0_csc0_28_), .Y(u0_u0__abc_72207_new_n483_));
OR2X2 OR2X2_1758 ( .A(u0_u0__abc_72207_new_n361__bF_buf1), .B(\wb_data_i[28] ), .Y(u0_u0__abc_72207_new_n484_));
OR2X2 OR2X2_1759 ( .A(u0_u0__0init_req_we_0_0_bF_buf0_), .B(u0_csc0_29_), .Y(u0_u0__abc_72207_new_n487_));
OR2X2 OR2X2_176 ( .A(u0__abc_76628_new_n1290_), .B(u0__abc_76628_new_n1292_), .Y(u0__abc_76628_new_n1293_));
OR2X2 OR2X2_1760 ( .A(u0_u0__abc_72207_new_n361__bF_buf0), .B(\wb_data_i[29] ), .Y(u0_u0__abc_72207_new_n488_));
OR2X2 OR2X2_1761 ( .A(u0_u0__0init_req_we_0_0_bF_buf4_), .B(u0_csc0_30_), .Y(u0_u0__abc_72207_new_n491_));
OR2X2 OR2X2_1762 ( .A(u0_u0__abc_72207_new_n361__bF_buf4), .B(\wb_data_i[30] ), .Y(u0_u0__abc_72207_new_n492_));
OR2X2 OR2X2_1763 ( .A(u0_u0__0init_req_we_0_0_bF_buf3_), .B(u0_csc0_31_), .Y(u0_u0__abc_72207_new_n495_));
OR2X2 OR2X2_1764 ( .A(u0_u0__abc_72207_new_n361__bF_buf3), .B(\wb_data_i[31] ), .Y(u0_u0__abc_72207_new_n496_));
OR2X2 OR2X2_1765 ( .A(u0_u0__abc_72207_new_n504_), .B(u0_u0__abc_72207_new_n503_), .Y(u0_u0__abc_72207_new_n505_));
OR2X2 OR2X2_1766 ( .A(u0_u0__abc_72207_new_n505_), .B(u0_u0__abc_72207_new_n502_), .Y(u0_u0__abc_72207_new_n506_));
OR2X2 OR2X2_1767 ( .A(u0_u0__abc_72207_new_n511_), .B(u0_u0__abc_72207_new_n508_), .Y(u0_u0__abc_72207_new_n512_));
OR2X2 OR2X2_1768 ( .A(u0_u0__abc_72207_new_n512_), .B(u0_u0__abc_72207_new_n507_), .Y(u0_u0__abc_72207_new_n513_));
OR2X2 OR2X2_1769 ( .A(u0_u0__abc_72207_new_n519_), .B(u0_u0__abc_72207_new_n516_), .Y(u0_u0__abc_72207_new_n520_));
OR2X2 OR2X2_177 ( .A(u0__abc_76628_new_n1197__bF_buf1), .B(u0_tms0_4_), .Y(u0__abc_76628_new_n1294_));
OR2X2 OR2X2_1770 ( .A(u0_u0__abc_72207_new_n520_), .B(u0_u0__abc_72207_new_n515_), .Y(u0_u0__abc_72207_new_n521_));
OR2X2 OR2X2_1771 ( .A(u0_u0__abc_72207_new_n527_), .B(u0_u0__abc_72207_new_n524_), .Y(u0_u0__abc_72207_new_n528_));
OR2X2 OR2X2_1772 ( .A(u0_u0__abc_72207_new_n528_), .B(u0_u0__abc_72207_new_n523_), .Y(u0_u0__abc_72207_new_n529_));
OR2X2 OR2X2_1773 ( .A(u0_u0__abc_72207_new_n535_), .B(u0_u0__abc_72207_new_n532_), .Y(u0_u0__abc_72207_new_n536_));
OR2X2 OR2X2_1774 ( .A(u0_u0__abc_72207_new_n536_), .B(u0_u0__abc_72207_new_n531_), .Y(u0_u0__abc_72207_new_n537_));
OR2X2 OR2X2_1775 ( .A(u0_u0__abc_72207_new_n539_), .B(u0_u0__abc_72207_new_n540_), .Y(u0_u0__abc_72207_new_n541_));
OR2X2 OR2X2_1776 ( .A(u0_u0__abc_72207_new_n542_), .B(u0_u0__abc_72207_new_n538_), .Y(u0_u0__abc_72207_new_n543_));
OR2X2 OR2X2_1777 ( .A(u0_u0__abc_72207_new_n547_), .B(u0_u0__abc_72207_new_n548_), .Y(u0_u0__abc_72207_new_n549_));
OR2X2 OR2X2_1778 ( .A(u0_u0__abc_72207_new_n550_), .B(u0_u0__abc_72207_new_n546_), .Y(u0_u0__abc_72207_new_n551_));
OR2X2 OR2X2_1779 ( .A(u0_u0__abc_72207_new_n554_), .B(u0_u0__abc_72207_new_n555_), .Y(u0_u0__abc_72207_new_n556_));
OR2X2 OR2X2_178 ( .A(u0__abc_76628_new_n1296_), .B(u0__abc_76628_new_n1274_), .Y(u0__0sp_tms_31_0__4_));
OR2X2 OR2X2_1780 ( .A(u0_u0__abc_72207_new_n557_), .B(u0_u0__abc_72207_new_n553_), .Y(u0_u0__abc_72207_new_n558_));
OR2X2 OR2X2_1781 ( .A(u0_u0_inited), .B(u0_init_ack0), .Y(u0_u0__0inited_0_0_));
OR2X2 OR2X2_1782 ( .A(u0_u0__abc_72207_new_n573_), .B(u0_u0__abc_72207_new_n569_), .Y(u0_u0__0init_req_0_0_));
OR2X2 OR2X2_1783 ( .A(u0_csc1_2_), .B(u0_csc1_1_), .Y(u0_u1__abc_72579_new_n201_));
OR2X2 OR2X2_1784 ( .A(u0_u1__abc_72579_new_n201_), .B(u0_csc1_3_), .Y(u0_u1__abc_72579_new_n202_));
OR2X2 OR2X2_1785 ( .A(u0_u1__abc_72579_new_n209_), .B(u0_u1__abc_72579_new_n205_), .Y(u0_u1__0lmr_req_0_0_));
OR2X2 OR2X2_1786 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf7_), .B(u0_tms1_0_), .Y(u0_u1__abc_72579_new_n218_));
OR2X2 OR2X2_1787 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf5_), .B(u0_tms1_1_), .Y(u0_u1__abc_72579_new_n225_));
OR2X2 OR2X2_1788 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms1_2_), .Y(u0_u1__abc_72579_new_n231_));
OR2X2 OR2X2_1789 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms1_3_), .Y(u0_u1__abc_72579_new_n237_));
OR2X2 OR2X2_179 ( .A(u0__abc_76628_new_n1177__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n1300_));
OR2X2 OR2X2_1790 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf7_), .B(u0_tms1_4_), .Y(u0_u1__abc_72579_new_n243_));
OR2X2 OR2X2_1791 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf5_), .B(u0_tms1_5_), .Y(u0_u1__abc_72579_new_n249_));
OR2X2 OR2X2_1792 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms1_6_), .Y(u0_u1__abc_72579_new_n255_));
OR2X2 OR2X2_1793 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms1_7_), .Y(u0_u1__abc_72579_new_n261_));
OR2X2 OR2X2_1794 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf7_), .B(u0_tms1_8_), .Y(u0_u1__abc_72579_new_n267_));
OR2X2 OR2X2_1795 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf5_), .B(u0_tms1_9_), .Y(u0_u1__abc_72579_new_n273_));
OR2X2 OR2X2_1796 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms1_10_), .Y(u0_u1__abc_72579_new_n279_));
OR2X2 OR2X2_1797 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms1_11_), .Y(u0_u1__abc_72579_new_n285_));
OR2X2 OR2X2_1798 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf7_), .B(u0_tms1_12_), .Y(u0_u1__abc_72579_new_n291_));
OR2X2 OR2X2_1799 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf5_), .B(u0_tms1_13_), .Y(u0_u1__abc_72579_new_n297_));
OR2X2 OR2X2_18 ( .A(_abc_85006_new_n245_), .B(cs_need_rfr_3_), .Y(_abc_85006_new_n264_));
OR2X2 OR2X2_180 ( .A(spec_req_cs_6_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1301_));
OR2X2 OR2X2_1800 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms1_14_), .Y(u0_u1__abc_72579_new_n303_));
OR2X2 OR2X2_1801 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms1_15_), .Y(u0_u1__abc_72579_new_n309_));
OR2X2 OR2X2_1802 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf7_), .B(u0_tms1_16_), .Y(u0_u1__abc_72579_new_n315_));
OR2X2 OR2X2_1803 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf5_), .B(u0_tms1_17_), .Y(u0_u1__abc_72579_new_n321_));
OR2X2 OR2X2_1804 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms1_18_), .Y(u0_u1__abc_72579_new_n327_));
OR2X2 OR2X2_1805 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms1_19_), .Y(u0_u1__abc_72579_new_n333_));
OR2X2 OR2X2_1806 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf7_), .B(u0_tms1_20_), .Y(u0_u1__abc_72579_new_n339_));
OR2X2 OR2X2_1807 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf5_), .B(u0_tms1_21_), .Y(u0_u1__abc_72579_new_n345_));
OR2X2 OR2X2_1808 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms1_22_), .Y(u0_u1__abc_72579_new_n351_));
OR2X2 OR2X2_1809 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms1_23_), .Y(u0_u1__abc_72579_new_n357_));
OR2X2 OR2X2_181 ( .A(u0__abc_76628_new_n1303_), .B(u0__abc_76628_new_n1299_), .Y(u0__abc_76628_new_n1304_));
OR2X2 OR2X2_1810 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf7_), .B(u0_tms1_24_), .Y(u0_u1__abc_72579_new_n363_));
OR2X2 OR2X2_1811 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf5_), .B(u0_tms1_25_), .Y(u0_u1__abc_72579_new_n369_));
OR2X2 OR2X2_1812 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms1_26_), .Y(u0_u1__abc_72579_new_n375_));
OR2X2 OR2X2_1813 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms1_27_), .Y(u0_u1__abc_72579_new_n381_));
OR2X2 OR2X2_1814 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf7_), .B(u0_tms1_28_), .Y(u0_u1__abc_72579_new_n387_));
OR2X2 OR2X2_1815 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf5_), .B(u0_tms1_29_), .Y(u0_u1__abc_72579_new_n393_));
OR2X2 OR2X2_1816 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf3_), .B(u0_tms1_30_), .Y(u0_u1__abc_72579_new_n399_));
OR2X2 OR2X2_1817 ( .A(u0_u1__0lmr_req_we_0_0_bF_buf1_), .B(u0_tms1_31_), .Y(u0_u1__abc_72579_new_n405_));
OR2X2 OR2X2_1818 ( .A(u0_u1__0init_req_we_0_0_bF_buf7_), .B(u0_csc1_0_), .Y(u0_u1__abc_72579_new_n413_));
OR2X2 OR2X2_1819 ( .A(u0_u1__0init_req_we_0_0_bF_buf5_), .B(u0_csc1_1_), .Y(u0_u1__abc_72579_new_n418_));
OR2X2 OR2X2_182 ( .A(u0__abc_76628_new_n1305_), .B(u0__abc_76628_new_n1306_), .Y(u0__abc_76628_new_n1307_));
OR2X2 OR2X2_1820 ( .A(u0_u1__0init_req_we_0_0_bF_buf3_), .B(u0_csc1_2_), .Y(u0_u1__abc_72579_new_n423_));
OR2X2 OR2X2_1821 ( .A(u0_u1__0init_req_we_0_0_bF_buf1_), .B(u0_csc1_3_), .Y(u0_u1__abc_72579_new_n428_));
OR2X2 OR2X2_1822 ( .A(u0_u1__0init_req_we_0_0_bF_buf7_), .B(u0_csc1_4_), .Y(u0_u1__abc_72579_new_n433_));
OR2X2 OR2X2_1823 ( .A(u0_u1__0init_req_we_0_0_bF_buf5_), .B(u0_csc1_5_), .Y(u0_u1__abc_72579_new_n438_));
OR2X2 OR2X2_1824 ( .A(u0_u1__0init_req_we_0_0_bF_buf3_), .B(u0_csc1_6_), .Y(u0_u1__abc_72579_new_n443_));
OR2X2 OR2X2_1825 ( .A(u0_u1__0init_req_we_0_0_bF_buf1_), .B(u0_csc1_7_), .Y(u0_u1__abc_72579_new_n448_));
OR2X2 OR2X2_1826 ( .A(u0_u1__0init_req_we_0_0_bF_buf7_), .B(u0_csc1_8_), .Y(u0_u1__abc_72579_new_n453_));
OR2X2 OR2X2_1827 ( .A(u0_u1__0init_req_we_0_0_bF_buf5_), .B(u0_csc1_9_), .Y(u0_u1__abc_72579_new_n458_));
OR2X2 OR2X2_1828 ( .A(u0_u1__0init_req_we_0_0_bF_buf3_), .B(u0_csc1_10_), .Y(u0_u1__abc_72579_new_n463_));
OR2X2 OR2X2_1829 ( .A(u0_u1__0init_req_we_0_0_bF_buf1_), .B(u0_csc1_11_), .Y(u0_u1__abc_72579_new_n468_));
OR2X2 OR2X2_183 ( .A(u0__abc_76628_new_n1308_), .B(u0__abc_76628_new_n1309_), .Y(u0__abc_76628_new_n1310_));
OR2X2 OR2X2_1830 ( .A(u0_u1__0init_req_we_0_0_bF_buf7_), .B(u0_csc1_12_), .Y(u0_u1__abc_72579_new_n473_));
OR2X2 OR2X2_1831 ( .A(u0_u1__0init_req_we_0_0_bF_buf5_), .B(u0_csc1_13_), .Y(u0_u1__abc_72579_new_n478_));
OR2X2 OR2X2_1832 ( .A(u0_u1__0init_req_we_0_0_bF_buf3_), .B(u0_csc1_14_), .Y(u0_u1__abc_72579_new_n483_));
OR2X2 OR2X2_1833 ( .A(u0_u1__0init_req_we_0_0_bF_buf1_), .B(u0_csc1_15_), .Y(u0_u1__abc_72579_new_n488_));
OR2X2 OR2X2_1834 ( .A(u0_u1__0init_req_we_0_0_bF_buf7_), .B(u0_csc1_16_), .Y(u0_u1__abc_72579_new_n493_));
OR2X2 OR2X2_1835 ( .A(u0_u1__0init_req_we_0_0_bF_buf5_), .B(u0_csc1_17_), .Y(u0_u1__abc_72579_new_n498_));
OR2X2 OR2X2_1836 ( .A(u0_u1__0init_req_we_0_0_bF_buf3_), .B(u0_csc1_18_), .Y(u0_u1__abc_72579_new_n503_));
OR2X2 OR2X2_1837 ( .A(u0_u1__0init_req_we_0_0_bF_buf1_), .B(u0_csc1_19_), .Y(u0_u1__abc_72579_new_n508_));
OR2X2 OR2X2_1838 ( .A(u0_u1__0init_req_we_0_0_bF_buf7_), .B(u0_csc1_20_), .Y(u0_u1__abc_72579_new_n513_));
OR2X2 OR2X2_1839 ( .A(u0_u1__0init_req_we_0_0_bF_buf5_), .B(u0_csc1_21_), .Y(u0_u1__abc_72579_new_n518_));
OR2X2 OR2X2_184 ( .A(u0__abc_76628_new_n1311_), .B(u0__abc_76628_new_n1312_), .Y(u0__abc_76628_new_n1313_));
OR2X2 OR2X2_1840 ( .A(u0_u1__0init_req_we_0_0_bF_buf3_), .B(u0_csc1_22_), .Y(u0_u1__abc_72579_new_n523_));
OR2X2 OR2X2_1841 ( .A(u0_u1__0init_req_we_0_0_bF_buf1_), .B(u0_csc1_23_), .Y(u0_u1__abc_72579_new_n528_));
OR2X2 OR2X2_1842 ( .A(u0_u1__0init_req_we_0_0_bF_buf7_), .B(u0_csc1_24_), .Y(u0_u1__abc_72579_new_n533_));
OR2X2 OR2X2_1843 ( .A(u0_u1__0init_req_we_0_0_bF_buf5_), .B(u0_csc1_25_), .Y(u0_u1__abc_72579_new_n538_));
OR2X2 OR2X2_1844 ( .A(u0_u1__0init_req_we_0_0_bF_buf3_), .B(u0_csc1_26_), .Y(u0_u1__abc_72579_new_n543_));
OR2X2 OR2X2_1845 ( .A(u0_u1__0init_req_we_0_0_bF_buf1_), .B(u0_csc1_27_), .Y(u0_u1__abc_72579_new_n548_));
OR2X2 OR2X2_1846 ( .A(u0_u1__0init_req_we_0_0_bF_buf7_), .B(u0_csc1_28_), .Y(u0_u1__abc_72579_new_n553_));
OR2X2 OR2X2_1847 ( .A(u0_u1__0init_req_we_0_0_bF_buf5_), .B(u0_csc1_29_), .Y(u0_u1__abc_72579_new_n558_));
OR2X2 OR2X2_1848 ( .A(u0_u1__0init_req_we_0_0_bF_buf3_), .B(u0_csc1_30_), .Y(u0_u1__abc_72579_new_n563_));
OR2X2 OR2X2_1849 ( .A(u0_u1__0init_req_we_0_0_bF_buf1_), .B(u0_csc1_31_), .Y(u0_u1__abc_72579_new_n568_));
OR2X2 OR2X2_185 ( .A(u0__abc_76628_new_n1315_), .B(spec_req_cs_0_bF_buf3_), .Y(u0__abc_76628_new_n1316_));
OR2X2 OR2X2_1850 ( .A(u0_u1__abc_72579_new_n578_), .B(u0_u1__abc_72579_new_n577_), .Y(u0_u1__abc_72579_new_n579_));
OR2X2 OR2X2_1851 ( .A(u0_u1__abc_72579_new_n579_), .B(u0_u1__abc_72579_new_n576_), .Y(u0_u1__abc_72579_new_n580_));
OR2X2 OR2X2_1852 ( .A(u0_u1__abc_72579_new_n585_), .B(u0_u1__abc_72579_new_n582_), .Y(u0_u1__abc_72579_new_n586_));
OR2X2 OR2X2_1853 ( .A(u0_u1__abc_72579_new_n586_), .B(u0_u1__abc_72579_new_n581_), .Y(u0_u1__abc_72579_new_n587_));
OR2X2 OR2X2_1854 ( .A(u0_u1__abc_72579_new_n593_), .B(u0_u1__abc_72579_new_n590_), .Y(u0_u1__abc_72579_new_n594_));
OR2X2 OR2X2_1855 ( .A(u0_u1__abc_72579_new_n594_), .B(u0_u1__abc_72579_new_n589_), .Y(u0_u1__abc_72579_new_n595_));
OR2X2 OR2X2_1856 ( .A(u0_u1__abc_72579_new_n601_), .B(u0_u1__abc_72579_new_n598_), .Y(u0_u1__abc_72579_new_n602_));
OR2X2 OR2X2_1857 ( .A(u0_u1__abc_72579_new_n602_), .B(u0_u1__abc_72579_new_n597_), .Y(u0_u1__abc_72579_new_n603_));
OR2X2 OR2X2_1858 ( .A(u0_u1__abc_72579_new_n606_), .B(u0_u1__abc_72579_new_n607_), .Y(u0_u1__abc_72579_new_n608_));
OR2X2 OR2X2_1859 ( .A(u0_u1__abc_72579_new_n609_), .B(u0_u1__abc_72579_new_n605_), .Y(u0_u1__abc_72579_new_n610_));
OR2X2 OR2X2_186 ( .A(u0__abc_76628_new_n1314_), .B(u0__abc_76628_new_n1316_), .Y(u0__abc_76628_new_n1317_));
OR2X2 OR2X2_1860 ( .A(u0_u1__abc_72579_new_n613_), .B(u0_u1__abc_72579_new_n614_), .Y(u0_u1__abc_72579_new_n615_));
OR2X2 OR2X2_1861 ( .A(u0_u1__abc_72579_new_n616_), .B(u0_u1__abc_72579_new_n612_), .Y(u0_u1__abc_72579_new_n617_));
OR2X2 OR2X2_1862 ( .A(u0_u1__abc_72579_new_n621_), .B(u0_u1__abc_72579_new_n622_), .Y(u0_u1__abc_72579_new_n623_));
OR2X2 OR2X2_1863 ( .A(u0_u1__abc_72579_new_n624_), .B(u0_u1__abc_72579_new_n620_), .Y(u0_u1__abc_72579_new_n625_));
OR2X2 OR2X2_1864 ( .A(u0_u1__abc_72579_new_n628_), .B(u0_u1__abc_72579_new_n629_), .Y(u0_u1__abc_72579_new_n630_));
OR2X2 OR2X2_1865 ( .A(u0_u1__abc_72579_new_n631_), .B(u0_u1__abc_72579_new_n627_), .Y(u0_u1__abc_72579_new_n632_));
OR2X2 OR2X2_1866 ( .A(u0_u1_inited), .B(u0_init_ack1), .Y(u0_u1__0inited_0_0_));
OR2X2 OR2X2_1867 ( .A(u0_u1__abc_72579_new_n647_), .B(u0_u1__abc_72579_new_n643_), .Y(u0_u1__0init_req_0_0_));
OR2X2 OR2X2_1868 ( .A(csc_s_5_), .B(csc_s_4_), .Y(u1__abc_73140_new_n258_));
OR2X2 OR2X2_1869 ( .A(csc_s_7_), .B(csc_s_6_), .Y(u1__abc_73140_new_n259_));
OR2X2 OR2X2_187 ( .A(u0__abc_76628_new_n1197__bF_buf0), .B(u0_tms0_5_), .Y(u0__abc_76628_new_n1318_));
OR2X2 OR2X2_1870 ( .A(u1__abc_73140_new_n258_), .B(u1__abc_73140_new_n259_), .Y(u1__abc_73140_new_n260_));
OR2X2 OR2X2_1871 ( .A(u1__abc_73140_new_n261_), .B(csc_s_5_), .Y(u1__abc_73140_new_n262_));
OR2X2 OR2X2_1872 ( .A(u1__abc_73140_new_n263_), .B(csc_s_7_), .Y(u1__abc_73140_new_n264_));
OR2X2 OR2X2_1873 ( .A(u1__abc_73140_new_n262_), .B(u1__abc_73140_new_n264_), .Y(u1__abc_73140_new_n265_));
OR2X2 OR2X2_1874 ( .A(u1__abc_73140_new_n274_), .B(u1__abc_73140_new_n278_), .Y(page_size_8_));
OR2X2 OR2X2_1875 ( .A(u1__abc_73140_new_n287_), .B(u1__abc_73140_new_n285_), .Y(u1__abc_73140_new_n288_));
OR2X2 OR2X2_1876 ( .A(u1__abc_73140_new_n288_), .B(u1__abc_73140_new_n284_), .Y(u1__abc_73140_new_n289_));
OR2X2 OR2X2_1877 ( .A(u1__abc_73140_new_n289_), .B(u1_bas_bF_buf3), .Y(u1__abc_73140_new_n290_));
OR2X2 OR2X2_1878 ( .A(u1__abc_73140_new_n291_), .B(u1__abc_73140_new_n292_), .Y(u1__abc_73140_new_n293_));
OR2X2 OR2X2_1879 ( .A(u1__abc_73140_new_n295_), .B(u1__abc_73140_new_n259_), .Y(u1__abc_73140_new_n296_));
OR2X2 OR2X2_188 ( .A(u0__abc_76628_new_n1320_), .B(u0__abc_76628_new_n1298_), .Y(u0__0sp_tms_31_0__5_));
OR2X2 OR2X2_1880 ( .A(u1__abc_73140_new_n274_), .B(u1__abc_73140_new_n300_), .Y(u1__abc_73140_new_n301_));
OR2X2 OR2X2_1881 ( .A(u1__abc_73140_new_n304_), .B(u1__abc_73140_new_n270_), .Y(u1__abc_73140_new_n311_));
OR2X2 OR2X2_1882 ( .A(u1__abc_73140_new_n316_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n317_));
OR2X2 OR2X2_1883 ( .A(u1__abc_73140_new_n313_), .B(u1__abc_73140_new_n317_), .Y(u1__abc_73140_new_n318_));
OR2X2 OR2X2_1884 ( .A(u1__abc_73140_new_n318_), .B(u1__abc_73140_new_n312_), .Y(u1__abc_73140_new_n319_));
OR2X2 OR2X2_1885 ( .A(u1__abc_73140_new_n319_), .B(u1__abc_73140_new_n310_), .Y(u1__abc_73140_new_n320_));
OR2X2 OR2X2_1886 ( .A(u1__abc_73140_new_n309_), .B(u1__abc_73140_new_n320_), .Y(u1__abc_73140_new_n321_));
OR2X2 OR2X2_1887 ( .A(u1__abc_73140_new_n323_), .B(u1__abc_73140_new_n283_), .Y(u1__0bank_adr_1_0__0_));
OR2X2 OR2X2_1888 ( .A(u1__abc_73140_new_n328_), .B(u1__abc_73140_new_n327_), .Y(u1__abc_73140_new_n329_));
OR2X2 OR2X2_1889 ( .A(u1__abc_73140_new_n329_), .B(u1__abc_73140_new_n326_), .Y(u1__abc_73140_new_n330_));
OR2X2 OR2X2_189 ( .A(u0__abc_76628_new_n1177__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n1324_));
OR2X2 OR2X2_1890 ( .A(u1__abc_73140_new_n330_), .B(u1_bas_bF_buf1), .Y(u1__abc_73140_new_n331_));
OR2X2 OR2X2_1891 ( .A(u1__abc_73140_new_n337_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n338_));
OR2X2 OR2X2_1892 ( .A(u1__abc_73140_new_n335_), .B(u1__abc_73140_new_n338_), .Y(u1__abc_73140_new_n339_));
OR2X2 OR2X2_1893 ( .A(u1__abc_73140_new_n339_), .B(u1__abc_73140_new_n334_), .Y(u1__abc_73140_new_n340_));
OR2X2 OR2X2_1894 ( .A(u1__abc_73140_new_n340_), .B(u1__abc_73140_new_n333_), .Y(u1__abc_73140_new_n341_));
OR2X2 OR2X2_1895 ( .A(u1__abc_73140_new_n332_), .B(u1__abc_73140_new_n341_), .Y(u1__abc_73140_new_n342_));
OR2X2 OR2X2_1896 ( .A(u1__abc_73140_new_n344_), .B(u1__abc_73140_new_n325_), .Y(u1__0bank_adr_1_0__1_));
OR2X2 OR2X2_1897 ( .A(u1__abc_73140_new_n349_), .B(u1__abc_73140_new_n348_), .Y(u1__abc_73140_new_n350_));
OR2X2 OR2X2_1898 ( .A(u1__abc_73140_new_n350_), .B(u1__abc_73140_new_n347_), .Y(u1__abc_73140_new_n351_));
OR2X2 OR2X2_1899 ( .A(u1__abc_73140_new_n351_), .B(u1_bas_bF_buf0), .Y(u1__abc_73140_new_n352_));
OR2X2 OR2X2_19 ( .A(_abc_85006_new_n240__bF_buf1), .B(spec_req_cs_4_bF_buf5_), .Y(_abc_85006_new_n266_));
OR2X2 OR2X2_190 ( .A(spec_req_cs_6_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1325_));
OR2X2 OR2X2_1900 ( .A(u1__abc_73140_new_n289_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n353_));
OR2X2 OR2X2_1901 ( .A(u1__abc_73140_new_n355_), .B(u1__abc_73140_new_n346_), .Y(u1__0row_adr_12_0__0_));
OR2X2 OR2X2_1902 ( .A(u1__abc_73140_new_n301_), .B(u1__abc_73140_new_n292_), .Y(u1__abc_73140_new_n358_));
OR2X2 OR2X2_1903 ( .A(u1__abc_73140_new_n368_), .B(u1__abc_73140_new_n367_), .Y(u1__abc_73140_new_n369_));
OR2X2 OR2X2_1904 ( .A(u1__abc_73140_new_n366_), .B(u1__abc_73140_new_n369_), .Y(u1__abc_73140_new_n370_));
OR2X2 OR2X2_1905 ( .A(u1__abc_73140_new_n365_), .B(u1__abc_73140_new_n370_), .Y(u1__abc_73140_new_n371_));
OR2X2 OR2X2_1906 ( .A(u1__abc_73140_new_n371_), .B(u1_bas_bF_buf3), .Y(u1__abc_73140_new_n372_));
OR2X2 OR2X2_1907 ( .A(u1__abc_73140_new_n330_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n373_));
OR2X2 OR2X2_1908 ( .A(u1__abc_73140_new_n375_), .B(u1__abc_73140_new_n357_), .Y(u1__0row_adr_12_0__1_));
OR2X2 OR2X2_1909 ( .A(u1__abc_73140_new_n351_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n378_));
OR2X2 OR2X2_191 ( .A(u0__abc_76628_new_n1327_), .B(u0__abc_76628_new_n1323_), .Y(u0__abc_76628_new_n1328_));
OR2X2 OR2X2_1910 ( .A(u1__abc_73140_new_n382_), .B(u1__abc_73140_new_n381_), .Y(u1__abc_73140_new_n383_));
OR2X2 OR2X2_1911 ( .A(u1__abc_73140_new_n380_), .B(u1__abc_73140_new_n383_), .Y(u1__abc_73140_new_n384_));
OR2X2 OR2X2_1912 ( .A(u1__abc_73140_new_n379_), .B(u1__abc_73140_new_n384_), .Y(u1__abc_73140_new_n385_));
OR2X2 OR2X2_1913 ( .A(u1__abc_73140_new_n385_), .B(u1_bas_bF_buf2), .Y(u1__abc_73140_new_n386_));
OR2X2 OR2X2_1914 ( .A(u1__abc_73140_new_n388_), .B(u1__abc_73140_new_n377_), .Y(u1__0row_adr_12_0__2_));
OR2X2 OR2X2_1915 ( .A(u1__abc_73140_new_n371_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n391_));
OR2X2 OR2X2_1916 ( .A(u1__abc_73140_new_n395_), .B(u1__abc_73140_new_n394_), .Y(u1__abc_73140_new_n396_));
OR2X2 OR2X2_1917 ( .A(u1__abc_73140_new_n393_), .B(u1__abc_73140_new_n396_), .Y(u1__abc_73140_new_n397_));
OR2X2 OR2X2_1918 ( .A(u1__abc_73140_new_n392_), .B(u1__abc_73140_new_n397_), .Y(u1__abc_73140_new_n398_));
OR2X2 OR2X2_1919 ( .A(u1__abc_73140_new_n398_), .B(u1_bas_bF_buf1), .Y(u1__abc_73140_new_n399_));
OR2X2 OR2X2_192 ( .A(u0__abc_76628_new_n1329_), .B(u0__abc_76628_new_n1330_), .Y(u0__abc_76628_new_n1331_));
OR2X2 OR2X2_1920 ( .A(u1__abc_73140_new_n401_), .B(u1__abc_73140_new_n390_), .Y(u1__0row_adr_12_0__3_));
OR2X2 OR2X2_1921 ( .A(u1__abc_73140_new_n407_), .B(u1__abc_73140_new_n406_), .Y(u1__abc_73140_new_n408_));
OR2X2 OR2X2_1922 ( .A(u1__abc_73140_new_n405_), .B(u1__abc_73140_new_n408_), .Y(u1__abc_73140_new_n409_));
OR2X2 OR2X2_1923 ( .A(u1__abc_73140_new_n404_), .B(u1__abc_73140_new_n409_), .Y(u1__abc_73140_new_n410_));
OR2X2 OR2X2_1924 ( .A(u1__abc_73140_new_n410_), .B(u1_bas_bF_buf0), .Y(u1__abc_73140_new_n411_));
OR2X2 OR2X2_1925 ( .A(u1__abc_73140_new_n385_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n412_));
OR2X2 OR2X2_1926 ( .A(u1__abc_73140_new_n414_), .B(u1__abc_73140_new_n403_), .Y(u1__0row_adr_12_0__4_));
OR2X2 OR2X2_1927 ( .A(u1__abc_73140_new_n398_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n417_));
OR2X2 OR2X2_1928 ( .A(u1__abc_73140_new_n421_), .B(u1__abc_73140_new_n420_), .Y(u1__abc_73140_new_n422_));
OR2X2 OR2X2_1929 ( .A(u1__abc_73140_new_n419_), .B(u1__abc_73140_new_n422_), .Y(u1__abc_73140_new_n423_));
OR2X2 OR2X2_193 ( .A(u0__abc_76628_new_n1332_), .B(u0__abc_76628_new_n1333_), .Y(u0__abc_76628_new_n1334_));
OR2X2 OR2X2_1930 ( .A(u1__abc_73140_new_n418_), .B(u1__abc_73140_new_n423_), .Y(u1__abc_73140_new_n424_));
OR2X2 OR2X2_1931 ( .A(u1__abc_73140_new_n424_), .B(u1_bas_bF_buf3), .Y(u1__abc_73140_new_n425_));
OR2X2 OR2X2_1932 ( .A(u1__abc_73140_new_n427_), .B(u1__abc_73140_new_n416_), .Y(u1__0row_adr_12_0__5_));
OR2X2 OR2X2_1933 ( .A(u1__abc_73140_new_n410_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n430_));
OR2X2 OR2X2_1934 ( .A(u1__abc_73140_new_n434_), .B(u1__abc_73140_new_n433_), .Y(u1__abc_73140_new_n435_));
OR2X2 OR2X2_1935 ( .A(u1__abc_73140_new_n432_), .B(u1__abc_73140_new_n435_), .Y(u1__abc_73140_new_n436_));
OR2X2 OR2X2_1936 ( .A(u1__abc_73140_new_n431_), .B(u1__abc_73140_new_n436_), .Y(u1__abc_73140_new_n437_));
OR2X2 OR2X2_1937 ( .A(u1__abc_73140_new_n437_), .B(u1_bas_bF_buf2), .Y(u1__abc_73140_new_n438_));
OR2X2 OR2X2_1938 ( .A(u1__abc_73140_new_n440_), .B(u1__abc_73140_new_n429_), .Y(u1__0row_adr_12_0__6_));
OR2X2 OR2X2_1939 ( .A(u1__abc_73140_new_n424_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n443_));
OR2X2 OR2X2_194 ( .A(u0__abc_76628_new_n1335_), .B(u0__abc_76628_new_n1336_), .Y(u0__abc_76628_new_n1337_));
OR2X2 OR2X2_1940 ( .A(u1__abc_73140_new_n445_), .B(u1__abc_73140_new_n446_), .Y(u1__abc_73140_new_n447_));
OR2X2 OR2X2_1941 ( .A(u1__abc_73140_new_n447_), .B(u1__abc_73140_new_n444_), .Y(u1__abc_73140_new_n448_));
OR2X2 OR2X2_1942 ( .A(u1__abc_73140_new_n448_), .B(u1_bas_bF_buf1), .Y(u1__abc_73140_new_n449_));
OR2X2 OR2X2_1943 ( .A(u1__abc_73140_new_n451_), .B(u1__abc_73140_new_n442_), .Y(u1__0row_adr_12_0__7_));
OR2X2 OR2X2_1944 ( .A(u1__abc_73140_new_n437_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n454_));
OR2X2 OR2X2_1945 ( .A(u1__abc_73140_new_n456_), .B(u1__abc_73140_new_n457_), .Y(u1__abc_73140_new_n458_));
OR2X2 OR2X2_1946 ( .A(u1__abc_73140_new_n458_), .B(u1__abc_73140_new_n455_), .Y(u1__abc_73140_new_n459_));
OR2X2 OR2X2_1947 ( .A(u1__abc_73140_new_n459_), .B(u1_bas_bF_buf0), .Y(u1__abc_73140_new_n460_));
OR2X2 OR2X2_1948 ( .A(u1__abc_73140_new_n462_), .B(u1__abc_73140_new_n453_), .Y(u1__0row_adr_12_0__8_));
OR2X2 OR2X2_1949 ( .A(u1__abc_73140_new_n448_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n465_));
OR2X2 OR2X2_195 ( .A(u0__abc_76628_new_n1339_), .B(spec_req_cs_0_bF_buf2_), .Y(u0__abc_76628_new_n1340_));
OR2X2 OR2X2_1950 ( .A(u1__abc_73140_new_n467_), .B(u1__abc_73140_new_n468_), .Y(u1__abc_73140_new_n469_));
OR2X2 OR2X2_1951 ( .A(u1__abc_73140_new_n471_), .B(u1__abc_73140_new_n470_), .Y(u1__abc_73140_new_n472_));
OR2X2 OR2X2_1952 ( .A(u1__abc_73140_new_n316_), .B(u1_bas_bF_buf3), .Y(u1__abc_73140_new_n473_));
OR2X2 OR2X2_1953 ( .A(u1__abc_73140_new_n472_), .B(u1__abc_73140_new_n473_), .Y(u1__abc_73140_new_n474_));
OR2X2 OR2X2_1954 ( .A(u1__abc_73140_new_n474_), .B(u1__abc_73140_new_n469_), .Y(u1__abc_73140_new_n475_));
OR2X2 OR2X2_1955 ( .A(u1__abc_73140_new_n475_), .B(u1__abc_73140_new_n466_), .Y(u1__abc_73140_new_n476_));
OR2X2 OR2X2_1956 ( .A(u1__abc_73140_new_n478_), .B(u1__abc_73140_new_n464_), .Y(u1__0row_adr_12_0__9_));
OR2X2 OR2X2_1957 ( .A(u1__abc_73140_new_n459_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n481_));
OR2X2 OR2X2_1958 ( .A(u1__abc_73140_new_n337_), .B(u1_bas_bF_buf2), .Y(u1__abc_73140_new_n484_));
OR2X2 OR2X2_1959 ( .A(u1__abc_73140_new_n484_), .B(u1__abc_73140_new_n483_), .Y(u1__abc_73140_new_n485_));
OR2X2 OR2X2_196 ( .A(u0__abc_76628_new_n1338_), .B(u0__abc_76628_new_n1340_), .Y(u0__abc_76628_new_n1341_));
OR2X2 OR2X2_1960 ( .A(u1__abc_73140_new_n486_), .B(u1__abc_73140_new_n488_), .Y(u1__abc_73140_new_n489_));
OR2X2 OR2X2_1961 ( .A(u1__abc_73140_new_n490_), .B(u1__abc_73140_new_n313_), .Y(u1__abc_73140_new_n491_));
OR2X2 OR2X2_1962 ( .A(u1__abc_73140_new_n491_), .B(u1__abc_73140_new_n489_), .Y(u1__abc_73140_new_n492_));
OR2X2 OR2X2_1963 ( .A(u1__abc_73140_new_n492_), .B(u1__abc_73140_new_n485_), .Y(u1__abc_73140_new_n493_));
OR2X2 OR2X2_1964 ( .A(u1__abc_73140_new_n493_), .B(u1__abc_73140_new_n482_), .Y(u1__abc_73140_new_n494_));
OR2X2 OR2X2_1965 ( .A(u1__abc_73140_new_n496_), .B(u1__abc_73140_new_n480_), .Y(u1__0row_adr_12_0__10_));
OR2X2 OR2X2_1966 ( .A(u1__abc_73140_new_n472_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n499_));
OR2X2 OR2X2_1967 ( .A(u1__abc_73140_new_n499_), .B(u1__abc_73140_new_n469_), .Y(u1__abc_73140_new_n500_));
OR2X2 OR2X2_1968 ( .A(u1__abc_73140_new_n500_), .B(u1__abc_73140_new_n466_), .Y(u1__abc_73140_new_n501_));
OR2X2 OR2X2_1969 ( .A(u1__abc_73140_new_n504_), .B(u1_bas_bF_buf1), .Y(u1__abc_73140_new_n505_));
OR2X2 OR2X2_197 ( .A(u0__abc_76628_new_n1197__bF_buf5), .B(u0_tms0_6_), .Y(u0__abc_76628_new_n1342_));
OR2X2 OR2X2_1970 ( .A(u1__abc_73140_new_n505_), .B(u1__abc_73140_new_n503_), .Y(u1__abc_73140_new_n506_));
OR2X2 OR2X2_1971 ( .A(u1__abc_73140_new_n506_), .B(u1__abc_73140_new_n502_), .Y(u1__abc_73140_new_n507_));
OR2X2 OR2X2_1972 ( .A(u1__abc_73140_new_n509_), .B(u1__abc_73140_new_n498_), .Y(u1__0row_adr_12_0__11_));
OR2X2 OR2X2_1973 ( .A(u1__abc_73140_new_n511_), .B(u1_bas_bF_buf0), .Y(u1__abc_73140_new_n512_));
OR2X2 OR2X2_1974 ( .A(u1__abc_73140_new_n513_), .B(u1__abc_73140_new_n515_), .Y(u1__abc_73140_new_n516_));
OR2X2 OR2X2_1975 ( .A(u1__abc_73140_new_n516_), .B(u1__abc_73140_new_n512_), .Y(u1__abc_73140_new_n517_));
OR2X2 OR2X2_1976 ( .A(u1__abc_73140_new_n483_), .B(u1__abc_73140_new_n314_), .Y(u1__abc_73140_new_n518_));
OR2X2 OR2X2_1977 ( .A(u1__abc_73140_new_n489_), .B(u1__abc_73140_new_n518_), .Y(u1__abc_73140_new_n519_));
OR2X2 OR2X2_1978 ( .A(u1__abc_73140_new_n520_), .B(u1__abc_73140_new_n282_), .Y(u1__abc_73140_new_n521_));
OR2X2 OR2X2_1979 ( .A(cs_le_bF_buf4), .B(row_adr_12_bF_buf3_), .Y(u1__abc_73140_new_n522_));
OR2X2 OR2X2_198 ( .A(u0__abc_76628_new_n1344_), .B(u0__abc_76628_new_n1322_), .Y(u0__0sp_tms_31_0__6_));
OR2X2 OR2X2_1980 ( .A(u1__abc_73140_new_n525_), .B(u1__abc_73140_new_n526_), .Y(u1__abc_73140_new_n527_));
OR2X2 OR2X2_1981 ( .A(u1__abc_73140_new_n528_), .B(\wb_addr_i[2] ), .Y(u1__abc_73140_new_n529_));
OR2X2 OR2X2_1982 ( .A(u1__abc_73140_new_n527_), .B(u1_col_adr_0_), .Y(u1__abc_73140_new_n530_));
OR2X2 OR2X2_1983 ( .A(u1__abc_73140_new_n528_), .B(\wb_addr_i[3] ), .Y(u1__abc_73140_new_n532_));
OR2X2 OR2X2_1984 ( .A(u1__abc_73140_new_n527_), .B(u1_col_adr_1_), .Y(u1__abc_73140_new_n533_));
OR2X2 OR2X2_1985 ( .A(u1__abc_73140_new_n528_), .B(\wb_addr_i[4] ), .Y(u1__abc_73140_new_n535_));
OR2X2 OR2X2_1986 ( .A(u1__abc_73140_new_n527_), .B(u1_col_adr_2_), .Y(u1__abc_73140_new_n536_));
OR2X2 OR2X2_1987 ( .A(u1__abc_73140_new_n528_), .B(\wb_addr_i[5] ), .Y(u1__abc_73140_new_n538_));
OR2X2 OR2X2_1988 ( .A(u1__abc_73140_new_n527_), .B(u1_col_adr_3_), .Y(u1__abc_73140_new_n539_));
OR2X2 OR2X2_1989 ( .A(u1__abc_73140_new_n528_), .B(\wb_addr_i[6] ), .Y(u1__abc_73140_new_n541_));
OR2X2 OR2X2_199 ( .A(u0__abc_76628_new_n1177__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n1348_));
OR2X2 OR2X2_1990 ( .A(u1__abc_73140_new_n527_), .B(u1_col_adr_4_), .Y(u1__abc_73140_new_n542_));
OR2X2 OR2X2_1991 ( .A(u1__abc_73140_new_n528_), .B(\wb_addr_i[7] ), .Y(u1__abc_73140_new_n544_));
OR2X2 OR2X2_1992 ( .A(u1__abc_73140_new_n527_), .B(u1_col_adr_5_), .Y(u1__abc_73140_new_n545_));
OR2X2 OR2X2_1993 ( .A(u1__abc_73140_new_n528_), .B(\wb_addr_i[8] ), .Y(u1__abc_73140_new_n547_));
OR2X2 OR2X2_1994 ( .A(u1__abc_73140_new_n527_), .B(u1_col_adr_6_), .Y(u1__abc_73140_new_n548_));
OR2X2 OR2X2_1995 ( .A(u1__abc_73140_new_n528_), .B(\wb_addr_i[9] ), .Y(u1__abc_73140_new_n550_));
OR2X2 OR2X2_1996 ( .A(u1__abc_73140_new_n527_), .B(u1_col_adr_7_), .Y(u1__abc_73140_new_n551_));
OR2X2 OR2X2_1997 ( .A(u1__abc_73140_new_n555_), .B(u1__abc_73140_new_n553_), .Y(u1__0col_adr_9_0__8_));
OR2X2 OR2X2_1998 ( .A(u1__abc_73140_new_n559_), .B(u1__abc_73140_new_n557_), .Y(u1__0col_adr_9_0__9_));
OR2X2 OR2X2_1999 ( .A(cs_le_bF_buf3), .B(wb_we_i), .Y(u1__abc_73140_new_n561_));
OR2X2 OR2X2_2 ( .A(susp_sel), .B(rfr_ack), .Y(_abc_85006_new_n237_));
OR2X2 OR2X2_20 ( .A(lmr_sel_bF_buf2), .B(cs_4_), .Y(_abc_85006_new_n267_));
OR2X2 OR2X2_200 ( .A(spec_req_cs_6_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1349_));
OR2X2 OR2X2_2000 ( .A(u1_acs_addr_0_), .B(next_adr_bF_buf4), .Y(u1__abc_73140_new_n562_));
OR2X2 OR2X2_2001 ( .A(u1__abc_73140_new_n563__bF_buf3), .B(u1_acs_addr_pl1_0_), .Y(u1__abc_73140_new_n564_));
OR2X2 OR2X2_2002 ( .A(u1__abc_73140_new_n565_), .B(u1__abc_73140_new_n561__bF_buf4), .Y(u1__abc_73140_new_n566_));
OR2X2 OR2X2_2003 ( .A(u1__abc_73140_new_n571_), .B(u1__abc_73140_new_n570__bF_buf3), .Y(u1__abc_73140_new_n572_));
OR2X2 OR2X2_2004 ( .A(u1__abc_73140_new_n572_), .B(u1__abc_73140_new_n569_), .Y(u1__abc_73140_new_n573_));
OR2X2 OR2X2_2005 ( .A(u1__abc_73140_new_n573_), .B(u1__abc_73140_new_n568_), .Y(u1__abc_73140_new_n574_));
OR2X2 OR2X2_2006 ( .A(next_adr_bF_buf2), .B(u1_acs_addr_1_), .Y(u1__abc_73140_new_n576_));
OR2X2 OR2X2_2007 ( .A(u1__abc_73140_new_n563__bF_buf2), .B(u1_acs_addr_pl1_1_), .Y(u1__abc_73140_new_n577_));
OR2X2 OR2X2_2008 ( .A(u1__abc_73140_new_n578_), .B(u1__abc_73140_new_n561__bF_buf2), .Y(u1__abc_73140_new_n579_));
OR2X2 OR2X2_2009 ( .A(u1__abc_73140_new_n582_), .B(u1__abc_73140_new_n570__bF_buf2), .Y(u1__abc_73140_new_n583_));
OR2X2 OR2X2_201 ( .A(u0__abc_76628_new_n1351_), .B(u0__abc_76628_new_n1347_), .Y(u0__abc_76628_new_n1352_));
OR2X2 OR2X2_2010 ( .A(u1__abc_73140_new_n583_), .B(u1__abc_73140_new_n581_), .Y(u1__abc_73140_new_n584_));
OR2X2 OR2X2_2011 ( .A(u1__abc_73140_new_n584_), .B(u1__abc_73140_new_n580_), .Y(u1__abc_73140_new_n585_));
OR2X2 OR2X2_2012 ( .A(next_adr_bF_buf1), .B(u1_acs_addr_2_), .Y(u1__abc_73140_new_n587_));
OR2X2 OR2X2_2013 ( .A(u1__abc_73140_new_n563__bF_buf1), .B(u1_acs_addr_pl1_2_), .Y(u1__abc_73140_new_n588_));
OR2X2 OR2X2_2014 ( .A(u1__abc_73140_new_n589_), .B(u1__abc_73140_new_n561__bF_buf1), .Y(u1__abc_73140_new_n590_));
OR2X2 OR2X2_2015 ( .A(u1__abc_73140_new_n593_), .B(u1__abc_73140_new_n570__bF_buf1), .Y(u1__abc_73140_new_n594_));
OR2X2 OR2X2_2016 ( .A(u1__abc_73140_new_n594_), .B(u1__abc_73140_new_n592_), .Y(u1__abc_73140_new_n595_));
OR2X2 OR2X2_2017 ( .A(u1__abc_73140_new_n595_), .B(u1__abc_73140_new_n591_), .Y(u1__abc_73140_new_n596_));
OR2X2 OR2X2_2018 ( .A(next_adr_bF_buf0), .B(u1_acs_addr_3_), .Y(u1__abc_73140_new_n598_));
OR2X2 OR2X2_2019 ( .A(u1__abc_73140_new_n563__bF_buf0), .B(u1_acs_addr_pl1_3_), .Y(u1__abc_73140_new_n599_));
OR2X2 OR2X2_202 ( .A(u0__abc_76628_new_n1353_), .B(u0__abc_76628_new_n1354_), .Y(u0__abc_76628_new_n1355_));
OR2X2 OR2X2_2020 ( .A(u1__abc_73140_new_n600_), .B(u1__abc_73140_new_n561__bF_buf0), .Y(u1__abc_73140_new_n601_));
OR2X2 OR2X2_2021 ( .A(u1__abc_73140_new_n604_), .B(u1__abc_73140_new_n570__bF_buf0), .Y(u1__abc_73140_new_n605_));
OR2X2 OR2X2_2022 ( .A(u1__abc_73140_new_n605_), .B(u1__abc_73140_new_n603_), .Y(u1__abc_73140_new_n606_));
OR2X2 OR2X2_2023 ( .A(u1__abc_73140_new_n606_), .B(u1__abc_73140_new_n602_), .Y(u1__abc_73140_new_n607_));
OR2X2 OR2X2_2024 ( .A(next_adr_bF_buf4), .B(u1_acs_addr_4_), .Y(u1__abc_73140_new_n609_));
OR2X2 OR2X2_2025 ( .A(u1__abc_73140_new_n563__bF_buf3), .B(u1_acs_addr_pl1_4_), .Y(u1__abc_73140_new_n610_));
OR2X2 OR2X2_2026 ( .A(u1__abc_73140_new_n611_), .B(u1__abc_73140_new_n561__bF_buf4), .Y(u1__abc_73140_new_n612_));
OR2X2 OR2X2_2027 ( .A(u1__abc_73140_new_n615_), .B(u1__abc_73140_new_n570__bF_buf3), .Y(u1__abc_73140_new_n616_));
OR2X2 OR2X2_2028 ( .A(u1__abc_73140_new_n616_), .B(u1__abc_73140_new_n614_), .Y(u1__abc_73140_new_n617_));
OR2X2 OR2X2_2029 ( .A(u1__abc_73140_new_n617_), .B(u1__abc_73140_new_n613_), .Y(u1__abc_73140_new_n618_));
OR2X2 OR2X2_203 ( .A(u0__abc_76628_new_n1356_), .B(u0__abc_76628_new_n1357_), .Y(u0__abc_76628_new_n1358_));
OR2X2 OR2X2_2030 ( .A(next_adr_bF_buf3), .B(u1_acs_addr_5_), .Y(u1__abc_73140_new_n620_));
OR2X2 OR2X2_2031 ( .A(u1__abc_73140_new_n563__bF_buf2), .B(u1_acs_addr_pl1_5_), .Y(u1__abc_73140_new_n621_));
OR2X2 OR2X2_2032 ( .A(u1__abc_73140_new_n622_), .B(u1__abc_73140_new_n561__bF_buf3), .Y(u1__abc_73140_new_n623_));
OR2X2 OR2X2_2033 ( .A(u1__abc_73140_new_n626_), .B(u1__abc_73140_new_n570__bF_buf2), .Y(u1__abc_73140_new_n627_));
OR2X2 OR2X2_2034 ( .A(u1__abc_73140_new_n627_), .B(u1__abc_73140_new_n625_), .Y(u1__abc_73140_new_n628_));
OR2X2 OR2X2_2035 ( .A(u1__abc_73140_new_n628_), .B(u1__abc_73140_new_n624_), .Y(u1__abc_73140_new_n629_));
OR2X2 OR2X2_2036 ( .A(next_adr_bF_buf2), .B(u1_acs_addr_6_), .Y(u1__abc_73140_new_n631_));
OR2X2 OR2X2_2037 ( .A(u1__abc_73140_new_n563__bF_buf1), .B(u1_acs_addr_pl1_6_), .Y(u1__abc_73140_new_n632_));
OR2X2 OR2X2_2038 ( .A(u1__abc_73140_new_n633_), .B(u1__abc_73140_new_n561__bF_buf2), .Y(u1__abc_73140_new_n634_));
OR2X2 OR2X2_2039 ( .A(u1__abc_73140_new_n637_), .B(u1__abc_73140_new_n570__bF_buf1), .Y(u1__abc_73140_new_n638_));
OR2X2 OR2X2_204 ( .A(u0__abc_76628_new_n1359_), .B(u0__abc_76628_new_n1360_), .Y(u0__abc_76628_new_n1361_));
OR2X2 OR2X2_2040 ( .A(u1__abc_73140_new_n638_), .B(u1__abc_73140_new_n636_), .Y(u1__abc_73140_new_n639_));
OR2X2 OR2X2_2041 ( .A(u1__abc_73140_new_n639_), .B(u1__abc_73140_new_n635_), .Y(u1__abc_73140_new_n640_));
OR2X2 OR2X2_2042 ( .A(next_adr_bF_buf1), .B(u1_acs_addr_7_), .Y(u1__abc_73140_new_n642_));
OR2X2 OR2X2_2043 ( .A(u1__abc_73140_new_n563__bF_buf0), .B(u1_acs_addr_pl1_7_), .Y(u1__abc_73140_new_n643_));
OR2X2 OR2X2_2044 ( .A(u1__abc_73140_new_n644_), .B(u1__abc_73140_new_n561__bF_buf1), .Y(u1__abc_73140_new_n645_));
OR2X2 OR2X2_2045 ( .A(u1__abc_73140_new_n648_), .B(u1__abc_73140_new_n570__bF_buf0), .Y(u1__abc_73140_new_n649_));
OR2X2 OR2X2_2046 ( .A(u1__abc_73140_new_n649_), .B(u1__abc_73140_new_n647_), .Y(u1__abc_73140_new_n650_));
OR2X2 OR2X2_2047 ( .A(u1__abc_73140_new_n650_), .B(u1__abc_73140_new_n646_), .Y(u1__abc_73140_new_n651_));
OR2X2 OR2X2_2048 ( .A(next_adr_bF_buf0), .B(u1_acs_addr_8_), .Y(u1__abc_73140_new_n653_));
OR2X2 OR2X2_2049 ( .A(u1__abc_73140_new_n563__bF_buf3), .B(u1_acs_addr_pl1_8_), .Y(u1__abc_73140_new_n654_));
OR2X2 OR2X2_205 ( .A(u0__abc_76628_new_n1363_), .B(spec_req_cs_0_bF_buf1_), .Y(u0__abc_76628_new_n1364_));
OR2X2 OR2X2_2050 ( .A(u1__abc_73140_new_n655_), .B(u1__abc_73140_new_n561__bF_buf0), .Y(u1__abc_73140_new_n656_));
OR2X2 OR2X2_2051 ( .A(u1__abc_73140_new_n659_), .B(u1__abc_73140_new_n570__bF_buf3), .Y(u1__abc_73140_new_n660_));
OR2X2 OR2X2_2052 ( .A(u1__abc_73140_new_n660_), .B(u1__abc_73140_new_n658_), .Y(u1__abc_73140_new_n661_));
OR2X2 OR2X2_2053 ( .A(u1__abc_73140_new_n661_), .B(u1__abc_73140_new_n657_), .Y(u1__abc_73140_new_n662_));
OR2X2 OR2X2_2054 ( .A(next_adr_bF_buf4), .B(u1_acs_addr_9_), .Y(u1__abc_73140_new_n664_));
OR2X2 OR2X2_2055 ( .A(u1__abc_73140_new_n563__bF_buf2), .B(u1_acs_addr_pl1_9_), .Y(u1__abc_73140_new_n665_));
OR2X2 OR2X2_2056 ( .A(u1__abc_73140_new_n666_), .B(u1__abc_73140_new_n561__bF_buf4), .Y(u1__abc_73140_new_n667_));
OR2X2 OR2X2_2057 ( .A(u1__abc_73140_new_n670_), .B(u1__abc_73140_new_n570__bF_buf2), .Y(u1__abc_73140_new_n671_));
OR2X2 OR2X2_2058 ( .A(u1__abc_73140_new_n671_), .B(u1__abc_73140_new_n669_), .Y(u1__abc_73140_new_n672_));
OR2X2 OR2X2_2059 ( .A(u1__abc_73140_new_n672_), .B(u1__abc_73140_new_n668_), .Y(u1__abc_73140_new_n673_));
OR2X2 OR2X2_206 ( .A(u0__abc_76628_new_n1362_), .B(u0__abc_76628_new_n1364_), .Y(u0__abc_76628_new_n1365_));
OR2X2 OR2X2_2060 ( .A(next_adr_bF_buf3), .B(u1_acs_addr_10_), .Y(u1__abc_73140_new_n675_));
OR2X2 OR2X2_2061 ( .A(u1__abc_73140_new_n563__bF_buf1), .B(u1_acs_addr_pl1_10_), .Y(u1__abc_73140_new_n676_));
OR2X2 OR2X2_2062 ( .A(u1__abc_73140_new_n677_), .B(u1__abc_73140_new_n561__bF_buf3), .Y(u1__abc_73140_new_n678_));
OR2X2 OR2X2_2063 ( .A(u1__abc_73140_new_n681_), .B(u1__abc_73140_new_n570__bF_buf1), .Y(u1__abc_73140_new_n682_));
OR2X2 OR2X2_2064 ( .A(u1__abc_73140_new_n682_), .B(u1__abc_73140_new_n680_), .Y(u1__abc_73140_new_n683_));
OR2X2 OR2X2_2065 ( .A(u1__abc_73140_new_n683_), .B(u1__abc_73140_new_n679_), .Y(u1__abc_73140_new_n684_));
OR2X2 OR2X2_2066 ( .A(next_adr_bF_buf2), .B(u1_acs_addr_11_), .Y(u1__abc_73140_new_n686_));
OR2X2 OR2X2_2067 ( .A(u1__abc_73140_new_n563__bF_buf0), .B(u1_acs_addr_pl1_11_), .Y(u1__abc_73140_new_n687_));
OR2X2 OR2X2_2068 ( .A(u1__abc_73140_new_n688_), .B(u1__abc_73140_new_n561__bF_buf2), .Y(u1__abc_73140_new_n689_));
OR2X2 OR2X2_2069 ( .A(u1__abc_73140_new_n692_), .B(u1__abc_73140_new_n570__bF_buf0), .Y(u1__abc_73140_new_n693_));
OR2X2 OR2X2_207 ( .A(u0__abc_76628_new_n1197__bF_buf4), .B(u0_tms0_7_), .Y(u0__abc_76628_new_n1366_));
OR2X2 OR2X2_2070 ( .A(u1__abc_73140_new_n693_), .B(u1__abc_73140_new_n691_), .Y(u1__abc_73140_new_n694_));
OR2X2 OR2X2_2071 ( .A(u1__abc_73140_new_n694_), .B(u1__abc_73140_new_n690_), .Y(u1__abc_73140_new_n695_));
OR2X2 OR2X2_2072 ( .A(next_adr_bF_buf1), .B(u1_acs_addr_12_), .Y(u1__abc_73140_new_n697_));
OR2X2 OR2X2_2073 ( .A(u1__abc_73140_new_n563__bF_buf3), .B(u1_acs_addr_pl1_12_), .Y(u1__abc_73140_new_n698_));
OR2X2 OR2X2_2074 ( .A(u1__abc_73140_new_n699_), .B(u1__abc_73140_new_n561__bF_buf1), .Y(u1__abc_73140_new_n700_));
OR2X2 OR2X2_2075 ( .A(u1__abc_73140_new_n703_), .B(u1__abc_73140_new_n570__bF_buf3), .Y(u1__abc_73140_new_n704_));
OR2X2 OR2X2_2076 ( .A(u1__abc_73140_new_n704_), .B(u1__abc_73140_new_n702_), .Y(u1__abc_73140_new_n705_));
OR2X2 OR2X2_2077 ( .A(u1__abc_73140_new_n705_), .B(u1__abc_73140_new_n701_), .Y(u1__abc_73140_new_n706_));
OR2X2 OR2X2_2078 ( .A(next_adr_bF_buf0), .B(u1_acs_addr_13_), .Y(u1__abc_73140_new_n708_));
OR2X2 OR2X2_2079 ( .A(u1__abc_73140_new_n563__bF_buf2), .B(u1_acs_addr_pl1_13_), .Y(u1__abc_73140_new_n709_));
OR2X2 OR2X2_208 ( .A(u0__abc_76628_new_n1368_), .B(u0__abc_76628_new_n1346_), .Y(u0__0sp_tms_31_0__7_));
OR2X2 OR2X2_2080 ( .A(u1__abc_73140_new_n710_), .B(u1__abc_73140_new_n561__bF_buf0), .Y(u1__abc_73140_new_n711_));
OR2X2 OR2X2_2081 ( .A(u1__abc_73140_new_n714_), .B(u1__abc_73140_new_n570__bF_buf2), .Y(u1__abc_73140_new_n715_));
OR2X2 OR2X2_2082 ( .A(u1__abc_73140_new_n715_), .B(u1__abc_73140_new_n713_), .Y(u1__abc_73140_new_n716_));
OR2X2 OR2X2_2083 ( .A(u1__abc_73140_new_n716_), .B(u1__abc_73140_new_n712_), .Y(u1__abc_73140_new_n717_));
OR2X2 OR2X2_2084 ( .A(next_adr_bF_buf4), .B(u1_acs_addr_14_), .Y(u1__abc_73140_new_n719_));
OR2X2 OR2X2_2085 ( .A(u1__abc_73140_new_n563__bF_buf1), .B(u1_acs_addr_pl1_14_), .Y(u1__abc_73140_new_n720_));
OR2X2 OR2X2_2086 ( .A(u1__abc_73140_new_n721_), .B(u1__abc_73140_new_n561__bF_buf4), .Y(u1__abc_73140_new_n722_));
OR2X2 OR2X2_2087 ( .A(u1__abc_73140_new_n725_), .B(u1__abc_73140_new_n570__bF_buf1), .Y(u1__abc_73140_new_n726_));
OR2X2 OR2X2_2088 ( .A(u1__abc_73140_new_n726_), .B(u1__abc_73140_new_n724_), .Y(u1__abc_73140_new_n727_));
OR2X2 OR2X2_2089 ( .A(u1__abc_73140_new_n727_), .B(u1__abc_73140_new_n723_), .Y(u1__abc_73140_new_n728_));
OR2X2 OR2X2_209 ( .A(u0__abc_76628_new_n1177__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n1372_));
OR2X2 OR2X2_2090 ( .A(next_adr_bF_buf3), .B(u1_acs_addr_15_), .Y(u1__abc_73140_new_n730_));
OR2X2 OR2X2_2091 ( .A(u1__abc_73140_new_n563__bF_buf0), .B(u1_acs_addr_pl1_15_), .Y(u1__abc_73140_new_n731_));
OR2X2 OR2X2_2092 ( .A(u1__abc_73140_new_n732_), .B(u1__abc_73140_new_n561__bF_buf3), .Y(u1__abc_73140_new_n733_));
OR2X2 OR2X2_2093 ( .A(u1__abc_73140_new_n736_), .B(u1__abc_73140_new_n570__bF_buf0), .Y(u1__abc_73140_new_n737_));
OR2X2 OR2X2_2094 ( .A(u1__abc_73140_new_n737_), .B(u1__abc_73140_new_n735_), .Y(u1__abc_73140_new_n738_));
OR2X2 OR2X2_2095 ( .A(u1__abc_73140_new_n738_), .B(u1__abc_73140_new_n734_), .Y(u1__abc_73140_new_n739_));
OR2X2 OR2X2_2096 ( .A(next_adr_bF_buf2), .B(u1_acs_addr_16_), .Y(u1__abc_73140_new_n741_));
OR2X2 OR2X2_2097 ( .A(u1__abc_73140_new_n563__bF_buf3), .B(u1_acs_addr_pl1_16_), .Y(u1__abc_73140_new_n742_));
OR2X2 OR2X2_2098 ( .A(u1__abc_73140_new_n743_), .B(u1__abc_73140_new_n561__bF_buf2), .Y(u1__abc_73140_new_n744_));
OR2X2 OR2X2_2099 ( .A(u1__abc_73140_new_n747_), .B(u1__abc_73140_new_n570__bF_buf3), .Y(u1__abc_73140_new_n748_));
OR2X2 OR2X2_21 ( .A(_abc_85006_new_n268_), .B(_abc_85006_new_n237_), .Y(_abc_85006_new_n269_));
OR2X2 OR2X2_210 ( .A(spec_req_cs_6_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1373_));
OR2X2 OR2X2_2100 ( .A(u1__abc_73140_new_n748_), .B(u1__abc_73140_new_n746_), .Y(u1__abc_73140_new_n749_));
OR2X2 OR2X2_2101 ( .A(u1__abc_73140_new_n749_), .B(u1__abc_73140_new_n745_), .Y(u1__abc_73140_new_n750_));
OR2X2 OR2X2_2102 ( .A(next_adr_bF_buf1), .B(u1_acs_addr_17_), .Y(u1__abc_73140_new_n752_));
OR2X2 OR2X2_2103 ( .A(u1__abc_73140_new_n563__bF_buf2), .B(u1_acs_addr_pl1_17_), .Y(u1__abc_73140_new_n753_));
OR2X2 OR2X2_2104 ( .A(u1__abc_73140_new_n754_), .B(u1__abc_73140_new_n561__bF_buf1), .Y(u1__abc_73140_new_n755_));
OR2X2 OR2X2_2105 ( .A(u1__abc_73140_new_n758_), .B(u1__abc_73140_new_n570__bF_buf2), .Y(u1__abc_73140_new_n759_));
OR2X2 OR2X2_2106 ( .A(u1__abc_73140_new_n759_), .B(u1__abc_73140_new_n757_), .Y(u1__abc_73140_new_n760_));
OR2X2 OR2X2_2107 ( .A(u1__abc_73140_new_n760_), .B(u1__abc_73140_new_n756_), .Y(u1__abc_73140_new_n761_));
OR2X2 OR2X2_2108 ( .A(next_adr_bF_buf0), .B(u1_acs_addr_18_), .Y(u1__abc_73140_new_n763_));
OR2X2 OR2X2_2109 ( .A(u1__abc_73140_new_n563__bF_buf1), .B(u1_acs_addr_pl1_18_), .Y(u1__abc_73140_new_n764_));
OR2X2 OR2X2_211 ( .A(u0__abc_76628_new_n1375_), .B(u0__abc_76628_new_n1371_), .Y(u0__abc_76628_new_n1376_));
OR2X2 OR2X2_2110 ( .A(u1__abc_73140_new_n765_), .B(u1__abc_73140_new_n561__bF_buf0), .Y(u1__abc_73140_new_n766_));
OR2X2 OR2X2_2111 ( .A(u1__abc_73140_new_n769_), .B(u1__abc_73140_new_n570__bF_buf1), .Y(u1__abc_73140_new_n770_));
OR2X2 OR2X2_2112 ( .A(u1__abc_73140_new_n770_), .B(u1__abc_73140_new_n768_), .Y(u1__abc_73140_new_n771_));
OR2X2 OR2X2_2113 ( .A(u1__abc_73140_new_n771_), .B(u1__abc_73140_new_n767_), .Y(u1__abc_73140_new_n772_));
OR2X2 OR2X2_2114 ( .A(next_adr_bF_buf4), .B(u1_acs_addr_19_), .Y(u1__abc_73140_new_n774_));
OR2X2 OR2X2_2115 ( .A(u1__abc_73140_new_n563__bF_buf0), .B(u1_acs_addr_pl1_19_), .Y(u1__abc_73140_new_n775_));
OR2X2 OR2X2_2116 ( .A(u1__abc_73140_new_n776_), .B(u1__abc_73140_new_n561__bF_buf4), .Y(u1__abc_73140_new_n777_));
OR2X2 OR2X2_2117 ( .A(u1__abc_73140_new_n779_), .B(u1__abc_73140_new_n570__bF_buf0), .Y(u1__abc_73140_new_n780_));
OR2X2 OR2X2_2118 ( .A(u1__abc_73140_new_n780_), .B(u1__abc_73140_new_n315_), .Y(u1__abc_73140_new_n781_));
OR2X2 OR2X2_2119 ( .A(u1__abc_73140_new_n781_), .B(u1__abc_73140_new_n778_), .Y(u1__abc_73140_new_n782_));
OR2X2 OR2X2_212 ( .A(u0__abc_76628_new_n1377_), .B(u0__abc_76628_new_n1378_), .Y(u0__abc_76628_new_n1379_));
OR2X2 OR2X2_2120 ( .A(next_adr_bF_buf3), .B(u1_acs_addr_20_), .Y(u1__abc_73140_new_n784_));
OR2X2 OR2X2_2121 ( .A(u1__abc_73140_new_n563__bF_buf3), .B(u1_acs_addr_pl1_20_), .Y(u1__abc_73140_new_n785_));
OR2X2 OR2X2_2122 ( .A(u1__abc_73140_new_n786_), .B(u1__abc_73140_new_n561__bF_buf3), .Y(u1__abc_73140_new_n787_));
OR2X2 OR2X2_2123 ( .A(u1__abc_73140_new_n789_), .B(u1__abc_73140_new_n570__bF_buf3), .Y(u1__abc_73140_new_n790_));
OR2X2 OR2X2_2124 ( .A(u1__abc_73140_new_n790_), .B(u1__abc_73140_new_n336_), .Y(u1__abc_73140_new_n791_));
OR2X2 OR2X2_2125 ( .A(u1__abc_73140_new_n791_), .B(u1__abc_73140_new_n788_), .Y(u1__abc_73140_new_n792_));
OR2X2 OR2X2_2126 ( .A(next_adr_bF_buf2), .B(u1_acs_addr_21_), .Y(u1__abc_73140_new_n794_));
OR2X2 OR2X2_2127 ( .A(u1__abc_73140_new_n563__bF_buf2), .B(u1_acs_addr_pl1_21_), .Y(u1__abc_73140_new_n795_));
OR2X2 OR2X2_2128 ( .A(u1__abc_73140_new_n796_), .B(u1__abc_73140_new_n561__bF_buf2), .Y(u1__abc_73140_new_n797_));
OR2X2 OR2X2_2129 ( .A(u1__abc_73140_new_n800_), .B(u1__abc_73140_new_n570__bF_buf2), .Y(u1__abc_73140_new_n801_));
OR2X2 OR2X2_213 ( .A(u0__abc_76628_new_n1380_), .B(u0__abc_76628_new_n1381_), .Y(u0__abc_76628_new_n1382_));
OR2X2 OR2X2_2130 ( .A(u1__abc_73140_new_n801_), .B(u1__abc_73140_new_n799_), .Y(u1__abc_73140_new_n802_));
OR2X2 OR2X2_2131 ( .A(u1__abc_73140_new_n802_), .B(u1__abc_73140_new_n798_), .Y(u1__abc_73140_new_n803_));
OR2X2 OR2X2_2132 ( .A(next_adr_bF_buf1), .B(u1_acs_addr_22_), .Y(u1__abc_73140_new_n805_));
OR2X2 OR2X2_2133 ( .A(u1__abc_73140_new_n563__bF_buf1), .B(u1_acs_addr_pl1_22_), .Y(u1__abc_73140_new_n806_));
OR2X2 OR2X2_2134 ( .A(u1__abc_73140_new_n807_), .B(u1__abc_73140_new_n561__bF_buf1), .Y(u1__abc_73140_new_n808_));
OR2X2 OR2X2_2135 ( .A(u1__abc_73140_new_n487_), .B(u1__abc_73140_new_n570__bF_buf1), .Y(u1__abc_73140_new_n810_));
OR2X2 OR2X2_2136 ( .A(u1__abc_73140_new_n810_), .B(u1__abc_73140_new_n514_), .Y(u1__abc_73140_new_n811_));
OR2X2 OR2X2_2137 ( .A(u1__abc_73140_new_n811_), .B(u1__abc_73140_new_n809_), .Y(u1__abc_73140_new_n812_));
OR2X2 OR2X2_2138 ( .A(next_adr_bF_buf0), .B(u1_acs_addr_23_), .Y(u1__abc_73140_new_n814_));
OR2X2 OR2X2_2139 ( .A(u1__abc_73140_new_n563__bF_buf0), .B(u1_acs_addr_pl1_23_), .Y(u1__abc_73140_new_n815_));
OR2X2 OR2X2_214 ( .A(u0__abc_76628_new_n1383_), .B(u0__abc_76628_new_n1384_), .Y(u0__abc_76628_new_n1385_));
OR2X2 OR2X2_2140 ( .A(u1__abc_73140_new_n816_), .B(u1__abc_73140_new_n561__bF_buf0), .Y(u1__abc_73140_new_n817_));
OR2X2 OR2X2_2141 ( .A(u1__abc_73140_new_n820_), .B(u1__abc_73140_new_n570__bF_buf0), .Y(u1__abc_73140_new_n821_));
OR2X2 OR2X2_2142 ( .A(u1__abc_73140_new_n821_), .B(u1__abc_73140_new_n819_), .Y(u1__abc_73140_new_n822_));
OR2X2 OR2X2_2143 ( .A(u1__abc_73140_new_n822_), .B(u1__abc_73140_new_n818_), .Y(u1__abc_73140_new_n823_));
OR2X2 OR2X2_2144 ( .A(wb_stb_i_bF_buf2), .B(u1_sram_addr_0_), .Y(u1__abc_73140_new_n825_));
OR2X2 OR2X2_2145 ( .A(u1__abc_73140_new_n826__bF_buf3), .B(\wb_addr_i[2] ), .Y(u1__abc_73140_new_n827_));
OR2X2 OR2X2_2146 ( .A(wb_stb_i_bF_buf0), .B(u1_sram_addr_1_), .Y(u1__abc_73140_new_n829_));
OR2X2 OR2X2_2147 ( .A(u1__abc_73140_new_n826__bF_buf2), .B(\wb_addr_i[3] ), .Y(u1__abc_73140_new_n830_));
OR2X2 OR2X2_2148 ( .A(wb_stb_i_bF_buf5), .B(u1_sram_addr_2_), .Y(u1__abc_73140_new_n832_));
OR2X2 OR2X2_2149 ( .A(u1__abc_73140_new_n826__bF_buf1), .B(\wb_addr_i[4] ), .Y(u1__abc_73140_new_n833_));
OR2X2 OR2X2_215 ( .A(u0__abc_76628_new_n1387_), .B(spec_req_cs_0_bF_buf0_), .Y(u0__abc_76628_new_n1388_));
OR2X2 OR2X2_2150 ( .A(wb_stb_i_bF_buf4), .B(u1_sram_addr_3_), .Y(u1__abc_73140_new_n835_));
OR2X2 OR2X2_2151 ( .A(u1__abc_73140_new_n826__bF_buf0), .B(\wb_addr_i[5] ), .Y(u1__abc_73140_new_n836_));
OR2X2 OR2X2_2152 ( .A(wb_stb_i_bF_buf3), .B(u1_sram_addr_4_), .Y(u1__abc_73140_new_n838_));
OR2X2 OR2X2_2153 ( .A(u1__abc_73140_new_n826__bF_buf3), .B(\wb_addr_i[6] ), .Y(u1__abc_73140_new_n839_));
OR2X2 OR2X2_2154 ( .A(wb_stb_i_bF_buf2), .B(u1_sram_addr_5_), .Y(u1__abc_73140_new_n841_));
OR2X2 OR2X2_2155 ( .A(u1__abc_73140_new_n826__bF_buf2), .B(\wb_addr_i[7] ), .Y(u1__abc_73140_new_n842_));
OR2X2 OR2X2_2156 ( .A(wb_stb_i_bF_buf1), .B(u1_sram_addr_6_), .Y(u1__abc_73140_new_n844_));
OR2X2 OR2X2_2157 ( .A(u1__abc_73140_new_n826__bF_buf1), .B(\wb_addr_i[8] ), .Y(u1__abc_73140_new_n845_));
OR2X2 OR2X2_2158 ( .A(wb_stb_i_bF_buf0), .B(u1_sram_addr_7_), .Y(u1__abc_73140_new_n847_));
OR2X2 OR2X2_2159 ( .A(u1__abc_73140_new_n826__bF_buf0), .B(\wb_addr_i[9] ), .Y(u1__abc_73140_new_n848_));
OR2X2 OR2X2_216 ( .A(u0__abc_76628_new_n1386_), .B(u0__abc_76628_new_n1388_), .Y(u0__abc_76628_new_n1389_));
OR2X2 OR2X2_2160 ( .A(wb_stb_i_bF_buf5), .B(u1_sram_addr_8_), .Y(u1__abc_73140_new_n850_));
OR2X2 OR2X2_2161 ( .A(u1__abc_73140_new_n826__bF_buf3), .B(\wb_addr_i[10] ), .Y(u1__abc_73140_new_n851_));
OR2X2 OR2X2_2162 ( .A(wb_stb_i_bF_buf4), .B(u1_sram_addr_9_), .Y(u1__abc_73140_new_n853_));
OR2X2 OR2X2_2163 ( .A(u1__abc_73140_new_n826__bF_buf2), .B(\wb_addr_i[11] ), .Y(u1__abc_73140_new_n854_));
OR2X2 OR2X2_2164 ( .A(wb_stb_i_bF_buf3), .B(u1_sram_addr_10_), .Y(u1__abc_73140_new_n856_));
OR2X2 OR2X2_2165 ( .A(u1__abc_73140_new_n826__bF_buf1), .B(\wb_addr_i[12] ), .Y(u1__abc_73140_new_n857_));
OR2X2 OR2X2_2166 ( .A(wb_stb_i_bF_buf2), .B(u1_sram_addr_11_), .Y(u1__abc_73140_new_n859_));
OR2X2 OR2X2_2167 ( .A(u1__abc_73140_new_n826__bF_buf0), .B(\wb_addr_i[13] ), .Y(u1__abc_73140_new_n860_));
OR2X2 OR2X2_2168 ( .A(wb_stb_i_bF_buf1), .B(u1_sram_addr_12_), .Y(u1__abc_73140_new_n862_));
OR2X2 OR2X2_2169 ( .A(u1__abc_73140_new_n826__bF_buf3), .B(\wb_addr_i[14] ), .Y(u1__abc_73140_new_n863_));
OR2X2 OR2X2_217 ( .A(u0__abc_76628_new_n1197__bF_buf3), .B(u0_tms0_8_), .Y(u0__abc_76628_new_n1390_));
OR2X2 OR2X2_2170 ( .A(wb_stb_i_bF_buf0), .B(u1_sram_addr_13_), .Y(u1__abc_73140_new_n865_));
OR2X2 OR2X2_2171 ( .A(u1__abc_73140_new_n826__bF_buf2), .B(\wb_addr_i[15] ), .Y(u1__abc_73140_new_n866_));
OR2X2 OR2X2_2172 ( .A(wb_stb_i_bF_buf5), .B(u1_sram_addr_14_), .Y(u1__abc_73140_new_n868_));
OR2X2 OR2X2_2173 ( .A(u1__abc_73140_new_n826__bF_buf1), .B(\wb_addr_i[16] ), .Y(u1__abc_73140_new_n869_));
OR2X2 OR2X2_2174 ( .A(wb_stb_i_bF_buf4), .B(u1_sram_addr_15_), .Y(u1__abc_73140_new_n871_));
OR2X2 OR2X2_2175 ( .A(u1__abc_73140_new_n826__bF_buf0), .B(\wb_addr_i[17] ), .Y(u1__abc_73140_new_n872_));
OR2X2 OR2X2_2176 ( .A(wb_stb_i_bF_buf3), .B(u1_sram_addr_16_), .Y(u1__abc_73140_new_n874_));
OR2X2 OR2X2_2177 ( .A(u1__abc_73140_new_n826__bF_buf3), .B(\wb_addr_i[18] ), .Y(u1__abc_73140_new_n875_));
OR2X2 OR2X2_2178 ( .A(wb_stb_i_bF_buf2), .B(u1_sram_addr_17_), .Y(u1__abc_73140_new_n877_));
OR2X2 OR2X2_2179 ( .A(u1__abc_73140_new_n826__bF_buf2), .B(\wb_addr_i[19] ), .Y(u1__abc_73140_new_n878_));
OR2X2 OR2X2_218 ( .A(u0__abc_76628_new_n1392_), .B(u0__abc_76628_new_n1370_), .Y(u0__0sp_tms_31_0__8_));
OR2X2 OR2X2_2180 ( .A(wb_stb_i_bF_buf1), .B(u1_sram_addr_18_), .Y(u1__abc_73140_new_n880_));
OR2X2 OR2X2_2181 ( .A(u1__abc_73140_new_n826__bF_buf1), .B(\wb_addr_i[20] ), .Y(u1__abc_73140_new_n881_));
OR2X2 OR2X2_2182 ( .A(wb_stb_i_bF_buf0), .B(u1_sram_addr_19_), .Y(u1__abc_73140_new_n883_));
OR2X2 OR2X2_2183 ( .A(u1__abc_73140_new_n826__bF_buf0), .B(\wb_addr_i[21] ), .Y(u1__abc_73140_new_n884_));
OR2X2 OR2X2_2184 ( .A(wb_stb_i_bF_buf5), .B(u1_sram_addr_20_), .Y(u1__abc_73140_new_n886_));
OR2X2 OR2X2_2185 ( .A(u1__abc_73140_new_n826__bF_buf3), .B(\wb_addr_i[22] ), .Y(u1__abc_73140_new_n887_));
OR2X2 OR2X2_2186 ( .A(wb_stb_i_bF_buf4), .B(u1_sram_addr_21_), .Y(u1__abc_73140_new_n889_));
OR2X2 OR2X2_2187 ( .A(u1__abc_73140_new_n826__bF_buf2), .B(\wb_addr_i[23] ), .Y(u1__abc_73140_new_n890_));
OR2X2 OR2X2_2188 ( .A(wb_stb_i_bF_buf3), .B(u1_sram_addr_22_), .Y(u1__abc_73140_new_n892_));
OR2X2 OR2X2_2189 ( .A(u1__abc_73140_new_n826__bF_buf1), .B(\wb_addr_i[24] ), .Y(u1__abc_73140_new_n893_));
OR2X2 OR2X2_219 ( .A(u0__abc_76628_new_n1177__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n1396_));
OR2X2 OR2X2_2190 ( .A(wb_stb_i_bF_buf2), .B(u1_sram_addr_23_), .Y(u1__abc_73140_new_n895_));
OR2X2 OR2X2_2191 ( .A(u1__abc_73140_new_n826__bF_buf0), .B(\wb_addr_i[25] ), .Y(u1__abc_73140_new_n896_));
OR2X2 OR2X2_2192 ( .A(csc_s_3_), .B(csc_s_1_), .Y(u1__abc_73140_new_n898_));
OR2X2 OR2X2_2193 ( .A(csc_s_3_), .B(csc_s_2_), .Y(u1__abc_73140_new_n901_));
OR2X2 OR2X2_2194 ( .A(u1__abc_73140_new_n904__bF_buf4), .B(\wb_addr_i[2] ), .Y(u1__abc_73140_new_n905_));
OR2X2 OR2X2_2195 ( .A(u1__abc_73140_new_n906__bF_buf3), .B(u1_sram_addr_0_), .Y(u1__abc_73140_new_n907_));
OR2X2 OR2X2_2196 ( .A(u1__abc_73140_new_n908_), .B(u1__abc_73140_new_n900__bF_buf4), .Y(u1__abc_73140_new_n909_));
OR2X2 OR2X2_2197 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_0_), .Y(u1__abc_73140_new_n914_));
OR2X2 OR2X2_2198 ( .A(u1__abc_73140_new_n919_), .B(tms_s_0_), .Y(u1__abc_73140_new_n920_));
OR2X2 OR2X2_2199 ( .A(u1__abc_73140_new_n921_), .B(row_adr_0_bF_buf2_), .Y(u1__abc_73140_new_n922_));
OR2X2 OR2X2_22 ( .A(_abc_85006_new_n245_), .B(cs_need_rfr_4_), .Y(_abc_85006_new_n270_));
OR2X2 OR2X2_220 ( .A(spec_req_cs_6_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1397_));
OR2X2 OR2X2_2200 ( .A(u1_col_adr_0_), .B(row_sel), .Y(u1__abc_73140_new_n923_));
OR2X2 OR2X2_2201 ( .A(u1__abc_73140_new_n924_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n925_));
OR2X2 OR2X2_2202 ( .A(u1__abc_73140_new_n916_), .B(u1__abc_73140_new_n927_), .Y(mc_addr_d_0_));
OR2X2 OR2X2_2203 ( .A(u1__abc_73140_new_n904__bF_buf2), .B(\wb_addr_i[3] ), .Y(u1__abc_73140_new_n929_));
OR2X2 OR2X2_2204 ( .A(u1__abc_73140_new_n906__bF_buf2), .B(u1_sram_addr_1_), .Y(u1__abc_73140_new_n930_));
OR2X2 OR2X2_2205 ( .A(u1__abc_73140_new_n931_), .B(u1__abc_73140_new_n900__bF_buf2), .Y(u1__abc_73140_new_n932_));
OR2X2 OR2X2_2206 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_1_), .Y(u1__abc_73140_new_n933_));
OR2X2 OR2X2_2207 ( .A(u1__abc_73140_new_n919_), .B(tms_s_1_), .Y(u1__abc_73140_new_n936_));
OR2X2 OR2X2_2208 ( .A(u1__abc_73140_new_n921_), .B(row_adr_1_bF_buf2_), .Y(u1__abc_73140_new_n937_));
OR2X2 OR2X2_2209 ( .A(u1_col_adr_1_), .B(row_sel), .Y(u1__abc_73140_new_n938_));
OR2X2 OR2X2_221 ( .A(u0__abc_76628_new_n1399_), .B(u0__abc_76628_new_n1395_), .Y(u0__abc_76628_new_n1400_));
OR2X2 OR2X2_2210 ( .A(u1__abc_73140_new_n939_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n940_));
OR2X2 OR2X2_2211 ( .A(u1__abc_73140_new_n935_), .B(u1__abc_73140_new_n942_), .Y(mc_addr_d_1_));
OR2X2 OR2X2_2212 ( .A(u1__abc_73140_new_n904__bF_buf1), .B(\wb_addr_i[4] ), .Y(u1__abc_73140_new_n944_));
OR2X2 OR2X2_2213 ( .A(u1__abc_73140_new_n906__bF_buf1), .B(u1_sram_addr_2_), .Y(u1__abc_73140_new_n945_));
OR2X2 OR2X2_2214 ( .A(u1__abc_73140_new_n946_), .B(u1__abc_73140_new_n900__bF_buf1), .Y(u1__abc_73140_new_n947_));
OR2X2 OR2X2_2215 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_2_), .Y(u1__abc_73140_new_n948_));
OR2X2 OR2X2_2216 ( .A(u1__abc_73140_new_n919_), .B(tms_s_2_), .Y(u1__abc_73140_new_n951_));
OR2X2 OR2X2_2217 ( .A(u1__abc_73140_new_n921_), .B(row_adr_2_bF_buf2_), .Y(u1__abc_73140_new_n952_));
OR2X2 OR2X2_2218 ( .A(u1_col_adr_2_), .B(row_sel), .Y(u1__abc_73140_new_n953_));
OR2X2 OR2X2_2219 ( .A(u1__abc_73140_new_n954_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n955_));
OR2X2 OR2X2_222 ( .A(u0__abc_76628_new_n1401_), .B(u0__abc_76628_new_n1402_), .Y(u0__abc_76628_new_n1403_));
OR2X2 OR2X2_2220 ( .A(u1__abc_73140_new_n950_), .B(u1__abc_73140_new_n957_), .Y(mc_addr_d_2_));
OR2X2 OR2X2_2221 ( .A(u1__abc_73140_new_n904__bF_buf0), .B(\wb_addr_i[5] ), .Y(u1__abc_73140_new_n959_));
OR2X2 OR2X2_2222 ( .A(u1__abc_73140_new_n906__bF_buf0), .B(u1_sram_addr_3_), .Y(u1__abc_73140_new_n960_));
OR2X2 OR2X2_2223 ( .A(u1__abc_73140_new_n961_), .B(u1__abc_73140_new_n900__bF_buf0), .Y(u1__abc_73140_new_n962_));
OR2X2 OR2X2_2224 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_3_), .Y(u1__abc_73140_new_n963_));
OR2X2 OR2X2_2225 ( .A(u1__abc_73140_new_n919_), .B(tms_s_3_), .Y(u1__abc_73140_new_n966_));
OR2X2 OR2X2_2226 ( .A(u1__abc_73140_new_n921_), .B(row_adr_3_bF_buf2_), .Y(u1__abc_73140_new_n967_));
OR2X2 OR2X2_2227 ( .A(u1_col_adr_3_), .B(row_sel), .Y(u1__abc_73140_new_n968_));
OR2X2 OR2X2_2228 ( .A(u1__abc_73140_new_n969_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n970_));
OR2X2 OR2X2_2229 ( .A(u1__abc_73140_new_n965_), .B(u1__abc_73140_new_n972_), .Y(mc_addr_d_3_));
OR2X2 OR2X2_223 ( .A(u0__abc_76628_new_n1404_), .B(u0__abc_76628_new_n1405_), .Y(u0__abc_76628_new_n1406_));
OR2X2 OR2X2_2230 ( .A(u1__abc_73140_new_n904__bF_buf4), .B(\wb_addr_i[6] ), .Y(u1__abc_73140_new_n974_));
OR2X2 OR2X2_2231 ( .A(u1__abc_73140_new_n906__bF_buf3), .B(u1_sram_addr_4_), .Y(u1__abc_73140_new_n975_));
OR2X2 OR2X2_2232 ( .A(u1__abc_73140_new_n976_), .B(u1__abc_73140_new_n900__bF_buf4), .Y(u1__abc_73140_new_n977_));
OR2X2 OR2X2_2233 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_4_), .Y(u1__abc_73140_new_n978_));
OR2X2 OR2X2_2234 ( .A(u1__abc_73140_new_n919_), .B(tms_s_4_), .Y(u1__abc_73140_new_n981_));
OR2X2 OR2X2_2235 ( .A(u1__abc_73140_new_n921_), .B(row_adr_4_bF_buf2_), .Y(u1__abc_73140_new_n982_));
OR2X2 OR2X2_2236 ( .A(u1_col_adr_4_), .B(row_sel), .Y(u1__abc_73140_new_n983_));
OR2X2 OR2X2_2237 ( .A(u1__abc_73140_new_n984_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n985_));
OR2X2 OR2X2_2238 ( .A(u1__abc_73140_new_n980_), .B(u1__abc_73140_new_n987_), .Y(mc_addr_d_4_));
OR2X2 OR2X2_2239 ( .A(u1__abc_73140_new_n904__bF_buf3), .B(\wb_addr_i[7] ), .Y(u1__abc_73140_new_n989_));
OR2X2 OR2X2_224 ( .A(u0__abc_76628_new_n1407_), .B(u0__abc_76628_new_n1408_), .Y(u0__abc_76628_new_n1409_));
OR2X2 OR2X2_2240 ( .A(u1__abc_73140_new_n906__bF_buf2), .B(u1_sram_addr_5_), .Y(u1__abc_73140_new_n990_));
OR2X2 OR2X2_2241 ( .A(u1__abc_73140_new_n991_), .B(u1__abc_73140_new_n900__bF_buf3), .Y(u1__abc_73140_new_n992_));
OR2X2 OR2X2_2242 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_5_), .Y(u1__abc_73140_new_n993_));
OR2X2 OR2X2_2243 ( .A(u1__abc_73140_new_n919_), .B(tms_s_5_), .Y(u1__abc_73140_new_n996_));
OR2X2 OR2X2_2244 ( .A(u1__abc_73140_new_n921_), .B(row_adr_5_bF_buf2_), .Y(u1__abc_73140_new_n997_));
OR2X2 OR2X2_2245 ( .A(u1_col_adr_5_), .B(row_sel), .Y(u1__abc_73140_new_n998_));
OR2X2 OR2X2_2246 ( .A(u1__abc_73140_new_n999_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n1000_));
OR2X2 OR2X2_2247 ( .A(u1__abc_73140_new_n995_), .B(u1__abc_73140_new_n1002_), .Y(mc_addr_d_5_));
OR2X2 OR2X2_2248 ( .A(u1__abc_73140_new_n904__bF_buf2), .B(\wb_addr_i[8] ), .Y(u1__abc_73140_new_n1004_));
OR2X2 OR2X2_2249 ( .A(u1__abc_73140_new_n906__bF_buf1), .B(u1_sram_addr_6_), .Y(u1__abc_73140_new_n1005_));
OR2X2 OR2X2_225 ( .A(u0__abc_76628_new_n1411_), .B(spec_req_cs_0_bF_buf5_), .Y(u0__abc_76628_new_n1412_));
OR2X2 OR2X2_2250 ( .A(u1__abc_73140_new_n1006_), .B(u1__abc_73140_new_n900__bF_buf2), .Y(u1__abc_73140_new_n1007_));
OR2X2 OR2X2_2251 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_6_), .Y(u1__abc_73140_new_n1008_));
OR2X2 OR2X2_2252 ( .A(u1__abc_73140_new_n919_), .B(tms_s_6_), .Y(u1__abc_73140_new_n1011_));
OR2X2 OR2X2_2253 ( .A(u1__abc_73140_new_n921_), .B(row_adr_6_bF_buf2_), .Y(u1__abc_73140_new_n1012_));
OR2X2 OR2X2_2254 ( .A(u1_col_adr_6_), .B(row_sel), .Y(u1__abc_73140_new_n1013_));
OR2X2 OR2X2_2255 ( .A(u1__abc_73140_new_n1014_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n1015_));
OR2X2 OR2X2_2256 ( .A(u1__abc_73140_new_n1010_), .B(u1__abc_73140_new_n1017_), .Y(mc_addr_d_6_));
OR2X2 OR2X2_2257 ( .A(u1__abc_73140_new_n904__bF_buf1), .B(\wb_addr_i[9] ), .Y(u1__abc_73140_new_n1019_));
OR2X2 OR2X2_2258 ( .A(u1__abc_73140_new_n906__bF_buf0), .B(u1_sram_addr_7_), .Y(u1__abc_73140_new_n1020_));
OR2X2 OR2X2_2259 ( .A(u1__abc_73140_new_n1021_), .B(u1__abc_73140_new_n900__bF_buf1), .Y(u1__abc_73140_new_n1022_));
OR2X2 OR2X2_226 ( .A(u0__abc_76628_new_n1410_), .B(u0__abc_76628_new_n1412_), .Y(u0__abc_76628_new_n1413_));
OR2X2 OR2X2_2260 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_7_), .Y(u1__abc_73140_new_n1023_));
OR2X2 OR2X2_2261 ( .A(u1__abc_73140_new_n919_), .B(tms_s_7_), .Y(u1__abc_73140_new_n1026_));
OR2X2 OR2X2_2262 ( .A(u1__abc_73140_new_n921_), .B(row_adr_7_bF_buf2_), .Y(u1__abc_73140_new_n1027_));
OR2X2 OR2X2_2263 ( .A(u1_col_adr_7_), .B(row_sel), .Y(u1__abc_73140_new_n1028_));
OR2X2 OR2X2_2264 ( .A(u1__abc_73140_new_n1029_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n1030_));
OR2X2 OR2X2_2265 ( .A(u1__abc_73140_new_n1025_), .B(u1__abc_73140_new_n1032_), .Y(mc_addr_d_7_));
OR2X2 OR2X2_2266 ( .A(u1__abc_73140_new_n904__bF_buf0), .B(\wb_addr_i[10] ), .Y(u1__abc_73140_new_n1034_));
OR2X2 OR2X2_2267 ( .A(u1__abc_73140_new_n906__bF_buf3), .B(u1_sram_addr_8_), .Y(u1__abc_73140_new_n1035_));
OR2X2 OR2X2_2268 ( .A(u1__abc_73140_new_n1036_), .B(u1__abc_73140_new_n900__bF_buf0), .Y(u1__abc_73140_new_n1037_));
OR2X2 OR2X2_2269 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_8_), .Y(u1__abc_73140_new_n1038_));
OR2X2 OR2X2_227 ( .A(u0__abc_76628_new_n1197__bF_buf2), .B(u0_tms0_9_), .Y(u0__abc_76628_new_n1414_));
OR2X2 OR2X2_2270 ( .A(u1__abc_73140_new_n919_), .B(tms_s_8_), .Y(u1__abc_73140_new_n1041_));
OR2X2 OR2X2_2271 ( .A(u1__abc_73140_new_n921_), .B(row_adr_8_bF_buf2_), .Y(u1__abc_73140_new_n1042_));
OR2X2 OR2X2_2272 ( .A(u1_col_adr_8_), .B(row_sel), .Y(u1__abc_73140_new_n1043_));
OR2X2 OR2X2_2273 ( .A(u1__abc_73140_new_n1044_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n1045_));
OR2X2 OR2X2_2274 ( .A(u1__abc_73140_new_n1040_), .B(u1__abc_73140_new_n1047_), .Y(mc_addr_d_8_));
OR2X2 OR2X2_2275 ( .A(u1__abc_73140_new_n904__bF_buf4), .B(\wb_addr_i[11] ), .Y(u1__abc_73140_new_n1049_));
OR2X2 OR2X2_2276 ( .A(u1__abc_73140_new_n906__bF_buf2), .B(u1_sram_addr_9_), .Y(u1__abc_73140_new_n1050_));
OR2X2 OR2X2_2277 ( .A(u1__abc_73140_new_n1051_), .B(u1__abc_73140_new_n900__bF_buf4), .Y(u1__abc_73140_new_n1052_));
OR2X2 OR2X2_2278 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_9_), .Y(u1__abc_73140_new_n1053_));
OR2X2 OR2X2_2279 ( .A(u1__abc_73140_new_n919_), .B(tms_s_9_), .Y(u1__abc_73140_new_n1056_));
OR2X2 OR2X2_228 ( .A(u0__abc_76628_new_n1416_), .B(u0__abc_76628_new_n1394_), .Y(u0__0sp_tms_31_0__9_));
OR2X2 OR2X2_2280 ( .A(u1__abc_73140_new_n921_), .B(row_adr_9_bF_buf2_), .Y(u1__abc_73140_new_n1057_));
OR2X2 OR2X2_2281 ( .A(u1_col_adr_9_), .B(row_sel), .Y(u1__abc_73140_new_n1058_));
OR2X2 OR2X2_2282 ( .A(u1__abc_73140_new_n1059_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n1060_));
OR2X2 OR2X2_2283 ( .A(u1__abc_73140_new_n1055_), .B(u1__abc_73140_new_n1062_), .Y(mc_addr_d_9_));
OR2X2 OR2X2_2284 ( .A(u1__abc_73140_new_n904__bF_buf3), .B(\wb_addr_i[13] ), .Y(u1__abc_73140_new_n1064_));
OR2X2 OR2X2_2285 ( .A(u1__abc_73140_new_n906__bF_buf1), .B(u1_sram_addr_11_), .Y(u1__abc_73140_new_n1065_));
OR2X2 OR2X2_2286 ( .A(u1__abc_73140_new_n1066_), .B(u1__abc_73140_new_n900__bF_buf3), .Y(u1__abc_73140_new_n1067_));
OR2X2 OR2X2_2287 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_11_), .Y(u1__abc_73140_new_n1068_));
OR2X2 OR2X2_2288 ( .A(u1__abc_73140_new_n919_), .B(tms_s_11_), .Y(u1__abc_73140_new_n1071_));
OR2X2 OR2X2_2289 ( .A(u1__abc_73140_new_n918_), .B(u1__abc_73140_new_n1072_), .Y(u1__abc_73140_new_n1073_));
OR2X2 OR2X2_229 ( .A(u0__abc_76628_new_n1177__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n1420_));
OR2X2 OR2X2_2290 ( .A(u1__abc_73140_new_n1070_), .B(u1__abc_73140_new_n1075_), .Y(mc_addr_d_11_));
OR2X2 OR2X2_2291 ( .A(u1__abc_73140_new_n904__bF_buf2), .B(\wb_addr_i[14] ), .Y(u1__abc_73140_new_n1077_));
OR2X2 OR2X2_2292 ( .A(u1__abc_73140_new_n906__bF_buf0), .B(u1_sram_addr_12_), .Y(u1__abc_73140_new_n1078_));
OR2X2 OR2X2_2293 ( .A(u1__abc_73140_new_n1079_), .B(u1__abc_73140_new_n900__bF_buf2), .Y(u1__abc_73140_new_n1080_));
OR2X2 OR2X2_2294 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_12_), .Y(u1__abc_73140_new_n1081_));
OR2X2 OR2X2_2295 ( .A(u1__abc_73140_new_n919_), .B(tms_s_12_), .Y(u1__abc_73140_new_n1084_));
OR2X2 OR2X2_2296 ( .A(u1__abc_73140_new_n918_), .B(u1__abc_73140_new_n1085_), .Y(u1__abc_73140_new_n1086_));
OR2X2 OR2X2_2297 ( .A(u1__abc_73140_new_n1083_), .B(u1__abc_73140_new_n1088_), .Y(mc_addr_d_12_));
OR2X2 OR2X2_2298 ( .A(u1__abc_73140_new_n904__bF_buf1), .B(\wb_addr_i[15] ), .Y(u1__abc_73140_new_n1090_));
OR2X2 OR2X2_2299 ( .A(u1__abc_73140_new_n906__bF_buf3), .B(u1_sram_addr_13_), .Y(u1__abc_73140_new_n1091_));
OR2X2 OR2X2_23 ( .A(_abc_85006_new_n240__bF_buf0), .B(spec_req_cs_5_bF_buf5_), .Y(_abc_85006_new_n272_));
OR2X2 OR2X2_230 ( .A(spec_req_cs_6_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1421_));
OR2X2 OR2X2_2300 ( .A(u1__abc_73140_new_n1092_), .B(u1__abc_73140_new_n900__bF_buf1), .Y(u1__abc_73140_new_n1093_));
OR2X2 OR2X2_2301 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_13_), .Y(u1__abc_73140_new_n1094_));
OR2X2 OR2X2_2302 ( .A(u1__abc_73140_new_n1096_), .B(u1__abc_73140_new_n1097_), .Y(mc_addr_d_13_));
OR2X2 OR2X2_2303 ( .A(u1__abc_73140_new_n904__bF_buf0), .B(\wb_addr_i[16] ), .Y(u1__abc_73140_new_n1099_));
OR2X2 OR2X2_2304 ( .A(u1__abc_73140_new_n906__bF_buf2), .B(u1_sram_addr_14_), .Y(u1__abc_73140_new_n1100_));
OR2X2 OR2X2_2305 ( .A(u1__abc_73140_new_n1101_), .B(u1__abc_73140_new_n900__bF_buf0), .Y(u1__abc_73140_new_n1102_));
OR2X2 OR2X2_2306 ( .A(u1__abc_73140_new_n913_), .B(u1_acs_addr_14_), .Y(u1__abc_73140_new_n1103_));
OR2X2 OR2X2_2307 ( .A(u1__abc_73140_new_n1105_), .B(u1__abc_73140_new_n1106_), .Y(mc_addr_d_14_));
OR2X2 OR2X2_2308 ( .A(u1__abc_73140_new_n1109_), .B(u1__abc_73140_new_n900__bF_buf4), .Y(u1__abc_73140_new_n1110_));
OR2X2 OR2X2_2309 ( .A(u1__abc_73140_new_n1110_), .B(u1__abc_73140_new_n1108_), .Y(u1__abc_73140_new_n1111_));
OR2X2 OR2X2_231 ( .A(u0__abc_76628_new_n1423_), .B(u0__abc_76628_new_n1419_), .Y(u0__abc_76628_new_n1424_));
OR2X2 OR2X2_2310 ( .A(u1__abc_73140_new_n898_), .B(u1_acs_addr_15_), .Y(u1__abc_73140_new_n1112_));
OR2X2 OR2X2_2311 ( .A(u1__abc_73140_new_n1116_), .B(u1__abc_73140_new_n900__bF_buf3), .Y(u1__abc_73140_new_n1117_));
OR2X2 OR2X2_2312 ( .A(u1__abc_73140_new_n1117_), .B(u1__abc_73140_new_n1115_), .Y(u1__abc_73140_new_n1118_));
OR2X2 OR2X2_2313 ( .A(u1__abc_73140_new_n898_), .B(u1_acs_addr_16_), .Y(u1__abc_73140_new_n1119_));
OR2X2 OR2X2_2314 ( .A(u1__abc_73140_new_n1123_), .B(u1__abc_73140_new_n900__bF_buf2), .Y(u1__abc_73140_new_n1124_));
OR2X2 OR2X2_2315 ( .A(u1__abc_73140_new_n1124_), .B(u1__abc_73140_new_n1122_), .Y(u1__abc_73140_new_n1125_));
OR2X2 OR2X2_2316 ( .A(u1__abc_73140_new_n898_), .B(u1_acs_addr_17_), .Y(u1__abc_73140_new_n1126_));
OR2X2 OR2X2_2317 ( .A(u1__abc_73140_new_n1130_), .B(u1__abc_73140_new_n900__bF_buf1), .Y(u1__abc_73140_new_n1131_));
OR2X2 OR2X2_2318 ( .A(u1__abc_73140_new_n1131_), .B(u1__abc_73140_new_n1129_), .Y(u1__abc_73140_new_n1132_));
OR2X2 OR2X2_2319 ( .A(u1__abc_73140_new_n898_), .B(u1_acs_addr_18_), .Y(u1__abc_73140_new_n1133_));
OR2X2 OR2X2_232 ( .A(u0__abc_76628_new_n1425_), .B(u0__abc_76628_new_n1426_), .Y(u0__abc_76628_new_n1427_));
OR2X2 OR2X2_2320 ( .A(u1__abc_73140_new_n1137_), .B(u1__abc_73140_new_n900__bF_buf0), .Y(u1__abc_73140_new_n1138_));
OR2X2 OR2X2_2321 ( .A(u1__abc_73140_new_n1138_), .B(u1__abc_73140_new_n1136_), .Y(u1__abc_73140_new_n1139_));
OR2X2 OR2X2_2322 ( .A(u1__abc_73140_new_n898_), .B(u1_acs_addr_19_), .Y(u1__abc_73140_new_n1140_));
OR2X2 OR2X2_2323 ( .A(u1__abc_73140_new_n1144_), .B(u1__abc_73140_new_n900__bF_buf4), .Y(u1__abc_73140_new_n1145_));
OR2X2 OR2X2_2324 ( .A(u1__abc_73140_new_n1145_), .B(u1__abc_73140_new_n1143_), .Y(u1__abc_73140_new_n1146_));
OR2X2 OR2X2_2325 ( .A(u1__abc_73140_new_n898_), .B(u1_acs_addr_20_), .Y(u1__abc_73140_new_n1147_));
OR2X2 OR2X2_2326 ( .A(u1__abc_73140_new_n1151_), .B(u1__abc_73140_new_n900__bF_buf3), .Y(u1__abc_73140_new_n1152_));
OR2X2 OR2X2_2327 ( .A(u1__abc_73140_new_n1152_), .B(u1__abc_73140_new_n1150_), .Y(u1__abc_73140_new_n1153_));
OR2X2 OR2X2_2328 ( .A(u1__abc_73140_new_n898_), .B(u1_acs_addr_21_), .Y(u1__abc_73140_new_n1154_));
OR2X2 OR2X2_2329 ( .A(u1__abc_73140_new_n1158_), .B(u1__abc_73140_new_n900__bF_buf2), .Y(u1__abc_73140_new_n1159_));
OR2X2 OR2X2_233 ( .A(u0__abc_76628_new_n1428_), .B(u0__abc_76628_new_n1429_), .Y(u0__abc_76628_new_n1430_));
OR2X2 OR2X2_2330 ( .A(u1__abc_73140_new_n1159_), .B(u1__abc_73140_new_n1157_), .Y(u1__abc_73140_new_n1160_));
OR2X2 OR2X2_2331 ( .A(u1__abc_73140_new_n898_), .B(u1_acs_addr_22_), .Y(u1__abc_73140_new_n1161_));
OR2X2 OR2X2_2332 ( .A(u1__abc_73140_new_n1165_), .B(u1__abc_73140_new_n1164_), .Y(u1__abc_73140_new_n1166_));
OR2X2 OR2X2_2333 ( .A(u1__abc_73140_new_n1166_), .B(u1__abc_73140_new_n900__bF_buf1), .Y(u1__abc_73140_new_n1167_));
OR2X2 OR2X2_2334 ( .A(u1__abc_73140_new_n898_), .B(u1_acs_addr_23_), .Y(u1__abc_73140_new_n1168_));
OR2X2 OR2X2_2335 ( .A(u1__abc_73140_new_n906__bF_buf0), .B(u1_sram_addr_10_), .Y(u1__abc_73140_new_n1171_));
OR2X2 OR2X2_2336 ( .A(u1__abc_73140_new_n904__bF_buf0), .B(\wb_addr_i[12] ), .Y(u1__abc_73140_new_n1172_));
OR2X2 OR2X2_2337 ( .A(u1__abc_73140_new_n1173_), .B(u1__abc_73140_new_n900__bF_buf0), .Y(u1__abc_73140_new_n1174_));
OR2X2 OR2X2_2338 ( .A(u1__abc_73140_new_n898_), .B(u1_acs_addr_10_), .Y(u1__abc_73140_new_n1175_));
OR2X2 OR2X2_2339 ( .A(u1__abc_73140_new_n921_), .B(row_adr_10_bF_buf2_), .Y(u1__abc_73140_new_n1178_));
OR2X2 OR2X2_234 ( .A(u0__abc_76628_new_n1431_), .B(u0__abc_76628_new_n1432_), .Y(u0__abc_76628_new_n1433_));
OR2X2 OR2X2_2340 ( .A(row_sel), .B(cmd_a10), .Y(u1__abc_73140_new_n1179_));
OR2X2 OR2X2_2341 ( .A(u1__abc_73140_new_n1180_), .B(u1__abc_73140_new_n918_), .Y(u1__abc_73140_new_n1181_));
OR2X2 OR2X2_2342 ( .A(u1__abc_73140_new_n919_), .B(tms_s_10_), .Y(u1__abc_73140_new_n1182_));
OR2X2 OR2X2_2343 ( .A(u1__abc_73140_new_n1184_), .B(rfr_ack), .Y(u1__abc_73140_new_n1185_));
OR2X2 OR2X2_2344 ( .A(u1__abc_73140_new_n1177_), .B(u1__abc_73140_new_n1185_), .Y(mc_addr_d_10_));
OR2X2 OR2X2_2345 ( .A(u1_acs_addr_0_), .B(u1_acs_addr_1_), .Y(u1_u0__abc_73035_new_n53_));
OR2X2 OR2X2_2346 ( .A(u1_u0__abc_73035_new_n51_), .B(u1_acs_addr_2_), .Y(u1_u0__abc_73035_new_n57_));
OR2X2 OR2X2_2347 ( .A(u1_u0__abc_73035_new_n55_), .B(u1_acs_addr_3_), .Y(u1_u0__abc_73035_new_n61_));
OR2X2 OR2X2_2348 ( .A(u1_u0__abc_73035_new_n59_), .B(u1_acs_addr_4_), .Y(u1_u0__abc_73035_new_n65_));
OR2X2 OR2X2_2349 ( .A(u1_u0__abc_73035_new_n63_), .B(u1_acs_addr_5_), .Y(u1_u0__abc_73035_new_n67_));
OR2X2 OR2X2_235 ( .A(u0__abc_76628_new_n1435_), .B(spec_req_cs_0_bF_buf4_), .Y(u0__abc_76628_new_n1436_));
OR2X2 OR2X2_2350 ( .A(u1_u0__abc_73035_new_n69_), .B(u1_acs_addr_6_), .Y(u1_u0__abc_73035_new_n74_));
OR2X2 OR2X2_2351 ( .A(u1_u0__abc_73035_new_n72_), .B(u1_acs_addr_7_), .Y(u1_u0__abc_73035_new_n76_));
OR2X2 OR2X2_2352 ( .A(u1_u0__abc_73035_new_n79_), .B(u1_acs_addr_8_), .Y(u1_u0__abc_73035_new_n84_));
OR2X2 OR2X2_2353 ( .A(u1_u0__abc_73035_new_n82_), .B(u1_acs_addr_9_), .Y(u1_u0__abc_73035_new_n86_));
OR2X2 OR2X2_2354 ( .A(u1_u0__abc_73035_new_n88_), .B(u1_acs_addr_10_), .Y(u1_u0__abc_73035_new_n93_));
OR2X2 OR2X2_2355 ( .A(u1_u0__abc_73035_new_n91_), .B(u1_acs_addr_11_), .Y(u1_u0__abc_73035_new_n99_));
OR2X2 OR2X2_2356 ( .A(u1_u0__abc_73035_new_n102_), .B(u1_acs_addr_13_), .Y(u1_u0__abc_73035_new_n105_));
OR2X2 OR2X2_2357 ( .A(u1_u0__abc_73035_new_n103_), .B(u1_acs_addr_14_), .Y(u1_u0__abc_73035_new_n109_));
OR2X2 OR2X2_2358 ( .A(u1_u0__abc_73035_new_n107_), .B(u1_acs_addr_15_), .Y(u1_u0__abc_73035_new_n111_));
OR2X2 OR2X2_2359 ( .A(u1_u0__abc_73035_new_n113_), .B(u1_acs_addr_16_), .Y(u1_u0__abc_73035_new_n118_));
OR2X2 OR2X2_236 ( .A(u0__abc_76628_new_n1434_), .B(u0__abc_76628_new_n1436_), .Y(u0__abc_76628_new_n1437_));
OR2X2 OR2X2_2360 ( .A(u1_u0__abc_73035_new_n116_), .B(u1_acs_addr_17_), .Y(u1_u0__abc_73035_new_n120_));
OR2X2 OR2X2_2361 ( .A(u1_u0__abc_73035_new_n122_), .B(u1_acs_addr_18_), .Y(u1_u0__abc_73035_new_n127_));
OR2X2 OR2X2_2362 ( .A(u1_u0__abc_73035_new_n125_), .B(u1_acs_addr_19_), .Y(u1_u0__abc_73035_new_n129_));
OR2X2 OR2X2_2363 ( .A(u1_u0__abc_73035_new_n132_), .B(u1_acs_addr_20_), .Y(u1_u0__abc_73035_new_n137_));
OR2X2 OR2X2_2364 ( .A(u1_u0__abc_73035_new_n135_), .B(u1_acs_addr_21_), .Y(u1_u0__abc_73035_new_n139_));
OR2X2 OR2X2_2365 ( .A(u1_u0__abc_73035_new_n141_), .B(u1_acs_addr_22_), .Y(u1_u0__abc_73035_new_n146_));
OR2X2 OR2X2_2366 ( .A(u1_u0__abc_73035_new_n144_), .B(u1_acs_addr_23_), .Y(u1_u0__abc_73035_new_n148_));
OR2X2 OR2X2_2367 ( .A(u1_u0_inc_next), .B(u1_acs_addr_12_), .Y(u1_u0__abc_73035_new_n153_));
OR2X2 OR2X2_2368 ( .A(u2__abc_75448_new_n80_), .B(rfr_ack), .Y(u2_bank_clr_all_0));
OR2X2 OR2X2_2369 ( .A(u2__abc_75448_new_n82_), .B(rfr_ack), .Y(u2_bank_clr_all_1));
OR2X2 OR2X2_237 ( .A(u0__abc_76628_new_n1197__bF_buf1), .B(u0_tms0_10_), .Y(u0__abc_76628_new_n1438_));
OR2X2 OR2X2_2370 ( .A(u2__abc_75448_new_n96_), .B(u2__abc_75448_new_n97_), .Y(u2__abc_75448_new_n98_));
OR2X2 OR2X2_2371 ( .A(u2__abc_75448_new_n99_), .B(u2__abc_75448_new_n100_), .Y(u2__abc_75448_new_n101_));
OR2X2 OR2X2_2372 ( .A(u2__abc_75448_new_n98_), .B(u2__abc_75448_new_n101_), .Y(u2__abc_75448_new_n102_));
OR2X2 OR2X2_2373 ( .A(u2__abc_75448_new_n103_), .B(u2__abc_75448_new_n104_), .Y(u2__abc_75448_new_n105_));
OR2X2 OR2X2_2374 ( .A(u2__abc_75448_new_n106_), .B(u2__abc_75448_new_n107_), .Y(u2__abc_75448_new_n108_));
OR2X2 OR2X2_2375 ( .A(u2__abc_75448_new_n105_), .B(u2__abc_75448_new_n108_), .Y(u2__abc_75448_new_n109_));
OR2X2 OR2X2_2376 ( .A(u2__abc_75448_new_n102_), .B(u2__abc_75448_new_n109_), .Y(u2__0bank_open_0_0_));
OR2X2 OR2X2_2377 ( .A(u2__abc_75448_new_n111_), .B(u2__abc_75448_new_n112_), .Y(u2__abc_75448_new_n113_));
OR2X2 OR2X2_2378 ( .A(u2__abc_75448_new_n114_), .B(u2__abc_75448_new_n115_), .Y(u2__abc_75448_new_n116_));
OR2X2 OR2X2_2379 ( .A(u2__abc_75448_new_n113_), .B(u2__abc_75448_new_n116_), .Y(u2__abc_75448_new_n117_));
OR2X2 OR2X2_238 ( .A(u0__abc_76628_new_n1440_), .B(u0__abc_76628_new_n1418_), .Y(u0__0sp_tms_31_0__10_));
OR2X2 OR2X2_2380 ( .A(u2__abc_75448_new_n118_), .B(u2__abc_75448_new_n119_), .Y(u2__abc_75448_new_n120_));
OR2X2 OR2X2_2381 ( .A(u2__abc_75448_new_n121_), .B(u2__abc_75448_new_n122_), .Y(u2__abc_75448_new_n123_));
OR2X2 OR2X2_2382 ( .A(u2__abc_75448_new_n120_), .B(u2__abc_75448_new_n123_), .Y(u2__abc_75448_new_n124_));
OR2X2 OR2X2_2383 ( .A(u2__abc_75448_new_n117_), .B(u2__abc_75448_new_n124_), .Y(u2__0row_same_0_0_));
OR2X2 OR2X2_2384 ( .A(u2_u0__abc_74955_new_n137__bF_buf4), .B(u2_u0_b3_last_row_0_), .Y(u2_u0__abc_74955_new_n138_));
OR2X2 OR2X2_2385 ( .A(u2_u0__abc_74955_new_n137__bF_buf2), .B(u2_u0_b3_last_row_1_), .Y(u2_u0__abc_74955_new_n143_));
OR2X2 OR2X2_2386 ( .A(u2_u0__abc_74955_new_n137__bF_buf0), .B(u2_u0_b3_last_row_2_), .Y(u2_u0__abc_74955_new_n148_));
OR2X2 OR2X2_2387 ( .A(u2_u0__abc_74955_new_n137__bF_buf3), .B(u2_u0_b3_last_row_3_), .Y(u2_u0__abc_74955_new_n153_));
OR2X2 OR2X2_2388 ( .A(u2_u0__abc_74955_new_n137__bF_buf1), .B(u2_u0_b3_last_row_4_), .Y(u2_u0__abc_74955_new_n158_));
OR2X2 OR2X2_2389 ( .A(u2_u0__abc_74955_new_n137__bF_buf4), .B(u2_u0_b3_last_row_5_), .Y(u2_u0__abc_74955_new_n163_));
OR2X2 OR2X2_239 ( .A(u0__abc_76628_new_n1177__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n1444_));
OR2X2 OR2X2_2390 ( .A(u2_u0__abc_74955_new_n137__bF_buf2), .B(u2_u0_b3_last_row_6_), .Y(u2_u0__abc_74955_new_n168_));
OR2X2 OR2X2_2391 ( .A(u2_u0__abc_74955_new_n137__bF_buf0), .B(u2_u0_b3_last_row_7_), .Y(u2_u0__abc_74955_new_n173_));
OR2X2 OR2X2_2392 ( .A(u2_u0__abc_74955_new_n137__bF_buf3), .B(u2_u0_b3_last_row_8_), .Y(u2_u0__abc_74955_new_n178_));
OR2X2 OR2X2_2393 ( .A(u2_u0__abc_74955_new_n137__bF_buf1), .B(u2_u0_b3_last_row_9_), .Y(u2_u0__abc_74955_new_n183_));
OR2X2 OR2X2_2394 ( .A(u2_u0__abc_74955_new_n137__bF_buf4), .B(u2_u0_b3_last_row_10_), .Y(u2_u0__abc_74955_new_n188_));
OR2X2 OR2X2_2395 ( .A(u2_u0__abc_74955_new_n137__bF_buf2), .B(u2_u0_b3_last_row_11_), .Y(u2_u0__abc_74955_new_n193_));
OR2X2 OR2X2_2396 ( .A(u2_u0__abc_74955_new_n137__bF_buf0), .B(u2_u0_b3_last_row_12_), .Y(u2_u0__abc_74955_new_n198_));
OR2X2 OR2X2_2397 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_0_), .Y(u2_u0__abc_74955_new_n207_));
OR2X2 OR2X2_2398 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_0_bF_buf0_), .Y(u2_u0__abc_74955_new_n209_));
OR2X2 OR2X2_2399 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_1_), .Y(u2_u0__abc_74955_new_n211_));
OR2X2 OR2X2_24 ( .A(lmr_sel_bF_buf1), .B(cs_5_), .Y(_abc_85006_new_n273_));
OR2X2 OR2X2_240 ( .A(spec_req_cs_6_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1445_));
OR2X2 OR2X2_2400 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_1_bF_buf0_), .Y(u2_u0__abc_74955_new_n212_));
OR2X2 OR2X2_2401 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_2_), .Y(u2_u0__abc_74955_new_n214_));
OR2X2 OR2X2_2402 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_2_bF_buf0_), .Y(u2_u0__abc_74955_new_n215_));
OR2X2 OR2X2_2403 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_3_), .Y(u2_u0__abc_74955_new_n217_));
OR2X2 OR2X2_2404 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_3_bF_buf0_), .Y(u2_u0__abc_74955_new_n218_));
OR2X2 OR2X2_2405 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_4_), .Y(u2_u0__abc_74955_new_n220_));
OR2X2 OR2X2_2406 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_4_bF_buf0_), .Y(u2_u0__abc_74955_new_n221_));
OR2X2 OR2X2_2407 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_5_), .Y(u2_u0__abc_74955_new_n223_));
OR2X2 OR2X2_2408 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_5_bF_buf0_), .Y(u2_u0__abc_74955_new_n224_));
OR2X2 OR2X2_2409 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_6_), .Y(u2_u0__abc_74955_new_n226_));
OR2X2 OR2X2_241 ( .A(u0__abc_76628_new_n1447_), .B(u0__abc_76628_new_n1443_), .Y(u0__abc_76628_new_n1448_));
OR2X2 OR2X2_2410 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_6_bF_buf0_), .Y(u2_u0__abc_74955_new_n227_));
OR2X2 OR2X2_2411 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_7_), .Y(u2_u0__abc_74955_new_n229_));
OR2X2 OR2X2_2412 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_7_bF_buf0_), .Y(u2_u0__abc_74955_new_n230_));
OR2X2 OR2X2_2413 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_8_), .Y(u2_u0__abc_74955_new_n232_));
OR2X2 OR2X2_2414 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_8_bF_buf0_), .Y(u2_u0__abc_74955_new_n233_));
OR2X2 OR2X2_2415 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_9_), .Y(u2_u0__abc_74955_new_n235_));
OR2X2 OR2X2_2416 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_9_bF_buf0_), .Y(u2_u0__abc_74955_new_n236_));
OR2X2 OR2X2_2417 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_10_), .Y(u2_u0__abc_74955_new_n238_));
OR2X2 OR2X2_2418 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_10_bF_buf0_), .Y(u2_u0__abc_74955_new_n239_));
OR2X2 OR2X2_2419 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_11_), .Y(u2_u0__abc_74955_new_n241_));
OR2X2 OR2X2_242 ( .A(u0__abc_76628_new_n1449_), .B(u0__abc_76628_new_n1450_), .Y(u0__abc_76628_new_n1451_));
OR2X2 OR2X2_2420 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_11_bF_buf0_), .Y(u2_u0__abc_74955_new_n242_));
OR2X2 OR2X2_2421 ( .A(u2_u0__abc_74955_new_n206_), .B(u2_u0_b0_last_row_12_), .Y(u2_u0__abc_74955_new_n244_));
OR2X2 OR2X2_2422 ( .A(u2_u0__abc_74955_new_n208_), .B(row_adr_12_bF_buf0_), .Y(u2_u0__abc_74955_new_n245_));
OR2X2 OR2X2_2423 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_0_), .Y(u2_u0__abc_74955_new_n249_));
OR2X2 OR2X2_2424 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_0_bF_buf3_), .Y(u2_u0__abc_74955_new_n251_));
OR2X2 OR2X2_2425 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_1_), .Y(u2_u0__abc_74955_new_n253_));
OR2X2 OR2X2_2426 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_1_bF_buf3_), .Y(u2_u0__abc_74955_new_n254_));
OR2X2 OR2X2_2427 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_2_), .Y(u2_u0__abc_74955_new_n256_));
OR2X2 OR2X2_2428 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_2_bF_buf3_), .Y(u2_u0__abc_74955_new_n257_));
OR2X2 OR2X2_2429 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_3_), .Y(u2_u0__abc_74955_new_n259_));
OR2X2 OR2X2_243 ( .A(u0__abc_76628_new_n1452_), .B(u0__abc_76628_new_n1453_), .Y(u0__abc_76628_new_n1454_));
OR2X2 OR2X2_2430 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_3_bF_buf3_), .Y(u2_u0__abc_74955_new_n260_));
OR2X2 OR2X2_2431 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_4_), .Y(u2_u0__abc_74955_new_n262_));
OR2X2 OR2X2_2432 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_4_bF_buf3_), .Y(u2_u0__abc_74955_new_n263_));
OR2X2 OR2X2_2433 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_5_), .Y(u2_u0__abc_74955_new_n265_));
OR2X2 OR2X2_2434 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_5_bF_buf3_), .Y(u2_u0__abc_74955_new_n266_));
OR2X2 OR2X2_2435 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_6_), .Y(u2_u0__abc_74955_new_n268_));
OR2X2 OR2X2_2436 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_6_bF_buf3_), .Y(u2_u0__abc_74955_new_n269_));
OR2X2 OR2X2_2437 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_7_), .Y(u2_u0__abc_74955_new_n271_));
OR2X2 OR2X2_2438 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_7_bF_buf3_), .Y(u2_u0__abc_74955_new_n272_));
OR2X2 OR2X2_2439 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_8_), .Y(u2_u0__abc_74955_new_n274_));
OR2X2 OR2X2_244 ( .A(u0__abc_76628_new_n1455_), .B(u0__abc_76628_new_n1456_), .Y(u0__abc_76628_new_n1457_));
OR2X2 OR2X2_2440 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_8_bF_buf3_), .Y(u2_u0__abc_74955_new_n275_));
OR2X2 OR2X2_2441 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_9_), .Y(u2_u0__abc_74955_new_n277_));
OR2X2 OR2X2_2442 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_9_bF_buf3_), .Y(u2_u0__abc_74955_new_n278_));
OR2X2 OR2X2_2443 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_10_), .Y(u2_u0__abc_74955_new_n280_));
OR2X2 OR2X2_2444 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_10_bF_buf3_), .Y(u2_u0__abc_74955_new_n281_));
OR2X2 OR2X2_2445 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_11_), .Y(u2_u0__abc_74955_new_n283_));
OR2X2 OR2X2_2446 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_11_bF_buf3_), .Y(u2_u0__abc_74955_new_n284_));
OR2X2 OR2X2_2447 ( .A(u2_u0__abc_74955_new_n248_), .B(u2_u0_b1_last_row_12_), .Y(u2_u0__abc_74955_new_n286_));
OR2X2 OR2X2_2448 ( .A(u2_u0__abc_74955_new_n250_), .B(row_adr_12_bF_buf3_), .Y(u2_u0__abc_74955_new_n287_));
OR2X2 OR2X2_2449 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_0_), .Y(u2_u0__abc_74955_new_n291_));
OR2X2 OR2X2_245 ( .A(u0__abc_76628_new_n1459_), .B(spec_req_cs_0_bF_buf3_), .Y(u0__abc_76628_new_n1460_));
OR2X2 OR2X2_2450 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_0_bF_buf2_), .Y(u2_u0__abc_74955_new_n293_));
OR2X2 OR2X2_2451 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_1_), .Y(u2_u0__abc_74955_new_n295_));
OR2X2 OR2X2_2452 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_1_bF_buf2_), .Y(u2_u0__abc_74955_new_n296_));
OR2X2 OR2X2_2453 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_2_), .Y(u2_u0__abc_74955_new_n298_));
OR2X2 OR2X2_2454 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_2_bF_buf2_), .Y(u2_u0__abc_74955_new_n299_));
OR2X2 OR2X2_2455 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_3_), .Y(u2_u0__abc_74955_new_n301_));
OR2X2 OR2X2_2456 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_3_bF_buf2_), .Y(u2_u0__abc_74955_new_n302_));
OR2X2 OR2X2_2457 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_4_), .Y(u2_u0__abc_74955_new_n304_));
OR2X2 OR2X2_2458 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_4_bF_buf2_), .Y(u2_u0__abc_74955_new_n305_));
OR2X2 OR2X2_2459 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_5_), .Y(u2_u0__abc_74955_new_n307_));
OR2X2 OR2X2_246 ( .A(u0__abc_76628_new_n1458_), .B(u0__abc_76628_new_n1460_), .Y(u0__abc_76628_new_n1461_));
OR2X2 OR2X2_2460 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_5_bF_buf2_), .Y(u2_u0__abc_74955_new_n308_));
OR2X2 OR2X2_2461 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_6_), .Y(u2_u0__abc_74955_new_n310_));
OR2X2 OR2X2_2462 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_6_bF_buf2_), .Y(u2_u0__abc_74955_new_n311_));
OR2X2 OR2X2_2463 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_7_), .Y(u2_u0__abc_74955_new_n313_));
OR2X2 OR2X2_2464 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_7_bF_buf2_), .Y(u2_u0__abc_74955_new_n314_));
OR2X2 OR2X2_2465 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_8_), .Y(u2_u0__abc_74955_new_n316_));
OR2X2 OR2X2_2466 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_8_bF_buf2_), .Y(u2_u0__abc_74955_new_n317_));
OR2X2 OR2X2_2467 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_9_), .Y(u2_u0__abc_74955_new_n319_));
OR2X2 OR2X2_2468 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_9_bF_buf2_), .Y(u2_u0__abc_74955_new_n320_));
OR2X2 OR2X2_2469 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_10_), .Y(u2_u0__abc_74955_new_n322_));
OR2X2 OR2X2_247 ( .A(u0__abc_76628_new_n1197__bF_buf0), .B(u0_tms0_11_), .Y(u0__abc_76628_new_n1462_));
OR2X2 OR2X2_2470 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_10_bF_buf2_), .Y(u2_u0__abc_74955_new_n323_));
OR2X2 OR2X2_2471 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_11_), .Y(u2_u0__abc_74955_new_n325_));
OR2X2 OR2X2_2472 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_11_bF_buf2_), .Y(u2_u0__abc_74955_new_n326_));
OR2X2 OR2X2_2473 ( .A(u2_u0__abc_74955_new_n290_), .B(u2_u0_b2_last_row_12_), .Y(u2_u0__abc_74955_new_n328_));
OR2X2 OR2X2_2474 ( .A(u2_u0__abc_74955_new_n292_), .B(row_adr_12_bF_buf2_), .Y(u2_u0__abc_74955_new_n329_));
OR2X2 OR2X2_2475 ( .A(u2_u0__abc_74955_new_n179_), .B(u2_u0_b3_last_row_8_), .Y(u2_u0__abc_74955_new_n331_));
OR2X2 OR2X2_2476 ( .A(u2_u0__abc_74955_new_n332_), .B(row_adr_9_bF_buf1_), .Y(u2_u0__abc_74955_new_n333_));
OR2X2 OR2X2_2477 ( .A(u2_u0__abc_74955_new_n334_), .B(row_adr_8_bF_buf1_), .Y(u2_u0__abc_74955_new_n335_));
OR2X2 OR2X2_2478 ( .A(u2_u0__abc_74955_new_n184_), .B(u2_u0_b3_last_row_9_), .Y(u2_u0__abc_74955_new_n338_));
OR2X2 OR2X2_2479 ( .A(u2_u0__abc_74955_new_n339_), .B(row_adr_11_bF_buf1_), .Y(u2_u0__abc_74955_new_n340_));
OR2X2 OR2X2_248 ( .A(u0__abc_76628_new_n1464_), .B(u0__abc_76628_new_n1442_), .Y(u0__0sp_tms_31_0__11_));
OR2X2 OR2X2_2480 ( .A(u2_u0__abc_74955_new_n342_), .B(row_adr_4_bF_buf1_), .Y(u2_u0__abc_74955_new_n343_));
OR2X2 OR2X2_2481 ( .A(u2_u0__abc_74955_new_n194_), .B(u2_u0_b3_last_row_11_), .Y(u2_u0__abc_74955_new_n344_));
OR2X2 OR2X2_2482 ( .A(u2_u0__abc_74955_new_n349_), .B(u2_u0__abc_74955_new_n350_), .Y(u2_u0__abc_74955_new_n351_));
OR2X2 OR2X2_2483 ( .A(u2_u0__abc_74955_new_n144_), .B(u2_u0_b3_last_row_1_), .Y(u2_u0__abc_74955_new_n352_));
OR2X2 OR2X2_2484 ( .A(u2_u0__abc_74955_new_n355_), .B(row_adr_7_bF_buf1_), .Y(u2_u0__abc_74955_new_n356_));
OR2X2 OR2X2_2485 ( .A(u2_u0__abc_74955_new_n174_), .B(u2_u0_b3_last_row_7_), .Y(u2_u0__abc_74955_new_n357_));
OR2X2 OR2X2_2486 ( .A(u2_u0__abc_74955_new_n359_), .B(row_adr_5_bF_buf1_), .Y(u2_u0__abc_74955_new_n360_));
OR2X2 OR2X2_2487 ( .A(u2_u0__abc_74955_new_n164_), .B(u2_u0_b3_last_row_5_), .Y(u2_u0__abc_74955_new_n361_));
OR2X2 OR2X2_2488 ( .A(u2_u0__abc_74955_new_n199_), .B(u2_u0_b3_last_row_12_), .Y(u2_u0__abc_74955_new_n366_));
OR2X2 OR2X2_2489 ( .A(u2_u0__abc_74955_new_n367_), .B(row_adr_12_bF_buf1_), .Y(u2_u0__abc_74955_new_n368_));
OR2X2 OR2X2_249 ( .A(u0__abc_76628_new_n1177__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n1468_));
OR2X2 OR2X2_2490 ( .A(u2_u0__abc_74955_new_n189_), .B(u2_u0_b3_last_row_10_), .Y(u2_u0__abc_74955_new_n370_));
OR2X2 OR2X2_2491 ( .A(u2_u0__abc_74955_new_n371_), .B(row_adr_10_bF_buf1_), .Y(u2_u0__abc_74955_new_n372_));
OR2X2 OR2X2_2492 ( .A(u2_u0__abc_74955_new_n375_), .B(row_adr_3_bF_buf1_), .Y(u2_u0__abc_74955_new_n376_));
OR2X2 OR2X2_2493 ( .A(u2_u0__abc_74955_new_n154_), .B(u2_u0_b3_last_row_3_), .Y(u2_u0__abc_74955_new_n377_));
OR2X2 OR2X2_2494 ( .A(u2_u0__abc_74955_new_n379_), .B(row_adr_1_bF_buf1_), .Y(u2_u0__abc_74955_new_n380_));
OR2X2 OR2X2_2495 ( .A(u2_u0__abc_74955_new_n149_), .B(u2_u0_b3_last_row_2_), .Y(u2_u0__abc_74955_new_n381_));
OR2X2 OR2X2_2496 ( .A(u2_u0__abc_74955_new_n159_), .B(u2_u0_b3_last_row_4_), .Y(u2_u0__abc_74955_new_n384_));
OR2X2 OR2X2_2497 ( .A(u2_u0__abc_74955_new_n385_), .B(row_adr_6_bF_buf1_), .Y(u2_u0__abc_74955_new_n386_));
OR2X2 OR2X2_2498 ( .A(u2_u0__abc_74955_new_n388_), .B(row_adr_2_bF_buf1_), .Y(u2_u0__abc_74955_new_n389_));
OR2X2 OR2X2_2499 ( .A(u2_u0__abc_74955_new_n169_), .B(u2_u0_b3_last_row_6_), .Y(u2_u0__abc_74955_new_n390_));
OR2X2 OR2X2_25 ( .A(_abc_85006_new_n274_), .B(_abc_85006_new_n237_), .Y(_abc_85006_new_n275_));
OR2X2 OR2X2_250 ( .A(spec_req_cs_6_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1469_));
OR2X2 OR2X2_2500 ( .A(u2_u0__abc_74955_new_n144_), .B(u2_u0_b1_last_row_1_), .Y(u2_u0__abc_74955_new_n396_));
OR2X2 OR2X2_2501 ( .A(u2_u0__abc_74955_new_n139_), .B(u2_u0_b1_last_row_0_), .Y(u2_u0__abc_74955_new_n397_));
OR2X2 OR2X2_2502 ( .A(u2_u0__abc_74955_new_n399_), .B(row_adr_0_bF_buf0_), .Y(u2_u0__abc_74955_new_n400_));
OR2X2 OR2X2_2503 ( .A(u2_u0__abc_74955_new_n159_), .B(u2_u0_b1_last_row_4_), .Y(u2_u0__abc_74955_new_n402_));
OR2X2 OR2X2_2504 ( .A(u2_u0__abc_74955_new_n403_), .B(row_adr_4_bF_buf0_), .Y(u2_u0__abc_74955_new_n404_));
OR2X2 OR2X2_2505 ( .A(u2_u0__abc_74955_new_n164_), .B(u2_u0_b1_last_row_5_), .Y(u2_u0__abc_74955_new_n406_));
OR2X2 OR2X2_2506 ( .A(u2_u0__abc_74955_new_n407_), .B(row_adr_3_bF_buf0_), .Y(u2_u0__abc_74955_new_n408_));
OR2X2 OR2X2_2507 ( .A(u2_u0__abc_74955_new_n179_), .B(u2_u0_b1_last_row_8_), .Y(u2_u0__abc_74955_new_n412_));
OR2X2 OR2X2_2508 ( .A(u2_u0__abc_74955_new_n413_), .B(row_adr_8_bF_buf0_), .Y(u2_u0__abc_74955_new_n414_));
OR2X2 OR2X2_2509 ( .A(u2_u0__abc_74955_new_n169_), .B(u2_u0_b1_last_row_6_), .Y(u2_u0__abc_74955_new_n416_));
OR2X2 OR2X2_251 ( .A(u0__abc_76628_new_n1471_), .B(u0__abc_76628_new_n1467_), .Y(u0__abc_76628_new_n1472_));
OR2X2 OR2X2_2510 ( .A(u2_u0__abc_74955_new_n417_), .B(row_adr_6_bF_buf0_), .Y(u2_u0__abc_74955_new_n418_));
OR2X2 OR2X2_2511 ( .A(u2_u0__abc_74955_new_n199_), .B(u2_u0_b1_last_row_12_), .Y(u2_u0__abc_74955_new_n421_));
OR2X2 OR2X2_2512 ( .A(u2_u0__abc_74955_new_n422_), .B(row_adr_12_bF_buf0_), .Y(u2_u0__abc_74955_new_n423_));
OR2X2 OR2X2_2513 ( .A(u2_u0__abc_74955_new_n425_), .B(row_adr_11_bF_buf0_), .Y(u2_u0__abc_74955_new_n426_));
OR2X2 OR2X2_2514 ( .A(u2_u0__abc_74955_new_n431_), .B(row_adr_2_bF_buf0_), .Y(u2_u0__abc_74955_new_n432_));
OR2X2 OR2X2_2515 ( .A(u2_u0__abc_74955_new_n149_), .B(u2_u0_b1_last_row_2_), .Y(u2_u0__abc_74955_new_n433_));
OR2X2 OR2X2_2516 ( .A(u2_u0__abc_74955_new_n435_), .B(row_adr_1_bF_buf0_), .Y(u2_u0__abc_74955_new_n436_));
OR2X2 OR2X2_2517 ( .A(u2_u0__abc_74955_new_n154_), .B(u2_u0_b1_last_row_3_), .Y(u2_u0__abc_74955_new_n437_));
OR2X2 OR2X2_2518 ( .A(u2_u0__abc_74955_new_n440_), .B(row_adr_10_bF_buf0_), .Y(u2_u0__abc_74955_new_n441_));
OR2X2 OR2X2_2519 ( .A(u2_u0__abc_74955_new_n189_), .B(u2_u0_b1_last_row_10_), .Y(u2_u0__abc_74955_new_n442_));
OR2X2 OR2X2_252 ( .A(u0__abc_76628_new_n1473_), .B(u0__abc_76628_new_n1474_), .Y(u0__abc_76628_new_n1475_));
OR2X2 OR2X2_2520 ( .A(u2_u0__abc_74955_new_n444_), .B(row_adr_9_bF_buf0_), .Y(u2_u0__abc_74955_new_n445_));
OR2X2 OR2X2_2521 ( .A(u2_u0__abc_74955_new_n194_), .B(u2_u0_b1_last_row_11_), .Y(u2_u0__abc_74955_new_n446_));
OR2X2 OR2X2_2522 ( .A(u2_u0__abc_74955_new_n184_), .B(u2_u0_b1_last_row_9_), .Y(u2_u0__abc_74955_new_n449_));
OR2X2 OR2X2_2523 ( .A(u2_u0__abc_74955_new_n450_), .B(row_adr_7_bF_buf0_), .Y(u2_u0__abc_74955_new_n451_));
OR2X2 OR2X2_2524 ( .A(u2_u0__abc_74955_new_n174_), .B(u2_u0_b1_last_row_7_), .Y(u2_u0__abc_74955_new_n453_));
OR2X2 OR2X2_2525 ( .A(u2_u0__abc_74955_new_n454_), .B(row_adr_5_bF_buf0_), .Y(u2_u0__abc_74955_new_n455_));
OR2X2 OR2X2_2526 ( .A(u2_u0__abc_74955_new_n395_), .B(u2_u0__abc_74955_new_n460_), .Y(u2_u0__abc_74955_new_n461_));
OR2X2 OR2X2_2527 ( .A(u2_u0__abc_74955_new_n462_), .B(row_adr_9_bF_buf3_), .Y(u2_u0__abc_74955_new_n463_));
OR2X2 OR2X2_2528 ( .A(u2_u0__abc_74955_new_n194_), .B(u2_u0_b0_last_row_11_), .Y(u2_u0__abc_74955_new_n464_));
OR2X2 OR2X2_2529 ( .A(u2_u0__abc_74955_new_n184_), .B(u2_u0_b0_last_row_9_), .Y(u2_u0__abc_74955_new_n465_));
OR2X2 OR2X2_253 ( .A(u0__abc_76628_new_n1476_), .B(u0__abc_76628_new_n1477_), .Y(u0__abc_76628_new_n1478_));
OR2X2 OR2X2_2530 ( .A(u2_u0__abc_74955_new_n154_), .B(u2_u0_b0_last_row_3_), .Y(u2_u0__abc_74955_new_n468_));
OR2X2 OR2X2_2531 ( .A(u2_u0__abc_74955_new_n469_), .B(row_adr_12_bF_buf3_), .Y(u2_u0__abc_74955_new_n470_));
OR2X2 OR2X2_2532 ( .A(u2_u0__abc_74955_new_n472_), .B(row_adr_3_bF_buf3_), .Y(u2_u0__abc_74955_new_n473_));
OR2X2 OR2X2_2533 ( .A(u2_u0__abc_74955_new_n179_), .B(u2_u0_b0_last_row_8_), .Y(u2_u0__abc_74955_new_n474_));
OR2X2 OR2X2_2534 ( .A(u2_u0__abc_74955_new_n477_), .B(row_adr_2_bF_buf3_), .Y(u2_u0__abc_74955_new_n478_));
OR2X2 OR2X2_2535 ( .A(u2_u0__abc_74955_new_n479_), .B(row_adr_6_bF_buf3_), .Y(u2_u0__abc_74955_new_n480_));
OR2X2 OR2X2_2536 ( .A(u2_u0__abc_74955_new_n169_), .B(u2_u0_b0_last_row_6_), .Y(u2_u0__abc_74955_new_n482_));
OR2X2 OR2X2_2537 ( .A(u2_u0__abc_74955_new_n199_), .B(u2_u0_b0_last_row_12_), .Y(u2_u0__abc_74955_new_n483_));
OR2X2 OR2X2_2538 ( .A(u2_u0__abc_74955_new_n489_), .B(u2_u0__abc_74955_new_n490_), .Y(u2_u0__abc_74955_new_n491_));
OR2X2 OR2X2_2539 ( .A(u2_u0__abc_74955_new_n492_), .B(row_adr_1_bF_buf3_), .Y(u2_u0__abc_74955_new_n493_));
OR2X2 OR2X2_254 ( .A(u0__abc_76628_new_n1479_), .B(u0__abc_76628_new_n1480_), .Y(u0__abc_76628_new_n1481_));
OR2X2 OR2X2_2540 ( .A(u2_u0__abc_74955_new_n144_), .B(u2_u0_b0_last_row_1_), .Y(u2_u0__abc_74955_new_n494_));
OR2X2 OR2X2_2541 ( .A(u2_u0__abc_74955_new_n164_), .B(u2_u0_b0_last_row_5_), .Y(u2_u0__abc_74955_new_n497_));
OR2X2 OR2X2_2542 ( .A(u2_u0__abc_74955_new_n498_), .B(row_adr_5_bF_buf3_), .Y(u2_u0__abc_74955_new_n499_));
OR2X2 OR2X2_2543 ( .A(u2_u0__abc_74955_new_n501_), .B(row_adr_8_bF_buf3_), .Y(u2_u0__abc_74955_new_n502_));
OR2X2 OR2X2_2544 ( .A(u2_u0__abc_74955_new_n506_), .B(row_adr_4_bF_buf3_), .Y(u2_u0__abc_74955_new_n507_));
OR2X2 OR2X2_2545 ( .A(u2_u0__abc_74955_new_n508_), .B(row_adr_11_bF_buf3_), .Y(u2_u0__abc_74955_new_n509_));
OR2X2 OR2X2_2546 ( .A(u2_u0__abc_74955_new_n149_), .B(u2_u0_b0_last_row_2_), .Y(u2_u0__abc_74955_new_n511_));
OR2X2 OR2X2_2547 ( .A(u2_u0__abc_74955_new_n159_), .B(u2_u0_b0_last_row_4_), .Y(u2_u0__abc_74955_new_n512_));
OR2X2 OR2X2_2548 ( .A(u2_u0__abc_74955_new_n174_), .B(u2_u0_b0_last_row_7_), .Y(u2_u0__abc_74955_new_n515_));
OR2X2 OR2X2_2549 ( .A(u2_u0__abc_74955_new_n516_), .B(row_adr_7_bF_buf3_), .Y(u2_u0__abc_74955_new_n517_));
OR2X2 OR2X2_255 ( .A(u0__abc_76628_new_n1483_), .B(spec_req_cs_0_bF_buf2_), .Y(u0__abc_76628_new_n1484_));
OR2X2 OR2X2_2550 ( .A(u2_u0__abc_74955_new_n189_), .B(u2_u0_b0_last_row_10_), .Y(u2_u0__abc_74955_new_n519_));
OR2X2 OR2X2_2551 ( .A(u2_u0__abc_74955_new_n520_), .B(row_adr_10_bF_buf3_), .Y(u2_u0__abc_74955_new_n521_));
OR2X2 OR2X2_2552 ( .A(u2_u0__abc_74955_new_n527_), .B(row_adr_8_bF_buf2_), .Y(u2_u0__abc_74955_new_n528_));
OR2X2 OR2X2_2553 ( .A(u2_u0__abc_74955_new_n184_), .B(u2_u0_b2_last_row_9_), .Y(u2_u0__abc_74955_new_n529_));
OR2X2 OR2X2_2554 ( .A(u2_u0__abc_74955_new_n179_), .B(u2_u0_b2_last_row_8_), .Y(u2_u0__abc_74955_new_n530_));
OR2X2 OR2X2_2555 ( .A(u2_u0__abc_74955_new_n533_), .B(row_adr_9_bF_buf2_), .Y(u2_u0__abc_74955_new_n534_));
OR2X2 OR2X2_2556 ( .A(u2_u0__abc_74955_new_n194_), .B(u2_u0_b2_last_row_11_), .Y(u2_u0__abc_74955_new_n535_));
OR2X2 OR2X2_2557 ( .A(u2_u0__abc_74955_new_n537_), .B(row_adr_11_bF_buf2_), .Y(u2_u0__abc_74955_new_n538_));
OR2X2 OR2X2_2558 ( .A(u2_u0__abc_74955_new_n159_), .B(u2_u0_b2_last_row_4_), .Y(u2_u0__abc_74955_new_n539_));
OR2X2 OR2X2_2559 ( .A(u2_u0__abc_74955_new_n174_), .B(u2_u0_b2_last_row_7_), .Y(u2_u0__abc_74955_new_n543_));
OR2X2 OR2X2_256 ( .A(u0__abc_76628_new_n1482_), .B(u0__abc_76628_new_n1484_), .Y(u0__abc_76628_new_n1485_));
OR2X2 OR2X2_2560 ( .A(u2_u0__abc_74955_new_n544_), .B(row_adr_7_bF_buf2_), .Y(u2_u0__abc_74955_new_n545_));
OR2X2 OR2X2_2561 ( .A(u2_u0__abc_74955_new_n149_), .B(u2_u0_b2_last_row_2_), .Y(u2_u0__abc_74955_new_n547_));
OR2X2 OR2X2_2562 ( .A(u2_u0__abc_74955_new_n548_), .B(row_adr_6_bF_buf2_), .Y(u2_u0__abc_74955_new_n549_));
OR2X2 OR2X2_2563 ( .A(u2_u0__abc_74955_new_n154_), .B(u2_u0_b2_last_row_3_), .Y(u2_u0__abc_74955_new_n552_));
OR2X2 OR2X2_2564 ( .A(u2_u0__abc_74955_new_n553_), .B(row_adr_3_bF_buf2_), .Y(u2_u0__abc_74955_new_n554_));
OR2X2 OR2X2_2565 ( .A(u2_u0__abc_74955_new_n144_), .B(u2_u0_b2_last_row_1_), .Y(u2_u0__abc_74955_new_n556_));
OR2X2 OR2X2_2566 ( .A(u2_u0__abc_74955_new_n557_), .B(row_adr_2_bF_buf2_), .Y(u2_u0__abc_74955_new_n558_));
OR2X2 OR2X2_2567 ( .A(u2_u0__abc_74955_new_n563_), .B(row_adr_12_bF_buf2_), .Y(u2_u0__abc_74955_new_n564_));
OR2X2 OR2X2_2568 ( .A(u2_u0__abc_74955_new_n199_), .B(u2_u0_b2_last_row_12_), .Y(u2_u0__abc_74955_new_n565_));
OR2X2 OR2X2_2569 ( .A(u2_u0__abc_74955_new_n567_), .B(row_adr_10_bF_buf2_), .Y(u2_u0__abc_74955_new_n568_));
OR2X2 OR2X2_257 ( .A(u0__abc_76628_new_n1197__bF_buf5), .B(u0_tms0_12_), .Y(u0__abc_76628_new_n1486_));
OR2X2 OR2X2_2570 ( .A(u2_u0__abc_74955_new_n189_), .B(u2_u0_b2_last_row_10_), .Y(u2_u0__abc_74955_new_n569_));
OR2X2 OR2X2_2571 ( .A(u2_u0__abc_74955_new_n169_), .B(u2_u0_b2_last_row_6_), .Y(u2_u0__abc_74955_new_n572_));
OR2X2 OR2X2_2572 ( .A(u2_u0__abc_74955_new_n573_), .B(row_adr_4_bF_buf2_), .Y(u2_u0__abc_74955_new_n574_));
OR2X2 OR2X2_2573 ( .A(u2_u0__abc_74955_new_n164_), .B(u2_u0_b2_last_row_5_), .Y(u2_u0__abc_74955_new_n576_));
OR2X2 OR2X2_2574 ( .A(u2_u0__abc_74955_new_n577_), .B(row_adr_5_bF_buf2_), .Y(u2_u0__abc_74955_new_n578_));
OR2X2 OR2X2_2575 ( .A(u2_u0__abc_74955_new_n139_), .B(u2_u0_b2_last_row_0_), .Y(u2_u0__abc_74955_new_n581_));
OR2X2 OR2X2_2576 ( .A(u2_u0__abc_74955_new_n582_), .B(row_adr_0_bF_buf2_), .Y(u2_u0__abc_74955_new_n583_));
OR2X2 OR2X2_2577 ( .A(u2_u0__abc_74955_new_n585_), .B(row_adr_1_bF_buf2_), .Y(u2_u0__abc_74955_new_n586_));
OR2X2 OR2X2_2578 ( .A(u2_u0__abc_74955_new_n526_), .B(u2_u0__abc_74955_new_n591_), .Y(u2_u0__abc_74955_new_n592_));
OR2X2 OR2X2_2579 ( .A(u2_u0__abc_74955_new_n461_), .B(u2_u0__abc_74955_new_n592_), .Y(u2_row_same_0));
OR2X2 OR2X2_258 ( .A(u0__abc_76628_new_n1488_), .B(u0__abc_76628_new_n1466_), .Y(u0__0sp_tms_31_0__12_));
OR2X2 OR2X2_2580 ( .A(u2_u0__abc_74955_new_n594_), .B(u2_u0__abc_74955_new_n595_), .Y(u2_u0__abc_74955_new_n596_));
OR2X2 OR2X2_2581 ( .A(u2_u0__abc_74955_new_n597_), .B(u2_u0__abc_74955_new_n598_), .Y(u2_u0__abc_74955_new_n599_));
OR2X2 OR2X2_2582 ( .A(u2_u0__abc_74955_new_n599_), .B(u2_u0__abc_74955_new_n596_), .Y(u2_bank_open_0));
OR2X2 OR2X2_2583 ( .A(u2_u0__abc_74955_new_n602_), .B(u2_u0__abc_74955_new_n601_), .Y(u2_u0__abc_74955_new_n603_));
OR2X2 OR2X2_2584 ( .A(u2_u0__abc_74955_new_n606_), .B(u2_u0__abc_74955_new_n290_), .Y(u2_u0__0bank2_open_0_0_));
OR2X2 OR2X2_2585 ( .A(u2_u0__abc_74955_new_n611_), .B(u2_u0__abc_74955_new_n137__bF_buf3), .Y(u2_u0__0bank3_open_0_0_));
OR2X2 OR2X2_2586 ( .A(u2_u0__abc_74955_new_n616_), .B(u2_u0__abc_74955_new_n601_), .Y(u2_u0__abc_74955_new_n617_));
OR2X2 OR2X2_2587 ( .A(u2_u0__abc_74955_new_n619_), .B(u2_u0__abc_74955_new_n248_), .Y(u2_u0__0bank1_open_0_0_));
OR2X2 OR2X2_2588 ( .A(u2_u0__abc_74955_new_n621_), .B(u2_u0__abc_74955_new_n601_), .Y(u2_u0__abc_74955_new_n622_));
OR2X2 OR2X2_2589 ( .A(u2_u0__abc_74955_new_n624_), .B(u2_u0__abc_74955_new_n206_), .Y(u2_u0__0bank0_open_0_0_));
OR2X2 OR2X2_259 ( .A(u0__abc_76628_new_n1177__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n1492_));
OR2X2 OR2X2_2590 ( .A(u2_u1__abc_74955_new_n137__bF_buf4), .B(u2_u1_b3_last_row_0_), .Y(u2_u1__abc_74955_new_n138_));
OR2X2 OR2X2_2591 ( .A(u2_u1__abc_74955_new_n137__bF_buf2), .B(u2_u1_b3_last_row_1_), .Y(u2_u1__abc_74955_new_n143_));
OR2X2 OR2X2_2592 ( .A(u2_u1__abc_74955_new_n137__bF_buf0), .B(u2_u1_b3_last_row_2_), .Y(u2_u1__abc_74955_new_n148_));
OR2X2 OR2X2_2593 ( .A(u2_u1__abc_74955_new_n137__bF_buf3), .B(u2_u1_b3_last_row_3_), .Y(u2_u1__abc_74955_new_n153_));
OR2X2 OR2X2_2594 ( .A(u2_u1__abc_74955_new_n137__bF_buf1), .B(u2_u1_b3_last_row_4_), .Y(u2_u1__abc_74955_new_n158_));
OR2X2 OR2X2_2595 ( .A(u2_u1__abc_74955_new_n137__bF_buf4), .B(u2_u1_b3_last_row_5_), .Y(u2_u1__abc_74955_new_n163_));
OR2X2 OR2X2_2596 ( .A(u2_u1__abc_74955_new_n137__bF_buf2), .B(u2_u1_b3_last_row_6_), .Y(u2_u1__abc_74955_new_n168_));
OR2X2 OR2X2_2597 ( .A(u2_u1__abc_74955_new_n137__bF_buf0), .B(u2_u1_b3_last_row_7_), .Y(u2_u1__abc_74955_new_n173_));
OR2X2 OR2X2_2598 ( .A(u2_u1__abc_74955_new_n137__bF_buf3), .B(u2_u1_b3_last_row_8_), .Y(u2_u1__abc_74955_new_n178_));
OR2X2 OR2X2_2599 ( .A(u2_u1__abc_74955_new_n137__bF_buf1), .B(u2_u1_b3_last_row_9_), .Y(u2_u1__abc_74955_new_n183_));
OR2X2 OR2X2_26 ( .A(_abc_85006_new_n245_), .B(cs_need_rfr_5_), .Y(_abc_85006_new_n276_));
OR2X2 OR2X2_260 ( .A(spec_req_cs_6_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1493_));
OR2X2 OR2X2_2600 ( .A(u2_u1__abc_74955_new_n137__bF_buf4), .B(u2_u1_b3_last_row_10_), .Y(u2_u1__abc_74955_new_n188_));
OR2X2 OR2X2_2601 ( .A(u2_u1__abc_74955_new_n137__bF_buf2), .B(u2_u1_b3_last_row_11_), .Y(u2_u1__abc_74955_new_n193_));
OR2X2 OR2X2_2602 ( .A(u2_u1__abc_74955_new_n137__bF_buf0), .B(u2_u1_b3_last_row_12_), .Y(u2_u1__abc_74955_new_n198_));
OR2X2 OR2X2_2603 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_0_), .Y(u2_u1__abc_74955_new_n207_));
OR2X2 OR2X2_2604 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_0_bF_buf0_), .Y(u2_u1__abc_74955_new_n209_));
OR2X2 OR2X2_2605 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_1_), .Y(u2_u1__abc_74955_new_n211_));
OR2X2 OR2X2_2606 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_1_bF_buf0_), .Y(u2_u1__abc_74955_new_n212_));
OR2X2 OR2X2_2607 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_2_), .Y(u2_u1__abc_74955_new_n214_));
OR2X2 OR2X2_2608 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_2_bF_buf0_), .Y(u2_u1__abc_74955_new_n215_));
OR2X2 OR2X2_2609 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_3_), .Y(u2_u1__abc_74955_new_n217_));
OR2X2 OR2X2_261 ( .A(u0__abc_76628_new_n1495_), .B(u0__abc_76628_new_n1491_), .Y(u0__abc_76628_new_n1496_));
OR2X2 OR2X2_2610 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_3_bF_buf0_), .Y(u2_u1__abc_74955_new_n218_));
OR2X2 OR2X2_2611 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_4_), .Y(u2_u1__abc_74955_new_n220_));
OR2X2 OR2X2_2612 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_4_bF_buf0_), .Y(u2_u1__abc_74955_new_n221_));
OR2X2 OR2X2_2613 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_5_), .Y(u2_u1__abc_74955_new_n223_));
OR2X2 OR2X2_2614 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_5_bF_buf0_), .Y(u2_u1__abc_74955_new_n224_));
OR2X2 OR2X2_2615 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_6_), .Y(u2_u1__abc_74955_new_n226_));
OR2X2 OR2X2_2616 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_6_bF_buf0_), .Y(u2_u1__abc_74955_new_n227_));
OR2X2 OR2X2_2617 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_7_), .Y(u2_u1__abc_74955_new_n229_));
OR2X2 OR2X2_2618 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_7_bF_buf0_), .Y(u2_u1__abc_74955_new_n230_));
OR2X2 OR2X2_2619 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_8_), .Y(u2_u1__abc_74955_new_n232_));
OR2X2 OR2X2_262 ( .A(u0__abc_76628_new_n1497_), .B(u0__abc_76628_new_n1498_), .Y(u0__abc_76628_new_n1499_));
OR2X2 OR2X2_2620 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_8_bF_buf0_), .Y(u2_u1__abc_74955_new_n233_));
OR2X2 OR2X2_2621 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_9_), .Y(u2_u1__abc_74955_new_n235_));
OR2X2 OR2X2_2622 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_9_bF_buf0_), .Y(u2_u1__abc_74955_new_n236_));
OR2X2 OR2X2_2623 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_10_), .Y(u2_u1__abc_74955_new_n238_));
OR2X2 OR2X2_2624 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_10_bF_buf0_), .Y(u2_u1__abc_74955_new_n239_));
OR2X2 OR2X2_2625 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_11_), .Y(u2_u1__abc_74955_new_n241_));
OR2X2 OR2X2_2626 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_11_bF_buf0_), .Y(u2_u1__abc_74955_new_n242_));
OR2X2 OR2X2_2627 ( .A(u2_u1__abc_74955_new_n206_), .B(u2_u1_b0_last_row_12_), .Y(u2_u1__abc_74955_new_n244_));
OR2X2 OR2X2_2628 ( .A(u2_u1__abc_74955_new_n208_), .B(row_adr_12_bF_buf0_), .Y(u2_u1__abc_74955_new_n245_));
OR2X2 OR2X2_2629 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_0_), .Y(u2_u1__abc_74955_new_n249_));
OR2X2 OR2X2_263 ( .A(u0__abc_76628_new_n1500_), .B(u0__abc_76628_new_n1501_), .Y(u0__abc_76628_new_n1502_));
OR2X2 OR2X2_2630 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_0_bF_buf3_), .Y(u2_u1__abc_74955_new_n251_));
OR2X2 OR2X2_2631 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_1_), .Y(u2_u1__abc_74955_new_n253_));
OR2X2 OR2X2_2632 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_1_bF_buf3_), .Y(u2_u1__abc_74955_new_n254_));
OR2X2 OR2X2_2633 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_2_), .Y(u2_u1__abc_74955_new_n256_));
OR2X2 OR2X2_2634 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_2_bF_buf3_), .Y(u2_u1__abc_74955_new_n257_));
OR2X2 OR2X2_2635 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_3_), .Y(u2_u1__abc_74955_new_n259_));
OR2X2 OR2X2_2636 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_3_bF_buf3_), .Y(u2_u1__abc_74955_new_n260_));
OR2X2 OR2X2_2637 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_4_), .Y(u2_u1__abc_74955_new_n262_));
OR2X2 OR2X2_2638 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_4_bF_buf3_), .Y(u2_u1__abc_74955_new_n263_));
OR2X2 OR2X2_2639 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_5_), .Y(u2_u1__abc_74955_new_n265_));
OR2X2 OR2X2_264 ( .A(u0__abc_76628_new_n1503_), .B(u0__abc_76628_new_n1504_), .Y(u0__abc_76628_new_n1505_));
OR2X2 OR2X2_2640 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_5_bF_buf3_), .Y(u2_u1__abc_74955_new_n266_));
OR2X2 OR2X2_2641 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_6_), .Y(u2_u1__abc_74955_new_n268_));
OR2X2 OR2X2_2642 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_6_bF_buf3_), .Y(u2_u1__abc_74955_new_n269_));
OR2X2 OR2X2_2643 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_7_), .Y(u2_u1__abc_74955_new_n271_));
OR2X2 OR2X2_2644 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_7_bF_buf3_), .Y(u2_u1__abc_74955_new_n272_));
OR2X2 OR2X2_2645 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_8_), .Y(u2_u1__abc_74955_new_n274_));
OR2X2 OR2X2_2646 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_8_bF_buf3_), .Y(u2_u1__abc_74955_new_n275_));
OR2X2 OR2X2_2647 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_9_), .Y(u2_u1__abc_74955_new_n277_));
OR2X2 OR2X2_2648 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_9_bF_buf3_), .Y(u2_u1__abc_74955_new_n278_));
OR2X2 OR2X2_2649 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_10_), .Y(u2_u1__abc_74955_new_n280_));
OR2X2 OR2X2_265 ( .A(u0__abc_76628_new_n1507_), .B(spec_req_cs_0_bF_buf1_), .Y(u0__abc_76628_new_n1508_));
OR2X2 OR2X2_2650 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_10_bF_buf3_), .Y(u2_u1__abc_74955_new_n281_));
OR2X2 OR2X2_2651 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_11_), .Y(u2_u1__abc_74955_new_n283_));
OR2X2 OR2X2_2652 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_11_bF_buf3_), .Y(u2_u1__abc_74955_new_n284_));
OR2X2 OR2X2_2653 ( .A(u2_u1__abc_74955_new_n248_), .B(u2_u1_b1_last_row_12_), .Y(u2_u1__abc_74955_new_n286_));
OR2X2 OR2X2_2654 ( .A(u2_u1__abc_74955_new_n250_), .B(row_adr_12_bF_buf3_), .Y(u2_u1__abc_74955_new_n287_));
OR2X2 OR2X2_2655 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_0_), .Y(u2_u1__abc_74955_new_n291_));
OR2X2 OR2X2_2656 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_0_bF_buf2_), .Y(u2_u1__abc_74955_new_n293_));
OR2X2 OR2X2_2657 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_1_), .Y(u2_u1__abc_74955_new_n295_));
OR2X2 OR2X2_2658 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_1_bF_buf2_), .Y(u2_u1__abc_74955_new_n296_));
OR2X2 OR2X2_2659 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_2_), .Y(u2_u1__abc_74955_new_n298_));
OR2X2 OR2X2_266 ( .A(u0__abc_76628_new_n1506_), .B(u0__abc_76628_new_n1508_), .Y(u0__abc_76628_new_n1509_));
OR2X2 OR2X2_2660 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_2_bF_buf2_), .Y(u2_u1__abc_74955_new_n299_));
OR2X2 OR2X2_2661 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_3_), .Y(u2_u1__abc_74955_new_n301_));
OR2X2 OR2X2_2662 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_3_bF_buf2_), .Y(u2_u1__abc_74955_new_n302_));
OR2X2 OR2X2_2663 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_4_), .Y(u2_u1__abc_74955_new_n304_));
OR2X2 OR2X2_2664 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_4_bF_buf2_), .Y(u2_u1__abc_74955_new_n305_));
OR2X2 OR2X2_2665 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_5_), .Y(u2_u1__abc_74955_new_n307_));
OR2X2 OR2X2_2666 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_5_bF_buf2_), .Y(u2_u1__abc_74955_new_n308_));
OR2X2 OR2X2_2667 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_6_), .Y(u2_u1__abc_74955_new_n310_));
OR2X2 OR2X2_2668 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_6_bF_buf2_), .Y(u2_u1__abc_74955_new_n311_));
OR2X2 OR2X2_2669 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_7_), .Y(u2_u1__abc_74955_new_n313_));
OR2X2 OR2X2_267 ( .A(u0__abc_76628_new_n1197__bF_buf4), .B(u0_tms0_13_), .Y(u0__abc_76628_new_n1510_));
OR2X2 OR2X2_2670 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_7_bF_buf2_), .Y(u2_u1__abc_74955_new_n314_));
OR2X2 OR2X2_2671 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_8_), .Y(u2_u1__abc_74955_new_n316_));
OR2X2 OR2X2_2672 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_8_bF_buf2_), .Y(u2_u1__abc_74955_new_n317_));
OR2X2 OR2X2_2673 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_9_), .Y(u2_u1__abc_74955_new_n319_));
OR2X2 OR2X2_2674 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_9_bF_buf2_), .Y(u2_u1__abc_74955_new_n320_));
OR2X2 OR2X2_2675 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_10_), .Y(u2_u1__abc_74955_new_n322_));
OR2X2 OR2X2_2676 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_10_bF_buf2_), .Y(u2_u1__abc_74955_new_n323_));
OR2X2 OR2X2_2677 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_11_), .Y(u2_u1__abc_74955_new_n325_));
OR2X2 OR2X2_2678 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_11_bF_buf2_), .Y(u2_u1__abc_74955_new_n326_));
OR2X2 OR2X2_2679 ( .A(u2_u1__abc_74955_new_n290_), .B(u2_u1_b2_last_row_12_), .Y(u2_u1__abc_74955_new_n328_));
OR2X2 OR2X2_268 ( .A(u0__abc_76628_new_n1512_), .B(u0__abc_76628_new_n1490_), .Y(u0__0sp_tms_31_0__13_));
OR2X2 OR2X2_2680 ( .A(u2_u1__abc_74955_new_n292_), .B(row_adr_12_bF_buf2_), .Y(u2_u1__abc_74955_new_n329_));
OR2X2 OR2X2_2681 ( .A(u2_u1__abc_74955_new_n179_), .B(u2_u1_b3_last_row_8_), .Y(u2_u1__abc_74955_new_n331_));
OR2X2 OR2X2_2682 ( .A(u2_u1__abc_74955_new_n332_), .B(row_adr_9_bF_buf1_), .Y(u2_u1__abc_74955_new_n333_));
OR2X2 OR2X2_2683 ( .A(u2_u1__abc_74955_new_n334_), .B(row_adr_8_bF_buf1_), .Y(u2_u1__abc_74955_new_n335_));
OR2X2 OR2X2_2684 ( .A(u2_u1__abc_74955_new_n184_), .B(u2_u1_b3_last_row_9_), .Y(u2_u1__abc_74955_new_n338_));
OR2X2 OR2X2_2685 ( .A(u2_u1__abc_74955_new_n339_), .B(row_adr_11_bF_buf1_), .Y(u2_u1__abc_74955_new_n340_));
OR2X2 OR2X2_2686 ( .A(u2_u1__abc_74955_new_n342_), .B(row_adr_4_bF_buf1_), .Y(u2_u1__abc_74955_new_n343_));
OR2X2 OR2X2_2687 ( .A(u2_u1__abc_74955_new_n194_), .B(u2_u1_b3_last_row_11_), .Y(u2_u1__abc_74955_new_n344_));
OR2X2 OR2X2_2688 ( .A(u2_u1__abc_74955_new_n349_), .B(u2_u1__abc_74955_new_n350_), .Y(u2_u1__abc_74955_new_n351_));
OR2X2 OR2X2_2689 ( .A(u2_u1__abc_74955_new_n144_), .B(u2_u1_b3_last_row_1_), .Y(u2_u1__abc_74955_new_n352_));
OR2X2 OR2X2_269 ( .A(u0__abc_76628_new_n1177__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n1516_));
OR2X2 OR2X2_2690 ( .A(u2_u1__abc_74955_new_n355_), .B(row_adr_7_bF_buf1_), .Y(u2_u1__abc_74955_new_n356_));
OR2X2 OR2X2_2691 ( .A(u2_u1__abc_74955_new_n174_), .B(u2_u1_b3_last_row_7_), .Y(u2_u1__abc_74955_new_n357_));
OR2X2 OR2X2_2692 ( .A(u2_u1__abc_74955_new_n359_), .B(row_adr_5_bF_buf1_), .Y(u2_u1__abc_74955_new_n360_));
OR2X2 OR2X2_2693 ( .A(u2_u1__abc_74955_new_n164_), .B(u2_u1_b3_last_row_5_), .Y(u2_u1__abc_74955_new_n361_));
OR2X2 OR2X2_2694 ( .A(u2_u1__abc_74955_new_n199_), .B(u2_u1_b3_last_row_12_), .Y(u2_u1__abc_74955_new_n366_));
OR2X2 OR2X2_2695 ( .A(u2_u1__abc_74955_new_n367_), .B(row_adr_12_bF_buf1_), .Y(u2_u1__abc_74955_new_n368_));
OR2X2 OR2X2_2696 ( .A(u2_u1__abc_74955_new_n189_), .B(u2_u1_b3_last_row_10_), .Y(u2_u1__abc_74955_new_n370_));
OR2X2 OR2X2_2697 ( .A(u2_u1__abc_74955_new_n371_), .B(row_adr_10_bF_buf1_), .Y(u2_u1__abc_74955_new_n372_));
OR2X2 OR2X2_2698 ( .A(u2_u1__abc_74955_new_n375_), .B(row_adr_3_bF_buf1_), .Y(u2_u1__abc_74955_new_n376_));
OR2X2 OR2X2_2699 ( .A(u2_u1__abc_74955_new_n154_), .B(u2_u1_b3_last_row_3_), .Y(u2_u1__abc_74955_new_n377_));
OR2X2 OR2X2_27 ( .A(_abc_85006_new_n240__bF_buf5), .B(spec_req_cs_6_bF_buf5_), .Y(_abc_85006_new_n278_));
OR2X2 OR2X2_270 ( .A(spec_req_cs_6_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1517_));
OR2X2 OR2X2_2700 ( .A(u2_u1__abc_74955_new_n379_), .B(row_adr_1_bF_buf1_), .Y(u2_u1__abc_74955_new_n380_));
OR2X2 OR2X2_2701 ( .A(u2_u1__abc_74955_new_n149_), .B(u2_u1_b3_last_row_2_), .Y(u2_u1__abc_74955_new_n381_));
OR2X2 OR2X2_2702 ( .A(u2_u1__abc_74955_new_n159_), .B(u2_u1_b3_last_row_4_), .Y(u2_u1__abc_74955_new_n384_));
OR2X2 OR2X2_2703 ( .A(u2_u1__abc_74955_new_n385_), .B(row_adr_6_bF_buf1_), .Y(u2_u1__abc_74955_new_n386_));
OR2X2 OR2X2_2704 ( .A(u2_u1__abc_74955_new_n388_), .B(row_adr_2_bF_buf1_), .Y(u2_u1__abc_74955_new_n389_));
OR2X2 OR2X2_2705 ( .A(u2_u1__abc_74955_new_n169_), .B(u2_u1_b3_last_row_6_), .Y(u2_u1__abc_74955_new_n390_));
OR2X2 OR2X2_2706 ( .A(u2_u1__abc_74955_new_n144_), .B(u2_u1_b1_last_row_1_), .Y(u2_u1__abc_74955_new_n396_));
OR2X2 OR2X2_2707 ( .A(u2_u1__abc_74955_new_n139_), .B(u2_u1_b1_last_row_0_), .Y(u2_u1__abc_74955_new_n397_));
OR2X2 OR2X2_2708 ( .A(u2_u1__abc_74955_new_n399_), .B(row_adr_0_bF_buf0_), .Y(u2_u1__abc_74955_new_n400_));
OR2X2 OR2X2_2709 ( .A(u2_u1__abc_74955_new_n159_), .B(u2_u1_b1_last_row_4_), .Y(u2_u1__abc_74955_new_n402_));
OR2X2 OR2X2_271 ( .A(u0__abc_76628_new_n1519_), .B(u0__abc_76628_new_n1515_), .Y(u0__abc_76628_new_n1520_));
OR2X2 OR2X2_2710 ( .A(u2_u1__abc_74955_new_n403_), .B(row_adr_4_bF_buf0_), .Y(u2_u1__abc_74955_new_n404_));
OR2X2 OR2X2_2711 ( .A(u2_u1__abc_74955_new_n164_), .B(u2_u1_b1_last_row_5_), .Y(u2_u1__abc_74955_new_n406_));
OR2X2 OR2X2_2712 ( .A(u2_u1__abc_74955_new_n407_), .B(row_adr_3_bF_buf0_), .Y(u2_u1__abc_74955_new_n408_));
OR2X2 OR2X2_2713 ( .A(u2_u1__abc_74955_new_n179_), .B(u2_u1_b1_last_row_8_), .Y(u2_u1__abc_74955_new_n412_));
OR2X2 OR2X2_2714 ( .A(u2_u1__abc_74955_new_n413_), .B(row_adr_8_bF_buf0_), .Y(u2_u1__abc_74955_new_n414_));
OR2X2 OR2X2_2715 ( .A(u2_u1__abc_74955_new_n169_), .B(u2_u1_b1_last_row_6_), .Y(u2_u1__abc_74955_new_n416_));
OR2X2 OR2X2_2716 ( .A(u2_u1__abc_74955_new_n417_), .B(row_adr_6_bF_buf0_), .Y(u2_u1__abc_74955_new_n418_));
OR2X2 OR2X2_2717 ( .A(u2_u1__abc_74955_new_n199_), .B(u2_u1_b1_last_row_12_), .Y(u2_u1__abc_74955_new_n421_));
OR2X2 OR2X2_2718 ( .A(u2_u1__abc_74955_new_n422_), .B(row_adr_12_bF_buf0_), .Y(u2_u1__abc_74955_new_n423_));
OR2X2 OR2X2_2719 ( .A(u2_u1__abc_74955_new_n425_), .B(row_adr_11_bF_buf0_), .Y(u2_u1__abc_74955_new_n426_));
OR2X2 OR2X2_272 ( .A(u0__abc_76628_new_n1521_), .B(u0__abc_76628_new_n1522_), .Y(u0__abc_76628_new_n1523_));
OR2X2 OR2X2_2720 ( .A(u2_u1__abc_74955_new_n431_), .B(row_adr_2_bF_buf0_), .Y(u2_u1__abc_74955_new_n432_));
OR2X2 OR2X2_2721 ( .A(u2_u1__abc_74955_new_n149_), .B(u2_u1_b1_last_row_2_), .Y(u2_u1__abc_74955_new_n433_));
OR2X2 OR2X2_2722 ( .A(u2_u1__abc_74955_new_n435_), .B(row_adr_1_bF_buf0_), .Y(u2_u1__abc_74955_new_n436_));
OR2X2 OR2X2_2723 ( .A(u2_u1__abc_74955_new_n154_), .B(u2_u1_b1_last_row_3_), .Y(u2_u1__abc_74955_new_n437_));
OR2X2 OR2X2_2724 ( .A(u2_u1__abc_74955_new_n440_), .B(row_adr_10_bF_buf0_), .Y(u2_u1__abc_74955_new_n441_));
OR2X2 OR2X2_2725 ( .A(u2_u1__abc_74955_new_n189_), .B(u2_u1_b1_last_row_10_), .Y(u2_u1__abc_74955_new_n442_));
OR2X2 OR2X2_2726 ( .A(u2_u1__abc_74955_new_n444_), .B(row_adr_9_bF_buf0_), .Y(u2_u1__abc_74955_new_n445_));
OR2X2 OR2X2_2727 ( .A(u2_u1__abc_74955_new_n194_), .B(u2_u1_b1_last_row_11_), .Y(u2_u1__abc_74955_new_n446_));
OR2X2 OR2X2_2728 ( .A(u2_u1__abc_74955_new_n184_), .B(u2_u1_b1_last_row_9_), .Y(u2_u1__abc_74955_new_n449_));
OR2X2 OR2X2_2729 ( .A(u2_u1__abc_74955_new_n450_), .B(row_adr_7_bF_buf0_), .Y(u2_u1__abc_74955_new_n451_));
OR2X2 OR2X2_273 ( .A(u0__abc_76628_new_n1524_), .B(u0__abc_76628_new_n1525_), .Y(u0__abc_76628_new_n1526_));
OR2X2 OR2X2_2730 ( .A(u2_u1__abc_74955_new_n174_), .B(u2_u1_b1_last_row_7_), .Y(u2_u1__abc_74955_new_n453_));
OR2X2 OR2X2_2731 ( .A(u2_u1__abc_74955_new_n454_), .B(row_adr_5_bF_buf0_), .Y(u2_u1__abc_74955_new_n455_));
OR2X2 OR2X2_2732 ( .A(u2_u1__abc_74955_new_n395_), .B(u2_u1__abc_74955_new_n460_), .Y(u2_u1__abc_74955_new_n461_));
OR2X2 OR2X2_2733 ( .A(u2_u1__abc_74955_new_n462_), .B(row_adr_9_bF_buf3_), .Y(u2_u1__abc_74955_new_n463_));
OR2X2 OR2X2_2734 ( .A(u2_u1__abc_74955_new_n194_), .B(u2_u1_b0_last_row_11_), .Y(u2_u1__abc_74955_new_n464_));
OR2X2 OR2X2_2735 ( .A(u2_u1__abc_74955_new_n184_), .B(u2_u1_b0_last_row_9_), .Y(u2_u1__abc_74955_new_n465_));
OR2X2 OR2X2_2736 ( .A(u2_u1__abc_74955_new_n154_), .B(u2_u1_b0_last_row_3_), .Y(u2_u1__abc_74955_new_n468_));
OR2X2 OR2X2_2737 ( .A(u2_u1__abc_74955_new_n469_), .B(row_adr_12_bF_buf3_), .Y(u2_u1__abc_74955_new_n470_));
OR2X2 OR2X2_2738 ( .A(u2_u1__abc_74955_new_n472_), .B(row_adr_3_bF_buf3_), .Y(u2_u1__abc_74955_new_n473_));
OR2X2 OR2X2_2739 ( .A(u2_u1__abc_74955_new_n179_), .B(u2_u1_b0_last_row_8_), .Y(u2_u1__abc_74955_new_n474_));
OR2X2 OR2X2_274 ( .A(u0__abc_76628_new_n1527_), .B(u0__abc_76628_new_n1528_), .Y(u0__abc_76628_new_n1529_));
OR2X2 OR2X2_2740 ( .A(u2_u1__abc_74955_new_n477_), .B(row_adr_2_bF_buf3_), .Y(u2_u1__abc_74955_new_n478_));
OR2X2 OR2X2_2741 ( .A(u2_u1__abc_74955_new_n479_), .B(row_adr_6_bF_buf3_), .Y(u2_u1__abc_74955_new_n480_));
OR2X2 OR2X2_2742 ( .A(u2_u1__abc_74955_new_n169_), .B(u2_u1_b0_last_row_6_), .Y(u2_u1__abc_74955_new_n482_));
OR2X2 OR2X2_2743 ( .A(u2_u1__abc_74955_new_n199_), .B(u2_u1_b0_last_row_12_), .Y(u2_u1__abc_74955_new_n483_));
OR2X2 OR2X2_2744 ( .A(u2_u1__abc_74955_new_n489_), .B(u2_u1__abc_74955_new_n490_), .Y(u2_u1__abc_74955_new_n491_));
OR2X2 OR2X2_2745 ( .A(u2_u1__abc_74955_new_n492_), .B(row_adr_1_bF_buf3_), .Y(u2_u1__abc_74955_new_n493_));
OR2X2 OR2X2_2746 ( .A(u2_u1__abc_74955_new_n144_), .B(u2_u1_b0_last_row_1_), .Y(u2_u1__abc_74955_new_n494_));
OR2X2 OR2X2_2747 ( .A(u2_u1__abc_74955_new_n164_), .B(u2_u1_b0_last_row_5_), .Y(u2_u1__abc_74955_new_n497_));
OR2X2 OR2X2_2748 ( .A(u2_u1__abc_74955_new_n498_), .B(row_adr_5_bF_buf3_), .Y(u2_u1__abc_74955_new_n499_));
OR2X2 OR2X2_2749 ( .A(u2_u1__abc_74955_new_n501_), .B(row_adr_8_bF_buf3_), .Y(u2_u1__abc_74955_new_n502_));
OR2X2 OR2X2_275 ( .A(u0__abc_76628_new_n1531_), .B(spec_req_cs_0_bF_buf0_), .Y(u0__abc_76628_new_n1532_));
OR2X2 OR2X2_2750 ( .A(u2_u1__abc_74955_new_n506_), .B(row_adr_4_bF_buf3_), .Y(u2_u1__abc_74955_new_n507_));
OR2X2 OR2X2_2751 ( .A(u2_u1__abc_74955_new_n508_), .B(row_adr_11_bF_buf3_), .Y(u2_u1__abc_74955_new_n509_));
OR2X2 OR2X2_2752 ( .A(u2_u1__abc_74955_new_n149_), .B(u2_u1_b0_last_row_2_), .Y(u2_u1__abc_74955_new_n511_));
OR2X2 OR2X2_2753 ( .A(u2_u1__abc_74955_new_n159_), .B(u2_u1_b0_last_row_4_), .Y(u2_u1__abc_74955_new_n512_));
OR2X2 OR2X2_2754 ( .A(u2_u1__abc_74955_new_n174_), .B(u2_u1_b0_last_row_7_), .Y(u2_u1__abc_74955_new_n515_));
OR2X2 OR2X2_2755 ( .A(u2_u1__abc_74955_new_n516_), .B(row_adr_7_bF_buf3_), .Y(u2_u1__abc_74955_new_n517_));
OR2X2 OR2X2_2756 ( .A(u2_u1__abc_74955_new_n189_), .B(u2_u1_b0_last_row_10_), .Y(u2_u1__abc_74955_new_n519_));
OR2X2 OR2X2_2757 ( .A(u2_u1__abc_74955_new_n520_), .B(row_adr_10_bF_buf3_), .Y(u2_u1__abc_74955_new_n521_));
OR2X2 OR2X2_2758 ( .A(u2_u1__abc_74955_new_n527_), .B(row_adr_8_bF_buf2_), .Y(u2_u1__abc_74955_new_n528_));
OR2X2 OR2X2_2759 ( .A(u2_u1__abc_74955_new_n184_), .B(u2_u1_b2_last_row_9_), .Y(u2_u1__abc_74955_new_n529_));
OR2X2 OR2X2_276 ( .A(u0__abc_76628_new_n1530_), .B(u0__abc_76628_new_n1532_), .Y(u0__abc_76628_new_n1533_));
OR2X2 OR2X2_2760 ( .A(u2_u1__abc_74955_new_n179_), .B(u2_u1_b2_last_row_8_), .Y(u2_u1__abc_74955_new_n530_));
OR2X2 OR2X2_2761 ( .A(u2_u1__abc_74955_new_n533_), .B(row_adr_9_bF_buf2_), .Y(u2_u1__abc_74955_new_n534_));
OR2X2 OR2X2_2762 ( .A(u2_u1__abc_74955_new_n194_), .B(u2_u1_b2_last_row_11_), .Y(u2_u1__abc_74955_new_n535_));
OR2X2 OR2X2_2763 ( .A(u2_u1__abc_74955_new_n537_), .B(row_adr_11_bF_buf2_), .Y(u2_u1__abc_74955_new_n538_));
OR2X2 OR2X2_2764 ( .A(u2_u1__abc_74955_new_n159_), .B(u2_u1_b2_last_row_4_), .Y(u2_u1__abc_74955_new_n539_));
OR2X2 OR2X2_2765 ( .A(u2_u1__abc_74955_new_n174_), .B(u2_u1_b2_last_row_7_), .Y(u2_u1__abc_74955_new_n543_));
OR2X2 OR2X2_2766 ( .A(u2_u1__abc_74955_new_n544_), .B(row_adr_7_bF_buf2_), .Y(u2_u1__abc_74955_new_n545_));
OR2X2 OR2X2_2767 ( .A(u2_u1__abc_74955_new_n149_), .B(u2_u1_b2_last_row_2_), .Y(u2_u1__abc_74955_new_n547_));
OR2X2 OR2X2_2768 ( .A(u2_u1__abc_74955_new_n548_), .B(row_adr_6_bF_buf2_), .Y(u2_u1__abc_74955_new_n549_));
OR2X2 OR2X2_2769 ( .A(u2_u1__abc_74955_new_n154_), .B(u2_u1_b2_last_row_3_), .Y(u2_u1__abc_74955_new_n552_));
OR2X2 OR2X2_277 ( .A(u0__abc_76628_new_n1197__bF_buf3), .B(u0_tms0_14_), .Y(u0__abc_76628_new_n1534_));
OR2X2 OR2X2_2770 ( .A(u2_u1__abc_74955_new_n553_), .B(row_adr_3_bF_buf2_), .Y(u2_u1__abc_74955_new_n554_));
OR2X2 OR2X2_2771 ( .A(u2_u1__abc_74955_new_n144_), .B(u2_u1_b2_last_row_1_), .Y(u2_u1__abc_74955_new_n556_));
OR2X2 OR2X2_2772 ( .A(u2_u1__abc_74955_new_n557_), .B(row_adr_2_bF_buf2_), .Y(u2_u1__abc_74955_new_n558_));
OR2X2 OR2X2_2773 ( .A(u2_u1__abc_74955_new_n563_), .B(row_adr_12_bF_buf2_), .Y(u2_u1__abc_74955_new_n564_));
OR2X2 OR2X2_2774 ( .A(u2_u1__abc_74955_new_n199_), .B(u2_u1_b2_last_row_12_), .Y(u2_u1__abc_74955_new_n565_));
OR2X2 OR2X2_2775 ( .A(u2_u1__abc_74955_new_n567_), .B(row_adr_10_bF_buf2_), .Y(u2_u1__abc_74955_new_n568_));
OR2X2 OR2X2_2776 ( .A(u2_u1__abc_74955_new_n189_), .B(u2_u1_b2_last_row_10_), .Y(u2_u1__abc_74955_new_n569_));
OR2X2 OR2X2_2777 ( .A(u2_u1__abc_74955_new_n169_), .B(u2_u1_b2_last_row_6_), .Y(u2_u1__abc_74955_new_n572_));
OR2X2 OR2X2_2778 ( .A(u2_u1__abc_74955_new_n573_), .B(row_adr_4_bF_buf2_), .Y(u2_u1__abc_74955_new_n574_));
OR2X2 OR2X2_2779 ( .A(u2_u1__abc_74955_new_n164_), .B(u2_u1_b2_last_row_5_), .Y(u2_u1__abc_74955_new_n576_));
OR2X2 OR2X2_278 ( .A(u0__abc_76628_new_n1536_), .B(u0__abc_76628_new_n1514_), .Y(u0__0sp_tms_31_0__14_));
OR2X2 OR2X2_2780 ( .A(u2_u1__abc_74955_new_n577_), .B(row_adr_5_bF_buf2_), .Y(u2_u1__abc_74955_new_n578_));
OR2X2 OR2X2_2781 ( .A(u2_u1__abc_74955_new_n139_), .B(u2_u1_b2_last_row_0_), .Y(u2_u1__abc_74955_new_n581_));
OR2X2 OR2X2_2782 ( .A(u2_u1__abc_74955_new_n582_), .B(row_adr_0_bF_buf2_), .Y(u2_u1__abc_74955_new_n583_));
OR2X2 OR2X2_2783 ( .A(u2_u1__abc_74955_new_n585_), .B(row_adr_1_bF_buf2_), .Y(u2_u1__abc_74955_new_n586_));
OR2X2 OR2X2_2784 ( .A(u2_u1__abc_74955_new_n526_), .B(u2_u1__abc_74955_new_n591_), .Y(u2_u1__abc_74955_new_n592_));
OR2X2 OR2X2_2785 ( .A(u2_u1__abc_74955_new_n461_), .B(u2_u1__abc_74955_new_n592_), .Y(u2_row_same_1));
OR2X2 OR2X2_2786 ( .A(u2_u1__abc_74955_new_n594_), .B(u2_u1__abc_74955_new_n595_), .Y(u2_u1__abc_74955_new_n596_));
OR2X2 OR2X2_2787 ( .A(u2_u1__abc_74955_new_n597_), .B(u2_u1__abc_74955_new_n598_), .Y(u2_u1__abc_74955_new_n599_));
OR2X2 OR2X2_2788 ( .A(u2_u1__abc_74955_new_n599_), .B(u2_u1__abc_74955_new_n596_), .Y(u2_bank_open_1));
OR2X2 OR2X2_2789 ( .A(u2_u1__abc_74955_new_n602_), .B(u2_u1__abc_74955_new_n601_), .Y(u2_u1__abc_74955_new_n603_));
OR2X2 OR2X2_279 ( .A(u0__abc_76628_new_n1177__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n1540_));
OR2X2 OR2X2_2790 ( .A(u2_u1__abc_74955_new_n606_), .B(u2_u1__abc_74955_new_n290_), .Y(u2_u1__0bank2_open_0_0_));
OR2X2 OR2X2_2791 ( .A(u2_u1__abc_74955_new_n611_), .B(u2_u1__abc_74955_new_n137__bF_buf3), .Y(u2_u1__0bank3_open_0_0_));
OR2X2 OR2X2_2792 ( .A(u2_u1__abc_74955_new_n616_), .B(u2_u1__abc_74955_new_n601_), .Y(u2_u1__abc_74955_new_n617_));
OR2X2 OR2X2_2793 ( .A(u2_u1__abc_74955_new_n619_), .B(u2_u1__abc_74955_new_n248_), .Y(u2_u1__0bank1_open_0_0_));
OR2X2 OR2X2_2794 ( .A(u2_u1__abc_74955_new_n621_), .B(u2_u1__abc_74955_new_n601_), .Y(u2_u1__abc_74955_new_n622_));
OR2X2 OR2X2_2795 ( .A(u2_u1__abc_74955_new_n624_), .B(u2_u1__abc_74955_new_n206_), .Y(u2_u1__0bank0_open_0_0_));
OR2X2 OR2X2_2796 ( .A(csc_2_), .B(csc_3_), .Y(u3__abc_74070_new_n275_));
OR2X2 OR2X2_2797 ( .A(csc_1_), .B(mem_ack_r), .Y(u3__abc_74070_new_n276_));
OR2X2 OR2X2_2798 ( .A(u3__abc_74070_new_n275__bF_buf4), .B(u3__abc_74070_new_n276_), .Y(u3__abc_74070_new_n277_));
OR2X2 OR2X2_2799 ( .A(u3__abc_74070_new_n277__bF_buf5), .B(mc_dp_od_0_), .Y(u3__abc_74070_new_n278_));
OR2X2 OR2X2_28 ( .A(lmr_sel_bF_buf0), .B(cs_6_), .Y(_abc_85006_new_n279_));
OR2X2 OR2X2_280 ( .A(spec_req_cs_6_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1541_));
OR2X2 OR2X2_2800 ( .A(\wb_data_i[3] ), .B(\wb_data_i[2] ), .Y(u3__abc_74070_new_n280_));
OR2X2 OR2X2_2801 ( .A(u3__abc_74070_new_n285_), .B(\wb_data_i[0] ), .Y(u3__abc_74070_new_n286_));
OR2X2 OR2X2_2802 ( .A(u3__abc_74070_new_n287_), .B(\wb_data_i[1] ), .Y(u3__abc_74070_new_n288_));
OR2X2 OR2X2_2803 ( .A(u3__abc_74070_new_n284_), .B(u3__abc_74070_new_n289_), .Y(u3__abc_74070_new_n292_));
OR2X2 OR2X2_2804 ( .A(\wb_data_i[7] ), .B(\wb_data_i[6] ), .Y(u3__abc_74070_new_n295_));
OR2X2 OR2X2_2805 ( .A(u3__abc_74070_new_n300_), .B(\wb_data_i[4] ), .Y(u3__abc_74070_new_n301_));
OR2X2 OR2X2_2806 ( .A(u3__abc_74070_new_n302_), .B(\wb_data_i[5] ), .Y(u3__abc_74070_new_n303_));
OR2X2 OR2X2_2807 ( .A(u3__abc_74070_new_n306_), .B(u3__abc_74070_new_n307_), .Y(u3__abc_74070_new_n308_));
OR2X2 OR2X2_2808 ( .A(u3__abc_74070_new_n294_), .B(u3__abc_74070_new_n309_), .Y(u3__abc_74070_new_n310_));
OR2X2 OR2X2_2809 ( .A(u3__abc_74070_new_n293_), .B(u3__abc_74070_new_n308_), .Y(u3__abc_74070_new_n311_));
OR2X2 OR2X2_281 ( .A(u0__abc_76628_new_n1543_), .B(u0__abc_76628_new_n1539_), .Y(u0__abc_76628_new_n1544_));
OR2X2 OR2X2_2810 ( .A(u3__abc_74070_new_n312_), .B(u3__abc_74070_new_n279__bF_buf5), .Y(u3__abc_74070_new_n313_));
OR2X2 OR2X2_2811 ( .A(u3__abc_74070_new_n277__bF_buf3), .B(mc_dp_od_1_), .Y(u3__abc_74070_new_n315_));
OR2X2 OR2X2_2812 ( .A(\wb_data_i[11] ), .B(\wb_data_i[10] ), .Y(u3__abc_74070_new_n316_));
OR2X2 OR2X2_2813 ( .A(u3__abc_74070_new_n320_), .B(\wb_data_i[8] ), .Y(u3__abc_74070_new_n321_));
OR2X2 OR2X2_2814 ( .A(u3__abc_74070_new_n322_), .B(\wb_data_i[9] ), .Y(u3__abc_74070_new_n323_));
OR2X2 OR2X2_2815 ( .A(u3__abc_74070_new_n325_), .B(u3__abc_74070_new_n319_), .Y(u3__abc_74070_new_n328_));
OR2X2 OR2X2_2816 ( .A(\wb_data_i[15] ), .B(\wb_data_i[14] ), .Y(u3__abc_74070_new_n331_));
OR2X2 OR2X2_2817 ( .A(u3__abc_74070_new_n336_), .B(\wb_data_i[12] ), .Y(u3__abc_74070_new_n337_));
OR2X2 OR2X2_2818 ( .A(u3__abc_74070_new_n338_), .B(\wb_data_i[13] ), .Y(u3__abc_74070_new_n339_));
OR2X2 OR2X2_2819 ( .A(u3__abc_74070_new_n342_), .B(u3__abc_74070_new_n343_), .Y(u3__abc_74070_new_n344_));
OR2X2 OR2X2_282 ( .A(u0__abc_76628_new_n1545_), .B(u0__abc_76628_new_n1546_), .Y(u0__abc_76628_new_n1547_));
OR2X2 OR2X2_2820 ( .A(u3__abc_74070_new_n330_), .B(u3__abc_74070_new_n345_), .Y(u3__abc_74070_new_n346_));
OR2X2 OR2X2_2821 ( .A(u3__abc_74070_new_n329_), .B(u3__abc_74070_new_n344_), .Y(u3__abc_74070_new_n347_));
OR2X2 OR2X2_2822 ( .A(u3__abc_74070_new_n348_), .B(u3__abc_74070_new_n279__bF_buf4), .Y(u3__abc_74070_new_n349_));
OR2X2 OR2X2_2823 ( .A(\wb_data_i[19] ), .B(\wb_data_i[18] ), .Y(u3__abc_74070_new_n351_));
OR2X2 OR2X2_2824 ( .A(u3__abc_74070_new_n355_), .B(\wb_data_i[16] ), .Y(u3__abc_74070_new_n356_));
OR2X2 OR2X2_2825 ( .A(u3__abc_74070_new_n357_), .B(\wb_data_i[17] ), .Y(u3__abc_74070_new_n358_));
OR2X2 OR2X2_2826 ( .A(u3__abc_74070_new_n360_), .B(u3__abc_74070_new_n354_), .Y(u3__abc_74070_new_n363_));
OR2X2 OR2X2_2827 ( .A(\wb_data_i[23] ), .B(\wb_data_i[22] ), .Y(u3__abc_74070_new_n365_));
OR2X2 OR2X2_2828 ( .A(u3__abc_74070_new_n370_), .B(\wb_data_i[20] ), .Y(u3__abc_74070_new_n371_));
OR2X2 OR2X2_2829 ( .A(u3__abc_74070_new_n372_), .B(\wb_data_i[21] ), .Y(u3__abc_74070_new_n373_));
OR2X2 OR2X2_283 ( .A(u0__abc_76628_new_n1548_), .B(u0__abc_76628_new_n1549_), .Y(u0__abc_76628_new_n1550_));
OR2X2 OR2X2_2830 ( .A(u3__abc_74070_new_n376_), .B(u3__abc_74070_new_n377_), .Y(u3__abc_74070_new_n378_));
OR2X2 OR2X2_2831 ( .A(u3__abc_74070_new_n382_), .B(u3__abc_74070_new_n380_), .Y(u3__abc_74070_new_n383_));
OR2X2 OR2X2_2832 ( .A(u3__abc_74070_new_n384_), .B(u3__abc_74070_new_n385_), .Y(u3__0mc_dp_o_3_0__2_));
OR2X2 OR2X2_2833 ( .A(\wb_data_i[27] ), .B(\wb_data_i[26] ), .Y(u3__abc_74070_new_n387_));
OR2X2 OR2X2_2834 ( .A(u3__abc_74070_new_n391_), .B(\wb_data_i[24] ), .Y(u3__abc_74070_new_n392_));
OR2X2 OR2X2_2835 ( .A(u3__abc_74070_new_n393_), .B(\wb_data_i[25] ), .Y(u3__abc_74070_new_n394_));
OR2X2 OR2X2_2836 ( .A(u3__abc_74070_new_n396_), .B(u3__abc_74070_new_n390_), .Y(u3__abc_74070_new_n399_));
OR2X2 OR2X2_2837 ( .A(\wb_data_i[31] ), .B(\wb_data_i[30] ), .Y(u3__abc_74070_new_n401_));
OR2X2 OR2X2_2838 ( .A(u3__abc_74070_new_n406_), .B(\wb_data_i[28] ), .Y(u3__abc_74070_new_n407_));
OR2X2 OR2X2_2839 ( .A(u3__abc_74070_new_n408_), .B(\wb_data_i[29] ), .Y(u3__abc_74070_new_n409_));
OR2X2 OR2X2_284 ( .A(u0__abc_76628_new_n1551_), .B(u0__abc_76628_new_n1552_), .Y(u0__abc_76628_new_n1553_));
OR2X2 OR2X2_2840 ( .A(u3__abc_74070_new_n412_), .B(u3__abc_74070_new_n413_), .Y(u3__abc_74070_new_n414_));
OR2X2 OR2X2_2841 ( .A(u3__abc_74070_new_n418_), .B(u3__abc_74070_new_n416_), .Y(u3__abc_74070_new_n419_));
OR2X2 OR2X2_2842 ( .A(u3__abc_74070_new_n420_), .B(u3__abc_74070_new_n421_), .Y(u3__0mc_dp_o_3_0__3_));
OR2X2 OR2X2_2843 ( .A(u3_byte2_0_), .B(pack_le2), .Y(u3__abc_74070_new_n423_));
OR2X2 OR2X2_2844 ( .A(u3__abc_74070_new_n424_), .B(mc_data_ir_0_), .Y(u3__abc_74070_new_n425_));
OR2X2 OR2X2_2845 ( .A(pack_le2), .B(u3_byte2_1_), .Y(u3__abc_74070_new_n427_));
OR2X2 OR2X2_2846 ( .A(u3__abc_74070_new_n424_), .B(mc_data_ir_1_), .Y(u3__abc_74070_new_n428_));
OR2X2 OR2X2_2847 ( .A(pack_le2), .B(u3_byte2_2_), .Y(u3__abc_74070_new_n430_));
OR2X2 OR2X2_2848 ( .A(u3__abc_74070_new_n424_), .B(mc_data_ir_2_), .Y(u3__abc_74070_new_n431_));
OR2X2 OR2X2_2849 ( .A(pack_le2), .B(u3_byte2_3_), .Y(u3__abc_74070_new_n433_));
OR2X2 OR2X2_285 ( .A(u0__abc_76628_new_n1555_), .B(spec_req_cs_0_bF_buf5_), .Y(u0__abc_76628_new_n1556_));
OR2X2 OR2X2_2850 ( .A(u3__abc_74070_new_n424_), .B(mc_data_ir_3_), .Y(u3__abc_74070_new_n434_));
OR2X2 OR2X2_2851 ( .A(pack_le2), .B(u3_byte2_4_), .Y(u3__abc_74070_new_n436_));
OR2X2 OR2X2_2852 ( .A(u3__abc_74070_new_n424_), .B(mc_data_ir_4_), .Y(u3__abc_74070_new_n437_));
OR2X2 OR2X2_2853 ( .A(pack_le2), .B(u3_byte2_5_), .Y(u3__abc_74070_new_n439_));
OR2X2 OR2X2_2854 ( .A(u3__abc_74070_new_n424_), .B(mc_data_ir_5_), .Y(u3__abc_74070_new_n440_));
OR2X2 OR2X2_2855 ( .A(pack_le2), .B(u3_byte2_6_), .Y(u3__abc_74070_new_n442_));
OR2X2 OR2X2_2856 ( .A(u3__abc_74070_new_n424_), .B(mc_data_ir_6_), .Y(u3__abc_74070_new_n443_));
OR2X2 OR2X2_2857 ( .A(pack_le2), .B(u3_byte2_7_), .Y(u3__abc_74070_new_n445_));
OR2X2 OR2X2_2858 ( .A(u3__abc_74070_new_n424_), .B(mc_data_ir_7_), .Y(u3__abc_74070_new_n446_));
OR2X2 OR2X2_2859 ( .A(u3__abc_74070_new_n454_), .B(mc_data_ir_8_), .Y(u3__abc_74070_new_n455_));
OR2X2 OR2X2_286 ( .A(u0__abc_76628_new_n1554_), .B(u0__abc_76628_new_n1556_), .Y(u0__abc_76628_new_n1557_));
OR2X2 OR2X2_2860 ( .A(u3__abc_74070_new_n453_), .B(u3_byte1_0_), .Y(u3__abc_74070_new_n456_));
OR2X2 OR2X2_2861 ( .A(u3__abc_74070_new_n457_), .B(u3__abc_74070_new_n451_), .Y(u3__abc_74070_new_n458_));
OR2X2 OR2X2_2862 ( .A(u3__abc_74070_new_n459_), .B(mc_data_ir_0_), .Y(u3__abc_74070_new_n460_));
OR2X2 OR2X2_2863 ( .A(u3__abc_74070_new_n454_), .B(mc_data_ir_9_), .Y(u3__abc_74070_new_n462_));
OR2X2 OR2X2_2864 ( .A(u3__abc_74070_new_n453_), .B(u3_byte1_1_), .Y(u3__abc_74070_new_n463_));
OR2X2 OR2X2_2865 ( .A(u3__abc_74070_new_n464_), .B(u3__abc_74070_new_n451_), .Y(u3__abc_74070_new_n465_));
OR2X2 OR2X2_2866 ( .A(u3__abc_74070_new_n459_), .B(mc_data_ir_1_), .Y(u3__abc_74070_new_n466_));
OR2X2 OR2X2_2867 ( .A(u3__abc_74070_new_n454_), .B(mc_data_ir_10_), .Y(u3__abc_74070_new_n468_));
OR2X2 OR2X2_2868 ( .A(u3__abc_74070_new_n453_), .B(u3_byte1_2_), .Y(u3__abc_74070_new_n469_));
OR2X2 OR2X2_2869 ( .A(u3__abc_74070_new_n470_), .B(u3__abc_74070_new_n451_), .Y(u3__abc_74070_new_n471_));
OR2X2 OR2X2_287 ( .A(u0__abc_76628_new_n1197__bF_buf2), .B(u0_tms0_15_), .Y(u0__abc_76628_new_n1558_));
OR2X2 OR2X2_2870 ( .A(u3__abc_74070_new_n459_), .B(mc_data_ir_2_), .Y(u3__abc_74070_new_n472_));
OR2X2 OR2X2_2871 ( .A(u3__abc_74070_new_n454_), .B(mc_data_ir_11_), .Y(u3__abc_74070_new_n474_));
OR2X2 OR2X2_2872 ( .A(u3__abc_74070_new_n453_), .B(u3_byte1_3_), .Y(u3__abc_74070_new_n475_));
OR2X2 OR2X2_2873 ( .A(u3__abc_74070_new_n476_), .B(u3__abc_74070_new_n451_), .Y(u3__abc_74070_new_n477_));
OR2X2 OR2X2_2874 ( .A(u3__abc_74070_new_n459_), .B(mc_data_ir_3_), .Y(u3__abc_74070_new_n478_));
OR2X2 OR2X2_2875 ( .A(u3__abc_74070_new_n454_), .B(mc_data_ir_12_), .Y(u3__abc_74070_new_n480_));
OR2X2 OR2X2_2876 ( .A(u3__abc_74070_new_n453_), .B(u3_byte1_4_), .Y(u3__abc_74070_new_n481_));
OR2X2 OR2X2_2877 ( .A(u3__abc_74070_new_n482_), .B(u3__abc_74070_new_n451_), .Y(u3__abc_74070_new_n483_));
OR2X2 OR2X2_2878 ( .A(u3__abc_74070_new_n459_), .B(mc_data_ir_4_), .Y(u3__abc_74070_new_n484_));
OR2X2 OR2X2_2879 ( .A(u3__abc_74070_new_n454_), .B(mc_data_ir_13_), .Y(u3__abc_74070_new_n486_));
OR2X2 OR2X2_288 ( .A(u0__abc_76628_new_n1560_), .B(u0__abc_76628_new_n1538_), .Y(u0__0sp_tms_31_0__15_));
OR2X2 OR2X2_2880 ( .A(u3__abc_74070_new_n453_), .B(u3_byte1_5_), .Y(u3__abc_74070_new_n487_));
OR2X2 OR2X2_2881 ( .A(u3__abc_74070_new_n488_), .B(u3__abc_74070_new_n451_), .Y(u3__abc_74070_new_n489_));
OR2X2 OR2X2_2882 ( .A(u3__abc_74070_new_n459_), .B(mc_data_ir_5_), .Y(u3__abc_74070_new_n490_));
OR2X2 OR2X2_2883 ( .A(u3__abc_74070_new_n454_), .B(mc_data_ir_14_), .Y(u3__abc_74070_new_n492_));
OR2X2 OR2X2_2884 ( .A(u3__abc_74070_new_n453_), .B(u3_byte1_6_), .Y(u3__abc_74070_new_n493_));
OR2X2 OR2X2_2885 ( .A(u3__abc_74070_new_n494_), .B(u3__abc_74070_new_n451_), .Y(u3__abc_74070_new_n495_));
OR2X2 OR2X2_2886 ( .A(u3__abc_74070_new_n459_), .B(mc_data_ir_6_), .Y(u3__abc_74070_new_n496_));
OR2X2 OR2X2_2887 ( .A(u3__abc_74070_new_n454_), .B(mc_data_ir_15_), .Y(u3__abc_74070_new_n498_));
OR2X2 OR2X2_2888 ( .A(u3__abc_74070_new_n453_), .B(u3_byte1_7_), .Y(u3__abc_74070_new_n499_));
OR2X2 OR2X2_2889 ( .A(u3__abc_74070_new_n500_), .B(u3__abc_74070_new_n451_), .Y(u3__abc_74070_new_n501_));
OR2X2 OR2X2_289 ( .A(u0__abc_76628_new_n1177__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n1564_));
OR2X2 OR2X2_2890 ( .A(u3__abc_74070_new_n459_), .B(mc_data_ir_7_), .Y(u3__abc_74070_new_n502_));
OR2X2 OR2X2_2891 ( .A(pack_le0), .B(u3_byte0_0_), .Y(u3__abc_74070_new_n504_));
OR2X2 OR2X2_2892 ( .A(u3__abc_74070_new_n505_), .B(mc_data_ir_0_), .Y(u3__abc_74070_new_n506_));
OR2X2 OR2X2_2893 ( .A(pack_le0), .B(u3_byte0_1_), .Y(u3__abc_74070_new_n508_));
OR2X2 OR2X2_2894 ( .A(u3__abc_74070_new_n505_), .B(mc_data_ir_1_), .Y(u3__abc_74070_new_n509_));
OR2X2 OR2X2_2895 ( .A(pack_le0), .B(u3_byte0_2_), .Y(u3__abc_74070_new_n511_));
OR2X2 OR2X2_2896 ( .A(u3__abc_74070_new_n505_), .B(mc_data_ir_2_), .Y(u3__abc_74070_new_n512_));
OR2X2 OR2X2_2897 ( .A(pack_le0), .B(u3_byte0_3_), .Y(u3__abc_74070_new_n514_));
OR2X2 OR2X2_2898 ( .A(u3__abc_74070_new_n505_), .B(mc_data_ir_3_), .Y(u3__abc_74070_new_n515_));
OR2X2 OR2X2_2899 ( .A(pack_le0), .B(u3_byte0_4_), .Y(u3__abc_74070_new_n517_));
OR2X2 OR2X2_29 ( .A(_abc_85006_new_n280_), .B(_abc_85006_new_n237_), .Y(_abc_85006_new_n281_));
OR2X2 OR2X2_290 ( .A(spec_req_cs_6_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1565_));
OR2X2 OR2X2_2900 ( .A(u3__abc_74070_new_n505_), .B(mc_data_ir_4_), .Y(u3__abc_74070_new_n518_));
OR2X2 OR2X2_2901 ( .A(pack_le0), .B(u3_byte0_5_), .Y(u3__abc_74070_new_n520_));
OR2X2 OR2X2_2902 ( .A(u3__abc_74070_new_n505_), .B(mc_data_ir_5_), .Y(u3__abc_74070_new_n521_));
OR2X2 OR2X2_2903 ( .A(pack_le0), .B(u3_byte0_6_), .Y(u3__abc_74070_new_n523_));
OR2X2 OR2X2_2904 ( .A(u3__abc_74070_new_n505_), .B(mc_data_ir_6_), .Y(u3__abc_74070_new_n524_));
OR2X2 OR2X2_2905 ( .A(pack_le0), .B(u3_byte0_7_), .Y(u3__abc_74070_new_n526_));
OR2X2 OR2X2_2906 ( .A(u3__abc_74070_new_n505_), .B(mc_data_ir_7_), .Y(u3__abc_74070_new_n527_));
OR2X2 OR2X2_2907 ( .A(u3__abc_74070_new_n279__bF_buf1), .B(\wb_data_i[0] ), .Y(u3__abc_74070_new_n529_));
OR2X2 OR2X2_2908 ( .A(u3__abc_74070_new_n277__bF_buf0), .B(mc_data_od_0_), .Y(u3__abc_74070_new_n530_));
OR2X2 OR2X2_2909 ( .A(u3__abc_74070_new_n279__bF_buf0), .B(\wb_data_i[1] ), .Y(u3__abc_74070_new_n532_));
OR2X2 OR2X2_291 ( .A(u0__abc_76628_new_n1567_), .B(u0__abc_76628_new_n1563_), .Y(u0__abc_76628_new_n1568_));
OR2X2 OR2X2_2910 ( .A(u3__abc_74070_new_n277__bF_buf5), .B(mc_data_od_1_), .Y(u3__abc_74070_new_n533_));
OR2X2 OR2X2_2911 ( .A(u3__abc_74070_new_n279__bF_buf5), .B(\wb_data_i[2] ), .Y(u3__abc_74070_new_n535_));
OR2X2 OR2X2_2912 ( .A(u3__abc_74070_new_n277__bF_buf4), .B(mc_data_od_2_), .Y(u3__abc_74070_new_n536_));
OR2X2 OR2X2_2913 ( .A(u3__abc_74070_new_n279__bF_buf4), .B(\wb_data_i[3] ), .Y(u3__abc_74070_new_n538_));
OR2X2 OR2X2_2914 ( .A(u3__abc_74070_new_n277__bF_buf3), .B(mc_data_od_3_), .Y(u3__abc_74070_new_n539_));
OR2X2 OR2X2_2915 ( .A(u3__abc_74070_new_n279__bF_buf3), .B(\wb_data_i[4] ), .Y(u3__abc_74070_new_n541_));
OR2X2 OR2X2_2916 ( .A(u3__abc_74070_new_n277__bF_buf2), .B(mc_data_od_4_), .Y(u3__abc_74070_new_n542_));
OR2X2 OR2X2_2917 ( .A(u3__abc_74070_new_n279__bF_buf2), .B(\wb_data_i[5] ), .Y(u3__abc_74070_new_n544_));
OR2X2 OR2X2_2918 ( .A(u3__abc_74070_new_n277__bF_buf1), .B(mc_data_od_5_), .Y(u3__abc_74070_new_n545_));
OR2X2 OR2X2_2919 ( .A(u3__abc_74070_new_n279__bF_buf1), .B(\wb_data_i[6] ), .Y(u3__abc_74070_new_n547_));
OR2X2 OR2X2_292 ( .A(u0__abc_76628_new_n1569_), .B(u0__abc_76628_new_n1570_), .Y(u0__abc_76628_new_n1571_));
OR2X2 OR2X2_2920 ( .A(u3__abc_74070_new_n277__bF_buf0), .B(mc_data_od_6_), .Y(u3__abc_74070_new_n548_));
OR2X2 OR2X2_2921 ( .A(u3__abc_74070_new_n279__bF_buf0), .B(\wb_data_i[7] ), .Y(u3__abc_74070_new_n550_));
OR2X2 OR2X2_2922 ( .A(u3__abc_74070_new_n277__bF_buf5), .B(mc_data_od_7_), .Y(u3__abc_74070_new_n551_));
OR2X2 OR2X2_2923 ( .A(u3__abc_74070_new_n279__bF_buf5), .B(\wb_data_i[8] ), .Y(u3__abc_74070_new_n553_));
OR2X2 OR2X2_2924 ( .A(u3__abc_74070_new_n277__bF_buf4), .B(mc_data_od_8_), .Y(u3__abc_74070_new_n554_));
OR2X2 OR2X2_2925 ( .A(u3__abc_74070_new_n279__bF_buf4), .B(\wb_data_i[9] ), .Y(u3__abc_74070_new_n556_));
OR2X2 OR2X2_2926 ( .A(u3__abc_74070_new_n277__bF_buf3), .B(mc_data_od_9_), .Y(u3__abc_74070_new_n557_));
OR2X2 OR2X2_2927 ( .A(u3__abc_74070_new_n279__bF_buf3), .B(\wb_data_i[10] ), .Y(u3__abc_74070_new_n559_));
OR2X2 OR2X2_2928 ( .A(u3__abc_74070_new_n277__bF_buf2), .B(mc_data_od_10_), .Y(u3__abc_74070_new_n560_));
OR2X2 OR2X2_2929 ( .A(u3__abc_74070_new_n279__bF_buf2), .B(\wb_data_i[11] ), .Y(u3__abc_74070_new_n562_));
OR2X2 OR2X2_293 ( .A(u0__abc_76628_new_n1572_), .B(u0__abc_76628_new_n1573_), .Y(u0__abc_76628_new_n1574_));
OR2X2 OR2X2_2930 ( .A(u3__abc_74070_new_n277__bF_buf1), .B(mc_data_od_11_), .Y(u3__abc_74070_new_n563_));
OR2X2 OR2X2_2931 ( .A(u3__abc_74070_new_n279__bF_buf1), .B(\wb_data_i[12] ), .Y(u3__abc_74070_new_n565_));
OR2X2 OR2X2_2932 ( .A(u3__abc_74070_new_n277__bF_buf0), .B(mc_data_od_12_), .Y(u3__abc_74070_new_n566_));
OR2X2 OR2X2_2933 ( .A(u3__abc_74070_new_n279__bF_buf0), .B(\wb_data_i[13] ), .Y(u3__abc_74070_new_n568_));
OR2X2 OR2X2_2934 ( .A(u3__abc_74070_new_n277__bF_buf5), .B(mc_data_od_13_), .Y(u3__abc_74070_new_n569_));
OR2X2 OR2X2_2935 ( .A(u3__abc_74070_new_n279__bF_buf5), .B(\wb_data_i[14] ), .Y(u3__abc_74070_new_n571_));
OR2X2 OR2X2_2936 ( .A(u3__abc_74070_new_n277__bF_buf4), .B(mc_data_od_14_), .Y(u3__abc_74070_new_n572_));
OR2X2 OR2X2_2937 ( .A(u3__abc_74070_new_n279__bF_buf4), .B(\wb_data_i[15] ), .Y(u3__abc_74070_new_n574_));
OR2X2 OR2X2_2938 ( .A(u3__abc_74070_new_n277__bF_buf3), .B(mc_data_od_15_), .Y(u3__abc_74070_new_n575_));
OR2X2 OR2X2_2939 ( .A(u3__abc_74070_new_n279__bF_buf3), .B(\wb_data_i[16] ), .Y(u3__abc_74070_new_n577_));
OR2X2 OR2X2_294 ( .A(u0__abc_76628_new_n1575_), .B(u0__abc_76628_new_n1576_), .Y(u0__abc_76628_new_n1577_));
OR2X2 OR2X2_2940 ( .A(u3__abc_74070_new_n277__bF_buf2), .B(mc_data_od_16_), .Y(u3__abc_74070_new_n578_));
OR2X2 OR2X2_2941 ( .A(u3__abc_74070_new_n279__bF_buf2), .B(\wb_data_i[17] ), .Y(u3__abc_74070_new_n580_));
OR2X2 OR2X2_2942 ( .A(u3__abc_74070_new_n277__bF_buf1), .B(mc_data_od_17_), .Y(u3__abc_74070_new_n581_));
OR2X2 OR2X2_2943 ( .A(u3__abc_74070_new_n279__bF_buf1), .B(\wb_data_i[18] ), .Y(u3__abc_74070_new_n583_));
OR2X2 OR2X2_2944 ( .A(u3__abc_74070_new_n277__bF_buf0), .B(mc_data_od_18_), .Y(u3__abc_74070_new_n584_));
OR2X2 OR2X2_2945 ( .A(u3__abc_74070_new_n279__bF_buf0), .B(\wb_data_i[19] ), .Y(u3__abc_74070_new_n586_));
OR2X2 OR2X2_2946 ( .A(u3__abc_74070_new_n277__bF_buf5), .B(mc_data_od_19_), .Y(u3__abc_74070_new_n587_));
OR2X2 OR2X2_2947 ( .A(u3__abc_74070_new_n279__bF_buf5), .B(\wb_data_i[20] ), .Y(u3__abc_74070_new_n589_));
OR2X2 OR2X2_2948 ( .A(u3__abc_74070_new_n277__bF_buf4), .B(mc_data_od_20_), .Y(u3__abc_74070_new_n590_));
OR2X2 OR2X2_2949 ( .A(u3__abc_74070_new_n279__bF_buf4), .B(\wb_data_i[21] ), .Y(u3__abc_74070_new_n592_));
OR2X2 OR2X2_295 ( .A(u0__abc_76628_new_n1579_), .B(spec_req_cs_0_bF_buf4_), .Y(u0__abc_76628_new_n1580_));
OR2X2 OR2X2_2950 ( .A(u3__abc_74070_new_n277__bF_buf3), .B(mc_data_od_21_), .Y(u3__abc_74070_new_n593_));
OR2X2 OR2X2_2951 ( .A(u3__abc_74070_new_n279__bF_buf3), .B(\wb_data_i[22] ), .Y(u3__abc_74070_new_n595_));
OR2X2 OR2X2_2952 ( .A(u3__abc_74070_new_n277__bF_buf2), .B(mc_data_od_22_), .Y(u3__abc_74070_new_n596_));
OR2X2 OR2X2_2953 ( .A(u3__abc_74070_new_n279__bF_buf2), .B(\wb_data_i[23] ), .Y(u3__abc_74070_new_n598_));
OR2X2 OR2X2_2954 ( .A(u3__abc_74070_new_n277__bF_buf1), .B(mc_data_od_23_), .Y(u3__abc_74070_new_n599_));
OR2X2 OR2X2_2955 ( .A(u3__abc_74070_new_n279__bF_buf1), .B(\wb_data_i[24] ), .Y(u3__abc_74070_new_n601_));
OR2X2 OR2X2_2956 ( .A(u3__abc_74070_new_n277__bF_buf0), .B(mc_data_od_24_), .Y(u3__abc_74070_new_n602_));
OR2X2 OR2X2_2957 ( .A(u3__abc_74070_new_n279__bF_buf0), .B(\wb_data_i[25] ), .Y(u3__abc_74070_new_n604_));
OR2X2 OR2X2_2958 ( .A(u3__abc_74070_new_n277__bF_buf5), .B(mc_data_od_25_), .Y(u3__abc_74070_new_n605_));
OR2X2 OR2X2_2959 ( .A(u3__abc_74070_new_n279__bF_buf5), .B(\wb_data_i[26] ), .Y(u3__abc_74070_new_n607_));
OR2X2 OR2X2_296 ( .A(u0__abc_76628_new_n1578_), .B(u0__abc_76628_new_n1580_), .Y(u0__abc_76628_new_n1581_));
OR2X2 OR2X2_2960 ( .A(u3__abc_74070_new_n277__bF_buf4), .B(mc_data_od_26_), .Y(u3__abc_74070_new_n608_));
OR2X2 OR2X2_2961 ( .A(u3__abc_74070_new_n279__bF_buf4), .B(\wb_data_i[27] ), .Y(u3__abc_74070_new_n610_));
OR2X2 OR2X2_2962 ( .A(u3__abc_74070_new_n277__bF_buf3), .B(mc_data_od_27_), .Y(u3__abc_74070_new_n611_));
OR2X2 OR2X2_2963 ( .A(u3__abc_74070_new_n279__bF_buf3), .B(\wb_data_i[28] ), .Y(u3__abc_74070_new_n613_));
OR2X2 OR2X2_2964 ( .A(u3__abc_74070_new_n277__bF_buf2), .B(mc_data_od_28_), .Y(u3__abc_74070_new_n614_));
OR2X2 OR2X2_2965 ( .A(u3__abc_74070_new_n279__bF_buf2), .B(\wb_data_i[29] ), .Y(u3__abc_74070_new_n616_));
OR2X2 OR2X2_2966 ( .A(u3__abc_74070_new_n277__bF_buf1), .B(mc_data_od_29_), .Y(u3__abc_74070_new_n617_));
OR2X2 OR2X2_2967 ( .A(u3__abc_74070_new_n279__bF_buf1), .B(\wb_data_i[30] ), .Y(u3__abc_74070_new_n619_));
OR2X2 OR2X2_2968 ( .A(u3__abc_74070_new_n277__bF_buf0), .B(mc_data_od_30_), .Y(u3__abc_74070_new_n620_));
OR2X2 OR2X2_2969 ( .A(u3__abc_74070_new_n279__bF_buf0), .B(\wb_data_i[31] ), .Y(u3__abc_74070_new_n622_));
OR2X2 OR2X2_297 ( .A(u0__abc_76628_new_n1197__bF_buf1), .B(u0_tms0_16_), .Y(u0__abc_76628_new_n1582_));
OR2X2 OR2X2_2970 ( .A(u3__abc_74070_new_n277__bF_buf5), .B(mc_data_od_31_), .Y(u3__abc_74070_new_n623_));
OR2X2 OR2X2_2971 ( .A(csc_5_bF_buf1_), .B(u3_byte0_0_), .Y(u3__abc_74070_new_n626_));
OR2X2 OR2X2_2972 ( .A(u3__abc_74070_new_n449__bF_buf1), .B(mc_data_ir_0_), .Y(u3__abc_74070_new_n627_));
OR2X2 OR2X2_2973 ( .A(u3__abc_74070_new_n628_), .B(u3__abc_74070_new_n625__bF_buf4), .Y(u3__abc_74070_new_n629_));
OR2X2 OR2X2_2974 ( .A(u3__abc_74070_new_n275__bF_buf2), .B(u3_rd_fifo_out_0_), .Y(u3__abc_74070_new_n630_));
OR2X2 OR2X2_2975 ( .A(csc_5_bF_buf0_), .B(u3_byte0_1_), .Y(u3__abc_74070_new_n632_));
OR2X2 OR2X2_2976 ( .A(u3__abc_74070_new_n449__bF_buf0), .B(mc_data_ir_1_), .Y(u3__abc_74070_new_n633_));
OR2X2 OR2X2_2977 ( .A(u3__abc_74070_new_n634_), .B(u3__abc_74070_new_n625__bF_buf3), .Y(u3__abc_74070_new_n635_));
OR2X2 OR2X2_2978 ( .A(u3__abc_74070_new_n275__bF_buf1), .B(u3_rd_fifo_out_1_), .Y(u3__abc_74070_new_n636_));
OR2X2 OR2X2_2979 ( .A(csc_5_bF_buf4_), .B(u3_byte0_2_), .Y(u3__abc_74070_new_n638_));
OR2X2 OR2X2_298 ( .A(u0__abc_76628_new_n1584_), .B(u0__abc_76628_new_n1562_), .Y(u0__0sp_tms_31_0__16_));
OR2X2 OR2X2_2980 ( .A(u3__abc_74070_new_n449__bF_buf3), .B(mc_data_ir_2_), .Y(u3__abc_74070_new_n639_));
OR2X2 OR2X2_2981 ( .A(u3__abc_74070_new_n640_), .B(u3__abc_74070_new_n625__bF_buf2), .Y(u3__abc_74070_new_n641_));
OR2X2 OR2X2_2982 ( .A(u3__abc_74070_new_n275__bF_buf0), .B(u3_rd_fifo_out_2_), .Y(u3__abc_74070_new_n642_));
OR2X2 OR2X2_2983 ( .A(csc_5_bF_buf3_), .B(u3_byte0_3_), .Y(u3__abc_74070_new_n644_));
OR2X2 OR2X2_2984 ( .A(u3__abc_74070_new_n449__bF_buf2), .B(mc_data_ir_3_), .Y(u3__abc_74070_new_n645_));
OR2X2 OR2X2_2985 ( .A(u3__abc_74070_new_n646_), .B(u3__abc_74070_new_n625__bF_buf1), .Y(u3__abc_74070_new_n647_));
OR2X2 OR2X2_2986 ( .A(u3__abc_74070_new_n275__bF_buf4), .B(u3_rd_fifo_out_3_), .Y(u3__abc_74070_new_n648_));
OR2X2 OR2X2_2987 ( .A(csc_5_bF_buf2_), .B(u3_byte0_4_), .Y(u3__abc_74070_new_n650_));
OR2X2 OR2X2_2988 ( .A(u3__abc_74070_new_n449__bF_buf1), .B(mc_data_ir_4_), .Y(u3__abc_74070_new_n651_));
OR2X2 OR2X2_2989 ( .A(u3__abc_74070_new_n652_), .B(u3__abc_74070_new_n625__bF_buf0), .Y(u3__abc_74070_new_n653_));
OR2X2 OR2X2_299 ( .A(u0__abc_76628_new_n1177__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n1588_));
OR2X2 OR2X2_2990 ( .A(u3__abc_74070_new_n275__bF_buf3), .B(u3_rd_fifo_out_4_), .Y(u3__abc_74070_new_n654_));
OR2X2 OR2X2_2991 ( .A(csc_5_bF_buf1_), .B(u3_byte0_5_), .Y(u3__abc_74070_new_n656_));
OR2X2 OR2X2_2992 ( .A(u3__abc_74070_new_n449__bF_buf0), .B(mc_data_ir_5_), .Y(u3__abc_74070_new_n657_));
OR2X2 OR2X2_2993 ( .A(u3__abc_74070_new_n658_), .B(u3__abc_74070_new_n625__bF_buf4), .Y(u3__abc_74070_new_n659_));
OR2X2 OR2X2_2994 ( .A(u3__abc_74070_new_n275__bF_buf2), .B(u3_rd_fifo_out_5_), .Y(u3__abc_74070_new_n660_));
OR2X2 OR2X2_2995 ( .A(csc_5_bF_buf0_), .B(u3_byte0_6_), .Y(u3__abc_74070_new_n662_));
OR2X2 OR2X2_2996 ( .A(u3__abc_74070_new_n449__bF_buf3), .B(mc_data_ir_6_), .Y(u3__abc_74070_new_n663_));
OR2X2 OR2X2_2997 ( .A(u3__abc_74070_new_n664_), .B(u3__abc_74070_new_n625__bF_buf3), .Y(u3__abc_74070_new_n665_));
OR2X2 OR2X2_2998 ( .A(u3__abc_74070_new_n275__bF_buf1), .B(u3_rd_fifo_out_6_), .Y(u3__abc_74070_new_n666_));
OR2X2 OR2X2_2999 ( .A(csc_5_bF_buf4_), .B(u3_byte0_7_), .Y(u3__abc_74070_new_n668_));
OR2X2 OR2X2_3 ( .A(_abc_85006_new_n240__bF_buf5), .B(spec_req_cs_0_bF_buf5_), .Y(_abc_85006_new_n241_));
OR2X2 OR2X2_30 ( .A(_abc_85006_new_n245_), .B(cs_need_rfr_6_), .Y(_abc_85006_new_n282_));
OR2X2 OR2X2_300 ( .A(spec_req_cs_6_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1589_));
OR2X2 OR2X2_3000 ( .A(u3__abc_74070_new_n449__bF_buf2), .B(mc_data_ir_7_), .Y(u3__abc_74070_new_n669_));
OR2X2 OR2X2_3001 ( .A(u3__abc_74070_new_n670_), .B(u3__abc_74070_new_n625__bF_buf2), .Y(u3__abc_74070_new_n671_));
OR2X2 OR2X2_3002 ( .A(u3__abc_74070_new_n275__bF_buf0), .B(u3_rd_fifo_out_7_), .Y(u3__abc_74070_new_n672_));
OR2X2 OR2X2_3003 ( .A(csc_5_bF_buf3_), .B(u3_byte1_0_), .Y(u3__abc_74070_new_n674_));
OR2X2 OR2X2_3004 ( .A(u3__abc_74070_new_n449__bF_buf1), .B(mc_data_ir_8_), .Y(u3__abc_74070_new_n675_));
OR2X2 OR2X2_3005 ( .A(u3__abc_74070_new_n676_), .B(u3__abc_74070_new_n625__bF_buf1), .Y(u3__abc_74070_new_n677_));
OR2X2 OR2X2_3006 ( .A(u3__abc_74070_new_n275__bF_buf4), .B(u3_rd_fifo_out_8_), .Y(u3__abc_74070_new_n678_));
OR2X2 OR2X2_3007 ( .A(csc_5_bF_buf2_), .B(u3_byte1_1_), .Y(u3__abc_74070_new_n680_));
OR2X2 OR2X2_3008 ( .A(u3__abc_74070_new_n449__bF_buf0), .B(mc_data_ir_9_), .Y(u3__abc_74070_new_n681_));
OR2X2 OR2X2_3009 ( .A(u3__abc_74070_new_n682_), .B(u3__abc_74070_new_n625__bF_buf0), .Y(u3__abc_74070_new_n683_));
OR2X2 OR2X2_301 ( .A(u0__abc_76628_new_n1591_), .B(u0__abc_76628_new_n1587_), .Y(u0__abc_76628_new_n1592_));
OR2X2 OR2X2_3010 ( .A(u3__abc_74070_new_n275__bF_buf3), .B(u3_rd_fifo_out_9_), .Y(u3__abc_74070_new_n684_));
OR2X2 OR2X2_3011 ( .A(csc_5_bF_buf1_), .B(u3_byte1_2_), .Y(u3__abc_74070_new_n686_));
OR2X2 OR2X2_3012 ( .A(u3__abc_74070_new_n449__bF_buf3), .B(mc_data_ir_10_), .Y(u3__abc_74070_new_n687_));
OR2X2 OR2X2_3013 ( .A(u3__abc_74070_new_n688_), .B(u3__abc_74070_new_n625__bF_buf4), .Y(u3__abc_74070_new_n689_));
OR2X2 OR2X2_3014 ( .A(u3__abc_74070_new_n275__bF_buf2), .B(u3_rd_fifo_out_10_), .Y(u3__abc_74070_new_n690_));
OR2X2 OR2X2_3015 ( .A(csc_5_bF_buf0_), .B(u3_byte1_3_), .Y(u3__abc_74070_new_n692_));
OR2X2 OR2X2_3016 ( .A(u3__abc_74070_new_n449__bF_buf2), .B(mc_data_ir_11_), .Y(u3__abc_74070_new_n693_));
OR2X2 OR2X2_3017 ( .A(u3__abc_74070_new_n694_), .B(u3__abc_74070_new_n625__bF_buf3), .Y(u3__abc_74070_new_n695_));
OR2X2 OR2X2_3018 ( .A(u3__abc_74070_new_n275__bF_buf1), .B(u3_rd_fifo_out_11_), .Y(u3__abc_74070_new_n696_));
OR2X2 OR2X2_3019 ( .A(csc_5_bF_buf4_), .B(u3_byte1_4_), .Y(u3__abc_74070_new_n698_));
OR2X2 OR2X2_302 ( .A(u0__abc_76628_new_n1593_), .B(u0__abc_76628_new_n1594_), .Y(u0__abc_76628_new_n1595_));
OR2X2 OR2X2_3020 ( .A(u3__abc_74070_new_n449__bF_buf1), .B(mc_data_ir_12_), .Y(u3__abc_74070_new_n699_));
OR2X2 OR2X2_3021 ( .A(u3__abc_74070_new_n700_), .B(u3__abc_74070_new_n625__bF_buf2), .Y(u3__abc_74070_new_n701_));
OR2X2 OR2X2_3022 ( .A(u3__abc_74070_new_n275__bF_buf0), .B(u3_rd_fifo_out_12_), .Y(u3__abc_74070_new_n702_));
OR2X2 OR2X2_3023 ( .A(csc_5_bF_buf3_), .B(u3_byte1_5_), .Y(u3__abc_74070_new_n704_));
OR2X2 OR2X2_3024 ( .A(u3__abc_74070_new_n449__bF_buf0), .B(mc_data_ir_13_), .Y(u3__abc_74070_new_n705_));
OR2X2 OR2X2_3025 ( .A(u3__abc_74070_new_n706_), .B(u3__abc_74070_new_n625__bF_buf1), .Y(u3__abc_74070_new_n707_));
OR2X2 OR2X2_3026 ( .A(u3__abc_74070_new_n275__bF_buf4), .B(u3_rd_fifo_out_13_), .Y(u3__abc_74070_new_n708_));
OR2X2 OR2X2_3027 ( .A(csc_5_bF_buf2_), .B(u3_byte1_6_), .Y(u3__abc_74070_new_n710_));
OR2X2 OR2X2_3028 ( .A(u3__abc_74070_new_n449__bF_buf3), .B(mc_data_ir_14_), .Y(u3__abc_74070_new_n711_));
OR2X2 OR2X2_3029 ( .A(u3__abc_74070_new_n712_), .B(u3__abc_74070_new_n625__bF_buf0), .Y(u3__abc_74070_new_n713_));
OR2X2 OR2X2_303 ( .A(u0__abc_76628_new_n1596_), .B(u0__abc_76628_new_n1597_), .Y(u0__abc_76628_new_n1598_));
OR2X2 OR2X2_3030 ( .A(u3__abc_74070_new_n275__bF_buf3), .B(u3_rd_fifo_out_14_), .Y(u3__abc_74070_new_n714_));
OR2X2 OR2X2_3031 ( .A(csc_5_bF_buf1_), .B(u3_byte1_7_), .Y(u3__abc_74070_new_n716_));
OR2X2 OR2X2_3032 ( .A(u3__abc_74070_new_n449__bF_buf2), .B(mc_data_ir_15_), .Y(u3__abc_74070_new_n717_));
OR2X2 OR2X2_3033 ( .A(u3__abc_74070_new_n718_), .B(u3__abc_74070_new_n625__bF_buf4), .Y(u3__abc_74070_new_n719_));
OR2X2 OR2X2_3034 ( .A(u3__abc_74070_new_n275__bF_buf2), .B(u3_rd_fifo_out_15_), .Y(u3__abc_74070_new_n720_));
OR2X2 OR2X2_3035 ( .A(u3__abc_74070_new_n722_), .B(u3__abc_74070_new_n723_), .Y(u3__abc_74070_new_n724_));
OR2X2 OR2X2_3036 ( .A(u3__abc_74070_new_n725_), .B(u3__abc_74070_new_n625__bF_buf3), .Y(u3__abc_74070_new_n726_));
OR2X2 OR2X2_3037 ( .A(u3__abc_74070_new_n726_), .B(u3__abc_74070_new_n724_), .Y(u3__abc_74070_new_n727_));
OR2X2 OR2X2_3038 ( .A(u3__abc_74070_new_n275__bF_buf1), .B(u3_rd_fifo_out_16_), .Y(u3__abc_74070_new_n728_));
OR2X2 OR2X2_3039 ( .A(u3__abc_74070_new_n730_), .B(u3__abc_74070_new_n731_), .Y(u3__abc_74070_new_n732_));
OR2X2 OR2X2_304 ( .A(u0__abc_76628_new_n1599_), .B(u0__abc_76628_new_n1600_), .Y(u0__abc_76628_new_n1601_));
OR2X2 OR2X2_3040 ( .A(u3__abc_74070_new_n733_), .B(u3__abc_74070_new_n625__bF_buf2), .Y(u3__abc_74070_new_n734_));
OR2X2 OR2X2_3041 ( .A(u3__abc_74070_new_n734_), .B(u3__abc_74070_new_n732_), .Y(u3__abc_74070_new_n735_));
OR2X2 OR2X2_3042 ( .A(u3__abc_74070_new_n275__bF_buf0), .B(u3_rd_fifo_out_17_), .Y(u3__abc_74070_new_n736_));
OR2X2 OR2X2_3043 ( .A(u3__abc_74070_new_n738_), .B(u3__abc_74070_new_n739_), .Y(u3__abc_74070_new_n740_));
OR2X2 OR2X2_3044 ( .A(u3__abc_74070_new_n741_), .B(u3__abc_74070_new_n625__bF_buf1), .Y(u3__abc_74070_new_n742_));
OR2X2 OR2X2_3045 ( .A(u3__abc_74070_new_n742_), .B(u3__abc_74070_new_n740_), .Y(u3__abc_74070_new_n743_));
OR2X2 OR2X2_3046 ( .A(u3__abc_74070_new_n275__bF_buf4), .B(u3_rd_fifo_out_18_), .Y(u3__abc_74070_new_n744_));
OR2X2 OR2X2_3047 ( .A(u3__abc_74070_new_n746_), .B(u3__abc_74070_new_n747_), .Y(u3__abc_74070_new_n748_));
OR2X2 OR2X2_3048 ( .A(u3__abc_74070_new_n749_), .B(u3__abc_74070_new_n625__bF_buf0), .Y(u3__abc_74070_new_n750_));
OR2X2 OR2X2_3049 ( .A(u3__abc_74070_new_n750_), .B(u3__abc_74070_new_n748_), .Y(u3__abc_74070_new_n751_));
OR2X2 OR2X2_305 ( .A(u0__abc_76628_new_n1603_), .B(spec_req_cs_0_bF_buf3_), .Y(u0__abc_76628_new_n1604_));
OR2X2 OR2X2_3050 ( .A(u3__abc_74070_new_n275__bF_buf3), .B(u3_rd_fifo_out_19_), .Y(u3__abc_74070_new_n752_));
OR2X2 OR2X2_3051 ( .A(u3__abc_74070_new_n754_), .B(u3__abc_74070_new_n755_), .Y(u3__abc_74070_new_n756_));
OR2X2 OR2X2_3052 ( .A(u3__abc_74070_new_n757_), .B(u3__abc_74070_new_n625__bF_buf4), .Y(u3__abc_74070_new_n758_));
OR2X2 OR2X2_3053 ( .A(u3__abc_74070_new_n758_), .B(u3__abc_74070_new_n756_), .Y(u3__abc_74070_new_n759_));
OR2X2 OR2X2_3054 ( .A(u3__abc_74070_new_n275__bF_buf2), .B(u3_rd_fifo_out_20_), .Y(u3__abc_74070_new_n760_));
OR2X2 OR2X2_3055 ( .A(u3__abc_74070_new_n762_), .B(u3__abc_74070_new_n763_), .Y(u3__abc_74070_new_n764_));
OR2X2 OR2X2_3056 ( .A(u3__abc_74070_new_n765_), .B(u3__abc_74070_new_n625__bF_buf3), .Y(u3__abc_74070_new_n766_));
OR2X2 OR2X2_3057 ( .A(u3__abc_74070_new_n766_), .B(u3__abc_74070_new_n764_), .Y(u3__abc_74070_new_n767_));
OR2X2 OR2X2_3058 ( .A(u3__abc_74070_new_n275__bF_buf1), .B(u3_rd_fifo_out_21_), .Y(u3__abc_74070_new_n768_));
OR2X2 OR2X2_3059 ( .A(u3__abc_74070_new_n770_), .B(u3__abc_74070_new_n771_), .Y(u3__abc_74070_new_n772_));
OR2X2 OR2X2_306 ( .A(u0__abc_76628_new_n1602_), .B(u0__abc_76628_new_n1604_), .Y(u0__abc_76628_new_n1605_));
OR2X2 OR2X2_3060 ( .A(u3__abc_74070_new_n773_), .B(u3__abc_74070_new_n625__bF_buf2), .Y(u3__abc_74070_new_n774_));
OR2X2 OR2X2_3061 ( .A(u3__abc_74070_new_n774_), .B(u3__abc_74070_new_n772_), .Y(u3__abc_74070_new_n775_));
OR2X2 OR2X2_3062 ( .A(u3__abc_74070_new_n275__bF_buf0), .B(u3_rd_fifo_out_22_), .Y(u3__abc_74070_new_n776_));
OR2X2 OR2X2_3063 ( .A(u3__abc_74070_new_n778_), .B(u3__abc_74070_new_n779_), .Y(u3__abc_74070_new_n780_));
OR2X2 OR2X2_3064 ( .A(u3__abc_74070_new_n781_), .B(u3__abc_74070_new_n625__bF_buf1), .Y(u3__abc_74070_new_n782_));
OR2X2 OR2X2_3065 ( .A(u3__abc_74070_new_n782_), .B(u3__abc_74070_new_n780_), .Y(u3__abc_74070_new_n783_));
OR2X2 OR2X2_3066 ( .A(u3__abc_74070_new_n275__bF_buf4), .B(u3_rd_fifo_out_23_), .Y(u3__abc_74070_new_n784_));
OR2X2 OR2X2_3067 ( .A(u3__abc_74070_new_n786_), .B(u3__abc_74070_new_n787_), .Y(u3__abc_74070_new_n788_));
OR2X2 OR2X2_3068 ( .A(u3__abc_74070_new_n789_), .B(u3__abc_74070_new_n625__bF_buf0), .Y(u3__abc_74070_new_n790_));
OR2X2 OR2X2_3069 ( .A(u3__abc_74070_new_n790_), .B(u3__abc_74070_new_n788_), .Y(u3__abc_74070_new_n791_));
OR2X2 OR2X2_307 ( .A(u0__abc_76628_new_n1197__bF_buf0), .B(u0_tms0_17_), .Y(u0__abc_76628_new_n1606_));
OR2X2 OR2X2_3070 ( .A(u3__abc_74070_new_n275__bF_buf3), .B(u3_rd_fifo_out_24_), .Y(u3__abc_74070_new_n792_));
OR2X2 OR2X2_3071 ( .A(u3__abc_74070_new_n794_), .B(u3__abc_74070_new_n795_), .Y(u3__abc_74070_new_n796_));
OR2X2 OR2X2_3072 ( .A(u3__abc_74070_new_n797_), .B(u3__abc_74070_new_n625__bF_buf4), .Y(u3__abc_74070_new_n798_));
OR2X2 OR2X2_3073 ( .A(u3__abc_74070_new_n798_), .B(u3__abc_74070_new_n796_), .Y(u3__abc_74070_new_n799_));
OR2X2 OR2X2_3074 ( .A(u3__abc_74070_new_n275__bF_buf2), .B(u3_rd_fifo_out_25_), .Y(u3__abc_74070_new_n800_));
OR2X2 OR2X2_3075 ( .A(u3__abc_74070_new_n802_), .B(u3__abc_74070_new_n803_), .Y(u3__abc_74070_new_n804_));
OR2X2 OR2X2_3076 ( .A(u3__abc_74070_new_n805_), .B(u3__abc_74070_new_n625__bF_buf3), .Y(u3__abc_74070_new_n806_));
OR2X2 OR2X2_3077 ( .A(u3__abc_74070_new_n806_), .B(u3__abc_74070_new_n804_), .Y(u3__abc_74070_new_n807_));
OR2X2 OR2X2_3078 ( .A(u3__abc_74070_new_n275__bF_buf1), .B(u3_rd_fifo_out_26_), .Y(u3__abc_74070_new_n808_));
OR2X2 OR2X2_3079 ( .A(u3__abc_74070_new_n810_), .B(u3__abc_74070_new_n811_), .Y(u3__abc_74070_new_n812_));
OR2X2 OR2X2_308 ( .A(u0__abc_76628_new_n1608_), .B(u0__abc_76628_new_n1586_), .Y(u0__0sp_tms_31_0__17_));
OR2X2 OR2X2_3080 ( .A(u3__abc_74070_new_n813_), .B(u3__abc_74070_new_n625__bF_buf2), .Y(u3__abc_74070_new_n814_));
OR2X2 OR2X2_3081 ( .A(u3__abc_74070_new_n814_), .B(u3__abc_74070_new_n812_), .Y(u3__abc_74070_new_n815_));
OR2X2 OR2X2_3082 ( .A(u3__abc_74070_new_n275__bF_buf0), .B(u3_rd_fifo_out_27_), .Y(u3__abc_74070_new_n816_));
OR2X2 OR2X2_3083 ( .A(u3__abc_74070_new_n818_), .B(u3__abc_74070_new_n819_), .Y(u3__abc_74070_new_n820_));
OR2X2 OR2X2_3084 ( .A(u3__abc_74070_new_n821_), .B(u3__abc_74070_new_n625__bF_buf1), .Y(u3__abc_74070_new_n822_));
OR2X2 OR2X2_3085 ( .A(u3__abc_74070_new_n822_), .B(u3__abc_74070_new_n820_), .Y(u3__abc_74070_new_n823_));
OR2X2 OR2X2_3086 ( .A(u3__abc_74070_new_n275__bF_buf4), .B(u3_rd_fifo_out_28_), .Y(u3__abc_74070_new_n824_));
OR2X2 OR2X2_3087 ( .A(u3__abc_74070_new_n826_), .B(u3__abc_74070_new_n827_), .Y(u3__abc_74070_new_n828_));
OR2X2 OR2X2_3088 ( .A(u3__abc_74070_new_n829_), .B(u3__abc_74070_new_n625__bF_buf0), .Y(u3__abc_74070_new_n830_));
OR2X2 OR2X2_3089 ( .A(u3__abc_74070_new_n830_), .B(u3__abc_74070_new_n828_), .Y(u3__abc_74070_new_n831_));
OR2X2 OR2X2_309 ( .A(u0__abc_76628_new_n1177__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n1612_));
OR2X2 OR2X2_3090 ( .A(u3__abc_74070_new_n275__bF_buf3), .B(u3_rd_fifo_out_29_), .Y(u3__abc_74070_new_n832_));
OR2X2 OR2X2_3091 ( .A(u3__abc_74070_new_n834_), .B(u3__abc_74070_new_n835_), .Y(u3__abc_74070_new_n836_));
OR2X2 OR2X2_3092 ( .A(u3__abc_74070_new_n837_), .B(u3__abc_74070_new_n625__bF_buf4), .Y(u3__abc_74070_new_n838_));
OR2X2 OR2X2_3093 ( .A(u3__abc_74070_new_n838_), .B(u3__abc_74070_new_n836_), .Y(u3__abc_74070_new_n839_));
OR2X2 OR2X2_3094 ( .A(u3__abc_74070_new_n275__bF_buf2), .B(u3_rd_fifo_out_30_), .Y(u3__abc_74070_new_n840_));
OR2X2 OR2X2_3095 ( .A(u3__abc_74070_new_n842_), .B(u3__abc_74070_new_n843_), .Y(u3__abc_74070_new_n844_));
OR2X2 OR2X2_3096 ( .A(u3__abc_74070_new_n845_), .B(u3__abc_74070_new_n625__bF_buf3), .Y(u3__abc_74070_new_n846_));
OR2X2 OR2X2_3097 ( .A(u3__abc_74070_new_n846_), .B(u3__abc_74070_new_n844_), .Y(u3__abc_74070_new_n847_));
OR2X2 OR2X2_3098 ( .A(u3__abc_74070_new_n275__bF_buf1), .B(u3_rd_fifo_out_31_), .Y(u3__abc_74070_new_n848_));
OR2X2 OR2X2_3099 ( .A(u3__abc_74070_new_n851_), .B(u3__abc_74070_new_n850_), .Y(u3_rd_fifo_clr));
OR2X2 OR2X2_31 ( .A(_abc_85006_new_n240__bF_buf4), .B(spec_req_cs_7_), .Y(_abc_85006_new_n284_));
OR2X2 OR2X2_310 ( .A(spec_req_cs_6_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1613_));
OR2X2 OR2X2_3100 ( .A(u3_rd_fifo_out_22_), .B(u3_rd_fifo_out_23_), .Y(u3__abc_74070_new_n854_));
OR2X2 OR2X2_3101 ( .A(u3__abc_74070_new_n858_), .B(u3_rd_fifo_out_17_), .Y(u3__abc_74070_new_n859_));
OR2X2 OR2X2_3102 ( .A(u3__abc_74070_new_n860_), .B(u3_rd_fifo_out_16_), .Y(u3__abc_74070_new_n861_));
OR2X2 OR2X2_3103 ( .A(u3__abc_74070_new_n865_), .B(u3__abc_74070_new_n866_), .Y(u3__abc_74070_new_n867_));
OR2X2 OR2X2_3104 ( .A(u3__abc_74070_new_n868_), .B(u3__abc_74070_new_n863_), .Y(u3__abc_74070_new_n869_));
OR2X2 OR2X2_3105 ( .A(u3__abc_74070_new_n867_), .B(u3__abc_74070_new_n864_), .Y(u3__abc_74070_new_n872_));
OR2X2 OR2X2_3106 ( .A(u3__abc_74070_new_n862_), .B(u3_rd_fifo_out_34_), .Y(u3__abc_74070_new_n873_));
OR2X2 OR2X2_3107 ( .A(u3__abc_74070_new_n870_), .B(u3__abc_74070_new_n875_), .Y(u3__abc_74070_new_n876_));
OR2X2 OR2X2_3108 ( .A(u3_rd_fifo_out_20_), .B(u3_rd_fifo_out_21_), .Y(u3__abc_74070_new_n878_));
OR2X2 OR2X2_3109 ( .A(u3__abc_74070_new_n882_), .B(u3_rd_fifo_out_18_), .Y(u3__abc_74070_new_n885_));
OR2X2 OR2X2_311 ( .A(u0__abc_76628_new_n1615_), .B(u0__abc_76628_new_n1611_), .Y(u0__abc_76628_new_n1616_));
OR2X2 OR2X2_3110 ( .A(u3__abc_74070_new_n886_), .B(u3__abc_74070_new_n881_), .Y(u3__abc_74070_new_n887_));
OR2X2 OR2X2_3111 ( .A(u3__abc_74070_new_n889_), .B(u3__abc_74070_new_n888_), .Y(u3__abc_74070_new_n890_));
OR2X2 OR2X2_3112 ( .A(u3__abc_74070_new_n877_), .B(u3__abc_74070_new_n892_), .Y(u3__abc_74070_new_n893_));
OR2X2 OR2X2_3113 ( .A(u3__abc_74070_new_n876_), .B(u3__abc_74070_new_n891_), .Y(u3__abc_74070_new_n894_));
OR2X2 OR2X2_3114 ( .A(u3_rd_fifo_out_30_), .B(u3_rd_fifo_out_31_), .Y(u3__abc_74070_new_n897_));
OR2X2 OR2X2_3115 ( .A(u3__abc_74070_new_n903_), .B(u3__abc_74070_new_n904_), .Y(u3__abc_74070_new_n905_));
OR2X2 OR2X2_3116 ( .A(u3_rd_fifo_out_24_), .B(u3_rd_fifo_out_25_), .Y(u3__abc_74070_new_n908_));
OR2X2 OR2X2_3117 ( .A(u3__abc_74070_new_n906_), .B(u3__abc_74070_new_n911_), .Y(u3__abc_74070_new_n912_));
OR2X2 OR2X2_3118 ( .A(u3__abc_74070_new_n910_), .B(u3__abc_74070_new_n907_), .Y(u3__abc_74070_new_n915_));
OR2X2 OR2X2_3119 ( .A(u3__abc_74070_new_n905_), .B(u3_rd_fifo_out_35_), .Y(u3__abc_74070_new_n916_));
OR2X2 OR2X2_312 ( .A(u0__abc_76628_new_n1617_), .B(u0__abc_76628_new_n1618_), .Y(u0__abc_76628_new_n1619_));
OR2X2 OR2X2_3120 ( .A(u3__abc_74070_new_n913_), .B(u3__abc_74070_new_n918_), .Y(u3__abc_74070_new_n919_));
OR2X2 OR2X2_3121 ( .A(u3_rd_fifo_out_28_), .B(u3_rd_fifo_out_29_), .Y(u3__abc_74070_new_n921_));
OR2X2 OR2X2_3122 ( .A(u3__abc_74070_new_n925_), .B(u3_rd_fifo_out_26_), .Y(u3__abc_74070_new_n928_));
OR2X2 OR2X2_3123 ( .A(u3__abc_74070_new_n929_), .B(u3__abc_74070_new_n924_), .Y(u3__abc_74070_new_n930_));
OR2X2 OR2X2_3124 ( .A(u3__abc_74070_new_n932_), .B(u3__abc_74070_new_n931_), .Y(u3__abc_74070_new_n933_));
OR2X2 OR2X2_3125 ( .A(u3__abc_74070_new_n920_), .B(u3__abc_74070_new_n935_), .Y(u3__abc_74070_new_n936_));
OR2X2 OR2X2_3126 ( .A(u3__abc_74070_new_n919_), .B(u3__abc_74070_new_n934_), .Y(u3__abc_74070_new_n937_));
OR2X2 OR2X2_3127 ( .A(u3__abc_74070_new_n896_), .B(u3__abc_74070_new_n939_), .Y(u3__abc_74070_new_n940_));
OR2X2 OR2X2_3128 ( .A(u3_rd_fifo_out_14_), .B(u3_rd_fifo_out_15_), .Y(u3__abc_74070_new_n941_));
OR2X2 OR2X2_3129 ( .A(u3_rd_fifo_out_8_), .B(u3_rd_fifo_out_9_), .Y(u3__abc_74070_new_n947_));
OR2X2 OR2X2_313 ( .A(u0__abc_76628_new_n1620_), .B(u0__abc_76628_new_n1621_), .Y(u0__abc_76628_new_n1622_));
OR2X2 OR2X2_3130 ( .A(u3__abc_74070_new_n950_), .B(u3__abc_74070_new_n946_), .Y(u3__abc_74070_new_n951_));
OR2X2 OR2X2_3131 ( .A(u3__abc_74070_new_n954_), .B(u3__abc_74070_new_n948_), .Y(u3__abc_74070_new_n955_));
OR2X2 OR2X2_3132 ( .A(u3__abc_74070_new_n955_), .B(u3_rd_fifo_out_33_), .Y(u3__abc_74070_new_n956_));
OR2X2 OR2X2_3133 ( .A(u3__abc_74070_new_n957_), .B(u3__abc_74070_new_n945_), .Y(u3__abc_74070_new_n958_));
OR2X2 OR2X2_3134 ( .A(u3__abc_74070_new_n959_), .B(u3__abc_74070_new_n960_), .Y(u3__abc_74070_new_n961_));
OR2X2 OR2X2_3135 ( .A(u3__abc_74070_new_n961_), .B(u3__abc_74070_new_n944_), .Y(u3__abc_74070_new_n962_));
OR2X2 OR2X2_3136 ( .A(u3_rd_fifo_out_12_), .B(u3_rd_fifo_out_13_), .Y(u3__abc_74070_new_n965_));
OR2X2 OR2X2_3137 ( .A(u3__abc_74070_new_n970_), .B(u3_rd_fifo_out_10_), .Y(u3__abc_74070_new_n973_));
OR2X2 OR2X2_3138 ( .A(u3__abc_74070_new_n976_), .B(u3__abc_74070_new_n977_), .Y(u3__abc_74070_new_n978_));
OR2X2 OR2X2_3139 ( .A(u3__abc_74070_new_n964_), .B(u3__abc_74070_new_n979_), .Y(u3__abc_74070_new_n980_));
OR2X2 OR2X2_314 ( .A(u0__abc_76628_new_n1623_), .B(u0__abc_76628_new_n1624_), .Y(u0__abc_76628_new_n1625_));
OR2X2 OR2X2_3140 ( .A(u3__abc_74070_new_n963_), .B(u3__abc_74070_new_n978_), .Y(u3__abc_74070_new_n981_));
OR2X2 OR2X2_3141 ( .A(u3_rd_fifo_out_6_), .B(u3_rd_fifo_out_7_), .Y(u3__abc_74070_new_n984_));
OR2X2 OR2X2_3142 ( .A(u3_rd_fifo_out_0_), .B(u3_rd_fifo_out_1_), .Y(u3__abc_74070_new_n990_));
OR2X2 OR2X2_3143 ( .A(u3__abc_74070_new_n993_), .B(u3__abc_74070_new_n989_), .Y(u3__abc_74070_new_n994_));
OR2X2 OR2X2_3144 ( .A(u3__abc_74070_new_n995_), .B(u3_rd_fifo_out_1_), .Y(u3__abc_74070_new_n996_));
OR2X2 OR2X2_3145 ( .A(u3__abc_74070_new_n997_), .B(u3_rd_fifo_out_0_), .Y(u3__abc_74070_new_n998_));
OR2X2 OR2X2_3146 ( .A(u3__abc_74070_new_n999_), .B(u3_rd_fifo_out_32_), .Y(u3__abc_74070_new_n1000_));
OR2X2 OR2X2_3147 ( .A(u3__abc_74070_new_n1001_), .B(u3__abc_74070_new_n988_), .Y(u3__abc_74070_new_n1002_));
OR2X2 OR2X2_3148 ( .A(u3__abc_74070_new_n1003_), .B(u3__abc_74070_new_n1004_), .Y(u3__abc_74070_new_n1005_));
OR2X2 OR2X2_3149 ( .A(u3__abc_74070_new_n1005_), .B(u3__abc_74070_new_n987_), .Y(u3__abc_74070_new_n1006_));
OR2X2 OR2X2_315 ( .A(u0__abc_76628_new_n1627_), .B(spec_req_cs_0_bF_buf2_), .Y(u0__abc_76628_new_n1628_));
OR2X2 OR2X2_3150 ( .A(u3_rd_fifo_out_4_), .B(u3_rd_fifo_out_5_), .Y(u3__abc_74070_new_n1009_));
OR2X2 OR2X2_3151 ( .A(u3__abc_74070_new_n1014_), .B(u3_rd_fifo_out_2_), .Y(u3__abc_74070_new_n1017_));
OR2X2 OR2X2_3152 ( .A(u3__abc_74070_new_n1020_), .B(u3__abc_74070_new_n1021_), .Y(u3__abc_74070_new_n1022_));
OR2X2 OR2X2_3153 ( .A(u3__abc_74070_new_n1008_), .B(u3__abc_74070_new_n1023_), .Y(u3__abc_74070_new_n1024_));
OR2X2 OR2X2_3154 ( .A(u3__abc_74070_new_n1007_), .B(u3__abc_74070_new_n1022_), .Y(u3__abc_74070_new_n1025_));
OR2X2 OR2X2_3155 ( .A(u3__abc_74070_new_n983_), .B(u3__abc_74070_new_n1027_), .Y(u3__abc_74070_new_n1028_));
OR2X2 OR2X2_3156 ( .A(u3__abc_74070_new_n940_), .B(u3__abc_74070_new_n1028_), .Y(u3__abc_74070_new_n1029_));
OR2X2 OR2X2_3157 ( .A(u3_u0__abc_75526_new_n382__bF_buf7), .B(u3_u0_r1_0_), .Y(u3_u0__abc_75526_new_n383_));
OR2X2 OR2X2_3158 ( .A(u3_u0__abc_75526_new_n382__bF_buf5), .B(u3_u0_r1_1_), .Y(u3_u0__abc_75526_new_n388_));
OR2X2 OR2X2_3159 ( .A(u3_u0__abc_75526_new_n382__bF_buf3), .B(u3_u0_r1_2_), .Y(u3_u0__abc_75526_new_n393_));
OR2X2 OR2X2_316 ( .A(u0__abc_76628_new_n1626_), .B(u0__abc_76628_new_n1628_), .Y(u0__abc_76628_new_n1629_));
OR2X2 OR2X2_3160 ( .A(u3_u0__abc_75526_new_n382__bF_buf1), .B(u3_u0_r1_3_), .Y(u3_u0__abc_75526_new_n398_));
OR2X2 OR2X2_3161 ( .A(u3_u0__abc_75526_new_n382__bF_buf7), .B(u3_u0_r1_4_), .Y(u3_u0__abc_75526_new_n403_));
OR2X2 OR2X2_3162 ( .A(u3_u0__abc_75526_new_n382__bF_buf5), .B(u3_u0_r1_5_), .Y(u3_u0__abc_75526_new_n408_));
OR2X2 OR2X2_3163 ( .A(u3_u0__abc_75526_new_n382__bF_buf3), .B(u3_u0_r1_6_), .Y(u3_u0__abc_75526_new_n413_));
OR2X2 OR2X2_3164 ( .A(u3_u0__abc_75526_new_n382__bF_buf1), .B(u3_u0_r1_7_), .Y(u3_u0__abc_75526_new_n418_));
OR2X2 OR2X2_3165 ( .A(u3_u0__abc_75526_new_n382__bF_buf7), .B(u3_u0_r1_8_), .Y(u3_u0__abc_75526_new_n423_));
OR2X2 OR2X2_3166 ( .A(u3_u0__abc_75526_new_n382__bF_buf5), .B(u3_u0_r1_9_), .Y(u3_u0__abc_75526_new_n428_));
OR2X2 OR2X2_3167 ( .A(u3_u0__abc_75526_new_n382__bF_buf3), .B(u3_u0_r1_10_), .Y(u3_u0__abc_75526_new_n433_));
OR2X2 OR2X2_3168 ( .A(u3_u0__abc_75526_new_n382__bF_buf1), .B(u3_u0_r1_11_), .Y(u3_u0__abc_75526_new_n438_));
OR2X2 OR2X2_3169 ( .A(u3_u0__abc_75526_new_n382__bF_buf7), .B(u3_u0_r1_12_), .Y(u3_u0__abc_75526_new_n443_));
OR2X2 OR2X2_317 ( .A(u0__abc_76628_new_n1197__bF_buf5), .B(u0_tms0_18_), .Y(u0__abc_76628_new_n1630_));
OR2X2 OR2X2_3170 ( .A(u3_u0__abc_75526_new_n382__bF_buf5), .B(u3_u0_r1_13_), .Y(u3_u0__abc_75526_new_n448_));
OR2X2 OR2X2_3171 ( .A(u3_u0__abc_75526_new_n382__bF_buf3), .B(u3_u0_r1_14_), .Y(u3_u0__abc_75526_new_n453_));
OR2X2 OR2X2_3172 ( .A(u3_u0__abc_75526_new_n382__bF_buf1), .B(u3_u0_r1_15_), .Y(u3_u0__abc_75526_new_n458_));
OR2X2 OR2X2_3173 ( .A(u3_u0__abc_75526_new_n382__bF_buf7), .B(u3_u0_r1_16_), .Y(u3_u0__abc_75526_new_n463_));
OR2X2 OR2X2_3174 ( .A(u3_u0__abc_75526_new_n382__bF_buf5), .B(u3_u0_r1_17_), .Y(u3_u0__abc_75526_new_n468_));
OR2X2 OR2X2_3175 ( .A(u3_u0__abc_75526_new_n382__bF_buf3), .B(u3_u0_r1_18_), .Y(u3_u0__abc_75526_new_n473_));
OR2X2 OR2X2_3176 ( .A(u3_u0__abc_75526_new_n382__bF_buf1), .B(u3_u0_r1_19_), .Y(u3_u0__abc_75526_new_n478_));
OR2X2 OR2X2_3177 ( .A(u3_u0__abc_75526_new_n382__bF_buf7), .B(u3_u0_r1_20_), .Y(u3_u0__abc_75526_new_n483_));
OR2X2 OR2X2_3178 ( .A(u3_u0__abc_75526_new_n382__bF_buf5), .B(u3_u0_r1_21_), .Y(u3_u0__abc_75526_new_n488_));
OR2X2 OR2X2_3179 ( .A(u3_u0__abc_75526_new_n382__bF_buf3), .B(u3_u0_r1_22_), .Y(u3_u0__abc_75526_new_n493_));
OR2X2 OR2X2_318 ( .A(u0__abc_76628_new_n1632_), .B(u0__abc_76628_new_n1610_), .Y(u0__0sp_tms_31_0__18_));
OR2X2 OR2X2_3180 ( .A(u3_u0__abc_75526_new_n382__bF_buf1), .B(u3_u0_r1_23_), .Y(u3_u0__abc_75526_new_n498_));
OR2X2 OR2X2_3181 ( .A(u3_u0__abc_75526_new_n382__bF_buf7), .B(u3_u0_r1_24_), .Y(u3_u0__abc_75526_new_n503_));
OR2X2 OR2X2_3182 ( .A(u3_u0__abc_75526_new_n382__bF_buf5), .B(u3_u0_r1_25_), .Y(u3_u0__abc_75526_new_n508_));
OR2X2 OR2X2_3183 ( .A(u3_u0__abc_75526_new_n382__bF_buf3), .B(u3_u0_r1_26_), .Y(u3_u0__abc_75526_new_n513_));
OR2X2 OR2X2_3184 ( .A(u3_u0__abc_75526_new_n382__bF_buf1), .B(u3_u0_r1_27_), .Y(u3_u0__abc_75526_new_n518_));
OR2X2 OR2X2_3185 ( .A(u3_u0__abc_75526_new_n382__bF_buf7), .B(u3_u0_r1_28_), .Y(u3_u0__abc_75526_new_n523_));
OR2X2 OR2X2_3186 ( .A(u3_u0__abc_75526_new_n382__bF_buf5), .B(u3_u0_r1_29_), .Y(u3_u0__abc_75526_new_n528_));
OR2X2 OR2X2_3187 ( .A(u3_u0__abc_75526_new_n382__bF_buf3), .B(u3_u0_r1_30_), .Y(u3_u0__abc_75526_new_n533_));
OR2X2 OR2X2_3188 ( .A(u3_u0__abc_75526_new_n382__bF_buf1), .B(u3_u0_r1_31_), .Y(u3_u0__abc_75526_new_n538_));
OR2X2 OR2X2_3189 ( .A(u3_u0__abc_75526_new_n382__bF_buf7), .B(u3_u0_r1_32_), .Y(u3_u0__abc_75526_new_n543_));
OR2X2 OR2X2_319 ( .A(u0__abc_76628_new_n1177__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n1636_));
OR2X2 OR2X2_3190 ( .A(u3_u0__abc_75526_new_n382__bF_buf5), .B(u3_u0_r1_33_), .Y(u3_u0__abc_75526_new_n548_));
OR2X2 OR2X2_3191 ( .A(u3_u0__abc_75526_new_n382__bF_buf3), .B(u3_u0_r1_34_), .Y(u3_u0__abc_75526_new_n553_));
OR2X2 OR2X2_3192 ( .A(u3_u0__abc_75526_new_n382__bF_buf1), .B(u3_u0_r1_35_), .Y(u3_u0__abc_75526_new_n558_));
OR2X2 OR2X2_3193 ( .A(u3_u0__abc_75526_new_n563__bF_buf7), .B(u3_u0_r3_0_), .Y(u3_u0__abc_75526_new_n564_));
OR2X2 OR2X2_3194 ( .A(u3_u0__abc_75526_new_n563__bF_buf5), .B(u3_u0_r3_1_), .Y(u3_u0__abc_75526_new_n568_));
OR2X2 OR2X2_3195 ( .A(u3_u0__abc_75526_new_n563__bF_buf3), .B(u3_u0_r3_2_), .Y(u3_u0__abc_75526_new_n572_));
OR2X2 OR2X2_3196 ( .A(u3_u0__abc_75526_new_n563__bF_buf1), .B(u3_u0_r3_3_), .Y(u3_u0__abc_75526_new_n576_));
OR2X2 OR2X2_3197 ( .A(u3_u0__abc_75526_new_n563__bF_buf7), .B(u3_u0_r3_4_), .Y(u3_u0__abc_75526_new_n580_));
OR2X2 OR2X2_3198 ( .A(u3_u0__abc_75526_new_n563__bF_buf5), .B(u3_u0_r3_5_), .Y(u3_u0__abc_75526_new_n584_));
OR2X2 OR2X2_3199 ( .A(u3_u0__abc_75526_new_n563__bF_buf3), .B(u3_u0_r3_6_), .Y(u3_u0__abc_75526_new_n588_));
OR2X2 OR2X2_32 ( .A(lmr_sel_bF_buf6), .B(cs_7_), .Y(_abc_85006_new_n285_));
OR2X2 OR2X2_320 ( .A(spec_req_cs_6_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1637_));
OR2X2 OR2X2_3200 ( .A(u3_u0__abc_75526_new_n563__bF_buf1), .B(u3_u0_r3_7_), .Y(u3_u0__abc_75526_new_n592_));
OR2X2 OR2X2_3201 ( .A(u3_u0__abc_75526_new_n563__bF_buf7), .B(u3_u0_r3_8_), .Y(u3_u0__abc_75526_new_n596_));
OR2X2 OR2X2_3202 ( .A(u3_u0__abc_75526_new_n563__bF_buf5), .B(u3_u0_r3_9_), .Y(u3_u0__abc_75526_new_n600_));
OR2X2 OR2X2_3203 ( .A(u3_u0__abc_75526_new_n563__bF_buf3), .B(u3_u0_r3_10_), .Y(u3_u0__abc_75526_new_n604_));
OR2X2 OR2X2_3204 ( .A(u3_u0__abc_75526_new_n563__bF_buf1), .B(u3_u0_r3_11_), .Y(u3_u0__abc_75526_new_n608_));
OR2X2 OR2X2_3205 ( .A(u3_u0__abc_75526_new_n563__bF_buf7), .B(u3_u0_r3_12_), .Y(u3_u0__abc_75526_new_n612_));
OR2X2 OR2X2_3206 ( .A(u3_u0__abc_75526_new_n563__bF_buf5), .B(u3_u0_r3_13_), .Y(u3_u0__abc_75526_new_n616_));
OR2X2 OR2X2_3207 ( .A(u3_u0__abc_75526_new_n563__bF_buf3), .B(u3_u0_r3_14_), .Y(u3_u0__abc_75526_new_n620_));
OR2X2 OR2X2_3208 ( .A(u3_u0__abc_75526_new_n563__bF_buf1), .B(u3_u0_r3_15_), .Y(u3_u0__abc_75526_new_n624_));
OR2X2 OR2X2_3209 ( .A(u3_u0__abc_75526_new_n563__bF_buf7), .B(u3_u0_r3_16_), .Y(u3_u0__abc_75526_new_n628_));
OR2X2 OR2X2_321 ( .A(u0__abc_76628_new_n1639_), .B(u0__abc_76628_new_n1635_), .Y(u0__abc_76628_new_n1640_));
OR2X2 OR2X2_3210 ( .A(u3_u0__abc_75526_new_n563__bF_buf5), .B(u3_u0_r3_17_), .Y(u3_u0__abc_75526_new_n632_));
OR2X2 OR2X2_3211 ( .A(u3_u0__abc_75526_new_n563__bF_buf3), .B(u3_u0_r3_18_), .Y(u3_u0__abc_75526_new_n636_));
OR2X2 OR2X2_3212 ( .A(u3_u0__abc_75526_new_n563__bF_buf1), .B(u3_u0_r3_19_), .Y(u3_u0__abc_75526_new_n640_));
OR2X2 OR2X2_3213 ( .A(u3_u0__abc_75526_new_n563__bF_buf7), .B(u3_u0_r3_20_), .Y(u3_u0__abc_75526_new_n644_));
OR2X2 OR2X2_3214 ( .A(u3_u0__abc_75526_new_n563__bF_buf5), .B(u3_u0_r3_21_), .Y(u3_u0__abc_75526_new_n648_));
OR2X2 OR2X2_3215 ( .A(u3_u0__abc_75526_new_n563__bF_buf3), .B(u3_u0_r3_22_), .Y(u3_u0__abc_75526_new_n652_));
OR2X2 OR2X2_3216 ( .A(u3_u0__abc_75526_new_n563__bF_buf1), .B(u3_u0_r3_23_), .Y(u3_u0__abc_75526_new_n656_));
OR2X2 OR2X2_3217 ( .A(u3_u0__abc_75526_new_n563__bF_buf7), .B(u3_u0_r3_24_), .Y(u3_u0__abc_75526_new_n660_));
OR2X2 OR2X2_3218 ( .A(u3_u0__abc_75526_new_n563__bF_buf5), .B(u3_u0_r3_25_), .Y(u3_u0__abc_75526_new_n664_));
OR2X2 OR2X2_3219 ( .A(u3_u0__abc_75526_new_n563__bF_buf3), .B(u3_u0_r3_26_), .Y(u3_u0__abc_75526_new_n668_));
OR2X2 OR2X2_322 ( .A(u0__abc_76628_new_n1641_), .B(u0__abc_76628_new_n1642_), .Y(u0__abc_76628_new_n1643_));
OR2X2 OR2X2_3220 ( .A(u3_u0__abc_75526_new_n563__bF_buf1), .B(u3_u0_r3_27_), .Y(u3_u0__abc_75526_new_n672_));
OR2X2 OR2X2_3221 ( .A(u3_u0__abc_75526_new_n563__bF_buf7), .B(u3_u0_r3_28_), .Y(u3_u0__abc_75526_new_n676_));
OR2X2 OR2X2_3222 ( .A(u3_u0__abc_75526_new_n563__bF_buf5), .B(u3_u0_r3_29_), .Y(u3_u0__abc_75526_new_n680_));
OR2X2 OR2X2_3223 ( .A(u3_u0__abc_75526_new_n563__bF_buf3), .B(u3_u0_r3_30_), .Y(u3_u0__abc_75526_new_n684_));
OR2X2 OR2X2_3224 ( .A(u3_u0__abc_75526_new_n563__bF_buf1), .B(u3_u0_r3_31_), .Y(u3_u0__abc_75526_new_n688_));
OR2X2 OR2X2_3225 ( .A(u3_u0__abc_75526_new_n563__bF_buf7), .B(u3_u0_r3_32_), .Y(u3_u0__abc_75526_new_n692_));
OR2X2 OR2X2_3226 ( .A(u3_u0__abc_75526_new_n563__bF_buf5), .B(u3_u0_r3_33_), .Y(u3_u0__abc_75526_new_n696_));
OR2X2 OR2X2_3227 ( .A(u3_u0__abc_75526_new_n563__bF_buf3), .B(u3_u0_r3_34_), .Y(u3_u0__abc_75526_new_n700_));
OR2X2 OR2X2_3228 ( .A(u3_u0__abc_75526_new_n563__bF_buf1), .B(u3_u0_r3_35_), .Y(u3_u0__abc_75526_new_n704_));
OR2X2 OR2X2_3229 ( .A(u3_u0__abc_75526_new_n708__bF_buf7), .B(u3_u0_r2_0_), .Y(u3_u0__abc_75526_new_n709_));
OR2X2 OR2X2_323 ( .A(u0__abc_76628_new_n1644_), .B(u0__abc_76628_new_n1645_), .Y(u0__abc_76628_new_n1646_));
OR2X2 OR2X2_3230 ( .A(u3_u0__abc_75526_new_n708__bF_buf5), .B(u3_u0_r2_1_), .Y(u3_u0__abc_75526_new_n713_));
OR2X2 OR2X2_3231 ( .A(u3_u0__abc_75526_new_n708__bF_buf3), .B(u3_u0_r2_2_), .Y(u3_u0__abc_75526_new_n717_));
OR2X2 OR2X2_3232 ( .A(u3_u0__abc_75526_new_n708__bF_buf1), .B(u3_u0_r2_3_), .Y(u3_u0__abc_75526_new_n721_));
OR2X2 OR2X2_3233 ( .A(u3_u0__abc_75526_new_n708__bF_buf7), .B(u3_u0_r2_4_), .Y(u3_u0__abc_75526_new_n725_));
OR2X2 OR2X2_3234 ( .A(u3_u0__abc_75526_new_n708__bF_buf5), .B(u3_u0_r2_5_), .Y(u3_u0__abc_75526_new_n729_));
OR2X2 OR2X2_3235 ( .A(u3_u0__abc_75526_new_n708__bF_buf3), .B(u3_u0_r2_6_), .Y(u3_u0__abc_75526_new_n733_));
OR2X2 OR2X2_3236 ( .A(u3_u0__abc_75526_new_n708__bF_buf1), .B(u3_u0_r2_7_), .Y(u3_u0__abc_75526_new_n737_));
OR2X2 OR2X2_3237 ( .A(u3_u0__abc_75526_new_n708__bF_buf7), .B(u3_u0_r2_8_), .Y(u3_u0__abc_75526_new_n741_));
OR2X2 OR2X2_3238 ( .A(u3_u0__abc_75526_new_n708__bF_buf5), .B(u3_u0_r2_9_), .Y(u3_u0__abc_75526_new_n745_));
OR2X2 OR2X2_3239 ( .A(u3_u0__abc_75526_new_n708__bF_buf3), .B(u3_u0_r2_10_), .Y(u3_u0__abc_75526_new_n749_));
OR2X2 OR2X2_324 ( .A(u0__abc_76628_new_n1647_), .B(u0__abc_76628_new_n1648_), .Y(u0__abc_76628_new_n1649_));
OR2X2 OR2X2_3240 ( .A(u3_u0__abc_75526_new_n708__bF_buf1), .B(u3_u0_r2_11_), .Y(u3_u0__abc_75526_new_n753_));
OR2X2 OR2X2_3241 ( .A(u3_u0__abc_75526_new_n708__bF_buf7), .B(u3_u0_r2_12_), .Y(u3_u0__abc_75526_new_n757_));
OR2X2 OR2X2_3242 ( .A(u3_u0__abc_75526_new_n708__bF_buf5), .B(u3_u0_r2_13_), .Y(u3_u0__abc_75526_new_n761_));
OR2X2 OR2X2_3243 ( .A(u3_u0__abc_75526_new_n708__bF_buf3), .B(u3_u0_r2_14_), .Y(u3_u0__abc_75526_new_n765_));
OR2X2 OR2X2_3244 ( .A(u3_u0__abc_75526_new_n708__bF_buf1), .B(u3_u0_r2_15_), .Y(u3_u0__abc_75526_new_n769_));
OR2X2 OR2X2_3245 ( .A(u3_u0__abc_75526_new_n708__bF_buf7), .B(u3_u0_r2_16_), .Y(u3_u0__abc_75526_new_n773_));
OR2X2 OR2X2_3246 ( .A(u3_u0__abc_75526_new_n708__bF_buf5), .B(u3_u0_r2_17_), .Y(u3_u0__abc_75526_new_n777_));
OR2X2 OR2X2_3247 ( .A(u3_u0__abc_75526_new_n708__bF_buf3), .B(u3_u0_r2_18_), .Y(u3_u0__abc_75526_new_n781_));
OR2X2 OR2X2_3248 ( .A(u3_u0__abc_75526_new_n708__bF_buf1), .B(u3_u0_r2_19_), .Y(u3_u0__abc_75526_new_n785_));
OR2X2 OR2X2_3249 ( .A(u3_u0__abc_75526_new_n708__bF_buf7), .B(u3_u0_r2_20_), .Y(u3_u0__abc_75526_new_n789_));
OR2X2 OR2X2_325 ( .A(u0__abc_76628_new_n1651_), .B(spec_req_cs_0_bF_buf1_), .Y(u0__abc_76628_new_n1652_));
OR2X2 OR2X2_3250 ( .A(u3_u0__abc_75526_new_n708__bF_buf5), .B(u3_u0_r2_21_), .Y(u3_u0__abc_75526_new_n793_));
OR2X2 OR2X2_3251 ( .A(u3_u0__abc_75526_new_n708__bF_buf3), .B(u3_u0_r2_22_), .Y(u3_u0__abc_75526_new_n797_));
OR2X2 OR2X2_3252 ( .A(u3_u0__abc_75526_new_n708__bF_buf1), .B(u3_u0_r2_23_), .Y(u3_u0__abc_75526_new_n801_));
OR2X2 OR2X2_3253 ( .A(u3_u0__abc_75526_new_n708__bF_buf7), .B(u3_u0_r2_24_), .Y(u3_u0__abc_75526_new_n805_));
OR2X2 OR2X2_3254 ( .A(u3_u0__abc_75526_new_n708__bF_buf5), .B(u3_u0_r2_25_), .Y(u3_u0__abc_75526_new_n809_));
OR2X2 OR2X2_3255 ( .A(u3_u0__abc_75526_new_n708__bF_buf3), .B(u3_u0_r2_26_), .Y(u3_u0__abc_75526_new_n813_));
OR2X2 OR2X2_3256 ( .A(u3_u0__abc_75526_new_n708__bF_buf1), .B(u3_u0_r2_27_), .Y(u3_u0__abc_75526_new_n817_));
OR2X2 OR2X2_3257 ( .A(u3_u0__abc_75526_new_n708__bF_buf7), .B(u3_u0_r2_28_), .Y(u3_u0__abc_75526_new_n821_));
OR2X2 OR2X2_3258 ( .A(u3_u0__abc_75526_new_n708__bF_buf5), .B(u3_u0_r2_29_), .Y(u3_u0__abc_75526_new_n825_));
OR2X2 OR2X2_3259 ( .A(u3_u0__abc_75526_new_n708__bF_buf3), .B(u3_u0_r2_30_), .Y(u3_u0__abc_75526_new_n829_));
OR2X2 OR2X2_326 ( .A(u0__abc_76628_new_n1650_), .B(u0__abc_76628_new_n1652_), .Y(u0__abc_76628_new_n1653_));
OR2X2 OR2X2_3260 ( .A(u3_u0__abc_75526_new_n708__bF_buf1), .B(u3_u0_r2_31_), .Y(u3_u0__abc_75526_new_n833_));
OR2X2 OR2X2_3261 ( .A(u3_u0__abc_75526_new_n708__bF_buf7), .B(u3_u0_r2_32_), .Y(u3_u0__abc_75526_new_n837_));
OR2X2 OR2X2_3262 ( .A(u3_u0__abc_75526_new_n708__bF_buf5), .B(u3_u0_r2_33_), .Y(u3_u0__abc_75526_new_n841_));
OR2X2 OR2X2_3263 ( .A(u3_u0__abc_75526_new_n708__bF_buf3), .B(u3_u0_r2_34_), .Y(u3_u0__abc_75526_new_n845_));
OR2X2 OR2X2_3264 ( .A(u3_u0__abc_75526_new_n708__bF_buf1), .B(u3_u0_r2_35_), .Y(u3_u0__abc_75526_new_n849_));
OR2X2 OR2X2_3265 ( .A(u3_u0__abc_75526_new_n855_), .B(u3_rd_fifo_clr), .Y(u3_u0__abc_75526_new_n856_));
OR2X2 OR2X2_3266 ( .A(u3_u0__abc_75526_new_n856_), .B(u3_u0__abc_75526_new_n854_), .Y(u3_u0__0rd_adr_3_0__0_));
OR2X2 OR2X2_3267 ( .A(u3_u0__abc_75526_new_n860_), .B(u3_u0__abc_75526_new_n859_), .Y(u3_u0__abc_75526_new_n861_));
OR2X2 OR2X2_3268 ( .A(u3_u0__abc_75526_new_n864_), .B(u3_u0__abc_75526_new_n863_), .Y(u3_u0__abc_75526_new_n865_));
OR2X2 OR2X2_3269 ( .A(u3_u0__abc_75526_new_n868_), .B(u3_u0__abc_75526_new_n867_), .Y(u3_u0__abc_75526_new_n869_));
OR2X2 OR2X2_327 ( .A(u0__abc_76628_new_n1197__bF_buf4), .B(u0_tms0_19_), .Y(u0__abc_76628_new_n1654_));
OR2X2 OR2X2_3270 ( .A(u3_u0__abc_75526_new_n563__bF_buf7), .B(u3_rd_fifo_clr), .Y(u3_u0__abc_75526_new_n873_));
OR2X2 OR2X2_3271 ( .A(u3_u0__abc_75526_new_n873_), .B(u3_u0__abc_75526_new_n872_), .Y(u3_u0__0wr_adr_3_0__0_));
OR2X2 OR2X2_3272 ( .A(u3_u0__abc_75526_new_n875_), .B(u3_u0__abc_75526_new_n876__bF_buf7), .Y(u3_u0__abc_75526_new_n877_));
OR2X2 OR2X2_3273 ( .A(u3_u0__abc_75526_new_n879_), .B(u3_u0__abc_75526_new_n382__bF_buf7), .Y(u3_u0__abc_75526_new_n880_));
OR2X2 OR2X2_3274 ( .A(u3_u0__abc_75526_new_n882_), .B(u3_u0__abc_75526_new_n708__bF_buf7), .Y(u3_u0__abc_75526_new_n883_));
OR2X2 OR2X2_3275 ( .A(u3_u0__abc_75526_new_n876__bF_buf6), .B(u3_u0_r0_0_), .Y(u3_u0__abc_75526_new_n885_));
OR2X2 OR2X2_3276 ( .A(u3_u0__abc_75526_new_n876__bF_buf4), .B(u3_u0_r0_1_), .Y(u3_u0__abc_75526_new_n889_));
OR2X2 OR2X2_3277 ( .A(u3_u0__abc_75526_new_n876__bF_buf2), .B(u3_u0_r0_2_), .Y(u3_u0__abc_75526_new_n893_));
OR2X2 OR2X2_3278 ( .A(u3_u0__abc_75526_new_n876__bF_buf0), .B(u3_u0_r0_3_), .Y(u3_u0__abc_75526_new_n897_));
OR2X2 OR2X2_3279 ( .A(u3_u0__abc_75526_new_n876__bF_buf6), .B(u3_u0_r0_4_), .Y(u3_u0__abc_75526_new_n901_));
OR2X2 OR2X2_328 ( .A(u0__abc_76628_new_n1656_), .B(u0__abc_76628_new_n1634_), .Y(u0__0sp_tms_31_0__19_));
OR2X2 OR2X2_3280 ( .A(u3_u0__abc_75526_new_n876__bF_buf4), .B(u3_u0_r0_5_), .Y(u3_u0__abc_75526_new_n905_));
OR2X2 OR2X2_3281 ( .A(u3_u0__abc_75526_new_n876__bF_buf2), .B(u3_u0_r0_6_), .Y(u3_u0__abc_75526_new_n909_));
OR2X2 OR2X2_3282 ( .A(u3_u0__abc_75526_new_n876__bF_buf0), .B(u3_u0_r0_7_), .Y(u3_u0__abc_75526_new_n913_));
OR2X2 OR2X2_3283 ( .A(u3_u0__abc_75526_new_n876__bF_buf6), .B(u3_u0_r0_8_), .Y(u3_u0__abc_75526_new_n917_));
OR2X2 OR2X2_3284 ( .A(u3_u0__abc_75526_new_n876__bF_buf4), .B(u3_u0_r0_9_), .Y(u3_u0__abc_75526_new_n921_));
OR2X2 OR2X2_3285 ( .A(u3_u0__abc_75526_new_n876__bF_buf2), .B(u3_u0_r0_10_), .Y(u3_u0__abc_75526_new_n925_));
OR2X2 OR2X2_3286 ( .A(u3_u0__abc_75526_new_n876__bF_buf0), .B(u3_u0_r0_11_), .Y(u3_u0__abc_75526_new_n929_));
OR2X2 OR2X2_3287 ( .A(u3_u0__abc_75526_new_n876__bF_buf6), .B(u3_u0_r0_12_), .Y(u3_u0__abc_75526_new_n933_));
OR2X2 OR2X2_3288 ( .A(u3_u0__abc_75526_new_n876__bF_buf4), .B(u3_u0_r0_13_), .Y(u3_u0__abc_75526_new_n937_));
OR2X2 OR2X2_3289 ( .A(u3_u0__abc_75526_new_n876__bF_buf2), .B(u3_u0_r0_14_), .Y(u3_u0__abc_75526_new_n941_));
OR2X2 OR2X2_329 ( .A(u0__abc_76628_new_n1177__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n1660_));
OR2X2 OR2X2_3290 ( .A(u3_u0__abc_75526_new_n876__bF_buf0), .B(u3_u0_r0_15_), .Y(u3_u0__abc_75526_new_n945_));
OR2X2 OR2X2_3291 ( .A(u3_u0__abc_75526_new_n876__bF_buf6), .B(u3_u0_r0_16_), .Y(u3_u0__abc_75526_new_n949_));
OR2X2 OR2X2_3292 ( .A(u3_u0__abc_75526_new_n876__bF_buf4), .B(u3_u0_r0_17_), .Y(u3_u0__abc_75526_new_n953_));
OR2X2 OR2X2_3293 ( .A(u3_u0__abc_75526_new_n876__bF_buf2), .B(u3_u0_r0_18_), .Y(u3_u0__abc_75526_new_n957_));
OR2X2 OR2X2_3294 ( .A(u3_u0__abc_75526_new_n876__bF_buf0), .B(u3_u0_r0_19_), .Y(u3_u0__abc_75526_new_n961_));
OR2X2 OR2X2_3295 ( .A(u3_u0__abc_75526_new_n876__bF_buf6), .B(u3_u0_r0_20_), .Y(u3_u0__abc_75526_new_n965_));
OR2X2 OR2X2_3296 ( .A(u3_u0__abc_75526_new_n876__bF_buf4), .B(u3_u0_r0_21_), .Y(u3_u0__abc_75526_new_n969_));
OR2X2 OR2X2_3297 ( .A(u3_u0__abc_75526_new_n876__bF_buf2), .B(u3_u0_r0_22_), .Y(u3_u0__abc_75526_new_n973_));
OR2X2 OR2X2_3298 ( .A(u3_u0__abc_75526_new_n876__bF_buf0), .B(u3_u0_r0_23_), .Y(u3_u0__abc_75526_new_n977_));
OR2X2 OR2X2_3299 ( .A(u3_u0__abc_75526_new_n876__bF_buf6), .B(u3_u0_r0_24_), .Y(u3_u0__abc_75526_new_n981_));
OR2X2 OR2X2_33 ( .A(_abc_85006_new_n286_), .B(_abc_85006_new_n237_), .Y(_abc_85006_new_n287_));
OR2X2 OR2X2_330 ( .A(spec_req_cs_6_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1661_));
OR2X2 OR2X2_3300 ( .A(u3_u0__abc_75526_new_n876__bF_buf4), .B(u3_u0_r0_25_), .Y(u3_u0__abc_75526_new_n985_));
OR2X2 OR2X2_3301 ( .A(u3_u0__abc_75526_new_n876__bF_buf2), .B(u3_u0_r0_26_), .Y(u3_u0__abc_75526_new_n989_));
OR2X2 OR2X2_3302 ( .A(u3_u0__abc_75526_new_n876__bF_buf0), .B(u3_u0_r0_27_), .Y(u3_u0__abc_75526_new_n993_));
OR2X2 OR2X2_3303 ( .A(u3_u0__abc_75526_new_n876__bF_buf6), .B(u3_u0_r0_28_), .Y(u3_u0__abc_75526_new_n997_));
OR2X2 OR2X2_3304 ( .A(u3_u0__abc_75526_new_n876__bF_buf4), .B(u3_u0_r0_29_), .Y(u3_u0__abc_75526_new_n1001_));
OR2X2 OR2X2_3305 ( .A(u3_u0__abc_75526_new_n876__bF_buf2), .B(u3_u0_r0_30_), .Y(u3_u0__abc_75526_new_n1005_));
OR2X2 OR2X2_3306 ( .A(u3_u0__abc_75526_new_n876__bF_buf0), .B(u3_u0_r0_31_), .Y(u3_u0__abc_75526_new_n1009_));
OR2X2 OR2X2_3307 ( .A(u3_u0__abc_75526_new_n876__bF_buf6), .B(u3_u0_r0_32_), .Y(u3_u0__abc_75526_new_n1013_));
OR2X2 OR2X2_3308 ( .A(u3_u0__abc_75526_new_n876__bF_buf4), .B(u3_u0_r0_33_), .Y(u3_u0__abc_75526_new_n1017_));
OR2X2 OR2X2_3309 ( .A(u3_u0__abc_75526_new_n876__bF_buf2), .B(u3_u0_r0_34_), .Y(u3_u0__abc_75526_new_n1021_));
OR2X2 OR2X2_331 ( .A(u0__abc_76628_new_n1663_), .B(u0__abc_76628_new_n1659_), .Y(u0__abc_76628_new_n1664_));
OR2X2 OR2X2_3310 ( .A(u3_u0__abc_75526_new_n876__bF_buf0), .B(u3_u0_r0_35_), .Y(u3_u0__abc_75526_new_n1025_));
OR2X2 OR2X2_3311 ( .A(u3_u0_rd_adr_0_), .B(u3_u0_rd_adr_3_), .Y(u3_u0__abc_75526_new_n1036_));
OR2X2 OR2X2_3312 ( .A(u3_u0__abc_75526_new_n1030_), .B(u3_u0_rd_adr_2_), .Y(u3_u0__abc_75526_new_n1037_));
OR2X2 OR2X2_3313 ( .A(u3_u0__abc_75526_new_n1037_), .B(u3_u0__abc_75526_new_n1036_), .Y(u3_u0__abc_75526_new_n1038_));
OR2X2 OR2X2_3314 ( .A(u3_u0_rd_adr_0_), .B(u3_u0_rd_adr_1_), .Y(u3_u0__abc_75526_new_n1039_));
OR2X2 OR2X2_3315 ( .A(u3_u0__abc_75526_new_n1032_), .B(u3_u0_rd_adr_3_), .Y(u3_u0__abc_75526_new_n1040_));
OR2X2 OR2X2_3316 ( .A(u3_u0__abc_75526_new_n1040_), .B(u3_u0__abc_75526_new_n1039_), .Y(u3_u0__abc_75526_new_n1041_));
OR2X2 OR2X2_3317 ( .A(u3_u0__abc_75526_new_n1050_), .B(u3_u0__abc_75526_new_n1053_), .Y(u3_u0__abc_75526_new_n1054_));
OR2X2 OR2X2_3318 ( .A(u3_u0__abc_75526_new_n1054_), .B(u3_u0__abc_75526_new_n1045_), .Y(u3_u0__abc_75526_new_n1055_));
OR2X2 OR2X2_3319 ( .A(u3_u0__abc_75526_new_n1055_), .B(u3_u0__abc_75526_new_n1044_), .Y(u3_rd_fifo_out_0_));
OR2X2 OR2X2_332 ( .A(u0__abc_76628_new_n1665_), .B(u0__abc_76628_new_n1666_), .Y(u0__abc_76628_new_n1667_));
OR2X2 OR2X2_3320 ( .A(u3_u0__abc_75526_new_n1059_), .B(u3_u0__abc_75526_new_n1060_), .Y(u3_u0__abc_75526_new_n1061_));
OR2X2 OR2X2_3321 ( .A(u3_u0__abc_75526_new_n1061_), .B(u3_u0__abc_75526_new_n1058_), .Y(u3_u0__abc_75526_new_n1062_));
OR2X2 OR2X2_3322 ( .A(u3_u0__abc_75526_new_n1062_), .B(u3_u0__abc_75526_new_n1057_), .Y(u3_rd_fifo_out_1_));
OR2X2 OR2X2_3323 ( .A(u3_u0__abc_75526_new_n1066_), .B(u3_u0__abc_75526_new_n1067_), .Y(u3_u0__abc_75526_new_n1068_));
OR2X2 OR2X2_3324 ( .A(u3_u0__abc_75526_new_n1068_), .B(u3_u0__abc_75526_new_n1065_), .Y(u3_u0__abc_75526_new_n1069_));
OR2X2 OR2X2_3325 ( .A(u3_u0__abc_75526_new_n1069_), .B(u3_u0__abc_75526_new_n1064_), .Y(u3_rd_fifo_out_2_));
OR2X2 OR2X2_3326 ( .A(u3_u0__abc_75526_new_n1073_), .B(u3_u0__abc_75526_new_n1074_), .Y(u3_u0__abc_75526_new_n1075_));
OR2X2 OR2X2_3327 ( .A(u3_u0__abc_75526_new_n1075_), .B(u3_u0__abc_75526_new_n1072_), .Y(u3_u0__abc_75526_new_n1076_));
OR2X2 OR2X2_3328 ( .A(u3_u0__abc_75526_new_n1076_), .B(u3_u0__abc_75526_new_n1071_), .Y(u3_rd_fifo_out_3_));
OR2X2 OR2X2_3329 ( .A(u3_u0__abc_75526_new_n1080_), .B(u3_u0__abc_75526_new_n1081_), .Y(u3_u0__abc_75526_new_n1082_));
OR2X2 OR2X2_333 ( .A(u0__abc_76628_new_n1668_), .B(u0__abc_76628_new_n1669_), .Y(u0__abc_76628_new_n1670_));
OR2X2 OR2X2_3330 ( .A(u3_u0__abc_75526_new_n1082_), .B(u3_u0__abc_75526_new_n1079_), .Y(u3_u0__abc_75526_new_n1083_));
OR2X2 OR2X2_3331 ( .A(u3_u0__abc_75526_new_n1083_), .B(u3_u0__abc_75526_new_n1078_), .Y(u3_rd_fifo_out_4_));
OR2X2 OR2X2_3332 ( .A(u3_u0__abc_75526_new_n1087_), .B(u3_u0__abc_75526_new_n1088_), .Y(u3_u0__abc_75526_new_n1089_));
OR2X2 OR2X2_3333 ( .A(u3_u0__abc_75526_new_n1089_), .B(u3_u0__abc_75526_new_n1086_), .Y(u3_u0__abc_75526_new_n1090_));
OR2X2 OR2X2_3334 ( .A(u3_u0__abc_75526_new_n1090_), .B(u3_u0__abc_75526_new_n1085_), .Y(u3_rd_fifo_out_5_));
OR2X2 OR2X2_3335 ( .A(u3_u0__abc_75526_new_n1094_), .B(u3_u0__abc_75526_new_n1095_), .Y(u3_u0__abc_75526_new_n1096_));
OR2X2 OR2X2_3336 ( .A(u3_u0__abc_75526_new_n1096_), .B(u3_u0__abc_75526_new_n1093_), .Y(u3_u0__abc_75526_new_n1097_));
OR2X2 OR2X2_3337 ( .A(u3_u0__abc_75526_new_n1097_), .B(u3_u0__abc_75526_new_n1092_), .Y(u3_rd_fifo_out_6_));
OR2X2 OR2X2_3338 ( .A(u3_u0__abc_75526_new_n1101_), .B(u3_u0__abc_75526_new_n1102_), .Y(u3_u0__abc_75526_new_n1103_));
OR2X2 OR2X2_3339 ( .A(u3_u0__abc_75526_new_n1103_), .B(u3_u0__abc_75526_new_n1100_), .Y(u3_u0__abc_75526_new_n1104_));
OR2X2 OR2X2_334 ( .A(u0__abc_76628_new_n1671_), .B(u0__abc_76628_new_n1672_), .Y(u0__abc_76628_new_n1673_));
OR2X2 OR2X2_3340 ( .A(u3_u0__abc_75526_new_n1104_), .B(u3_u0__abc_75526_new_n1099_), .Y(u3_rd_fifo_out_7_));
OR2X2 OR2X2_3341 ( .A(u3_u0__abc_75526_new_n1108_), .B(u3_u0__abc_75526_new_n1109_), .Y(u3_u0__abc_75526_new_n1110_));
OR2X2 OR2X2_3342 ( .A(u3_u0__abc_75526_new_n1110_), .B(u3_u0__abc_75526_new_n1107_), .Y(u3_u0__abc_75526_new_n1111_));
OR2X2 OR2X2_3343 ( .A(u3_u0__abc_75526_new_n1111_), .B(u3_u0__abc_75526_new_n1106_), .Y(u3_rd_fifo_out_8_));
OR2X2 OR2X2_3344 ( .A(u3_u0__abc_75526_new_n1115_), .B(u3_u0__abc_75526_new_n1116_), .Y(u3_u0__abc_75526_new_n1117_));
OR2X2 OR2X2_3345 ( .A(u3_u0__abc_75526_new_n1117_), .B(u3_u0__abc_75526_new_n1114_), .Y(u3_u0__abc_75526_new_n1118_));
OR2X2 OR2X2_3346 ( .A(u3_u0__abc_75526_new_n1118_), .B(u3_u0__abc_75526_new_n1113_), .Y(u3_rd_fifo_out_9_));
OR2X2 OR2X2_3347 ( .A(u3_u0__abc_75526_new_n1122_), .B(u3_u0__abc_75526_new_n1123_), .Y(u3_u0__abc_75526_new_n1124_));
OR2X2 OR2X2_3348 ( .A(u3_u0__abc_75526_new_n1124_), .B(u3_u0__abc_75526_new_n1121_), .Y(u3_u0__abc_75526_new_n1125_));
OR2X2 OR2X2_3349 ( .A(u3_u0__abc_75526_new_n1125_), .B(u3_u0__abc_75526_new_n1120_), .Y(u3_rd_fifo_out_10_));
OR2X2 OR2X2_335 ( .A(u0__abc_76628_new_n1675_), .B(spec_req_cs_0_bF_buf0_), .Y(u0__abc_76628_new_n1676_));
OR2X2 OR2X2_3350 ( .A(u3_u0__abc_75526_new_n1129_), .B(u3_u0__abc_75526_new_n1130_), .Y(u3_u0__abc_75526_new_n1131_));
OR2X2 OR2X2_3351 ( .A(u3_u0__abc_75526_new_n1131_), .B(u3_u0__abc_75526_new_n1128_), .Y(u3_u0__abc_75526_new_n1132_));
OR2X2 OR2X2_3352 ( .A(u3_u0__abc_75526_new_n1132_), .B(u3_u0__abc_75526_new_n1127_), .Y(u3_rd_fifo_out_11_));
OR2X2 OR2X2_3353 ( .A(u3_u0__abc_75526_new_n1136_), .B(u3_u0__abc_75526_new_n1137_), .Y(u3_u0__abc_75526_new_n1138_));
OR2X2 OR2X2_3354 ( .A(u3_u0__abc_75526_new_n1138_), .B(u3_u0__abc_75526_new_n1135_), .Y(u3_u0__abc_75526_new_n1139_));
OR2X2 OR2X2_3355 ( .A(u3_u0__abc_75526_new_n1139_), .B(u3_u0__abc_75526_new_n1134_), .Y(u3_rd_fifo_out_12_));
OR2X2 OR2X2_3356 ( .A(u3_u0__abc_75526_new_n1143_), .B(u3_u0__abc_75526_new_n1144_), .Y(u3_u0__abc_75526_new_n1145_));
OR2X2 OR2X2_3357 ( .A(u3_u0__abc_75526_new_n1145_), .B(u3_u0__abc_75526_new_n1142_), .Y(u3_u0__abc_75526_new_n1146_));
OR2X2 OR2X2_3358 ( .A(u3_u0__abc_75526_new_n1146_), .B(u3_u0__abc_75526_new_n1141_), .Y(u3_rd_fifo_out_13_));
OR2X2 OR2X2_3359 ( .A(u3_u0__abc_75526_new_n1150_), .B(u3_u0__abc_75526_new_n1151_), .Y(u3_u0__abc_75526_new_n1152_));
OR2X2 OR2X2_336 ( .A(u0__abc_76628_new_n1674_), .B(u0__abc_76628_new_n1676_), .Y(u0__abc_76628_new_n1677_));
OR2X2 OR2X2_3360 ( .A(u3_u0__abc_75526_new_n1152_), .B(u3_u0__abc_75526_new_n1149_), .Y(u3_u0__abc_75526_new_n1153_));
OR2X2 OR2X2_3361 ( .A(u3_u0__abc_75526_new_n1153_), .B(u3_u0__abc_75526_new_n1148_), .Y(u3_rd_fifo_out_14_));
OR2X2 OR2X2_3362 ( .A(u3_u0__abc_75526_new_n1157_), .B(u3_u0__abc_75526_new_n1158_), .Y(u3_u0__abc_75526_new_n1159_));
OR2X2 OR2X2_3363 ( .A(u3_u0__abc_75526_new_n1159_), .B(u3_u0__abc_75526_new_n1156_), .Y(u3_u0__abc_75526_new_n1160_));
OR2X2 OR2X2_3364 ( .A(u3_u0__abc_75526_new_n1160_), .B(u3_u0__abc_75526_new_n1155_), .Y(u3_rd_fifo_out_15_));
OR2X2 OR2X2_3365 ( .A(u3_u0__abc_75526_new_n1164_), .B(u3_u0__abc_75526_new_n1165_), .Y(u3_u0__abc_75526_new_n1166_));
OR2X2 OR2X2_3366 ( .A(u3_u0__abc_75526_new_n1166_), .B(u3_u0__abc_75526_new_n1163_), .Y(u3_u0__abc_75526_new_n1167_));
OR2X2 OR2X2_3367 ( .A(u3_u0__abc_75526_new_n1167_), .B(u3_u0__abc_75526_new_n1162_), .Y(u3_rd_fifo_out_16_));
OR2X2 OR2X2_3368 ( .A(u3_u0__abc_75526_new_n1171_), .B(u3_u0__abc_75526_new_n1172_), .Y(u3_u0__abc_75526_new_n1173_));
OR2X2 OR2X2_3369 ( .A(u3_u0__abc_75526_new_n1173_), .B(u3_u0__abc_75526_new_n1170_), .Y(u3_u0__abc_75526_new_n1174_));
OR2X2 OR2X2_337 ( .A(u0__abc_76628_new_n1197__bF_buf3), .B(u0_tms0_20_), .Y(u0__abc_76628_new_n1678_));
OR2X2 OR2X2_3370 ( .A(u3_u0__abc_75526_new_n1174_), .B(u3_u0__abc_75526_new_n1169_), .Y(u3_rd_fifo_out_17_));
OR2X2 OR2X2_3371 ( .A(u3_u0__abc_75526_new_n1178_), .B(u3_u0__abc_75526_new_n1179_), .Y(u3_u0__abc_75526_new_n1180_));
OR2X2 OR2X2_3372 ( .A(u3_u0__abc_75526_new_n1180_), .B(u3_u0__abc_75526_new_n1177_), .Y(u3_u0__abc_75526_new_n1181_));
OR2X2 OR2X2_3373 ( .A(u3_u0__abc_75526_new_n1181_), .B(u3_u0__abc_75526_new_n1176_), .Y(u3_rd_fifo_out_18_));
OR2X2 OR2X2_3374 ( .A(u3_u0__abc_75526_new_n1185_), .B(u3_u0__abc_75526_new_n1186_), .Y(u3_u0__abc_75526_new_n1187_));
OR2X2 OR2X2_3375 ( .A(u3_u0__abc_75526_new_n1187_), .B(u3_u0__abc_75526_new_n1184_), .Y(u3_u0__abc_75526_new_n1188_));
OR2X2 OR2X2_3376 ( .A(u3_u0__abc_75526_new_n1188_), .B(u3_u0__abc_75526_new_n1183_), .Y(u3_rd_fifo_out_19_));
OR2X2 OR2X2_3377 ( .A(u3_u0__abc_75526_new_n1192_), .B(u3_u0__abc_75526_new_n1193_), .Y(u3_u0__abc_75526_new_n1194_));
OR2X2 OR2X2_3378 ( .A(u3_u0__abc_75526_new_n1194_), .B(u3_u0__abc_75526_new_n1191_), .Y(u3_u0__abc_75526_new_n1195_));
OR2X2 OR2X2_3379 ( .A(u3_u0__abc_75526_new_n1195_), .B(u3_u0__abc_75526_new_n1190_), .Y(u3_rd_fifo_out_20_));
OR2X2 OR2X2_338 ( .A(u0__abc_76628_new_n1680_), .B(u0__abc_76628_new_n1658_), .Y(u0__0sp_tms_31_0__20_));
OR2X2 OR2X2_3380 ( .A(u3_u0__abc_75526_new_n1199_), .B(u3_u0__abc_75526_new_n1200_), .Y(u3_u0__abc_75526_new_n1201_));
OR2X2 OR2X2_3381 ( .A(u3_u0__abc_75526_new_n1201_), .B(u3_u0__abc_75526_new_n1198_), .Y(u3_u0__abc_75526_new_n1202_));
OR2X2 OR2X2_3382 ( .A(u3_u0__abc_75526_new_n1202_), .B(u3_u0__abc_75526_new_n1197_), .Y(u3_rd_fifo_out_21_));
OR2X2 OR2X2_3383 ( .A(u3_u0__abc_75526_new_n1206_), .B(u3_u0__abc_75526_new_n1207_), .Y(u3_u0__abc_75526_new_n1208_));
OR2X2 OR2X2_3384 ( .A(u3_u0__abc_75526_new_n1208_), .B(u3_u0__abc_75526_new_n1205_), .Y(u3_u0__abc_75526_new_n1209_));
OR2X2 OR2X2_3385 ( .A(u3_u0__abc_75526_new_n1209_), .B(u3_u0__abc_75526_new_n1204_), .Y(u3_rd_fifo_out_22_));
OR2X2 OR2X2_3386 ( .A(u3_u0__abc_75526_new_n1213_), .B(u3_u0__abc_75526_new_n1214_), .Y(u3_u0__abc_75526_new_n1215_));
OR2X2 OR2X2_3387 ( .A(u3_u0__abc_75526_new_n1215_), .B(u3_u0__abc_75526_new_n1212_), .Y(u3_u0__abc_75526_new_n1216_));
OR2X2 OR2X2_3388 ( .A(u3_u0__abc_75526_new_n1216_), .B(u3_u0__abc_75526_new_n1211_), .Y(u3_rd_fifo_out_23_));
OR2X2 OR2X2_3389 ( .A(u3_u0__abc_75526_new_n1220_), .B(u3_u0__abc_75526_new_n1221_), .Y(u3_u0__abc_75526_new_n1222_));
OR2X2 OR2X2_339 ( .A(u0__abc_76628_new_n1177__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n1684_));
OR2X2 OR2X2_3390 ( .A(u3_u0__abc_75526_new_n1222_), .B(u3_u0__abc_75526_new_n1219_), .Y(u3_u0__abc_75526_new_n1223_));
OR2X2 OR2X2_3391 ( .A(u3_u0__abc_75526_new_n1223_), .B(u3_u0__abc_75526_new_n1218_), .Y(u3_rd_fifo_out_24_));
OR2X2 OR2X2_3392 ( .A(u3_u0__abc_75526_new_n1227_), .B(u3_u0__abc_75526_new_n1228_), .Y(u3_u0__abc_75526_new_n1229_));
OR2X2 OR2X2_3393 ( .A(u3_u0__abc_75526_new_n1229_), .B(u3_u0__abc_75526_new_n1226_), .Y(u3_u0__abc_75526_new_n1230_));
OR2X2 OR2X2_3394 ( .A(u3_u0__abc_75526_new_n1230_), .B(u3_u0__abc_75526_new_n1225_), .Y(u3_rd_fifo_out_25_));
OR2X2 OR2X2_3395 ( .A(u3_u0__abc_75526_new_n1234_), .B(u3_u0__abc_75526_new_n1235_), .Y(u3_u0__abc_75526_new_n1236_));
OR2X2 OR2X2_3396 ( .A(u3_u0__abc_75526_new_n1236_), .B(u3_u0__abc_75526_new_n1233_), .Y(u3_u0__abc_75526_new_n1237_));
OR2X2 OR2X2_3397 ( .A(u3_u0__abc_75526_new_n1237_), .B(u3_u0__abc_75526_new_n1232_), .Y(u3_rd_fifo_out_26_));
OR2X2 OR2X2_3398 ( .A(u3_u0__abc_75526_new_n1241_), .B(u3_u0__abc_75526_new_n1242_), .Y(u3_u0__abc_75526_new_n1243_));
OR2X2 OR2X2_3399 ( .A(u3_u0__abc_75526_new_n1243_), .B(u3_u0__abc_75526_new_n1240_), .Y(u3_u0__abc_75526_new_n1244_));
OR2X2 OR2X2_34 ( .A(_abc_85006_new_n245_), .B(cs_need_rfr_7_), .Y(_abc_85006_new_n288_));
OR2X2 OR2X2_340 ( .A(spec_req_cs_6_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1685_));
OR2X2 OR2X2_3400 ( .A(u3_u0__abc_75526_new_n1244_), .B(u3_u0__abc_75526_new_n1239_), .Y(u3_rd_fifo_out_27_));
OR2X2 OR2X2_3401 ( .A(u3_u0__abc_75526_new_n1248_), .B(u3_u0__abc_75526_new_n1249_), .Y(u3_u0__abc_75526_new_n1250_));
OR2X2 OR2X2_3402 ( .A(u3_u0__abc_75526_new_n1250_), .B(u3_u0__abc_75526_new_n1247_), .Y(u3_u0__abc_75526_new_n1251_));
OR2X2 OR2X2_3403 ( .A(u3_u0__abc_75526_new_n1251_), .B(u3_u0__abc_75526_new_n1246_), .Y(u3_rd_fifo_out_28_));
OR2X2 OR2X2_3404 ( .A(u3_u0__abc_75526_new_n1255_), .B(u3_u0__abc_75526_new_n1256_), .Y(u3_u0__abc_75526_new_n1257_));
OR2X2 OR2X2_3405 ( .A(u3_u0__abc_75526_new_n1257_), .B(u3_u0__abc_75526_new_n1254_), .Y(u3_u0__abc_75526_new_n1258_));
OR2X2 OR2X2_3406 ( .A(u3_u0__abc_75526_new_n1258_), .B(u3_u0__abc_75526_new_n1253_), .Y(u3_rd_fifo_out_29_));
OR2X2 OR2X2_3407 ( .A(u3_u0__abc_75526_new_n1262_), .B(u3_u0__abc_75526_new_n1263_), .Y(u3_u0__abc_75526_new_n1264_));
OR2X2 OR2X2_3408 ( .A(u3_u0__abc_75526_new_n1264_), .B(u3_u0__abc_75526_new_n1261_), .Y(u3_u0__abc_75526_new_n1265_));
OR2X2 OR2X2_3409 ( .A(u3_u0__abc_75526_new_n1265_), .B(u3_u0__abc_75526_new_n1260_), .Y(u3_rd_fifo_out_30_));
OR2X2 OR2X2_341 ( .A(u0__abc_76628_new_n1687_), .B(u0__abc_76628_new_n1683_), .Y(u0__abc_76628_new_n1688_));
OR2X2 OR2X2_3410 ( .A(u3_u0__abc_75526_new_n1269_), .B(u3_u0__abc_75526_new_n1270_), .Y(u3_u0__abc_75526_new_n1271_));
OR2X2 OR2X2_3411 ( .A(u3_u0__abc_75526_new_n1271_), .B(u3_u0__abc_75526_new_n1268_), .Y(u3_u0__abc_75526_new_n1272_));
OR2X2 OR2X2_3412 ( .A(u3_u0__abc_75526_new_n1272_), .B(u3_u0__abc_75526_new_n1267_), .Y(u3_rd_fifo_out_31_));
OR2X2 OR2X2_3413 ( .A(u3_u0__abc_75526_new_n1276_), .B(u3_u0__abc_75526_new_n1277_), .Y(u3_u0__abc_75526_new_n1278_));
OR2X2 OR2X2_3414 ( .A(u3_u0__abc_75526_new_n1278_), .B(u3_u0__abc_75526_new_n1275_), .Y(u3_u0__abc_75526_new_n1279_));
OR2X2 OR2X2_3415 ( .A(u3_u0__abc_75526_new_n1279_), .B(u3_u0__abc_75526_new_n1274_), .Y(u3_rd_fifo_out_32_));
OR2X2 OR2X2_3416 ( .A(u3_u0__abc_75526_new_n1283_), .B(u3_u0__abc_75526_new_n1284_), .Y(u3_u0__abc_75526_new_n1285_));
OR2X2 OR2X2_3417 ( .A(u3_u0__abc_75526_new_n1285_), .B(u3_u0__abc_75526_new_n1282_), .Y(u3_u0__abc_75526_new_n1286_));
OR2X2 OR2X2_3418 ( .A(u3_u0__abc_75526_new_n1286_), .B(u3_u0__abc_75526_new_n1281_), .Y(u3_rd_fifo_out_33_));
OR2X2 OR2X2_3419 ( .A(u3_u0__abc_75526_new_n1290_), .B(u3_u0__abc_75526_new_n1291_), .Y(u3_u0__abc_75526_new_n1292_));
OR2X2 OR2X2_342 ( .A(u0__abc_76628_new_n1689_), .B(u0__abc_76628_new_n1690_), .Y(u0__abc_76628_new_n1691_));
OR2X2 OR2X2_3420 ( .A(u3_u0__abc_75526_new_n1292_), .B(u3_u0__abc_75526_new_n1289_), .Y(u3_u0__abc_75526_new_n1293_));
OR2X2 OR2X2_3421 ( .A(u3_u0__abc_75526_new_n1293_), .B(u3_u0__abc_75526_new_n1288_), .Y(u3_rd_fifo_out_34_));
OR2X2 OR2X2_3422 ( .A(u3_u0__abc_75526_new_n1297_), .B(u3_u0__abc_75526_new_n1298_), .Y(u3_u0__abc_75526_new_n1299_));
OR2X2 OR2X2_3423 ( .A(u3_u0__abc_75526_new_n1299_), .B(u3_u0__abc_75526_new_n1296_), .Y(u3_u0__abc_75526_new_n1300_));
OR2X2 OR2X2_3424 ( .A(u3_u0__abc_75526_new_n1300_), .B(u3_u0__abc_75526_new_n1295_), .Y(u3_rd_fifo_out_35_));
OR2X2 OR2X2_3425 ( .A(cs_need_rfr_2_), .B(cs_need_rfr_3_), .Y(u4__abc_76448_new_n65_));
OR2X2 OR2X2_3426 ( .A(cs_need_rfr_0_), .B(cs_need_rfr_1_), .Y(u4__abc_76448_new_n66_));
OR2X2 OR2X2_3427 ( .A(u4__abc_76448_new_n65_), .B(u4__abc_76448_new_n66_), .Y(u4__abc_76448_new_n67_));
OR2X2 OR2X2_3428 ( .A(cs_need_rfr_6_), .B(cs_need_rfr_7_), .Y(u4__abc_76448_new_n68_));
OR2X2 OR2X2_3429 ( .A(cs_need_rfr_4_), .B(cs_need_rfr_5_), .Y(u4__abc_76448_new_n69_));
OR2X2 OR2X2_343 ( .A(u0__abc_76628_new_n1692_), .B(u0__abc_76628_new_n1693_), .Y(u0__abc_76628_new_n1694_));
OR2X2 OR2X2_3430 ( .A(u4__abc_76448_new_n68_), .B(u4__abc_76448_new_n69_), .Y(u4__abc_76448_new_n70_));
OR2X2 OR2X2_3431 ( .A(u4__abc_76448_new_n67_), .B(u4__abc_76448_new_n70_), .Y(u4__0rfr_en_0_0_));
OR2X2 OR2X2_3432 ( .A(u4_ps_cnt_3_), .B(rfr_ps_val_3_), .Y(u4__abc_76448_new_n72_));
OR2X2 OR2X2_3433 ( .A(u4_ps_cnt_2_), .B(rfr_ps_val_2_), .Y(u4__abc_76448_new_n76_));
OR2X2 OR2X2_3434 ( .A(u4__abc_76448_new_n75_), .B(u4__abc_76448_new_n79_), .Y(u4__abc_76448_new_n80_));
OR2X2 OR2X2_3435 ( .A(u4_ps_cnt_7_), .B(rfr_ps_val_7_), .Y(u4__abc_76448_new_n81_));
OR2X2 OR2X2_3436 ( .A(u4_ps_cnt_6_), .B(rfr_ps_val_6_), .Y(u4__abc_76448_new_n85_));
OR2X2 OR2X2_3437 ( .A(u4__abc_76448_new_n84_), .B(u4__abc_76448_new_n88_), .Y(u4__abc_76448_new_n89_));
OR2X2 OR2X2_3438 ( .A(u4__abc_76448_new_n80_), .B(u4__abc_76448_new_n89_), .Y(u4__abc_76448_new_n90_));
OR2X2 OR2X2_3439 ( .A(u4__abc_76448_new_n92_), .B(u4__abc_76448_new_n94_), .Y(u4__abc_76448_new_n95_));
OR2X2 OR2X2_344 ( .A(u0__abc_76628_new_n1695_), .B(u0__abc_76628_new_n1696_), .Y(u0__abc_76628_new_n1697_));
OR2X2 OR2X2_3440 ( .A(u4__abc_76448_new_n97_), .B(u4__abc_76448_new_n99_), .Y(u4__abc_76448_new_n100_));
OR2X2 OR2X2_3441 ( .A(u4__abc_76448_new_n95_), .B(u4__abc_76448_new_n100_), .Y(u4__abc_76448_new_n101_));
OR2X2 OR2X2_3442 ( .A(u4__abc_76448_new_n103_), .B(u4__abc_76448_new_n105_), .Y(u4__abc_76448_new_n106_));
OR2X2 OR2X2_3443 ( .A(u4__abc_76448_new_n108_), .B(u4__abc_76448_new_n110_), .Y(u4__abc_76448_new_n111_));
OR2X2 OR2X2_3444 ( .A(u4__abc_76448_new_n106_), .B(u4__abc_76448_new_n111_), .Y(u4__abc_76448_new_n112_));
OR2X2 OR2X2_3445 ( .A(u4__abc_76448_new_n112_), .B(u4__abc_76448_new_n101_), .Y(u4__abc_76448_new_n113_));
OR2X2 OR2X2_3446 ( .A(u4__abc_76448_new_n113_), .B(u4__abc_76448_new_n90_), .Y(u4__abc_76448_new_n114_));
OR2X2 OR2X2_3447 ( .A(u4_rfr_clr), .B(rfr_req), .Y(u4__abc_76448_new_n117_));
OR2X2 OR2X2_3448 ( .A(u4_rfr_ce), .B(u4_rfr_cnt_0_), .Y(u4__abc_76448_new_n121_));
OR2X2 OR2X2_3449 ( .A(u4__abc_76448_new_n119_), .B(u4_rfr_cnt_1_), .Y(u4__abc_76448_new_n126_));
OR2X2 OR2X2_345 ( .A(u0__abc_76628_new_n1699_), .B(spec_req_cs_0_bF_buf5_), .Y(u0__abc_76628_new_n1700_));
OR2X2 OR2X2_3450 ( .A(u4__abc_76448_new_n124_), .B(u4_rfr_cnt_2_), .Y(u4__abc_76448_new_n133_));
OR2X2 OR2X2_3451 ( .A(u4__abc_76448_new_n131_), .B(u4_rfr_cnt_3_), .Y(u4__abc_76448_new_n139_));
OR2X2 OR2X2_3452 ( .A(u4__abc_76448_new_n137_), .B(u4_rfr_cnt_4_), .Y(u4__abc_76448_new_n142_));
OR2X2 OR2X2_3453 ( .A(u4__abc_76448_new_n145_), .B(u4_rfr_cnt_5_), .Y(u4__abc_76448_new_n152_));
OR2X2 OR2X2_3454 ( .A(u4__abc_76448_new_n150_), .B(u4_rfr_cnt_6_), .Y(u4__abc_76448_new_n155_));
OR2X2 OR2X2_3455 ( .A(u4__abc_76448_new_n157_), .B(u4_rfr_cnt_7_), .Y(u4__abc_76448_new_n163_));
OR2X2 OR2X2_3456 ( .A(u4__abc_76448_new_n114_), .B(u4__abc_76448_new_n176_), .Y(u4__abc_76448_new_n177_));
OR2X2 OR2X2_3457 ( .A(u4_ps_cnt_0_), .B(u4_rfr_en), .Y(u4__abc_76448_new_n181_));
OR2X2 OR2X2_3458 ( .A(u4__abc_76448_new_n179_), .B(u4_ps_cnt_1_), .Y(u4__abc_76448_new_n186_));
OR2X2 OR2X2_3459 ( .A(u4__abc_76448_new_n184_), .B(u4_ps_cnt_2_), .Y(u4__abc_76448_new_n189_));
OR2X2 OR2X2_346 ( .A(u0__abc_76628_new_n1698_), .B(u0__abc_76628_new_n1700_), .Y(u0__abc_76628_new_n1701_));
OR2X2 OR2X2_3460 ( .A(u4__abc_76448_new_n190_), .B(u4_ps_cnt_3_), .Y(u4__abc_76448_new_n194_));
OR2X2 OR2X2_3461 ( .A(u4__abc_76448_new_n195_), .B(u4_ps_cnt_4_), .Y(u4__abc_76448_new_n199_));
OR2X2 OR2X2_3462 ( .A(u4__abc_76448_new_n200_), .B(u4_ps_cnt_5_), .Y(u4__abc_76448_new_n208_));
OR2X2 OR2X2_3463 ( .A(u4__abc_76448_new_n213_), .B(u4__abc_76448_new_n212_), .Y(u4__abc_76448_new_n214_));
OR2X2 OR2X2_3464 ( .A(u4__abc_76448_new_n216_), .B(u4_ps_cnt_7_), .Y(u4__abc_76448_new_n219_));
OR2X2 OR2X2_3465 ( .A(u4__abc_76448_new_n223_), .B(u4_rfr_cnt_3_), .Y(u4__abc_76448_new_n224_));
OR2X2 OR2X2_3466 ( .A(u4__abc_76448_new_n223_), .B(u4_rfr_cnt_1_), .Y(u4__abc_76448_new_n227_));
OR2X2 OR2X2_3467 ( .A(u4__abc_76448_new_n226_), .B(u4__abc_76448_new_n230_), .Y(u4__abc_76448_new_n231_));
OR2X2 OR2X2_3468 ( .A(u4__abc_76448_new_n223_), .B(u4_rfr_cnt_5_), .Y(u4__abc_76448_new_n233_));
OR2X2 OR2X2_3469 ( .A(u4__abc_76448_new_n235_), .B(u4__abc_76448_new_n223_), .Y(u4__abc_76448_new_n236_));
OR2X2 OR2X2_347 ( .A(u0__abc_76628_new_n1197__bF_buf2), .B(u0_tms0_21_), .Y(u0__abc_76628_new_n1702_));
OR2X2 OR2X2_3470 ( .A(u4__abc_76448_new_n237_), .B(u4__abc_76448_new_n234_), .Y(u4__abc_76448_new_n238_));
OR2X2 OR2X2_3471 ( .A(u4__abc_76448_new_n232_), .B(u4__abc_76448_new_n240_), .Y(u4__abc_76448_new_n241_));
OR2X2 OR2X2_3472 ( .A(u5_burst_cnt_9_), .B(u5_burst_cnt_8_), .Y(u5__abc_81276_new_n381_));
OR2X2 OR2X2_3473 ( .A(u5__abc_81276_new_n537_), .B(u5__abc_81276_new_n530_), .Y(u5__abc_81276_new_n538_));
OR2X2 OR2X2_3474 ( .A(u5__abc_81276_new_n538_), .B(u5__abc_81276_new_n516_), .Y(u5_suspended_d));
OR2X2 OR2X2_3475 ( .A(u5__abc_81276_new_n656_), .B(u5__abc_81276_new_n657_), .Y(u5__abc_81276_new_n658_));
OR2X2 OR2X2_3476 ( .A(u5__abc_81276_new_n678_), .B(u5__abc_81276_new_n685_), .Y(u5__abc_81276_new_n686_));
OR2X2 OR2X2_3477 ( .A(u5__abc_81276_new_n767_), .B(u5__abc_81276_new_n761_), .Y(u5__abc_81276_new_n768_));
OR2X2 OR2X2_3478 ( .A(u5_state_19_), .B(u5_state_18_), .Y(u5__abc_81276_new_n917_));
OR2X2 OR2X2_3479 ( .A(u5_state_17_), .B(u5_state_16_), .Y(u5__abc_81276_new_n918_));
OR2X2 OR2X2_348 ( .A(u0__abc_76628_new_n1704_), .B(u0__abc_76628_new_n1682_), .Y(u0__0sp_tms_31_0__21_));
OR2X2 OR2X2_3480 ( .A(u5__abc_81276_new_n917_), .B(u5__abc_81276_new_n918_), .Y(u5__abc_81276_new_n919_));
OR2X2 OR2X2_3481 ( .A(u5__abc_81276_new_n492_), .B(u5_state_20_), .Y(u5__abc_81276_new_n920_));
OR2X2 OR2X2_3482 ( .A(u5__abc_81276_new_n919_), .B(u5__abc_81276_new_n920_), .Y(u5__abc_81276_new_n921_));
OR2X2 OR2X2_3483 ( .A(u5__abc_81276_new_n967_), .B(u5__abc_81276_new_n974_), .Y(u5__abc_81276_new_n975_));
OR2X2 OR2X2_3484 ( .A(u5__abc_81276_new_n982_), .B(u5__abc_81276_new_n989_), .Y(u5__abc_81276_new_n990_));
OR2X2 OR2X2_3485 ( .A(u5__abc_81276_new_n990_), .B(u5__abc_81276_new_n975_), .Y(u5__abc_81276_new_n991_));
OR2X2 OR2X2_3486 ( .A(u5__abc_81276_new_n1060_), .B(u5__abc_81276_new_n1067_), .Y(u5__abc_81276_new_n1068_));
OR2X2 OR2X2_3487 ( .A(u5__abc_81276_new_n1093_), .B(u5__abc_81276_new_n1098_), .Y(dv));
OR2X2 OR2X2_3488 ( .A(u5__abc_81276_new_n402_), .B(u5_state_54_), .Y(u5__abc_81276_new_n1188_));
OR2X2 OR2X2_3489 ( .A(u5__abc_81276_new_n656_), .B(u5__abc_81276_new_n1188_), .Y(u5__abc_81276_new_n1189_));
OR2X2 OR2X2_349 ( .A(u0__abc_76628_new_n1177__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n1708_));
OR2X2 OR2X2_3490 ( .A(u5__abc_81276_new_n1189_), .B(u5__abc_81276_new_n1187_), .Y(u5__abc_81276_new_n1190_));
OR2X2 OR2X2_3491 ( .A(u5__abc_81276_new_n1190_), .B(u5__abc_81276_new_n1186_), .Y(u5__abc_81276_new_n1191_));
OR2X2 OR2X2_3492 ( .A(u5__abc_81276_new_n1185_), .B(u5__abc_81276_new_n1191_), .Y(u5__abc_81276_new_n1192_));
OR2X2 OR2X2_3493 ( .A(u5__abc_81276_new_n1192_), .B(u5__abc_81276_new_n1183_), .Y(u5__abc_81276_new_n1193_));
OR2X2 OR2X2_3494 ( .A(u5__abc_81276_new_n395_), .B(u5_state_59_), .Y(u5__abc_81276_new_n1220_));
OR2X2 OR2X2_3495 ( .A(u5__abc_81276_new_n656_), .B(u5__abc_81276_new_n1220_), .Y(u5__abc_81276_new_n1221_));
OR2X2 OR2X2_3496 ( .A(u5__abc_81276_new_n1221_), .B(u5__abc_81276_new_n1219_), .Y(u5__abc_81276_new_n1222_));
OR2X2 OR2X2_3497 ( .A(u5__abc_81276_new_n1218_), .B(u5__abc_81276_new_n1222_), .Y(u5__abc_81276_new_n1223_));
OR2X2 OR2X2_3498 ( .A(u5__abc_81276_new_n1223_), .B(u5__abc_81276_new_n1217_), .Y(u5__abc_81276_new_n1224_));
OR2X2 OR2X2_3499 ( .A(u5__abc_81276_new_n1224_), .B(u5__abc_81276_new_n1183_), .Y(u5__abc_81276_new_n1225_));
OR2X2 OR2X2_35 ( .A(_abc_85006_new_n240__bF_buf3), .B(sp_tms_0_), .Y(_abc_85006_new_n290_));
OR2X2 OR2X2_350 ( .A(spec_req_cs_6_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1709_));
OR2X2 OR2X2_3500 ( .A(u5__abc_81276_new_n921_), .B(u5__abc_81276_new_n658_), .Y(u5__abc_81276_new_n1395_));
OR2X2 OR2X2_3501 ( .A(u5__abc_81276_new_n1395_), .B(u5__abc_81276_new_n1394_), .Y(u5__abc_81276_new_n1396_));
OR2X2 OR2X2_3502 ( .A(u5__abc_81276_new_n1396_), .B(u5__abc_81276_new_n1393_), .Y(u5__abc_81276_new_n1397_));
OR2X2 OR2X2_3503 ( .A(u5__abc_81276_new_n1397_), .B(u5__abc_81276_new_n1392_), .Y(u5__abc_81276_new_n1398_));
OR2X2 OR2X2_3504 ( .A(u5__abc_81276_new_n1530_), .B(u5__abc_81276_new_n1528_), .Y(u5__abc_81276_new_n1531_));
OR2X2 OR2X2_3505 ( .A(u5__abc_81276_new_n1527_), .B(u5__abc_81276_new_n1531_), .Y(u5_rfr_ack_d));
OR2X2 OR2X2_3506 ( .A(obct_cs_2_), .B(obct_cs_3_), .Y(u5__abc_81276_new_n1540_));
OR2X2 OR2X2_3507 ( .A(obct_cs_0_), .B(obct_cs_1_), .Y(u5__abc_81276_new_n1541_));
OR2X2 OR2X2_3508 ( .A(u5__abc_81276_new_n1540_), .B(u5__abc_81276_new_n1541_), .Y(u5__abc_81276_new_n1542_));
OR2X2 OR2X2_3509 ( .A(obct_cs_6_), .B(obct_cs_7_), .Y(u5__abc_81276_new_n1543_));
OR2X2 OR2X2_351 ( .A(u0__abc_76628_new_n1711_), .B(u0__abc_76628_new_n1707_), .Y(u0__abc_76628_new_n1712_));
OR2X2 OR2X2_3510 ( .A(obct_cs_4_), .B(obct_cs_5_), .Y(u5__abc_81276_new_n1544_));
OR2X2 OR2X2_3511 ( .A(u5__abc_81276_new_n1543_), .B(u5__abc_81276_new_n1544_), .Y(u5__abc_81276_new_n1545_));
OR2X2 OR2X2_3512 ( .A(u5__abc_81276_new_n1542_), .B(u5__abc_81276_new_n1545_), .Y(u5__abc_81276_new_n1546_));
OR2X2 OR2X2_3513 ( .A(u5__abc_81276_new_n1561_), .B(u5__abc_81276_new_n1539_), .Y(u5__abc_81276_new_n1562_));
OR2X2 OR2X2_3514 ( .A(u5__abc_81276_new_n1609_), .B(tms_s_9_), .Y(u5__abc_81276_new_n1610_));
OR2X2 OR2X2_3515 ( .A(u5__abc_81276_new_n1616_), .B(u5_cke_r), .Y(u5__abc_81276_new_n1619_));
OR2X2 OR2X2_3516 ( .A(u5__abc_81276_new_n1624_), .B(u5__abc_81276_new_n1611_), .Y(u5__abc_81276_new_n1625_));
OR2X2 OR2X2_3517 ( .A(u5__abc_81276_new_n1634_), .B(u5__abc_81276_new_n1563_), .Y(u5_cmd_0_));
OR2X2 OR2X2_3518 ( .A(u5__abc_81276_new_n1638_), .B(u5__abc_81276_new_n1636_), .Y(u5_we_));
OR2X2 OR2X2_3519 ( .A(u5__abc_81276_new_n1640_), .B(u5__abc_81276_new_n994_), .Y(u5__abc_81276_new_n1641_));
OR2X2 OR2X2_352 ( .A(u0__abc_76628_new_n1713_), .B(u0__abc_76628_new_n1714_), .Y(u0__abc_76628_new_n1715_));
OR2X2 OR2X2_3520 ( .A(u5__abc_81276_new_n1526__bF_buf1), .B(u5__abc_81276_new_n1641_), .Y(u5__abc_81276_new_n1642_));
OR2X2 OR2X2_3521 ( .A(u5__abc_81276_new_n1648_), .B(u5__abc_81276_new_n1652_), .Y(u5__abc_81276_new_n1653_));
OR2X2 OR2X2_3522 ( .A(u5__abc_81276_new_n1656_), .B(u5__abc_81276_new_n624_), .Y(u5__abc_81276_new_n1657_));
OR2X2 OR2X2_3523 ( .A(u5__abc_81276_new_n1654_), .B(u5__abc_81276_new_n1657_), .Y(u5__abc_81276_new_n1658_));
OR2X2 OR2X2_3524 ( .A(u5__abc_81276_new_n1653_), .B(u5__abc_81276_new_n1658_), .Y(u5__abc_81276_new_n1659_));
OR2X2 OR2X2_3525 ( .A(u5__abc_81276_new_n1643_), .B(u5__abc_81276_new_n1659_), .Y(u5__abc_81276_new_n1660_));
OR2X2 OR2X2_3526 ( .A(u5__abc_81276_new_n1642_), .B(u5__abc_81276_new_n1660_), .Y(u5_cmd_1_));
OR2X2 OR2X2_3527 ( .A(u5__abc_81276_new_n1663_), .B(u5__abc_81276_new_n1662_), .Y(cas_));
OR2X2 OR2X2_3528 ( .A(u5__abc_81276_new_n1673_), .B(u5__abc_81276_new_n1642_), .Y(u5_cmd_2_));
OR2X2 OR2X2_3529 ( .A(u5__abc_81276_new_n1676_), .B(u5__abc_81276_new_n1675_), .Y(ras_));
OR2X2 OR2X2_353 ( .A(u0__abc_76628_new_n1716_), .B(u0__abc_76628_new_n1717_), .Y(u0__abc_76628_new_n1718_));
OR2X2 OR2X2_3530 ( .A(rfr_ack), .B(susp_sel), .Y(u5__abc_81276_new_n1678_));
OR2X2 OR2X2_3531 ( .A(u5_rfr_ack_d), .B(u5__abc_81276_new_n1681_), .Y(u5__abc_81276_new_n1682_));
OR2X2 OR2X2_3532 ( .A(u5__abc_81276_new_n1682__bF_buf4), .B(tms_s_19_), .Y(u5__abc_81276_new_n1683_));
OR2X2 OR2X2_3533 ( .A(tms_s_16_), .B(tms_s_17_), .Y(u5__abc_81276_new_n1684_));
OR2X2 OR2X2_3534 ( .A(u5__abc_81276_new_n1684_), .B(tms_s_18_), .Y(u5__abc_81276_new_n1685_));
OR2X2 OR2X2_3535 ( .A(u5__abc_81276_new_n1683_), .B(u5__abc_81276_new_n1685_), .Y(u5__abc_81276_new_n1686_));
OR2X2 OR2X2_3536 ( .A(u5__abc_81276_new_n1690_), .B(csc_s_3_), .Y(u5__abc_81276_new_n1691_));
OR2X2 OR2X2_3537 ( .A(u5__abc_81276_new_n1368_), .B(u5__abc_81276_new_n1351_), .Y(u5__abc_81276_new_n1701_));
OR2X2 OR2X2_3538 ( .A(u5__abc_81276_new_n1701_), .B(u5__abc_81276_new_n1702_), .Y(u5__abc_81276_new_n1703_));
OR2X2 OR2X2_3539 ( .A(u5__abc_81276_new_n1703_), .B(u5__abc_81276_new_n1700_), .Y(u5__abc_81276_new_n1704_));
OR2X2 OR2X2_354 ( .A(u0__abc_76628_new_n1719_), .B(u0__abc_76628_new_n1720_), .Y(u0__abc_76628_new_n1721_));
OR2X2 OR2X2_3540 ( .A(u5__abc_81276_new_n1707_), .B(u5__abc_81276_new_n1709_), .Y(u5__abc_81276_new_n1710_));
OR2X2 OR2X2_3541 ( .A(u5__abc_81276_new_n1710_), .B(u5__abc_81276_new_n1705_), .Y(u5__abc_81276_new_n1711_));
OR2X2 OR2X2_3542 ( .A(u5__abc_81276_new_n1621_), .B(u5__abc_81276_new_n1611_), .Y(u5__abc_81276_new_n1714_));
OR2X2 OR2X2_3543 ( .A(u5__abc_81276_new_n1715_), .B(u5__abc_81276_new_n1713_), .Y(u5__abc_81276_new_n1716_));
OR2X2 OR2X2_3544 ( .A(u5__abc_81276_new_n1711_), .B(u5__abc_81276_new_n1716_), .Y(u5__abc_81276_new_n1717_));
OR2X2 OR2X2_3545 ( .A(u5__abc_81276_new_n1717_), .B(u5__abc_81276_new_n1704_), .Y(u5__abc_81276_new_n1718_));
OR2X2 OR2X2_3546 ( .A(u5__abc_81276_new_n1653_), .B(u5__abc_81276_new_n1640_), .Y(u5__abc_81276_new_n1719_));
OR2X2 OR2X2_3547 ( .A(u5__abc_81276_new_n1718_), .B(u5__abc_81276_new_n1719_), .Y(u5__abc_81276_new_n1720_));
OR2X2 OR2X2_3548 ( .A(u5__abc_81276_new_n1698_), .B(u5__abc_81276_new_n1720_), .Y(u5__abc_81276_new_n1721_));
OR2X2 OR2X2_3549 ( .A(u5__abc_81276_new_n1721_), .B(u5__abc_81276_new_n1696_), .Y(u5__abc_81276_new_n1722_));
OR2X2 OR2X2_355 ( .A(u0__abc_76628_new_n1723_), .B(spec_req_cs_0_bF_buf4_), .Y(u0__abc_76628_new_n1724_));
OR2X2 OR2X2_3550 ( .A(u5__abc_81276_new_n1687_), .B(u5__abc_81276_new_n1722_), .Y(u5_cmd_3_));
OR2X2 OR2X2_3551 ( .A(u5__abc_81276_new_n1725_), .B(u5__abc_81276_new_n1724_), .Y(cs_en));
OR2X2 OR2X2_3552 ( .A(u5__abc_81276_new_n1692_), .B(u5__abc_81276_new_n1727_), .Y(u5__abc_81276_new_n1728_));
OR2X2 OR2X2_3553 ( .A(u5__abc_81276_new_n1731_), .B(u5__abc_81276_new_n994_), .Y(u5__abc_81276_new_n1732_));
OR2X2 OR2X2_3554 ( .A(u5__abc_81276_new_n1733_), .B(u5__abc_81276_new_n1734_), .Y(u5__abc_81276_new_n1735_));
OR2X2 OR2X2_3555 ( .A(u5__abc_81276_new_n1732_), .B(u5__abc_81276_new_n1735_), .Y(u5__abc_81276_new_n1736_));
OR2X2 OR2X2_3556 ( .A(u5__abc_81276_new_n1736_), .B(u5__abc_81276_new_n1652_), .Y(u5__abc_81276_new_n1737_));
OR2X2 OR2X2_3557 ( .A(u5__abc_81276_new_n1730_), .B(u5__abc_81276_new_n1737_), .Y(u5__abc_81276_new_n1738_));
OR2X2 OR2X2_3558 ( .A(u5__abc_81276_new_n1687_), .B(u5__abc_81276_new_n1738_), .Y(u5_data_oe_d));
OR2X2 OR2X2_3559 ( .A(u5__abc_81276_new_n1741_), .B(u5__abc_81276_new_n1740_), .Y(u5__0data_oe_0_0_));
OR2X2 OR2X2_356 ( .A(u0__abc_76628_new_n1722_), .B(u0__abc_76628_new_n1724_), .Y(u0__abc_76628_new_n1725_));
OR2X2 OR2X2_3560 ( .A(u5_ack_cnt_1_), .B(u5_ack_cnt_0_), .Y(u5__abc_81276_new_n1817_));
OR2X2 OR2X2_3561 ( .A(u5__abc_81276_new_n1682__bF_buf3), .B(u5__abc_81276_new_n1834_), .Y(u5__abc_81276_new_n1835_));
OR2X2 OR2X2_3562 ( .A(u5__abc_81276_new_n1839_), .B(u5__abc_81276_new_n1842_), .Y(u5__abc_81276_new_n1843_));
OR2X2 OR2X2_3563 ( .A(u5__abc_81276_new_n1845_), .B(u5__abc_81276_new_n1712_), .Y(u5__abc_81276_new_n1846_));
OR2X2 OR2X2_3564 ( .A(u5__abc_81276_new_n1853_), .B(u5__abc_81276_new_n1854_), .Y(u5__abc_81276_new_n1855_));
OR2X2 OR2X2_3565 ( .A(u5__abc_81276_new_n1850_), .B(u5__abc_81276_new_n1855_), .Y(u5__abc_81276_new_n1856_));
OR2X2 OR2X2_3566 ( .A(u5__abc_81276_new_n1856_), .B(u5__abc_81276_new_n1848_), .Y(u5__abc_81276_new_n1857_));
OR2X2 OR2X2_3567 ( .A(u5__abc_81276_new_n1844_), .B(u5__abc_81276_new_n1860_), .Y(u5__abc_81276_new_n1861_));
OR2X2 OR2X2_3568 ( .A(u5__abc_81276_new_n1861_), .B(u5__abc_81276_new_n1833_), .Y(u5__abc_81276_new_n1862_));
OR2X2 OR2X2_3569 ( .A(u5__abc_81276_new_n1864_), .B(u5__0no_wb_cycle_0_0_), .Y(u5__abc_81276_new_n1865_));
OR2X2 OR2X2_357 ( .A(u0__abc_76628_new_n1197__bF_buf1), .B(u0_tms0_22_), .Y(u0__abc_76628_new_n1726_));
OR2X2 OR2X2_3570 ( .A(u5__abc_81276_new_n1867_), .B(u5_wb_stb_first), .Y(u5__abc_81276_new_n1868_));
OR2X2 OR2X2_3571 ( .A(u5__abc_81276_new_n1965_), .B(u5__abc_81276_new_n656_), .Y(u5__abc_81276_new_n1966_));
OR2X2 OR2X2_3572 ( .A(u5__abc_81276_new_n1971_), .B(u5__abc_81276_new_n1974_), .Y(u5__abc_81276_new_n1975_));
OR2X2 OR2X2_3573 ( .A(u5__abc_81276_new_n1982_), .B(u5__abc_81276_new_n1987_), .Y(u5__abc_81276_new_n1988_));
OR2X2 OR2X2_3574 ( .A(u5__abc_81276_new_n1996_), .B(u5__abc_81276_new_n2001_), .Y(u5__abc_81276_new_n2002_));
OR2X2 OR2X2_3575 ( .A(u5__abc_81276_new_n2008_), .B(u5__abc_81276_new_n2012_), .Y(u5__abc_81276_new_n2013_));
OR2X2 OR2X2_3576 ( .A(u5__abc_81276_new_n2027_), .B(u5__abc_81276_new_n2021_), .Y(u5__abc_81276_new_n2028_));
OR2X2 OR2X2_3577 ( .A(u5__abc_81276_new_n2035_), .B(u5__abc_81276_new_n2040_), .Y(u5__abc_81276_new_n2041_));
OR2X2 OR2X2_3578 ( .A(u5__abc_81276_new_n2048_), .B(u5__abc_81276_new_n2051_), .Y(u5__abc_81276_new_n2052_));
OR2X2 OR2X2_3579 ( .A(u5__abc_81276_new_n2066_), .B(u5__abc_81276_new_n656_), .Y(u5__abc_81276_new_n2067_));
OR2X2 OR2X2_358 ( .A(u0__abc_76628_new_n1728_), .B(u0__abc_76628_new_n1706_), .Y(u0__0sp_tms_31_0__22_));
OR2X2 OR2X2_3580 ( .A(u5__abc_81276_new_n2074_), .B(u5__abc_81276_new_n2079_), .Y(u5__abc_81276_new_n2080_));
OR2X2 OR2X2_3581 ( .A(u5__abc_81276_new_n2087_), .B(u5__abc_81276_new_n2092_), .Y(u5__abc_81276_new_n2093_));
OR2X2 OR2X2_3582 ( .A(u5__abc_81276_new_n2101_), .B(u5__abc_81276_new_n2106_), .Y(u5__abc_81276_new_n2107_));
OR2X2 OR2X2_3583 ( .A(u5__abc_81276_new_n2114_), .B(u5__abc_81276_new_n2119_), .Y(u5__abc_81276_new_n2120_));
OR2X2 OR2X2_3584 ( .A(u5__abc_81276_new_n2131_), .B(u5__abc_81276_new_n2136_), .Y(u5__abc_81276_new_n2137_));
OR2X2 OR2X2_3585 ( .A(u5__abc_81276_new_n2143_), .B(u5__abc_81276_new_n2148_), .Y(u5__abc_81276_new_n2149_));
OR2X2 OR2X2_3586 ( .A(u5__abc_81276_new_n2138_), .B(u5__abc_81276_new_n2150_), .Y(u5__abc_81276_new_n2151_));
OR2X2 OR2X2_3587 ( .A(u5__abc_81276_new_n2154_), .B(u5__abc_81276_new_n2157_), .Y(u5__abc_81276_new_n2158_));
OR2X2 OR2X2_3588 ( .A(u5__abc_81276_new_n2162_), .B(u5__abc_81276_new_n2165_), .Y(u5__abc_81276_new_n2166_));
OR2X2 OR2X2_3589 ( .A(u5__abc_81276_new_n2159_), .B(u5__abc_81276_new_n2167_), .Y(u5__abc_81276_new_n2168_));
OR2X2 OR2X2_359 ( .A(u0__abc_76628_new_n1177__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n1732_));
OR2X2 OR2X2_3590 ( .A(u5__abc_81276_new_n2151_), .B(u5__abc_81276_new_n2168_), .Y(u5__abc_81276_new_n2169_));
OR2X2 OR2X2_3591 ( .A(u5__abc_81276_new_n2170_), .B(u5__abc_81276_new_n2173_), .Y(u5__abc_81276_new_n2174_));
OR2X2 OR2X2_3592 ( .A(u5__abc_81276_new_n2178_), .B(u5__abc_81276_new_n2181_), .Y(u5__abc_81276_new_n2182_));
OR2X2 OR2X2_3593 ( .A(u5__abc_81276_new_n2175_), .B(u5__abc_81276_new_n2183_), .Y(u5__abc_81276_new_n2184_));
OR2X2 OR2X2_3594 ( .A(u5__abc_81276_new_n2187_), .B(u5__abc_81276_new_n2190_), .Y(u5__abc_81276_new_n2191_));
OR2X2 OR2X2_3595 ( .A(u5__abc_81276_new_n2195_), .B(u5__abc_81276_new_n2198_), .Y(u5__abc_81276_new_n2199_));
OR2X2 OR2X2_3596 ( .A(u5__abc_81276_new_n2192_), .B(u5__abc_81276_new_n2200_), .Y(u5__abc_81276_new_n2201_));
OR2X2 OR2X2_3597 ( .A(u5__abc_81276_new_n2184_), .B(u5__abc_81276_new_n2201_), .Y(u5__abc_81276_new_n2202_));
OR2X2 OR2X2_3598 ( .A(u5__abc_81276_new_n2202_), .B(u5__abc_81276_new_n2169_), .Y(u5__abc_81276_new_n2203_));
OR2X2 OR2X2_3599 ( .A(u5__abc_81276_new_n949_), .B(u5__abc_81276_new_n993_), .Y(u5__abc_81276_new_n2204_));
OR2X2 OR2X2_36 ( .A(lmr_sel_bF_buf5), .B(tms_0_), .Y(_abc_85006_new_n291_));
OR2X2 OR2X2_360 ( .A(spec_req_cs_6_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1733_));
OR2X2 OR2X2_3600 ( .A(u5__abc_81276_new_n2206_), .B(u5__abc_81276_new_n2211_), .Y(u5__abc_81276_new_n2212_));
OR2X2 OR2X2_3601 ( .A(u5__abc_81276_new_n2213_), .B(u5__abc_81276_new_n2205_), .Y(u5__abc_81276_new_n2214_));
OR2X2 OR2X2_3602 ( .A(u5__abc_81276_new_n2219_), .B(u5__abc_81276_new_n2224_), .Y(u5__abc_81276_new_n2225_));
OR2X2 OR2X2_3603 ( .A(u5__abc_81276_new_n2231_), .B(u5__abc_81276_new_n2236_), .Y(u5__abc_81276_new_n2237_));
OR2X2 OR2X2_3604 ( .A(u5__abc_81276_new_n2226_), .B(u5__abc_81276_new_n2238_), .Y(u5__abc_81276_new_n2239_));
OR2X2 OR2X2_3605 ( .A(u5__abc_81276_new_n2239_), .B(u5__abc_81276_new_n2214_), .Y(u5__abc_81276_new_n2240_));
OR2X2 OR2X2_3606 ( .A(u5__abc_81276_new_n2250_), .B(u5__abc_81276_new_n2244_), .Y(u5__abc_81276_new_n2251_));
OR2X2 OR2X2_3607 ( .A(u5__abc_81276_new_n2257_), .B(u5__abc_81276_new_n2262_), .Y(u5__abc_81276_new_n2263_));
OR2X2 OR2X2_3608 ( .A(u5__abc_81276_new_n2252_), .B(u5__abc_81276_new_n2264_), .Y(u5__abc_81276_new_n2265_));
OR2X2 OR2X2_3609 ( .A(u5__abc_81276_new_n2270_), .B(u5__abc_81276_new_n2275_), .Y(u5__abc_81276_new_n2276_));
OR2X2 OR2X2_361 ( .A(u0__abc_76628_new_n1735_), .B(u0__abc_76628_new_n1731_), .Y(u0__abc_76628_new_n1736_));
OR2X2 OR2X2_3610 ( .A(u5__abc_81276_new_n2283_), .B(u5__abc_81276_new_n2288_), .Y(u5__abc_81276_new_n2289_));
OR2X2 OR2X2_3611 ( .A(u5__abc_81276_new_n2290_), .B(u5__abc_81276_new_n2277_), .Y(u5__abc_81276_new_n2291_));
OR2X2 OR2X2_3612 ( .A(u5__abc_81276_new_n2265_), .B(u5__abc_81276_new_n2291_), .Y(u5__abc_81276_new_n2292_));
OR2X2 OR2X2_3613 ( .A(u5__abc_81276_new_n2292_), .B(u5__abc_81276_new_n2240_), .Y(u5__abc_81276_new_n2293_));
OR2X2 OR2X2_3614 ( .A(u5__abc_81276_new_n2203_), .B(u5__abc_81276_new_n2293_), .Y(u5__abc_81276_new_n2294_));
OR2X2 OR2X2_3615 ( .A(u5__abc_81276_new_n1922_), .B(u5__abc_81276_new_n2300_), .Y(u5__0ap_en_0_0_));
OR2X2 OR2X2_3616 ( .A(u5__abc_81276_new_n2322_), .B(u5__abc_81276_new_n2320_), .Y(u5__abc_81276_new_n2323_));
OR2X2 OR2X2_3617 ( .A(u5__abc_81276_new_n2319_), .B(u5__abc_81276_new_n2330_), .Y(u5__abc_81276_new_n2331_));
OR2X2 OR2X2_3618 ( .A(u5__abc_81276_new_n2333_), .B(u5__abc_81276_new_n2332_), .Y(u5__abc_81276_new_n2334_));
OR2X2 OR2X2_3619 ( .A(u5__abc_81276_new_n2337_), .B(u5__abc_81276_new_n2335_), .Y(u5__abc_81276_new_n2338_));
OR2X2 OR2X2_362 ( .A(u0__abc_76628_new_n1737_), .B(u0__abc_76628_new_n1738_), .Y(u0__abc_76628_new_n1739_));
OR2X2 OR2X2_3620 ( .A(u5__abc_81276_new_n2339_), .B(u5__abc_81276_new_n2331_), .Y(u5__abc_81276_new_n2340_));
OR2X2 OR2X2_3621 ( .A(u5__abc_81276_new_n2344_), .B(u5__abc_81276_new_n1526__bF_buf1), .Y(u5__abc_81276_new_n2345_));
OR2X2 OR2X2_3622 ( .A(u5__abc_81276_new_n2343_), .B(u5__abc_81276_new_n2345_), .Y(u5__abc_81276_new_n2346_));
OR2X2 OR2X2_3623 ( .A(u5__abc_81276_new_n2347_), .B(u5__abc_81276_new_n2323_), .Y(u5__abc_81276_new_n2348_));
OR2X2 OR2X2_3624 ( .A(u5__abc_81276_new_n2353_), .B(u5__abc_81276_new_n2351_), .Y(u5__abc_81276_new_n2354_));
OR2X2 OR2X2_3625 ( .A(u5__abc_81276_new_n2357_), .B(u5__abc_81276_new_n2307_), .Y(u5__abc_81276_new_n2358_));
OR2X2 OR2X2_3626 ( .A(u5__abc_81276_new_n2356_), .B(u5__abc_81276_new_n2358_), .Y(u5__abc_81276_new_n2359_));
OR2X2 OR2X2_3627 ( .A(u5__abc_81276_new_n2355_), .B(u5__abc_81276_new_n2359_), .Y(u5__0burst_cnt_10_0__2_));
OR2X2 OR2X2_3628 ( .A(u5__abc_81276_new_n2363_), .B(u5__abc_81276_new_n1526__bF_buf3), .Y(u5__abc_81276_new_n2364_));
OR2X2 OR2X2_3629 ( .A(u5__abc_81276_new_n2362_), .B(u5__abc_81276_new_n2364_), .Y(u5__abc_81276_new_n2365_));
OR2X2 OR2X2_363 ( .A(u0__abc_76628_new_n1740_), .B(u0__abc_76628_new_n1741_), .Y(u0__abc_76628_new_n1742_));
OR2X2 OR2X2_3630 ( .A(u5__abc_81276_new_n2310_), .B(1'h0), .Y(u5__abc_81276_new_n2366_));
OR2X2 OR2X2_3631 ( .A(u5__abc_81276_new_n2367_), .B(u5__abc_81276_new_n2299_), .Y(u5__abc_81276_new_n2368_));
OR2X2 OR2X2_3632 ( .A(u5__abc_81276_new_n2371_), .B(u5__abc_81276_new_n2299_), .Y(u5__abc_81276_new_n2372_));
OR2X2 OR2X2_3633 ( .A(u5__abc_81276_new_n2374_), .B(u5__abc_81276_new_n2375_), .Y(u5__abc_81276_new_n2376_));
OR2X2 OR2X2_3634 ( .A(u5__abc_81276_new_n2376_), .B(u5__abc_81276_new_n2298_), .Y(u5__abc_81276_new_n2377_));
OR2X2 OR2X2_3635 ( .A(u5__abc_81276_new_n2382_), .B(u5__abc_81276_new_n1526__bF_buf2), .Y(u5__abc_81276_new_n2383_));
OR2X2 OR2X2_3636 ( .A(u5__abc_81276_new_n2383_), .B(u5__abc_81276_new_n2380_), .Y(u5__abc_81276_new_n2384_));
OR2X2 OR2X2_3637 ( .A(u5__abc_81276_new_n2385_), .B(u5__abc_81276_new_n2299_), .Y(u5__abc_81276_new_n2386_));
OR2X2 OR2X2_3638 ( .A(u5__abc_81276_new_n2381_), .B(u5_burst_cnt_5_), .Y(u5__abc_81276_new_n2389_));
OR2X2 OR2X2_3639 ( .A(u5__abc_81276_new_n2391_), .B(u5__abc_81276_new_n1526__bF_buf1), .Y(u5__abc_81276_new_n2392_));
OR2X2 OR2X2_364 ( .A(u0__abc_76628_new_n1743_), .B(u0__abc_76628_new_n1744_), .Y(u0__abc_76628_new_n1745_));
OR2X2 OR2X2_3640 ( .A(u5__abc_81276_new_n2392_), .B(u5__abc_81276_new_n2390_), .Y(u5__abc_81276_new_n2393_));
OR2X2 OR2X2_3641 ( .A(u5__abc_81276_new_n2394_), .B(u5__abc_81276_new_n2299_), .Y(u5__abc_81276_new_n2395_));
OR2X2 OR2X2_3642 ( .A(u5__abc_81276_new_n2399_), .B(u5_burst_cnt_7_), .Y(u5__abc_81276_new_n2400_));
OR2X2 OR2X2_3643 ( .A(u5__abc_81276_new_n2401_), .B(u5__abc_81276_new_n376_), .Y(u5__abc_81276_new_n2402_));
OR2X2 OR2X2_3644 ( .A(u5__abc_81276_new_n2336_), .B(u5__abc_81276_new_n2403_), .Y(u5__abc_81276_new_n2404_));
OR2X2 OR2X2_3645 ( .A(u5__abc_81276_new_n2334_), .B(u5_burst_cnt_7_), .Y(u5__abc_81276_new_n2405_));
OR2X2 OR2X2_3646 ( .A(u5__abc_81276_new_n2406_), .B(u5__abc_81276_new_n2298_), .Y(u5__abc_81276_new_n2407_));
OR2X2 OR2X2_3647 ( .A(u5__abc_81276_new_n2408_), .B(u5__abc_81276_new_n2299_), .Y(u5__abc_81276_new_n2409_));
OR2X2 OR2X2_3648 ( .A(u5__abc_81276_new_n2416_), .B(u5__abc_81276_new_n1526__bF_buf0), .Y(u5__abc_81276_new_n2417_));
OR2X2 OR2X2_3649 ( .A(u5__abc_81276_new_n2417_), .B(u5__abc_81276_new_n2414_), .Y(u5__abc_81276_new_n2418_));
OR2X2 OR2X2_365 ( .A(u0__abc_76628_new_n1747_), .B(spec_req_cs_0_bF_buf3_), .Y(u0__abc_76628_new_n1748_));
OR2X2 OR2X2_3650 ( .A(u5__abc_81276_new_n2419_), .B(u5__abc_81276_new_n2299_), .Y(u5__abc_81276_new_n2420_));
OR2X2 OR2X2_3651 ( .A(u5__abc_81276_new_n2425_), .B(u5__abc_81276_new_n1526__bF_buf3), .Y(u5__abc_81276_new_n2426_));
OR2X2 OR2X2_3652 ( .A(u5__abc_81276_new_n2424_), .B(u5__abc_81276_new_n2426_), .Y(u5__abc_81276_new_n2427_));
OR2X2 OR2X2_3653 ( .A(u5__abc_81276_new_n2428_), .B(u5__abc_81276_new_n2299_), .Y(u5__abc_81276_new_n2429_));
OR2X2 OR2X2_3654 ( .A(u5__abc_81276_new_n2433_), .B(u5_burst_cnt_10_), .Y(u5__abc_81276_new_n2434_));
OR2X2 OR2X2_3655 ( .A(u5__abc_81276_new_n2435_), .B(u5__abc_81276_new_n380_), .Y(u5__abc_81276_new_n2436_));
OR2X2 OR2X2_3656 ( .A(u5__abc_81276_new_n2336_), .B(u5__abc_81276_new_n2437_), .Y(u5__abc_81276_new_n2438_));
OR2X2 OR2X2_3657 ( .A(u5__abc_81276_new_n2334_), .B(u5_burst_cnt_10_), .Y(u5__abc_81276_new_n2439_));
OR2X2 OR2X2_3658 ( .A(u5__abc_81276_new_n2440_), .B(u5__abc_81276_new_n1526__bF_buf2), .Y(u5__abc_81276_new_n2441_));
OR2X2 OR2X2_3659 ( .A(u5__abc_81276_new_n2442_), .B(u5__abc_81276_new_n2299_), .Y(u5__abc_81276_new_n2443_));
OR2X2 OR2X2_366 ( .A(u0__abc_76628_new_n1746_), .B(u0__abc_76628_new_n1748_), .Y(u0__abc_76628_new_n1749_));
OR2X2 OR2X2_3660 ( .A(u5__abc_81276_new_n2465_), .B(u5__abc_81276_new_n2463_), .Y(u5__abc_81276_new_n2466_));
OR2X2 OR2X2_3661 ( .A(u5__abc_81276_new_n2463_), .B(u5__abc_81276_new_n1116_), .Y(u5__abc_81276_new_n2477_));
OR2X2 OR2X2_3662 ( .A(u5__abc_81276_new_n2481_), .B(u5__abc_81276_new_n2482_), .Y(u5__abc_81276_new_n2483_));
OR2X2 OR2X2_3663 ( .A(u5__abc_81276_new_n2482_), .B(u5_ir_cnt_3_), .Y(u5__abc_81276_new_n2487_));
OR2X2 OR2X2_3664 ( .A(u5__abc_81276_new_n2500_), .B(u5__abc_81276_new_n1648_), .Y(u5__abc_81276_new_n2501_));
OR2X2 OR2X2_3665 ( .A(u5__abc_81276_new_n1682__bF_buf1), .B(tms_s_4_), .Y(u5__abc_81276_new_n2509_));
OR2X2 OR2X2_3666 ( .A(u5__abc_81276_new_n2509_), .B(u5__abc_81276_new_n2516_), .Y(u5__abc_81276_new_n2517_));
OR2X2 OR2X2_3667 ( .A(u5__abc_81276_new_n1682__bF_buf0), .B(tms_s_24_), .Y(u5__abc_81276_new_n2518_));
OR2X2 OR2X2_3668 ( .A(u5__abc_81276_new_n2518_), .B(u5__abc_81276_new_n2528_), .Y(u5__abc_81276_new_n2529_));
OR2X2 OR2X2_3669 ( .A(u5_timer_is_zero), .B(u5_mc_le), .Y(u5__abc_81276_new_n2539_));
OR2X2 OR2X2_367 ( .A(u0__abc_76628_new_n1197__bF_buf0), .B(u0_tms0_23_), .Y(u0__abc_76628_new_n1750_));
OR2X2 OR2X2_3670 ( .A(u5__abc_81276_new_n2541_), .B(u5__abc_81276_new_n2542_), .Y(u5__abc_81276_new_n2543_));
OR2X2 OR2X2_3671 ( .A(u5__abc_81276_new_n2538_), .B(u5__abc_81276_new_n2543_), .Y(u5__abc_81276_new_n2544_));
OR2X2 OR2X2_3672 ( .A(u5__abc_81276_new_n2551_), .B(u5__abc_81276_new_n2544_), .Y(u5__abc_81276_new_n2552_));
OR2X2 OR2X2_3673 ( .A(u5__abc_81276_new_n2553_), .B(u5__abc_81276_new_n2515_), .Y(u5__abc_81276_new_n2554_));
OR2X2 OR2X2_3674 ( .A(u5__abc_81276_new_n2555_), .B(u5__abc_81276_new_n2508_), .Y(u5__abc_81276_new_n2556_));
OR2X2 OR2X2_3675 ( .A(u5__abc_81276_new_n1682__bF_buf4), .B(tms_s_17_), .Y(u5__abc_81276_new_n2557_));
OR2X2 OR2X2_3676 ( .A(u5__abc_81276_new_n2557_), .B(u5__abc_81276_new_n2558_), .Y(u5__abc_81276_new_n2559_));
OR2X2 OR2X2_3677 ( .A(u5__abc_81276_new_n2560_), .B(u5__abc_81276_new_n2501_), .Y(u5__abc_81276_new_n2561_));
OR2X2 OR2X2_3678 ( .A(u5__abc_81276_new_n1682__bF_buf3), .B(tms_s_20_), .Y(u5__abc_81276_new_n2562_));
OR2X2 OR2X2_3679 ( .A(u5__abc_81276_new_n2562_), .B(u5__abc_81276_new_n2563_), .Y(u5__abc_81276_new_n2564_));
OR2X2 OR2X2_368 ( .A(u0__abc_76628_new_n1752_), .B(u0__abc_76628_new_n1730_), .Y(u0__0sp_tms_31_0__23_));
OR2X2 OR2X2_3680 ( .A(u5__abc_81276_new_n2562_), .B(tms_s_15_), .Y(u5__abc_81276_new_n2573_));
OR2X2 OR2X2_3681 ( .A(u5__abc_81276_new_n1682__bF_buf2), .B(tms_s_15_), .Y(u5__abc_81276_new_n2574_));
OR2X2 OR2X2_3682 ( .A(u5__abc_81276_new_n1561_), .B(u5__abc_81276_new_n2581_), .Y(u5__abc_81276_new_n2582_));
OR2X2 OR2X2_3683 ( .A(u5__abc_81276_new_n2582_), .B(u5__abc_81276_new_n2579_), .Y(u5__abc_81276_new_n2583_));
OR2X2 OR2X2_3684 ( .A(u5__abc_81276_new_n2578_), .B(u5__abc_81276_new_n2609_), .Y(u5__abc_81276_new_n2610_));
OR2X2 OR2X2_3685 ( .A(u5__abc_81276_new_n2572_), .B(u5__abc_81276_new_n2610_), .Y(u5__abc_81276_new_n2611_));
OR2X2 OR2X2_3686 ( .A(u5__abc_81276_new_n2638_), .B(u5__abc_81276_new_n2612_), .Y(u5__abc_81276_new_n2639_));
OR2X2 OR2X2_3687 ( .A(u5__abc_81276_new_n2313_), .B(u5__abc_81276_new_n2654_), .Y(u5__abc_81276_new_n2655_));
OR2X2 OR2X2_3688 ( .A(u5__abc_81276_new_n2582_), .B(u5__abc_81276_new_n2658_), .Y(u5__abc_81276_new_n2659_));
OR2X2 OR2X2_3689 ( .A(u5__abc_81276_new_n1682__bF_buf1), .B(tms_s_8_), .Y(u5__abc_81276_new_n2669_));
OR2X2 OR2X2_369 ( .A(u0__abc_76628_new_n1177__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n1756_));
OR2X2 OR2X2_3690 ( .A(u5__abc_81276_new_n2670_), .B(u5__abc_81276_new_n2668_), .Y(u5__abc_81276_new_n2671_));
OR2X2 OR2X2_3691 ( .A(u5__abc_81276_new_n2657_), .B(u5__abc_81276_new_n2671_), .Y(u5__abc_81276_new_n2672_));
OR2X2 OR2X2_3692 ( .A(u5__abc_81276_new_n1682__bF_buf0), .B(tms_s_12_), .Y(u5__abc_81276_new_n2674_));
OR2X2 OR2X2_3693 ( .A(u5__abc_81276_new_n2674_), .B(u5__abc_81276_new_n2673_), .Y(u5__abc_81276_new_n2675_));
OR2X2 OR2X2_3694 ( .A(u5__abc_81276_new_n1682__bF_buf4), .B(tms_s_13_), .Y(u5__abc_81276_new_n2677_));
OR2X2 OR2X2_3695 ( .A(u5__abc_81276_new_n2677_), .B(u5__abc_81276_new_n2673_), .Y(u5__abc_81276_new_n2678_));
OR2X2 OR2X2_3696 ( .A(u5__abc_81276_new_n1682__bF_buf3), .B(tms_s_18_), .Y(u5__abc_81276_new_n2679_));
OR2X2 OR2X2_3697 ( .A(u5__abc_81276_new_n2679_), .B(u5__abc_81276_new_n2558_), .Y(u5__abc_81276_new_n2680_));
OR2X2 OR2X2_3698 ( .A(u5__abc_81276_new_n1682__bF_buf2), .B(tms_s_5_), .Y(u5__abc_81276_new_n2681_));
OR2X2 OR2X2_3699 ( .A(u5__abc_81276_new_n2681_), .B(u5__abc_81276_new_n2516_), .Y(u5__abc_81276_new_n2682_));
OR2X2 OR2X2_37 ( .A(_abc_85006_new_n240__bF_buf2), .B(sp_tms_1_), .Y(_abc_85006_new_n293_));
OR2X2 OR2X2_370 ( .A(spec_req_cs_6_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n1757_));
OR2X2 OR2X2_3700 ( .A(u5__abc_81276_new_n1682__bF_buf1), .B(tms_s_25_), .Y(u5__abc_81276_new_n2683_));
OR2X2 OR2X2_3701 ( .A(u5__abc_81276_new_n2683_), .B(u5__abc_81276_new_n2528_), .Y(u5__abc_81276_new_n2684_));
OR2X2 OR2X2_3702 ( .A(u5__abc_81276_new_n2686_), .B(u5__abc_81276_new_n2687_), .Y(u5__abc_81276_new_n2688_));
OR2X2 OR2X2_3703 ( .A(u5__abc_81276_new_n2691_), .B(u5__abc_81276_new_n2688_), .Y(u5__abc_81276_new_n2692_));
OR2X2 OR2X2_3704 ( .A(u5__abc_81276_new_n2693_), .B(u5__abc_81276_new_n2515_), .Y(u5__abc_81276_new_n2694_));
OR2X2 OR2X2_3705 ( .A(u5__abc_81276_new_n2695_), .B(u5__abc_81276_new_n2508_), .Y(u5__abc_81276_new_n2696_));
OR2X2 OR2X2_3706 ( .A(u5__abc_81276_new_n2697_), .B(u5__abc_81276_new_n2501_), .Y(u5__abc_81276_new_n2698_));
OR2X2 OR2X2_3707 ( .A(u5__abc_81276_new_n1682__bF_buf0), .B(tms_s_21_), .Y(u5__abc_81276_new_n2699_));
OR2X2 OR2X2_3708 ( .A(u5__abc_81276_new_n2699_), .B(u5__abc_81276_new_n2563_), .Y(u5__abc_81276_new_n2700_));
OR2X2 OR2X2_3709 ( .A(u5__abc_81276_new_n1682__bF_buf4), .B(tms_s_16_), .Y(u5__abc_81276_new_n2703_));
OR2X2 OR2X2_371 ( .A(u0__abc_76628_new_n1759_), .B(u0__abc_76628_new_n1755_), .Y(u0__abc_76628_new_n1760_));
OR2X2 OR2X2_3710 ( .A(u5__abc_81276_new_n2699_), .B(tms_s_16_), .Y(u5__abc_81276_new_n2706_));
OR2X2 OR2X2_3711 ( .A(u5__abc_81276_new_n2707_), .B(u5__abc_81276_new_n2575_), .Y(u5__abc_81276_new_n2708_));
OR2X2 OR2X2_3712 ( .A(u5__abc_81276_new_n2709_), .B(u5__abc_81276_new_n2704_), .Y(u5__abc_81276_new_n2710_));
OR2X2 OR2X2_3713 ( .A(u5__abc_81276_new_n2710_), .B(u5__abc_81276_new_n2576_), .Y(u5__abc_81276_new_n2711_));
OR2X2 OR2X2_3714 ( .A(u5__abc_81276_new_n2713_), .B(u5__abc_81276_new_n2609_), .Y(u5__abc_81276_new_n2714_));
OR2X2 OR2X2_3715 ( .A(u5__abc_81276_new_n2702_), .B(u5__abc_81276_new_n2714_), .Y(u5__abc_81276_new_n2715_));
OR2X2 OR2X2_3716 ( .A(u5__abc_81276_new_n2315_), .B(u5__abc_81276_new_n2654_), .Y(u5__abc_81276_new_n2716_));
OR2X2 OR2X2_3717 ( .A(u5__abc_81276_new_n1682__bF_buf3), .B(tms_s_9_), .Y(u5__abc_81276_new_n2719_));
OR2X2 OR2X2_3718 ( .A(u5__abc_81276_new_n2720_), .B(u5__abc_81276_new_n2668_), .Y(u5__abc_81276_new_n2721_));
OR2X2 OR2X2_3719 ( .A(u5__abc_81276_new_n2718_), .B(u5__abc_81276_new_n2721_), .Y(u5__abc_81276_new_n2722_));
OR2X2 OR2X2_372 ( .A(u0__abc_76628_new_n1761_), .B(u0__abc_76628_new_n1762_), .Y(u0__abc_76628_new_n1763_));
OR2X2 OR2X2_3720 ( .A(u5__abc_81276_new_n2311_), .B(u5__abc_81276_new_n2654_), .Y(u5__abc_81276_new_n2724_));
OR2X2 OR2X2_3721 ( .A(u5__abc_81276_new_n1682__bF_buf2), .B(tms_s_22_), .Y(u5__abc_81276_new_n2725_));
OR2X2 OR2X2_3722 ( .A(u5__abc_81276_new_n2726_), .B(u5__abc_81276_new_n2704_), .Y(u5__abc_81276_new_n2727_));
OR2X2 OR2X2_3723 ( .A(u5__abc_81276_new_n2727_), .B(u5__abc_81276_new_n2725_), .Y(u5__abc_81276_new_n2728_));
OR2X2 OR2X2_3724 ( .A(u5__abc_81276_new_n2730_), .B(u5__abc_81276_new_n2729_), .Y(u5__abc_81276_new_n2731_));
OR2X2 OR2X2_3725 ( .A(u5__abc_81276_new_n2734_), .B(u5__abc_81276_new_n2501_), .Y(u5__abc_81276_new_n2735_));
OR2X2 OR2X2_3726 ( .A(u5__abc_81276_new_n2743_), .B(u5__abc_81276_new_n1955_), .Y(u5__abc_81276_new_n2744_));
OR2X2 OR2X2_3727 ( .A(u5__abc_81276_new_n1941_), .B(u5__abc_81276_new_n2746_), .Y(u5__abc_81276_new_n2747_));
OR2X2 OR2X2_3728 ( .A(u5__abc_81276_new_n2767_), .B(u5__abc_81276_new_n2768_), .Y(u5__abc_81276_new_n2769_));
OR2X2 OR2X2_3729 ( .A(u5__abc_81276_new_n1682__bF_buf1), .B(tms_s_26_), .Y(u5__abc_81276_new_n2781_));
OR2X2 OR2X2_373 ( .A(u0__abc_76628_new_n1764_), .B(u0__abc_76628_new_n1765_), .Y(u0__abc_76628_new_n1766_));
OR2X2 OR2X2_3730 ( .A(u5__abc_81276_new_n2784_), .B(u5__abc_81276_new_n2785_), .Y(u5__abc_81276_new_n2786_));
OR2X2 OR2X2_3731 ( .A(u5__abc_81276_new_n2538_), .B(u5__abc_81276_new_n2786_), .Y(u5__abc_81276_new_n2787_));
OR2X2 OR2X2_3732 ( .A(u5__abc_81276_new_n2782_), .B(u5__abc_81276_new_n2788_), .Y(u5__abc_81276_new_n2789_));
OR2X2 OR2X2_3733 ( .A(u5__abc_81276_new_n2791_), .B(u5__abc_81276_new_n2735_), .Y(u5__abc_81276_new_n2792_));
OR2X2 OR2X2_3734 ( .A(u5__abc_81276_new_n2725_), .B(u5__abc_81276_new_n2563_), .Y(u5__abc_81276_new_n2793_));
OR2X2 OR2X2_3735 ( .A(u5__abc_81276_new_n2795_), .B(u5__abc_81276_new_n2609_), .Y(u5__abc_81276_new_n2796_));
OR2X2 OR2X2_3736 ( .A(u5__abc_81276_new_n2733_), .B(u5__abc_81276_new_n2796_), .Y(u5__abc_81276_new_n2797_));
OR2X2 OR2X2_3737 ( .A(u5__abc_81276_new_n1682__bF_buf0), .B(tms_s_10_), .Y(u5__abc_81276_new_n2800_));
OR2X2 OR2X2_3738 ( .A(u5__abc_81276_new_n2801_), .B(u5__abc_81276_new_n2668_), .Y(u5__abc_81276_new_n2802_));
OR2X2 OR2X2_3739 ( .A(u5__abc_81276_new_n2799_), .B(u5__abc_81276_new_n2802_), .Y(u5__abc_81276_new_n2803_));
OR2X2 OR2X2_374 ( .A(u0__abc_76628_new_n1767_), .B(u0__abc_76628_new_n1768_), .Y(u0__abc_76628_new_n1769_));
OR2X2 OR2X2_3740 ( .A(u5__abc_81276_new_n1682__bF_buf4), .B(tms_s_14_), .Y(u5__abc_81276_new_n2804_));
OR2X2 OR2X2_3741 ( .A(u5__abc_81276_new_n2804_), .B(u5__abc_81276_new_n2673_), .Y(u5__abc_81276_new_n2805_));
OR2X2 OR2X2_3742 ( .A(u5__abc_81276_new_n2574_), .B(u5__abc_81276_new_n2673_), .Y(u5__abc_81276_new_n2807_));
OR2X2 OR2X2_3743 ( .A(u5__abc_81276_new_n1682__bF_buf3), .B(tms_s_23_), .Y(u5__abc_81276_new_n2808_));
OR2X2 OR2X2_3744 ( .A(u5__abc_81276_new_n2731_), .B(u5__abc_81276_new_n2809_), .Y(u5__abc_81276_new_n2810_));
OR2X2 OR2X2_3745 ( .A(u5__abc_81276_new_n2811_), .B(u5__abc_81276_new_n2808_), .Y(u5__abc_81276_new_n2812_));
OR2X2 OR2X2_3746 ( .A(u5__abc_81276_new_n1682__bF_buf2), .B(tms_s_27_), .Y(u5__abc_81276_new_n2816_));
OR2X2 OR2X2_3747 ( .A(u5__abc_81276_new_n2820_), .B(u5__abc_81276_new_n2818_), .Y(u5__abc_81276_new_n2821_));
OR2X2 OR2X2_3748 ( .A(u5__abc_81276_new_n2817_), .B(u5__abc_81276_new_n2822_), .Y(u5__abc_81276_new_n2823_));
OR2X2 OR2X2_3749 ( .A(u5__abc_81276_new_n2849_), .B(u5__abc_81276_new_n2815_), .Y(u5__abc_81276_new_n2850_));
OR2X2 OR2X2_375 ( .A(u0__abc_76628_new_n1771_), .B(spec_req_cs_0_bF_buf2_), .Y(u0__abc_76628_new_n1772_));
OR2X2 OR2X2_3750 ( .A(u5__abc_81276_new_n2851_), .B(u5__abc_81276_new_n2609_), .Y(u5__abc_81276_new_n2852_));
OR2X2 OR2X2_3751 ( .A(u5__abc_81276_new_n2814_), .B(u5__abc_81276_new_n2852_), .Y(u5__abc_81276_new_n2853_));
OR2X2 OR2X2_3752 ( .A(u5__abc_81276_new_n1682__bF_buf1), .B(tms_s_3_), .Y(u5__abc_81276_new_n2854_));
OR2X2 OR2X2_3753 ( .A(u5__abc_81276_new_n2854_), .B(u5__abc_81276_new_n2654_), .Y(u5__abc_81276_new_n2855_));
OR2X2 OR2X2_3754 ( .A(u5__abc_81276_new_n1682__bF_buf0), .B(tms_s_11_), .Y(u5__abc_81276_new_n2858_));
OR2X2 OR2X2_3755 ( .A(u5__abc_81276_new_n2859_), .B(u5__abc_81276_new_n2668_), .Y(u5__abc_81276_new_n2860_));
OR2X2 OR2X2_3756 ( .A(u5__abc_81276_new_n2857_), .B(u5__abc_81276_new_n2860_), .Y(u5__abc_81276_new_n2861_));
OR2X2 OR2X2_3757 ( .A(u5__abc_81276_new_n2875_), .B(u5__abc_81276_new_n2873_), .Y(u5__abc_81276_new_n2876_));
OR2X2 OR2X2_3758 ( .A(u5__abc_81276_new_n2879_), .B(u5__abc_81276_new_n2880_), .Y(u5__abc_81276_new_n2881_));
OR2X2 OR2X2_3759 ( .A(u5__abc_81276_new_n2885_), .B(u5__abc_81276_new_n2883_), .Y(u5__abc_81276_new_n2886_));
OR2X2 OR2X2_376 ( .A(u0__abc_76628_new_n1770_), .B(u0__abc_76628_new_n1772_), .Y(u0__abc_76628_new_n1773_));
OR2X2 OR2X2_3760 ( .A(u5__abc_81276_new_n2888_), .B(u5__abc_81276_new_n2653_), .Y(u5__abc_81276_new_n2889_));
OR2X2 OR2X2_3761 ( .A(u5__abc_81276_new_n2681_), .B(u5__abc_81276_new_n2654_), .Y(u5__abc_81276_new_n2890_));
OR2X2 OR2X2_3762 ( .A(u5__abc_81276_new_n2894_), .B(u5__abc_81276_new_n2896_), .Y(u5__abc_81276_new_n2897_));
OR2X2 OR2X2_3763 ( .A(u5__abc_81276_new_n2898_), .B(u5__abc_81276_new_n2653_), .Y(u5__abc_81276_new_n2899_));
OR2X2 OR2X2_3764 ( .A(u5__abc_81276_new_n1682__bF_buf4), .B(tms_s_6_), .Y(u5__abc_81276_new_n2900_));
OR2X2 OR2X2_3765 ( .A(u5__abc_81276_new_n2900_), .B(u5__abc_81276_new_n2654_), .Y(u5__abc_81276_new_n2901_));
OR2X2 OR2X2_3766 ( .A(u5__abc_81276_new_n2906_), .B(u5__abc_81276_new_n2653_), .Y(u5__abc_81276_new_n2907_));
OR2X2 OR2X2_3767 ( .A(u5__abc_81276_new_n1682__bF_buf3), .B(tms_s_7_), .Y(u5__abc_81276_new_n2908_));
OR2X2 OR2X2_3768 ( .A(u5__abc_81276_new_n2908_), .B(u5__abc_81276_new_n2654_), .Y(u5__abc_81276_new_n2909_));
OR2X2 OR2X2_3769 ( .A(u5__abc_81276_new_n2562_), .B(u5__abc_81276_new_n2920_), .Y(u5__abc_81276_new_n2921_));
OR2X2 OR2X2_377 ( .A(u0__abc_76628_new_n1197__bF_buf5), .B(u0_tms0_24_), .Y(u0__abc_76628_new_n1774_));
OR2X2 OR2X2_3770 ( .A(u5_timer2_1_), .B(u5_timer2_0_), .Y(u5__abc_81276_new_n2935_));
OR2X2 OR2X2_3771 ( .A(u5__abc_81276_new_n2935_), .B(u5_timer2_2_), .Y(u5__abc_81276_new_n2936_));
OR2X2 OR2X2_3772 ( .A(u5__abc_81276_new_n2936_), .B(u5_timer2_3_), .Y(u5__abc_81276_new_n2937_));
OR2X2 OR2X2_3773 ( .A(u5__abc_81276_new_n2937_), .B(u5_timer2_4_), .Y(u5__abc_81276_new_n2938_));
OR2X2 OR2X2_3774 ( .A(u5__abc_81276_new_n2938_), .B(u5_timer2_5_), .Y(u5__abc_81276_new_n2939_));
OR2X2 OR2X2_3775 ( .A(u5__abc_81276_new_n2939_), .B(u5_timer2_6_), .Y(u5__abc_81276_new_n2940_));
OR2X2 OR2X2_3776 ( .A(u5__abc_81276_new_n2940_), .B(u5_timer2_7_), .Y(u5__abc_81276_new_n2941_));
OR2X2 OR2X2_3777 ( .A(u5__abc_81276_new_n2941_), .B(u5_timer2_8_), .Y(u5__abc_81276_new_n2942_));
OR2X2 OR2X2_3778 ( .A(u5__abc_81276_new_n2948_), .B(u5__abc_81276_new_n2943_), .Y(u5__abc_81276_new_n2949_));
OR2X2 OR2X2_3779 ( .A(u5__abc_81276_new_n2933_), .B(u5__abc_81276_new_n2949_), .Y(u5__abc_81276_new_n2950_));
OR2X2 OR2X2_378 ( .A(u0__abc_76628_new_n1776_), .B(u0__abc_76628_new_n1754_), .Y(u0__0sp_tms_31_0__24_));
OR2X2 OR2X2_3780 ( .A(u5__abc_81276_new_n2960_), .B(u5__abc_81276_new_n2954_), .Y(u5__abc_81276_new_n2961_));
OR2X2 OR2X2_3781 ( .A(u5__abc_81276_new_n2952_), .B(u5__abc_81276_new_n2961_), .Y(u5__abc_81276_new_n2962_));
OR2X2 OR2X2_3782 ( .A(u5__abc_81276_new_n2967_), .B(u5__abc_81276_new_n2912_), .Y(u5__abc_81276_new_n2968_));
OR2X2 OR2X2_3783 ( .A(u5__abc_81276_new_n2674_), .B(u5__abc_81276_new_n2970_), .Y(u5__abc_81276_new_n2971_));
OR2X2 OR2X2_3784 ( .A(u5__abc_81276_new_n2973_), .B(u5__abc_81276_new_n2913_), .Y(u5__0timer2_8_0__0_));
OR2X2 OR2X2_3785 ( .A(u5__abc_81276_new_n782_), .B(u5__abc_81276_new_n761_), .Y(u5__abc_81276_new_n2996_));
OR2X2 OR2X2_3786 ( .A(u5__abc_81276_new_n3011_), .B(u5__abc_81276_new_n3012_), .Y(u5__abc_81276_new_n3013_));
OR2X2 OR2X2_3787 ( .A(u5__abc_81276_new_n3015_), .B(u5__abc_81276_new_n2992_), .Y(u5__abc_81276_new_n3016_));
OR2X2 OR2X2_3788 ( .A(u5__abc_81276_new_n2987_), .B(u5__abc_81276_new_n3016_), .Y(u5__abc_81276_new_n3017_));
OR2X2 OR2X2_3789 ( .A(u5__abc_81276_new_n2669_), .B(u5__abc_81276_new_n3018_), .Y(u5__abc_81276_new_n3019_));
OR2X2 OR2X2_379 ( .A(u0__abc_76628_new_n1177__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n1780_));
OR2X2 OR2X2_3790 ( .A(u5__abc_81276_new_n3020_), .B(u5__abc_81276_new_n2986_), .Y(u5__abc_81276_new_n3021_));
OR2X2 OR2X2_3791 ( .A(u5__abc_81276_new_n2699_), .B(u5__abc_81276_new_n3022_), .Y(u5__abc_81276_new_n3023_));
OR2X2 OR2X2_3792 ( .A(u5__abc_81276_new_n3026_), .B(u5__abc_81276_new_n2961_), .Y(u5__abc_81276_new_n3027_));
OR2X2 OR2X2_3793 ( .A(u5__abc_81276_new_n3025_), .B(u5__abc_81276_new_n3027_), .Y(u5__abc_81276_new_n3028_));
OR2X2 OR2X2_3794 ( .A(u5__abc_81276_new_n3030_), .B(u5__abc_81276_new_n3029_), .Y(u5__abc_81276_new_n3031_));
OR2X2 OR2X2_3795 ( .A(u5__abc_81276_new_n3032_), .B(u5__abc_81276_new_n2975_), .Y(u5__0timer2_8_0__1_));
OR2X2 OR2X2_3796 ( .A(u5__abc_81276_new_n2679_), .B(u5__abc_81276_new_n3034_), .Y(u5__abc_81276_new_n3035_));
OR2X2 OR2X2_3797 ( .A(u5__abc_81276_new_n2725_), .B(u5__abc_81276_new_n2920_), .Y(u5__abc_81276_new_n3036_));
OR2X2 OR2X2_3798 ( .A(u5__abc_81276_new_n2719_), .B(u5__abc_81276_new_n2931_), .Y(u5__abc_81276_new_n3037_));
OR2X2 OR2X2_3799 ( .A(u5__abc_81276_new_n3039_), .B(u5__abc_81276_new_n3040_), .Y(u5__abc_81276_new_n3041_));
OR2X2 OR2X2_38 ( .A(lmr_sel_bF_buf4), .B(tms_1_), .Y(_abc_85006_new_n294_));
OR2X2 OR2X2_380 ( .A(spec_req_cs_6_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n1781_));
OR2X2 OR2X2_3800 ( .A(u5__abc_81276_new_n3043_), .B(u5__abc_81276_new_n2992_), .Y(u5__abc_81276_new_n3044_));
OR2X2 OR2X2_3801 ( .A(u5__abc_81276_new_n3038_), .B(u5__abc_81276_new_n3044_), .Y(u5__abc_81276_new_n3045_));
OR2X2 OR2X2_3802 ( .A(u5__abc_81276_new_n3046_), .B(u5__abc_81276_new_n2919_), .Y(u5__abc_81276_new_n3047_));
OR2X2 OR2X2_3803 ( .A(u5__abc_81276_new_n3048_), .B(u5__abc_81276_new_n2925_), .Y(u5__abc_81276_new_n3049_));
OR2X2 OR2X2_3804 ( .A(u5__abc_81276_new_n2557_), .B(u5__abc_81276_new_n2926_), .Y(u5__abc_81276_new_n3050_));
OR2X2 OR2X2_3805 ( .A(u5__abc_81276_new_n2804_), .B(u5__abc_81276_new_n2968_), .Y(u5__abc_81276_new_n3054_));
OR2X2 OR2X2_3806 ( .A(u5__abc_81276_new_n3052_), .B(u5__abc_81276_new_n3055_), .Y(u5__abc_81276_new_n3056_));
OR2X2 OR2X2_3807 ( .A(u5__abc_81276_new_n3059_), .B(u5__abc_81276_new_n3029_), .Y(u5__abc_81276_new_n3060_));
OR2X2 OR2X2_3808 ( .A(u5__abc_81276_new_n3062_), .B(u5__abc_81276_new_n3063_), .Y(u5__abc_81276_new_n3064_));
OR2X2 OR2X2_3809 ( .A(u5__abc_81276_new_n3066_), .B(u5__abc_81276_new_n2992_), .Y(u5__abc_81276_new_n3067_));
OR2X2 OR2X2_381 ( .A(u0__abc_76628_new_n1783_), .B(u0__abc_76628_new_n1779_), .Y(u0__abc_76628_new_n1784_));
OR2X2 OR2X2_3810 ( .A(u5__abc_81276_new_n3061_), .B(u5__abc_81276_new_n3067_), .Y(u5__abc_81276_new_n3068_));
OR2X2 OR2X2_3811 ( .A(u5__abc_81276_new_n2800_), .B(u5__abc_81276_new_n3018_), .Y(u5__abc_81276_new_n3069_));
OR2X2 OR2X2_3812 ( .A(u5__abc_81276_new_n3070_), .B(u5__abc_81276_new_n2986_), .Y(u5__abc_81276_new_n3071_));
OR2X2 OR2X2_3813 ( .A(u5__abc_81276_new_n2808_), .B(u5__abc_81276_new_n3022_), .Y(u5__abc_81276_new_n3072_));
OR2X2 OR2X2_3814 ( .A(u5__abc_81276_new_n3075_), .B(u5__abc_81276_new_n2961_), .Y(u5__abc_81276_new_n3076_));
OR2X2 OR2X2_3815 ( .A(u5__abc_81276_new_n3074_), .B(u5__abc_81276_new_n3076_), .Y(u5__abc_81276_new_n3077_));
OR2X2 OR2X2_3816 ( .A(u5__abc_81276_new_n3078_), .B(u5__abc_81276_new_n3058_), .Y(u5__0timer2_8_0__3_));
OR2X2 OR2X2_3817 ( .A(u5__abc_81276_new_n3082_), .B(u5__abc_81276_new_n3083_), .Y(u5__abc_81276_new_n3084_));
OR2X2 OR2X2_3818 ( .A(u5__abc_81276_new_n3086_), .B(u5__abc_81276_new_n2992_), .Y(u5__abc_81276_new_n3087_));
OR2X2 OR2X2_3819 ( .A(u5__abc_81276_new_n3081_), .B(u5__abc_81276_new_n3087_), .Y(u5__abc_81276_new_n3088_));
OR2X2 OR2X2_382 ( .A(u0__abc_76628_new_n1785_), .B(u0__abc_76628_new_n1786_), .Y(u0__abc_76628_new_n1787_));
OR2X2 OR2X2_3820 ( .A(u5__abc_81276_new_n2858_), .B(u5__abc_81276_new_n3018_), .Y(u5__abc_81276_new_n3089_));
OR2X2 OR2X2_3821 ( .A(u5__abc_81276_new_n3090_), .B(u5__abc_81276_new_n2986_), .Y(u5__abc_81276_new_n3091_));
OR2X2 OR2X2_3822 ( .A(u5__abc_81276_new_n2518_), .B(u5__abc_81276_new_n3022_), .Y(u5__abc_81276_new_n3092_));
OR2X2 OR2X2_3823 ( .A(u5__abc_81276_new_n3094_), .B(u5__abc_81276_new_n3095_), .Y(u5__abc_81276_new_n3096_));
OR2X2 OR2X2_3824 ( .A(u5__abc_81276_new_n3097_), .B(u5__abc_81276_new_n3080_), .Y(u5__0timer2_8_0__4_));
OR2X2 OR2X2_3825 ( .A(u5__abc_81276_new_n2509_), .B(u5__abc_81276_new_n3100_), .Y(u5__abc_81276_new_n3101_));
OR2X2 OR2X2_3826 ( .A(u5__abc_81276_new_n3102_), .B(u5__abc_81276_new_n3103_), .Y(u5__abc_81276_new_n3104_));
OR2X2 OR2X2_3827 ( .A(u5__abc_81276_new_n2948_), .B(u5__abc_81276_new_n3105_), .Y(u5__abc_81276_new_n3106_));
OR2X2 OR2X2_3828 ( .A(u5__abc_81276_new_n3108_), .B(u5__abc_81276_new_n2919_), .Y(u5__abc_81276_new_n3109_));
OR2X2 OR2X2_3829 ( .A(u5__abc_81276_new_n2683_), .B(u5__abc_81276_new_n2920_), .Y(u5__abc_81276_new_n3110_));
OR2X2 OR2X2_383 ( .A(u0__abc_76628_new_n1788_), .B(u0__abc_76628_new_n1789_), .Y(u0__abc_76628_new_n1790_));
OR2X2 OR2X2_3830 ( .A(u5__abc_81276_new_n3113_), .B(u5__abc_81276_new_n3099_), .Y(u5__0timer2_8_0__5_));
OR2X2 OR2X2_3831 ( .A(u5__abc_81276_new_n3117_), .B(u5__abc_81276_new_n3118_), .Y(u5__abc_81276_new_n3119_));
OR2X2 OR2X2_3832 ( .A(u5__abc_81276_new_n3116_), .B(u5__abc_81276_new_n3121_), .Y(u5__abc_81276_new_n3122_));
OR2X2 OR2X2_3833 ( .A(u5__abc_81276_new_n3124_), .B(u5__abc_81276_new_n3115_), .Y(u5__0timer2_8_0__6_));
OR2X2 OR2X2_3834 ( .A(u5__abc_81276_new_n3129_), .B(u5__abc_81276_new_n3130_), .Y(u5__abc_81276_new_n3131_));
OR2X2 OR2X2_3835 ( .A(u5__abc_81276_new_n3127_), .B(u5__abc_81276_new_n3132_), .Y(u5__abc_81276_new_n3133_));
OR2X2 OR2X2_3836 ( .A(u5__abc_81276_new_n3134_), .B(u5__abc_81276_new_n3126_), .Y(u5__0timer2_8_0__7_));
OR2X2 OR2X2_3837 ( .A(u5__abc_81276_new_n3137_), .B(u5__abc_81276_new_n3139_), .Y(u5__abc_81276_new_n3140_));
OR2X2 OR2X2_3838 ( .A(u5__abc_81276_new_n3141_), .B(u5__abc_81276_new_n3136_), .Y(u5__0timer2_8_0__8_));
OR2X2 OR2X2_3839 ( .A(dv), .B(u5__abc_81276_new_n1829_), .Y(u5__abc_81276_new_n3145_));
OR2X2 OR2X2_384 ( .A(u0__abc_76628_new_n1791_), .B(u0__abc_76628_new_n1792_), .Y(u0__abc_76628_new_n1793_));
OR2X2 OR2X2_3840 ( .A(u5__abc_81276_new_n3146_), .B(u5__abc_81276_new_n3144_), .Y(u5__abc_81276_new_n3147_));
OR2X2 OR2X2_3841 ( .A(u5__abc_81276_new_n3148_), .B(u5__abc_81276_new_n3143_), .Y(u5__abc_81276_new_n3149_));
OR2X2 OR2X2_3842 ( .A(u5__abc_81276_new_n3147_), .B(u5_ack_cnt_0_), .Y(u5__abc_81276_new_n3151_));
OR2X2 OR2X2_3843 ( .A(u5__abc_81276_new_n3146_), .B(u5_ack_cnt_1_), .Y(u5__abc_81276_new_n3154_));
OR2X2 OR2X2_3844 ( .A(u5__abc_81276_new_n1818_), .B(u5__abc_81276_new_n3155_), .Y(u5__abc_81276_new_n3156_));
OR2X2 OR2X2_3845 ( .A(u5__abc_81276_new_n3145_), .B(u5__abc_81276_new_n3156_), .Y(u5__abc_81276_new_n3157_));
OR2X2 OR2X2_3846 ( .A(u5__abc_81276_new_n3158_), .B(u5__abc_81276_new_n3144_), .Y(u5__abc_81276_new_n3159_));
OR2X2 OR2X2_3847 ( .A(u5__abc_81276_new_n3164_), .B(u5__abc_81276_new_n3165_), .Y(u5__abc_81276_new_n3166_));
OR2X2 OR2X2_3848 ( .A(u5__abc_81276_new_n3167_), .B(u5__abc_81276_new_n1816_), .Y(u5__abc_81276_new_n3168_));
OR2X2 OR2X2_3849 ( .A(u5__abc_81276_new_n3166_), .B(u5_ack_cnt_2_), .Y(u5__abc_81276_new_n3169_));
OR2X2 OR2X2_385 ( .A(u0__abc_76628_new_n1795_), .B(spec_req_cs_0_bF_buf1_), .Y(u0__abc_76628_new_n1796_));
OR2X2 OR2X2_3850 ( .A(u5__abc_81276_new_n3145_), .B(u5__abc_81276_new_n3172_), .Y(u5__abc_81276_new_n3173_));
OR2X2 OR2X2_3851 ( .A(u5__abc_81276_new_n3174_), .B(u5__abc_81276_new_n3144_), .Y(u5__abc_81276_new_n3175_));
OR2X2 OR2X2_3852 ( .A(u5__abc_81276_new_n3176_), .B(u5__abc_81276_new_n1815_), .Y(u5__abc_81276_new_n3179_));
OR2X2 OR2X2_3853 ( .A(u5_mc_le), .B(u5_cmd_asserted_bF_buf0), .Y(u5__abc_81276_new_n3185_));
OR2X2 OR2X2_3854 ( .A(u5__0mc_le_0_0_), .B(u5_cmd_asserted2), .Y(u5__abc_81276_new_n3186_));
OR2X2 OR2X2_3855 ( .A(u5__abc_81276_new_n3189_), .B(u5__abc_81276_new_n3188_), .Y(u5__0cmd_asserted_0_0_));
OR2X2 OR2X2_3856 ( .A(u5_mc_le), .B(u5_mc_adv_r1), .Y(u5__abc_81276_new_n3191_));
OR2X2 OR2X2_3857 ( .A(u5__0mc_le_0_0_), .B(u5_mc_adv_r), .Y(u5__abc_81276_new_n3192_));
OR2X2 OR2X2_3858 ( .A(u5__abc_81276_new_n3194_), .B(u5__abc_81276_new_n1536_), .Y(u5__abc_81276_new_n3195_));
OR2X2 OR2X2_3859 ( .A(u5__abc_81276_new_n3204_), .B(u5__abc_81276_new_n3203_), .Y(u5__0mc_adv_r1_0_0_));
OR2X2 OR2X2_386 ( .A(u0__abc_76628_new_n1794_), .B(u0__abc_76628_new_n1796_), .Y(u0__abc_76628_new_n1797_));
OR2X2 OR2X2_3860 ( .A(u5__abc_81276_new_n1155_), .B(u5__abc_81276_new_n1518_), .Y(u5__abc_81276_new_n3206_));
OR2X2 OR2X2_3861 ( .A(u5__abc_81276_new_n3208_), .B(u5_cmd_asserted2), .Y(u5__abc_81276_new_n3209_));
OR2X2 OR2X2_3862 ( .A(u5__abc_81276_new_n1549_), .B(u5__abc_81276_new_n3209_), .Y(u5__abc_81276_new_n3210_));
OR2X2 OR2X2_3863 ( .A(u5__abc_81276_new_n3211_), .B(u5_wb_wait), .Y(u5__abc_81276_new_n3212_));
OR2X2 OR2X2_3864 ( .A(u5__abc_81276_new_n3215__bF_buf4), .B(u5__abc_81276_new_n3207_), .Y(u5__abc_81276_new_n3216_));
OR2X2 OR2X2_3865 ( .A(u5__abc_81276_new_n1552_), .B(u5_cs_le_r), .Y(u5__abc_81276_new_n3219_));
OR2X2 OR2X2_3866 ( .A(u5__abc_81276_new_n3220_), .B(u5__abc_81276_new_n1708_), .Y(u5__abc_81276_new_n3221_));
OR2X2 OR2X2_3867 ( .A(u5__abc_81276_new_n3223_), .B(u5_state_1_), .Y(u5__abc_81276_new_n3224_));
OR2X2 OR2X2_3868 ( .A(u5__abc_81276_new_n3218_), .B(u5__abc_81276_new_n3225_), .Y(u5__abc_81276_new_n3226_));
OR2X2 OR2X2_3869 ( .A(u5_state_1_), .B(u5_tmr_done_bF_buf2), .Y(u5__abc_81276_new_n3227_));
OR2X2 OR2X2_387 ( .A(u0__abc_76628_new_n1197__bF_buf4), .B(u0_tms0_25_), .Y(u0__abc_76628_new_n1798_));
OR2X2 OR2X2_3870 ( .A(u5__abc_81276_new_n3232_), .B(u5__abc_81276_new_n3229_), .Y(u5__abc_81276_new_n3233_));
OR2X2 OR2X2_3871 ( .A(u5__abc_81276_new_n3234_), .B(u5__abc_81276_new_n1231_), .Y(u5__abc_81276_new_n3235_));
OR2X2 OR2X2_3872 ( .A(u5__abc_81276_new_n3228_), .B(u5__abc_81276_new_n3235_), .Y(u5__abc_81276_new_n3236_));
OR2X2 OR2X2_3873 ( .A(u5__abc_81276_new_n3236_), .B(u5__abc_81276_new_n3226_), .Y(u5_next_state_1_));
OR2X2 OR2X2_3874 ( .A(u5__abc_81276_new_n3243_), .B(u5_state_2_), .Y(u5__abc_81276_new_n3244_));
OR2X2 OR2X2_3875 ( .A(u5__abc_81276_new_n3239_), .B(u5__abc_81276_new_n3244_), .Y(u5__abc_81276_new_n3245_));
OR2X2 OR2X2_3876 ( .A(u5__abc_81276_new_n3248_), .B(u5__abc_81276_new_n3249_), .Y(u5__abc_81276_new_n3250_));
OR2X2 OR2X2_3877 ( .A(u5__abc_81276_new_n3247_), .B(u5__abc_81276_new_n3250_), .Y(u5__abc_81276_new_n3251_));
OR2X2 OR2X2_3878 ( .A(u5__abc_81276_new_n1620_), .B(u5_state_2_), .Y(u5__abc_81276_new_n3252_));
OR2X2 OR2X2_3879 ( .A(u5__abc_81276_new_n3216_), .B(u5__abc_81276_new_n3255_), .Y(u5__abc_81276_new_n3256_));
OR2X2 OR2X2_388 ( .A(u0__abc_76628_new_n1800_), .B(u0__abc_76628_new_n1778_), .Y(u0__0sp_tms_31_0__25_));
OR2X2 OR2X2_3880 ( .A(u5_state_2_), .B(u5_cmd_asserted_bF_buf1), .Y(u5__abc_81276_new_n3258_));
OR2X2 OR2X2_3881 ( .A(u5__abc_81276_new_n1701_), .B(u5__abc_81276_new_n1510_), .Y(u5__abc_81276_new_n3259_));
OR2X2 OR2X2_3882 ( .A(u5__abc_81276_new_n3208_), .B(u5_state_2_), .Y(u5__abc_81276_new_n3261_));
OR2X2 OR2X2_3883 ( .A(u5__abc_81276_new_n3262_), .B(u5__abc_81276_new_n1132_), .Y(u5__abc_81276_new_n3263_));
OR2X2 OR2X2_3884 ( .A(u5__abc_81276_new_n3263_), .B(u5__abc_81276_new_n1627_), .Y(u5__abc_81276_new_n3264_));
OR2X2 OR2X2_3885 ( .A(u5__abc_81276_new_n3267_), .B(u5_state_2_), .Y(u5__abc_81276_new_n3268_));
OR2X2 OR2X2_3886 ( .A(u5__abc_81276_new_n3230_), .B(u5_state_2_), .Y(u5__abc_81276_new_n3274_));
OR2X2 OR2X2_3887 ( .A(u5__abc_81276_new_n3273_), .B(u5__abc_81276_new_n3277_), .Y(u5__abc_81276_new_n3278_));
OR2X2 OR2X2_3888 ( .A(u5__abc_81276_new_n3264_), .B(u5__abc_81276_new_n3278_), .Y(u5__abc_81276_new_n3279_));
OR2X2 OR2X2_3889 ( .A(u5__abc_81276_new_n3279_), .B(u5__abc_81276_new_n3260_), .Y(u5__abc_81276_new_n3280_));
OR2X2 OR2X2_389 ( .A(u0__abc_76628_new_n1177__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n1804_));
OR2X2 OR2X2_3890 ( .A(u5__abc_81276_new_n3257_), .B(u5__abc_81276_new_n3280_), .Y(u5__abc_81276_new_n3281_));
OR2X2 OR2X2_3891 ( .A(u5__abc_81276_new_n3285_), .B(u5__abc_81276_new_n2953__bF_buf1), .Y(u5__abc_81276_new_n3286_));
OR2X2 OR2X2_3892 ( .A(u5__abc_81276_new_n3282_), .B(u5__abc_81276_new_n3286_), .Y(u5__abc_81276_new_n3287_));
OR2X2 OR2X2_3893 ( .A(u5__abc_81276_new_n3289_), .B(u5__abc_81276_new_n3281_), .Y(u5__abc_81276_new_n3290_));
OR2X2 OR2X2_3894 ( .A(u5__abc_81276_new_n3254_), .B(u5__abc_81276_new_n3290_), .Y(u5_next_state_2_));
OR2X2 OR2X2_3895 ( .A(u5__abc_81276_new_n1848_), .B(u5__abc_81276_new_n3296_), .Y(u5__abc_81276_new_n3297_));
OR2X2 OR2X2_3896 ( .A(u5__abc_81276_new_n3293_), .B(u5__abc_81276_new_n3297_), .Y(u5_next_state_3_));
OR2X2 OR2X2_3897 ( .A(u5__abc_81276_new_n1549_), .B(u5__abc_81276_new_n3300_), .Y(u5__abc_81276_new_n3301_));
OR2X2 OR2X2_3898 ( .A(u5__abc_81276_new_n3310_), .B(u5__abc_81276_new_n3309_), .Y(u5__abc_81276_new_n3311_));
OR2X2 OR2X2_3899 ( .A(u5__abc_81276_new_n3312_), .B(rfr_req), .Y(u5__abc_81276_new_n3313_));
OR2X2 OR2X2_39 ( .A(_abc_85006_new_n240__bF_buf1), .B(sp_tms_2_), .Y(_abc_85006_new_n296_));
OR2X2 OR2X2_390 ( .A(spec_req_cs_6_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n1805_));
OR2X2 OR2X2_3900 ( .A(u5__abc_81276_new_n3314_), .B(u5__abc_81276_new_n3315_), .Y(u5_next_state_4_));
OR2X2 OR2X2_3901 ( .A(u5__abc_81276_new_n3215__bF_buf3), .B(u5__abc_81276_new_n3317_), .Y(u5__abc_81276_new_n3318_));
OR2X2 OR2X2_3902 ( .A(u5_state_5_), .B(u5_cmd_asserted_bF_buf0), .Y(u5__abc_81276_new_n3320_));
OR2X2 OR2X2_3903 ( .A(u5__abc_81276_new_n3319_), .B(u5__abc_81276_new_n3321_), .Y(u5_next_state_5_));
OR2X2 OR2X2_3904 ( .A(u5__abc_81276_new_n3328_), .B(u5__abc_81276_new_n3211_), .Y(u5__abc_81276_new_n3329_));
OR2X2 OR2X2_3905 ( .A(u5__abc_81276_new_n3331_), .B(u5_state_6_), .Y(u5__abc_81276_new_n3332_));
OR2X2 OR2X2_3906 ( .A(u5_state_6_), .B(u5_tmr_done_bF_buf3), .Y(u5__abc_81276_new_n3338_));
OR2X2 OR2X2_3907 ( .A(u5__abc_81276_new_n3340_), .B(u5__abc_81276_new_n3343_), .Y(u5__abc_81276_new_n3344_));
OR2X2 OR2X2_3908 ( .A(u5__abc_81276_new_n3335_), .B(u5__abc_81276_new_n3344_), .Y(u5_next_state_6_));
OR2X2 OR2X2_3909 ( .A(u5_state_7_), .B(u5_cmd_asserted_bF_buf3), .Y(u5__abc_81276_new_n3350_));
OR2X2 OR2X2_391 ( .A(u0__abc_76628_new_n1807_), .B(u0__abc_76628_new_n1803_), .Y(u0__abc_76628_new_n1808_));
OR2X2 OR2X2_3910 ( .A(u5__abc_81276_new_n3351_), .B(u5__abc_81276_new_n3358_), .Y(u5__abc_81276_new_n3359_));
OR2X2 OR2X2_3911 ( .A(u5__abc_81276_new_n3349_), .B(u5__abc_81276_new_n3359_), .Y(u5_next_state_7_));
OR2X2 OR2X2_3912 ( .A(u5__abc_81276_new_n3364_), .B(u5__abc_81276_new_n3363_), .Y(u5__abc_81276_new_n3365_));
OR2X2 OR2X2_3913 ( .A(u5__abc_81276_new_n3211_), .B(u5__abc_81276_new_n3368_), .Y(u5__abc_81276_new_n3369_));
OR2X2 OR2X2_3914 ( .A(u5__abc_81276_new_n3369_), .B(u5__abc_81276_new_n3366_), .Y(u5__abc_81276_new_n3370_));
OR2X2 OR2X2_3915 ( .A(u5__abc_81276_new_n1549_), .B(u5_state_8_), .Y(u5__abc_81276_new_n3371_));
OR2X2 OR2X2_3916 ( .A(u5__abc_81276_new_n3377_), .B(u5__abc_81276_new_n3367_), .Y(u5__abc_81276_new_n3378_));
OR2X2 OR2X2_3917 ( .A(u5__abc_81276_new_n3373_), .B(u5__abc_81276_new_n3379_), .Y(u5_next_state_8_));
OR2X2 OR2X2_3918 ( .A(u5__abc_81276_new_n3381_), .B(u5_state_9_), .Y(u5__abc_81276_new_n3382_));
OR2X2 OR2X2_3919 ( .A(u5__abc_81276_new_n3211_), .B(u5__abc_81276_new_n3384_), .Y(u5__abc_81276_new_n3385_));
OR2X2 OR2X2_392 ( .A(u0__abc_76628_new_n1809_), .B(u0__abc_76628_new_n1810_), .Y(u0__abc_76628_new_n1811_));
OR2X2 OR2X2_3920 ( .A(u5__abc_81276_new_n3385_), .B(u5__abc_81276_new_n3383_), .Y(u5__abc_81276_new_n3386_));
OR2X2 OR2X2_3921 ( .A(u5__abc_81276_new_n3354_), .B(u5_state_9_), .Y(u5__abc_81276_new_n3393_));
OR2X2 OR2X2_3922 ( .A(u5__abc_81276_new_n1693_), .B(u5__abc_81276_new_n3383_), .Y(u5__abc_81276_new_n3396_));
OR2X2 OR2X2_3923 ( .A(u5__abc_81276_new_n3395_), .B(u5__abc_81276_new_n3397_), .Y(u5__abc_81276_new_n3398_));
OR2X2 OR2X2_3924 ( .A(u5__abc_81276_new_n3398_), .B(u5__abc_81276_new_n3392_), .Y(u5__abc_81276_new_n3399_));
OR2X2 OR2X2_3925 ( .A(u5__abc_81276_new_n3388_), .B(u5__abc_81276_new_n3400_), .Y(u5_next_state_9_));
OR2X2 OR2X2_3926 ( .A(u5__abc_81276_new_n3404_), .B(u5__abc_81276_new_n3405_), .Y(u5__abc_81276_new_n3406_));
OR2X2 OR2X2_3927 ( .A(u5__abc_81276_new_n3403_), .B(u5__abc_81276_new_n3406_), .Y(u5_next_state_10_));
OR2X2 OR2X2_3928 ( .A(u5__abc_81276_new_n3239_), .B(u5_wb_cycle), .Y(u5__abc_81276_new_n3409_));
OR2X2 OR2X2_3929 ( .A(u5_state_11_), .B(u5_tmr_done_bF_buf1), .Y(u5__abc_81276_new_n3417_));
OR2X2 OR2X2_393 ( .A(u0__abc_76628_new_n1812_), .B(u0__abc_76628_new_n1813_), .Y(u0__abc_76628_new_n1814_));
OR2X2 OR2X2_3930 ( .A(u5__abc_81276_new_n3416_), .B(u5__abc_81276_new_n3418_), .Y(u5__abc_81276_new_n3419_));
OR2X2 OR2X2_3931 ( .A(u5__abc_81276_new_n3414_), .B(u5__abc_81276_new_n3419_), .Y(u5_next_state_11_));
OR2X2 OR2X2_3932 ( .A(u5__abc_81276_new_n3239_), .B(u5_state_12_), .Y(u5__abc_81276_new_n3421_));
OR2X2 OR2X2_3933 ( .A(u5__abc_81276_new_n3424_), .B(u5__abc_81276_new_n3427_), .Y(u5__abc_81276_new_n3428_));
OR2X2 OR2X2_3934 ( .A(u5__abc_81276_new_n3422_), .B(u5__abc_81276_new_n3428_), .Y(u5_next_state_12_));
OR2X2 OR2X2_3935 ( .A(u5__abc_81276_new_n1733_), .B(u5__abc_81276_new_n3433_), .Y(u5__abc_81276_new_n3434_));
OR2X2 OR2X2_3936 ( .A(u5__abc_81276_new_n3434_), .B(u5__abc_81276_new_n3432_), .Y(u5__abc_81276_new_n3435_));
OR2X2 OR2X2_3937 ( .A(u5__abc_81276_new_n3431_), .B(u5__abc_81276_new_n3435_), .Y(u5_next_state_13_));
OR2X2 OR2X2_3938 ( .A(u5__abc_81276_new_n3437_), .B(u5__abc_81276_new_n2953__bF_buf0), .Y(u5__abc_81276_new_n3438_));
OR2X2 OR2X2_3939 ( .A(u5_state_14_), .B(u5_cmd_asserted_bF_buf1), .Y(u5__abc_81276_new_n3439_));
OR2X2 OR2X2_394 ( .A(u0__abc_76628_new_n1815_), .B(u0__abc_76628_new_n1816_), .Y(u0__abc_76628_new_n1817_));
OR2X2 OR2X2_3940 ( .A(u5__abc_81276_new_n3449_), .B(u5__abc_81276_new_n3248_), .Y(u5__abc_81276_new_n3450_));
OR2X2 OR2X2_3941 ( .A(u5__abc_81276_new_n3451_), .B(u5__abc_81276_new_n3445_), .Y(u5__abc_81276_new_n3452_));
OR2X2 OR2X2_3942 ( .A(u5__abc_81276_new_n3444_), .B(u5__abc_81276_new_n3452_), .Y(u5_next_state_14_));
OR2X2 OR2X2_3943 ( .A(u5__abc_81276_new_n3381_), .B(u5_state_15_), .Y(u5__abc_81276_new_n3455_));
OR2X2 OR2X2_3944 ( .A(u5__abc_81276_new_n3385_), .B(u5__abc_81276_new_n3456_), .Y(u5__abc_81276_new_n3457_));
OR2X2 OR2X2_3945 ( .A(u5__abc_81276_new_n3461_), .B(u5__abc_81276_new_n3460_), .Y(u5__abc_81276_new_n3462_));
OR2X2 OR2X2_3946 ( .A(u5__abc_81276_new_n3459_), .B(u5__abc_81276_new_n3463_), .Y(u5__abc_81276_new_n3464_));
OR2X2 OR2X2_3947 ( .A(u5__abc_81276_new_n3464_), .B(u5__abc_81276_new_n3454_), .Y(u5__abc_81276_new_n3465_));
OR2X2 OR2X2_3948 ( .A(u5__abc_81276_new_n1552_), .B(u5_state_15_), .Y(u5__abc_81276_new_n3466_));
OR2X2 OR2X2_3949 ( .A(u5__abc_81276_new_n3467_), .B(u5__abc_81276_new_n3410_), .Y(u5__abc_81276_new_n3468_));
OR2X2 OR2X2_395 ( .A(u0__abc_76628_new_n1819_), .B(spec_req_cs_0_bF_buf0_), .Y(u0__abc_76628_new_n1820_));
OR2X2 OR2X2_3950 ( .A(u5__abc_81276_new_n3469_), .B(u5__abc_81276_new_n3465_), .Y(u5__abc_81276_new_n3470_));
OR2X2 OR2X2_3951 ( .A(u5__abc_81276_new_n3472_), .B(u5__abc_81276_new_n1615_), .Y(u5__abc_81276_new_n3473_));
OR2X2 OR2X2_3952 ( .A(u5__abc_81276_new_n3474_), .B(u5__abc_81276_new_n3248_), .Y(u5__abc_81276_new_n3475_));
OR2X2 OR2X2_3953 ( .A(u5__abc_81276_new_n3476_), .B(u5__abc_81276_new_n3470_), .Y(u5_next_state_15_));
OR2X2 OR2X2_3954 ( .A(u5__abc_81276_new_n3479_), .B(u5__abc_81276_new_n2953__bF_buf1), .Y(u5__abc_81276_new_n3480_));
OR2X2 OR2X2_3955 ( .A(u5__abc_81276_new_n3487_), .B(u5__abc_81276_new_n3270_), .Y(u5__abc_81276_new_n3488_));
OR2X2 OR2X2_3956 ( .A(u5_state_16_), .B(u5_cmd_asserted_bF_buf3), .Y(u5__abc_81276_new_n3490_));
OR2X2 OR2X2_3957 ( .A(u5__abc_81276_new_n3489_), .B(u5__abc_81276_new_n3491_), .Y(u5__abc_81276_new_n3492_));
OR2X2 OR2X2_3958 ( .A(u5__abc_81276_new_n3492_), .B(u5__abc_81276_new_n3486_), .Y(u5__abc_81276_new_n3493_));
OR2X2 OR2X2_3959 ( .A(u5__abc_81276_new_n3484_), .B(u5__abc_81276_new_n3493_), .Y(u5__abc_81276_new_n3494_));
OR2X2 OR2X2_396 ( .A(u0__abc_76628_new_n1818_), .B(u0__abc_76628_new_n1820_), .Y(u0__abc_76628_new_n1821_));
OR2X2 OR2X2_3960 ( .A(u5__abc_81276_new_n3482_), .B(u5__abc_81276_new_n3494_), .Y(u5__abc_81276_new_n3495_));
OR2X2 OR2X2_3961 ( .A(u5__abc_81276_new_n3240_), .B(u5__abc_81276_new_n3497_), .Y(u5__abc_81276_new_n3498_));
OR2X2 OR2X2_3962 ( .A(u5__abc_81276_new_n3500_), .B(u5__abc_81276_new_n3248_), .Y(u5__abc_81276_new_n3501_));
OR2X2 OR2X2_3963 ( .A(u5__abc_81276_new_n3502_), .B(u5__abc_81276_new_n3495_), .Y(u5_next_state_16_));
OR2X2 OR2X2_3964 ( .A(u5__abc_81276_new_n3259_), .B(u5__abc_81276_new_n3507_), .Y(u5__abc_81276_new_n3508_));
OR2X2 OR2X2_3965 ( .A(u5_state_17_), .B(u5_tmr_done_bF_buf0), .Y(u5__abc_81276_new_n3510_));
OR2X2 OR2X2_3966 ( .A(u5__abc_81276_new_n3511_), .B(u5__abc_81276_new_n530_), .Y(u5__abc_81276_new_n3512_));
OR2X2 OR2X2_3967 ( .A(u5__abc_81276_new_n3514_), .B(u5__abc_81276_new_n3336_), .Y(u5__abc_81276_new_n3515_));
OR2X2 OR2X2_3968 ( .A(u5__abc_81276_new_n3513_), .B(u5__abc_81276_new_n3516_), .Y(u5__abc_81276_new_n3517_));
OR2X2 OR2X2_3969 ( .A(u5__abc_81276_new_n3509_), .B(u5__abc_81276_new_n3517_), .Y(u5__abc_81276_new_n3518_));
OR2X2 OR2X2_397 ( .A(u0__abc_76628_new_n1197__bF_buf3), .B(u0_tms0_26_), .Y(u0__abc_76628_new_n1822_));
OR2X2 OR2X2_3970 ( .A(u5__abc_81276_new_n3505_), .B(u5__abc_81276_new_n3518_), .Y(u5_next_state_17_));
OR2X2 OR2X2_3971 ( .A(u5__abc_81276_new_n3521_), .B(u5__abc_81276_new_n1550_), .Y(u5__abc_81276_new_n3522_));
OR2X2 OR2X2_3972 ( .A(u5__abc_81276_new_n3523_), .B(u5__abc_81276_new_n3524_), .Y(u5_next_state_18_));
OR2X2 OR2X2_3973 ( .A(u5_state_19_), .B(u5_cmd_asserted_bF_buf2), .Y(u5__abc_81276_new_n3531_));
OR2X2 OR2X2_3974 ( .A(u5__abc_81276_new_n3530_), .B(u5__abc_81276_new_n3532_), .Y(u5__abc_81276_new_n3533_));
OR2X2 OR2X2_3975 ( .A(u5__abc_81276_new_n3528_), .B(u5__abc_81276_new_n3533_), .Y(u5_next_state_19_));
OR2X2 OR2X2_3976 ( .A(u5_state_20_), .B(u5_tmr_done_bF_buf3), .Y(u5__abc_81276_new_n3539_));
OR2X2 OR2X2_3977 ( .A(u5__abc_81276_new_n3542_), .B(u5__abc_81276_new_n3540_), .Y(u5__abc_81276_new_n3543_));
OR2X2 OR2X2_3978 ( .A(u5__abc_81276_new_n3538_), .B(u5__abc_81276_new_n3543_), .Y(u5_next_state_20_));
OR2X2 OR2X2_3979 ( .A(u5__abc_81276_new_n3545_), .B(init_req), .Y(u5__abc_81276_new_n3546_));
OR2X2 OR2X2_398 ( .A(u0__abc_76628_new_n1824_), .B(u0__abc_76628_new_n1802_), .Y(u0__0sp_tms_31_0__26_));
OR2X2 OR2X2_3980 ( .A(u5__abc_81276_new_n3552_), .B(u5__abc_81276_new_n3550_), .Y(u5__abc_81276_new_n3553_));
OR2X2 OR2X2_3981 ( .A(u5__abc_81276_new_n3549_), .B(u5__abc_81276_new_n3553_), .Y(u5_next_state_22_));
OR2X2 OR2X2_3982 ( .A(u5_state_23_), .B(u5_cmd_asserted_bF_buf1), .Y(u5__abc_81276_new_n3557_));
OR2X2 OR2X2_3983 ( .A(u5__abc_81276_new_n3558_), .B(u5__abc_81276_new_n3560_), .Y(u5__abc_81276_new_n3561_));
OR2X2 OR2X2_3984 ( .A(u5__abc_81276_new_n3556_), .B(u5__abc_81276_new_n3561_), .Y(u5_next_state_23_));
OR2X2 OR2X2_3985 ( .A(u5__abc_81276_new_n1363_), .B(u5__abc_81276_new_n3566_), .Y(u5__abc_81276_new_n3567_));
OR2X2 OR2X2_3986 ( .A(u5__abc_81276_new_n546_), .B(u5__abc_81276_new_n646_), .Y(u5__abc_81276_new_n3568_));
OR2X2 OR2X2_3987 ( .A(u5_state_24_), .B(u5_tmr_done_bF_buf1), .Y(u5__abc_81276_new_n3569_));
OR2X2 OR2X2_3988 ( .A(u5__abc_81276_new_n3571_), .B(u5__abc_81276_new_n3572_), .Y(u5__abc_81276_new_n3573_));
OR2X2 OR2X2_3989 ( .A(u5__abc_81276_new_n3564_), .B(u5__abc_81276_new_n3573_), .Y(u5_next_state_24_));
OR2X2 OR2X2_399 ( .A(u0__abc_76628_new_n1177__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n1828_));
OR2X2 OR2X2_3990 ( .A(u5_state_25_), .B(u5_cmd_asserted_bF_buf0), .Y(u5__abc_81276_new_n3577_));
OR2X2 OR2X2_3991 ( .A(u5__abc_81276_new_n3578_), .B(u5__abc_81276_new_n3580_), .Y(u5__abc_81276_new_n3581_));
OR2X2 OR2X2_3992 ( .A(u5__abc_81276_new_n3576_), .B(u5__abc_81276_new_n3581_), .Y(u5_next_state_25_));
OR2X2 OR2X2_3993 ( .A(u5__abc_81276_new_n3585_), .B(u5__abc_81276_new_n3565_), .Y(u5__abc_81276_new_n3586_));
OR2X2 OR2X2_3994 ( .A(u5__abc_81276_new_n3589_), .B(u5__abc_81276_new_n3587_), .Y(u5__abc_81276_new_n3590_));
OR2X2 OR2X2_3995 ( .A(u5__abc_81276_new_n3584_), .B(u5__abc_81276_new_n3590_), .Y(u5_next_state_26_));
OR2X2 OR2X2_3996 ( .A(u5__abc_81276_new_n3593_), .B(u5__abc_81276_new_n1553_), .Y(u5__abc_81276_new_n3594_));
OR2X2 OR2X2_3997 ( .A(u5__abc_81276_new_n3595_), .B(u5__abc_81276_new_n3596_), .Y(u5_next_state_27_));
OR2X2 OR2X2_3998 ( .A(u5_state_28_), .B(u5_cmd_asserted_bF_buf3), .Y(u5__abc_81276_new_n3600_));
OR2X2 OR2X2_3999 ( .A(u5__abc_81276_new_n3511_), .B(u5__abc_81276_new_n3601_), .Y(u5__abc_81276_new_n3602_));
OR2X2 OR2X2_4 ( .A(lmr_sel_bF_buf6), .B(cs_0_), .Y(_abc_85006_new_n242_));
OR2X2 OR2X2_40 ( .A(lmr_sel_bF_buf3), .B(tms_2_), .Y(_abc_85006_new_n297_));
OR2X2 OR2X2_400 ( .A(spec_req_cs_6_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n1829_));
OR2X2 OR2X2_4000 ( .A(u5__abc_81276_new_n3599_), .B(u5__abc_81276_new_n3602_), .Y(u5_next_state_28_));
OR2X2 OR2X2_4001 ( .A(u5_state_29_), .B(u5_tmr_done_bF_buf0), .Y(u5__abc_81276_new_n3606_));
OR2X2 OR2X2_4002 ( .A(u5__abc_81276_new_n3607_), .B(u5__abc_81276_new_n3609_), .Y(u5__abc_81276_new_n3610_));
OR2X2 OR2X2_4003 ( .A(u5__abc_81276_new_n3605_), .B(u5__abc_81276_new_n3610_), .Y(u5_next_state_29_));
OR2X2 OR2X2_4004 ( .A(u5_state_30_), .B(u5_cmd_asserted_bF_buf2), .Y(u5__abc_81276_new_n3614_));
OR2X2 OR2X2_4005 ( .A(u5__abc_81276_new_n3615_), .B(u5__abc_81276_new_n3618_), .Y(u5__abc_81276_new_n3619_));
OR2X2 OR2X2_4006 ( .A(u5__abc_81276_new_n3613_), .B(u5__abc_81276_new_n3619_), .Y(u5_next_state_30_));
OR2X2 OR2X2_4007 ( .A(u5_state_31_), .B(u5_resume_req_r), .Y(u5__abc_81276_new_n3623_));
OR2X2 OR2X2_4008 ( .A(u5__abc_81276_new_n3622_), .B(u5__abc_81276_new_n3624_), .Y(u5_next_state_31_));
OR2X2 OR2X2_4009 ( .A(u5__abc_81276_new_n3629_), .B(u5__abc_81276_new_n537_), .Y(u5__abc_81276_new_n3630_));
OR2X2 OR2X2_401 ( .A(u0__abc_76628_new_n1831_), .B(u0__abc_76628_new_n1827_), .Y(u0__abc_76628_new_n1832_));
OR2X2 OR2X2_4010 ( .A(u5__abc_81276_new_n3627_), .B(u5__abc_81276_new_n3630_), .Y(u5_next_state_32_));
OR2X2 OR2X2_4011 ( .A(u5__abc_81276_new_n3632_), .B(u5_state_33_), .Y(u5__abc_81276_new_n3633_));
OR2X2 OR2X2_4012 ( .A(u5__abc_81276_new_n3636_), .B(u5__abc_81276_new_n1390_), .Y(u5_next_state_34_));
OR2X2 OR2X2_4013 ( .A(u5__abc_81276_new_n3639_), .B(u5__abc_81276_new_n1421_), .Y(u5__abc_81276_new_n3640_));
OR2X2 OR2X2_4014 ( .A(u5__abc_81276_new_n3638_), .B(u5__abc_81276_new_n3640_), .Y(u5_next_state_35_));
OR2X2 OR2X2_4015 ( .A(u5__abc_81276_new_n3211_), .B(u5__abc_81276_new_n3645_), .Y(u5__abc_81276_new_n3646_));
OR2X2 OR2X2_4016 ( .A(u5__abc_81276_new_n3643_), .B(u5__abc_81276_new_n3646_), .Y(u5__abc_81276_new_n3647_));
OR2X2 OR2X2_4017 ( .A(u5__abc_81276_new_n1549_), .B(u5_state_36_), .Y(u5__abc_81276_new_n3648_));
OR2X2 OR2X2_4018 ( .A(u5__abc_81276_new_n3655_), .B(u5__abc_81276_new_n1342_), .Y(u5__abc_81276_new_n3656_));
OR2X2 OR2X2_4019 ( .A(u5__abc_81276_new_n3652_), .B(u5__abc_81276_new_n3656_), .Y(u5_next_state_37_));
OR2X2 OR2X2_402 ( .A(u0__abc_76628_new_n1833_), .B(u0__abc_76628_new_n1834_), .Y(u0__abc_76628_new_n1835_));
OR2X2 OR2X2_4020 ( .A(u5_state_38_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3660_));
OR2X2 OR2X2_4021 ( .A(u5__abc_81276_new_n3658_), .B(u5__abc_81276_new_n3664_), .Y(u5_next_state_38_));
OR2X2 OR2X2_4022 ( .A(u5_state_39_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3667_));
OR2X2 OR2X2_4023 ( .A(u5__abc_81276_new_n3668_), .B(u5__abc_81276_new_n775_), .Y(u5__abc_81276_new_n3669_));
OR2X2 OR2X2_4024 ( .A(u5__abc_81276_new_n3666_), .B(u5__abc_81276_new_n3669_), .Y(u5_next_state_39_));
OR2X2 OR2X2_4025 ( .A(u5__abc_81276_new_n3671_), .B(u5__abc_81276_new_n1247_), .Y(u5_next_state_40_));
OR2X2 OR2X2_4026 ( .A(u5__abc_81276_new_n1751_), .B(u5__abc_81276_new_n1708_), .Y(u5__abc_81276_new_n3674_));
OR2X2 OR2X2_4027 ( .A(u5_state_41_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3675_));
OR2X2 OR2X2_4028 ( .A(u5__abc_81276_new_n3673_), .B(u5__abc_81276_new_n3677_), .Y(u5_next_state_41_));
OR2X2 OR2X2_4029 ( .A(u5__abc_81276_new_n3681_), .B(u5__abc_81276_new_n1329_), .Y(u5__abc_81276_new_n3682_));
OR2X2 OR2X2_403 ( .A(u0__abc_76628_new_n1836_), .B(u0__abc_76628_new_n1837_), .Y(u0__abc_76628_new_n1838_));
OR2X2 OR2X2_4030 ( .A(u5__abc_81276_new_n3679_), .B(u5__abc_81276_new_n3682_), .Y(u5_next_state_42_));
OR2X2 OR2X2_4031 ( .A(u5__abc_81276_new_n3684_), .B(u5_state_43_), .Y(u5__abc_81276_new_n3685_));
OR2X2 OR2X2_4032 ( .A(u5__abc_81276_new_n3215__bF_buf3), .B(u5__abc_81276_new_n1323_), .Y(u5__abc_81276_new_n3686_));
OR2X2 OR2X2_4033 ( .A(u5__abc_81276_new_n3688_), .B(u5__abc_81276_new_n3690_), .Y(u5__abc_81276_new_n3691_));
OR2X2 OR2X2_4034 ( .A(u5__abc_81276_new_n3691_), .B(u5__abc_81276_new_n791_), .Y(u5_next_state_44_));
OR2X2 OR2X2_4035 ( .A(u5_state_45_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3694_));
OR2X2 OR2X2_4036 ( .A(u5__abc_81276_new_n3695_), .B(u5__abc_81276_new_n1708_), .Y(u5__abc_81276_new_n3696_));
OR2X2 OR2X2_4037 ( .A(u5__abc_81276_new_n3697_), .B(u5__abc_81276_new_n1296_), .Y(u5__abc_81276_new_n3698_));
OR2X2 OR2X2_4038 ( .A(u5__abc_81276_new_n3693_), .B(u5__abc_81276_new_n3699_), .Y(u5_next_state_45_));
OR2X2 OR2X2_4039 ( .A(u5__abc_81276_new_n3703_), .B(u5__abc_81276_new_n1315_), .Y(u5__abc_81276_new_n3704_));
OR2X2 OR2X2_404 ( .A(u0__abc_76628_new_n1839_), .B(u0__abc_76628_new_n1840_), .Y(u0__abc_76628_new_n1841_));
OR2X2 OR2X2_4040 ( .A(u5__abc_81276_new_n3701_), .B(u5__abc_81276_new_n3704_), .Y(u5_next_state_46_));
OR2X2 OR2X2_4041 ( .A(u5__abc_81276_new_n3706_), .B(u5__abc_81276_new_n3708_), .Y(u5__abc_81276_new_n3709_));
OR2X2 OR2X2_4042 ( .A(u5__abc_81276_new_n3713_), .B(u5__abc_81276_new_n727_), .Y(u5__abc_81276_new_n3714_));
OR2X2 OR2X2_4043 ( .A(u5__abc_81276_new_n3714_), .B(u5__abc_81276_new_n3712_), .Y(u5_next_state_48_));
OR2X2 OR2X2_4044 ( .A(u5__abc_81276_new_n3716_), .B(u5_state_49_), .Y(u5__abc_81276_new_n3717_));
OR2X2 OR2X2_4045 ( .A(u5__abc_81276_new_n3215__bF_buf3), .B(u5__abc_81276_new_n1287_), .Y(u5__abc_81276_new_n3718_));
OR2X2 OR2X2_4046 ( .A(u5__abc_81276_new_n1709_), .B(u5__abc_81276_new_n1281_), .Y(u5__abc_81276_new_n3721_));
OR2X2 OR2X2_4047 ( .A(u5__abc_81276_new_n3720_), .B(u5__abc_81276_new_n3721_), .Y(u5_next_state_50_));
OR2X2 OR2X2_4048 ( .A(u5__abc_81276_new_n3723_), .B(u5_state_51_), .Y(u5__abc_81276_new_n3724_));
OR2X2 OR2X2_4049 ( .A(u5__abc_81276_new_n3215__bF_buf1), .B(u5__abc_81276_new_n1270_), .Y(u5__abc_81276_new_n3725_));
OR2X2 OR2X2_405 ( .A(u0__abc_76628_new_n1843_), .B(spec_req_cs_0_bF_buf5_), .Y(u0__abc_76628_new_n1844_));
OR2X2 OR2X2_4050 ( .A(u5__abc_81276_new_n3727_), .B(u5__abc_81276_new_n3729_), .Y(u5__abc_81276_new_n3730_));
OR2X2 OR2X2_4051 ( .A(u5__abc_81276_new_n1536_), .B(u5_state_52_), .Y(u5__abc_81276_new_n3732_));
OR2X2 OR2X2_4052 ( .A(u5__abc_81276_new_n3734_), .B(u5__abc_81276_new_n3736_), .Y(u5__abc_81276_new_n3737_));
OR2X2 OR2X2_4053 ( .A(u5__abc_81276_new_n3731_), .B(u5__abc_81276_new_n3737_), .Y(u5_next_state_52_));
OR2X2 OR2X2_4054 ( .A(u5_state_53_), .B(u5_cmd_asserted_bF_buf1), .Y(u5__abc_81276_new_n3741_));
OR2X2 OR2X2_4055 ( .A(u5__abc_81276_new_n3740_), .B(u5__abc_81276_new_n3742_), .Y(u5__abc_81276_new_n3743_));
OR2X2 OR2X2_4056 ( .A(u5__abc_81276_new_n3739_), .B(u5__abc_81276_new_n3743_), .Y(u5_next_state_53_));
OR2X2 OR2X2_4057 ( .A(u5__abc_81276_new_n3747_), .B(u5_state_54_), .Y(u5__abc_81276_new_n3748_));
OR2X2 OR2X2_4058 ( .A(u5__abc_81276_new_n3215__bF_buf4), .B(u5__abc_81276_new_n1206_), .Y(u5__abc_81276_new_n3749_));
OR2X2 OR2X2_4059 ( .A(u5__abc_81276_new_n3746_), .B(u5__abc_81276_new_n3750_), .Y(u5_next_state_54_));
OR2X2 OR2X2_406 ( .A(u0__abc_76628_new_n1842_), .B(u0__abc_76628_new_n1844_), .Y(u0__abc_76628_new_n1845_));
OR2X2 OR2X2_4060 ( .A(u5__abc_81276_new_n3752_), .B(u5_state_55_), .Y(u5__abc_81276_new_n3753_));
OR2X2 OR2X2_4061 ( .A(u5__abc_81276_new_n3381_), .B(u5_state_55_), .Y(u5__abc_81276_new_n3755_));
OR2X2 OR2X2_4062 ( .A(u5__abc_81276_new_n3385_), .B(u5__abc_81276_new_n3756_), .Y(u5__abc_81276_new_n3757_));
OR2X2 OR2X2_4063 ( .A(u5__abc_81276_new_n3759_), .B(u5__abc_81276_new_n3762_), .Y(u5__abc_81276_new_n3763_));
OR2X2 OR2X2_4064 ( .A(u5__abc_81276_new_n3754_), .B(u5__abc_81276_new_n3763_), .Y(u5_next_state_55_));
OR2X2 OR2X2_4065 ( .A(u5__abc_81276_new_n3381_), .B(u5_state_56_), .Y(u5__abc_81276_new_n3765_));
OR2X2 OR2X2_4066 ( .A(u5__abc_81276_new_n3385_), .B(u5__abc_81276_new_n3766_), .Y(u5__abc_81276_new_n3767_));
OR2X2 OR2X2_4067 ( .A(u5__abc_81276_new_n1820_), .B(u5_state_56_), .Y(u5__abc_81276_new_n3771_));
OR2X2 OR2X2_4068 ( .A(u5__abc_81276_new_n3773_), .B(u5__abc_81276_new_n3770_), .Y(u5__abc_81276_new_n3774_));
OR2X2 OR2X2_4069 ( .A(u5__abc_81276_new_n3769_), .B(u5__abc_81276_new_n3774_), .Y(u5_next_state_56_));
OR2X2 OR2X2_407 ( .A(u0__abc_76628_new_n1197__bF_buf2), .B(u0_tms0_27_), .Y(u0__abc_76628_new_n1846_));
OR2X2 OR2X2_4070 ( .A(u5__abc_81276_new_n3440_), .B(u5_state_57_), .Y(u5__abc_81276_new_n3781_));
OR2X2 OR2X2_4071 ( .A(u5__abc_81276_new_n3783_), .B(u5__abc_81276_new_n3784_), .Y(u5__abc_81276_new_n3785_));
OR2X2 OR2X2_4072 ( .A(u5__abc_81276_new_n3785_), .B(u5__abc_81276_new_n3778_), .Y(u5__abc_81276_new_n3786_));
OR2X2 OR2X2_4073 ( .A(u5__abc_81276_new_n3776_), .B(u5__abc_81276_new_n3786_), .Y(u5_next_state_57_));
OR2X2 OR2X2_4074 ( .A(u5__abc_81276_new_n3789_), .B(u5__abc_81276_new_n3788_), .Y(u5__abc_81276_new_n3790_));
OR2X2 OR2X2_4075 ( .A(u5__abc_81276_new_n3794_), .B(u5__abc_81276_new_n1734_), .Y(u5__abc_81276_new_n3795_));
OR2X2 OR2X2_4076 ( .A(u5__abc_81276_new_n3791_), .B(u5__abc_81276_new_n3795_), .Y(u5_next_state_58_));
OR2X2 OR2X2_4077 ( .A(u5__abc_81276_new_n3798_), .B(u5__abc_81276_new_n3779_), .Y(u5__abc_81276_new_n3799_));
OR2X2 OR2X2_4078 ( .A(u5__abc_81276_new_n3800_), .B(u5__abc_81276_new_n3801_), .Y(u5__abc_81276_new_n3802_));
OR2X2 OR2X2_4079 ( .A(u5__abc_81276_new_n3797_), .B(u5__abc_81276_new_n3802_), .Y(u5_next_state_59_));
OR2X2 OR2X2_408 ( .A(u0__abc_76628_new_n1848_), .B(u0__abc_76628_new_n1826_), .Y(u0__0sp_tms_31_0__27_));
OR2X2 OR2X2_4080 ( .A(u5__abc_81276_new_n3804_), .B(u5__abc_81276_new_n3806_), .Y(u5__abc_81276_new_n3807_));
OR2X2 OR2X2_4081 ( .A(u5__abc_81276_new_n3808_), .B(u5__abc_81276_new_n3812_), .Y(u5_next_state_60_));
OR2X2 OR2X2_4082 ( .A(u5__abc_81276_new_n3817_), .B(mc_ack_r), .Y(u5__abc_81276_new_n3818_));
OR2X2 OR2X2_4083 ( .A(u5__abc_81276_new_n3816_), .B(u5__abc_81276_new_n3819_), .Y(u5__abc_81276_new_n3820_));
OR2X2 OR2X2_4084 ( .A(u5__abc_81276_new_n3814_), .B(u5__abc_81276_new_n3820_), .Y(u5_next_state_61_));
OR2X2 OR2X2_4085 ( .A(u5__abc_81276_new_n3822_), .B(u5_state_62_), .Y(u5__abc_81276_new_n3823_));
OR2X2 OR2X2_4086 ( .A(u5__abc_81276_new_n3215__bF_buf0), .B(u5__abc_81276_new_n1141_), .Y(u5__abc_81276_new_n3824_));
OR2X2 OR2X2_4087 ( .A(u5__abc_81276_new_n3827_), .B(u5__abc_81276_new_n3826_), .Y(u5__abc_81276_new_n3828_));
OR2X2 OR2X2_4088 ( .A(u5__abc_81276_new_n3829_), .B(u5__abc_81276_new_n3830_), .Y(u5_next_state_63_));
OR2X2 OR2X2_4089 ( .A(u5__abc_81276_new_n3833_), .B(mc_ack_r), .Y(u5__abc_81276_new_n3834_));
OR2X2 OR2X2_409 ( .A(u0__abc_76628_new_n1177__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n1974_));
OR2X2 OR2X2_4090 ( .A(u5__abc_81276_new_n1713_), .B(u5__abc_81276_new_n3835_), .Y(u5__abc_81276_new_n3836_));
OR2X2 OR2X2_4091 ( .A(u5__abc_81276_new_n3832_), .B(u5__abc_81276_new_n3836_), .Y(u5_next_state_64_));
OR2X2 OR2X2_4092 ( .A(u5_state_65_), .B(u5_tmr2_done), .Y(u5__abc_81276_new_n3838_));
OR2X2 OR2X2_4093 ( .A(u5__abc_81276_new_n3839_), .B(u5__abc_81276_new_n3841_), .Y(u5__abc_81276_new_n3842_));
OR2X2 OR2X2_4094 ( .A(u5__abc_81276_new_n3856_), .B(u5__abc_81276_new_n1536_), .Y(u5__abc_81276_new_n3857_));
OR2X2 OR2X2_4095 ( .A(u5__abc_81276_new_n3855_), .B(u5_cke_r), .Y(u5__abc_81276_new_n3858_));
OR2X2 OR2X2_4096 ( .A(u5__abc_81276_new_n1094_), .B(u5_cke_r), .Y(u5__abc_81276_new_n3862_));
OR2X2 OR2X2_4097 ( .A(u5__abc_81276_new_n1536_), .B(u5_cnt), .Y(u5__abc_81276_new_n3863_));
OR2X2 OR2X2_4098 ( .A(u5__abc_81276_new_n3861_), .B(u5__abc_81276_new_n3873_), .Y(u5_cke_d));
OR2X2 OR2X2_4099 ( .A(u5__abc_81276_new_n3883_), .B(u5__abc_81276_new_n3875_), .Y(u5_lmr_ack_d));
OR2X2 OR2X2_41 ( .A(_abc_85006_new_n240__bF_buf0), .B(sp_tms_3_), .Y(_abc_85006_new_n299_));
OR2X2 OR2X2_410 ( .A(spec_req_cs_6_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n1975_));
OR2X2 OR2X2_4100 ( .A(u5__abc_81276_new_n3885_), .B(u5__abc_81276_new_n1849_), .Y(u5__abc_81276_new_n3886_));
OR2X2 OR2X2_4101 ( .A(u5__abc_81276_new_n3886_), .B(u5__abc_81276_new_n3784_), .Y(u5__abc_81276_new_n3887_));
OR2X2 OR2X2_4102 ( .A(u5__abc_81276_new_n3887_), .B(u5__abc_81276_new_n3778_), .Y(u5__abc_81276_new_n3888_));
OR2X2 OR2X2_4103 ( .A(u5__abc_81276_new_n1696_), .B(u5__abc_81276_new_n3888_), .Y(mc_adsc_d));
OR2X2 OR2X2_4104 ( .A(u5__abc_81276_new_n3903_), .B(u5__abc_81276_new_n3895_), .Y(mc_bg_d));
OR2X2 OR2X2_4105 ( .A(u5__abc_81276_new_n3906_), .B(u5__abc_81276_new_n3905_), .Y(u5__abc_81276_new_n3907_));
OR2X2 OR2X2_4106 ( .A(u5__abc_81276_new_n3912_), .B(u5__abc_81276_new_n1231_), .Y(u5__abc_81276_new_n3913_));
OR2X2 OR2X2_4107 ( .A(u5__abc_81276_new_n3913_), .B(u5__abc_81276_new_n3911_), .Y(u5__abc_81276_new_n3914_));
OR2X2 OR2X2_4108 ( .A(u5__abc_81276_new_n3550_), .B(u5__abc_81276_new_n1421_), .Y(u5__abc_81276_new_n3919_));
OR2X2 OR2X2_4109 ( .A(u5__abc_81276_new_n1428_), .B(u5__abc_81276_new_n1510_), .Y(u5__abc_81276_new_n3920_));
OR2X2 OR2X2_411 ( .A(u0__abc_76628_new_n1977_), .B(u0__abc_76628_new_n1973_), .Y(u0__abc_76628_new_n1978_));
OR2X2 OR2X2_4110 ( .A(u5__abc_81276_new_n3919_), .B(u5__abc_81276_new_n3920_), .Y(u5__abc_81276_new_n3921_));
OR2X2 OR2X2_4111 ( .A(u5__abc_81276_new_n3921_), .B(u5__abc_81276_new_n3918_), .Y(u5__abc_81276_new_n3922_));
OR2X2 OR2X2_4112 ( .A(u5__abc_81276_new_n3922_), .B(u5__abc_81276_new_n3734_), .Y(u5__abc_81276_new_n3923_));
OR2X2 OR2X2_4113 ( .A(u5__abc_81276_new_n3923_), .B(u5__abc_81276_new_n3915_), .Y(u5__abc_81276_new_n3924_));
OR2X2 OR2X2_4114 ( .A(u5__abc_81276_new_n3909_), .B(u5__abc_81276_new_n3924_), .Y(u5__abc_81276_new_n3925_));
OR2X2 OR2X2_4115 ( .A(u5__abc_81276_new_n3925_), .B(u5__abc_81276_new_n3908_), .Y(cs_le_d));
OR2X2 OR2X2_4116 ( .A(u5__abc_81276_new_n3210_), .B(u5__abc_81276_new_n3927_), .Y(u5__abc_81276_new_n3928_));
OR2X2 OR2X2_4117 ( .A(u5__abc_81276_new_n1368_), .B(u5__abc_81276_new_n1433_), .Y(u5__abc_81276_new_n3934_));
OR2X2 OR2X2_4118 ( .A(u5__abc_81276_new_n3933_), .B(u5__abc_81276_new_n3934_), .Y(u5__abc_81276_new_n3935_));
OR2X2 OR2X2_4119 ( .A(u5__abc_81276_new_n3935_), .B(u5__abc_81276_new_n3932_), .Y(u5__abc_81276_new_n3936_));
OR2X2 OR2X2_412 ( .A(u0__abc_76628_new_n1979_), .B(u0__abc_76628_new_n1980_), .Y(u0__abc_76628_new_n1981_));
OR2X2 OR2X2_4120 ( .A(u5__abc_81276_new_n3937_), .B(u5__abc_81276_new_n3639_), .Y(u5__abc_81276_new_n3938_));
OR2X2 OR2X2_4121 ( .A(u5__abc_81276_new_n3936_), .B(u5__abc_81276_new_n3938_), .Y(u5__abc_81276_new_n3939_));
OR2X2 OR2X2_4122 ( .A(u5__abc_81276_new_n3940_), .B(u5__abc_81276_new_n3941_), .Y(u5__abc_81276_new_n3942_));
OR2X2 OR2X2_4123 ( .A(u5__abc_81276_new_n3939_), .B(u5__abc_81276_new_n3942_), .Y(u5__abc_81276_new_n3943_));
OR2X2 OR2X2_4124 ( .A(u5__abc_81276_new_n3943_), .B(u5__abc_81276_new_n3931_), .Y(u5__abc_81276_new_n3944_));
OR2X2 OR2X2_4125 ( .A(u5__abc_81276_new_n3944_), .B(u5__abc_81276_new_n3930_), .Y(u5__abc_81276_new_n3945_));
OR2X2 OR2X2_4126 ( .A(u5__abc_81276_new_n3945_), .B(u5__abc_81276_new_n3929_), .Y(u5_mc_c_oe_d));
OR2X2 OR2X2_4127 ( .A(u5__abc_81276_new_n3954_), .B(u5__abc_81276_new_n1701_), .Y(u5__abc_81276_new_n3955_));
OR2X2 OR2X2_4128 ( .A(u5__abc_81276_new_n3953_), .B(u5__abc_81276_new_n3955_), .Y(bank_clr_all));
OR2X2 OR2X2_4129 ( .A(u5__abc_81276_new_n3963_), .B(u5__abc_81276_new_n1702_), .Y(bank_clr));
OR2X2 OR2X2_413 ( .A(u0__abc_76628_new_n1982_), .B(u0__abc_76628_new_n1983_), .Y(u0__abc_76628_new_n1984_));
OR2X2 OR2X2_4130 ( .A(u5__abc_81276_new_n1323_), .B(u5__abc_81276_new_n1296_), .Y(u5__abc_81276_new_n3976_));
OR2X2 OR2X2_4131 ( .A(u5__abc_81276_new_n3975_), .B(u5__abc_81276_new_n3977_), .Y(next_adr));
OR2X2 OR2X2_4132 ( .A(u5__abc_81276_new_n3982_), .B(u5__abc_81276_new_n3352_), .Y(row_sel));
OR2X2 OR2X2_4133 ( .A(u5__abc_81276_new_n3995_), .B(u5__abc_81276_new_n3238_), .Y(u5__abc_81276_new_n4003_));
OR2X2 OR2X2_4134 ( .A(u5__abc_81276_new_n1613_), .B(u5_kro), .Y(u5__abc_81276_new_n4004_));
OR2X2 OR2X2_4135 ( .A(u5__abc_81276_new_n4007_), .B(u5__abc_81276_new_n4004_), .Y(u5__abc_81276_new_n4008_));
OR2X2 OR2X2_4136 ( .A(u5__abc_81276_new_n1537_), .B(u5_ap_en), .Y(u5__abc_81276_new_n4010_));
OR2X2 OR2X2_4137 ( .A(u5__abc_81276_new_n4009_), .B(u5__abc_81276_new_n4014_), .Y(u5__abc_81276_new_n4015_));
OR2X2 OR2X2_4138 ( .A(u5__abc_81276_new_n4047_), .B(u5__abc_81276_new_n1536_), .Y(u5__abc_81276_new_n4048_));
OR2X2 OR2X2_4139 ( .A(u5__abc_81276_new_n4046_), .B(_auto_iopadmap_cc_368_execute_85453), .Y(u5__abc_81276_new_n4049_));
OR2X2 OR2X2_414 ( .A(u0__abc_76628_new_n1985_), .B(u0__abc_76628_new_n1986_), .Y(u0__abc_76628_new_n1987_));
OR2X2 OR2X2_4140 ( .A(u5__abc_81276_new_n4053_), .B(u5__abc_81276_new_n4054_), .Y(u5__abc_81276_new_n4055_));
OR2X2 OR2X2_4141 ( .A(u5__abc_81276_new_n4055_), .B(u5__abc_81276_new_n3940_), .Y(u5__abc_81276_new_n4056_));
OR2X2 OR2X2_4142 ( .A(u5__abc_81276_new_n4056_), .B(u5__abc_81276_new_n4052_), .Y(u5__abc_81276_new_n4057_));
OR2X2 OR2X2_4143 ( .A(u5__abc_81276_new_n4057_), .B(u5__abc_81276_new_n3930_), .Y(u5__abc_81276_new_n4058_));
OR2X2 OR2X2_4144 ( .A(u5__abc_81276_new_n4051_), .B(u5__abc_81276_new_n4058_), .Y(u5__abc_81276_new_n4059_));
OR2X2 OR2X2_4145 ( .A(u5__abc_81276_new_n4074_), .B(u5__abc_81276_new_n4075_), .Y(u5__abc_81276_new_n4076_));
OR2X2 OR2X2_4146 ( .A(u5__abc_81276_new_n4076_), .B(u5__abc_81276_new_n4073_), .Y(u5__abc_81276_new_n4077_));
OR2X2 OR2X2_4147 ( .A(u5__abc_81276_new_n4077_), .B(u5__abc_81276_new_n4072_), .Y(u5__abc_81276_new_n4078_));
OR2X2 OR2X2_4148 ( .A(u5__abc_81276_new_n4071_), .B(u5__abc_81276_new_n4078_), .Y(u5__abc_81276_new_n4079_));
OR2X2 OR2X2_4149 ( .A(u5__abc_81276_new_n4070_), .B(u5__abc_81276_new_n4080_), .Y(u5__0susp_sel_r_0_0_));
OR2X2 OR2X2_415 ( .A(u0__abc_76628_new_n1989_), .B(spec_req_cs_0_bF_buf4_), .Y(u0__abc_76628_new_n1990_));
OR2X2 OR2X2_4150 ( .A(u5__abc_81276_new_n1689_), .B(u5__abc_81276_new_n4084_), .Y(u5__0wb_cycle_0_0_));
OR2X2 OR2X2_4151 ( .A(u5__abc_81276_new_n1822_), .B(u1_wb_write_go), .Y(u5__abc_81276_new_n4086_));
OR2X2 OR2X2_4152 ( .A(u5__abc_81276_new_n4088_), .B(u5__abc_81276_new_n4087_), .Y(u5__abc_81276_new_n4089_));
OR2X2 OR2X2_4153 ( .A(u5__abc_81276_new_n4090_), .B(u5__abc_81276_new_n4091_), .Y(u5__0wr_cycle_0_0_));
OR2X2 OR2X2_4154 ( .A(u6__abc_85257_new_n139_), .B(u6__abc_85257_new_n134_), .Y(u6__abc_85257_new_n140_));
OR2X2 OR2X2_4155 ( .A(u6__abc_85257_new_n147_), .B(u6__abc_85257_new_n152_), .Y(u6__0wb_ack_o_0_0_));
OR2X2 OR2X2_4156 ( .A(u6__abc_85257_new_n145__bF_buf4), .B(rf_dout_0_), .Y(u6__abc_85257_new_n154_));
OR2X2 OR2X2_4157 ( .A(u6__abc_85257_new_n155__bF_buf4), .B(mem_dout_0_), .Y(u6__abc_85257_new_n156_));
OR2X2 OR2X2_4158 ( .A(u6__abc_85257_new_n145__bF_buf2), .B(rf_dout_1_), .Y(u6__abc_85257_new_n158_));
OR2X2 OR2X2_4159 ( .A(u6__abc_85257_new_n155__bF_buf3), .B(mem_dout_1_), .Y(u6__abc_85257_new_n159_));
OR2X2 OR2X2_416 ( .A(u0__abc_76628_new_n1988_), .B(u0__abc_76628_new_n1990_), .Y(u0__abc_76628_new_n1991_));
OR2X2 OR2X2_4160 ( .A(u6__abc_85257_new_n145__bF_buf1), .B(rf_dout_2_), .Y(u6__abc_85257_new_n161_));
OR2X2 OR2X2_4161 ( .A(u6__abc_85257_new_n155__bF_buf2), .B(mem_dout_2_), .Y(u6__abc_85257_new_n162_));
OR2X2 OR2X2_4162 ( .A(u6__abc_85257_new_n145__bF_buf0), .B(rf_dout_3_), .Y(u6__abc_85257_new_n164_));
OR2X2 OR2X2_4163 ( .A(u6__abc_85257_new_n155__bF_buf1), .B(mem_dout_3_), .Y(u6__abc_85257_new_n165_));
OR2X2 OR2X2_4164 ( .A(u6__abc_85257_new_n145__bF_buf5), .B(rf_dout_4_), .Y(u6__abc_85257_new_n167_));
OR2X2 OR2X2_4165 ( .A(u6__abc_85257_new_n155__bF_buf0), .B(mem_dout_4_), .Y(u6__abc_85257_new_n168_));
OR2X2 OR2X2_4166 ( .A(u6__abc_85257_new_n145__bF_buf4), .B(rf_dout_5_), .Y(u6__abc_85257_new_n170_));
OR2X2 OR2X2_4167 ( .A(u6__abc_85257_new_n155__bF_buf4), .B(mem_dout_5_), .Y(u6__abc_85257_new_n171_));
OR2X2 OR2X2_4168 ( .A(u6__abc_85257_new_n145__bF_buf3), .B(rf_dout_6_), .Y(u6__abc_85257_new_n173_));
OR2X2 OR2X2_4169 ( .A(u6__abc_85257_new_n155__bF_buf3), .B(mem_dout_6_), .Y(u6__abc_85257_new_n174_));
OR2X2 OR2X2_417 ( .A(u0__abc_76628_new_n1197__bF_buf1), .B(u0_csc0_1_), .Y(u0__abc_76628_new_n1992_));
OR2X2 OR2X2_4170 ( .A(u6__abc_85257_new_n145__bF_buf2), .B(rf_dout_7_), .Y(u6__abc_85257_new_n176_));
OR2X2 OR2X2_4171 ( .A(u6__abc_85257_new_n155__bF_buf2), .B(mem_dout_7_), .Y(u6__abc_85257_new_n177_));
OR2X2 OR2X2_4172 ( .A(u6__abc_85257_new_n145__bF_buf1), .B(rf_dout_8_), .Y(u6__abc_85257_new_n179_));
OR2X2 OR2X2_4173 ( .A(u6__abc_85257_new_n155__bF_buf1), .B(mem_dout_8_), .Y(u6__abc_85257_new_n180_));
OR2X2 OR2X2_4174 ( .A(u6__abc_85257_new_n145__bF_buf0), .B(rf_dout_9_), .Y(u6__abc_85257_new_n182_));
OR2X2 OR2X2_4175 ( .A(u6__abc_85257_new_n155__bF_buf0), .B(mem_dout_9_), .Y(u6__abc_85257_new_n183_));
OR2X2 OR2X2_4176 ( .A(u6__abc_85257_new_n145__bF_buf5), .B(rf_dout_10_), .Y(u6__abc_85257_new_n185_));
OR2X2 OR2X2_4177 ( .A(u6__abc_85257_new_n155__bF_buf4), .B(mem_dout_10_), .Y(u6__abc_85257_new_n186_));
OR2X2 OR2X2_4178 ( .A(u6__abc_85257_new_n145__bF_buf4), .B(rf_dout_11_), .Y(u6__abc_85257_new_n188_));
OR2X2 OR2X2_4179 ( .A(u6__abc_85257_new_n155__bF_buf3), .B(mem_dout_11_), .Y(u6__abc_85257_new_n189_));
OR2X2 OR2X2_418 ( .A(u0__abc_76628_new_n1994_), .B(u0__abc_76628_new_n1972_), .Y(u0__0sp_csc_31_0__1_));
OR2X2 OR2X2_4180 ( .A(u6__abc_85257_new_n145__bF_buf3), .B(rf_dout_12_), .Y(u6__abc_85257_new_n191_));
OR2X2 OR2X2_4181 ( .A(u6__abc_85257_new_n155__bF_buf2), .B(mem_dout_12_), .Y(u6__abc_85257_new_n192_));
OR2X2 OR2X2_4182 ( .A(u6__abc_85257_new_n145__bF_buf2), .B(rf_dout_13_), .Y(u6__abc_85257_new_n194_));
OR2X2 OR2X2_4183 ( .A(u6__abc_85257_new_n155__bF_buf1), .B(mem_dout_13_), .Y(u6__abc_85257_new_n195_));
OR2X2 OR2X2_4184 ( .A(u6__abc_85257_new_n145__bF_buf1), .B(rf_dout_14_), .Y(u6__abc_85257_new_n197_));
OR2X2 OR2X2_4185 ( .A(u6__abc_85257_new_n155__bF_buf0), .B(mem_dout_14_), .Y(u6__abc_85257_new_n198_));
OR2X2 OR2X2_4186 ( .A(u6__abc_85257_new_n145__bF_buf0), .B(rf_dout_15_), .Y(u6__abc_85257_new_n200_));
OR2X2 OR2X2_4187 ( .A(u6__abc_85257_new_n155__bF_buf4), .B(mem_dout_15_), .Y(u6__abc_85257_new_n201_));
OR2X2 OR2X2_4188 ( .A(u6__abc_85257_new_n145__bF_buf5), .B(rf_dout_16_), .Y(u6__abc_85257_new_n203_));
OR2X2 OR2X2_4189 ( .A(u6__abc_85257_new_n155__bF_buf3), .B(mem_dout_16_), .Y(u6__abc_85257_new_n204_));
OR2X2 OR2X2_419 ( .A(u0__abc_76628_new_n1177__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n1998_));
OR2X2 OR2X2_4190 ( .A(u6__abc_85257_new_n145__bF_buf4), .B(rf_dout_17_), .Y(u6__abc_85257_new_n206_));
OR2X2 OR2X2_4191 ( .A(u6__abc_85257_new_n155__bF_buf2), .B(mem_dout_17_), .Y(u6__abc_85257_new_n207_));
OR2X2 OR2X2_4192 ( .A(u6__abc_85257_new_n145__bF_buf3), .B(rf_dout_18_), .Y(u6__abc_85257_new_n209_));
OR2X2 OR2X2_4193 ( .A(u6__abc_85257_new_n155__bF_buf1), .B(mem_dout_18_), .Y(u6__abc_85257_new_n210_));
OR2X2 OR2X2_4194 ( .A(u6__abc_85257_new_n145__bF_buf2), .B(rf_dout_19_), .Y(u6__abc_85257_new_n212_));
OR2X2 OR2X2_4195 ( .A(u6__abc_85257_new_n155__bF_buf0), .B(mem_dout_19_), .Y(u6__abc_85257_new_n213_));
OR2X2 OR2X2_4196 ( .A(u6__abc_85257_new_n145__bF_buf1), .B(rf_dout_20_), .Y(u6__abc_85257_new_n215_));
OR2X2 OR2X2_4197 ( .A(u6__abc_85257_new_n155__bF_buf4), .B(mem_dout_20_), .Y(u6__abc_85257_new_n216_));
OR2X2 OR2X2_4198 ( .A(u6__abc_85257_new_n145__bF_buf0), .B(rf_dout_21_), .Y(u6__abc_85257_new_n218_));
OR2X2 OR2X2_4199 ( .A(u6__abc_85257_new_n155__bF_buf3), .B(mem_dout_21_), .Y(u6__abc_85257_new_n219_));
OR2X2 OR2X2_42 ( .A(lmr_sel_bF_buf2), .B(tms_3_), .Y(_abc_85006_new_n300_));
OR2X2 OR2X2_420 ( .A(spec_req_cs_6_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n1999_));
OR2X2 OR2X2_4200 ( .A(u6__abc_85257_new_n145__bF_buf5), .B(rf_dout_22_), .Y(u6__abc_85257_new_n221_));
OR2X2 OR2X2_4201 ( .A(u6__abc_85257_new_n155__bF_buf2), .B(mem_dout_22_), .Y(u6__abc_85257_new_n222_));
OR2X2 OR2X2_4202 ( .A(u6__abc_85257_new_n145__bF_buf4), .B(rf_dout_23_), .Y(u6__abc_85257_new_n224_));
OR2X2 OR2X2_4203 ( .A(u6__abc_85257_new_n155__bF_buf1), .B(mem_dout_23_), .Y(u6__abc_85257_new_n225_));
OR2X2 OR2X2_4204 ( .A(u6__abc_85257_new_n145__bF_buf3), .B(rf_dout_24_), .Y(u6__abc_85257_new_n227_));
OR2X2 OR2X2_4205 ( .A(u6__abc_85257_new_n155__bF_buf0), .B(mem_dout_24_), .Y(u6__abc_85257_new_n228_));
OR2X2 OR2X2_4206 ( .A(u6__abc_85257_new_n145__bF_buf2), .B(rf_dout_25_), .Y(u6__abc_85257_new_n230_));
OR2X2 OR2X2_4207 ( .A(u6__abc_85257_new_n155__bF_buf4), .B(mem_dout_25_), .Y(u6__abc_85257_new_n231_));
OR2X2 OR2X2_4208 ( .A(u6__abc_85257_new_n145__bF_buf1), .B(rf_dout_26_), .Y(u6__abc_85257_new_n233_));
OR2X2 OR2X2_4209 ( .A(u6__abc_85257_new_n155__bF_buf3), .B(mem_dout_26_), .Y(u6__abc_85257_new_n234_));
OR2X2 OR2X2_421 ( .A(u0__abc_76628_new_n2001_), .B(u0__abc_76628_new_n1997_), .Y(u0__abc_76628_new_n2002_));
OR2X2 OR2X2_4210 ( .A(u6__abc_85257_new_n145__bF_buf0), .B(rf_dout_27_), .Y(u6__abc_85257_new_n236_));
OR2X2 OR2X2_4211 ( .A(u6__abc_85257_new_n155__bF_buf2), .B(mem_dout_27_), .Y(u6__abc_85257_new_n237_));
OR2X2 OR2X2_4212 ( .A(u6__abc_85257_new_n145__bF_buf5), .B(rf_dout_28_), .Y(u6__abc_85257_new_n239_));
OR2X2 OR2X2_4213 ( .A(u6__abc_85257_new_n155__bF_buf1), .B(mem_dout_28_), .Y(u6__abc_85257_new_n240_));
OR2X2 OR2X2_4214 ( .A(u6__abc_85257_new_n145__bF_buf4), .B(rf_dout_29_), .Y(u6__abc_85257_new_n242_));
OR2X2 OR2X2_4215 ( .A(u6__abc_85257_new_n155__bF_buf0), .B(mem_dout_29_), .Y(u6__abc_85257_new_n243_));
OR2X2 OR2X2_4216 ( .A(u6__abc_85257_new_n145__bF_buf3), .B(rf_dout_30_), .Y(u6__abc_85257_new_n245_));
OR2X2 OR2X2_4217 ( .A(u6__abc_85257_new_n155__bF_buf4), .B(mem_dout_30_), .Y(u6__abc_85257_new_n246_));
OR2X2 OR2X2_4218 ( .A(u6__abc_85257_new_n145__bF_buf2), .B(rf_dout_31_), .Y(u6__abc_85257_new_n248_));
OR2X2 OR2X2_4219 ( .A(u6__abc_85257_new_n155__bF_buf3), .B(mem_dout_31_), .Y(u6__abc_85257_new_n249_));
OR2X2 OR2X2_422 ( .A(u0__abc_76628_new_n2003_), .B(u0__abc_76628_new_n2004_), .Y(u0__abc_76628_new_n2005_));
OR2X2 OR2X2_4220 ( .A(u6__abc_85257_new_n252_), .B(u6__abc_85257_new_n251_), .Y(u6__0wr_hold_0_0_));
OR2X2 OR2X2_4221 ( .A(u6__abc_85257_new_n259_), .B(u6_read_go_r), .Y(u6__abc_85257_new_n260_));
OR2X2 OR2X2_4222 ( .A(u6__abc_85257_new_n268_), .B(u6_write_go_r), .Y(u6__abc_85257_new_n269_));
OR2X2 OR2X2_4223 ( .A(u6__abc_85257_new_n271_), .B(wb_we_i), .Y(u6__abc_85257_new_n272_));
OR2X2 OR2X2_4224 ( .A(u6__abc_85257_new_n280_), .B(u6__abc_85257_new_n283_), .Y(u5_wb_first));
OR2X2 OR2X2_4225 ( .A(u3_wb_read_go), .B(u1_wb_write_go), .Y(u6__abc_85257_new_n288_));
OR2X2 OR2X2_4226 ( .A(u6__abc_85257_new_n291_), .B(_auto_iopadmap_cc_368_execute_85558), .Y(u6__0rmw_en_0_0_));
OR2X2 OR2X2_4227 ( .A(u6__abc_85257_new_n280_), .B(u6__abc_85257_new_n283_), .Y(u6__0wb_first_r_0_0_));
OR2X2 OR2X2_4228 ( .A(u7__abc_74830_new_n78_), .B(u1_wr_cycle), .Y(u7__abc_74830_new_n79_));
OR2X2 OR2X2_4229 ( .A(u7__abc_74830_new_n80_), .B(susp_sel), .Y(u7__abc_74830_new_n81_));
OR2X2 OR2X2_423 ( .A(u0__abc_76628_new_n2006_), .B(u0__abc_76628_new_n2007_), .Y(u0__abc_76628_new_n2008_));
OR2X2 OR2X2_4230 ( .A(u7__abc_74830_new_n81_), .B(u7__abc_74830_new_n76_), .Y(u7__0mc_dqm_3_0__0_));
OR2X2 OR2X2_4231 ( .A(u7__abc_74830_new_n81_), .B(u7__abc_74830_new_n84_), .Y(u7__0mc_dqm_3_0__1_));
OR2X2 OR2X2_4232 ( .A(u7__abc_74830_new_n81_), .B(u7__abc_74830_new_n87_), .Y(u7__0mc_dqm_3_0__2_));
OR2X2 OR2X2_4233 ( .A(u7__abc_74830_new_n81_), .B(u7__abc_74830_new_n90_), .Y(u7__0mc_dqm_3_0__3_));
OR2X2 OR2X2_4234 ( .A(u7__abc_74830_new_n95_), .B(u7__abc_74830_new_n93_), .Y(u7__0mc_dqm_r_3_0__0_));
OR2X2 OR2X2_4235 ( .A(u7__abc_74830_new_n98_), .B(u7__abc_74830_new_n97_), .Y(u7__0mc_dqm_r_3_0__1_));
OR2X2 OR2X2_4236 ( .A(u7__abc_74830_new_n101_), .B(u7__abc_74830_new_n100_), .Y(u7__0mc_dqm_r_3_0__2_));
OR2X2 OR2X2_4237 ( .A(u7__abc_74830_new_n104_), .B(u7__abc_74830_new_n103_), .Y(u7__0mc_dqm_r_3_0__3_));
OR2X2 OR2X2_4238 ( .A(susp_sel), .B(rfr_ack), .Y(u7__abc_74830_new_n106_));
OR2X2 OR2X2_4239 ( .A(u7__abc_74830_new_n108_), .B(lmr_sel_bF_buf2), .Y(u7__abc_74830_new_n109_));
OR2X2 OR2X2_424 ( .A(u0__abc_76628_new_n2009_), .B(u0__abc_76628_new_n2010_), .Y(u0__abc_76628_new_n2011_));
OR2X2 OR2X2_4240 ( .A(u7__abc_74830_new_n116_), .B(u7__abc_74830_new_n114_), .Y(u7__abc_74830_new_n117_));
OR2X2 OR2X2_4241 ( .A(u7__abc_74830_new_n113_), .B(u7__abc_74830_new_n117_), .Y(u7__0mc_cs__0_0_));
OR2X2 OR2X2_4242 ( .A(u7__abc_74830_new_n119_), .B(lmr_sel_bF_buf0), .Y(u7__abc_74830_new_n120_));
OR2X2 OR2X2_4243 ( .A(u7__abc_74830_new_n126_), .B(u7__abc_74830_new_n114_), .Y(u7__abc_74830_new_n127_));
OR2X2 OR2X2_4244 ( .A(u7__abc_74830_new_n124_), .B(u7__abc_74830_new_n127_), .Y(u7__0mc_cs__1_1_));
OR2X2 OR2X2_4245 ( .A(u7__abc_74830_new_n129_), .B(lmr_sel_bF_buf5), .Y(u7__abc_74830_new_n130_));
OR2X2 OR2X2_4246 ( .A(u7__abc_74830_new_n136_), .B(u7__abc_74830_new_n114_), .Y(u7__abc_74830_new_n137_));
OR2X2 OR2X2_4247 ( .A(u7__abc_74830_new_n134_), .B(u7__abc_74830_new_n137_), .Y(u7__0mc_cs__2_2_));
OR2X2 OR2X2_4248 ( .A(u7__abc_74830_new_n139_), .B(lmr_sel_bF_buf3), .Y(u7__abc_74830_new_n140_));
OR2X2 OR2X2_4249 ( .A(u7__abc_74830_new_n146_), .B(u7__abc_74830_new_n114_), .Y(u7__abc_74830_new_n147_));
OR2X2 OR2X2_425 ( .A(u0__abc_76628_new_n2013_), .B(spec_req_cs_0_bF_buf3_), .Y(u0__abc_76628_new_n2014_));
OR2X2 OR2X2_4250 ( .A(u7__abc_74830_new_n144_), .B(u7__abc_74830_new_n147_), .Y(u7__0mc_cs__3_3_));
OR2X2 OR2X2_4251 ( .A(u7__abc_74830_new_n149_), .B(lmr_sel_bF_buf1), .Y(u7__abc_74830_new_n150_));
OR2X2 OR2X2_4252 ( .A(u7__abc_74830_new_n156_), .B(u7__abc_74830_new_n114_), .Y(u7__abc_74830_new_n157_));
OR2X2 OR2X2_4253 ( .A(u7__abc_74830_new_n154_), .B(u7__abc_74830_new_n157_), .Y(u7__0mc_cs__4_4_));
OR2X2 OR2X2_4254 ( .A(u7__abc_74830_new_n159_), .B(lmr_sel_bF_buf6), .Y(u7__abc_74830_new_n160_));
OR2X2 OR2X2_4255 ( .A(u7__abc_74830_new_n166_), .B(u7__abc_74830_new_n114_), .Y(u7__abc_74830_new_n167_));
OR2X2 OR2X2_4256 ( .A(u7__abc_74830_new_n164_), .B(u7__abc_74830_new_n167_), .Y(u7__0mc_cs__5_5_));
OR2X2 OR2X2_4257 ( .A(u7__abc_74830_new_n169_), .B(lmr_sel_bF_buf4), .Y(u7__abc_74830_new_n170_));
OR2X2 OR2X2_4258 ( .A(u7__abc_74830_new_n176_), .B(u7__abc_74830_new_n114_), .Y(u7__abc_74830_new_n177_));
OR2X2 OR2X2_4259 ( .A(u7__abc_74830_new_n174_), .B(u7__abc_74830_new_n177_), .Y(u7__0mc_cs__6_6_));
OR2X2 OR2X2_426 ( .A(u0__abc_76628_new_n2012_), .B(u0__abc_76628_new_n2014_), .Y(u0__abc_76628_new_n2015_));
OR2X2 OR2X2_4260 ( .A(u7__abc_74830_new_n179_), .B(lmr_sel_bF_buf2), .Y(u7__abc_74830_new_n180_));
OR2X2 OR2X2_4261 ( .A(u7__abc_74830_new_n186_), .B(u7__abc_74830_new_n114_), .Y(u7__abc_74830_new_n187_));
OR2X2 OR2X2_4262 ( .A(u7__abc_74830_new_n184_), .B(u7__abc_74830_new_n187_), .Y(u7__0mc_cs__7_7_));
OR2X2 OR2X2_4263 ( .A(susp_sel), .B(oe_), .Y(u7__0mc_oe__0_0_));
OR2X2 OR2X2_427 ( .A(u0__abc_76628_new_n1197__bF_buf0), .B(u0_csc0_2_), .Y(u0__abc_76628_new_n2016_));
OR2X2 OR2X2_428 ( .A(u0__abc_76628_new_n2018_), .B(u0__abc_76628_new_n1996_), .Y(u0__0sp_csc_31_0__2_));
OR2X2 OR2X2_429 ( .A(u0__abc_76628_new_n1177__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n2022_));
OR2X2 OR2X2_43 ( .A(_abc_85006_new_n240__bF_buf5), .B(sp_tms_4_), .Y(_abc_85006_new_n302_));
OR2X2 OR2X2_430 ( .A(spec_req_cs_6_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n2023_));
OR2X2 OR2X2_431 ( .A(u0__abc_76628_new_n2025_), .B(u0__abc_76628_new_n2021_), .Y(u0__abc_76628_new_n2026_));
OR2X2 OR2X2_432 ( .A(u0__abc_76628_new_n2027_), .B(u0__abc_76628_new_n2028_), .Y(u0__abc_76628_new_n2029_));
OR2X2 OR2X2_433 ( .A(u0__abc_76628_new_n2030_), .B(u0__abc_76628_new_n2031_), .Y(u0__abc_76628_new_n2032_));
OR2X2 OR2X2_434 ( .A(u0__abc_76628_new_n2033_), .B(u0__abc_76628_new_n2034_), .Y(u0__abc_76628_new_n2035_));
OR2X2 OR2X2_435 ( .A(u0__abc_76628_new_n2037_), .B(spec_req_cs_0_bF_buf2_), .Y(u0__abc_76628_new_n2038_));
OR2X2 OR2X2_436 ( .A(u0__abc_76628_new_n2036_), .B(u0__abc_76628_new_n2038_), .Y(u0__abc_76628_new_n2039_));
OR2X2 OR2X2_437 ( .A(u0__abc_76628_new_n1197__bF_buf5), .B(u0_csc0_3_), .Y(u0__abc_76628_new_n2040_));
OR2X2 OR2X2_438 ( .A(u0__abc_76628_new_n2042_), .B(u0__abc_76628_new_n2020_), .Y(u0__0sp_csc_31_0__3_));
OR2X2 OR2X2_439 ( .A(u0__abc_76628_new_n1177__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n2046_));
OR2X2 OR2X2_44 ( .A(lmr_sel_bF_buf1), .B(tms_4_), .Y(_abc_85006_new_n303_));
OR2X2 OR2X2_440 ( .A(spec_req_cs_6_bF_buf1_), .B(1'h0), .Y(u0__abc_76628_new_n2047_));
OR2X2 OR2X2_441 ( .A(u0__abc_76628_new_n2049_), .B(u0__abc_76628_new_n2045_), .Y(u0__abc_76628_new_n2050_));
OR2X2 OR2X2_442 ( .A(u0__abc_76628_new_n2051_), .B(u0__abc_76628_new_n2052_), .Y(u0__abc_76628_new_n2053_));
OR2X2 OR2X2_443 ( .A(u0__abc_76628_new_n2054_), .B(u0__abc_76628_new_n2055_), .Y(u0__abc_76628_new_n2056_));
OR2X2 OR2X2_444 ( .A(u0__abc_76628_new_n2057_), .B(u0__abc_76628_new_n2058_), .Y(u0__abc_76628_new_n2059_));
OR2X2 OR2X2_445 ( .A(u0__abc_76628_new_n2061_), .B(spec_req_cs_0_bF_buf1_), .Y(u0__abc_76628_new_n2062_));
OR2X2 OR2X2_446 ( .A(u0__abc_76628_new_n2060_), .B(u0__abc_76628_new_n2062_), .Y(u0__abc_76628_new_n2063_));
OR2X2 OR2X2_447 ( .A(u0__abc_76628_new_n1197__bF_buf4), .B(u0_csc0_4_), .Y(u0__abc_76628_new_n2064_));
OR2X2 OR2X2_448 ( .A(u0__abc_76628_new_n2066_), .B(u0__abc_76628_new_n2044_), .Y(u0__0sp_csc_31_0__4_));
OR2X2 OR2X2_449 ( .A(u0__abc_76628_new_n1177__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n2070_));
OR2X2 OR2X2_45 ( .A(_abc_85006_new_n240__bF_buf4), .B(sp_tms_5_), .Y(_abc_85006_new_n305_));
OR2X2 OR2X2_450 ( .A(spec_req_cs_6_bF_buf0_), .B(1'h0), .Y(u0__abc_76628_new_n2071_));
OR2X2 OR2X2_451 ( .A(u0__abc_76628_new_n2073_), .B(u0__abc_76628_new_n2069_), .Y(u0__abc_76628_new_n2074_));
OR2X2 OR2X2_452 ( .A(u0__abc_76628_new_n2075_), .B(u0__abc_76628_new_n2076_), .Y(u0__abc_76628_new_n2077_));
OR2X2 OR2X2_453 ( .A(u0__abc_76628_new_n2078_), .B(u0__abc_76628_new_n2079_), .Y(u0__abc_76628_new_n2080_));
OR2X2 OR2X2_454 ( .A(u0__abc_76628_new_n2081_), .B(u0__abc_76628_new_n2082_), .Y(u0__abc_76628_new_n2083_));
OR2X2 OR2X2_455 ( .A(u0__abc_76628_new_n2085_), .B(spec_req_cs_0_bF_buf0_), .Y(u0__abc_76628_new_n2086_));
OR2X2 OR2X2_456 ( .A(u0__abc_76628_new_n2084_), .B(u0__abc_76628_new_n2086_), .Y(u0__abc_76628_new_n2087_));
OR2X2 OR2X2_457 ( .A(u0__abc_76628_new_n1197__bF_buf3), .B(u0_csc0_5_), .Y(u0__abc_76628_new_n2088_));
OR2X2 OR2X2_458 ( .A(u0__abc_76628_new_n2090_), .B(u0__abc_76628_new_n2068_), .Y(u0__0sp_csc_31_0__5_));
OR2X2 OR2X2_459 ( .A(u0__abc_76628_new_n1177__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n2094_));
OR2X2 OR2X2_46 ( .A(lmr_sel_bF_buf0), .B(tms_5_), .Y(_abc_85006_new_n306_));
OR2X2 OR2X2_460 ( .A(spec_req_cs_6_bF_buf5_), .B(1'h0), .Y(u0__abc_76628_new_n2095_));
OR2X2 OR2X2_461 ( .A(u0__abc_76628_new_n2097_), .B(u0__abc_76628_new_n2093_), .Y(u0__abc_76628_new_n2098_));
OR2X2 OR2X2_462 ( .A(u0__abc_76628_new_n2099_), .B(u0__abc_76628_new_n2100_), .Y(u0__abc_76628_new_n2101_));
OR2X2 OR2X2_463 ( .A(u0__abc_76628_new_n2102_), .B(u0__abc_76628_new_n2103_), .Y(u0__abc_76628_new_n2104_));
OR2X2 OR2X2_464 ( .A(u0__abc_76628_new_n2105_), .B(u0__abc_76628_new_n2106_), .Y(u0__abc_76628_new_n2107_));
OR2X2 OR2X2_465 ( .A(u0__abc_76628_new_n2109_), .B(spec_req_cs_0_bF_buf5_), .Y(u0__abc_76628_new_n2110_));
OR2X2 OR2X2_466 ( .A(u0__abc_76628_new_n2108_), .B(u0__abc_76628_new_n2110_), .Y(u0__abc_76628_new_n2111_));
OR2X2 OR2X2_467 ( .A(u0__abc_76628_new_n1197__bF_buf2), .B(u0_csc0_6_), .Y(u0__abc_76628_new_n2112_));
OR2X2 OR2X2_468 ( .A(u0__abc_76628_new_n2114_), .B(u0__abc_76628_new_n2092_), .Y(u0__0sp_csc_31_0__6_));
OR2X2 OR2X2_469 ( .A(u0__abc_76628_new_n1177__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n2118_));
OR2X2 OR2X2_47 ( .A(_abc_85006_new_n240__bF_buf3), .B(sp_tms_6_), .Y(_abc_85006_new_n308_));
OR2X2 OR2X2_470 ( .A(spec_req_cs_6_bF_buf4_), .B(1'h0), .Y(u0__abc_76628_new_n2119_));
OR2X2 OR2X2_471 ( .A(u0__abc_76628_new_n2121_), .B(u0__abc_76628_new_n2117_), .Y(u0__abc_76628_new_n2122_));
OR2X2 OR2X2_472 ( .A(u0__abc_76628_new_n2123_), .B(u0__abc_76628_new_n2124_), .Y(u0__abc_76628_new_n2125_));
OR2X2 OR2X2_473 ( .A(u0__abc_76628_new_n2126_), .B(u0__abc_76628_new_n2127_), .Y(u0__abc_76628_new_n2128_));
OR2X2 OR2X2_474 ( .A(u0__abc_76628_new_n2129_), .B(u0__abc_76628_new_n2130_), .Y(u0__abc_76628_new_n2131_));
OR2X2 OR2X2_475 ( .A(u0__abc_76628_new_n2133_), .B(spec_req_cs_0_bF_buf4_), .Y(u0__abc_76628_new_n2134_));
OR2X2 OR2X2_476 ( .A(u0__abc_76628_new_n2132_), .B(u0__abc_76628_new_n2134_), .Y(u0__abc_76628_new_n2135_));
OR2X2 OR2X2_477 ( .A(u0__abc_76628_new_n1197__bF_buf1), .B(u0_csc0_7_), .Y(u0__abc_76628_new_n2136_));
OR2X2 OR2X2_478 ( .A(u0__abc_76628_new_n2138_), .B(u0__abc_76628_new_n2116_), .Y(u0__0sp_csc_31_0__7_));
OR2X2 OR2X2_479 ( .A(u0__abc_76628_new_n1177__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n2166_));
OR2X2 OR2X2_48 ( .A(lmr_sel_bF_buf6), .B(tms_6_), .Y(_abc_85006_new_n309_));
OR2X2 OR2X2_480 ( .A(spec_req_cs_6_bF_buf3_), .B(1'h0), .Y(u0__abc_76628_new_n2167_));
OR2X2 OR2X2_481 ( .A(u0__abc_76628_new_n2169_), .B(u0__abc_76628_new_n2165_), .Y(u0__abc_76628_new_n2170_));
OR2X2 OR2X2_482 ( .A(u0__abc_76628_new_n2171_), .B(u0__abc_76628_new_n2172_), .Y(u0__abc_76628_new_n2173_));
OR2X2 OR2X2_483 ( .A(u0__abc_76628_new_n2174_), .B(u0__abc_76628_new_n2175_), .Y(u0__abc_76628_new_n2176_));
OR2X2 OR2X2_484 ( .A(u0__abc_76628_new_n2177_), .B(u0__abc_76628_new_n2178_), .Y(u0__abc_76628_new_n2179_));
OR2X2 OR2X2_485 ( .A(u0__abc_76628_new_n2181_), .B(spec_req_cs_0_bF_buf3_), .Y(u0__abc_76628_new_n2182_));
OR2X2 OR2X2_486 ( .A(u0__abc_76628_new_n2180_), .B(u0__abc_76628_new_n2182_), .Y(u0__abc_76628_new_n2183_));
OR2X2 OR2X2_487 ( .A(u0__abc_76628_new_n1197__bF_buf0), .B(u0_csc0_9_), .Y(u0__abc_76628_new_n2184_));
OR2X2 OR2X2_488 ( .A(u0__abc_76628_new_n2186_), .B(u0__abc_76628_new_n2164_), .Y(u0__0sp_csc_31_0__9_));
OR2X2 OR2X2_489 ( .A(u0__abc_76628_new_n1177__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n2190_));
OR2X2 OR2X2_49 ( .A(_abc_85006_new_n240__bF_buf2), .B(sp_tms_7_), .Y(_abc_85006_new_n311_));
OR2X2 OR2X2_490 ( .A(spec_req_cs_6_bF_buf2_), .B(1'h0), .Y(u0__abc_76628_new_n2191_));
OR2X2 OR2X2_491 ( .A(u0__abc_76628_new_n2193_), .B(u0__abc_76628_new_n2189_), .Y(u0__abc_76628_new_n2194_));
OR2X2 OR2X2_492 ( .A(u0__abc_76628_new_n2195_), .B(u0__abc_76628_new_n2196_), .Y(u0__abc_76628_new_n2197_));
OR2X2 OR2X2_493 ( .A(u0__abc_76628_new_n2198_), .B(u0__abc_76628_new_n2199_), .Y(u0__abc_76628_new_n2200_));
OR2X2 OR2X2_494 ( .A(u0__abc_76628_new_n2201_), .B(u0__abc_76628_new_n2202_), .Y(u0__abc_76628_new_n2203_));
OR2X2 OR2X2_495 ( .A(u0__abc_76628_new_n2205_), .B(spec_req_cs_0_bF_buf2_), .Y(u0__abc_76628_new_n2206_));
OR2X2 OR2X2_496 ( .A(u0__abc_76628_new_n2204_), .B(u0__abc_76628_new_n2206_), .Y(u0__abc_76628_new_n2207_));
OR2X2 OR2X2_497 ( .A(u0__abc_76628_new_n1197__bF_buf5), .B(u0_csc0_10_), .Y(u0__abc_76628_new_n2208_));
OR2X2 OR2X2_498 ( .A(u0__abc_76628_new_n2210_), .B(u0__abc_76628_new_n2188_), .Y(u0__0sp_csc_31_0__10_));
OR2X2 OR2X2_499 ( .A(u0__abc_76628_new_n2722__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n2723_));
OR2X2 OR2X2_5 ( .A(_abc_85006_new_n243_), .B(_abc_85006_new_n237_), .Y(_abc_85006_new_n244_));
OR2X2 OR2X2_50 ( .A(lmr_sel_bF_buf5), .B(tms_7_), .Y(_abc_85006_new_n312_));
OR2X2 OR2X2_500 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2725_));
OR2X2 OR2X2_501 ( .A(u0__abc_76628_new_n2727_), .B(u0__abc_76628_new_n2721_), .Y(u0__abc_76628_new_n2728_));
OR2X2 OR2X2_502 ( .A(u0__abc_76628_new_n2729_), .B(u0__abc_76628_new_n2730_), .Y(u0__abc_76628_new_n2731_));
OR2X2 OR2X2_503 ( .A(u0__abc_76628_new_n2732_), .B(u0__abc_76628_new_n2733_), .Y(u0__abc_76628_new_n2734_));
OR2X2 OR2X2_504 ( .A(u0__abc_76628_new_n2735_), .B(u0__abc_76628_new_n2736_), .Y(u0__abc_76628_new_n2737_));
OR2X2 OR2X2_505 ( .A(u0__abc_76628_new_n2739_), .B(u0_cs0_bF_buf5), .Y(u0__abc_76628_new_n2740_));
OR2X2 OR2X2_506 ( .A(u0__abc_76628_new_n2738_), .B(u0__abc_76628_new_n2740_), .Y(u0__abc_76628_new_n2741_));
OR2X2 OR2X2_507 ( .A(u0__abc_76628_new_n2742__bF_buf5), .B(u0_tms0_0_), .Y(u0__abc_76628_new_n2743_));
OR2X2 OR2X2_508 ( .A(u0__abc_76628_new_n2745_), .B(u0__abc_76628_new_n2716_), .Y(u0__0tms_31_0__0_));
OR2X2 OR2X2_509 ( .A(u0__abc_76628_new_n2722__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n2749_));
OR2X2 OR2X2_51 ( .A(_abc_85006_new_n240__bF_buf1), .B(sp_tms_8_), .Y(_abc_85006_new_n314_));
OR2X2 OR2X2_510 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2750_));
OR2X2 OR2X2_511 ( .A(u0__abc_76628_new_n2752_), .B(u0__abc_76628_new_n2748_), .Y(u0__abc_76628_new_n2753_));
OR2X2 OR2X2_512 ( .A(u0__abc_76628_new_n2754_), .B(u0__abc_76628_new_n2755_), .Y(u0__abc_76628_new_n2756_));
OR2X2 OR2X2_513 ( .A(u0__abc_76628_new_n2757_), .B(u0__abc_76628_new_n2758_), .Y(u0__abc_76628_new_n2759_));
OR2X2 OR2X2_514 ( .A(u0__abc_76628_new_n2760_), .B(u0__abc_76628_new_n2761_), .Y(u0__abc_76628_new_n2762_));
OR2X2 OR2X2_515 ( .A(u0__abc_76628_new_n2764_), .B(u0_cs0_bF_buf3), .Y(u0__abc_76628_new_n2765_));
OR2X2 OR2X2_516 ( .A(u0__abc_76628_new_n2763_), .B(u0__abc_76628_new_n2765_), .Y(u0__abc_76628_new_n2766_));
OR2X2 OR2X2_517 ( .A(u0__abc_76628_new_n2742__bF_buf4), .B(u0_tms0_1_), .Y(u0__abc_76628_new_n2767_));
OR2X2 OR2X2_518 ( .A(u0__abc_76628_new_n2769_), .B(u0__abc_76628_new_n2747_), .Y(u0__0tms_31_0__1_));
OR2X2 OR2X2_519 ( .A(u0__abc_76628_new_n2722__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n2773_));
OR2X2 OR2X2_52 ( .A(lmr_sel_bF_buf4), .B(tms_8_), .Y(_abc_85006_new_n315_));
OR2X2 OR2X2_520 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2774_));
OR2X2 OR2X2_521 ( .A(u0__abc_76628_new_n2776_), .B(u0__abc_76628_new_n2772_), .Y(u0__abc_76628_new_n2777_));
OR2X2 OR2X2_522 ( .A(u0__abc_76628_new_n2778_), .B(u0__abc_76628_new_n2779_), .Y(u0__abc_76628_new_n2780_));
OR2X2 OR2X2_523 ( .A(u0__abc_76628_new_n2781_), .B(u0__abc_76628_new_n2782_), .Y(u0__abc_76628_new_n2783_));
OR2X2 OR2X2_524 ( .A(u0__abc_76628_new_n2784_), .B(u0__abc_76628_new_n2785_), .Y(u0__abc_76628_new_n2786_));
OR2X2 OR2X2_525 ( .A(u0__abc_76628_new_n2788_), .B(u0_cs0_bF_buf2), .Y(u0__abc_76628_new_n2789_));
OR2X2 OR2X2_526 ( .A(u0__abc_76628_new_n2787_), .B(u0__abc_76628_new_n2789_), .Y(u0__abc_76628_new_n2790_));
OR2X2 OR2X2_527 ( .A(u0__abc_76628_new_n2742__bF_buf3), .B(u0_tms0_2_), .Y(u0__abc_76628_new_n2791_));
OR2X2 OR2X2_528 ( .A(u0__abc_76628_new_n2793_), .B(u0__abc_76628_new_n2771_), .Y(u0__0tms_31_0__2_));
OR2X2 OR2X2_529 ( .A(u0__abc_76628_new_n2722__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n2797_));
OR2X2 OR2X2_53 ( .A(_abc_85006_new_n240__bF_buf0), .B(sp_tms_9_), .Y(_abc_85006_new_n317_));
OR2X2 OR2X2_530 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2798_));
OR2X2 OR2X2_531 ( .A(u0__abc_76628_new_n2800_), .B(u0__abc_76628_new_n2796_), .Y(u0__abc_76628_new_n2801_));
OR2X2 OR2X2_532 ( .A(u0__abc_76628_new_n2802_), .B(u0__abc_76628_new_n2803_), .Y(u0__abc_76628_new_n2804_));
OR2X2 OR2X2_533 ( .A(u0__abc_76628_new_n2805_), .B(u0__abc_76628_new_n2806_), .Y(u0__abc_76628_new_n2807_));
OR2X2 OR2X2_534 ( .A(u0__abc_76628_new_n2808_), .B(u0__abc_76628_new_n2809_), .Y(u0__abc_76628_new_n2810_));
OR2X2 OR2X2_535 ( .A(u0__abc_76628_new_n2812_), .B(u0_cs0_bF_buf1), .Y(u0__abc_76628_new_n2813_));
OR2X2 OR2X2_536 ( .A(u0__abc_76628_new_n2811_), .B(u0__abc_76628_new_n2813_), .Y(u0__abc_76628_new_n2814_));
OR2X2 OR2X2_537 ( .A(u0__abc_76628_new_n2742__bF_buf2), .B(u0_tms0_3_), .Y(u0__abc_76628_new_n2815_));
OR2X2 OR2X2_538 ( .A(u0__abc_76628_new_n2817_), .B(u0__abc_76628_new_n2795_), .Y(u0__0tms_31_0__3_));
OR2X2 OR2X2_539 ( .A(u0__abc_76628_new_n2722__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n2821_));
OR2X2 OR2X2_54 ( .A(lmr_sel_bF_buf3), .B(tms_9_), .Y(_abc_85006_new_n318_));
OR2X2 OR2X2_540 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2822_));
OR2X2 OR2X2_541 ( .A(u0__abc_76628_new_n2824_), .B(u0__abc_76628_new_n2820_), .Y(u0__abc_76628_new_n2825_));
OR2X2 OR2X2_542 ( .A(u0__abc_76628_new_n2826_), .B(u0__abc_76628_new_n2827_), .Y(u0__abc_76628_new_n2828_));
OR2X2 OR2X2_543 ( .A(u0__abc_76628_new_n2829_), .B(u0__abc_76628_new_n2830_), .Y(u0__abc_76628_new_n2831_));
OR2X2 OR2X2_544 ( .A(u0__abc_76628_new_n2832_), .B(u0__abc_76628_new_n2833_), .Y(u0__abc_76628_new_n2834_));
OR2X2 OR2X2_545 ( .A(u0__abc_76628_new_n2836_), .B(u0_cs0_bF_buf0), .Y(u0__abc_76628_new_n2837_));
OR2X2 OR2X2_546 ( .A(u0__abc_76628_new_n2835_), .B(u0__abc_76628_new_n2837_), .Y(u0__abc_76628_new_n2838_));
OR2X2 OR2X2_547 ( .A(u0__abc_76628_new_n2742__bF_buf1), .B(u0_tms0_4_), .Y(u0__abc_76628_new_n2839_));
OR2X2 OR2X2_548 ( .A(u0__abc_76628_new_n2841_), .B(u0__abc_76628_new_n2819_), .Y(u0__0tms_31_0__4_));
OR2X2 OR2X2_549 ( .A(u0__abc_76628_new_n2722__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n2845_));
OR2X2 OR2X2_55 ( .A(_abc_85006_new_n240__bF_buf5), .B(sp_tms_10_), .Y(_abc_85006_new_n320_));
OR2X2 OR2X2_550 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2846_));
OR2X2 OR2X2_551 ( .A(u0__abc_76628_new_n2848_), .B(u0__abc_76628_new_n2844_), .Y(u0__abc_76628_new_n2849_));
OR2X2 OR2X2_552 ( .A(u0__abc_76628_new_n2850_), .B(u0__abc_76628_new_n2851_), .Y(u0__abc_76628_new_n2852_));
OR2X2 OR2X2_553 ( .A(u0__abc_76628_new_n2853_), .B(u0__abc_76628_new_n2854_), .Y(u0__abc_76628_new_n2855_));
OR2X2 OR2X2_554 ( .A(u0__abc_76628_new_n2856_), .B(u0__abc_76628_new_n2857_), .Y(u0__abc_76628_new_n2858_));
OR2X2 OR2X2_555 ( .A(u0__abc_76628_new_n2860_), .B(u0_cs0_bF_buf5), .Y(u0__abc_76628_new_n2861_));
OR2X2 OR2X2_556 ( .A(u0__abc_76628_new_n2859_), .B(u0__abc_76628_new_n2861_), .Y(u0__abc_76628_new_n2862_));
OR2X2 OR2X2_557 ( .A(u0__abc_76628_new_n2742__bF_buf0), .B(u0_tms0_5_), .Y(u0__abc_76628_new_n2863_));
OR2X2 OR2X2_558 ( .A(u0__abc_76628_new_n2865_), .B(u0__abc_76628_new_n2843_), .Y(u0__0tms_31_0__5_));
OR2X2 OR2X2_559 ( .A(u0__abc_76628_new_n2722__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n2869_));
OR2X2 OR2X2_56 ( .A(lmr_sel_bF_buf2), .B(tms_10_), .Y(_abc_85006_new_n321_));
OR2X2 OR2X2_560 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2870_));
OR2X2 OR2X2_561 ( .A(u0__abc_76628_new_n2872_), .B(u0__abc_76628_new_n2868_), .Y(u0__abc_76628_new_n2873_));
OR2X2 OR2X2_562 ( .A(u0__abc_76628_new_n2874_), .B(u0__abc_76628_new_n2875_), .Y(u0__abc_76628_new_n2876_));
OR2X2 OR2X2_563 ( .A(u0__abc_76628_new_n2877_), .B(u0__abc_76628_new_n2878_), .Y(u0__abc_76628_new_n2879_));
OR2X2 OR2X2_564 ( .A(u0__abc_76628_new_n2880_), .B(u0__abc_76628_new_n2881_), .Y(u0__abc_76628_new_n2882_));
OR2X2 OR2X2_565 ( .A(u0__abc_76628_new_n2884_), .B(u0_cs0_bF_buf4), .Y(u0__abc_76628_new_n2885_));
OR2X2 OR2X2_566 ( .A(u0__abc_76628_new_n2883_), .B(u0__abc_76628_new_n2885_), .Y(u0__abc_76628_new_n2886_));
OR2X2 OR2X2_567 ( .A(u0__abc_76628_new_n2742__bF_buf5), .B(u0_tms0_6_), .Y(u0__abc_76628_new_n2887_));
OR2X2 OR2X2_568 ( .A(u0__abc_76628_new_n2889_), .B(u0__abc_76628_new_n2867_), .Y(u0__0tms_31_0__6_));
OR2X2 OR2X2_569 ( .A(u0__abc_76628_new_n2722__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n2893_));
OR2X2 OR2X2_57 ( .A(_abc_85006_new_n240__bF_buf4), .B(sp_tms_11_), .Y(_abc_85006_new_n323_));
OR2X2 OR2X2_570 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2894_));
OR2X2 OR2X2_571 ( .A(u0__abc_76628_new_n2896_), .B(u0__abc_76628_new_n2892_), .Y(u0__abc_76628_new_n2897_));
OR2X2 OR2X2_572 ( .A(u0__abc_76628_new_n2898_), .B(u0__abc_76628_new_n2899_), .Y(u0__abc_76628_new_n2900_));
OR2X2 OR2X2_573 ( .A(u0__abc_76628_new_n2901_), .B(u0__abc_76628_new_n2902_), .Y(u0__abc_76628_new_n2903_));
OR2X2 OR2X2_574 ( .A(u0__abc_76628_new_n2904_), .B(u0__abc_76628_new_n2905_), .Y(u0__abc_76628_new_n2906_));
OR2X2 OR2X2_575 ( .A(u0__abc_76628_new_n2908_), .B(u0_cs0_bF_buf3), .Y(u0__abc_76628_new_n2909_));
OR2X2 OR2X2_576 ( .A(u0__abc_76628_new_n2907_), .B(u0__abc_76628_new_n2909_), .Y(u0__abc_76628_new_n2910_));
OR2X2 OR2X2_577 ( .A(u0__abc_76628_new_n2742__bF_buf4), .B(u0_tms0_7_), .Y(u0__abc_76628_new_n2911_));
OR2X2 OR2X2_578 ( .A(u0__abc_76628_new_n2913_), .B(u0__abc_76628_new_n2891_), .Y(u0__0tms_31_0__7_));
OR2X2 OR2X2_579 ( .A(u0__abc_76628_new_n2722__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n2917_));
OR2X2 OR2X2_58 ( .A(lmr_sel_bF_buf1), .B(tms_11_), .Y(_abc_85006_new_n324_));
OR2X2 OR2X2_580 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2918_));
OR2X2 OR2X2_581 ( .A(u0__abc_76628_new_n2920_), .B(u0__abc_76628_new_n2916_), .Y(u0__abc_76628_new_n2921_));
OR2X2 OR2X2_582 ( .A(u0__abc_76628_new_n2922_), .B(u0__abc_76628_new_n2923_), .Y(u0__abc_76628_new_n2924_));
OR2X2 OR2X2_583 ( .A(u0__abc_76628_new_n2925_), .B(u0__abc_76628_new_n2926_), .Y(u0__abc_76628_new_n2927_));
OR2X2 OR2X2_584 ( .A(u0__abc_76628_new_n2928_), .B(u0__abc_76628_new_n2929_), .Y(u0__abc_76628_new_n2930_));
OR2X2 OR2X2_585 ( .A(u0__abc_76628_new_n2932_), .B(u0_cs0_bF_buf2), .Y(u0__abc_76628_new_n2933_));
OR2X2 OR2X2_586 ( .A(u0__abc_76628_new_n2931_), .B(u0__abc_76628_new_n2933_), .Y(u0__abc_76628_new_n2934_));
OR2X2 OR2X2_587 ( .A(u0__abc_76628_new_n2742__bF_buf3), .B(u0_tms0_8_), .Y(u0__abc_76628_new_n2935_));
OR2X2 OR2X2_588 ( .A(u0__abc_76628_new_n2937_), .B(u0__abc_76628_new_n2915_), .Y(u0__0tms_31_0__8_));
OR2X2 OR2X2_589 ( .A(u0__abc_76628_new_n2722__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n2941_));
OR2X2 OR2X2_59 ( .A(_abc_85006_new_n240__bF_buf3), .B(sp_tms_12_), .Y(_abc_85006_new_n326_));
OR2X2 OR2X2_590 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2942_));
OR2X2 OR2X2_591 ( .A(u0__abc_76628_new_n2944_), .B(u0__abc_76628_new_n2940_), .Y(u0__abc_76628_new_n2945_));
OR2X2 OR2X2_592 ( .A(u0__abc_76628_new_n2946_), .B(u0__abc_76628_new_n2947_), .Y(u0__abc_76628_new_n2948_));
OR2X2 OR2X2_593 ( .A(u0__abc_76628_new_n2949_), .B(u0__abc_76628_new_n2950_), .Y(u0__abc_76628_new_n2951_));
OR2X2 OR2X2_594 ( .A(u0__abc_76628_new_n2952_), .B(u0__abc_76628_new_n2953_), .Y(u0__abc_76628_new_n2954_));
OR2X2 OR2X2_595 ( .A(u0__abc_76628_new_n2956_), .B(u0_cs0_bF_buf1), .Y(u0__abc_76628_new_n2957_));
OR2X2 OR2X2_596 ( .A(u0__abc_76628_new_n2955_), .B(u0__abc_76628_new_n2957_), .Y(u0__abc_76628_new_n2958_));
OR2X2 OR2X2_597 ( .A(u0__abc_76628_new_n2742__bF_buf2), .B(u0_tms0_9_), .Y(u0__abc_76628_new_n2959_));
OR2X2 OR2X2_598 ( .A(u0__abc_76628_new_n2961_), .B(u0__abc_76628_new_n2939_), .Y(u0__0tms_31_0__9_));
OR2X2 OR2X2_599 ( .A(u0__abc_76628_new_n2722__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n2965_));
OR2X2 OR2X2_6 ( .A(_abc_85006_new_n245_), .B(cs_need_rfr_0_), .Y(_abc_85006_new_n246_));
OR2X2 OR2X2_60 ( .A(lmr_sel_bF_buf0), .B(tms_12_), .Y(_abc_85006_new_n327_));
OR2X2 OR2X2_600 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2966_));
OR2X2 OR2X2_601 ( .A(u0__abc_76628_new_n2968_), .B(u0__abc_76628_new_n2964_), .Y(u0__abc_76628_new_n2969_));
OR2X2 OR2X2_602 ( .A(u0__abc_76628_new_n2970_), .B(u0__abc_76628_new_n2971_), .Y(u0__abc_76628_new_n2972_));
OR2X2 OR2X2_603 ( .A(u0__abc_76628_new_n2973_), .B(u0__abc_76628_new_n2974_), .Y(u0__abc_76628_new_n2975_));
OR2X2 OR2X2_604 ( .A(u0__abc_76628_new_n2976_), .B(u0__abc_76628_new_n2977_), .Y(u0__abc_76628_new_n2978_));
OR2X2 OR2X2_605 ( .A(u0__abc_76628_new_n2980_), .B(u0_cs0_bF_buf0), .Y(u0__abc_76628_new_n2981_));
OR2X2 OR2X2_606 ( .A(u0__abc_76628_new_n2979_), .B(u0__abc_76628_new_n2981_), .Y(u0__abc_76628_new_n2982_));
OR2X2 OR2X2_607 ( .A(u0__abc_76628_new_n2742__bF_buf1), .B(u0_tms0_10_), .Y(u0__abc_76628_new_n2983_));
OR2X2 OR2X2_608 ( .A(u0__abc_76628_new_n2985_), .B(u0__abc_76628_new_n2963_), .Y(u0__0tms_31_0__10_));
OR2X2 OR2X2_609 ( .A(u0__abc_76628_new_n2722__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n2989_));
OR2X2 OR2X2_61 ( .A(_abc_85006_new_n240__bF_buf2), .B(sp_tms_13_), .Y(_abc_85006_new_n329_));
OR2X2 OR2X2_610 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n2990_));
OR2X2 OR2X2_611 ( .A(u0__abc_76628_new_n2992_), .B(u0__abc_76628_new_n2988_), .Y(u0__abc_76628_new_n2993_));
OR2X2 OR2X2_612 ( .A(u0__abc_76628_new_n2994_), .B(u0__abc_76628_new_n2995_), .Y(u0__abc_76628_new_n2996_));
OR2X2 OR2X2_613 ( .A(u0__abc_76628_new_n2997_), .B(u0__abc_76628_new_n2998_), .Y(u0__abc_76628_new_n2999_));
OR2X2 OR2X2_614 ( .A(u0__abc_76628_new_n3000_), .B(u0__abc_76628_new_n3001_), .Y(u0__abc_76628_new_n3002_));
OR2X2 OR2X2_615 ( .A(u0__abc_76628_new_n3004_), .B(u0_cs0_bF_buf5), .Y(u0__abc_76628_new_n3005_));
OR2X2 OR2X2_616 ( .A(u0__abc_76628_new_n3003_), .B(u0__abc_76628_new_n3005_), .Y(u0__abc_76628_new_n3006_));
OR2X2 OR2X2_617 ( .A(u0__abc_76628_new_n2742__bF_buf0), .B(u0_tms0_11_), .Y(u0__abc_76628_new_n3007_));
OR2X2 OR2X2_618 ( .A(u0__abc_76628_new_n3009_), .B(u0__abc_76628_new_n2987_), .Y(u0__0tms_31_0__11_));
OR2X2 OR2X2_619 ( .A(u0__abc_76628_new_n2722__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n3013_));
OR2X2 OR2X2_62 ( .A(lmr_sel_bF_buf6), .B(tms_13_), .Y(_abc_85006_new_n330_));
OR2X2 OR2X2_620 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3014_));
OR2X2 OR2X2_621 ( .A(u0__abc_76628_new_n3016_), .B(u0__abc_76628_new_n3012_), .Y(u0__abc_76628_new_n3017_));
OR2X2 OR2X2_622 ( .A(u0__abc_76628_new_n3018_), .B(u0__abc_76628_new_n3019_), .Y(u0__abc_76628_new_n3020_));
OR2X2 OR2X2_623 ( .A(u0__abc_76628_new_n3021_), .B(u0__abc_76628_new_n3022_), .Y(u0__abc_76628_new_n3023_));
OR2X2 OR2X2_624 ( .A(u0__abc_76628_new_n3024_), .B(u0__abc_76628_new_n3025_), .Y(u0__abc_76628_new_n3026_));
OR2X2 OR2X2_625 ( .A(u0__abc_76628_new_n3028_), .B(u0_cs0_bF_buf4), .Y(u0__abc_76628_new_n3029_));
OR2X2 OR2X2_626 ( .A(u0__abc_76628_new_n3027_), .B(u0__abc_76628_new_n3029_), .Y(u0__abc_76628_new_n3030_));
OR2X2 OR2X2_627 ( .A(u0__abc_76628_new_n2742__bF_buf5), .B(u0_tms0_12_), .Y(u0__abc_76628_new_n3031_));
OR2X2 OR2X2_628 ( .A(u0__abc_76628_new_n3033_), .B(u0__abc_76628_new_n3011_), .Y(u0__0tms_31_0__12_));
OR2X2 OR2X2_629 ( .A(u0__abc_76628_new_n2722__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n3037_));
OR2X2 OR2X2_63 ( .A(_abc_85006_new_n240__bF_buf1), .B(sp_tms_14_), .Y(_abc_85006_new_n332_));
OR2X2 OR2X2_630 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3038_));
OR2X2 OR2X2_631 ( .A(u0__abc_76628_new_n3040_), .B(u0__abc_76628_new_n3036_), .Y(u0__abc_76628_new_n3041_));
OR2X2 OR2X2_632 ( .A(u0__abc_76628_new_n3042_), .B(u0__abc_76628_new_n3043_), .Y(u0__abc_76628_new_n3044_));
OR2X2 OR2X2_633 ( .A(u0__abc_76628_new_n3045_), .B(u0__abc_76628_new_n3046_), .Y(u0__abc_76628_new_n3047_));
OR2X2 OR2X2_634 ( .A(u0__abc_76628_new_n3048_), .B(u0__abc_76628_new_n3049_), .Y(u0__abc_76628_new_n3050_));
OR2X2 OR2X2_635 ( .A(u0__abc_76628_new_n3052_), .B(u0_cs0_bF_buf3), .Y(u0__abc_76628_new_n3053_));
OR2X2 OR2X2_636 ( .A(u0__abc_76628_new_n3051_), .B(u0__abc_76628_new_n3053_), .Y(u0__abc_76628_new_n3054_));
OR2X2 OR2X2_637 ( .A(u0__abc_76628_new_n2742__bF_buf4), .B(u0_tms0_13_), .Y(u0__abc_76628_new_n3055_));
OR2X2 OR2X2_638 ( .A(u0__abc_76628_new_n3057_), .B(u0__abc_76628_new_n3035_), .Y(u0__0tms_31_0__13_));
OR2X2 OR2X2_639 ( .A(u0__abc_76628_new_n2722__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n3061_));
OR2X2 OR2X2_64 ( .A(lmr_sel_bF_buf5), .B(tms_14_), .Y(_abc_85006_new_n333_));
OR2X2 OR2X2_640 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3062_));
OR2X2 OR2X2_641 ( .A(u0__abc_76628_new_n3064_), .B(u0__abc_76628_new_n3060_), .Y(u0__abc_76628_new_n3065_));
OR2X2 OR2X2_642 ( .A(u0__abc_76628_new_n3066_), .B(u0__abc_76628_new_n3067_), .Y(u0__abc_76628_new_n3068_));
OR2X2 OR2X2_643 ( .A(u0__abc_76628_new_n3069_), .B(u0__abc_76628_new_n3070_), .Y(u0__abc_76628_new_n3071_));
OR2X2 OR2X2_644 ( .A(u0__abc_76628_new_n3072_), .B(u0__abc_76628_new_n3073_), .Y(u0__abc_76628_new_n3074_));
OR2X2 OR2X2_645 ( .A(u0__abc_76628_new_n3076_), .B(u0_cs0_bF_buf2), .Y(u0__abc_76628_new_n3077_));
OR2X2 OR2X2_646 ( .A(u0__abc_76628_new_n3075_), .B(u0__abc_76628_new_n3077_), .Y(u0__abc_76628_new_n3078_));
OR2X2 OR2X2_647 ( .A(u0__abc_76628_new_n2742__bF_buf3), .B(u0_tms0_14_), .Y(u0__abc_76628_new_n3079_));
OR2X2 OR2X2_648 ( .A(u0__abc_76628_new_n3081_), .B(u0__abc_76628_new_n3059_), .Y(u0__0tms_31_0__14_));
OR2X2 OR2X2_649 ( .A(u0__abc_76628_new_n2722__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n3085_));
OR2X2 OR2X2_65 ( .A(_abc_85006_new_n240__bF_buf0), .B(sp_tms_15_), .Y(_abc_85006_new_n335_));
OR2X2 OR2X2_650 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3086_));
OR2X2 OR2X2_651 ( .A(u0__abc_76628_new_n3088_), .B(u0__abc_76628_new_n3084_), .Y(u0__abc_76628_new_n3089_));
OR2X2 OR2X2_652 ( .A(u0__abc_76628_new_n3090_), .B(u0__abc_76628_new_n3091_), .Y(u0__abc_76628_new_n3092_));
OR2X2 OR2X2_653 ( .A(u0__abc_76628_new_n3093_), .B(u0__abc_76628_new_n3094_), .Y(u0__abc_76628_new_n3095_));
OR2X2 OR2X2_654 ( .A(u0__abc_76628_new_n3096_), .B(u0__abc_76628_new_n3097_), .Y(u0__abc_76628_new_n3098_));
OR2X2 OR2X2_655 ( .A(u0__abc_76628_new_n3100_), .B(u0_cs0_bF_buf1), .Y(u0__abc_76628_new_n3101_));
OR2X2 OR2X2_656 ( .A(u0__abc_76628_new_n3099_), .B(u0__abc_76628_new_n3101_), .Y(u0__abc_76628_new_n3102_));
OR2X2 OR2X2_657 ( .A(u0__abc_76628_new_n2742__bF_buf2), .B(u0_tms0_15_), .Y(u0__abc_76628_new_n3103_));
OR2X2 OR2X2_658 ( .A(u0__abc_76628_new_n3105_), .B(u0__abc_76628_new_n3083_), .Y(u0__0tms_31_0__15_));
OR2X2 OR2X2_659 ( .A(u0__abc_76628_new_n2722__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n3109_));
OR2X2 OR2X2_66 ( .A(lmr_sel_bF_buf4), .B(tms_15_), .Y(_abc_85006_new_n336_));
OR2X2 OR2X2_660 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3110_));
OR2X2 OR2X2_661 ( .A(u0__abc_76628_new_n3112_), .B(u0__abc_76628_new_n3108_), .Y(u0__abc_76628_new_n3113_));
OR2X2 OR2X2_662 ( .A(u0__abc_76628_new_n3114_), .B(u0__abc_76628_new_n3115_), .Y(u0__abc_76628_new_n3116_));
OR2X2 OR2X2_663 ( .A(u0__abc_76628_new_n3117_), .B(u0__abc_76628_new_n3118_), .Y(u0__abc_76628_new_n3119_));
OR2X2 OR2X2_664 ( .A(u0__abc_76628_new_n3120_), .B(u0__abc_76628_new_n3121_), .Y(u0__abc_76628_new_n3122_));
OR2X2 OR2X2_665 ( .A(u0__abc_76628_new_n3124_), .B(u0_cs0_bF_buf0), .Y(u0__abc_76628_new_n3125_));
OR2X2 OR2X2_666 ( .A(u0__abc_76628_new_n3123_), .B(u0__abc_76628_new_n3125_), .Y(u0__abc_76628_new_n3126_));
OR2X2 OR2X2_667 ( .A(u0__abc_76628_new_n2742__bF_buf1), .B(u0_tms0_16_), .Y(u0__abc_76628_new_n3127_));
OR2X2 OR2X2_668 ( .A(u0__abc_76628_new_n3129_), .B(u0__abc_76628_new_n3107_), .Y(u0__0tms_31_0__16_));
OR2X2 OR2X2_669 ( .A(u0__abc_76628_new_n2722__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n3133_));
OR2X2 OR2X2_67 ( .A(_abc_85006_new_n240__bF_buf5), .B(sp_tms_16_), .Y(_abc_85006_new_n338_));
OR2X2 OR2X2_670 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3134_));
OR2X2 OR2X2_671 ( .A(u0__abc_76628_new_n3136_), .B(u0__abc_76628_new_n3132_), .Y(u0__abc_76628_new_n3137_));
OR2X2 OR2X2_672 ( .A(u0__abc_76628_new_n3138_), .B(u0__abc_76628_new_n3139_), .Y(u0__abc_76628_new_n3140_));
OR2X2 OR2X2_673 ( .A(u0__abc_76628_new_n3141_), .B(u0__abc_76628_new_n3142_), .Y(u0__abc_76628_new_n3143_));
OR2X2 OR2X2_674 ( .A(u0__abc_76628_new_n3144_), .B(u0__abc_76628_new_n3145_), .Y(u0__abc_76628_new_n3146_));
OR2X2 OR2X2_675 ( .A(u0__abc_76628_new_n3148_), .B(u0_cs0_bF_buf5), .Y(u0__abc_76628_new_n3149_));
OR2X2 OR2X2_676 ( .A(u0__abc_76628_new_n3147_), .B(u0__abc_76628_new_n3149_), .Y(u0__abc_76628_new_n3150_));
OR2X2 OR2X2_677 ( .A(u0__abc_76628_new_n2742__bF_buf0), .B(u0_tms0_17_), .Y(u0__abc_76628_new_n3151_));
OR2X2 OR2X2_678 ( .A(u0__abc_76628_new_n3153_), .B(u0__abc_76628_new_n3131_), .Y(u0__0tms_31_0__17_));
OR2X2 OR2X2_679 ( .A(u0__abc_76628_new_n2722__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n3157_));
OR2X2 OR2X2_68 ( .A(lmr_sel_bF_buf3), .B(tms_16_), .Y(_abc_85006_new_n339_));
OR2X2 OR2X2_680 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3158_));
OR2X2 OR2X2_681 ( .A(u0__abc_76628_new_n3160_), .B(u0__abc_76628_new_n3156_), .Y(u0__abc_76628_new_n3161_));
OR2X2 OR2X2_682 ( .A(u0__abc_76628_new_n3162_), .B(u0__abc_76628_new_n3163_), .Y(u0__abc_76628_new_n3164_));
OR2X2 OR2X2_683 ( .A(u0__abc_76628_new_n3165_), .B(u0__abc_76628_new_n3166_), .Y(u0__abc_76628_new_n3167_));
OR2X2 OR2X2_684 ( .A(u0__abc_76628_new_n3168_), .B(u0__abc_76628_new_n3169_), .Y(u0__abc_76628_new_n3170_));
OR2X2 OR2X2_685 ( .A(u0__abc_76628_new_n3172_), .B(u0_cs0_bF_buf4), .Y(u0__abc_76628_new_n3173_));
OR2X2 OR2X2_686 ( .A(u0__abc_76628_new_n3171_), .B(u0__abc_76628_new_n3173_), .Y(u0__abc_76628_new_n3174_));
OR2X2 OR2X2_687 ( .A(u0__abc_76628_new_n2742__bF_buf5), .B(u0_tms0_18_), .Y(u0__abc_76628_new_n3175_));
OR2X2 OR2X2_688 ( .A(u0__abc_76628_new_n3177_), .B(u0__abc_76628_new_n3155_), .Y(u0__0tms_31_0__18_));
OR2X2 OR2X2_689 ( .A(u0__abc_76628_new_n2722__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n3181_));
OR2X2 OR2X2_69 ( .A(_abc_85006_new_n240__bF_buf4), .B(sp_tms_17_), .Y(_abc_85006_new_n341_));
OR2X2 OR2X2_690 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3182_));
OR2X2 OR2X2_691 ( .A(u0__abc_76628_new_n3184_), .B(u0__abc_76628_new_n3180_), .Y(u0__abc_76628_new_n3185_));
OR2X2 OR2X2_692 ( .A(u0__abc_76628_new_n3186_), .B(u0__abc_76628_new_n3187_), .Y(u0__abc_76628_new_n3188_));
OR2X2 OR2X2_693 ( .A(u0__abc_76628_new_n3189_), .B(u0__abc_76628_new_n3190_), .Y(u0__abc_76628_new_n3191_));
OR2X2 OR2X2_694 ( .A(u0__abc_76628_new_n3192_), .B(u0__abc_76628_new_n3193_), .Y(u0__abc_76628_new_n3194_));
OR2X2 OR2X2_695 ( .A(u0__abc_76628_new_n3196_), .B(u0_cs0_bF_buf3), .Y(u0__abc_76628_new_n3197_));
OR2X2 OR2X2_696 ( .A(u0__abc_76628_new_n3195_), .B(u0__abc_76628_new_n3197_), .Y(u0__abc_76628_new_n3198_));
OR2X2 OR2X2_697 ( .A(u0__abc_76628_new_n2742__bF_buf4), .B(u0_tms0_19_), .Y(u0__abc_76628_new_n3199_));
OR2X2 OR2X2_698 ( .A(u0__abc_76628_new_n3201_), .B(u0__abc_76628_new_n3179_), .Y(u0__0tms_31_0__19_));
OR2X2 OR2X2_699 ( .A(u0__abc_76628_new_n2722__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n3205_));
OR2X2 OR2X2_7 ( .A(_abc_85006_new_n240__bF_buf4), .B(spec_req_cs_1_bF_buf5_), .Y(_abc_85006_new_n248_));
OR2X2 OR2X2_70 ( .A(lmr_sel_bF_buf2), .B(tms_17_), .Y(_abc_85006_new_n342_));
OR2X2 OR2X2_700 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3206_));
OR2X2 OR2X2_701 ( .A(u0__abc_76628_new_n3208_), .B(u0__abc_76628_new_n3204_), .Y(u0__abc_76628_new_n3209_));
OR2X2 OR2X2_702 ( .A(u0__abc_76628_new_n3210_), .B(u0__abc_76628_new_n3211_), .Y(u0__abc_76628_new_n3212_));
OR2X2 OR2X2_703 ( .A(u0__abc_76628_new_n3213_), .B(u0__abc_76628_new_n3214_), .Y(u0__abc_76628_new_n3215_));
OR2X2 OR2X2_704 ( .A(u0__abc_76628_new_n3216_), .B(u0__abc_76628_new_n3217_), .Y(u0__abc_76628_new_n3218_));
OR2X2 OR2X2_705 ( .A(u0__abc_76628_new_n3220_), .B(u0_cs0_bF_buf2), .Y(u0__abc_76628_new_n3221_));
OR2X2 OR2X2_706 ( .A(u0__abc_76628_new_n3219_), .B(u0__abc_76628_new_n3221_), .Y(u0__abc_76628_new_n3222_));
OR2X2 OR2X2_707 ( .A(u0__abc_76628_new_n2742__bF_buf3), .B(u0_tms0_20_), .Y(u0__abc_76628_new_n3223_));
OR2X2 OR2X2_708 ( .A(u0__abc_76628_new_n3225_), .B(u0__abc_76628_new_n3203_), .Y(u0__0tms_31_0__20_));
OR2X2 OR2X2_709 ( .A(u0__abc_76628_new_n2722__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n3229_));
OR2X2 OR2X2_71 ( .A(_abc_85006_new_n240__bF_buf3), .B(sp_tms_18_), .Y(_abc_85006_new_n344_));
OR2X2 OR2X2_710 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3230_));
OR2X2 OR2X2_711 ( .A(u0__abc_76628_new_n3232_), .B(u0__abc_76628_new_n3228_), .Y(u0__abc_76628_new_n3233_));
OR2X2 OR2X2_712 ( .A(u0__abc_76628_new_n3234_), .B(u0__abc_76628_new_n3235_), .Y(u0__abc_76628_new_n3236_));
OR2X2 OR2X2_713 ( .A(u0__abc_76628_new_n3237_), .B(u0__abc_76628_new_n3238_), .Y(u0__abc_76628_new_n3239_));
OR2X2 OR2X2_714 ( .A(u0__abc_76628_new_n3240_), .B(u0__abc_76628_new_n3241_), .Y(u0__abc_76628_new_n3242_));
OR2X2 OR2X2_715 ( .A(u0__abc_76628_new_n3244_), .B(u0_cs0_bF_buf1), .Y(u0__abc_76628_new_n3245_));
OR2X2 OR2X2_716 ( .A(u0__abc_76628_new_n3243_), .B(u0__abc_76628_new_n3245_), .Y(u0__abc_76628_new_n3246_));
OR2X2 OR2X2_717 ( .A(u0__abc_76628_new_n2742__bF_buf2), .B(u0_tms0_21_), .Y(u0__abc_76628_new_n3247_));
OR2X2 OR2X2_718 ( .A(u0__abc_76628_new_n3249_), .B(u0__abc_76628_new_n3227_), .Y(u0__0tms_31_0__21_));
OR2X2 OR2X2_719 ( .A(u0__abc_76628_new_n2722__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n3253_));
OR2X2 OR2X2_72 ( .A(lmr_sel_bF_buf1), .B(tms_18_), .Y(_abc_85006_new_n345_));
OR2X2 OR2X2_720 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3254_));
OR2X2 OR2X2_721 ( .A(u0__abc_76628_new_n3256_), .B(u0__abc_76628_new_n3252_), .Y(u0__abc_76628_new_n3257_));
OR2X2 OR2X2_722 ( .A(u0__abc_76628_new_n3258_), .B(u0__abc_76628_new_n3259_), .Y(u0__abc_76628_new_n3260_));
OR2X2 OR2X2_723 ( .A(u0__abc_76628_new_n3261_), .B(u0__abc_76628_new_n3262_), .Y(u0__abc_76628_new_n3263_));
OR2X2 OR2X2_724 ( .A(u0__abc_76628_new_n3264_), .B(u0__abc_76628_new_n3265_), .Y(u0__abc_76628_new_n3266_));
OR2X2 OR2X2_725 ( .A(u0__abc_76628_new_n3268_), .B(u0_cs0_bF_buf0), .Y(u0__abc_76628_new_n3269_));
OR2X2 OR2X2_726 ( .A(u0__abc_76628_new_n3267_), .B(u0__abc_76628_new_n3269_), .Y(u0__abc_76628_new_n3270_));
OR2X2 OR2X2_727 ( .A(u0__abc_76628_new_n2742__bF_buf1), .B(u0_tms0_22_), .Y(u0__abc_76628_new_n3271_));
OR2X2 OR2X2_728 ( .A(u0__abc_76628_new_n3273_), .B(u0__abc_76628_new_n3251_), .Y(u0__0tms_31_0__22_));
OR2X2 OR2X2_729 ( .A(u0__abc_76628_new_n2722__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n3277_));
OR2X2 OR2X2_73 ( .A(_abc_85006_new_n240__bF_buf2), .B(sp_tms_19_), .Y(_abc_85006_new_n347_));
OR2X2 OR2X2_730 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3278_));
OR2X2 OR2X2_731 ( .A(u0__abc_76628_new_n3280_), .B(u0__abc_76628_new_n3276_), .Y(u0__abc_76628_new_n3281_));
OR2X2 OR2X2_732 ( .A(u0__abc_76628_new_n3282_), .B(u0__abc_76628_new_n3283_), .Y(u0__abc_76628_new_n3284_));
OR2X2 OR2X2_733 ( .A(u0__abc_76628_new_n3285_), .B(u0__abc_76628_new_n3286_), .Y(u0__abc_76628_new_n3287_));
OR2X2 OR2X2_734 ( .A(u0__abc_76628_new_n3288_), .B(u0__abc_76628_new_n3289_), .Y(u0__abc_76628_new_n3290_));
OR2X2 OR2X2_735 ( .A(u0__abc_76628_new_n3292_), .B(u0_cs0_bF_buf5), .Y(u0__abc_76628_new_n3293_));
OR2X2 OR2X2_736 ( .A(u0__abc_76628_new_n3291_), .B(u0__abc_76628_new_n3293_), .Y(u0__abc_76628_new_n3294_));
OR2X2 OR2X2_737 ( .A(u0__abc_76628_new_n2742__bF_buf0), .B(u0_tms0_23_), .Y(u0__abc_76628_new_n3295_));
OR2X2 OR2X2_738 ( .A(u0__abc_76628_new_n3297_), .B(u0__abc_76628_new_n3275_), .Y(u0__0tms_31_0__23_));
OR2X2 OR2X2_739 ( .A(u0__abc_76628_new_n2722__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n3301_));
OR2X2 OR2X2_74 ( .A(lmr_sel_bF_buf0), .B(tms_19_), .Y(_abc_85006_new_n348_));
OR2X2 OR2X2_740 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3302_));
OR2X2 OR2X2_741 ( .A(u0__abc_76628_new_n3304_), .B(u0__abc_76628_new_n3300_), .Y(u0__abc_76628_new_n3305_));
OR2X2 OR2X2_742 ( .A(u0__abc_76628_new_n3306_), .B(u0__abc_76628_new_n3307_), .Y(u0__abc_76628_new_n3308_));
OR2X2 OR2X2_743 ( .A(u0__abc_76628_new_n3309_), .B(u0__abc_76628_new_n3310_), .Y(u0__abc_76628_new_n3311_));
OR2X2 OR2X2_744 ( .A(u0__abc_76628_new_n3312_), .B(u0__abc_76628_new_n3313_), .Y(u0__abc_76628_new_n3314_));
OR2X2 OR2X2_745 ( .A(u0__abc_76628_new_n3316_), .B(u0_cs0_bF_buf4), .Y(u0__abc_76628_new_n3317_));
OR2X2 OR2X2_746 ( .A(u0__abc_76628_new_n3315_), .B(u0__abc_76628_new_n3317_), .Y(u0__abc_76628_new_n3318_));
OR2X2 OR2X2_747 ( .A(u0__abc_76628_new_n2742__bF_buf5), .B(u0_tms0_24_), .Y(u0__abc_76628_new_n3319_));
OR2X2 OR2X2_748 ( .A(u0__abc_76628_new_n3321_), .B(u0__abc_76628_new_n3299_), .Y(u0__0tms_31_0__24_));
OR2X2 OR2X2_749 ( .A(u0__abc_76628_new_n2722__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n3325_));
OR2X2 OR2X2_75 ( .A(_abc_85006_new_n240__bF_buf1), .B(sp_tms_20_), .Y(_abc_85006_new_n350_));
OR2X2 OR2X2_750 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3326_));
OR2X2 OR2X2_751 ( .A(u0__abc_76628_new_n3328_), .B(u0__abc_76628_new_n3324_), .Y(u0__abc_76628_new_n3329_));
OR2X2 OR2X2_752 ( .A(u0__abc_76628_new_n3330_), .B(u0__abc_76628_new_n3331_), .Y(u0__abc_76628_new_n3332_));
OR2X2 OR2X2_753 ( .A(u0__abc_76628_new_n3333_), .B(u0__abc_76628_new_n3334_), .Y(u0__abc_76628_new_n3335_));
OR2X2 OR2X2_754 ( .A(u0__abc_76628_new_n3336_), .B(u0__abc_76628_new_n3337_), .Y(u0__abc_76628_new_n3338_));
OR2X2 OR2X2_755 ( .A(u0__abc_76628_new_n3340_), .B(u0_cs0_bF_buf3), .Y(u0__abc_76628_new_n3341_));
OR2X2 OR2X2_756 ( .A(u0__abc_76628_new_n3339_), .B(u0__abc_76628_new_n3341_), .Y(u0__abc_76628_new_n3342_));
OR2X2 OR2X2_757 ( .A(u0__abc_76628_new_n2742__bF_buf4), .B(u0_tms0_25_), .Y(u0__abc_76628_new_n3343_));
OR2X2 OR2X2_758 ( .A(u0__abc_76628_new_n3345_), .B(u0__abc_76628_new_n3323_), .Y(u0__0tms_31_0__25_));
OR2X2 OR2X2_759 ( .A(u0__abc_76628_new_n2722__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n3349_));
OR2X2 OR2X2_76 ( .A(lmr_sel_bF_buf6), .B(tms_20_), .Y(_abc_85006_new_n351_));
OR2X2 OR2X2_760 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3350_));
OR2X2 OR2X2_761 ( .A(u0__abc_76628_new_n3352_), .B(u0__abc_76628_new_n3348_), .Y(u0__abc_76628_new_n3353_));
OR2X2 OR2X2_762 ( .A(u0__abc_76628_new_n3354_), .B(u0__abc_76628_new_n3355_), .Y(u0__abc_76628_new_n3356_));
OR2X2 OR2X2_763 ( .A(u0__abc_76628_new_n3357_), .B(u0__abc_76628_new_n3358_), .Y(u0__abc_76628_new_n3359_));
OR2X2 OR2X2_764 ( .A(u0__abc_76628_new_n3360_), .B(u0__abc_76628_new_n3361_), .Y(u0__abc_76628_new_n3362_));
OR2X2 OR2X2_765 ( .A(u0__abc_76628_new_n3364_), .B(u0_cs0_bF_buf2), .Y(u0__abc_76628_new_n3365_));
OR2X2 OR2X2_766 ( .A(u0__abc_76628_new_n3363_), .B(u0__abc_76628_new_n3365_), .Y(u0__abc_76628_new_n3366_));
OR2X2 OR2X2_767 ( .A(u0__abc_76628_new_n2742__bF_buf3), .B(u0_tms0_26_), .Y(u0__abc_76628_new_n3367_));
OR2X2 OR2X2_768 ( .A(u0__abc_76628_new_n3369_), .B(u0__abc_76628_new_n3347_), .Y(u0__0tms_31_0__26_));
OR2X2 OR2X2_769 ( .A(u0__abc_76628_new_n2722__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n3373_));
OR2X2 OR2X2_77 ( .A(_abc_85006_new_n240__bF_buf0), .B(sp_tms_21_), .Y(_abc_85006_new_n353_));
OR2X2 OR2X2_770 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3374_));
OR2X2 OR2X2_771 ( .A(u0__abc_76628_new_n3376_), .B(u0__abc_76628_new_n3372_), .Y(u0__abc_76628_new_n3377_));
OR2X2 OR2X2_772 ( .A(u0__abc_76628_new_n3378_), .B(u0__abc_76628_new_n3379_), .Y(u0__abc_76628_new_n3380_));
OR2X2 OR2X2_773 ( .A(u0__abc_76628_new_n3381_), .B(u0__abc_76628_new_n3382_), .Y(u0__abc_76628_new_n3383_));
OR2X2 OR2X2_774 ( .A(u0__abc_76628_new_n3384_), .B(u0__abc_76628_new_n3385_), .Y(u0__abc_76628_new_n3386_));
OR2X2 OR2X2_775 ( .A(u0__abc_76628_new_n3388_), .B(u0_cs0_bF_buf1), .Y(u0__abc_76628_new_n3389_));
OR2X2 OR2X2_776 ( .A(u0__abc_76628_new_n3387_), .B(u0__abc_76628_new_n3389_), .Y(u0__abc_76628_new_n3390_));
OR2X2 OR2X2_777 ( .A(u0__abc_76628_new_n2742__bF_buf2), .B(u0_tms0_27_), .Y(u0__abc_76628_new_n3391_));
OR2X2 OR2X2_778 ( .A(u0__abc_76628_new_n3393_), .B(u0__abc_76628_new_n3371_), .Y(u0__0tms_31_0__27_));
OR2X2 OR2X2_779 ( .A(u0__abc_76628_new_n2722__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n3517_));
OR2X2 OR2X2_78 ( .A(lmr_sel_bF_buf5), .B(tms_21_), .Y(_abc_85006_new_n354_));
OR2X2 OR2X2_780 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3518_));
OR2X2 OR2X2_781 ( .A(u0__abc_76628_new_n3520_), .B(u0__abc_76628_new_n3516_), .Y(u0__abc_76628_new_n3521_));
OR2X2 OR2X2_782 ( .A(u0__abc_76628_new_n3522_), .B(u0__abc_76628_new_n3523_), .Y(u0__abc_76628_new_n3524_));
OR2X2 OR2X2_783 ( .A(u0__abc_76628_new_n3525_), .B(u0__abc_76628_new_n3526_), .Y(u0__abc_76628_new_n3527_));
OR2X2 OR2X2_784 ( .A(u0__abc_76628_new_n3528_), .B(u0__abc_76628_new_n3529_), .Y(u0__abc_76628_new_n3530_));
OR2X2 OR2X2_785 ( .A(u0__abc_76628_new_n3532_), .B(u0_cs0_bF_buf0), .Y(u0__abc_76628_new_n3533_));
OR2X2 OR2X2_786 ( .A(u0__abc_76628_new_n3531_), .B(u0__abc_76628_new_n3533_), .Y(u0__abc_76628_new_n3534_));
OR2X2 OR2X2_787 ( .A(u0__abc_76628_new_n2742__bF_buf1), .B(u0_csc0_1_), .Y(u0__abc_76628_new_n3535_));
OR2X2 OR2X2_788 ( .A(u0__abc_76628_new_n3537_), .B(u0__abc_76628_new_n3515_), .Y(u0__0csc_31_0__1_));
OR2X2 OR2X2_789 ( .A(u0__abc_76628_new_n2722__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n3541_));
OR2X2 OR2X2_79 ( .A(_abc_85006_new_n240__bF_buf5), .B(sp_tms_22_), .Y(_abc_85006_new_n356_));
OR2X2 OR2X2_790 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3542_));
OR2X2 OR2X2_791 ( .A(u0__abc_76628_new_n3544_), .B(u0__abc_76628_new_n3540_), .Y(u0__abc_76628_new_n3545_));
OR2X2 OR2X2_792 ( .A(u0__abc_76628_new_n3546_), .B(u0__abc_76628_new_n3547_), .Y(u0__abc_76628_new_n3548_));
OR2X2 OR2X2_793 ( .A(u0__abc_76628_new_n3549_), .B(u0__abc_76628_new_n3550_), .Y(u0__abc_76628_new_n3551_));
OR2X2 OR2X2_794 ( .A(u0__abc_76628_new_n3552_), .B(u0__abc_76628_new_n3553_), .Y(u0__abc_76628_new_n3554_));
OR2X2 OR2X2_795 ( .A(u0__abc_76628_new_n3556_), .B(u0_cs0_bF_buf5), .Y(u0__abc_76628_new_n3557_));
OR2X2 OR2X2_796 ( .A(u0__abc_76628_new_n3555_), .B(u0__abc_76628_new_n3557_), .Y(u0__abc_76628_new_n3558_));
OR2X2 OR2X2_797 ( .A(u0__abc_76628_new_n2742__bF_buf0), .B(u0_csc0_2_), .Y(u0__abc_76628_new_n3559_));
OR2X2 OR2X2_798 ( .A(u0__abc_76628_new_n3561_), .B(u0__abc_76628_new_n3539_), .Y(u0__0csc_31_0__2_));
OR2X2 OR2X2_799 ( .A(u0__abc_76628_new_n2722__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n3565_));
OR2X2 OR2X2_8 ( .A(lmr_sel_bF_buf5), .B(cs_1_), .Y(_abc_85006_new_n249_));
OR2X2 OR2X2_80 ( .A(lmr_sel_bF_buf4), .B(tms_22_), .Y(_abc_85006_new_n357_));
OR2X2 OR2X2_800 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3566_));
OR2X2 OR2X2_801 ( .A(u0__abc_76628_new_n3568_), .B(u0__abc_76628_new_n3564_), .Y(u0__abc_76628_new_n3569_));
OR2X2 OR2X2_802 ( .A(u0__abc_76628_new_n3570_), .B(u0__abc_76628_new_n3571_), .Y(u0__abc_76628_new_n3572_));
OR2X2 OR2X2_803 ( .A(u0__abc_76628_new_n3573_), .B(u0__abc_76628_new_n3574_), .Y(u0__abc_76628_new_n3575_));
OR2X2 OR2X2_804 ( .A(u0__abc_76628_new_n3576_), .B(u0__abc_76628_new_n3577_), .Y(u0__abc_76628_new_n3578_));
OR2X2 OR2X2_805 ( .A(u0__abc_76628_new_n3580_), .B(u0_cs0_bF_buf4), .Y(u0__abc_76628_new_n3581_));
OR2X2 OR2X2_806 ( .A(u0__abc_76628_new_n3579_), .B(u0__abc_76628_new_n3581_), .Y(u0__abc_76628_new_n3582_));
OR2X2 OR2X2_807 ( .A(u0__abc_76628_new_n2742__bF_buf5), .B(u0_csc0_3_), .Y(u0__abc_76628_new_n3583_));
OR2X2 OR2X2_808 ( .A(u0__abc_76628_new_n3585_), .B(u0__abc_76628_new_n3563_), .Y(u0__0csc_31_0__3_));
OR2X2 OR2X2_809 ( .A(u0__abc_76628_new_n2722__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n3589_));
OR2X2 OR2X2_81 ( .A(_abc_85006_new_n240__bF_buf4), .B(sp_tms_23_), .Y(_abc_85006_new_n359_));
OR2X2 OR2X2_810 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3590_));
OR2X2 OR2X2_811 ( .A(u0__abc_76628_new_n3592_), .B(u0__abc_76628_new_n3588_), .Y(u0__abc_76628_new_n3593_));
OR2X2 OR2X2_812 ( .A(u0__abc_76628_new_n3594_), .B(u0__abc_76628_new_n3595_), .Y(u0__abc_76628_new_n3596_));
OR2X2 OR2X2_813 ( .A(u0__abc_76628_new_n3597_), .B(u0__abc_76628_new_n3598_), .Y(u0__abc_76628_new_n3599_));
OR2X2 OR2X2_814 ( .A(u0__abc_76628_new_n3600_), .B(u0__abc_76628_new_n3601_), .Y(u0__abc_76628_new_n3602_));
OR2X2 OR2X2_815 ( .A(u0__abc_76628_new_n3604_), .B(u0_cs0_bF_buf3), .Y(u0__abc_76628_new_n3605_));
OR2X2 OR2X2_816 ( .A(u0__abc_76628_new_n3603_), .B(u0__abc_76628_new_n3605_), .Y(u0__abc_76628_new_n3606_));
OR2X2 OR2X2_817 ( .A(u0__abc_76628_new_n2742__bF_buf4), .B(u0_csc0_4_), .Y(u0__abc_76628_new_n3607_));
OR2X2 OR2X2_818 ( .A(u0__abc_76628_new_n3609_), .B(u0__abc_76628_new_n3587_), .Y(u0__0csc_31_0__4_));
OR2X2 OR2X2_819 ( .A(u0__abc_76628_new_n2722__bF_buf3), .B(1'h0), .Y(u0__abc_76628_new_n3613_));
OR2X2 OR2X2_82 ( .A(lmr_sel_bF_buf3), .B(tms_23_), .Y(_abc_85006_new_n360_));
OR2X2 OR2X2_820 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3614_));
OR2X2 OR2X2_821 ( .A(u0__abc_76628_new_n3616_), .B(u0__abc_76628_new_n3612_), .Y(u0__abc_76628_new_n3617_));
OR2X2 OR2X2_822 ( .A(u0__abc_76628_new_n3618_), .B(u0__abc_76628_new_n3619_), .Y(u0__abc_76628_new_n3620_));
OR2X2 OR2X2_823 ( .A(u0__abc_76628_new_n3621_), .B(u0__abc_76628_new_n3622_), .Y(u0__abc_76628_new_n3623_));
OR2X2 OR2X2_824 ( .A(u0__abc_76628_new_n3624_), .B(u0__abc_76628_new_n3625_), .Y(u0__abc_76628_new_n3626_));
OR2X2 OR2X2_825 ( .A(u0__abc_76628_new_n3628_), .B(u0_cs0_bF_buf2), .Y(u0__abc_76628_new_n3629_));
OR2X2 OR2X2_826 ( .A(u0__abc_76628_new_n3627_), .B(u0__abc_76628_new_n3629_), .Y(u0__abc_76628_new_n3630_));
OR2X2 OR2X2_827 ( .A(u0__abc_76628_new_n2742__bF_buf3), .B(u0_csc0_5_), .Y(u0__abc_76628_new_n3631_));
OR2X2 OR2X2_828 ( .A(u0__abc_76628_new_n3633_), .B(u0__abc_76628_new_n3611_), .Y(u0__0csc_31_0__5_));
OR2X2 OR2X2_829 ( .A(u0__abc_76628_new_n2722__bF_buf2), .B(1'h0), .Y(u0__abc_76628_new_n3637_));
OR2X2 OR2X2_83 ( .A(_abc_85006_new_n240__bF_buf3), .B(sp_tms_24_), .Y(_abc_85006_new_n362_));
OR2X2 OR2X2_830 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3638_));
OR2X2 OR2X2_831 ( .A(u0__abc_76628_new_n3640_), .B(u0__abc_76628_new_n3636_), .Y(u0__abc_76628_new_n3641_));
OR2X2 OR2X2_832 ( .A(u0__abc_76628_new_n3642_), .B(u0__abc_76628_new_n3643_), .Y(u0__abc_76628_new_n3644_));
OR2X2 OR2X2_833 ( .A(u0__abc_76628_new_n3645_), .B(u0__abc_76628_new_n3646_), .Y(u0__abc_76628_new_n3647_));
OR2X2 OR2X2_834 ( .A(u0__abc_76628_new_n3648_), .B(u0__abc_76628_new_n3649_), .Y(u0__abc_76628_new_n3650_));
OR2X2 OR2X2_835 ( .A(u0__abc_76628_new_n3652_), .B(u0_cs0_bF_buf1), .Y(u0__abc_76628_new_n3653_));
OR2X2 OR2X2_836 ( .A(u0__abc_76628_new_n3651_), .B(u0__abc_76628_new_n3653_), .Y(u0__abc_76628_new_n3654_));
OR2X2 OR2X2_837 ( .A(u0__abc_76628_new_n2742__bF_buf2), .B(u0_csc0_6_), .Y(u0__abc_76628_new_n3655_));
OR2X2 OR2X2_838 ( .A(u0__abc_76628_new_n3657_), .B(u0__abc_76628_new_n3635_), .Y(u0__0csc_31_0__6_));
OR2X2 OR2X2_839 ( .A(u0__abc_76628_new_n2722__bF_buf1), .B(1'h0), .Y(u0__abc_76628_new_n3661_));
OR2X2 OR2X2_84 ( .A(lmr_sel_bF_buf2), .B(tms_24_), .Y(_abc_85006_new_n363_));
OR2X2 OR2X2_840 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3662_));
OR2X2 OR2X2_841 ( .A(u0__abc_76628_new_n3664_), .B(u0__abc_76628_new_n3660_), .Y(u0__abc_76628_new_n3665_));
OR2X2 OR2X2_842 ( .A(u0__abc_76628_new_n3666_), .B(u0__abc_76628_new_n3667_), .Y(u0__abc_76628_new_n3668_));
OR2X2 OR2X2_843 ( .A(u0__abc_76628_new_n3669_), .B(u0__abc_76628_new_n3670_), .Y(u0__abc_76628_new_n3671_));
OR2X2 OR2X2_844 ( .A(u0__abc_76628_new_n3672_), .B(u0__abc_76628_new_n3673_), .Y(u0__abc_76628_new_n3674_));
OR2X2 OR2X2_845 ( .A(u0__abc_76628_new_n3676_), .B(u0_cs0_bF_buf0), .Y(u0__abc_76628_new_n3677_));
OR2X2 OR2X2_846 ( .A(u0__abc_76628_new_n3675_), .B(u0__abc_76628_new_n3677_), .Y(u0__abc_76628_new_n3678_));
OR2X2 OR2X2_847 ( .A(u0__abc_76628_new_n2742__bF_buf1), .B(u0_csc0_7_), .Y(u0__abc_76628_new_n3679_));
OR2X2 OR2X2_848 ( .A(u0__abc_76628_new_n3681_), .B(u0__abc_76628_new_n3659_), .Y(u0__0csc_31_0__7_));
OR2X2 OR2X2_849 ( .A(u0__abc_76628_new_n2722__bF_buf0), .B(1'h0), .Y(u0__abc_76628_new_n3709_));
OR2X2 OR2X2_85 ( .A(_abc_85006_new_n240__bF_buf2), .B(sp_tms_25_), .Y(_abc_85006_new_n365_));
OR2X2 OR2X2_850 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3710_));
OR2X2 OR2X2_851 ( .A(u0__abc_76628_new_n3712_), .B(u0__abc_76628_new_n3708_), .Y(u0__abc_76628_new_n3713_));
OR2X2 OR2X2_852 ( .A(u0__abc_76628_new_n3714_), .B(u0__abc_76628_new_n3715_), .Y(u0__abc_76628_new_n3716_));
OR2X2 OR2X2_853 ( .A(u0__abc_76628_new_n3717_), .B(u0__abc_76628_new_n3718_), .Y(u0__abc_76628_new_n3719_));
OR2X2 OR2X2_854 ( .A(u0__abc_76628_new_n3720_), .B(u0__abc_76628_new_n3721_), .Y(u0__abc_76628_new_n3722_));
OR2X2 OR2X2_855 ( .A(u0__abc_76628_new_n3724_), .B(u0_cs0_bF_buf5), .Y(u0__abc_76628_new_n3725_));
OR2X2 OR2X2_856 ( .A(u0__abc_76628_new_n3723_), .B(u0__abc_76628_new_n3725_), .Y(u0__abc_76628_new_n3726_));
OR2X2 OR2X2_857 ( .A(u0__abc_76628_new_n2742__bF_buf0), .B(u0_csc0_9_), .Y(u0__abc_76628_new_n3727_));
OR2X2 OR2X2_858 ( .A(u0__abc_76628_new_n3729_), .B(u0__abc_76628_new_n3707_), .Y(u0__0csc_31_0__9_));
OR2X2 OR2X2_859 ( .A(u0__abc_76628_new_n2722__bF_buf5), .B(1'h0), .Y(u0__abc_76628_new_n3733_));
OR2X2 OR2X2_86 ( .A(lmr_sel_bF_buf1), .B(tms_25_), .Y(_abc_85006_new_n366_));
OR2X2 OR2X2_860 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3734_));
OR2X2 OR2X2_861 ( .A(u0__abc_76628_new_n3736_), .B(u0__abc_76628_new_n3732_), .Y(u0__abc_76628_new_n3737_));
OR2X2 OR2X2_862 ( .A(u0__abc_76628_new_n3738_), .B(u0__abc_76628_new_n3739_), .Y(u0__abc_76628_new_n3740_));
OR2X2 OR2X2_863 ( .A(u0__abc_76628_new_n3741_), .B(u0__abc_76628_new_n3742_), .Y(u0__abc_76628_new_n3743_));
OR2X2 OR2X2_864 ( .A(u0__abc_76628_new_n3744_), .B(u0__abc_76628_new_n3745_), .Y(u0__abc_76628_new_n3746_));
OR2X2 OR2X2_865 ( .A(u0__abc_76628_new_n3748_), .B(u0_cs0_bF_buf4), .Y(u0__abc_76628_new_n3749_));
OR2X2 OR2X2_866 ( .A(u0__abc_76628_new_n3747_), .B(u0__abc_76628_new_n3749_), .Y(u0__abc_76628_new_n3750_));
OR2X2 OR2X2_867 ( .A(u0__abc_76628_new_n2742__bF_buf5), .B(u0_csc0_10_), .Y(u0__abc_76628_new_n3751_));
OR2X2 OR2X2_868 ( .A(u0__abc_76628_new_n3753_), .B(u0__abc_76628_new_n3731_), .Y(u0__0csc_31_0__10_));
OR2X2 OR2X2_869 ( .A(u0__abc_76628_new_n2722__bF_buf4), .B(1'h0), .Y(u0__abc_76628_new_n3757_));
OR2X2 OR2X2_87 ( .A(_abc_85006_new_n240__bF_buf1), .B(sp_tms_26_), .Y(_abc_85006_new_n368_));
OR2X2 OR2X2_870 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n3758_));
OR2X2 OR2X2_871 ( .A(u0__abc_76628_new_n3760_), .B(u0__abc_76628_new_n3756_), .Y(u0__abc_76628_new_n3761_));
OR2X2 OR2X2_872 ( .A(u0__abc_76628_new_n3762_), .B(u0__abc_76628_new_n3763_), .Y(u0__abc_76628_new_n3764_));
OR2X2 OR2X2_873 ( .A(u0__abc_76628_new_n3765_), .B(u0__abc_76628_new_n3766_), .Y(u0__abc_76628_new_n3767_));
OR2X2 OR2X2_874 ( .A(u0__abc_76628_new_n3768_), .B(u0__abc_76628_new_n3769_), .Y(u0__abc_76628_new_n3770_));
OR2X2 OR2X2_875 ( .A(u0__abc_76628_new_n3772_), .B(u0_cs0_bF_buf3), .Y(u0__abc_76628_new_n3773_));
OR2X2 OR2X2_876 ( .A(u0__abc_76628_new_n3771_), .B(u0__abc_76628_new_n3773_), .Y(u0__abc_76628_new_n3774_));
OR2X2 OR2X2_877 ( .A(u0__abc_76628_new_n2742__bF_buf4), .B(u0_csc0_11_), .Y(u0__abc_76628_new_n3775_));
OR2X2 OR2X2_878 ( .A(u0__abc_76628_new_n3777_), .B(u0__abc_76628_new_n3755_), .Y(u0__0csc_31_0__11_));
OR2X2 OR2X2_879 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n4260_));
OR2X2 OR2X2_88 ( .A(lmr_sel_bF_buf0), .B(tms_26_), .Y(_abc_85006_new_n369_));
OR2X2 OR2X2_880 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n4261_));
OR2X2 OR2X2_881 ( .A(u0__abc_76628_new_n4260_), .B(u0__abc_76628_new_n4261_), .Y(u0__abc_76628_new_n4262_));
OR2X2 OR2X2_882 ( .A(1'h0), .B(1'h0), .Y(u0__abc_76628_new_n4263_));
OR2X2 OR2X2_883 ( .A(u0_u1_wp_err), .B(u0_u0_wp_err), .Y(u0__abc_76628_new_n4264_));
OR2X2 OR2X2_884 ( .A(u0__abc_76628_new_n4263_), .B(u0__abc_76628_new_n4264_), .Y(u0__abc_76628_new_n4265_));
OR2X2 OR2X2_885 ( .A(u0__abc_76628_new_n4262_), .B(u0__abc_76628_new_n4265_), .Y(u0__abc_76628_new_n4266_));
OR2X2 OR2X2_886 ( .A(u0__abc_76628_new_n4267_), .B(u0__abc_76628_new_n4270_), .Y(u0__0wp_err_0_0_));
OR2X2 OR2X2_887 ( .A(cs_le_bF_buf3), .B(cs_0_), .Y(u0__abc_76628_new_n4272_));
OR2X2 OR2X2_888 ( .A(u0__abc_76628_new_n4273_), .B(u0_cs0_bF_buf2), .Y(u0__abc_76628_new_n4274_));
OR2X2 OR2X2_889 ( .A(cs_le_bF_buf1), .B(cs_1_), .Y(u0__abc_76628_new_n4276_));
OR2X2 OR2X2_89 ( .A(_abc_85006_new_n240__bF_buf0), .B(sp_tms_27_), .Y(_abc_85006_new_n371_));
OR2X2 OR2X2_890 ( .A(u0__abc_76628_new_n4273_), .B(u0_cs1_bF_buf2), .Y(u0__abc_76628_new_n4277_));
OR2X2 OR2X2_891 ( .A(cs_le_bF_buf0), .B(cs_2_), .Y(u0__abc_76628_new_n4279_));
OR2X2 OR2X2_892 ( .A(u0__abc_76628_new_n4273_), .B(1'h0), .Y(u0__abc_76628_new_n4280_));
OR2X2 OR2X2_893 ( .A(cs_le_bF_buf4), .B(cs_3_), .Y(u0__abc_76628_new_n4282_));
OR2X2 OR2X2_894 ( .A(u0__abc_76628_new_n4273_), .B(1'h0), .Y(u0__abc_76628_new_n4283_));
OR2X2 OR2X2_895 ( .A(cs_le_bF_buf3), .B(cs_4_), .Y(u0__abc_76628_new_n4285_));
OR2X2 OR2X2_896 ( .A(u0__abc_76628_new_n4273_), .B(1'h0), .Y(u0__abc_76628_new_n4286_));
OR2X2 OR2X2_897 ( .A(cs_le_bF_buf2), .B(cs_5_), .Y(u0__abc_76628_new_n4288_));
OR2X2 OR2X2_898 ( .A(u0__abc_76628_new_n4273_), .B(1'h0), .Y(u0__abc_76628_new_n4289_));
OR2X2 OR2X2_899 ( .A(cs_le_bF_buf1), .B(cs_6_), .Y(u0__abc_76628_new_n4291_));
OR2X2 OR2X2_9 ( .A(_abc_85006_new_n250_), .B(_abc_85006_new_n237_), .Y(_abc_85006_new_n251_));
OR2X2 OR2X2_90 ( .A(lmr_sel_bF_buf6), .B(tms_27_), .Y(_abc_85006_new_n372_));
OR2X2 OR2X2_900 ( .A(u0__abc_76628_new_n4273_), .B(1'h0), .Y(u0__abc_76628_new_n4292_));
OR2X2 OR2X2_901 ( .A(cs_le_bF_buf0), .B(cs_7_), .Y(u0__abc_76628_new_n4294_));
OR2X2 OR2X2_902 ( .A(u0__abc_76628_new_n4273_), .B(1'h0), .Y(u0__abc_76628_new_n4295_));
OR2X2 OR2X2_903 ( .A(_auto_iopadmap_cc_368_execute_85523_0_), .B(u0_rst_r3_bF_buf4), .Y(u0__abc_76628_new_n4297_));
OR2X2 OR2X2_904 ( .A(u0__abc_76628_new_n4298__bF_buf4), .B(mc_data_ir_0_), .Y(u0__abc_76628_new_n4299_));
OR2X2 OR2X2_905 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_1_), .Y(u0__abc_76628_new_n4301_));
OR2X2 OR2X2_906 ( .A(u0__abc_76628_new_n4298__bF_buf3), .B(mc_data_ir_1_), .Y(u0__abc_76628_new_n4302_));
OR2X2 OR2X2_907 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_2_), .Y(u0__abc_76628_new_n4304_));
OR2X2 OR2X2_908 ( .A(u0__abc_76628_new_n4298__bF_buf2), .B(mc_data_ir_2_), .Y(u0__abc_76628_new_n4305_));
OR2X2 OR2X2_909 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_3_), .Y(u0__abc_76628_new_n4307_));
OR2X2 OR2X2_91 ( .A(_abc_85006_new_n240__bF_buf5), .B(sp_csc_1_), .Y(_abc_85006_new_n389_));
OR2X2 OR2X2_910 ( .A(u0__abc_76628_new_n4298__bF_buf1), .B(mc_data_ir_3_), .Y(u0__abc_76628_new_n4308_));
OR2X2 OR2X2_911 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_4_), .Y(u0__abc_76628_new_n4310_));
OR2X2 OR2X2_912 ( .A(u0__abc_76628_new_n4298__bF_buf0), .B(mc_data_ir_4_), .Y(u0__abc_76628_new_n4311_));
OR2X2 OR2X2_913 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_5_), .Y(u0__abc_76628_new_n4313_));
OR2X2 OR2X2_914 ( .A(u0__abc_76628_new_n4298__bF_buf4), .B(mc_data_ir_5_), .Y(u0__abc_76628_new_n4314_));
OR2X2 OR2X2_915 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_6_), .Y(u0__abc_76628_new_n4316_));
OR2X2 OR2X2_916 ( .A(u0__abc_76628_new_n4298__bF_buf3), .B(mc_data_ir_6_), .Y(u0__abc_76628_new_n4317_));
OR2X2 OR2X2_917 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_7_), .Y(u0__abc_76628_new_n4319_));
OR2X2 OR2X2_918 ( .A(u0__abc_76628_new_n4298__bF_buf2), .B(mc_data_ir_7_), .Y(u0__abc_76628_new_n4320_));
OR2X2 OR2X2_919 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_8_), .Y(u0__abc_76628_new_n4322_));
OR2X2 OR2X2_92 ( .A(lmr_sel_bF_buf5), .B(csc_1_), .Y(_abc_85006_new_n390_));
OR2X2 OR2X2_920 ( .A(u0__abc_76628_new_n4298__bF_buf1), .B(mc_data_ir_8_), .Y(u0__abc_76628_new_n4323_));
OR2X2 OR2X2_921 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_9_), .Y(u0__abc_76628_new_n4325_));
OR2X2 OR2X2_922 ( .A(u0__abc_76628_new_n4298__bF_buf0), .B(mc_data_ir_9_), .Y(u0__abc_76628_new_n4326_));
OR2X2 OR2X2_923 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_10_), .Y(u0__abc_76628_new_n4328_));
OR2X2 OR2X2_924 ( .A(u0__abc_76628_new_n4298__bF_buf4), .B(mc_data_ir_10_), .Y(u0__abc_76628_new_n4329_));
OR2X2 OR2X2_925 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_11_), .Y(u0__abc_76628_new_n4331_));
OR2X2 OR2X2_926 ( .A(u0__abc_76628_new_n4298__bF_buf3), .B(mc_data_ir_11_), .Y(u0__abc_76628_new_n4332_));
OR2X2 OR2X2_927 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_12_), .Y(u0__abc_76628_new_n4334_));
OR2X2 OR2X2_928 ( .A(u0__abc_76628_new_n4298__bF_buf2), .B(mc_data_ir_12_), .Y(u0__abc_76628_new_n4335_));
OR2X2 OR2X2_929 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_13_), .Y(u0__abc_76628_new_n4337_));
OR2X2 OR2X2_93 ( .A(_abc_85006_new_n240__bF_buf4), .B(sp_csc_2_), .Y(_abc_85006_new_n392_));
OR2X2 OR2X2_930 ( .A(u0__abc_76628_new_n4298__bF_buf1), .B(mc_data_ir_13_), .Y(u0__abc_76628_new_n4338_));
OR2X2 OR2X2_931 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_14_), .Y(u0__abc_76628_new_n4340_));
OR2X2 OR2X2_932 ( .A(u0__abc_76628_new_n4298__bF_buf0), .B(mc_data_ir_14_), .Y(u0__abc_76628_new_n4341_));
OR2X2 OR2X2_933 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_15_), .Y(u0__abc_76628_new_n4343_));
OR2X2 OR2X2_934 ( .A(u0__abc_76628_new_n4298__bF_buf4), .B(mc_data_ir_15_), .Y(u0__abc_76628_new_n4344_));
OR2X2 OR2X2_935 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_16_), .Y(u0__abc_76628_new_n4346_));
OR2X2 OR2X2_936 ( .A(u0__abc_76628_new_n4298__bF_buf3), .B(mc_data_ir_16_), .Y(u0__abc_76628_new_n4347_));
OR2X2 OR2X2_937 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_17_), .Y(u0__abc_76628_new_n4349_));
OR2X2 OR2X2_938 ( .A(u0__abc_76628_new_n4298__bF_buf2), .B(mc_data_ir_17_), .Y(u0__abc_76628_new_n4350_));
OR2X2 OR2X2_939 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_18_), .Y(u0__abc_76628_new_n4352_));
OR2X2 OR2X2_94 ( .A(lmr_sel_bF_buf4), .B(csc_2_), .Y(_abc_85006_new_n393_));
OR2X2 OR2X2_940 ( .A(u0__abc_76628_new_n4298__bF_buf1), .B(mc_data_ir_18_), .Y(u0__abc_76628_new_n4353_));
OR2X2 OR2X2_941 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_19_), .Y(u0__abc_76628_new_n4355_));
OR2X2 OR2X2_942 ( .A(u0__abc_76628_new_n4298__bF_buf0), .B(mc_data_ir_19_), .Y(u0__abc_76628_new_n4356_));
OR2X2 OR2X2_943 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_20_), .Y(u0__abc_76628_new_n4358_));
OR2X2 OR2X2_944 ( .A(u0__abc_76628_new_n4298__bF_buf4), .B(mc_data_ir_20_), .Y(u0__abc_76628_new_n4359_));
OR2X2 OR2X2_945 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_21_), .Y(u0__abc_76628_new_n4361_));
OR2X2 OR2X2_946 ( .A(u0__abc_76628_new_n4298__bF_buf3), .B(mc_data_ir_21_), .Y(u0__abc_76628_new_n4362_));
OR2X2 OR2X2_947 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_22_), .Y(u0__abc_76628_new_n4364_));
OR2X2 OR2X2_948 ( .A(u0__abc_76628_new_n4298__bF_buf2), .B(mc_data_ir_22_), .Y(u0__abc_76628_new_n4365_));
OR2X2 OR2X2_949 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_23_), .Y(u0__abc_76628_new_n4367_));
OR2X2 OR2X2_95 ( .A(_abc_85006_new_n240__bF_buf3), .B(sp_csc_3_), .Y(_abc_85006_new_n395_));
OR2X2 OR2X2_950 ( .A(u0__abc_76628_new_n4298__bF_buf1), .B(mc_data_ir_23_), .Y(u0__abc_76628_new_n4368_));
OR2X2 OR2X2_951 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_24_), .Y(u0__abc_76628_new_n4370_));
OR2X2 OR2X2_952 ( .A(u0__abc_76628_new_n4298__bF_buf0), .B(mc_data_ir_24_), .Y(u0__abc_76628_new_n4371_));
OR2X2 OR2X2_953 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_25_), .Y(u0__abc_76628_new_n4373_));
OR2X2 OR2X2_954 ( .A(u0__abc_76628_new_n4298__bF_buf4), .B(mc_data_ir_25_), .Y(u0__abc_76628_new_n4374_));
OR2X2 OR2X2_955 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_26_), .Y(u0__abc_76628_new_n4376_));
OR2X2 OR2X2_956 ( .A(u0__abc_76628_new_n4298__bF_buf3), .B(mc_data_ir_26_), .Y(u0__abc_76628_new_n4377_));
OR2X2 OR2X2_957 ( .A(u0_rst_r3_bF_buf1), .B(_auto_iopadmap_cc_368_execute_85523_27_), .Y(u0__abc_76628_new_n4379_));
OR2X2 OR2X2_958 ( .A(u0__abc_76628_new_n4298__bF_buf2), .B(mc_data_ir_27_), .Y(u0__abc_76628_new_n4380_));
OR2X2 OR2X2_959 ( .A(u0_rst_r3_bF_buf0), .B(_auto_iopadmap_cc_368_execute_85523_28_), .Y(u0__abc_76628_new_n4382_));
OR2X2 OR2X2_96 ( .A(lmr_sel_bF_buf3), .B(csc_3_), .Y(_abc_85006_new_n396_));
OR2X2 OR2X2_960 ( .A(u0__abc_76628_new_n4298__bF_buf1), .B(mc_data_ir_28_), .Y(u0__abc_76628_new_n4383_));
OR2X2 OR2X2_961 ( .A(u0_rst_r3_bF_buf4), .B(_auto_iopadmap_cc_368_execute_85523_29_), .Y(u0__abc_76628_new_n4385_));
OR2X2 OR2X2_962 ( .A(u0__abc_76628_new_n4298__bF_buf0), .B(mc_data_ir_29_), .Y(u0__abc_76628_new_n4386_));
OR2X2 OR2X2_963 ( .A(u0_rst_r3_bF_buf3), .B(_auto_iopadmap_cc_368_execute_85523_30_), .Y(u0__abc_76628_new_n4388_));
OR2X2 OR2X2_964 ( .A(u0__abc_76628_new_n4298__bF_buf4), .B(mc_data_ir_30_), .Y(u0__abc_76628_new_n4389_));
OR2X2 OR2X2_965 ( .A(u0_rst_r3_bF_buf2), .B(_auto_iopadmap_cc_368_execute_85523_31_), .Y(u0__abc_76628_new_n4391_));
OR2X2 OR2X2_966 ( .A(u0__abc_76628_new_n4298__bF_buf3), .B(mc_data_ir_31_), .Y(u0__abc_76628_new_n4392_));
OR2X2 OR2X2_967 ( .A(u0_wb_addr_r_5_), .B(u0_wb_addr_r_4_), .Y(u0__abc_76628_new_n4394_));
OR2X2 OR2X2_968 ( .A(u0__abc_76628_new_n4394_), .B(u0_wb_addr_r_6_), .Y(u0__abc_76628_new_n4395_));
OR2X2 OR2X2_969 ( .A(u0__abc_76628_new_n4397_), .B(u0_wb_addr_r_2_), .Y(u0__abc_76628_new_n4398_));
OR2X2 OR2X2_97 ( .A(_abc_85006_new_n240__bF_buf2), .B(sp_csc_4_), .Y(_abc_85006_new_n398_));
OR2X2 OR2X2_970 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_0_), .Y(u0__abc_76628_new_n4402_));
OR2X2 OR2X2_971 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[0] ), .Y(u0__abc_76628_new_n4404_));
OR2X2 OR2X2_972 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_1_), .Y(u0__abc_76628_new_n4406_));
OR2X2 OR2X2_973 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[1] ), .Y(u0__abc_76628_new_n4407_));
OR2X2 OR2X2_974 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_2_), .Y(u0__abc_76628_new_n4409_));
OR2X2 OR2X2_975 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[2] ), .Y(u0__abc_76628_new_n4410_));
OR2X2 OR2X2_976 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_3_), .Y(u0__abc_76628_new_n4412_));
OR2X2 OR2X2_977 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[3] ), .Y(u0__abc_76628_new_n4413_));
OR2X2 OR2X2_978 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_4_), .Y(u0__abc_76628_new_n4415_));
OR2X2 OR2X2_979 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[4] ), .Y(u0__abc_76628_new_n4416_));
OR2X2 OR2X2_98 ( .A(lmr_sel_bF_buf2), .B(csc_4_), .Y(_abc_85006_new_n399_));
OR2X2 OR2X2_980 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_5_), .Y(u0__abc_76628_new_n4418_));
OR2X2 OR2X2_981 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[5] ), .Y(u0__abc_76628_new_n4419_));
OR2X2 OR2X2_982 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_6_), .Y(u0__abc_76628_new_n4421_));
OR2X2 OR2X2_983 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[6] ), .Y(u0__abc_76628_new_n4422_));
OR2X2 OR2X2_984 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_7_), .Y(u0__abc_76628_new_n4424_));
OR2X2 OR2X2_985 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[7] ), .Y(u0__abc_76628_new_n4425_));
OR2X2 OR2X2_986 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_8_), .Y(u0__abc_76628_new_n4427_));
OR2X2 OR2X2_987 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[8] ), .Y(u0__abc_76628_new_n4428_));
OR2X2 OR2X2_988 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_9_), .Y(u0__abc_76628_new_n4430_));
OR2X2 OR2X2_989 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[9] ), .Y(u0__abc_76628_new_n4431_));
OR2X2 OR2X2_99 ( .A(_abc_85006_new_n240__bF_buf1), .B(sp_csc_5_), .Y(_abc_85006_new_n401_));
OR2X2 OR2X2_990 ( .A(u0__abc_76628_new_n4401_), .B(u0_csc_mask_10_), .Y(u0__abc_76628_new_n4433_));
OR2X2 OR2X2_991 ( .A(u0__abc_76628_new_n4403_), .B(\wb_data_i[10] ), .Y(u0__abc_76628_new_n4434_));
OR2X2 OR2X2_992 ( .A(u0__abc_76628_new_n4398_), .B(u0_wb_addr_r_3_), .Y(u0__abc_76628_new_n4436_));
OR2X2 OR2X2_993 ( .A(u0__abc_76628_new_n4436_), .B(u0__abc_76628_new_n4395_), .Y(u0__abc_76628_new_n4437_));
OR2X2 OR2X2_994 ( .A(u0__abc_76628_new_n4438__bF_buf3), .B(u0_csr_1_), .Y(u0__abc_76628_new_n4439_));
OR2X2 OR2X2_995 ( .A(u0__abc_76628_new_n4437__bF_buf2), .B(\wb_data_i[1] ), .Y(u0__abc_76628_new_n4440_));
OR2X2 OR2X2_996 ( .A(u0__abc_76628_new_n4438__bF_buf2), .B(fs), .Y(u0__abc_76628_new_n4442_));
OR2X2 OR2X2_997 ( .A(u0__abc_76628_new_n4437__bF_buf1), .B(\wb_data_i[2] ), .Y(u0__abc_76628_new_n4443_));
OR2X2 OR2X2_998 ( .A(u0__abc_76628_new_n4438__bF_buf1), .B(u0_csr_3_), .Y(u0__abc_76628_new_n4445_));
OR2X2 OR2X2_999 ( .A(u0__abc_76628_new_n4437__bF_buf0), .B(\wb_data_i[3] ), .Y(u0__abc_76628_new_n4446_));


endmodule