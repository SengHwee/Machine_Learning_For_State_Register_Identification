module b10_reset(clock, RESET_G, nRESET_G, R_BUTTON, G_BUTTON, KEY, START, TEST, RTS, RTR, V_IN_3_, V_IN_2_, V_IN_1_, V_IN_0_, CTS_REG, CTR_REG, V_OUT_REG_3_, V_OUT_REG_2_, V_OUT_REG_1_, V_OUT_REG_0_);
  output CTR_REG;
  output CTS_REG;
  input G_BUTTON;
  input KEY;
  wire LAST_G_REG;
  wire LAST_R_REG;
  input RESET_G;
  input RTR;
  input RTS;
  input R_BUTTON;
  wire SIGN_REG_3_;
  input START;
  wire STATO_REG_0_;
  wire STATO_REG_1_;
  wire STATO_REG_2_;
  wire STATO_REG_3_;
  input TEST;
  wire VOTO0_REG;
  wire VOTO1_REG;
  wire VOTO2_REG;
  wire VOTO3_REG;
  input V_IN_0_;
  input V_IN_1_;
  input V_IN_2_;
  input V_IN_3_;
  output V_OUT_REG_0_;
  output V_OUT_REG_1_;
  output V_OUT_REG_2_;
  output V_OUT_REG_3_;
  wire _abc_1116_n100_1;
  wire _abc_1116_n101;
  wire _abc_1116_n102_1;
  wire _abc_1116_n103;
  wire _abc_1116_n104;
  wire _abc_1116_n105;
  wire _abc_1116_n106;
  wire _abc_1116_n107;
  wire _abc_1116_n108;
  wire _abc_1116_n109;
  wire _abc_1116_n110_1;
  wire _abc_1116_n111;
  wire _abc_1116_n112;
  wire _abc_1116_n113_1;
  wire _abc_1116_n114;
  wire _abc_1116_n115_1;
  wire _abc_1116_n116;
  wire _abc_1116_n117;
  wire _abc_1116_n118;
  wire _abc_1116_n120;
  wire _abc_1116_n121;
  wire _abc_1116_n122;
  wire _abc_1116_n123;
  wire _abc_1116_n124_1;
  wire _abc_1116_n125;
  wire _abc_1116_n126;
  wire _abc_1116_n127;
  wire _abc_1116_n128;
  wire _abc_1116_n129;
  wire _abc_1116_n130;
  wire _abc_1116_n131;
  wire _abc_1116_n132;
  wire _abc_1116_n133_1;
  wire _abc_1116_n134_1;
  wire _abc_1116_n135;
  wire _abc_1116_n137;
  wire _abc_1116_n138_1;
  wire _abc_1116_n139;
  wire _abc_1116_n140_1;
  wire _abc_1116_n141;
  wire _abc_1116_n142;
  wire _abc_1116_n143;
  wire _abc_1116_n144;
  wire _abc_1116_n146_1;
  wire _abc_1116_n147;
  wire _abc_1116_n148_1;
  wire _abc_1116_n149;
  wire _abc_1116_n150;
  wire _abc_1116_n151;
  wire _abc_1116_n152;
  wire _abc_1116_n153;
  wire _abc_1116_n155_1;
  wire _abc_1116_n156_1;
  wire _abc_1116_n157;
  wire _abc_1116_n158;
  wire _abc_1116_n160;
  wire _abc_1116_n161;
  wire _abc_1116_n162;
  wire _abc_1116_n164;
  wire _abc_1116_n165;
  wire _abc_1116_n166;
  wire _abc_1116_n168;
  wire _abc_1116_n169;
  wire _abc_1116_n170_1;
  wire _abc_1116_n172;
  wire _abc_1116_n173;
  wire _abc_1116_n174;
  wire _abc_1116_n175;
  wire _abc_1116_n176;
  wire _abc_1116_n177;
  wire _abc_1116_n178;
  wire _abc_1116_n179;
  wire _abc_1116_n180;
  wire _abc_1116_n181;
  wire _abc_1116_n182;
  wire _abc_1116_n183;
  wire _abc_1116_n184;
  wire _abc_1116_n185;
  wire _abc_1116_n186;
  wire _abc_1116_n187;
  wire _abc_1116_n188;
  wire _abc_1116_n189;
  wire _abc_1116_n190;
  wire _abc_1116_n191;
  wire _abc_1116_n192;
  wire _abc_1116_n193;
  wire _abc_1116_n194;
  wire _abc_1116_n195;
  wire _abc_1116_n196;
  wire _abc_1116_n197;
  wire _abc_1116_n198;
  wire _abc_1116_n200;
  wire _abc_1116_n201;
  wire _abc_1116_n202;
  wire _abc_1116_n203;
  wire _abc_1116_n204;
  wire _abc_1116_n205;
  wire _abc_1116_n206;
  wire _abc_1116_n207;
  wire _abc_1116_n208;
  wire _abc_1116_n209;
  wire _abc_1116_n210;
  wire _abc_1116_n211;
  wire _abc_1116_n212;
  wire _abc_1116_n213;
  wire _abc_1116_n214;
  wire _abc_1116_n215;
  wire _abc_1116_n216;
  wire _abc_1116_n217;
  wire _abc_1116_n219;
  wire _abc_1116_n220;
  wire _abc_1116_n221;
  wire _abc_1116_n222;
  wire _abc_1116_n223;
  wire _abc_1116_n225;
  wire _abc_1116_n226;
  wire _abc_1116_n227;
  wire _abc_1116_n228;
  wire _abc_1116_n229;
  wire _abc_1116_n230;
  wire _abc_1116_n231;
  wire _abc_1116_n232;
  wire _abc_1116_n233;
  wire _abc_1116_n234;
  wire _abc_1116_n235;
  wire _abc_1116_n236;
  wire _abc_1116_n237;
  wire _abc_1116_n239;
  wire _abc_1116_n240;
  wire _abc_1116_n241;
  wire _abc_1116_n243;
  wire _abc_1116_n244;
  wire _abc_1116_n245;
  wire _abc_1116_n246;
  wire _abc_1116_n247;
  wire _abc_1116_n248;
  wire _abc_1116_n249;
  wire _abc_1116_n250;
  wire _abc_1116_n251;
  wire _abc_1116_n252;
  wire _abc_1116_n253;
  wire _abc_1116_n254;
  wire _abc_1116_n255;
  wire _abc_1116_n256;
  wire _abc_1116_n257;
  wire _abc_1116_n258;
  wire _abc_1116_n259;
  wire _abc_1116_n260;
  wire _abc_1116_n262;
  wire _abc_1116_n263;
  wire _abc_1116_n264;
  wire _abc_1116_n265;
  wire _abc_1116_n266;
  wire _abc_1116_n267;
  wire _abc_1116_n268;
  wire _abc_1116_n269;
  wire _abc_1116_n270;
  wire _abc_1116_n271;
  wire _abc_1116_n272;
  wire _abc_1116_n273;
  wire _abc_1116_n274;
  wire _abc_1116_n47;
  wire _abc_1116_n48_1;
  wire _abc_1116_n49;
  wire _abc_1116_n50;
  wire _abc_1116_n51;
  wire _abc_1116_n52;
  wire _abc_1116_n53;
  wire _abc_1116_n54;
  wire _abc_1116_n55;
  wire _abc_1116_n56;
  wire _abc_1116_n57;
  wire _abc_1116_n58;
  wire _abc_1116_n59;
  wire _abc_1116_n60;
  wire _abc_1116_n61_1;
  wire _abc_1116_n62;
  wire _abc_1116_n64;
  wire _abc_1116_n65_1;
  wire _abc_1116_n66;
  wire _abc_1116_n67_1;
  wire _abc_1116_n68;
  wire _abc_1116_n69_1;
  wire _abc_1116_n70;
  wire _abc_1116_n71;
  wire _abc_1116_n72;
  wire _abc_1116_n73;
  wire _abc_1116_n74;
  wire _abc_1116_n75;
  wire _abc_1116_n77;
  wire _abc_1116_n78;
  wire _abc_1116_n79;
  wire _abc_1116_n80;
  wire _abc_1116_n81_1;
  wire _abc_1116_n82;
  wire _abc_1116_n83;
  wire _abc_1116_n84;
  wire _abc_1116_n85;
  wire _abc_1116_n86;
  wire _abc_1116_n87_1;
  wire _abc_1116_n88;
  wire _abc_1116_n89_1;
  wire _abc_1116_n90;
  wire _abc_1116_n91_1;
  wire _abc_1116_n92;
  wire _abc_1116_n93_1;
  wire _abc_1116_n94;
  wire _abc_1116_n95_1;
  wire _abc_1116_n96;
  wire _abc_1116_n97_1;
  wire _abc_1116_n98;
  wire _abc_1116_n99_1;
  input clock;
  wire clock_bF_buf0;
  wire clock_bF_buf1;
  wire clock_bF_buf2;
  wire clock_bF_buf3;
  wire n100;
  wire n105;
  wire n109;
  wire n114;
  wire n40;
  wire n45;
  wire n50;
  wire n55;
  wire n60;
  wire n65;
  wire n69;
  wire n73;
  wire n77;
  wire n81;
  wire n86;
  wire n91;
  wire n95;
  input nRESET_G;
  AND2X2 AND2X2_1 ( .A(_abc_1116_n47), .B(STATO_REG_2_), .Y(_abc_1116_n48_1) );
  AND2X2 AND2X2_10 ( .A(_abc_1116_n69_1), .B(_abc_1116_n64), .Y(_abc_1116_n70) );
  AND2X2 AND2X2_100 ( .A(_abc_1116_n253), .B(STATO_REG_3_), .Y(_abc_1116_n254) );
  AND2X2 AND2X2_101 ( .A(_abc_1116_n254), .B(STATO_REG_1_), .Y(_abc_1116_n255) );
  AND2X2 AND2X2_102 ( .A(_abc_1116_n250), .B(_abc_1116_n257), .Y(_abc_1116_n258) );
  AND2X2 AND2X2_103 ( .A(_abc_1116_n249), .B(VOTO0_REG), .Y(_abc_1116_n259) );
  AND2X2 AND2X2_104 ( .A(_abc_1116_n60), .B(STATO_REG_3_), .Y(_abc_1116_n262) );
  AND2X2 AND2X2_105 ( .A(_abc_1116_n263), .B(RTR), .Y(_abc_1116_n264) );
  AND2X2 AND2X2_106 ( .A(_abc_1116_n267), .B(CTS_REG), .Y(_abc_1116_n268) );
  AND2X2 AND2X2_107 ( .A(_abc_1116_n68), .B(_abc_1116_n60), .Y(_abc_1116_n269) );
  AND2X2 AND2X2_108 ( .A(_abc_1116_n270), .B(RTR), .Y(_abc_1116_n271) );
  AND2X2 AND2X2_109 ( .A(_abc_1116_n55), .B(_abc_1116_n87_1), .Y(_abc_1116_n272) );
  AND2X2 AND2X2_11 ( .A(_abc_1116_n70), .B(_abc_1116_n54), .Y(_abc_1116_n71) );
  AND2X2 AND2X2_12 ( .A(_abc_1116_n72), .B(SIGN_REG_3_), .Y(_abc_1116_n73) );
  AND2X2 AND2X2_13 ( .A(STATO_REG_0_), .B(STATO_REG_3_), .Y(_abc_1116_n74) );
  AND2X2 AND2X2_14 ( .A(_abc_1116_n54), .B(RTR), .Y(_abc_1116_n77) );
  AND2X2 AND2X2_15 ( .A(_abc_1116_n65_1), .B(STATO_REG_3_), .Y(_abc_1116_n79) );
  AND2X2 AND2X2_16 ( .A(_abc_1116_n52), .B(_abc_1116_n79), .Y(_abc_1116_n80) );
  AND2X2 AND2X2_17 ( .A(_abc_1116_n80), .B(_abc_1116_n78), .Y(_abc_1116_n81_1) );
  AND2X2 AND2X2_18 ( .A(V_IN_3_), .B(V_IN_1_), .Y(_abc_1116_n82) );
  AND2X2 AND2X2_19 ( .A(V_IN_0_), .B(V_IN_2_), .Y(_abc_1116_n83) );
  AND2X2 AND2X2_2 ( .A(STATO_REG_1_), .B(STATO_REG_2_), .Y(_abc_1116_n51) );
  AND2X2 AND2X2_20 ( .A(_abc_1116_n82), .B(_abc_1116_n83), .Y(_abc_1116_n84) );
  AND2X2 AND2X2_21 ( .A(_abc_1116_n84), .B(_abc_1116_n74), .Y(_abc_1116_n85) );
  AND2X2 AND2X2_22 ( .A(_abc_1116_n65_1), .B(STATO_REG_2_), .Y(_abc_1116_n87_1) );
  AND2X2 AND2X2_23 ( .A(_abc_1116_n77), .B(_abc_1116_n87_1), .Y(_abc_1116_n88) );
  AND2X2 AND2X2_24 ( .A(STATO_REG_1_), .B(STATO_REG_0_), .Y(_abc_1116_n91_1) );
  AND2X2 AND2X2_25 ( .A(_abc_1116_n92), .B(STATO_REG_2_), .Y(_abc_1116_n93_1) );
  AND2X2 AND2X2_26 ( .A(_abc_1116_n93_1), .B(_abc_1116_n91_1), .Y(_abc_1116_n94) );
  AND2X2 AND2X2_27 ( .A(_abc_1116_n67_1), .B(START), .Y(_abc_1116_n96) );
  AND2X2 AND2X2_28 ( .A(_abc_1116_n66), .B(STATO_REG_0_), .Y(_abc_1116_n97_1) );
  AND2X2 AND2X2_29 ( .A(_abc_1116_n96), .B(_abc_1116_n97_1), .Y(_abc_1116_n98) );
  AND2X2 AND2X2_3 ( .A(_abc_1116_n52), .B(_abc_1116_n50), .Y(_abc_1116_n53) );
  AND2X2 AND2X2_30 ( .A(_abc_1116_n99_1), .B(STATO_REG_1_), .Y(_abc_1116_n100_1) );
  AND2X2 AND2X2_31 ( .A(_abc_1116_n68), .B(_abc_1116_n100_1), .Y(_abc_1116_n101) );
  AND2X2 AND2X2_32 ( .A(_abc_1116_n105), .B(_abc_1116_n106), .Y(_abc_1116_n107) );
  AND2X2 AND2X2_33 ( .A(_abc_1116_n109), .B(_abc_1116_n57), .Y(_abc_1116_n110_1) );
  AND2X2 AND2X2_34 ( .A(_abc_1116_n110_1), .B(_abc_1116_n108), .Y(_abc_1116_n111) );
  AND2X2 AND2X2_35 ( .A(_abc_1116_n111), .B(STATO_REG_1_), .Y(_abc_1116_n112) );
  AND2X2 AND2X2_36 ( .A(_abc_1116_n65_1), .B(_abc_1116_n66), .Y(_abc_1116_n113_1) );
  AND2X2 AND2X2_37 ( .A(_abc_1116_n113_1), .B(STATO_REG_1_), .Y(_abc_1116_n114) );
  AND2X2 AND2X2_38 ( .A(_abc_1116_n87_1), .B(STATO_REG_1_), .Y(_abc_1116_n115_1) );
  AND2X2 AND2X2_39 ( .A(_abc_1116_n120), .B(VOTO1_REG), .Y(_abc_1116_n121) );
  AND2X2 AND2X2_4 ( .A(_abc_1116_n54), .B(STATO_REG_3_), .Y(_abc_1116_n55) );
  AND2X2 AND2X2_40 ( .A(_abc_1116_n125), .B(_abc_1116_n65_1), .Y(_abc_1116_n126) );
  AND2X2 AND2X2_41 ( .A(_abc_1116_n128), .B(STATO_REG_2_), .Y(_abc_1116_n129) );
  AND2X2 AND2X2_42 ( .A(_abc_1116_n130), .B(_abc_1116_n131), .Y(_abc_1116_n132) );
  AND2X2 AND2X2_43 ( .A(_abc_1116_n133_1), .B(STATO_REG_1_), .Y(_abc_1116_n134_1) );
  AND2X2 AND2X2_44 ( .A(_abc_1116_n137), .B(STATO_REG_3_), .Y(_abc_1116_n138_1) );
  AND2X2 AND2X2_45 ( .A(_abc_1116_n87_1), .B(_abc_1116_n54), .Y(_abc_1116_n139) );
  AND2X2 AND2X2_46 ( .A(_abc_1116_n140_1), .B(_abc_1116_n139), .Y(_abc_1116_n141) );
  AND2X2 AND2X2_47 ( .A(_abc_1116_n105), .B(_abc_1116_n142), .Y(_abc_1116_n143) );
  AND2X2 AND2X2_48 ( .A(_abc_1116_n54), .B(_abc_1116_n65_1), .Y(_abc_1116_n146_1) );
  AND2X2 AND2X2_49 ( .A(_abc_1116_n147), .B(_abc_1116_n146_1), .Y(_abc_1116_n148_1) );
  AND2X2 AND2X2_5 ( .A(_abc_1116_n57), .B(CTR_REG), .Y(_abc_1116_n58) );
  AND2X2 AND2X2_50 ( .A(_abc_1116_n105), .B(_abc_1116_n150), .Y(_abc_1116_n151) );
  AND2X2 AND2X2_51 ( .A(_abc_1116_n111), .B(STATO_REG_0_), .Y(_abc_1116_n152) );
  AND2X2 AND2X2_52 ( .A(_abc_1116_n155_1), .B(V_OUT_REG_3_), .Y(_abc_1116_n156_1) );
  AND2X2 AND2X2_53 ( .A(_abc_1116_n88), .B(VOTO3_REG), .Y(_abc_1116_n157) );
  AND2X2 AND2X2_54 ( .A(_abc_1116_n155_1), .B(V_OUT_REG_2_), .Y(_abc_1116_n160) );
  AND2X2 AND2X2_55 ( .A(_abc_1116_n88), .B(VOTO2_REG), .Y(_abc_1116_n161) );
  AND2X2 AND2X2_56 ( .A(_abc_1116_n155_1), .B(V_OUT_REG_1_), .Y(_abc_1116_n164) );
  AND2X2 AND2X2_57 ( .A(_abc_1116_n88), .B(VOTO1_REG), .Y(_abc_1116_n165) );
  AND2X2 AND2X2_58 ( .A(_abc_1116_n155_1), .B(V_OUT_REG_0_), .Y(_abc_1116_n168) );
  AND2X2 AND2X2_59 ( .A(_abc_1116_n88), .B(VOTO0_REG), .Y(_abc_1116_n169) );
  AND2X2 AND2X2_6 ( .A(_abc_1116_n54), .B(STATO_REG_0_), .Y(_abc_1116_n60) );
  AND2X2 AND2X2_60 ( .A(_abc_1116_n113_1), .B(_abc_1116_n96), .Y(_abc_1116_n172) );
  AND2X2 AND2X2_61 ( .A(_abc_1116_n174), .B(G_BUTTON), .Y(_abc_1116_n175) );
  AND2X2 AND2X2_62 ( .A(_abc_1116_n176), .B(_abc_1116_n172), .Y(_abc_1116_n177) );
  AND2X2 AND2X2_63 ( .A(_abc_1116_n60), .B(_abc_1116_n96), .Y(_abc_1116_n179) );
  AND2X2 AND2X2_64 ( .A(_abc_1116_n57), .B(_abc_1116_n182), .Y(_abc_1116_n183) );
  AND2X2 AND2X2_65 ( .A(_abc_1116_n183), .B(_abc_1116_n180), .Y(_abc_1116_n184) );
  AND2X2 AND2X2_66 ( .A(_abc_1116_n184), .B(_abc_1116_n178), .Y(_abc_1116_n185) );
  AND2X2 AND2X2_67 ( .A(STATO_REG_1_), .B(KEY), .Y(_abc_1116_n188) );
  AND2X2 AND2X2_68 ( .A(_abc_1116_n188), .B(_abc_1116_n67_1), .Y(_abc_1116_n189) );
  AND2X2 AND2X2_69 ( .A(_abc_1116_n189), .B(_abc_1116_n187), .Y(_abc_1116_n190) );
  AND2X2 AND2X2_7 ( .A(_abc_1116_n48_1), .B(_abc_1116_n60), .Y(_abc_1116_n61_1) );
  AND2X2 AND2X2_70 ( .A(_abc_1116_n115_1), .B(_abc_1116_n66), .Y(_abc_1116_n192) );
  AND2X2 AND2X2_71 ( .A(_abc_1116_n193), .B(V_IN_1_), .Y(_abc_1116_n194) );
  AND2X2 AND2X2_72 ( .A(_abc_1116_n186), .B(_abc_1116_n195), .Y(_abc_1116_n196) );
  AND2X2 AND2X2_73 ( .A(_abc_1116_n185), .B(VOTO1_REG), .Y(_abc_1116_n197) );
  AND2X2 AND2X2_74 ( .A(_abc_1116_n173), .B(START), .Y(_abc_1116_n200) );
  AND2X2 AND2X2_75 ( .A(_abc_1116_n201), .B(_abc_1116_n68), .Y(_abc_1116_n202) );
  AND2X2 AND2X2_76 ( .A(_abc_1116_n184), .B(_abc_1116_n203), .Y(_abc_1116_n204) );
  AND2X2 AND2X2_77 ( .A(_abc_1116_n193), .B(V_IN_3_), .Y(_abc_1116_n206) );
  AND2X2 AND2X2_78 ( .A(_abc_1116_n187), .B(VOTO0_REG), .Y(_abc_1116_n207) );
  AND2X2 AND2X2_79 ( .A(_abc_1116_n211), .B(_abc_1116_n91_1), .Y(_abc_1116_n212) );
  AND2X2 AND2X2_8 ( .A(_abc_1116_n66), .B(_abc_1116_n67_1), .Y(_abc_1116_n68) );
  AND2X2 AND2X2_80 ( .A(_abc_1116_n212), .B(_abc_1116_n210), .Y(_abc_1116_n213) );
  AND2X2 AND2X2_81 ( .A(_abc_1116_n205), .B(_abc_1116_n214), .Y(_abc_1116_n215) );
  AND2X2 AND2X2_82 ( .A(_abc_1116_n204), .B(VOTO3_REG), .Y(_abc_1116_n216) );
  AND2X2 AND2X2_83 ( .A(_abc_1116_n172), .B(_abc_1116_n188), .Y(_abc_1116_n219) );
  AND2X2 AND2X2_84 ( .A(_abc_1116_n220), .B(LAST_R_REG), .Y(_abc_1116_n221) );
  AND2X2 AND2X2_85 ( .A(_abc_1116_n219), .B(R_BUTTON), .Y(_abc_1116_n222) );
  AND2X2 AND2X2_86 ( .A(_abc_1116_n225), .B(R_BUTTON), .Y(_abc_1116_n226) );
  AND2X2 AND2X2_87 ( .A(_abc_1116_n227), .B(_abc_1116_n172), .Y(_abc_1116_n228) );
  AND2X2 AND2X2_88 ( .A(_abc_1116_n184), .B(_abc_1116_n229), .Y(_abc_1116_n230) );
  AND2X2 AND2X2_89 ( .A(_abc_1116_n189), .B(_abc_1116_n123), .Y(_abc_1116_n232) );
  AND2X2 AND2X2_9 ( .A(_abc_1116_n68), .B(_abc_1116_n65_1), .Y(_abc_1116_n69_1) );
  AND2X2 AND2X2_90 ( .A(_abc_1116_n193), .B(V_IN_2_), .Y(_abc_1116_n233) );
  AND2X2 AND2X2_91 ( .A(_abc_1116_n231), .B(_abc_1116_n234), .Y(_abc_1116_n235) );
  AND2X2 AND2X2_92 ( .A(_abc_1116_n230), .B(VOTO2_REG), .Y(_abc_1116_n236) );
  AND2X2 AND2X2_93 ( .A(_abc_1116_n220), .B(LAST_G_REG), .Y(_abc_1116_n239) );
  AND2X2 AND2X2_94 ( .A(_abc_1116_n219), .B(G_BUTTON), .Y(_abc_1116_n240) );
  AND2X2 AND2X2_95 ( .A(_abc_1116_n67_1), .B(STATO_REG_1_), .Y(_abc_1116_n245) );
  AND2X2 AND2X2_96 ( .A(_abc_1116_n247), .B(_abc_1116_n244), .Y(_abc_1116_n248) );
  AND2X2 AND2X2_97 ( .A(_abc_1116_n183), .B(_abc_1116_n248), .Y(_abc_1116_n249) );
  AND2X2 AND2X2_98 ( .A(_abc_1116_n193), .B(V_IN_0_), .Y(_abc_1116_n251) );
  AND2X2 AND2X2_99 ( .A(_abc_1116_n69_1), .B(_abc_1116_n188), .Y(_abc_1116_n252) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n105), .Q(CTS_REG) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(n55), .Q(STATO_REG_1_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(n60), .Q(STATO_REG_0_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(n81), .Q(SIGN_REG_3_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(n86), .Q(VOTO1_REG) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(n95), .Q(VOTO3_REG) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(n100), .Q(LAST_R_REG) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(n109), .Q(VOTO2_REG) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(n114), .Q(LAST_G_REG) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n91), .Q(CTR_REG) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n65), .Q(V_OUT_REG_3_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n69), .Q(V_OUT_REG_2_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n73), .Q(V_OUT_REG_1_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n77), .Q(V_OUT_REG_0_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n40), .Q(VOTO0_REG) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n45), .Q(STATO_REG_3_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(n50), .Q(STATO_REG_2_) );
  INVX1 INVX1_1 ( .A(RTS), .Y(_abc_1116_n47) );
  INVX1 INVX1_10 ( .A(START), .Y(_abc_1116_n99_1) );
  INVX1 INVX1_11 ( .A(_abc_1116_n89_1), .Y(_abc_1116_n108) );
  INVX1 INVX1_12 ( .A(_abc_1116_n103), .Y(_abc_1116_n109) );
  INVX1 INVX1_13 ( .A(VOTO0_REG), .Y(_abc_1116_n120) );
  INVX1 INVX1_14 ( .A(_abc_1116_n121), .Y(_abc_1116_n122) );
  INVX1 INVX1_15 ( .A(VOTO2_REG), .Y(_abc_1116_n123) );
  INVX1 INVX1_16 ( .A(_abc_1116_n79), .Y(_abc_1116_n130) );
  INVX1 INVX1_17 ( .A(_abc_1116_n97_1), .Y(_abc_1116_n131) );
  INVX1 INVX1_18 ( .A(_abc_1116_n132), .Y(_abc_1116_n133_1) );
  INVX1 INVX1_19 ( .A(_abc_1116_n125), .Y(_abc_1116_n140_1) );
  INVX1 INVX1_2 ( .A(_abc_1116_n51), .Y(_abc_1116_n52) );
  INVX1 INVX1_20 ( .A(_abc_1116_n88), .Y(_abc_1116_n155_1) );
  INVX1 INVX1_21 ( .A(KEY), .Y(_abc_1116_n173) );
  INVX1 INVX1_22 ( .A(LAST_G_REG), .Y(_abc_1116_n174) );
  INVX1 INVX1_23 ( .A(_abc_1116_n177), .Y(_abc_1116_n178) );
  INVX1 INVX1_24 ( .A(_abc_1116_n179), .Y(_abc_1116_n180) );
  INVX1 INVX1_25 ( .A(_abc_1116_n74), .Y(_abc_1116_n181) );
  INVX1 INVX1_26 ( .A(_abc_1116_n185), .Y(_abc_1116_n186) );
  INVX1 INVX1_27 ( .A(VOTO1_REG), .Y(_abc_1116_n187) );
  INVX1 INVX1_28 ( .A(_abc_1116_n182), .Y(_abc_1116_n191) );
  INVX1 INVX1_29 ( .A(_abc_1116_n202), .Y(_abc_1116_n203) );
  INVX1 INVX1_3 ( .A(TEST), .Y(_abc_1116_n64) );
  INVX1 INVX1_30 ( .A(_abc_1116_n204), .Y(_abc_1116_n205) );
  INVX1 INVX1_31 ( .A(_abc_1116_n208), .Y(_abc_1116_n209) );
  INVX1 INVX1_32 ( .A(_abc_1116_n219), .Y(_abc_1116_n220) );
  INVX1 INVX1_33 ( .A(LAST_R_REG), .Y(_abc_1116_n225) );
  INVX1 INVX1_34 ( .A(_abc_1116_n228), .Y(_abc_1116_n229) );
  INVX1 INVX1_35 ( .A(_abc_1116_n230), .Y(_abc_1116_n231) );
  INVX1 INVX1_36 ( .A(_abc_1116_n96), .Y(_abc_1116_n243) );
  INVX1 INVX1_37 ( .A(_abc_1116_n245), .Y(_abc_1116_n246) );
  INVX1 INVX1_38 ( .A(_abc_1116_n249), .Y(_abc_1116_n250) );
  INVX1 INVX1_39 ( .A(SIGN_REG_3_), .Y(_abc_1116_n253) );
  INVX1 INVX1_4 ( .A(STATO_REG_3_), .Y(_abc_1116_n66) );
  INVX1 INVX1_40 ( .A(_abc_1116_n113_1), .Y(_abc_1116_n263) );
  INVX1 INVX1_5 ( .A(STATO_REG_2_), .Y(_abc_1116_n67_1) );
  INVX1 INVX1_6 ( .A(_abc_1116_n71), .Y(_abc_1116_n72) );
  INVX1 INVX1_7 ( .A(_abc_1116_n77), .Y(_abc_1116_n78) );
  INVX1 INVX1_8 ( .A(_abc_1116_n57), .Y(_abc_1116_n90) );
  INVX1 INVX1_9 ( .A(RTR), .Y(_abc_1116_n92) );
  INVX2 INVX2_1 ( .A(STATO_REG_1_), .Y(_abc_1116_n54) );
  INVX2 INVX2_2 ( .A(STATO_REG_0_), .Y(_abc_1116_n65_1) );
  INVX4 INVX4_1 ( .A(nRESET_G), .Y(_abc_1116_n59) );
  OR2X2 OR2X2_1 ( .A(_abc_1116_n48_1), .B(STATO_REG_0_), .Y(_abc_1116_n49) );
  OR2X2 OR2X2_10 ( .A(_abc_1116_n86), .B(_abc_1116_n88), .Y(_abc_1116_n89_1) );
  OR2X2 OR2X2_11 ( .A(_abc_1116_n61_1), .B(_abc_1116_n94), .Y(_abc_1116_n95_1) );
  OR2X2 OR2X2_12 ( .A(_abc_1116_n98), .B(_abc_1116_n101), .Y(_abc_1116_n102_1) );
  OR2X2 OR2X2_13 ( .A(_abc_1116_n102_1), .B(_abc_1116_n95_1), .Y(_abc_1116_n103) );
  OR2X2 OR2X2_14 ( .A(_abc_1116_n90), .B(_abc_1116_n103), .Y(_abc_1116_n104) );
  OR2X2 OR2X2_15 ( .A(_abc_1116_n104), .B(_abc_1116_n89_1), .Y(_abc_1116_n105) );
  OR2X2 OR2X2_16 ( .A(_abc_1116_n60), .B(_abc_1116_n74), .Y(_abc_1116_n106) );
  OR2X2 OR2X2_17 ( .A(_abc_1116_n115_1), .B(_abc_1116_n59), .Y(_abc_1116_n116) );
  OR2X2 OR2X2_18 ( .A(_abc_1116_n116), .B(_abc_1116_n114), .Y(_abc_1116_n117) );
  OR2X2 OR2X2_19 ( .A(_abc_1116_n112), .B(_abc_1116_n117), .Y(_abc_1116_n118) );
  OR2X2 OR2X2_2 ( .A(STATO_REG_1_), .B(STATO_REG_2_), .Y(_abc_1116_n50) );
  OR2X2 OR2X2_20 ( .A(_abc_1116_n118), .B(_abc_1116_n107), .Y(n55) );
  OR2X2 OR2X2_21 ( .A(_abc_1116_n123), .B(VOTO3_REG), .Y(_abc_1116_n124_1) );
  OR2X2 OR2X2_22 ( .A(_abc_1116_n122), .B(_abc_1116_n124_1), .Y(_abc_1116_n125) );
  OR2X2 OR2X2_23 ( .A(_abc_1116_n126), .B(_abc_1116_n60), .Y(_abc_1116_n127) );
  OR2X2 OR2X2_24 ( .A(_abc_1116_n111), .B(_abc_1116_n127), .Y(_abc_1116_n128) );
  OR2X2 OR2X2_25 ( .A(_abc_1116_n134_1), .B(_abc_1116_n116), .Y(_abc_1116_n135) );
  OR2X2 OR2X2_26 ( .A(_abc_1116_n129), .B(_abc_1116_n135), .Y(n50) );
  OR2X2 OR2X2_27 ( .A(_abc_1116_n111), .B(STATO_REG_0_), .Y(_abc_1116_n137) );
  OR2X2 OR2X2_28 ( .A(_abc_1116_n141), .B(_abc_1116_n71), .Y(_abc_1116_n142) );
  OR2X2 OR2X2_29 ( .A(_abc_1116_n143), .B(_abc_1116_n59), .Y(_abc_1116_n144) );
  OR2X2 OR2X2_3 ( .A(_abc_1116_n53), .B(_abc_1116_n55), .Y(_abc_1116_n56) );
  OR2X2 OR2X2_30 ( .A(_abc_1116_n144), .B(_abc_1116_n138_1), .Y(n45) );
  OR2X2 OR2X2_31 ( .A(_abc_1116_n125), .B(STATO_REG_3_), .Y(_abc_1116_n147) );
  OR2X2 OR2X2_32 ( .A(_abc_1116_n69_1), .B(_abc_1116_n115_1), .Y(_abc_1116_n149) );
  OR2X2 OR2X2_33 ( .A(_abc_1116_n148_1), .B(_abc_1116_n149), .Y(_abc_1116_n150) );
  OR2X2 OR2X2_34 ( .A(_abc_1116_n152), .B(_abc_1116_n59), .Y(_abc_1116_n153) );
  OR2X2 OR2X2_35 ( .A(_abc_1116_n153), .B(_abc_1116_n151), .Y(n60) );
  OR2X2 OR2X2_36 ( .A(_abc_1116_n157), .B(_abc_1116_n59), .Y(_abc_1116_n158) );
  OR2X2 OR2X2_37 ( .A(_abc_1116_n158), .B(_abc_1116_n156_1), .Y(n65) );
  OR2X2 OR2X2_38 ( .A(_abc_1116_n161), .B(_abc_1116_n59), .Y(_abc_1116_n162) );
  OR2X2 OR2X2_39 ( .A(_abc_1116_n162), .B(_abc_1116_n160), .Y(n69) );
  OR2X2 OR2X2_4 ( .A(_abc_1116_n56), .B(_abc_1116_n49), .Y(_abc_1116_n57) );
  OR2X2 OR2X2_40 ( .A(_abc_1116_n165), .B(_abc_1116_n59), .Y(_abc_1116_n166) );
  OR2X2 OR2X2_41 ( .A(_abc_1116_n166), .B(_abc_1116_n164), .Y(n73) );
  OR2X2 OR2X2_42 ( .A(_abc_1116_n169), .B(_abc_1116_n59), .Y(_abc_1116_n170_1) );
  OR2X2 OR2X2_43 ( .A(_abc_1116_n170_1), .B(_abc_1116_n168), .Y(n77) );
  OR2X2 OR2X2_44 ( .A(_abc_1116_n175), .B(_abc_1116_n173), .Y(_abc_1116_n176) );
  OR2X2 OR2X2_45 ( .A(_abc_1116_n181), .B(_abc_1116_n50), .Y(_abc_1116_n182) );
  OR2X2 OR2X2_46 ( .A(_abc_1116_n192), .B(_abc_1116_n191), .Y(_abc_1116_n193) );
  OR2X2 OR2X2_47 ( .A(_abc_1116_n194), .B(_abc_1116_n190), .Y(_abc_1116_n195) );
  OR2X2 OR2X2_48 ( .A(_abc_1116_n197), .B(_abc_1116_n59), .Y(_abc_1116_n198) );
  OR2X2 OR2X2_49 ( .A(_abc_1116_n198), .B(_abc_1116_n196), .Y(n86) );
  OR2X2 OR2X2_5 ( .A(_abc_1116_n61_1), .B(_abc_1116_n59), .Y(_abc_1116_n62) );
  OR2X2 OR2X2_50 ( .A(_abc_1116_n200), .B(_abc_1116_n91_1), .Y(_abc_1116_n201) );
  OR2X2 OR2X2_51 ( .A(_abc_1116_n121), .B(_abc_1116_n207), .Y(_abc_1116_n208) );
  OR2X2 OR2X2_52 ( .A(_abc_1116_n209), .B(_abc_1116_n123), .Y(_abc_1116_n210) );
  OR2X2 OR2X2_53 ( .A(_abc_1116_n208), .B(VOTO2_REG), .Y(_abc_1116_n211) );
  OR2X2 OR2X2_54 ( .A(_abc_1116_n213), .B(_abc_1116_n206), .Y(_abc_1116_n214) );
  OR2X2 OR2X2_55 ( .A(_abc_1116_n216), .B(_abc_1116_n59), .Y(_abc_1116_n217) );
  OR2X2 OR2X2_56 ( .A(_abc_1116_n217), .B(_abc_1116_n215), .Y(n95) );
  OR2X2 OR2X2_57 ( .A(_abc_1116_n222), .B(_abc_1116_n59), .Y(_abc_1116_n223) );
  OR2X2 OR2X2_58 ( .A(_abc_1116_n223), .B(_abc_1116_n221), .Y(n100) );
  OR2X2 OR2X2_59 ( .A(_abc_1116_n226), .B(_abc_1116_n173), .Y(_abc_1116_n227) );
  OR2X2 OR2X2_6 ( .A(_abc_1116_n58), .B(_abc_1116_n62), .Y(n91) );
  OR2X2 OR2X2_60 ( .A(_abc_1116_n233), .B(_abc_1116_n232), .Y(_abc_1116_n234) );
  OR2X2 OR2X2_61 ( .A(_abc_1116_n236), .B(_abc_1116_n59), .Y(_abc_1116_n237) );
  OR2X2 OR2X2_62 ( .A(_abc_1116_n237), .B(_abc_1116_n235), .Y(n109) );
  OR2X2 OR2X2_63 ( .A(_abc_1116_n240), .B(_abc_1116_n59), .Y(_abc_1116_n241) );
  OR2X2 OR2X2_64 ( .A(_abc_1116_n241), .B(_abc_1116_n239), .Y(n114) );
  OR2X2 OR2X2_65 ( .A(_abc_1116_n243), .B(STATO_REG_3_), .Y(_abc_1116_n244) );
  OR2X2 OR2X2_66 ( .A(_abc_1116_n132), .B(_abc_1116_n246), .Y(_abc_1116_n247) );
  OR2X2 OR2X2_67 ( .A(_abc_1116_n252), .B(_abc_1116_n255), .Y(_abc_1116_n256) );
  OR2X2 OR2X2_68 ( .A(_abc_1116_n251), .B(_abc_1116_n256), .Y(_abc_1116_n257) );
  OR2X2 OR2X2_69 ( .A(_abc_1116_n259), .B(_abc_1116_n59), .Y(_abc_1116_n260) );
  OR2X2 OR2X2_7 ( .A(_abc_1116_n74), .B(_abc_1116_n59), .Y(_abc_1116_n75) );
  OR2X2 OR2X2_70 ( .A(_abc_1116_n260), .B(_abc_1116_n258), .Y(n40) );
  OR2X2 OR2X2_71 ( .A(_abc_1116_n264), .B(_abc_1116_n262), .Y(_abc_1116_n265) );
  OR2X2 OR2X2_72 ( .A(_abc_1116_n53), .B(_abc_1116_n87_1), .Y(_abc_1116_n266) );
  OR2X2 OR2X2_73 ( .A(_abc_1116_n265), .B(_abc_1116_n266), .Y(_abc_1116_n267) );
  OR2X2 OR2X2_74 ( .A(_abc_1116_n269), .B(_abc_1116_n139), .Y(_abc_1116_n270) );
  OR2X2 OR2X2_75 ( .A(_abc_1116_n272), .B(_abc_1116_n59), .Y(_abc_1116_n273) );
  OR2X2 OR2X2_76 ( .A(_abc_1116_n271), .B(_abc_1116_n273), .Y(_abc_1116_n274) );
  OR2X2 OR2X2_77 ( .A(_abc_1116_n268), .B(_abc_1116_n274), .Y(n105) );
  OR2X2 OR2X2_8 ( .A(_abc_1116_n73), .B(_abc_1116_n75), .Y(n81) );
  OR2X2 OR2X2_9 ( .A(_abc_1116_n81_1), .B(_abc_1116_n85), .Y(_abc_1116_n86) );
endmodule