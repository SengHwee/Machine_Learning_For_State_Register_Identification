module b02_reset(clock, RESET_G, nRESET_G, LINEA, U_REG);
  input LINEA;
  input RESET_G;
  wire STATO_REG_0_;
  wire STATO_REG_1_;
  wire STATO_REG_2_;
  output U_REG;
  wire _abc_181_n10_1;
  wire _abc_181_n11;
  wire _abc_181_n12;
  wire _abc_181_n13;
  wire _abc_181_n15_1;
  wire _abc_181_n16;
  wire _abc_181_n17;
  wire _abc_181_n18;
  wire _abc_181_n19;
  wire _abc_181_n20;
  wire _abc_181_n21_1;
  wire _abc_181_n22;
  wire _abc_181_n23;
  wire _abc_181_n25_1;
  wire _abc_181_n26;
  wire _abc_181_n27;
  wire _abc_181_n28;
  wire _abc_181_n29;
  wire _abc_181_n30;
  wire _abc_181_n31;
  wire _abc_181_n33;
  wire _abc_181_n34;
  wire _abc_181_n35;
  wire _abc_181_n36;
  wire _abc_181_n37;
  wire _abc_181_n38;
  input clock;
  wire n10;
  wire n14;
  wire n19;
  wire n24;
  input nRESET_G;
  AND2X2 AND2X2_1 ( .A(_abc_181_n10_1), .B(nRESET_G), .Y(_abc_181_n11) );
  AND2X2 AND2X2_10 ( .A(_abc_181_n12), .B(_abc_181_n25_1), .Y(_abc_181_n33) );
  AND2X2 AND2X2_11 ( .A(_abc_181_n34), .B(STATO_REG_0_), .Y(_abc_181_n35) );
  AND2X2 AND2X2_12 ( .A(_abc_181_n15_1), .B(STATO_REG_1_), .Y(_abc_181_n36) );
  AND2X2 AND2X2_13 ( .A(_abc_181_n36), .B(_abc_181_n10_1), .Y(_abc_181_n37) );
  AND2X2 AND2X2_2 ( .A(_abc_181_n12), .B(STATO_REG_2_), .Y(_abc_181_n13) );
  AND2X2 AND2X2_3 ( .A(_abc_181_n11), .B(_abc_181_n13), .Y(n10) );
  AND2X2 AND2X2_4 ( .A(_abc_181_n15_1), .B(LINEA), .Y(_abc_181_n16) );
  AND2X2 AND2X2_5 ( .A(_abc_181_n17), .B(_abc_181_n12), .Y(_abc_181_n18) );
  AND2X2 AND2X2_6 ( .A(_abc_181_n21_1), .B(_abc_181_n10_1), .Y(_abc_181_n22) );
  AND2X2 AND2X2_7 ( .A(_abc_181_n25_1), .B(STATO_REG_2_), .Y(_abc_181_n26) );
  AND2X2 AND2X2_8 ( .A(_abc_181_n20), .B(STATO_REG_0_), .Y(_abc_181_n29) );
  AND2X2 AND2X2_9 ( .A(_abc_181_n28), .B(_abc_181_n30), .Y(_abc_181_n31) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n10), .Q(U_REG) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n14), .Q(STATO_REG_2_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n19), .Q(STATO_REG_1_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n24), .Q(STATO_REG_0_) );
  INVX1 INVX1_1 ( .A(STATO_REG_0_), .Y(_abc_181_n10_1) );
  INVX1 INVX1_2 ( .A(STATO_REG_1_), .Y(_abc_181_n12) );
  INVX1 INVX1_3 ( .A(STATO_REG_2_), .Y(_abc_181_n15_1) );
  INVX1 INVX1_4 ( .A(nRESET_G), .Y(_abc_181_n19) );
  INVX1 INVX1_5 ( .A(_abc_181_n20), .Y(_abc_181_n21_1) );
  INVX1 INVX1_6 ( .A(LINEA), .Y(_abc_181_n25_1) );
  OR2X2 OR2X2_1 ( .A(_abc_181_n16), .B(_abc_181_n10_1), .Y(_abc_181_n17) );
  OR2X2 OR2X2_10 ( .A(_abc_181_n37), .B(_abc_181_n19), .Y(_abc_181_n38) );
  OR2X2 OR2X2_11 ( .A(_abc_181_n35), .B(_abc_181_n38), .Y(n19) );
  OR2X2 OR2X2_2 ( .A(STATO_REG_2_), .B(LINEA), .Y(_abc_181_n20) );
  OR2X2 OR2X2_3 ( .A(_abc_181_n22), .B(_abc_181_n19), .Y(_abc_181_n23) );
  OR2X2 OR2X2_4 ( .A(_abc_181_n23), .B(_abc_181_n18), .Y(n24) );
  OR2X2 OR2X2_5 ( .A(_abc_181_n16), .B(STATO_REG_0_), .Y(_abc_181_n27) );
  OR2X2 OR2X2_6 ( .A(_abc_181_n27), .B(_abc_181_n26), .Y(_abc_181_n28) );
  OR2X2 OR2X2_7 ( .A(_abc_181_n29), .B(STATO_REG_1_), .Y(_abc_181_n30) );
  OR2X2 OR2X2_8 ( .A(_abc_181_n31), .B(_abc_181_n19), .Y(n14) );
  OR2X2 OR2X2_9 ( .A(_abc_181_n33), .B(STATO_REG_2_), .Y(_abc_181_n34) );
endmodule