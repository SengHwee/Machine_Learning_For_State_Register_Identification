module MEMORY_INTERFACE(clock, resetn, \rs1[0] , \rs1[1] , \rs1[2] , \rs1[3] , \rs1[4] , \rs1[5] , \rs1[6] , \rs1[7] , \rs1[8] , \rs1[9] , \rs1[10] , \rs1[11] , \rs1[12] , \rs1[13] , \rs1[14] , \rs1[15] , \rs1[16] , \rs1[17] , \rs1[18] , \rs1[19] , \rs1[20] , \rs1[21] , \rs1[22] , \rs1[23] , \rs1[24] , \rs1[25] , \rs1[26] , \rs1[27] , \rs1[28] , \rs1[29] , \rs1[30] , \rs1[31] , \rs2[0] , \rs2[1] , \rs2[2] , \rs2[3] , \rs2[4] , \rs2[5] , \rs2[6] , \rs2[7] , \rs2[8] , \rs2[9] , \rs2[10] , \rs2[11] , \rs2[12] , \rs2[13] , \rs2[14] , \rs2[15] , \rs2[16] , \rs2[17] , \rs2[18] , \rs2[19] , \rs2[20] , \rs2[21] , \rs2[22] , \rs2[23] , \rs2[24] , \rs2[25] , \rs2[26] , \rs2[27] , \rs2[28] , \rs2[29] , \rs2[30] , \rs2[31] , \Rdata_mem[0] , \Rdata_mem[1] , \Rdata_mem[2] , \Rdata_mem[3] , \Rdata_mem[4] , \Rdata_mem[5] , \Rdata_mem[6] , \Rdata_mem[7] , \Rdata_mem[8] , \Rdata_mem[9] , \Rdata_mem[10] , \Rdata_mem[11] , \Rdata_mem[12] , \Rdata_mem[13] , \Rdata_mem[14] , \Rdata_mem[15] , \Rdata_mem[16] , \Rdata_mem[17] , \Rdata_mem[18] , \Rdata_mem[19] , \Rdata_mem[20] , \Rdata_mem[21] , \Rdata_mem[22] , \Rdata_mem[23] , \Rdata_mem[24] , \Rdata_mem[25] , \Rdata_mem[26] , \Rdata_mem[27] , \Rdata_mem[28] , \Rdata_mem[29] , \Rdata_mem[30] , \Rdata_mem[31] , ARready, Rvalid, AWready, Wready, Bvalid, \imm[0] , \imm[1] , \imm[2] , \imm[3] , \imm[4] , \imm[5] , \imm[6] , \imm[7] , \imm[8] , \imm[9] , \imm[10] , \imm[11] , \imm[12] , \imm[13] , \imm[14] , \imm[15] , \imm[16] , \imm[17] , \imm[18] , \imm[19] , \imm[20] , \imm[21] , \imm[22] , \imm[23] , \imm[24] , \imm[25] , \imm[26] , \imm[27] , \imm[28] , \imm[29] , \imm[30] , \imm[31] , \W_R[0] , \W_R[1] , \wordsize[0] , \wordsize[1] , enable, \pc[0] , \pc[1] , \pc[2] , \pc[3] , \pc[4] , \pc[5] , \pc[6] , \pc[7] , \pc[8] , \pc[9] , \pc[10] , \pc[11] , \pc[12] , \pc[13] , \pc[14] , \pc[15] , \pc[16] , \pc[17] , \pc[18] , \pc[19] , \pc[20] , \pc[21] , \pc[22] , \pc[23] , \pc[24] , \pc[25] , \pc[26] , \pc[27] , \pc[28] , \pc[29] , \pc[30] , \pc[31] , signo, busy, done, align, \AWdata[0] , \AWdata[1] , \AWdata[2] , \AWdata[3] , \AWdata[4] , \AWdata[5] , \AWdata[6] , \AWdata[7] , \AWdata[8] , \AWdata[9] , \AWdata[10] , \AWdata[11] , \AWdata[12] , \AWdata[13] , \AWdata[14] , \AWdata[15] , \AWdata[16] , \AWdata[17] , \AWdata[18] , \AWdata[19] , \AWdata[20] , \AWdata[21] , \AWdata[22] , \AWdata[23] , \AWdata[24] , \AWdata[25] , \AWdata[26] , \AWdata[27] , \AWdata[28] , \AWdata[29] , \AWdata[30] , \AWdata[31] , \ARdata[0] , \ARdata[1] , \ARdata[2] , \ARdata[3] , \ARdata[4] , \ARdata[5] , \ARdata[6] , \ARdata[7] , \ARdata[8] , \ARdata[9] , \ARdata[10] , \ARdata[11] , \ARdata[12] , \ARdata[13] , \ARdata[14] , \ARdata[15] , \ARdata[16] , \ARdata[17] , \ARdata[18] , \ARdata[19] , \ARdata[20] , \ARdata[21] , \ARdata[22] , \ARdata[23] , \ARdata[24] , \ARdata[25] , \ARdata[26] , \ARdata[27] , \ARdata[28] , \ARdata[29] , \ARdata[30] , \ARdata[31] , \Wdata[0] , \Wdata[1] , \Wdata[2] , \Wdata[3] , \Wdata[4] , \Wdata[5] , \Wdata[6] , \Wdata[7] , \Wdata[8] , \Wdata[9] , \Wdata[10] , \Wdata[11] , \Wdata[12] , \Wdata[13] , \Wdata[14] , \Wdata[15] , \Wdata[16] , \Wdata[17] , \Wdata[18] , \Wdata[19] , \Wdata[20] , \Wdata[21] , \Wdata[22] , \Wdata[23] , \Wdata[24] , \Wdata[25] , \Wdata[26] , \Wdata[27] , \Wdata[28] , \Wdata[29] , \Wdata[30] , \Wdata[31] , \rd[0] , \rd[1] , \rd[2] , \rd[3] , \rd[4] , \rd[5] , \rd[6] , \rd[7] , \rd[8] , \rd[9] , \rd[10] , \rd[11] , \rd[12] , \rd[13] , \rd[14] , \rd[15] , \rd[16] , \rd[17] , \rd[18] , \rd[19] , \rd[20] , \rd[21] , \rd[22] , \rd[23] , \rd[24] , \rd[25] , \rd[26] , \rd[27] , \rd[28] , \rd[29] , \rd[30] , \rd[31] , \inst[0] , \inst[1] , \inst[2] , \inst[3] , \inst[4] , \inst[5] , \inst[6] , \inst[7] , \inst[8] , \inst[9] , \inst[10] , \inst[11] , \inst[12] , \inst[13] , \inst[14] , \inst[15] , \inst[16] , \inst[17] , \inst[18] , \inst[19] , \inst[20] , \inst[21] , \inst[22] , \inst[23] , \inst[24] , \inst[25] , \inst[26] , \inst[27] , \inst[28] , \inst[29] , \inst[30] , \inst[31] , ARvalid, RReady, AWvalid, Wvalid, \arprot[0] , \arprot[1] , \arprot[2] , \awprot[0] , \awprot[1] , \awprot[2] , Bready, \Wstrb[0] , \Wstrb[1] , \Wstrb[2] , \Wstrb[3] , rd_en);

output \ARdata[0] ;
output \ARdata[10] ;
output \ARdata[11] ;
output \ARdata[12] ;
output \ARdata[13] ;
output \ARdata[14] ;
output \ARdata[15] ;
output \ARdata[16] ;
output \ARdata[17] ;
output \ARdata[18] ;
output \ARdata[19] ;
output \ARdata[1] ;
output \ARdata[20] ;
output \ARdata[21] ;
output \ARdata[22] ;
output \ARdata[23] ;
output \ARdata[24] ;
output \ARdata[25] ;
output \ARdata[26] ;
output \ARdata[27] ;
output \ARdata[28] ;
output \ARdata[29] ;
output \ARdata[2] ;
output \ARdata[30] ;
output \ARdata[31] ;
output \ARdata[3] ;
output \ARdata[4] ;
output \ARdata[5] ;
output \ARdata[6] ;
output \ARdata[7] ;
output \ARdata[8] ;
output \ARdata[9] ;
input ARready;
output ARvalid;
output \AWdata[0] ;
output \AWdata[10] ;
output \AWdata[11] ;
output \AWdata[12] ;
output \AWdata[13] ;
output \AWdata[14] ;
output \AWdata[15] ;
output \AWdata[16] ;
output \AWdata[17] ;
output \AWdata[18] ;
output \AWdata[19] ;
output \AWdata[1] ;
output \AWdata[20] ;
output \AWdata[21] ;
output \AWdata[22] ;
output \AWdata[23] ;
output \AWdata[24] ;
output \AWdata[25] ;
output \AWdata[26] ;
output \AWdata[27] ;
output \AWdata[28] ;
output \AWdata[29] ;
output \AWdata[2] ;
output \AWdata[30] ;
output \AWdata[31] ;
output \AWdata[3] ;
output \AWdata[4] ;
output \AWdata[5] ;
output \AWdata[6] ;
output \AWdata[7] ;
output \AWdata[8] ;
output \AWdata[9] ;
input AWready;
output AWvalid;
output Bready;
input Bvalid;
output RReady;
input \Rdata_mem[0] ;
input \Rdata_mem[10] ;
input \Rdata_mem[11] ;
input \Rdata_mem[12] ;
input \Rdata_mem[13] ;
input \Rdata_mem[14] ;
input \Rdata_mem[15] ;
input \Rdata_mem[16] ;
input \Rdata_mem[17] ;
input \Rdata_mem[18] ;
input \Rdata_mem[19] ;
input \Rdata_mem[1] ;
input \Rdata_mem[20] ;
input \Rdata_mem[21] ;
input \Rdata_mem[22] ;
input \Rdata_mem[23] ;
input \Rdata_mem[24] ;
input \Rdata_mem[25] ;
input \Rdata_mem[26] ;
input \Rdata_mem[27] ;
input \Rdata_mem[28] ;
input \Rdata_mem[29] ;
input \Rdata_mem[2] ;
input \Rdata_mem[30] ;
input \Rdata_mem[31] ;
input \Rdata_mem[3] ;
input \Rdata_mem[4] ;
input \Rdata_mem[5] ;
input \Rdata_mem[6] ;
input \Rdata_mem[7] ;
input \Rdata_mem[8] ;
input \Rdata_mem[9] ;
input Rvalid;
input \W_R[0] ;
input \W_R[1] ;
wire W_R_1_bF_buf0_; 
wire W_R_1_bF_buf1_; 
wire W_R_1_bF_buf2_; 
wire W_R_1_bF_buf3_; 
wire W_R_1_bF_buf4_; 
wire W_R_1_bF_buf5_; 
output \Wdata[0] ;
output \Wdata[10] ;
output \Wdata[11] ;
output \Wdata[12] ;
output \Wdata[13] ;
output \Wdata[14] ;
output \Wdata[15] ;
output \Wdata[16] ;
output \Wdata[17] ;
output \Wdata[18] ;
output \Wdata[19] ;
output \Wdata[1] ;
output \Wdata[20] ;
output \Wdata[21] ;
output \Wdata[22] ;
output \Wdata[23] ;
output \Wdata[24] ;
output \Wdata[25] ;
output \Wdata[26] ;
output \Wdata[27] ;
output \Wdata[28] ;
output \Wdata[29] ;
output \Wdata[2] ;
output \Wdata[30] ;
output \Wdata[31] ;
output \Wdata[3] ;
output \Wdata[4] ;
output \Wdata[5] ;
output \Wdata[6] ;
output \Wdata[7] ;
output \Wdata[8] ;
output \Wdata[9] ;
input Wready;
output \Wstrb[0] ;
output \Wstrb[1] ;
output \Wstrb[2] ;
output \Wstrb[3] ;
output Wvalid;
wire _0Wdata_31_0__0_; 
wire _0Wdata_31_0__10_; 
wire _0Wdata_31_0__11_; 
wire _0Wdata_31_0__12_; 
wire _0Wdata_31_0__13_; 
wire _0Wdata_31_0__14_; 
wire _0Wdata_31_0__15_; 
wire _0Wdata_31_0__16_; 
wire _0Wdata_31_0__17_; 
wire _0Wdata_31_0__18_; 
wire _0Wdata_31_0__19_; 
wire _0Wdata_31_0__1_; 
wire _0Wdata_31_0__20_; 
wire _0Wdata_31_0__21_; 
wire _0Wdata_31_0__22_; 
wire _0Wdata_31_0__23_; 
wire _0Wdata_31_0__24_; 
wire _0Wdata_31_0__25_; 
wire _0Wdata_31_0__26_; 
wire _0Wdata_31_0__27_; 
wire _0Wdata_31_0__28_; 
wire _0Wdata_31_0__29_; 
wire _0Wdata_31_0__2_; 
wire _0Wdata_31_0__30_; 
wire _0Wdata_31_0__31_; 
wire _0Wdata_31_0__3_; 
wire _0Wdata_31_0__4_; 
wire _0Wdata_31_0__5_; 
wire _0Wdata_31_0__6_; 
wire _0Wdata_31_0__7_; 
wire _0Wdata_31_0__8_; 
wire _0Wdata_31_0__9_; 
wire _0Wstrb_3_0__0_; 
wire _0Wstrb_3_0__1_; 
wire _0Wstrb_3_0__2_; 
wire _0Wstrb_3_0__3_; 
wire _0inst_31_0__0_; 
wire _0inst_31_0__10_; 
wire _0inst_31_0__11_; 
wire _0inst_31_0__12_; 
wire _0inst_31_0__13_; 
wire _0inst_31_0__14_; 
wire _0inst_31_0__15_; 
wire _0inst_31_0__16_; 
wire _0inst_31_0__17_; 
wire _0inst_31_0__18_; 
wire _0inst_31_0__19_; 
wire _0inst_31_0__1_; 
wire _0inst_31_0__20_; 
wire _0inst_31_0__21_; 
wire _0inst_31_0__22_; 
wire _0inst_31_0__23_; 
wire _0inst_31_0__24_; 
wire _0inst_31_0__25_; 
wire _0inst_31_0__26_; 
wire _0inst_31_0__27_; 
wire _0inst_31_0__28_; 
wire _0inst_31_0__29_; 
wire _0inst_31_0__2_; 
wire _0inst_31_0__30_; 
wire _0inst_31_0__31_; 
wire _0inst_31_0__3_; 
wire _0inst_31_0__4_; 
wire _0inst_31_0__5_; 
wire _0inst_31_0__6_; 
wire _0inst_31_0__7_; 
wire _0inst_31_0__8_; 
wire _0inst_31_0__9_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_0_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_1_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_2_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_3_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_4_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_5_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_6_; 
wire _abc_4635_new_n1000_; 
wire _abc_4635_new_n1001_; 
wire _abc_4635_new_n1002_; 
wire _abc_4635_new_n1003_; 
wire _abc_4635_new_n1004_; 
wire _abc_4635_new_n1006_; 
wire _abc_4635_new_n1007_; 
wire _abc_4635_new_n1008_; 
wire _abc_4635_new_n1009_; 
wire _abc_4635_new_n1010_; 
wire _abc_4635_new_n1011_; 
wire _abc_4635_new_n1012_; 
wire _abc_4635_new_n1013_; 
wire _abc_4635_new_n1014_; 
wire _abc_4635_new_n1015_; 
wire _abc_4635_new_n1016_; 
wire _abc_4635_new_n1017_; 
wire _abc_4635_new_n1019_; 
wire _abc_4635_new_n1020_; 
wire _abc_4635_new_n1021_; 
wire _abc_4635_new_n1022_; 
wire _abc_4635_new_n1023_; 
wire _abc_4635_new_n1024_; 
wire _abc_4635_new_n1025_; 
wire _abc_4635_new_n1026_; 
wire _abc_4635_new_n1027_; 
wire _abc_4635_new_n1028_; 
wire _abc_4635_new_n1029_; 
wire _abc_4635_new_n1030_; 
wire _abc_4635_new_n1031_; 
wire _abc_4635_new_n1032_; 
wire _abc_4635_new_n1033_; 
wire _abc_4635_new_n1035_; 
wire _abc_4635_new_n1036_; 
wire _abc_4635_new_n1037_; 
wire _abc_4635_new_n1038_; 
wire _abc_4635_new_n1039_; 
wire _abc_4635_new_n1040_; 
wire _abc_4635_new_n1041_; 
wire _abc_4635_new_n1042_; 
wire _abc_4635_new_n1043_; 
wire _abc_4635_new_n1044_; 
wire _abc_4635_new_n1045_; 
wire _abc_4635_new_n1046_; 
wire _abc_4635_new_n1048_; 
wire _abc_4635_new_n1049_; 
wire _abc_4635_new_n1050_; 
wire _abc_4635_new_n1051_; 
wire _abc_4635_new_n1052_; 
wire _abc_4635_new_n1053_; 
wire _abc_4635_new_n1054_; 
wire _abc_4635_new_n1055_; 
wire _abc_4635_new_n1056_; 
wire _abc_4635_new_n1057_; 
wire _abc_4635_new_n1058_; 
wire _abc_4635_new_n1059_; 
wire _abc_4635_new_n1060_; 
wire _abc_4635_new_n1061_; 
wire _abc_4635_new_n1062_; 
wire _abc_4635_new_n1064_; 
wire _abc_4635_new_n1065_; 
wire _abc_4635_new_n1066_; 
wire _abc_4635_new_n1067_; 
wire _abc_4635_new_n1068_; 
wire _abc_4635_new_n1069_; 
wire _abc_4635_new_n1070_; 
wire _abc_4635_new_n1071_; 
wire _abc_4635_new_n1072_; 
wire _abc_4635_new_n1073_; 
wire _abc_4635_new_n1074_; 
wire _abc_4635_new_n1075_; 
wire _abc_4635_new_n1077_; 
wire _abc_4635_new_n1078_; 
wire _abc_4635_new_n1079_; 
wire _abc_4635_new_n1080_; 
wire _abc_4635_new_n1081_; 
wire _abc_4635_new_n1082_; 
wire _abc_4635_new_n1083_; 
wire _abc_4635_new_n1084_; 
wire _abc_4635_new_n1085_; 
wire _abc_4635_new_n1086_; 
wire _abc_4635_new_n1087_; 
wire _abc_4635_new_n1088_; 
wire _abc_4635_new_n1089_; 
wire _abc_4635_new_n1090_; 
wire _abc_4635_new_n1091_; 
wire _abc_4635_new_n1092_; 
wire _abc_4635_new_n1093_; 
wire _abc_4635_new_n1094_; 
wire _abc_4635_new_n1096_; 
wire _abc_4635_new_n1097_; 
wire _abc_4635_new_n1098_; 
wire _abc_4635_new_n1099_; 
wire _abc_4635_new_n1100_; 
wire _abc_4635_new_n1101_; 
wire _abc_4635_new_n1102_; 
wire _abc_4635_new_n1103_; 
wire _abc_4635_new_n1104_; 
wire _abc_4635_new_n1105_; 
wire _abc_4635_new_n1106_; 
wire _abc_4635_new_n1107_; 
wire _abc_4635_new_n1109_; 
wire _abc_4635_new_n1110_; 
wire _abc_4635_new_n1111_; 
wire _abc_4635_new_n1112_; 
wire _abc_4635_new_n1113_; 
wire _abc_4635_new_n1114_; 
wire _abc_4635_new_n1115_; 
wire _abc_4635_new_n1116_; 
wire _abc_4635_new_n1117_; 
wire _abc_4635_new_n1118_; 
wire _abc_4635_new_n1119_; 
wire _abc_4635_new_n1120_; 
wire _abc_4635_new_n1121_; 
wire _abc_4635_new_n1122_; 
wire _abc_4635_new_n1123_; 
wire _abc_4635_new_n1125_; 
wire _abc_4635_new_n1126_; 
wire _abc_4635_new_n1127_; 
wire _abc_4635_new_n1128_; 
wire _abc_4635_new_n1129_; 
wire _abc_4635_new_n1130_; 
wire _abc_4635_new_n1131_; 
wire _abc_4635_new_n1132_; 
wire _abc_4635_new_n1133_; 
wire _abc_4635_new_n1134_; 
wire _abc_4635_new_n1135_; 
wire _abc_4635_new_n1136_; 
wire _abc_4635_new_n1138_; 
wire _abc_4635_new_n1139_; 
wire _abc_4635_new_n1140_; 
wire _abc_4635_new_n1141_; 
wire _abc_4635_new_n1142_; 
wire _abc_4635_new_n1143_; 
wire _abc_4635_new_n1144_; 
wire _abc_4635_new_n1145_; 
wire _abc_4635_new_n1146_; 
wire _abc_4635_new_n1147_; 
wire _abc_4635_new_n1148_; 
wire _abc_4635_new_n1149_; 
wire _abc_4635_new_n1150_; 
wire _abc_4635_new_n1151_; 
wire _abc_4635_new_n1152_; 
wire _abc_4635_new_n1153_; 
wire _abc_4635_new_n1154_; 
wire _abc_4635_new_n1155_; 
wire _abc_4635_new_n1157_; 
wire _abc_4635_new_n1158_; 
wire _abc_4635_new_n1159_; 
wire _abc_4635_new_n1160_; 
wire _abc_4635_new_n1161_; 
wire _abc_4635_new_n1162_; 
wire _abc_4635_new_n1163_; 
wire _abc_4635_new_n1164_; 
wire _abc_4635_new_n1165_; 
wire _abc_4635_new_n1166_; 
wire _abc_4635_new_n1167_; 
wire _abc_4635_new_n1168_; 
wire _abc_4635_new_n1170_; 
wire _abc_4635_new_n1171_; 
wire _abc_4635_new_n1172_; 
wire _abc_4635_new_n1173_; 
wire _abc_4635_new_n1174_; 
wire _abc_4635_new_n1175_; 
wire _abc_4635_new_n1176_; 
wire _abc_4635_new_n1177_; 
wire _abc_4635_new_n1178_; 
wire _abc_4635_new_n1179_; 
wire _abc_4635_new_n1180_; 
wire _abc_4635_new_n1181_; 
wire _abc_4635_new_n1182_; 
wire _abc_4635_new_n1183_; 
wire _abc_4635_new_n1184_; 
wire _abc_4635_new_n1185_; 
wire _abc_4635_new_n1187_; 
wire _abc_4635_new_n1188_; 
wire _abc_4635_new_n1189_; 
wire _abc_4635_new_n1190_; 
wire _abc_4635_new_n1191_; 
wire _abc_4635_new_n1192_; 
wire _abc_4635_new_n1193_; 
wire _abc_4635_new_n1194_; 
wire _abc_4635_new_n1195_; 
wire _abc_4635_new_n1196_; 
wire _abc_4635_new_n1197_; 
wire _abc_4635_new_n1198_; 
wire _abc_4635_new_n1200_; 
wire _abc_4635_new_n1201_; 
wire _abc_4635_new_n1202_; 
wire _abc_4635_new_n1203_; 
wire _abc_4635_new_n1204_; 
wire _abc_4635_new_n1205_; 
wire _abc_4635_new_n1206_; 
wire _abc_4635_new_n1207_; 
wire _abc_4635_new_n1208_; 
wire _abc_4635_new_n1209_; 
wire _abc_4635_new_n1210_; 
wire _abc_4635_new_n1211_; 
wire _abc_4635_new_n1212_; 
wire _abc_4635_new_n1213_; 
wire _abc_4635_new_n1214_; 
wire _abc_4635_new_n1215_; 
wire _abc_4635_new_n1216_; 
wire _abc_4635_new_n1217_; 
wire _abc_4635_new_n1218_; 
wire _abc_4635_new_n1219_; 
wire _abc_4635_new_n1220_; 
wire _abc_4635_new_n1222_; 
wire _abc_4635_new_n1223_; 
wire _abc_4635_new_n1224_; 
wire _abc_4635_new_n1225_; 
wire _abc_4635_new_n1226_; 
wire _abc_4635_new_n1227_; 
wire _abc_4635_new_n1228_; 
wire _abc_4635_new_n1229_; 
wire _abc_4635_new_n1230_; 
wire _abc_4635_new_n1231_; 
wire _abc_4635_new_n1232_; 
wire _abc_4635_new_n1233_; 
wire _abc_4635_new_n1235_; 
wire _abc_4635_new_n1236_; 
wire _abc_4635_new_n1237_; 
wire _abc_4635_new_n1238_; 
wire _abc_4635_new_n1239_; 
wire _abc_4635_new_n1240_; 
wire _abc_4635_new_n1241_; 
wire _abc_4635_new_n1242_; 
wire _abc_4635_new_n1243_; 
wire _abc_4635_new_n1244_; 
wire _abc_4635_new_n1245_; 
wire _abc_4635_new_n1246_; 
wire _abc_4635_new_n1247_; 
wire _abc_4635_new_n1248_; 
wire _abc_4635_new_n1249_; 
wire _abc_4635_new_n1250_; 
wire _abc_4635_new_n1252_; 
wire _abc_4635_new_n1253_; 
wire _abc_4635_new_n1254_; 
wire _abc_4635_new_n1255_; 
wire _abc_4635_new_n1256_; 
wire _abc_4635_new_n1257_; 
wire _abc_4635_new_n1258_; 
wire _abc_4635_new_n1259_; 
wire _abc_4635_new_n1260_; 
wire _abc_4635_new_n1261_; 
wire _abc_4635_new_n1262_; 
wire _abc_4635_new_n1263_; 
wire _abc_4635_new_n1265_; 
wire _abc_4635_new_n1266_; 
wire _abc_4635_new_n1267_; 
wire _abc_4635_new_n1268_; 
wire _abc_4635_new_n1269_; 
wire _abc_4635_new_n1270_; 
wire _abc_4635_new_n1271_; 
wire _abc_4635_new_n1272_; 
wire _abc_4635_new_n1273_; 
wire _abc_4635_new_n1274_; 
wire _abc_4635_new_n1275_; 
wire _abc_4635_new_n1276_; 
wire _abc_4635_new_n1277_; 
wire _abc_4635_new_n1278_; 
wire _abc_4635_new_n1279_; 
wire _abc_4635_new_n1280_; 
wire _abc_4635_new_n1281_; 
wire _abc_4635_new_n1282_; 
wire _abc_4635_new_n1284_; 
wire _abc_4635_new_n1285_; 
wire _abc_4635_new_n1286_; 
wire _abc_4635_new_n1287_; 
wire _abc_4635_new_n1288_; 
wire _abc_4635_new_n1289_; 
wire _abc_4635_new_n1290_; 
wire _abc_4635_new_n1291_; 
wire _abc_4635_new_n1292_; 
wire _abc_4635_new_n1293_; 
wire _abc_4635_new_n1294_; 
wire _abc_4635_new_n1295_; 
wire _abc_4635_new_n1297_; 
wire _abc_4635_new_n1298_; 
wire _abc_4635_new_n1299_; 
wire _abc_4635_new_n1300_; 
wire _abc_4635_new_n1301_; 
wire _abc_4635_new_n1302_; 
wire _abc_4635_new_n1303_; 
wire _abc_4635_new_n1304_; 
wire _abc_4635_new_n1305_; 
wire _abc_4635_new_n1306_; 
wire _abc_4635_new_n1307_; 
wire _abc_4635_new_n1308_; 
wire _abc_4635_new_n1309_; 
wire _abc_4635_new_n1310_; 
wire _abc_4635_new_n1311_; 
wire _abc_4635_new_n1312_; 
wire _abc_4635_new_n1314_; 
wire _abc_4635_new_n1315_; 
wire _abc_4635_new_n1316_; 
wire _abc_4635_new_n1317_; 
wire _abc_4635_new_n1318_; 
wire _abc_4635_new_n1319_; 
wire _abc_4635_new_n1320_; 
wire _abc_4635_new_n1321_; 
wire _abc_4635_new_n1322_; 
wire _abc_4635_new_n1323_; 
wire _abc_4635_new_n1324_; 
wire _abc_4635_new_n1325_; 
wire _abc_4635_new_n1327_; 
wire _abc_4635_new_n1328_; 
wire _abc_4635_new_n1329_; 
wire _abc_4635_new_n1330_; 
wire _abc_4635_new_n1331_; 
wire _abc_4635_new_n1332_; 
wire _abc_4635_new_n1333_; 
wire _abc_4635_new_n1334_; 
wire _abc_4635_new_n1335_; 
wire _abc_4635_new_n1336_; 
wire _abc_4635_new_n1337_; 
wire _abc_4635_new_n1338_; 
wire _abc_4635_new_n1339_; 
wire _abc_4635_new_n1340_; 
wire _abc_4635_new_n1341_; 
wire _abc_4635_new_n1342_; 
wire _abc_4635_new_n1343_; 
wire _abc_4635_new_n1344_; 
wire _abc_4635_new_n1345_; 
wire _abc_4635_new_n1346_; 
wire _abc_4635_new_n1347_; 
wire _abc_4635_new_n1349_; 
wire _abc_4635_new_n1350_; 
wire _abc_4635_new_n1351_; 
wire _abc_4635_new_n1352_; 
wire _abc_4635_new_n1353_; 
wire _abc_4635_new_n1354_; 
wire _abc_4635_new_n1355_; 
wire _abc_4635_new_n1356_; 
wire _abc_4635_new_n1357_; 
wire _abc_4635_new_n1358_; 
wire _abc_4635_new_n1359_; 
wire _abc_4635_new_n1360_; 
wire _abc_4635_new_n1362_; 
wire _abc_4635_new_n1363_; 
wire _abc_4635_new_n1364_; 
wire _abc_4635_new_n1365_; 
wire _abc_4635_new_n1366_; 
wire _abc_4635_new_n1367_; 
wire _abc_4635_new_n1368_; 
wire _abc_4635_new_n1369_; 
wire _abc_4635_new_n1370_; 
wire _abc_4635_new_n1371_; 
wire _abc_4635_new_n1372_; 
wire _abc_4635_new_n1373_; 
wire _abc_4635_new_n1374_; 
wire _abc_4635_new_n1375_; 
wire _abc_4635_new_n1376_; 
wire _abc_4635_new_n1377_; 
wire _abc_4635_new_n1379_; 
wire _abc_4635_new_n1380_; 
wire _abc_4635_new_n1381_; 
wire _abc_4635_new_n1382_; 
wire _abc_4635_new_n1383_; 
wire _abc_4635_new_n1384_; 
wire _abc_4635_new_n1385_; 
wire _abc_4635_new_n1386_; 
wire _abc_4635_new_n1387_; 
wire _abc_4635_new_n1388_; 
wire _abc_4635_new_n1389_; 
wire _abc_4635_new_n1390_; 
wire _abc_4635_new_n1392_; 
wire _abc_4635_new_n1393_; 
wire _abc_4635_new_n1394_; 
wire _abc_4635_new_n1395_; 
wire _abc_4635_new_n1396_; 
wire _abc_4635_new_n1397_; 
wire _abc_4635_new_n1398_; 
wire _abc_4635_new_n1399_; 
wire _abc_4635_new_n1400_; 
wire _abc_4635_new_n1401_; 
wire _abc_4635_new_n1402_; 
wire _abc_4635_new_n1403_; 
wire _abc_4635_new_n1404_; 
wire _abc_4635_new_n1405_; 
wire _abc_4635_new_n1406_; 
wire _abc_4635_new_n1407_; 
wire _abc_4635_new_n1408_; 
wire _abc_4635_new_n1409_; 
wire _abc_4635_new_n1411_; 
wire _abc_4635_new_n1412_; 
wire _abc_4635_new_n1413_; 
wire _abc_4635_new_n1414_; 
wire _abc_4635_new_n1415_; 
wire _abc_4635_new_n1416_; 
wire _abc_4635_new_n1417_; 
wire _abc_4635_new_n1418_; 
wire _abc_4635_new_n1419_; 
wire _abc_4635_new_n1420_; 
wire _abc_4635_new_n1421_; 
wire _abc_4635_new_n1422_; 
wire _abc_4635_new_n1424_; 
wire _abc_4635_new_n1425_; 
wire _abc_4635_new_n1426_; 
wire _abc_4635_new_n1427_; 
wire _abc_4635_new_n1428_; 
wire _abc_4635_new_n1429_; 
wire _abc_4635_new_n1430_; 
wire _abc_4635_new_n1431_; 
wire _abc_4635_new_n1432_; 
wire _abc_4635_new_n1433_; 
wire _abc_4635_new_n1434_; 
wire _abc_4635_new_n1435_; 
wire _abc_4635_new_n1436_; 
wire _abc_4635_new_n1437_; 
wire _abc_4635_new_n1438_; 
wire _abc_4635_new_n1439_; 
wire _abc_4635_new_n1440_; 
wire _abc_4635_new_n1441_; 
wire _abc_4635_new_n1442_; 
wire _abc_4635_new_n1443_; 
wire _abc_4635_new_n1444_; 
wire _abc_4635_new_n1445_; 
wire _abc_4635_new_n1446_; 
wire _abc_4635_new_n1447_; 
wire _abc_4635_new_n1448_; 
wire _abc_4635_new_n1449_; 
wire _abc_4635_new_n1450_; 
wire _abc_4635_new_n1451_; 
wire _abc_4635_new_n1452_; 
wire _abc_4635_new_n1453_; 
wire _abc_4635_new_n1454_; 
wire _abc_4635_new_n1455_; 
wire _abc_4635_new_n1456_; 
wire _abc_4635_new_n1457_; 
wire _abc_4635_new_n1458_; 
wire _abc_4635_new_n1459_; 
wire _abc_4635_new_n1460_; 
wire _abc_4635_new_n1461_; 
wire _abc_4635_new_n1462_; 
wire _abc_4635_new_n1463_; 
wire _abc_4635_new_n1464_; 
wire _abc_4635_new_n1466_; 
wire _abc_4635_new_n1467_; 
wire _abc_4635_new_n1468_; 
wire _abc_4635_new_n1469_; 
wire _abc_4635_new_n1470_; 
wire _abc_4635_new_n1471_; 
wire _abc_4635_new_n1472_; 
wire _abc_4635_new_n1473_; 
wire _abc_4635_new_n1474_; 
wire _abc_4635_new_n1475_; 
wire _abc_4635_new_n1476_; 
wire _abc_4635_new_n1477_; 
wire _abc_4635_new_n1478_; 
wire _abc_4635_new_n1479_; 
wire _abc_4635_new_n1482_; 
wire _abc_4635_new_n1483_; 
wire _abc_4635_new_n1484_; 
wire _abc_4635_new_n1486_; 
wire _abc_4635_new_n361_; 
wire _abc_4635_new_n362_; 
wire _abc_4635_new_n363_; 
wire _abc_4635_new_n364_; 
wire _abc_4635_new_n365_; 
wire _abc_4635_new_n366_; 
wire _abc_4635_new_n367_; 
wire _abc_4635_new_n368_; 
wire _abc_4635_new_n369_; 
wire _abc_4635_new_n370_; 
wire _abc_4635_new_n371_; 
wire _abc_4635_new_n372_; 
wire _abc_4635_new_n373_; 
wire _abc_4635_new_n374_; 
wire _abc_4635_new_n375_; 
wire _abc_4635_new_n376_; 
wire _abc_4635_new_n377_; 
wire _abc_4635_new_n378_; 
wire _abc_4635_new_n379_; 
wire _abc_4635_new_n380_; 
wire _abc_4635_new_n381_; 
wire _abc_4635_new_n382_; 
wire _abc_4635_new_n383_; 
wire _abc_4635_new_n384_; 
wire _abc_4635_new_n385_; 
wire _abc_4635_new_n386_; 
wire _abc_4635_new_n387_; 
wire _abc_4635_new_n389_; 
wire _abc_4635_new_n390_; 
wire _abc_4635_new_n391_; 
wire _abc_4635_new_n392_; 
wire _abc_4635_new_n393_; 
wire _abc_4635_new_n394_; 
wire _abc_4635_new_n395_; 
wire _abc_4635_new_n397_; 
wire _abc_4635_new_n398_; 
wire _abc_4635_new_n399_; 
wire _abc_4635_new_n401_; 
wire _abc_4635_new_n402_; 
wire _abc_4635_new_n403_; 
wire _abc_4635_new_n404_; 
wire _abc_4635_new_n405_; 
wire _abc_4635_new_n406_; 
wire _abc_4635_new_n407_; 
wire _abc_4635_new_n408_; 
wire _abc_4635_new_n409_; 
wire _abc_4635_new_n410_; 
wire _abc_4635_new_n411_; 
wire _abc_4635_new_n412_; 
wire _abc_4635_new_n413_; 
wire _abc_4635_new_n414_; 
wire _abc_4635_new_n415_; 
wire _abc_4635_new_n416_; 
wire _abc_4635_new_n417_; 
wire _abc_4635_new_n419_; 
wire _abc_4635_new_n420_; 
wire _abc_4635_new_n421_; 
wire _abc_4635_new_n422_; 
wire _abc_4635_new_n423_; 
wire _abc_4635_new_n425_; 
wire _abc_4635_new_n426_; 
wire _abc_4635_new_n428_; 
wire _abc_4635_new_n429_; 
wire _abc_4635_new_n430_; 
wire _abc_4635_new_n431_; 
wire _abc_4635_new_n433_; 
wire _abc_4635_new_n434_; 
wire _abc_4635_new_n435_; 
wire _abc_4635_new_n436_; 
wire _abc_4635_new_n437_; 
wire _abc_4635_new_n438_; 
wire _abc_4635_new_n439_; 
wire _abc_4635_new_n440_; 
wire _abc_4635_new_n441_; 
wire _abc_4635_new_n442_; 
wire _abc_4635_new_n443_; 
wire _abc_4635_new_n444_; 
wire _abc_4635_new_n445_; 
wire _abc_4635_new_n446_; 
wire _abc_4635_new_n447_; 
wire _abc_4635_new_n448_; 
wire _abc_4635_new_n449_; 
wire _abc_4635_new_n450_; 
wire _abc_4635_new_n451_; 
wire _abc_4635_new_n452_; 
wire _abc_4635_new_n453_; 
wire _abc_4635_new_n454_; 
wire _abc_4635_new_n457_; 
wire _abc_4635_new_n458_; 
wire _abc_4635_new_n459_; 
wire _abc_4635_new_n460_; 
wire _abc_4635_new_n461_; 
wire _abc_4635_new_n462_; 
wire _abc_4635_new_n463_; 
wire _abc_4635_new_n464_; 
wire _abc_4635_new_n465_; 
wire _abc_4635_new_n466_; 
wire _abc_4635_new_n467_; 
wire _abc_4635_new_n468_; 
wire _abc_4635_new_n469_; 
wire _abc_4635_new_n470_; 
wire _abc_4635_new_n471_; 
wire _abc_4635_new_n472_; 
wire _abc_4635_new_n472__bF_buf0; 
wire _abc_4635_new_n472__bF_buf1; 
wire _abc_4635_new_n472__bF_buf2; 
wire _abc_4635_new_n472__bF_buf3; 
wire _abc_4635_new_n473_; 
wire _abc_4635_new_n474_; 
wire _abc_4635_new_n475_; 
wire _abc_4635_new_n476_; 
wire _abc_4635_new_n477_; 
wire _abc_4635_new_n478_; 
wire _abc_4635_new_n479_; 
wire _abc_4635_new_n480_; 
wire _abc_4635_new_n480__bF_buf0; 
wire _abc_4635_new_n480__bF_buf1; 
wire _abc_4635_new_n480__bF_buf2; 
wire _abc_4635_new_n480__bF_buf3; 
wire _abc_4635_new_n480__bF_buf4; 
wire _abc_4635_new_n481_; 
wire _abc_4635_new_n482_; 
wire _abc_4635_new_n483_; 
wire _abc_4635_new_n484_; 
wire _abc_4635_new_n485_; 
wire _abc_4635_new_n485__bF_buf0; 
wire _abc_4635_new_n485__bF_buf1; 
wire _abc_4635_new_n485__bF_buf2; 
wire _abc_4635_new_n485__bF_buf3; 
wire _abc_4635_new_n485__bF_buf4; 
wire _abc_4635_new_n486_; 
wire _abc_4635_new_n487_; 
wire _abc_4635_new_n489_; 
wire _abc_4635_new_n490_; 
wire _abc_4635_new_n491_; 
wire _abc_4635_new_n493_; 
wire _abc_4635_new_n493__bF_buf0; 
wire _abc_4635_new_n493__bF_buf1; 
wire _abc_4635_new_n493__bF_buf2; 
wire _abc_4635_new_n493__bF_buf3; 
wire _abc_4635_new_n494_; 
wire _abc_4635_new_n495_; 
wire _abc_4635_new_n496_; 
wire _abc_4635_new_n498_; 
wire _abc_4635_new_n499_; 
wire _abc_4635_new_n509_; 
wire _abc_4635_new_n510_; 
wire _abc_4635_new_n511_; 
wire _abc_4635_new_n511__bF_buf0; 
wire _abc_4635_new_n511__bF_buf1; 
wire _abc_4635_new_n511__bF_buf2; 
wire _abc_4635_new_n511__bF_buf3; 
wire _abc_4635_new_n511__bF_buf4; 
wire _abc_4635_new_n511__bF_buf5; 
wire _abc_4635_new_n511__bF_buf6; 
wire _abc_4635_new_n512_; 
wire _abc_4635_new_n513_; 
wire _abc_4635_new_n514_; 
wire _abc_4635_new_n516_; 
wire _abc_4635_new_n517_; 
wire _abc_4635_new_n518_; 
wire _abc_4635_new_n519_; 
wire _abc_4635_new_n521_; 
wire _abc_4635_new_n522_; 
wire _abc_4635_new_n523_; 
wire _abc_4635_new_n524_; 
wire _abc_4635_new_n526_; 
wire _abc_4635_new_n527_; 
wire _abc_4635_new_n528_; 
wire _abc_4635_new_n529_; 
wire _abc_4635_new_n531_; 
wire _abc_4635_new_n532_; 
wire _abc_4635_new_n533_; 
wire _abc_4635_new_n534_; 
wire _abc_4635_new_n536_; 
wire _abc_4635_new_n537_; 
wire _abc_4635_new_n538_; 
wire _abc_4635_new_n539_; 
wire _abc_4635_new_n541_; 
wire _abc_4635_new_n542_; 
wire _abc_4635_new_n543_; 
wire _abc_4635_new_n544_; 
wire _abc_4635_new_n546_; 
wire _abc_4635_new_n547_; 
wire _abc_4635_new_n548_; 
wire _abc_4635_new_n549_; 
wire _abc_4635_new_n551_; 
wire _abc_4635_new_n552_; 
wire _abc_4635_new_n554_; 
wire _abc_4635_new_n555_; 
wire _abc_4635_new_n557_; 
wire _abc_4635_new_n558_; 
wire _abc_4635_new_n560_; 
wire _abc_4635_new_n561_; 
wire _abc_4635_new_n563_; 
wire _abc_4635_new_n564_; 
wire _abc_4635_new_n566_; 
wire _abc_4635_new_n567_; 
wire _abc_4635_new_n569_; 
wire _abc_4635_new_n570_; 
wire _abc_4635_new_n572_; 
wire _abc_4635_new_n573_; 
wire _abc_4635_new_n575_; 
wire _abc_4635_new_n576_; 
wire _abc_4635_new_n577_; 
wire _abc_4635_new_n578_; 
wire _abc_4635_new_n580_; 
wire _abc_4635_new_n581_; 
wire _abc_4635_new_n582_; 
wire _abc_4635_new_n583_; 
wire _abc_4635_new_n585_; 
wire _abc_4635_new_n586_; 
wire _abc_4635_new_n587_; 
wire _abc_4635_new_n588_; 
wire _abc_4635_new_n590_; 
wire _abc_4635_new_n591_; 
wire _abc_4635_new_n592_; 
wire _abc_4635_new_n593_; 
wire _abc_4635_new_n595_; 
wire _abc_4635_new_n596_; 
wire _abc_4635_new_n597_; 
wire _abc_4635_new_n598_; 
wire _abc_4635_new_n600_; 
wire _abc_4635_new_n601_; 
wire _abc_4635_new_n602_; 
wire _abc_4635_new_n603_; 
wire _abc_4635_new_n605_; 
wire _abc_4635_new_n606_; 
wire _abc_4635_new_n607_; 
wire _abc_4635_new_n608_; 
wire _abc_4635_new_n610_; 
wire _abc_4635_new_n611_; 
wire _abc_4635_new_n612_; 
wire _abc_4635_new_n613_; 
wire _abc_4635_new_n615_; 
wire _abc_4635_new_n616_; 
wire _abc_4635_new_n616__bF_buf0; 
wire _abc_4635_new_n616__bF_buf1; 
wire _abc_4635_new_n616__bF_buf2; 
wire _abc_4635_new_n616__bF_buf3; 
wire _abc_4635_new_n616__bF_buf4; 
wire _abc_4635_new_n617_; 
wire _abc_4635_new_n618_; 
wire _abc_4635_new_n618__bF_buf0; 
wire _abc_4635_new_n618__bF_buf1; 
wire _abc_4635_new_n618__bF_buf2; 
wire _abc_4635_new_n618__bF_buf3; 
wire _abc_4635_new_n618__bF_buf4; 
wire _abc_4635_new_n619_; 
wire _abc_4635_new_n620_; 
wire _abc_4635_new_n622_; 
wire _abc_4635_new_n623_; 
wire _abc_4635_new_n624_; 
wire _abc_4635_new_n626_; 
wire _abc_4635_new_n627_; 
wire _abc_4635_new_n628_; 
wire _abc_4635_new_n630_; 
wire _abc_4635_new_n631_; 
wire _abc_4635_new_n632_; 
wire _abc_4635_new_n634_; 
wire _abc_4635_new_n635_; 
wire _abc_4635_new_n636_; 
wire _abc_4635_new_n638_; 
wire _abc_4635_new_n639_; 
wire _abc_4635_new_n640_; 
wire _abc_4635_new_n642_; 
wire _abc_4635_new_n643_; 
wire _abc_4635_new_n644_; 
wire _abc_4635_new_n646_; 
wire _abc_4635_new_n647_; 
wire _abc_4635_new_n648_; 
wire _abc_4635_new_n650_; 
wire _abc_4635_new_n651_; 
wire _abc_4635_new_n652_; 
wire _abc_4635_new_n654_; 
wire _abc_4635_new_n655_; 
wire _abc_4635_new_n656_; 
wire _abc_4635_new_n658_; 
wire _abc_4635_new_n659_; 
wire _abc_4635_new_n660_; 
wire _abc_4635_new_n662_; 
wire _abc_4635_new_n663_; 
wire _abc_4635_new_n664_; 
wire _abc_4635_new_n666_; 
wire _abc_4635_new_n667_; 
wire _abc_4635_new_n668_; 
wire _abc_4635_new_n670_; 
wire _abc_4635_new_n671_; 
wire _abc_4635_new_n672_; 
wire _abc_4635_new_n674_; 
wire _abc_4635_new_n675_; 
wire _abc_4635_new_n676_; 
wire _abc_4635_new_n678_; 
wire _abc_4635_new_n679_; 
wire _abc_4635_new_n680_; 
wire _abc_4635_new_n682_; 
wire _abc_4635_new_n683_; 
wire _abc_4635_new_n684_; 
wire _abc_4635_new_n686_; 
wire _abc_4635_new_n687_; 
wire _abc_4635_new_n688_; 
wire _abc_4635_new_n690_; 
wire _abc_4635_new_n691_; 
wire _abc_4635_new_n692_; 
wire _abc_4635_new_n694_; 
wire _abc_4635_new_n695_; 
wire _abc_4635_new_n696_; 
wire _abc_4635_new_n698_; 
wire _abc_4635_new_n699_; 
wire _abc_4635_new_n700_; 
wire _abc_4635_new_n702_; 
wire _abc_4635_new_n703_; 
wire _abc_4635_new_n704_; 
wire _abc_4635_new_n706_; 
wire _abc_4635_new_n707_; 
wire _abc_4635_new_n708_; 
wire _abc_4635_new_n710_; 
wire _abc_4635_new_n711_; 
wire _abc_4635_new_n712_; 
wire _abc_4635_new_n714_; 
wire _abc_4635_new_n715_; 
wire _abc_4635_new_n716_; 
wire _abc_4635_new_n718_; 
wire _abc_4635_new_n719_; 
wire _abc_4635_new_n720_; 
wire _abc_4635_new_n722_; 
wire _abc_4635_new_n723_; 
wire _abc_4635_new_n724_; 
wire _abc_4635_new_n726_; 
wire _abc_4635_new_n727_; 
wire _abc_4635_new_n728_; 
wire _abc_4635_new_n730_; 
wire _abc_4635_new_n731_; 
wire _abc_4635_new_n732_; 
wire _abc_4635_new_n734_; 
wire _abc_4635_new_n735_; 
wire _abc_4635_new_n736_; 
wire _abc_4635_new_n738_; 
wire _abc_4635_new_n739_; 
wire _abc_4635_new_n740_; 
wire _abc_4635_new_n742_; 
wire _abc_4635_new_n743_; 
wire _abc_4635_new_n744_; 
wire _abc_4635_new_n746_; 
wire _abc_4635_new_n747_; 
wire _abc_4635_new_n748_; 
wire _abc_4635_new_n749_; 
wire _abc_4635_new_n750_; 
wire _abc_4635_new_n751_; 
wire _abc_4635_new_n753_; 
wire _abc_4635_new_n753__bF_buf0; 
wire _abc_4635_new_n753__bF_buf1; 
wire _abc_4635_new_n753__bF_buf2; 
wire _abc_4635_new_n753__bF_buf3; 
wire _abc_4635_new_n753__bF_buf4; 
wire _abc_4635_new_n754_; 
wire _abc_4635_new_n754__bF_buf0; 
wire _abc_4635_new_n754__bF_buf1; 
wire _abc_4635_new_n754__bF_buf2; 
wire _abc_4635_new_n754__bF_buf3; 
wire _abc_4635_new_n754__bF_buf4; 
wire _abc_4635_new_n755_; 
wire _abc_4635_new_n756_; 
wire _abc_4635_new_n757_; 
wire _abc_4635_new_n758_; 
wire _abc_4635_new_n759_; 
wire _abc_4635_new_n760_; 
wire _abc_4635_new_n761_; 
wire _abc_4635_new_n762_; 
wire _abc_4635_new_n763_; 
wire _abc_4635_new_n764_; 
wire _abc_4635_new_n765_; 
wire _abc_4635_new_n766_; 
wire _abc_4635_new_n767_; 
wire _abc_4635_new_n768_; 
wire _abc_4635_new_n769_; 
wire _abc_4635_new_n770_; 
wire _abc_4635_new_n772_; 
wire _abc_4635_new_n773_; 
wire _abc_4635_new_n774_; 
wire _abc_4635_new_n775_; 
wire _abc_4635_new_n776_; 
wire _abc_4635_new_n777_; 
wire _abc_4635_new_n778_; 
wire _abc_4635_new_n779_; 
wire _abc_4635_new_n780_; 
wire _abc_4635_new_n781_; 
wire _abc_4635_new_n782_; 
wire _abc_4635_new_n783_; 
wire _abc_4635_new_n784_; 
wire _abc_4635_new_n785_; 
wire _abc_4635_new_n786_; 
wire _abc_4635_new_n787_; 
wire _abc_4635_new_n789_; 
wire _abc_4635_new_n790_; 
wire _abc_4635_new_n791_; 
wire _abc_4635_new_n792_; 
wire _abc_4635_new_n793_; 
wire _abc_4635_new_n794_; 
wire _abc_4635_new_n795_; 
wire _abc_4635_new_n796_; 
wire _abc_4635_new_n797_; 
wire _abc_4635_new_n798_; 
wire _abc_4635_new_n799_; 
wire _abc_4635_new_n800_; 
wire _abc_4635_new_n801_; 
wire _abc_4635_new_n802_; 
wire _abc_4635_new_n803_; 
wire _abc_4635_new_n804_; 
wire _abc_4635_new_n806_; 
wire _abc_4635_new_n807_; 
wire _abc_4635_new_n808_; 
wire _abc_4635_new_n809_; 
wire _abc_4635_new_n810_; 
wire _abc_4635_new_n811_; 
wire _abc_4635_new_n812_; 
wire _abc_4635_new_n813_; 
wire _abc_4635_new_n814_; 
wire _abc_4635_new_n815_; 
wire _abc_4635_new_n816_; 
wire _abc_4635_new_n817_; 
wire _abc_4635_new_n818_; 
wire _abc_4635_new_n819_; 
wire _abc_4635_new_n820_; 
wire _abc_4635_new_n821_; 
wire _abc_4635_new_n823_; 
wire _abc_4635_new_n824_; 
wire _abc_4635_new_n825_; 
wire _abc_4635_new_n826_; 
wire _abc_4635_new_n827_; 
wire _abc_4635_new_n828_; 
wire _abc_4635_new_n829_; 
wire _abc_4635_new_n830_; 
wire _abc_4635_new_n831_; 
wire _abc_4635_new_n832_; 
wire _abc_4635_new_n833_; 
wire _abc_4635_new_n834_; 
wire _abc_4635_new_n835_; 
wire _abc_4635_new_n836_; 
wire _abc_4635_new_n837_; 
wire _abc_4635_new_n838_; 
wire _abc_4635_new_n840_; 
wire _abc_4635_new_n841_; 
wire _abc_4635_new_n842_; 
wire _abc_4635_new_n843_; 
wire _abc_4635_new_n844_; 
wire _abc_4635_new_n845_; 
wire _abc_4635_new_n846_; 
wire _abc_4635_new_n847_; 
wire _abc_4635_new_n848_; 
wire _abc_4635_new_n849_; 
wire _abc_4635_new_n850_; 
wire _abc_4635_new_n851_; 
wire _abc_4635_new_n852_; 
wire _abc_4635_new_n853_; 
wire _abc_4635_new_n854_; 
wire _abc_4635_new_n855_; 
wire _abc_4635_new_n857_; 
wire _abc_4635_new_n858_; 
wire _abc_4635_new_n859_; 
wire _abc_4635_new_n860_; 
wire _abc_4635_new_n861_; 
wire _abc_4635_new_n862_; 
wire _abc_4635_new_n863_; 
wire _abc_4635_new_n864_; 
wire _abc_4635_new_n865_; 
wire _abc_4635_new_n866_; 
wire _abc_4635_new_n867_; 
wire _abc_4635_new_n868_; 
wire _abc_4635_new_n869_; 
wire _abc_4635_new_n870_; 
wire _abc_4635_new_n871_; 
wire _abc_4635_new_n872_; 
wire _abc_4635_new_n874_; 
wire _abc_4635_new_n875_; 
wire _abc_4635_new_n876_; 
wire _abc_4635_new_n877_; 
wire _abc_4635_new_n878_; 
wire _abc_4635_new_n879_; 
wire _abc_4635_new_n880_; 
wire _abc_4635_new_n881_; 
wire _abc_4635_new_n882_; 
wire _abc_4635_new_n883_; 
wire _abc_4635_new_n884_; 
wire _abc_4635_new_n885_; 
wire _abc_4635_new_n886_; 
wire _abc_4635_new_n887_; 
wire _abc_4635_new_n888_; 
wire _abc_4635_new_n889_; 
wire _abc_4635_new_n890_; 
wire _abc_4635_new_n891_; 
wire _abc_4635_new_n893_; 
wire _abc_4635_new_n894_; 
wire _abc_4635_new_n895_; 
wire _abc_4635_new_n896_; 
wire _abc_4635_new_n897_; 
wire _abc_4635_new_n898_; 
wire _abc_4635_new_n900_; 
wire _abc_4635_new_n901_; 
wire _abc_4635_new_n902_; 
wire _abc_4635_new_n903_; 
wire _abc_4635_new_n905_; 
wire _abc_4635_new_n906_; 
wire _abc_4635_new_n907_; 
wire _abc_4635_new_n908_; 
wire _abc_4635_new_n910_; 
wire _abc_4635_new_n911_; 
wire _abc_4635_new_n912_; 
wire _abc_4635_new_n913_; 
wire _abc_4635_new_n915_; 
wire _abc_4635_new_n916_; 
wire _abc_4635_new_n917_; 
wire _abc_4635_new_n918_; 
wire _abc_4635_new_n920_; 
wire _abc_4635_new_n921_; 
wire _abc_4635_new_n922_; 
wire _abc_4635_new_n923_; 
wire _abc_4635_new_n925_; 
wire _abc_4635_new_n926_; 
wire _abc_4635_new_n927_; 
wire _abc_4635_new_n928_; 
wire _abc_4635_new_n930_; 
wire _abc_4635_new_n931_; 
wire _abc_4635_new_n932_; 
wire _abc_4635_new_n933_; 
wire _abc_4635_new_n934_; 
wire _abc_4635_new_n935_; 
wire _abc_4635_new_n936_; 
wire _abc_4635_new_n938_; 
wire _abc_4635_new_n939_; 
wire _abc_4635_new_n940_; 
wire _abc_4635_new_n941_; 
wire _abc_4635_new_n943_; 
wire _abc_4635_new_n944_; 
wire _abc_4635_new_n946_; 
wire _abc_4635_new_n947_; 
wire _abc_4635_new_n949_; 
wire _abc_4635_new_n950_; 
wire _abc_4635_new_n952_; 
wire _abc_4635_new_n953_; 
wire _abc_4635_new_n955_; 
wire _abc_4635_new_n956_; 
wire _abc_4635_new_n958_; 
wire _abc_4635_new_n959_; 
wire _abc_4635_new_n961_; 
wire _abc_4635_new_n962_; 
wire _abc_4635_new_n964_; 
wire _abc_4635_new_n965_; 
wire _abc_4635_new_n967_; 
wire _abc_4635_new_n968_; 
wire _abc_4635_new_n970_; 
wire _abc_4635_new_n971_; 
wire _abc_4635_new_n973_; 
wire _abc_4635_new_n974_; 
wire _abc_4635_new_n976_; 
wire _abc_4635_new_n977_; 
wire _abc_4635_new_n979_; 
wire _abc_4635_new_n980_; 
wire _abc_4635_new_n982_; 
wire _abc_4635_new_n983_; 
wire _abc_4635_new_n985_; 
wire _abc_4635_new_n986_; 
wire _abc_4635_new_n988_; 
wire _abc_4635_new_n989_; 
wire _abc_4635_new_n991_; 
wire _abc_4635_new_n992_; 
wire _abc_4635_new_n994_; 
wire _abc_4635_new_n995_; 
wire _abc_4635_new_n996_; 
wire _abc_4635_new_n997_; 
wire _abc_4635_new_n998_; 
wire _abc_4635_new_n999_; 
wire _auto_iopadmap_cc_368_execute_5767_0_; 
wire _auto_iopadmap_cc_368_execute_5767_10_; 
wire _auto_iopadmap_cc_368_execute_5767_11_; 
wire _auto_iopadmap_cc_368_execute_5767_12_; 
wire _auto_iopadmap_cc_368_execute_5767_13_; 
wire _auto_iopadmap_cc_368_execute_5767_14_; 
wire _auto_iopadmap_cc_368_execute_5767_15_; 
wire _auto_iopadmap_cc_368_execute_5767_16_; 
wire _auto_iopadmap_cc_368_execute_5767_17_; 
wire _auto_iopadmap_cc_368_execute_5767_18_; 
wire _auto_iopadmap_cc_368_execute_5767_19_; 
wire _auto_iopadmap_cc_368_execute_5767_1_; 
wire _auto_iopadmap_cc_368_execute_5767_20_; 
wire _auto_iopadmap_cc_368_execute_5767_21_; 
wire _auto_iopadmap_cc_368_execute_5767_22_; 
wire _auto_iopadmap_cc_368_execute_5767_23_; 
wire _auto_iopadmap_cc_368_execute_5767_24_; 
wire _auto_iopadmap_cc_368_execute_5767_25_; 
wire _auto_iopadmap_cc_368_execute_5767_26_; 
wire _auto_iopadmap_cc_368_execute_5767_27_; 
wire _auto_iopadmap_cc_368_execute_5767_28_; 
wire _auto_iopadmap_cc_368_execute_5767_29_; 
wire _auto_iopadmap_cc_368_execute_5767_2_; 
wire _auto_iopadmap_cc_368_execute_5767_30_; 
wire _auto_iopadmap_cc_368_execute_5767_31_; 
wire _auto_iopadmap_cc_368_execute_5767_3_; 
wire _auto_iopadmap_cc_368_execute_5767_4_; 
wire _auto_iopadmap_cc_368_execute_5767_5_; 
wire _auto_iopadmap_cc_368_execute_5767_6_; 
wire _auto_iopadmap_cc_368_execute_5767_7_; 
wire _auto_iopadmap_cc_368_execute_5767_8_; 
wire _auto_iopadmap_cc_368_execute_5767_9_; 
wire _auto_iopadmap_cc_368_execute_5800; 
wire _auto_iopadmap_cc_368_execute_5835; 
wire _auto_iopadmap_cc_368_execute_5837; 
wire _auto_iopadmap_cc_368_execute_5839; 
wire _auto_iopadmap_cc_368_execute_5841_0_; 
wire _auto_iopadmap_cc_368_execute_5841_10_; 
wire _auto_iopadmap_cc_368_execute_5841_11_; 
wire _auto_iopadmap_cc_368_execute_5841_12_; 
wire _auto_iopadmap_cc_368_execute_5841_13_; 
wire _auto_iopadmap_cc_368_execute_5841_14_; 
wire _auto_iopadmap_cc_368_execute_5841_15_; 
wire _auto_iopadmap_cc_368_execute_5841_16_; 
wire _auto_iopadmap_cc_368_execute_5841_17_; 
wire _auto_iopadmap_cc_368_execute_5841_18_; 
wire _auto_iopadmap_cc_368_execute_5841_19_; 
wire _auto_iopadmap_cc_368_execute_5841_1_; 
wire _auto_iopadmap_cc_368_execute_5841_20_; 
wire _auto_iopadmap_cc_368_execute_5841_21_; 
wire _auto_iopadmap_cc_368_execute_5841_22_; 
wire _auto_iopadmap_cc_368_execute_5841_23_; 
wire _auto_iopadmap_cc_368_execute_5841_24_; 
wire _auto_iopadmap_cc_368_execute_5841_25_; 
wire _auto_iopadmap_cc_368_execute_5841_26_; 
wire _auto_iopadmap_cc_368_execute_5841_27_; 
wire _auto_iopadmap_cc_368_execute_5841_28_; 
wire _auto_iopadmap_cc_368_execute_5841_29_; 
wire _auto_iopadmap_cc_368_execute_5841_2_; 
wire _auto_iopadmap_cc_368_execute_5841_30_; 
wire _auto_iopadmap_cc_368_execute_5841_31_; 
wire _auto_iopadmap_cc_368_execute_5841_3_; 
wire _auto_iopadmap_cc_368_execute_5841_4_; 
wire _auto_iopadmap_cc_368_execute_5841_5_; 
wire _auto_iopadmap_cc_368_execute_5841_6_; 
wire _auto_iopadmap_cc_368_execute_5841_7_; 
wire _auto_iopadmap_cc_368_execute_5841_8_; 
wire _auto_iopadmap_cc_368_execute_5841_9_; 
wire _auto_iopadmap_cc_368_execute_5874_0_; 
wire _auto_iopadmap_cc_368_execute_5874_1_; 
wire _auto_iopadmap_cc_368_execute_5874_2_; 
wire _auto_iopadmap_cc_368_execute_5874_3_; 
wire _auto_iopadmap_cc_368_execute_5879; 
wire _auto_iopadmap_cc_368_execute_5881; 
wire _auto_iopadmap_cc_368_execute_5890; 
wire _auto_iopadmap_cc_368_execute_5892; 
wire _auto_iopadmap_cc_368_execute_5894_0_; 
wire _auto_iopadmap_cc_368_execute_5894_10_; 
wire _auto_iopadmap_cc_368_execute_5894_11_; 
wire _auto_iopadmap_cc_368_execute_5894_12_; 
wire _auto_iopadmap_cc_368_execute_5894_13_; 
wire _auto_iopadmap_cc_368_execute_5894_14_; 
wire _auto_iopadmap_cc_368_execute_5894_15_; 
wire _auto_iopadmap_cc_368_execute_5894_16_; 
wire _auto_iopadmap_cc_368_execute_5894_17_; 
wire _auto_iopadmap_cc_368_execute_5894_18_; 
wire _auto_iopadmap_cc_368_execute_5894_19_; 
wire _auto_iopadmap_cc_368_execute_5894_1_; 
wire _auto_iopadmap_cc_368_execute_5894_20_; 
wire _auto_iopadmap_cc_368_execute_5894_21_; 
wire _auto_iopadmap_cc_368_execute_5894_22_; 
wire _auto_iopadmap_cc_368_execute_5894_23_; 
wire _auto_iopadmap_cc_368_execute_5894_24_; 
wire _auto_iopadmap_cc_368_execute_5894_25_; 
wire _auto_iopadmap_cc_368_execute_5894_26_; 
wire _auto_iopadmap_cc_368_execute_5894_27_; 
wire _auto_iopadmap_cc_368_execute_5894_28_; 
wire _auto_iopadmap_cc_368_execute_5894_29_; 
wire _auto_iopadmap_cc_368_execute_5894_2_; 
wire _auto_iopadmap_cc_368_execute_5894_30_; 
wire _auto_iopadmap_cc_368_execute_5894_31_; 
wire _auto_iopadmap_cc_368_execute_5894_3_; 
wire _auto_iopadmap_cc_368_execute_5894_4_; 
wire _auto_iopadmap_cc_368_execute_5894_5_; 
wire _auto_iopadmap_cc_368_execute_5894_6_; 
wire _auto_iopadmap_cc_368_execute_5894_7_; 
wire _auto_iopadmap_cc_368_execute_5894_8_; 
wire _auto_iopadmap_cc_368_execute_5894_9_; 
wire _auto_iopadmap_cc_368_execute_5927_0_; 
wire _auto_iopadmap_cc_368_execute_5927_10_; 
wire _auto_iopadmap_cc_368_execute_5927_11_; 
wire _auto_iopadmap_cc_368_execute_5927_12_; 
wire _auto_iopadmap_cc_368_execute_5927_13_; 
wire _auto_iopadmap_cc_368_execute_5927_14_; 
wire _auto_iopadmap_cc_368_execute_5927_15_; 
wire _auto_iopadmap_cc_368_execute_5927_16_; 
wire _auto_iopadmap_cc_368_execute_5927_17_; 
wire _auto_iopadmap_cc_368_execute_5927_18_; 
wire _auto_iopadmap_cc_368_execute_5927_19_; 
wire _auto_iopadmap_cc_368_execute_5927_1_; 
wire _auto_iopadmap_cc_368_execute_5927_20_; 
wire _auto_iopadmap_cc_368_execute_5927_21_; 
wire _auto_iopadmap_cc_368_execute_5927_22_; 
wire _auto_iopadmap_cc_368_execute_5927_23_; 
wire _auto_iopadmap_cc_368_execute_5927_24_; 
wire _auto_iopadmap_cc_368_execute_5927_25_; 
wire _auto_iopadmap_cc_368_execute_5927_26_; 
wire _auto_iopadmap_cc_368_execute_5927_27_; 
wire _auto_iopadmap_cc_368_execute_5927_28_; 
wire _auto_iopadmap_cc_368_execute_5927_29_; 
wire _auto_iopadmap_cc_368_execute_5927_2_; 
wire _auto_iopadmap_cc_368_execute_5927_30_; 
wire _auto_iopadmap_cc_368_execute_5927_31_; 
wire _auto_iopadmap_cc_368_execute_5927_3_; 
wire _auto_iopadmap_cc_368_execute_5927_4_; 
wire _auto_iopadmap_cc_368_execute_5927_5_; 
wire _auto_iopadmap_cc_368_execute_5927_6_; 
wire _auto_iopadmap_cc_368_execute_5927_7_; 
wire _auto_iopadmap_cc_368_execute_5927_8_; 
wire _auto_iopadmap_cc_368_execute_5927_9_; 
wire _auto_iopadmap_cc_368_execute_5960; 
output align;
output \arprot[0] ;
output \arprot[1] ;
output \arprot[2] ;
output \awprot[0] ;
output \awprot[1] ;
output \awprot[2] ;
output busy;
input clock;
wire clock_bF_buf0; 
wire clock_bF_buf1; 
wire clock_bF_buf2; 
wire clock_bF_buf3; 
wire clock_bF_buf4; 
wire clock_bF_buf5; 
wire clock_bF_buf6; 
wire clock_bF_buf7; 
output done;
wire en_instr; 
input enable;
input \imm[0] ;
input \imm[10] ;
input \imm[11] ;
input \imm[12] ;
input \imm[13] ;
input \imm[14] ;
input \imm[15] ;
input \imm[16] ;
input \imm[17] ;
input \imm[18] ;
input \imm[19] ;
input \imm[1] ;
input \imm[20] ;
input \imm[21] ;
input \imm[22] ;
input \imm[23] ;
input \imm[24] ;
input \imm[25] ;
input \imm[26] ;
input \imm[27] ;
input \imm[28] ;
input \imm[29] ;
input \imm[2] ;
input \imm[30] ;
input \imm[31] ;
input \imm[3] ;
input \imm[4] ;
input \imm[5] ;
input \imm[6] ;
input \imm[7] ;
input \imm[8] ;
input \imm[9] ;
output \inst[0] ;
output \inst[10] ;
output \inst[11] ;
output \inst[12] ;
output \inst[13] ;
output \inst[14] ;
output \inst[15] ;
output \inst[16] ;
output \inst[17] ;
output \inst[18] ;
output \inst[19] ;
output \inst[1] ;
output \inst[20] ;
output \inst[21] ;
output \inst[22] ;
output \inst[23] ;
output \inst[24] ;
output \inst[25] ;
output \inst[26] ;
output \inst[27] ;
output \inst[28] ;
output \inst[29] ;
output \inst[2] ;
output \inst[30] ;
output \inst[31] ;
output \inst[3] ;
output \inst[4] ;
output \inst[5] ;
output \inst[6] ;
output \inst[7] ;
output \inst[8] ;
output \inst[9] ;
input \pc[0] ;
input \pc[10] ;
input \pc[11] ;
input \pc[12] ;
input \pc[13] ;
input \pc[14] ;
input \pc[15] ;
input \pc[16] ;
input \pc[17] ;
input \pc[18] ;
input \pc[19] ;
input \pc[1] ;
input \pc[20] ;
input \pc[21] ;
input \pc[22] ;
input \pc[23] ;
input \pc[24] ;
input \pc[25] ;
input \pc[26] ;
input \pc[27] ;
input \pc[28] ;
input \pc[29] ;
input \pc[2] ;
input \pc[30] ;
input \pc[31] ;
input \pc[3] ;
input \pc[4] ;
input \pc[5] ;
input \pc[6] ;
input \pc[7] ;
input \pc[8] ;
input \pc[9] ;
output \rd[0] ;
output \rd[10] ;
output \rd[11] ;
output \rd[12] ;
output \rd[13] ;
output \rd[14] ;
output \rd[15] ;
output \rd[16] ;
output \rd[17] ;
output \rd[18] ;
output \rd[19] ;
output \rd[1] ;
output \rd[20] ;
output \rd[21] ;
output \rd[22] ;
output \rd[23] ;
output \rd[24] ;
output \rd[25] ;
output \rd[26] ;
output \rd[27] ;
output \rd[28] ;
output \rd[29] ;
output \rd[2] ;
output \rd[30] ;
output \rd[31] ;
output \rd[3] ;
output \rd[4] ;
output \rd[5] ;
output \rd[6] ;
output \rd[7] ;
output \rd[8] ;
output \rd[9] ;
output rd_en;
input resetn;
wire resetn_bF_buf0; 
wire resetn_bF_buf1; 
wire resetn_bF_buf2; 
wire resetn_bF_buf3; 
wire resetn_bF_buf4; 
wire resetn_bF_buf5; 
input \rs1[0] ;
input \rs1[10] ;
input \rs1[11] ;
input \rs1[12] ;
input \rs1[13] ;
input \rs1[14] ;
input \rs1[15] ;
input \rs1[16] ;
input \rs1[17] ;
input \rs1[18] ;
input \rs1[19] ;
input \rs1[1] ;
input \rs1[20] ;
input \rs1[21] ;
input \rs1[22] ;
input \rs1[23] ;
input \rs1[24] ;
input \rs1[25] ;
input \rs1[26] ;
input \rs1[27] ;
input \rs1[28] ;
input \rs1[29] ;
input \rs1[2] ;
input \rs1[30] ;
input \rs1[31] ;
input \rs1[3] ;
input \rs1[4] ;
input \rs1[5] ;
input \rs1[6] ;
input \rs1[7] ;
input \rs1[8] ;
input \rs1[9] ;
input \rs2[0] ;
input \rs2[10] ;
input \rs2[11] ;
input \rs2[12] ;
input \rs2[13] ;
input \rs2[14] ;
input \rs2[15] ;
input \rs2[16] ;
input \rs2[17] ;
input \rs2[18] ;
input \rs2[19] ;
input \rs2[1] ;
input \rs2[20] ;
input \rs2[21] ;
input \rs2[22] ;
input \rs2[23] ;
input \rs2[24] ;
input \rs2[25] ;
input \rs2[26] ;
input \rs2[27] ;
input \rs2[28] ;
input \rs2[29] ;
input \rs2[2] ;
input \rs2[30] ;
input \rs2[31] ;
input \rs2[3] ;
input \rs2[4] ;
input \rs2[5] ;
input \rs2[6] ;
input \rs2[7] ;
input \rs2[8] ;
input \rs2[9] ;
input signo;
wire state_0_; 
wire state_1_; 
wire state_2_; 
wire state_3_; 
wire state_4_; 
wire state_5_; 
wire state_6_; 
input \wordsize[0] ;
input \wordsize[1] ;
AND2X2 AND2X2_1 ( .A(Wready), .B(state_3_), .Y(_abc_4635_new_n362_));
AND2X2 AND2X2_10 ( .A(_abc_4635_new_n378_), .B(resetn_bF_buf3), .Y(_abc_4635_new_n379_));
AND2X2 AND2X2_100 ( .A(_abc_4635_new_n531_), .B(_abc_4635_new_n457_), .Y(_abc_4635_new_n532_));
AND2X2 AND2X2_101 ( .A(_abc_4635_new_n512_), .B(\rs2[12] ), .Y(_abc_4635_new_n533_));
AND2X2 AND2X2_102 ( .A(_abc_4635_new_n534_), .B(_abc_4635_new_n485__bF_buf4), .Y(_0Wdata_31_0__12_));
AND2X2 AND2X2_103 ( .A(_abc_4635_new_n458_), .B(\rs2[5] ), .Y(_abc_4635_new_n536_));
AND2X2 AND2X2_104 ( .A(_abc_4635_new_n536_), .B(_abc_4635_new_n457_), .Y(_abc_4635_new_n537_));
AND2X2 AND2X2_105 ( .A(_abc_4635_new_n512_), .B(\rs2[13] ), .Y(_abc_4635_new_n538_));
AND2X2 AND2X2_106 ( .A(_abc_4635_new_n539_), .B(_abc_4635_new_n485__bF_buf3), .Y(_0Wdata_31_0__13_));
AND2X2 AND2X2_107 ( .A(_abc_4635_new_n458_), .B(\rs2[6] ), .Y(_abc_4635_new_n541_));
AND2X2 AND2X2_108 ( .A(_abc_4635_new_n541_), .B(_abc_4635_new_n457_), .Y(_abc_4635_new_n542_));
AND2X2 AND2X2_109 ( .A(_abc_4635_new_n512_), .B(\rs2[14] ), .Y(_abc_4635_new_n543_));
AND2X2 AND2X2_11 ( .A(enable), .B(state_0_), .Y(_abc_4635_new_n381_));
AND2X2 AND2X2_110 ( .A(_abc_4635_new_n544_), .B(_abc_4635_new_n485__bF_buf2), .Y(_0Wdata_31_0__14_));
AND2X2 AND2X2_111 ( .A(_abc_4635_new_n458_), .B(\rs2[7] ), .Y(_abc_4635_new_n546_));
AND2X2 AND2X2_112 ( .A(_abc_4635_new_n546_), .B(_abc_4635_new_n457_), .Y(_abc_4635_new_n547_));
AND2X2 AND2X2_113 ( .A(_abc_4635_new_n512_), .B(\rs2[15] ), .Y(_abc_4635_new_n548_));
AND2X2 AND2X2_114 ( .A(_abc_4635_new_n549_), .B(_abc_4635_new_n485__bF_buf1), .Y(_0Wdata_31_0__15_));
AND2X2 AND2X2_115 ( .A(_abc_4635_new_n511__bF_buf5), .B(\rs2[16] ), .Y(_abc_4635_new_n551_));
AND2X2 AND2X2_116 ( .A(_abc_4635_new_n552_), .B(_abc_4635_new_n485__bF_buf0), .Y(_0Wdata_31_0__16_));
AND2X2 AND2X2_117 ( .A(_abc_4635_new_n511__bF_buf4), .B(\rs2[17] ), .Y(_abc_4635_new_n554_));
AND2X2 AND2X2_118 ( .A(_abc_4635_new_n555_), .B(_abc_4635_new_n485__bF_buf4), .Y(_0Wdata_31_0__17_));
AND2X2 AND2X2_119 ( .A(_abc_4635_new_n511__bF_buf3), .B(\rs2[18] ), .Y(_abc_4635_new_n557_));
AND2X2 AND2X2_12 ( .A(_abc_4635_new_n380_), .B(_abc_4635_new_n381_), .Y(_abc_4635_new_n382_));
AND2X2 AND2X2_120 ( .A(_abc_4635_new_n558_), .B(_abc_4635_new_n485__bF_buf3), .Y(_0Wdata_31_0__18_));
AND2X2 AND2X2_121 ( .A(_abc_4635_new_n511__bF_buf2), .B(\rs2[19] ), .Y(_abc_4635_new_n560_));
AND2X2 AND2X2_122 ( .A(_abc_4635_new_n561_), .B(_abc_4635_new_n485__bF_buf2), .Y(_0Wdata_31_0__19_));
AND2X2 AND2X2_123 ( .A(_abc_4635_new_n511__bF_buf1), .B(\rs2[20] ), .Y(_abc_4635_new_n563_));
AND2X2 AND2X2_124 ( .A(_abc_4635_new_n564_), .B(_abc_4635_new_n485__bF_buf1), .Y(_0Wdata_31_0__20_));
AND2X2 AND2X2_125 ( .A(_abc_4635_new_n511__bF_buf0), .B(\rs2[21] ), .Y(_abc_4635_new_n566_));
AND2X2 AND2X2_126 ( .A(_abc_4635_new_n567_), .B(_abc_4635_new_n485__bF_buf0), .Y(_0Wdata_31_0__21_));
AND2X2 AND2X2_127 ( .A(_abc_4635_new_n511__bF_buf6), .B(\rs2[22] ), .Y(_abc_4635_new_n569_));
AND2X2 AND2X2_128 ( .A(_abc_4635_new_n570_), .B(_abc_4635_new_n485__bF_buf4), .Y(_0Wdata_31_0__22_));
AND2X2 AND2X2_129 ( .A(_abc_4635_new_n511__bF_buf5), .B(\rs2[23] ), .Y(_abc_4635_new_n572_));
AND2X2 AND2X2_13 ( .A(_abc_4635_new_n379_), .B(_abc_4635_new_n382_), .Y(_abc_4635_new_n383_));
AND2X2 AND2X2_130 ( .A(_abc_4635_new_n573_), .B(_abc_4635_new_n485__bF_buf3), .Y(_0Wdata_31_0__23_));
AND2X2 AND2X2_131 ( .A(_abc_4635_new_n480__bF_buf2), .B(\rs2[8] ), .Y(_abc_4635_new_n575_));
AND2X2 AND2X2_132 ( .A(_abc_4635_new_n511__bF_buf4), .B(\rs2[24] ), .Y(_abc_4635_new_n577_));
AND2X2 AND2X2_133 ( .A(_abc_4635_new_n578_), .B(_abc_4635_new_n485__bF_buf2), .Y(_0Wdata_31_0__24_));
AND2X2 AND2X2_134 ( .A(_abc_4635_new_n480__bF_buf1), .B(\rs2[9] ), .Y(_abc_4635_new_n580_));
AND2X2 AND2X2_135 ( .A(_abc_4635_new_n511__bF_buf3), .B(\rs2[25] ), .Y(_abc_4635_new_n582_));
AND2X2 AND2X2_136 ( .A(_abc_4635_new_n583_), .B(_abc_4635_new_n485__bF_buf1), .Y(_0Wdata_31_0__25_));
AND2X2 AND2X2_137 ( .A(_abc_4635_new_n480__bF_buf0), .B(\rs2[10] ), .Y(_abc_4635_new_n585_));
AND2X2 AND2X2_138 ( .A(_abc_4635_new_n511__bF_buf2), .B(\rs2[26] ), .Y(_abc_4635_new_n587_));
AND2X2 AND2X2_139 ( .A(_abc_4635_new_n588_), .B(_abc_4635_new_n485__bF_buf0), .Y(_0Wdata_31_0__26_));
AND2X2 AND2X2_14 ( .A(_abc_4635_new_n383_), .B(_abc_4635_new_n375_), .Y(_abc_4635_new_n384_));
AND2X2 AND2X2_140 ( .A(_abc_4635_new_n480__bF_buf4), .B(\rs2[11] ), .Y(_abc_4635_new_n590_));
AND2X2 AND2X2_141 ( .A(_abc_4635_new_n511__bF_buf1), .B(\rs2[27] ), .Y(_abc_4635_new_n592_));
AND2X2 AND2X2_142 ( .A(_abc_4635_new_n593_), .B(_abc_4635_new_n485__bF_buf4), .Y(_0Wdata_31_0__27_));
AND2X2 AND2X2_143 ( .A(_abc_4635_new_n480__bF_buf3), .B(\rs2[12] ), .Y(_abc_4635_new_n595_));
AND2X2 AND2X2_144 ( .A(_abc_4635_new_n511__bF_buf0), .B(\rs2[28] ), .Y(_abc_4635_new_n597_));
AND2X2 AND2X2_145 ( .A(_abc_4635_new_n598_), .B(_abc_4635_new_n485__bF_buf3), .Y(_0Wdata_31_0__28_));
AND2X2 AND2X2_146 ( .A(_abc_4635_new_n480__bF_buf2), .B(\rs2[13] ), .Y(_abc_4635_new_n600_));
AND2X2 AND2X2_147 ( .A(_abc_4635_new_n511__bF_buf6), .B(\rs2[29] ), .Y(_abc_4635_new_n602_));
AND2X2 AND2X2_148 ( .A(_abc_4635_new_n603_), .B(_abc_4635_new_n485__bF_buf2), .Y(_0Wdata_31_0__29_));
AND2X2 AND2X2_149 ( .A(_abc_4635_new_n480__bF_buf1), .B(\rs2[14] ), .Y(_abc_4635_new_n605_));
AND2X2 AND2X2_15 ( .A(_abc_4635_new_n385_), .B(_abc_4635_new_n367_), .Y(_abc_4635_new_n386_));
AND2X2 AND2X2_150 ( .A(_abc_4635_new_n511__bF_buf5), .B(\rs2[30] ), .Y(_abc_4635_new_n607_));
AND2X2 AND2X2_151 ( .A(_abc_4635_new_n608_), .B(_abc_4635_new_n485__bF_buf1), .Y(_0Wdata_31_0__30_));
AND2X2 AND2X2_152 ( .A(_abc_4635_new_n480__bF_buf0), .B(\rs2[15] ), .Y(_abc_4635_new_n610_));
AND2X2 AND2X2_153 ( .A(_abc_4635_new_n511__bF_buf4), .B(\rs2[31] ), .Y(_abc_4635_new_n612_));
AND2X2 AND2X2_154 ( .A(_abc_4635_new_n613_), .B(_abc_4635_new_n485__bF_buf0), .Y(_0Wdata_31_0__31_));
AND2X2 AND2X2_155 ( .A(_abc_4635_new_n411_), .B(resetn_bF_buf1), .Y(_abc_4635_new_n615_));
AND2X2 AND2X2_156 ( .A(_abc_4635_new_n615_), .B(W_R_1_bF_buf4_), .Y(_abc_4635_new_n616_));
AND2X2 AND2X2_157 ( .A(_abc_4635_new_n616__bF_buf4), .B(\Rdata_mem[0] ), .Y(_abc_4635_new_n617_));
AND2X2 AND2X2_158 ( .A(_abc_4635_new_n618__bF_buf4), .B(_auto_iopadmap_cc_368_execute_5894_0_), .Y(_abc_4635_new_n619_));
AND2X2 AND2X2_159 ( .A(_abc_4635_new_n620_), .B(resetn_bF_buf0), .Y(_0inst_31_0__0_));
AND2X2 AND2X2_16 ( .A(_abc_4635_new_n387_), .B(_abc_4635_new_n361_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_1_));
AND2X2 AND2X2_160 ( .A(_abc_4635_new_n616__bF_buf2), .B(\Rdata_mem[1] ), .Y(_abc_4635_new_n622_));
AND2X2 AND2X2_161 ( .A(_abc_4635_new_n618__bF_buf3), .B(_auto_iopadmap_cc_368_execute_5894_1_), .Y(_abc_4635_new_n623_));
AND2X2 AND2X2_162 ( .A(_abc_4635_new_n624_), .B(resetn_bF_buf5), .Y(_0inst_31_0__1_));
AND2X2 AND2X2_163 ( .A(_abc_4635_new_n616__bF_buf1), .B(\Rdata_mem[2] ), .Y(_abc_4635_new_n626_));
AND2X2 AND2X2_164 ( .A(_abc_4635_new_n618__bF_buf2), .B(_auto_iopadmap_cc_368_execute_5894_2_), .Y(_abc_4635_new_n627_));
AND2X2 AND2X2_165 ( .A(_abc_4635_new_n628_), .B(resetn_bF_buf4), .Y(_0inst_31_0__2_));
AND2X2 AND2X2_166 ( .A(_abc_4635_new_n616__bF_buf0), .B(\Rdata_mem[3] ), .Y(_abc_4635_new_n630_));
AND2X2 AND2X2_167 ( .A(_abc_4635_new_n618__bF_buf1), .B(_auto_iopadmap_cc_368_execute_5894_3_), .Y(_abc_4635_new_n631_));
AND2X2 AND2X2_168 ( .A(_abc_4635_new_n632_), .B(resetn_bF_buf3), .Y(_0inst_31_0__3_));
AND2X2 AND2X2_169 ( .A(_abc_4635_new_n616__bF_buf4), .B(\Rdata_mem[4] ), .Y(_abc_4635_new_n634_));
AND2X2 AND2X2_17 ( .A(ARready), .B(Rvalid), .Y(_abc_4635_new_n390_));
AND2X2 AND2X2_170 ( .A(_abc_4635_new_n618__bF_buf0), .B(_auto_iopadmap_cc_368_execute_5894_4_), .Y(_abc_4635_new_n635_));
AND2X2 AND2X2_171 ( .A(_abc_4635_new_n636_), .B(resetn_bF_buf2), .Y(_0inst_31_0__4_));
AND2X2 AND2X2_172 ( .A(_abc_4635_new_n616__bF_buf3), .B(\Rdata_mem[5] ), .Y(_abc_4635_new_n638_));
AND2X2 AND2X2_173 ( .A(_abc_4635_new_n618__bF_buf4), .B(_auto_iopadmap_cc_368_execute_5894_5_), .Y(_abc_4635_new_n639_));
AND2X2 AND2X2_174 ( .A(_abc_4635_new_n640_), .B(resetn_bF_buf1), .Y(_0inst_31_0__5_));
AND2X2 AND2X2_175 ( .A(_abc_4635_new_n616__bF_buf2), .B(\Rdata_mem[6] ), .Y(_abc_4635_new_n642_));
AND2X2 AND2X2_176 ( .A(_abc_4635_new_n618__bF_buf3), .B(_auto_iopadmap_cc_368_execute_5894_6_), .Y(_abc_4635_new_n643_));
AND2X2 AND2X2_177 ( .A(_abc_4635_new_n644_), .B(resetn_bF_buf0), .Y(_0inst_31_0__6_));
AND2X2 AND2X2_178 ( .A(_abc_4635_new_n616__bF_buf1), .B(\Rdata_mem[7] ), .Y(_abc_4635_new_n646_));
AND2X2 AND2X2_179 ( .A(_abc_4635_new_n618__bF_buf2), .B(_auto_iopadmap_cc_368_execute_5894_7_), .Y(_abc_4635_new_n647_));
AND2X2 AND2X2_18 ( .A(_abc_4635_new_n391_), .B(state_2_), .Y(_abc_4635_new_n392_));
AND2X2 AND2X2_180 ( .A(_abc_4635_new_n648_), .B(resetn_bF_buf5), .Y(_0inst_31_0__7_));
AND2X2 AND2X2_181 ( .A(_abc_4635_new_n616__bF_buf0), .B(\Rdata_mem[8] ), .Y(_abc_4635_new_n650_));
AND2X2 AND2X2_182 ( .A(_abc_4635_new_n618__bF_buf1), .B(_auto_iopadmap_cc_368_execute_5894_8_), .Y(_abc_4635_new_n651_));
AND2X2 AND2X2_183 ( .A(_abc_4635_new_n652_), .B(resetn_bF_buf4), .Y(_0inst_31_0__8_));
AND2X2 AND2X2_184 ( .A(_abc_4635_new_n616__bF_buf4), .B(\Rdata_mem[9] ), .Y(_abc_4635_new_n654_));
AND2X2 AND2X2_185 ( .A(_abc_4635_new_n618__bF_buf0), .B(_auto_iopadmap_cc_368_execute_5894_9_), .Y(_abc_4635_new_n655_));
AND2X2 AND2X2_186 ( .A(_abc_4635_new_n656_), .B(resetn_bF_buf3), .Y(_0inst_31_0__9_));
AND2X2 AND2X2_187 ( .A(_abc_4635_new_n616__bF_buf3), .B(\Rdata_mem[10] ), .Y(_abc_4635_new_n658_));
AND2X2 AND2X2_188 ( .A(_abc_4635_new_n618__bF_buf4), .B(_auto_iopadmap_cc_368_execute_5894_10_), .Y(_abc_4635_new_n659_));
AND2X2 AND2X2_189 ( .A(_abc_4635_new_n660_), .B(resetn_bF_buf2), .Y(_0inst_31_0__10_));
AND2X2 AND2X2_19 ( .A(_abc_4635_new_n376_), .B(_abc_4635_new_n381_), .Y(_abc_4635_new_n393_));
AND2X2 AND2X2_190 ( .A(_abc_4635_new_n616__bF_buf2), .B(\Rdata_mem[11] ), .Y(_abc_4635_new_n662_));
AND2X2 AND2X2_191 ( .A(_abc_4635_new_n618__bF_buf3), .B(_auto_iopadmap_cc_368_execute_5894_11_), .Y(_abc_4635_new_n663_));
AND2X2 AND2X2_192 ( .A(_abc_4635_new_n664_), .B(resetn_bF_buf1), .Y(_0inst_31_0__11_));
AND2X2 AND2X2_193 ( .A(_abc_4635_new_n616__bF_buf1), .B(\Rdata_mem[12] ), .Y(_abc_4635_new_n666_));
AND2X2 AND2X2_194 ( .A(_abc_4635_new_n618__bF_buf2), .B(_auto_iopadmap_cc_368_execute_5894_12_), .Y(_abc_4635_new_n667_));
AND2X2 AND2X2_195 ( .A(_abc_4635_new_n668_), .B(resetn_bF_buf0), .Y(_0inst_31_0__12_));
AND2X2 AND2X2_196 ( .A(_abc_4635_new_n616__bF_buf0), .B(\Rdata_mem[13] ), .Y(_abc_4635_new_n670_));
AND2X2 AND2X2_197 ( .A(_abc_4635_new_n618__bF_buf1), .B(_auto_iopadmap_cc_368_execute_5894_13_), .Y(_abc_4635_new_n671_));
AND2X2 AND2X2_198 ( .A(_abc_4635_new_n672_), .B(resetn_bF_buf5), .Y(_0inst_31_0__13_));
AND2X2 AND2X2_199 ( .A(_abc_4635_new_n616__bF_buf4), .B(\Rdata_mem[14] ), .Y(_abc_4635_new_n674_));
AND2X2 AND2X2_2 ( .A(state_6_), .B(AWready), .Y(_abc_4635_new_n363_));
AND2X2 AND2X2_20 ( .A(_abc_4635_new_n394_), .B(resetn_bF_buf2), .Y(_abc_4635_new_n395_));
AND2X2 AND2X2_200 ( .A(_abc_4635_new_n618__bF_buf0), .B(_auto_iopadmap_cc_368_execute_5894_14_), .Y(_abc_4635_new_n675_));
AND2X2 AND2X2_201 ( .A(_abc_4635_new_n676_), .B(resetn_bF_buf4), .Y(_0inst_31_0__14_));
AND2X2 AND2X2_202 ( .A(_abc_4635_new_n616__bF_buf3), .B(\Rdata_mem[15] ), .Y(_abc_4635_new_n678_));
AND2X2 AND2X2_203 ( .A(_abc_4635_new_n618__bF_buf4), .B(_auto_iopadmap_cc_368_execute_5894_15_), .Y(_abc_4635_new_n679_));
AND2X2 AND2X2_204 ( .A(_abc_4635_new_n680_), .B(resetn_bF_buf3), .Y(_0inst_31_0__15_));
AND2X2 AND2X2_205 ( .A(_abc_4635_new_n616__bF_buf2), .B(\Rdata_mem[16] ), .Y(_abc_4635_new_n682_));
AND2X2 AND2X2_206 ( .A(_abc_4635_new_n618__bF_buf3), .B(_auto_iopadmap_cc_368_execute_5894_16_), .Y(_abc_4635_new_n683_));
AND2X2 AND2X2_207 ( .A(_abc_4635_new_n684_), .B(resetn_bF_buf2), .Y(_0inst_31_0__16_));
AND2X2 AND2X2_208 ( .A(_abc_4635_new_n616__bF_buf1), .B(\Rdata_mem[17] ), .Y(_abc_4635_new_n686_));
AND2X2 AND2X2_209 ( .A(_abc_4635_new_n618__bF_buf2), .B(_auto_iopadmap_cc_368_execute_5894_17_), .Y(_abc_4635_new_n687_));
AND2X2 AND2X2_21 ( .A(_abc_4635_new_n395_), .B(_abc_4635_new_n389_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_2_));
AND2X2 AND2X2_210 ( .A(_abc_4635_new_n688_), .B(resetn_bF_buf1), .Y(_0inst_31_0__17_));
AND2X2 AND2X2_211 ( .A(_abc_4635_new_n616__bF_buf0), .B(\Rdata_mem[18] ), .Y(_abc_4635_new_n690_));
AND2X2 AND2X2_212 ( .A(_abc_4635_new_n618__bF_buf1), .B(_auto_iopadmap_cc_368_execute_5894_18_), .Y(_abc_4635_new_n691_));
AND2X2 AND2X2_213 ( .A(_abc_4635_new_n692_), .B(resetn_bF_buf0), .Y(_0inst_31_0__18_));
AND2X2 AND2X2_214 ( .A(_abc_4635_new_n616__bF_buf4), .B(\Rdata_mem[19] ), .Y(_abc_4635_new_n694_));
AND2X2 AND2X2_215 ( .A(_abc_4635_new_n618__bF_buf0), .B(_auto_iopadmap_cc_368_execute_5894_19_), .Y(_abc_4635_new_n695_));
AND2X2 AND2X2_216 ( .A(_abc_4635_new_n696_), .B(resetn_bF_buf5), .Y(_0inst_31_0__19_));
AND2X2 AND2X2_217 ( .A(_abc_4635_new_n616__bF_buf3), .B(\Rdata_mem[20] ), .Y(_abc_4635_new_n698_));
AND2X2 AND2X2_218 ( .A(_abc_4635_new_n618__bF_buf4), .B(_auto_iopadmap_cc_368_execute_5894_20_), .Y(_abc_4635_new_n699_));
AND2X2 AND2X2_219 ( .A(_abc_4635_new_n700_), .B(resetn_bF_buf4), .Y(_0inst_31_0__20_));
AND2X2 AND2X2_22 ( .A(state_6_), .B(resetn_bF_buf1), .Y(_abc_4635_new_n397_));
AND2X2 AND2X2_220 ( .A(_abc_4635_new_n616__bF_buf2), .B(\Rdata_mem[21] ), .Y(_abc_4635_new_n702_));
AND2X2 AND2X2_221 ( .A(_abc_4635_new_n618__bF_buf3), .B(_auto_iopadmap_cc_368_execute_5894_21_), .Y(_abc_4635_new_n703_));
AND2X2 AND2X2_222 ( .A(_abc_4635_new_n704_), .B(resetn_bF_buf3), .Y(_0inst_31_0__21_));
AND2X2 AND2X2_223 ( .A(_abc_4635_new_n616__bF_buf1), .B(\Rdata_mem[22] ), .Y(_abc_4635_new_n706_));
AND2X2 AND2X2_224 ( .A(_abc_4635_new_n618__bF_buf2), .B(_auto_iopadmap_cc_368_execute_5894_22_), .Y(_abc_4635_new_n707_));
AND2X2 AND2X2_225 ( .A(_abc_4635_new_n708_), .B(resetn_bF_buf2), .Y(_0inst_31_0__22_));
AND2X2 AND2X2_226 ( .A(_abc_4635_new_n616__bF_buf0), .B(\Rdata_mem[23] ), .Y(_abc_4635_new_n710_));
AND2X2 AND2X2_227 ( .A(_abc_4635_new_n618__bF_buf1), .B(_auto_iopadmap_cc_368_execute_5894_23_), .Y(_abc_4635_new_n711_));
AND2X2 AND2X2_228 ( .A(_abc_4635_new_n712_), .B(resetn_bF_buf1), .Y(_0inst_31_0__23_));
AND2X2 AND2X2_229 ( .A(_abc_4635_new_n616__bF_buf4), .B(\Rdata_mem[24] ), .Y(_abc_4635_new_n714_));
AND2X2 AND2X2_23 ( .A(_abc_4635_new_n385_), .B(Wready), .Y(_abc_4635_new_n398_));
AND2X2 AND2X2_230 ( .A(_abc_4635_new_n618__bF_buf0), .B(_auto_iopadmap_cc_368_execute_5894_24_), .Y(_abc_4635_new_n715_));
AND2X2 AND2X2_231 ( .A(_abc_4635_new_n716_), .B(resetn_bF_buf0), .Y(_0inst_31_0__24_));
AND2X2 AND2X2_232 ( .A(_abc_4635_new_n616__bF_buf3), .B(\Rdata_mem[25] ), .Y(_abc_4635_new_n718_));
AND2X2 AND2X2_233 ( .A(_abc_4635_new_n618__bF_buf4), .B(_auto_iopadmap_cc_368_execute_5894_25_), .Y(_abc_4635_new_n719_));
AND2X2 AND2X2_234 ( .A(_abc_4635_new_n720_), .B(resetn_bF_buf5), .Y(_0inst_31_0__25_));
AND2X2 AND2X2_235 ( .A(_abc_4635_new_n616__bF_buf2), .B(\Rdata_mem[26] ), .Y(_abc_4635_new_n722_));
AND2X2 AND2X2_236 ( .A(_abc_4635_new_n618__bF_buf3), .B(_auto_iopadmap_cc_368_execute_5894_26_), .Y(_abc_4635_new_n723_));
AND2X2 AND2X2_237 ( .A(_abc_4635_new_n724_), .B(resetn_bF_buf4), .Y(_0inst_31_0__26_));
AND2X2 AND2X2_238 ( .A(_abc_4635_new_n616__bF_buf1), .B(\Rdata_mem[27] ), .Y(_abc_4635_new_n726_));
AND2X2 AND2X2_239 ( .A(_abc_4635_new_n618__bF_buf2), .B(_auto_iopadmap_cc_368_execute_5894_27_), .Y(_abc_4635_new_n727_));
AND2X2 AND2X2_24 ( .A(_abc_4635_new_n399_), .B(_abc_4635_new_n373_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_6_));
AND2X2 AND2X2_240 ( .A(_abc_4635_new_n728_), .B(resetn_bF_buf3), .Y(_0inst_31_0__27_));
AND2X2 AND2X2_241 ( .A(_abc_4635_new_n616__bF_buf0), .B(\Rdata_mem[28] ), .Y(_abc_4635_new_n730_));
AND2X2 AND2X2_242 ( .A(_abc_4635_new_n618__bF_buf1), .B(_auto_iopadmap_cc_368_execute_5894_28_), .Y(_abc_4635_new_n731_));
AND2X2 AND2X2_243 ( .A(_abc_4635_new_n732_), .B(resetn_bF_buf2), .Y(_0inst_31_0__28_));
AND2X2 AND2X2_244 ( .A(_abc_4635_new_n616__bF_buf4), .B(\Rdata_mem[29] ), .Y(_abc_4635_new_n734_));
AND2X2 AND2X2_245 ( .A(_abc_4635_new_n618__bF_buf0), .B(_auto_iopadmap_cc_368_execute_5894_29_), .Y(_abc_4635_new_n735_));
AND2X2 AND2X2_246 ( .A(_abc_4635_new_n736_), .B(resetn_bF_buf1), .Y(_0inst_31_0__29_));
AND2X2 AND2X2_247 ( .A(_abc_4635_new_n616__bF_buf3), .B(\Rdata_mem[30] ), .Y(_abc_4635_new_n738_));
AND2X2 AND2X2_248 ( .A(_abc_4635_new_n618__bF_buf4), .B(_auto_iopadmap_cc_368_execute_5894_30_), .Y(_abc_4635_new_n739_));
AND2X2 AND2X2_249 ( .A(_abc_4635_new_n740_), .B(resetn_bF_buf0), .Y(_0inst_31_0__30_));
AND2X2 AND2X2_25 ( .A(Bvalid), .B(AWready), .Y(_abc_4635_new_n402_));
AND2X2 AND2X2_250 ( .A(_abc_4635_new_n616__bF_buf2), .B(\Rdata_mem[31] ), .Y(_abc_4635_new_n742_));
AND2X2 AND2X2_251 ( .A(_abc_4635_new_n618__bF_buf3), .B(_auto_iopadmap_cc_368_execute_5894_31_), .Y(_abc_4635_new_n743_));
AND2X2 AND2X2_252 ( .A(_abc_4635_new_n744_), .B(resetn_bF_buf5), .Y(_0inst_31_0__31_));
AND2X2 AND2X2_253 ( .A(_abc_4635_new_n476_), .B(_abc_4635_new_n511__bF_buf3), .Y(_abc_4635_new_n746_));
AND2X2 AND2X2_254 ( .A(_abc_4635_new_n475_), .B(_abc_4635_new_n480__bF_buf4), .Y(_abc_4635_new_n747_));
AND2X2 AND2X2_255 ( .A(_abc_4635_new_n753__bF_buf4), .B(\W_R[0] ), .Y(_abc_4635_new_n754_));
AND2X2 AND2X2_256 ( .A(_abc_4635_new_n755_), .B(_abc_4635_new_n475_), .Y(_abc_4635_new_n756_));
AND2X2 AND2X2_257 ( .A(_abc_4635_new_n757_), .B(_abc_4635_new_n758_), .Y(_abc_4635_new_n759_));
AND2X2 AND2X2_258 ( .A(_abc_4635_new_n759_), .B(_abc_4635_new_n474_), .Y(_abc_4635_new_n760_));
AND2X2 AND2X2_259 ( .A(_abc_4635_new_n459_), .B(\Rdata_mem[0] ), .Y(_abc_4635_new_n762_));
AND2X2 AND2X2_26 ( .A(_abc_4635_new_n402_), .B(Wready), .Y(_abc_4635_new_n403_));
AND2X2 AND2X2_260 ( .A(_abc_4635_new_n761_), .B(_abc_4635_new_n763_), .Y(_abc_4635_new_n764_));
AND2X2 AND2X2_261 ( .A(_abc_4635_new_n511__bF_buf2), .B(\Rdata_mem[0] ), .Y(_abc_4635_new_n765_));
AND2X2 AND2X2_262 ( .A(_abc_4635_new_n755_), .B(_abc_4635_new_n480__bF_buf3), .Y(_abc_4635_new_n767_));
AND2X2 AND2X2_263 ( .A(_abc_4635_new_n767_), .B(_abc_4635_new_n766_), .Y(_abc_4635_new_n768_));
AND2X2 AND2X2_264 ( .A(_abc_4635_new_n770_), .B(_abc_4635_new_n754__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_5927_0_));
AND2X2 AND2X2_265 ( .A(_abc_4635_new_n772_), .B(_abc_4635_new_n773_), .Y(_abc_4635_new_n774_));
AND2X2 AND2X2_266 ( .A(_abc_4635_new_n774_), .B(_abc_4635_new_n474_), .Y(_abc_4635_new_n775_));
AND2X2 AND2X2_267 ( .A(_abc_4635_new_n776_), .B(_abc_4635_new_n475_), .Y(_abc_4635_new_n777_));
AND2X2 AND2X2_268 ( .A(_abc_4635_new_n459_), .B(\Rdata_mem[1] ), .Y(_abc_4635_new_n779_));
AND2X2 AND2X2_269 ( .A(_abc_4635_new_n778_), .B(_abc_4635_new_n780_), .Y(_abc_4635_new_n781_));
AND2X2 AND2X2_27 ( .A(_abc_4635_new_n403_), .B(_abc_4635_new_n380_), .Y(_abc_4635_new_n404_));
AND2X2 AND2X2_270 ( .A(_abc_4635_new_n511__bF_buf1), .B(\Rdata_mem[1] ), .Y(_abc_4635_new_n782_));
AND2X2 AND2X2_271 ( .A(_abc_4635_new_n776_), .B(_abc_4635_new_n480__bF_buf2), .Y(_abc_4635_new_n784_));
AND2X2 AND2X2_272 ( .A(_abc_4635_new_n784_), .B(_abc_4635_new_n783_), .Y(_abc_4635_new_n785_));
AND2X2 AND2X2_273 ( .A(_abc_4635_new_n787_), .B(_abc_4635_new_n754__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_5927_1_));
AND2X2 AND2X2_274 ( .A(_abc_4635_new_n789_), .B(_abc_4635_new_n790_), .Y(_abc_4635_new_n791_));
AND2X2 AND2X2_275 ( .A(_abc_4635_new_n791_), .B(_abc_4635_new_n474_), .Y(_abc_4635_new_n792_));
AND2X2 AND2X2_276 ( .A(_abc_4635_new_n793_), .B(_abc_4635_new_n475_), .Y(_abc_4635_new_n794_));
AND2X2 AND2X2_277 ( .A(_abc_4635_new_n459_), .B(\Rdata_mem[2] ), .Y(_abc_4635_new_n796_));
AND2X2 AND2X2_278 ( .A(_abc_4635_new_n795_), .B(_abc_4635_new_n797_), .Y(_abc_4635_new_n798_));
AND2X2 AND2X2_279 ( .A(_abc_4635_new_n511__bF_buf0), .B(\Rdata_mem[2] ), .Y(_abc_4635_new_n799_));
AND2X2 AND2X2_28 ( .A(_abc_4635_new_n405_), .B(state_0_), .Y(_abc_4635_new_n406_));
AND2X2 AND2X2_280 ( .A(_abc_4635_new_n793_), .B(_abc_4635_new_n480__bF_buf1), .Y(_abc_4635_new_n801_));
AND2X2 AND2X2_281 ( .A(_abc_4635_new_n801_), .B(_abc_4635_new_n800_), .Y(_abc_4635_new_n802_));
AND2X2 AND2X2_282 ( .A(_abc_4635_new_n804_), .B(_abc_4635_new_n754__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_5927_2_));
AND2X2 AND2X2_283 ( .A(_abc_4635_new_n806_), .B(_abc_4635_new_n807_), .Y(_abc_4635_new_n808_));
AND2X2 AND2X2_284 ( .A(_abc_4635_new_n808_), .B(_abc_4635_new_n474_), .Y(_abc_4635_new_n809_));
AND2X2 AND2X2_285 ( .A(_abc_4635_new_n810_), .B(_abc_4635_new_n475_), .Y(_abc_4635_new_n811_));
AND2X2 AND2X2_286 ( .A(_abc_4635_new_n459_), .B(\Rdata_mem[3] ), .Y(_abc_4635_new_n813_));
AND2X2 AND2X2_287 ( .A(_abc_4635_new_n812_), .B(_abc_4635_new_n814_), .Y(_abc_4635_new_n815_));
AND2X2 AND2X2_288 ( .A(_abc_4635_new_n511__bF_buf6), .B(\Rdata_mem[3] ), .Y(_abc_4635_new_n816_));
AND2X2 AND2X2_289 ( .A(_abc_4635_new_n810_), .B(_abc_4635_new_n480__bF_buf0), .Y(_abc_4635_new_n818_));
AND2X2 AND2X2_29 ( .A(_abc_4635_new_n393_), .B(_abc_4635_new_n390_), .Y(_abc_4635_new_n407_));
AND2X2 AND2X2_290 ( .A(_abc_4635_new_n818_), .B(_abc_4635_new_n817_), .Y(_abc_4635_new_n819_));
AND2X2 AND2X2_291 ( .A(_abc_4635_new_n821_), .B(_abc_4635_new_n754__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_5927_3_));
AND2X2 AND2X2_292 ( .A(_abc_4635_new_n823_), .B(_abc_4635_new_n475_), .Y(_abc_4635_new_n824_));
AND2X2 AND2X2_293 ( .A(_abc_4635_new_n825_), .B(_abc_4635_new_n826_), .Y(_abc_4635_new_n827_));
AND2X2 AND2X2_294 ( .A(_abc_4635_new_n827_), .B(_abc_4635_new_n474_), .Y(_abc_4635_new_n828_));
AND2X2 AND2X2_295 ( .A(_abc_4635_new_n459_), .B(\Rdata_mem[4] ), .Y(_abc_4635_new_n830_));
AND2X2 AND2X2_296 ( .A(_abc_4635_new_n829_), .B(_abc_4635_new_n831_), .Y(_abc_4635_new_n832_));
AND2X2 AND2X2_297 ( .A(_abc_4635_new_n511__bF_buf5), .B(\Rdata_mem[4] ), .Y(_abc_4635_new_n833_));
AND2X2 AND2X2_298 ( .A(_abc_4635_new_n823_), .B(_abc_4635_new_n480__bF_buf4), .Y(_abc_4635_new_n835_));
AND2X2 AND2X2_299 ( .A(_abc_4635_new_n835_), .B(_abc_4635_new_n834_), .Y(_abc_4635_new_n836_));
AND2X2 AND2X2_3 ( .A(_abc_4635_new_n365_), .B(resetn_bF_buf5), .Y(_abc_4635_new_n366_));
AND2X2 AND2X2_30 ( .A(_abc_4635_new_n390_), .B(state_2_), .Y(_abc_4635_new_n408_));
AND2X2 AND2X2_300 ( .A(_abc_4635_new_n838_), .B(_abc_4635_new_n754__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_5927_4_));
AND2X2 AND2X2_301 ( .A(_abc_4635_new_n840_), .B(_abc_4635_new_n475_), .Y(_abc_4635_new_n841_));
AND2X2 AND2X2_302 ( .A(_abc_4635_new_n842_), .B(_abc_4635_new_n843_), .Y(_abc_4635_new_n844_));
AND2X2 AND2X2_303 ( .A(_abc_4635_new_n844_), .B(_abc_4635_new_n474_), .Y(_abc_4635_new_n845_));
AND2X2 AND2X2_304 ( .A(_abc_4635_new_n459_), .B(\Rdata_mem[5] ), .Y(_abc_4635_new_n847_));
AND2X2 AND2X2_305 ( .A(_abc_4635_new_n846_), .B(_abc_4635_new_n848_), .Y(_abc_4635_new_n849_));
AND2X2 AND2X2_306 ( .A(_abc_4635_new_n511__bF_buf4), .B(\Rdata_mem[5] ), .Y(_abc_4635_new_n850_));
AND2X2 AND2X2_307 ( .A(_abc_4635_new_n840_), .B(_abc_4635_new_n480__bF_buf3), .Y(_abc_4635_new_n852_));
AND2X2 AND2X2_308 ( .A(_abc_4635_new_n852_), .B(_abc_4635_new_n851_), .Y(_abc_4635_new_n853_));
AND2X2 AND2X2_309 ( .A(_abc_4635_new_n855_), .B(_abc_4635_new_n754__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_5927_5_));
AND2X2 AND2X2_31 ( .A(Rvalid), .B(state_5_), .Y(_abc_4635_new_n409_));
AND2X2 AND2X2_310 ( .A(_abc_4635_new_n857_), .B(_abc_4635_new_n858_), .Y(_abc_4635_new_n859_));
AND2X2 AND2X2_311 ( .A(_abc_4635_new_n859_), .B(_abc_4635_new_n474_), .Y(_abc_4635_new_n860_));
AND2X2 AND2X2_312 ( .A(_abc_4635_new_n861_), .B(_abc_4635_new_n475_), .Y(_abc_4635_new_n862_));
AND2X2 AND2X2_313 ( .A(_abc_4635_new_n459_), .B(\Rdata_mem[6] ), .Y(_abc_4635_new_n864_));
AND2X2 AND2X2_314 ( .A(_abc_4635_new_n863_), .B(_abc_4635_new_n865_), .Y(_abc_4635_new_n866_));
AND2X2 AND2X2_315 ( .A(_abc_4635_new_n511__bF_buf3), .B(\Rdata_mem[6] ), .Y(_abc_4635_new_n867_));
AND2X2 AND2X2_316 ( .A(_abc_4635_new_n861_), .B(_abc_4635_new_n480__bF_buf2), .Y(_abc_4635_new_n869_));
AND2X2 AND2X2_317 ( .A(_abc_4635_new_n869_), .B(_abc_4635_new_n868_), .Y(_abc_4635_new_n870_));
AND2X2 AND2X2_318 ( .A(_abc_4635_new_n872_), .B(_abc_4635_new_n754__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_5927_6_));
AND2X2 AND2X2_319 ( .A(_abc_4635_new_n472__bF_buf1), .B(_abc_4635_new_n474_), .Y(_abc_4635_new_n874_));
AND2X2 AND2X2_32 ( .A(_abc_4635_new_n365_), .B(Bvalid), .Y(_abc_4635_new_n412_));
AND2X2 AND2X2_320 ( .A(_abc_4635_new_n874_), .B(\Rdata_mem[15] ), .Y(_abc_4635_new_n875_));
AND2X2 AND2X2_321 ( .A(_abc_4635_new_n493__bF_buf3), .B(_abc_4635_new_n475_), .Y(_abc_4635_new_n876_));
AND2X2 AND2X2_322 ( .A(_abc_4635_new_n876_), .B(\Rdata_mem[23] ), .Y(_abc_4635_new_n877_));
AND2X2 AND2X2_323 ( .A(_abc_4635_new_n493__bF_buf2), .B(_abc_4635_new_n474_), .Y(_abc_4635_new_n879_));
AND2X2 AND2X2_324 ( .A(_abc_4635_new_n879_), .B(\Rdata_mem[31] ), .Y(_abc_4635_new_n880_));
AND2X2 AND2X2_325 ( .A(_abc_4635_new_n476_), .B(\Rdata_mem[7] ), .Y(_abc_4635_new_n881_));
AND2X2 AND2X2_326 ( .A(_abc_4635_new_n883_), .B(_abc_4635_new_n459_), .Y(_abc_4635_new_n884_));
AND2X2 AND2X2_327 ( .A(_abc_4635_new_n511__bF_buf2), .B(\Rdata_mem[7] ), .Y(_abc_4635_new_n885_));
AND2X2 AND2X2_328 ( .A(_abc_4635_new_n887_), .B(_abc_4635_new_n480__bF_buf1), .Y(_abc_4635_new_n888_));
AND2X2 AND2X2_329 ( .A(_abc_4635_new_n888_), .B(_abc_4635_new_n886_), .Y(_abc_4635_new_n889_));
AND2X2 AND2X2_33 ( .A(_abc_4635_new_n403_), .B(_abc_4635_new_n371_), .Y(_abc_4635_new_n414_));
AND2X2 AND2X2_330 ( .A(_abc_4635_new_n891_), .B(_abc_4635_new_n754__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_5927_7_));
AND2X2 AND2X2_331 ( .A(_abc_4635_new_n459_), .B(signo), .Y(_abc_4635_new_n893_));
AND2X2 AND2X2_332 ( .A(_abc_4635_new_n883_), .B(_abc_4635_new_n893_), .Y(_abc_4635_new_n894_));
AND2X2 AND2X2_333 ( .A(_abc_4635_new_n511__bF_buf1), .B(\Rdata_mem[8] ), .Y(_abc_4635_new_n895_));
AND2X2 AND2X2_334 ( .A(_abc_4635_new_n759_), .B(_abc_4635_new_n480__bF_buf0), .Y(_abc_4635_new_n896_));
AND2X2 AND2X2_335 ( .A(_abc_4635_new_n898_), .B(_abc_4635_new_n754__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_5927_8_));
AND2X2 AND2X2_336 ( .A(_abc_4635_new_n511__bF_buf0), .B(\Rdata_mem[9] ), .Y(_abc_4635_new_n900_));
AND2X2 AND2X2_337 ( .A(_abc_4635_new_n774_), .B(_abc_4635_new_n480__bF_buf4), .Y(_abc_4635_new_n901_));
AND2X2 AND2X2_338 ( .A(_abc_4635_new_n903_), .B(_abc_4635_new_n754__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_5927_9_));
AND2X2 AND2X2_339 ( .A(_abc_4635_new_n511__bF_buf6), .B(\Rdata_mem[10] ), .Y(_abc_4635_new_n905_));
AND2X2 AND2X2_34 ( .A(_abc_4635_new_n383_), .B(_abc_4635_new_n369_), .Y(_abc_4635_new_n419_));
AND2X2 AND2X2_340 ( .A(_abc_4635_new_n791_), .B(_abc_4635_new_n480__bF_buf3), .Y(_abc_4635_new_n906_));
AND2X2 AND2X2_341 ( .A(_abc_4635_new_n908_), .B(_abc_4635_new_n754__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_5927_10_));
AND2X2 AND2X2_342 ( .A(_abc_4635_new_n511__bF_buf5), .B(\Rdata_mem[11] ), .Y(_abc_4635_new_n910_));
AND2X2 AND2X2_343 ( .A(_abc_4635_new_n808_), .B(_abc_4635_new_n480__bF_buf2), .Y(_abc_4635_new_n911_));
AND2X2 AND2X2_344 ( .A(_abc_4635_new_n913_), .B(_abc_4635_new_n754__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_5927_11_));
AND2X2 AND2X2_345 ( .A(_abc_4635_new_n511__bF_buf4), .B(\Rdata_mem[12] ), .Y(_abc_4635_new_n915_));
AND2X2 AND2X2_346 ( .A(_abc_4635_new_n827_), .B(_abc_4635_new_n480__bF_buf1), .Y(_abc_4635_new_n916_));
AND2X2 AND2X2_347 ( .A(_abc_4635_new_n918_), .B(_abc_4635_new_n754__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_5927_12_));
AND2X2 AND2X2_348 ( .A(_abc_4635_new_n511__bF_buf3), .B(\Rdata_mem[13] ), .Y(_abc_4635_new_n920_));
AND2X2 AND2X2_349 ( .A(_abc_4635_new_n844_), .B(_abc_4635_new_n480__bF_buf0), .Y(_abc_4635_new_n921_));
AND2X2 AND2X2_35 ( .A(_abc_4635_new_n368_), .B(resetn_bF_buf5), .Y(_abc_4635_new_n420_));
AND2X2 AND2X2_350 ( .A(_abc_4635_new_n923_), .B(_abc_4635_new_n754__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_5927_13_));
AND2X2 AND2X2_351 ( .A(_abc_4635_new_n511__bF_buf2), .B(\Rdata_mem[14] ), .Y(_abc_4635_new_n925_));
AND2X2 AND2X2_352 ( .A(_abc_4635_new_n859_), .B(_abc_4635_new_n480__bF_buf4), .Y(_abc_4635_new_n926_));
AND2X2 AND2X2_353 ( .A(_abc_4635_new_n928_), .B(_abc_4635_new_n754__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_5927_14_));
AND2X2 AND2X2_354 ( .A(_abc_4635_new_n511__bF_buf1), .B(\Rdata_mem[15] ), .Y(_abc_4635_new_n930_));
AND2X2 AND2X2_355 ( .A(_abc_4635_new_n932_), .B(_abc_4635_new_n480__bF_buf3), .Y(_abc_4635_new_n933_));
AND2X2 AND2X2_356 ( .A(_abc_4635_new_n933_), .B(_abc_4635_new_n931_), .Y(_abc_4635_new_n934_));
AND2X2 AND2X2_357 ( .A(_abc_4635_new_n936_), .B(_abc_4635_new_n754__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_5927_15_));
AND2X2 AND2X2_358 ( .A(_abc_4635_new_n511__bF_buf0), .B(\Rdata_mem[16] ), .Y(_abc_4635_new_n938_));
AND2X2 AND2X2_359 ( .A(_abc_4635_new_n934_), .B(signo), .Y(_abc_4635_new_n939_));
AND2X2 AND2X2_36 ( .A(AWready), .B(state_4_), .Y(_abc_4635_new_n421_));
AND2X2 AND2X2_360 ( .A(_abc_4635_new_n941_), .B(_abc_4635_new_n754__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_5927_16_));
AND2X2 AND2X2_361 ( .A(_abc_4635_new_n511__bF_buf6), .B(\Rdata_mem[17] ), .Y(_abc_4635_new_n943_));
AND2X2 AND2X2_362 ( .A(_abc_4635_new_n944_), .B(_abc_4635_new_n754__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_5927_17_));
AND2X2 AND2X2_363 ( .A(_abc_4635_new_n511__bF_buf5), .B(\Rdata_mem[18] ), .Y(_abc_4635_new_n946_));
AND2X2 AND2X2_364 ( .A(_abc_4635_new_n947_), .B(_abc_4635_new_n754__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_5927_18_));
AND2X2 AND2X2_365 ( .A(_abc_4635_new_n511__bF_buf4), .B(\Rdata_mem[19] ), .Y(_abc_4635_new_n949_));
AND2X2 AND2X2_366 ( .A(_abc_4635_new_n950_), .B(_abc_4635_new_n754__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_5927_19_));
AND2X2 AND2X2_367 ( .A(_abc_4635_new_n511__bF_buf3), .B(\Rdata_mem[20] ), .Y(_abc_4635_new_n952_));
AND2X2 AND2X2_368 ( .A(_abc_4635_new_n953_), .B(_abc_4635_new_n754__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_5927_20_));
AND2X2 AND2X2_369 ( .A(_abc_4635_new_n511__bF_buf2), .B(\Rdata_mem[21] ), .Y(_abc_4635_new_n955_));
AND2X2 AND2X2_37 ( .A(_abc_4635_new_n422_), .B(_abc_4635_new_n420_), .Y(_abc_4635_new_n423_));
AND2X2 AND2X2_370 ( .A(_abc_4635_new_n956_), .B(_abc_4635_new_n754__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_5927_21_));
AND2X2 AND2X2_371 ( .A(_abc_4635_new_n511__bF_buf1), .B(\Rdata_mem[22] ), .Y(_abc_4635_new_n958_));
AND2X2 AND2X2_372 ( .A(_abc_4635_new_n959_), .B(_abc_4635_new_n754__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_5927_22_));
AND2X2 AND2X2_373 ( .A(_abc_4635_new_n511__bF_buf0), .B(\Rdata_mem[23] ), .Y(_abc_4635_new_n961_));
AND2X2 AND2X2_374 ( .A(_abc_4635_new_n962_), .B(_abc_4635_new_n754__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_5927_23_));
AND2X2 AND2X2_375 ( .A(_abc_4635_new_n511__bF_buf6), .B(\Rdata_mem[24] ), .Y(_abc_4635_new_n964_));
AND2X2 AND2X2_376 ( .A(_abc_4635_new_n965_), .B(_abc_4635_new_n754__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_5927_24_));
AND2X2 AND2X2_377 ( .A(_abc_4635_new_n511__bF_buf5), .B(\Rdata_mem[25] ), .Y(_abc_4635_new_n967_));
AND2X2 AND2X2_378 ( .A(_abc_4635_new_n968_), .B(_abc_4635_new_n754__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_5927_25_));
AND2X2 AND2X2_379 ( .A(_abc_4635_new_n511__bF_buf4), .B(\Rdata_mem[26] ), .Y(_abc_4635_new_n970_));
AND2X2 AND2X2_38 ( .A(_abc_4635_new_n425_), .B(resetn_bF_buf4), .Y(_abc_4635_new_n426_));
AND2X2 AND2X2_380 ( .A(_abc_4635_new_n971_), .B(_abc_4635_new_n754__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_5927_26_));
AND2X2 AND2X2_381 ( .A(_abc_4635_new_n511__bF_buf3), .B(\Rdata_mem[27] ), .Y(_abc_4635_new_n973_));
AND2X2 AND2X2_382 ( .A(_abc_4635_new_n974_), .B(_abc_4635_new_n754__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_5927_27_));
AND2X2 AND2X2_383 ( .A(_abc_4635_new_n511__bF_buf2), .B(\Rdata_mem[28] ), .Y(_abc_4635_new_n976_));
AND2X2 AND2X2_384 ( .A(_abc_4635_new_n977_), .B(_abc_4635_new_n754__bF_buf1), .Y(_auto_iopadmap_cc_368_execute_5927_28_));
AND2X2 AND2X2_385 ( .A(_abc_4635_new_n511__bF_buf1), .B(\Rdata_mem[29] ), .Y(_abc_4635_new_n979_));
AND2X2 AND2X2_386 ( .A(_abc_4635_new_n980_), .B(_abc_4635_new_n754__bF_buf0), .Y(_auto_iopadmap_cc_368_execute_5927_29_));
AND2X2 AND2X2_387 ( .A(_abc_4635_new_n511__bF_buf0), .B(\Rdata_mem[30] ), .Y(_abc_4635_new_n982_));
AND2X2 AND2X2_388 ( .A(_abc_4635_new_n983_), .B(_abc_4635_new_n754__bF_buf4), .Y(_auto_iopadmap_cc_368_execute_5927_30_));
AND2X2 AND2X2_389 ( .A(_abc_4635_new_n511__bF_buf6), .B(\Rdata_mem[31] ), .Y(_abc_4635_new_n985_));
AND2X2 AND2X2_39 ( .A(_abc_4635_new_n426_), .B(_abc_4635_new_n374_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_4_));
AND2X2 AND2X2_390 ( .A(_abc_4635_new_n986_), .B(_abc_4635_new_n754__bF_buf3), .Y(_auto_iopadmap_cc_368_execute_5927_31_));
AND2X2 AND2X2_391 ( .A(_abc_4635_new_n988_), .B(_abc_4635_new_n989_), .Y(_auto_iopadmap_cc_368_execute_5767_0_));
AND2X2 AND2X2_392 ( .A(_abc_4635_new_n991_), .B(_abc_4635_new_n992_), .Y(_auto_iopadmap_cc_368_execute_5767_1_));
AND2X2 AND2X2_393 ( .A(\imm[2] ), .B(\rs1[2] ), .Y(_abc_4635_new_n995_));
AND2X2 AND2X2_394 ( .A(_abc_4635_new_n996_), .B(_abc_4635_new_n997_), .Y(_abc_4635_new_n998_));
AND2X2 AND2X2_395 ( .A(_abc_4635_new_n994_), .B(_abc_4635_new_n998_), .Y(_abc_4635_new_n999_));
AND2X2 AND2X2_396 ( .A(_abc_4635_new_n1000_), .B(_abc_4635_new_n1001_), .Y(_abc_4635_new_n1002_));
AND2X2 AND2X2_397 ( .A(_abc_4635_new_n1003_), .B(_abc_4635_new_n1004_), .Y(_auto_iopadmap_cc_368_execute_5767_2_));
AND2X2 AND2X2_398 ( .A(_abc_4635_new_n1000_), .B(_abc_4635_new_n996_), .Y(_abc_4635_new_n1006_));
AND2X2 AND2X2_399 ( .A(\imm[3] ), .B(\rs1[3] ), .Y(_abc_4635_new_n1008_));
AND2X2 AND2X2_4 ( .A(AWready), .B(Wready), .Y(_abc_4635_new_n367_));
AND2X2 AND2X2_40 ( .A(resetn_bF_buf3), .B(state_5_), .Y(_abc_4635_new_n429_));
AND2X2 AND2X2_400 ( .A(_abc_4635_new_n1009_), .B(_abc_4635_new_n1007_), .Y(_abc_4635_new_n1010_));
AND2X2 AND2X2_401 ( .A(_abc_4635_new_n1014_), .B(_abc_4635_new_n1012_), .Y(_abc_4635_new_n1015_));
AND2X2 AND2X2_402 ( .A(_abc_4635_new_n1016_), .B(_abc_4635_new_n1017_), .Y(_auto_iopadmap_cc_368_execute_5767_3_));
AND2X2 AND2X2_403 ( .A(_abc_4635_new_n998_), .B(_abc_4635_new_n1010_), .Y(_abc_4635_new_n1019_));
AND2X2 AND2X2_404 ( .A(_abc_4635_new_n994_), .B(_abc_4635_new_n1019_), .Y(_abc_4635_new_n1020_));
AND2X2 AND2X2_405 ( .A(_abc_4635_new_n1007_), .B(_abc_4635_new_n995_), .Y(_abc_4635_new_n1021_));
AND2X2 AND2X2_406 ( .A(\imm[4] ), .B(\rs1[4] ), .Y(_abc_4635_new_n1025_));
AND2X2 AND2X2_407 ( .A(_abc_4635_new_n1026_), .B(_abc_4635_new_n1024_), .Y(_abc_4635_new_n1027_));
AND2X2 AND2X2_408 ( .A(_abc_4635_new_n1023_), .B(_abc_4635_new_n1027_), .Y(_abc_4635_new_n1028_));
AND2X2 AND2X2_409 ( .A(_abc_4635_new_n1029_), .B(_abc_4635_new_n1030_), .Y(_abc_4635_new_n1031_));
AND2X2 AND2X2_41 ( .A(_abc_4635_new_n395_), .B(ARready), .Y(_abc_4635_new_n430_));
AND2X2 AND2X2_410 ( .A(_abc_4635_new_n1032_), .B(_abc_4635_new_n1033_), .Y(_auto_iopadmap_cc_368_execute_5767_4_));
AND2X2 AND2X2_411 ( .A(_abc_4635_new_n1029_), .B(_abc_4635_new_n1026_), .Y(_abc_4635_new_n1035_));
AND2X2 AND2X2_412 ( .A(\imm[5] ), .B(\rs1[5] ), .Y(_abc_4635_new_n1038_));
AND2X2 AND2X2_413 ( .A(_abc_4635_new_n1039_), .B(_abc_4635_new_n1037_), .Y(_abc_4635_new_n1040_));
AND2X2 AND2X2_414 ( .A(_abc_4635_new_n1041_), .B(_abc_4635_new_n1043_), .Y(_abc_4635_new_n1044_));
AND2X2 AND2X2_415 ( .A(_abc_4635_new_n1045_), .B(_abc_4635_new_n1046_), .Y(_auto_iopadmap_cc_368_execute_5767_5_));
AND2X2 AND2X2_416 ( .A(W_R_1_bF_buf1_), .B(\pc[6] ), .Y(_abc_4635_new_n1048_));
AND2X2 AND2X2_417 ( .A(_abc_4635_new_n1049_), .B(_abc_4635_new_n1037_), .Y(_abc_4635_new_n1050_));
AND2X2 AND2X2_418 ( .A(_abc_4635_new_n1027_), .B(_abc_4635_new_n1040_), .Y(_abc_4635_new_n1051_));
AND2X2 AND2X2_419 ( .A(_abc_4635_new_n1023_), .B(_abc_4635_new_n1051_), .Y(_abc_4635_new_n1052_));
AND2X2 AND2X2_42 ( .A(_abc_4635_new_n431_), .B(_abc_4635_new_n428_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_5_));
AND2X2 AND2X2_420 ( .A(\imm[6] ), .B(\rs1[6] ), .Y(_abc_4635_new_n1054_));
AND2X2 AND2X2_421 ( .A(_abc_4635_new_n1055_), .B(_abc_4635_new_n1056_), .Y(_abc_4635_new_n1057_));
AND2X2 AND2X2_422 ( .A(_abc_4635_new_n1053_), .B(_abc_4635_new_n1057_), .Y(_abc_4635_new_n1059_));
AND2X2 AND2X2_423 ( .A(_abc_4635_new_n1060_), .B(_abc_4635_new_n1058_), .Y(_abc_4635_new_n1061_));
AND2X2 AND2X2_424 ( .A(_abc_4635_new_n1061_), .B(_abc_4635_new_n753__bF_buf2), .Y(_abc_4635_new_n1062_));
AND2X2 AND2X2_425 ( .A(_abc_4635_new_n1060_), .B(_abc_4635_new_n1055_), .Y(_abc_4635_new_n1065_));
AND2X2 AND2X2_426 ( .A(\imm[7] ), .B(\rs1[7] ), .Y(_abc_4635_new_n1067_));
AND2X2 AND2X2_427 ( .A(_abc_4635_new_n1068_), .B(_abc_4635_new_n1066_), .Y(_abc_4635_new_n1069_));
AND2X2 AND2X2_428 ( .A(_abc_4635_new_n1073_), .B(_abc_4635_new_n1071_), .Y(_abc_4635_new_n1074_));
AND2X2 AND2X2_429 ( .A(_abc_4635_new_n1075_), .B(_abc_4635_new_n1064_), .Y(_auto_iopadmap_cc_368_execute_5767_7_));
AND2X2 AND2X2_43 ( .A(_abc_4635_new_n377_), .B(_abc_4635_new_n390_), .Y(_abc_4635_new_n434_));
AND2X2 AND2X2_430 ( .A(W_R_1_bF_buf5_), .B(\pc[8] ), .Y(_abc_4635_new_n1077_));
AND2X2 AND2X2_431 ( .A(_abc_4635_new_n1057_), .B(_abc_4635_new_n1069_), .Y(_abc_4635_new_n1078_));
AND2X2 AND2X2_432 ( .A(_abc_4635_new_n1051_), .B(_abc_4635_new_n1078_), .Y(_abc_4635_new_n1079_));
AND2X2 AND2X2_433 ( .A(_abc_4635_new_n1023_), .B(_abc_4635_new_n1079_), .Y(_abc_4635_new_n1080_));
AND2X2 AND2X2_434 ( .A(_abc_4635_new_n1078_), .B(_abc_4635_new_n1050_), .Y(_abc_4635_new_n1081_));
AND2X2 AND2X2_435 ( .A(_abc_4635_new_n1066_), .B(_abc_4635_new_n1054_), .Y(_abc_4635_new_n1082_));
AND2X2 AND2X2_436 ( .A(\imm[8] ), .B(\rs1[8] ), .Y(_abc_4635_new_n1086_));
AND2X2 AND2X2_437 ( .A(_abc_4635_new_n1087_), .B(_abc_4635_new_n1088_), .Y(_abc_4635_new_n1089_));
AND2X2 AND2X2_438 ( .A(_abc_4635_new_n1085_), .B(_abc_4635_new_n1089_), .Y(_abc_4635_new_n1091_));
AND2X2 AND2X2_439 ( .A(_abc_4635_new_n1092_), .B(_abc_4635_new_n1090_), .Y(_abc_4635_new_n1093_));
AND2X2 AND2X2_44 ( .A(_abc_4635_new_n428_), .B(state_5_), .Y(_abc_4635_new_n440_));
AND2X2 AND2X2_440 ( .A(_abc_4635_new_n1093_), .B(_abc_4635_new_n753__bF_buf0), .Y(_abc_4635_new_n1094_));
AND2X2 AND2X2_441 ( .A(_abc_4635_new_n1092_), .B(_abc_4635_new_n1087_), .Y(_abc_4635_new_n1096_));
AND2X2 AND2X2_442 ( .A(\imm[9] ), .B(\rs1[9] ), .Y(_abc_4635_new_n1099_));
AND2X2 AND2X2_443 ( .A(_abc_4635_new_n1100_), .B(_abc_4635_new_n1098_), .Y(_abc_4635_new_n1101_));
AND2X2 AND2X2_444 ( .A(_abc_4635_new_n1102_), .B(_abc_4635_new_n1104_), .Y(_abc_4635_new_n1105_));
AND2X2 AND2X2_445 ( .A(_abc_4635_new_n1106_), .B(_abc_4635_new_n1107_), .Y(_auto_iopadmap_cc_368_execute_5767_9_));
AND2X2 AND2X2_446 ( .A(W_R_1_bF_buf3_), .B(\pc[10] ), .Y(_abc_4635_new_n1109_));
AND2X2 AND2X2_447 ( .A(_abc_4635_new_n1110_), .B(_abc_4635_new_n1098_), .Y(_abc_4635_new_n1111_));
AND2X2 AND2X2_448 ( .A(_abc_4635_new_n1089_), .B(_abc_4635_new_n1101_), .Y(_abc_4635_new_n1112_));
AND2X2 AND2X2_449 ( .A(_abc_4635_new_n1085_), .B(_abc_4635_new_n1112_), .Y(_abc_4635_new_n1113_));
AND2X2 AND2X2_45 ( .A(_abc_4635_new_n441_), .B(_abc_4635_new_n443_), .Y(_abc_4635_new_n444_));
AND2X2 AND2X2_450 ( .A(\imm[10] ), .B(\rs1[10] ), .Y(_abc_4635_new_n1115_));
AND2X2 AND2X2_451 ( .A(_abc_4635_new_n1116_), .B(_abc_4635_new_n1117_), .Y(_abc_4635_new_n1118_));
AND2X2 AND2X2_452 ( .A(_abc_4635_new_n1114_), .B(_abc_4635_new_n1118_), .Y(_abc_4635_new_n1120_));
AND2X2 AND2X2_453 ( .A(_abc_4635_new_n1121_), .B(_abc_4635_new_n1119_), .Y(_abc_4635_new_n1122_));
AND2X2 AND2X2_454 ( .A(_abc_4635_new_n1122_), .B(_abc_4635_new_n753__bF_buf3), .Y(_abc_4635_new_n1123_));
AND2X2 AND2X2_455 ( .A(_abc_4635_new_n1121_), .B(_abc_4635_new_n1116_), .Y(_abc_4635_new_n1125_));
AND2X2 AND2X2_456 ( .A(\imm[11] ), .B(\rs1[11] ), .Y(_abc_4635_new_n1128_));
AND2X2 AND2X2_457 ( .A(_abc_4635_new_n1129_), .B(_abc_4635_new_n1127_), .Y(_abc_4635_new_n1130_));
AND2X2 AND2X2_458 ( .A(_abc_4635_new_n1126_), .B(_abc_4635_new_n1131_), .Y(_abc_4635_new_n1132_));
AND2X2 AND2X2_459 ( .A(_abc_4635_new_n1125_), .B(_abc_4635_new_n1130_), .Y(_abc_4635_new_n1133_));
AND2X2 AND2X2_46 ( .A(_abc_4635_new_n439_), .B(_abc_4635_new_n444_), .Y(_abc_4635_new_n445_));
AND2X2 AND2X2_460 ( .A(_abc_4635_new_n1134_), .B(_abc_4635_new_n753__bF_buf2), .Y(_abc_4635_new_n1135_));
AND2X2 AND2X2_461 ( .A(W_R_1_bF_buf2_), .B(\pc[11] ), .Y(_abc_4635_new_n1136_));
AND2X2 AND2X2_462 ( .A(W_R_1_bF_buf1_), .B(\pc[12] ), .Y(_abc_4635_new_n1138_));
AND2X2 AND2X2_463 ( .A(_abc_4635_new_n1118_), .B(_abc_4635_new_n1130_), .Y(_abc_4635_new_n1139_));
AND2X2 AND2X2_464 ( .A(_abc_4635_new_n1139_), .B(_abc_4635_new_n1111_), .Y(_abc_4635_new_n1140_));
AND2X2 AND2X2_465 ( .A(_abc_4635_new_n1127_), .B(_abc_4635_new_n1115_), .Y(_abc_4635_new_n1141_));
AND2X2 AND2X2_466 ( .A(_abc_4635_new_n1112_), .B(_abc_4635_new_n1139_), .Y(_abc_4635_new_n1144_));
AND2X2 AND2X2_467 ( .A(_abc_4635_new_n1085_), .B(_abc_4635_new_n1144_), .Y(_abc_4635_new_n1145_));
AND2X2 AND2X2_468 ( .A(\imm[12] ), .B(\rs1[12] ), .Y(_abc_4635_new_n1148_));
AND2X2 AND2X2_469 ( .A(_abc_4635_new_n1149_), .B(_abc_4635_new_n1147_), .Y(_abc_4635_new_n1150_));
AND2X2 AND2X2_47 ( .A(Bvalid), .B(Wready), .Y(_abc_4635_new_n447_));
AND2X2 AND2X2_470 ( .A(_abc_4635_new_n1146_), .B(_abc_4635_new_n1150_), .Y(_abc_4635_new_n1152_));
AND2X2 AND2X2_471 ( .A(_abc_4635_new_n1153_), .B(_abc_4635_new_n1151_), .Y(_abc_4635_new_n1154_));
AND2X2 AND2X2_472 ( .A(_abc_4635_new_n1154_), .B(_abc_4635_new_n753__bF_buf1), .Y(_abc_4635_new_n1155_));
AND2X2 AND2X2_473 ( .A(_abc_4635_new_n1153_), .B(_abc_4635_new_n1149_), .Y(_abc_4635_new_n1157_));
AND2X2 AND2X2_474 ( .A(\imm[13] ), .B(\rs1[13] ), .Y(_abc_4635_new_n1159_));
AND2X2 AND2X2_475 ( .A(_abc_4635_new_n1160_), .B(_abc_4635_new_n1158_), .Y(_abc_4635_new_n1161_));
AND2X2 AND2X2_476 ( .A(_abc_4635_new_n1157_), .B(_abc_4635_new_n1161_), .Y(_abc_4635_new_n1162_));
AND2X2 AND2X2_477 ( .A(_abc_4635_new_n1163_), .B(_abc_4635_new_n1164_), .Y(_abc_4635_new_n1165_));
AND2X2 AND2X2_478 ( .A(_abc_4635_new_n1166_), .B(_abc_4635_new_n753__bF_buf0), .Y(_abc_4635_new_n1167_));
AND2X2 AND2X2_479 ( .A(W_R_1_bF_buf0_), .B(\pc[13] ), .Y(_abc_4635_new_n1168_));
AND2X2 AND2X2_48 ( .A(_abc_4635_new_n448_), .B(_abc_4635_new_n450_), .Y(_abc_4635_new_n451_));
AND2X2 AND2X2_480 ( .A(W_R_1_bF_buf5_), .B(\pc[14] ), .Y(_abc_4635_new_n1170_));
AND2X2 AND2X2_481 ( .A(_abc_4635_new_n1171_), .B(_abc_4635_new_n1160_), .Y(_abc_4635_new_n1172_));
AND2X2 AND2X2_482 ( .A(_abc_4635_new_n1150_), .B(_abc_4635_new_n1161_), .Y(_abc_4635_new_n1174_));
AND2X2 AND2X2_483 ( .A(_abc_4635_new_n1146_), .B(_abc_4635_new_n1174_), .Y(_abc_4635_new_n1175_));
AND2X2 AND2X2_484 ( .A(\imm[14] ), .B(\rs1[14] ), .Y(_abc_4635_new_n1177_));
AND2X2 AND2X2_485 ( .A(_abc_4635_new_n1178_), .B(_abc_4635_new_n1179_), .Y(_abc_4635_new_n1180_));
AND2X2 AND2X2_486 ( .A(_abc_4635_new_n1176_), .B(_abc_4635_new_n1180_), .Y(_abc_4635_new_n1182_));
AND2X2 AND2X2_487 ( .A(_abc_4635_new_n1183_), .B(_abc_4635_new_n1181_), .Y(_abc_4635_new_n1184_));
AND2X2 AND2X2_488 ( .A(_abc_4635_new_n1184_), .B(_abc_4635_new_n753__bF_buf4), .Y(_abc_4635_new_n1185_));
AND2X2 AND2X2_489 ( .A(_abc_4635_new_n1183_), .B(_abc_4635_new_n1178_), .Y(_abc_4635_new_n1188_));
AND2X2 AND2X2_49 ( .A(_abc_4635_new_n445_), .B(_abc_4635_new_n451_), .Y(_abc_4635_new_n452_));
AND2X2 AND2X2_490 ( .A(\imm[15] ), .B(\rs1[15] ), .Y(_abc_4635_new_n1190_));
AND2X2 AND2X2_491 ( .A(_abc_4635_new_n1191_), .B(_abc_4635_new_n1189_), .Y(_abc_4635_new_n1192_));
AND2X2 AND2X2_492 ( .A(_abc_4635_new_n1196_), .B(_abc_4635_new_n1194_), .Y(_abc_4635_new_n1197_));
AND2X2 AND2X2_493 ( .A(_abc_4635_new_n1198_), .B(_abc_4635_new_n1187_), .Y(_auto_iopadmap_cc_368_execute_5767_15_));
AND2X2 AND2X2_494 ( .A(W_R_1_bF_buf3_), .B(\pc[16] ), .Y(_abc_4635_new_n1200_));
AND2X2 AND2X2_495 ( .A(_abc_4635_new_n1180_), .B(_abc_4635_new_n1192_), .Y(_abc_4635_new_n1201_));
AND2X2 AND2X2_496 ( .A(_abc_4635_new_n1174_), .B(_abc_4635_new_n1201_), .Y(_abc_4635_new_n1202_));
AND2X2 AND2X2_497 ( .A(_abc_4635_new_n1144_), .B(_abc_4635_new_n1202_), .Y(_abc_4635_new_n1203_));
AND2X2 AND2X2_498 ( .A(_abc_4635_new_n1085_), .B(_abc_4635_new_n1203_), .Y(_abc_4635_new_n1204_));
AND2X2 AND2X2_499 ( .A(_abc_4635_new_n1143_), .B(_abc_4635_new_n1202_), .Y(_abc_4635_new_n1205_));
AND2X2 AND2X2_5 ( .A(_abc_4635_new_n368_), .B(AWready), .Y(_abc_4635_new_n369_));
AND2X2 AND2X2_50 ( .A(_abc_4635_new_n452_), .B(_abc_4635_new_n438_), .Y(_abc_4635_new_n453_));
AND2X2 AND2X2_500 ( .A(_abc_4635_new_n1189_), .B(_abc_4635_new_n1177_), .Y(_abc_4635_new_n1206_));
AND2X2 AND2X2_501 ( .A(_abc_4635_new_n1173_), .B(_abc_4635_new_n1201_), .Y(_abc_4635_new_n1208_));
AND2X2 AND2X2_502 ( .A(\imm[16] ), .B(\rs1[16] ), .Y(_abc_4635_new_n1213_));
AND2X2 AND2X2_503 ( .A(_abc_4635_new_n1214_), .B(_abc_4635_new_n1212_), .Y(_abc_4635_new_n1215_));
AND2X2 AND2X2_504 ( .A(_abc_4635_new_n1211_), .B(_abc_4635_new_n1215_), .Y(_abc_4635_new_n1217_));
AND2X2 AND2X2_505 ( .A(_abc_4635_new_n1218_), .B(_abc_4635_new_n1216_), .Y(_abc_4635_new_n1219_));
AND2X2 AND2X2_506 ( .A(_abc_4635_new_n1219_), .B(_abc_4635_new_n753__bF_buf2), .Y(_abc_4635_new_n1220_));
AND2X2 AND2X2_507 ( .A(_abc_4635_new_n1218_), .B(_abc_4635_new_n1214_), .Y(_abc_4635_new_n1222_));
AND2X2 AND2X2_508 ( .A(\imm[17] ), .B(\rs1[17] ), .Y(_abc_4635_new_n1224_));
AND2X2 AND2X2_509 ( .A(_abc_4635_new_n1225_), .B(_abc_4635_new_n1226_), .Y(_abc_4635_new_n1227_));
AND2X2 AND2X2_51 ( .A(_abc_4635_new_n453_), .B(_abc_4635_new_n436_), .Y(_abc_4635_new_n454_));
AND2X2 AND2X2_510 ( .A(_abc_4635_new_n1228_), .B(_abc_4635_new_n1230_), .Y(_abc_4635_new_n1231_));
AND2X2 AND2X2_511 ( .A(_abc_4635_new_n1232_), .B(_abc_4635_new_n1233_), .Y(_auto_iopadmap_cc_368_execute_5767_17_));
AND2X2 AND2X2_512 ( .A(W_R_1_bF_buf1_), .B(\pc[18] ), .Y(_abc_4635_new_n1235_));
AND2X2 AND2X2_513 ( .A(_abc_4635_new_n1236_), .B(_abc_4635_new_n1225_), .Y(_abc_4635_new_n1237_));
AND2X2 AND2X2_514 ( .A(_abc_4635_new_n1215_), .B(_abc_4635_new_n1227_), .Y(_abc_4635_new_n1239_));
AND2X2 AND2X2_515 ( .A(_abc_4635_new_n1211_), .B(_abc_4635_new_n1239_), .Y(_abc_4635_new_n1240_));
AND2X2 AND2X2_516 ( .A(\imm[18] ), .B(\rs1[18] ), .Y(_abc_4635_new_n1242_));
AND2X2 AND2X2_517 ( .A(_abc_4635_new_n1243_), .B(_abc_4635_new_n1244_), .Y(_abc_4635_new_n1245_));
AND2X2 AND2X2_518 ( .A(_abc_4635_new_n1241_), .B(_abc_4635_new_n1245_), .Y(_abc_4635_new_n1247_));
AND2X2 AND2X2_519 ( .A(_abc_4635_new_n1248_), .B(_abc_4635_new_n1246_), .Y(_abc_4635_new_n1249_));
AND2X2 AND2X2_52 ( .A(_abc_4635_new_n457_), .B(_abc_4635_new_n458_), .Y(_abc_4635_new_n459_));
AND2X2 AND2X2_520 ( .A(_abc_4635_new_n1249_), .B(_abc_4635_new_n753__bF_buf0), .Y(_abc_4635_new_n1250_));
AND2X2 AND2X2_521 ( .A(_abc_4635_new_n1248_), .B(_abc_4635_new_n1243_), .Y(_abc_4635_new_n1253_));
AND2X2 AND2X2_522 ( .A(\imm[19] ), .B(\rs1[19] ), .Y(_abc_4635_new_n1254_));
AND2X2 AND2X2_523 ( .A(_abc_4635_new_n1255_), .B(_abc_4635_new_n1256_), .Y(_abc_4635_new_n1257_));
AND2X2 AND2X2_524 ( .A(_abc_4635_new_n1261_), .B(_abc_4635_new_n1259_), .Y(_abc_4635_new_n1262_));
AND2X2 AND2X2_525 ( .A(_abc_4635_new_n1263_), .B(_abc_4635_new_n1252_), .Y(_auto_iopadmap_cc_368_execute_5767_19_));
AND2X2 AND2X2_526 ( .A(W_R_1_bF_buf5_), .B(\pc[20] ), .Y(_abc_4635_new_n1265_));
AND2X2 AND2X2_527 ( .A(_abc_4635_new_n1245_), .B(_abc_4635_new_n1257_), .Y(_abc_4635_new_n1266_));
AND2X2 AND2X2_528 ( .A(_abc_4635_new_n1238_), .B(_abc_4635_new_n1266_), .Y(_abc_4635_new_n1267_));
AND2X2 AND2X2_529 ( .A(_abc_4635_new_n1256_), .B(_abc_4635_new_n1242_), .Y(_abc_4635_new_n1268_));
AND2X2 AND2X2_53 ( .A(\imm[0] ), .B(\rs1[0] ), .Y(_abc_4635_new_n460_));
AND2X2 AND2X2_530 ( .A(_abc_4635_new_n1239_), .B(_abc_4635_new_n1266_), .Y(_abc_4635_new_n1271_));
AND2X2 AND2X2_531 ( .A(_abc_4635_new_n1211_), .B(_abc_4635_new_n1271_), .Y(_abc_4635_new_n1272_));
AND2X2 AND2X2_532 ( .A(\imm[20] ), .B(\rs1[20] ), .Y(_abc_4635_new_n1274_));
AND2X2 AND2X2_533 ( .A(_abc_4635_new_n1275_), .B(_abc_4635_new_n1276_), .Y(_abc_4635_new_n1277_));
AND2X2 AND2X2_534 ( .A(_abc_4635_new_n1273_), .B(_abc_4635_new_n1277_), .Y(_abc_4635_new_n1279_));
AND2X2 AND2X2_535 ( .A(_abc_4635_new_n1280_), .B(_abc_4635_new_n1278_), .Y(_abc_4635_new_n1281_));
AND2X2 AND2X2_536 ( .A(_abc_4635_new_n1281_), .B(_abc_4635_new_n753__bF_buf3), .Y(_abc_4635_new_n1282_));
AND2X2 AND2X2_537 ( .A(_abc_4635_new_n1280_), .B(_abc_4635_new_n1275_), .Y(_abc_4635_new_n1284_));
AND2X2 AND2X2_538 ( .A(\imm[21] ), .B(\rs1[21] ), .Y(_abc_4635_new_n1286_));
AND2X2 AND2X2_539 ( .A(_abc_4635_new_n1287_), .B(_abc_4635_new_n1288_), .Y(_abc_4635_new_n1289_));
AND2X2 AND2X2_54 ( .A(\imm[1] ), .B(\rs1[1] ), .Y(_abc_4635_new_n462_));
AND2X2 AND2X2_540 ( .A(_abc_4635_new_n1290_), .B(_abc_4635_new_n1292_), .Y(_abc_4635_new_n1293_));
AND2X2 AND2X2_541 ( .A(_abc_4635_new_n1294_), .B(_abc_4635_new_n1295_), .Y(_auto_iopadmap_cc_368_execute_5767_21_));
AND2X2 AND2X2_542 ( .A(W_R_1_bF_buf3_), .B(\pc[22] ), .Y(_abc_4635_new_n1297_));
AND2X2 AND2X2_543 ( .A(_abc_4635_new_n1298_), .B(_abc_4635_new_n1287_), .Y(_abc_4635_new_n1299_));
AND2X2 AND2X2_544 ( .A(_abc_4635_new_n1277_), .B(_abc_4635_new_n1289_), .Y(_abc_4635_new_n1301_));
AND2X2 AND2X2_545 ( .A(_abc_4635_new_n1273_), .B(_abc_4635_new_n1301_), .Y(_abc_4635_new_n1302_));
AND2X2 AND2X2_546 ( .A(\imm[22] ), .B(\rs1[22] ), .Y(_abc_4635_new_n1304_));
AND2X2 AND2X2_547 ( .A(_abc_4635_new_n1305_), .B(_abc_4635_new_n1306_), .Y(_abc_4635_new_n1307_));
AND2X2 AND2X2_548 ( .A(_abc_4635_new_n1303_), .B(_abc_4635_new_n1307_), .Y(_abc_4635_new_n1309_));
AND2X2 AND2X2_549 ( .A(_abc_4635_new_n1310_), .B(_abc_4635_new_n1308_), .Y(_abc_4635_new_n1311_));
AND2X2 AND2X2_55 ( .A(_abc_4635_new_n463_), .B(_abc_4635_new_n461_), .Y(_abc_4635_new_n464_));
AND2X2 AND2X2_550 ( .A(_abc_4635_new_n1311_), .B(_abc_4635_new_n753__bF_buf1), .Y(_abc_4635_new_n1312_));
AND2X2 AND2X2_551 ( .A(_abc_4635_new_n1310_), .B(_abc_4635_new_n1305_), .Y(_abc_4635_new_n1315_));
AND2X2 AND2X2_552 ( .A(\imm[23] ), .B(\rs1[23] ), .Y(_abc_4635_new_n1316_));
AND2X2 AND2X2_553 ( .A(_abc_4635_new_n1317_), .B(_abc_4635_new_n1318_), .Y(_abc_4635_new_n1319_));
AND2X2 AND2X2_554 ( .A(_abc_4635_new_n1323_), .B(_abc_4635_new_n1321_), .Y(_abc_4635_new_n1324_));
AND2X2 AND2X2_555 ( .A(_abc_4635_new_n1325_), .B(_abc_4635_new_n1314_), .Y(_auto_iopadmap_cc_368_execute_5767_23_));
AND2X2 AND2X2_556 ( .A(W_R_1_bF_buf1_), .B(\pc[24] ), .Y(_abc_4635_new_n1327_));
AND2X2 AND2X2_557 ( .A(_abc_4635_new_n1307_), .B(_abc_4635_new_n1319_), .Y(_abc_4635_new_n1328_));
AND2X2 AND2X2_558 ( .A(_abc_4635_new_n1301_), .B(_abc_4635_new_n1328_), .Y(_abc_4635_new_n1329_));
AND2X2 AND2X2_559 ( .A(_abc_4635_new_n1271_), .B(_abc_4635_new_n1329_), .Y(_abc_4635_new_n1330_));
AND2X2 AND2X2_56 ( .A(_abc_4635_new_n464_), .B(_abc_4635_new_n460_), .Y(_abc_4635_new_n465_));
AND2X2 AND2X2_560 ( .A(_abc_4635_new_n1211_), .B(_abc_4635_new_n1330_), .Y(_abc_4635_new_n1331_));
AND2X2 AND2X2_561 ( .A(_abc_4635_new_n1270_), .B(_abc_4635_new_n1329_), .Y(_abc_4635_new_n1332_));
AND2X2 AND2X2_562 ( .A(_abc_4635_new_n1300_), .B(_abc_4635_new_n1328_), .Y(_abc_4635_new_n1333_));
AND2X2 AND2X2_563 ( .A(_abc_4635_new_n1318_), .B(_abc_4635_new_n1304_), .Y(_abc_4635_new_n1334_));
AND2X2 AND2X2_564 ( .A(\imm[24] ), .B(\rs1[24] ), .Y(_abc_4635_new_n1339_));
AND2X2 AND2X2_565 ( .A(_abc_4635_new_n1340_), .B(_abc_4635_new_n1341_), .Y(_abc_4635_new_n1342_));
AND2X2 AND2X2_566 ( .A(_abc_4635_new_n1338_), .B(_abc_4635_new_n1342_), .Y(_abc_4635_new_n1344_));
AND2X2 AND2X2_567 ( .A(_abc_4635_new_n1345_), .B(_abc_4635_new_n1343_), .Y(_abc_4635_new_n1346_));
AND2X2 AND2X2_568 ( .A(_abc_4635_new_n1346_), .B(_abc_4635_new_n753__bF_buf4), .Y(_abc_4635_new_n1347_));
AND2X2 AND2X2_569 ( .A(_abc_4635_new_n1345_), .B(_abc_4635_new_n1340_), .Y(_abc_4635_new_n1349_));
AND2X2 AND2X2_57 ( .A(_abc_4635_new_n467_), .B(_abc_4635_new_n468_), .Y(_abc_4635_new_n469_));
AND2X2 AND2X2_570 ( .A(\imm[25] ), .B(\rs1[25] ), .Y(_abc_4635_new_n1351_));
AND2X2 AND2X2_571 ( .A(_abc_4635_new_n1352_), .B(_abc_4635_new_n1353_), .Y(_abc_4635_new_n1354_));
AND2X2 AND2X2_572 ( .A(_abc_4635_new_n1355_), .B(_abc_4635_new_n1357_), .Y(_abc_4635_new_n1358_));
AND2X2 AND2X2_573 ( .A(_abc_4635_new_n1359_), .B(_abc_4635_new_n1360_), .Y(_auto_iopadmap_cc_368_execute_5767_25_));
AND2X2 AND2X2_574 ( .A(W_R_1_bF_buf5_), .B(\pc[26] ), .Y(_abc_4635_new_n1362_));
AND2X2 AND2X2_575 ( .A(_abc_4635_new_n1363_), .B(_abc_4635_new_n1352_), .Y(_abc_4635_new_n1364_));
AND2X2 AND2X2_576 ( .A(_abc_4635_new_n1342_), .B(_abc_4635_new_n1354_), .Y(_abc_4635_new_n1366_));
AND2X2 AND2X2_577 ( .A(_abc_4635_new_n1338_), .B(_abc_4635_new_n1366_), .Y(_abc_4635_new_n1367_));
AND2X2 AND2X2_578 ( .A(\imm[26] ), .B(\rs1[26] ), .Y(_abc_4635_new_n1369_));
AND2X2 AND2X2_579 ( .A(_abc_4635_new_n1370_), .B(_abc_4635_new_n1371_), .Y(_abc_4635_new_n1372_));
AND2X2 AND2X2_58 ( .A(_abc_4635_new_n470_), .B(_abc_4635_new_n466_), .Y(_abc_4635_new_n471_));
AND2X2 AND2X2_580 ( .A(_abc_4635_new_n1368_), .B(_abc_4635_new_n1372_), .Y(_abc_4635_new_n1374_));
AND2X2 AND2X2_581 ( .A(_abc_4635_new_n1375_), .B(_abc_4635_new_n1373_), .Y(_abc_4635_new_n1376_));
AND2X2 AND2X2_582 ( .A(_abc_4635_new_n1376_), .B(_abc_4635_new_n753__bF_buf2), .Y(_abc_4635_new_n1377_));
AND2X2 AND2X2_583 ( .A(_abc_4635_new_n1375_), .B(_abc_4635_new_n1370_), .Y(_abc_4635_new_n1380_));
AND2X2 AND2X2_584 ( .A(\imm[27] ), .B(\rs1[27] ), .Y(_abc_4635_new_n1382_));
AND2X2 AND2X2_585 ( .A(_abc_4635_new_n1383_), .B(_abc_4635_new_n1381_), .Y(_abc_4635_new_n1384_));
AND2X2 AND2X2_586 ( .A(_abc_4635_new_n1388_), .B(_abc_4635_new_n1386_), .Y(_abc_4635_new_n1389_));
AND2X2 AND2X2_587 ( .A(_abc_4635_new_n1390_), .B(_abc_4635_new_n1379_), .Y(_auto_iopadmap_cc_368_execute_5767_27_));
AND2X2 AND2X2_588 ( .A(W_R_1_bF_buf3_), .B(\pc[28] ), .Y(_abc_4635_new_n1392_));
AND2X2 AND2X2_589 ( .A(_abc_4635_new_n1372_), .B(_abc_4635_new_n1384_), .Y(_abc_4635_new_n1393_));
AND2X2 AND2X2_59 ( .A(_abc_4635_new_n466_), .B(_abc_4635_new_n473_), .Y(_abc_4635_new_n474_));
AND2X2 AND2X2_590 ( .A(_abc_4635_new_n1366_), .B(_abc_4635_new_n1393_), .Y(_abc_4635_new_n1394_));
AND2X2 AND2X2_591 ( .A(_abc_4635_new_n1338_), .B(_abc_4635_new_n1394_), .Y(_abc_4635_new_n1395_));
AND2X2 AND2X2_592 ( .A(_abc_4635_new_n1365_), .B(_abc_4635_new_n1393_), .Y(_abc_4635_new_n1396_));
AND2X2 AND2X2_593 ( .A(_abc_4635_new_n1381_), .B(_abc_4635_new_n1369_), .Y(_abc_4635_new_n1397_));
AND2X2 AND2X2_594 ( .A(\imm[28] ), .B(\rs1[28] ), .Y(_abc_4635_new_n1402_));
AND2X2 AND2X2_595 ( .A(_abc_4635_new_n1403_), .B(_abc_4635_new_n1401_), .Y(_abc_4635_new_n1404_));
AND2X2 AND2X2_596 ( .A(_abc_4635_new_n1400_), .B(_abc_4635_new_n1404_), .Y(_abc_4635_new_n1406_));
AND2X2 AND2X2_597 ( .A(_abc_4635_new_n1407_), .B(_abc_4635_new_n1405_), .Y(_abc_4635_new_n1408_));
AND2X2 AND2X2_598 ( .A(_abc_4635_new_n1408_), .B(_abc_4635_new_n753__bF_buf0), .Y(_abc_4635_new_n1409_));
AND2X2 AND2X2_599 ( .A(_abc_4635_new_n1407_), .B(_abc_4635_new_n1403_), .Y(_abc_4635_new_n1411_));
AND2X2 AND2X2_6 ( .A(resetn_bF_buf4), .B(state_4_), .Y(_abc_4635_new_n371_));
AND2X2 AND2X2_60 ( .A(_abc_4635_new_n472__bF_buf3), .B(_abc_4635_new_n475_), .Y(_abc_4635_new_n476_));
AND2X2 AND2X2_600 ( .A(\imm[29] ), .B(\rs1[29] ), .Y(_abc_4635_new_n1414_));
AND2X2 AND2X2_601 ( .A(_abc_4635_new_n1415_), .B(_abc_4635_new_n1413_), .Y(_abc_4635_new_n1416_));
AND2X2 AND2X2_602 ( .A(_abc_4635_new_n1417_), .B(_abc_4635_new_n1419_), .Y(_abc_4635_new_n1420_));
AND2X2 AND2X2_603 ( .A(_abc_4635_new_n1421_), .B(_abc_4635_new_n1422_), .Y(_auto_iopadmap_cc_368_execute_5767_29_));
AND2X2 AND2X2_604 ( .A(W_R_1_bF_buf1_), .B(\pc[30] ), .Y(_abc_4635_new_n1424_));
AND2X2 AND2X2_605 ( .A(_abc_4635_new_n1404_), .B(_abc_4635_new_n1416_), .Y(_abc_4635_new_n1425_));
AND2X2 AND2X2_606 ( .A(_abc_4635_new_n1400_), .B(_abc_4635_new_n1425_), .Y(_abc_4635_new_n1426_));
AND2X2 AND2X2_607 ( .A(_abc_4635_new_n1413_), .B(_abc_4635_new_n1402_), .Y(_abc_4635_new_n1427_));
AND2X2 AND2X2_608 ( .A(\imm[30] ), .B(\rs1[30] ), .Y(_abc_4635_new_n1431_));
AND2X2 AND2X2_609 ( .A(_abc_4635_new_n1432_), .B(_abc_4635_new_n1430_), .Y(_abc_4635_new_n1433_));
AND2X2 AND2X2_61 ( .A(_abc_4635_new_n477_), .B(_abc_4635_new_n459_), .Y(_abc_4635_new_n478_));
AND2X2 AND2X2_610 ( .A(_abc_4635_new_n1435_), .B(_abc_4635_new_n463_), .Y(_abc_4635_new_n1436_));
AND2X2 AND2X2_611 ( .A(_abc_4635_new_n1438_), .B(_abc_4635_new_n1439_), .Y(_abc_4635_new_n1440_));
AND2X2 AND2X2_612 ( .A(_abc_4635_new_n1442_), .B(_abc_4635_new_n1443_), .Y(_abc_4635_new_n1444_));
AND2X2 AND2X2_613 ( .A(_abc_4635_new_n1446_), .B(_abc_4635_new_n1447_), .Y(_abc_4635_new_n1448_));
AND2X2 AND2X2_614 ( .A(_abc_4635_new_n1450_), .B(_abc_4635_new_n1451_), .Y(_abc_4635_new_n1452_));
AND2X2 AND2X2_615 ( .A(_abc_4635_new_n1454_), .B(_abc_4635_new_n1455_), .Y(_abc_4635_new_n1456_));
AND2X2 AND2X2_616 ( .A(_abc_4635_new_n1458_), .B(_abc_4635_new_n1459_), .Y(_abc_4635_new_n1460_));
AND2X2 AND2X2_617 ( .A(_abc_4635_new_n1462_), .B(_abc_4635_new_n1434_), .Y(_abc_4635_new_n1463_));
AND2X2 AND2X2_618 ( .A(_abc_4635_new_n1463_), .B(_abc_4635_new_n753__bF_buf3), .Y(_abc_4635_new_n1464_));
AND2X2 AND2X2_619 ( .A(_abc_4635_new_n1429_), .B(_abc_4635_new_n1433_), .Y(_abc_4635_new_n1466_));
AND2X2 AND2X2_62 ( .A(_abc_4635_new_n458_), .B(\wordsize[0] ), .Y(_abc_4635_new_n480_));
AND2X2 AND2X2_620 ( .A(_abc_4635_new_n1469_), .B(_abc_4635_new_n1471_), .Y(_abc_4635_new_n1472_));
AND2X2 AND2X2_621 ( .A(_abc_4635_new_n1462_), .B(_abc_4635_new_n1432_), .Y(_abc_4635_new_n1475_));
AND2X2 AND2X2_622 ( .A(_abc_4635_new_n1476_), .B(_abc_4635_new_n1474_), .Y(_abc_4635_new_n1477_));
AND2X2 AND2X2_623 ( .A(_abc_4635_new_n1478_), .B(_abc_4635_new_n1479_), .Y(_auto_iopadmap_cc_368_execute_5767_31_));
AND2X2 AND2X2_624 ( .A(_abc_4635_new_n615_), .B(_abc_4635_new_n754__bF_buf2), .Y(_auto_iopadmap_cc_368_execute_5960));
AND2X2 AND2X2_625 ( .A(_abc_4635_new_n1484_), .B(resetn_bF_buf4), .Y(_auto_iopadmap_cc_368_execute_5837));
AND2X2 AND2X2_626 ( .A(_abc_4635_new_n1486_), .B(resetn_bF_buf3), .Y(_auto_iopadmap_cc_368_execute_5800));
AND2X2 AND2X2_627 ( .A(_abc_4635_new_n1483_), .B(resetn_bF_buf2), .Y(_auto_iopadmap_cc_368_execute_5879));
AND2X2 AND2X2_63 ( .A(\wordsize[0] ), .B(\wordsize[1] ), .Y(_abc_4635_new_n483_));
AND2X2 AND2X2_64 ( .A(_abc_4635_new_n380_), .B(resetn_bF_buf2), .Y(_abc_4635_new_n485_));
AND2X2 AND2X2_65 ( .A(_abc_4635_new_n485__bF_buf4), .B(_abc_4635_new_n484_), .Y(_abc_4635_new_n486_));
AND2X2 AND2X2_66 ( .A(_abc_4635_new_n482_), .B(_abc_4635_new_n486_), .Y(_abc_4635_new_n487_));
AND2X2 AND2X2_67 ( .A(_abc_4635_new_n479_), .B(_abc_4635_new_n487_), .Y(_0Wstrb_3_0__0_));
AND2X2 AND2X2_68 ( .A(_abc_4635_new_n472__bF_buf1), .B(_abc_4635_new_n489_), .Y(_abc_4635_new_n490_));
AND2X2 AND2X2_69 ( .A(_abc_4635_new_n491_), .B(_abc_4635_new_n486_), .Y(_0Wstrb_3_0__1_));
AND2X2 AND2X2_7 ( .A(_abc_4635_new_n370_), .B(_abc_4635_new_n371_), .Y(_abc_4635_new_n372_));
AND2X2 AND2X2_70 ( .A(_abc_4635_new_n493__bF_buf3), .B(_abc_4635_new_n494_), .Y(_abc_4635_new_n495_));
AND2X2 AND2X2_71 ( .A(_abc_4635_new_n496_), .B(_abc_4635_new_n486_), .Y(_0Wstrb_3_0__2_));
AND2X2 AND2X2_72 ( .A(_abc_4635_new_n493__bF_buf2), .B(_abc_4635_new_n489_), .Y(_abc_4635_new_n498_));
AND2X2 AND2X2_73 ( .A(_abc_4635_new_n499_), .B(_abc_4635_new_n486_), .Y(_0Wstrb_3_0__3_));
AND2X2 AND2X2_74 ( .A(_abc_4635_new_n486_), .B(\rs2[0] ), .Y(_0Wdata_31_0__0_));
AND2X2 AND2X2_75 ( .A(_abc_4635_new_n486_), .B(\rs2[1] ), .Y(_0Wdata_31_0__1_));
AND2X2 AND2X2_76 ( .A(_abc_4635_new_n486_), .B(\rs2[2] ), .Y(_0Wdata_31_0__2_));
AND2X2 AND2X2_77 ( .A(_abc_4635_new_n486_), .B(\rs2[3] ), .Y(_0Wdata_31_0__3_));
AND2X2 AND2X2_78 ( .A(_abc_4635_new_n486_), .B(\rs2[4] ), .Y(_0Wdata_31_0__4_));
AND2X2 AND2X2_79 ( .A(_abc_4635_new_n486_), .B(\rs2[5] ), .Y(_0Wdata_31_0__5_));
AND2X2 AND2X2_8 ( .A(_abc_4635_new_n373_), .B(_abc_4635_new_n368_), .Y(_abc_4635_new_n374_));
AND2X2 AND2X2_80 ( .A(_abc_4635_new_n486_), .B(\rs2[6] ), .Y(_0Wdata_31_0__6_));
AND2X2 AND2X2_81 ( .A(_abc_4635_new_n486_), .B(\rs2[7] ), .Y(_0Wdata_31_0__7_));
AND2X2 AND2X2_82 ( .A(_abc_4635_new_n458_), .B(\rs2[0] ), .Y(_abc_4635_new_n509_));
AND2X2 AND2X2_83 ( .A(_abc_4635_new_n509_), .B(_abc_4635_new_n457_), .Y(_abc_4635_new_n510_));
AND2X2 AND2X2_84 ( .A(_abc_4635_new_n457_), .B(\wordsize[1] ), .Y(_abc_4635_new_n511_));
AND2X2 AND2X2_85 ( .A(_abc_4635_new_n512_), .B(\rs2[8] ), .Y(_abc_4635_new_n513_));
AND2X2 AND2X2_86 ( .A(_abc_4635_new_n514_), .B(_abc_4635_new_n485__bF_buf3), .Y(_0Wdata_31_0__8_));
AND2X2 AND2X2_87 ( .A(_abc_4635_new_n458_), .B(\rs2[1] ), .Y(_abc_4635_new_n516_));
AND2X2 AND2X2_88 ( .A(_abc_4635_new_n516_), .B(_abc_4635_new_n457_), .Y(_abc_4635_new_n517_));
AND2X2 AND2X2_89 ( .A(_abc_4635_new_n512_), .B(\rs2[9] ), .Y(_abc_4635_new_n518_));
AND2X2 AND2X2_9 ( .A(_abc_4635_new_n376_), .B(enable), .Y(_abc_4635_new_n377_));
AND2X2 AND2X2_90 ( .A(_abc_4635_new_n519_), .B(_abc_4635_new_n485__bF_buf2), .Y(_0Wdata_31_0__9_));
AND2X2 AND2X2_91 ( .A(_abc_4635_new_n458_), .B(\rs2[2] ), .Y(_abc_4635_new_n521_));
AND2X2 AND2X2_92 ( .A(_abc_4635_new_n521_), .B(_abc_4635_new_n457_), .Y(_abc_4635_new_n522_));
AND2X2 AND2X2_93 ( .A(_abc_4635_new_n512_), .B(\rs2[10] ), .Y(_abc_4635_new_n523_));
AND2X2 AND2X2_94 ( .A(_abc_4635_new_n524_), .B(_abc_4635_new_n485__bF_buf1), .Y(_0Wdata_31_0__10_));
AND2X2 AND2X2_95 ( .A(_abc_4635_new_n458_), .B(\rs2[3] ), .Y(_abc_4635_new_n526_));
AND2X2 AND2X2_96 ( .A(_abc_4635_new_n526_), .B(_abc_4635_new_n457_), .Y(_abc_4635_new_n527_));
AND2X2 AND2X2_97 ( .A(_abc_4635_new_n512_), .B(\rs2[11] ), .Y(_abc_4635_new_n528_));
AND2X2 AND2X2_98 ( .A(_abc_4635_new_n529_), .B(_abc_4635_new_n485__bF_buf0), .Y(_0Wdata_31_0__11_));
AND2X2 AND2X2_99 ( .A(_abc_4635_new_n458_), .B(\rs2[4] ), .Y(_abc_4635_new_n531_));
BUFX2 BUFX2_1 ( .A(_abc_4635_new_n485_), .Y(_abc_4635_new_n485__bF_buf4));
BUFX2 BUFX2_10 ( .A(_auto_iopadmap_cc_368_execute_5767_0_), .Y(\ARdata[0] ));
BUFX2 BUFX2_100 ( .A(_auto_iopadmap_cc_368_execute_5841_22_), .Y(\Wdata[22] ));
BUFX2 BUFX2_101 ( .A(_auto_iopadmap_cc_368_execute_5841_23_), .Y(\Wdata[23] ));
BUFX2 BUFX2_102 ( .A(_auto_iopadmap_cc_368_execute_5841_24_), .Y(\Wdata[24] ));
BUFX2 BUFX2_103 ( .A(_auto_iopadmap_cc_368_execute_5841_25_), .Y(\Wdata[25] ));
BUFX2 BUFX2_104 ( .A(_auto_iopadmap_cc_368_execute_5841_26_), .Y(\Wdata[26] ));
BUFX2 BUFX2_105 ( .A(_auto_iopadmap_cc_368_execute_5841_27_), .Y(\Wdata[27] ));
BUFX2 BUFX2_106 ( .A(_auto_iopadmap_cc_368_execute_5841_28_), .Y(\Wdata[28] ));
BUFX2 BUFX2_107 ( .A(_auto_iopadmap_cc_368_execute_5841_29_), .Y(\Wdata[29] ));
BUFX2 BUFX2_108 ( .A(_auto_iopadmap_cc_368_execute_5841_30_), .Y(\Wdata[30] ));
BUFX2 BUFX2_109 ( .A(_auto_iopadmap_cc_368_execute_5841_31_), .Y(\Wdata[31] ));
BUFX2 BUFX2_11 ( .A(_auto_iopadmap_cc_368_execute_5767_1_), .Y(\ARdata[1] ));
BUFX2 BUFX2_110 ( .A(_auto_iopadmap_cc_368_execute_5874_0_), .Y(\Wstrb[0] ));
BUFX2 BUFX2_111 ( .A(_auto_iopadmap_cc_368_execute_5874_1_), .Y(\Wstrb[1] ));
BUFX2 BUFX2_112 ( .A(_auto_iopadmap_cc_368_execute_5874_2_), .Y(\Wstrb[2] ));
BUFX2 BUFX2_113 ( .A(_auto_iopadmap_cc_368_execute_5874_3_), .Y(\Wstrb[3] ));
BUFX2 BUFX2_114 ( .A(_auto_iopadmap_cc_368_execute_5879), .Y(Wvalid));
BUFX2 BUFX2_115 ( .A(_auto_iopadmap_cc_368_execute_5881), .Y(align));
BUFX2 BUFX2_116 ( .A(1'h0), .Y(\arprot[0] ));
BUFX2 BUFX2_117 ( .A(1'h0), .Y(\arprot[1] ));
BUFX2 BUFX2_118 ( .A(1'h0), .Y(\awprot[0] ));
BUFX2 BUFX2_119 ( .A(1'h0), .Y(\awprot[1] ));
BUFX2 BUFX2_12 ( .A(_auto_iopadmap_cc_368_execute_5767_2_), .Y(\ARdata[2] ));
BUFX2 BUFX2_120 ( .A(1'h0), .Y(\awprot[2] ));
BUFX2 BUFX2_121 ( .A(_auto_iopadmap_cc_368_execute_5890), .Y(busy));
BUFX2 BUFX2_122 ( .A(_auto_iopadmap_cc_368_execute_5892), .Y(done));
BUFX2 BUFX2_123 ( .A(_auto_iopadmap_cc_368_execute_5894_0_), .Y(\inst[0] ));
BUFX2 BUFX2_124 ( .A(_auto_iopadmap_cc_368_execute_5894_1_), .Y(\inst[1] ));
BUFX2 BUFX2_125 ( .A(_auto_iopadmap_cc_368_execute_5894_2_), .Y(\inst[2] ));
BUFX2 BUFX2_126 ( .A(_auto_iopadmap_cc_368_execute_5894_3_), .Y(\inst[3] ));
BUFX2 BUFX2_127 ( .A(_auto_iopadmap_cc_368_execute_5894_4_), .Y(\inst[4] ));
BUFX2 BUFX2_128 ( .A(_auto_iopadmap_cc_368_execute_5894_5_), .Y(\inst[5] ));
BUFX2 BUFX2_129 ( .A(_auto_iopadmap_cc_368_execute_5894_6_), .Y(\inst[6] ));
BUFX2 BUFX2_13 ( .A(_auto_iopadmap_cc_368_execute_5767_3_), .Y(\ARdata[3] ));
BUFX2 BUFX2_130 ( .A(_auto_iopadmap_cc_368_execute_5894_7_), .Y(\inst[7] ));
BUFX2 BUFX2_131 ( .A(_auto_iopadmap_cc_368_execute_5894_8_), .Y(\inst[8] ));
BUFX2 BUFX2_132 ( .A(_auto_iopadmap_cc_368_execute_5894_9_), .Y(\inst[9] ));
BUFX2 BUFX2_133 ( .A(_auto_iopadmap_cc_368_execute_5894_10_), .Y(\inst[10] ));
BUFX2 BUFX2_134 ( .A(_auto_iopadmap_cc_368_execute_5894_11_), .Y(\inst[11] ));
BUFX2 BUFX2_135 ( .A(_auto_iopadmap_cc_368_execute_5894_12_), .Y(\inst[12] ));
BUFX2 BUFX2_136 ( .A(_auto_iopadmap_cc_368_execute_5894_13_), .Y(\inst[13] ));
BUFX2 BUFX2_137 ( .A(_auto_iopadmap_cc_368_execute_5894_14_), .Y(\inst[14] ));
BUFX2 BUFX2_138 ( .A(_auto_iopadmap_cc_368_execute_5894_15_), .Y(\inst[15] ));
BUFX2 BUFX2_139 ( .A(_auto_iopadmap_cc_368_execute_5894_16_), .Y(\inst[16] ));
BUFX2 BUFX2_14 ( .A(_auto_iopadmap_cc_368_execute_5767_4_), .Y(\ARdata[4] ));
BUFX2 BUFX2_140 ( .A(_auto_iopadmap_cc_368_execute_5894_17_), .Y(\inst[17] ));
BUFX2 BUFX2_141 ( .A(_auto_iopadmap_cc_368_execute_5894_18_), .Y(\inst[18] ));
BUFX2 BUFX2_142 ( .A(_auto_iopadmap_cc_368_execute_5894_19_), .Y(\inst[19] ));
BUFX2 BUFX2_143 ( .A(_auto_iopadmap_cc_368_execute_5894_20_), .Y(\inst[20] ));
BUFX2 BUFX2_144 ( .A(_auto_iopadmap_cc_368_execute_5894_21_), .Y(\inst[21] ));
BUFX2 BUFX2_145 ( .A(_auto_iopadmap_cc_368_execute_5894_22_), .Y(\inst[22] ));
BUFX2 BUFX2_146 ( .A(_auto_iopadmap_cc_368_execute_5894_23_), .Y(\inst[23] ));
BUFX2 BUFX2_147 ( .A(_auto_iopadmap_cc_368_execute_5894_24_), .Y(\inst[24] ));
BUFX2 BUFX2_148 ( .A(_auto_iopadmap_cc_368_execute_5894_25_), .Y(\inst[25] ));
BUFX2 BUFX2_149 ( .A(_auto_iopadmap_cc_368_execute_5894_26_), .Y(\inst[26] ));
BUFX2 BUFX2_15 ( .A(_auto_iopadmap_cc_368_execute_5767_5_), .Y(\ARdata[5] ));
BUFX2 BUFX2_150 ( .A(_auto_iopadmap_cc_368_execute_5894_27_), .Y(\inst[27] ));
BUFX2 BUFX2_151 ( .A(_auto_iopadmap_cc_368_execute_5894_28_), .Y(\inst[28] ));
BUFX2 BUFX2_152 ( .A(_auto_iopadmap_cc_368_execute_5894_29_), .Y(\inst[29] ));
BUFX2 BUFX2_153 ( .A(_auto_iopadmap_cc_368_execute_5894_30_), .Y(\inst[30] ));
BUFX2 BUFX2_154 ( .A(_auto_iopadmap_cc_368_execute_5894_31_), .Y(\inst[31] ));
BUFX2 BUFX2_155 ( .A(_auto_iopadmap_cc_368_execute_5927_0_), .Y(\rd[0] ));
BUFX2 BUFX2_156 ( .A(_auto_iopadmap_cc_368_execute_5927_1_), .Y(\rd[1] ));
BUFX2 BUFX2_157 ( .A(_auto_iopadmap_cc_368_execute_5927_2_), .Y(\rd[2] ));
BUFX2 BUFX2_158 ( .A(_auto_iopadmap_cc_368_execute_5927_3_), .Y(\rd[3] ));
BUFX2 BUFX2_159 ( .A(_auto_iopadmap_cc_368_execute_5927_4_), .Y(\rd[4] ));
BUFX2 BUFX2_16 ( .A(_auto_iopadmap_cc_368_execute_5767_6_), .Y(\ARdata[6] ));
BUFX2 BUFX2_160 ( .A(_auto_iopadmap_cc_368_execute_5927_5_), .Y(\rd[5] ));
BUFX2 BUFX2_161 ( .A(_auto_iopadmap_cc_368_execute_5927_6_), .Y(\rd[6] ));
BUFX2 BUFX2_162 ( .A(_auto_iopadmap_cc_368_execute_5927_7_), .Y(\rd[7] ));
BUFX2 BUFX2_163 ( .A(_auto_iopadmap_cc_368_execute_5927_8_), .Y(\rd[8] ));
BUFX2 BUFX2_164 ( .A(_auto_iopadmap_cc_368_execute_5927_9_), .Y(\rd[9] ));
BUFX2 BUFX2_165 ( .A(_auto_iopadmap_cc_368_execute_5927_10_), .Y(\rd[10] ));
BUFX2 BUFX2_166 ( .A(_auto_iopadmap_cc_368_execute_5927_11_), .Y(\rd[11] ));
BUFX2 BUFX2_167 ( .A(_auto_iopadmap_cc_368_execute_5927_12_), .Y(\rd[12] ));
BUFX2 BUFX2_168 ( .A(_auto_iopadmap_cc_368_execute_5927_13_), .Y(\rd[13] ));
BUFX2 BUFX2_169 ( .A(_auto_iopadmap_cc_368_execute_5927_14_), .Y(\rd[14] ));
BUFX2 BUFX2_17 ( .A(_auto_iopadmap_cc_368_execute_5767_7_), .Y(\ARdata[7] ));
BUFX2 BUFX2_170 ( .A(_auto_iopadmap_cc_368_execute_5927_15_), .Y(\rd[15] ));
BUFX2 BUFX2_171 ( .A(_auto_iopadmap_cc_368_execute_5927_16_), .Y(\rd[16] ));
BUFX2 BUFX2_172 ( .A(_auto_iopadmap_cc_368_execute_5927_17_), .Y(\rd[17] ));
BUFX2 BUFX2_173 ( .A(_auto_iopadmap_cc_368_execute_5927_18_), .Y(\rd[18] ));
BUFX2 BUFX2_174 ( .A(_auto_iopadmap_cc_368_execute_5927_19_), .Y(\rd[19] ));
BUFX2 BUFX2_175 ( .A(_auto_iopadmap_cc_368_execute_5927_20_), .Y(\rd[20] ));
BUFX2 BUFX2_176 ( .A(_auto_iopadmap_cc_368_execute_5927_21_), .Y(\rd[21] ));
BUFX2 BUFX2_177 ( .A(_auto_iopadmap_cc_368_execute_5927_22_), .Y(\rd[22] ));
BUFX2 BUFX2_178 ( .A(_auto_iopadmap_cc_368_execute_5927_23_), .Y(\rd[23] ));
BUFX2 BUFX2_179 ( .A(_auto_iopadmap_cc_368_execute_5927_24_), .Y(\rd[24] ));
BUFX2 BUFX2_18 ( .A(_auto_iopadmap_cc_368_execute_5767_8_), .Y(\ARdata[8] ));
BUFX2 BUFX2_180 ( .A(_auto_iopadmap_cc_368_execute_5927_25_), .Y(\rd[25] ));
BUFX2 BUFX2_181 ( .A(_auto_iopadmap_cc_368_execute_5927_26_), .Y(\rd[26] ));
BUFX2 BUFX2_182 ( .A(_auto_iopadmap_cc_368_execute_5927_27_), .Y(\rd[27] ));
BUFX2 BUFX2_183 ( .A(_auto_iopadmap_cc_368_execute_5927_28_), .Y(\rd[28] ));
BUFX2 BUFX2_184 ( .A(_auto_iopadmap_cc_368_execute_5927_29_), .Y(\rd[29] ));
BUFX2 BUFX2_185 ( .A(_auto_iopadmap_cc_368_execute_5927_30_), .Y(\rd[30] ));
BUFX2 BUFX2_186 ( .A(_auto_iopadmap_cc_368_execute_5927_31_), .Y(\rd[31] ));
BUFX2 BUFX2_187 ( .A(_auto_iopadmap_cc_368_execute_5960), .Y(rd_en));
BUFX2 BUFX2_188 ( .A(en_instr), .Y(\arprot[2] ));
BUFX2 BUFX2_19 ( .A(_auto_iopadmap_cc_368_execute_5767_9_), .Y(\ARdata[9] ));
BUFX2 BUFX2_2 ( .A(_abc_4635_new_n485_), .Y(_abc_4635_new_n485__bF_buf3));
BUFX2 BUFX2_20 ( .A(_auto_iopadmap_cc_368_execute_5767_10_), .Y(\ARdata[10] ));
BUFX2 BUFX2_21 ( .A(_auto_iopadmap_cc_368_execute_5767_11_), .Y(\ARdata[11] ));
BUFX2 BUFX2_22 ( .A(_auto_iopadmap_cc_368_execute_5767_12_), .Y(\ARdata[12] ));
BUFX2 BUFX2_23 ( .A(_auto_iopadmap_cc_368_execute_5767_13_), .Y(\ARdata[13] ));
BUFX2 BUFX2_24 ( .A(_auto_iopadmap_cc_368_execute_5767_14_), .Y(\ARdata[14] ));
BUFX2 BUFX2_25 ( .A(_auto_iopadmap_cc_368_execute_5767_15_), .Y(\ARdata[15] ));
BUFX2 BUFX2_26 ( .A(_auto_iopadmap_cc_368_execute_5767_16_), .Y(\ARdata[16] ));
BUFX2 BUFX2_27 ( .A(_auto_iopadmap_cc_368_execute_5767_17_), .Y(\ARdata[17] ));
BUFX2 BUFX2_28 ( .A(_auto_iopadmap_cc_368_execute_5767_18_), .Y(\ARdata[18] ));
BUFX2 BUFX2_29 ( .A(_auto_iopadmap_cc_368_execute_5767_19_), .Y(\ARdata[19] ));
BUFX2 BUFX2_3 ( .A(_abc_4635_new_n485_), .Y(_abc_4635_new_n485__bF_buf2));
BUFX2 BUFX2_30 ( .A(_auto_iopadmap_cc_368_execute_5767_20_), .Y(\ARdata[20] ));
BUFX2 BUFX2_31 ( .A(_auto_iopadmap_cc_368_execute_5767_21_), .Y(\ARdata[21] ));
BUFX2 BUFX2_32 ( .A(_auto_iopadmap_cc_368_execute_5767_22_), .Y(\ARdata[22] ));
BUFX2 BUFX2_33 ( .A(_auto_iopadmap_cc_368_execute_5767_23_), .Y(\ARdata[23] ));
BUFX2 BUFX2_34 ( .A(_auto_iopadmap_cc_368_execute_5767_24_), .Y(\ARdata[24] ));
BUFX2 BUFX2_35 ( .A(_auto_iopadmap_cc_368_execute_5767_25_), .Y(\ARdata[25] ));
BUFX2 BUFX2_36 ( .A(_auto_iopadmap_cc_368_execute_5767_26_), .Y(\ARdata[26] ));
BUFX2 BUFX2_37 ( .A(_auto_iopadmap_cc_368_execute_5767_27_), .Y(\ARdata[27] ));
BUFX2 BUFX2_38 ( .A(_auto_iopadmap_cc_368_execute_5767_28_), .Y(\ARdata[28] ));
BUFX2 BUFX2_39 ( .A(_auto_iopadmap_cc_368_execute_5767_29_), .Y(\ARdata[29] ));
BUFX2 BUFX2_4 ( .A(_abc_4635_new_n485_), .Y(_abc_4635_new_n485__bF_buf1));
BUFX2 BUFX2_40 ( .A(_auto_iopadmap_cc_368_execute_5767_30_), .Y(\ARdata[30] ));
BUFX2 BUFX2_41 ( .A(_auto_iopadmap_cc_368_execute_5767_31_), .Y(\ARdata[31] ));
BUFX2 BUFX2_42 ( .A(_auto_iopadmap_cc_368_execute_5800), .Y(ARvalid));
BUFX2 BUFX2_43 ( .A(_auto_iopadmap_cc_368_execute_5767_0_), .Y(\AWdata[0] ));
BUFX2 BUFX2_44 ( .A(_auto_iopadmap_cc_368_execute_5767_1_), .Y(\AWdata[1] ));
BUFX2 BUFX2_45 ( .A(_auto_iopadmap_cc_368_execute_5767_2_), .Y(\AWdata[2] ));
BUFX2 BUFX2_46 ( .A(_auto_iopadmap_cc_368_execute_5767_3_), .Y(\AWdata[3] ));
BUFX2 BUFX2_47 ( .A(_auto_iopadmap_cc_368_execute_5767_4_), .Y(\AWdata[4] ));
BUFX2 BUFX2_48 ( .A(_auto_iopadmap_cc_368_execute_5767_5_), .Y(\AWdata[5] ));
BUFX2 BUFX2_49 ( .A(_auto_iopadmap_cc_368_execute_5767_6_), .Y(\AWdata[6] ));
BUFX2 BUFX2_5 ( .A(_abc_4635_new_n485_), .Y(_abc_4635_new_n485__bF_buf0));
BUFX2 BUFX2_50 ( .A(_auto_iopadmap_cc_368_execute_5767_7_), .Y(\AWdata[7] ));
BUFX2 BUFX2_51 ( .A(_auto_iopadmap_cc_368_execute_5767_8_), .Y(\AWdata[8] ));
BUFX2 BUFX2_52 ( .A(_auto_iopadmap_cc_368_execute_5767_9_), .Y(\AWdata[9] ));
BUFX2 BUFX2_53 ( .A(_auto_iopadmap_cc_368_execute_5767_10_), .Y(\AWdata[10] ));
BUFX2 BUFX2_54 ( .A(_auto_iopadmap_cc_368_execute_5767_11_), .Y(\AWdata[11] ));
BUFX2 BUFX2_55 ( .A(_auto_iopadmap_cc_368_execute_5767_12_), .Y(\AWdata[12] ));
BUFX2 BUFX2_56 ( .A(_auto_iopadmap_cc_368_execute_5767_13_), .Y(\AWdata[13] ));
BUFX2 BUFX2_57 ( .A(_auto_iopadmap_cc_368_execute_5767_14_), .Y(\AWdata[14] ));
BUFX2 BUFX2_58 ( .A(_auto_iopadmap_cc_368_execute_5767_15_), .Y(\AWdata[15] ));
BUFX2 BUFX2_59 ( .A(_auto_iopadmap_cc_368_execute_5767_16_), .Y(\AWdata[16] ));
BUFX2 BUFX2_6 ( .A(_abc_4635_new_n480_), .Y(_abc_4635_new_n480__bF_buf2));
BUFX2 BUFX2_60 ( .A(_auto_iopadmap_cc_368_execute_5767_17_), .Y(\AWdata[17] ));
BUFX2 BUFX2_61 ( .A(_auto_iopadmap_cc_368_execute_5767_18_), .Y(\AWdata[18] ));
BUFX2 BUFX2_62 ( .A(_auto_iopadmap_cc_368_execute_5767_19_), .Y(\AWdata[19] ));
BUFX2 BUFX2_63 ( .A(_auto_iopadmap_cc_368_execute_5767_20_), .Y(\AWdata[20] ));
BUFX2 BUFX2_64 ( .A(_auto_iopadmap_cc_368_execute_5767_21_), .Y(\AWdata[21] ));
BUFX2 BUFX2_65 ( .A(_auto_iopadmap_cc_368_execute_5767_22_), .Y(\AWdata[22] ));
BUFX2 BUFX2_66 ( .A(_auto_iopadmap_cc_368_execute_5767_23_), .Y(\AWdata[23] ));
BUFX2 BUFX2_67 ( .A(_auto_iopadmap_cc_368_execute_5767_24_), .Y(\AWdata[24] ));
BUFX2 BUFX2_68 ( .A(_auto_iopadmap_cc_368_execute_5767_25_), .Y(\AWdata[25] ));
BUFX2 BUFX2_69 ( .A(_auto_iopadmap_cc_368_execute_5767_26_), .Y(\AWdata[26] ));
BUFX2 BUFX2_7 ( .A(_abc_4635_new_n480_), .Y(_abc_4635_new_n480__bF_buf1));
BUFX2 BUFX2_70 ( .A(_auto_iopadmap_cc_368_execute_5767_27_), .Y(\AWdata[27] ));
BUFX2 BUFX2_71 ( .A(_auto_iopadmap_cc_368_execute_5767_28_), .Y(\AWdata[28] ));
BUFX2 BUFX2_72 ( .A(_auto_iopadmap_cc_368_execute_5767_29_), .Y(\AWdata[29] ));
BUFX2 BUFX2_73 ( .A(_auto_iopadmap_cc_368_execute_5767_30_), .Y(\AWdata[30] ));
BUFX2 BUFX2_74 ( .A(_auto_iopadmap_cc_368_execute_5767_31_), .Y(\AWdata[31] ));
BUFX2 BUFX2_75 ( .A(_auto_iopadmap_cc_368_execute_5835), .Y(AWvalid));
BUFX2 BUFX2_76 ( .A(_auto_iopadmap_cc_368_execute_5837), .Y(Bready));
BUFX2 BUFX2_77 ( .A(_auto_iopadmap_cc_368_execute_5839), .Y(RReady));
BUFX2 BUFX2_78 ( .A(_auto_iopadmap_cc_368_execute_5841_0_), .Y(\Wdata[0] ));
BUFX2 BUFX2_79 ( .A(_auto_iopadmap_cc_368_execute_5841_1_), .Y(\Wdata[1] ));
BUFX2 BUFX2_8 ( .A(_abc_4635_new_n480_), .Y(_abc_4635_new_n480__bF_buf0));
BUFX2 BUFX2_80 ( .A(_auto_iopadmap_cc_368_execute_5841_2_), .Y(\Wdata[2] ));
BUFX2 BUFX2_81 ( .A(_auto_iopadmap_cc_368_execute_5841_3_), .Y(\Wdata[3] ));
BUFX2 BUFX2_82 ( .A(_auto_iopadmap_cc_368_execute_5841_4_), .Y(\Wdata[4] ));
BUFX2 BUFX2_83 ( .A(_auto_iopadmap_cc_368_execute_5841_5_), .Y(\Wdata[5] ));
BUFX2 BUFX2_84 ( .A(_auto_iopadmap_cc_368_execute_5841_6_), .Y(\Wdata[6] ));
BUFX2 BUFX2_85 ( .A(_auto_iopadmap_cc_368_execute_5841_7_), .Y(\Wdata[7] ));
BUFX2 BUFX2_86 ( .A(_auto_iopadmap_cc_368_execute_5841_8_), .Y(\Wdata[8] ));
BUFX2 BUFX2_87 ( .A(_auto_iopadmap_cc_368_execute_5841_9_), .Y(\Wdata[9] ));
BUFX2 BUFX2_88 ( .A(_auto_iopadmap_cc_368_execute_5841_10_), .Y(\Wdata[10] ));
BUFX2 BUFX2_89 ( .A(_auto_iopadmap_cc_368_execute_5841_11_), .Y(\Wdata[11] ));
BUFX2 BUFX2_9 ( .A(W_R_1_bF_buf5_), .Y(en_instr));
BUFX2 BUFX2_90 ( .A(_auto_iopadmap_cc_368_execute_5841_12_), .Y(\Wdata[12] ));
BUFX2 BUFX2_91 ( .A(_auto_iopadmap_cc_368_execute_5841_13_), .Y(\Wdata[13] ));
BUFX2 BUFX2_92 ( .A(_auto_iopadmap_cc_368_execute_5841_14_), .Y(\Wdata[14] ));
BUFX2 BUFX2_93 ( .A(_auto_iopadmap_cc_368_execute_5841_15_), .Y(\Wdata[15] ));
BUFX2 BUFX2_94 ( .A(_auto_iopadmap_cc_368_execute_5841_16_), .Y(\Wdata[16] ));
BUFX2 BUFX2_95 ( .A(_auto_iopadmap_cc_368_execute_5841_17_), .Y(\Wdata[17] ));
BUFX2 BUFX2_96 ( .A(_auto_iopadmap_cc_368_execute_5841_18_), .Y(\Wdata[18] ));
BUFX2 BUFX2_97 ( .A(_auto_iopadmap_cc_368_execute_5841_19_), .Y(\Wdata[19] ));
BUFX2 BUFX2_98 ( .A(_auto_iopadmap_cc_368_execute_5841_20_), .Y(\Wdata[20] ));
BUFX2 BUFX2_99 ( .A(_auto_iopadmap_cc_368_execute_5841_21_), .Y(\Wdata[21] ));
BUFX4 BUFX4_1 ( .A(clock), .Y(clock_bF_buf7));
BUFX4 BUFX4_10 ( .A(_abc_4635_new_n493_), .Y(_abc_4635_new_n493__bF_buf2));
BUFX4 BUFX4_11 ( .A(_abc_4635_new_n493_), .Y(_abc_4635_new_n493__bF_buf1));
BUFX4 BUFX4_12 ( .A(_abc_4635_new_n493_), .Y(_abc_4635_new_n493__bF_buf0));
BUFX4 BUFX4_13 ( .A(_abc_4635_new_n511_), .Y(_abc_4635_new_n511__bF_buf6));
BUFX4 BUFX4_14 ( .A(_abc_4635_new_n511_), .Y(_abc_4635_new_n511__bF_buf5));
BUFX4 BUFX4_15 ( .A(_abc_4635_new_n511_), .Y(_abc_4635_new_n511__bF_buf4));
BUFX4 BUFX4_16 ( .A(_abc_4635_new_n511_), .Y(_abc_4635_new_n511__bF_buf3));
BUFX4 BUFX4_17 ( .A(_abc_4635_new_n511_), .Y(_abc_4635_new_n511__bF_buf2));
BUFX4 BUFX4_18 ( .A(_abc_4635_new_n511_), .Y(_abc_4635_new_n511__bF_buf1));
BUFX4 BUFX4_19 ( .A(_abc_4635_new_n511_), .Y(_abc_4635_new_n511__bF_buf0));
BUFX4 BUFX4_2 ( .A(clock), .Y(clock_bF_buf6));
BUFX4 BUFX4_20 ( .A(_abc_4635_new_n472_), .Y(_abc_4635_new_n472__bF_buf3));
BUFX4 BUFX4_21 ( .A(_abc_4635_new_n472_), .Y(_abc_4635_new_n472__bF_buf2));
BUFX4 BUFX4_22 ( .A(_abc_4635_new_n472_), .Y(_abc_4635_new_n472__bF_buf1));
BUFX4 BUFX4_23 ( .A(_abc_4635_new_n472_), .Y(_abc_4635_new_n472__bF_buf0));
BUFX4 BUFX4_24 ( .A(_abc_4635_new_n754_), .Y(_abc_4635_new_n754__bF_buf4));
BUFX4 BUFX4_25 ( .A(_abc_4635_new_n754_), .Y(_abc_4635_new_n754__bF_buf3));
BUFX4 BUFX4_26 ( .A(_abc_4635_new_n754_), .Y(_abc_4635_new_n754__bF_buf2));
BUFX4 BUFX4_27 ( .A(_abc_4635_new_n754_), .Y(_abc_4635_new_n754__bF_buf1));
BUFX4 BUFX4_28 ( .A(_abc_4635_new_n754_), .Y(_abc_4635_new_n754__bF_buf0));
BUFX4 BUFX4_29 ( .A(\W_R[1] ), .Y(W_R_1_bF_buf5_));
BUFX4 BUFX4_3 ( .A(clock), .Y(clock_bF_buf5));
BUFX4 BUFX4_30 ( .A(\W_R[1] ), .Y(W_R_1_bF_buf4_));
BUFX4 BUFX4_31 ( .A(\W_R[1] ), .Y(W_R_1_bF_buf3_));
BUFX4 BUFX4_32 ( .A(\W_R[1] ), .Y(W_R_1_bF_buf2_));
BUFX4 BUFX4_33 ( .A(\W_R[1] ), .Y(W_R_1_bF_buf1_));
BUFX4 BUFX4_34 ( .A(\W_R[1] ), .Y(W_R_1_bF_buf0_));
BUFX4 BUFX4_35 ( .A(_abc_4635_new_n616_), .Y(_abc_4635_new_n616__bF_buf4));
BUFX4 BUFX4_36 ( .A(_abc_4635_new_n616_), .Y(_abc_4635_new_n616__bF_buf3));
BUFX4 BUFX4_37 ( .A(_abc_4635_new_n616_), .Y(_abc_4635_new_n616__bF_buf2));
BUFX4 BUFX4_38 ( .A(_abc_4635_new_n616_), .Y(_abc_4635_new_n616__bF_buf1));
BUFX4 BUFX4_39 ( .A(_abc_4635_new_n616_), .Y(_abc_4635_new_n616__bF_buf0));
BUFX4 BUFX4_4 ( .A(clock), .Y(clock_bF_buf4));
BUFX4 BUFX4_40 ( .A(resetn), .Y(resetn_bF_buf5));
BUFX4 BUFX4_41 ( .A(resetn), .Y(resetn_bF_buf4));
BUFX4 BUFX4_42 ( .A(resetn), .Y(resetn_bF_buf3));
BUFX4 BUFX4_43 ( .A(resetn), .Y(resetn_bF_buf2));
BUFX4 BUFX4_44 ( .A(resetn), .Y(resetn_bF_buf1));
BUFX4 BUFX4_45 ( .A(resetn), .Y(resetn_bF_buf0));
BUFX4 BUFX4_46 ( .A(_abc_4635_new_n480_), .Y(_abc_4635_new_n480__bF_buf4));
BUFX4 BUFX4_47 ( .A(_abc_4635_new_n480_), .Y(_abc_4635_new_n480__bF_buf3));
BUFX4 BUFX4_48 ( .A(_abc_4635_new_n753_), .Y(_abc_4635_new_n753__bF_buf4));
BUFX4 BUFX4_49 ( .A(_abc_4635_new_n753_), .Y(_abc_4635_new_n753__bF_buf3));
BUFX4 BUFX4_5 ( .A(clock), .Y(clock_bF_buf3));
BUFX4 BUFX4_50 ( .A(_abc_4635_new_n753_), .Y(_abc_4635_new_n753__bF_buf2));
BUFX4 BUFX4_51 ( .A(_abc_4635_new_n753_), .Y(_abc_4635_new_n753__bF_buf1));
BUFX4 BUFX4_52 ( .A(_abc_4635_new_n753_), .Y(_abc_4635_new_n753__bF_buf0));
BUFX4 BUFX4_53 ( .A(_abc_4635_new_n618_), .Y(_abc_4635_new_n618__bF_buf4));
BUFX4 BUFX4_54 ( .A(_abc_4635_new_n618_), .Y(_abc_4635_new_n618__bF_buf3));
BUFX4 BUFX4_55 ( .A(_abc_4635_new_n618_), .Y(_abc_4635_new_n618__bF_buf2));
BUFX4 BUFX4_56 ( .A(_abc_4635_new_n618_), .Y(_abc_4635_new_n618__bF_buf1));
BUFX4 BUFX4_57 ( .A(_abc_4635_new_n618_), .Y(_abc_4635_new_n618__bF_buf0));
BUFX4 BUFX4_6 ( .A(clock), .Y(clock_bF_buf2));
BUFX4 BUFX4_7 ( .A(clock), .Y(clock_bF_buf1));
BUFX4 BUFX4_8 ( .A(clock), .Y(clock_bF_buf0));
BUFX4 BUFX4_9 ( .A(_abc_4635_new_n493_), .Y(_abc_4635_new_n493__bF_buf3));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock_bF_buf7), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_0_), .Q(state_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock_bF_buf6), .D(_0Wdata_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_5841_2_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock_bF_buf5), .D(_0Wdata_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_5841_3_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock_bF_buf4), .D(_0Wdata_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_5841_4_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock_bF_buf3), .D(_0Wdata_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_5841_5_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock_bF_buf2), .D(_0Wdata_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_5841_6_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock_bF_buf1), .D(_0Wdata_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_5841_7_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock_bF_buf0), .D(_0Wdata_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_5841_8_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock_bF_buf7), .D(_0Wdata_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_5841_9_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock_bF_buf6), .D(_0Wdata_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_5841_10_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock_bF_buf5), .D(_0Wdata_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_5841_11_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock_bF_buf6), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_1_), .Q(state_1_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock_bF_buf4), .D(_0Wdata_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_5841_12_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock_bF_buf3), .D(_0Wdata_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_5841_13_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock_bF_buf2), .D(_0Wdata_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_5841_14_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock_bF_buf1), .D(_0Wdata_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_5841_15_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock_bF_buf0), .D(_0Wdata_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_5841_16_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock_bF_buf7), .D(_0Wdata_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_5841_17_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock_bF_buf6), .D(_0Wdata_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_5841_18_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock_bF_buf5), .D(_0Wdata_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_5841_19_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock_bF_buf4), .D(_0Wdata_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_5841_20_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock_bF_buf3), .D(_0Wdata_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_5841_21_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock_bF_buf5), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_2_), .Q(state_2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock_bF_buf2), .D(_0Wdata_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_5841_22_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock_bF_buf1), .D(_0Wdata_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_5841_23_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock_bF_buf0), .D(_0Wdata_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_5841_24_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clock_bF_buf7), .D(_0Wdata_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_5841_25_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clock_bF_buf6), .D(_0Wdata_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_5841_26_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clock_bF_buf5), .D(_0Wdata_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_5841_27_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clock_bF_buf4), .D(_0Wdata_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_5841_28_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clock_bF_buf3), .D(_0Wdata_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_5841_29_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clock_bF_buf2), .D(_0Wdata_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_5841_30_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clock_bF_buf1), .D(_0Wdata_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_5841_31_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock_bF_buf4), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_3_), .Q(state_3_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clock_bF_buf0), .D(_0inst_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_5894_0_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clock_bF_buf7), .D(_0inst_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_5894_1_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clock_bF_buf6), .D(_0inst_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_5894_2_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clock_bF_buf5), .D(_0inst_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_5894_3_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clock_bF_buf4), .D(_0inst_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_5894_4_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clock_bF_buf3), .D(_0inst_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_5894_5_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clock_bF_buf2), .D(_0inst_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_5894_6_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clock_bF_buf1), .D(_0inst_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_5894_7_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clock_bF_buf0), .D(_0inst_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_5894_8_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock_bF_buf7), .D(_0inst_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_5894_9_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock_bF_buf3), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_4_), .Q(state_4_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock_bF_buf6), .D(_0inst_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_5894_10_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock_bF_buf5), .D(_0inst_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_5894_11_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clock_bF_buf4), .D(_0inst_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_5894_12_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clock_bF_buf3), .D(_0inst_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_5894_13_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clock_bF_buf2), .D(_0inst_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_5894_14_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clock_bF_buf1), .D(_0inst_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_5894_15_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clock_bF_buf0), .D(_0inst_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_5894_16_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clock_bF_buf7), .D(_0inst_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_5894_17_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clock_bF_buf6), .D(_0inst_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_5894_18_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clock_bF_buf5), .D(_0inst_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_5894_19_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock_bF_buf2), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_5_), .Q(state_5_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clock_bF_buf4), .D(_0inst_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_5894_20_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clock_bF_buf3), .D(_0inst_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_5894_21_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clock_bF_buf2), .D(_0inst_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_5894_22_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clock_bF_buf1), .D(_0inst_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_5894_23_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clock_bF_buf0), .D(_0inst_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_5894_24_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clock_bF_buf7), .D(_0inst_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_5894_25_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clock_bF_buf6), .D(_0inst_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_5894_26_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clock_bF_buf5), .D(_0inst_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_5894_27_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clock_bF_buf4), .D(_0inst_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_5894_28_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clock_bF_buf3), .D(_0inst_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_5894_29_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock_bF_buf1), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_6_), .Q(state_6_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clock_bF_buf2), .D(_0inst_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_5894_30_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clock_bF_buf1), .D(_0inst_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_5894_31_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clock_bF_buf0), .D(_0Wstrb_3_0__0_), .Q(_auto_iopadmap_cc_368_execute_5874_0_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clock_bF_buf7), .D(_0Wstrb_3_0__1_), .Q(_auto_iopadmap_cc_368_execute_5874_1_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clock_bF_buf6), .D(_0Wstrb_3_0__2_), .Q(_auto_iopadmap_cc_368_execute_5874_2_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clock_bF_buf5), .D(_0Wstrb_3_0__3_), .Q(_auto_iopadmap_cc_368_execute_5874_3_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock_bF_buf0), .D(_0Wdata_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_5841_0_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock_bF_buf7), .D(_0Wdata_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_5841_1_));
INVX1 INVX1_1 ( .A(Bvalid), .Y(_abc_4635_new_n361_));
INVX1 INVX1_10 ( .A(enable), .Y(_abc_4635_new_n401_));
INVX1 INVX1_100 ( .A(_abc_4635_new_n1406_), .Y(_abc_4635_new_n1407_));
INVX1 INVX1_101 ( .A(_abc_4635_new_n1411_), .Y(_abc_4635_new_n1412_));
INVX1 INVX1_102 ( .A(_abc_4635_new_n1414_), .Y(_abc_4635_new_n1415_));
INVX1 INVX1_103 ( .A(_abc_4635_new_n1416_), .Y(_abc_4635_new_n1418_));
INVX1 INVX1_104 ( .A(_abc_4635_new_n1431_), .Y(_abc_4635_new_n1432_));
INVX1 INVX1_105 ( .A(_abc_4635_new_n1019_), .Y(_abc_4635_new_n1437_));
INVX1 INVX1_106 ( .A(_abc_4635_new_n1022_), .Y(_abc_4635_new_n1439_));
INVX1 INVX1_107 ( .A(_abc_4635_new_n1079_), .Y(_abc_4635_new_n1441_));
INVX1 INVX1_108 ( .A(_abc_4635_new_n1084_), .Y(_abc_4635_new_n1443_));
INVX1 INVX1_109 ( .A(_abc_4635_new_n1203_), .Y(_abc_4635_new_n1445_));
INVX1 INVX1_11 ( .A(resetn_bF_buf0), .Y(_abc_4635_new_n413_));
INVX1 INVX1_110 ( .A(_abc_4635_new_n1210_), .Y(_abc_4635_new_n1447_));
INVX1 INVX1_111 ( .A(_abc_4635_new_n1330_), .Y(_abc_4635_new_n1449_));
INVX1 INVX1_112 ( .A(_abc_4635_new_n1337_), .Y(_abc_4635_new_n1451_));
INVX1 INVX1_113 ( .A(_abc_4635_new_n1394_), .Y(_abc_4635_new_n1453_));
INVX1 INVX1_114 ( .A(_abc_4635_new_n1399_), .Y(_abc_4635_new_n1455_));
INVX1 INVX1_115 ( .A(_abc_4635_new_n1425_), .Y(_abc_4635_new_n1457_));
INVX1 INVX1_116 ( .A(_abc_4635_new_n1428_), .Y(_abc_4635_new_n1459_));
INVX1 INVX1_117 ( .A(_abc_4635_new_n1433_), .Y(_abc_4635_new_n1461_));
INVX1 INVX1_118 ( .A(\imm[31] ), .Y(_abc_4635_new_n1468_));
INVX1 INVX1_119 ( .A(\rs1[31] ), .Y(_abc_4635_new_n1470_));
INVX1 INVX1_12 ( .A(Rvalid), .Y(_abc_4635_new_n428_));
INVX1 INVX1_120 ( .A(_abc_4635_new_n1472_), .Y(_abc_4635_new_n1473_));
INVX1 INVX1_13 ( .A(state_0_), .Y(_abc_4635_new_n433_));
INVX1 INVX1_14 ( .A(state_4_), .Y(_abc_4635_new_n437_));
INVX1 INVX1_15 ( .A(_abc_4635_new_n392_), .Y(_abc_4635_new_n439_));
INVX1 INVX1_16 ( .A(_abc_4635_new_n440_), .Y(_abc_4635_new_n441_));
INVX1 INVX1_17 ( .A(state_1_), .Y(_abc_4635_new_n442_));
INVX1 INVX1_18 ( .A(state_3_), .Y(_abc_4635_new_n446_));
INVX1 INVX1_19 ( .A(state_6_), .Y(_abc_4635_new_n449_));
INVX1 INVX1_2 ( .A(Wready), .Y(_abc_4635_new_n368_));
INVX1 INVX1_20 ( .A(_auto_iopadmap_cc_368_execute_5892), .Y(_auto_iopadmap_cc_368_execute_5890));
INVX1 INVX1_21 ( .A(_abc_4635_new_n462_), .Y(_abc_4635_new_n463_));
INVX1 INVX1_22 ( .A(_abc_4635_new_n460_), .Y(_abc_4635_new_n466_));
INVX1 INVX1_23 ( .A(\imm[1] ), .Y(_abc_4635_new_n467_));
INVX1 INVX1_24 ( .A(\rs1[1] ), .Y(_abc_4635_new_n468_));
INVX1 INVX1_25 ( .A(_abc_4635_new_n476_), .Y(_abc_4635_new_n477_));
INVX1 INVX1_26 ( .A(_abc_4635_new_n478_), .Y(_abc_4635_new_n479_));
INVX1 INVX1_27 ( .A(_abc_4635_new_n480__bF_buf4), .Y(_abc_4635_new_n481_));
INVX1 INVX1_28 ( .A(_abc_4635_new_n483_), .Y(_abc_4635_new_n484_));
INVX1 INVX1_29 ( .A(_abc_4635_new_n512_), .Y(_abc_4635_new_n749_));
INVX1 INVX1_3 ( .A(_abc_4635_new_n369_), .Y(_abc_4635_new_n370_));
INVX1 INVX1_30 ( .A(_abc_4635_new_n995_), .Y(_abc_4635_new_n996_));
INVX1 INVX1_31 ( .A(_abc_4635_new_n999_), .Y(_abc_4635_new_n1000_));
INVX1 INVX1_32 ( .A(_abc_4635_new_n1008_), .Y(_abc_4635_new_n1009_));
INVX1 INVX1_33 ( .A(_abc_4635_new_n1010_), .Y(_abc_4635_new_n1011_));
INVX1 INVX1_34 ( .A(_abc_4635_new_n1006_), .Y(_abc_4635_new_n1013_));
INVX1 INVX1_35 ( .A(_abc_4635_new_n1025_), .Y(_abc_4635_new_n1026_));
INVX1 INVX1_36 ( .A(_abc_4635_new_n1028_), .Y(_abc_4635_new_n1029_));
INVX1 INVX1_37 ( .A(_abc_4635_new_n1035_), .Y(_abc_4635_new_n1036_));
INVX1 INVX1_38 ( .A(_abc_4635_new_n1038_), .Y(_abc_4635_new_n1039_));
INVX1 INVX1_39 ( .A(_abc_4635_new_n1040_), .Y(_abc_4635_new_n1042_));
INVX1 INVX1_4 ( .A(AWready), .Y(_abc_4635_new_n373_));
INVX1 INVX1_40 ( .A(_abc_4635_new_n1054_), .Y(_abc_4635_new_n1055_));
INVX1 INVX1_41 ( .A(_abc_4635_new_n1059_), .Y(_abc_4635_new_n1060_));
INVX1 INVX1_42 ( .A(_abc_4635_new_n1067_), .Y(_abc_4635_new_n1068_));
INVX1 INVX1_43 ( .A(_abc_4635_new_n1069_), .Y(_abc_4635_new_n1070_));
INVX1 INVX1_44 ( .A(_abc_4635_new_n1065_), .Y(_abc_4635_new_n1072_));
INVX1 INVX1_45 ( .A(_abc_4635_new_n1086_), .Y(_abc_4635_new_n1087_));
INVX1 INVX1_46 ( .A(_abc_4635_new_n1091_), .Y(_abc_4635_new_n1092_));
INVX1 INVX1_47 ( .A(_abc_4635_new_n1096_), .Y(_abc_4635_new_n1097_));
INVX1 INVX1_48 ( .A(_abc_4635_new_n1099_), .Y(_abc_4635_new_n1100_));
INVX1 INVX1_49 ( .A(_abc_4635_new_n1101_), .Y(_abc_4635_new_n1103_));
INVX1 INVX1_5 ( .A(_abc_4635_new_n374_), .Y(_abc_4635_new_n375_));
INVX1 INVX1_50 ( .A(_abc_4635_new_n1115_), .Y(_abc_4635_new_n1116_));
INVX1 INVX1_51 ( .A(_abc_4635_new_n1120_), .Y(_abc_4635_new_n1121_));
INVX1 INVX1_52 ( .A(_abc_4635_new_n1125_), .Y(_abc_4635_new_n1126_));
INVX1 INVX1_53 ( .A(_abc_4635_new_n1128_), .Y(_abc_4635_new_n1129_));
INVX1 INVX1_54 ( .A(_abc_4635_new_n1130_), .Y(_abc_4635_new_n1131_));
INVX1 INVX1_55 ( .A(_abc_4635_new_n1148_), .Y(_abc_4635_new_n1149_));
INVX1 INVX1_56 ( .A(_abc_4635_new_n1152_), .Y(_abc_4635_new_n1153_));
INVX1 INVX1_57 ( .A(_abc_4635_new_n1159_), .Y(_abc_4635_new_n1160_));
INVX1 INVX1_58 ( .A(_abc_4635_new_n1157_), .Y(_abc_4635_new_n1163_));
INVX1 INVX1_59 ( .A(_abc_4635_new_n1161_), .Y(_abc_4635_new_n1164_));
INVX1 INVX1_6 ( .A(_abc_4635_new_n377_), .Y(_abc_4635_new_n378_));
INVX1 INVX1_60 ( .A(_abc_4635_new_n1172_), .Y(_abc_4635_new_n1173_));
INVX1 INVX1_61 ( .A(_abc_4635_new_n1177_), .Y(_abc_4635_new_n1178_));
INVX1 INVX1_62 ( .A(_abc_4635_new_n1182_), .Y(_abc_4635_new_n1183_));
INVX1 INVX1_63 ( .A(_abc_4635_new_n1190_), .Y(_abc_4635_new_n1191_));
INVX1 INVX1_64 ( .A(_abc_4635_new_n1192_), .Y(_abc_4635_new_n1193_));
INVX1 INVX1_65 ( .A(_abc_4635_new_n1188_), .Y(_abc_4635_new_n1195_));
INVX1 INVX1_66 ( .A(_abc_4635_new_n1213_), .Y(_abc_4635_new_n1214_));
INVX1 INVX1_67 ( .A(_abc_4635_new_n1217_), .Y(_abc_4635_new_n1218_));
INVX1 INVX1_68 ( .A(_abc_4635_new_n1222_), .Y(_abc_4635_new_n1223_));
INVX1 INVX1_69 ( .A(_abc_4635_new_n1224_), .Y(_abc_4635_new_n1225_));
INVX1 INVX1_7 ( .A(_abc_4635_new_n376_), .Y(_abc_4635_new_n380_));
INVX1 INVX1_70 ( .A(_abc_4635_new_n1227_), .Y(_abc_4635_new_n1229_));
INVX1 INVX1_71 ( .A(_abc_4635_new_n1237_), .Y(_abc_4635_new_n1238_));
INVX1 INVX1_72 ( .A(_abc_4635_new_n1242_), .Y(_abc_4635_new_n1243_));
INVX1 INVX1_73 ( .A(_abc_4635_new_n1247_), .Y(_abc_4635_new_n1248_));
INVX1 INVX1_74 ( .A(_abc_4635_new_n1254_), .Y(_abc_4635_new_n1255_));
INVX1 INVX1_75 ( .A(_abc_4635_new_n1257_), .Y(_abc_4635_new_n1258_));
INVX1 INVX1_76 ( .A(_abc_4635_new_n1253_), .Y(_abc_4635_new_n1260_));
INVX1 INVX1_77 ( .A(_abc_4635_new_n1274_), .Y(_abc_4635_new_n1275_));
INVX1 INVX1_78 ( .A(_abc_4635_new_n1279_), .Y(_abc_4635_new_n1280_));
INVX1 INVX1_79 ( .A(_abc_4635_new_n1284_), .Y(_abc_4635_new_n1285_));
INVX1 INVX1_8 ( .A(ARready), .Y(_abc_4635_new_n389_));
INVX1 INVX1_80 ( .A(_abc_4635_new_n1286_), .Y(_abc_4635_new_n1287_));
INVX1 INVX1_81 ( .A(_abc_4635_new_n1289_), .Y(_abc_4635_new_n1291_));
INVX1 INVX1_82 ( .A(_abc_4635_new_n1299_), .Y(_abc_4635_new_n1300_));
INVX1 INVX1_83 ( .A(_abc_4635_new_n1304_), .Y(_abc_4635_new_n1305_));
INVX1 INVX1_84 ( .A(_abc_4635_new_n1309_), .Y(_abc_4635_new_n1310_));
INVX1 INVX1_85 ( .A(_abc_4635_new_n1316_), .Y(_abc_4635_new_n1317_));
INVX1 INVX1_86 ( .A(_abc_4635_new_n1319_), .Y(_abc_4635_new_n1320_));
INVX1 INVX1_87 ( .A(_abc_4635_new_n1315_), .Y(_abc_4635_new_n1322_));
INVX1 INVX1_88 ( .A(_abc_4635_new_n1339_), .Y(_abc_4635_new_n1340_));
INVX1 INVX1_89 ( .A(_abc_4635_new_n1344_), .Y(_abc_4635_new_n1345_));
INVX1 INVX1_9 ( .A(_abc_4635_new_n390_), .Y(_abc_4635_new_n391_));
INVX1 INVX1_90 ( .A(_abc_4635_new_n1349_), .Y(_abc_4635_new_n1350_));
INVX1 INVX1_91 ( .A(_abc_4635_new_n1351_), .Y(_abc_4635_new_n1352_));
INVX1 INVX1_92 ( .A(_abc_4635_new_n1354_), .Y(_abc_4635_new_n1356_));
INVX1 INVX1_93 ( .A(_abc_4635_new_n1364_), .Y(_abc_4635_new_n1365_));
INVX1 INVX1_94 ( .A(_abc_4635_new_n1369_), .Y(_abc_4635_new_n1370_));
INVX1 INVX1_95 ( .A(_abc_4635_new_n1374_), .Y(_abc_4635_new_n1375_));
INVX1 INVX1_96 ( .A(_abc_4635_new_n1382_), .Y(_abc_4635_new_n1383_));
INVX1 INVX1_97 ( .A(_abc_4635_new_n1384_), .Y(_abc_4635_new_n1385_));
INVX1 INVX1_98 ( .A(_abc_4635_new_n1380_), .Y(_abc_4635_new_n1387_));
INVX1 INVX1_99 ( .A(_abc_4635_new_n1402_), .Y(_abc_4635_new_n1403_));
INVX2 INVX2_1 ( .A(\wordsize[0] ), .Y(_abc_4635_new_n457_));
INVX4 INVX4_1 ( .A(\wordsize[1] ), .Y(_abc_4635_new_n458_));
INVX4 INVX4_2 ( .A(_abc_4635_new_n474_), .Y(_abc_4635_new_n475_));
INVX8 INVX8_1 ( .A(_abc_4635_new_n472__bF_buf0), .Y(_abc_4635_new_n493_));
INVX8 INVX8_2 ( .A(_abc_4635_new_n616__bF_buf3), .Y(_abc_4635_new_n618_));
INVX8 INVX8_3 ( .A(W_R_1_bF_buf2_), .Y(_abc_4635_new_n753_));
OR2X2 OR2X2_1 ( .A(_abc_4635_new_n363_), .B(state_1_), .Y(_abc_4635_new_n364_));
OR2X2 OR2X2_10 ( .A(_abc_4635_new_n407_), .B(_abc_4635_new_n410_), .Y(_abc_4635_new_n411_));
OR2X2 OR2X2_100 ( .A(_abc_4635_new_n743_), .B(_abc_4635_new_n742_), .Y(_abc_4635_new_n744_));
OR2X2 OR2X2_101 ( .A(_abc_4635_new_n401_), .B(W_R_1_bF_buf3_), .Y(_abc_4635_new_n748_));
OR2X2 OR2X2_102 ( .A(_abc_4635_new_n749_), .B(_abc_4635_new_n748_), .Y(_abc_4635_new_n750_));
OR2X2 OR2X2_103 ( .A(_abc_4635_new_n750_), .B(_abc_4635_new_n747_), .Y(_abc_4635_new_n751_));
OR2X2 OR2X2_104 ( .A(_abc_4635_new_n746_), .B(_abc_4635_new_n751_), .Y(_auto_iopadmap_cc_368_execute_5881));
OR2X2 OR2X2_105 ( .A(_abc_4635_new_n472__bF_buf3), .B(\Rdata_mem[16] ), .Y(_abc_4635_new_n755_));
OR2X2 OR2X2_106 ( .A(_abc_4635_new_n493__bF_buf1), .B(\Rdata_mem[8] ), .Y(_abc_4635_new_n757_));
OR2X2 OR2X2_107 ( .A(_abc_4635_new_n472__bF_buf2), .B(\Rdata_mem[24] ), .Y(_abc_4635_new_n758_));
OR2X2 OR2X2_108 ( .A(_abc_4635_new_n760_), .B(_abc_4635_new_n756_), .Y(_abc_4635_new_n761_));
OR2X2 OR2X2_109 ( .A(_abc_4635_new_n478_), .B(_abc_4635_new_n762_), .Y(_abc_4635_new_n763_));
OR2X2 OR2X2_11 ( .A(_abc_4635_new_n414_), .B(_abc_4635_new_n413_), .Y(_abc_4635_new_n415_));
OR2X2 OR2X2_110 ( .A(_abc_4635_new_n493__bF_buf0), .B(\Rdata_mem[0] ), .Y(_abc_4635_new_n766_));
OR2X2 OR2X2_111 ( .A(_abc_4635_new_n768_), .B(_abc_4635_new_n765_), .Y(_abc_4635_new_n769_));
OR2X2 OR2X2_112 ( .A(_abc_4635_new_n764_), .B(_abc_4635_new_n769_), .Y(_abc_4635_new_n770_));
OR2X2 OR2X2_113 ( .A(_abc_4635_new_n493__bF_buf3), .B(\Rdata_mem[9] ), .Y(_abc_4635_new_n772_));
OR2X2 OR2X2_114 ( .A(_abc_4635_new_n472__bF_buf1), .B(\Rdata_mem[25] ), .Y(_abc_4635_new_n773_));
OR2X2 OR2X2_115 ( .A(_abc_4635_new_n472__bF_buf0), .B(\Rdata_mem[17] ), .Y(_abc_4635_new_n776_));
OR2X2 OR2X2_116 ( .A(_abc_4635_new_n775_), .B(_abc_4635_new_n777_), .Y(_abc_4635_new_n778_));
OR2X2 OR2X2_117 ( .A(_abc_4635_new_n478_), .B(_abc_4635_new_n779_), .Y(_abc_4635_new_n780_));
OR2X2 OR2X2_118 ( .A(_abc_4635_new_n493__bF_buf2), .B(\Rdata_mem[1] ), .Y(_abc_4635_new_n783_));
OR2X2 OR2X2_119 ( .A(_abc_4635_new_n785_), .B(_abc_4635_new_n782_), .Y(_abc_4635_new_n786_));
OR2X2 OR2X2_12 ( .A(_abc_4635_new_n412_), .B(_abc_4635_new_n415_), .Y(_abc_4635_new_n416_));
OR2X2 OR2X2_120 ( .A(_abc_4635_new_n781_), .B(_abc_4635_new_n786_), .Y(_abc_4635_new_n787_));
OR2X2 OR2X2_121 ( .A(_abc_4635_new_n493__bF_buf1), .B(\Rdata_mem[10] ), .Y(_abc_4635_new_n789_));
OR2X2 OR2X2_122 ( .A(_abc_4635_new_n472__bF_buf3), .B(\Rdata_mem[26] ), .Y(_abc_4635_new_n790_));
OR2X2 OR2X2_123 ( .A(_abc_4635_new_n472__bF_buf2), .B(\Rdata_mem[18] ), .Y(_abc_4635_new_n793_));
OR2X2 OR2X2_124 ( .A(_abc_4635_new_n792_), .B(_abc_4635_new_n794_), .Y(_abc_4635_new_n795_));
OR2X2 OR2X2_125 ( .A(_abc_4635_new_n478_), .B(_abc_4635_new_n796_), .Y(_abc_4635_new_n797_));
OR2X2 OR2X2_126 ( .A(_abc_4635_new_n493__bF_buf0), .B(\Rdata_mem[2] ), .Y(_abc_4635_new_n800_));
OR2X2 OR2X2_127 ( .A(_abc_4635_new_n802_), .B(_abc_4635_new_n799_), .Y(_abc_4635_new_n803_));
OR2X2 OR2X2_128 ( .A(_abc_4635_new_n798_), .B(_abc_4635_new_n803_), .Y(_abc_4635_new_n804_));
OR2X2 OR2X2_129 ( .A(_abc_4635_new_n493__bF_buf3), .B(\Rdata_mem[11] ), .Y(_abc_4635_new_n806_));
OR2X2 OR2X2_13 ( .A(_abc_4635_new_n416_), .B(_abc_4635_new_n411_), .Y(_abc_4635_new_n417_));
OR2X2 OR2X2_130 ( .A(_abc_4635_new_n472__bF_buf1), .B(\Rdata_mem[27] ), .Y(_abc_4635_new_n807_));
OR2X2 OR2X2_131 ( .A(_abc_4635_new_n472__bF_buf0), .B(\Rdata_mem[19] ), .Y(_abc_4635_new_n810_));
OR2X2 OR2X2_132 ( .A(_abc_4635_new_n809_), .B(_abc_4635_new_n811_), .Y(_abc_4635_new_n812_));
OR2X2 OR2X2_133 ( .A(_abc_4635_new_n478_), .B(_abc_4635_new_n813_), .Y(_abc_4635_new_n814_));
OR2X2 OR2X2_134 ( .A(_abc_4635_new_n493__bF_buf2), .B(\Rdata_mem[3] ), .Y(_abc_4635_new_n817_));
OR2X2 OR2X2_135 ( .A(_abc_4635_new_n819_), .B(_abc_4635_new_n816_), .Y(_abc_4635_new_n820_));
OR2X2 OR2X2_136 ( .A(_abc_4635_new_n815_), .B(_abc_4635_new_n820_), .Y(_abc_4635_new_n821_));
OR2X2 OR2X2_137 ( .A(_abc_4635_new_n472__bF_buf3), .B(\Rdata_mem[20] ), .Y(_abc_4635_new_n823_));
OR2X2 OR2X2_138 ( .A(_abc_4635_new_n493__bF_buf1), .B(\Rdata_mem[12] ), .Y(_abc_4635_new_n825_));
OR2X2 OR2X2_139 ( .A(_abc_4635_new_n472__bF_buf2), .B(\Rdata_mem[28] ), .Y(_abc_4635_new_n826_));
OR2X2 OR2X2_14 ( .A(_abc_4635_new_n417_), .B(_abc_4635_new_n406_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_0_));
OR2X2 OR2X2_140 ( .A(_abc_4635_new_n828_), .B(_abc_4635_new_n824_), .Y(_abc_4635_new_n829_));
OR2X2 OR2X2_141 ( .A(_abc_4635_new_n478_), .B(_abc_4635_new_n830_), .Y(_abc_4635_new_n831_));
OR2X2 OR2X2_142 ( .A(_abc_4635_new_n493__bF_buf0), .B(\Rdata_mem[4] ), .Y(_abc_4635_new_n834_));
OR2X2 OR2X2_143 ( .A(_abc_4635_new_n836_), .B(_abc_4635_new_n833_), .Y(_abc_4635_new_n837_));
OR2X2 OR2X2_144 ( .A(_abc_4635_new_n832_), .B(_abc_4635_new_n837_), .Y(_abc_4635_new_n838_));
OR2X2 OR2X2_145 ( .A(_abc_4635_new_n472__bF_buf1), .B(\Rdata_mem[21] ), .Y(_abc_4635_new_n840_));
OR2X2 OR2X2_146 ( .A(_abc_4635_new_n493__bF_buf3), .B(\Rdata_mem[13] ), .Y(_abc_4635_new_n842_));
OR2X2 OR2X2_147 ( .A(_abc_4635_new_n472__bF_buf0), .B(\Rdata_mem[29] ), .Y(_abc_4635_new_n843_));
OR2X2 OR2X2_148 ( .A(_abc_4635_new_n845_), .B(_abc_4635_new_n841_), .Y(_abc_4635_new_n846_));
OR2X2 OR2X2_149 ( .A(_abc_4635_new_n478_), .B(_abc_4635_new_n847_), .Y(_abc_4635_new_n848_));
OR2X2 OR2X2_15 ( .A(_abc_4635_new_n421_), .B(state_3_), .Y(_abc_4635_new_n422_));
OR2X2 OR2X2_150 ( .A(_abc_4635_new_n493__bF_buf2), .B(\Rdata_mem[5] ), .Y(_abc_4635_new_n851_));
OR2X2 OR2X2_151 ( .A(_abc_4635_new_n853_), .B(_abc_4635_new_n850_), .Y(_abc_4635_new_n854_));
OR2X2 OR2X2_152 ( .A(_abc_4635_new_n849_), .B(_abc_4635_new_n854_), .Y(_abc_4635_new_n855_));
OR2X2 OR2X2_153 ( .A(_abc_4635_new_n493__bF_buf1), .B(\Rdata_mem[14] ), .Y(_abc_4635_new_n857_));
OR2X2 OR2X2_154 ( .A(_abc_4635_new_n472__bF_buf3), .B(\Rdata_mem[30] ), .Y(_abc_4635_new_n858_));
OR2X2 OR2X2_155 ( .A(_abc_4635_new_n472__bF_buf2), .B(\Rdata_mem[22] ), .Y(_abc_4635_new_n861_));
OR2X2 OR2X2_156 ( .A(_abc_4635_new_n860_), .B(_abc_4635_new_n862_), .Y(_abc_4635_new_n863_));
OR2X2 OR2X2_157 ( .A(_abc_4635_new_n478_), .B(_abc_4635_new_n864_), .Y(_abc_4635_new_n865_));
OR2X2 OR2X2_158 ( .A(_abc_4635_new_n493__bF_buf0), .B(\Rdata_mem[6] ), .Y(_abc_4635_new_n868_));
OR2X2 OR2X2_159 ( .A(_abc_4635_new_n870_), .B(_abc_4635_new_n867_), .Y(_abc_4635_new_n871_));
OR2X2 OR2X2_16 ( .A(_abc_4635_new_n419_), .B(_abc_4635_new_n423_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_3_));
OR2X2 OR2X2_160 ( .A(_abc_4635_new_n866_), .B(_abc_4635_new_n871_), .Y(_abc_4635_new_n872_));
OR2X2 OR2X2_161 ( .A(_abc_4635_new_n877_), .B(_abc_4635_new_n875_), .Y(_abc_4635_new_n878_));
OR2X2 OR2X2_162 ( .A(_abc_4635_new_n880_), .B(_abc_4635_new_n881_), .Y(_abc_4635_new_n882_));
OR2X2 OR2X2_163 ( .A(_abc_4635_new_n878_), .B(_abc_4635_new_n882_), .Y(_abc_4635_new_n883_));
OR2X2 OR2X2_164 ( .A(_abc_4635_new_n493__bF_buf1), .B(\Rdata_mem[7] ), .Y(_abc_4635_new_n886_));
OR2X2 OR2X2_165 ( .A(_abc_4635_new_n472__bF_buf0), .B(\Rdata_mem[23] ), .Y(_abc_4635_new_n887_));
OR2X2 OR2X2_166 ( .A(_abc_4635_new_n889_), .B(_abc_4635_new_n885_), .Y(_abc_4635_new_n890_));
OR2X2 OR2X2_167 ( .A(_abc_4635_new_n884_), .B(_abc_4635_new_n890_), .Y(_abc_4635_new_n891_));
OR2X2 OR2X2_168 ( .A(_abc_4635_new_n896_), .B(_abc_4635_new_n895_), .Y(_abc_4635_new_n897_));
OR2X2 OR2X2_169 ( .A(_abc_4635_new_n894_), .B(_abc_4635_new_n897_), .Y(_abc_4635_new_n898_));
OR2X2 OR2X2_17 ( .A(_abc_4635_new_n382_), .B(state_4_), .Y(_abc_4635_new_n425_));
OR2X2 OR2X2_170 ( .A(_abc_4635_new_n901_), .B(_abc_4635_new_n900_), .Y(_abc_4635_new_n902_));
OR2X2 OR2X2_171 ( .A(_abc_4635_new_n894_), .B(_abc_4635_new_n902_), .Y(_abc_4635_new_n903_));
OR2X2 OR2X2_172 ( .A(_abc_4635_new_n906_), .B(_abc_4635_new_n905_), .Y(_abc_4635_new_n907_));
OR2X2 OR2X2_173 ( .A(_abc_4635_new_n894_), .B(_abc_4635_new_n907_), .Y(_abc_4635_new_n908_));
OR2X2 OR2X2_174 ( .A(_abc_4635_new_n911_), .B(_abc_4635_new_n910_), .Y(_abc_4635_new_n912_));
OR2X2 OR2X2_175 ( .A(_abc_4635_new_n894_), .B(_abc_4635_new_n912_), .Y(_abc_4635_new_n913_));
OR2X2 OR2X2_176 ( .A(_abc_4635_new_n916_), .B(_abc_4635_new_n915_), .Y(_abc_4635_new_n917_));
OR2X2 OR2X2_177 ( .A(_abc_4635_new_n894_), .B(_abc_4635_new_n917_), .Y(_abc_4635_new_n918_));
OR2X2 OR2X2_178 ( .A(_abc_4635_new_n921_), .B(_abc_4635_new_n920_), .Y(_abc_4635_new_n922_));
OR2X2 OR2X2_179 ( .A(_abc_4635_new_n894_), .B(_abc_4635_new_n922_), .Y(_abc_4635_new_n923_));
OR2X2 OR2X2_18 ( .A(_abc_4635_new_n430_), .B(_abc_4635_new_n429_), .Y(_abc_4635_new_n431_));
OR2X2 OR2X2_180 ( .A(_abc_4635_new_n926_), .B(_abc_4635_new_n925_), .Y(_abc_4635_new_n927_));
OR2X2 OR2X2_181 ( .A(_abc_4635_new_n894_), .B(_abc_4635_new_n927_), .Y(_abc_4635_new_n928_));
OR2X2 OR2X2_182 ( .A(_abc_4635_new_n472__bF_buf3), .B(\Rdata_mem[31] ), .Y(_abc_4635_new_n931_));
OR2X2 OR2X2_183 ( .A(_abc_4635_new_n493__bF_buf0), .B(\Rdata_mem[15] ), .Y(_abc_4635_new_n932_));
OR2X2 OR2X2_184 ( .A(_abc_4635_new_n934_), .B(_abc_4635_new_n930_), .Y(_abc_4635_new_n935_));
OR2X2 OR2X2_185 ( .A(_abc_4635_new_n894_), .B(_abc_4635_new_n935_), .Y(_abc_4635_new_n936_));
OR2X2 OR2X2_186 ( .A(_abc_4635_new_n894_), .B(_abc_4635_new_n939_), .Y(_abc_4635_new_n940_));
OR2X2 OR2X2_187 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n938_), .Y(_abc_4635_new_n941_));
OR2X2 OR2X2_188 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n943_), .Y(_abc_4635_new_n944_));
OR2X2 OR2X2_189 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n946_), .Y(_abc_4635_new_n947_));
OR2X2 OR2X2_19 ( .A(_abc_4635_new_n434_), .B(_abc_4635_new_n433_), .Y(_abc_4635_new_n435_));
OR2X2 OR2X2_190 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n949_), .Y(_abc_4635_new_n950_));
OR2X2 OR2X2_191 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n952_), .Y(_abc_4635_new_n953_));
OR2X2 OR2X2_192 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n955_), .Y(_abc_4635_new_n956_));
OR2X2 OR2X2_193 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n958_), .Y(_abc_4635_new_n959_));
OR2X2 OR2X2_194 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n961_), .Y(_abc_4635_new_n962_));
OR2X2 OR2X2_195 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n964_), .Y(_abc_4635_new_n965_));
OR2X2 OR2X2_196 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n967_), .Y(_abc_4635_new_n968_));
OR2X2 OR2X2_197 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n970_), .Y(_abc_4635_new_n971_));
OR2X2 OR2X2_198 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n973_), .Y(_abc_4635_new_n974_));
OR2X2 OR2X2_199 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n976_), .Y(_abc_4635_new_n977_));
OR2X2 OR2X2_2 ( .A(_abc_4635_new_n364_), .B(_abc_4635_new_n362_), .Y(_abc_4635_new_n365_));
OR2X2 OR2X2_20 ( .A(_abc_4635_new_n435_), .B(_abc_4635_new_n405_), .Y(_abc_4635_new_n436_));
OR2X2 OR2X2_200 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n979_), .Y(_abc_4635_new_n980_));
OR2X2 OR2X2_201 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n982_), .Y(_abc_4635_new_n983_));
OR2X2 OR2X2_202 ( .A(_abc_4635_new_n940_), .B(_abc_4635_new_n985_), .Y(_abc_4635_new_n986_));
OR2X2 OR2X2_203 ( .A(_abc_4635_new_n474_), .B(W_R_1_bF_buf1_), .Y(_abc_4635_new_n988_));
OR2X2 OR2X2_204 ( .A(_abc_4635_new_n753__bF_buf3), .B(\pc[0] ), .Y(_abc_4635_new_n989_));
OR2X2 OR2X2_205 ( .A(_abc_4635_new_n493__bF_buf3), .B(W_R_1_bF_buf0_), .Y(_abc_4635_new_n991_));
OR2X2 OR2X2_206 ( .A(_abc_4635_new_n753__bF_buf2), .B(\pc[1] ), .Y(_abc_4635_new_n992_));
OR2X2 OR2X2_207 ( .A(_abc_4635_new_n465_), .B(_abc_4635_new_n462_), .Y(_abc_4635_new_n994_));
OR2X2 OR2X2_208 ( .A(\imm[2] ), .B(\rs1[2] ), .Y(_abc_4635_new_n997_));
OR2X2 OR2X2_209 ( .A(_abc_4635_new_n994_), .B(_abc_4635_new_n998_), .Y(_abc_4635_new_n1001_));
OR2X2 OR2X2_21 ( .A(_abc_4635_new_n403_), .B(_abc_4635_new_n437_), .Y(_abc_4635_new_n438_));
OR2X2 OR2X2_210 ( .A(_abc_4635_new_n1002_), .B(W_R_1_bF_buf5_), .Y(_abc_4635_new_n1003_));
OR2X2 OR2X2_211 ( .A(_abc_4635_new_n753__bF_buf1), .B(\pc[2] ), .Y(_abc_4635_new_n1004_));
OR2X2 OR2X2_212 ( .A(\imm[3] ), .B(\rs1[3] ), .Y(_abc_4635_new_n1007_));
OR2X2 OR2X2_213 ( .A(_abc_4635_new_n1006_), .B(_abc_4635_new_n1011_), .Y(_abc_4635_new_n1012_));
OR2X2 OR2X2_214 ( .A(_abc_4635_new_n1013_), .B(_abc_4635_new_n1010_), .Y(_abc_4635_new_n1014_));
OR2X2 OR2X2_215 ( .A(_abc_4635_new_n1015_), .B(W_R_1_bF_buf4_), .Y(_abc_4635_new_n1016_));
OR2X2 OR2X2_216 ( .A(_abc_4635_new_n753__bF_buf0), .B(\pc[3] ), .Y(_abc_4635_new_n1017_));
OR2X2 OR2X2_217 ( .A(_abc_4635_new_n1021_), .B(_abc_4635_new_n1008_), .Y(_abc_4635_new_n1022_));
OR2X2 OR2X2_218 ( .A(_abc_4635_new_n1020_), .B(_abc_4635_new_n1022_), .Y(_abc_4635_new_n1023_));
OR2X2 OR2X2_219 ( .A(\imm[4] ), .B(\rs1[4] ), .Y(_abc_4635_new_n1024_));
OR2X2 OR2X2_22 ( .A(_abc_4635_new_n442_), .B(Bvalid), .Y(_abc_4635_new_n443_));
OR2X2 OR2X2_220 ( .A(_abc_4635_new_n1023_), .B(_abc_4635_new_n1027_), .Y(_abc_4635_new_n1030_));
OR2X2 OR2X2_221 ( .A(_abc_4635_new_n1031_), .B(W_R_1_bF_buf3_), .Y(_abc_4635_new_n1032_));
OR2X2 OR2X2_222 ( .A(_abc_4635_new_n753__bF_buf4), .B(\pc[4] ), .Y(_abc_4635_new_n1033_));
OR2X2 OR2X2_223 ( .A(\imm[5] ), .B(\rs1[5] ), .Y(_abc_4635_new_n1037_));
OR2X2 OR2X2_224 ( .A(_abc_4635_new_n1036_), .B(_abc_4635_new_n1040_), .Y(_abc_4635_new_n1041_));
OR2X2 OR2X2_225 ( .A(_abc_4635_new_n1035_), .B(_abc_4635_new_n1042_), .Y(_abc_4635_new_n1043_));
OR2X2 OR2X2_226 ( .A(_abc_4635_new_n1044_), .B(W_R_1_bF_buf2_), .Y(_abc_4635_new_n1045_));
OR2X2 OR2X2_227 ( .A(_abc_4635_new_n753__bF_buf3), .B(\pc[5] ), .Y(_abc_4635_new_n1046_));
OR2X2 OR2X2_228 ( .A(_abc_4635_new_n1025_), .B(_abc_4635_new_n1038_), .Y(_abc_4635_new_n1049_));
OR2X2 OR2X2_229 ( .A(_abc_4635_new_n1052_), .B(_abc_4635_new_n1050_), .Y(_abc_4635_new_n1053_));
OR2X2 OR2X2_23 ( .A(_abc_4635_new_n447_), .B(_abc_4635_new_n446_), .Y(_abc_4635_new_n448_));
OR2X2 OR2X2_230 ( .A(\imm[6] ), .B(\rs1[6] ), .Y(_abc_4635_new_n1056_));
OR2X2 OR2X2_231 ( .A(_abc_4635_new_n1053_), .B(_abc_4635_new_n1057_), .Y(_abc_4635_new_n1058_));
OR2X2 OR2X2_232 ( .A(_abc_4635_new_n1062_), .B(_abc_4635_new_n1048_), .Y(_auto_iopadmap_cc_368_execute_5767_6_));
OR2X2 OR2X2_233 ( .A(_abc_4635_new_n753__bF_buf1), .B(\pc[7] ), .Y(_abc_4635_new_n1064_));
OR2X2 OR2X2_234 ( .A(\imm[7] ), .B(\rs1[7] ), .Y(_abc_4635_new_n1066_));
OR2X2 OR2X2_235 ( .A(_abc_4635_new_n1065_), .B(_abc_4635_new_n1070_), .Y(_abc_4635_new_n1071_));
OR2X2 OR2X2_236 ( .A(_abc_4635_new_n1072_), .B(_abc_4635_new_n1069_), .Y(_abc_4635_new_n1073_));
OR2X2 OR2X2_237 ( .A(_abc_4635_new_n1074_), .B(W_R_1_bF_buf0_), .Y(_abc_4635_new_n1075_));
OR2X2 OR2X2_238 ( .A(_abc_4635_new_n1082_), .B(_abc_4635_new_n1067_), .Y(_abc_4635_new_n1083_));
OR2X2 OR2X2_239 ( .A(_abc_4635_new_n1081_), .B(_abc_4635_new_n1083_), .Y(_abc_4635_new_n1084_));
OR2X2 OR2X2_24 ( .A(_abc_4635_new_n402_), .B(_abc_4635_new_n449_), .Y(_abc_4635_new_n450_));
OR2X2 OR2X2_240 ( .A(_abc_4635_new_n1080_), .B(_abc_4635_new_n1084_), .Y(_abc_4635_new_n1085_));
OR2X2 OR2X2_241 ( .A(\imm[8] ), .B(\rs1[8] ), .Y(_abc_4635_new_n1088_));
OR2X2 OR2X2_242 ( .A(_abc_4635_new_n1085_), .B(_abc_4635_new_n1089_), .Y(_abc_4635_new_n1090_));
OR2X2 OR2X2_243 ( .A(_abc_4635_new_n1094_), .B(_abc_4635_new_n1077_), .Y(_auto_iopadmap_cc_368_execute_5767_8_));
OR2X2 OR2X2_244 ( .A(\imm[9] ), .B(\rs1[9] ), .Y(_abc_4635_new_n1098_));
OR2X2 OR2X2_245 ( .A(_abc_4635_new_n1097_), .B(_abc_4635_new_n1101_), .Y(_abc_4635_new_n1102_));
OR2X2 OR2X2_246 ( .A(_abc_4635_new_n1096_), .B(_abc_4635_new_n1103_), .Y(_abc_4635_new_n1104_));
OR2X2 OR2X2_247 ( .A(_abc_4635_new_n1105_), .B(W_R_1_bF_buf4_), .Y(_abc_4635_new_n1106_));
OR2X2 OR2X2_248 ( .A(_abc_4635_new_n753__bF_buf4), .B(\pc[9] ), .Y(_abc_4635_new_n1107_));
OR2X2 OR2X2_249 ( .A(_abc_4635_new_n1086_), .B(_abc_4635_new_n1099_), .Y(_abc_4635_new_n1110_));
OR2X2 OR2X2_25 ( .A(_abc_4635_new_n454_), .B(_abc_4635_new_n413_), .Y(_auto_iopadmap_cc_368_execute_5892));
OR2X2 OR2X2_250 ( .A(_abc_4635_new_n1113_), .B(_abc_4635_new_n1111_), .Y(_abc_4635_new_n1114_));
OR2X2 OR2X2_251 ( .A(\imm[10] ), .B(\rs1[10] ), .Y(_abc_4635_new_n1117_));
OR2X2 OR2X2_252 ( .A(_abc_4635_new_n1114_), .B(_abc_4635_new_n1118_), .Y(_abc_4635_new_n1119_));
OR2X2 OR2X2_253 ( .A(_abc_4635_new_n1123_), .B(_abc_4635_new_n1109_), .Y(_auto_iopadmap_cc_368_execute_5767_10_));
OR2X2 OR2X2_254 ( .A(\imm[11] ), .B(\rs1[11] ), .Y(_abc_4635_new_n1127_));
OR2X2 OR2X2_255 ( .A(_abc_4635_new_n1132_), .B(_abc_4635_new_n1133_), .Y(_abc_4635_new_n1134_));
OR2X2 OR2X2_256 ( .A(_abc_4635_new_n1135_), .B(_abc_4635_new_n1136_), .Y(_auto_iopadmap_cc_368_execute_5767_11_));
OR2X2 OR2X2_257 ( .A(_abc_4635_new_n1141_), .B(_abc_4635_new_n1128_), .Y(_abc_4635_new_n1142_));
OR2X2 OR2X2_258 ( .A(_abc_4635_new_n1140_), .B(_abc_4635_new_n1142_), .Y(_abc_4635_new_n1143_));
OR2X2 OR2X2_259 ( .A(_abc_4635_new_n1145_), .B(_abc_4635_new_n1143_), .Y(_abc_4635_new_n1146_));
OR2X2 OR2X2_26 ( .A(\imm[1] ), .B(\rs1[1] ), .Y(_abc_4635_new_n461_));
OR2X2 OR2X2_260 ( .A(\imm[12] ), .B(\rs1[12] ), .Y(_abc_4635_new_n1147_));
OR2X2 OR2X2_261 ( .A(_abc_4635_new_n1146_), .B(_abc_4635_new_n1150_), .Y(_abc_4635_new_n1151_));
OR2X2 OR2X2_262 ( .A(_abc_4635_new_n1155_), .B(_abc_4635_new_n1138_), .Y(_auto_iopadmap_cc_368_execute_5767_12_));
OR2X2 OR2X2_263 ( .A(\imm[13] ), .B(\rs1[13] ), .Y(_abc_4635_new_n1158_));
OR2X2 OR2X2_264 ( .A(_abc_4635_new_n1165_), .B(_abc_4635_new_n1162_), .Y(_abc_4635_new_n1166_));
OR2X2 OR2X2_265 ( .A(_abc_4635_new_n1167_), .B(_abc_4635_new_n1168_), .Y(_auto_iopadmap_cc_368_execute_5767_13_));
OR2X2 OR2X2_266 ( .A(_abc_4635_new_n1164_), .B(_abc_4635_new_n1149_), .Y(_abc_4635_new_n1171_));
OR2X2 OR2X2_267 ( .A(_abc_4635_new_n1175_), .B(_abc_4635_new_n1173_), .Y(_abc_4635_new_n1176_));
OR2X2 OR2X2_268 ( .A(\imm[14] ), .B(\rs1[14] ), .Y(_abc_4635_new_n1179_));
OR2X2 OR2X2_269 ( .A(_abc_4635_new_n1176_), .B(_abc_4635_new_n1180_), .Y(_abc_4635_new_n1181_));
OR2X2 OR2X2_27 ( .A(_abc_4635_new_n469_), .B(_abc_4635_new_n462_), .Y(_abc_4635_new_n470_));
OR2X2 OR2X2_270 ( .A(_abc_4635_new_n1185_), .B(_abc_4635_new_n1170_), .Y(_auto_iopadmap_cc_368_execute_5767_14_));
OR2X2 OR2X2_271 ( .A(_abc_4635_new_n753__bF_buf3), .B(\pc[15] ), .Y(_abc_4635_new_n1187_));
OR2X2 OR2X2_272 ( .A(\imm[15] ), .B(\rs1[15] ), .Y(_abc_4635_new_n1189_));
OR2X2 OR2X2_273 ( .A(_abc_4635_new_n1188_), .B(_abc_4635_new_n1193_), .Y(_abc_4635_new_n1194_));
OR2X2 OR2X2_274 ( .A(_abc_4635_new_n1195_), .B(_abc_4635_new_n1192_), .Y(_abc_4635_new_n1196_));
OR2X2 OR2X2_275 ( .A(_abc_4635_new_n1197_), .B(W_R_1_bF_buf4_), .Y(_abc_4635_new_n1198_));
OR2X2 OR2X2_276 ( .A(_abc_4635_new_n1206_), .B(_abc_4635_new_n1190_), .Y(_abc_4635_new_n1207_));
OR2X2 OR2X2_277 ( .A(_abc_4635_new_n1208_), .B(_abc_4635_new_n1207_), .Y(_abc_4635_new_n1209_));
OR2X2 OR2X2_278 ( .A(_abc_4635_new_n1209_), .B(_abc_4635_new_n1205_), .Y(_abc_4635_new_n1210_));
OR2X2 OR2X2_279 ( .A(_abc_4635_new_n1204_), .B(_abc_4635_new_n1210_), .Y(_abc_4635_new_n1211_));
OR2X2 OR2X2_28 ( .A(_abc_4635_new_n471_), .B(_abc_4635_new_n465_), .Y(_abc_4635_new_n472_));
OR2X2 OR2X2_280 ( .A(\imm[16] ), .B(\rs1[16] ), .Y(_abc_4635_new_n1212_));
OR2X2 OR2X2_281 ( .A(_abc_4635_new_n1211_), .B(_abc_4635_new_n1215_), .Y(_abc_4635_new_n1216_));
OR2X2 OR2X2_282 ( .A(_abc_4635_new_n1220_), .B(_abc_4635_new_n1200_), .Y(_auto_iopadmap_cc_368_execute_5767_16_));
OR2X2 OR2X2_283 ( .A(\imm[17] ), .B(\rs1[17] ), .Y(_abc_4635_new_n1226_));
OR2X2 OR2X2_284 ( .A(_abc_4635_new_n1223_), .B(_abc_4635_new_n1227_), .Y(_abc_4635_new_n1228_));
OR2X2 OR2X2_285 ( .A(_abc_4635_new_n1222_), .B(_abc_4635_new_n1229_), .Y(_abc_4635_new_n1230_));
OR2X2 OR2X2_286 ( .A(_abc_4635_new_n1231_), .B(W_R_1_bF_buf2_), .Y(_abc_4635_new_n1232_));
OR2X2 OR2X2_287 ( .A(_abc_4635_new_n753__bF_buf1), .B(\pc[17] ), .Y(_abc_4635_new_n1233_));
OR2X2 OR2X2_288 ( .A(_abc_4635_new_n1229_), .B(_abc_4635_new_n1214_), .Y(_abc_4635_new_n1236_));
OR2X2 OR2X2_289 ( .A(_abc_4635_new_n1240_), .B(_abc_4635_new_n1238_), .Y(_abc_4635_new_n1241_));
OR2X2 OR2X2_29 ( .A(\imm[0] ), .B(\rs1[0] ), .Y(_abc_4635_new_n473_));
OR2X2 OR2X2_290 ( .A(\imm[18] ), .B(\rs1[18] ), .Y(_abc_4635_new_n1244_));
OR2X2 OR2X2_291 ( .A(_abc_4635_new_n1241_), .B(_abc_4635_new_n1245_), .Y(_abc_4635_new_n1246_));
OR2X2 OR2X2_292 ( .A(_abc_4635_new_n1250_), .B(_abc_4635_new_n1235_), .Y(_auto_iopadmap_cc_368_execute_5767_18_));
OR2X2 OR2X2_293 ( .A(_abc_4635_new_n753__bF_buf4), .B(\pc[19] ), .Y(_abc_4635_new_n1252_));
OR2X2 OR2X2_294 ( .A(\imm[19] ), .B(\rs1[19] ), .Y(_abc_4635_new_n1256_));
OR2X2 OR2X2_295 ( .A(_abc_4635_new_n1253_), .B(_abc_4635_new_n1258_), .Y(_abc_4635_new_n1259_));
OR2X2 OR2X2_296 ( .A(_abc_4635_new_n1260_), .B(_abc_4635_new_n1257_), .Y(_abc_4635_new_n1261_));
OR2X2 OR2X2_297 ( .A(_abc_4635_new_n1262_), .B(W_R_1_bF_buf0_), .Y(_abc_4635_new_n1263_));
OR2X2 OR2X2_298 ( .A(_abc_4635_new_n1268_), .B(_abc_4635_new_n1254_), .Y(_abc_4635_new_n1269_));
OR2X2 OR2X2_299 ( .A(_abc_4635_new_n1267_), .B(_abc_4635_new_n1269_), .Y(_abc_4635_new_n1270_));
OR2X2 OR2X2_3 ( .A(\W_R[0] ), .B(W_R_1_bF_buf5_), .Y(_abc_4635_new_n376_));
OR2X2 OR2X2_30 ( .A(_abc_4635_new_n472__bF_buf2), .B(_abc_4635_new_n481_), .Y(_abc_4635_new_n482_));
OR2X2 OR2X2_300 ( .A(_abc_4635_new_n1272_), .B(_abc_4635_new_n1270_), .Y(_abc_4635_new_n1273_));
OR2X2 OR2X2_301 ( .A(\imm[20] ), .B(\rs1[20] ), .Y(_abc_4635_new_n1276_));
OR2X2 OR2X2_302 ( .A(_abc_4635_new_n1273_), .B(_abc_4635_new_n1277_), .Y(_abc_4635_new_n1278_));
OR2X2 OR2X2_303 ( .A(_abc_4635_new_n1282_), .B(_abc_4635_new_n1265_), .Y(_auto_iopadmap_cc_368_execute_5767_20_));
OR2X2 OR2X2_304 ( .A(\imm[21] ), .B(\rs1[21] ), .Y(_abc_4635_new_n1288_));
OR2X2 OR2X2_305 ( .A(_abc_4635_new_n1285_), .B(_abc_4635_new_n1289_), .Y(_abc_4635_new_n1290_));
OR2X2 OR2X2_306 ( .A(_abc_4635_new_n1284_), .B(_abc_4635_new_n1291_), .Y(_abc_4635_new_n1292_));
OR2X2 OR2X2_307 ( .A(_abc_4635_new_n1293_), .B(W_R_1_bF_buf4_), .Y(_abc_4635_new_n1294_));
OR2X2 OR2X2_308 ( .A(_abc_4635_new_n753__bF_buf2), .B(\pc[21] ), .Y(_abc_4635_new_n1295_));
OR2X2 OR2X2_309 ( .A(_abc_4635_new_n1291_), .B(_abc_4635_new_n1275_), .Y(_abc_4635_new_n1298_));
OR2X2 OR2X2_31 ( .A(_abc_4635_new_n474_), .B(\wordsize[0] ), .Y(_abc_4635_new_n489_));
OR2X2 OR2X2_310 ( .A(_abc_4635_new_n1302_), .B(_abc_4635_new_n1300_), .Y(_abc_4635_new_n1303_));
OR2X2 OR2X2_311 ( .A(\imm[22] ), .B(\rs1[22] ), .Y(_abc_4635_new_n1306_));
OR2X2 OR2X2_312 ( .A(_abc_4635_new_n1303_), .B(_abc_4635_new_n1307_), .Y(_abc_4635_new_n1308_));
OR2X2 OR2X2_313 ( .A(_abc_4635_new_n1312_), .B(_abc_4635_new_n1297_), .Y(_auto_iopadmap_cc_368_execute_5767_22_));
OR2X2 OR2X2_314 ( .A(_abc_4635_new_n753__bF_buf0), .B(\pc[23] ), .Y(_abc_4635_new_n1314_));
OR2X2 OR2X2_315 ( .A(\imm[23] ), .B(\rs1[23] ), .Y(_abc_4635_new_n1318_));
OR2X2 OR2X2_316 ( .A(_abc_4635_new_n1315_), .B(_abc_4635_new_n1320_), .Y(_abc_4635_new_n1321_));
OR2X2 OR2X2_317 ( .A(_abc_4635_new_n1322_), .B(_abc_4635_new_n1319_), .Y(_abc_4635_new_n1323_));
OR2X2 OR2X2_318 ( .A(_abc_4635_new_n1324_), .B(W_R_1_bF_buf2_), .Y(_abc_4635_new_n1325_));
OR2X2 OR2X2_319 ( .A(_abc_4635_new_n1334_), .B(_abc_4635_new_n1316_), .Y(_abc_4635_new_n1335_));
OR2X2 OR2X2_32 ( .A(_abc_4635_new_n490_), .B(\wordsize[1] ), .Y(_abc_4635_new_n491_));
OR2X2 OR2X2_320 ( .A(_abc_4635_new_n1333_), .B(_abc_4635_new_n1335_), .Y(_abc_4635_new_n1336_));
OR2X2 OR2X2_321 ( .A(_abc_4635_new_n1332_), .B(_abc_4635_new_n1336_), .Y(_abc_4635_new_n1337_));
OR2X2 OR2X2_322 ( .A(_abc_4635_new_n1331_), .B(_abc_4635_new_n1337_), .Y(_abc_4635_new_n1338_));
OR2X2 OR2X2_323 ( .A(\imm[24] ), .B(\rs1[24] ), .Y(_abc_4635_new_n1341_));
OR2X2 OR2X2_324 ( .A(_abc_4635_new_n1338_), .B(_abc_4635_new_n1342_), .Y(_abc_4635_new_n1343_));
OR2X2 OR2X2_325 ( .A(_abc_4635_new_n1347_), .B(_abc_4635_new_n1327_), .Y(_auto_iopadmap_cc_368_execute_5767_24_));
OR2X2 OR2X2_326 ( .A(\imm[25] ), .B(\rs1[25] ), .Y(_abc_4635_new_n1353_));
OR2X2 OR2X2_327 ( .A(_abc_4635_new_n1350_), .B(_abc_4635_new_n1354_), .Y(_abc_4635_new_n1355_));
OR2X2 OR2X2_328 ( .A(_abc_4635_new_n1349_), .B(_abc_4635_new_n1356_), .Y(_abc_4635_new_n1357_));
OR2X2 OR2X2_329 ( .A(_abc_4635_new_n1358_), .B(W_R_1_bF_buf0_), .Y(_abc_4635_new_n1359_));
OR2X2 OR2X2_33 ( .A(_abc_4635_new_n475_), .B(\wordsize[0] ), .Y(_abc_4635_new_n494_));
OR2X2 OR2X2_330 ( .A(_abc_4635_new_n753__bF_buf3), .B(\pc[25] ), .Y(_abc_4635_new_n1360_));
OR2X2 OR2X2_331 ( .A(_abc_4635_new_n1356_), .B(_abc_4635_new_n1340_), .Y(_abc_4635_new_n1363_));
OR2X2 OR2X2_332 ( .A(_abc_4635_new_n1367_), .B(_abc_4635_new_n1365_), .Y(_abc_4635_new_n1368_));
OR2X2 OR2X2_333 ( .A(\imm[26] ), .B(\rs1[26] ), .Y(_abc_4635_new_n1371_));
OR2X2 OR2X2_334 ( .A(_abc_4635_new_n1368_), .B(_abc_4635_new_n1372_), .Y(_abc_4635_new_n1373_));
OR2X2 OR2X2_335 ( .A(_abc_4635_new_n1377_), .B(_abc_4635_new_n1362_), .Y(_auto_iopadmap_cc_368_execute_5767_26_));
OR2X2 OR2X2_336 ( .A(_abc_4635_new_n753__bF_buf1), .B(\pc[27] ), .Y(_abc_4635_new_n1379_));
OR2X2 OR2X2_337 ( .A(\imm[27] ), .B(\rs1[27] ), .Y(_abc_4635_new_n1381_));
OR2X2 OR2X2_338 ( .A(_abc_4635_new_n1380_), .B(_abc_4635_new_n1385_), .Y(_abc_4635_new_n1386_));
OR2X2 OR2X2_339 ( .A(_abc_4635_new_n1387_), .B(_abc_4635_new_n1384_), .Y(_abc_4635_new_n1388_));
OR2X2 OR2X2_34 ( .A(_abc_4635_new_n495_), .B(\wordsize[1] ), .Y(_abc_4635_new_n496_));
OR2X2 OR2X2_340 ( .A(_abc_4635_new_n1389_), .B(W_R_1_bF_buf4_), .Y(_abc_4635_new_n1390_));
OR2X2 OR2X2_341 ( .A(_abc_4635_new_n1397_), .B(_abc_4635_new_n1382_), .Y(_abc_4635_new_n1398_));
OR2X2 OR2X2_342 ( .A(_abc_4635_new_n1396_), .B(_abc_4635_new_n1398_), .Y(_abc_4635_new_n1399_));
OR2X2 OR2X2_343 ( .A(_abc_4635_new_n1395_), .B(_abc_4635_new_n1399_), .Y(_abc_4635_new_n1400_));
OR2X2 OR2X2_344 ( .A(\imm[28] ), .B(\rs1[28] ), .Y(_abc_4635_new_n1401_));
OR2X2 OR2X2_345 ( .A(_abc_4635_new_n1400_), .B(_abc_4635_new_n1404_), .Y(_abc_4635_new_n1405_));
OR2X2 OR2X2_346 ( .A(_abc_4635_new_n1409_), .B(_abc_4635_new_n1392_), .Y(_auto_iopadmap_cc_368_execute_5767_28_));
OR2X2 OR2X2_347 ( .A(\imm[29] ), .B(\rs1[29] ), .Y(_abc_4635_new_n1413_));
OR2X2 OR2X2_348 ( .A(_abc_4635_new_n1412_), .B(_abc_4635_new_n1416_), .Y(_abc_4635_new_n1417_));
OR2X2 OR2X2_349 ( .A(_abc_4635_new_n1411_), .B(_abc_4635_new_n1418_), .Y(_abc_4635_new_n1419_));
OR2X2 OR2X2_35 ( .A(_abc_4635_new_n498_), .B(\wordsize[1] ), .Y(_abc_4635_new_n499_));
OR2X2 OR2X2_350 ( .A(_abc_4635_new_n1420_), .B(W_R_1_bF_buf2_), .Y(_abc_4635_new_n1421_));
OR2X2 OR2X2_351 ( .A(_abc_4635_new_n753__bF_buf4), .B(\pc[29] ), .Y(_abc_4635_new_n1422_));
OR2X2 OR2X2_352 ( .A(_abc_4635_new_n1427_), .B(_abc_4635_new_n1414_), .Y(_abc_4635_new_n1428_));
OR2X2 OR2X2_353 ( .A(_abc_4635_new_n1426_), .B(_abc_4635_new_n1428_), .Y(_abc_4635_new_n1429_));
OR2X2 OR2X2_354 ( .A(\imm[30] ), .B(\rs1[30] ), .Y(_abc_4635_new_n1430_));
OR2X2 OR2X2_355 ( .A(_abc_4635_new_n1429_), .B(_abc_4635_new_n1433_), .Y(_abc_4635_new_n1434_));
OR2X2 OR2X2_356 ( .A(_abc_4635_new_n470_), .B(_abc_4635_new_n466_), .Y(_abc_4635_new_n1435_));
OR2X2 OR2X2_357 ( .A(_abc_4635_new_n1436_), .B(_abc_4635_new_n1437_), .Y(_abc_4635_new_n1438_));
OR2X2 OR2X2_358 ( .A(_abc_4635_new_n1440_), .B(_abc_4635_new_n1441_), .Y(_abc_4635_new_n1442_));
OR2X2 OR2X2_359 ( .A(_abc_4635_new_n1444_), .B(_abc_4635_new_n1445_), .Y(_abc_4635_new_n1446_));
OR2X2 OR2X2_36 ( .A(_abc_4635_new_n480__bF_buf3), .B(_abc_4635_new_n511__bF_buf6), .Y(_abc_4635_new_n512_));
OR2X2 OR2X2_360 ( .A(_abc_4635_new_n1448_), .B(_abc_4635_new_n1449_), .Y(_abc_4635_new_n1450_));
OR2X2 OR2X2_361 ( .A(_abc_4635_new_n1452_), .B(_abc_4635_new_n1453_), .Y(_abc_4635_new_n1454_));
OR2X2 OR2X2_362 ( .A(_abc_4635_new_n1456_), .B(_abc_4635_new_n1457_), .Y(_abc_4635_new_n1458_));
OR2X2 OR2X2_363 ( .A(_abc_4635_new_n1460_), .B(_abc_4635_new_n1461_), .Y(_abc_4635_new_n1462_));
OR2X2 OR2X2_364 ( .A(_abc_4635_new_n1464_), .B(_abc_4635_new_n1424_), .Y(_auto_iopadmap_cc_368_execute_5767_30_));
OR2X2 OR2X2_365 ( .A(_abc_4635_new_n1466_), .B(_abc_4635_new_n1431_), .Y(_abc_4635_new_n1467_));
OR2X2 OR2X2_366 ( .A(_abc_4635_new_n1468_), .B(\rs1[31] ), .Y(_abc_4635_new_n1469_));
OR2X2 OR2X2_367 ( .A(_abc_4635_new_n1470_), .B(\imm[31] ), .Y(_abc_4635_new_n1471_));
OR2X2 OR2X2_368 ( .A(_abc_4635_new_n1467_), .B(_abc_4635_new_n1473_), .Y(_abc_4635_new_n1474_));
OR2X2 OR2X2_369 ( .A(_abc_4635_new_n1475_), .B(_abc_4635_new_n1472_), .Y(_abc_4635_new_n1476_));
OR2X2 OR2X2_37 ( .A(_abc_4635_new_n513_), .B(_abc_4635_new_n510_), .Y(_abc_4635_new_n514_));
OR2X2 OR2X2_370 ( .A(_abc_4635_new_n1477_), .B(W_R_1_bF_buf0_), .Y(_abc_4635_new_n1478_));
OR2X2 OR2X2_371 ( .A(_abc_4635_new_n753__bF_buf2), .B(\pc[31] ), .Y(_abc_4635_new_n1479_));
OR2X2 OR2X2_372 ( .A(state_6_), .B(state_1_), .Y(_abc_4635_new_n1482_));
OR2X2 OR2X2_373 ( .A(_abc_4635_new_n425_), .B(state_3_), .Y(_abc_4635_new_n1483_));
OR2X2 OR2X2_374 ( .A(_abc_4635_new_n1483_), .B(_abc_4635_new_n1482_), .Y(_abc_4635_new_n1484_));
OR2X2 OR2X2_375 ( .A(_abc_4635_new_n393_), .B(state_2_), .Y(_abc_4635_new_n1486_));
OR2X2 OR2X2_376 ( .A(_auto_iopadmap_cc_368_execute_5800), .B(_abc_4635_new_n429_), .Y(_auto_iopadmap_cc_368_execute_5839));
OR2X2 OR2X2_377 ( .A(_abc_4635_new_n426_), .B(_abc_4635_new_n397_), .Y(_auto_iopadmap_cc_368_execute_5835));
OR2X2 OR2X2_38 ( .A(_abc_4635_new_n518_), .B(_abc_4635_new_n517_), .Y(_abc_4635_new_n519_));
OR2X2 OR2X2_39 ( .A(_abc_4635_new_n523_), .B(_abc_4635_new_n522_), .Y(_abc_4635_new_n524_));
OR2X2 OR2X2_4 ( .A(_abc_4635_new_n384_), .B(_abc_4635_new_n372_), .Y(_abc_4635_new_n385_));
OR2X2 OR2X2_40 ( .A(_abc_4635_new_n528_), .B(_abc_4635_new_n527_), .Y(_abc_4635_new_n529_));
OR2X2 OR2X2_41 ( .A(_abc_4635_new_n533_), .B(_abc_4635_new_n532_), .Y(_abc_4635_new_n534_));
OR2X2 OR2X2_42 ( .A(_abc_4635_new_n538_), .B(_abc_4635_new_n537_), .Y(_abc_4635_new_n539_));
OR2X2 OR2X2_43 ( .A(_abc_4635_new_n543_), .B(_abc_4635_new_n542_), .Y(_abc_4635_new_n544_));
OR2X2 OR2X2_44 ( .A(_abc_4635_new_n548_), .B(_abc_4635_new_n547_), .Y(_abc_4635_new_n549_));
OR2X2 OR2X2_45 ( .A(_abc_4635_new_n551_), .B(_abc_4635_new_n509_), .Y(_abc_4635_new_n552_));
OR2X2 OR2X2_46 ( .A(_abc_4635_new_n554_), .B(_abc_4635_new_n516_), .Y(_abc_4635_new_n555_));
OR2X2 OR2X2_47 ( .A(_abc_4635_new_n557_), .B(_abc_4635_new_n521_), .Y(_abc_4635_new_n558_));
OR2X2 OR2X2_48 ( .A(_abc_4635_new_n560_), .B(_abc_4635_new_n526_), .Y(_abc_4635_new_n561_));
OR2X2 OR2X2_49 ( .A(_abc_4635_new_n563_), .B(_abc_4635_new_n531_), .Y(_abc_4635_new_n564_));
OR2X2 OR2X2_5 ( .A(_abc_4635_new_n386_), .B(_abc_4635_new_n366_), .Y(_abc_4635_new_n387_));
OR2X2 OR2X2_50 ( .A(_abc_4635_new_n566_), .B(_abc_4635_new_n536_), .Y(_abc_4635_new_n567_));
OR2X2 OR2X2_51 ( .A(_abc_4635_new_n569_), .B(_abc_4635_new_n541_), .Y(_abc_4635_new_n570_));
OR2X2 OR2X2_52 ( .A(_abc_4635_new_n572_), .B(_abc_4635_new_n546_), .Y(_abc_4635_new_n573_));
OR2X2 OR2X2_53 ( .A(_abc_4635_new_n510_), .B(_abc_4635_new_n575_), .Y(_abc_4635_new_n576_));
OR2X2 OR2X2_54 ( .A(_abc_4635_new_n576_), .B(_abc_4635_new_n577_), .Y(_abc_4635_new_n578_));
OR2X2 OR2X2_55 ( .A(_abc_4635_new_n517_), .B(_abc_4635_new_n580_), .Y(_abc_4635_new_n581_));
OR2X2 OR2X2_56 ( .A(_abc_4635_new_n581_), .B(_abc_4635_new_n582_), .Y(_abc_4635_new_n583_));
OR2X2 OR2X2_57 ( .A(_abc_4635_new_n522_), .B(_abc_4635_new_n585_), .Y(_abc_4635_new_n586_));
OR2X2 OR2X2_58 ( .A(_abc_4635_new_n586_), .B(_abc_4635_new_n587_), .Y(_abc_4635_new_n588_));
OR2X2 OR2X2_59 ( .A(_abc_4635_new_n527_), .B(_abc_4635_new_n590_), .Y(_abc_4635_new_n591_));
OR2X2 OR2X2_6 ( .A(_abc_4635_new_n392_), .B(_abc_4635_new_n393_), .Y(_abc_4635_new_n394_));
OR2X2 OR2X2_60 ( .A(_abc_4635_new_n591_), .B(_abc_4635_new_n592_), .Y(_abc_4635_new_n593_));
OR2X2 OR2X2_61 ( .A(_abc_4635_new_n532_), .B(_abc_4635_new_n595_), .Y(_abc_4635_new_n596_));
OR2X2 OR2X2_62 ( .A(_abc_4635_new_n596_), .B(_abc_4635_new_n597_), .Y(_abc_4635_new_n598_));
OR2X2 OR2X2_63 ( .A(_abc_4635_new_n537_), .B(_abc_4635_new_n600_), .Y(_abc_4635_new_n601_));
OR2X2 OR2X2_64 ( .A(_abc_4635_new_n601_), .B(_abc_4635_new_n602_), .Y(_abc_4635_new_n603_));
OR2X2 OR2X2_65 ( .A(_abc_4635_new_n542_), .B(_abc_4635_new_n605_), .Y(_abc_4635_new_n606_));
OR2X2 OR2X2_66 ( .A(_abc_4635_new_n606_), .B(_abc_4635_new_n607_), .Y(_abc_4635_new_n608_));
OR2X2 OR2X2_67 ( .A(_abc_4635_new_n547_), .B(_abc_4635_new_n610_), .Y(_abc_4635_new_n611_));
OR2X2 OR2X2_68 ( .A(_abc_4635_new_n611_), .B(_abc_4635_new_n612_), .Y(_abc_4635_new_n613_));
OR2X2 OR2X2_69 ( .A(_abc_4635_new_n619_), .B(_abc_4635_new_n617_), .Y(_abc_4635_new_n620_));
OR2X2 OR2X2_7 ( .A(_abc_4635_new_n398_), .B(_abc_4635_new_n397_), .Y(_abc_4635_new_n399_));
OR2X2 OR2X2_70 ( .A(_abc_4635_new_n623_), .B(_abc_4635_new_n622_), .Y(_abc_4635_new_n624_));
OR2X2 OR2X2_71 ( .A(_abc_4635_new_n627_), .B(_abc_4635_new_n626_), .Y(_abc_4635_new_n628_));
OR2X2 OR2X2_72 ( .A(_abc_4635_new_n631_), .B(_abc_4635_new_n630_), .Y(_abc_4635_new_n632_));
OR2X2 OR2X2_73 ( .A(_abc_4635_new_n635_), .B(_abc_4635_new_n634_), .Y(_abc_4635_new_n636_));
OR2X2 OR2X2_74 ( .A(_abc_4635_new_n639_), .B(_abc_4635_new_n638_), .Y(_abc_4635_new_n640_));
OR2X2 OR2X2_75 ( .A(_abc_4635_new_n643_), .B(_abc_4635_new_n642_), .Y(_abc_4635_new_n644_));
OR2X2 OR2X2_76 ( .A(_abc_4635_new_n647_), .B(_abc_4635_new_n646_), .Y(_abc_4635_new_n648_));
OR2X2 OR2X2_77 ( .A(_abc_4635_new_n651_), .B(_abc_4635_new_n650_), .Y(_abc_4635_new_n652_));
OR2X2 OR2X2_78 ( .A(_abc_4635_new_n655_), .B(_abc_4635_new_n654_), .Y(_abc_4635_new_n656_));
OR2X2 OR2X2_79 ( .A(_abc_4635_new_n659_), .B(_abc_4635_new_n658_), .Y(_abc_4635_new_n660_));
OR2X2 OR2X2_8 ( .A(_abc_4635_new_n404_), .B(_abc_4635_new_n401_), .Y(_abc_4635_new_n405_));
OR2X2 OR2X2_80 ( .A(_abc_4635_new_n663_), .B(_abc_4635_new_n662_), .Y(_abc_4635_new_n664_));
OR2X2 OR2X2_81 ( .A(_abc_4635_new_n667_), .B(_abc_4635_new_n666_), .Y(_abc_4635_new_n668_));
OR2X2 OR2X2_82 ( .A(_abc_4635_new_n671_), .B(_abc_4635_new_n670_), .Y(_abc_4635_new_n672_));
OR2X2 OR2X2_83 ( .A(_abc_4635_new_n675_), .B(_abc_4635_new_n674_), .Y(_abc_4635_new_n676_));
OR2X2 OR2X2_84 ( .A(_abc_4635_new_n679_), .B(_abc_4635_new_n678_), .Y(_abc_4635_new_n680_));
OR2X2 OR2X2_85 ( .A(_abc_4635_new_n683_), .B(_abc_4635_new_n682_), .Y(_abc_4635_new_n684_));
OR2X2 OR2X2_86 ( .A(_abc_4635_new_n687_), .B(_abc_4635_new_n686_), .Y(_abc_4635_new_n688_));
OR2X2 OR2X2_87 ( .A(_abc_4635_new_n691_), .B(_abc_4635_new_n690_), .Y(_abc_4635_new_n692_));
OR2X2 OR2X2_88 ( .A(_abc_4635_new_n695_), .B(_abc_4635_new_n694_), .Y(_abc_4635_new_n696_));
OR2X2 OR2X2_89 ( .A(_abc_4635_new_n699_), .B(_abc_4635_new_n698_), .Y(_abc_4635_new_n700_));
OR2X2 OR2X2_9 ( .A(_abc_4635_new_n408_), .B(_abc_4635_new_n409_), .Y(_abc_4635_new_n410_));
OR2X2 OR2X2_90 ( .A(_abc_4635_new_n703_), .B(_abc_4635_new_n702_), .Y(_abc_4635_new_n704_));
OR2X2 OR2X2_91 ( .A(_abc_4635_new_n707_), .B(_abc_4635_new_n706_), .Y(_abc_4635_new_n708_));
OR2X2 OR2X2_92 ( .A(_abc_4635_new_n711_), .B(_abc_4635_new_n710_), .Y(_abc_4635_new_n712_));
OR2X2 OR2X2_93 ( .A(_abc_4635_new_n715_), .B(_abc_4635_new_n714_), .Y(_abc_4635_new_n716_));
OR2X2 OR2X2_94 ( .A(_abc_4635_new_n719_), .B(_abc_4635_new_n718_), .Y(_abc_4635_new_n720_));
OR2X2 OR2X2_95 ( .A(_abc_4635_new_n723_), .B(_abc_4635_new_n722_), .Y(_abc_4635_new_n724_));
OR2X2 OR2X2_96 ( .A(_abc_4635_new_n727_), .B(_abc_4635_new_n726_), .Y(_abc_4635_new_n728_));
OR2X2 OR2X2_97 ( .A(_abc_4635_new_n731_), .B(_abc_4635_new_n730_), .Y(_abc_4635_new_n732_));
OR2X2 OR2X2_98 ( .A(_abc_4635_new_n735_), .B(_abc_4635_new_n734_), .Y(_abc_4635_new_n736_));
OR2X2 OR2X2_99 ( .A(_abc_4635_new_n739_), .B(_abc_4635_new_n738_), .Y(_abc_4635_new_n740_));


endmodule