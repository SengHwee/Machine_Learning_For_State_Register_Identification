module MEMORY_INTERFACE(clock, resetn, \rs1[0] , \rs1[1] , \rs1[2] , \rs1[3] , \rs1[4] , \rs1[5] , \rs1[6] , \rs1[7] , \rs1[8] , \rs1[9] , \rs1[10] , \rs1[11] , \rs1[12] , \rs1[13] , \rs1[14] , \rs1[15] , \rs1[16] , \rs1[17] , \rs1[18] , \rs1[19] , \rs1[20] , \rs1[21] , \rs1[22] , \rs1[23] , \rs1[24] , \rs1[25] , \rs1[26] , \rs1[27] , \rs1[28] , \rs1[29] , \rs1[30] , \rs1[31] , \rs2[0] , \rs2[1] , \rs2[2] , \rs2[3] , \rs2[4] , \rs2[5] , \rs2[6] , \rs2[7] , \rs2[8] , \rs2[9] , \rs2[10] , \rs2[11] , \rs2[12] , \rs2[13] , \rs2[14] , \rs2[15] , \rs2[16] , \rs2[17] , \rs2[18] , \rs2[19] , \rs2[20] , \rs2[21] , \rs2[22] , \rs2[23] , \rs2[24] , \rs2[25] , \rs2[26] , \rs2[27] , \rs2[28] , \rs2[29] , \rs2[30] , \rs2[31] , \Rdata_mem[0] , \Rdata_mem[1] , \Rdata_mem[2] , \Rdata_mem[3] , \Rdata_mem[4] , \Rdata_mem[5] , \Rdata_mem[6] , \Rdata_mem[7] , \Rdata_mem[8] , \Rdata_mem[9] , \Rdata_mem[10] , \Rdata_mem[11] , \Rdata_mem[12] , \Rdata_mem[13] , \Rdata_mem[14] , \Rdata_mem[15] , \Rdata_mem[16] , \Rdata_mem[17] , \Rdata_mem[18] , \Rdata_mem[19] , \Rdata_mem[20] , \Rdata_mem[21] , \Rdata_mem[22] , \Rdata_mem[23] , \Rdata_mem[24] , \Rdata_mem[25] , \Rdata_mem[26] , \Rdata_mem[27] , \Rdata_mem[28] , \Rdata_mem[29] , \Rdata_mem[30] , \Rdata_mem[31] , ARready, Rvalid, AWready, Wready, Bvalid, \imm[0] , \imm[1] , \imm[2] , \imm[3] , \imm[4] , \imm[5] , \imm[6] , \imm[7] , \imm[8] , \imm[9] , \imm[10] , \imm[11] , \imm[12] , \imm[13] , \imm[14] , \imm[15] , \imm[16] , \imm[17] , \imm[18] , \imm[19] , \imm[20] , \imm[21] , \imm[22] , \imm[23] , \imm[24] , \imm[25] , \imm[26] , \imm[27] , \imm[28] , \imm[29] , \imm[30] , \imm[31] , \W_R[0] , \W_R[1] , \wordsize[0] , \wordsize[1] , enable, \pc[0] , \pc[1] , \pc[2] , \pc[3] , \pc[4] , \pc[5] , \pc[6] , \pc[7] , \pc[8] , \pc[9] , \pc[10] , \pc[11] , \pc[12] , \pc[13] , \pc[14] , \pc[15] , \pc[16] , \pc[17] , \pc[18] , \pc[19] , \pc[20] , \pc[21] , \pc[22] , \pc[23] , \pc[24] , \pc[25] , \pc[26] , \pc[27] , \pc[28] , \pc[29] , \pc[30] , \pc[31] , signo, busy, done, align, \AWdata[0] , \AWdata[1] , \AWdata[2] , \AWdata[3] , \AWdata[4] , \AWdata[5] , \AWdata[6] , \AWdata[7] , \AWdata[8] , \AWdata[9] , \AWdata[10] , \AWdata[11] , \AWdata[12] , \AWdata[13] , \AWdata[14] , \AWdata[15] , \AWdata[16] , \AWdata[17] , \AWdata[18] , \AWdata[19] , \AWdata[20] , \AWdata[21] , \AWdata[22] , \AWdata[23] , \AWdata[24] , \AWdata[25] , \AWdata[26] , \AWdata[27] , \AWdata[28] , \AWdata[29] , \AWdata[30] , \AWdata[31] , \ARdata[0] , \ARdata[1] , \ARdata[2] , \ARdata[3] , \ARdata[4] , \ARdata[5] , \ARdata[6] , \ARdata[7] , \ARdata[8] , \ARdata[9] , \ARdata[10] , \ARdata[11] , \ARdata[12] , \ARdata[13] , \ARdata[14] , \ARdata[15] , \ARdata[16] , \ARdata[17] , \ARdata[18] , \ARdata[19] , \ARdata[20] , \ARdata[21] , \ARdata[22] , \ARdata[23] , \ARdata[24] , \ARdata[25] , \ARdata[26] , \ARdata[27] , \ARdata[28] , \ARdata[29] , \ARdata[30] , \ARdata[31] , \Wdata[0] , \Wdata[1] , \Wdata[2] , \Wdata[3] , \Wdata[4] , \Wdata[5] , \Wdata[6] , \Wdata[7] , \Wdata[8] , \Wdata[9] , \Wdata[10] , \Wdata[11] , \Wdata[12] , \Wdata[13] , \Wdata[14] , \Wdata[15] , \Wdata[16] , \Wdata[17] , \Wdata[18] , \Wdata[19] , \Wdata[20] , \Wdata[21] , \Wdata[22] , \Wdata[23] , \Wdata[24] , \Wdata[25] , \Wdata[26] , \Wdata[27] , \Wdata[28] , \Wdata[29] , \Wdata[30] , \Wdata[31] , \rd[0] , \rd[1] , \rd[2] , \rd[3] , \rd[4] , \rd[5] , \rd[6] , \rd[7] , \rd[8] , \rd[9] , \rd[10] , \rd[11] , \rd[12] , \rd[13] , \rd[14] , \rd[15] , \rd[16] , \rd[17] , \rd[18] , \rd[19] , \rd[20] , \rd[21] , \rd[22] , \rd[23] , \rd[24] , \rd[25] , \rd[26] , \rd[27] , \rd[28] , \rd[29] , \rd[30] , \rd[31] , \inst[0] , \inst[1] , \inst[2] , \inst[3] , \inst[4] , \inst[5] , \inst[6] , \inst[7] , \inst[8] , \inst[9] , \inst[10] , \inst[11] , \inst[12] , \inst[13] , \inst[14] , \inst[15] , \inst[16] , \inst[17] , \inst[18] , \inst[19] , \inst[20] , \inst[21] , \inst[22] , \inst[23] , \inst[24] , \inst[25] , \inst[26] , \inst[27] , \inst[28] , \inst[29] , \inst[30] , \inst[31] , ARvalid, RReady, AWvalid, Wvalid, \arprot[0] , \arprot[1] , \arprot[2] , \awprot[0] , \awprot[1] , \awprot[2] , Bready, \Wstrb[0] , \Wstrb[1] , \Wstrb[2] , \Wstrb[3] , rd_en);

output \ARdata[0] ;
output \ARdata[10] ;
output \ARdata[11] ;
output \ARdata[12] ;
output \ARdata[13] ;
output \ARdata[14] ;
output \ARdata[15] ;
output \ARdata[16] ;
output \ARdata[17] ;
output \ARdata[18] ;
output \ARdata[19] ;
output \ARdata[1] ;
output \ARdata[20] ;
output \ARdata[21] ;
output \ARdata[22] ;
output \ARdata[23] ;
output \ARdata[24] ;
output \ARdata[25] ;
output \ARdata[26] ;
output \ARdata[27] ;
output \ARdata[28] ;
output \ARdata[29] ;
output \ARdata[2] ;
output \ARdata[30] ;
output \ARdata[31] ;
output \ARdata[3] ;
output \ARdata[4] ;
output \ARdata[5] ;
output \ARdata[6] ;
output \ARdata[7] ;
output \ARdata[8] ;
output \ARdata[9] ;
input ARready;
output ARvalid;
output \AWdata[0] ;
output \AWdata[10] ;
output \AWdata[11] ;
output \AWdata[12] ;
output \AWdata[13] ;
output \AWdata[14] ;
output \AWdata[15] ;
output \AWdata[16] ;
output \AWdata[17] ;
output \AWdata[18] ;
output \AWdata[19] ;
output \AWdata[1] ;
output \AWdata[20] ;
output \AWdata[21] ;
output \AWdata[22] ;
output \AWdata[23] ;
output \AWdata[24] ;
output \AWdata[25] ;
output \AWdata[26] ;
output \AWdata[27] ;
output \AWdata[28] ;
output \AWdata[29] ;
output \AWdata[2] ;
output \AWdata[30] ;
output \AWdata[31] ;
output \AWdata[3] ;
output \AWdata[4] ;
output \AWdata[5] ;
output \AWdata[6] ;
output \AWdata[7] ;
output \AWdata[8] ;
output \AWdata[9] ;
input AWready;
output AWvalid;
output Bready;
input Bvalid;
output RReady;
input \Rdata_mem[0] ;
input \Rdata_mem[10] ;
input \Rdata_mem[11] ;
input \Rdata_mem[12] ;
input \Rdata_mem[13] ;
input \Rdata_mem[14] ;
input \Rdata_mem[15] ;
input \Rdata_mem[16] ;
input \Rdata_mem[17] ;
input \Rdata_mem[18] ;
input \Rdata_mem[19] ;
input \Rdata_mem[1] ;
input \Rdata_mem[20] ;
input \Rdata_mem[21] ;
input \Rdata_mem[22] ;
input \Rdata_mem[23] ;
input \Rdata_mem[24] ;
input \Rdata_mem[25] ;
input \Rdata_mem[26] ;
input \Rdata_mem[27] ;
input \Rdata_mem[28] ;
input \Rdata_mem[29] ;
input \Rdata_mem[2] ;
input \Rdata_mem[30] ;
input \Rdata_mem[31] ;
input \Rdata_mem[3] ;
input \Rdata_mem[4] ;
input \Rdata_mem[5] ;
input \Rdata_mem[6] ;
input \Rdata_mem[7] ;
input \Rdata_mem[8] ;
input \Rdata_mem[9] ;
input Rvalid;
input \W_R[0] ;
input \W_R[1] ;
output \Wdata[0] ;
output \Wdata[10] ;
output \Wdata[11] ;
output \Wdata[12] ;
output \Wdata[13] ;
output \Wdata[14] ;
output \Wdata[15] ;
output \Wdata[16] ;
output \Wdata[17] ;
output \Wdata[18] ;
output \Wdata[19] ;
output \Wdata[1] ;
output \Wdata[20] ;
output \Wdata[21] ;
output \Wdata[22] ;
output \Wdata[23] ;
output \Wdata[24] ;
output \Wdata[25] ;
output \Wdata[26] ;
output \Wdata[27] ;
output \Wdata[28] ;
output \Wdata[29] ;
output \Wdata[2] ;
output \Wdata[30] ;
output \Wdata[31] ;
output \Wdata[3] ;
output \Wdata[4] ;
output \Wdata[5] ;
output \Wdata[6] ;
output \Wdata[7] ;
output \Wdata[8] ;
output \Wdata[9] ;
input Wready;
output \Wstrb[0] ;
output \Wstrb[1] ;
output \Wstrb[2] ;
output \Wstrb[3] ;
output Wvalid;
wire _0Wdata_31_0__0_; 
wire _0Wdata_31_0__10_; 
wire _0Wdata_31_0__11_; 
wire _0Wdata_31_0__12_; 
wire _0Wdata_31_0__13_; 
wire _0Wdata_31_0__14_; 
wire _0Wdata_31_0__15_; 
wire _0Wdata_31_0__16_; 
wire _0Wdata_31_0__17_; 
wire _0Wdata_31_0__18_; 
wire _0Wdata_31_0__19_; 
wire _0Wdata_31_0__1_; 
wire _0Wdata_31_0__20_; 
wire _0Wdata_31_0__21_; 
wire _0Wdata_31_0__22_; 
wire _0Wdata_31_0__23_; 
wire _0Wdata_31_0__24_; 
wire _0Wdata_31_0__25_; 
wire _0Wdata_31_0__26_; 
wire _0Wdata_31_0__27_; 
wire _0Wdata_31_0__28_; 
wire _0Wdata_31_0__29_; 
wire _0Wdata_31_0__2_; 
wire _0Wdata_31_0__30_; 
wire _0Wdata_31_0__31_; 
wire _0Wdata_31_0__3_; 
wire _0Wdata_31_0__4_; 
wire _0Wdata_31_0__5_; 
wire _0Wdata_31_0__6_; 
wire _0Wdata_31_0__7_; 
wire _0Wdata_31_0__8_; 
wire _0Wdata_31_0__9_; 
wire _0Wstrb_3_0__0_; 
wire _0Wstrb_3_0__1_; 
wire _0Wstrb_3_0__2_; 
wire _0Wstrb_3_0__3_; 
wire _0inst_31_0__0_; 
wire _0inst_31_0__10_; 
wire _0inst_31_0__11_; 
wire _0inst_31_0__12_; 
wire _0inst_31_0__13_; 
wire _0inst_31_0__14_; 
wire _0inst_31_0__15_; 
wire _0inst_31_0__16_; 
wire _0inst_31_0__17_; 
wire _0inst_31_0__18_; 
wire _0inst_31_0__19_; 
wire _0inst_31_0__1_; 
wire _0inst_31_0__20_; 
wire _0inst_31_0__21_; 
wire _0inst_31_0__22_; 
wire _0inst_31_0__23_; 
wire _0inst_31_0__24_; 
wire _0inst_31_0__25_; 
wire _0inst_31_0__26_; 
wire _0inst_31_0__27_; 
wire _0inst_31_0__28_; 
wire _0inst_31_0__29_; 
wire _0inst_31_0__2_; 
wire _0inst_31_0__30_; 
wire _0inst_31_0__31_; 
wire _0inst_31_0__3_; 
wire _0inst_31_0__4_; 
wire _0inst_31_0__5_; 
wire _0inst_31_0__6_; 
wire _0inst_31_0__7_; 
wire _0inst_31_0__8_; 
wire _0inst_31_0__9_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_0_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_1_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_2_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_3_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_4_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_5_; 
wire _abc_3813_auto_fsm_map_cc_170_map_fsm_1372_6_; 
wire _abc_4635_new_n1000_; 
wire _abc_4635_new_n1001_; 
wire _abc_4635_new_n1003_; 
wire _abc_4635_new_n1004_; 
wire _abc_4635_new_n1005_; 
wire _abc_4635_new_n1006_; 
wire _abc_4635_new_n1007_; 
wire _abc_4635_new_n1008_; 
wire _abc_4635_new_n1009_; 
wire _abc_4635_new_n1010_; 
wire _abc_4635_new_n1012_; 
wire _abc_4635_new_n1013_; 
wire _abc_4635_new_n1014_; 
wire _abc_4635_new_n1015_; 
wire _abc_4635_new_n1016_; 
wire _abc_4635_new_n1017_; 
wire _abc_4635_new_n1018_; 
wire _abc_4635_new_n1019_; 
wire _abc_4635_new_n1020_; 
wire _abc_4635_new_n1021_; 
wire _abc_4635_new_n1022_; 
wire _abc_4635_new_n1023_; 
wire _abc_4635_new_n1024_; 
wire _abc_4635_new_n1025_; 
wire _abc_4635_new_n1026_; 
wire _abc_4635_new_n1027_; 
wire _abc_4635_new_n1028_; 
wire _abc_4635_new_n1029_; 
wire _abc_4635_new_n1030_; 
wire _abc_4635_new_n1031_; 
wire _abc_4635_new_n1032_; 
wire _abc_4635_new_n1033_; 
wire _abc_4635_new_n1034_; 
wire _abc_4635_new_n1036_; 
wire _abc_4635_new_n1037_; 
wire _abc_4635_new_n1038_; 
wire _abc_4635_new_n1039_; 
wire _abc_4635_new_n1040_; 
wire _abc_4635_new_n1041_; 
wire _abc_4635_new_n1043_; 
wire _abc_4635_new_n1044_; 
wire _abc_4635_new_n1045_; 
wire _abc_4635_new_n1046_; 
wire _abc_4635_new_n1047_; 
wire _abc_4635_new_n1048_; 
wire _abc_4635_new_n1049_; 
wire _abc_4635_new_n1050_; 
wire _abc_4635_new_n1051_; 
wire _abc_4635_new_n1052_; 
wire _abc_4635_new_n1053_; 
wire _abc_4635_new_n1054_; 
wire _abc_4635_new_n1056_; 
wire _abc_4635_new_n1057_; 
wire _abc_4635_new_n1058_; 
wire _abc_4635_new_n1059_; 
wire _abc_4635_new_n1060_; 
wire _abc_4635_new_n1061_; 
wire _abc_4635_new_n1062_; 
wire _abc_4635_new_n1064_; 
wire _abc_4635_new_n1065_; 
wire _abc_4635_new_n1066_; 
wire _abc_4635_new_n1067_; 
wire _abc_4635_new_n1068_; 
wire _abc_4635_new_n1069_; 
wire _abc_4635_new_n1070_; 
wire _abc_4635_new_n1071_; 
wire _abc_4635_new_n1072_; 
wire _abc_4635_new_n1073_; 
wire _abc_4635_new_n1074_; 
wire _abc_4635_new_n1075_; 
wire _abc_4635_new_n1076_; 
wire _abc_4635_new_n1077_; 
wire _abc_4635_new_n1078_; 
wire _abc_4635_new_n1079_; 
wire _abc_4635_new_n1080_; 
wire _abc_4635_new_n1082_; 
wire _abc_4635_new_n1083_; 
wire _abc_4635_new_n1084_; 
wire _abc_4635_new_n1085_; 
wire _abc_4635_new_n1086_; 
wire _abc_4635_new_n1087_; 
wire _abc_4635_new_n1088_; 
wire _abc_4635_new_n1090_; 
wire _abc_4635_new_n1091_; 
wire _abc_4635_new_n1092_; 
wire _abc_4635_new_n1093_; 
wire _abc_4635_new_n1094_; 
wire _abc_4635_new_n1095_; 
wire _abc_4635_new_n1096_; 
wire _abc_4635_new_n1097_; 
wire _abc_4635_new_n1098_; 
wire _abc_4635_new_n1099_; 
wire _abc_4635_new_n1100_; 
wire _abc_4635_new_n1101_; 
wire _abc_4635_new_n1102_; 
wire _abc_4635_new_n1103_; 
wire _abc_4635_new_n1104_; 
wire _abc_4635_new_n1106_; 
wire _abc_4635_new_n1107_; 
wire _abc_4635_new_n1108_; 
wire _abc_4635_new_n1109_; 
wire _abc_4635_new_n1110_; 
wire _abc_4635_new_n1111_; 
wire _abc_4635_new_n1112_; 
wire _abc_4635_new_n1115_; 
wire _abc_4635_new_n1116_; 
wire _abc_4635_new_n1117_; 
wire _abc_4635_new_n1119_; 
wire _abc_4635_new_n361_; 
wire _abc_4635_new_n362_; 
wire _abc_4635_new_n363_; 
wire _abc_4635_new_n364_; 
wire _abc_4635_new_n365_; 
wire _abc_4635_new_n366_; 
wire _abc_4635_new_n367_; 
wire _abc_4635_new_n368_; 
wire _abc_4635_new_n369_; 
wire _abc_4635_new_n370_; 
wire _abc_4635_new_n371_; 
wire _abc_4635_new_n372_; 
wire _abc_4635_new_n373_; 
wire _abc_4635_new_n374_; 
wire _abc_4635_new_n375_; 
wire _abc_4635_new_n376_; 
wire _abc_4635_new_n377_; 
wire _abc_4635_new_n378_; 
wire _abc_4635_new_n379_; 
wire _abc_4635_new_n380_; 
wire _abc_4635_new_n382_; 
wire _abc_4635_new_n383_; 
wire _abc_4635_new_n384_; 
wire _abc_4635_new_n385_; 
wire _abc_4635_new_n386_; 
wire _abc_4635_new_n387_; 
wire _abc_4635_new_n388_; 
wire _abc_4635_new_n389_; 
wire _abc_4635_new_n390_; 
wire _abc_4635_new_n392_; 
wire _abc_4635_new_n393_; 
wire _abc_4635_new_n395_; 
wire _abc_4635_new_n396_; 
wire _abc_4635_new_n397_; 
wire _abc_4635_new_n398_; 
wire _abc_4635_new_n399_; 
wire _abc_4635_new_n400_; 
wire _abc_4635_new_n401_; 
wire _abc_4635_new_n402_; 
wire _abc_4635_new_n403_; 
wire _abc_4635_new_n404_; 
wire _abc_4635_new_n405_; 
wire _abc_4635_new_n406_; 
wire _abc_4635_new_n408_; 
wire _abc_4635_new_n409_; 
wire _abc_4635_new_n410_; 
wire _abc_4635_new_n412_; 
wire _abc_4635_new_n413_; 
wire _abc_4635_new_n415_; 
wire _abc_4635_new_n416_; 
wire _abc_4635_new_n418_; 
wire _abc_4635_new_n419_; 
wire _abc_4635_new_n420_; 
wire _abc_4635_new_n421_; 
wire _abc_4635_new_n422_; 
wire _abc_4635_new_n423_; 
wire _abc_4635_new_n424_; 
wire _abc_4635_new_n425_; 
wire _abc_4635_new_n426_; 
wire _abc_4635_new_n427_; 
wire _abc_4635_new_n428_; 
wire _abc_4635_new_n429_; 
wire _abc_4635_new_n432_; 
wire _abc_4635_new_n433_; 
wire _abc_4635_new_n434_; 
wire _abc_4635_new_n435_; 
wire _abc_4635_new_n436_; 
wire _abc_4635_new_n437_; 
wire _abc_4635_new_n438_; 
wire _abc_4635_new_n439_; 
wire _abc_4635_new_n440_; 
wire _abc_4635_new_n441_; 
wire _abc_4635_new_n442_; 
wire _abc_4635_new_n443_; 
wire _abc_4635_new_n444_; 
wire _abc_4635_new_n445_; 
wire _abc_4635_new_n446_; 
wire _abc_4635_new_n447_; 
wire _abc_4635_new_n448_; 
wire _abc_4635_new_n449_; 
wire _abc_4635_new_n450_; 
wire _abc_4635_new_n451_; 
wire _abc_4635_new_n453_; 
wire _abc_4635_new_n454_; 
wire _abc_4635_new_n456_; 
wire _abc_4635_new_n457_; 
wire _abc_4635_new_n458_; 
wire _abc_4635_new_n460_; 
wire _abc_4635_new_n462_; 
wire _abc_4635_new_n464_; 
wire _abc_4635_new_n466_; 
wire _abc_4635_new_n468_; 
wire _abc_4635_new_n470_; 
wire _abc_4635_new_n472_; 
wire _abc_4635_new_n474_; 
wire _abc_4635_new_n476_; 
wire _abc_4635_new_n478_; 
wire _abc_4635_new_n479_; 
wire _abc_4635_new_n480_; 
wire _abc_4635_new_n481_; 
wire _abc_4635_new_n483_; 
wire _abc_4635_new_n484_; 
wire _abc_4635_new_n486_; 
wire _abc_4635_new_n487_; 
wire _abc_4635_new_n489_; 
wire _abc_4635_new_n490_; 
wire _abc_4635_new_n492_; 
wire _abc_4635_new_n493_; 
wire _abc_4635_new_n495_; 
wire _abc_4635_new_n496_; 
wire _abc_4635_new_n498_; 
wire _abc_4635_new_n499_; 
wire _abc_4635_new_n501_; 
wire _abc_4635_new_n502_; 
wire _abc_4635_new_n504_; 
wire _abc_4635_new_n506_; 
wire _abc_4635_new_n508_; 
wire _abc_4635_new_n510_; 
wire _abc_4635_new_n512_; 
wire _abc_4635_new_n514_; 
wire _abc_4635_new_n516_; 
wire _abc_4635_new_n518_; 
wire _abc_4635_new_n520_; 
wire _abc_4635_new_n522_; 
wire _abc_4635_new_n524_; 
wire _abc_4635_new_n526_; 
wire _abc_4635_new_n528_; 
wire _abc_4635_new_n530_; 
wire _abc_4635_new_n532_; 
wire _abc_4635_new_n534_; 
wire _abc_4635_new_n536_; 
wire _abc_4635_new_n537_; 
wire _abc_4635_new_n538_; 
wire _abc_4635_new_n539_; 
wire _abc_4635_new_n541_; 
wire _abc_4635_new_n542_; 
wire _abc_4635_new_n544_; 
wire _abc_4635_new_n545_; 
wire _abc_4635_new_n547_; 
wire _abc_4635_new_n548_; 
wire _abc_4635_new_n550_; 
wire _abc_4635_new_n551_; 
wire _abc_4635_new_n553_; 
wire _abc_4635_new_n554_; 
wire _abc_4635_new_n556_; 
wire _abc_4635_new_n557_; 
wire _abc_4635_new_n559_; 
wire _abc_4635_new_n560_; 
wire _abc_4635_new_n562_; 
wire _abc_4635_new_n563_; 
wire _abc_4635_new_n565_; 
wire _abc_4635_new_n566_; 
wire _abc_4635_new_n568_; 
wire _abc_4635_new_n569_; 
wire _abc_4635_new_n571_; 
wire _abc_4635_new_n572_; 
wire _abc_4635_new_n574_; 
wire _abc_4635_new_n575_; 
wire _abc_4635_new_n577_; 
wire _abc_4635_new_n578_; 
wire _abc_4635_new_n580_; 
wire _abc_4635_new_n581_; 
wire _abc_4635_new_n583_; 
wire _abc_4635_new_n584_; 
wire _abc_4635_new_n586_; 
wire _abc_4635_new_n587_; 
wire _abc_4635_new_n589_; 
wire _abc_4635_new_n590_; 
wire _abc_4635_new_n592_; 
wire _abc_4635_new_n593_; 
wire _abc_4635_new_n595_; 
wire _abc_4635_new_n596_; 
wire _abc_4635_new_n598_; 
wire _abc_4635_new_n599_; 
wire _abc_4635_new_n601_; 
wire _abc_4635_new_n602_; 
wire _abc_4635_new_n604_; 
wire _abc_4635_new_n605_; 
wire _abc_4635_new_n607_; 
wire _abc_4635_new_n608_; 
wire _abc_4635_new_n610_; 
wire _abc_4635_new_n611_; 
wire _abc_4635_new_n613_; 
wire _abc_4635_new_n614_; 
wire _abc_4635_new_n616_; 
wire _abc_4635_new_n617_; 
wire _abc_4635_new_n619_; 
wire _abc_4635_new_n620_; 
wire _abc_4635_new_n622_; 
wire _abc_4635_new_n623_; 
wire _abc_4635_new_n625_; 
wire _abc_4635_new_n626_; 
wire _abc_4635_new_n628_; 
wire _abc_4635_new_n629_; 
wire _abc_4635_new_n631_; 
wire _abc_4635_new_n632_; 
wire _abc_4635_new_n634_; 
wire _abc_4635_new_n635_; 
wire _abc_4635_new_n636_; 
wire _abc_4635_new_n637_; 
wire _abc_4635_new_n639_; 
wire _abc_4635_new_n640_; 
wire _abc_4635_new_n641_; 
wire _abc_4635_new_n642_; 
wire _abc_4635_new_n643_; 
wire _abc_4635_new_n644_; 
wire _abc_4635_new_n645_; 
wire _abc_4635_new_n646_; 
wire _abc_4635_new_n647_; 
wire _abc_4635_new_n648_; 
wire _abc_4635_new_n649_; 
wire _abc_4635_new_n651_; 
wire _abc_4635_new_n652_; 
wire _abc_4635_new_n653_; 
wire _abc_4635_new_n654_; 
wire _abc_4635_new_n655_; 
wire _abc_4635_new_n656_; 
wire _abc_4635_new_n657_; 
wire _abc_4635_new_n658_; 
wire _abc_4635_new_n659_; 
wire _abc_4635_new_n661_; 
wire _abc_4635_new_n662_; 
wire _abc_4635_new_n663_; 
wire _abc_4635_new_n664_; 
wire _abc_4635_new_n665_; 
wire _abc_4635_new_n666_; 
wire _abc_4635_new_n667_; 
wire _abc_4635_new_n668_; 
wire _abc_4635_new_n669_; 
wire _abc_4635_new_n671_; 
wire _abc_4635_new_n672_; 
wire _abc_4635_new_n673_; 
wire _abc_4635_new_n674_; 
wire _abc_4635_new_n675_; 
wire _abc_4635_new_n676_; 
wire _abc_4635_new_n677_; 
wire _abc_4635_new_n678_; 
wire _abc_4635_new_n679_; 
wire _abc_4635_new_n681_; 
wire _abc_4635_new_n682_; 
wire _abc_4635_new_n683_; 
wire _abc_4635_new_n684_; 
wire _abc_4635_new_n685_; 
wire _abc_4635_new_n686_; 
wire _abc_4635_new_n688_; 
wire _abc_4635_new_n689_; 
wire _abc_4635_new_n690_; 
wire _abc_4635_new_n691_; 
wire _abc_4635_new_n692_; 
wire _abc_4635_new_n693_; 
wire _abc_4635_new_n695_; 
wire _abc_4635_new_n696_; 
wire _abc_4635_new_n697_; 
wire _abc_4635_new_n698_; 
wire _abc_4635_new_n699_; 
wire _abc_4635_new_n700_; 
wire _abc_4635_new_n701_; 
wire _abc_4635_new_n702_; 
wire _abc_4635_new_n703_; 
wire _abc_4635_new_n705_; 
wire _abc_4635_new_n706_; 
wire _abc_4635_new_n707_; 
wire _abc_4635_new_n708_; 
wire _abc_4635_new_n709_; 
wire _abc_4635_new_n710_; 
wire _abc_4635_new_n711_; 
wire _abc_4635_new_n712_; 
wire _abc_4635_new_n713_; 
wire _abc_4635_new_n714_; 
wire _abc_4635_new_n715_; 
wire _abc_4635_new_n717_; 
wire _abc_4635_new_n718_; 
wire _abc_4635_new_n719_; 
wire _abc_4635_new_n720_; 
wire _abc_4635_new_n722_; 
wire _abc_4635_new_n723_; 
wire _abc_4635_new_n725_; 
wire _abc_4635_new_n726_; 
wire _abc_4635_new_n728_; 
wire _abc_4635_new_n729_; 
wire _abc_4635_new_n731_; 
wire _abc_4635_new_n732_; 
wire _abc_4635_new_n734_; 
wire _abc_4635_new_n735_; 
wire _abc_4635_new_n737_; 
wire _abc_4635_new_n738_; 
wire _abc_4635_new_n740_; 
wire _abc_4635_new_n741_; 
wire _abc_4635_new_n743_; 
wire _abc_4635_new_n744_; 
wire _abc_4635_new_n746_; 
wire _abc_4635_new_n748_; 
wire _abc_4635_new_n750_; 
wire _abc_4635_new_n752_; 
wire _abc_4635_new_n754_; 
wire _abc_4635_new_n756_; 
wire _abc_4635_new_n758_; 
wire _abc_4635_new_n760_; 
wire _abc_4635_new_n762_; 
wire _abc_4635_new_n764_; 
wire _abc_4635_new_n766_; 
wire _abc_4635_new_n768_; 
wire _abc_4635_new_n770_; 
wire _abc_4635_new_n772_; 
wire _abc_4635_new_n774_; 
wire _abc_4635_new_n776_; 
wire _abc_4635_new_n778_; 
wire _abc_4635_new_n780_; 
wire _abc_4635_new_n781_; 
wire _abc_4635_new_n782_; 
wire _abc_4635_new_n783_; 
wire _abc_4635_new_n784_; 
wire _abc_4635_new_n785_; 
wire _abc_4635_new_n787_; 
wire _abc_4635_new_n788_; 
wire _abc_4635_new_n789_; 
wire _abc_4635_new_n790_; 
wire _abc_4635_new_n791_; 
wire _abc_4635_new_n792_; 
wire _abc_4635_new_n794_; 
wire _abc_4635_new_n795_; 
wire _abc_4635_new_n796_; 
wire _abc_4635_new_n797_; 
wire _abc_4635_new_n798_; 
wire _abc_4635_new_n799_; 
wire _abc_4635_new_n800_; 
wire _abc_4635_new_n801_; 
wire _abc_4635_new_n802_; 
wire _abc_4635_new_n804_; 
wire _abc_4635_new_n805_; 
wire _abc_4635_new_n806_; 
wire _abc_4635_new_n807_; 
wire _abc_4635_new_n808_; 
wire _abc_4635_new_n809_; 
wire _abc_4635_new_n810_; 
wire _abc_4635_new_n811_; 
wire _abc_4635_new_n813_; 
wire _abc_4635_new_n814_; 
wire _abc_4635_new_n815_; 
wire _abc_4635_new_n816_; 
wire _abc_4635_new_n817_; 
wire _abc_4635_new_n818_; 
wire _abc_4635_new_n819_; 
wire _abc_4635_new_n820_; 
wire _abc_4635_new_n821_; 
wire _abc_4635_new_n822_; 
wire _abc_4635_new_n823_; 
wire _abc_4635_new_n825_; 
wire _abc_4635_new_n826_; 
wire _abc_4635_new_n827_; 
wire _abc_4635_new_n828_; 
wire _abc_4635_new_n829_; 
wire _abc_4635_new_n830_; 
wire _abc_4635_new_n831_; 
wire _abc_4635_new_n832_; 
wire _abc_4635_new_n834_; 
wire _abc_4635_new_n835_; 
wire _abc_4635_new_n836_; 
wire _abc_4635_new_n837_; 
wire _abc_4635_new_n838_; 
wire _abc_4635_new_n839_; 
wire _abc_4635_new_n840_; 
wire _abc_4635_new_n841_; 
wire _abc_4635_new_n842_; 
wire _abc_4635_new_n843_; 
wire _abc_4635_new_n845_; 
wire _abc_4635_new_n846_; 
wire _abc_4635_new_n847_; 
wire _abc_4635_new_n848_; 
wire _abc_4635_new_n849_; 
wire _abc_4635_new_n850_; 
wire _abc_4635_new_n851_; 
wire _abc_4635_new_n853_; 
wire _abc_4635_new_n854_; 
wire _abc_4635_new_n855_; 
wire _abc_4635_new_n856_; 
wire _abc_4635_new_n857_; 
wire _abc_4635_new_n858_; 
wire _abc_4635_new_n859_; 
wire _abc_4635_new_n860_; 
wire _abc_4635_new_n861_; 
wire _abc_4635_new_n862_; 
wire _abc_4635_new_n863_; 
wire _abc_4635_new_n865_; 
wire _abc_4635_new_n866_; 
wire _abc_4635_new_n867_; 
wire _abc_4635_new_n868_; 
wire _abc_4635_new_n869_; 
wire _abc_4635_new_n870_; 
wire _abc_4635_new_n872_; 
wire _abc_4635_new_n873_; 
wire _abc_4635_new_n874_; 
wire _abc_4635_new_n875_; 
wire _abc_4635_new_n876_; 
wire _abc_4635_new_n877_; 
wire _abc_4635_new_n878_; 
wire _abc_4635_new_n879_; 
wire _abc_4635_new_n880_; 
wire _abc_4635_new_n881_; 
wire _abc_4635_new_n882_; 
wire _abc_4635_new_n883_; 
wire _abc_4635_new_n884_; 
wire _abc_4635_new_n885_; 
wire _abc_4635_new_n886_; 
wire _abc_4635_new_n887_; 
wire _abc_4635_new_n888_; 
wire _abc_4635_new_n889_; 
wire _abc_4635_new_n890_; 
wire _abc_4635_new_n891_; 
wire _abc_4635_new_n892_; 
wire _abc_4635_new_n893_; 
wire _abc_4635_new_n894_; 
wire _abc_4635_new_n896_; 
wire _abc_4635_new_n897_; 
wire _abc_4635_new_n898_; 
wire _abc_4635_new_n899_; 
wire _abc_4635_new_n900_; 
wire _abc_4635_new_n901_; 
wire _abc_4635_new_n902_; 
wire _abc_4635_new_n904_; 
wire _abc_4635_new_n905_; 
wire _abc_4635_new_n906_; 
wire _abc_4635_new_n907_; 
wire _abc_4635_new_n908_; 
wire _abc_4635_new_n909_; 
wire _abc_4635_new_n910_; 
wire _abc_4635_new_n911_; 
wire _abc_4635_new_n912_; 
wire _abc_4635_new_n913_; 
wire _abc_4635_new_n914_; 
wire _abc_4635_new_n916_; 
wire _abc_4635_new_n917_; 
wire _abc_4635_new_n918_; 
wire _abc_4635_new_n919_; 
wire _abc_4635_new_n920_; 
wire _abc_4635_new_n921_; 
wire _abc_4635_new_n923_; 
wire _abc_4635_new_n924_; 
wire _abc_4635_new_n925_; 
wire _abc_4635_new_n926_; 
wire _abc_4635_new_n927_; 
wire _abc_4635_new_n928_; 
wire _abc_4635_new_n929_; 
wire _abc_4635_new_n930_; 
wire _abc_4635_new_n931_; 
wire _abc_4635_new_n932_; 
wire _abc_4635_new_n933_; 
wire _abc_4635_new_n934_; 
wire _abc_4635_new_n935_; 
wire _abc_4635_new_n937_; 
wire _abc_4635_new_n938_; 
wire _abc_4635_new_n939_; 
wire _abc_4635_new_n940_; 
wire _abc_4635_new_n941_; 
wire _abc_4635_new_n943_; 
wire _abc_4635_new_n944_; 
wire _abc_4635_new_n945_; 
wire _abc_4635_new_n946_; 
wire _abc_4635_new_n947_; 
wire _abc_4635_new_n948_; 
wire _abc_4635_new_n949_; 
wire _abc_4635_new_n950_; 
wire _abc_4635_new_n951_; 
wire _abc_4635_new_n952_; 
wire _abc_4635_new_n953_; 
wire _abc_4635_new_n954_; 
wire _abc_4635_new_n955_; 
wire _abc_4635_new_n956_; 
wire _abc_4635_new_n957_; 
wire _abc_4635_new_n959_; 
wire _abc_4635_new_n960_; 
wire _abc_4635_new_n961_; 
wire _abc_4635_new_n962_; 
wire _abc_4635_new_n963_; 
wire _abc_4635_new_n964_; 
wire _abc_4635_new_n966_; 
wire _abc_4635_new_n967_; 
wire _abc_4635_new_n968_; 
wire _abc_4635_new_n969_; 
wire _abc_4635_new_n970_; 
wire _abc_4635_new_n971_; 
wire _abc_4635_new_n972_; 
wire _abc_4635_new_n973_; 
wire _abc_4635_new_n974_; 
wire _abc_4635_new_n975_; 
wire _abc_4635_new_n976_; 
wire _abc_4635_new_n977_; 
wire _abc_4635_new_n978_; 
wire _abc_4635_new_n980_; 
wire _abc_4635_new_n981_; 
wire _abc_4635_new_n982_; 
wire _abc_4635_new_n983_; 
wire _abc_4635_new_n984_; 
wire _abc_4635_new_n985_; 
wire _abc_4635_new_n987_; 
wire _abc_4635_new_n988_; 
wire _abc_4635_new_n989_; 
wire _abc_4635_new_n990_; 
wire _abc_4635_new_n991_; 
wire _abc_4635_new_n992_; 
wire _abc_4635_new_n993_; 
wire _abc_4635_new_n994_; 
wire _abc_4635_new_n995_; 
wire _abc_4635_new_n996_; 
wire _abc_4635_new_n997_; 
wire _abc_4635_new_n998_; 
wire _abc_4635_new_n999_; 
output align;
output \arprot[0] ;
output \arprot[1] ;
output \arprot[2] ;
output \awprot[0] ;
output \awprot[1] ;
output \awprot[2] ;
output busy;
input clock;
output done;
wire en_instr; 
input enable;
input \imm[0] ;
input \imm[10] ;
input \imm[11] ;
input \imm[12] ;
input \imm[13] ;
input \imm[14] ;
input \imm[15] ;
input \imm[16] ;
input \imm[17] ;
input \imm[18] ;
input \imm[19] ;
input \imm[1] ;
input \imm[20] ;
input \imm[21] ;
input \imm[22] ;
input \imm[23] ;
input \imm[24] ;
input \imm[25] ;
input \imm[26] ;
input \imm[27] ;
input \imm[28] ;
input \imm[29] ;
input \imm[2] ;
input \imm[30] ;
input \imm[31] ;
input \imm[3] ;
input \imm[4] ;
input \imm[5] ;
input \imm[6] ;
input \imm[7] ;
input \imm[8] ;
input \imm[9] ;
output \inst[0] ;
output \inst[10] ;
output \inst[11] ;
output \inst[12] ;
output \inst[13] ;
output \inst[14] ;
output \inst[15] ;
output \inst[16] ;
output \inst[17] ;
output \inst[18] ;
output \inst[19] ;
output \inst[1] ;
output \inst[20] ;
output \inst[21] ;
output \inst[22] ;
output \inst[23] ;
output \inst[24] ;
output \inst[25] ;
output \inst[26] ;
output \inst[27] ;
output \inst[28] ;
output \inst[29] ;
output \inst[2] ;
output \inst[30] ;
output \inst[31] ;
output \inst[3] ;
output \inst[4] ;
output \inst[5] ;
output \inst[6] ;
output \inst[7] ;
output \inst[8] ;
output \inst[9] ;
input \pc[0] ;
input \pc[10] ;
input \pc[11] ;
input \pc[12] ;
input \pc[13] ;
input \pc[14] ;
input \pc[15] ;
input \pc[16] ;
input \pc[17] ;
input \pc[18] ;
input \pc[19] ;
input \pc[1] ;
input \pc[20] ;
input \pc[21] ;
input \pc[22] ;
input \pc[23] ;
input \pc[24] ;
input \pc[25] ;
input \pc[26] ;
input \pc[27] ;
input \pc[28] ;
input \pc[29] ;
input \pc[2] ;
input \pc[30] ;
input \pc[31] ;
input \pc[3] ;
input \pc[4] ;
input \pc[5] ;
input \pc[6] ;
input \pc[7] ;
input \pc[8] ;
input \pc[9] ;
output \rd[0] ;
output \rd[10] ;
output \rd[11] ;
output \rd[12] ;
output \rd[13] ;
output \rd[14] ;
output \rd[15] ;
output \rd[16] ;
output \rd[17] ;
output \rd[18] ;
output \rd[19] ;
output \rd[1] ;
output \rd[20] ;
output \rd[21] ;
output \rd[22] ;
output \rd[23] ;
output \rd[24] ;
output \rd[25] ;
output \rd[26] ;
output \rd[27] ;
output \rd[28] ;
output \rd[29] ;
output \rd[2] ;
output \rd[30] ;
output \rd[31] ;
output \rd[3] ;
output \rd[4] ;
output \rd[5] ;
output \rd[6] ;
output \rd[7] ;
output \rd[8] ;
output \rd[9] ;
output rd_en;
input resetn;
input \rs1[0] ;
input \rs1[10] ;
input \rs1[11] ;
input \rs1[12] ;
input \rs1[13] ;
input \rs1[14] ;
input \rs1[15] ;
input \rs1[16] ;
input \rs1[17] ;
input \rs1[18] ;
input \rs1[19] ;
input \rs1[1] ;
input \rs1[20] ;
input \rs1[21] ;
input \rs1[22] ;
input \rs1[23] ;
input \rs1[24] ;
input \rs1[25] ;
input \rs1[26] ;
input \rs1[27] ;
input \rs1[28] ;
input \rs1[29] ;
input \rs1[2] ;
input \rs1[30] ;
input \rs1[31] ;
input \rs1[3] ;
input \rs1[4] ;
input \rs1[5] ;
input \rs1[6] ;
input \rs1[7] ;
input \rs1[8] ;
input \rs1[9] ;
input \rs2[0] ;
input \rs2[10] ;
input \rs2[11] ;
input \rs2[12] ;
input \rs2[13] ;
input \rs2[14] ;
input \rs2[15] ;
input \rs2[16] ;
input \rs2[17] ;
input \rs2[18] ;
input \rs2[19] ;
input \rs2[1] ;
input \rs2[20] ;
input \rs2[21] ;
input \rs2[22] ;
input \rs2[23] ;
input \rs2[24] ;
input \rs2[25] ;
input \rs2[26] ;
input \rs2[27] ;
input \rs2[28] ;
input \rs2[29] ;
input \rs2[2] ;
input \rs2[30] ;
input \rs2[31] ;
input \rs2[3] ;
input \rs2[4] ;
input \rs2[5] ;
input \rs2[6] ;
input \rs2[7] ;
input \rs2[8] ;
input \rs2[9] ;
input signo;
wire state_0_; 
wire state_1_; 
wire state_2_; 
wire state_3_; 
wire state_4_; 
wire state_5_; 
wire state_6_; 
input \wordsize[0] ;
input \wordsize[1] ;
AND2X2 AND2X2_1 ( .A(_abc_4635_new_n393_), .B(_abc_4635_new_n367_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_6_));
AND2X2 AND2X2_10 ( .A(_abc_4635_new_n758_), .B(_abc_4635_new_n641_), .Y(\rd[23] ));
AND2X2 AND2X2_11 ( .A(\rs1[2] ), .B(\imm[2] ), .Y(_abc_4635_new_n781_));
AND2X2 AND2X2_12 ( .A(\rs1[3] ), .B(\imm[3] ), .Y(_abc_4635_new_n789_));
AND2X2 AND2X2_13 ( .A(\rs1[4] ), .B(\imm[4] ), .Y(_abc_4635_new_n799_));
AND2X2 AND2X2_14 ( .A(\rs1[5] ), .B(\imm[5] ), .Y(_abc_4635_new_n808_));
AND2X2 AND2X2_15 ( .A(\rs1[6] ), .B(\imm[6] ), .Y(_abc_4635_new_n818_));
AND2X2 AND2X2_16 ( .A(\rs1[7] ), .B(\imm[7] ), .Y(_abc_4635_new_n829_));
AND2X2 AND2X2_17 ( .A(\rs1[8] ), .B(\imm[8] ), .Y(_abc_4635_new_n840_));
AND2X2 AND2X2_18 ( .A(\rs1[9] ), .B(\imm[9] ), .Y(_abc_4635_new_n848_));
AND2X2 AND2X2_19 ( .A(\rs1[10] ), .B(\imm[10] ), .Y(_abc_4635_new_n858_));
AND2X2 AND2X2_2 ( .A(_abc_4635_new_n649_), .B(_abc_4635_new_n641_), .Y(\rd[0] ));
AND2X2 AND2X2_20 ( .A(\rs1[11] ), .B(\imm[11] ), .Y(_abc_4635_new_n867_));
AND2X2 AND2X2_21 ( .A(\rs1[13] ), .B(\imm[13] ), .Y(_abc_4635_new_n899_));
AND2X2 AND2X2_22 ( .A(\rs1[14] ), .B(\imm[14] ), .Y(_abc_4635_new_n911_));
AND2X2 AND2X2_23 ( .A(\rs1[15] ), .B(\imm[15] ), .Y(_abc_4635_new_n918_));
AND2X2 AND2X2_24 ( .A(_abc_4635_new_n934_), .B(_abc_4635_new_n939_), .Y(_abc_4635_new_n949_));
AND2X2 AND2X2_25 ( .A(_abc_4635_new_n950_), .B(_abc_4635_new_n955_), .Y(_abc_4635_new_n956_));
AND2X2 AND2X2_26 ( .A(\rs1[19] ), .B(\imm[19] ), .Y(_abc_4635_new_n960_));
AND2X2 AND2X2_27 ( .A(_abc_4635_new_n973_), .B(_abc_4635_new_n976_), .Y(_abc_4635_new_n977_));
AND2X2 AND2X2_28 ( .A(\rs1[23] ), .B(\imm[23] ), .Y(_abc_4635_new_n1005_));
AND2X2 AND2X2_29 ( .A(_abc_4635_new_n1004_), .B(_abc_4635_new_n1007_), .Y(_abc_4635_new_n1008_));
AND2X2 AND2X2_3 ( .A(_abc_4635_new_n659_), .B(_abc_4635_new_n641_), .Y(\rd[1] ));
AND2X2 AND2X2_30 ( .A(_abc_4635_new_n1013_), .B(_abc_4635_new_n990_), .Y(_abc_4635_new_n1014_));
AND2X2 AND2X2_31 ( .A(_abc_4635_new_n888_), .B(_abc_4635_new_n925_), .Y(_abc_4635_new_n1028_));
AND2X2 AND2X2_32 ( .A(\rs1[25] ), .B(\imm[25] ), .Y(_abc_4635_new_n1037_));
AND2X2 AND2X2_33 ( .A(_abc_4635_new_n1096_), .B(_abc_4635_new_n1097_), .Y(_abc_4635_new_n1098_));
AND2X2 AND2X2_34 ( .A(_abc_4635_new_n537_), .B(_abc_4635_new_n641_), .Y(rd_en));
AND2X2 AND2X2_4 ( .A(_abc_4635_new_n669_), .B(_abc_4635_new_n641_), .Y(\rd[2] ));
AND2X2 AND2X2_5 ( .A(_abc_4635_new_n679_), .B(_abc_4635_new_n641_), .Y(\rd[3] ));
AND2X2 AND2X2_6 ( .A(_abc_4635_new_n686_), .B(_abc_4635_new_n641_), .Y(\rd[4] ));
AND2X2 AND2X2_7 ( .A(_abc_4635_new_n693_), .B(_abc_4635_new_n641_), .Y(\rd[5] ));
AND2X2 AND2X2_8 ( .A(_abc_4635_new_n703_), .B(_abc_4635_new_n641_), .Y(\rd[6] ));
AND2X2 AND2X2_9 ( .A(_abc_4635_new_n432_), .B(signo), .Y(_abc_4635_new_n717_));
AOI21X1 AOI21X1_1 ( .A(state_6_), .B(AWready), .C(state_1_), .Y(_abc_4635_new_n363_));
AOI21X1 AOI21X1_10 ( .A(_abc_4635_new_n486_), .B(_abc_4635_new_n487_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__10_));
AOI21X1 AOI21X1_100 ( .A(_abc_4635_new_n795_), .B(_abc_4635_new_n781_), .C(_abc_4635_new_n789_), .Y(_abc_4635_new_n796_));
AOI21X1 AOI21X1_101 ( .A(_abc_4635_new_n814_), .B(_abc_4635_new_n799_), .C(_abc_4635_new_n808_), .Y(_abc_4635_new_n815_));
AOI21X1 AOI21X1_102 ( .A(_abc_4635_new_n830_), .B(_abc_4635_new_n818_), .C(_abc_4635_new_n829_), .Y(_abc_4635_new_n837_));
AOI21X1 AOI21X1_103 ( .A(_abc_4635_new_n836_), .B(_abc_4635_new_n797_), .C(_abc_4635_new_n838_), .Y(_abc_4635_new_n839_));
AOI21X1 AOI21X1_104 ( .A(_abc_4635_new_n854_), .B(_abc_4635_new_n840_), .C(_abc_4635_new_n848_), .Y(_abc_4635_new_n855_));
AOI21X1 AOI21X1_105 ( .A(_abc_4635_new_n857_), .B(_abc_4635_new_n860_), .C(_abc_4635_new_n858_), .Y(_abc_4635_new_n865_));
AOI21X1 AOI21X1_106 ( .A(_abc_4635_new_n868_), .B(_abc_4635_new_n858_), .C(_abc_4635_new_n867_), .Y(_abc_4635_new_n874_));
AOI21X1 AOI21X1_107 ( .A(_abc_4635_new_n882_), .B(_abc_4635_new_n883_), .C(_abc_4635_new_n884_), .Y(_abc_4635_new_n885_));
AOI21X1 AOI21X1_108 ( .A(_abc_4635_new_n794_), .B(_abc_4635_new_n796_), .C(_abc_4635_new_n886_), .Y(_abc_4635_new_n887_));
AOI21X1 AOI21X1_109 ( .A(_abc_4635_new_n910_), .B(_abc_4635_new_n913_), .C(_abc_4635_new_n911_), .Y(_abc_4635_new_n916_));
AOI21X1 AOI21X1_11 ( .A(_abc_4635_new_n489_), .B(_abc_4635_new_n490_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__11_));
AOI21X1 AOI21X1_110 ( .A(_abc_4635_new_n919_), .B(_abc_4635_new_n911_), .C(_abc_4635_new_n918_), .Y(_abc_4635_new_n927_));
AOI21X1 AOI21X1_111 ( .A(_abc_4635_new_n875_), .B(_abc_4635_new_n925_), .C(_abc_4635_new_n928_), .Y(_abc_4635_new_n929_));
AOI21X1 AOI21X1_112 ( .A(_abc_4635_new_n930_), .B(_abc_4635_new_n949_), .C(_abc_4635_new_n948_), .Y(_abc_4635_new_n950_));
AOI21X1 AOI21X1_113 ( .A(_abc_4635_new_n962_), .B(_abc_4635_new_n952_), .C(_abc_4635_new_n960_), .Y(_abc_4635_new_n968_));
AOI21X1 AOI21X1_114 ( .A(_abc_4635_new_n930_), .B(_abc_4635_new_n972_), .C(_abc_4635_new_n969_), .Y(_abc_4635_new_n973_));
AOI21X1 AOI21X1_115 ( .A(_abc_4635_new_n930_), .B(_abc_4635_new_n1016_), .C(_abc_4635_new_n1021_), .Y(_abc_4635_new_n1022_));
AOI21X1 AOI21X1_116 ( .A(_abc_4635_new_n1029_), .B(_abc_4635_new_n929_), .C(_abc_4635_new_n1030_), .Y(_abc_4635_new_n1031_));
AOI21X1 AOI21X1_117 ( .A(_abc_4635_new_n1039_), .B(_abc_4635_new_n1025_), .C(_abc_4635_new_n1037_), .Y(_abc_4635_new_n1044_));
AOI21X1 AOI21X1_118 ( .A(_abc_4635_new_n1072_), .B(_abc_4635_new_n1092_), .C(_abc_4635_new_n1094_), .Y(_abc_4635_new_n1095_));
AOI21X1 AOI21X1_119 ( .A(_abc_4635_new_n1101_), .B(_abc_4635_new_n1071_), .C(_abc_4635_new_n1091_), .Y(_abc_4635_new_n1102_));
AOI21X1 AOI21X1_12 ( .A(_abc_4635_new_n492_), .B(_abc_4635_new_n493_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__12_));
AOI21X1 AOI21X1_120 ( .A(_abc_4635_new_n1117_), .B(_abc_4635_new_n1115_), .C(_abc_4635_new_n366_), .Y(Bready));
AOI21X1 AOI21X1_13 ( .A(_abc_4635_new_n495_), .B(_abc_4635_new_n496_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__13_));
AOI21X1 AOI21X1_14 ( .A(_abc_4635_new_n498_), .B(_abc_4635_new_n499_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__14_));
AOI21X1 AOI21X1_15 ( .A(_abc_4635_new_n501_), .B(_abc_4635_new_n502_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__15_));
AOI21X1 AOI21X1_16 ( .A(_abc_4635_new_n481_), .B(_abc_4635_new_n520_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__24_));
AOI21X1 AOI21X1_17 ( .A(_abc_4635_new_n484_), .B(_abc_4635_new_n522_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__25_));
AOI21X1 AOI21X1_18 ( .A(_abc_4635_new_n487_), .B(_abc_4635_new_n524_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__26_));
AOI21X1 AOI21X1_19 ( .A(_abc_4635_new_n490_), .B(_abc_4635_new_n526_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__27_));
AOI21X1 AOI21X1_2 ( .A(Bvalid), .B(_abc_4635_new_n364_), .C(_abc_4635_new_n405_), .Y(_abc_4635_new_n406_));
AOI21X1 AOI21X1_20 ( .A(_abc_4635_new_n493_), .B(_abc_4635_new_n528_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__28_));
AOI21X1 AOI21X1_21 ( .A(_abc_4635_new_n496_), .B(_abc_4635_new_n530_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__29_));
AOI21X1 AOI21X1_22 ( .A(_abc_4635_new_n499_), .B(_abc_4635_new_n532_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__30_));
AOI21X1 AOI21X1_23 ( .A(_abc_4635_new_n502_), .B(_abc_4635_new_n534_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__31_));
AOI21X1 AOI21X1_24 ( .A(_abc_4635_new_n536_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n539_), .Y(_0inst_31_0__0_));
AOI21X1 AOI21X1_25 ( .A(_abc_4635_new_n541_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n542_), .Y(_0inst_31_0__1_));
AOI21X1 AOI21X1_26 ( .A(_abc_4635_new_n544_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n545_), .Y(_0inst_31_0__2_));
AOI21X1 AOI21X1_27 ( .A(_abc_4635_new_n547_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n548_), .Y(_0inst_31_0__3_));
AOI21X1 AOI21X1_28 ( .A(_abc_4635_new_n550_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n551_), .Y(_0inst_31_0__4_));
AOI21X1 AOI21X1_29 ( .A(_abc_4635_new_n553_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n554_), .Y(_0inst_31_0__5_));
AOI21X1 AOI21X1_3 ( .A(state_4_), .B(_abc_4635_new_n396_), .C(_abc_4635_new_n427_), .Y(_abc_4635_new_n428_));
AOI21X1 AOI21X1_30 ( .A(_abc_4635_new_n556_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n557_), .Y(_0inst_31_0__6_));
AOI21X1 AOI21X1_31 ( .A(_abc_4635_new_n559_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n560_), .Y(_0inst_31_0__7_));
AOI21X1 AOI21X1_32 ( .A(_abc_4635_new_n562_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n563_), .Y(_0inst_31_0__8_));
AOI21X1 AOI21X1_33 ( .A(_abc_4635_new_n565_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n566_), .Y(_0inst_31_0__9_));
AOI21X1 AOI21X1_34 ( .A(_abc_4635_new_n568_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n569_), .Y(_0inst_31_0__10_));
AOI21X1 AOI21X1_35 ( .A(_abc_4635_new_n571_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n572_), .Y(_0inst_31_0__11_));
AOI21X1 AOI21X1_36 ( .A(_abc_4635_new_n574_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n575_), .Y(_0inst_31_0__12_));
AOI21X1 AOI21X1_37 ( .A(_abc_4635_new_n577_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n578_), .Y(_0inst_31_0__13_));
AOI21X1 AOI21X1_38 ( .A(_abc_4635_new_n580_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n581_), .Y(_0inst_31_0__14_));
AOI21X1 AOI21X1_39 ( .A(_abc_4635_new_n583_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n584_), .Y(_0inst_31_0__15_));
AOI21X1 AOI21X1_4 ( .A(_abc_4635_new_n432_), .B(_abc_4635_new_n443_), .C(_abc_4635_new_n451_), .Y(_0Wstrb_3_0__0_));
AOI21X1 AOI21X1_40 ( .A(_abc_4635_new_n586_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n587_), .Y(_0inst_31_0__16_));
AOI21X1 AOI21X1_41 ( .A(_abc_4635_new_n589_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n590_), .Y(_0inst_31_0__17_));
AOI21X1 AOI21X1_42 ( .A(_abc_4635_new_n592_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n593_), .Y(_0inst_31_0__18_));
AOI21X1 AOI21X1_43 ( .A(_abc_4635_new_n595_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n596_), .Y(_0inst_31_0__19_));
AOI21X1 AOI21X1_44 ( .A(_abc_4635_new_n598_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n599_), .Y(_0inst_31_0__20_));
AOI21X1 AOI21X1_45 ( .A(_abc_4635_new_n601_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n602_), .Y(_0inst_31_0__21_));
AOI21X1 AOI21X1_46 ( .A(_abc_4635_new_n604_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n605_), .Y(_0inst_31_0__22_));
AOI21X1 AOI21X1_47 ( .A(_abc_4635_new_n607_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n608_), .Y(_0inst_31_0__23_));
AOI21X1 AOI21X1_48 ( .A(_abc_4635_new_n610_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n611_), .Y(_0inst_31_0__24_));
AOI21X1 AOI21X1_49 ( .A(_abc_4635_new_n613_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n614_), .Y(_0inst_31_0__25_));
AOI21X1 AOI21X1_5 ( .A(_abc_4635_new_n454_), .B(_abc_4635_new_n448_), .C(_abc_4635_new_n450_), .Y(_0Wstrb_3_0__1_));
AOI21X1 AOI21X1_50 ( .A(_abc_4635_new_n616_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n617_), .Y(_0inst_31_0__26_));
AOI21X1 AOI21X1_51 ( .A(_abc_4635_new_n619_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n620_), .Y(_0inst_31_0__27_));
AOI21X1 AOI21X1_52 ( .A(_abc_4635_new_n622_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n623_), .Y(_0inst_31_0__28_));
AOI21X1 AOI21X1_53 ( .A(_abc_4635_new_n625_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n626_), .Y(_0inst_31_0__29_));
AOI21X1 AOI21X1_54 ( .A(_abc_4635_new_n628_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n629_), .Y(_0inst_31_0__30_));
AOI21X1 AOI21X1_55 ( .A(_abc_4635_new_n631_), .B(_abc_4635_new_n538_), .C(_abc_4635_new_n632_), .Y(_0inst_31_0__31_));
AOI21X1 AOI21X1_56 ( .A(_abc_4635_new_n457_), .B(_abc_4635_new_n445_), .C(_abc_4635_new_n636_), .Y(_abc_4635_new_n637_));
AOI21X1 AOI21X1_57 ( .A(_abc_4635_new_n655_), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n656_), .Y(_abc_4635_new_n657_));
AOI21X1 AOI21X1_58 ( .A(\Rdata_mem[1] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n657_), .Y(_abc_4635_new_n658_));
AOI21X1 AOI21X1_59 ( .A(_abc_4635_new_n665_), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n666_), .Y(_abc_4635_new_n667_));
AOI21X1 AOI21X1_6 ( .A(_abc_4635_new_n458_), .B(_abc_4635_new_n448_), .C(_abc_4635_new_n450_), .Y(_0Wstrb_3_0__2_));
AOI21X1 AOI21X1_60 ( .A(\Rdata_mem[2] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n667_), .Y(_abc_4635_new_n668_));
AOI21X1 AOI21X1_61 ( .A(_abc_4635_new_n675_), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n676_), .Y(_abc_4635_new_n677_));
AOI21X1 AOI21X1_62 ( .A(\Rdata_mem[3] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n677_), .Y(_abc_4635_new_n678_));
AOI21X1 AOI21X1_63 ( .A(_abc_4635_new_n699_), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n700_), .Y(_abc_4635_new_n701_));
AOI21X1 AOI21X1_64 ( .A(\Rdata_mem[6] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n701_), .Y(_abc_4635_new_n702_));
AOI21X1 AOI21X1_65 ( .A(_abc_4635_new_n456_), .B(_abc_4635_new_n705_), .C(_abc_4635_new_n446_), .Y(_abc_4635_new_n706_));
AOI21X1 AOI21X1_66 ( .A(_abc_4635_new_n715_), .B(_abc_4635_new_n707_), .C(_abc_4635_new_n640_), .Y(\rd[7] ));
AOI21X1 AOI21X1_67 ( .A(\Rdata_mem[8] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n719_), .Y(_abc_4635_new_n720_));
AOI21X1 AOI21X1_68 ( .A(_abc_4635_new_n718_), .B(_abc_4635_new_n720_), .C(_abc_4635_new_n640_), .Y(\rd[8] ));
AOI21X1 AOI21X1_69 ( .A(\Rdata_mem[9] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n722_), .Y(_abc_4635_new_n723_));
AOI21X1 AOI21X1_7 ( .A(_abc_4635_new_n460_), .B(_abc_4635_new_n448_), .C(_abc_4635_new_n450_), .Y(_0Wstrb_3_0__3_));
AOI21X1 AOI21X1_70 ( .A(_abc_4635_new_n718_), .B(_abc_4635_new_n723_), .C(_abc_4635_new_n640_), .Y(\rd[9] ));
AOI21X1 AOI21X1_71 ( .A(\Rdata_mem[10] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n725_), .Y(_abc_4635_new_n726_));
AOI21X1 AOI21X1_72 ( .A(_abc_4635_new_n718_), .B(_abc_4635_new_n726_), .C(_abc_4635_new_n640_), .Y(\rd[10] ));
AOI21X1 AOI21X1_73 ( .A(\Rdata_mem[11] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n728_), .Y(_abc_4635_new_n729_));
AOI21X1 AOI21X1_74 ( .A(_abc_4635_new_n718_), .B(_abc_4635_new_n729_), .C(_abc_4635_new_n640_), .Y(\rd[11] ));
AOI21X1 AOI21X1_75 ( .A(\Rdata_mem[12] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n731_), .Y(_abc_4635_new_n732_));
AOI21X1 AOI21X1_76 ( .A(_abc_4635_new_n718_), .B(_abc_4635_new_n732_), .C(_abc_4635_new_n640_), .Y(\rd[12] ));
AOI21X1 AOI21X1_77 ( .A(\Rdata_mem[13] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n734_), .Y(_abc_4635_new_n735_));
AOI21X1 AOI21X1_78 ( .A(_abc_4635_new_n718_), .B(_abc_4635_new_n735_), .C(_abc_4635_new_n640_), .Y(\rd[13] ));
AOI21X1 AOI21X1_79 ( .A(\Rdata_mem[14] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n737_), .Y(_abc_4635_new_n738_));
AOI21X1 AOI21X1_8 ( .A(_abc_4635_new_n480_), .B(_abc_4635_new_n481_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__8_));
AOI21X1 AOI21X1_80 ( .A(_abc_4635_new_n718_), .B(_abc_4635_new_n738_), .C(_abc_4635_new_n640_), .Y(\rd[14] ));
AOI21X1 AOI21X1_81 ( .A(_abc_4635_new_n712_), .B(_abc_4635_new_n711_), .C(_abc_4635_new_n446_), .Y(_abc_4635_new_n740_));
AOI21X1 AOI21X1_82 ( .A(\Rdata_mem[15] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n740_), .Y(_abc_4635_new_n741_));
AOI21X1 AOI21X1_83 ( .A(_abc_4635_new_n718_), .B(_abc_4635_new_n741_), .C(_abc_4635_new_n640_), .Y(\rd[15] ));
AOI21X1 AOI21X1_84 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n743_), .C(_abc_4635_new_n640_), .Y(\rd[16] ));
AOI21X1 AOI21X1_85 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n746_), .C(_abc_4635_new_n640_), .Y(\rd[17] ));
AOI21X1 AOI21X1_86 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n748_), .C(_abc_4635_new_n640_), .Y(\rd[18] ));
AOI21X1 AOI21X1_87 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n750_), .C(_abc_4635_new_n640_), .Y(\rd[19] ));
AOI21X1 AOI21X1_88 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n752_), .C(_abc_4635_new_n640_), .Y(\rd[20] ));
AOI21X1 AOI21X1_89 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n754_), .C(_abc_4635_new_n640_), .Y(\rd[21] ));
AOI21X1 AOI21X1_9 ( .A(_abc_4635_new_n483_), .B(_abc_4635_new_n484_), .C(_abc_4635_new_n478_), .Y(_0Wdata_31_0__9_));
AOI21X1 AOI21X1_90 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n756_), .C(_abc_4635_new_n640_), .Y(\rd[22] ));
AOI21X1 AOI21X1_91 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n760_), .C(_abc_4635_new_n640_), .Y(\rd[24] ));
AOI21X1 AOI21X1_92 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n762_), .C(_abc_4635_new_n640_), .Y(\rd[25] ));
AOI21X1 AOI21X1_93 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n764_), .C(_abc_4635_new_n640_), .Y(\rd[26] ));
AOI21X1 AOI21X1_94 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n766_), .C(_abc_4635_new_n640_), .Y(\rd[27] ));
AOI21X1 AOI21X1_95 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n768_), .C(_abc_4635_new_n640_), .Y(\rd[28] ));
AOI21X1 AOI21X1_96 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n770_), .C(_abc_4635_new_n640_), .Y(\rd[29] ));
AOI21X1 AOI21X1_97 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n772_), .C(_abc_4635_new_n640_), .Y(\rd[30] ));
AOI21X1 AOI21X1_98 ( .A(_abc_4635_new_n744_), .B(_abc_4635_new_n774_), .C(_abc_4635_new_n640_), .Y(\rd[31] ));
AOI21X1 AOI21X1_99 ( .A(_abc_4635_new_n780_), .B(_abc_4635_new_n783_), .C(_abc_4635_new_n781_), .Y(_abc_4635_new_n787_));
AOI22X1 AOI22X1_1 ( .A(state_4_), .B(_abc_4635_new_n369_), .C(_abc_4635_new_n370_), .D(_abc_4635_new_n377_), .Y(_abc_4635_new_n378_));
AOI22X1 AOI22X1_10 ( .A(\rs2[7] ), .B(_abc_4635_new_n432_), .C(\rs2[15] ), .D(_abc_4635_new_n445_), .Y(_abc_4635_new_n502_));
AOI22X1 AOI22X1_11 ( .A(_abc_4635_new_n448_), .B(\rs2[0] ), .C(\rs2[16] ), .D(_abc_4635_new_n479_), .Y(_abc_4635_new_n504_));
AOI22X1 AOI22X1_12 ( .A(_abc_4635_new_n448_), .B(\rs2[1] ), .C(\rs2[17] ), .D(_abc_4635_new_n479_), .Y(_abc_4635_new_n506_));
AOI22X1 AOI22X1_13 ( .A(_abc_4635_new_n448_), .B(\rs2[2] ), .C(\rs2[18] ), .D(_abc_4635_new_n479_), .Y(_abc_4635_new_n508_));
AOI22X1 AOI22X1_14 ( .A(_abc_4635_new_n448_), .B(\rs2[3] ), .C(\rs2[19] ), .D(_abc_4635_new_n479_), .Y(_abc_4635_new_n510_));
AOI22X1 AOI22X1_15 ( .A(_abc_4635_new_n448_), .B(\rs2[4] ), .C(\rs2[20] ), .D(_abc_4635_new_n479_), .Y(_abc_4635_new_n512_));
AOI22X1 AOI22X1_16 ( .A(_abc_4635_new_n448_), .B(\rs2[5] ), .C(\rs2[21] ), .D(_abc_4635_new_n479_), .Y(_abc_4635_new_n514_));
AOI22X1 AOI22X1_17 ( .A(_abc_4635_new_n448_), .B(\rs2[6] ), .C(\rs2[22] ), .D(_abc_4635_new_n479_), .Y(_abc_4635_new_n516_));
AOI22X1 AOI22X1_18 ( .A(_abc_4635_new_n448_), .B(\rs2[7] ), .C(\rs2[23] ), .D(_abc_4635_new_n479_), .Y(_abc_4635_new_n518_));
AOI22X1 AOI22X1_19 ( .A(\Rdata_mem[16] ), .B(_abc_4635_new_n447_), .C(\Rdata_mem[0] ), .D(_abc_4635_new_n647_), .Y(_abc_4635_new_n648_));
AOI22X1 AOI22X1_2 ( .A(Rvalid), .B(_abc_4635_new_n402_), .C(_abc_4635_new_n399_), .D(_abc_4635_new_n389_), .Y(_abc_4635_new_n403_));
AOI22X1 AOI22X1_20 ( .A(\Rdata_mem[20] ), .B(_abc_4635_new_n447_), .C(\Rdata_mem[4] ), .D(_abc_4635_new_n647_), .Y(_abc_4635_new_n685_));
AOI22X1 AOI22X1_21 ( .A(\Rdata_mem[21] ), .B(_abc_4635_new_n447_), .C(\Rdata_mem[5] ), .D(_abc_4635_new_n647_), .Y(_abc_4635_new_n692_));
AOI22X1 AOI22X1_22 ( .A(\Rdata_mem[7] ), .B(_abc_4635_new_n441_), .C(\Rdata_mem[23] ), .D(_abc_4635_new_n443_), .Y(_abc_4635_new_n708_));
AOI22X1 AOI22X1_23 ( .A(\Rdata_mem[7] ), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n432_), .D(_abc_4635_new_n714_), .Y(_abc_4635_new_n715_));
AOI22X1 AOI22X1_24 ( .A(signo), .B(_abc_4635_new_n740_), .C(_abc_4635_new_n717_), .D(_abc_4635_new_n714_), .Y(_abc_4635_new_n744_));
AOI22X1 AOI22X1_3 ( .A(\rs2[0] ), .B(_abc_4635_new_n432_), .C(\rs2[8] ), .D(_abc_4635_new_n445_), .Y(_abc_4635_new_n481_));
AOI22X1 AOI22X1_4 ( .A(\rs2[1] ), .B(_abc_4635_new_n432_), .C(\rs2[9] ), .D(_abc_4635_new_n445_), .Y(_abc_4635_new_n484_));
AOI22X1 AOI22X1_5 ( .A(\rs2[2] ), .B(_abc_4635_new_n432_), .C(\rs2[10] ), .D(_abc_4635_new_n445_), .Y(_abc_4635_new_n487_));
AOI22X1 AOI22X1_6 ( .A(\rs2[3] ), .B(_abc_4635_new_n432_), .C(\rs2[11] ), .D(_abc_4635_new_n445_), .Y(_abc_4635_new_n490_));
AOI22X1 AOI22X1_7 ( .A(\rs2[4] ), .B(_abc_4635_new_n432_), .C(\rs2[12] ), .D(_abc_4635_new_n445_), .Y(_abc_4635_new_n493_));
AOI22X1 AOI22X1_8 ( .A(\rs2[5] ), .B(_abc_4635_new_n432_), .C(\rs2[13] ), .D(_abc_4635_new_n445_), .Y(_abc_4635_new_n496_));
AOI22X1 AOI22X1_9 ( .A(\rs2[6] ), .B(_abc_4635_new_n432_), .C(\rs2[14] ), .D(_abc_4635_new_n445_), .Y(_abc_4635_new_n499_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_0_), .Q(state_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(_0Wdata_31_0__2_), .Q(\Wdata[2] ));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(_0Wdata_31_0__3_), .Q(\Wdata[3] ));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(_0Wdata_31_0__4_), .Q(\Wdata[4] ));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(_0Wdata_31_0__5_), .Q(\Wdata[5] ));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(_0Wdata_31_0__6_), .Q(\Wdata[6] ));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(_0Wdata_31_0__7_), .Q(\Wdata[7] ));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(_0Wdata_31_0__8_), .Q(\Wdata[8] ));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(_0Wdata_31_0__9_), .Q(\Wdata[9] ));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(_0Wdata_31_0__10_), .Q(\Wdata[10] ));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(_0Wdata_31_0__11_), .Q(\Wdata[11] ));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_1_), .Q(state_1_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(_0Wdata_31_0__12_), .Q(\Wdata[12] ));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(_0Wdata_31_0__13_), .Q(\Wdata[13] ));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(_0Wdata_31_0__14_), .Q(\Wdata[14] ));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(_0Wdata_31_0__15_), .Q(\Wdata[15] ));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(_0Wdata_31_0__16_), .Q(\Wdata[16] ));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(_0Wdata_31_0__17_), .Q(\Wdata[17] ));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(_0Wdata_31_0__18_), .Q(\Wdata[18] ));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(_0Wdata_31_0__19_), .Q(\Wdata[19] ));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(_0Wdata_31_0__20_), .Q(\Wdata[20] ));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock), .D(_0Wdata_31_0__21_), .Q(\Wdata[21] ));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_2_), .Q(state_2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock), .D(_0Wdata_31_0__22_), .Q(\Wdata[22] ));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock), .D(_0Wdata_31_0__23_), .Q(\Wdata[23] ));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock), .D(_0Wdata_31_0__24_), .Q(\Wdata[24] ));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clock), .D(_0Wdata_31_0__25_), .Q(\Wdata[25] ));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clock), .D(_0Wdata_31_0__26_), .Q(\Wdata[26] ));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clock), .D(_0Wdata_31_0__27_), .Q(\Wdata[27] ));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clock), .D(_0Wdata_31_0__28_), .Q(\Wdata[28] ));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clock), .D(_0Wdata_31_0__29_), .Q(\Wdata[29] ));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clock), .D(_0Wdata_31_0__30_), .Q(\Wdata[30] ));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clock), .D(_0Wdata_31_0__31_), .Q(\Wdata[31] ));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_3_), .Q(state_3_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clock), .D(_0inst_31_0__0_), .Q(\inst[0] ));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clock), .D(_0inst_31_0__1_), .Q(\inst[1] ));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clock), .D(_0inst_31_0__2_), .Q(\inst[2] ));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clock), .D(_0inst_31_0__3_), .Q(\inst[3] ));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clock), .D(_0inst_31_0__4_), .Q(\inst[4] ));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clock), .D(_0inst_31_0__5_), .Q(\inst[5] ));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clock), .D(_0inst_31_0__6_), .Q(\inst[6] ));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clock), .D(_0inst_31_0__7_), .Q(\inst[7] ));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clock), .D(_0inst_31_0__8_), .Q(\inst[8] ));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock), .D(_0inst_31_0__9_), .Q(\inst[9] ));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_4_), .Q(state_4_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock), .D(_0inst_31_0__10_), .Q(\inst[10] ));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock), .D(_0inst_31_0__11_), .Q(\inst[11] ));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clock), .D(_0inst_31_0__12_), .Q(\inst[12] ));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clock), .D(_0inst_31_0__13_), .Q(\inst[13] ));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clock), .D(_0inst_31_0__14_), .Q(\inst[14] ));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clock), .D(_0inst_31_0__15_), .Q(\inst[15] ));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clock), .D(_0inst_31_0__16_), .Q(\inst[16] ));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clock), .D(_0inst_31_0__17_), .Q(\inst[17] ));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clock), .D(_0inst_31_0__18_), .Q(\inst[18] ));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clock), .D(_0inst_31_0__19_), .Q(\inst[19] ));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_5_), .Q(state_5_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clock), .D(_0inst_31_0__20_), .Q(\inst[20] ));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clock), .D(_0inst_31_0__21_), .Q(\inst[21] ));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clock), .D(_0inst_31_0__22_), .Q(\inst[22] ));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clock), .D(_0inst_31_0__23_), .Q(\inst[23] ));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clock), .D(_0inst_31_0__24_), .Q(\inst[24] ));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clock), .D(_0inst_31_0__25_), .Q(\inst[25] ));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clock), .D(_0inst_31_0__26_), .Q(\inst[26] ));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clock), .D(_0inst_31_0__27_), .Q(\inst[27] ));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clock), .D(_0inst_31_0__28_), .Q(\inst[28] ));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clock), .D(_0inst_31_0__29_), .Q(\inst[29] ));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_6_), .Q(state_6_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clock), .D(_0inst_31_0__30_), .Q(\inst[30] ));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clock), .D(_0inst_31_0__31_), .Q(\inst[31] ));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clock), .D(_0Wstrb_3_0__0_), .Q(\Wstrb[0] ));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clock), .D(_0Wstrb_3_0__1_), .Q(\Wstrb[1] ));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clock), .D(_0Wstrb_3_0__2_), .Q(\Wstrb[2] ));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clock), .D(_0Wstrb_3_0__3_), .Q(\Wstrb[3] ));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(_0Wdata_31_0__0_), .Q(\Wdata[0] ));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(_0Wdata_31_0__1_), .Q(\Wdata[1] ));
INVX1 INVX1_1 ( .A(Wready), .Y(_abc_4635_new_n361_));
INVX1 INVX1_10 ( .A(_abc_4635_new_n384_), .Y(_abc_4635_new_n385_));
INVX1 INVX1_100 ( .A(_abc_4635_new_n990_), .Y(_abc_4635_new_n991_));
INVX1 INVX1_101 ( .A(\rs1[22] ), .Y(_abc_4635_new_n994_));
INVX1 INVX1_102 ( .A(\imm[22] ), .Y(_abc_4635_new_n995_));
INVX1 INVX1_103 ( .A(_abc_4635_new_n997_), .Y(_abc_4635_new_n998_));
INVX1 INVX1_104 ( .A(\pc[23] ), .Y(_abc_4635_new_n1003_));
INVX1 INVX1_105 ( .A(_abc_4635_new_n1014_), .Y(_abc_4635_new_n1015_));
INVX1 INVX1_106 ( .A(\rs1[24] ), .Y(_abc_4635_new_n1023_));
INVX1 INVX1_107 ( .A(\imm[24] ), .Y(_abc_4635_new_n1024_));
INVX1 INVX1_108 ( .A(\rs1[26] ), .Y(_abc_4635_new_n1047_));
INVX1 INVX1_109 ( .A(\imm[26] ), .Y(_abc_4635_new_n1048_));
INVX1 INVX1_11 ( .A(_abc_4635_new_n386_), .Y(_abc_4635_new_n387_));
INVX1 INVX1_110 ( .A(_abc_4635_new_n1058_), .Y(_abc_4635_new_n1059_));
INVX1 INVX1_111 ( .A(_abc_4635_new_n1066_), .Y(_abc_4635_new_n1067_));
INVX1 INVX1_112 ( .A(_abc_4635_new_n1049_), .Y(_abc_4635_new_n1069_));
INVX1 INVX1_113 ( .A(\rs1[28] ), .Y(_abc_4635_new_n1074_));
INVX1 INVX1_114 ( .A(\imm[28] ), .Y(_abc_4635_new_n1075_));
INVX1 INVX1_115 ( .A(_abc_4635_new_n1084_), .Y(_abc_4635_new_n1085_));
INVX1 INVX1_116 ( .A(_abc_4635_new_n1091_), .Y(_abc_4635_new_n1092_));
INVX1 INVX1_117 ( .A(_abc_4635_new_n1076_), .Y(_abc_4635_new_n1093_));
INVX1 INVX1_118 ( .A(_abc_4635_new_n1098_), .Y(_abc_4635_new_n1099_));
INVX1 INVX1_119 ( .A(_abc_4635_new_n1107_), .Y(_abc_4635_new_n1110_));
INVX1 INVX1_12 ( .A(_abc_4635_new_n388_), .Y(_abc_4635_new_n389_));
INVX1 INVX1_120 ( .A(_abc_4635_new_n1119_), .Y(ARvalid));
INVX1 INVX1_13 ( .A(state_6_), .Y(_abc_4635_new_n392_));
INVX1 INVX1_14 ( .A(state_2_), .Y(_abc_4635_new_n400_));
INVX1 INVX1_15 ( .A(state_5_), .Y(_abc_4635_new_n401_));
INVX1 INVX1_16 ( .A(state_4_), .Y(_abc_4635_new_n404_));
INVX1 INVX1_17 ( .A(_abc_4635_new_n376_), .Y(_abc_4635_new_n412_));
INVX1 INVX1_18 ( .A(_abc_4635_new_n399_), .Y(_abc_4635_new_n418_));
INVX1 INVX1_19 ( .A(state_1_), .Y(_abc_4635_new_n421_));
INVX1 INVX1_2 ( .A(state_3_), .Y(_abc_4635_new_n362_));
INVX1 INVX1_20 ( .A(_abc_4635_new_n423_), .Y(_abc_4635_new_n424_));
INVX1 INVX1_21 ( .A(_abc_4635_new_n428_), .Y(_abc_4635_new_n429_));
INVX1 INVX1_22 ( .A(done), .Y(busy));
INVX1 INVX1_23 ( .A(_abc_4635_new_n433_), .Y(_abc_4635_new_n434_));
INVX1 INVX1_24 ( .A(_abc_4635_new_n436_), .Y(_abc_4635_new_n437_));
INVX1 INVX1_25 ( .A(\wordsize[0] ), .Y(_abc_4635_new_n444_));
INVX1 INVX1_26 ( .A(_abc_4635_new_n445_), .Y(_abc_4635_new_n446_));
INVX1 INVX1_27 ( .A(\wordsize[1] ), .Y(_abc_4635_new_n448_));
INVX1 INVX1_28 ( .A(_abc_4635_new_n441_), .Y(_abc_4635_new_n456_));
INVX1 INVX1_29 ( .A(_abc_4635_new_n453_), .Y(_abc_4635_new_n457_));
INVX1 INVX1_3 ( .A(resetn), .Y(_abc_4635_new_n366_));
INVX1 INVX1_30 ( .A(\rs2[0] ), .Y(_abc_4635_new_n462_));
INVX1 INVX1_31 ( .A(\rs2[1] ), .Y(_abc_4635_new_n464_));
INVX1 INVX1_32 ( .A(\rs2[2] ), .Y(_abc_4635_new_n466_));
INVX1 INVX1_33 ( .A(\rs2[3] ), .Y(_abc_4635_new_n468_));
INVX1 INVX1_34 ( .A(\rs2[4] ), .Y(_abc_4635_new_n470_));
INVX1 INVX1_35 ( .A(\rs2[5] ), .Y(_abc_4635_new_n472_));
INVX1 INVX1_36 ( .A(\rs2[6] ), .Y(_abc_4635_new_n474_));
INVX1 INVX1_37 ( .A(\rs2[7] ), .Y(_abc_4635_new_n476_));
INVX1 INVX1_38 ( .A(_abc_4635_new_n449_), .Y(_abc_4635_new_n478_));
INVX1 INVX1_39 ( .A(\inst[0] ), .Y(_abc_4635_new_n536_));
INVX1 INVX1_4 ( .A(AWready), .Y(_abc_4635_new_n367_));
INVX1 INVX1_40 ( .A(\inst[1] ), .Y(_abc_4635_new_n541_));
INVX1 INVX1_41 ( .A(\inst[2] ), .Y(_abc_4635_new_n544_));
INVX1 INVX1_42 ( .A(\inst[3] ), .Y(_abc_4635_new_n547_));
INVX1 INVX1_43 ( .A(\inst[4] ), .Y(_abc_4635_new_n550_));
INVX1 INVX1_44 ( .A(\inst[5] ), .Y(_abc_4635_new_n553_));
INVX1 INVX1_45 ( .A(\inst[6] ), .Y(_abc_4635_new_n556_));
INVX1 INVX1_46 ( .A(\inst[7] ), .Y(_abc_4635_new_n559_));
INVX1 INVX1_47 ( .A(\inst[8] ), .Y(_abc_4635_new_n562_));
INVX1 INVX1_48 ( .A(\inst[9] ), .Y(_abc_4635_new_n565_));
INVX1 INVX1_49 ( .A(\inst[10] ), .Y(_abc_4635_new_n568_));
INVX1 INVX1_5 ( .A(enable), .Y(_abc_4635_new_n371_));
INVX1 INVX1_50 ( .A(\inst[11] ), .Y(_abc_4635_new_n571_));
INVX1 INVX1_51 ( .A(\inst[12] ), .Y(_abc_4635_new_n574_));
INVX1 INVX1_52 ( .A(\inst[13] ), .Y(_abc_4635_new_n577_));
INVX1 INVX1_53 ( .A(\inst[14] ), .Y(_abc_4635_new_n580_));
INVX1 INVX1_54 ( .A(\inst[15] ), .Y(_abc_4635_new_n583_));
INVX1 INVX1_55 ( .A(\inst[16] ), .Y(_abc_4635_new_n586_));
INVX1 INVX1_56 ( .A(\inst[17] ), .Y(_abc_4635_new_n589_));
INVX1 INVX1_57 ( .A(\inst[18] ), .Y(_abc_4635_new_n592_));
INVX1 INVX1_58 ( .A(\inst[19] ), .Y(_abc_4635_new_n595_));
INVX1 INVX1_59 ( .A(\inst[20] ), .Y(_abc_4635_new_n598_));
INVX1 INVX1_6 ( .A(_abc_4635_new_n372_), .Y(_abc_4635_new_n374_));
INVX1 INVX1_60 ( .A(\inst[21] ), .Y(_abc_4635_new_n601_));
INVX1 INVX1_61 ( .A(\inst[22] ), .Y(_abc_4635_new_n604_));
INVX1 INVX1_62 ( .A(\inst[23] ), .Y(_abc_4635_new_n607_));
INVX1 INVX1_63 ( .A(\inst[24] ), .Y(_abc_4635_new_n610_));
INVX1 INVX1_64 ( .A(\inst[25] ), .Y(_abc_4635_new_n613_));
INVX1 INVX1_65 ( .A(\inst[26] ), .Y(_abc_4635_new_n616_));
INVX1 INVX1_66 ( .A(\inst[27] ), .Y(_abc_4635_new_n619_));
INVX1 INVX1_67 ( .A(\inst[28] ), .Y(_abc_4635_new_n622_));
INVX1 INVX1_68 ( .A(\inst[29] ), .Y(_abc_4635_new_n625_));
INVX1 INVX1_69 ( .A(\inst[30] ), .Y(_abc_4635_new_n628_));
INVX1 INVX1_7 ( .A(Bvalid), .Y(_abc_4635_new_n379_));
INVX1 INVX1_70 ( .A(\inst[31] ), .Y(_abc_4635_new_n631_));
INVX1 INVX1_71 ( .A(_abc_4635_new_n479_), .Y(_abc_4635_new_n634_));
INVX1 INVX1_72 ( .A(\W_R[1] ), .Y(_abc_4635_new_n639_));
INVX1 INVX1_73 ( .A(_abc_4635_new_n640_), .Y(_abc_4635_new_n641_));
INVX1 INVX1_74 ( .A(_abc_4635_new_n432_), .Y(_abc_4635_new_n642_));
INVX1 INVX1_75 ( .A(\Rdata_mem[1] ), .Y(_abc_4635_new_n655_));
INVX1 INVX1_76 ( .A(\Rdata_mem[2] ), .Y(_abc_4635_new_n665_));
INVX1 INVX1_77 ( .A(\Rdata_mem[3] ), .Y(_abc_4635_new_n675_));
INVX1 INVX1_78 ( .A(\Rdata_mem[6] ), .Y(_abc_4635_new_n699_));
INVX1 INVX1_79 ( .A(\Rdata_mem[23] ), .Y(_abc_4635_new_n705_));
INVX1 INVX1_8 ( .A(ARready), .Y(_abc_4635_new_n382_));
INVX1 INVX1_80 ( .A(_abc_4635_new_n443_), .Y(_abc_4635_new_n710_));
INVX1 INVX1_81 ( .A(_abc_4635_new_n788_), .Y(_abc_4635_new_n795_));
INVX1 INVX1_82 ( .A(_abc_4635_new_n797_), .Y(_abc_4635_new_n804_));
INVX1 INVX1_83 ( .A(\rs1[6] ), .Y(_abc_4635_new_n825_));
INVX1 INVX1_84 ( .A(\imm[6] ), .Y(_abc_4635_new_n826_));
INVX1 INVX1_85 ( .A(_abc_4635_new_n840_), .Y(_abc_4635_new_n845_));
INVX1 INVX1_86 ( .A(_abc_4635_new_n875_), .Y(_abc_4635_new_n876_));
INVX1 INVX1_87 ( .A(_abc_4635_new_n890_), .Y(_abc_4635_new_n905_));
INVX1 INVX1_88 ( .A(_abc_4635_new_n899_), .Y(_abc_4635_new_n906_));
INVX1 INVX1_89 ( .A(_abc_4635_new_n907_), .Y(_abc_4635_new_n908_));
INVX1 INVX1_9 ( .A(Rvalid), .Y(_abc_4635_new_n383_));
INVX1 INVX1_90 ( .A(_abc_4635_new_n932_), .Y(_abc_4635_new_n933_));
INVX1 INVX1_91 ( .A(_abc_4635_new_n930_), .Y(_abc_4635_new_n937_));
INVX1 INVX1_92 ( .A(\rs1[17] ), .Y(_abc_4635_new_n944_));
INVX1 INVX1_93 ( .A(\imm[17] ), .Y(_abc_4635_new_n945_));
INVX1 INVX1_94 ( .A(_abc_4635_new_n947_), .Y(_abc_4635_new_n948_));
INVX1 INVX1_95 ( .A(_abc_4635_new_n951_), .Y(_abc_4635_new_n952_));
INVX1 INVX1_96 ( .A(_abc_4635_new_n954_), .Y(_abc_4635_new_n955_));
INVX1 INVX1_97 ( .A(_abc_4635_new_n967_), .Y(_abc_4635_new_n970_));
INVX1 INVX1_98 ( .A(_abc_4635_new_n971_), .Y(_abc_4635_new_n972_));
INVX1 INVX1_99 ( .A(_abc_4635_new_n988_), .Y(_abc_4635_new_n989_));
MUX2X1 MUX2X1_1 ( .A(\Rdata_mem[8] ), .B(\Rdata_mem[24] ), .S(_abc_4635_new_n441_), .Y(_abc_4635_new_n644_));
MUX2X1 MUX2X1_2 ( .A(\Rdata_mem[9] ), .B(\Rdata_mem[25] ), .S(_abc_4635_new_n441_), .Y(_abc_4635_new_n651_));
MUX2X1 MUX2X1_3 ( .A(\Rdata_mem[10] ), .B(\Rdata_mem[26] ), .S(_abc_4635_new_n441_), .Y(_abc_4635_new_n661_));
MUX2X1 MUX2X1_4 ( .A(\Rdata_mem[11] ), .B(\Rdata_mem[27] ), .S(_abc_4635_new_n441_), .Y(_abc_4635_new_n671_));
MUX2X1 MUX2X1_5 ( .A(\Rdata_mem[12] ), .B(\Rdata_mem[28] ), .S(_abc_4635_new_n441_), .Y(_abc_4635_new_n682_));
MUX2X1 MUX2X1_6 ( .A(\Rdata_mem[13] ), .B(\Rdata_mem[29] ), .S(_abc_4635_new_n441_), .Y(_abc_4635_new_n689_));
MUX2X1 MUX2X1_7 ( .A(\Rdata_mem[14] ), .B(\Rdata_mem[30] ), .S(_abc_4635_new_n441_), .Y(_abc_4635_new_n695_));
NAND2X1 NAND2X1_1 ( .A(resetn), .B(_abc_4635_new_n364_), .Y(_abc_4635_new_n365_));
NAND2X1 NAND2X1_10 ( .A(state_5_), .B(_abc_4635_new_n383_), .Y(_abc_4635_new_n416_));
NAND2X1 NAND2X1_100 ( .A(_abc_4635_new_n974_), .B(_abc_4635_new_n975_), .Y(_abc_4635_new_n976_));
NAND2X1 NAND2X1_101 ( .A(\rs1[21] ), .B(\imm[21] ), .Y(_abc_4635_new_n981_));
NAND2X1 NAND2X1_102 ( .A(_abc_4635_new_n981_), .B(_abc_4635_new_n982_), .Y(_abc_4635_new_n983_));
NAND2X1 NAND2X1_103 ( .A(\W_R[1] ), .B(\pc[21] ), .Y(_abc_4635_new_n985_));
NAND2X1 NAND2X1_104 ( .A(\W_R[1] ), .B(\pc[22] ), .Y(_abc_4635_new_n987_));
NAND2X1 NAND2X1_105 ( .A(\rs1[22] ), .B(\imm[22] ), .Y(_abc_4635_new_n993_));
NAND2X1 NAND2X1_106 ( .A(_abc_4635_new_n994_), .B(_abc_4635_new_n995_), .Y(_abc_4635_new_n996_));
NAND2X1 NAND2X1_107 ( .A(_abc_4635_new_n993_), .B(_abc_4635_new_n996_), .Y(_abc_4635_new_n997_));
NAND2X1 NAND2X1_108 ( .A(_abc_4635_new_n998_), .B(_abc_4635_new_n992_), .Y(_abc_4635_new_n1000_));
NAND2X1 NAND2X1_109 ( .A(_abc_4635_new_n639_), .B(_abc_4635_new_n1000_), .Y(_abc_4635_new_n1001_));
NAND2X1 NAND2X1_11 ( .A(\rs1[0] ), .B(\imm[0] ), .Y(_abc_4635_new_n433_));
NAND2X1 NAND2X1_110 ( .A(\W_R[1] ), .B(\pc[24] ), .Y(_abc_4635_new_n1012_));
NAND2X1 NAND2X1_111 ( .A(_abc_4635_new_n969_), .B(_abc_4635_new_n1014_), .Y(_abc_4635_new_n1017_));
NAND2X1 NAND2X1_112 ( .A(_abc_4635_new_n988_), .B(_abc_4635_new_n1013_), .Y(_abc_4635_new_n1018_));
NAND2X1 NAND2X1_113 ( .A(_abc_4635_new_n1014_), .B(_abc_4635_new_n972_), .Y(_abc_4635_new_n1030_));
NAND2X1 NAND2X1_114 ( .A(_abc_4635_new_n1027_), .B(_abc_4635_new_n1033_), .Y(_abc_4635_new_n1034_));
NAND2X1 NAND2X1_115 ( .A(\W_R[1] ), .B(\pc[25] ), .Y(_abc_4635_new_n1041_));
NAND2X1 NAND2X1_116 ( .A(\W_R[1] ), .B(\pc[26] ), .Y(_abc_4635_new_n1043_));
NAND2X1 NAND2X1_117 ( .A(_abc_4635_new_n1039_), .B(_abc_4635_new_n1032_), .Y(_abc_4635_new_n1045_));
NAND2X1 NAND2X1_118 ( .A(_abc_4635_new_n1051_), .B(_abc_4635_new_n1046_), .Y(_abc_4635_new_n1053_));
NAND2X1 NAND2X1_119 ( .A(_abc_4635_new_n639_), .B(_abc_4635_new_n1053_), .Y(_abc_4635_new_n1054_));
NAND2X1 NAND2X1_12 ( .A(\rs1[1] ), .B(\imm[1] ), .Y(_abc_4635_new_n436_));
NAND2X1 NAND2X1_120 ( .A(\rs1[27] ), .B(\imm[27] ), .Y(_abc_4635_new_n1058_));
NAND2X1 NAND2X1_121 ( .A(\W_R[1] ), .B(\pc[27] ), .Y(_abc_4635_new_n1062_));
NAND2X1 NAND2X1_122 ( .A(\W_R[1] ), .B(\pc[28] ), .Y(_abc_4635_new_n1064_));
NAND2X1 NAND2X1_123 ( .A(_abc_4635_new_n1060_), .B(_abc_4635_new_n1051_), .Y(_abc_4635_new_n1065_));
NAND2X1 NAND2X1_124 ( .A(_abc_4635_new_n1077_), .B(_abc_4635_new_n1072_), .Y(_abc_4635_new_n1079_));
NAND2X1 NAND2X1_125 ( .A(_abc_4635_new_n639_), .B(_abc_4635_new_n1079_), .Y(_abc_4635_new_n1080_));
NAND2X1 NAND2X1_126 ( .A(\rs1[29] ), .B(\imm[29] ), .Y(_abc_4635_new_n1084_));
NAND2X1 NAND2X1_127 ( .A(\W_R[1] ), .B(\pc[29] ), .Y(_abc_4635_new_n1088_));
NAND2X1 NAND2X1_128 ( .A(\W_R[1] ), .B(\pc[30] ), .Y(_abc_4635_new_n1090_));
NAND2X1 NAND2X1_129 ( .A(_abc_4635_new_n1086_), .B(_abc_4635_new_n1077_), .Y(_abc_4635_new_n1091_));
NAND2X1 NAND2X1_13 ( .A(_abc_4635_new_n434_), .B(_abc_4635_new_n438_), .Y(_abc_4635_new_n439_));
NAND2X1 NAND2X1_130 ( .A(\rs1[30] ), .B(\imm[30] ), .Y(_abc_4635_new_n1097_));
NAND2X1 NAND2X1_131 ( .A(_abc_4635_new_n1099_), .B(_abc_4635_new_n1095_), .Y(_abc_4635_new_n1100_));
NAND2X1 NAND2X1_132 ( .A(_abc_4635_new_n1100_), .B(_abc_4635_new_n1103_), .Y(_abc_4635_new_n1104_));
NAND2X1 NAND2X1_133 ( .A(\W_R[1] ), .B(\pc[31] ), .Y(_abc_4635_new_n1106_));
NAND2X1 NAND2X1_134 ( .A(_abc_4635_new_n1110_), .B(_abc_4635_new_n1109_), .Y(_abc_4635_new_n1111_));
NAND2X1 NAND2X1_135 ( .A(_abc_4635_new_n1106_), .B(_abc_4635_new_n1112_), .Y(\ARdata[31] ));
NAND2X1 NAND2X1_136 ( .A(_abc_4635_new_n404_), .B(_abc_4635_new_n362_), .Y(_abc_4635_new_n1116_));
NAND2X1 NAND2X1_14 ( .A(_abc_4635_new_n440_), .B(_abc_4635_new_n439_), .Y(_abc_4635_new_n441_));
NAND2X1 NAND2X1_15 ( .A(\rs2[8] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n480_));
NAND2X1 NAND2X1_16 ( .A(\rs2[9] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n483_));
NAND2X1 NAND2X1_17 ( .A(\rs2[10] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n486_));
NAND2X1 NAND2X1_18 ( .A(\rs2[11] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n489_));
NAND2X1 NAND2X1_19 ( .A(\rs2[12] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n492_));
NAND2X1 NAND2X1_2 ( .A(_abc_4635_new_n367_), .B(_abc_4635_new_n361_), .Y(_abc_4635_new_n370_));
NAND2X1 NAND2X1_20 ( .A(\rs2[13] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n495_));
NAND2X1 NAND2X1_21 ( .A(\rs2[14] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n498_));
NAND2X1 NAND2X1_22 ( .A(\rs2[15] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n501_));
NAND2X1 NAND2X1_23 ( .A(\rs2[24] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n520_));
NAND2X1 NAND2X1_24 ( .A(\rs2[25] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n522_));
NAND2X1 NAND2X1_25 ( .A(\rs2[26] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n524_));
NAND2X1 NAND2X1_26 ( .A(\rs2[27] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n526_));
NAND2X1 NAND2X1_27 ( .A(\rs2[28] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n528_));
NAND2X1 NAND2X1_28 ( .A(\rs2[29] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n530_));
NAND2X1 NAND2X1_29 ( .A(\rs2[30] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n532_));
NAND2X1 NAND2X1_3 ( .A(state_0_), .B(_abc_4635_new_n375_), .Y(_abc_4635_new_n376_));
NAND2X1 NAND2X1_30 ( .A(\rs2[31] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n534_));
NAND2X1 NAND2X1_31 ( .A(\W_R[1] ), .B(_abc_4635_new_n537_), .Y(_abc_4635_new_n538_));
NAND2X1 NAND2X1_32 ( .A(\W_R[0] ), .B(_abc_4635_new_n639_), .Y(_abc_4635_new_n640_));
NAND2X1 NAND2X1_33 ( .A(\Rdata_mem[15] ), .B(_abc_4635_new_n441_), .Y(_abc_4635_new_n711_));
NAND2X1 NAND2X1_34 ( .A(\Rdata_mem[31] ), .B(_abc_4635_new_n456_), .Y(_abc_4635_new_n712_));
NAND2X1 NAND2X1_35 ( .A(\Rdata_mem[16] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n743_));
NAND2X1 NAND2X1_36 ( .A(\Rdata_mem[17] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n746_));
NAND2X1 NAND2X1_37 ( .A(\Rdata_mem[18] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n748_));
NAND2X1 NAND2X1_38 ( .A(\Rdata_mem[19] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n750_));
NAND2X1 NAND2X1_39 ( .A(\Rdata_mem[20] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n752_));
NAND2X1 NAND2X1_4 ( .A(state_0_), .B(_abc_4635_new_n387_), .Y(_abc_4635_new_n388_));
NAND2X1 NAND2X1_40 ( .A(\Rdata_mem[21] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n754_));
NAND2X1 NAND2X1_41 ( .A(\Rdata_mem[22] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n756_));
NAND2X1 NAND2X1_42 ( .A(\Rdata_mem[24] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n760_));
NAND2X1 NAND2X1_43 ( .A(\Rdata_mem[25] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n762_));
NAND2X1 NAND2X1_44 ( .A(\Rdata_mem[26] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n764_));
NAND2X1 NAND2X1_45 ( .A(\Rdata_mem[27] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n766_));
NAND2X1 NAND2X1_46 ( .A(\Rdata_mem[28] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n768_));
NAND2X1 NAND2X1_47 ( .A(\Rdata_mem[29] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n770_));
NAND2X1 NAND2X1_48 ( .A(\Rdata_mem[30] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n772_));
NAND2X1 NAND2X1_49 ( .A(\Rdata_mem[31] ), .B(_abc_4635_new_n479_), .Y(_abc_4635_new_n774_));
NAND2X1 NAND2X1_5 ( .A(Wready), .B(_abc_4635_new_n395_), .Y(_abc_4635_new_n396_));
NAND2X1 NAND2X1_50 ( .A(\W_R[1] ), .B(\pc[0] ), .Y(_abc_4635_new_n776_));
NAND2X1 NAND2X1_51 ( .A(\W_R[1] ), .B(\pc[1] ), .Y(_abc_4635_new_n778_));
NAND2X1 NAND2X1_52 ( .A(\W_R[1] ), .B(\pc[2] ), .Y(_abc_4635_new_n785_));
NAND2X1 NAND2X1_53 ( .A(\W_R[1] ), .B(\pc[3] ), .Y(_abc_4635_new_n792_));
NAND2X1 NAND2X1_54 ( .A(_abc_4635_new_n796_), .B(_abc_4635_new_n794_), .Y(_abc_4635_new_n797_));
NAND2X1 NAND2X1_55 ( .A(\W_R[1] ), .B(\pc[4] ), .Y(_abc_4635_new_n802_));
NAND2X1 NAND2X1_56 ( .A(\rs1[4] ), .B(\imm[4] ), .Y(_abc_4635_new_n805_));
NAND2X1 NAND2X1_57 ( .A(\W_R[1] ), .B(\pc[5] ), .Y(_abc_4635_new_n811_));
NAND2X1 NAND2X1_58 ( .A(\W_R[1] ), .B(\pc[6] ), .Y(_abc_4635_new_n813_));
NAND2X1 NAND2X1_59 ( .A(_abc_4635_new_n800_), .B(_abc_4635_new_n809_), .Y(_abc_4635_new_n816_));
NAND2X1 NAND2X1_6 ( .A(state_0_), .B(_abc_4635_new_n397_), .Y(_abc_4635_new_n398_));
NAND2X1 NAND2X1_60 ( .A(_abc_4635_new_n820_), .B(_abc_4635_new_n817_), .Y(_abc_4635_new_n822_));
NAND2X1 NAND2X1_61 ( .A(_abc_4635_new_n639_), .B(_abc_4635_new_n822_), .Y(_abc_4635_new_n823_));
NAND2X1 NAND2X1_62 ( .A(\W_R[1] ), .B(\pc[7] ), .Y(_abc_4635_new_n832_));
NAND2X1 NAND2X1_63 ( .A(\W_R[1] ), .B(\pc[8] ), .Y(_abc_4635_new_n834_));
NAND2X1 NAND2X1_64 ( .A(_abc_4635_new_n820_), .B(_abc_4635_new_n830_), .Y(_abc_4635_new_n835_));
NAND2X1 NAND2X1_65 ( .A(\W_R[1] ), .B(\pc[9] ), .Y(_abc_4635_new_n851_));
NAND2X1 NAND2X1_66 ( .A(\W_R[1] ), .B(\pc[10] ), .Y(_abc_4635_new_n853_));
NAND2X1 NAND2X1_67 ( .A(_abc_4635_new_n842_), .B(_abc_4635_new_n849_), .Y(_abc_4635_new_n856_));
NAND2X1 NAND2X1_68 ( .A(_abc_4635_new_n860_), .B(_abc_4635_new_n857_), .Y(_abc_4635_new_n862_));
NAND2X1 NAND2X1_69 ( .A(_abc_4635_new_n639_), .B(_abc_4635_new_n862_), .Y(_abc_4635_new_n863_));
NAND2X1 NAND2X1_7 ( .A(_abc_4635_new_n368_), .B(_abc_4635_new_n377_), .Y(_abc_4635_new_n408_));
NAND2X1 NAND2X1_70 ( .A(\W_R[1] ), .B(\pc[11] ), .Y(_abc_4635_new_n870_));
NAND2X1 NAND2X1_71 ( .A(\W_R[1] ), .B(\pc[12] ), .Y(_abc_4635_new_n872_));
NAND2X1 NAND2X1_72 ( .A(_abc_4635_new_n860_), .B(_abc_4635_new_n868_), .Y(_abc_4635_new_n873_));
NAND2X1 NAND2X1_73 ( .A(_abc_4635_new_n805_), .B(_abc_4635_new_n877_), .Y(_abc_4635_new_n878_));
NAND2X1 NAND2X1_74 ( .A(\rs1[5] ), .B(\imm[5] ), .Y(_abc_4635_new_n879_));
NAND2X1 NAND2X1_75 ( .A(_abc_4635_new_n879_), .B(_abc_4635_new_n814_), .Y(_abc_4635_new_n880_));
NAND2X1 NAND2X1_76 ( .A(\rs1[6] ), .B(_abc_4635_new_n826_), .Y(_abc_4635_new_n882_));
NAND2X1 NAND2X1_77 ( .A(\imm[6] ), .B(_abc_4635_new_n825_), .Y(_abc_4635_new_n883_));
NAND2X1 NAND2X1_78 ( .A(_abc_4635_new_n885_), .B(_abc_4635_new_n881_), .Y(_abc_4635_new_n886_));
NAND2X1 NAND2X1_79 ( .A(_abc_4635_new_n876_), .B(_abc_4635_new_n889_), .Y(_abc_4635_new_n890_));
NAND2X1 NAND2X1_8 ( .A(resetn), .B(_abc_4635_new_n409_), .Y(_abc_4635_new_n410_));
NAND2X1 NAND2X1_80 ( .A(_abc_4635_new_n891_), .B(_abc_4635_new_n890_), .Y(_abc_4635_new_n893_));
NAND2X1 NAND2X1_81 ( .A(_abc_4635_new_n639_), .B(_abc_4635_new_n893_), .Y(_abc_4635_new_n894_));
NAND2X1 NAND2X1_82 ( .A(\rs1[12] ), .B(\imm[12] ), .Y(_abc_4635_new_n896_));
NAND2X1 NAND2X1_83 ( .A(_abc_4635_new_n896_), .B(_abc_4635_new_n893_), .Y(_abc_4635_new_n897_));
NAND2X1 NAND2X1_84 ( .A(\W_R[1] ), .B(\pc[13] ), .Y(_abc_4635_new_n902_));
NAND2X1 NAND2X1_85 ( .A(\W_R[1] ), .B(\pc[14] ), .Y(_abc_4635_new_n904_));
NAND2X1 NAND2X1_86 ( .A(_abc_4635_new_n900_), .B(_abc_4635_new_n891_), .Y(_abc_4635_new_n909_));
NAND2X1 NAND2X1_87 ( .A(\W_R[1] ), .B(\pc[15] ), .Y(_abc_4635_new_n921_));
NAND2X1 NAND2X1_88 ( .A(\W_R[1] ), .B(\pc[16] ), .Y(_abc_4635_new_n923_));
NAND2X1 NAND2X1_89 ( .A(_abc_4635_new_n913_), .B(_abc_4635_new_n919_), .Y(_abc_4635_new_n924_));
NAND2X1 NAND2X1_9 ( .A(ARready), .B(_abc_4635_new_n383_), .Y(_abc_4635_new_n415_));
NAND2X1 NAND2X1_90 ( .A(_abc_4635_new_n888_), .B(_abc_4635_new_n925_), .Y(_abc_4635_new_n926_));
NAND2X1 NAND2X1_91 ( .A(\rs1[16] ), .B(\imm[16] ), .Y(_abc_4635_new_n932_));
NAND2X1 NAND2X1_92 ( .A(\W_R[1] ), .B(\pc[17] ), .Y(_abc_4635_new_n941_));
NAND2X1 NAND2X1_93 ( .A(\W_R[1] ), .B(\pc[18] ), .Y(_abc_4635_new_n943_));
NAND2X1 NAND2X1_94 ( .A(\rs1[18] ), .B(\imm[18] ), .Y(_abc_4635_new_n951_));
NAND2X1 NAND2X1_95 ( .A(\W_R[1] ), .B(\pc[19] ), .Y(_abc_4635_new_n964_));
NAND2X1 NAND2X1_96 ( .A(\W_R[1] ), .B(\pc[20] ), .Y(_abc_4635_new_n966_));
NAND2X1 NAND2X1_97 ( .A(_abc_4635_new_n962_), .B(_abc_4635_new_n954_), .Y(_abc_4635_new_n967_));
NAND2X1 NAND2X1_98 ( .A(_abc_4635_new_n949_), .B(_abc_4635_new_n970_), .Y(_abc_4635_new_n971_));
NAND2X1 NAND2X1_99 ( .A(\rs1[20] ), .B(\imm[20] ), .Y(_abc_4635_new_n974_));
NAND3X1 NAND3X1_1 ( .A(AWready), .B(Wready), .C(_abc_4635_new_n379_), .Y(_abc_4635_new_n380_));
NAND3X1 NAND3X1_2 ( .A(_abc_4635_new_n398_), .B(_abc_4635_new_n403_), .C(_abc_4635_new_n406_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_0_));
NAND3X1 NAND3X1_3 ( .A(_abc_4635_new_n783_), .B(_abc_4635_new_n780_), .C(_abc_4635_new_n790_), .Y(_abc_4635_new_n794_));
NAND3X1 NAND3X1_4 ( .A(_abc_4635_new_n1018_), .B(_abc_4635_new_n1020_), .C(_abc_4635_new_n1017_), .Y(_abc_4635_new_n1021_));
NAND3X1 NAND3X1_5 ( .A(_abc_4635_new_n1097_), .B(_abc_4635_new_n1107_), .C(_abc_4635_new_n1103_), .Y(_abc_4635_new_n1108_));
NAND3X1 NAND3X1_6 ( .A(_abc_4635_new_n639_), .B(_abc_4635_new_n1108_), .C(_abc_4635_new_n1111_), .Y(_abc_4635_new_n1112_));
NOR2X1 NOR2X1_1 ( .A(Wready), .B(_abc_4635_new_n367_), .Y(_abc_4635_new_n368_));
NOR2X1 NOR2X1_10 ( .A(_abc_4635_new_n419_), .B(_abc_4635_new_n397_), .Y(_abc_4635_new_n420_));
NOR2X1 NOR2X1_100 ( .A(\rs1[26] ), .B(\imm[26] ), .Y(_abc_4635_new_n1050_));
NOR2X1 NOR2X1_101 ( .A(_abc_4635_new_n1050_), .B(_abc_4635_new_n1049_), .Y(_abc_4635_new_n1051_));
NOR2X1 NOR2X1_102 ( .A(_abc_4635_new_n1051_), .B(_abc_4635_new_n1046_), .Y(_abc_4635_new_n1052_));
NOR2X1 NOR2X1_103 ( .A(\rs1[27] ), .B(\imm[27] ), .Y(_abc_4635_new_n1057_));
NOR2X1 NOR2X1_104 ( .A(_abc_4635_new_n1057_), .B(_abc_4635_new_n1059_), .Y(_abc_4635_new_n1060_));
NOR2X1 NOR2X1_105 ( .A(_abc_4635_new_n1065_), .B(_abc_4635_new_n1045_), .Y(_abc_4635_new_n1066_));
NOR2X1 NOR2X1_106 ( .A(_abc_4635_new_n1044_), .B(_abc_4635_new_n1065_), .Y(_abc_4635_new_n1068_));
NOR2X1 NOR2X1_107 ( .A(_abc_4635_new_n1070_), .B(_abc_4635_new_n1068_), .Y(_abc_4635_new_n1071_));
NOR2X1 NOR2X1_108 ( .A(\rs1[28] ), .B(\imm[28] ), .Y(_abc_4635_new_n1073_));
NOR2X1 NOR2X1_109 ( .A(_abc_4635_new_n1074_), .B(_abc_4635_new_n1075_), .Y(_abc_4635_new_n1076_));
NOR2X1 NOR2X1_11 ( .A(_abc_4635_new_n422_), .B(_abc_4635_new_n385_), .Y(_abc_4635_new_n423_));
NOR2X1 NOR2X1_110 ( .A(_abc_4635_new_n1073_), .B(_abc_4635_new_n1076_), .Y(_abc_4635_new_n1077_));
NOR2X1 NOR2X1_111 ( .A(_abc_4635_new_n1077_), .B(_abc_4635_new_n1072_), .Y(_abc_4635_new_n1078_));
NOR2X1 NOR2X1_112 ( .A(\rs1[29] ), .B(\imm[29] ), .Y(_abc_4635_new_n1083_));
NOR2X1 NOR2X1_113 ( .A(_abc_4635_new_n1083_), .B(_abc_4635_new_n1085_), .Y(_abc_4635_new_n1086_));
NOR2X1 NOR2X1_114 ( .A(state_6_), .B(state_1_), .Y(_abc_4635_new_n1115_));
NOR2X1 NOR2X1_115 ( .A(_abc_4635_new_n1116_), .B(_abc_4635_new_n412_), .Y(_abc_4635_new_n1117_));
NOR2X1 NOR2X1_116 ( .A(_abc_4635_new_n366_), .B(_abc_4635_new_n1117_), .Y(Wvalid));
NOR2X1 NOR2X1_12 ( .A(\wordsize[0] ), .B(\wordsize[1] ), .Y(_abc_4635_new_n432_));
NOR2X1 NOR2X1_13 ( .A(\rs1[1] ), .B(\imm[1] ), .Y(_abc_4635_new_n435_));
NOR2X1 NOR2X1_14 ( .A(_abc_4635_new_n435_), .B(_abc_4635_new_n437_), .Y(_abc_4635_new_n438_));
NOR2X1 NOR2X1_15 ( .A(\rs1[0] ), .B(\imm[0] ), .Y(_abc_4635_new_n442_));
NOR2X1 NOR2X1_16 ( .A(\wordsize[1] ), .B(_abc_4635_new_n444_), .Y(_abc_4635_new_n445_));
NOR2X1 NOR2X1_17 ( .A(_abc_4635_new_n446_), .B(_abc_4635_new_n441_), .Y(_abc_4635_new_n447_));
NOR2X1 NOR2X1_18 ( .A(_abc_4635_new_n366_), .B(_abc_4635_new_n374_), .Y(_abc_4635_new_n449_));
NOR2X1 NOR2X1_19 ( .A(_abc_4635_new_n442_), .B(_abc_4635_new_n434_), .Y(_abc_4635_new_n453_));
NOR2X1 NOR2X1_2 ( .A(_abc_4635_new_n366_), .B(_abc_4635_new_n368_), .Y(_abc_4635_new_n369_));
NOR2X1 NOR2X1_20 ( .A(_abc_4635_new_n462_), .B(_abc_4635_new_n450_), .Y(_0Wdata_31_0__0_));
NOR2X1 NOR2X1_21 ( .A(_abc_4635_new_n464_), .B(_abc_4635_new_n450_), .Y(_0Wdata_31_0__1_));
NOR2X1 NOR2X1_22 ( .A(_abc_4635_new_n466_), .B(_abc_4635_new_n450_), .Y(_0Wdata_31_0__2_));
NOR2X1 NOR2X1_23 ( .A(_abc_4635_new_n468_), .B(_abc_4635_new_n450_), .Y(_0Wdata_31_0__3_));
NOR2X1 NOR2X1_24 ( .A(_abc_4635_new_n470_), .B(_abc_4635_new_n450_), .Y(_0Wdata_31_0__4_));
NOR2X1 NOR2X1_25 ( .A(_abc_4635_new_n472_), .B(_abc_4635_new_n450_), .Y(_0Wdata_31_0__5_));
NOR2X1 NOR2X1_26 ( .A(_abc_4635_new_n474_), .B(_abc_4635_new_n450_), .Y(_0Wdata_31_0__6_));
NOR2X1 NOR2X1_27 ( .A(_abc_4635_new_n476_), .B(_abc_4635_new_n450_), .Y(_0Wdata_31_0__7_));
NOR2X1 NOR2X1_28 ( .A(\wordsize[0] ), .B(_abc_4635_new_n448_), .Y(_abc_4635_new_n479_));
NOR2X1 NOR2X1_29 ( .A(_abc_4635_new_n504_), .B(_abc_4635_new_n478_), .Y(_0Wdata_31_0__16_));
NOR2X1 NOR2X1_3 ( .A(\W_R[0] ), .B(\W_R[1] ), .Y(_abc_4635_new_n372_));
NOR2X1 NOR2X1_30 ( .A(_abc_4635_new_n506_), .B(_abc_4635_new_n478_), .Y(_0Wdata_31_0__17_));
NOR2X1 NOR2X1_31 ( .A(_abc_4635_new_n508_), .B(_abc_4635_new_n478_), .Y(_0Wdata_31_0__18_));
NOR2X1 NOR2X1_32 ( .A(_abc_4635_new_n510_), .B(_abc_4635_new_n478_), .Y(_0Wdata_31_0__19_));
NOR2X1 NOR2X1_33 ( .A(_abc_4635_new_n512_), .B(_abc_4635_new_n478_), .Y(_0Wdata_31_0__20_));
NOR2X1 NOR2X1_34 ( .A(_abc_4635_new_n514_), .B(_abc_4635_new_n478_), .Y(_0Wdata_31_0__21_));
NOR2X1 NOR2X1_35 ( .A(_abc_4635_new_n516_), .B(_abc_4635_new_n478_), .Y(_0Wdata_31_0__22_));
NOR2X1 NOR2X1_36 ( .A(_abc_4635_new_n518_), .B(_abc_4635_new_n478_), .Y(_0Wdata_31_0__23_));
NOR2X1 NOR2X1_37 ( .A(_abc_4635_new_n366_), .B(_abc_4635_new_n403_), .Y(_abc_4635_new_n537_));
NOR2X1 NOR2X1_38 ( .A(\W_R[1] ), .B(_abc_4635_new_n371_), .Y(_abc_4635_new_n635_));
NOR2X1 NOR2X1_39 ( .A(_abc_4635_new_n453_), .B(_abc_4635_new_n708_), .Y(_abc_4635_new_n709_));
NOR2X1 NOR2X1_4 ( .A(_abc_4635_new_n371_), .B(_abc_4635_new_n374_), .Y(_abc_4635_new_n375_));
NOR2X1 NOR2X1_40 ( .A(_abc_4635_new_n446_), .B(_abc_4635_new_n644_), .Y(_abc_4635_new_n719_));
NOR2X1 NOR2X1_41 ( .A(_abc_4635_new_n446_), .B(_abc_4635_new_n651_), .Y(_abc_4635_new_n722_));
NOR2X1 NOR2X1_42 ( .A(_abc_4635_new_n446_), .B(_abc_4635_new_n661_), .Y(_abc_4635_new_n725_));
NOR2X1 NOR2X1_43 ( .A(_abc_4635_new_n446_), .B(_abc_4635_new_n671_), .Y(_abc_4635_new_n728_));
NOR2X1 NOR2X1_44 ( .A(_abc_4635_new_n446_), .B(_abc_4635_new_n682_), .Y(_abc_4635_new_n731_));
NOR2X1 NOR2X1_45 ( .A(_abc_4635_new_n446_), .B(_abc_4635_new_n689_), .Y(_abc_4635_new_n734_));
NOR2X1 NOR2X1_46 ( .A(_abc_4635_new_n446_), .B(_abc_4635_new_n695_), .Y(_abc_4635_new_n737_));
NOR2X1 NOR2X1_47 ( .A(\rs1[2] ), .B(\imm[2] ), .Y(_abc_4635_new_n782_));
NOR2X1 NOR2X1_48 ( .A(_abc_4635_new_n782_), .B(_abc_4635_new_n781_), .Y(_abc_4635_new_n783_));
NOR2X1 NOR2X1_49 ( .A(\rs1[3] ), .B(\imm[3] ), .Y(_abc_4635_new_n788_));
NOR2X1 NOR2X1_5 ( .A(_abc_4635_new_n373_), .B(_abc_4635_new_n376_), .Y(_abc_4635_new_n377_));
NOR2X1 NOR2X1_50 ( .A(_abc_4635_new_n788_), .B(_abc_4635_new_n789_), .Y(_abc_4635_new_n790_));
NOR2X1 NOR2X1_51 ( .A(\rs1[4] ), .B(\imm[4] ), .Y(_abc_4635_new_n798_));
NOR2X1 NOR2X1_52 ( .A(_abc_4635_new_n798_), .B(_abc_4635_new_n799_), .Y(_abc_4635_new_n800_));
NOR2X1 NOR2X1_53 ( .A(\rs1[5] ), .B(\imm[5] ), .Y(_abc_4635_new_n807_));
NOR2X1 NOR2X1_54 ( .A(_abc_4635_new_n807_), .B(_abc_4635_new_n808_), .Y(_abc_4635_new_n809_));
NOR2X1 NOR2X1_55 ( .A(\rs1[6] ), .B(\imm[6] ), .Y(_abc_4635_new_n819_));
NOR2X1 NOR2X1_56 ( .A(_abc_4635_new_n819_), .B(_abc_4635_new_n818_), .Y(_abc_4635_new_n820_));
NOR2X1 NOR2X1_57 ( .A(_abc_4635_new_n820_), .B(_abc_4635_new_n817_), .Y(_abc_4635_new_n821_));
NOR2X1 NOR2X1_58 ( .A(\rs1[7] ), .B(\imm[7] ), .Y(_abc_4635_new_n828_));
NOR2X1 NOR2X1_59 ( .A(_abc_4635_new_n828_), .B(_abc_4635_new_n829_), .Y(_abc_4635_new_n830_));
NOR2X1 NOR2X1_6 ( .A(ARready), .B(_abc_4635_new_n390_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_2_));
NOR2X1 NOR2X1_60 ( .A(_abc_4635_new_n816_), .B(_abc_4635_new_n835_), .Y(_abc_4635_new_n836_));
NOR2X1 NOR2X1_61 ( .A(\rs1[8] ), .B(\imm[8] ), .Y(_abc_4635_new_n841_));
NOR2X1 NOR2X1_62 ( .A(_abc_4635_new_n841_), .B(_abc_4635_new_n840_), .Y(_abc_4635_new_n842_));
NOR2X1 NOR2X1_63 ( .A(\rs1[9] ), .B(\imm[9] ), .Y(_abc_4635_new_n847_));
NOR2X1 NOR2X1_64 ( .A(_abc_4635_new_n847_), .B(_abc_4635_new_n848_), .Y(_abc_4635_new_n849_));
NOR2X1 NOR2X1_65 ( .A(\rs1[10] ), .B(\imm[10] ), .Y(_abc_4635_new_n859_));
NOR2X1 NOR2X1_66 ( .A(_abc_4635_new_n859_), .B(_abc_4635_new_n858_), .Y(_abc_4635_new_n860_));
NOR2X1 NOR2X1_67 ( .A(_abc_4635_new_n860_), .B(_abc_4635_new_n857_), .Y(_abc_4635_new_n861_));
NOR2X1 NOR2X1_68 ( .A(\rs1[11] ), .B(\imm[11] ), .Y(_abc_4635_new_n866_));
NOR2X1 NOR2X1_69 ( .A(_abc_4635_new_n866_), .B(_abc_4635_new_n867_), .Y(_abc_4635_new_n868_));
NOR2X1 NOR2X1_7 ( .A(_abc_4635_new_n379_), .B(_abc_4635_new_n367_), .Y(_abc_4635_new_n395_));
NOR2X1 NOR2X1_70 ( .A(_abc_4635_new_n878_), .B(_abc_4635_new_n880_), .Y(_abc_4635_new_n881_));
NOR2X1 NOR2X1_71 ( .A(_abc_4635_new_n856_), .B(_abc_4635_new_n873_), .Y(_abc_4635_new_n888_));
NOR2X1 NOR2X1_72 ( .A(_abc_4635_new_n891_), .B(_abc_4635_new_n890_), .Y(_abc_4635_new_n892_));
NOR2X1 NOR2X1_73 ( .A(\rs1[13] ), .B(\imm[13] ), .Y(_abc_4635_new_n898_));
NOR2X1 NOR2X1_74 ( .A(_abc_4635_new_n898_), .B(_abc_4635_new_n899_), .Y(_abc_4635_new_n900_));
NOR2X1 NOR2X1_75 ( .A(\rs1[14] ), .B(\imm[14] ), .Y(_abc_4635_new_n912_));
NOR2X1 NOR2X1_76 ( .A(_abc_4635_new_n912_), .B(_abc_4635_new_n911_), .Y(_abc_4635_new_n913_));
NOR2X1 NOR2X1_77 ( .A(\rs1[15] ), .B(\imm[15] ), .Y(_abc_4635_new_n917_));
NOR2X1 NOR2X1_78 ( .A(_abc_4635_new_n917_), .B(_abc_4635_new_n918_), .Y(_abc_4635_new_n919_));
NOR2X1 NOR2X1_79 ( .A(_abc_4635_new_n909_), .B(_abc_4635_new_n924_), .Y(_abc_4635_new_n925_));
NOR2X1 NOR2X1_8 ( .A(_abc_4635_new_n382_), .B(_abc_4635_new_n383_), .Y(_abc_4635_new_n399_));
NOR2X1 NOR2X1_80 ( .A(\rs1[16] ), .B(\imm[16] ), .Y(_abc_4635_new_n931_));
NOR2X1 NOR2X1_81 ( .A(_abc_4635_new_n931_), .B(_abc_4635_new_n933_), .Y(_abc_4635_new_n934_));
NOR2X1 NOR2X1_82 ( .A(\rs1[18] ), .B(\imm[18] ), .Y(_abc_4635_new_n953_));
NOR2X1 NOR2X1_83 ( .A(_abc_4635_new_n953_), .B(_abc_4635_new_n952_), .Y(_abc_4635_new_n954_));
NOR2X1 NOR2X1_84 ( .A(\rs1[19] ), .B(\imm[19] ), .Y(_abc_4635_new_n961_));
NOR2X1 NOR2X1_85 ( .A(_abc_4635_new_n961_), .B(_abc_4635_new_n960_), .Y(_abc_4635_new_n962_));
NOR2X1 NOR2X1_86 ( .A(_abc_4635_new_n976_), .B(_abc_4635_new_n983_), .Y(_abc_4635_new_n990_));
NOR2X1 NOR2X1_87 ( .A(_abc_4635_new_n998_), .B(_abc_4635_new_n992_), .Y(_abc_4635_new_n999_));
NOR2X1 NOR2X1_88 ( .A(\rs1[23] ), .B(\imm[23] ), .Y(_abc_4635_new_n1006_));
NOR2X1 NOR2X1_89 ( .A(_abc_4635_new_n1007_), .B(_abc_4635_new_n1004_), .Y(_abc_4635_new_n1009_));
NOR2X1 NOR2X1_9 ( .A(_abc_4635_new_n370_), .B(_abc_4635_new_n413_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_4_));
NOR2X1 NOR2X1_90 ( .A(_abc_4635_new_n997_), .B(_abc_4635_new_n1007_), .Y(_abc_4635_new_n1013_));
NOR2X1 NOR2X1_91 ( .A(_abc_4635_new_n971_), .B(_abc_4635_new_n1015_), .Y(_abc_4635_new_n1016_));
NOR2X1 NOR2X1_92 ( .A(_abc_4635_new_n993_), .B(_abc_4635_new_n1006_), .Y(_abc_4635_new_n1019_));
NOR2X1 NOR2X1_93 ( .A(_abc_4635_new_n1005_), .B(_abc_4635_new_n1019_), .Y(_abc_4635_new_n1020_));
NOR2X1 NOR2X1_94 ( .A(_abc_4635_new_n1023_), .B(_abc_4635_new_n1024_), .Y(_abc_4635_new_n1025_));
NOR2X1 NOR2X1_95 ( .A(\rs1[24] ), .B(\imm[24] ), .Y(_abc_4635_new_n1026_));
NOR2X1 NOR2X1_96 ( .A(_abc_4635_new_n1026_), .B(_abc_4635_new_n1025_), .Y(_abc_4635_new_n1032_));
NOR2X1 NOR2X1_97 ( .A(\rs1[25] ), .B(\imm[25] ), .Y(_abc_4635_new_n1038_));
NOR2X1 NOR2X1_98 ( .A(_abc_4635_new_n1038_), .B(_abc_4635_new_n1037_), .Y(_abc_4635_new_n1039_));
NOR2X1 NOR2X1_99 ( .A(_abc_4635_new_n1047_), .B(_abc_4635_new_n1048_), .Y(_abc_4635_new_n1049_));
OAI21X1 OAI21X1_1 ( .A(_abc_4635_new_n361_), .B(_abc_4635_new_n362_), .C(_abc_4635_new_n363_), .Y(_abc_4635_new_n364_));
OAI21X1 OAI21X1_10 ( .A(Wready), .B(_abc_4635_new_n410_), .C(_abc_4635_new_n408_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_3_));
OAI21X1 OAI21X1_100 ( .A(\W_R[1] ), .B(_abc_4635_new_n810_), .C(_abc_4635_new_n811_), .Y(\ARdata[5] ));
OAI21X1 OAI21X1_101 ( .A(_abc_4635_new_n816_), .B(_abc_4635_new_n804_), .C(_abc_4635_new_n815_), .Y(_abc_4635_new_n817_));
OAI21X1 OAI21X1_102 ( .A(_abc_4635_new_n821_), .B(_abc_4635_new_n823_), .C(_abc_4635_new_n813_), .Y(\ARdata[6] ));
OAI21X1 OAI21X1_103 ( .A(_abc_4635_new_n825_), .B(_abc_4635_new_n826_), .C(_abc_4635_new_n822_), .Y(_abc_4635_new_n827_));
OAI21X1 OAI21X1_104 ( .A(\W_R[1] ), .B(_abc_4635_new_n831_), .C(_abc_4635_new_n832_), .Y(\ARdata[7] ));
OAI21X1 OAI21X1_105 ( .A(_abc_4635_new_n815_), .B(_abc_4635_new_n835_), .C(_abc_4635_new_n837_), .Y(_abc_4635_new_n838_));
OAI21X1 OAI21X1_106 ( .A(\W_R[1] ), .B(_abc_4635_new_n843_), .C(_abc_4635_new_n834_), .Y(\ARdata[8] ));
OAI21X1 OAI21X1_107 ( .A(_abc_4635_new_n841_), .B(_abc_4635_new_n839_), .C(_abc_4635_new_n845_), .Y(_abc_4635_new_n846_));
OAI21X1 OAI21X1_108 ( .A(\W_R[1] ), .B(_abc_4635_new_n850_), .C(_abc_4635_new_n851_), .Y(\ARdata[9] ));
OAI21X1 OAI21X1_109 ( .A(_abc_4635_new_n856_), .B(_abc_4635_new_n839_), .C(_abc_4635_new_n855_), .Y(_abc_4635_new_n857_));
OAI21X1 OAI21X1_11 ( .A(state_4_), .B(_abc_4635_new_n412_), .C(resetn), .Y(_abc_4635_new_n413_));
OAI21X1 OAI21X1_110 ( .A(_abc_4635_new_n861_), .B(_abc_4635_new_n863_), .C(_abc_4635_new_n853_), .Y(\ARdata[10] ));
OAI21X1 OAI21X1_111 ( .A(\W_R[1] ), .B(_abc_4635_new_n869_), .C(_abc_4635_new_n870_), .Y(\ARdata[11] ));
OAI21X1 OAI21X1_112 ( .A(_abc_4635_new_n855_), .B(_abc_4635_new_n873_), .C(_abc_4635_new_n874_), .Y(_abc_4635_new_n875_));
OAI21X1 OAI21X1_113 ( .A(_abc_4635_new_n838_), .B(_abc_4635_new_n887_), .C(_abc_4635_new_n888_), .Y(_abc_4635_new_n889_));
OAI21X1 OAI21X1_114 ( .A(_abc_4635_new_n892_), .B(_abc_4635_new_n894_), .C(_abc_4635_new_n872_), .Y(\ARdata[12] ));
OAI21X1 OAI21X1_115 ( .A(\W_R[1] ), .B(_abc_4635_new_n901_), .C(_abc_4635_new_n902_), .Y(\ARdata[13] ));
OAI21X1 OAI21X1_116 ( .A(_abc_4635_new_n896_), .B(_abc_4635_new_n898_), .C(_abc_4635_new_n906_), .Y(_abc_4635_new_n907_));
OAI21X1 OAI21X1_117 ( .A(_abc_4635_new_n909_), .B(_abc_4635_new_n905_), .C(_abc_4635_new_n908_), .Y(_abc_4635_new_n910_));
OAI21X1 OAI21X1_118 ( .A(\W_R[1] ), .B(_abc_4635_new_n914_), .C(_abc_4635_new_n904_), .Y(\ARdata[14] ));
OAI21X1 OAI21X1_119 ( .A(\W_R[1] ), .B(_abc_4635_new_n920_), .C(_abc_4635_new_n921_), .Y(\ARdata[15] ));
OAI21X1 OAI21X1_12 ( .A(_abc_4635_new_n386_), .B(_abc_4635_new_n418_), .C(state_0_), .Y(_abc_4635_new_n419_));
OAI21X1 OAI21X1_120 ( .A(_abc_4635_new_n924_), .B(_abc_4635_new_n908_), .C(_abc_4635_new_n927_), .Y(_abc_4635_new_n928_));
OAI21X1 OAI21X1_121 ( .A(_abc_4635_new_n926_), .B(_abc_4635_new_n839_), .C(_abc_4635_new_n929_), .Y(_abc_4635_new_n930_));
OAI21X1 OAI21X1_122 ( .A(\W_R[1] ), .B(_abc_4635_new_n935_), .C(_abc_4635_new_n923_), .Y(\ARdata[16] ));
OAI21X1 OAI21X1_123 ( .A(_abc_4635_new_n931_), .B(_abc_4635_new_n937_), .C(_abc_4635_new_n932_), .Y(_abc_4635_new_n938_));
OAI21X1 OAI21X1_124 ( .A(\W_R[1] ), .B(_abc_4635_new_n940_), .C(_abc_4635_new_n941_), .Y(\ARdata[17] ));
OAI21X1 OAI21X1_125 ( .A(_abc_4635_new_n944_), .B(_abc_4635_new_n945_), .C(_abc_4635_new_n932_), .Y(_abc_4635_new_n946_));
OAI21X1 OAI21X1_126 ( .A(\rs1[17] ), .B(\imm[17] ), .C(_abc_4635_new_n946_), .Y(_abc_4635_new_n947_));
OAI21X1 OAI21X1_127 ( .A(_abc_4635_new_n955_), .B(_abc_4635_new_n950_), .C(_abc_4635_new_n639_), .Y(_abc_4635_new_n957_));
OAI21X1 OAI21X1_128 ( .A(_abc_4635_new_n956_), .B(_abc_4635_new_n957_), .C(_abc_4635_new_n943_), .Y(\ARdata[18] ));
OAI21X1 OAI21X1_129 ( .A(_abc_4635_new_n953_), .B(_abc_4635_new_n950_), .C(_abc_4635_new_n951_), .Y(_abc_4635_new_n959_));
OAI21X1 OAI21X1_13 ( .A(Bvalid), .B(_abc_4635_new_n421_), .C(_abc_4635_new_n416_), .Y(_abc_4635_new_n422_));
OAI21X1 OAI21X1_130 ( .A(\W_R[1] ), .B(_abc_4635_new_n963_), .C(_abc_4635_new_n964_), .Y(\ARdata[19] ));
OAI21X1 OAI21X1_131 ( .A(_abc_4635_new_n947_), .B(_abc_4635_new_n967_), .C(_abc_4635_new_n968_), .Y(_abc_4635_new_n969_));
OAI21X1 OAI21X1_132 ( .A(_abc_4635_new_n976_), .B(_abc_4635_new_n973_), .C(_abc_4635_new_n639_), .Y(_abc_4635_new_n978_));
OAI21X1 OAI21X1_133 ( .A(_abc_4635_new_n977_), .B(_abc_4635_new_n978_), .C(_abc_4635_new_n966_), .Y(\ARdata[20] ));
OAI21X1 OAI21X1_134 ( .A(_abc_4635_new_n976_), .B(_abc_4635_new_n973_), .C(_abc_4635_new_n974_), .Y(_abc_4635_new_n980_));
OAI21X1 OAI21X1_135 ( .A(\W_R[1] ), .B(_abc_4635_new_n984_), .C(_abc_4635_new_n985_), .Y(\ARdata[21] ));
OAI21X1 OAI21X1_136 ( .A(_abc_4635_new_n974_), .B(_abc_4635_new_n983_), .C(_abc_4635_new_n981_), .Y(_abc_4635_new_n988_));
OAI21X1 OAI21X1_137 ( .A(_abc_4635_new_n991_), .B(_abc_4635_new_n973_), .C(_abc_4635_new_n989_), .Y(_abc_4635_new_n992_));
OAI21X1 OAI21X1_138 ( .A(_abc_4635_new_n999_), .B(_abc_4635_new_n1001_), .C(_abc_4635_new_n987_), .Y(\ARdata[22] ));
OAI21X1 OAI21X1_139 ( .A(_abc_4635_new_n994_), .B(_abc_4635_new_n995_), .C(_abc_4635_new_n1000_), .Y(_abc_4635_new_n1004_));
OAI21X1 OAI21X1_14 ( .A(_abc_4635_new_n379_), .B(_abc_4635_new_n361_), .C(state_3_), .Y(_abc_4635_new_n425_));
OAI21X1 OAI21X1_140 ( .A(_abc_4635_new_n1009_), .B(_abc_4635_new_n1008_), .C(_abc_4635_new_n639_), .Y(_abc_4635_new_n1010_));
OAI21X1 OAI21X1_141 ( .A(_abc_4635_new_n639_), .B(_abc_4635_new_n1003_), .C(_abc_4635_new_n1010_), .Y(\ARdata[23] ));
OAI21X1 OAI21X1_142 ( .A(_abc_4635_new_n1025_), .B(_abc_4635_new_n1026_), .C(_abc_4635_new_n1022_), .Y(_abc_4635_new_n1027_));
OAI21X1 OAI21X1_143 ( .A(_abc_4635_new_n838_), .B(_abc_4635_new_n887_), .C(_abc_4635_new_n1028_), .Y(_abc_4635_new_n1029_));
OAI21X1 OAI21X1_144 ( .A(_abc_4635_new_n1021_), .B(_abc_4635_new_n1031_), .C(_abc_4635_new_n1032_), .Y(_abc_4635_new_n1033_));
OAI21X1 OAI21X1_145 ( .A(\W_R[1] ), .B(_abc_4635_new_n1034_), .C(_abc_4635_new_n1012_), .Y(\ARdata[24] ));
OAI21X1 OAI21X1_146 ( .A(_abc_4635_new_n1023_), .B(_abc_4635_new_n1024_), .C(_abc_4635_new_n1033_), .Y(_abc_4635_new_n1036_));
OAI21X1 OAI21X1_147 ( .A(\W_R[1] ), .B(_abc_4635_new_n1040_), .C(_abc_4635_new_n1041_), .Y(\ARdata[25] ));
OAI21X1 OAI21X1_148 ( .A(_abc_4635_new_n1045_), .B(_abc_4635_new_n1022_), .C(_abc_4635_new_n1044_), .Y(_abc_4635_new_n1046_));
OAI21X1 OAI21X1_149 ( .A(_abc_4635_new_n1052_), .B(_abc_4635_new_n1054_), .C(_abc_4635_new_n1043_), .Y(\ARdata[26] ));
OAI21X1 OAI21X1_15 ( .A(_abc_4635_new_n392_), .B(_abc_4635_new_n395_), .C(_abc_4635_new_n425_), .Y(_abc_4635_new_n426_));
OAI21X1 OAI21X1_150 ( .A(_abc_4635_new_n1047_), .B(_abc_4635_new_n1048_), .C(_abc_4635_new_n1053_), .Y(_abc_4635_new_n1056_));
OAI21X1 OAI21X1_151 ( .A(\W_R[1] ), .B(_abc_4635_new_n1061_), .C(_abc_4635_new_n1062_), .Y(\ARdata[27] ));
OAI21X1 OAI21X1_152 ( .A(_abc_4635_new_n1057_), .B(_abc_4635_new_n1069_), .C(_abc_4635_new_n1058_), .Y(_abc_4635_new_n1070_));
OAI21X1 OAI21X1_153 ( .A(_abc_4635_new_n1067_), .B(_abc_4635_new_n1022_), .C(_abc_4635_new_n1071_), .Y(_abc_4635_new_n1072_));
OAI21X1 OAI21X1_154 ( .A(_abc_4635_new_n1078_), .B(_abc_4635_new_n1080_), .C(_abc_4635_new_n1064_), .Y(\ARdata[28] ));
OAI21X1 OAI21X1_155 ( .A(_abc_4635_new_n1074_), .B(_abc_4635_new_n1075_), .C(_abc_4635_new_n1079_), .Y(_abc_4635_new_n1082_));
OAI21X1 OAI21X1_156 ( .A(\W_R[1] ), .B(_abc_4635_new_n1087_), .C(_abc_4635_new_n1088_), .Y(\ARdata[29] ));
OAI21X1 OAI21X1_157 ( .A(_abc_4635_new_n1083_), .B(_abc_4635_new_n1093_), .C(_abc_4635_new_n1084_), .Y(_abc_4635_new_n1094_));
OAI21X1 OAI21X1_158 ( .A(_abc_4635_new_n1021_), .B(_abc_4635_new_n1031_), .C(_abc_4635_new_n1066_), .Y(_abc_4635_new_n1101_));
OAI21X1 OAI21X1_159 ( .A(_abc_4635_new_n1094_), .B(_abc_4635_new_n1102_), .C(_abc_4635_new_n1098_), .Y(_abc_4635_new_n1103_));
OAI21X1 OAI21X1_16 ( .A(_abc_4635_new_n420_), .B(_abc_4635_new_n429_), .C(resetn), .Y(done));
OAI21X1 OAI21X1_160 ( .A(\W_R[1] ), .B(_abc_4635_new_n1104_), .C(_abc_4635_new_n1090_), .Y(\ARdata[30] ));
OAI21X1 OAI21X1_161 ( .A(_abc_4635_new_n1099_), .B(_abc_4635_new_n1095_), .C(_abc_4635_new_n1097_), .Y(_abc_4635_new_n1109_));
OAI21X1 OAI21X1_162 ( .A(state_2_), .B(_abc_4635_new_n389_), .C(resetn), .Y(_abc_4635_new_n1119_));
OAI21X1 OAI21X1_163 ( .A(_abc_4635_new_n366_), .B(_abc_4635_new_n401_), .C(_abc_4635_new_n1119_), .Y(RReady));
OAI21X1 OAI21X1_164 ( .A(_abc_4635_new_n392_), .B(_abc_4635_new_n366_), .C(_abc_4635_new_n413_), .Y(AWvalid));
OAI21X1 OAI21X1_17 ( .A(_abc_4635_new_n435_), .B(_abc_4635_new_n437_), .C(_abc_4635_new_n433_), .Y(_abc_4635_new_n440_));
OAI21X1 OAI21X1_18 ( .A(_abc_4635_new_n434_), .B(_abc_4635_new_n442_), .C(_abc_4635_new_n441_), .Y(_abc_4635_new_n443_));
OAI21X1 OAI21X1_19 ( .A(_abc_4635_new_n444_), .B(_abc_4635_new_n448_), .C(_abc_4635_new_n449_), .Y(_abc_4635_new_n450_));
OAI21X1 OAI21X1_2 ( .A(_abc_4635_new_n371_), .B(_abc_4635_new_n372_), .C(resetn), .Y(_abc_4635_new_n373_));
OAI21X1 OAI21X1_20 ( .A(\wordsize[0] ), .B(_abc_4635_new_n453_), .C(_abc_4635_new_n441_), .Y(_abc_4635_new_n454_));
OAI21X1 OAI21X1_21 ( .A(\wordsize[0] ), .B(_abc_4635_new_n457_), .C(_abc_4635_new_n456_), .Y(_abc_4635_new_n458_));
OAI21X1 OAI21X1_22 ( .A(\wordsize[0] ), .B(_abc_4635_new_n453_), .C(_abc_4635_new_n456_), .Y(_abc_4635_new_n460_));
OAI21X1 OAI21X1_23 ( .A(\Rdata_mem[0] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n539_));
OAI21X1 OAI21X1_24 ( .A(\Rdata_mem[1] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n542_));
OAI21X1 OAI21X1_25 ( .A(\Rdata_mem[2] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n545_));
OAI21X1 OAI21X1_26 ( .A(\Rdata_mem[3] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n548_));
OAI21X1 OAI21X1_27 ( .A(\Rdata_mem[4] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n551_));
OAI21X1 OAI21X1_28 ( .A(\Rdata_mem[5] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n554_));
OAI21X1 OAI21X1_29 ( .A(\Rdata_mem[6] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n557_));
OAI21X1 OAI21X1_3 ( .A(_abc_4635_new_n382_), .B(_abc_4635_new_n383_), .C(state_2_), .Y(_abc_4635_new_n384_));
OAI21X1 OAI21X1_30 ( .A(\Rdata_mem[7] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n560_));
OAI21X1 OAI21X1_31 ( .A(\Rdata_mem[8] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n563_));
OAI21X1 OAI21X1_32 ( .A(\Rdata_mem[9] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n566_));
OAI21X1 OAI21X1_33 ( .A(\Rdata_mem[10] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n569_));
OAI21X1 OAI21X1_34 ( .A(\Rdata_mem[11] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n572_));
OAI21X1 OAI21X1_35 ( .A(\Rdata_mem[12] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n575_));
OAI21X1 OAI21X1_36 ( .A(\Rdata_mem[13] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n578_));
OAI21X1 OAI21X1_37 ( .A(\Rdata_mem[14] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n581_));
OAI21X1 OAI21X1_38 ( .A(\Rdata_mem[15] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n584_));
OAI21X1 OAI21X1_39 ( .A(\Rdata_mem[16] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n587_));
OAI21X1 OAI21X1_4 ( .A(\W_R[0] ), .B(\W_R[1] ), .C(enable), .Y(_abc_4635_new_n386_));
OAI21X1 OAI21X1_40 ( .A(\Rdata_mem[17] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n590_));
OAI21X1 OAI21X1_41 ( .A(\Rdata_mem[18] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n593_));
OAI21X1 OAI21X1_42 ( .A(\Rdata_mem[19] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n596_));
OAI21X1 OAI21X1_43 ( .A(\Rdata_mem[20] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n599_));
OAI21X1 OAI21X1_44 ( .A(\Rdata_mem[21] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n602_));
OAI21X1 OAI21X1_45 ( .A(\Rdata_mem[22] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n605_));
OAI21X1 OAI21X1_46 ( .A(\Rdata_mem[23] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n608_));
OAI21X1 OAI21X1_47 ( .A(\Rdata_mem[24] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n611_));
OAI21X1 OAI21X1_48 ( .A(\Rdata_mem[25] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n614_));
OAI21X1 OAI21X1_49 ( .A(\Rdata_mem[26] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n617_));
OAI21X1 OAI21X1_5 ( .A(_abc_4635_new_n385_), .B(_abc_4635_new_n389_), .C(resetn), .Y(_abc_4635_new_n390_));
OAI21X1 OAI21X1_50 ( .A(\Rdata_mem[27] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n620_));
OAI21X1 OAI21X1_51 ( .A(\Rdata_mem[28] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n623_));
OAI21X1 OAI21X1_52 ( .A(\Rdata_mem[29] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n626_));
OAI21X1 OAI21X1_53 ( .A(\Rdata_mem[30] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n629_));
OAI21X1 OAI21X1_54 ( .A(\Rdata_mem[31] ), .B(_abc_4635_new_n538_), .C(resetn), .Y(_abc_4635_new_n632_));
OAI21X1 OAI21X1_55 ( .A(_abc_4635_new_n445_), .B(_abc_4635_new_n479_), .C(_abc_4635_new_n635_), .Y(_abc_4635_new_n636_));
OAI21X1 OAI21X1_56 ( .A(_abc_4635_new_n634_), .B(_abc_4635_new_n443_), .C(_abc_4635_new_n637_), .Y(align));
OAI21X1 OAI21X1_57 ( .A(\Rdata_mem[16] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n457_), .Y(_abc_4635_new_n643_));
OAI21X1 OAI21X1_58 ( .A(_abc_4635_new_n457_), .B(_abc_4635_new_n644_), .C(_abc_4635_new_n643_), .Y(_abc_4635_new_n645_));
OAI21X1 OAI21X1_59 ( .A(\Rdata_mem[0] ), .B(_abc_4635_new_n443_), .C(_abc_4635_new_n645_), .Y(_abc_4635_new_n646_));
OAI21X1 OAI21X1_6 ( .A(_abc_4635_new_n374_), .B(_abc_4635_new_n396_), .C(enable), .Y(_abc_4635_new_n397_));
OAI21X1 OAI21X1_60 ( .A(_abc_4635_new_n446_), .B(_abc_4635_new_n456_), .C(_abc_4635_new_n634_), .Y(_abc_4635_new_n647_));
OAI21X1 OAI21X1_61 ( .A(_abc_4635_new_n642_), .B(_abc_4635_new_n646_), .C(_abc_4635_new_n648_), .Y(_abc_4635_new_n649_));
OAI21X1 OAI21X1_62 ( .A(\Rdata_mem[17] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n457_), .Y(_abc_4635_new_n652_));
OAI21X1 OAI21X1_63 ( .A(_abc_4635_new_n457_), .B(_abc_4635_new_n651_), .C(_abc_4635_new_n652_), .Y(_abc_4635_new_n653_));
OAI21X1 OAI21X1_64 ( .A(\Rdata_mem[1] ), .B(_abc_4635_new_n443_), .C(_abc_4635_new_n653_), .Y(_abc_4635_new_n654_));
OAI21X1 OAI21X1_65 ( .A(\Rdata_mem[17] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n445_), .Y(_abc_4635_new_n656_));
OAI21X1 OAI21X1_66 ( .A(_abc_4635_new_n642_), .B(_abc_4635_new_n654_), .C(_abc_4635_new_n658_), .Y(_abc_4635_new_n659_));
OAI21X1 OAI21X1_67 ( .A(\Rdata_mem[18] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n457_), .Y(_abc_4635_new_n662_));
OAI21X1 OAI21X1_68 ( .A(_abc_4635_new_n457_), .B(_abc_4635_new_n661_), .C(_abc_4635_new_n662_), .Y(_abc_4635_new_n663_));
OAI21X1 OAI21X1_69 ( .A(\Rdata_mem[2] ), .B(_abc_4635_new_n443_), .C(_abc_4635_new_n663_), .Y(_abc_4635_new_n664_));
OAI21X1 OAI21X1_7 ( .A(_abc_4635_new_n400_), .B(_abc_4635_new_n382_), .C(_abc_4635_new_n401_), .Y(_abc_4635_new_n402_));
OAI21X1 OAI21X1_70 ( .A(\Rdata_mem[18] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n445_), .Y(_abc_4635_new_n666_));
OAI21X1 OAI21X1_71 ( .A(_abc_4635_new_n642_), .B(_abc_4635_new_n664_), .C(_abc_4635_new_n668_), .Y(_abc_4635_new_n669_));
OAI21X1 OAI21X1_72 ( .A(\Rdata_mem[19] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n457_), .Y(_abc_4635_new_n672_));
OAI21X1 OAI21X1_73 ( .A(_abc_4635_new_n457_), .B(_abc_4635_new_n671_), .C(_abc_4635_new_n672_), .Y(_abc_4635_new_n673_));
OAI21X1 OAI21X1_74 ( .A(\Rdata_mem[3] ), .B(_abc_4635_new_n443_), .C(_abc_4635_new_n673_), .Y(_abc_4635_new_n674_));
OAI21X1 OAI21X1_75 ( .A(\Rdata_mem[19] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n445_), .Y(_abc_4635_new_n676_));
OAI21X1 OAI21X1_76 ( .A(_abc_4635_new_n642_), .B(_abc_4635_new_n674_), .C(_abc_4635_new_n678_), .Y(_abc_4635_new_n679_));
OAI21X1 OAI21X1_77 ( .A(\Rdata_mem[20] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n457_), .Y(_abc_4635_new_n681_));
OAI21X1 OAI21X1_78 ( .A(_abc_4635_new_n457_), .B(_abc_4635_new_n682_), .C(_abc_4635_new_n681_), .Y(_abc_4635_new_n683_));
OAI21X1 OAI21X1_79 ( .A(\Rdata_mem[4] ), .B(_abc_4635_new_n443_), .C(_abc_4635_new_n683_), .Y(_abc_4635_new_n684_));
OAI21X1 OAI21X1_8 ( .A(_abc_4635_new_n404_), .B(_abc_4635_new_n396_), .C(resetn), .Y(_abc_4635_new_n405_));
OAI21X1 OAI21X1_80 ( .A(_abc_4635_new_n642_), .B(_abc_4635_new_n684_), .C(_abc_4635_new_n685_), .Y(_abc_4635_new_n686_));
OAI21X1 OAI21X1_81 ( .A(\Rdata_mem[21] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n457_), .Y(_abc_4635_new_n688_));
OAI21X1 OAI21X1_82 ( .A(_abc_4635_new_n457_), .B(_abc_4635_new_n689_), .C(_abc_4635_new_n688_), .Y(_abc_4635_new_n690_));
OAI21X1 OAI21X1_83 ( .A(\Rdata_mem[5] ), .B(_abc_4635_new_n443_), .C(_abc_4635_new_n690_), .Y(_abc_4635_new_n691_));
OAI21X1 OAI21X1_84 ( .A(_abc_4635_new_n642_), .B(_abc_4635_new_n691_), .C(_abc_4635_new_n692_), .Y(_abc_4635_new_n693_));
OAI21X1 OAI21X1_85 ( .A(\Rdata_mem[22] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n457_), .Y(_abc_4635_new_n696_));
OAI21X1 OAI21X1_86 ( .A(_abc_4635_new_n457_), .B(_abc_4635_new_n695_), .C(_abc_4635_new_n696_), .Y(_abc_4635_new_n697_));
OAI21X1 OAI21X1_87 ( .A(\Rdata_mem[6] ), .B(_abc_4635_new_n443_), .C(_abc_4635_new_n697_), .Y(_abc_4635_new_n698_));
OAI21X1 OAI21X1_88 ( .A(\Rdata_mem[22] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n445_), .Y(_abc_4635_new_n700_));
OAI21X1 OAI21X1_89 ( .A(_abc_4635_new_n642_), .B(_abc_4635_new_n698_), .C(_abc_4635_new_n702_), .Y(_abc_4635_new_n703_));
OAI21X1 OAI21X1_9 ( .A(_abc_4635_new_n367_), .B(_abc_4635_new_n404_), .C(_abc_4635_new_n362_), .Y(_abc_4635_new_n409_));
OAI21X1 OAI21X1_90 ( .A(\Rdata_mem[7] ), .B(_abc_4635_new_n456_), .C(_abc_4635_new_n706_), .Y(_abc_4635_new_n707_));
OAI21X1 OAI21X1_91 ( .A(_abc_4635_new_n713_), .B(_abc_4635_new_n709_), .C(_abc_4635_new_n717_), .Y(_abc_4635_new_n718_));
OAI21X1 OAI21X1_92 ( .A(_abc_4635_new_n705_), .B(_abc_4635_new_n634_), .C(_abc_4635_new_n744_), .Y(_abc_4635_new_n758_));
OAI21X1 OAI21X1_93 ( .A(\W_R[1] ), .B(_abc_4635_new_n457_), .C(_abc_4635_new_n776_), .Y(\ARdata[0] ));
OAI21X1 OAI21X1_94 ( .A(\W_R[1] ), .B(_abc_4635_new_n441_), .C(_abc_4635_new_n778_), .Y(\ARdata[1] ));
OAI21X1 OAI21X1_95 ( .A(_abc_4635_new_n433_), .B(_abc_4635_new_n435_), .C(_abc_4635_new_n436_), .Y(_abc_4635_new_n780_));
OAI21X1 OAI21X1_96 ( .A(\W_R[1] ), .B(_abc_4635_new_n784_), .C(_abc_4635_new_n785_), .Y(\ARdata[2] ));
OAI21X1 OAI21X1_97 ( .A(\W_R[1] ), .B(_abc_4635_new_n791_), .C(_abc_4635_new_n792_), .Y(\ARdata[3] ));
OAI21X1 OAI21X1_98 ( .A(\W_R[1] ), .B(_abc_4635_new_n801_), .C(_abc_4635_new_n802_), .Y(\ARdata[4] ));
OAI21X1 OAI21X1_99 ( .A(_abc_4635_new_n798_), .B(_abc_4635_new_n804_), .C(_abc_4635_new_n805_), .Y(_abc_4635_new_n806_));
OAI22X1 OAI22X1_1 ( .A(Bvalid), .B(_abc_4635_new_n365_), .C(_abc_4635_new_n380_), .D(_abc_4635_new_n378_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_1_));
OAI22X1 OAI22X1_2 ( .A(_abc_4635_new_n392_), .B(_abc_4635_new_n366_), .C(_abc_4635_new_n361_), .D(_abc_4635_new_n378_), .Y(_abc_4635_new_n393_));
OAI22X1 OAI22X1_3 ( .A(_abc_4635_new_n366_), .B(_abc_4635_new_n416_), .C(_abc_4635_new_n415_), .D(_abc_4635_new_n390_), .Y(_abc_3813_auto_fsm_map_cc_170_map_fsm_1372_5_));
OAI22X1 OAI22X1_4 ( .A(_abc_4635_new_n457_), .B(_abc_4635_new_n712_), .C(_abc_4635_new_n711_), .D(_abc_4635_new_n710_), .Y(_abc_4635_new_n713_));
OR2X2 OR2X2_1 ( .A(_abc_4635_new_n424_), .B(_abc_4635_new_n426_), .Y(_abc_4635_new_n427_));
OR2X2 OR2X2_10 ( .A(\rs1[30] ), .B(\imm[30] ), .Y(_abc_4635_new_n1096_));
OR2X2 OR2X2_2 ( .A(_abc_4635_new_n447_), .B(_abc_4635_new_n450_), .Y(_abc_4635_new_n451_));
OR2X2 OR2X2_3 ( .A(_abc_4635_new_n709_), .B(_abc_4635_new_n713_), .Y(_abc_4635_new_n714_));
OR2X2 OR2X2_4 ( .A(\rs1[5] ), .B(\imm[5] ), .Y(_abc_4635_new_n814_));
OR2X2 OR2X2_5 ( .A(\rs1[9] ), .B(\imm[9] ), .Y(_abc_4635_new_n854_));
OR2X2 OR2X2_6 ( .A(\rs1[4] ), .B(\imm[4] ), .Y(_abc_4635_new_n877_));
OR2X2 OR2X2_7 ( .A(\rs1[20] ), .B(\imm[20] ), .Y(_abc_4635_new_n975_));
OR2X2 OR2X2_8 ( .A(\rs1[21] ), .B(\imm[21] ), .Y(_abc_4635_new_n982_));
OR2X2 OR2X2_9 ( .A(_abc_4635_new_n1005_), .B(_abc_4635_new_n1006_), .Y(_abc_4635_new_n1007_));
XNOR2X1 XNOR2X1_1 ( .A(_abc_4635_new_n780_), .B(_abc_4635_new_n783_), .Y(_abc_4635_new_n784_));
XNOR2X1 XNOR2X1_10 ( .A(_abc_4635_new_n938_), .B(_abc_4635_new_n939_), .Y(_abc_4635_new_n940_));
XNOR2X1 XNOR2X1_11 ( .A(_abc_4635_new_n959_), .B(_abc_4635_new_n962_), .Y(_abc_4635_new_n963_));
XNOR2X1 XNOR2X1_12 ( .A(_abc_4635_new_n1036_), .B(_abc_4635_new_n1039_), .Y(_abc_4635_new_n1040_));
XNOR2X1 XNOR2X1_13 ( .A(_abc_4635_new_n1056_), .B(_abc_4635_new_n1060_), .Y(_abc_4635_new_n1061_));
XNOR2X1 XNOR2X1_14 ( .A(_abc_4635_new_n1082_), .B(_abc_4635_new_n1086_), .Y(_abc_4635_new_n1087_));
XNOR2X1 XNOR2X1_15 ( .A(\rs1[31] ), .B(\imm[31] ), .Y(_abc_4635_new_n1107_));
XNOR2X1 XNOR2X1_2 ( .A(_abc_4635_new_n797_), .B(_abc_4635_new_n800_), .Y(_abc_4635_new_n801_));
XNOR2X1 XNOR2X1_3 ( .A(_abc_4635_new_n806_), .B(_abc_4635_new_n809_), .Y(_abc_4635_new_n810_));
XNOR2X1 XNOR2X1_4 ( .A(_abc_4635_new_n827_), .B(_abc_4635_new_n830_), .Y(_abc_4635_new_n831_));
XNOR2X1 XNOR2X1_5 ( .A(_abc_4635_new_n846_), .B(_abc_4635_new_n849_), .Y(_abc_4635_new_n850_));
XNOR2X1 XNOR2X1_6 ( .A(\rs1[7] ), .B(\imm[7] ), .Y(_abc_4635_new_n884_));
XNOR2X1 XNOR2X1_7 ( .A(_abc_4635_new_n897_), .B(_abc_4635_new_n900_), .Y(_abc_4635_new_n901_));
XNOR2X1 XNOR2X1_8 ( .A(_abc_4635_new_n910_), .B(_abc_4635_new_n913_), .Y(_abc_4635_new_n914_));
XNOR2X1 XNOR2X1_9 ( .A(_abc_4635_new_n930_), .B(_abc_4635_new_n934_), .Y(_abc_4635_new_n935_));
XOR2X1 XOR2X1_1 ( .A(_abc_4635_new_n787_), .B(_abc_4635_new_n790_), .Y(_abc_4635_new_n791_));
XOR2X1 XOR2X1_2 ( .A(_abc_4635_new_n839_), .B(_abc_4635_new_n842_), .Y(_abc_4635_new_n843_));
XOR2X1 XOR2X1_3 ( .A(_abc_4635_new_n865_), .B(_abc_4635_new_n868_), .Y(_abc_4635_new_n869_));
XOR2X1 XOR2X1_4 ( .A(\rs1[12] ), .B(\imm[12] ), .Y(_abc_4635_new_n891_));
XOR2X1 XOR2X1_5 ( .A(_abc_4635_new_n916_), .B(_abc_4635_new_n919_), .Y(_abc_4635_new_n920_));
XOR2X1 XOR2X1_6 ( .A(\rs1[17] ), .B(\imm[17] ), .Y(_abc_4635_new_n939_));
XOR2X1 XOR2X1_7 ( .A(_abc_4635_new_n980_), .B(_abc_4635_new_n983_), .Y(_abc_4635_new_n984_));

assign \arprot[0]  = 1'h0;
assign \arprot[1]  = 1'h0;
assign \awprot[0]  = 1'h0;
assign \awprot[1]  = 1'h0;
assign \awprot[2]  = 1'h0;

endmodule