module b14_reset(clock, RESET_G, nRESET_G, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, ADDR_REG_19_, ADDR_REG_18_, ADDR_REG_17_, ADDR_REG_16_, ADDR_REG_15_, ADDR_REG_14_, ADDR_REG_13_, ADDR_REG_12_, ADDR_REG_11_, ADDR_REG_10_, ADDR_REG_9_, ADDR_REG_8_, ADDR_REG_7_, ADDR_REG_6_, ADDR_REG_5_, ADDR_REG_4_, ADDR_REG_3_, ADDR_REG_2_, ADDR_REG_1_, ADDR_REG_0_, DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_, DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_, DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_, DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_, DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_, DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_, DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_, DATAO_REG_1_, DATAO_REG_0_, RD_REG, WR_REG);

output ADDR_REG_0_;
output ADDR_REG_10_;
output ADDR_REG_11_;
output ADDR_REG_12_;
output ADDR_REG_13_;
output ADDR_REG_14_;
output ADDR_REG_15_;
output ADDR_REG_16_;
output ADDR_REG_17_;
output ADDR_REG_18_;
output ADDR_REG_19_;
output ADDR_REG_1_;
output ADDR_REG_2_;
output ADDR_REG_3_;
output ADDR_REG_4_;
output ADDR_REG_5_;
output ADDR_REG_6_;
output ADDR_REG_7_;
output ADDR_REG_8_;
output ADDR_REG_9_;
wire B_REG; 
input DATAI_0_;
input DATAI_10_;
input DATAI_11_;
input DATAI_12_;
input DATAI_13_;
input DATAI_14_;
input DATAI_15_;
input DATAI_16_;
input DATAI_17_;
input DATAI_18_;
input DATAI_19_;
input DATAI_1_;
input DATAI_20_;
input DATAI_21_;
input DATAI_22_;
input DATAI_23_;
input DATAI_24_;
input DATAI_25_;
input DATAI_26_;
input DATAI_27_;
input DATAI_28_;
input DATAI_29_;
input DATAI_2_;
input DATAI_30_;
input DATAI_31_;
input DATAI_3_;
input DATAI_4_;
input DATAI_5_;
input DATAI_6_;
input DATAI_7_;
input DATAI_8_;
input DATAI_9_;
output DATAO_REG_0_;
output DATAO_REG_10_;
output DATAO_REG_11_;
output DATAO_REG_12_;
output DATAO_REG_13_;
output DATAO_REG_14_;
output DATAO_REG_15_;
output DATAO_REG_16_;
output DATAO_REG_17_;
output DATAO_REG_18_;
output DATAO_REG_19_;
output DATAO_REG_1_;
output DATAO_REG_20_;
output DATAO_REG_21_;
output DATAO_REG_22_;
output DATAO_REG_23_;
output DATAO_REG_24_;
output DATAO_REG_25_;
output DATAO_REG_26_;
output DATAO_REG_27_;
output DATAO_REG_28_;
output DATAO_REG_29_;
output DATAO_REG_2_;
output DATAO_REG_30_;
output DATAO_REG_31_;
output DATAO_REG_3_;
output DATAO_REG_4_;
output DATAO_REG_5_;
output DATAO_REG_6_;
output DATAO_REG_7_;
output DATAO_REG_8_;
output DATAO_REG_9_;
wire D_REG_0_; 
wire D_REG_10_; 
wire D_REG_11_; 
wire D_REG_12_; 
wire D_REG_13_; 
wire D_REG_14_; 
wire D_REG_15_; 
wire D_REG_16_; 
wire D_REG_17_; 
wire D_REG_18_; 
wire D_REG_19_; 
wire D_REG_1_; 
wire D_REG_20_; 
wire D_REG_21_; 
wire D_REG_22_; 
wire D_REG_23_; 
wire D_REG_24_; 
wire D_REG_25_; 
wire D_REG_26_; 
wire D_REG_27_; 
wire D_REG_28_; 
wire D_REG_29_; 
wire D_REG_2_; 
wire D_REG_30_; 
wire D_REG_31_; 
wire D_REG_3_; 
wire D_REG_4_; 
wire D_REG_5_; 
wire D_REG_6_; 
wire D_REG_7_; 
wire D_REG_8_; 
wire D_REG_9_; 
wire IR_REG_0_; 
wire IR_REG_10_; 
wire IR_REG_11_; 
wire IR_REG_12_; 
wire IR_REG_13_; 
wire IR_REG_14_; 
wire IR_REG_15_; 
wire IR_REG_16_; 
wire IR_REG_17_; 
wire IR_REG_18_; 
wire IR_REG_19_; 
wire IR_REG_1_; 
wire IR_REG_20_; 
wire IR_REG_21_; 
wire IR_REG_22_; 
wire IR_REG_23_; 
wire IR_REG_24_; 
wire IR_REG_25_; 
wire IR_REG_26_; 
wire IR_REG_27_; 
wire IR_REG_28_; 
wire IR_REG_29_; 
wire IR_REG_2_; 
wire IR_REG_30_; 
wire IR_REG_31_; 
wire IR_REG_3_; 
wire IR_REG_4_; 
wire IR_REG_5_; 
wire IR_REG_6_; 
wire IR_REG_7_; 
wire IR_REG_8_; 
wire IR_REG_9_; 
output RD_REG;
wire REG0_REG_0_; 
wire REG0_REG_10_; 
wire REG0_REG_11_; 
wire REG0_REG_12_; 
wire REG0_REG_13_; 
wire REG0_REG_14_; 
wire REG0_REG_15_; 
wire REG0_REG_16_; 
wire REG0_REG_17_; 
wire REG0_REG_18_; 
wire REG0_REG_19_; 
wire REG0_REG_1_; 
wire REG0_REG_20_; 
wire REG0_REG_21_; 
wire REG0_REG_22_; 
wire REG0_REG_23_; 
wire REG0_REG_24_; 
wire REG0_REG_25_; 
wire REG0_REG_26_; 
wire REG0_REG_27_; 
wire REG0_REG_28_; 
wire REG0_REG_29_; 
wire REG0_REG_2_; 
wire REG0_REG_30_; 
wire REG0_REG_31_; 
wire REG0_REG_3_; 
wire REG0_REG_4_; 
wire REG0_REG_5_; 
wire REG0_REG_6_; 
wire REG0_REG_7_; 
wire REG0_REG_8_; 
wire REG0_REG_9_; 
wire REG1_REG_0_; 
wire REG1_REG_10_; 
wire REG1_REG_11_; 
wire REG1_REG_12_; 
wire REG1_REG_13_; 
wire REG1_REG_14_; 
wire REG1_REG_15_; 
wire REG1_REG_16_; 
wire REG1_REG_17_; 
wire REG1_REG_18_; 
wire REG1_REG_19_; 
wire REG1_REG_1_; 
wire REG1_REG_20_; 
wire REG1_REG_21_; 
wire REG1_REG_22_; 
wire REG1_REG_23_; 
wire REG1_REG_24_; 
wire REG1_REG_25_; 
wire REG1_REG_26_; 
wire REG1_REG_27_; 
wire REG1_REG_28_; 
wire REG1_REG_29_; 
wire REG1_REG_2_; 
wire REG1_REG_30_; 
wire REG1_REG_31_; 
wire REG1_REG_3_; 
wire REG1_REG_4_; 
wire REG1_REG_5_; 
wire REG1_REG_6_; 
wire REG1_REG_7_; 
wire REG1_REG_8_; 
wire REG1_REG_9_; 
wire REG2_REG_0_; 
wire REG2_REG_10_; 
wire REG2_REG_11_; 
wire REG2_REG_12_; 
wire REG2_REG_13_; 
wire REG2_REG_14_; 
wire REG2_REG_15_; 
wire REG2_REG_16_; 
wire REG2_REG_17_; 
wire REG2_REG_18_; 
wire REG2_REG_19_; 
wire REG2_REG_1_; 
wire REG2_REG_20_; 
wire REG2_REG_21_; 
wire REG2_REG_22_; 
wire REG2_REG_23_; 
wire REG2_REG_24_; 
wire REG2_REG_25_; 
wire REG2_REG_26_; 
wire REG2_REG_27_; 
wire REG2_REG_28_; 
wire REG2_REG_29_; 
wire REG2_REG_2_; 
wire REG2_REG_30_; 
wire REG2_REG_31_; 
wire REG2_REG_3_; 
wire REG2_REG_4_; 
wire REG2_REG_5_; 
wire REG2_REG_6_; 
wire REG2_REG_7_; 
wire REG2_REG_8_; 
wire REG2_REG_9_; 
wire REG3_REG_0_; 
wire REG3_REG_10_; 
wire REG3_REG_11_; 
wire REG3_REG_12_; 
wire REG3_REG_13_; 
wire REG3_REG_14_; 
wire REG3_REG_15_; 
wire REG3_REG_16_; 
wire REG3_REG_17_; 
wire REG3_REG_18_; 
wire REG3_REG_19_; 
wire REG3_REG_1_; 
wire REG3_REG_20_; 
wire REG3_REG_21_; 
wire REG3_REG_22_; 
wire REG3_REG_23_; 
wire REG3_REG_24_; 
wire REG3_REG_25_; 
wire REG3_REG_26_; 
wire REG3_REG_27_; 
wire REG3_REG_28_; 
wire REG3_REG_2_; 
wire REG3_REG_3_; 
wire REG3_REG_4_; 
wire REG3_REG_5_; 
wire REG3_REG_6_; 
wire REG3_REG_7_; 
wire REG3_REG_8_; 
wire REG3_REG_9_; 
input RESET_G;
wire STATE_REG; 
output WR_REG;
wire _abc_40319_new_n1000_; 
wire _abc_40319_new_n1001_; 
wire _abc_40319_new_n1002_; 
wire _abc_40319_new_n1003_; 
wire _abc_40319_new_n1004_; 
wire _abc_40319_new_n1005_; 
wire _abc_40319_new_n1006_; 
wire _abc_40319_new_n1007_; 
wire _abc_40319_new_n1008_; 
wire _abc_40319_new_n1009_; 
wire _abc_40319_new_n1010_; 
wire _abc_40319_new_n1011_; 
wire _abc_40319_new_n1012_; 
wire _abc_40319_new_n1013_; 
wire _abc_40319_new_n1014_; 
wire _abc_40319_new_n1015_; 
wire _abc_40319_new_n1017_; 
wire _abc_40319_new_n1018_; 
wire _abc_40319_new_n1019_; 
wire _abc_40319_new_n1020_; 
wire _abc_40319_new_n1021_; 
wire _abc_40319_new_n1022_; 
wire _abc_40319_new_n1023_; 
wire _abc_40319_new_n1024_; 
wire _abc_40319_new_n1025_; 
wire _abc_40319_new_n1026_; 
wire _abc_40319_new_n1027_; 
wire _abc_40319_new_n1028_; 
wire _abc_40319_new_n1029_; 
wire _abc_40319_new_n1030_; 
wire _abc_40319_new_n1031_; 
wire _abc_40319_new_n1032_; 
wire _abc_40319_new_n1033_; 
wire _abc_40319_new_n1034_; 
wire _abc_40319_new_n1035_; 
wire _abc_40319_new_n1036_; 
wire _abc_40319_new_n1037_; 
wire _abc_40319_new_n1038_; 
wire _abc_40319_new_n1039_; 
wire _abc_40319_new_n1040_; 
wire _abc_40319_new_n1041_; 
wire _abc_40319_new_n1042_; 
wire _abc_40319_new_n1043_; 
wire _abc_40319_new_n1044_; 
wire _abc_40319_new_n1045_; 
wire _abc_40319_new_n1046_; 
wire _abc_40319_new_n1047_; 
wire _abc_40319_new_n1048_; 
wire _abc_40319_new_n1049_; 
wire _abc_40319_new_n1050_; 
wire _abc_40319_new_n1051_; 
wire _abc_40319_new_n1052_; 
wire _abc_40319_new_n1053_; 
wire _abc_40319_new_n1054_; 
wire _abc_40319_new_n1055_; 
wire _abc_40319_new_n1056_; 
wire _abc_40319_new_n1057_; 
wire _abc_40319_new_n1058_; 
wire _abc_40319_new_n1059_; 
wire _abc_40319_new_n1060_; 
wire _abc_40319_new_n1061_; 
wire _abc_40319_new_n1062_; 
wire _abc_40319_new_n1063_; 
wire _abc_40319_new_n1064_; 
wire _abc_40319_new_n1065_; 
wire _abc_40319_new_n1066_; 
wire _abc_40319_new_n1067_; 
wire _abc_40319_new_n1068_; 
wire _abc_40319_new_n1069_; 
wire _abc_40319_new_n1070_; 
wire _abc_40319_new_n1071_; 
wire _abc_40319_new_n1072_; 
wire _abc_40319_new_n1073_; 
wire _abc_40319_new_n1074_; 
wire _abc_40319_new_n1075_; 
wire _abc_40319_new_n1076_; 
wire _abc_40319_new_n1077_; 
wire _abc_40319_new_n1078_; 
wire _abc_40319_new_n1079_; 
wire _abc_40319_new_n1080_; 
wire _abc_40319_new_n1081_; 
wire _abc_40319_new_n1082_; 
wire _abc_40319_new_n1083_; 
wire _abc_40319_new_n1084_; 
wire _abc_40319_new_n1085_; 
wire _abc_40319_new_n1086_; 
wire _abc_40319_new_n1087_; 
wire _abc_40319_new_n1088_; 
wire _abc_40319_new_n1089_; 
wire _abc_40319_new_n1090_; 
wire _abc_40319_new_n1091_; 
wire _abc_40319_new_n1092_; 
wire _abc_40319_new_n1093_; 
wire _abc_40319_new_n1094_; 
wire _abc_40319_new_n1095_; 
wire _abc_40319_new_n1096_; 
wire _abc_40319_new_n1097_; 
wire _abc_40319_new_n1098_; 
wire _abc_40319_new_n1099_; 
wire _abc_40319_new_n1100_; 
wire _abc_40319_new_n1101_; 
wire _abc_40319_new_n1102_; 
wire _abc_40319_new_n1103_; 
wire _abc_40319_new_n1104_; 
wire _abc_40319_new_n1105_; 
wire _abc_40319_new_n1106_; 
wire _abc_40319_new_n1107_; 
wire _abc_40319_new_n1108_; 
wire _abc_40319_new_n1109_; 
wire _abc_40319_new_n1110_; 
wire _abc_40319_new_n1111_; 
wire _abc_40319_new_n1112_; 
wire _abc_40319_new_n1113_; 
wire _abc_40319_new_n1114_; 
wire _abc_40319_new_n1115_; 
wire _abc_40319_new_n1116_; 
wire _abc_40319_new_n1117_; 
wire _abc_40319_new_n1118_; 
wire _abc_40319_new_n1119_; 
wire _abc_40319_new_n1120_; 
wire _abc_40319_new_n1121_; 
wire _abc_40319_new_n1122_; 
wire _abc_40319_new_n1123_; 
wire _abc_40319_new_n1124_; 
wire _abc_40319_new_n1125_; 
wire _abc_40319_new_n1126_; 
wire _abc_40319_new_n1127_; 
wire _abc_40319_new_n1128_; 
wire _abc_40319_new_n1129_; 
wire _abc_40319_new_n1130_; 
wire _abc_40319_new_n1131_; 
wire _abc_40319_new_n1132_; 
wire _abc_40319_new_n1133_; 
wire _abc_40319_new_n1134_; 
wire _abc_40319_new_n1135_; 
wire _abc_40319_new_n1136_; 
wire _abc_40319_new_n1137_; 
wire _abc_40319_new_n1138_; 
wire _abc_40319_new_n1139_; 
wire _abc_40319_new_n1140_; 
wire _abc_40319_new_n1141_; 
wire _abc_40319_new_n1142_; 
wire _abc_40319_new_n1143_; 
wire _abc_40319_new_n1144_; 
wire _abc_40319_new_n1145_; 
wire _abc_40319_new_n1146_; 
wire _abc_40319_new_n1147_; 
wire _abc_40319_new_n1148_; 
wire _abc_40319_new_n1149_; 
wire _abc_40319_new_n1150_; 
wire _abc_40319_new_n1151_; 
wire _abc_40319_new_n1152_; 
wire _abc_40319_new_n1153_; 
wire _abc_40319_new_n1154_; 
wire _abc_40319_new_n1155_; 
wire _abc_40319_new_n1156_; 
wire _abc_40319_new_n1157_; 
wire _abc_40319_new_n1158_; 
wire _abc_40319_new_n1159_; 
wire _abc_40319_new_n1160_; 
wire _abc_40319_new_n1161_; 
wire _abc_40319_new_n1162_; 
wire _abc_40319_new_n1163_; 
wire _abc_40319_new_n1164_; 
wire _abc_40319_new_n1165_; 
wire _abc_40319_new_n1166_; 
wire _abc_40319_new_n1167_; 
wire _abc_40319_new_n1168_; 
wire _abc_40319_new_n1169_; 
wire _abc_40319_new_n1170_; 
wire _abc_40319_new_n1171_; 
wire _abc_40319_new_n1172_; 
wire _abc_40319_new_n1173_; 
wire _abc_40319_new_n1174_; 
wire _abc_40319_new_n1175_; 
wire _abc_40319_new_n1176_; 
wire _abc_40319_new_n1177_; 
wire _abc_40319_new_n1178_; 
wire _abc_40319_new_n1179_; 
wire _abc_40319_new_n1180_; 
wire _abc_40319_new_n1181_; 
wire _abc_40319_new_n1182_; 
wire _abc_40319_new_n1183_; 
wire _abc_40319_new_n1184_; 
wire _abc_40319_new_n1185_; 
wire _abc_40319_new_n1186_; 
wire _abc_40319_new_n1187_; 
wire _abc_40319_new_n1188_; 
wire _abc_40319_new_n1189_; 
wire _abc_40319_new_n1190_; 
wire _abc_40319_new_n1191_; 
wire _abc_40319_new_n1192_; 
wire _abc_40319_new_n1193_; 
wire _abc_40319_new_n1194_; 
wire _abc_40319_new_n1195_; 
wire _abc_40319_new_n1196_; 
wire _abc_40319_new_n1197_; 
wire _abc_40319_new_n1198_; 
wire _abc_40319_new_n1199_; 
wire _abc_40319_new_n1200_; 
wire _abc_40319_new_n1201_; 
wire _abc_40319_new_n1202_; 
wire _abc_40319_new_n1203_; 
wire _abc_40319_new_n1204_; 
wire _abc_40319_new_n1205_; 
wire _abc_40319_new_n1206_; 
wire _abc_40319_new_n1207_; 
wire _abc_40319_new_n1208_; 
wire _abc_40319_new_n1209_; 
wire _abc_40319_new_n1210_; 
wire _abc_40319_new_n1211_; 
wire _abc_40319_new_n1212_; 
wire _abc_40319_new_n1213_; 
wire _abc_40319_new_n1214_; 
wire _abc_40319_new_n1215_; 
wire _abc_40319_new_n1216_; 
wire _abc_40319_new_n1217_; 
wire _abc_40319_new_n1218_; 
wire _abc_40319_new_n1219_; 
wire _abc_40319_new_n1220_; 
wire _abc_40319_new_n1221_; 
wire _abc_40319_new_n1222_; 
wire _abc_40319_new_n1223_; 
wire _abc_40319_new_n1224_; 
wire _abc_40319_new_n1225_; 
wire _abc_40319_new_n1226_; 
wire _abc_40319_new_n1227_; 
wire _abc_40319_new_n1228_; 
wire _abc_40319_new_n1229_; 
wire _abc_40319_new_n1230_; 
wire _abc_40319_new_n1231_; 
wire _abc_40319_new_n1232_; 
wire _abc_40319_new_n1233_; 
wire _abc_40319_new_n1234_; 
wire _abc_40319_new_n1235_; 
wire _abc_40319_new_n1236_; 
wire _abc_40319_new_n1237_; 
wire _abc_40319_new_n1238_; 
wire _abc_40319_new_n1239_; 
wire _abc_40319_new_n1240_; 
wire _abc_40319_new_n1241_; 
wire _abc_40319_new_n1242_; 
wire _abc_40319_new_n1243_; 
wire _abc_40319_new_n1244_; 
wire _abc_40319_new_n1245_; 
wire _abc_40319_new_n1246_; 
wire _abc_40319_new_n1247_; 
wire _abc_40319_new_n1248_; 
wire _abc_40319_new_n1249_; 
wire _abc_40319_new_n1250_; 
wire _abc_40319_new_n1251_; 
wire _abc_40319_new_n1252_; 
wire _abc_40319_new_n1253_; 
wire _abc_40319_new_n1254_; 
wire _abc_40319_new_n1255_; 
wire _abc_40319_new_n1256_; 
wire _abc_40319_new_n1257_; 
wire _abc_40319_new_n1258_; 
wire _abc_40319_new_n1259_; 
wire _abc_40319_new_n1260_; 
wire _abc_40319_new_n1261_; 
wire _abc_40319_new_n1262_; 
wire _abc_40319_new_n1263_; 
wire _abc_40319_new_n1264_; 
wire _abc_40319_new_n1265_; 
wire _abc_40319_new_n1266_; 
wire _abc_40319_new_n1267_; 
wire _abc_40319_new_n1268_; 
wire _abc_40319_new_n1269_; 
wire _abc_40319_new_n1270_; 
wire _abc_40319_new_n1271_; 
wire _abc_40319_new_n1272_; 
wire _abc_40319_new_n1273_; 
wire _abc_40319_new_n1274_; 
wire _abc_40319_new_n1275_; 
wire _abc_40319_new_n1276_; 
wire _abc_40319_new_n1277_; 
wire _abc_40319_new_n1278_; 
wire _abc_40319_new_n1279_; 
wire _abc_40319_new_n1280_; 
wire _abc_40319_new_n1281_; 
wire _abc_40319_new_n1282_; 
wire _abc_40319_new_n1283_; 
wire _abc_40319_new_n1284_; 
wire _abc_40319_new_n1285_; 
wire _abc_40319_new_n1286_; 
wire _abc_40319_new_n1287_; 
wire _abc_40319_new_n1288_; 
wire _abc_40319_new_n1289_; 
wire _abc_40319_new_n1290_; 
wire _abc_40319_new_n1291_; 
wire _abc_40319_new_n1292_; 
wire _abc_40319_new_n1293_; 
wire _abc_40319_new_n1294_; 
wire _abc_40319_new_n1295_; 
wire _abc_40319_new_n1296_; 
wire _abc_40319_new_n1297_; 
wire _abc_40319_new_n1298_; 
wire _abc_40319_new_n1299_; 
wire _abc_40319_new_n1300_; 
wire _abc_40319_new_n1301_; 
wire _abc_40319_new_n1302_; 
wire _abc_40319_new_n1303_; 
wire _abc_40319_new_n1304_; 
wire _abc_40319_new_n1305_; 
wire _abc_40319_new_n1306_; 
wire _abc_40319_new_n1307_; 
wire _abc_40319_new_n1308_; 
wire _abc_40319_new_n1309_; 
wire _abc_40319_new_n1310_; 
wire _abc_40319_new_n1311_; 
wire _abc_40319_new_n1312_; 
wire _abc_40319_new_n1313_; 
wire _abc_40319_new_n1314_; 
wire _abc_40319_new_n1315_; 
wire _abc_40319_new_n1316_; 
wire _abc_40319_new_n1317_; 
wire _abc_40319_new_n1318_; 
wire _abc_40319_new_n1319_; 
wire _abc_40319_new_n1320_; 
wire _abc_40319_new_n1321_; 
wire _abc_40319_new_n1322_; 
wire _abc_40319_new_n1323_; 
wire _abc_40319_new_n1324_; 
wire _abc_40319_new_n1325_; 
wire _abc_40319_new_n1326_; 
wire _abc_40319_new_n1327_; 
wire _abc_40319_new_n1328_; 
wire _abc_40319_new_n1329_; 
wire _abc_40319_new_n1330_; 
wire _abc_40319_new_n1331_; 
wire _abc_40319_new_n1332_; 
wire _abc_40319_new_n1333_; 
wire _abc_40319_new_n1334_; 
wire _abc_40319_new_n1335_; 
wire _abc_40319_new_n1336_; 
wire _abc_40319_new_n1337_; 
wire _abc_40319_new_n1338_; 
wire _abc_40319_new_n1339_; 
wire _abc_40319_new_n1340_; 
wire _abc_40319_new_n1341_; 
wire _abc_40319_new_n1342_; 
wire _abc_40319_new_n1343_; 
wire _abc_40319_new_n1344_; 
wire _abc_40319_new_n1345_; 
wire _abc_40319_new_n1346_; 
wire _abc_40319_new_n1347_; 
wire _abc_40319_new_n1348_; 
wire _abc_40319_new_n1349_; 
wire _abc_40319_new_n1350_; 
wire _abc_40319_new_n1351_; 
wire _abc_40319_new_n1352_; 
wire _abc_40319_new_n1353_; 
wire _abc_40319_new_n1354_; 
wire _abc_40319_new_n1355_; 
wire _abc_40319_new_n1356_; 
wire _abc_40319_new_n1357_; 
wire _abc_40319_new_n1358_; 
wire _abc_40319_new_n1359_; 
wire _abc_40319_new_n1360_; 
wire _abc_40319_new_n1361_; 
wire _abc_40319_new_n1362_; 
wire _abc_40319_new_n1363_; 
wire _abc_40319_new_n1364_; 
wire _abc_40319_new_n1365_; 
wire _abc_40319_new_n1366_; 
wire _abc_40319_new_n1367_; 
wire _abc_40319_new_n1368_; 
wire _abc_40319_new_n1369_; 
wire _abc_40319_new_n1370_; 
wire _abc_40319_new_n1371_; 
wire _abc_40319_new_n1372_; 
wire _abc_40319_new_n1373_; 
wire _abc_40319_new_n1374_; 
wire _abc_40319_new_n1375_; 
wire _abc_40319_new_n1376_; 
wire _abc_40319_new_n1377_; 
wire _abc_40319_new_n1378_; 
wire _abc_40319_new_n1379_; 
wire _abc_40319_new_n1380_; 
wire _abc_40319_new_n1381_; 
wire _abc_40319_new_n1382_; 
wire _abc_40319_new_n1383_; 
wire _abc_40319_new_n1384_; 
wire _abc_40319_new_n1385_; 
wire _abc_40319_new_n1386_; 
wire _abc_40319_new_n1387_; 
wire _abc_40319_new_n1388_; 
wire _abc_40319_new_n1389_; 
wire _abc_40319_new_n1390_; 
wire _abc_40319_new_n1391_; 
wire _abc_40319_new_n1392_; 
wire _abc_40319_new_n1393_; 
wire _abc_40319_new_n1394_; 
wire _abc_40319_new_n1395_; 
wire _abc_40319_new_n1396_; 
wire _abc_40319_new_n1397_; 
wire _abc_40319_new_n1398_; 
wire _abc_40319_new_n1399_; 
wire _abc_40319_new_n1400_; 
wire _abc_40319_new_n1401_; 
wire _abc_40319_new_n1402_; 
wire _abc_40319_new_n1403_; 
wire _abc_40319_new_n1404_; 
wire _abc_40319_new_n1405_; 
wire _abc_40319_new_n1406_; 
wire _abc_40319_new_n1407_; 
wire _abc_40319_new_n1408_; 
wire _abc_40319_new_n1409_; 
wire _abc_40319_new_n1410_; 
wire _abc_40319_new_n1411_; 
wire _abc_40319_new_n1412_; 
wire _abc_40319_new_n1413_; 
wire _abc_40319_new_n1414_; 
wire _abc_40319_new_n1415_; 
wire _abc_40319_new_n1416_; 
wire _abc_40319_new_n1417_; 
wire _abc_40319_new_n1418_; 
wire _abc_40319_new_n1419_; 
wire _abc_40319_new_n1420_; 
wire _abc_40319_new_n1421_; 
wire _abc_40319_new_n1422_; 
wire _abc_40319_new_n1423_; 
wire _abc_40319_new_n1424_; 
wire _abc_40319_new_n1425_; 
wire _abc_40319_new_n1426_; 
wire _abc_40319_new_n1427_; 
wire _abc_40319_new_n1428_; 
wire _abc_40319_new_n1429_; 
wire _abc_40319_new_n1430_; 
wire _abc_40319_new_n1431_; 
wire _abc_40319_new_n1432_; 
wire _abc_40319_new_n1433_; 
wire _abc_40319_new_n1434_; 
wire _abc_40319_new_n1435_; 
wire _abc_40319_new_n1436_; 
wire _abc_40319_new_n1437_; 
wire _abc_40319_new_n1438_; 
wire _abc_40319_new_n1439_; 
wire _abc_40319_new_n1440_; 
wire _abc_40319_new_n1441_; 
wire _abc_40319_new_n1442_; 
wire _abc_40319_new_n1443_; 
wire _abc_40319_new_n1444_; 
wire _abc_40319_new_n1445_; 
wire _abc_40319_new_n1446_; 
wire _abc_40319_new_n1447_; 
wire _abc_40319_new_n1448_; 
wire _abc_40319_new_n1449_; 
wire _abc_40319_new_n1450_; 
wire _abc_40319_new_n1451_; 
wire _abc_40319_new_n1452_; 
wire _abc_40319_new_n1453_; 
wire _abc_40319_new_n1454_; 
wire _abc_40319_new_n1455_; 
wire _abc_40319_new_n1456_; 
wire _abc_40319_new_n1457_; 
wire _abc_40319_new_n1458_; 
wire _abc_40319_new_n1459_; 
wire _abc_40319_new_n1460_; 
wire _abc_40319_new_n1461_; 
wire _abc_40319_new_n1462_; 
wire _abc_40319_new_n1463_; 
wire _abc_40319_new_n1464_; 
wire _abc_40319_new_n1465_; 
wire _abc_40319_new_n1466_; 
wire _abc_40319_new_n1467_; 
wire _abc_40319_new_n1468_; 
wire _abc_40319_new_n1469_; 
wire _abc_40319_new_n1470_; 
wire _abc_40319_new_n1471_; 
wire _abc_40319_new_n1472_; 
wire _abc_40319_new_n1473_; 
wire _abc_40319_new_n1474_; 
wire _abc_40319_new_n1475_; 
wire _abc_40319_new_n1476_; 
wire _abc_40319_new_n1477_; 
wire _abc_40319_new_n1478_; 
wire _abc_40319_new_n1479_; 
wire _abc_40319_new_n1480_; 
wire _abc_40319_new_n1481_; 
wire _abc_40319_new_n1482_; 
wire _abc_40319_new_n1483_; 
wire _abc_40319_new_n1484_; 
wire _abc_40319_new_n1485_; 
wire _abc_40319_new_n1486_; 
wire _abc_40319_new_n1487_; 
wire _abc_40319_new_n1488_; 
wire _abc_40319_new_n1489_; 
wire _abc_40319_new_n1490_; 
wire _abc_40319_new_n1491_; 
wire _abc_40319_new_n1492_; 
wire _abc_40319_new_n1493_; 
wire _abc_40319_new_n1494_; 
wire _abc_40319_new_n1495_; 
wire _abc_40319_new_n1496_; 
wire _abc_40319_new_n1497_; 
wire _abc_40319_new_n1498_; 
wire _abc_40319_new_n1499_; 
wire _abc_40319_new_n1500_; 
wire _abc_40319_new_n1501_; 
wire _abc_40319_new_n1502_; 
wire _abc_40319_new_n1503_; 
wire _abc_40319_new_n1504_; 
wire _abc_40319_new_n1505_; 
wire _abc_40319_new_n1506_; 
wire _abc_40319_new_n1507_; 
wire _abc_40319_new_n1508_; 
wire _abc_40319_new_n1509_; 
wire _abc_40319_new_n1510_; 
wire _abc_40319_new_n1512_; 
wire _abc_40319_new_n1513_; 
wire _abc_40319_new_n1514_; 
wire _abc_40319_new_n1515_; 
wire _abc_40319_new_n1516_; 
wire _abc_40319_new_n1517_; 
wire _abc_40319_new_n1518_; 
wire _abc_40319_new_n1519_; 
wire _abc_40319_new_n1520_; 
wire _abc_40319_new_n1521_; 
wire _abc_40319_new_n1522_; 
wire _abc_40319_new_n1523_; 
wire _abc_40319_new_n1525_; 
wire _abc_40319_new_n1526_; 
wire _abc_40319_new_n1527_; 
wire _abc_40319_new_n1528_; 
wire _abc_40319_new_n1529_; 
wire _abc_40319_new_n1530_; 
wire _abc_40319_new_n1531_; 
wire _abc_40319_new_n1532_; 
wire _abc_40319_new_n1533_; 
wire _abc_40319_new_n1534_; 
wire _abc_40319_new_n1536_; 
wire _abc_40319_new_n1537_; 
wire _abc_40319_new_n1538_; 
wire _abc_40319_new_n1539_; 
wire _abc_40319_new_n1540_; 
wire _abc_40319_new_n1541_; 
wire _abc_40319_new_n1542_; 
wire _abc_40319_new_n1543_; 
wire _abc_40319_new_n1544_; 
wire _abc_40319_new_n1545_; 
wire _abc_40319_new_n1547_; 
wire _abc_40319_new_n1548_; 
wire _abc_40319_new_n1549_; 
wire _abc_40319_new_n1550_; 
wire _abc_40319_new_n1551_; 
wire _abc_40319_new_n1552_; 
wire _abc_40319_new_n1553_; 
wire _abc_40319_new_n1554_; 
wire _abc_40319_new_n1555_; 
wire _abc_40319_new_n1556_; 
wire _abc_40319_new_n1557_; 
wire _abc_40319_new_n1558_; 
wire _abc_40319_new_n1559_; 
wire _abc_40319_new_n1560_; 
wire _abc_40319_new_n1561_; 
wire _abc_40319_new_n1563_; 
wire _abc_40319_new_n1564_; 
wire _abc_40319_new_n1565_; 
wire _abc_40319_new_n1566_; 
wire _abc_40319_new_n1567_; 
wire _abc_40319_new_n1568_; 
wire _abc_40319_new_n1569_; 
wire _abc_40319_new_n1570_; 
wire _abc_40319_new_n1571_; 
wire _abc_40319_new_n1572_; 
wire _abc_40319_new_n1573_; 
wire _abc_40319_new_n1574_; 
wire _abc_40319_new_n1575_; 
wire _abc_40319_new_n1577_; 
wire _abc_40319_new_n1578_; 
wire _abc_40319_new_n1579_; 
wire _abc_40319_new_n1580_; 
wire _abc_40319_new_n1581_; 
wire _abc_40319_new_n1582_; 
wire _abc_40319_new_n1583_; 
wire _abc_40319_new_n1584_; 
wire _abc_40319_new_n1585_; 
wire _abc_40319_new_n1586_; 
wire _abc_40319_new_n1587_; 
wire _abc_40319_new_n1588_; 
wire _abc_40319_new_n1589_; 
wire _abc_40319_new_n1590_; 
wire _abc_40319_new_n1591_; 
wire _abc_40319_new_n1592_; 
wire _abc_40319_new_n1593_; 
wire _abc_40319_new_n1594_; 
wire _abc_40319_new_n1595_; 
wire _abc_40319_new_n1596_; 
wire _abc_40319_new_n1597_; 
wire _abc_40319_new_n1598_; 
wire _abc_40319_new_n1599_; 
wire _abc_40319_new_n1600_; 
wire _abc_40319_new_n1601_; 
wire _abc_40319_new_n1602_; 
wire _abc_40319_new_n1603_; 
wire _abc_40319_new_n1604_; 
wire _abc_40319_new_n1605_; 
wire _abc_40319_new_n1607_; 
wire _abc_40319_new_n1608_; 
wire _abc_40319_new_n1609_; 
wire _abc_40319_new_n1610_; 
wire _abc_40319_new_n1611_; 
wire _abc_40319_new_n1612_; 
wire _abc_40319_new_n1613_; 
wire _abc_40319_new_n1614_; 
wire _abc_40319_new_n1615_; 
wire _abc_40319_new_n1616_; 
wire _abc_40319_new_n1617_; 
wire _abc_40319_new_n1618_; 
wire _abc_40319_new_n1619_; 
wire _abc_40319_new_n1621_; 
wire _abc_40319_new_n1622_; 
wire _abc_40319_new_n1623_; 
wire _abc_40319_new_n1624_; 
wire _abc_40319_new_n1625_; 
wire _abc_40319_new_n1626_; 
wire _abc_40319_new_n1627_; 
wire _abc_40319_new_n1628_; 
wire _abc_40319_new_n1630_; 
wire _abc_40319_new_n1631_; 
wire _abc_40319_new_n1632_; 
wire _abc_40319_new_n1633_; 
wire _abc_40319_new_n1634_; 
wire _abc_40319_new_n1635_; 
wire _abc_40319_new_n1636_; 
wire _abc_40319_new_n1637_; 
wire _abc_40319_new_n1638_; 
wire _abc_40319_new_n1639_; 
wire _abc_40319_new_n1640_; 
wire _abc_40319_new_n1641_; 
wire _abc_40319_new_n1642_; 
wire _abc_40319_new_n1643_; 
wire _abc_40319_new_n1645_; 
wire _abc_40319_new_n1646_; 
wire _abc_40319_new_n1647_; 
wire _abc_40319_new_n1648_; 
wire _abc_40319_new_n1649_; 
wire _abc_40319_new_n1650_; 
wire _abc_40319_new_n1651_; 
wire _abc_40319_new_n1652_; 
wire _abc_40319_new_n1653_; 
wire _abc_40319_new_n1654_; 
wire _abc_40319_new_n1655_; 
wire _abc_40319_new_n1656_; 
wire _abc_40319_new_n1657_; 
wire _abc_40319_new_n1658_; 
wire _abc_40319_new_n1660_; 
wire _abc_40319_new_n1661_; 
wire _abc_40319_new_n1662_; 
wire _abc_40319_new_n1663_; 
wire _abc_40319_new_n1664_; 
wire _abc_40319_new_n1665_; 
wire _abc_40319_new_n1666_; 
wire _abc_40319_new_n1667_; 
wire _abc_40319_new_n1668_; 
wire _abc_40319_new_n1669_; 
wire _abc_40319_new_n1670_; 
wire _abc_40319_new_n1671_; 
wire _abc_40319_new_n1673_; 
wire _abc_40319_new_n1674_; 
wire _abc_40319_new_n1675_; 
wire _abc_40319_new_n1676_; 
wire _abc_40319_new_n1677_; 
wire _abc_40319_new_n1678_; 
wire _abc_40319_new_n1679_; 
wire _abc_40319_new_n1680_; 
wire _abc_40319_new_n1681_; 
wire _abc_40319_new_n1682_; 
wire _abc_40319_new_n1683_; 
wire _abc_40319_new_n1685_; 
wire _abc_40319_new_n1686_; 
wire _abc_40319_new_n1687_; 
wire _abc_40319_new_n1688_; 
wire _abc_40319_new_n1689_; 
wire _abc_40319_new_n1690_; 
wire _abc_40319_new_n1691_; 
wire _abc_40319_new_n1692_; 
wire _abc_40319_new_n1694_; 
wire _abc_40319_new_n1695_; 
wire _abc_40319_new_n1696_; 
wire _abc_40319_new_n1697_; 
wire _abc_40319_new_n1698_; 
wire _abc_40319_new_n1699_; 
wire _abc_40319_new_n1700_; 
wire _abc_40319_new_n1701_; 
wire _abc_40319_new_n1702_; 
wire _abc_40319_new_n1703_; 
wire _abc_40319_new_n1704_; 
wire _abc_40319_new_n1705_; 
wire _abc_40319_new_n1707_; 
wire _abc_40319_new_n1708_; 
wire _abc_40319_new_n1709_; 
wire _abc_40319_new_n1710_; 
wire _abc_40319_new_n1711_; 
wire _abc_40319_new_n1712_; 
wire _abc_40319_new_n1713_; 
wire _abc_40319_new_n1714_; 
wire _abc_40319_new_n1715_; 
wire _abc_40319_new_n1716_; 
wire _abc_40319_new_n1717_; 
wire _abc_40319_new_n1719_; 
wire _abc_40319_new_n1720_; 
wire _abc_40319_new_n1721_; 
wire _abc_40319_new_n1722_; 
wire _abc_40319_new_n1723_; 
wire _abc_40319_new_n1724_; 
wire _abc_40319_new_n1725_; 
wire _abc_40319_new_n1726_; 
wire _abc_40319_new_n1727_; 
wire _abc_40319_new_n1728_; 
wire _abc_40319_new_n1729_; 
wire _abc_40319_new_n1730_; 
wire _abc_40319_new_n1732_; 
wire _abc_40319_new_n1733_; 
wire _abc_40319_new_n1734_; 
wire _abc_40319_new_n1735_; 
wire _abc_40319_new_n1736_; 
wire _abc_40319_new_n1737_; 
wire _abc_40319_new_n1738_; 
wire _abc_40319_new_n1739_; 
wire _abc_40319_new_n1740_; 
wire _abc_40319_new_n1741_; 
wire _abc_40319_new_n1742_; 
wire _abc_40319_new_n1743_; 
wire _abc_40319_new_n1744_; 
wire _abc_40319_new_n1746_; 
wire _abc_40319_new_n1747_; 
wire _abc_40319_new_n1748_; 
wire _abc_40319_new_n1749_; 
wire _abc_40319_new_n1750_; 
wire _abc_40319_new_n1751_; 
wire _abc_40319_new_n1752_; 
wire _abc_40319_new_n1753_; 
wire _abc_40319_new_n1754_; 
wire _abc_40319_new_n1755_; 
wire _abc_40319_new_n1757_; 
wire _abc_40319_new_n1758_; 
wire _abc_40319_new_n1759_; 
wire _abc_40319_new_n1760_; 
wire _abc_40319_new_n1761_; 
wire _abc_40319_new_n1762_; 
wire _abc_40319_new_n1763_; 
wire _abc_40319_new_n1764_; 
wire _abc_40319_new_n1765_; 
wire _abc_40319_new_n1767_; 
wire _abc_40319_new_n1768_; 
wire _abc_40319_new_n1769_; 
wire _abc_40319_new_n1770_; 
wire _abc_40319_new_n1771_; 
wire _abc_40319_new_n1772_; 
wire _abc_40319_new_n1773_; 
wire _abc_40319_new_n1774_; 
wire _abc_40319_new_n1775_; 
wire _abc_40319_new_n1776_; 
wire _abc_40319_new_n1777_; 
wire _abc_40319_new_n1778_; 
wire _abc_40319_new_n1779_; 
wire _abc_40319_new_n1781_; 
wire _abc_40319_new_n1782_; 
wire _abc_40319_new_n1783_; 
wire _abc_40319_new_n1784_; 
wire _abc_40319_new_n1785_; 
wire _abc_40319_new_n1786_; 
wire _abc_40319_new_n1787_; 
wire _abc_40319_new_n1788_; 
wire _abc_40319_new_n1789_; 
wire _abc_40319_new_n1790_; 
wire _abc_40319_new_n1791_; 
wire _abc_40319_new_n1793_; 
wire _abc_40319_new_n1794_; 
wire _abc_40319_new_n1795_; 
wire _abc_40319_new_n1796_; 
wire _abc_40319_new_n1797_; 
wire _abc_40319_new_n1798_; 
wire _abc_40319_new_n1799_; 
wire _abc_40319_new_n1800_; 
wire _abc_40319_new_n1801_; 
wire _abc_40319_new_n1802_; 
wire _abc_40319_new_n1803_; 
wire _abc_40319_new_n1805_; 
wire _abc_40319_new_n1806_; 
wire _abc_40319_new_n1807_; 
wire _abc_40319_new_n1808_; 
wire _abc_40319_new_n1809_; 
wire _abc_40319_new_n1810_; 
wire _abc_40319_new_n1811_; 
wire _abc_40319_new_n1812_; 
wire _abc_40319_new_n1813_; 
wire _abc_40319_new_n1814_; 
wire _abc_40319_new_n1815_; 
wire _abc_40319_new_n1816_; 
wire _abc_40319_new_n1818_; 
wire _abc_40319_new_n1819_; 
wire _abc_40319_new_n1820_; 
wire _abc_40319_new_n1821_; 
wire _abc_40319_new_n1822_; 
wire _abc_40319_new_n1823_; 
wire _abc_40319_new_n1824_; 
wire _abc_40319_new_n1825_; 
wire _abc_40319_new_n1826_; 
wire _abc_40319_new_n1827_; 
wire _abc_40319_new_n1828_; 
wire _abc_40319_new_n1830_; 
wire _abc_40319_new_n1831_; 
wire _abc_40319_new_n1832_; 
wire _abc_40319_new_n1833_; 
wire _abc_40319_new_n1834_; 
wire _abc_40319_new_n1835_; 
wire _abc_40319_new_n1836_; 
wire _abc_40319_new_n1837_; 
wire _abc_40319_new_n1838_; 
wire _abc_40319_new_n1839_; 
wire _abc_40319_new_n1840_; 
wire _abc_40319_new_n1842_; 
wire _abc_40319_new_n1843_; 
wire _abc_40319_new_n1844_; 
wire _abc_40319_new_n1845_; 
wire _abc_40319_new_n1846_; 
wire _abc_40319_new_n1847_; 
wire _abc_40319_new_n1848_; 
wire _abc_40319_new_n1849_; 
wire _abc_40319_new_n1850_; 
wire _abc_40319_new_n1851_; 
wire _abc_40319_new_n1852_; 
wire _abc_40319_new_n1853_; 
wire _abc_40319_new_n1854_; 
wire _abc_40319_new_n1855_; 
wire _abc_40319_new_n1856_; 
wire _abc_40319_new_n1858_; 
wire _abc_40319_new_n1859_; 
wire _abc_40319_new_n1860_; 
wire _abc_40319_new_n1861_; 
wire _abc_40319_new_n1862_; 
wire _abc_40319_new_n1863_; 
wire _abc_40319_new_n1864_; 
wire _abc_40319_new_n1865_; 
wire _abc_40319_new_n1866_; 
wire _abc_40319_new_n1867_; 
wire _abc_40319_new_n1868_; 
wire _abc_40319_new_n1870_; 
wire _abc_40319_new_n1871_; 
wire _abc_40319_new_n1872_; 
wire _abc_40319_new_n1873_; 
wire _abc_40319_new_n1874_; 
wire _abc_40319_new_n1875_; 
wire _abc_40319_new_n1876_; 
wire _abc_40319_new_n1877_; 
wire _abc_40319_new_n1878_; 
wire _abc_40319_new_n1879_; 
wire _abc_40319_new_n1880_; 
wire _abc_40319_new_n1881_; 
wire _abc_40319_new_n1882_; 
wire _abc_40319_new_n1883_; 
wire _abc_40319_new_n1884_; 
wire _abc_40319_new_n1885_; 
wire _abc_40319_new_n1886_; 
wire _abc_40319_new_n1887_; 
wire _abc_40319_new_n1888_; 
wire _abc_40319_new_n1889_; 
wire _abc_40319_new_n1890_; 
wire _abc_40319_new_n1891_; 
wire _abc_40319_new_n1892_; 
wire _abc_40319_new_n1893_; 
wire _abc_40319_new_n1894_; 
wire _abc_40319_new_n1895_; 
wire _abc_40319_new_n1896_; 
wire _abc_40319_new_n1897_; 
wire _abc_40319_new_n1898_; 
wire _abc_40319_new_n1899_; 
wire _abc_40319_new_n1900_; 
wire _abc_40319_new_n1901_; 
wire _abc_40319_new_n1902_; 
wire _abc_40319_new_n1903_; 
wire _abc_40319_new_n1904_; 
wire _abc_40319_new_n1905_; 
wire _abc_40319_new_n1906_; 
wire _abc_40319_new_n1907_; 
wire _abc_40319_new_n1908_; 
wire _abc_40319_new_n1909_; 
wire _abc_40319_new_n1910_; 
wire _abc_40319_new_n1911_; 
wire _abc_40319_new_n1912_; 
wire _abc_40319_new_n1913_; 
wire _abc_40319_new_n1914_; 
wire _abc_40319_new_n1915_; 
wire _abc_40319_new_n1916_; 
wire _abc_40319_new_n1917_; 
wire _abc_40319_new_n1918_; 
wire _abc_40319_new_n1919_; 
wire _abc_40319_new_n1920_; 
wire _abc_40319_new_n1921_; 
wire _abc_40319_new_n1922_; 
wire _abc_40319_new_n1923_; 
wire _abc_40319_new_n1924_; 
wire _abc_40319_new_n1925_; 
wire _abc_40319_new_n1926_; 
wire _abc_40319_new_n1927_; 
wire _abc_40319_new_n1928_; 
wire _abc_40319_new_n1929_; 
wire _abc_40319_new_n1930_; 
wire _abc_40319_new_n1931_; 
wire _abc_40319_new_n1932_; 
wire _abc_40319_new_n1933_; 
wire _abc_40319_new_n1934_; 
wire _abc_40319_new_n1935_; 
wire _abc_40319_new_n1936_; 
wire _abc_40319_new_n1937_; 
wire _abc_40319_new_n1938_; 
wire _abc_40319_new_n1939_; 
wire _abc_40319_new_n1940_; 
wire _abc_40319_new_n1941_; 
wire _abc_40319_new_n1942_; 
wire _abc_40319_new_n1943_; 
wire _abc_40319_new_n1944_; 
wire _abc_40319_new_n1945_; 
wire _abc_40319_new_n1946_; 
wire _abc_40319_new_n1947_; 
wire _abc_40319_new_n1948_; 
wire _abc_40319_new_n1949_; 
wire _abc_40319_new_n1950_; 
wire _abc_40319_new_n1951_; 
wire _abc_40319_new_n1952_; 
wire _abc_40319_new_n1953_; 
wire _abc_40319_new_n1954_; 
wire _abc_40319_new_n1955_; 
wire _abc_40319_new_n1956_; 
wire _abc_40319_new_n1957_; 
wire _abc_40319_new_n1958_; 
wire _abc_40319_new_n1959_; 
wire _abc_40319_new_n1960_; 
wire _abc_40319_new_n1961_; 
wire _abc_40319_new_n1962_; 
wire _abc_40319_new_n1963_; 
wire _abc_40319_new_n1964_; 
wire _abc_40319_new_n1965_; 
wire _abc_40319_new_n1966_; 
wire _abc_40319_new_n1967_; 
wire _abc_40319_new_n1968_; 
wire _abc_40319_new_n1969_; 
wire _abc_40319_new_n1970_; 
wire _abc_40319_new_n1971_; 
wire _abc_40319_new_n1972_; 
wire _abc_40319_new_n1973_; 
wire _abc_40319_new_n1974_; 
wire _abc_40319_new_n1975_; 
wire _abc_40319_new_n1976_; 
wire _abc_40319_new_n1977_; 
wire _abc_40319_new_n1978_; 
wire _abc_40319_new_n1979_; 
wire _abc_40319_new_n1980_; 
wire _abc_40319_new_n1981_; 
wire _abc_40319_new_n1982_; 
wire _abc_40319_new_n1983_; 
wire _abc_40319_new_n1984_; 
wire _abc_40319_new_n1985_; 
wire _abc_40319_new_n1986_; 
wire _abc_40319_new_n1987_; 
wire _abc_40319_new_n1988_; 
wire _abc_40319_new_n1989_; 
wire _abc_40319_new_n1990_; 
wire _abc_40319_new_n1991_; 
wire _abc_40319_new_n1992_; 
wire _abc_40319_new_n1993_; 
wire _abc_40319_new_n1994_; 
wire _abc_40319_new_n1995_; 
wire _abc_40319_new_n1996_; 
wire _abc_40319_new_n1997_; 
wire _abc_40319_new_n1998_; 
wire _abc_40319_new_n1999_; 
wire _abc_40319_new_n2000_; 
wire _abc_40319_new_n2001_; 
wire _abc_40319_new_n2002_; 
wire _abc_40319_new_n2003_; 
wire _abc_40319_new_n2004_; 
wire _abc_40319_new_n2005_; 
wire _abc_40319_new_n2006_; 
wire _abc_40319_new_n2007_; 
wire _abc_40319_new_n2008_; 
wire _abc_40319_new_n2009_; 
wire _abc_40319_new_n2010_; 
wire _abc_40319_new_n2011_; 
wire _abc_40319_new_n2012_; 
wire _abc_40319_new_n2013_; 
wire _abc_40319_new_n2014_; 
wire _abc_40319_new_n2015_; 
wire _abc_40319_new_n2016_; 
wire _abc_40319_new_n2017_; 
wire _abc_40319_new_n2018_; 
wire _abc_40319_new_n2019_; 
wire _abc_40319_new_n2020_; 
wire _abc_40319_new_n2021_; 
wire _abc_40319_new_n2022_; 
wire _abc_40319_new_n2023_; 
wire _abc_40319_new_n2024_; 
wire _abc_40319_new_n2025_; 
wire _abc_40319_new_n2026_; 
wire _abc_40319_new_n2027_; 
wire _abc_40319_new_n2028_; 
wire _abc_40319_new_n2029_; 
wire _abc_40319_new_n2030_; 
wire _abc_40319_new_n2031_; 
wire _abc_40319_new_n2032_; 
wire _abc_40319_new_n2033_; 
wire _abc_40319_new_n2034_; 
wire _abc_40319_new_n2035_; 
wire _abc_40319_new_n2036_; 
wire _abc_40319_new_n2037_; 
wire _abc_40319_new_n2038_; 
wire _abc_40319_new_n2039_; 
wire _abc_40319_new_n2040_; 
wire _abc_40319_new_n2041_; 
wire _abc_40319_new_n2042_; 
wire _abc_40319_new_n2043_; 
wire _abc_40319_new_n2044_; 
wire _abc_40319_new_n2045_; 
wire _abc_40319_new_n2046_; 
wire _abc_40319_new_n2047_; 
wire _abc_40319_new_n2048_; 
wire _abc_40319_new_n2049_; 
wire _abc_40319_new_n2050_; 
wire _abc_40319_new_n2051_; 
wire _abc_40319_new_n2052_; 
wire _abc_40319_new_n2053_; 
wire _abc_40319_new_n2054_; 
wire _abc_40319_new_n2055_; 
wire _abc_40319_new_n2056_; 
wire _abc_40319_new_n2057_; 
wire _abc_40319_new_n2058_; 
wire _abc_40319_new_n2059_; 
wire _abc_40319_new_n2060_; 
wire _abc_40319_new_n2061_; 
wire _abc_40319_new_n2062_; 
wire _abc_40319_new_n2063_; 
wire _abc_40319_new_n2064_; 
wire _abc_40319_new_n2065_; 
wire _abc_40319_new_n2066_; 
wire _abc_40319_new_n2067_; 
wire _abc_40319_new_n2068_; 
wire _abc_40319_new_n2069_; 
wire _abc_40319_new_n2070_; 
wire _abc_40319_new_n2071_; 
wire _abc_40319_new_n2072_; 
wire _abc_40319_new_n2073_; 
wire _abc_40319_new_n2074_; 
wire _abc_40319_new_n2075_; 
wire _abc_40319_new_n2076_; 
wire _abc_40319_new_n2077_; 
wire _abc_40319_new_n2078_; 
wire _abc_40319_new_n2079_; 
wire _abc_40319_new_n2080_; 
wire _abc_40319_new_n2081_; 
wire _abc_40319_new_n2082_; 
wire _abc_40319_new_n2083_; 
wire _abc_40319_new_n2084_; 
wire _abc_40319_new_n2085_; 
wire _abc_40319_new_n2086_; 
wire _abc_40319_new_n2087_; 
wire _abc_40319_new_n2088_; 
wire _abc_40319_new_n2089_; 
wire _abc_40319_new_n2090_; 
wire _abc_40319_new_n2091_; 
wire _abc_40319_new_n2092_; 
wire _abc_40319_new_n2093_; 
wire _abc_40319_new_n2094_; 
wire _abc_40319_new_n2095_; 
wire _abc_40319_new_n2096_; 
wire _abc_40319_new_n2097_; 
wire _abc_40319_new_n2098_; 
wire _abc_40319_new_n2099_; 
wire _abc_40319_new_n2100_; 
wire _abc_40319_new_n2101_; 
wire _abc_40319_new_n2102_; 
wire _abc_40319_new_n2103_; 
wire _abc_40319_new_n2104_; 
wire _abc_40319_new_n2105_; 
wire _abc_40319_new_n2106_; 
wire _abc_40319_new_n2107_; 
wire _abc_40319_new_n2108_; 
wire _abc_40319_new_n2109_; 
wire _abc_40319_new_n2110_; 
wire _abc_40319_new_n2111_; 
wire _abc_40319_new_n2112_; 
wire _abc_40319_new_n2113_; 
wire _abc_40319_new_n2114_; 
wire _abc_40319_new_n2115_; 
wire _abc_40319_new_n2116_; 
wire _abc_40319_new_n2117_; 
wire _abc_40319_new_n2118_; 
wire _abc_40319_new_n2119_; 
wire _abc_40319_new_n2120_; 
wire _abc_40319_new_n2121_; 
wire _abc_40319_new_n2122_; 
wire _abc_40319_new_n2123_; 
wire _abc_40319_new_n2124_; 
wire _abc_40319_new_n2125_; 
wire _abc_40319_new_n2126_; 
wire _abc_40319_new_n2127_; 
wire _abc_40319_new_n2128_; 
wire _abc_40319_new_n2129_; 
wire _abc_40319_new_n2130_; 
wire _abc_40319_new_n2131_; 
wire _abc_40319_new_n2132_; 
wire _abc_40319_new_n2133_; 
wire _abc_40319_new_n2134_; 
wire _abc_40319_new_n2135_; 
wire _abc_40319_new_n2136_; 
wire _abc_40319_new_n2137_; 
wire _abc_40319_new_n2138_; 
wire _abc_40319_new_n2139_; 
wire _abc_40319_new_n2140_; 
wire _abc_40319_new_n2141_; 
wire _abc_40319_new_n2142_; 
wire _abc_40319_new_n2143_; 
wire _abc_40319_new_n2144_; 
wire _abc_40319_new_n2145_; 
wire _abc_40319_new_n2146_; 
wire _abc_40319_new_n2147_; 
wire _abc_40319_new_n2148_; 
wire _abc_40319_new_n2149_; 
wire _abc_40319_new_n2150_; 
wire _abc_40319_new_n2151_; 
wire _abc_40319_new_n2152_; 
wire _abc_40319_new_n2153_; 
wire _abc_40319_new_n2154_; 
wire _abc_40319_new_n2155_; 
wire _abc_40319_new_n2156_; 
wire _abc_40319_new_n2157_; 
wire _abc_40319_new_n2158_; 
wire _abc_40319_new_n2159_; 
wire _abc_40319_new_n2160_; 
wire _abc_40319_new_n2161_; 
wire _abc_40319_new_n2162_; 
wire _abc_40319_new_n2163_; 
wire _abc_40319_new_n2164_; 
wire _abc_40319_new_n2165_; 
wire _abc_40319_new_n2166_; 
wire _abc_40319_new_n2167_; 
wire _abc_40319_new_n2168_; 
wire _abc_40319_new_n2169_; 
wire _abc_40319_new_n2170_; 
wire _abc_40319_new_n2171_; 
wire _abc_40319_new_n2172_; 
wire _abc_40319_new_n2173_; 
wire _abc_40319_new_n2174_; 
wire _abc_40319_new_n2175_; 
wire _abc_40319_new_n2176_; 
wire _abc_40319_new_n2177_; 
wire _abc_40319_new_n2178_; 
wire _abc_40319_new_n2179_; 
wire _abc_40319_new_n2180_; 
wire _abc_40319_new_n2181_; 
wire _abc_40319_new_n2182_; 
wire _abc_40319_new_n2183_; 
wire _abc_40319_new_n2184_; 
wire _abc_40319_new_n2185_; 
wire _abc_40319_new_n2186_; 
wire _abc_40319_new_n2187_; 
wire _abc_40319_new_n2188_; 
wire _abc_40319_new_n2189_; 
wire _abc_40319_new_n2190_; 
wire _abc_40319_new_n2191_; 
wire _abc_40319_new_n2192_; 
wire _abc_40319_new_n2193_; 
wire _abc_40319_new_n2194_; 
wire _abc_40319_new_n2195_; 
wire _abc_40319_new_n2196_; 
wire _abc_40319_new_n2197_; 
wire _abc_40319_new_n2198_; 
wire _abc_40319_new_n2199_; 
wire _abc_40319_new_n2200_; 
wire _abc_40319_new_n2201_; 
wire _abc_40319_new_n2202_; 
wire _abc_40319_new_n2203_; 
wire _abc_40319_new_n2204_; 
wire _abc_40319_new_n2205_; 
wire _abc_40319_new_n2206_; 
wire _abc_40319_new_n2207_; 
wire _abc_40319_new_n2208_; 
wire _abc_40319_new_n2209_; 
wire _abc_40319_new_n2210_; 
wire _abc_40319_new_n2211_; 
wire _abc_40319_new_n2212_; 
wire _abc_40319_new_n2213_; 
wire _abc_40319_new_n2214_; 
wire _abc_40319_new_n2215_; 
wire _abc_40319_new_n2216_; 
wire _abc_40319_new_n2217_; 
wire _abc_40319_new_n2218_; 
wire _abc_40319_new_n2219_; 
wire _abc_40319_new_n2220_; 
wire _abc_40319_new_n2221_; 
wire _abc_40319_new_n2222_; 
wire _abc_40319_new_n2223_; 
wire _abc_40319_new_n2224_; 
wire _abc_40319_new_n2225_; 
wire _abc_40319_new_n2226_; 
wire _abc_40319_new_n2227_; 
wire _abc_40319_new_n2228_; 
wire _abc_40319_new_n2229_; 
wire _abc_40319_new_n2230_; 
wire _abc_40319_new_n2231_; 
wire _abc_40319_new_n2232_; 
wire _abc_40319_new_n2233_; 
wire _abc_40319_new_n2234_; 
wire _abc_40319_new_n2235_; 
wire _abc_40319_new_n2236_; 
wire _abc_40319_new_n2237_; 
wire _abc_40319_new_n2238_; 
wire _abc_40319_new_n2239_; 
wire _abc_40319_new_n2240_; 
wire _abc_40319_new_n2241_; 
wire _abc_40319_new_n2242_; 
wire _abc_40319_new_n2243_; 
wire _abc_40319_new_n2244_; 
wire _abc_40319_new_n2245_; 
wire _abc_40319_new_n2246_; 
wire _abc_40319_new_n2247_; 
wire _abc_40319_new_n2248_; 
wire _abc_40319_new_n2249_; 
wire _abc_40319_new_n2250_; 
wire _abc_40319_new_n2251_; 
wire _abc_40319_new_n2252_; 
wire _abc_40319_new_n2253_; 
wire _abc_40319_new_n2254_; 
wire _abc_40319_new_n2255_; 
wire _abc_40319_new_n2256_; 
wire _abc_40319_new_n2257_; 
wire _abc_40319_new_n2258_; 
wire _abc_40319_new_n2259_; 
wire _abc_40319_new_n2260_; 
wire _abc_40319_new_n2261_; 
wire _abc_40319_new_n2262_; 
wire _abc_40319_new_n2263_; 
wire _abc_40319_new_n2264_; 
wire _abc_40319_new_n2265_; 
wire _abc_40319_new_n2266_; 
wire _abc_40319_new_n2267_; 
wire _abc_40319_new_n2268_; 
wire _abc_40319_new_n2269_; 
wire _abc_40319_new_n2270_; 
wire _abc_40319_new_n2271_; 
wire _abc_40319_new_n2272_; 
wire _abc_40319_new_n2273_; 
wire _abc_40319_new_n2274_; 
wire _abc_40319_new_n2275_; 
wire _abc_40319_new_n2276_; 
wire _abc_40319_new_n2277_; 
wire _abc_40319_new_n2278_; 
wire _abc_40319_new_n2279_; 
wire _abc_40319_new_n2280_; 
wire _abc_40319_new_n2281_; 
wire _abc_40319_new_n2282_; 
wire _abc_40319_new_n2283_; 
wire _abc_40319_new_n2284_; 
wire _abc_40319_new_n2285_; 
wire _abc_40319_new_n2286_; 
wire _abc_40319_new_n2287_; 
wire _abc_40319_new_n2288_; 
wire _abc_40319_new_n2289_; 
wire _abc_40319_new_n2290_; 
wire _abc_40319_new_n2291_; 
wire _abc_40319_new_n2292_; 
wire _abc_40319_new_n2293_; 
wire _abc_40319_new_n2294_; 
wire _abc_40319_new_n2295_; 
wire _abc_40319_new_n2296_; 
wire _abc_40319_new_n2297_; 
wire _abc_40319_new_n2298_; 
wire _abc_40319_new_n2299_; 
wire _abc_40319_new_n2300_; 
wire _abc_40319_new_n2301_; 
wire _abc_40319_new_n2302_; 
wire _abc_40319_new_n2303_; 
wire _abc_40319_new_n2304_; 
wire _abc_40319_new_n2305_; 
wire _abc_40319_new_n2306_; 
wire _abc_40319_new_n2307_; 
wire _abc_40319_new_n2308_; 
wire _abc_40319_new_n2309_; 
wire _abc_40319_new_n2310_; 
wire _abc_40319_new_n2311_; 
wire _abc_40319_new_n2312_; 
wire _abc_40319_new_n2313_; 
wire _abc_40319_new_n2314_; 
wire _abc_40319_new_n2315_; 
wire _abc_40319_new_n2316_; 
wire _abc_40319_new_n2317_; 
wire _abc_40319_new_n2318_; 
wire _abc_40319_new_n2319_; 
wire _abc_40319_new_n2320_; 
wire _abc_40319_new_n2321_; 
wire _abc_40319_new_n2322_; 
wire _abc_40319_new_n2323_; 
wire _abc_40319_new_n2324_; 
wire _abc_40319_new_n2325_; 
wire _abc_40319_new_n2326_; 
wire _abc_40319_new_n2327_; 
wire _abc_40319_new_n2328_; 
wire _abc_40319_new_n2329_; 
wire _abc_40319_new_n2330_; 
wire _abc_40319_new_n2331_; 
wire _abc_40319_new_n2332_; 
wire _abc_40319_new_n2333_; 
wire _abc_40319_new_n2334_; 
wire _abc_40319_new_n2335_; 
wire _abc_40319_new_n2336_; 
wire _abc_40319_new_n2337_; 
wire _abc_40319_new_n2338_; 
wire _abc_40319_new_n2339_; 
wire _abc_40319_new_n2340_; 
wire _abc_40319_new_n2341_; 
wire _abc_40319_new_n2342_; 
wire _abc_40319_new_n2343_; 
wire _abc_40319_new_n2344_; 
wire _abc_40319_new_n2345_; 
wire _abc_40319_new_n2346_; 
wire _abc_40319_new_n2347_; 
wire _abc_40319_new_n2348_; 
wire _abc_40319_new_n2349_; 
wire _abc_40319_new_n2350_; 
wire _abc_40319_new_n2351_; 
wire _abc_40319_new_n2352_; 
wire _abc_40319_new_n2353_; 
wire _abc_40319_new_n2354_; 
wire _abc_40319_new_n2355_; 
wire _abc_40319_new_n2356_; 
wire _abc_40319_new_n2357_; 
wire _abc_40319_new_n2358_; 
wire _abc_40319_new_n2359_; 
wire _abc_40319_new_n2360_; 
wire _abc_40319_new_n2361_; 
wire _abc_40319_new_n2362_; 
wire _abc_40319_new_n2363_; 
wire _abc_40319_new_n2364_; 
wire _abc_40319_new_n2365_; 
wire _abc_40319_new_n2366_; 
wire _abc_40319_new_n2367_; 
wire _abc_40319_new_n2368_; 
wire _abc_40319_new_n2369_; 
wire _abc_40319_new_n2370_; 
wire _abc_40319_new_n2371_; 
wire _abc_40319_new_n2372_; 
wire _abc_40319_new_n2373_; 
wire _abc_40319_new_n2374_; 
wire _abc_40319_new_n2375_; 
wire _abc_40319_new_n2376_; 
wire _abc_40319_new_n2377_; 
wire _abc_40319_new_n2378_; 
wire _abc_40319_new_n2379_; 
wire _abc_40319_new_n2380_; 
wire _abc_40319_new_n2381_; 
wire _abc_40319_new_n2382_; 
wire _abc_40319_new_n2383_; 
wire _abc_40319_new_n2384_; 
wire _abc_40319_new_n2385_; 
wire _abc_40319_new_n2386_; 
wire _abc_40319_new_n2387_; 
wire _abc_40319_new_n2388_; 
wire _abc_40319_new_n2389_; 
wire _abc_40319_new_n2390_; 
wire _abc_40319_new_n2391_; 
wire _abc_40319_new_n2392_; 
wire _abc_40319_new_n2393_; 
wire _abc_40319_new_n2394_; 
wire _abc_40319_new_n2395_; 
wire _abc_40319_new_n2396_; 
wire _abc_40319_new_n2397_; 
wire _abc_40319_new_n2398_; 
wire _abc_40319_new_n2399_; 
wire _abc_40319_new_n2400_; 
wire _abc_40319_new_n2401_; 
wire _abc_40319_new_n2402_; 
wire _abc_40319_new_n2403_; 
wire _abc_40319_new_n2404_; 
wire _abc_40319_new_n2405_; 
wire _abc_40319_new_n2406_; 
wire _abc_40319_new_n2407_; 
wire _abc_40319_new_n2408_; 
wire _abc_40319_new_n2409_; 
wire _abc_40319_new_n2410_; 
wire _abc_40319_new_n2411_; 
wire _abc_40319_new_n2412_; 
wire _abc_40319_new_n2413_; 
wire _abc_40319_new_n2414_; 
wire _abc_40319_new_n2415_; 
wire _abc_40319_new_n2416_; 
wire _abc_40319_new_n2417_; 
wire _abc_40319_new_n2418_; 
wire _abc_40319_new_n2419_; 
wire _abc_40319_new_n2420_; 
wire _abc_40319_new_n2421_; 
wire _abc_40319_new_n2422_; 
wire _abc_40319_new_n2423_; 
wire _abc_40319_new_n2424_; 
wire _abc_40319_new_n2425_; 
wire _abc_40319_new_n2426_; 
wire _abc_40319_new_n2427_; 
wire _abc_40319_new_n2428_; 
wire _abc_40319_new_n2429_; 
wire _abc_40319_new_n2430_; 
wire _abc_40319_new_n2431_; 
wire _abc_40319_new_n2432_; 
wire _abc_40319_new_n2433_; 
wire _abc_40319_new_n2434_; 
wire _abc_40319_new_n2435_; 
wire _abc_40319_new_n2436_; 
wire _abc_40319_new_n2437_; 
wire _abc_40319_new_n2438_; 
wire _abc_40319_new_n2439_; 
wire _abc_40319_new_n2440_; 
wire _abc_40319_new_n2441_; 
wire _abc_40319_new_n2442_; 
wire _abc_40319_new_n2443_; 
wire _abc_40319_new_n2444_; 
wire _abc_40319_new_n2445_; 
wire _abc_40319_new_n2446_; 
wire _abc_40319_new_n2447_; 
wire _abc_40319_new_n2448_; 
wire _abc_40319_new_n2449_; 
wire _abc_40319_new_n2450_; 
wire _abc_40319_new_n2451_; 
wire _abc_40319_new_n2452_; 
wire _abc_40319_new_n2453_; 
wire _abc_40319_new_n2454_; 
wire _abc_40319_new_n2455_; 
wire _abc_40319_new_n2456_; 
wire _abc_40319_new_n2457_; 
wire _abc_40319_new_n2458_; 
wire _abc_40319_new_n2459_; 
wire _abc_40319_new_n2460_; 
wire _abc_40319_new_n2461_; 
wire _abc_40319_new_n2462_; 
wire _abc_40319_new_n2463_; 
wire _abc_40319_new_n2464_; 
wire _abc_40319_new_n2465_; 
wire _abc_40319_new_n2466_; 
wire _abc_40319_new_n2467_; 
wire _abc_40319_new_n2468_; 
wire _abc_40319_new_n2469_; 
wire _abc_40319_new_n2470_; 
wire _abc_40319_new_n2471_; 
wire _abc_40319_new_n2472_; 
wire _abc_40319_new_n2473_; 
wire _abc_40319_new_n2474_; 
wire _abc_40319_new_n2475_; 
wire _abc_40319_new_n2476_; 
wire _abc_40319_new_n2477_; 
wire _abc_40319_new_n2478_; 
wire _abc_40319_new_n2479_; 
wire _abc_40319_new_n2480_; 
wire _abc_40319_new_n2481_; 
wire _abc_40319_new_n2482_; 
wire _abc_40319_new_n2483_; 
wire _abc_40319_new_n2484_; 
wire _abc_40319_new_n2485_; 
wire _abc_40319_new_n2486_; 
wire _abc_40319_new_n2487_; 
wire _abc_40319_new_n2488_; 
wire _abc_40319_new_n2489_; 
wire _abc_40319_new_n2490_; 
wire _abc_40319_new_n2491_; 
wire _abc_40319_new_n2492_; 
wire _abc_40319_new_n2493_; 
wire _abc_40319_new_n2494_; 
wire _abc_40319_new_n2495_; 
wire _abc_40319_new_n2496_; 
wire _abc_40319_new_n2497_; 
wire _abc_40319_new_n2498_; 
wire _abc_40319_new_n2499_; 
wire _abc_40319_new_n2500_; 
wire _abc_40319_new_n2501_; 
wire _abc_40319_new_n2502_; 
wire _abc_40319_new_n2503_; 
wire _abc_40319_new_n2504_; 
wire _abc_40319_new_n2505_; 
wire _abc_40319_new_n2506_; 
wire _abc_40319_new_n2507_; 
wire _abc_40319_new_n2508_; 
wire _abc_40319_new_n2509_; 
wire _abc_40319_new_n2510_; 
wire _abc_40319_new_n2511_; 
wire _abc_40319_new_n2512_; 
wire _abc_40319_new_n2513_; 
wire _abc_40319_new_n2514_; 
wire _abc_40319_new_n2515_; 
wire _abc_40319_new_n2516_; 
wire _abc_40319_new_n2517_; 
wire _abc_40319_new_n2518_; 
wire _abc_40319_new_n2519_; 
wire _abc_40319_new_n2520_; 
wire _abc_40319_new_n2521_; 
wire _abc_40319_new_n2522_; 
wire _abc_40319_new_n2523_; 
wire _abc_40319_new_n2524_; 
wire _abc_40319_new_n2525_; 
wire _abc_40319_new_n2526_; 
wire _abc_40319_new_n2527_; 
wire _abc_40319_new_n2528_; 
wire _abc_40319_new_n2529_; 
wire _abc_40319_new_n2531_; 
wire _abc_40319_new_n2532_; 
wire _abc_40319_new_n2533_; 
wire _abc_40319_new_n2534_; 
wire _abc_40319_new_n2535_; 
wire _abc_40319_new_n2536_; 
wire _abc_40319_new_n2537_; 
wire _abc_40319_new_n2538_; 
wire _abc_40319_new_n2539_; 
wire _abc_40319_new_n2540_; 
wire _abc_40319_new_n2542_; 
wire _abc_40319_new_n2543_; 
wire _abc_40319_new_n2544_; 
wire _abc_40319_new_n2545_; 
wire _abc_40319_new_n2546_; 
wire _abc_40319_new_n2547_; 
wire _abc_40319_new_n2548_; 
wire _abc_40319_new_n2549_; 
wire _abc_40319_new_n2550_; 
wire _abc_40319_new_n2551_; 
wire _abc_40319_new_n2552_; 
wire _abc_40319_new_n2553_; 
wire _abc_40319_new_n2554_; 
wire _abc_40319_new_n2555_; 
wire _abc_40319_new_n2556_; 
wire _abc_40319_new_n2557_; 
wire _abc_40319_new_n2559_; 
wire _abc_40319_new_n2560_; 
wire _abc_40319_new_n2561_; 
wire _abc_40319_new_n2562_; 
wire _abc_40319_new_n2563_; 
wire _abc_40319_new_n2564_; 
wire _abc_40319_new_n2565_; 
wire _abc_40319_new_n2566_; 
wire _abc_40319_new_n2567_; 
wire _abc_40319_new_n2568_; 
wire _abc_40319_new_n2569_; 
wire _abc_40319_new_n2570_; 
wire _abc_40319_new_n2571_; 
wire _abc_40319_new_n2572_; 
wire _abc_40319_new_n2573_; 
wire _abc_40319_new_n2574_; 
wire _abc_40319_new_n2575_; 
wire _abc_40319_new_n2577_; 
wire _abc_40319_new_n2578_; 
wire _abc_40319_new_n2579_; 
wire _abc_40319_new_n2580_; 
wire _abc_40319_new_n2581_; 
wire _abc_40319_new_n2582_; 
wire _abc_40319_new_n2583_; 
wire _abc_40319_new_n2584_; 
wire _abc_40319_new_n2585_; 
wire _abc_40319_new_n2586_; 
wire _abc_40319_new_n2587_; 
wire _abc_40319_new_n2588_; 
wire _abc_40319_new_n2589_; 
wire _abc_40319_new_n2590_; 
wire _abc_40319_new_n2591_; 
wire _abc_40319_new_n2593_; 
wire _abc_40319_new_n2594_; 
wire _abc_40319_new_n2595_; 
wire _abc_40319_new_n2596_; 
wire _abc_40319_new_n2597_; 
wire _abc_40319_new_n2598_; 
wire _abc_40319_new_n2599_; 
wire _abc_40319_new_n2600_; 
wire _abc_40319_new_n2601_; 
wire _abc_40319_new_n2602_; 
wire _abc_40319_new_n2603_; 
wire _abc_40319_new_n2604_; 
wire _abc_40319_new_n2605_; 
wire _abc_40319_new_n2607_; 
wire _abc_40319_new_n2608_; 
wire _abc_40319_new_n2609_; 
wire _abc_40319_new_n2610_; 
wire _abc_40319_new_n2611_; 
wire _abc_40319_new_n2612_; 
wire _abc_40319_new_n2613_; 
wire _abc_40319_new_n2614_; 
wire _abc_40319_new_n2615_; 
wire _abc_40319_new_n2616_; 
wire _abc_40319_new_n2617_; 
wire _abc_40319_new_n2618_; 
wire _abc_40319_new_n2619_; 
wire _abc_40319_new_n2620_; 
wire _abc_40319_new_n2621_; 
wire _abc_40319_new_n2623_; 
wire _abc_40319_new_n2624_; 
wire _abc_40319_new_n2625_; 
wire _abc_40319_new_n2626_; 
wire _abc_40319_new_n2627_; 
wire _abc_40319_new_n2628_; 
wire _abc_40319_new_n2629_; 
wire _abc_40319_new_n2630_; 
wire _abc_40319_new_n2631_; 
wire _abc_40319_new_n2632_; 
wire _abc_40319_new_n2633_; 
wire _abc_40319_new_n2634_; 
wire _abc_40319_new_n2635_; 
wire _abc_40319_new_n2636_; 
wire _abc_40319_new_n2637_; 
wire _abc_40319_new_n2639_; 
wire _abc_40319_new_n2640_; 
wire _abc_40319_new_n2641_; 
wire _abc_40319_new_n2642_; 
wire _abc_40319_new_n2643_; 
wire _abc_40319_new_n2644_; 
wire _abc_40319_new_n2645_; 
wire _abc_40319_new_n2646_; 
wire _abc_40319_new_n2647_; 
wire _abc_40319_new_n2648_; 
wire _abc_40319_new_n2649_; 
wire _abc_40319_new_n2650_; 
wire _abc_40319_new_n2651_; 
wire _abc_40319_new_n2652_; 
wire _abc_40319_new_n2653_; 
wire _abc_40319_new_n2654_; 
wire _abc_40319_new_n2655_; 
wire _abc_40319_new_n2656_; 
wire _abc_40319_new_n2657_; 
wire _abc_40319_new_n2658_; 
wire _abc_40319_new_n2659_; 
wire _abc_40319_new_n2660_; 
wire _abc_40319_new_n2661_; 
wire _abc_40319_new_n2663_; 
wire _abc_40319_new_n2664_; 
wire _abc_40319_new_n2665_; 
wire _abc_40319_new_n2666_; 
wire _abc_40319_new_n2667_; 
wire _abc_40319_new_n2668_; 
wire _abc_40319_new_n2669_; 
wire _abc_40319_new_n2670_; 
wire _abc_40319_new_n2671_; 
wire _abc_40319_new_n2672_; 
wire _abc_40319_new_n2673_; 
wire _abc_40319_new_n2674_; 
wire _abc_40319_new_n2675_; 
wire _abc_40319_new_n2676_; 
wire _abc_40319_new_n2677_; 
wire _abc_40319_new_n2678_; 
wire _abc_40319_new_n2679_; 
wire _abc_40319_new_n2680_; 
wire _abc_40319_new_n2681_; 
wire _abc_40319_new_n2682_; 
wire _abc_40319_new_n2683_; 
wire _abc_40319_new_n2684_; 
wire _abc_40319_new_n2685_; 
wire _abc_40319_new_n2686_; 
wire _abc_40319_new_n2687_; 
wire _abc_40319_new_n2688_; 
wire _abc_40319_new_n2689_; 
wire _abc_40319_new_n2690_; 
wire _abc_40319_new_n2691_; 
wire _abc_40319_new_n2692_; 
wire _abc_40319_new_n2694_; 
wire _abc_40319_new_n2695_; 
wire _abc_40319_new_n2696_; 
wire _abc_40319_new_n2697_; 
wire _abc_40319_new_n2698_; 
wire _abc_40319_new_n2699_; 
wire _abc_40319_new_n2700_; 
wire _abc_40319_new_n2701_; 
wire _abc_40319_new_n2702_; 
wire _abc_40319_new_n2703_; 
wire _abc_40319_new_n2704_; 
wire _abc_40319_new_n2705_; 
wire _abc_40319_new_n2706_; 
wire _abc_40319_new_n2707_; 
wire _abc_40319_new_n2708_; 
wire _abc_40319_new_n2709_; 
wire _abc_40319_new_n2710_; 
wire _abc_40319_new_n2711_; 
wire _abc_40319_new_n2712_; 
wire _abc_40319_new_n2713_; 
wire _abc_40319_new_n2715_; 
wire _abc_40319_new_n2716_; 
wire _abc_40319_new_n2717_; 
wire _abc_40319_new_n2718_; 
wire _abc_40319_new_n2719_; 
wire _abc_40319_new_n2720_; 
wire _abc_40319_new_n2721_; 
wire _abc_40319_new_n2722_; 
wire _abc_40319_new_n2723_; 
wire _abc_40319_new_n2724_; 
wire _abc_40319_new_n2725_; 
wire _abc_40319_new_n2726_; 
wire _abc_40319_new_n2727_; 
wire _abc_40319_new_n2728_; 
wire _abc_40319_new_n2729_; 
wire _abc_40319_new_n2730_; 
wire _abc_40319_new_n2731_; 
wire _abc_40319_new_n2732_; 
wire _abc_40319_new_n2733_; 
wire _abc_40319_new_n2734_; 
wire _abc_40319_new_n2735_; 
wire _abc_40319_new_n2736_; 
wire _abc_40319_new_n2738_; 
wire _abc_40319_new_n2739_; 
wire _abc_40319_new_n2740_; 
wire _abc_40319_new_n2741_; 
wire _abc_40319_new_n2742_; 
wire _abc_40319_new_n2743_; 
wire _abc_40319_new_n2744_; 
wire _abc_40319_new_n2745_; 
wire _abc_40319_new_n2746_; 
wire _abc_40319_new_n2747_; 
wire _abc_40319_new_n2748_; 
wire _abc_40319_new_n2749_; 
wire _abc_40319_new_n2750_; 
wire _abc_40319_new_n2751_; 
wire _abc_40319_new_n2752_; 
wire _abc_40319_new_n2753_; 
wire _abc_40319_new_n2754_; 
wire _abc_40319_new_n2755_; 
wire _abc_40319_new_n2756_; 
wire _abc_40319_new_n2757_; 
wire _abc_40319_new_n2758_; 
wire _abc_40319_new_n2759_; 
wire _abc_40319_new_n2761_; 
wire _abc_40319_new_n2762_; 
wire _abc_40319_new_n2763_; 
wire _abc_40319_new_n2764_; 
wire _abc_40319_new_n2765_; 
wire _abc_40319_new_n2766_; 
wire _abc_40319_new_n2767_; 
wire _abc_40319_new_n2768_; 
wire _abc_40319_new_n2769_; 
wire _abc_40319_new_n2770_; 
wire _abc_40319_new_n2771_; 
wire _abc_40319_new_n2772_; 
wire _abc_40319_new_n2773_; 
wire _abc_40319_new_n2774_; 
wire _abc_40319_new_n2775_; 
wire _abc_40319_new_n2776_; 
wire _abc_40319_new_n2777_; 
wire _abc_40319_new_n2778_; 
wire _abc_40319_new_n2779_; 
wire _abc_40319_new_n2780_; 
wire _abc_40319_new_n2781_; 
wire _abc_40319_new_n2783_; 
wire _abc_40319_new_n2784_; 
wire _abc_40319_new_n2785_; 
wire _abc_40319_new_n2786_; 
wire _abc_40319_new_n2787_; 
wire _abc_40319_new_n2788_; 
wire _abc_40319_new_n2789_; 
wire _abc_40319_new_n2790_; 
wire _abc_40319_new_n2791_; 
wire _abc_40319_new_n2792_; 
wire _abc_40319_new_n2793_; 
wire _abc_40319_new_n2794_; 
wire _abc_40319_new_n2795_; 
wire _abc_40319_new_n2796_; 
wire _abc_40319_new_n2797_; 
wire _abc_40319_new_n2798_; 
wire _abc_40319_new_n2799_; 
wire _abc_40319_new_n2800_; 
wire _abc_40319_new_n2801_; 
wire _abc_40319_new_n2803_; 
wire _abc_40319_new_n2804_; 
wire _abc_40319_new_n2805_; 
wire _abc_40319_new_n2806_; 
wire _abc_40319_new_n2807_; 
wire _abc_40319_new_n2808_; 
wire _abc_40319_new_n2809_; 
wire _abc_40319_new_n2810_; 
wire _abc_40319_new_n2811_; 
wire _abc_40319_new_n2812_; 
wire _abc_40319_new_n2813_; 
wire _abc_40319_new_n2814_; 
wire _abc_40319_new_n2815_; 
wire _abc_40319_new_n2816_; 
wire _abc_40319_new_n2817_; 
wire _abc_40319_new_n2818_; 
wire _abc_40319_new_n2819_; 
wire _abc_40319_new_n2820_; 
wire _abc_40319_new_n2821_; 
wire _abc_40319_new_n2822_; 
wire _abc_40319_new_n2823_; 
wire _abc_40319_new_n2824_; 
wire _abc_40319_new_n2825_; 
wire _abc_40319_new_n2826_; 
wire _abc_40319_new_n2828_; 
wire _abc_40319_new_n2829_; 
wire _abc_40319_new_n2830_; 
wire _abc_40319_new_n2831_; 
wire _abc_40319_new_n2832_; 
wire _abc_40319_new_n2833_; 
wire _abc_40319_new_n2834_; 
wire _abc_40319_new_n2835_; 
wire _abc_40319_new_n2836_; 
wire _abc_40319_new_n2837_; 
wire _abc_40319_new_n2838_; 
wire _abc_40319_new_n2839_; 
wire _abc_40319_new_n2840_; 
wire _abc_40319_new_n2841_; 
wire _abc_40319_new_n2842_; 
wire _abc_40319_new_n2843_; 
wire _abc_40319_new_n2844_; 
wire _abc_40319_new_n2845_; 
wire _abc_40319_new_n2846_; 
wire _abc_40319_new_n2847_; 
wire _abc_40319_new_n2848_; 
wire _abc_40319_new_n2849_; 
wire _abc_40319_new_n2850_; 
wire _abc_40319_new_n2851_; 
wire _abc_40319_new_n2853_; 
wire _abc_40319_new_n2854_; 
wire _abc_40319_new_n2855_; 
wire _abc_40319_new_n2856_; 
wire _abc_40319_new_n2857_; 
wire _abc_40319_new_n2858_; 
wire _abc_40319_new_n2859_; 
wire _abc_40319_new_n2860_; 
wire _abc_40319_new_n2861_; 
wire _abc_40319_new_n2862_; 
wire _abc_40319_new_n2863_; 
wire _abc_40319_new_n2864_; 
wire _abc_40319_new_n2865_; 
wire _abc_40319_new_n2866_; 
wire _abc_40319_new_n2867_; 
wire _abc_40319_new_n2868_; 
wire _abc_40319_new_n2869_; 
wire _abc_40319_new_n2870_; 
wire _abc_40319_new_n2871_; 
wire _abc_40319_new_n2872_; 
wire _abc_40319_new_n2873_; 
wire _abc_40319_new_n2874_; 
wire _abc_40319_new_n2875_; 
wire _abc_40319_new_n2876_; 
wire _abc_40319_new_n2878_; 
wire _abc_40319_new_n2879_; 
wire _abc_40319_new_n2880_; 
wire _abc_40319_new_n2881_; 
wire _abc_40319_new_n2882_; 
wire _abc_40319_new_n2883_; 
wire _abc_40319_new_n2884_; 
wire _abc_40319_new_n2885_; 
wire _abc_40319_new_n2886_; 
wire _abc_40319_new_n2887_; 
wire _abc_40319_new_n2888_; 
wire _abc_40319_new_n2889_; 
wire _abc_40319_new_n2890_; 
wire _abc_40319_new_n2891_; 
wire _abc_40319_new_n2892_; 
wire _abc_40319_new_n2893_; 
wire _abc_40319_new_n2894_; 
wire _abc_40319_new_n2895_; 
wire _abc_40319_new_n2896_; 
wire _abc_40319_new_n2897_; 
wire _abc_40319_new_n2899_; 
wire _abc_40319_new_n2900_; 
wire _abc_40319_new_n2901_; 
wire _abc_40319_new_n2902_; 
wire _abc_40319_new_n2903_; 
wire _abc_40319_new_n2904_; 
wire _abc_40319_new_n2905_; 
wire _abc_40319_new_n2906_; 
wire _abc_40319_new_n2907_; 
wire _abc_40319_new_n2908_; 
wire _abc_40319_new_n2909_; 
wire _abc_40319_new_n2910_; 
wire _abc_40319_new_n2911_; 
wire _abc_40319_new_n2912_; 
wire _abc_40319_new_n2913_; 
wire _abc_40319_new_n2914_; 
wire _abc_40319_new_n2915_; 
wire _abc_40319_new_n2916_; 
wire _abc_40319_new_n2917_; 
wire _abc_40319_new_n2918_; 
wire _abc_40319_new_n2919_; 
wire _abc_40319_new_n2920_; 
wire _abc_40319_new_n2921_; 
wire _abc_40319_new_n2922_; 
wire _abc_40319_new_n2923_; 
wire _abc_40319_new_n2924_; 
wire _abc_40319_new_n2925_; 
wire _abc_40319_new_n2926_; 
wire _abc_40319_new_n2927_; 
wire _abc_40319_new_n2928_; 
wire _abc_40319_new_n2930_; 
wire _abc_40319_new_n2931_; 
wire _abc_40319_new_n2932_; 
wire _abc_40319_new_n2933_; 
wire _abc_40319_new_n2934_; 
wire _abc_40319_new_n2935_; 
wire _abc_40319_new_n2936_; 
wire _abc_40319_new_n2937_; 
wire _abc_40319_new_n2938_; 
wire _abc_40319_new_n2939_; 
wire _abc_40319_new_n2940_; 
wire _abc_40319_new_n2941_; 
wire _abc_40319_new_n2942_; 
wire _abc_40319_new_n2943_; 
wire _abc_40319_new_n2944_; 
wire _abc_40319_new_n2945_; 
wire _abc_40319_new_n2946_; 
wire _abc_40319_new_n2947_; 
wire _abc_40319_new_n2948_; 
wire _abc_40319_new_n2949_; 
wire _abc_40319_new_n2950_; 
wire _abc_40319_new_n2951_; 
wire _abc_40319_new_n2952_; 
wire _abc_40319_new_n2953_; 
wire _abc_40319_new_n2955_; 
wire _abc_40319_new_n2956_; 
wire _abc_40319_new_n2957_; 
wire _abc_40319_new_n2958_; 
wire _abc_40319_new_n2959_; 
wire _abc_40319_new_n2960_; 
wire _abc_40319_new_n2961_; 
wire _abc_40319_new_n2962_; 
wire _abc_40319_new_n2963_; 
wire _abc_40319_new_n2964_; 
wire _abc_40319_new_n2965_; 
wire _abc_40319_new_n2966_; 
wire _abc_40319_new_n2967_; 
wire _abc_40319_new_n2968_; 
wire _abc_40319_new_n2969_; 
wire _abc_40319_new_n2970_; 
wire _abc_40319_new_n2971_; 
wire _abc_40319_new_n2972_; 
wire _abc_40319_new_n2973_; 
wire _abc_40319_new_n2974_; 
wire _abc_40319_new_n2975_; 
wire _abc_40319_new_n2976_; 
wire _abc_40319_new_n2977_; 
wire _abc_40319_new_n2978_; 
wire _abc_40319_new_n2979_; 
wire _abc_40319_new_n2980_; 
wire _abc_40319_new_n2981_; 
wire _abc_40319_new_n2982_; 
wire _abc_40319_new_n2983_; 
wire _abc_40319_new_n2984_; 
wire _abc_40319_new_n2985_; 
wire _abc_40319_new_n2986_; 
wire _abc_40319_new_n2987_; 
wire _abc_40319_new_n2988_; 
wire _abc_40319_new_n2989_; 
wire _abc_40319_new_n2990_; 
wire _abc_40319_new_n2991_; 
wire _abc_40319_new_n2992_; 
wire _abc_40319_new_n2993_; 
wire _abc_40319_new_n2994_; 
wire _abc_40319_new_n2996_; 
wire _abc_40319_new_n2997_; 
wire _abc_40319_new_n2998_; 
wire _abc_40319_new_n2999_; 
wire _abc_40319_new_n3000_; 
wire _abc_40319_new_n3001_; 
wire _abc_40319_new_n3003_; 
wire _abc_40319_new_n3004_; 
wire _abc_40319_new_n3005_; 
wire _abc_40319_new_n3006_; 
wire _abc_40319_new_n3007_; 
wire _abc_40319_new_n3008_; 
wire _abc_40319_new_n3009_; 
wire _abc_40319_new_n3010_; 
wire _abc_40319_new_n3011_; 
wire _abc_40319_new_n3012_; 
wire _abc_40319_new_n3013_; 
wire _abc_40319_new_n3014_; 
wire _abc_40319_new_n3015_; 
wire _abc_40319_new_n3016_; 
wire _abc_40319_new_n3017_; 
wire _abc_40319_new_n3018_; 
wire _abc_40319_new_n3019_; 
wire _abc_40319_new_n3020_; 
wire _abc_40319_new_n3021_; 
wire _abc_40319_new_n3022_; 
wire _abc_40319_new_n3023_; 
wire _abc_40319_new_n3024_; 
wire _abc_40319_new_n3025_; 
wire _abc_40319_new_n3026_; 
wire _abc_40319_new_n3027_; 
wire _abc_40319_new_n3028_; 
wire _abc_40319_new_n3029_; 
wire _abc_40319_new_n3030_; 
wire _abc_40319_new_n3031_; 
wire _abc_40319_new_n3032_; 
wire _abc_40319_new_n3033_; 
wire _abc_40319_new_n3034_; 
wire _abc_40319_new_n3035_; 
wire _abc_40319_new_n3036_; 
wire _abc_40319_new_n3037_; 
wire _abc_40319_new_n3038_; 
wire _abc_40319_new_n3039_; 
wire _abc_40319_new_n3040_; 
wire _abc_40319_new_n3041_; 
wire _abc_40319_new_n3042_; 
wire _abc_40319_new_n3043_; 
wire _abc_40319_new_n3044_; 
wire _abc_40319_new_n3045_; 
wire _abc_40319_new_n3046_; 
wire _abc_40319_new_n3047_; 
wire _abc_40319_new_n3048_; 
wire _abc_40319_new_n3049_; 
wire _abc_40319_new_n3050_; 
wire _abc_40319_new_n3051_; 
wire _abc_40319_new_n3052_; 
wire _abc_40319_new_n3053_; 
wire _abc_40319_new_n3054_; 
wire _abc_40319_new_n3055_; 
wire _abc_40319_new_n3056_; 
wire _abc_40319_new_n3057_; 
wire _abc_40319_new_n3058_; 
wire _abc_40319_new_n3059_; 
wire _abc_40319_new_n3060_; 
wire _abc_40319_new_n3061_; 
wire _abc_40319_new_n3062_; 
wire _abc_40319_new_n3063_; 
wire _abc_40319_new_n3064_; 
wire _abc_40319_new_n3065_; 
wire _abc_40319_new_n3066_; 
wire _abc_40319_new_n3067_; 
wire _abc_40319_new_n3068_; 
wire _abc_40319_new_n3069_; 
wire _abc_40319_new_n3070_; 
wire _abc_40319_new_n3071_; 
wire _abc_40319_new_n3072_; 
wire _abc_40319_new_n3073_; 
wire _abc_40319_new_n3074_; 
wire _abc_40319_new_n3075_; 
wire _abc_40319_new_n3076_; 
wire _abc_40319_new_n3077_; 
wire _abc_40319_new_n3078_; 
wire _abc_40319_new_n3079_; 
wire _abc_40319_new_n3080_; 
wire _abc_40319_new_n3081_; 
wire _abc_40319_new_n3082_; 
wire _abc_40319_new_n3083_; 
wire _abc_40319_new_n3084_; 
wire _abc_40319_new_n3085_; 
wire _abc_40319_new_n3086_; 
wire _abc_40319_new_n3087_; 
wire _abc_40319_new_n3088_; 
wire _abc_40319_new_n3089_; 
wire _abc_40319_new_n3090_; 
wire _abc_40319_new_n3091_; 
wire _abc_40319_new_n3092_; 
wire _abc_40319_new_n3093_; 
wire _abc_40319_new_n3094_; 
wire _abc_40319_new_n3095_; 
wire _abc_40319_new_n3096_; 
wire _abc_40319_new_n3097_; 
wire _abc_40319_new_n3098_; 
wire _abc_40319_new_n3099_; 
wire _abc_40319_new_n3100_; 
wire _abc_40319_new_n3101_; 
wire _abc_40319_new_n3102_; 
wire _abc_40319_new_n3103_; 
wire _abc_40319_new_n3104_; 
wire _abc_40319_new_n3105_; 
wire _abc_40319_new_n3106_; 
wire _abc_40319_new_n3107_; 
wire _abc_40319_new_n3108_; 
wire _abc_40319_new_n3109_; 
wire _abc_40319_new_n3110_; 
wire _abc_40319_new_n3111_; 
wire _abc_40319_new_n3112_; 
wire _abc_40319_new_n3113_; 
wire _abc_40319_new_n3114_; 
wire _abc_40319_new_n3115_; 
wire _abc_40319_new_n3116_; 
wire _abc_40319_new_n3117_; 
wire _abc_40319_new_n3119_; 
wire _abc_40319_new_n3120_; 
wire _abc_40319_new_n3121_; 
wire _abc_40319_new_n3122_; 
wire _abc_40319_new_n3123_; 
wire _abc_40319_new_n3124_; 
wire _abc_40319_new_n3125_; 
wire _abc_40319_new_n3126_; 
wire _abc_40319_new_n3127_; 
wire _abc_40319_new_n3128_; 
wire _abc_40319_new_n3129_; 
wire _abc_40319_new_n3130_; 
wire _abc_40319_new_n3131_; 
wire _abc_40319_new_n3132_; 
wire _abc_40319_new_n3133_; 
wire _abc_40319_new_n3134_; 
wire _abc_40319_new_n3135_; 
wire _abc_40319_new_n3136_; 
wire _abc_40319_new_n3137_; 
wire _abc_40319_new_n3138_; 
wire _abc_40319_new_n3139_; 
wire _abc_40319_new_n3140_; 
wire _abc_40319_new_n3141_; 
wire _abc_40319_new_n3142_; 
wire _abc_40319_new_n3144_; 
wire _abc_40319_new_n3145_; 
wire _abc_40319_new_n3146_; 
wire _abc_40319_new_n3147_; 
wire _abc_40319_new_n3148_; 
wire _abc_40319_new_n3149_; 
wire _abc_40319_new_n3150_; 
wire _abc_40319_new_n3151_; 
wire _abc_40319_new_n3152_; 
wire _abc_40319_new_n3153_; 
wire _abc_40319_new_n3154_; 
wire _abc_40319_new_n3155_; 
wire _abc_40319_new_n3156_; 
wire _abc_40319_new_n3157_; 
wire _abc_40319_new_n3158_; 
wire _abc_40319_new_n3159_; 
wire _abc_40319_new_n3160_; 
wire _abc_40319_new_n3161_; 
wire _abc_40319_new_n3162_; 
wire _abc_40319_new_n3163_; 
wire _abc_40319_new_n3164_; 
wire _abc_40319_new_n3165_; 
wire _abc_40319_new_n3166_; 
wire _abc_40319_new_n3167_; 
wire _abc_40319_new_n3168_; 
wire _abc_40319_new_n3169_; 
wire _abc_40319_new_n3170_; 
wire _abc_40319_new_n3171_; 
wire _abc_40319_new_n3172_; 
wire _abc_40319_new_n3174_; 
wire _abc_40319_new_n3175_; 
wire _abc_40319_new_n3176_; 
wire _abc_40319_new_n3177_; 
wire _abc_40319_new_n3178_; 
wire _abc_40319_new_n3179_; 
wire _abc_40319_new_n3180_; 
wire _abc_40319_new_n3181_; 
wire _abc_40319_new_n3182_; 
wire _abc_40319_new_n3183_; 
wire _abc_40319_new_n3184_; 
wire _abc_40319_new_n3185_; 
wire _abc_40319_new_n3186_; 
wire _abc_40319_new_n3187_; 
wire _abc_40319_new_n3188_; 
wire _abc_40319_new_n3189_; 
wire _abc_40319_new_n3190_; 
wire _abc_40319_new_n3191_; 
wire _abc_40319_new_n3192_; 
wire _abc_40319_new_n3193_; 
wire _abc_40319_new_n3194_; 
wire _abc_40319_new_n3195_; 
wire _abc_40319_new_n3196_; 
wire _abc_40319_new_n3197_; 
wire _abc_40319_new_n3198_; 
wire _abc_40319_new_n3199_; 
wire _abc_40319_new_n3200_; 
wire _abc_40319_new_n3201_; 
wire _abc_40319_new_n3203_; 
wire _abc_40319_new_n3204_; 
wire _abc_40319_new_n3205_; 
wire _abc_40319_new_n3206_; 
wire _abc_40319_new_n3207_; 
wire _abc_40319_new_n3208_; 
wire _abc_40319_new_n3209_; 
wire _abc_40319_new_n3210_; 
wire _abc_40319_new_n3211_; 
wire _abc_40319_new_n3212_; 
wire _abc_40319_new_n3213_; 
wire _abc_40319_new_n3214_; 
wire _abc_40319_new_n3215_; 
wire _abc_40319_new_n3216_; 
wire _abc_40319_new_n3217_; 
wire _abc_40319_new_n3218_; 
wire _abc_40319_new_n3219_; 
wire _abc_40319_new_n3220_; 
wire _abc_40319_new_n3221_; 
wire _abc_40319_new_n3223_; 
wire _abc_40319_new_n3224_; 
wire _abc_40319_new_n3225_; 
wire _abc_40319_new_n3226_; 
wire _abc_40319_new_n3227_; 
wire _abc_40319_new_n3228_; 
wire _abc_40319_new_n3229_; 
wire _abc_40319_new_n3230_; 
wire _abc_40319_new_n3231_; 
wire _abc_40319_new_n3232_; 
wire _abc_40319_new_n3233_; 
wire _abc_40319_new_n3234_; 
wire _abc_40319_new_n3235_; 
wire _abc_40319_new_n3236_; 
wire _abc_40319_new_n3237_; 
wire _abc_40319_new_n3238_; 
wire _abc_40319_new_n3239_; 
wire _abc_40319_new_n3240_; 
wire _abc_40319_new_n3241_; 
wire _abc_40319_new_n3242_; 
wire _abc_40319_new_n3243_; 
wire _abc_40319_new_n3244_; 
wire _abc_40319_new_n3246_; 
wire _abc_40319_new_n3247_; 
wire _abc_40319_new_n3248_; 
wire _abc_40319_new_n3249_; 
wire _abc_40319_new_n3250_; 
wire _abc_40319_new_n3251_; 
wire _abc_40319_new_n3252_; 
wire _abc_40319_new_n3253_; 
wire _abc_40319_new_n3254_; 
wire _abc_40319_new_n3255_; 
wire _abc_40319_new_n3256_; 
wire _abc_40319_new_n3257_; 
wire _abc_40319_new_n3258_; 
wire _abc_40319_new_n3259_; 
wire _abc_40319_new_n3260_; 
wire _abc_40319_new_n3261_; 
wire _abc_40319_new_n3262_; 
wire _abc_40319_new_n3263_; 
wire _abc_40319_new_n3265_; 
wire _abc_40319_new_n3266_; 
wire _abc_40319_new_n3267_; 
wire _abc_40319_new_n3268_; 
wire _abc_40319_new_n3269_; 
wire _abc_40319_new_n3270_; 
wire _abc_40319_new_n3271_; 
wire _abc_40319_new_n3272_; 
wire _abc_40319_new_n3273_; 
wire _abc_40319_new_n3274_; 
wire _abc_40319_new_n3275_; 
wire _abc_40319_new_n3276_; 
wire _abc_40319_new_n3277_; 
wire _abc_40319_new_n3278_; 
wire _abc_40319_new_n3279_; 
wire _abc_40319_new_n3280_; 
wire _abc_40319_new_n3281_; 
wire _abc_40319_new_n3282_; 
wire _abc_40319_new_n3283_; 
wire _abc_40319_new_n3284_; 
wire _abc_40319_new_n3286_; 
wire _abc_40319_new_n3287_; 
wire _abc_40319_new_n3288_; 
wire _abc_40319_new_n3289_; 
wire _abc_40319_new_n3290_; 
wire _abc_40319_new_n3291_; 
wire _abc_40319_new_n3292_; 
wire _abc_40319_new_n3293_; 
wire _abc_40319_new_n3294_; 
wire _abc_40319_new_n3295_; 
wire _abc_40319_new_n3296_; 
wire _abc_40319_new_n3297_; 
wire _abc_40319_new_n3298_; 
wire _abc_40319_new_n3299_; 
wire _abc_40319_new_n3300_; 
wire _abc_40319_new_n3301_; 
wire _abc_40319_new_n3302_; 
wire _abc_40319_new_n3303_; 
wire _abc_40319_new_n3304_; 
wire _abc_40319_new_n3305_; 
wire _abc_40319_new_n3306_; 
wire _abc_40319_new_n3308_; 
wire _abc_40319_new_n3309_; 
wire _abc_40319_new_n3310_; 
wire _abc_40319_new_n3311_; 
wire _abc_40319_new_n3312_; 
wire _abc_40319_new_n3313_; 
wire _abc_40319_new_n3314_; 
wire _abc_40319_new_n3315_; 
wire _abc_40319_new_n3316_; 
wire _abc_40319_new_n3317_; 
wire _abc_40319_new_n3318_; 
wire _abc_40319_new_n3319_; 
wire _abc_40319_new_n3320_; 
wire _abc_40319_new_n3321_; 
wire _abc_40319_new_n3322_; 
wire _abc_40319_new_n3324_; 
wire _abc_40319_new_n3325_; 
wire _abc_40319_new_n3326_; 
wire _abc_40319_new_n3327_; 
wire _abc_40319_new_n3328_; 
wire _abc_40319_new_n3329_; 
wire _abc_40319_new_n3330_; 
wire _abc_40319_new_n3331_; 
wire _abc_40319_new_n3332_; 
wire _abc_40319_new_n3333_; 
wire _abc_40319_new_n3334_; 
wire _abc_40319_new_n3335_; 
wire _abc_40319_new_n3336_; 
wire _abc_40319_new_n3337_; 
wire _abc_40319_new_n3338_; 
wire _abc_40319_new_n3339_; 
wire _abc_40319_new_n3340_; 
wire _abc_40319_new_n3341_; 
wire _abc_40319_new_n3343_; 
wire _abc_40319_new_n3344_; 
wire _abc_40319_new_n3345_; 
wire _abc_40319_new_n3346_; 
wire _abc_40319_new_n3347_; 
wire _abc_40319_new_n3348_; 
wire _abc_40319_new_n3349_; 
wire _abc_40319_new_n3350_; 
wire _abc_40319_new_n3351_; 
wire _abc_40319_new_n3352_; 
wire _abc_40319_new_n3353_; 
wire _abc_40319_new_n3354_; 
wire _abc_40319_new_n3355_; 
wire _abc_40319_new_n3356_; 
wire _abc_40319_new_n3357_; 
wire _abc_40319_new_n3358_; 
wire _abc_40319_new_n3359_; 
wire _abc_40319_new_n3360_; 
wire _abc_40319_new_n3361_; 
wire _abc_40319_new_n3362_; 
wire _abc_40319_new_n3363_; 
wire _abc_40319_new_n3364_; 
wire _abc_40319_new_n3365_; 
wire _abc_40319_new_n3366_; 
wire _abc_40319_new_n3367_; 
wire _abc_40319_new_n3368_; 
wire _abc_40319_new_n3369_; 
wire _abc_40319_new_n3370_; 
wire _abc_40319_new_n3371_; 
wire _abc_40319_new_n3372_; 
wire _abc_40319_new_n3373_; 
wire _abc_40319_new_n3374_; 
wire _abc_40319_new_n3376_; 
wire _abc_40319_new_n3377_; 
wire _abc_40319_new_n3378_; 
wire _abc_40319_new_n3379_; 
wire _abc_40319_new_n3380_; 
wire _abc_40319_new_n3381_; 
wire _abc_40319_new_n3382_; 
wire _abc_40319_new_n3383_; 
wire _abc_40319_new_n3384_; 
wire _abc_40319_new_n3385_; 
wire _abc_40319_new_n3386_; 
wire _abc_40319_new_n3387_; 
wire _abc_40319_new_n3388_; 
wire _abc_40319_new_n3389_; 
wire _abc_40319_new_n3390_; 
wire _abc_40319_new_n3391_; 
wire _abc_40319_new_n3392_; 
wire _abc_40319_new_n3394_; 
wire _abc_40319_new_n3395_; 
wire _abc_40319_new_n3396_; 
wire _abc_40319_new_n3397_; 
wire _abc_40319_new_n3398_; 
wire _abc_40319_new_n3399_; 
wire _abc_40319_new_n3400_; 
wire _abc_40319_new_n3401_; 
wire _abc_40319_new_n3402_; 
wire _abc_40319_new_n3403_; 
wire _abc_40319_new_n3404_; 
wire _abc_40319_new_n3405_; 
wire _abc_40319_new_n3406_; 
wire _abc_40319_new_n3408_; 
wire _abc_40319_new_n3409_; 
wire _abc_40319_new_n3410_; 
wire _abc_40319_new_n3411_; 
wire _abc_40319_new_n3412_; 
wire _abc_40319_new_n3413_; 
wire _abc_40319_new_n3414_; 
wire _abc_40319_new_n3415_; 
wire _abc_40319_new_n3416_; 
wire _abc_40319_new_n3417_; 
wire _abc_40319_new_n3418_; 
wire _abc_40319_new_n3419_; 
wire _abc_40319_new_n3420_; 
wire _abc_40319_new_n3421_; 
wire _abc_40319_new_n3422_; 
wire _abc_40319_new_n3423_; 
wire _abc_40319_new_n3424_; 
wire _abc_40319_new_n3425_; 
wire _abc_40319_new_n3427_; 
wire _abc_40319_new_n3428_; 
wire _abc_40319_new_n3429_; 
wire _abc_40319_new_n3430_; 
wire _abc_40319_new_n3431_; 
wire _abc_40319_new_n3432_; 
wire _abc_40319_new_n3433_; 
wire _abc_40319_new_n3434_; 
wire _abc_40319_new_n3435_; 
wire _abc_40319_new_n3436_; 
wire _abc_40319_new_n3437_; 
wire _abc_40319_new_n3438_; 
wire _abc_40319_new_n3439_; 
wire _abc_40319_new_n3440_; 
wire _abc_40319_new_n3441_; 
wire _abc_40319_new_n3442_; 
wire _abc_40319_new_n3443_; 
wire _abc_40319_new_n3444_; 
wire _abc_40319_new_n3446_; 
wire _abc_40319_new_n3447_; 
wire _abc_40319_new_n3448_; 
wire _abc_40319_new_n3449_; 
wire _abc_40319_new_n3450_; 
wire _abc_40319_new_n3451_; 
wire _abc_40319_new_n3452_; 
wire _abc_40319_new_n3453_; 
wire _abc_40319_new_n3454_; 
wire _abc_40319_new_n3455_; 
wire _abc_40319_new_n3456_; 
wire _abc_40319_new_n3457_; 
wire _abc_40319_new_n3459_; 
wire _abc_40319_new_n3460_; 
wire _abc_40319_new_n3461_; 
wire _abc_40319_new_n3462_; 
wire _abc_40319_new_n3463_; 
wire _abc_40319_new_n3464_; 
wire _abc_40319_new_n3465_; 
wire _abc_40319_new_n3466_; 
wire _abc_40319_new_n3467_; 
wire _abc_40319_new_n3468_; 
wire _abc_40319_new_n3469_; 
wire _abc_40319_new_n3470_; 
wire _abc_40319_new_n3471_; 
wire _abc_40319_new_n3472_; 
wire _abc_40319_new_n3473_; 
wire _abc_40319_new_n3474_; 
wire _abc_40319_new_n3476_; 
wire _abc_40319_new_n3477_; 
wire _abc_40319_new_n3478_; 
wire _abc_40319_new_n3479_; 
wire _abc_40319_new_n3480_; 
wire _abc_40319_new_n3481_; 
wire _abc_40319_new_n3482_; 
wire _abc_40319_new_n3483_; 
wire _abc_40319_new_n3484_; 
wire _abc_40319_new_n3485_; 
wire _abc_40319_new_n3486_; 
wire _abc_40319_new_n3487_; 
wire _abc_40319_new_n3488_; 
wire _abc_40319_new_n3489_; 
wire _abc_40319_new_n3490_; 
wire _abc_40319_new_n3491_; 
wire _abc_40319_new_n3492_; 
wire _abc_40319_new_n3493_; 
wire _abc_40319_new_n3494_; 
wire _abc_40319_new_n3496_; 
wire _abc_40319_new_n3497_; 
wire _abc_40319_new_n3498_; 
wire _abc_40319_new_n3499_; 
wire _abc_40319_new_n3500_; 
wire _abc_40319_new_n3501_; 
wire _abc_40319_new_n3502_; 
wire _abc_40319_new_n3503_; 
wire _abc_40319_new_n3504_; 
wire _abc_40319_new_n3505_; 
wire _abc_40319_new_n3506_; 
wire _abc_40319_new_n3507_; 
wire _abc_40319_new_n3508_; 
wire _abc_40319_new_n3509_; 
wire _abc_40319_new_n3510_; 
wire _abc_40319_new_n3512_; 
wire _abc_40319_new_n3513_; 
wire _abc_40319_new_n3514_; 
wire _abc_40319_new_n3515_; 
wire _abc_40319_new_n3516_; 
wire _abc_40319_new_n3517_; 
wire _abc_40319_new_n3518_; 
wire _abc_40319_new_n3519_; 
wire _abc_40319_new_n3520_; 
wire _abc_40319_new_n3521_; 
wire _abc_40319_new_n3522_; 
wire _abc_40319_new_n3523_; 
wire _abc_40319_new_n3524_; 
wire _abc_40319_new_n3525_; 
wire _abc_40319_new_n3526_; 
wire _abc_40319_new_n3528_; 
wire _abc_40319_new_n3529_; 
wire _abc_40319_new_n3530_; 
wire _abc_40319_new_n3531_; 
wire _abc_40319_new_n3532_; 
wire _abc_40319_new_n3533_; 
wire _abc_40319_new_n3534_; 
wire _abc_40319_new_n3535_; 
wire _abc_40319_new_n3536_; 
wire _abc_40319_new_n3537_; 
wire _abc_40319_new_n3538_; 
wire _abc_40319_new_n3539_; 
wire _abc_40319_new_n3540_; 
wire _abc_40319_new_n3541_; 
wire _abc_40319_new_n3542_; 
wire _abc_40319_new_n3543_; 
wire _abc_40319_new_n3544_; 
wire _abc_40319_new_n3546_; 
wire _abc_40319_new_n3547_; 
wire _abc_40319_new_n3548_; 
wire _abc_40319_new_n3549_; 
wire _abc_40319_new_n3550_; 
wire _abc_40319_new_n3551_; 
wire _abc_40319_new_n3552_; 
wire _abc_40319_new_n3553_; 
wire _abc_40319_new_n3554_; 
wire _abc_40319_new_n3555_; 
wire _abc_40319_new_n3556_; 
wire _abc_40319_new_n3557_; 
wire _abc_40319_new_n3558_; 
wire _abc_40319_new_n3559_; 
wire _abc_40319_new_n3560_; 
wire _abc_40319_new_n3561_; 
wire _abc_40319_new_n3563_; 
wire _abc_40319_new_n3564_; 
wire _abc_40319_new_n3565_; 
wire _abc_40319_new_n3566_; 
wire _abc_40319_new_n3567_; 
wire _abc_40319_new_n3568_; 
wire _abc_40319_new_n3569_; 
wire _abc_40319_new_n3570_; 
wire _abc_40319_new_n3571_; 
wire _abc_40319_new_n3572_; 
wire _abc_40319_new_n3573_; 
wire _abc_40319_new_n3574_; 
wire _abc_40319_new_n3575_; 
wire _abc_40319_new_n3576_; 
wire _abc_40319_new_n3577_; 
wire _abc_40319_new_n3578_; 
wire _abc_40319_new_n3580_; 
wire _abc_40319_new_n3581_; 
wire _abc_40319_new_n3582_; 
wire _abc_40319_new_n3583_; 
wire _abc_40319_new_n3584_; 
wire _abc_40319_new_n3585_; 
wire _abc_40319_new_n3586_; 
wire _abc_40319_new_n3587_; 
wire _abc_40319_new_n3588_; 
wire _abc_40319_new_n3589_; 
wire _abc_40319_new_n3590_; 
wire _abc_40319_new_n3591_; 
wire _abc_40319_new_n3592_; 
wire _abc_40319_new_n3593_; 
wire _abc_40319_new_n3594_; 
wire _abc_40319_new_n3596_; 
wire _abc_40319_new_n3597_; 
wire _abc_40319_new_n3598_; 
wire _abc_40319_new_n3599_; 
wire _abc_40319_new_n3600_; 
wire _abc_40319_new_n3601_; 
wire _abc_40319_new_n3602_; 
wire _abc_40319_new_n3603_; 
wire _abc_40319_new_n3604_; 
wire _abc_40319_new_n3605_; 
wire _abc_40319_new_n3606_; 
wire _abc_40319_new_n3607_; 
wire _abc_40319_new_n3608_; 
wire _abc_40319_new_n3609_; 
wire _abc_40319_new_n3610_; 
wire _abc_40319_new_n3612_; 
wire _abc_40319_new_n3613_; 
wire _abc_40319_new_n3614_; 
wire _abc_40319_new_n3615_; 
wire _abc_40319_new_n3616_; 
wire _abc_40319_new_n3617_; 
wire _abc_40319_new_n3618_; 
wire _abc_40319_new_n3619_; 
wire _abc_40319_new_n3620_; 
wire _abc_40319_new_n3621_; 
wire _abc_40319_new_n3622_; 
wire _abc_40319_new_n3623_; 
wire _abc_40319_new_n3624_; 
wire _abc_40319_new_n3625_; 
wire _abc_40319_new_n3626_; 
wire _abc_40319_new_n3627_; 
wire _abc_40319_new_n3629_; 
wire _abc_40319_new_n3630_; 
wire _abc_40319_new_n3631_; 
wire _abc_40319_new_n3632_; 
wire _abc_40319_new_n3633_; 
wire _abc_40319_new_n3634_; 
wire _abc_40319_new_n3635_; 
wire _abc_40319_new_n3636_; 
wire _abc_40319_new_n3637_; 
wire _abc_40319_new_n3638_; 
wire _abc_40319_new_n3639_; 
wire _abc_40319_new_n3640_; 
wire _abc_40319_new_n3641_; 
wire _abc_40319_new_n3642_; 
wire _abc_40319_new_n3643_; 
wire _abc_40319_new_n3645_; 
wire _abc_40319_new_n3646_; 
wire _abc_40319_new_n3647_; 
wire _abc_40319_new_n3648_; 
wire _abc_40319_new_n3649_; 
wire _abc_40319_new_n3650_; 
wire _abc_40319_new_n3651_; 
wire _abc_40319_new_n3653_; 
wire _abc_40319_new_n3654_; 
wire _abc_40319_new_n3655_; 
wire _abc_40319_new_n3657_; 
wire _abc_40319_new_n3658_; 
wire _abc_40319_new_n3659_; 
wire _abc_40319_new_n3661_; 
wire _abc_40319_new_n3663_; 
wire _abc_40319_new_n3665_; 
wire _abc_40319_new_n3667_; 
wire _abc_40319_new_n3669_; 
wire _abc_40319_new_n3671_; 
wire _abc_40319_new_n3673_; 
wire _abc_40319_new_n3675_; 
wire _abc_40319_new_n3677_; 
wire _abc_40319_new_n3679_; 
wire _abc_40319_new_n3681_; 
wire _abc_40319_new_n3683_; 
wire _abc_40319_new_n3685_; 
wire _abc_40319_new_n3687_; 
wire _abc_40319_new_n3689_; 
wire _abc_40319_new_n3691_; 
wire _abc_40319_new_n3693_; 
wire _abc_40319_new_n3695_; 
wire _abc_40319_new_n3697_; 
wire _abc_40319_new_n3699_; 
wire _abc_40319_new_n3701_; 
wire _abc_40319_new_n3703_; 
wire _abc_40319_new_n3705_; 
wire _abc_40319_new_n3707_; 
wire _abc_40319_new_n3709_; 
wire _abc_40319_new_n3711_; 
wire _abc_40319_new_n3713_; 
wire _abc_40319_new_n3715_; 
wire _abc_40319_new_n3717_; 
wire _abc_40319_new_n3719_; 
wire _abc_40319_new_n3720_; 
wire _abc_40319_new_n3721_; 
wire _abc_40319_new_n3723_; 
wire _abc_40319_new_n3724_; 
wire _abc_40319_new_n3726_; 
wire _abc_40319_new_n3727_; 
wire _abc_40319_new_n3728_; 
wire _abc_40319_new_n3729_; 
wire _abc_40319_new_n3731_; 
wire _abc_40319_new_n3732_; 
wire _abc_40319_new_n3734_; 
wire _abc_40319_new_n3735_; 
wire _abc_40319_new_n3736_; 
wire _abc_40319_new_n3738_; 
wire _abc_40319_new_n3739_; 
wire _abc_40319_new_n3740_; 
wire _abc_40319_new_n3742_; 
wire _abc_40319_new_n3743_; 
wire _abc_40319_new_n3744_; 
wire _abc_40319_new_n3745_; 
wire _abc_40319_new_n3747_; 
wire _abc_40319_new_n3749_; 
wire _abc_40319_new_n3750_; 
wire _abc_40319_new_n3751_; 
wire _abc_40319_new_n3753_; 
wire _abc_40319_new_n3754_; 
wire _abc_40319_new_n3756_; 
wire _abc_40319_new_n3757_; 
wire _abc_40319_new_n3758_; 
wire _abc_40319_new_n3760_; 
wire _abc_40319_new_n3761_; 
wire _abc_40319_new_n3763_; 
wire _abc_40319_new_n3764_; 
wire _abc_40319_new_n3766_; 
wire _abc_40319_new_n3767_; 
wire _abc_40319_new_n3769_; 
wire _abc_40319_new_n3770_; 
wire _abc_40319_new_n3771_; 
wire _abc_40319_new_n3773_; 
wire _abc_40319_new_n3774_; 
wire _abc_40319_new_n3776_; 
wire _abc_40319_new_n3777_; 
wire _abc_40319_new_n3779_; 
wire _abc_40319_new_n3780_; 
wire _abc_40319_new_n3782_; 
wire _abc_40319_new_n3783_; 
wire _abc_40319_new_n3784_; 
wire _abc_40319_new_n3785_; 
wire _abc_40319_new_n3787_; 
wire _abc_40319_new_n3788_; 
wire _abc_40319_new_n3790_; 
wire _abc_40319_new_n3791_; 
wire _abc_40319_new_n3793_; 
wire _abc_40319_new_n3794_; 
wire _abc_40319_new_n3796_; 
wire _abc_40319_new_n3797_; 
wire _abc_40319_new_n3799_; 
wire _abc_40319_new_n3800_; 
wire _abc_40319_new_n3802_; 
wire _abc_40319_new_n3803_; 
wire _abc_40319_new_n3805_; 
wire _abc_40319_new_n3806_; 
wire _abc_40319_new_n3808_; 
wire _abc_40319_new_n3809_; 
wire _abc_40319_new_n3811_; 
wire _abc_40319_new_n3812_; 
wire _abc_40319_new_n3813_; 
wire _abc_40319_new_n3815_; 
wire _abc_40319_new_n3816_; 
wire _abc_40319_new_n3817_; 
wire _abc_40319_new_n3819_; 
wire _abc_40319_new_n3821_; 
wire _abc_40319_new_n3823_; 
wire _abc_40319_new_n3824_; 
wire _abc_40319_new_n3825_; 
wire _abc_40319_new_n3826_; 
wire _abc_40319_new_n3827_; 
wire _abc_40319_new_n3828_; 
wire _abc_40319_new_n3829_; 
wire _abc_40319_new_n3830_; 
wire _abc_40319_new_n3831_; 
wire _abc_40319_new_n3832_; 
wire _abc_40319_new_n3833_; 
wire _abc_40319_new_n3834_; 
wire _abc_40319_new_n3835_; 
wire _abc_40319_new_n3836_; 
wire _abc_40319_new_n3837_; 
wire _abc_40319_new_n3838_; 
wire _abc_40319_new_n3839_; 
wire _abc_40319_new_n3840_; 
wire _abc_40319_new_n3841_; 
wire _abc_40319_new_n3842_; 
wire _abc_40319_new_n3843_; 
wire _abc_40319_new_n3844_; 
wire _abc_40319_new_n3845_; 
wire _abc_40319_new_n3846_; 
wire _abc_40319_new_n3847_; 
wire _abc_40319_new_n3848_; 
wire _abc_40319_new_n3849_; 
wire _abc_40319_new_n3850_; 
wire _abc_40319_new_n3851_; 
wire _abc_40319_new_n3852_; 
wire _abc_40319_new_n3853_; 
wire _abc_40319_new_n3854_; 
wire _abc_40319_new_n3855_; 
wire _abc_40319_new_n3856_; 
wire _abc_40319_new_n3857_; 
wire _abc_40319_new_n3858_; 
wire _abc_40319_new_n3859_; 
wire _abc_40319_new_n3860_; 
wire _abc_40319_new_n3861_; 
wire _abc_40319_new_n3862_; 
wire _abc_40319_new_n3863_; 
wire _abc_40319_new_n3864_; 
wire _abc_40319_new_n3865_; 
wire _abc_40319_new_n3866_; 
wire _abc_40319_new_n3867_; 
wire _abc_40319_new_n3868_; 
wire _abc_40319_new_n3869_; 
wire _abc_40319_new_n3870_; 
wire _abc_40319_new_n3871_; 
wire _abc_40319_new_n3872_; 
wire _abc_40319_new_n3873_; 
wire _abc_40319_new_n3874_; 
wire _abc_40319_new_n3875_; 
wire _abc_40319_new_n3877_; 
wire _abc_40319_new_n3878_; 
wire _abc_40319_new_n3879_; 
wire _abc_40319_new_n3880_; 
wire _abc_40319_new_n3882_; 
wire _abc_40319_new_n3883_; 
wire _abc_40319_new_n3885_; 
wire _abc_40319_new_n3886_; 
wire _abc_40319_new_n3887_; 
wire _abc_40319_new_n3888_; 
wire _abc_40319_new_n3889_; 
wire _abc_40319_new_n3890_; 
wire _abc_40319_new_n3891_; 
wire _abc_40319_new_n3892_; 
wire _abc_40319_new_n3893_; 
wire _abc_40319_new_n3894_; 
wire _abc_40319_new_n3895_; 
wire _abc_40319_new_n3896_; 
wire _abc_40319_new_n3897_; 
wire _abc_40319_new_n3898_; 
wire _abc_40319_new_n3900_; 
wire _abc_40319_new_n3901_; 
wire _abc_40319_new_n3902_; 
wire _abc_40319_new_n3903_; 
wire _abc_40319_new_n3905_; 
wire _abc_40319_new_n3906_; 
wire _abc_40319_new_n3907_; 
wire _abc_40319_new_n3908_; 
wire _abc_40319_new_n3910_; 
wire _abc_40319_new_n3911_; 
wire _abc_40319_new_n3912_; 
wire _abc_40319_new_n3914_; 
wire _abc_40319_new_n3915_; 
wire _abc_40319_new_n3916_; 
wire _abc_40319_new_n3917_; 
wire _abc_40319_new_n3918_; 
wire _abc_40319_new_n3920_; 
wire _abc_40319_new_n3921_; 
wire _abc_40319_new_n3922_; 
wire _abc_40319_new_n3923_; 
wire _abc_40319_new_n3925_; 
wire _abc_40319_new_n3926_; 
wire _abc_40319_new_n3927_; 
wire _abc_40319_new_n3928_; 
wire _abc_40319_new_n3929_; 
wire _abc_40319_new_n3931_; 
wire _abc_40319_new_n3932_; 
wire _abc_40319_new_n3933_; 
wire _abc_40319_new_n3934_; 
wire _abc_40319_new_n3936_; 
wire _abc_40319_new_n3937_; 
wire _abc_40319_new_n3938_; 
wire _abc_40319_new_n3939_; 
wire _abc_40319_new_n3940_; 
wire _abc_40319_new_n3941_; 
wire _abc_40319_new_n3943_; 
wire _abc_40319_new_n3944_; 
wire _abc_40319_new_n3945_; 
wire _abc_40319_new_n3946_; 
wire _abc_40319_new_n3947_; 
wire _abc_40319_new_n3949_; 
wire _abc_40319_new_n3950_; 
wire _abc_40319_new_n3951_; 
wire _abc_40319_new_n3952_; 
wire _abc_40319_new_n3953_; 
wire _abc_40319_new_n3955_; 
wire _abc_40319_new_n3956_; 
wire _abc_40319_new_n3957_; 
wire _abc_40319_new_n3958_; 
wire _abc_40319_new_n3960_; 
wire _abc_40319_new_n3961_; 
wire _abc_40319_new_n3962_; 
wire _abc_40319_new_n3963_; 
wire _abc_40319_new_n3964_; 
wire _abc_40319_new_n3965_; 
wire _abc_40319_new_n3967_; 
wire _abc_40319_new_n3968_; 
wire _abc_40319_new_n3969_; 
wire _abc_40319_new_n3970_; 
wire _abc_40319_new_n3972_; 
wire _abc_40319_new_n3973_; 
wire _abc_40319_new_n3974_; 
wire _abc_40319_new_n3975_; 
wire _abc_40319_new_n3977_; 
wire _abc_40319_new_n3978_; 
wire _abc_40319_new_n3979_; 
wire _abc_40319_new_n3980_; 
wire _abc_40319_new_n3982_; 
wire _abc_40319_new_n3983_; 
wire _abc_40319_new_n3984_; 
wire _abc_40319_new_n3985_; 
wire _abc_40319_new_n3986_; 
wire _abc_40319_new_n3988_; 
wire _abc_40319_new_n3989_; 
wire _abc_40319_new_n3990_; 
wire _abc_40319_new_n3991_; 
wire _abc_40319_new_n3992_; 
wire _abc_40319_new_n3994_; 
wire _abc_40319_new_n3995_; 
wire _abc_40319_new_n3996_; 
wire _abc_40319_new_n3997_; 
wire _abc_40319_new_n3998_; 
wire _abc_40319_new_n3999_; 
wire _abc_40319_new_n4001_; 
wire _abc_40319_new_n4002_; 
wire _abc_40319_new_n4003_; 
wire _abc_40319_new_n4004_; 
wire _abc_40319_new_n4005_; 
wire _abc_40319_new_n4007_; 
wire _abc_40319_new_n4008_; 
wire _abc_40319_new_n4009_; 
wire _abc_40319_new_n4010_; 
wire _abc_40319_new_n4011_; 
wire _abc_40319_new_n4013_; 
wire _abc_40319_new_n4014_; 
wire _abc_40319_new_n4015_; 
wire _abc_40319_new_n4016_; 
wire _abc_40319_new_n4017_; 
wire _abc_40319_new_n4018_; 
wire _abc_40319_new_n4020_; 
wire _abc_40319_new_n4021_; 
wire _abc_40319_new_n4022_; 
wire _abc_40319_new_n4023_; 
wire _abc_40319_new_n4024_; 
wire _abc_40319_new_n4025_; 
wire _abc_40319_new_n4026_; 
wire _abc_40319_new_n4028_; 
wire _abc_40319_new_n4029_; 
wire _abc_40319_new_n4030_; 
wire _abc_40319_new_n4031_; 
wire _abc_40319_new_n4032_; 
wire _abc_40319_new_n4034_; 
wire _abc_40319_new_n4035_; 
wire _abc_40319_new_n4036_; 
wire _abc_40319_new_n4037_; 
wire _abc_40319_new_n4038_; 
wire _abc_40319_new_n4040_; 
wire _abc_40319_new_n4041_; 
wire _abc_40319_new_n4042_; 
wire _abc_40319_new_n4043_; 
wire _abc_40319_new_n4044_; 
wire _abc_40319_new_n4046_; 
wire _abc_40319_new_n4047_; 
wire _abc_40319_new_n4048_; 
wire _abc_40319_new_n4049_; 
wire _abc_40319_new_n4050_; 
wire _abc_40319_new_n4052_; 
wire _abc_40319_new_n4053_; 
wire _abc_40319_new_n4054_; 
wire _abc_40319_new_n4055_; 
wire _abc_40319_new_n4056_; 
wire _abc_40319_new_n4057_; 
wire _abc_40319_new_n4058_; 
wire _abc_40319_new_n4059_; 
wire _abc_40319_new_n4061_; 
wire _abc_40319_new_n4062_; 
wire _abc_40319_new_n4063_; 
wire _abc_40319_new_n4064_; 
wire _abc_40319_new_n4065_; 
wire _abc_40319_new_n4066_; 
wire _abc_40319_new_n4068_; 
wire _abc_40319_new_n4069_; 
wire _abc_40319_new_n4070_; 
wire _abc_40319_new_n4071_; 
wire _abc_40319_new_n4072_; 
wire _abc_40319_new_n4073_; 
wire _abc_40319_new_n4075_; 
wire _abc_40319_new_n4076_; 
wire _abc_40319_new_n4077_; 
wire _abc_40319_new_n4079_; 
wire _abc_40319_new_n4080_; 
wire _abc_40319_new_n4081_; 
wire _abc_40319_new_n4082_; 
wire _abc_40319_new_n4084_; 
wire _abc_40319_new_n4085_; 
wire _abc_40319_new_n4086_; 
wire _abc_40319_new_n4087_; 
wire _abc_40319_new_n4089_; 
wire _abc_40319_new_n4091_; 
wire _abc_40319_new_n4092_; 
wire _abc_40319_new_n4094_; 
wire _abc_40319_new_n4096_; 
wire _abc_40319_new_n4098_; 
wire _abc_40319_new_n4100_; 
wire _abc_40319_new_n4102_; 
wire _abc_40319_new_n4104_; 
wire _abc_40319_new_n4106_; 
wire _abc_40319_new_n4108_; 
wire _abc_40319_new_n4110_; 
wire _abc_40319_new_n4112_; 
wire _abc_40319_new_n4114_; 
wire _abc_40319_new_n4116_; 
wire _abc_40319_new_n4118_; 
wire _abc_40319_new_n4119_; 
wire _abc_40319_new_n4121_; 
wire _abc_40319_new_n4122_; 
wire _abc_40319_new_n4124_; 
wire _abc_40319_new_n4126_; 
wire _abc_40319_new_n4128_; 
wire _abc_40319_new_n4129_; 
wire _abc_40319_new_n4131_; 
wire _abc_40319_new_n4133_; 
wire _abc_40319_new_n4134_; 
wire _abc_40319_new_n4136_; 
wire _abc_40319_new_n4138_; 
wire _abc_40319_new_n4140_; 
wire _abc_40319_new_n4142_; 
wire _abc_40319_new_n4144_; 
wire _abc_40319_new_n4146_; 
wire _abc_40319_new_n4148_; 
wire _abc_40319_new_n4150_; 
wire _abc_40319_new_n4151_; 
wire _abc_40319_new_n4153_; 
wire _abc_40319_new_n4155_; 
wire _abc_40319_new_n4156_; 
wire _abc_40319_new_n4158_; 
wire _abc_40319_new_n4159_; 
wire _abc_40319_new_n4161_; 
wire _abc_40319_new_n4163_; 
wire _abc_40319_new_n4165_; 
wire _abc_40319_new_n4167_; 
wire _abc_40319_new_n4169_; 
wire _abc_40319_new_n4171_; 
wire _abc_40319_new_n4173_; 
wire _abc_40319_new_n4175_; 
wire _abc_40319_new_n4177_; 
wire _abc_40319_new_n4179_; 
wire _abc_40319_new_n4181_; 
wire _abc_40319_new_n4183_; 
wire _abc_40319_new_n4185_; 
wire _abc_40319_new_n4187_; 
wire _abc_40319_new_n4189_; 
wire _abc_40319_new_n4191_; 
wire _abc_40319_new_n4193_; 
wire _abc_40319_new_n4195_; 
wire _abc_40319_new_n4197_; 
wire _abc_40319_new_n4199_; 
wire _abc_40319_new_n4201_; 
wire _abc_40319_new_n4203_; 
wire _abc_40319_new_n4205_; 
wire _abc_40319_new_n4207_; 
wire _abc_40319_new_n4209_; 
wire _abc_40319_new_n4211_; 
wire _abc_40319_new_n4213_; 
wire _abc_40319_new_n4215_; 
wire _abc_40319_new_n4217_; 
wire _abc_40319_new_n4219_; 
wire _abc_40319_new_n4221_; 
wire _abc_40319_new_n523_; 
wire _abc_40319_new_n524_; 
wire _abc_40319_new_n525_; 
wire _abc_40319_new_n526_; 
wire _abc_40319_new_n527_; 
wire _abc_40319_new_n528_; 
wire _abc_40319_new_n529_; 
wire _abc_40319_new_n530_; 
wire _abc_40319_new_n531_; 
wire _abc_40319_new_n532_; 
wire _abc_40319_new_n533_; 
wire _abc_40319_new_n534_; 
wire _abc_40319_new_n535_; 
wire _abc_40319_new_n536_; 
wire _abc_40319_new_n537_; 
wire _abc_40319_new_n538_; 
wire _abc_40319_new_n539_; 
wire _abc_40319_new_n540_; 
wire _abc_40319_new_n541_; 
wire _abc_40319_new_n542_; 
wire _abc_40319_new_n543_; 
wire _abc_40319_new_n544_; 
wire _abc_40319_new_n545_; 
wire _abc_40319_new_n546_; 
wire _abc_40319_new_n547_; 
wire _abc_40319_new_n548_; 
wire _abc_40319_new_n549_; 
wire _abc_40319_new_n550_; 
wire _abc_40319_new_n551_; 
wire _abc_40319_new_n552_; 
wire _abc_40319_new_n553_; 
wire _abc_40319_new_n554_; 
wire _abc_40319_new_n555_; 
wire _abc_40319_new_n556_; 
wire _abc_40319_new_n557_; 
wire _abc_40319_new_n558_; 
wire _abc_40319_new_n559_; 
wire _abc_40319_new_n560_; 
wire _abc_40319_new_n561_; 
wire _abc_40319_new_n562_; 
wire _abc_40319_new_n563_; 
wire _abc_40319_new_n564_; 
wire _abc_40319_new_n565_; 
wire _abc_40319_new_n566_; 
wire _abc_40319_new_n567_; 
wire _abc_40319_new_n568_; 
wire _abc_40319_new_n569_; 
wire _abc_40319_new_n570_; 
wire _abc_40319_new_n571_; 
wire _abc_40319_new_n572_; 
wire _abc_40319_new_n573_; 
wire _abc_40319_new_n574_; 
wire _abc_40319_new_n575_; 
wire _abc_40319_new_n576_; 
wire _abc_40319_new_n577_; 
wire _abc_40319_new_n578_; 
wire _abc_40319_new_n579_; 
wire _abc_40319_new_n580_; 
wire _abc_40319_new_n581_; 
wire _abc_40319_new_n582_; 
wire _abc_40319_new_n583_; 
wire _abc_40319_new_n586_; 
wire _abc_40319_new_n587_; 
wire _abc_40319_new_n588_; 
wire _abc_40319_new_n589_; 
wire _abc_40319_new_n590_; 
wire _abc_40319_new_n591_; 
wire _abc_40319_new_n592_; 
wire _abc_40319_new_n593_; 
wire _abc_40319_new_n594_; 
wire _abc_40319_new_n595_; 
wire _abc_40319_new_n596_; 
wire _abc_40319_new_n597_; 
wire _abc_40319_new_n598_; 
wire _abc_40319_new_n599_; 
wire _abc_40319_new_n600_; 
wire _abc_40319_new_n601_; 
wire _abc_40319_new_n602_; 
wire _abc_40319_new_n603_; 
wire _abc_40319_new_n604_; 
wire _abc_40319_new_n605_; 
wire _abc_40319_new_n606_; 
wire _abc_40319_new_n607_; 
wire _abc_40319_new_n608_; 
wire _abc_40319_new_n609_; 
wire _abc_40319_new_n610_; 
wire _abc_40319_new_n611_; 
wire _abc_40319_new_n612_; 
wire _abc_40319_new_n613_; 
wire _abc_40319_new_n614_; 
wire _abc_40319_new_n615_; 
wire _abc_40319_new_n616_; 
wire _abc_40319_new_n617_; 
wire _abc_40319_new_n618_; 
wire _abc_40319_new_n619_; 
wire _abc_40319_new_n620_; 
wire _abc_40319_new_n622_; 
wire _abc_40319_new_n623_; 
wire _abc_40319_new_n624_; 
wire _abc_40319_new_n625_; 
wire _abc_40319_new_n626_; 
wire _abc_40319_new_n627_; 
wire _abc_40319_new_n628_; 
wire _abc_40319_new_n629_; 
wire _abc_40319_new_n630_; 
wire _abc_40319_new_n631_; 
wire _abc_40319_new_n632_; 
wire _abc_40319_new_n633_; 
wire _abc_40319_new_n634_; 
wire _abc_40319_new_n635_; 
wire _abc_40319_new_n636_; 
wire _abc_40319_new_n637_; 
wire _abc_40319_new_n638_; 
wire _abc_40319_new_n639_; 
wire _abc_40319_new_n640_; 
wire _abc_40319_new_n641_; 
wire _abc_40319_new_n642_; 
wire _abc_40319_new_n643_; 
wire _abc_40319_new_n644_; 
wire _abc_40319_new_n645_; 
wire _abc_40319_new_n646_; 
wire _abc_40319_new_n647_; 
wire _abc_40319_new_n648_; 
wire _abc_40319_new_n649_; 
wire _abc_40319_new_n650_; 
wire _abc_40319_new_n651_; 
wire _abc_40319_new_n652_; 
wire _abc_40319_new_n653_; 
wire _abc_40319_new_n654_; 
wire _abc_40319_new_n655_; 
wire _abc_40319_new_n656_; 
wire _abc_40319_new_n657_; 
wire _abc_40319_new_n658_; 
wire _abc_40319_new_n659_; 
wire _abc_40319_new_n660_; 
wire _abc_40319_new_n661_; 
wire _abc_40319_new_n662_; 
wire _abc_40319_new_n663_; 
wire _abc_40319_new_n664_; 
wire _abc_40319_new_n665_; 
wire _abc_40319_new_n666_; 
wire _abc_40319_new_n667_; 
wire _abc_40319_new_n668_; 
wire _abc_40319_new_n669_; 
wire _abc_40319_new_n670_; 
wire _abc_40319_new_n671_; 
wire _abc_40319_new_n672_; 
wire _abc_40319_new_n673_; 
wire _abc_40319_new_n674_; 
wire _abc_40319_new_n675_; 
wire _abc_40319_new_n676_; 
wire _abc_40319_new_n677_; 
wire _abc_40319_new_n678_; 
wire _abc_40319_new_n679_; 
wire _abc_40319_new_n680_; 
wire _abc_40319_new_n681_; 
wire _abc_40319_new_n682_; 
wire _abc_40319_new_n683_; 
wire _abc_40319_new_n684_; 
wire _abc_40319_new_n685_; 
wire _abc_40319_new_n686_; 
wire _abc_40319_new_n687_; 
wire _abc_40319_new_n688_; 
wire _abc_40319_new_n689_; 
wire _abc_40319_new_n690_; 
wire _abc_40319_new_n691_; 
wire _abc_40319_new_n692_; 
wire _abc_40319_new_n693_; 
wire _abc_40319_new_n694_; 
wire _abc_40319_new_n695_; 
wire _abc_40319_new_n696_; 
wire _abc_40319_new_n697_; 
wire _abc_40319_new_n698_; 
wire _abc_40319_new_n699_; 
wire _abc_40319_new_n700_; 
wire _abc_40319_new_n701_; 
wire _abc_40319_new_n702_; 
wire _abc_40319_new_n703_; 
wire _abc_40319_new_n704_; 
wire _abc_40319_new_n705_; 
wire _abc_40319_new_n706_; 
wire _abc_40319_new_n707_; 
wire _abc_40319_new_n708_; 
wire _abc_40319_new_n709_; 
wire _abc_40319_new_n710_; 
wire _abc_40319_new_n711_; 
wire _abc_40319_new_n712_; 
wire _abc_40319_new_n713_; 
wire _abc_40319_new_n714_; 
wire _abc_40319_new_n715_; 
wire _abc_40319_new_n716_; 
wire _abc_40319_new_n717_; 
wire _abc_40319_new_n718_; 
wire _abc_40319_new_n719_; 
wire _abc_40319_new_n720_; 
wire _abc_40319_new_n721_; 
wire _abc_40319_new_n722_; 
wire _abc_40319_new_n723_; 
wire _abc_40319_new_n724_; 
wire _abc_40319_new_n725_; 
wire _abc_40319_new_n726_; 
wire _abc_40319_new_n727_; 
wire _abc_40319_new_n728_; 
wire _abc_40319_new_n729_; 
wire _abc_40319_new_n730_; 
wire _abc_40319_new_n731_; 
wire _abc_40319_new_n732_; 
wire _abc_40319_new_n733_; 
wire _abc_40319_new_n734_; 
wire _abc_40319_new_n735_; 
wire _abc_40319_new_n736_; 
wire _abc_40319_new_n737_; 
wire _abc_40319_new_n738_; 
wire _abc_40319_new_n739_; 
wire _abc_40319_new_n740_; 
wire _abc_40319_new_n741_; 
wire _abc_40319_new_n742_; 
wire _abc_40319_new_n743_; 
wire _abc_40319_new_n744_; 
wire _abc_40319_new_n745_; 
wire _abc_40319_new_n746_; 
wire _abc_40319_new_n747_; 
wire _abc_40319_new_n748_; 
wire _abc_40319_new_n749_; 
wire _abc_40319_new_n750_; 
wire _abc_40319_new_n751_; 
wire _abc_40319_new_n752_; 
wire _abc_40319_new_n753_; 
wire _abc_40319_new_n754_; 
wire _abc_40319_new_n755_; 
wire _abc_40319_new_n756_; 
wire _abc_40319_new_n757_; 
wire _abc_40319_new_n758_; 
wire _abc_40319_new_n759_; 
wire _abc_40319_new_n760_; 
wire _abc_40319_new_n761_; 
wire _abc_40319_new_n762_; 
wire _abc_40319_new_n763_; 
wire _abc_40319_new_n764_; 
wire _abc_40319_new_n765_; 
wire _abc_40319_new_n766_; 
wire _abc_40319_new_n767_; 
wire _abc_40319_new_n768_; 
wire _abc_40319_new_n769_; 
wire _abc_40319_new_n770_; 
wire _abc_40319_new_n771_; 
wire _abc_40319_new_n772_; 
wire _abc_40319_new_n773_; 
wire _abc_40319_new_n774_; 
wire _abc_40319_new_n775_; 
wire _abc_40319_new_n776_; 
wire _abc_40319_new_n777_; 
wire _abc_40319_new_n778_; 
wire _abc_40319_new_n779_; 
wire _abc_40319_new_n780_; 
wire _abc_40319_new_n781_; 
wire _abc_40319_new_n782_; 
wire _abc_40319_new_n783_; 
wire _abc_40319_new_n784_; 
wire _abc_40319_new_n785_; 
wire _abc_40319_new_n786_; 
wire _abc_40319_new_n787_; 
wire _abc_40319_new_n788_; 
wire _abc_40319_new_n789_; 
wire _abc_40319_new_n790_; 
wire _abc_40319_new_n791_; 
wire _abc_40319_new_n792_; 
wire _abc_40319_new_n793_; 
wire _abc_40319_new_n794_; 
wire _abc_40319_new_n795_; 
wire _abc_40319_new_n796_; 
wire _abc_40319_new_n797_; 
wire _abc_40319_new_n798_; 
wire _abc_40319_new_n799_; 
wire _abc_40319_new_n800_; 
wire _abc_40319_new_n801_; 
wire _abc_40319_new_n802_; 
wire _abc_40319_new_n803_; 
wire _abc_40319_new_n804_; 
wire _abc_40319_new_n805_; 
wire _abc_40319_new_n806_; 
wire _abc_40319_new_n807_; 
wire _abc_40319_new_n808_; 
wire _abc_40319_new_n809_; 
wire _abc_40319_new_n810_; 
wire _abc_40319_new_n811_; 
wire _abc_40319_new_n812_; 
wire _abc_40319_new_n813_; 
wire _abc_40319_new_n814_; 
wire _abc_40319_new_n815_; 
wire _abc_40319_new_n816_; 
wire _abc_40319_new_n817_; 
wire _abc_40319_new_n818_; 
wire _abc_40319_new_n819_; 
wire _abc_40319_new_n820_; 
wire _abc_40319_new_n821_; 
wire _abc_40319_new_n822_; 
wire _abc_40319_new_n823_; 
wire _abc_40319_new_n824_; 
wire _abc_40319_new_n825_; 
wire _abc_40319_new_n826_; 
wire _abc_40319_new_n827_; 
wire _abc_40319_new_n828_; 
wire _abc_40319_new_n829_; 
wire _abc_40319_new_n830_; 
wire _abc_40319_new_n831_; 
wire _abc_40319_new_n832_; 
wire _abc_40319_new_n833_; 
wire _abc_40319_new_n834_; 
wire _abc_40319_new_n835_; 
wire _abc_40319_new_n836_; 
wire _abc_40319_new_n837_; 
wire _abc_40319_new_n838_; 
wire _abc_40319_new_n839_; 
wire _abc_40319_new_n840_; 
wire _abc_40319_new_n841_; 
wire _abc_40319_new_n842_; 
wire _abc_40319_new_n843_; 
wire _abc_40319_new_n844_; 
wire _abc_40319_new_n845_; 
wire _abc_40319_new_n846_; 
wire _abc_40319_new_n847_; 
wire _abc_40319_new_n848_; 
wire _abc_40319_new_n849_; 
wire _abc_40319_new_n850_; 
wire _abc_40319_new_n851_; 
wire _abc_40319_new_n852_; 
wire _abc_40319_new_n853_; 
wire _abc_40319_new_n854_; 
wire _abc_40319_new_n855_; 
wire _abc_40319_new_n856_; 
wire _abc_40319_new_n857_; 
wire _abc_40319_new_n858_; 
wire _abc_40319_new_n859_; 
wire _abc_40319_new_n860_; 
wire _abc_40319_new_n861_; 
wire _abc_40319_new_n862_; 
wire _abc_40319_new_n863_; 
wire _abc_40319_new_n864_; 
wire _abc_40319_new_n865_; 
wire _abc_40319_new_n866_; 
wire _abc_40319_new_n867_; 
wire _abc_40319_new_n868_; 
wire _abc_40319_new_n869_; 
wire _abc_40319_new_n870_; 
wire _abc_40319_new_n871_; 
wire _abc_40319_new_n872_; 
wire _abc_40319_new_n873_; 
wire _abc_40319_new_n874_; 
wire _abc_40319_new_n875_; 
wire _abc_40319_new_n876_; 
wire _abc_40319_new_n877_; 
wire _abc_40319_new_n878_; 
wire _abc_40319_new_n879_; 
wire _abc_40319_new_n880_; 
wire _abc_40319_new_n881_; 
wire _abc_40319_new_n882_; 
wire _abc_40319_new_n883_; 
wire _abc_40319_new_n884_; 
wire _abc_40319_new_n885_; 
wire _abc_40319_new_n886_; 
wire _abc_40319_new_n887_; 
wire _abc_40319_new_n888_; 
wire _abc_40319_new_n889_; 
wire _abc_40319_new_n890_; 
wire _abc_40319_new_n891_; 
wire _abc_40319_new_n892_; 
wire _abc_40319_new_n893_; 
wire _abc_40319_new_n894_; 
wire _abc_40319_new_n895_; 
wire _abc_40319_new_n896_; 
wire _abc_40319_new_n897_; 
wire _abc_40319_new_n898_; 
wire _abc_40319_new_n899_; 
wire _abc_40319_new_n900_; 
wire _abc_40319_new_n901_; 
wire _abc_40319_new_n902_; 
wire _abc_40319_new_n903_; 
wire _abc_40319_new_n904_; 
wire _abc_40319_new_n905_; 
wire _abc_40319_new_n906_; 
wire _abc_40319_new_n907_; 
wire _abc_40319_new_n908_; 
wire _abc_40319_new_n909_; 
wire _abc_40319_new_n910_; 
wire _abc_40319_new_n911_; 
wire _abc_40319_new_n912_; 
wire _abc_40319_new_n913_; 
wire _abc_40319_new_n914_; 
wire _abc_40319_new_n915_; 
wire _abc_40319_new_n916_; 
wire _abc_40319_new_n917_; 
wire _abc_40319_new_n918_; 
wire _abc_40319_new_n919_; 
wire _abc_40319_new_n920_; 
wire _abc_40319_new_n921_; 
wire _abc_40319_new_n922_; 
wire _abc_40319_new_n923_; 
wire _abc_40319_new_n924_; 
wire _abc_40319_new_n925_; 
wire _abc_40319_new_n926_; 
wire _abc_40319_new_n927_; 
wire _abc_40319_new_n928_; 
wire _abc_40319_new_n929_; 
wire _abc_40319_new_n930_; 
wire _abc_40319_new_n931_; 
wire _abc_40319_new_n932_; 
wire _abc_40319_new_n933_; 
wire _abc_40319_new_n934_; 
wire _abc_40319_new_n935_; 
wire _abc_40319_new_n936_; 
wire _abc_40319_new_n937_; 
wire _abc_40319_new_n938_; 
wire _abc_40319_new_n939_; 
wire _abc_40319_new_n940_; 
wire _abc_40319_new_n941_; 
wire _abc_40319_new_n942_; 
wire _abc_40319_new_n943_; 
wire _abc_40319_new_n944_; 
wire _abc_40319_new_n945_; 
wire _abc_40319_new_n946_; 
wire _abc_40319_new_n947_; 
wire _abc_40319_new_n948_; 
wire _abc_40319_new_n949_; 
wire _abc_40319_new_n950_; 
wire _abc_40319_new_n951_; 
wire _abc_40319_new_n952_; 
wire _abc_40319_new_n953_; 
wire _abc_40319_new_n954_; 
wire _abc_40319_new_n955_; 
wire _abc_40319_new_n956_; 
wire _abc_40319_new_n957_; 
wire _abc_40319_new_n958_; 
wire _abc_40319_new_n959_; 
wire _abc_40319_new_n960_; 
wire _abc_40319_new_n961_; 
wire _abc_40319_new_n962_; 
wire _abc_40319_new_n963_; 
wire _abc_40319_new_n964_; 
wire _abc_40319_new_n965_; 
wire _abc_40319_new_n966_; 
wire _abc_40319_new_n967_; 
wire _abc_40319_new_n968_; 
wire _abc_40319_new_n969_; 
wire _abc_40319_new_n970_; 
wire _abc_40319_new_n971_; 
wire _abc_40319_new_n972_; 
wire _abc_40319_new_n973_; 
wire _abc_40319_new_n974_; 
wire _abc_40319_new_n975_; 
wire _abc_40319_new_n976_; 
wire _abc_40319_new_n977_; 
wire _abc_40319_new_n978_; 
wire _abc_40319_new_n979_; 
wire _abc_40319_new_n980_; 
wire _abc_40319_new_n981_; 
wire _abc_40319_new_n982_; 
wire _abc_40319_new_n983_; 
wire _abc_40319_new_n984_; 
wire _abc_40319_new_n985_; 
wire _abc_40319_new_n986_; 
wire _abc_40319_new_n987_; 
wire _abc_40319_new_n988_; 
wire _abc_40319_new_n989_; 
wire _abc_40319_new_n990_; 
wire _abc_40319_new_n991_; 
wire _abc_40319_new_n992_; 
wire _abc_40319_new_n993_; 
wire _abc_40319_new_n994_; 
wire _abc_40319_new_n995_; 
wire _abc_40319_new_n996_; 
wire _abc_40319_new_n997_; 
wire _abc_40319_new_n998_; 
wire _abc_40319_new_n999_; 
input clock;
wire n1002; 
wire n1006; 
wire n1010; 
wire n1014; 
wire n1018; 
wire n1022; 
wire n1026; 
wire n1030; 
wire n1034; 
wire n1038; 
wire n1042; 
wire n1046; 
wire n1050; 
wire n1054; 
wire n1058; 
wire n1062; 
wire n1066; 
wire n1070; 
wire n1074; 
wire n1078; 
wire n1082; 
wire n1086; 
wire n1090; 
wire n1094; 
wire n1098; 
wire n1102; 
wire n1106; 
wire n1110; 
wire n1114; 
wire n1118; 
wire n1122; 
wire n1126; 
wire n1130; 
wire n1134; 
wire n1138; 
wire n1142; 
wire n1146; 
wire n1150; 
wire n1154; 
wire n1158; 
wire n1162; 
wire n1166; 
wire n1170; 
wire n1174; 
wire n1178; 
wire n1182; 
wire n1186; 
wire n1191; 
wire n1196; 
wire n1201; 
wire n1206; 
wire n1211; 
wire n1216; 
wire n1221; 
wire n1226; 
wire n1231; 
wire n1236; 
wire n1241; 
wire n1246; 
wire n1251; 
wire n1256; 
wire n1261; 
wire n1266; 
wire n1271; 
wire n1276; 
wire n1281; 
wire n1286; 
wire n1291; 
wire n1296; 
wire n1301; 
wire n1306; 
wire n1311; 
wire n1316; 
wire n1321; 
wire n1326; 
wire n1331; 
wire n1336; 
wire n1341; 
wire n1345; 
wire n178; 
wire n183; 
wire n188; 
wire n193; 
wire n198; 
wire n203; 
wire n208; 
wire n213; 
wire n218; 
wire n223; 
wire n228; 
wire n233; 
wire n238; 
wire n243; 
wire n248; 
wire n253; 
wire n258; 
wire n263; 
wire n268; 
wire n273; 
wire n278; 
wire n283; 
wire n288; 
wire n293; 
wire n298; 
wire n303; 
wire n308; 
wire n313; 
wire n318; 
wire n323; 
wire n328; 
wire n333; 
wire n338; 
wire n343; 
wire n348; 
wire n353; 
wire n358; 
wire n363; 
wire n368; 
wire n373; 
wire n378; 
wire n383; 
wire n388; 
wire n393; 
wire n398; 
wire n403; 
wire n408; 
wire n413; 
wire n418; 
wire n423; 
wire n428; 
wire n433; 
wire n438; 
wire n443; 
wire n448; 
wire n453; 
wire n458; 
wire n463; 
wire n468; 
wire n473; 
wire n478; 
wire n483; 
wire n488; 
wire n493; 
wire n498; 
wire n503; 
wire n508; 
wire n513; 
wire n518; 
wire n523; 
wire n528; 
wire n533; 
wire n538; 
wire n543; 
wire n548; 
wire n553; 
wire n558; 
wire n563; 
wire n568; 
wire n573; 
wire n578; 
wire n583; 
wire n588; 
wire n593; 
wire n598; 
wire n603; 
wire n608; 
wire n613; 
wire n618; 
wire n623; 
wire n628; 
wire n633; 
wire n638; 
wire n643; 
wire n648; 
wire n653; 
wire n658; 
wire n663; 
wire n668; 
wire n673; 
wire n678; 
wire n683; 
wire n688; 
wire n693; 
wire n698; 
wire n703; 
wire n708; 
wire n713; 
wire n718; 
wire n723; 
wire n728; 
wire n733; 
wire n738; 
wire n743; 
wire n748; 
wire n753; 
wire n758; 
wire n763; 
wire n768; 
wire n773; 
wire n778; 
wire n783; 
wire n788; 
wire n793; 
wire n798; 
wire n803; 
wire n808; 
wire n813; 
wire n818; 
wire n823; 
wire n828; 
wire n833; 
wire n838; 
wire n843; 
wire n848; 
wire n853; 
wire n858; 
wire n863; 
wire n868; 
wire n873; 
wire n878; 
wire n883; 
wire n888; 
wire n893; 
wire n898; 
wire n903; 
wire n908; 
wire n913; 
wire n918; 
wire n923; 
wire n928; 
wire n933; 
wire n938; 
wire n943; 
wire n948; 
wire n953; 
wire n958; 
wire n963; 
wire n968; 
wire n973; 
wire n978; 
wire n982; 
wire n986; 
wire n990; 
wire n994; 
wire n998; 
input nRESET_G;
AND2X2 AND2X2_1 ( .A(_abc_40319_new_n530_), .B(_abc_40319_new_n529_), .Y(_abc_40319_new_n551_));
AND2X2 AND2X2_10 ( .A(_abc_40319_new_n744_), .B(_abc_40319_new_n574_), .Y(_abc_40319_new_n745_));
AND2X2 AND2X2_100 ( .A(_abc_40319_new_n3617_), .B(_abc_40319_new_n3618_), .Y(_abc_40319_new_n3619_));
AND2X2 AND2X2_101 ( .A(_abc_40319_new_n3620_), .B(_abc_40319_new_n2962_), .Y(_abc_40319_new_n3636_));
AND2X2 AND2X2_102 ( .A(_abc_40319_new_n3642_), .B(_abc_40319_new_n3640_), .Y(_abc_40319_new_n3643_));
AND2X2 AND2X2_103 ( .A(_abc_40319_new_n3833_), .B(_abc_40319_new_n3831_), .Y(_abc_40319_new_n3834_));
AND2X2 AND2X2_104 ( .A(_abc_40319_new_n3855_), .B(_abc_40319_new_n3856_), .Y(_abc_40319_new_n3857_));
AND2X2 AND2X2_105 ( .A(_abc_40319_new_n3858_), .B(REG3_REG_13_), .Y(_abc_40319_new_n3859_));
AND2X2 AND2X2_106 ( .A(_abc_40319_new_n3865_), .B(REG3_REG_22_), .Y(_abc_40319_new_n3866_));
AND2X2 AND2X2_107 ( .A(_abc_40319_new_n3868_), .B(REG3_REG_26_), .Y(_abc_40319_new_n3869_));
AND2X2 AND2X2_108 ( .A(_abc_40319_new_n3902_), .B(nRESET_G), .Y(_abc_40319_new_n3903_));
AND2X2 AND2X2_109 ( .A(_abc_40319_new_n3637_), .B(_abc_40319_new_n3638_), .Y(_abc_40319_new_n3905_));
AND2X2 AND2X2_11 ( .A(_abc_40319_new_n574_), .B(_abc_40319_new_n750_), .Y(_abc_40319_new_n751_));
AND2X2 AND2X2_110 ( .A(_abc_40319_new_n3472_), .B(_abc_40319_new_n3963_), .Y(_abc_40319_new_n3964_));
AND2X2 AND2X2_111 ( .A(_abc_40319_new_n3985_), .B(nRESET_G), .Y(_abc_40319_new_n3986_));
AND2X2 AND2X2_112 ( .A(_abc_40319_new_n4086_), .B(nRESET_G), .Y(_abc_40319_new_n4087_));
AND2X2 AND2X2_113 ( .A(_abc_40319_new_n4118_), .B(nRESET_G), .Y(_abc_40319_new_n4119_));
AND2X2 AND2X2_114 ( .A(_abc_40319_new_n4121_), .B(nRESET_G), .Y(_abc_40319_new_n4122_));
AND2X2 AND2X2_115 ( .A(_abc_40319_new_n4128_), .B(nRESET_G), .Y(_abc_40319_new_n4129_));
AND2X2 AND2X2_12 ( .A(_abc_40319_new_n873_), .B(_abc_40319_new_n874_), .Y(_abc_40319_new_n875_));
AND2X2 AND2X2_13 ( .A(_abc_40319_new_n938_), .B(_abc_40319_new_n939_), .Y(_abc_40319_new_n940_));
AND2X2 AND2X2_14 ( .A(_abc_40319_new_n946_), .B(_abc_40319_new_n947_), .Y(_abc_40319_new_n948_));
AND2X2 AND2X2_15 ( .A(_abc_40319_new_n983_), .B(_abc_40319_new_n981_), .Y(_abc_40319_new_n984_));
AND2X2 AND2X2_16 ( .A(_abc_40319_new_n1033_), .B(REG3_REG_20_), .Y(_abc_40319_new_n1034_));
AND2X2 AND2X2_17 ( .A(_abc_40319_new_n1088_), .B(_abc_40319_new_n1092_), .Y(_abc_40319_new_n1093_));
AND2X2 AND2X2_18 ( .A(_abc_40319_new_n1106_), .B(_abc_40319_new_n1069_), .Y(_abc_40319_new_n1107_));
AND2X2 AND2X2_19 ( .A(_abc_40319_new_n1131_), .B(_abc_40319_new_n1132_), .Y(_abc_40319_new_n1133_));
AND2X2 AND2X2_2 ( .A(_abc_40319_new_n581_), .B(STATE_REG), .Y(_abc_40319_new_n582_));
AND2X2 AND2X2_20 ( .A(_abc_40319_new_n1167_), .B(_abc_40319_new_n1241_), .Y(_abc_40319_new_n1242_));
AND2X2 AND2X2_21 ( .A(_abc_40319_new_n1229_), .B(_abc_40319_new_n1254_), .Y(_abc_40319_new_n1255_));
AND2X2 AND2X2_22 ( .A(_abc_40319_new_n1268_), .B(_abc_40319_new_n1269_), .Y(_abc_40319_new_n1270_));
AND2X2 AND2X2_23 ( .A(_abc_40319_new_n1290_), .B(_abc_40319_new_n1291_), .Y(_abc_40319_new_n1292_));
AND2X2 AND2X2_24 ( .A(_abc_40319_new_n1299_), .B(_abc_40319_new_n1301_), .Y(_abc_40319_new_n1302_));
AND2X2 AND2X2_25 ( .A(_abc_40319_new_n1180_), .B(_abc_40319_new_n1329_), .Y(_abc_40319_new_n1330_));
AND2X2 AND2X2_26 ( .A(_abc_40319_new_n1346_), .B(_abc_40319_new_n1347_), .Y(_abc_40319_new_n1348_));
AND2X2 AND2X2_27 ( .A(_abc_40319_new_n1349_), .B(_abc_40319_new_n1351_), .Y(_abc_40319_new_n1352_));
AND2X2 AND2X2_28 ( .A(_abc_40319_new_n1364_), .B(_abc_40319_new_n1340_), .Y(_abc_40319_new_n1365_));
AND2X2 AND2X2_29 ( .A(_abc_40319_new_n1493_), .B(_abc_40319_new_n1053_), .Y(_abc_40319_new_n1494_));
AND2X2 AND2X2_3 ( .A(_abc_40319_new_n612_), .B(_abc_40319_new_n576_), .Y(_abc_40319_new_n613_));
AND2X2 AND2X2_30 ( .A(_abc_40319_new_n1522_), .B(_abc_40319_new_n1518_), .Y(_abc_40319_new_n1523_));
AND2X2 AND2X2_31 ( .A(_abc_40319_new_n1544_), .B(_abc_40319_new_n1540_), .Y(_abc_40319_new_n1545_));
AND2X2 AND2X2_32 ( .A(_abc_40319_new_n1427_), .B(_abc_40319_new_n1163_), .Y(_abc_40319_new_n1563_));
AND2X2 AND2X2_33 ( .A(_abc_40319_new_n1574_), .B(_abc_40319_new_n1569_), .Y(_abc_40319_new_n1575_));
AND2X2 AND2X2_34 ( .A(_abc_40319_new_n1488_), .B(_abc_40319_new_n1120_), .Y(_abc_40319_new_n1577_));
AND2X2 AND2X2_35 ( .A(_abc_40319_new_n1597_), .B(_abc_40319_new_n1593_), .Y(_abc_40319_new_n1598_));
AND2X2 AND2X2_36 ( .A(_abc_40319_new_n1600_), .B(_abc_40319_new_n1604_), .Y(_abc_40319_new_n1605_));
AND2X2 AND2X2_37 ( .A(_abc_40319_new_n1286_), .B(_abc_40319_new_n1285_), .Y(_abc_40319_new_n1610_));
AND2X2 AND2X2_38 ( .A(_abc_40319_new_n1638_), .B(_abc_40319_new_n676_), .Y(_abc_40319_new_n1639_));
AND2X2 AND2X2_39 ( .A(_abc_40319_new_n1648_), .B(_abc_40319_new_n1645_), .Y(_abc_40319_new_n1649_));
AND2X2 AND2X2_4 ( .A(_abc_40319_new_n641_), .B(_abc_40319_new_n642_), .Y(_abc_40319_new_n643_));
AND2X2 AND2X2_40 ( .A(_abc_40319_new_n1657_), .B(_abc_40319_new_n1653_), .Y(_abc_40319_new_n1658_));
AND2X2 AND2X2_41 ( .A(_abc_40319_new_n1660_), .B(_abc_40319_new_n1103_), .Y(_abc_40319_new_n1661_));
AND2X2 AND2X2_42 ( .A(_abc_40319_new_n1674_), .B(_abc_40319_new_n1676_), .Y(_abc_40319_new_n1677_));
AND2X2 AND2X2_43 ( .A(_abc_40319_new_n1696_), .B(_abc_40319_new_n1215_), .Y(_abc_40319_new_n1697_));
AND2X2 AND2X2_44 ( .A(_abc_40319_new_n870_), .B(_abc_40319_new_n934_), .Y(_abc_40319_new_n1719_));
AND2X2 AND2X2_45 ( .A(_abc_40319_new_n1732_), .B(_abc_40319_new_n1314_), .Y(_abc_40319_new_n1733_));
AND2X2 AND2X2_46 ( .A(_abc_40319_new_n1733_), .B(_abc_40319_new_n1316_), .Y(_abc_40319_new_n1734_));
AND2X2 AND2X2_47 ( .A(_abc_40319_new_n1743_), .B(_abc_40319_new_n1738_), .Y(_abc_40319_new_n1744_));
AND2X2 AND2X2_48 ( .A(_abc_40319_new_n1802_), .B(_abc_40319_new_n1798_), .Y(_abc_40319_new_n1803_));
AND2X2 AND2X2_49 ( .A(_abc_40319_new_n1422_), .B(_abc_40319_new_n1426_), .Y(_abc_40319_new_n1818_));
AND2X2 AND2X2_5 ( .A(_abc_40319_new_n573_), .B(_abc_40319_new_n560_), .Y(_abc_40319_new_n671_));
AND2X2 AND2X2_50 ( .A(_abc_40319_new_n937_), .B(_abc_40319_new_n1831_), .Y(_abc_40319_new_n1832_));
AND2X2 AND2X2_51 ( .A(_abc_40319_new_n1056_), .B(_abc_40319_new_n1059_), .Y(_abc_40319_new_n1852_));
AND2X2 AND2X2_52 ( .A(_abc_40319_new_n1851_), .B(_abc_40319_new_n1855_), .Y(_abc_40319_new_n1856_));
AND2X2 AND2X2_53 ( .A(_abc_40319_new_n1420_), .B(_abc_40319_new_n1265_), .Y(_abc_40319_new_n1858_));
AND2X2 AND2X2_54 ( .A(_abc_40319_new_n715_), .B(REG2_REG_31_), .Y(_abc_40319_new_n1878_));
AND2X2 AND2X2_55 ( .A(_abc_40319_new_n1899_), .B(_abc_40319_new_n1898_), .Y(_abc_40319_new_n1900_));
AND2X2 AND2X2_56 ( .A(_abc_40319_new_n1988_), .B(_abc_40319_new_n1989_), .Y(_abc_40319_new_n1995_));
AND2X2 AND2X2_57 ( .A(_abc_40319_new_n715_), .B(REG2_REG_30_), .Y(_abc_40319_new_n2098_));
AND2X2 AND2X2_58 ( .A(_abc_40319_new_n2197_), .B(_abc_40319_new_n2198_), .Y(_abc_40319_new_n2199_));
AND2X2 AND2X2_59 ( .A(_abc_40319_new_n2254_), .B(_abc_40319_new_n2139_), .Y(_abc_40319_new_n2255_));
AND2X2 AND2X2_6 ( .A(_abc_40319_new_n574_), .B(_abc_40319_new_n678_), .Y(_abc_40319_new_n679_));
AND2X2 AND2X2_60 ( .A(_abc_40319_new_n1902_), .B(_abc_40319_new_n1875_), .Y(_abc_40319_new_n2276_));
AND2X2 AND2X2_61 ( .A(_abc_40319_new_n2315_), .B(_abc_40319_new_n2123_), .Y(_abc_40319_new_n2316_));
AND2X2 AND2X2_62 ( .A(_abc_40319_new_n2248_), .B(_abc_40319_new_n2232_), .Y(_abc_40319_new_n2356_));
AND2X2 AND2X2_63 ( .A(_abc_40319_new_n2384_), .B(_abc_40319_new_n2221_), .Y(_abc_40319_new_n2385_));
AND2X2 AND2X2_64 ( .A(_abc_40319_new_n2434_), .B(_abc_40319_new_n2348_), .Y(_abc_40319_new_n2435_));
AND2X2 AND2X2_65 ( .A(_abc_40319_new_n2424_), .B(_abc_40319_new_n2436_), .Y(_abc_40319_new_n2437_));
AND2X2 AND2X2_66 ( .A(_abc_40319_new_n2469_), .B(_abc_40319_new_n2243_), .Y(_abc_40319_new_n2470_));
AND2X2 AND2X2_67 ( .A(_abc_40319_new_n2478_), .B(_abc_40319_new_n2467_), .Y(_abc_40319_new_n2479_));
AND2X2 AND2X2_68 ( .A(_abc_40319_new_n2322_), .B(_abc_40319_new_n2221_), .Y(_abc_40319_new_n2493_));
AND2X2 AND2X2_69 ( .A(_abc_40319_new_n2502_), .B(_abc_40319_new_n2131_), .Y(_abc_40319_new_n2503_));
AND2X2 AND2X2_7 ( .A(_abc_40319_new_n686_), .B(_abc_40319_new_n687_), .Y(_abc_40319_new_n688_));
AND2X2 AND2X2_70 ( .A(_abc_40319_new_n2269_), .B(_abc_40319_new_n2116_), .Y(_abc_40319_new_n2516_));
AND2X2 AND2X2_71 ( .A(_abc_40319_new_n2607_), .B(_abc_40319_new_n2593_), .Y(_abc_40319_new_n2608_));
AND2X2 AND2X2_72 ( .A(_abc_40319_new_n2629_), .B(_abc_40319_new_n2628_), .Y(_abc_40319_new_n2630_));
AND2X2 AND2X2_73 ( .A(_abc_40319_new_n2651_), .B(_abc_40319_new_n2655_), .Y(_abc_40319_new_n2656_));
AND2X2 AND2X2_74 ( .A(_abc_40319_new_n2666_), .B(_abc_40319_new_n2697_), .Y(_abc_40319_new_n2698_));
AND2X2 AND2X2_75 ( .A(_abc_40319_new_n2799_), .B(_abc_40319_new_n2798_), .Y(_abc_40319_new_n2800_));
AND2X2 AND2X2_76 ( .A(_abc_40319_new_n2796_), .B(_abc_40319_new_n2800_), .Y(_abc_40319_new_n2801_));
AND2X2 AND2X2_77 ( .A(_abc_40319_new_n2784_), .B(_abc_40319_new_n1322_), .Y(_abc_40319_new_n2805_));
AND2X2 AND2X2_78 ( .A(_abc_40319_new_n2803_), .B(_abc_40319_new_n1252_), .Y(_abc_40319_new_n2808_));
AND2X2 AND2X2_79 ( .A(_abc_40319_new_n2893_), .B(_abc_40319_new_n2896_), .Y(_abc_40319_new_n2897_));
AND2X2 AND2X2_8 ( .A(_abc_40319_new_n600_), .B(IR_REG_29_), .Y(_abc_40319_new_n713_));
AND2X2 AND2X2_80 ( .A(_abc_40319_new_n2952_), .B(_abc_40319_new_n2951_), .Y(_abc_40319_new_n2953_));
AND2X2 AND2X2_81 ( .A(_abc_40319_new_n2981_), .B(_abc_40319_new_n2983_), .Y(_abc_40319_new_n2984_));
AND2X2 AND2X2_82 ( .A(_abc_40319_new_n3083_), .B(_abc_40319_new_n3078_), .Y(_abc_40319_new_n3084_));
AND2X2 AND2X2_83 ( .A(_abc_40319_new_n3077_), .B(_abc_40319_new_n3084_), .Y(_abc_40319_new_n3085_));
AND2X2 AND2X2_84 ( .A(_abc_40319_new_n2504_), .B(_abc_40319_new_n2464_), .Y(_abc_40319_new_n3126_));
AND2X2 AND2X2_85 ( .A(_abc_40319_new_n3127_), .B(_abc_40319_new_n3119_), .Y(_abc_40319_new_n3128_));
AND2X2 AND2X2_86 ( .A(_abc_40319_new_n3162_), .B(_abc_40319_new_n3135_), .Y(_abc_40319_new_n3163_));
AND2X2 AND2X2_87 ( .A(_abc_40319_new_n3184_), .B(_abc_40319_new_n2129_), .Y(_abc_40319_new_n3185_));
AND2X2 AND2X2_88 ( .A(_abc_40319_new_n3161_), .B(_abc_40319_new_n3212_), .Y(_abc_40319_new_n3213_));
AND2X2 AND2X2_89 ( .A(_abc_40319_new_n3225_), .B(_abc_40319_new_n2976_), .Y(_abc_40319_new_n3226_));
AND2X2 AND2X2_9 ( .A(_abc_40319_new_n711_), .B(IR_REG_30_), .Y(_abc_40319_new_n718_));
AND2X2 AND2X2_90 ( .A(_abc_40319_new_n3250_), .B(_abc_40319_new_n3211_), .Y(_abc_40319_new_n3251_));
AND2X2 AND2X2_91 ( .A(_abc_40319_new_n3224_), .B(_abc_40319_new_n3276_), .Y(_abc_40319_new_n3277_));
AND2X2 AND2X2_92 ( .A(_abc_40319_new_n3333_), .B(_abc_40319_new_n3298_), .Y(_abc_40319_new_n3334_));
AND2X2 AND2X2_93 ( .A(_abc_40319_new_n3344_), .B(_abc_40319_new_n3101_), .Y(_abc_40319_new_n3345_));
AND2X2 AND2X2_94 ( .A(_abc_40319_new_n3332_), .B(_abc_40319_new_n3378_), .Y(_abc_40319_new_n3379_));
AND2X2 AND2X2_95 ( .A(_abc_40319_new_n3416_), .B(_abc_40319_new_n3377_), .Y(_abc_40319_new_n3417_));
AND2X2 AND2X2_96 ( .A(_abc_40319_new_n3460_), .B(_abc_40319_new_n2970_), .Y(_abc_40319_new_n3461_));
AND2X2 AND2X2_97 ( .A(_abc_40319_new_n2968_), .B(_abc_40319_new_n3536_), .Y(_abc_40319_new_n3537_));
AND2X2 AND2X2_98 ( .A(_abc_40319_new_n2966_), .B(_abc_40319_new_n3586_), .Y(_abc_40319_new_n3587_));
AND2X2 AND2X2_99 ( .A(_abc_40319_new_n2996_), .B(_abc_40319_new_n3587_), .Y(_abc_40319_new_n3588_));
AOI21X1 AOI21X1_1 ( .A(_abc_40319_new_n532_), .B(_abc_40319_new_n541_), .C(_abc_40319_new_n568_), .Y(_abc_40319_new_n578_));
AOI21X1 AOI21X1_10 ( .A(_abc_40319_new_n852_), .B(_abc_40319_new_n812_), .C(_abc_40319_new_n853_), .Y(_abc_40319_new_n854_));
AOI21X1 AOI21X1_100 ( .A(_abc_40319_new_n878_), .B(_abc_40319_new_n879_), .C(_abc_40319_new_n580_), .Y(_abc_40319_new_n1891_));
AOI21X1 AOI21X1_101 ( .A(_abc_40319_new_n841_), .B(_abc_40319_new_n840_), .C(_abc_40319_new_n580_), .Y(_abc_40319_new_n1911_));
AOI21X1 AOI21X1_102 ( .A(_abc_40319_new_n809_), .B(_abc_40319_new_n1874_), .C(_abc_40319_new_n1917_), .Y(_abc_40319_new_n1918_));
AOI21X1 AOI21X1_103 ( .A(_abc_40319_new_n1937_), .B(_abc_40319_new_n1936_), .C(_abc_40319_new_n1939_), .Y(_abc_40319_new_n1967_));
AOI21X1 AOI21X1_104 ( .A(_abc_40319_new_n1948_), .B(_abc_40319_new_n1947_), .C(_abc_40319_new_n1950_), .Y(_abc_40319_new_n1973_));
AOI21X1 AOI21X1_105 ( .A(_abc_40319_new_n1979_), .B(_abc_40319_new_n1984_), .C(_abc_40319_new_n1990_), .Y(_abc_40319_new_n1991_));
AOI21X1 AOI21X1_106 ( .A(_abc_40319_new_n1943_), .B(_abc_40319_new_n1970_), .C(_abc_40319_new_n1992_), .Y(_abc_40319_new_n1993_));
AOI21X1 AOI21X1_107 ( .A(_abc_40319_new_n1994_), .B(_abc_40319_new_n1995_), .C(_abc_40319_new_n2002_), .Y(_abc_40319_new_n2003_));
AOI21X1 AOI21X1_108 ( .A(_abc_40319_new_n1233_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n2006_), .Y(_abc_40319_new_n2007_));
AOI21X1 AOI21X1_109 ( .A(_abc_40319_new_n2007_), .B(_abc_40319_new_n2008_), .C(_abc_40319_new_n2005_), .Y(_abc_40319_new_n2009_));
AOI21X1 AOI21X1_11 ( .A(_abc_40319_new_n852_), .B(_abc_40319_new_n812_), .C(_abc_40319_new_n825_), .Y(_abc_40319_new_n864_));
AOI21X1 AOI21X1_110 ( .A(_abc_40319_new_n2010_), .B(_abc_40319_new_n2016_), .C(_abc_40319_new_n2020_), .Y(_abc_40319_new_n2021_));
AOI21X1 AOI21X1_111 ( .A(_abc_40319_new_n1157_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n2023_), .Y(_abc_40319_new_n2024_));
AOI21X1 AOI21X1_112 ( .A(_abc_40319_new_n2034_), .B(_abc_40319_new_n2039_), .C(_abc_40319_new_n2043_), .Y(_abc_40319_new_n2044_));
AOI21X1 AOI21X1_113 ( .A(_abc_40319_new_n1135_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n2046_), .Y(_abc_40319_new_n2047_));
AOI21X1 AOI21X1_114 ( .A(_abc_40319_new_n2055_), .B(_abc_40319_new_n2062_), .C(_abc_40319_new_n2066_), .Y(_abc_40319_new_n2067_));
AOI21X1 AOI21X1_115 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1018_), .C(_abc_40319_new_n2075_), .Y(_abc_40319_new_n2076_));
AOI21X1 AOI21X1_116 ( .A(_abc_40319_new_n2087_), .B(_abc_40319_new_n2093_), .C(_abc_40319_new_n2111_), .Y(_abc_40319_new_n2112_));
AOI21X1 AOI21X1_117 ( .A(_abc_40319_new_n840_), .B(_abc_40319_new_n841_), .C(_abc_40319_new_n1888_), .Y(_abc_40319_new_n2271_));
AOI21X1 AOI21X1_118 ( .A(_abc_40319_new_n830_), .B(_abc_40319_new_n831_), .C(_abc_40319_new_n1888_), .Y(_abc_40319_new_n2279_));
AOI21X1 AOI21X1_119 ( .A(_abc_40319_new_n2282_), .B(_abc_40319_new_n1921_), .C(_abc_40319_new_n1941_), .Y(_abc_40319_new_n2283_));
AOI21X1 AOI21X1_12 ( .A(_abc_40319_new_n858_), .B(_abc_40319_new_n833_), .C(_abc_40319_new_n868_), .Y(_abc_40319_new_n869_));
AOI21X1 AOI21X1_120 ( .A(_abc_40319_new_n1929_), .B(_abc_40319_new_n2284_), .C(_abc_40319_new_n2287_), .Y(_abc_40319_new_n2288_));
AOI21X1 AOI21X1_121 ( .A(_abc_40319_new_n2283_), .B(_abc_40319_new_n1923_), .C(_abc_40319_new_n2290_), .Y(_abc_40319_new_n2291_));
AOI21X1 AOI21X1_122 ( .A(_abc_40319_new_n2292_), .B(_abc_40319_new_n2009_), .C(_abc_40319_new_n2015_), .Y(_abc_40319_new_n2293_));
AOI21X1 AOI21X1_123 ( .A(_abc_40319_new_n2295_), .B(_abc_40319_new_n2033_), .C(_abc_40319_new_n2296_), .Y(_abc_40319_new_n2297_));
AOI21X1 AOI21X1_124 ( .A(_abc_40319_new_n2299_), .B(_abc_40319_new_n2054_), .C(_abc_40319_new_n2061_), .Y(_abc_40319_new_n2300_));
AOI21X1 AOI21X1_125 ( .A(_abc_40319_new_n2301_), .B(_abc_40319_new_n2078_), .C(_abc_40319_new_n2085_), .Y(_abc_40319_new_n2302_));
AOI21X1 AOI21X1_126 ( .A(_abc_40319_new_n2264_), .B(_abc_40319_new_n2088_), .C(_abc_40319_new_n2150_), .Y(_abc_40319_new_n2307_));
AOI21X1 AOI21X1_127 ( .A(_abc_40319_new_n1077_), .B(_abc_40319_new_n1070_), .C(_abc_40319_new_n2133_), .Y(_abc_40319_new_n2315_));
AOI21X1 AOI21X1_128 ( .A(_abc_40319_new_n2412_), .B(_abc_40319_new_n2118_), .C(_abc_40319_new_n2265_), .Y(_abc_40319_new_n2413_));
AOI21X1 AOI21X1_129 ( .A(_abc_40319_new_n2423_), .B(_abc_40319_new_n2357_), .C(_abc_40319_new_n2146_), .Y(_abc_40319_new_n2424_));
AOI21X1 AOI21X1_13 ( .A(_abc_40319_new_n834_), .B(_abc_40319_new_n859_), .C(_abc_40319_new_n869_), .Y(_abc_40319_new_n870_));
AOI21X1 AOI21X1_130 ( .A(_abc_40319_new_n2311_), .B(_abc_40319_new_n2435_), .C(_abc_40319_new_n2432_), .Y(_abc_40319_new_n2436_));
AOI21X1 AOI21X1_131 ( .A(_abc_40319_new_n2401_), .B(_abc_40319_new_n2311_), .C(_abc_40319_new_n2438_), .Y(_abc_40319_new_n2439_));
AOI21X1 AOI21X1_132 ( .A(_abc_40319_new_n2439_), .B(_abc_40319_new_n616_), .C(_abc_40319_new_n663_), .Y(_abc_40319_new_n2440_));
AOI21X1 AOI21X1_133 ( .A(_abc_40319_new_n1115_), .B(_abc_40319_new_n1108_), .C(_abc_40319_new_n2312_), .Y(_abc_40319_new_n2457_));
AOI21X1 AOI21X1_134 ( .A(_abc_40319_new_n2463_), .B(_abc_40319_new_n2128_), .C(_abc_40319_new_n2455_), .Y(_abc_40319_new_n2464_));
AOI21X1 AOI21X1_135 ( .A(_abc_40319_new_n944_), .B(_abc_40319_new_n959_), .C(_abc_40319_new_n2234_), .Y(_abc_40319_new_n2472_));
AOI21X1 AOI21X1_136 ( .A(_abc_40319_new_n2471_), .B(_abc_40319_new_n2474_), .C(_abc_40319_new_n2476_), .Y(_abc_40319_new_n2477_));
AOI21X1 AOI21X1_137 ( .A(_abc_40319_new_n2504_), .B(_abc_40319_new_n2464_), .C(_abc_40319_new_n2454_), .Y(_abc_40319_new_n2505_));
AOI21X1 AOI21X1_138 ( .A(_abc_40319_new_n2106_), .B(_abc_40319_new_n2097_), .C(_abc_40319_new_n2146_), .Y(_abc_40319_new_n2507_));
AOI21X1 AOI21X1_139 ( .A(_abc_40319_new_n2263_), .B(_abc_40319_new_n2507_), .C(_abc_40319_new_n2144_), .Y(_abc_40319_new_n2511_));
AOI21X1 AOI21X1_14 ( .A(_abc_40319_new_n852_), .B(_abc_40319_new_n812_), .C(_abc_40319_new_n895_), .Y(_abc_40319_new_n896_));
AOI21X1 AOI21X1_140 ( .A(_abc_40319_new_n2442_), .B(_abc_40319_new_n749_), .C(_abc_40319_new_n2521_), .Y(_abc_40319_new_n2522_));
AOI21X1 AOI21X1_141 ( .A(_abc_40319_new_n2528_), .B(B_REG), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n2529_));
AOI21X1 AOI21X1_142 ( .A(_abc_40319_new_n2523_), .B(_abc_40319_new_n2533_), .C(_abc_40319_new_n2536_), .Y(_abc_40319_new_n2537_));
AOI21X1 AOI21X1_143 ( .A(_abc_40319_new_n2539_), .B(ADDR_REG_0_), .C(_abc_40319_new_n1752_), .Y(_abc_40319_new_n2540_));
AOI21X1 AOI21X1_144 ( .A(_abc_40319_new_n2539_), .B(ADDR_REG_1_), .C(_abc_40319_new_n1625_), .Y(_abc_40319_new_n2557_));
AOI21X1 AOI21X1_145 ( .A(_abc_40319_new_n2539_), .B(ADDR_REG_2_), .C(_abc_40319_new_n1813_), .Y(_abc_40319_new_n2562_));
AOI21X1 AOI21X1_146 ( .A(_abc_40319_new_n875_), .B(_abc_40319_new_n2546_), .C(_abc_40319_new_n2545_), .Y(_abc_40319_new_n2564_));
AOI21X1 AOI21X1_147 ( .A(_abc_40319_new_n892_), .B(_abc_40319_new_n2551_), .C(_abc_40319_new_n2571_), .Y(_abc_40319_new_n2572_));
AOI21X1 AOI21X1_148 ( .A(_abc_40319_new_n2583_), .B(_abc_40319_new_n2584_), .C(_abc_40319_new_n821_), .Y(_abc_40319_new_n2585_));
AOI21X1 AOI21X1_149 ( .A(_abc_40319_new_n2524_), .B(_abc_40319_new_n2580_), .C(_abc_40319_new_n2589_), .Y(_abc_40319_new_n2590_));
AOI21X1 AOI21X1_15 ( .A(_abc_40319_new_n852_), .B(_abc_40319_new_n812_), .C(_abc_40319_new_n922_), .Y(_abc_40319_new_n923_));
AOI21X1 AOI21X1_150 ( .A(_abc_40319_new_n2539_), .B(ADDR_REG_3_), .C(_abc_40319_new_n1558_), .Y(_abc_40319_new_n2591_));
AOI21X1 AOI21X1_151 ( .A(_abc_40319_new_n2542_), .B(_abc_40319_new_n2603_), .C(_abc_40319_new_n1727_), .Y(_abc_40319_new_n2605_));
AOI21X1 AOI21X1_152 ( .A(_abc_40319_new_n2616_), .B(_abc_40319_new_n767_), .C(_abc_40319_new_n694_), .Y(_abc_40319_new_n2617_));
AOI21X1 AOI21X1_153 ( .A(_abc_40319_new_n2524_), .B(_abc_40319_new_n2610_), .C(_abc_40319_new_n2619_), .Y(_abc_40319_new_n2620_));
AOI21X1 AOI21X1_154 ( .A(_abc_40319_new_n2539_), .B(ADDR_REG_5_), .C(_abc_40319_new_n1689_), .Y(_abc_40319_new_n2621_));
AOI21X1 AOI21X1_155 ( .A(_abc_40319_new_n2624_), .B(_abc_40319_new_n2625_), .C(_abc_40319_new_n2626_), .Y(_abc_40319_new_n2627_));
AOI21X1 AOI21X1_156 ( .A(_abc_40319_new_n2631_), .B(_abc_40319_new_n2632_), .C(_abc_40319_new_n2525_), .Y(_abc_40319_new_n2633_));
AOI21X1 AOI21X1_157 ( .A(_abc_40319_new_n2539_), .B(ADDR_REG_6_), .C(_abc_40319_new_n1837_), .Y(_abc_40319_new_n2637_));
AOI21X1 AOI21X1_158 ( .A(_abc_40319_new_n2641_), .B(_abc_40319_new_n2645_), .C(_abc_40319_new_n2644_), .Y(_abc_40319_new_n2646_));
AOI21X1 AOI21X1_159 ( .A(_abc_40319_new_n2539_), .B(ADDR_REG_7_), .C(_abc_40319_new_n1012_), .Y(_abc_40319_new_n2661_));
AOI21X1 AOI21X1_16 ( .A(_abc_40319_new_n961_), .B(_abc_40319_new_n958_), .C(_abc_40319_new_n955_), .Y(_abc_40319_new_n962_));
AOI21X1 AOI21X1_160 ( .A(_abc_40319_new_n2684_), .B(_abc_40319_new_n1273_), .C(_abc_40319_new_n1616_), .Y(_abc_40319_new_n2685_));
AOI21X1 AOI21X1_161 ( .A(_abc_40319_new_n2687_), .B(_abc_40319_new_n2679_), .C(_abc_40319_new_n2691_), .Y(_abc_40319_new_n2692_));
AOI21X1 AOI21X1_162 ( .A(ADDR_REG_10_), .B(_abc_40319_new_n2539_), .C(_abc_40319_new_n2722_), .Y(_abc_40319_new_n2723_));
AOI21X1 AOI21X1_163 ( .A(_abc_40319_new_n2724_), .B(_abc_40319_new_n2726_), .C(_abc_40319_new_n2728_), .Y(_abc_40319_new_n2729_));
AOI21X1 AOI21X1_164 ( .A(_abc_40319_new_n2687_), .B(_abc_40319_new_n2720_), .C(_abc_40319_new_n2735_), .Y(_abc_40319_new_n2736_));
AOI21X1 AOI21X1_165 ( .A(_abc_40319_new_n2754_), .B(_abc_40319_new_n2733_), .C(_abc_40319_new_n2758_), .Y(_abc_40319_new_n2759_));
AOI21X1 AOI21X1_166 ( .A(_abc_40319_new_n2776_), .B(_abc_40319_new_n2733_), .C(_abc_40319_new_n2780_), .Y(_abc_40319_new_n2781_));
AOI21X1 AOI21X1_167 ( .A(_abc_40319_new_n2783_), .B(_abc_40319_new_n2762_), .C(_abc_40319_new_n1326_), .Y(_abc_40319_new_n2785_));
AOI21X1 AOI21X1_168 ( .A(_abc_40319_new_n2794_), .B(_abc_40319_new_n2791_), .C(_abc_40319_new_n2732_), .Y(_abc_40319_new_n2795_));
AOI21X1 AOI21X1_169 ( .A(_abc_40319_new_n2543_), .B(_abc_40319_new_n2797_), .C(_abc_40319_new_n1776_), .Y(_abc_40319_new_n2799_));
AOI21X1 AOI21X1_17 ( .A(_abc_40319_new_n937_), .B(_abc_40319_new_n963_), .C(_abc_40319_new_n962_), .Y(_abc_40319_new_n969_));
AOI21X1 AOI21X1_170 ( .A(_abc_40319_new_n1322_), .B(_abc_40319_new_n2784_), .C(_abc_40319_new_n2785_), .Y(_abc_40319_new_n2803_));
AOI21X1 AOI21X1_171 ( .A(_abc_40319_new_n2806_), .B(_abc_40319_new_n2804_), .C(_abc_40319_new_n1246_), .Y(_abc_40319_new_n2807_));
AOI21X1 AOI21X1_172 ( .A(ADDR_REG_14_), .B(_abc_40319_new_n2539_), .C(_abc_40319_new_n2821_), .Y(_abc_40319_new_n2822_));
AOI21X1 AOI21X1_173 ( .A(_abc_40319_new_n2825_), .B(_abc_40319_new_n2543_), .C(_abc_40319_new_n2823_), .Y(_abc_40319_new_n2826_));
AOI21X1 AOI21X1_174 ( .A(_abc_40319_new_n2806_), .B(_abc_40319_new_n1246_), .C(_abc_40319_new_n2808_), .Y(_abc_40319_new_n2830_));
AOI21X1 AOI21X1_175 ( .A(ADDR_REG_15_), .B(_abc_40319_new_n2539_), .C(_abc_40319_new_n2848_), .Y(_abc_40319_new_n2849_));
AOI21X1 AOI21X1_176 ( .A(_abc_40319_new_n2846_), .B(_abc_40319_new_n2543_), .C(_abc_40319_new_n2850_), .Y(_abc_40319_new_n2851_));
AOI21X1 AOI21X1_177 ( .A(_abc_40319_new_n2875_), .B(_abc_40319_new_n2543_), .C(_abc_40319_new_n2873_), .Y(_abc_40319_new_n2876_));
AOI21X1 AOI21X1_178 ( .A(_abc_40319_new_n2539_), .B(ADDR_REG_17_), .C(_abc_40319_new_n1702_), .Y(_abc_40319_new_n2894_));
AOI21X1 AOI21X1_179 ( .A(_abc_40319_new_n2890_), .B(_abc_40319_new_n2688_), .C(_abc_40319_new_n2895_), .Y(_abc_40319_new_n2896_));
AOI21X1 AOI21X1_18 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n698_), .C(_abc_40319_new_n1012_), .Y(_abc_40319_new_n1013_));
AOI21X1 AOI21X1_180 ( .A(_abc_40319_new_n2907_), .B(_abc_40319_new_n2913_), .C(_abc_40319_new_n694_), .Y(_abc_40319_new_n2914_));
AOI21X1 AOI21X1_181 ( .A(_abc_40319_new_n2920_), .B(_abc_40319_new_n2922_), .C(_abc_40319_new_n2923_), .Y(_abc_40319_new_n2924_));
AOI21X1 AOI21X1_182 ( .A(_abc_40319_new_n2542_), .B(_abc_40319_new_n2926_), .C(_abc_40319_new_n1825_), .Y(_abc_40319_new_n2927_));
AOI21X1 AOI21X1_183 ( .A(_abc_40319_new_n2934_), .B(_abc_40319_new_n2937_), .C(_abc_40319_new_n694_), .Y(_abc_40319_new_n2938_));
AOI21X1 AOI21X1_184 ( .A(_abc_40319_new_n2922_), .B(_abc_40319_new_n2919_), .C(_abc_40319_new_n2941_), .Y(_abc_40319_new_n2942_));
AOI21X1 AOI21X1_185 ( .A(_abc_40319_new_n2939_), .B(_abc_40319_new_n667_), .C(_abc_40319_new_n2943_), .Y(_abc_40319_new_n2944_));
AOI21X1 AOI21X1_186 ( .A(_abc_40319_new_n2684_), .B(_abc_40319_new_n667_), .C(_abc_40319_new_n1571_), .Y(_abc_40319_new_n2952_));
AOI21X1 AOI21X1_187 ( .A(B_REG), .B(_abc_40319_new_n694_), .C(_abc_40319_new_n2985_), .Y(_abc_40319_new_n2986_));
AOI21X1 AOI21X1_188 ( .A(_abc_40319_new_n1570_), .B(_abc_40319_new_n1759_), .C(_abc_40319_new_n3009_), .Y(_abc_40319_new_n3010_));
AOI21X1 AOI21X1_189 ( .A(_abc_40319_new_n1654_), .B(_abc_40319_new_n1796_), .C(_abc_40319_new_n2227_), .Y(_abc_40319_new_n3031_));
AOI21X1 AOI21X1_19 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n990_), .C(_abc_40319_new_n1014_), .Y(_abc_40319_new_n1015_));
AOI21X1 AOI21X1_190 ( .A(_abc_40319_new_n1352_), .B(_abc_40319_new_n1360_), .C(_abc_40319_new_n2229_), .Y(_abc_40319_new_n3034_));
AOI21X1 AOI21X1_191 ( .A(_abc_40319_new_n1726_), .B(_abc_40319_new_n1556_), .C(_abc_40319_new_n3040_), .Y(_abc_40319_new_n3041_));
AOI21X1 AOI21X1_192 ( .A(_abc_40319_new_n3041_), .B(_abc_40319_new_n3048_), .C(_abc_40319_new_n3051_), .Y(_abc_40319_new_n3052_));
AOI21X1 AOI21X1_193 ( .A(_abc_40319_new_n959_), .B(_abc_40319_new_n2246_), .C(_abc_40319_new_n2187_), .Y(_abc_40319_new_n3065_));
AOI21X1 AOI21X1_194 ( .A(_abc_40319_new_n3069_), .B(_abc_40319_new_n3030_), .C(_abc_40319_new_n2240_), .Y(_abc_40319_new_n3070_));
AOI21X1 AOI21X1_195 ( .A(_abc_40319_new_n1122_), .B(_abc_40319_new_n1137_), .C(_abc_40319_new_n3074_), .Y(_abc_40319_new_n3075_));
AOI21X1 AOI21X1_196 ( .A(_abc_40319_new_n3092_), .B(_abc_40319_new_n3079_), .C(_abc_40319_new_n3086_), .Y(_abc_40319_new_n3093_));
AOI21X1 AOI21X1_197 ( .A(_abc_40319_new_n3004_), .B(_abc_40319_new_n3005_), .C(_abc_40319_new_n3105_), .Y(_abc_40319_new_n3106_));
AOI21X1 AOI21X1_198 ( .A(_abc_40319_new_n1601_), .B(_abc_40319_new_n1008_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3112_));
AOI21X1 AOI21X1_199 ( .A(_abc_40319_new_n3111_), .B(_abc_40319_new_n2996_), .C(_abc_40319_new_n3113_), .Y(_abc_40319_new_n3114_));
AOI21X1 AOI21X1_2 ( .A(_abc_40319_new_n587_), .B(_abc_40319_new_n591_), .C(_abc_40319_new_n568_), .Y(_abc_40319_new_n592_));
AOI21X1 AOI21X1_20 ( .A(REG0_REG_27_), .B(_abc_40319_new_n724_), .C(_abc_40319_new_n1044_), .Y(_abc_40319_new_n1045_));
AOI21X1 AOI21X1_200 ( .A(_abc_40319_new_n2264_), .B(_abc_40319_new_n3108_), .C(_abc_40319_new_n3115_), .Y(_abc_40319_new_n3116_));
AOI21X1 AOI21X1_201 ( .A(_abc_40319_new_n3125_), .B(_abc_40319_new_n3101_), .C(_abc_40319_new_n3130_), .Y(_abc_40319_new_n3131_));
AOI21X1 AOI21X1_202 ( .A(_abc_40319_new_n1018_), .B(_abc_40319_new_n2991_), .C(_abc_40319_new_n3138_), .Y(_abc_40319_new_n3139_));
AOI21X1 AOI21X1_203 ( .A(_abc_40319_new_n1580_), .B(_abc_40319_new_n3108_), .C(_abc_40319_new_n3140_), .Y(_abc_40319_new_n3141_));
AOI21X1 AOI21X1_204 ( .A(_abc_40319_new_n3154_), .B(_abc_40319_new_n3101_), .C(_abc_40319_new_n3157_), .Y(_abc_40319_new_n3158_));
AOI21X1 AOI21X1_205 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1852_), .C(_abc_40319_new_n3167_), .Y(_abc_40319_new_n3168_));
AOI21X1 AOI21X1_206 ( .A(_abc_40319_new_n3163_), .B(_abc_40319_new_n2996_), .C(_abc_40319_new_n3169_), .Y(_abc_40319_new_n3170_));
AOI21X1 AOI21X1_207 ( .A(_abc_40319_new_n3180_), .B(_abc_40319_new_n2320_), .C(_abc_40319_new_n2410_), .Y(_abc_40319_new_n3181_));
AOI21X1 AOI21X1_208 ( .A(_abc_40319_new_n3101_), .B(_abc_40319_new_n3177_), .C(_abc_40319_new_n3187_), .Y(_abc_40319_new_n3188_));
AOI21X1 AOI21X1_209 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n3192_), .C(_abc_40319_new_n3196_), .Y(_abc_40319_new_n3197_));
AOI21X1 AOI21X1_21 ( .A(REG2_REG_26_), .B(_abc_40319_new_n715_), .C(_abc_40319_new_n1063_), .Y(_abc_40319_new_n1064_));
AOI21X1 AOI21X1_210 ( .A(_abc_40319_new_n3191_), .B(_abc_40319_new_n2996_), .C(_abc_40319_new_n3198_), .Y(_abc_40319_new_n3199_));
AOI21X1 AOI21X1_211 ( .A(_abc_40319_new_n1115_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3208_), .Y(_abc_40319_new_n3209_));
AOI21X1 AOI21X1_212 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1714_), .C(_abc_40319_new_n3216_), .Y(_abc_40319_new_n3217_));
AOI21X1 AOI21X1_213 ( .A(_abc_40319_new_n3213_), .B(_abc_40319_new_n2996_), .C(_abc_40319_new_n3218_), .Y(_abc_40319_new_n3219_));
AOI21X1 AOI21X1_214 ( .A(_abc_40319_new_n2498_), .B(_abc_40319_new_n2500_), .C(_abc_40319_new_n2458_), .Y(_abc_40319_new_n3230_));
AOI21X1 AOI21X1_215 ( .A(_abc_40319_new_n3230_), .B(_abc_40319_new_n2140_), .C(_abc_40319_new_n2142_), .Y(_abc_40319_new_n3231_));
AOI21X1 AOI21X1_216 ( .A(_abc_40319_new_n3237_), .B(_abc_40319_new_n3005_), .C(_abc_40319_new_n3239_), .Y(_abc_40319_new_n3240_));
AOI21X1 AOI21X1_217 ( .A(_abc_40319_new_n3240_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3241_), .Y(_abc_40319_new_n3242_));
AOI21X1 AOI21X1_218 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3229_), .C(_abc_40319_new_n3242_), .Y(_abc_40319_new_n3243_));
AOI21X1 AOI21X1_219 ( .A(_abc_40319_new_n3071_), .B(_abc_40319_new_n3073_), .C(_abc_40319_new_n3022_), .Y(_abc_40319_new_n3253_));
AOI21X1 AOI21X1_22 ( .A(REG1_REG_25_), .B(_abc_40319_new_n726_), .C(_abc_40319_new_n1075_), .Y(_abc_40319_new_n1076_));
AOI21X1 AOI21X1_220 ( .A(_abc_40319_new_n3005_), .B(_abc_40319_new_n3257_), .C(_abc_40319_new_n3259_), .Y(_abc_40319_new_n3260_));
AOI21X1 AOI21X1_221 ( .A(_abc_40319_new_n3265_), .B(_abc_40319_new_n3230_), .C(_abc_40319_new_n3270_), .Y(_abc_40319_new_n3271_));
AOI21X1 AOI21X1_222 ( .A(_abc_40319_new_n1452_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3271_), .Y(_abc_40319_new_n3272_));
AOI21X1 AOI21X1_223 ( .A(_abc_40319_new_n2960_), .B(_abc_40319_new_n3279_), .C(_abc_40319_new_n3278_), .Y(_abc_40319_new_n3280_));
AOI21X1 AOI21X1_224 ( .A(_abc_40319_new_n3277_), .B(_abc_40319_new_n2996_), .C(_abc_40319_new_n3281_), .Y(_abc_40319_new_n3282_));
AOI21X1 AOI21X1_225 ( .A(_abc_40319_new_n3291_), .B(_abc_40319_new_n2220_), .C(_abc_40319_new_n3155_), .Y(_abc_40319_new_n3292_));
AOI21X1 AOI21X1_226 ( .A(_abc_40319_new_n2960_), .B(_abc_40319_new_n3302_), .C(_abc_40319_new_n3303_), .Y(_abc_40319_new_n3304_));
AOI21X1 AOI21X1_227 ( .A(_abc_40319_new_n1469_), .B(_abc_40319_new_n3108_), .C(_abc_40319_new_n3305_), .Y(_abc_40319_new_n3306_));
AOI21X1 AOI21X1_228 ( .A(_abc_40319_new_n2170_), .B(_abc_40319_new_n2498_), .C(_abc_40319_new_n3309_), .Y(_abc_40319_new_n3310_));
AOI21X1 AOI21X1_229 ( .A(_abc_40319_new_n3308_), .B(_abc_40319_new_n3101_), .C(_abc_40319_new_n3310_), .Y(_abc_40319_new_n3311_));
AOI21X1 AOI21X1_23 ( .A(REG1_REG_24_), .B(_abc_40319_new_n726_), .C(_abc_40319_new_n1091_), .Y(_abc_40319_new_n1092_));
AOI21X1 AOI21X1_230 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1432_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3318_));
AOI21X1 AOI21X1_231 ( .A(REG2_REG_19_), .B(_abc_40319_new_n2990_), .C(_abc_40319_new_n3319_), .Y(_abc_40319_new_n3320_));
AOI21X1 AOI21X1_232 ( .A(_abc_40319_new_n3315_), .B(_abc_40319_new_n2996_), .C(_abc_40319_new_n3321_), .Y(_abc_40319_new_n3322_));
AOI21X1 AOI21X1_233 ( .A(_abc_40319_new_n3325_), .B(_abc_40319_new_n2164_), .C(_abc_40319_new_n3155_), .Y(_abc_40319_new_n3326_));
AOI21X1 AOI21X1_234 ( .A(_abc_40319_new_n3324_), .B(_abc_40319_new_n3101_), .C(_abc_40319_new_n3328_), .Y(_abc_40319_new_n3329_));
AOI21X1 AOI21X1_235 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1824_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3335_));
AOI21X1 AOI21X1_236 ( .A(REG2_REG_18_), .B(_abc_40319_new_n2990_), .C(_abc_40319_new_n3336_), .Y(_abc_40319_new_n3337_));
AOI21X1 AOI21X1_237 ( .A(_abc_40319_new_n3334_), .B(_abc_40319_new_n2996_), .C(_abc_40319_new_n3338_), .Y(_abc_40319_new_n3339_));
AOI21X1 AOI21X1_238 ( .A(_abc_40319_new_n3071_), .B(_abc_40319_new_n2197_), .C(_abc_40319_new_n3020_), .Y(_abc_40319_new_n3343_));
AOI21X1 AOI21X1_239 ( .A(_abc_40319_new_n3359_), .B(_abc_40319_new_n2484_), .C(_abc_40319_new_n3346_), .Y(_abc_40319_new_n3360_));
AOI21X1 AOI21X1_24 ( .A(REG0_REG_23_), .B(_abc_40319_new_n724_), .C(_abc_40319_new_n1113_), .Y(_abc_40319_new_n1114_));
AOI21X1 AOI21X1_240 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1205_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3370_));
AOI21X1 AOI21X1_241 ( .A(_abc_40319_new_n2991_), .B(_abc_40319_new_n1198_), .C(_abc_40319_new_n3371_), .Y(_abc_40319_new_n3372_));
AOI21X1 AOI21X1_242 ( .A(_abc_40319_new_n3367_), .B(_abc_40319_new_n2996_), .C(_abc_40319_new_n3373_), .Y(_abc_40319_new_n3374_));
AOI21X1 AOI21X1_243 ( .A(_abc_40319_new_n3383_), .B(_abc_40319_new_n2223_), .C(_abc_40319_new_n2330_), .Y(_abc_40319_new_n3384_));
AOI21X1 AOI21X1_244 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1255_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3420_));
AOI21X1 AOI21X1_245 ( .A(_abc_40319_new_n3417_), .B(_abc_40319_new_n2996_), .C(_abc_40319_new_n3422_), .Y(_abc_40319_new_n3423_));
AOI21X1 AOI21X1_246 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1330_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3442_));
AOI21X1 AOI21X1_247 ( .A(_abc_40319_new_n3431_), .B(_abc_40319_new_n3133_), .C(_abc_40319_new_n3443_), .Y(_abc_40319_new_n3444_));
AOI21X1 AOI21X1_248 ( .A(_abc_40319_new_n3469_), .B(_abc_40319_new_n3005_), .C(_abc_40319_new_n3471_), .Y(_abc_40319_new_n3472_));
AOI21X1 AOI21X1_249 ( .A(_abc_40319_new_n3053_), .B(_abc_40319_new_n3065_), .C(_abc_40319_new_n3061_), .Y(_abc_40319_new_n3477_));
AOI21X1 AOI21X1_25 ( .A(_abc_40319_new_n1204_), .B(_abc_40319_new_n1203_), .C(_abc_40319_new_n1031_), .Y(_abc_40319_new_n1205_));
AOI21X1 AOI21X1_250 ( .A(_abc_40319_new_n2990_), .B(REG2_REG_10_), .C(_abc_40319_new_n3487_), .Y(_abc_40319_new_n3488_));
AOI21X1 AOI21X1_251 ( .A(_abc_40319_new_n3481_), .B(_abc_40319_new_n3133_), .C(_abc_40319_new_n3493_), .Y(_abc_40319_new_n3494_));
AOI21X1 AOI21X1_252 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1302_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3506_));
AOI21X1 AOI21X1_253 ( .A(_abc_40319_new_n2960_), .B(_abc_40319_new_n3505_), .C(_abc_40319_new_n3507_), .Y(_abc_40319_new_n3508_));
AOI21X1 AOI21X1_254 ( .A(_abc_40319_new_n3498_), .B(_abc_40319_new_n3133_), .C(_abc_40319_new_n3509_), .Y(_abc_40319_new_n3510_));
AOI21X1 AOI21X1_255 ( .A(_abc_40319_new_n3005_), .B(_abc_40319_new_n3513_), .C(_abc_40319_new_n3516_), .Y(_abc_40319_new_n3517_));
AOI21X1 AOI21X1_256 ( .A(_abc_40319_new_n2990_), .B(REG2_REG_8_), .C(_abc_40319_new_n3523_), .Y(_abc_40319_new_n3524_));
AOI21X1 AOI21X1_257 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3514_), .C(_abc_40319_new_n3525_), .Y(_abc_40319_new_n3526_));
AOI21X1 AOI21X1_258 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n738_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3542_));
AOI21X1 AOI21X1_259 ( .A(_abc_40319_new_n3532_), .B(_abc_40319_new_n3133_), .C(_abc_40319_new_n3543_), .Y(_abc_40319_new_n3544_));
AOI21X1 AOI21X1_26 ( .A(_abc_40319_new_n1228_), .B(_abc_40319_new_n1229_), .C(_abc_40319_new_n1182_), .Y(_abc_40319_new_n1230_));
AOI21X1 AOI21X1_260 ( .A(_abc_40319_new_n3549_), .B(_abc_40319_new_n3005_), .C(_abc_40319_new_n3551_), .Y(_abc_40319_new_n3552_));
AOI21X1 AOI21X1_261 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n948_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3559_));
AOI21X1 AOI21X1_262 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3553_), .C(_abc_40319_new_n3560_), .Y(_abc_40319_new_n3561_));
AOI21X1 AOI21X1_263 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n806_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3574_));
AOI21X1 AOI21X1_264 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3567_), .C(_abc_40319_new_n3575_), .Y(_abc_40319_new_n3576_));
AOI21X1 AOI21X1_265 ( .A(REG2_REG_4_), .B(_abc_40319_new_n2990_), .C(_abc_40319_new_n3577_), .Y(_abc_40319_new_n3578_));
AOI21X1 AOI21X1_266 ( .A(_abc_40319_new_n3005_), .B(_abc_40319_new_n3580_), .C(_abc_40319_new_n3584_), .Y(_abc_40319_new_n3585_));
AOI21X1 AOI21X1_267 ( .A(_abc_40319_new_n2960_), .B(_abc_40319_new_n3589_), .C(_abc_40319_new_n3590_), .Y(_abc_40319_new_n3591_));
AOI21X1 AOI21X1_268 ( .A(REG2_REG_5_), .B(_abc_40319_new_n2990_), .C(_abc_40319_new_n3593_), .Y(_abc_40319_new_n3594_));
AOI21X1 AOI21X1_269 ( .A(_abc_40319_new_n2470_), .B(_abc_40319_new_n2155_), .C(_abc_40319_new_n3155_), .Y(_abc_40319_new_n3596_));
AOI21X1 AOI21X1_27 ( .A(_abc_40319_new_n1277_), .B(_abc_40319_new_n1279_), .C(_abc_40319_new_n1280_), .Y(_abc_40319_new_n1281_));
AOI21X1 AOI21X1_270 ( .A(_abc_40319_new_n2990_), .B(REG2_REG_3_), .C(_abc_40319_new_n3607_), .Y(_abc_40319_new_n3608_));
AOI21X1 AOI21X1_271 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3600_), .C(_abc_40319_new_n3609_), .Y(_abc_40319_new_n3610_));
AOI21X1 AOI21X1_272 ( .A(_abc_40319_new_n3613_), .B(_abc_40319_new_n2245_), .C(_abc_40319_new_n3155_), .Y(_abc_40319_new_n3614_));
AOI21X1 AOI21X1_273 ( .A(_abc_40319_new_n880_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3616_), .Y(_abc_40319_new_n3617_));
AOI21X1 AOI21X1_274 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n2962_), .C(_abc_40319_new_n3621_), .Y(_abc_40319_new_n3622_));
AOI21X1 AOI21X1_275 ( .A(_abc_40319_new_n1008_), .B(REG3_REG_2_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3625_));
AOI21X1 AOI21X1_276 ( .A(_abc_40319_new_n3624_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3626_), .Y(_abc_40319_new_n3627_));
AOI21X1 AOI21X1_277 ( .A(_abc_40319_new_n3631_), .B(_abc_40319_new_n1905_), .C(_abc_40319_new_n3155_), .Y(_abc_40319_new_n3632_));
AOI21X1 AOI21X1_278 ( .A(_abc_40319_new_n2990_), .B(REG2_REG_1_), .C(_abc_40319_new_n3641_), .Y(_abc_40319_new_n3642_));
AOI21X1 AOI21X1_279 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n2237_), .C(_abc_40319_new_n3650_), .Y(_abc_40319_new_n3651_));
AOI21X1 AOI21X1_28 ( .A(_abc_40319_new_n1282_), .B(_abc_40319_new_n1288_), .C(_abc_40319_new_n1312_), .Y(_abc_40319_new_n1313_));
AOI21X1 AOI21X1_280 ( .A(n1336), .B(DATAI_31_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3655_));
AOI21X1 AOI21X1_281 ( .A(_abc_40319_new_n772_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3724_));
AOI21X1 AOI21X1_282 ( .A(_abc_40319_new_n3720_), .B(IR_REG_26_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3734_));
AOI21X1 AOI21X1_283 ( .A(_abc_40319_new_n3720_), .B(IR_REG_25_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3738_));
AOI21X1 AOI21X1_284 ( .A(_abc_40319_new_n3720_), .B(IR_REG_24_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3743_));
AOI21X1 AOI21X1_285 ( .A(n1336), .B(DATAI_23_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3747_));
AOI21X1 AOI21X1_286 ( .A(_abc_40319_new_n3720_), .B(IR_REG_22_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3749_));
AOI21X1 AOI21X1_287 ( .A(_abc_40319_new_n613_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3754_));
AOI21X1 AOI21X1_288 ( .A(_abc_40319_new_n3720_), .B(IR_REG_20_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3756_));
AOI21X1 AOI21X1_289 ( .A(_abc_40319_new_n1144_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3764_));
AOI21X1 AOI21X1_29 ( .A(_abc_40319_new_n1314_), .B(_abc_40319_new_n1316_), .C(_abc_40319_new_n1313_), .Y(_abc_40319_new_n1317_));
AOI21X1 AOI21X1_290 ( .A(_abc_40319_new_n3770_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3771_));
AOI21X1 AOI21X1_291 ( .A(_abc_40319_new_n1242_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3777_));
AOI21X1 AOI21X1_292 ( .A(_abc_40319_new_n1292_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3794_));
AOI21X1 AOI21X1_293 ( .A(_abc_40319_new_n1270_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3797_));
AOI21X1 AOI21X1_294 ( .A(_abc_40319_new_n688_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3800_));
AOI21X1 AOI21X1_295 ( .A(_abc_40319_new_n940_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3803_));
AOI21X1 AOI21X1_296 ( .A(_abc_40319_new_n794_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3809_));
AOI21X1 AOI21X1_297 ( .A(_abc_40319_new_n3720_), .B(IR_REG_3_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3811_));
AOI21X1 AOI21X1_298 ( .A(n1336), .B(DATAI_1_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3819_));
AOI21X1 AOI21X1_299 ( .A(IR_REG_0_), .B(STATE_REG), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3821_));
AOI21X1 AOI21X1_3 ( .A(_abc_40319_new_n601_), .B(_abc_40319_new_n600_), .C(_abc_40319_new_n568_), .Y(_abc_40319_new_n602_));
AOI21X1 AOI21X1_30 ( .A(_abc_40319_new_n1488_), .B(_abc_40319_new_n1120_), .C(_abc_40319_new_n1491_), .Y(_abc_40319_new_n1492_));
AOI21X1 AOI21X1_300 ( .A(_abc_40319_new_n3844_), .B(_abc_40319_new_n3101_), .C(_abc_40319_new_n3850_), .Y(_abc_40319_new_n3851_));
AOI21X1 AOI21X1_301 ( .A(_abc_40319_new_n2960_), .B(_abc_40319_new_n3871_), .C(_abc_40319_new_n3872_), .Y(_abc_40319_new_n3873_));
AOI21X1 AOI21X1_302 ( .A(_abc_40319_new_n3857_), .B(_abc_40319_new_n2996_), .C(_abc_40319_new_n3874_), .Y(_abc_40319_new_n3875_));
AOI21X1 AOI21X1_303 ( .A(_abc_40319_new_n3878_), .B(_abc_40319_new_n629_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3883_));
AOI21X1 AOI21X1_304 ( .A(_abc_40319_new_n3287_), .B(_abc_40319_new_n3893_), .C(_abc_40319_new_n3302_), .Y(_abc_40319_new_n3894_));
AOI21X1 AOI21X1_305 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_20_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3898_));
AOI21X1 AOI21X1_306 ( .A(_abc_40319_new_n3907_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3908_));
AOI21X1 AOI21X1_307 ( .A(_abc_40319_new_n3911_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3912_));
AOI21X1 AOI21X1_308 ( .A(_abc_40319_new_n3600_), .B(_abc_40319_new_n3893_), .C(_abc_40319_new_n3603_), .Y(_abc_40319_new_n3915_));
AOI21X1 AOI21X1_309 ( .A(_abc_40319_new_n3917_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3918_));
AOI21X1 AOI21X1_31 ( .A(_abc_40319_new_n1498_), .B(_abc_40319_new_n1497_), .C(_abc_40319_new_n778_), .Y(_abc_40319_new_n1499_));
AOI21X1 AOI21X1_310 ( .A(_abc_40319_new_n3620_), .B(_abc_40319_new_n3571_), .C(_abc_40319_new_n3569_), .Y(_abc_40319_new_n3921_));
AOI21X1 AOI21X1_311 ( .A(_abc_40319_new_n3922_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3923_));
AOI21X1 AOI21X1_312 ( .A(_abc_40319_new_n3587_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n3589_), .Y(_abc_40319_new_n3926_));
AOI21X1 AOI21X1_313 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_5_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3929_));
AOI21X1 AOI21X1_314 ( .A(_abc_40319_new_n3554_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n3557_), .Y(_abc_40319_new_n3931_));
AOI21X1 AOI21X1_315 ( .A(_abc_40319_new_n3933_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3934_));
AOI21X1 AOI21X1_316 ( .A(_abc_40319_new_n3532_), .B(_abc_40319_new_n3893_), .C(_abc_40319_new_n3938_), .Y(_abc_40319_new_n3939_));
AOI21X1 AOI21X1_317 ( .A(_abc_40319_new_n3940_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3941_));
AOI21X1 AOI21X1_318 ( .A(_abc_40319_new_n3518_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n3520_), .Y(_abc_40319_new_n3944_));
AOI21X1 AOI21X1_319 ( .A(_abc_40319_new_n3514_), .B(_abc_40319_new_n3893_), .C(_abc_40319_new_n3521_), .Y(_abc_40319_new_n3945_));
AOI21X1 AOI21X1_32 ( .A(REG0_REG_28_), .B(_abc_40319_new_n724_), .C(_abc_40319_new_n1502_), .Y(_abc_40319_new_n1503_));
AOI21X1 AOI21X1_320 ( .A(_abc_40319_new_n3946_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3947_));
AOI21X1 AOI21X1_321 ( .A(_abc_40319_new_n3498_), .B(_abc_40319_new_n3893_), .C(_abc_40319_new_n3950_), .Y(_abc_40319_new_n3951_));
AOI21X1 AOI21X1_322 ( .A(_abc_40319_new_n3952_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3953_));
AOI21X1 AOI21X1_323 ( .A(_abc_40319_new_n3485_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n3489_), .Y(_abc_40319_new_n3955_));
AOI21X1 AOI21X1_324 ( .A(_abc_40319_new_n3481_), .B(_abc_40319_new_n3893_), .C(_abc_40319_new_n3491_), .Y(_abc_40319_new_n3956_));
AOI21X1 AOI21X1_325 ( .A(_abc_40319_new_n3957_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3958_));
AOI21X1 AOI21X1_326 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_11_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3965_));
AOI21X1 AOI21X1_327 ( .A(_abc_40319_new_n3969_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3970_));
AOI21X1 AOI21X1_328 ( .A(_abc_40319_new_n3436_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n3438_), .Y(_abc_40319_new_n3972_));
AOI21X1 AOI21X1_329 ( .A(_abc_40319_new_n3974_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3975_));
AOI21X1 AOI21X1_33 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n1018_), .C(_abc_40319_new_n1507_), .Y(_abc_40319_new_n1508_));
AOI21X1 AOI21X1_330 ( .A(_abc_40319_new_n3893_), .B(_abc_40319_new_n3410_), .C(_abc_40319_new_n3412_), .Y(_abc_40319_new_n3978_));
AOI21X1 AOI21X1_331 ( .A(_abc_40319_new_n3979_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3980_));
AOI21X1 AOI21X1_332 ( .A(_abc_40319_new_n3379_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n3988_), .Y(_abc_40319_new_n3989_));
AOI21X1 AOI21X1_333 ( .A(_abc_40319_new_n3367_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n3995_), .Y(_abc_40319_new_n3996_));
AOI21X1 AOI21X1_334 ( .A(_abc_40319_new_n3998_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n3999_));
AOI21X1 AOI21X1_335 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_18_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4005_));
AOI21X1 AOI21X1_336 ( .A(_abc_40319_new_n3315_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n3316_), .Y(_abc_40319_new_n4007_));
AOI21X1 AOI21X1_337 ( .A(_abc_40319_new_n3277_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n4014_), .Y(_abc_40319_new_n4015_));
AOI21X1 AOI21X1_338 ( .A(_abc_40319_new_n1115_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n4022_), .Y(_abc_40319_new_n4023_));
AOI21X1 AOI21X1_339 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_22_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4026_));
AOI21X1 AOI21X1_34 ( .A(_abc_40319_new_n1506_), .B(_abc_40319_new_n976_), .C(_abc_40319_new_n1509_), .Y(_abc_40319_new_n1510_));
AOI21X1 AOI21X1_340 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_23_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4032_));
AOI21X1 AOI21X1_341 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_24_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4038_));
AOI21X1 AOI21X1_342 ( .A(_abc_40319_new_n3191_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n3194_), .Y(_abc_40319_new_n4040_));
AOI21X1 AOI21X1_343 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_25_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4044_));
AOI21X1 AOI21X1_344 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_26_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4050_));
AOI21X1 AOI21X1_345 ( .A(_abc_40319_new_n3123_), .B(_abc_40319_new_n3124_), .C(_abc_40319_new_n1005_), .Y(_abc_40319_new_n4054_));
AOI21X1 AOI21X1_346 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_27_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4059_));
AOI21X1 AOI21X1_347 ( .A(_abc_40319_new_n2264_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n4062_), .Y(_abc_40319_new_n4063_));
AOI21X1 AOI21X1_348 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_28_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4066_));
AOI21X1 AOI21X1_349 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_29_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4073_));
AOI21X1 AOI21X1_35 ( .A(n1336), .B(REG3_REG_14_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n1520_));
AOI21X1 AOI21X1_350 ( .A(_abc_40319_new_n2997_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n4075_), .Y(_abc_40319_new_n4076_));
AOI21X1 AOI21X1_351 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_30_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4077_));
AOI21X1 AOI21X1_352 ( .A(_abc_40319_new_n2981_), .B(_abc_40319_new_n2983_), .C(_abc_40319_new_n3891_), .Y(_abc_40319_new_n4079_));
AOI21X1 AOI21X1_353 ( .A(_abc_40319_new_n3890_), .B(REG0_REG_31_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4082_));
AOI21X1 AOI21X1_354 ( .A(_abc_40319_new_n3907_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4089_));
AOI21X1 AOI21X1_355 ( .A(_abc_40319_new_n3911_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4092_));
AOI21X1 AOI21X1_356 ( .A(_abc_40319_new_n3917_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4094_));
AOI21X1 AOI21X1_357 ( .A(_abc_40319_new_n3922_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4096_));
AOI21X1 AOI21X1_358 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_5_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4098_));
AOI21X1 AOI21X1_359 ( .A(_abc_40319_new_n3933_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4100_));
AOI21X1 AOI21X1_36 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1255_), .C(_abc_40319_new_n1521_), .Y(_abc_40319_new_n1522_));
AOI21X1 AOI21X1_360 ( .A(_abc_40319_new_n3940_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4102_));
AOI21X1 AOI21X1_361 ( .A(_abc_40319_new_n3946_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4104_));
AOI21X1 AOI21X1_362 ( .A(_abc_40319_new_n3952_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4106_));
AOI21X1 AOI21X1_363 ( .A(_abc_40319_new_n3957_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4108_));
AOI21X1 AOI21X1_364 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_11_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4110_));
AOI21X1 AOI21X1_365 ( .A(_abc_40319_new_n3969_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4112_));
AOI21X1 AOI21X1_366 ( .A(_abc_40319_new_n3974_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4114_));
AOI21X1 AOI21X1_367 ( .A(_abc_40319_new_n3979_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4116_));
AOI21X1 AOI21X1_368 ( .A(_abc_40319_new_n3998_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4124_));
AOI21X1 AOI21X1_369 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_18_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4126_));
AOI21X1 AOI21X1_37 ( .A(_abc_40319_new_n1525_), .B(_abc_40319_new_n1526_), .C(_abc_40319_new_n677_), .Y(_abc_40319_new_n1527_));
AOI21X1 AOI21X1_370 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_20_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4131_));
AOI21X1 AOI21X1_371 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_21_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4134_));
AOI21X1 AOI21X1_372 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_22_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4136_));
AOI21X1 AOI21X1_373 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_23_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4138_));
AOI21X1 AOI21X1_374 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_24_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4140_));
AOI21X1 AOI21X1_375 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_25_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4142_));
AOI21X1 AOI21X1_376 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_26_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4144_));
AOI21X1 AOI21X1_377 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_27_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4146_));
AOI21X1 AOI21X1_378 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_28_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4148_));
AOI21X1 AOI21X1_379 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_29_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4151_));
AOI21X1 AOI21X1_38 ( .A(n1336), .B(REG3_REG_23_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n1532_));
AOI21X1 AOI21X1_380 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_30_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4153_));
AOI21X1 AOI21X1_381 ( .A(_abc_40319_new_n4084_), .B(REG1_REG_31_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4156_));
AOI21X1 AOI21X1_382 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_0_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4159_));
AOI21X1 AOI21X1_383 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_1_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4161_));
AOI21X1 AOI21X1_384 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_2_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4163_));
AOI21X1 AOI21X1_385 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_3_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4165_));
AOI21X1 AOI21X1_386 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_4_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4167_));
AOI21X1 AOI21X1_387 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_5_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4169_));
AOI21X1 AOI21X1_388 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_6_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4171_));
AOI21X1 AOI21X1_389 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_7_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4173_));
AOI21X1 AOI21X1_39 ( .A(n1336), .B(REG3_REG_10_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n1542_));
AOI21X1 AOI21X1_390 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_8_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4175_));
AOI21X1 AOI21X1_391 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_9_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4177_));
AOI21X1 AOI21X1_392 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_10_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4179_));
AOI21X1 AOI21X1_393 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_11_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4181_));
AOI21X1 AOI21X1_394 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_12_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4183_));
AOI21X1 AOI21X1_395 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_13_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4185_));
AOI21X1 AOI21X1_396 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_14_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4187_));
AOI21X1 AOI21X1_397 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_15_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4189_));
AOI21X1 AOI21X1_398 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_16_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4191_));
AOI21X1 AOI21X1_399 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_17_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4193_));
AOI21X1 AOI21X1_4 ( .A(_abc_40319_new_n681_), .B(_abc_40319_new_n682_), .C(_abc_40319_new_n671_), .Y(_abc_40319_new_n683_));
AOI21X1 AOI21X1_40 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1398_), .C(_abc_40319_new_n1543_), .Y(_abc_40319_new_n1544_));
AOI21X1 AOI21X1_400 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_18_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4195_));
AOI21X1 AOI21X1_401 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_19_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4197_));
AOI21X1 AOI21X1_402 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_20_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4199_));
AOI21X1 AOI21X1_403 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_21_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4201_));
AOI21X1 AOI21X1_404 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_22_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4203_));
AOI21X1 AOI21X1_405 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_23_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4205_));
AOI21X1 AOI21X1_406 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_24_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4207_));
AOI21X1 AOI21X1_407 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_25_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4209_));
AOI21X1 AOI21X1_408 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_26_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4211_));
AOI21X1 AOI21X1_409 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_27_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4213_));
AOI21X1 AOI21X1_41 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n826_), .C(_abc_40319_new_n1558_), .Y(_abc_40319_new_n1559_));
AOI21X1 AOI21X1_410 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_28_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4215_));
AOI21X1 AOI21X1_411 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_29_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4217_));
AOI21X1 AOI21X1_412 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_30_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4219_));
AOI21X1 AOI21X1_413 ( .A(_abc_40319_new_n583_), .B(DATAO_REG_31_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n4221_));
AOI21X1 AOI21X1_42 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1557_), .C(_abc_40319_new_n1560_), .Y(_abc_40319_new_n1561_));
AOI21X1 AOI21X1_43 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1432_), .C(_abc_40319_new_n1573_), .Y(_abc_40319_new_n1574_));
AOI21X1 AOI21X1_44 ( .A(REG0_REG_29_), .B(_abc_40319_new_n724_), .C(_abc_40319_new_n1596_), .Y(_abc_40319_new_n1597_));
AOI21X1 AOI21X1_45 ( .A(n1336), .B(REG3_REG_28_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n1602_));
AOI21X1 AOI21X1_46 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1601_), .C(_abc_40319_new_n1603_), .Y(_abc_40319_new_n1604_));
AOI21X1 AOI21X1_47 ( .A(_abc_40319_new_n1611_), .B(_abc_40319_new_n1608_), .C(_abc_40319_new_n677_), .Y(_abc_40319_new_n1612_));
AOI21X1 AOI21X1_48 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n1276_), .C(_abc_40319_new_n1616_), .Y(_abc_40319_new_n1617_));
AOI21X1 AOI21X1_49 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1614_), .C(_abc_40319_new_n1618_), .Y(_abc_40319_new_n1619_));
AOI21X1 AOI21X1_5 ( .A(_abc_40319_new_n695_), .B(IR_REG_31_), .C(_abc_40319_new_n593_), .Y(_abc_40319_new_n696_));
AOI21X1 AOI21X1_50 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n877_), .C(_abc_40319_new_n1625_), .Y(_abc_40319_new_n1626_));
AOI21X1 AOI21X1_51 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1623_), .C(_abc_40319_new_n1627_), .Y(_abc_40319_new_n1628_));
AOI21X1 AOI21X1_52 ( .A(_abc_40319_new_n978_), .B(_abc_40319_new_n1452_), .C(_abc_40319_new_n1630_), .Y(_abc_40319_new_n1631_));
AOI21X1 AOI21X1_53 ( .A(_abc_40319_new_n1634_), .B(_abc_40319_new_n1458_), .C(_abc_40319_new_n1483_), .Y(_abc_40319_new_n1635_));
AOI21X1 AOI21X1_54 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n1460_), .C(_abc_40319_new_n1640_), .Y(_abc_40319_new_n1641_));
AOI21X1 AOI21X1_55 ( .A(_abc_40319_new_n1639_), .B(_abc_40319_new_n1636_), .C(_abc_40319_new_n1642_), .Y(_abc_40319_new_n1643_));
AOI21X1 AOI21X1_56 ( .A(_abc_40319_new_n1647_), .B(_abc_40319_new_n1646_), .C(_abc_40319_new_n1411_), .Y(_abc_40319_new_n1648_));
AOI21X1 AOI21X1_57 ( .A(n1336), .B(REG3_REG_12_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n1655_));
AOI21X1 AOI21X1_58 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1357_), .C(_abc_40319_new_n1656_), .Y(_abc_40319_new_n1657_));
AOI21X1 AOI21X1_59 ( .A(_abc_40319_new_n1662_), .B(_abc_40319_new_n1489_), .C(_abc_40319_new_n1661_), .Y(_abc_40319_new_n1663_));
AOI21X1 AOI21X1_6 ( .A(_abc_40319_new_n716_), .B(_abc_40319_new_n719_), .C(_abc_40319_new_n723_), .Y(_abc_40319_new_n724_));
AOI21X1 AOI21X1_60 ( .A(_abc_40319_new_n1488_), .B(_abc_40319_new_n1120_), .C(_abc_40319_new_n1490_), .Y(_abc_40319_new_n1664_));
AOI21X1 AOI21X1_61 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n1080_), .C(_abc_40319_new_n1668_), .Y(_abc_40319_new_n1669_));
AOI21X1 AOI21X1_62 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1667_), .C(_abc_40319_new_n1670_), .Y(_abc_40319_new_n1671_));
AOI21X1 AOI21X1_63 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n1175_), .C(_abc_40319_new_n1680_), .Y(_abc_40319_new_n1681_));
AOI21X1 AOI21X1_64 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1679_), .C(_abc_40319_new_n1682_), .Y(_abc_40319_new_n1683_));
AOI21X1 AOI21X1_65 ( .A(_abc_40319_new_n1609_), .B(_abc_40319_new_n1685_), .C(_abc_40319_new_n677_), .Y(_abc_40319_new_n1686_));
AOI21X1 AOI21X1_66 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n769_), .C(_abc_40319_new_n1689_), .Y(_abc_40319_new_n1690_));
AOI21X1 AOI21X1_67 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1688_), .C(_abc_40319_new_n1691_), .Y(_abc_40319_new_n1692_));
AOI21X1 AOI21X1_68 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n1198_), .C(_abc_40319_new_n1702_), .Y(_abc_40319_new_n1703_));
AOI21X1 AOI21X1_69 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1701_), .C(_abc_40319_new_n1704_), .Y(_abc_40319_new_n1705_));
AOI21X1 AOI21X1_7 ( .A(_abc_40319_new_n560_), .B(_abc_40319_new_n573_), .C(_abc_40319_new_n681_), .Y(_abc_40319_new_n746_));
AOI21X1 AOI21X1_70 ( .A(_abc_40319_new_n1577_), .B(_abc_40319_new_n1707_), .C(_abc_40319_new_n677_), .Y(_abc_40319_new_n1708_));
AOI21X1 AOI21X1_71 ( .A(n1336), .B(REG3_REG_24_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n1715_));
AOI21X1 AOI21X1_72 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1714_), .C(_abc_40319_new_n1716_), .Y(_abc_40319_new_n1717_));
AOI21X1 AOI21X1_73 ( .A(_abc_40319_new_n1719_), .B(_abc_40319_new_n1720_), .C(_abc_40319_new_n677_), .Y(_abc_40319_new_n1721_));
AOI21X1 AOI21X1_74 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n806_), .C(_abc_40319_new_n1729_), .Y(_abc_40319_new_n1730_));
AOI21X1 AOI21X1_75 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1302_), .C(_abc_40319_new_n1742_), .Y(_abc_40319_new_n1743_));
AOI21X1 AOI21X1_76 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n914_), .C(_abc_40319_new_n1752_), .Y(_abc_40319_new_n1753_));
AOI21X1 AOI21X1_77 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1751_), .C(_abc_40319_new_n1754_), .Y(_abc_40319_new_n1755_));
AOI21X1 AOI21X1_78 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n1443_), .C(_abc_40319_new_n1762_), .Y(_abc_40319_new_n1763_));
AOI21X1 AOI21X1_79 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1761_), .C(_abc_40319_new_n1764_), .Y(_abc_40319_new_n1765_));
AOI21X1 AOI21X1_8 ( .A(_abc_40319_new_n761_), .B(_abc_40319_new_n756_), .C(_abc_40319_new_n741_), .Y(_abc_40319_new_n762_));
AOI21X1 AOI21X1_80 ( .A(_abc_40319_new_n1416_), .B(_abc_40319_new_n1340_), .C(_abc_40319_new_n1413_), .Y(_abc_40319_new_n1770_));
AOI21X1 AOI21X1_81 ( .A(_abc_40319_new_n978_), .B(_abc_40319_new_n1360_), .C(_abc_40319_new_n1773_), .Y(_abc_40319_new_n1774_));
AOI21X1 AOI21X1_82 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n1325_), .C(_abc_40319_new_n1776_), .Y(_abc_40319_new_n1777_));
AOI21X1 AOI21X1_83 ( .A(_abc_40319_new_n1781_), .B(_abc_40319_new_n1783_), .C(_abc_40319_new_n677_), .Y(_abc_40319_new_n1784_));
AOI21X1 AOI21X1_84 ( .A(n1336), .B(REG3_REG_22_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n1789_));
AOI21X1 AOI21X1_85 ( .A(n1336), .B(REG3_REG_11_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n1800_));
AOI21X1 AOI21X1_86 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1799_), .C(_abc_40319_new_n1801_), .Y(_abc_40319_new_n1802_));
AOI21X1 AOI21X1_87 ( .A(_abc_40319_new_n1551_), .B(_abc_40319_new_n1806_), .C(_abc_40319_new_n677_), .Y(_abc_40319_new_n1807_));
AOI21X1 AOI21X1_88 ( .A(_abc_40319_new_n1002_), .B(REG3_REG_2_), .C(_abc_40319_new_n1815_), .Y(_abc_40319_new_n1816_));
AOI21X1 AOI21X1_89 ( .A(_abc_40319_new_n1818_), .B(_abc_40319_new_n1819_), .C(_abc_40319_new_n677_), .Y(_abc_40319_new_n1820_));
AOI21X1 AOI21X1_9 ( .A(_abc_40319_new_n790_), .B(_abc_40319_new_n787_), .C(_abc_40319_new_n784_), .Y(_abc_40319_new_n791_));
AOI21X1 AOI21X1_90 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1824_), .C(_abc_40319_new_n1827_), .Y(_abc_40319_new_n1828_));
AOI21X1 AOI21X1_91 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n944_), .C(_abc_40319_new_n1837_), .Y(_abc_40319_new_n1838_));
AOI21X1 AOI21X1_92 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1836_), .C(_abc_40319_new_n1839_), .Y(_abc_40319_new_n1840_));
AOI21X1 AOI21X1_93 ( .A(_abc_40319_new_n1846_), .B(_abc_40319_new_n1069_), .C(_abc_40319_new_n1104_), .Y(_abc_40319_new_n1847_));
AOI21X1 AOI21X1_94 ( .A(n1336), .B(REG3_REG_26_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n1853_));
AOI21X1 AOI21X1_95 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1852_), .C(_abc_40319_new_n1854_), .Y(_abc_40319_new_n1855_));
AOI21X1 AOI21X1_96 ( .A(_abc_40319_new_n1858_), .B(_abc_40319_new_n1859_), .C(_abc_40319_new_n677_), .Y(_abc_40319_new_n1860_));
AOI21X1 AOI21X1_97 ( .A(n1336), .B(REG3_REG_15_), .C(_abc_40319_new_n619_), .Y(_abc_40319_new_n1866_));
AOI21X1 AOI21X1_98 ( .A(_abc_40319_new_n1002_), .B(_abc_40319_new_n1230_), .C(_abc_40319_new_n1867_), .Y(_abc_40319_new_n1868_));
AOI21X1 AOI21X1_99 ( .A(_abc_40319_new_n1889_), .B(_abc_40319_new_n838_), .C(_abc_40319_new_n1873_), .Y(_abc_40319_new_n1890_));
AOI22X1 AOI22X1_1 ( .A(_abc_40319_new_n572_), .B(_abc_40319_new_n623_), .C(_abc_40319_new_n655_), .D(_abc_40319_new_n627_), .Y(_abc_40319_new_n656_));
AOI22X1 AOI22X1_10 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n769_), .C(_abc_40319_new_n783_), .D(_abc_40319_new_n683_), .Y(_abc_40319_new_n784_));
AOI22X1 AOI22X1_100 ( .A(_abc_40319_new_n1017_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n1592_), .Y(_abc_40319_new_n2077_));
AOI22X1 AOI22X1_101 ( .A(_abc_40319_new_n2074_), .B(_abc_40319_new_n2070_), .C(_abc_40319_new_n2077_), .D(_abc_40319_new_n2076_), .Y(_abc_40319_new_n2078_));
AOI22X1 AOI22X1_102 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1582_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n1046_), .Y(_abc_40319_new_n2080_));
AOI22X1 AOI22X1_103 ( .A(_abc_40319_new_n1875_), .B(_abc_40319_new_n2088_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n1598_), .Y(_abc_40319_new_n2092_));
AOI22X1 AOI22X1_104 ( .A(_abc_40319_new_n2091_), .B(_abc_40319_new_n2092_), .C(_abc_40319_new_n2082_), .D(_abc_40319_new_n2084_), .Y(_abc_40319_new_n2093_));
AOI22X1 AOI22X1_105 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n2097_), .C(_abc_40319_new_n1875_), .D(_abc_40319_new_n2103_), .Y(_abc_40319_new_n2104_));
AOI22X1 AOI22X1_106 ( .A(_abc_40319_new_n1875_), .B(_abc_40319_new_n2097_), .C(_abc_40319_new_n609_), .D(_abc_40319_new_n2103_), .Y(_abc_40319_new_n2107_));
AOI22X1 AOI22X1_107 ( .A(_abc_40319_new_n2105_), .B(_abc_40319_new_n2109_), .C(_abc_40319_new_n2095_), .D(_abc_40319_new_n2094_), .Y(_abc_40319_new_n2110_));
AOI22X1 AOI22X1_108 ( .A(_abc_40319_new_n2274_), .B(_abc_40319_new_n579_), .C(_abc_40319_new_n1907_), .D(_abc_40319_new_n2277_), .Y(_abc_40319_new_n2278_));
AOI22X1 AOI22X1_109 ( .A(_abc_40319_new_n2272_), .B(_abc_40319_new_n1896_), .C(_abc_40319_new_n1914_), .D(_abc_40319_new_n2280_), .Y(_abc_40319_new_n2281_));
AOI22X1 AOI22X1_11 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n799_), .C(_abc_40319_new_n809_), .D(_abc_40319_new_n683_), .Y(_abc_40319_new_n810_));
AOI22X1 AOI22X1_110 ( .A(_abc_40319_new_n1885_), .B(_abc_40319_new_n1886_), .C(_abc_40319_new_n2305_), .D(_abc_40319_new_n2304_), .Y(_abc_40319_new_n2306_));
AOI22X1 AOI22X1_111 ( .A(_abc_40319_new_n2352_), .B(_abc_40319_new_n2367_), .C(_abc_40319_new_n2361_), .D(_abc_40319_new_n2357_), .Y(_abc_40319_new_n2368_));
AOI22X1 AOI22X1_112 ( .A(_abc_40319_new_n2320_), .B(_abc_40319_new_n2383_), .C(_abc_40319_new_n2385_), .D(_abc_40319_new_n2329_), .Y(_abc_40319_new_n2386_));
AOI22X1 AOI22X1_113 ( .A(_abc_40319_new_n2123_), .B(_abc_40319_new_n2393_), .C(_abc_40319_new_n2348_), .D(_abc_40319_new_n2396_), .Y(_abc_40319_new_n2397_));
AOI22X1 AOI22X1_114 ( .A(_abc_40319_new_n1018_), .B(_abc_40319_new_n1592_), .C(_abc_40319_new_n1582_), .D(_abc_40319_new_n1505_), .Y(_abc_40319_new_n2404_));
AOI22X1 AOI22X1_115 ( .A(_abc_40319_new_n2516_), .B(_abc_40319_new_n667_), .C(_abc_40319_new_n2514_), .D(_abc_40319_new_n2517_), .Y(_abc_40319_new_n2518_));
AOI22X1 AOI22X1_116 ( .A(_abc_40319_new_n580_), .B(_abc_40319_new_n608_), .C(_abc_40319_new_n1872_), .D(_abc_40319_new_n972_), .Y(_abc_40319_new_n2527_));
AOI22X1 AOI22X1_117 ( .A(_abc_40319_new_n871_), .B(_abc_40319_new_n907_), .C(_abc_40319_new_n2534_), .D(_abc_40319_new_n2535_), .Y(_abc_40319_new_n2536_));
AOI22X1 AOI22X1_118 ( .A(_abc_40319_new_n977_), .B(_abc_40319_new_n892_), .C(_abc_40319_new_n2523_), .D(_abc_40319_new_n2553_), .Y(_abc_40319_new_n2554_));
AOI22X1 AOI22X1_119 ( .A(_abc_40319_new_n977_), .B(_abc_40319_new_n796_), .C(_abc_40319_new_n2523_), .D(_abc_40319_new_n2601_), .Y(_abc_40319_new_n2602_));
AOI22X1 AOI22X1_12 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n809_), .C(_abc_40319_new_n799_), .D(_abc_40319_new_n813_), .Y(_abc_40319_new_n814_));
AOI22X1 AOI22X1_120 ( .A(ADDR_REG_4_), .B(_abc_40319_new_n2539_), .C(_abc_40319_new_n2603_), .D(_abc_40319_new_n2543_), .Y(_abc_40319_new_n2604_));
AOI22X1 AOI22X1_121 ( .A(_abc_40319_new_n2523_), .B(_abc_40319_new_n2706_), .C(_abc_40319_new_n2524_), .D(_abc_40319_new_n2699_), .Y(_abc_40319_new_n2707_));
AOI22X1 AOI22X1_122 ( .A(_abc_40319_new_n977_), .B(_abc_40319_new_n1390_), .C(_abc_40319_new_n2523_), .D(_abc_40319_new_n2720_), .Y(_abc_40319_new_n2721_));
AOI22X1 AOI22X1_123 ( .A(ADDR_REG_13_), .B(_abc_40319_new_n2539_), .C(_abc_40319_new_n2797_), .D(_abc_40319_new_n2542_), .Y(_abc_40319_new_n2798_));
AOI22X1 AOI22X1_124 ( .A(ADDR_REG_16_), .B(_abc_40319_new_n2539_), .C(_abc_40319_new_n2855_), .D(_abc_40319_new_n2684_), .Y(_abc_40319_new_n2872_));
AOI22X1 AOI22X1_125 ( .A(ADDR_REG_18_), .B(_abc_40319_new_n2539_), .C(_abc_40319_new_n2926_), .D(_abc_40319_new_n2543_), .Y(_abc_40319_new_n2928_));
AOI22X1 AOI22X1_126 ( .A(_abc_40319_new_n2205_), .B(_abc_40319_new_n3057_), .C(_abc_40319_new_n3061_), .D(_abc_40319_new_n3063_), .Y(_abc_40319_new_n3064_));
AOI22X1 AOI22X1_127 ( .A(_abc_40319_new_n1070_), .B(_abc_40319_new_n1078_), .C(_abc_40319_new_n1054_), .D(_abc_40319_new_n1496_), .Y(_abc_40319_new_n3081_));
AOI22X1 AOI22X1_128 ( .A(_abc_40319_new_n2135_), .B(_abc_40319_new_n2461_), .C(_abc_40319_new_n2502_), .D(_abc_40319_new_n2498_), .Y(_abc_40319_new_n3206_));
AOI22X1 AOI22X1_129 ( .A(_abc_40319_new_n1109_), .B(_abc_40319_new_n2991_), .C(_abc_40319_new_n2996_), .D(_abc_40319_new_n3226_), .Y(_abc_40319_new_n3227_));
AOI22X1 AOI22X1_13 ( .A(_abc_40319_new_n729_), .B(_abc_40319_new_n727_), .C(REG0_REG_3_), .D(_abc_40319_new_n724_), .Y(_abc_40319_new_n831_));
AOI22X1 AOI22X1_130 ( .A(_abc_40319_new_n3234_), .B(_abc_40319_new_n3235_), .C(_abc_40319_new_n2138_), .D(_abc_40319_new_n3233_), .Y(_abc_40319_new_n3236_));
AOI22X1 AOI22X1_131 ( .A(_abc_40319_new_n1123_), .B(_abc_40319_new_n2991_), .C(_abc_40319_new_n2996_), .D(_abc_40319_new_n3251_), .Y(_abc_40319_new_n3252_));
AOI22X1 AOI22X1_132 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3255_), .C(_abc_40319_new_n3256_), .D(_abc_40319_new_n3261_), .Y(_abc_40319_new_n3262_));
AOI22X1 AOI22X1_133 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1186_), .C(_abc_40319_new_n1209_), .D(_abc_40319_new_n3108_), .Y(_abc_40319_new_n3376_));
AOI22X1 AOI22X1_134 ( .A(_abc_40319_new_n1233_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3101_), .D(_abc_40319_new_n3386_), .Y(_abc_40319_new_n3387_));
AOI22X1 AOI22X1_135 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1230_), .C(_abc_40319_new_n1189_), .D(_abc_40319_new_n3108_), .Y(_abc_40319_new_n3394_));
AOI22X1 AOI22X1_136 ( .A(_abc_40319_new_n1259_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3101_), .D(_abc_40319_new_n3398_), .Y(_abc_40319_new_n3401_));
AOI22X1 AOI22X1_137 ( .A(_abc_40319_new_n1336_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3101_), .D(_abc_40319_new_n3410_), .Y(_abc_40319_new_n3411_));
AOI22X1 AOI22X1_138 ( .A(_abc_40319_new_n993_), .B(_abc_40319_new_n1248_), .C(_abc_40319_new_n3368_), .D(_abc_40319_new_n1233_), .Y(_abc_40319_new_n3418_));
AOI22X1 AOI22X1_139 ( .A(_abc_40319_new_n1360_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3101_), .D(_abc_40319_new_n3431_), .Y(_abc_40319_new_n3432_));
AOI22X1 AOI22X1_14 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n826_), .C(_abc_40319_new_n832_), .D(_abc_40319_new_n683_), .Y(_abc_40319_new_n833_));
AOI22X1 AOI22X1_140 ( .A(_abc_40319_new_n1352_), .B(_abc_40319_new_n2991_), .C(_abc_40319_new_n2996_), .D(_abc_40319_new_n3446_), .Y(_abc_40319_new_n3447_));
AOI22X1 AOI22X1_141 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1357_), .C(_abc_40319_new_n3133_), .D(_abc_40319_new_n3449_), .Y(_abc_40319_new_n3450_));
AOI22X1 AOI22X1_142 ( .A(_abc_40319_new_n1380_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3101_), .D(_abc_40319_new_n3449_), .Y(_abc_40319_new_n3453_));
AOI22X1 AOI22X1_143 ( .A(_abc_40319_new_n1371_), .B(_abc_40319_new_n2991_), .C(_abc_40319_new_n2996_), .D(_abc_40319_new_n3461_), .Y(_abc_40319_new_n3462_));
AOI22X1 AOI22X1_144 ( .A(_abc_40319_new_n1008_), .B(_abc_40319_new_n1799_), .C(_abc_40319_new_n3133_), .D(_abc_40319_new_n3463_), .Y(_abc_40319_new_n3464_));
AOI22X1 AOI22X1_145 ( .A(_abc_40319_new_n1309_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3101_), .D(_abc_40319_new_n3481_), .Y(_abc_40319_new_n3482_));
AOI22X1 AOI22X1_146 ( .A(_abc_40319_new_n987_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3101_), .D(_abc_40319_new_n3498_), .Y(_abc_40319_new_n3499_));
AOI22X1 AOI22X1_147 ( .A(_abc_40319_new_n954_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3101_), .D(_abc_40319_new_n3532_), .Y(_abc_40319_new_n3533_));
AOI22X1 AOI22X1_148 ( .A(_abc_40319_new_n698_), .B(_abc_40319_new_n993_), .C(_abc_40319_new_n987_), .D(_abc_40319_new_n3368_), .Y(_abc_40319_new_n3539_));
AOI22X1 AOI22X1_149 ( .A(_abc_40319_new_n832_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3101_), .D(_abc_40319_new_n3567_), .Y(_abc_40319_new_n3568_));
AOI22X1 AOI22X1_15 ( .A(REG3_REG_2_), .B(_abc_40319_new_n727_), .C(REG1_REG_2_), .D(_abc_40319_new_n726_), .Y(_abc_40319_new_n840_));
AOI22X1 AOI22X1_150 ( .A(_abc_40319_new_n799_), .B(_abc_40319_new_n993_), .C(_abc_40319_new_n783_), .D(_abc_40319_new_n3368_), .Y(_abc_40319_new_n3573_));
AOI22X1 AOI22X1_151 ( .A(_abc_40319_new_n842_), .B(_abc_40319_new_n3103_), .C(_abc_40319_new_n3101_), .D(_abc_40319_new_n3600_), .Y(_abc_40319_new_n3601_));
AOI22X1 AOI22X1_152 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n993_), .C(_abc_40319_new_n832_), .D(_abc_40319_new_n3368_), .Y(_abc_40319_new_n3618_));
AOI22X1 AOI22X1_153 ( .A(_abc_40319_new_n877_), .B(_abc_40319_new_n993_), .C(_abc_40319_new_n842_), .D(_abc_40319_new_n3368_), .Y(_abc_40319_new_n3638_));
AOI22X1 AOI22X1_154 ( .A(DATAI_30_), .B(n1336), .C(IR_REG_30_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3721_));
AOI22X1 AOI22X1_155 ( .A(DATAI_29_), .B(n1336), .C(IR_REG_29_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3723_));
AOI22X1 AOI22X1_156 ( .A(DATAI_27_), .B(n1336), .C(IR_REG_27_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3732_));
AOI22X1 AOI22X1_157 ( .A(DATAI_21_), .B(n1336), .C(IR_REG_21_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3753_));
AOI22X1 AOI22X1_158 ( .A(DATAI_19_), .B(n1336), .C(IR_REG_19_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3761_));
AOI22X1 AOI22X1_159 ( .A(DATAI_18_), .B(n1336), .C(IR_REG_18_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3763_));
AOI22X1 AOI22X1_16 ( .A(_abc_40319_new_n715_), .B(REG2_REG_2_), .C(REG0_REG_2_), .D(_abc_40319_new_n724_), .Y(_abc_40319_new_n841_));
AOI22X1 AOI22X1_160 ( .A(DATAI_17_), .B(n1336), .C(IR_REG_17_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3767_));
AOI22X1 AOI22X1_161 ( .A(DATAI_16_), .B(n1336), .C(IR_REG_16_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3769_));
AOI22X1 AOI22X1_162 ( .A(DATAI_15_), .B(n1336), .C(IR_REG_15_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3774_));
AOI22X1 AOI22X1_163 ( .A(DATAI_14_), .B(n1336), .C(IR_REG_14_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3776_));
AOI22X1 AOI22X1_164 ( .A(DATAI_13_), .B(n1336), .C(IR_REG_13_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3780_));
AOI22X1 AOI22X1_165 ( .A(DATAI_11_), .B(n1336), .C(IR_REG_11_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3788_));
AOI22X1 AOI22X1_166 ( .A(DATAI_10_), .B(n1336), .C(IR_REG_10_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3791_));
AOI22X1 AOI22X1_167 ( .A(DATAI_9_), .B(n1336), .C(IR_REG_9_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3793_));
AOI22X1 AOI22X1_168 ( .A(DATAI_8_), .B(n1336), .C(IR_REG_8_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3796_));
AOI22X1 AOI22X1_169 ( .A(DATAI_7_), .B(n1336), .C(IR_REG_7_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3799_));
AOI22X1 AOI22X1_17 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n839_), .C(_abc_40319_new_n842_), .D(_abc_40319_new_n683_), .Y(_abc_40319_new_n843_));
AOI22X1 AOI22X1_170 ( .A(DATAI_6_), .B(n1336), .C(IR_REG_6_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3802_));
AOI22X1 AOI22X1_171 ( .A(DATAI_5_), .B(n1336), .C(IR_REG_5_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3806_));
AOI22X1 AOI22X1_172 ( .A(DATAI_4_), .B(n1336), .C(IR_REG_4_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3808_));
AOI22X1 AOI22X1_173 ( .A(DATAI_2_), .B(n1336), .C(IR_REG_2_), .D(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3817_));
AOI22X1 AOI22X1_174 ( .A(_abc_40319_new_n3827_), .B(_abc_40319_new_n2267_), .C(_abc_40319_new_n1505_), .D(_abc_40319_new_n3828_), .Y(_abc_40319_new_n3829_));
AOI22X1 AOI22X1_175 ( .A(_abc_40319_new_n993_), .B(_abc_40319_new_n1371_), .C(_abc_40319_new_n3620_), .D(_abc_40319_new_n3461_), .Y(_abc_40319_new_n3960_));
AOI22X1 AOI22X1_176 ( .A(_abc_40319_new_n1360_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n3893_), .D(_abc_40319_new_n3463_), .Y(_abc_40319_new_n3961_));
AOI22X1 AOI22X1_177 ( .A(_abc_40319_new_n993_), .B(_abc_40319_new_n1352_), .C(_abc_40319_new_n3620_), .D(_abc_40319_new_n3446_), .Y(_abc_40319_new_n3967_));
AOI22X1 AOI22X1_178 ( .A(_abc_40319_new_n1336_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n3893_), .D(_abc_40319_new_n3449_), .Y(_abc_40319_new_n3968_));
AOI22X1 AOI22X1_179 ( .A(_abc_40319_new_n1259_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n3893_), .D(_abc_40319_new_n3431_), .Y(_abc_40319_new_n3973_));
AOI22X1 AOI22X1_18 ( .A(_abc_40319_new_n726_), .B(REG1_REG_1_), .C(REG0_REG_1_), .D(_abc_40319_new_n724_), .Y(_abc_40319_new_n878_));
AOI22X1 AOI22X1_180 ( .A(_abc_40319_new_n993_), .B(_abc_40319_new_n1223_), .C(_abc_40319_new_n3620_), .D(_abc_40319_new_n3395_), .Y(_abc_40319_new_n3982_));
AOI22X1 AOI22X1_181 ( .A(_abc_40319_new_n1189_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n3893_), .D(_abc_40319_new_n3398_), .Y(_abc_40319_new_n3983_));
AOI22X1 AOI22X1_182 ( .A(_abc_40319_new_n993_), .B(_abc_40319_new_n1148_), .C(_abc_40319_new_n3620_), .D(_abc_40319_new_n3334_), .Y(_abc_40319_new_n4001_));
AOI22X1 AOI22X1_183 ( .A(_abc_40319_new_n1437_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n3893_), .D(_abc_40319_new_n3324_), .Y(_abc_40319_new_n4002_));
AOI22X1 AOI22X1_184 ( .A(_abc_40319_new_n1452_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n3893_), .D(_abc_40319_new_n3308_), .Y(_abc_40319_new_n4008_));
AOI22X1 AOI22X1_185 ( .A(_abc_40319_new_n993_), .B(_abc_40319_new_n1109_), .C(_abc_40319_new_n3620_), .D(_abc_40319_new_n3226_), .Y(_abc_40319_new_n4028_));
AOI22X1 AOI22X1_186 ( .A(_abc_40319_new_n1094_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n3893_), .D(_abc_40319_new_n3229_), .Y(_abc_40319_new_n4029_));
AOI22X1 AOI22X1_187 ( .A(_abc_40319_new_n993_), .B(_abc_40319_new_n1085_), .C(_abc_40319_new_n3620_), .D(_abc_40319_new_n3213_), .Y(_abc_40319_new_n4034_));
AOI22X1 AOI22X1_188 ( .A(_abc_40319_new_n1077_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n3893_), .D(_abc_40319_new_n3204_), .Y(_abc_40319_new_n4035_));
AOI22X1 AOI22X1_189 ( .A(_abc_40319_new_n1065_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n3893_), .D(_abc_40319_new_n3177_), .Y(_abc_40319_new_n4041_));
AOI22X1 AOI22X1_19 ( .A(REG3_REG_1_), .B(_abc_40319_new_n727_), .C(REG2_REG_1_), .D(_abc_40319_new_n715_), .Y(_abc_40319_new_n879_));
AOI22X1 AOI22X1_190 ( .A(_abc_40319_new_n993_), .B(_abc_40319_new_n1055_), .C(_abc_40319_new_n3620_), .D(_abc_40319_new_n3163_), .Y(_abc_40319_new_n4046_));
AOI22X1 AOI22X1_191 ( .A(_abc_40319_new_n1046_), .B(_abc_40319_new_n3368_), .C(_abc_40319_new_n3893_), .D(_abc_40319_new_n3154_), .Y(_abc_40319_new_n4047_));
AOI22X1 AOI22X1_192 ( .A(_abc_40319_new_n993_), .B(_abc_40319_new_n1582_), .C(_abc_40319_new_n3620_), .D(_abc_40319_new_n3111_), .Y(_abc_40319_new_n4061_));
AOI22X1 AOI22X1_2 ( .A(_abc_40319_new_n707_), .B(_abc_40319_new_n708_), .C(_abc_40319_new_n709_), .D(_abc_40319_new_n714_), .Y(_abc_40319_new_n715_));
AOI22X1 AOI22X1_20 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n877_), .C(_abc_40319_new_n880_), .D(_abc_40319_new_n683_), .Y(_abc_40319_new_n881_));
AOI22X1 AOI22X1_21 ( .A(IR_REG_0_), .B(_abc_40319_new_n671_), .C(_abc_40319_new_n914_), .D(_abc_40319_new_n679_), .Y(_abc_40319_new_n915_));
AOI22X1 AOI22X1_22 ( .A(_abc_40319_new_n868_), .B(_abc_40319_new_n833_), .C(_abc_40319_new_n843_), .D(_abc_40319_new_n932_), .Y(_abc_40319_new_n933_));
AOI22X1 AOI22X1_23 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n944_), .C(_abc_40319_new_n954_), .D(_abc_40319_new_n683_), .Y(_abc_40319_new_n955_));
AOI22X1 AOI22X1_24 ( .A(_abc_40319_new_n727_), .B(_abc_40319_new_n984_), .C(REG1_REG_8_), .D(_abc_40319_new_n726_), .Y(_abc_40319_new_n985_));
AOI22X1 AOI22X1_25 ( .A(_abc_40319_new_n715_), .B(REG2_REG_8_), .C(REG0_REG_8_), .D(_abc_40319_new_n724_), .Y(_abc_40319_new_n986_));
AOI22X1 AOI22X1_26 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1018_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1046_), .Y(_abc_40319_new_n1047_));
AOI22X1 AOI22X1_27 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1018_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1046_), .Y(_abc_40319_new_n1048_));
AOI22X1 AOI22X1_28 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1055_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1065_), .Y(_abc_40319_new_n1066_));
AOI22X1 AOI22X1_29 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1055_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1065_), .Y(_abc_40319_new_n1067_));
AOI22X1 AOI22X1_3 ( .A(_abc_40319_new_n715_), .B(REG2_REG_7_), .C(REG0_REG_7_), .D(_abc_40319_new_n724_), .Y(_abc_40319_new_n725_));
AOI22X1 AOI22X1_30 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1080_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1077_), .Y(_abc_40319_new_n1081_));
AOI22X1 AOI22X1_31 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1085_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1094_), .Y(_abc_40319_new_n1095_));
AOI22X1 AOI22X1_32 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1109_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1115_), .Y(_abc_40319_new_n1116_));
AOI22X1 AOI22X1_33 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1109_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1115_), .Y(_abc_40319_new_n1117_));
AOI22X1 AOI22X1_34 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1123_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1135_), .Y(_abc_40319_new_n1136_));
AOI22X1 AOI22X1_35 ( .A(_abc_40319_new_n715_), .B(REG2_REG_18_), .C(REG0_REG_18_), .D(_abc_40319_new_n724_), .Y(_abc_40319_new_n1154_));
AOI22X1 AOI22X1_36 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1148_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1157_), .Y(_abc_40319_new_n1158_));
AOI22X1 AOI22X1_37 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1175_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1189_), .Y(_abc_40319_new_n1190_));
AOI22X1 AOI22X1_38 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1175_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1189_), .Y(_abc_40319_new_n1192_));
AOI22X1 AOI22X1_39 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1198_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1209_), .Y(_abc_40319_new_n1210_));
AOI22X1 AOI22X1_4 ( .A(_abc_40319_new_n721_), .B(_abc_40319_new_n722_), .C(_abc_40319_new_n716_), .D(_abc_40319_new_n719_), .Y(_abc_40319_new_n726_));
AOI22X1 AOI22X1_40 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1223_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1233_), .Y(_abc_40319_new_n1234_));
AOI22X1 AOI22X1_41 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1223_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1233_), .Y(_abc_40319_new_n1235_));
AOI22X1 AOI22X1_42 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1248_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1259_), .Y(_abc_40319_new_n1260_));
AOI22X1 AOI22X1_43 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1276_), .C(_abc_40319_new_n987_), .D(_abc_40319_new_n683_), .Y(_abc_40319_new_n1277_));
AOI22X1 AOI22X1_44 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n987_), .C(_abc_40319_new_n1276_), .D(_abc_40319_new_n813_), .Y(_abc_40319_new_n1278_));
AOI22X1 AOI22X1_45 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1309_), .C(_abc_40319_new_n1297_), .D(_abc_40319_new_n813_), .Y(_abc_40319_new_n1310_));
AOI22X1 AOI22X1_46 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1297_), .C(_abc_40319_new_n1309_), .D(_abc_40319_new_n683_), .Y(_abc_40319_new_n1315_));
AOI22X1 AOI22X1_47 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1325_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1336_), .Y(_abc_40319_new_n1337_));
AOI22X1 AOI22X1_48 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1325_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1336_), .Y(_abc_40319_new_n1338_));
AOI22X1 AOI22X1_49 ( .A(_abc_40319_new_n683_), .B(_abc_40319_new_n1360_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1352_), .Y(_abc_40319_new_n1361_));
AOI22X1 AOI22X1_5 ( .A(_abc_40319_new_n721_), .B(_abc_40319_new_n722_), .C(_abc_40319_new_n708_), .D(_abc_40319_new_n707_), .Y(_abc_40319_new_n727_));
AOI22X1 AOI22X1_50 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1360_), .C(_abc_40319_new_n813_), .D(_abc_40319_new_n1352_), .Y(_abc_40319_new_n1362_));
AOI22X1 AOI22X1_51 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1371_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1380_), .Y(_abc_40319_new_n1381_));
AOI22X1 AOI22X1_52 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1393_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1402_), .Y(_abc_40319_new_n1403_));
AOI22X1 AOI22X1_53 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1393_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1402_), .Y(_abc_40319_new_n1405_));
AOI22X1 AOI22X1_54 ( .A(_abc_40319_new_n1386_), .B(_abc_40319_new_n1409_), .C(_abc_40319_new_n1340_), .D(_abc_40319_new_n1417_), .Y(_abc_40319_new_n1418_));
AOI22X1 AOI22X1_55 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1429_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1437_), .Y(_abc_40319_new_n1438_));
AOI22X1 AOI22X1_56 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1429_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1437_), .Y(_abc_40319_new_n1440_));
AOI22X1 AOI22X1_57 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1443_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1452_), .Y(_abc_40319_new_n1453_));
AOI22X1 AOI22X1_58 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1443_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1452_), .Y(_abc_40319_new_n1455_));
AOI22X1 AOI22X1_59 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1460_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1469_), .Y(_abc_40319_new_n1470_));
AOI22X1 AOI22X1_6 ( .A(_abc_40319_new_n727_), .B(_abc_40319_new_n738_), .C(REG1_REG_7_), .D(_abc_40319_new_n726_), .Y(_abc_40319_new_n739_));
AOI22X1 AOI22X1_60 ( .A(_abc_40319_new_n813_), .B(_abc_40319_new_n1460_), .C(_abc_40319_new_n679_), .D(_abc_40319_new_n1469_), .Y(_abc_40319_new_n1472_));
AOI22X1 AOI22X1_61 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n1582_), .C(_abc_40319_new_n683_), .D(_abc_40319_new_n1580_), .Y(_abc_40319_new_n1583_));
AOI22X1 AOI22X1_62 ( .A(_abc_40319_new_n1579_), .B(_abc_40319_new_n1587_), .C(_abc_40319_new_n1588_), .D(_abc_40319_new_n1590_), .Y(_abc_40319_new_n1591_));
AOI22X1 AOI22X1_63 ( .A(_abc_40319_new_n1875_), .B(_abc_40319_new_n1877_), .C(_abc_40319_new_n1874_), .D(_abc_40319_new_n1883_), .Y(_abc_40319_new_n1884_));
AOI22X1 AOI22X1_64 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1877_), .C(_abc_40319_new_n1875_), .D(_abc_40319_new_n1883_), .Y(_abc_40319_new_n1886_));
AOI22X1 AOI22X1_65 ( .A(_abc_40319_new_n853_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n855_), .Y(_abc_40319_new_n1896_));
AOI22X1 AOI22X1_66 ( .A(_abc_40319_new_n715_), .B(REG2_REG_0_), .C(REG0_REG_0_), .D(_abc_40319_new_n724_), .Y(_abc_40319_new_n1903_));
AOI22X1 AOI22X1_67 ( .A(REG3_REG_0_), .B(_abc_40319_new_n727_), .C(REG1_REG_0_), .D(_abc_40319_new_n726_), .Y(_abc_40319_new_n1904_));
AOI22X1 AOI22X1_68 ( .A(_abc_40319_new_n1893_), .B(_abc_40319_new_n1897_), .C(_abc_40319_new_n580_), .D(_abc_40319_new_n1908_), .Y(_abc_40319_new_n1909_));
AOI22X1 AOI22X1_69 ( .A(_abc_40319_new_n825_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n865_), .Y(_abc_40319_new_n1914_));
AOI22X1 AOI22X1_7 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n698_), .C(_abc_40319_new_n740_), .D(_abc_40319_new_n683_), .Y(_abc_40319_new_n741_));
AOI22X1 AOI22X1_70 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n799_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n832_), .Y(_abc_40319_new_n1919_));
AOI22X1 AOI22X1_71 ( .A(_abc_40319_new_n1915_), .B(_abc_40319_new_n1913_), .C(_abc_40319_new_n1918_), .D(_abc_40319_new_n1920_), .Y(_abc_40319_new_n1921_));
AOI22X1 AOI22X1_72 ( .A(_abc_40319_new_n769_), .B(_abc_40319_new_n1874_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n809_), .Y(_abc_40319_new_n1937_));
AOI22X1 AOI22X1_73 ( .A(_abc_40319_new_n1938_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n788_), .Y(_abc_40319_new_n1939_));
AOI22X1 AOI22X1_74 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1297_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n987_), .Y(_abc_40319_new_n1949_));
AOI22X1 AOI22X1_75 ( .A(_abc_40319_new_n1308_), .B(_abc_40319_new_n1895_), .C(_abc_40319_new_n1875_), .D(_abc_40319_new_n1739_), .Y(_abc_40319_new_n1951_));
AOI22X1 AOI22X1_76 ( .A(_abc_40319_new_n1950_), .B(_abc_40319_new_n1952_), .C(_abc_40319_new_n1947_), .D(_abc_40319_new_n1948_), .Y(_abc_40319_new_n1953_));
AOI22X1 AOI22X1_77 ( .A(_abc_40319_new_n1927_), .B(_abc_40319_new_n1928_), .C(_abc_40319_new_n1962_), .D(_abc_40319_new_n1963_), .Y(_abc_40319_new_n1964_));
AOI22X1 AOI22X1_78 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1325_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n1360_), .Y(_abc_40319_new_n1975_));
AOI22X1 AOI22X1_79 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1248_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n1336_), .Y(_abc_40319_new_n1998_));
AOI22X1 AOI22X1_8 ( .A(_abc_40319_new_n749_), .B(_abc_40319_new_n608_), .C(_abc_40319_new_n610_), .D(_abc_40319_new_n748_), .Y(_abc_40319_new_n750_));
AOI22X1 AOI22X1_80 ( .A(_abc_40319_new_n1976_), .B(_abc_40319_new_n1977_), .C(_abc_40319_new_n2000_), .D(_abc_40319_new_n1999_), .Y(_abc_40319_new_n2001_));
AOI22X1 AOI22X1_81 ( .A(_abc_40319_new_n1865_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n1516_), .Y(_abc_40319_new_n2008_));
AOI22X1 AOI22X1_82 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1175_), .C(_abc_40319_new_n1875_), .D(_abc_40319_new_n1189_), .Y(_abc_40319_new_n2011_));
AOI22X1 AOI22X1_83 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1198_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n1189_), .Y(_abc_40319_new_n2017_));
AOI22X1 AOI22X1_84 ( .A(_abc_40319_new_n1159_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n1156_), .Y(_abc_40319_new_n2025_));
AOI22X1 AOI22X1_85 ( .A(_abc_40319_new_n1570_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n1759_), .Y(_abc_40319_new_n2032_));
AOI22X1 AOI22X1_86 ( .A(_abc_40319_new_n2024_), .B(_abc_40319_new_n2025_), .C(_abc_40319_new_n2031_), .D(_abc_40319_new_n2032_), .Y(_abc_40319_new_n2033_));
AOI22X1 AOI22X1_87 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1443_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n1437_), .Y(_abc_40319_new_n2036_));
AOI22X1 AOI22X1_88 ( .A(_abc_40319_new_n2037_), .B(_abc_40319_new_n2038_), .C(_abc_40319_new_n2030_), .D(_abc_40319_new_n2035_), .Y(_abc_40319_new_n2039_));
AOI22X1 AOI22X1_89 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1460_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n1452_), .Y(_abc_40319_new_n2040_));
AOI22X1 AOI22X1_9 ( .A(_abc_40319_new_n600_), .B(IR_REG_29_), .C(_abc_40319_new_n590_), .D(_abc_40319_new_n703_), .Y(_abc_40319_new_n772_));
AOI22X1 AOI22X1_90 ( .A(_abc_40319_new_n1122_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n1137_), .Y(_abc_40319_new_n2048_));
AOI22X1 AOI22X1_91 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1109_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n1135_), .Y(_abc_40319_new_n2050_));
AOI22X1 AOI22X1_92 ( .A(_abc_40319_new_n1108_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n1710_), .Y(_abc_40319_new_n2053_));
AOI22X1 AOI22X1_93 ( .A(_abc_40319_new_n2047_), .B(_abc_40319_new_n2048_), .C(_abc_40319_new_n2053_), .D(_abc_40319_new_n2052_), .Y(_abc_40319_new_n2054_));
AOI22X1 AOI22X1_94 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1085_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n1115_), .Y(_abc_40319_new_n2056_));
AOI22X1 AOI22X1_95 ( .A(_abc_40319_new_n1084_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n1093_), .Y(_abc_40319_new_n2058_));
AOI22X1 AOI22X1_96 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1080_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n1094_), .Y(_abc_40319_new_n2063_));
AOI22X1 AOI22X1_97 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1055_), .C(_abc_40319_new_n1870_), .D(_abc_40319_new_n1077_), .Y(_abc_40319_new_n2068_));
AOI22X1 AOI22X1_98 ( .A(_abc_40319_new_n1054_), .B(_abc_40319_new_n1875_), .C(_abc_40319_new_n1895_), .D(_abc_40319_new_n1496_), .Y(_abc_40319_new_n2070_));
AOI22X1 AOI22X1_99 ( .A(_abc_40319_new_n2064_), .B(_abc_40319_new_n2065_), .C(_abc_40319_new_n2069_), .D(_abc_40319_new_n2071_), .Y(_abc_40319_new_n2072_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n978), .Q(ADDR_REG_19_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(n1014), .Q(ADDR_REG_10_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(clock), .D(n403), .Q(D_REG_13_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(clock), .D(n408), .Q(D_REG_14_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(clock), .D(n413), .Q(D_REG_15_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(clock), .D(n418), .Q(D_REG_16_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(clock), .D(n423), .Q(D_REG_17_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(clock), .D(n428), .Q(D_REG_18_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(clock), .D(n433), .Q(D_REG_19_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(clock), .D(n438), .Q(D_REG_20_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(clock), .D(n443), .Q(D_REG_21_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(clock), .D(n448), .Q(D_REG_22_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(n1018), .Q(ADDR_REG_9_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(clock), .D(n453), .Q(D_REG_23_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(clock), .D(n458), .Q(D_REG_24_));
DFFPOSX1 DFFPOSX1_112 ( .CLK(clock), .D(n463), .Q(D_REG_25_));
DFFPOSX1 DFFPOSX1_113 ( .CLK(clock), .D(n468), .Q(D_REG_26_));
DFFPOSX1 DFFPOSX1_114 ( .CLK(clock), .D(n473), .Q(D_REG_27_));
DFFPOSX1 DFFPOSX1_115 ( .CLK(clock), .D(n478), .Q(D_REG_28_));
DFFPOSX1 DFFPOSX1_116 ( .CLK(clock), .D(n483), .Q(D_REG_29_));
DFFPOSX1 DFFPOSX1_117 ( .CLK(clock), .D(n488), .Q(D_REG_30_));
DFFPOSX1 DFFPOSX1_118 ( .CLK(clock), .D(n493), .Q(D_REG_31_));
DFFPOSX1 DFFPOSX1_119 ( .CLK(clock), .D(n498), .Q(REG0_REG_0_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(n1022), .Q(ADDR_REG_8_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(clock), .D(n503), .Q(REG0_REG_1_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(clock), .D(n508), .Q(REG0_REG_2_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(clock), .D(n513), .Q(REG0_REG_3_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(clock), .D(n518), .Q(REG0_REG_4_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(clock), .D(n523), .Q(REG0_REG_5_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(clock), .D(n528), .Q(REG0_REG_6_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(clock), .D(n533), .Q(REG0_REG_7_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(clock), .D(n538), .Q(REG0_REG_8_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(clock), .D(n543), .Q(REG0_REG_9_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(clock), .D(n548), .Q(REG0_REG_10_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(n1026), .Q(ADDR_REG_7_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(clock), .D(n553), .Q(REG0_REG_11_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(clock), .D(n558), .Q(REG0_REG_12_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(clock), .D(n563), .Q(REG0_REG_13_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(clock), .D(n568), .Q(REG0_REG_14_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(clock), .D(n573), .Q(REG0_REG_15_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(clock), .D(n578), .Q(REG0_REG_16_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(clock), .D(n583), .Q(REG0_REG_17_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(clock), .D(n588), .Q(REG0_REG_18_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(clock), .D(n593), .Q(REG0_REG_19_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(clock), .D(n598), .Q(REG0_REG_20_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(n1030), .Q(ADDR_REG_6_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(clock), .D(n603), .Q(REG0_REG_21_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(clock), .D(n608), .Q(REG0_REG_22_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(clock), .D(n613), .Q(REG0_REG_23_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(clock), .D(n618), .Q(REG0_REG_24_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(clock), .D(n623), .Q(REG0_REG_25_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(clock), .D(n628), .Q(REG0_REG_26_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(clock), .D(n633), .Q(REG0_REG_27_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(clock), .D(n638), .Q(REG0_REG_28_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(clock), .D(n643), .Q(REG0_REG_29_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(clock), .D(n648), .Q(REG0_REG_30_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(n1034), .Q(ADDR_REG_5_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(clock), .D(n653), .Q(REG0_REG_31_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(clock), .D(n658), .Q(REG1_REG_0_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(clock), .D(n663), .Q(REG1_REG_1_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(clock), .D(n668), .Q(REG1_REG_2_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(clock), .D(n673), .Q(REG1_REG_3_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(clock), .D(n678), .Q(REG1_REG_4_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(clock), .D(n683), .Q(REG1_REG_5_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(clock), .D(n688), .Q(REG1_REG_6_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(clock), .D(n693), .Q(REG1_REG_7_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(clock), .D(n698), .Q(REG1_REG_8_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(n1038), .Q(ADDR_REG_4_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(clock), .D(n703), .Q(REG1_REG_9_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(clock), .D(n708), .Q(REG1_REG_10_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(clock), .D(n713), .Q(REG1_REG_11_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(clock), .D(n718), .Q(REG1_REG_12_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(clock), .D(n723), .Q(REG1_REG_13_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(clock), .D(n728), .Q(REG1_REG_14_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(clock), .D(n733), .Q(REG1_REG_15_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(clock), .D(n738), .Q(REG1_REG_16_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(clock), .D(n743), .Q(REG1_REG_17_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(clock), .D(n748), .Q(REG1_REG_18_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(n1042), .Q(ADDR_REG_3_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(clock), .D(n753), .Q(REG1_REG_19_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(clock), .D(n758), .Q(REG1_REG_20_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(clock), .D(n763), .Q(REG1_REG_21_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(clock), .D(n768), .Q(REG1_REG_22_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(clock), .D(n773), .Q(REG1_REG_23_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(clock), .D(n778), .Q(REG1_REG_24_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(clock), .D(n783), .Q(REG1_REG_25_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(clock), .D(n788), .Q(REG1_REG_26_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(clock), .D(n793), .Q(REG1_REG_27_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(clock), .D(n798), .Q(REG1_REG_28_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(n1046), .Q(ADDR_REG_2_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(clock), .D(n803), .Q(REG1_REG_29_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(clock), .D(n808), .Q(REG1_REG_30_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(clock), .D(n813), .Q(REG1_REG_31_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(clock), .D(n818), .Q(REG2_REG_0_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(clock), .D(n823), .Q(REG2_REG_1_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(clock), .D(n828), .Q(REG2_REG_2_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(clock), .D(n833), .Q(REG2_REG_3_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(clock), .D(n838), .Q(REG2_REG_4_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(clock), .D(n843), .Q(REG2_REG_5_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(clock), .D(n848), .Q(REG2_REG_6_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(n1050), .Q(ADDR_REG_1_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(clock), .D(n853), .Q(REG2_REG_7_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(clock), .D(n858), .Q(REG2_REG_8_));
DFFPOSX1 DFFPOSX1_192 ( .CLK(clock), .D(n863), .Q(REG2_REG_9_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(clock), .D(n868), .Q(REG2_REG_10_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(clock), .D(n873), .Q(REG2_REG_11_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(clock), .D(n878), .Q(REG2_REG_12_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(clock), .D(n883), .Q(REG2_REG_13_));
DFFPOSX1 DFFPOSX1_197 ( .CLK(clock), .D(n888), .Q(REG2_REG_14_));
DFFPOSX1 DFFPOSX1_198 ( .CLK(clock), .D(n893), .Q(REG2_REG_15_));
DFFPOSX1 DFFPOSX1_199 ( .CLK(clock), .D(n898), .Q(REG2_REG_16_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n986), .Q(ADDR_REG_17_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(n1054), .Q(ADDR_REG_0_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(clock), .D(n903), .Q(REG2_REG_17_));
DFFPOSX1 DFFPOSX1_201 ( .CLK(clock), .D(n908), .Q(REG2_REG_18_));
DFFPOSX1 DFFPOSX1_202 ( .CLK(clock), .D(n913), .Q(REG2_REG_19_));
DFFPOSX1 DFFPOSX1_203 ( .CLK(clock), .D(n918), .Q(REG2_REG_20_));
DFFPOSX1 DFFPOSX1_204 ( .CLK(clock), .D(n923), .Q(REG2_REG_21_));
DFFPOSX1 DFFPOSX1_205 ( .CLK(clock), .D(n928), .Q(REG2_REG_22_));
DFFPOSX1 DFFPOSX1_206 ( .CLK(clock), .D(n933), .Q(REG2_REG_23_));
DFFPOSX1 DFFPOSX1_207 ( .CLK(clock), .D(n938), .Q(REG2_REG_24_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(clock), .D(n943), .Q(REG2_REG_25_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(clock), .D(n948), .Q(REG2_REG_26_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(n1182), .Q(DATAO_REG_31_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(clock), .D(n953), .Q(REG2_REG_27_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(clock), .D(n958), .Q(REG2_REG_28_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(clock), .D(n963), .Q(REG2_REG_29_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(clock), .D(n968), .Q(REG2_REG_30_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(clock), .D(n973), .Q(REG2_REG_31_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(clock), .D(n1186), .Q(B_REG));
DFFPOSX1 DFFPOSX1_216 ( .CLK(clock), .D(n1191), .Q(REG3_REG_15_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(clock), .D(n1196), .Q(REG3_REG_26_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(clock), .D(n1201), .Q(REG3_REG_6_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(clock), .D(n1206), .Q(REG3_REG_18_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(n1178), .Q(DATAO_REG_30_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(clock), .D(n1211), .Q(REG3_REG_2_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(clock), .D(n1216), .Q(REG3_REG_11_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(clock), .D(n1221), .Q(REG3_REG_22_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(clock), .D(n1226), .Q(REG3_REG_13_));
DFFPOSX1 DFFPOSX1_224 ( .CLK(clock), .D(n1231), .Q(REG3_REG_20_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(clock), .D(n1236), .Q(REG3_REG_0_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(clock), .D(n1241), .Q(REG3_REG_9_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(clock), .D(n1246), .Q(REG3_REG_4_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(clock), .D(n1251), .Q(REG3_REG_24_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(clock), .D(n1256), .Q(REG3_REG_17_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(n1174), .Q(DATAO_REG_29_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(clock), .D(n1261), .Q(REG3_REG_5_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(clock), .D(n1266), .Q(REG3_REG_16_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(clock), .D(n1271), .Q(REG3_REG_25_));
DFFPOSX1 DFFPOSX1_233 ( .CLK(clock), .D(n1276), .Q(REG3_REG_12_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(clock), .D(n1281), .Q(REG3_REG_21_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(clock), .D(n1286), .Q(REG3_REG_1_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(clock), .D(n1291), .Q(REG3_REG_8_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(clock), .D(n1296), .Q(REG3_REG_28_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(clock), .D(n1301), .Q(REG3_REG_19_));
DFFPOSX1 DFFPOSX1_239 ( .CLK(clock), .D(n1306), .Q(REG3_REG_3_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(n1170), .Q(DATAO_REG_28_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(clock), .D(n1311), .Q(REG3_REG_10_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(clock), .D(n1316), .Q(REG3_REG_23_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(clock), .D(n1321), .Q(REG3_REG_14_));
DFFPOSX1 DFFPOSX1_243 ( .CLK(clock), .D(n1326), .Q(REG3_REG_27_));
DFFPOSX1 DFFPOSX1_244 ( .CLK(clock), .D(n1331), .Q(REG3_REG_7_));
DFFPOSX1 DFFPOSX1_245 ( .CLK(clock), .D(n1336), .Q(STATE_REG));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(n1166), .Q(DATAO_REG_27_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(n1162), .Q(DATAO_REG_26_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(n1158), .Q(DATAO_REG_25_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(n1154), .Q(DATAO_REG_24_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock), .D(n1150), .Q(DATAO_REG_23_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n998), .Q(ADDR_REG_14_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock), .D(n1146), .Q(DATAO_REG_22_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock), .D(n1142), .Q(DATAO_REG_21_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock), .D(n1138), .Q(DATAO_REG_20_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clock), .D(n1134), .Q(DATAO_REG_19_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clock), .D(n1130), .Q(DATAO_REG_18_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clock), .D(n1126), .Q(DATAO_REG_17_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clock), .D(n1122), .Q(DATAO_REG_16_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clock), .D(n1118), .Q(DATAO_REG_15_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clock), .D(n1114), .Q(DATAO_REG_14_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clock), .D(n1110), .Q(DATAO_REG_13_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n990), .Q(ADDR_REG_16_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clock), .D(n1106), .Q(DATAO_REG_12_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clock), .D(n1102), .Q(DATAO_REG_11_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clock), .D(n1098), .Q(DATAO_REG_10_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clock), .D(n1094), .Q(DATAO_REG_9_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clock), .D(n1090), .Q(DATAO_REG_8_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clock), .D(n1086), .Q(DATAO_REG_7_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clock), .D(n1082), .Q(DATAO_REG_6_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clock), .D(n1078), .Q(DATAO_REG_5_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clock), .D(n1074), .Q(DATAO_REG_4_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock), .D(n1070), .Q(DATAO_REG_3_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n994), .Q(ADDR_REG_15_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock), .D(n1066), .Q(DATAO_REG_2_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock), .D(n1062), .Q(DATAO_REG_1_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clock), .D(n1058), .Q(DATAO_REG_0_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clock), .D(n1341), .Q(RD_REG));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clock), .D(n1345), .Q(WR_REG));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clock), .D(n178), .Q(IR_REG_0_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clock), .D(n183), .Q(IR_REG_1_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clock), .D(n188), .Q(IR_REG_2_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clock), .D(n193), .Q(IR_REG_3_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clock), .D(n198), .Q(IR_REG_4_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n982), .Q(ADDR_REG_18_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clock), .D(n203), .Q(IR_REG_5_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clock), .D(n208), .Q(IR_REG_6_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clock), .D(n213), .Q(IR_REG_7_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clock), .D(n218), .Q(IR_REG_8_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clock), .D(n223), .Q(IR_REG_9_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clock), .D(n228), .Q(IR_REG_10_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clock), .D(n233), .Q(IR_REG_11_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clock), .D(n238), .Q(IR_REG_12_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clock), .D(n243), .Q(IR_REG_13_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clock), .D(n248), .Q(IR_REG_14_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n1002), .Q(ADDR_REG_13_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clock), .D(n253), .Q(IR_REG_15_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clock), .D(n258), .Q(IR_REG_16_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clock), .D(n263), .Q(IR_REG_17_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clock), .D(n268), .Q(IR_REG_18_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clock), .D(n273), .Q(IR_REG_19_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clock), .D(n278), .Q(IR_REG_20_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clock), .D(n283), .Q(IR_REG_21_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clock), .D(n288), .Q(IR_REG_22_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clock), .D(n293), .Q(IR_REG_23_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clock), .D(n298), .Q(IR_REG_24_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n1006), .Q(ADDR_REG_12_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clock), .D(n303), .Q(IR_REG_25_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(clock), .D(n308), .Q(IR_REG_26_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(clock), .D(n313), .Q(IR_REG_27_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(clock), .D(n318), .Q(IR_REG_28_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(clock), .D(n323), .Q(IR_REG_29_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(clock), .D(n328), .Q(IR_REG_30_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(clock), .D(n333), .Q(IR_REG_31_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(clock), .D(n338), .Q(D_REG_0_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(clock), .D(n343), .Q(D_REG_1_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(clock), .D(n348), .Q(D_REG_2_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(n1010), .Q(ADDR_REG_11_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(clock), .D(n353), .Q(D_REG_3_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(clock), .D(n358), .Q(D_REG_4_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(clock), .D(n363), .Q(D_REG_5_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(clock), .D(n368), .Q(D_REG_6_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(clock), .D(n373), .Q(D_REG_7_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(clock), .D(n378), .Q(D_REG_8_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(clock), .D(n383), .Q(D_REG_9_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(clock), .D(n388), .Q(D_REG_10_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(clock), .D(n393), .Q(D_REG_11_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(clock), .D(n398), .Q(D_REG_12_));
INVX1 INVX1_1 ( .A(IR_REG_24_), .Y(_abc_40319_new_n523_));
INVX1 INVX1_10 ( .A(_abc_40319_new_n555_), .Y(_abc_40319_new_n556_));
INVX1 INVX1_100 ( .A(_abc_40319_new_n993_), .Y(_abc_40319_new_n994_));
INVX1 INVX1_101 ( .A(_abc_40319_new_n995_), .Y(_abc_40319_new_n996_));
INVX1 INVX1_102 ( .A(_abc_40319_new_n1000_), .Y(_abc_40319_new_n1001_));
INVX1 INVX1_103 ( .A(_abc_40319_new_n1002_), .Y(_abc_40319_new_n1003_));
INVX1 INVX1_104 ( .A(_abc_40319_new_n1006_), .Y(_abc_40319_new_n1007_));
INVX1 INVX1_105 ( .A(_abc_40319_new_n1008_), .Y(_abc_40319_new_n1009_));
INVX1 INVX1_106 ( .A(n1336), .Y(_abc_40319_new_n1011_));
INVX1 INVX1_107 ( .A(_abc_40319_new_n1017_), .Y(_abc_40319_new_n1018_));
INVX1 INVX1_108 ( .A(REG3_REG_26_), .Y(_abc_40319_new_n1019_));
INVX1 INVX1_109 ( .A(REG3_REG_27_), .Y(_abc_40319_new_n1020_));
INVX1 INVX1_11 ( .A(IR_REG_31_), .Y(_abc_40319_new_n568_));
INVX1 INVX1_110 ( .A(REG3_REG_23_), .Y(_abc_40319_new_n1021_));
INVX1 INVX1_111 ( .A(REG3_REG_19_), .Y(_abc_40319_new_n1022_));
INVX1 INVX1_112 ( .A(REG3_REG_10_), .Y(_abc_40319_new_n1023_));
INVX1 INVX1_113 ( .A(REG3_REG_11_), .Y(_abc_40319_new_n1024_));
INVX1 INVX1_114 ( .A(REG2_REG_27_), .Y(_abc_40319_new_n1042_));
INVX1 INVX1_115 ( .A(_abc_40319_new_n1051_), .Y(_abc_40319_new_n1052_));
INVX1 INVX1_116 ( .A(_abc_40319_new_n1054_), .Y(_abc_40319_new_n1055_));
INVX1 INVX1_117 ( .A(REG3_REG_25_), .Y(_abc_40319_new_n1057_));
INVX1 INVX1_118 ( .A(REG0_REG_26_), .Y(_abc_40319_new_n1061_));
INVX1 INVX1_119 ( .A(REG0_REG_25_), .Y(_abc_40319_new_n1073_));
INVX1 INVX1_12 ( .A(_abc_40319_new_n571_), .Y(_abc_40319_new_n572_));
INVX1 INVX1_120 ( .A(_abc_40319_new_n1077_), .Y(_abc_40319_new_n1078_));
INVX1 INVX1_121 ( .A(_abc_40319_new_n1070_), .Y(_abc_40319_new_n1080_));
INVX1 INVX1_122 ( .A(_abc_40319_new_n1084_), .Y(_abc_40319_new_n1085_));
INVX1 INVX1_123 ( .A(REG3_REG_24_), .Y(_abc_40319_new_n1086_));
INVX1 INVX1_124 ( .A(REG0_REG_24_), .Y(_abc_40319_new_n1089_));
INVX1 INVX1_125 ( .A(_abc_40319_new_n1093_), .Y(_abc_40319_new_n1094_));
INVX1 INVX1_126 ( .A(_abc_40319_new_n813_), .Y(_abc_40319_new_n1096_));
INVX1 INVX1_127 ( .A(_abc_40319_new_n1098_), .Y(_abc_40319_new_n1099_));
INVX1 INVX1_128 ( .A(_abc_40319_new_n1100_), .Y(_abc_40319_new_n1101_));
INVX1 INVX1_129 ( .A(_abc_40319_new_n1103_), .Y(_abc_40319_new_n1104_));
INVX1 INVX1_13 ( .A(IR_REG_23_), .Y(_abc_40319_new_n575_));
INVX1 INVX1_130 ( .A(_abc_40319_new_n1108_), .Y(_abc_40319_new_n1109_));
INVX1 INVX1_131 ( .A(REG2_REG_23_), .Y(_abc_40319_new_n1111_));
INVX1 INVX1_132 ( .A(_abc_40319_new_n1118_), .Y(_abc_40319_new_n1119_));
INVX1 INVX1_133 ( .A(_abc_40319_new_n1122_), .Y(_abc_40319_new_n1123_));
INVX1 INVX1_134 ( .A(REG3_REG_21_), .Y(_abc_40319_new_n1124_));
INVX1 INVX1_135 ( .A(REG3_REG_22_), .Y(_abc_40319_new_n1125_));
INVX1 INVX1_136 ( .A(REG0_REG_22_), .Y(_abc_40319_new_n1130_));
INVX1 INVX1_137 ( .A(_abc_40319_new_n1139_), .Y(_abc_40319_new_n1140_));
INVX1 INVX1_138 ( .A(_abc_40319_new_n1142_), .Y(_abc_40319_new_n1143_));
INVX1 INVX1_139 ( .A(REG1_REG_18_), .Y(_abc_40319_new_n1149_));
INVX1 INVX1_14 ( .A(_abc_40319_new_n582_), .Y(_abc_40319_new_n583_));
INVX1 INVX1_140 ( .A(REG3_REG_18_), .Y(_abc_40319_new_n1151_));
INVX1 INVX1_141 ( .A(_abc_40319_new_n1156_), .Y(_abc_40319_new_n1157_));
INVX1 INVX1_142 ( .A(_abc_40319_new_n1148_), .Y(_abc_40319_new_n1159_));
INVX1 INVX1_143 ( .A(_abc_40319_new_n1161_), .Y(_abc_40319_new_n1162_));
INVX1 INVX1_144 ( .A(_abc_40319_new_n1164_), .Y(_abc_40319_new_n1165_));
INVX1 INVX1_145 ( .A(_abc_40319_new_n1166_), .Y(_abc_40319_new_n1167_));
INVX1 INVX1_146 ( .A(_abc_40319_new_n1168_), .Y(_abc_40319_new_n1169_));
INVX1 INVX1_147 ( .A(REG2_REG_16_), .Y(_abc_40319_new_n1176_));
INVX1 INVX1_148 ( .A(REG1_REG_16_), .Y(_abc_40319_new_n1179_));
INVX1 INVX1_149 ( .A(REG3_REG_16_), .Y(_abc_40319_new_n1184_));
INVX1 INVX1_15 ( .A(IR_REG_26_), .Y(_abc_40319_new_n588_));
INVX1 INVX1_150 ( .A(_abc_40319_new_n1186_), .Y(_abc_40319_new_n1187_));
INVX1 INVX1_151 ( .A(_abc_40319_new_n1190_), .Y(_abc_40319_new_n1191_));
INVX1 INVX1_152 ( .A(REG1_REG_17_), .Y(_abc_40319_new_n1199_));
INVX1 INVX1_153 ( .A(REG0_REG_17_), .Y(_abc_40319_new_n1200_));
INVX1 INVX1_154 ( .A(REG2_REG_17_), .Y(_abc_40319_new_n1202_));
INVX1 INVX1_155 ( .A(REG3_REG_17_), .Y(_abc_40319_new_n1203_));
INVX1 INVX1_156 ( .A(_abc_40319_new_n1185_), .Y(_abc_40319_new_n1204_));
INVX1 INVX1_157 ( .A(_abc_40319_new_n1205_), .Y(_abc_40319_new_n1206_));
INVX1 INVX1_158 ( .A(_abc_40319_new_n1208_), .Y(_abc_40319_new_n1209_));
INVX1 INVX1_159 ( .A(_abc_40319_new_n1198_), .Y(_abc_40319_new_n1211_));
INVX1 INVX1_16 ( .A(IR_REG_18_), .Y(_abc_40319_new_n594_));
INVX1 INVX1_160 ( .A(_abc_40319_new_n1213_), .Y(_abc_40319_new_n1214_));
INVX1 INVX1_161 ( .A(_abc_40319_new_n1216_), .Y(_abc_40319_new_n1217_));
INVX1 INVX1_162 ( .A(REG1_REG_15_), .Y(_abc_40319_new_n1224_));
INVX1 INVX1_163 ( .A(REG2_REG_15_), .Y(_abc_40319_new_n1225_));
INVX1 INVX1_164 ( .A(REG0_REG_15_), .Y(_abc_40319_new_n1227_));
INVX1 INVX1_165 ( .A(REG3_REG_15_), .Y(_abc_40319_new_n1228_));
INVX1 INVX1_166 ( .A(_abc_40319_new_n1236_), .Y(_abc_40319_new_n1237_));
INVX1 INVX1_167 ( .A(_abc_40319_new_n1239_), .Y(_abc_40319_new_n1240_));
INVX1 INVX1_168 ( .A(_abc_40319_new_n1242_), .Y(_abc_40319_new_n1243_));
INVX1 INVX1_169 ( .A(_abc_40319_new_n1245_), .Y(_abc_40319_new_n1246_));
INVX1 INVX1_17 ( .A(_abc_40319_new_n608_), .Y(_abc_40319_new_n609_));
INVX1 INVX1_170 ( .A(REG2_REG_14_), .Y(_abc_40319_new_n1249_));
INVX1 INVX1_171 ( .A(REG0_REG_14_), .Y(_abc_40319_new_n1250_));
INVX1 INVX1_172 ( .A(REG1_REG_14_), .Y(_abc_40319_new_n1252_));
INVX1 INVX1_173 ( .A(REG3_REG_14_), .Y(_abc_40319_new_n1253_));
INVX1 INVX1_174 ( .A(_abc_40319_new_n1258_), .Y(_abc_40319_new_n1259_));
INVX1 INVX1_175 ( .A(_abc_40319_new_n1248_), .Y(_abc_40319_new_n1261_));
INVX1 INVX1_176 ( .A(_abc_40319_new_n1263_), .Y(_abc_40319_new_n1264_));
INVX1 INVX1_177 ( .A(_abc_40319_new_n1267_), .Y(_abc_40319_new_n1268_));
INVX1 INVX1_178 ( .A(_abc_40319_new_n1270_), .Y(_abc_40319_new_n1271_));
INVX1 INVX1_179 ( .A(_abc_40319_new_n1273_), .Y(_abc_40319_new_n1274_));
INVX1 INVX1_18 ( .A(_abc_40319_new_n615_), .Y(_abc_40319_new_n616_));
INVX1 INVX1_180 ( .A(IR_REG_9_), .Y(_abc_40319_new_n1289_));
INVX1 INVX1_181 ( .A(_abc_40319_new_n1294_), .Y(_abc_40319_new_n1295_));
INVX1 INVX1_182 ( .A(REG1_REG_9_), .Y(_abc_40319_new_n1298_));
INVX1 INVX1_183 ( .A(REG3_REG_9_), .Y(_abc_40319_new_n1300_));
INVX1 INVX1_184 ( .A(REG2_REG_9_), .Y(_abc_40319_new_n1305_));
INVX1 INVX1_185 ( .A(REG0_REG_9_), .Y(_abc_40319_new_n1306_));
INVX1 INVX1_186 ( .A(_abc_40319_new_n1308_), .Y(_abc_40319_new_n1309_));
INVX1 INVX1_187 ( .A(_abc_40319_new_n1311_), .Y(_abc_40319_new_n1312_));
INVX1 INVX1_188 ( .A(_abc_40319_new_n1315_), .Y(_abc_40319_new_n1316_));
INVX1 INVX1_189 ( .A(_abc_40319_new_n530_), .Y(_abc_40319_new_n1318_));
INVX1 INVX1_19 ( .A(STATE_REG), .Y(_abc_40319_new_n618_));
INVX1 INVX1_190 ( .A(_abc_40319_new_n1322_), .Y(_abc_40319_new_n1323_));
INVX1 INVX1_191 ( .A(REG1_REG_13_), .Y(_abc_40319_new_n1326_));
INVX1 INVX1_192 ( .A(REG3_REG_12_), .Y(_abc_40319_new_n1327_));
INVX1 INVX1_193 ( .A(REG3_REG_13_), .Y(_abc_40319_new_n1328_));
INVX1 INVX1_194 ( .A(_abc_40319_new_n1330_), .Y(_abc_40319_new_n1331_));
INVX1 INVX1_195 ( .A(REG2_REG_13_), .Y(_abc_40319_new_n1333_));
INVX1 INVX1_196 ( .A(REG0_REG_13_), .Y(_abc_40319_new_n1334_));
INVX1 INVX1_197 ( .A(_abc_40319_new_n603_), .Y(_abc_40319_new_n1341_));
INVX1 INVX1_198 ( .A(_abc_40319_new_n1343_), .Y(_abc_40319_new_n1344_));
INVX1 INVX1_199 ( .A(DATAI_12_), .Y(_abc_40319_new_n1350_));
INVX1 INVX1_2 ( .A(IR_REG_3_), .Y(_abc_40319_new_n524_));
INVX1 INVX1_20 ( .A(nRESET_G), .Y(_abc_40319_new_n619_));
INVX1 INVX1_200 ( .A(REG1_REG_12_), .Y(_abc_40319_new_n1353_));
INVX1 INVX1_201 ( .A(REG2_REG_12_), .Y(_abc_40319_new_n1354_));
INVX1 INVX1_202 ( .A(REG0_REG_12_), .Y(_abc_40319_new_n1356_));
INVX1 INVX1_203 ( .A(IR_REG_11_), .Y(_abc_40319_new_n1366_));
INVX1 INVX1_204 ( .A(_abc_40319_new_n1370_), .Y(_abc_40319_new_n1371_));
INVX1 INVX1_205 ( .A(REG1_REG_11_), .Y(_abc_40319_new_n1372_));
INVX1 INVX1_206 ( .A(REG2_REG_11_), .Y(_abc_40319_new_n1373_));
INVX1 INVX1_207 ( .A(_abc_40319_new_n1379_), .Y(_abc_40319_new_n1380_));
INVX1 INVX1_208 ( .A(_abc_40319_new_n1381_), .Y(_abc_40319_new_n1382_));
INVX1 INVX1_209 ( .A(_abc_40319_new_n1385_), .Y(_abc_40319_new_n1386_));
INVX1 INVX1_21 ( .A(_abc_40319_new_n567_), .Y(_abc_40319_new_n622_));
INVX1 INVX1_210 ( .A(_abc_40319_new_n1390_), .Y(_abc_40319_new_n1391_));
INVX1 INVX1_211 ( .A(REG1_REG_10_), .Y(_abc_40319_new_n1394_));
INVX1 INVX1_212 ( .A(REG0_REG_10_), .Y(_abc_40319_new_n1397_));
INVX1 INVX1_213 ( .A(_abc_40319_new_n1398_), .Y(_abc_40319_new_n1399_));
INVX1 INVX1_214 ( .A(_abc_40319_new_n1401_), .Y(_abc_40319_new_n1402_));
INVX1 INVX1_215 ( .A(_abc_40319_new_n1403_), .Y(_abc_40319_new_n1404_));
INVX1 INVX1_216 ( .A(_abc_40319_new_n1408_), .Y(_abc_40319_new_n1409_));
INVX1 INVX1_217 ( .A(_abc_40319_new_n1410_), .Y(_abc_40319_new_n1411_));
INVX1 INVX1_218 ( .A(_abc_40319_new_n1413_), .Y(_abc_40319_new_n1414_));
INVX1 INVX1_219 ( .A(_abc_40319_new_n1415_), .Y(_abc_40319_new_n1416_));
INVX1 INVX1_22 ( .A(_abc_40319_new_n560_), .Y(_abc_40319_new_n623_));
INVX1 INVX1_220 ( .A(_abc_40319_new_n1423_), .Y(_abc_40319_new_n1424_));
INVX1 INVX1_221 ( .A(REG1_REG_19_), .Y(_abc_40319_new_n1430_));
INVX1 INVX1_222 ( .A(_abc_40319_new_n1438_), .Y(_abc_40319_new_n1439_));
INVX1 INVX1_223 ( .A(_abc_40319_new_n1442_), .Y(_abc_40319_new_n1443_));
INVX1 INVX1_224 ( .A(REG3_REG_20_), .Y(_abc_40319_new_n1444_));
INVX1 INVX1_225 ( .A(_abc_40319_new_n1453_), .Y(_abc_40319_new_n1454_));
INVX1 INVX1_226 ( .A(_abc_40319_new_n1457_), .Y(_abc_40319_new_n1458_));
INVX1 INVX1_227 ( .A(_abc_40319_new_n1459_), .Y(_abc_40319_new_n1460_));
INVX1 INVX1_228 ( .A(_abc_40319_new_n1470_), .Y(_abc_40319_new_n1471_));
INVX1 INVX1_229 ( .A(_abc_40319_new_n1473_), .Y(_abc_40319_new_n1474_));
INVX1 INVX1_23 ( .A(_abc_40319_new_n627_), .Y(_abc_40319_new_n628_));
INVX1 INVX1_230 ( .A(_abc_40319_new_n1475_), .Y(_abc_40319_new_n1476_));
INVX1 INVX1_231 ( .A(_abc_40319_new_n1477_), .Y(_abc_40319_new_n1478_));
INVX1 INVX1_232 ( .A(_abc_40319_new_n1482_), .Y(_abc_40319_new_n1483_));
INVX1 INVX1_233 ( .A(_abc_40319_new_n1489_), .Y(_abc_40319_new_n1490_));
INVX1 INVX1_234 ( .A(_abc_40319_new_n1065_), .Y(_abc_40319_new_n1496_));
INVX1 INVX1_235 ( .A(REG2_REG_28_), .Y(_abc_40319_new_n1500_));
INVX1 INVX1_236 ( .A(_abc_40319_new_n1503_), .Y(_abc_40319_new_n1504_));
INVX1 INVX1_237 ( .A(_abc_40319_new_n1233_), .Y(_abc_40319_new_n1516_));
INVX1 INVX1_238 ( .A(_abc_40319_new_n1010_), .Y(_abc_40319_new_n1519_));
INVX1 INVX1_239 ( .A(_abc_40319_new_n1393_), .Y(_abc_40319_new_n1541_));
INVX1 INVX1_24 ( .A(D_REG_0_), .Y(_abc_40319_new_n655_));
INVX1 INVX1_240 ( .A(_abc_40319_new_n901_), .Y(_abc_40319_new_n1548_));
INVX1 INVX1_241 ( .A(_abc_40319_new_n1549_), .Y(_abc_40319_new_n1550_));
INVX1 INVX1_242 ( .A(_abc_40319_new_n932_), .Y(_abc_40319_new_n1552_));
INVX1 INVX1_243 ( .A(_abc_40319_new_n809_), .Y(_abc_40319_new_n1556_));
INVX1 INVX1_244 ( .A(_abc_40319_new_n1452_), .Y(_abc_40319_new_n1567_));
INVX1 INVX1_245 ( .A(_abc_40319_new_n1429_), .Y(_abc_40319_new_n1570_));
INVX1 INVX1_246 ( .A(_abc_40319_new_n1571_), .Y(_abc_40319_new_n1572_));
INVX1 INVX1_247 ( .A(_abc_40319_new_n1505_), .Y(_abc_40319_new_n1580_));
INVX1 INVX1_248 ( .A(_abc_40319_new_n1581_), .Y(_abc_40319_new_n1582_));
INVX1 INVX1_249 ( .A(_abc_40319_new_n1586_), .Y(_abc_40319_new_n1589_));
INVX1 INVX1_25 ( .A(_abc_40319_new_n658_), .Y(_abc_40319_new_n659_));
INVX1 INVX1_250 ( .A(_abc_40319_new_n1046_), .Y(_abc_40319_new_n1592_));
INVX1 INVX1_251 ( .A(REG2_REG_29_), .Y(_abc_40319_new_n1594_));
INVX1 INVX1_252 ( .A(_abc_40319_new_n1607_), .Y(_abc_40319_new_n1608_));
INVX1 INVX1_253 ( .A(_abc_40319_new_n984_), .Y(_abc_40319_new_n1615_));
INVX1 INVX1_254 ( .A(REG3_REG_1_), .Y(_abc_40319_new_n1624_));
INVX1 INVX1_255 ( .A(_abc_40319_new_n1352_), .Y(_abc_40319_new_n1654_));
INVX1 INVX1_256 ( .A(_abc_40319_new_n1673_), .Y(_abc_40319_new_n1674_));
INVX1 INVX1_257 ( .A(_abc_40319_new_n1425_), .Y(_abc_40319_new_n1696_));
INVX1 INVX1_258 ( .A(_abc_40319_new_n1189_), .Y(_abc_40319_new_n1700_));
INVX1 INVX1_259 ( .A(_abc_40319_new_n1115_), .Y(_abc_40319_new_n1710_));
INVX1 INVX1_26 ( .A(_abc_40319_new_n669_), .Y(_abc_40319_new_n670_));
INVX1 INVX1_260 ( .A(_abc_40319_new_n1713_), .Y(_abc_40319_new_n1714_));
INVX1 INVX1_261 ( .A(_abc_40319_new_n799_), .Y(_abc_40319_new_n1726_));
INVX1 INVX1_262 ( .A(_abc_40319_new_n1727_), .Y(_abc_40319_new_n1728_));
INVX1 INVX1_263 ( .A(_abc_40319_new_n1313_), .Y(_abc_40319_new_n1732_));
INVX1 INVX1_264 ( .A(_abc_40319_new_n1297_), .Y(_abc_40319_new_n1739_));
INVX1 INVX1_265 ( .A(_abc_40319_new_n1740_), .Y(_abc_40319_new_n1741_));
INVX1 INVX1_266 ( .A(_abc_40319_new_n1748_), .Y(_abc_40319_new_n1749_));
INVX1 INVX1_267 ( .A(REG3_REG_0_), .Y(_abc_40319_new_n1750_));
INVX1 INVX1_268 ( .A(_abc_40319_new_n1437_), .Y(_abc_40319_new_n1759_));
INVX1 INVX1_269 ( .A(_abc_40319_new_n1648_), .Y(_abc_40319_new_n1767_));
INVX1 INVX1_27 ( .A(_abc_40319_new_n672_), .Y(_abc_40319_new_n673_));
INVX1 INVX1_270 ( .A(_abc_40319_new_n1782_), .Y(_abc_40319_new_n1783_));
INVX1 INVX1_271 ( .A(_abc_40319_new_n1360_), .Y(_abc_40319_new_n1796_));
INVX1 INVX1_272 ( .A(_abc_40319_new_n1377_), .Y(_abc_40319_new_n1799_));
INVX1 INVX1_273 ( .A(REG3_REG_2_), .Y(_abc_40319_new_n1812_));
INVX1 INVX1_274 ( .A(_abc_40319_new_n1813_), .Y(_abc_40319_new_n1814_));
INVX1 INVX1_275 ( .A(_abc_40319_new_n1153_), .Y(_abc_40319_new_n1824_));
INVX1 INVX1_276 ( .A(_abc_40319_new_n1825_), .Y(_abc_40319_new_n1826_));
INVX1 INVX1_277 ( .A(_abc_40319_new_n963_), .Y(_abc_40319_new_n1830_));
INVX1 INVX1_278 ( .A(_abc_40319_new_n1102_), .Y(_abc_40319_new_n1846_));
INVX1 INVX1_279 ( .A(_abc_40319_new_n1223_), .Y(_abc_40319_new_n1865_));
INVX1 INVX1_28 ( .A(_abc_40319_new_n676_), .Y(_abc_40319_new_n677_));
INVX1 INVX1_280 ( .A(_abc_40319_new_n580_), .Y(_abc_40319_new_n1870_));
INVX1 INVX1_281 ( .A(_abc_40319_new_n1871_), .Y(_abc_40319_new_n1872_));
INVX1 INVX1_282 ( .A(_abc_40319_new_n1873_), .Y(_abc_40319_new_n1874_));
INVX1 INVX1_283 ( .A(_abc_40319_new_n1876_), .Y(_abc_40319_new_n1877_));
INVX1 INVX1_284 ( .A(REG0_REG_31_), .Y(_abc_40319_new_n1879_));
INVX1 INVX1_285 ( .A(_abc_40319_new_n1882_), .Y(_abc_40319_new_n1883_));
INVX1 INVX1_286 ( .A(_abc_40319_new_n1884_), .Y(_abc_40319_new_n1885_));
INVX1 INVX1_287 ( .A(_abc_40319_new_n1894_), .Y(_abc_40319_new_n1895_));
INVX1 INVX1_288 ( .A(_abc_40319_new_n1896_), .Y(_abc_40319_new_n1897_));
INVX1 INVX1_289 ( .A(_abc_40319_new_n1914_), .Y(_abc_40319_new_n1915_));
INVX1 INVX1_29 ( .A(IR_REG_7_), .Y(_abc_40319_new_n684_));
INVX1 INVX1_290 ( .A(_abc_40319_new_n769_), .Y(_abc_40319_new_n1938_));
INVX1 INVX1_291 ( .A(_abc_40319_new_n1941_), .Y(_abc_40319_new_n1942_));
INVX1 INVX1_292 ( .A(_abc_40319_new_n1951_), .Y(_abc_40319_new_n1952_));
INVX1 INVX1_293 ( .A(_abc_40319_new_n1953_), .Y(_abc_40319_new_n1954_));
INVX1 INVX1_294 ( .A(_abc_40319_new_n985_), .Y(_abc_40319_new_n1957_));
INVX1 INVX1_295 ( .A(_abc_40319_new_n986_), .Y(_abc_40319_new_n1958_));
INVX1 INVX1_296 ( .A(_abc_40319_new_n1967_), .Y(_abc_40319_new_n1968_));
INVX1 INVX1_297 ( .A(_abc_40319_new_n2003_), .Y(_abc_40319_new_n2004_));
INVX1 INVX1_298 ( .A(_abc_40319_new_n2015_), .Y(_abc_40319_new_n2016_));
INVX1 INVX1_299 ( .A(_abc_40319_new_n2030_), .Y(_abc_40319_new_n2031_));
INVX1 INVX1_3 ( .A(IR_REG_16_), .Y(_abc_40319_new_n533_));
INVX1 INVX1_30 ( .A(IR_REG_6_), .Y(_abc_40319_new_n685_));
INVX1 INVX1_300 ( .A(_abc_40319_new_n2032_), .Y(_abc_40319_new_n2035_));
INVX1 INVX1_301 ( .A(_abc_40319_new_n2051_), .Y(_abc_40319_new_n2052_));
INVX1 INVX1_302 ( .A(_abc_40319_new_n2058_), .Y(_abc_40319_new_n2059_));
INVX1 INVX1_303 ( .A(_abc_40319_new_n2061_), .Y(_abc_40319_new_n2062_));
INVX1 INVX1_304 ( .A(_abc_40319_new_n2070_), .Y(_abc_40319_new_n2071_));
INVX1 INVX1_305 ( .A(_abc_40319_new_n2072_), .Y(_abc_40319_new_n2073_));
INVX1 INVX1_306 ( .A(_abc_40319_new_n2069_), .Y(_abc_40319_new_n2074_));
INVX1 INVX1_307 ( .A(_abc_40319_new_n2081_), .Y(_abc_40319_new_n2082_));
INVX1 INVX1_308 ( .A(_abc_40319_new_n2083_), .Y(_abc_40319_new_n2084_));
INVX1 INVX1_309 ( .A(_abc_40319_new_n2085_), .Y(_abc_40319_new_n2086_));
INVX1 INVX1_31 ( .A(_abc_40319_new_n690_), .Y(_abc_40319_new_n691_));
INVX1 INVX1_310 ( .A(_abc_40319_new_n2091_), .Y(_abc_40319_new_n2094_));
INVX1 INVX1_311 ( .A(_abc_40319_new_n2092_), .Y(_abc_40319_new_n2095_));
INVX1 INVX1_312 ( .A(_abc_40319_new_n2096_), .Y(_abc_40319_new_n2097_));
INVX1 INVX1_313 ( .A(REG0_REG_30_), .Y(_abc_40319_new_n2099_));
INVX1 INVX1_314 ( .A(_abc_40319_new_n2102_), .Y(_abc_40319_new_n2103_));
INVX1 INVX1_315 ( .A(_abc_40319_new_n2104_), .Y(_abc_40319_new_n2105_));
INVX1 INVX1_316 ( .A(_abc_40319_new_n2108_), .Y(_abc_40319_new_n2109_));
INVX1 INVX1_317 ( .A(_abc_40319_new_n2110_), .Y(_abc_40319_new_n2111_));
INVX1 INVX1_318 ( .A(_abc_40319_new_n2116_), .Y(_abc_40319_new_n2117_));
INVX1 INVX1_319 ( .A(_abc_40319_new_n2120_), .Y(_abc_40319_new_n2121_));
INVX1 INVX1_32 ( .A(IR_REG_30_), .Y(_abc_40319_new_n699_));
INVX1 INVX1_320 ( .A(DATAI_26_), .Y(_abc_40319_new_n2122_));
INVX1 INVX1_321 ( .A(DATAI_25_), .Y(_abc_40319_new_n2126_));
INVX1 INVX1_322 ( .A(_abc_40319_new_n2129_), .Y(_abc_40319_new_n2130_));
INVX1 INVX1_323 ( .A(_abc_40319_new_n2131_), .Y(_abc_40319_new_n2132_));
INVX1 INVX1_324 ( .A(DATAI_23_), .Y(_abc_40319_new_n2136_));
INVX1 INVX1_325 ( .A(_abc_40319_new_n2138_), .Y(_abc_40319_new_n2139_));
INVX1 INVX1_326 ( .A(_abc_40319_new_n2140_), .Y(_abc_40319_new_n2141_));
INVX1 INVX1_327 ( .A(_abc_40319_new_n2145_), .Y(_abc_40319_new_n2146_));
INVX1 INVX1_328 ( .A(_abc_40319_new_n2149_), .Y(_abc_40319_new_n2150_));
INVX1 INVX1_329 ( .A(_abc_40319_new_n2152_), .Y(_abc_40319_new_n2153_));
INVX1 INVX1_33 ( .A(_abc_40319_new_n701_), .Y(_abc_40319_new_n705_));
INVX1 INVX1_330 ( .A(_abc_40319_new_n2162_), .Y(_abc_40319_new_n2163_));
INVX1 INVX1_331 ( .A(_abc_40319_new_n2164_), .Y(_abc_40319_new_n2165_));
INVX1 INVX1_332 ( .A(_abc_40319_new_n2167_), .Y(_abc_40319_new_n2168_));
INVX1 INVX1_333 ( .A(_abc_40319_new_n2169_), .Y(_abc_40319_new_n2170_));
INVX1 INVX1_334 ( .A(_abc_40319_new_n2173_), .Y(_abc_40319_new_n2174_));
INVX1 INVX1_335 ( .A(_abc_40319_new_n2178_), .Y(_abc_40319_new_n2179_));
INVX1 INVX1_336 ( .A(_abc_40319_new_n2183_), .Y(_abc_40319_new_n2184_));
INVX1 INVX1_337 ( .A(_abc_40319_new_n2185_), .Y(_abc_40319_new_n2186_));
INVX1 INVX1_338 ( .A(_abc_40319_new_n2187_), .Y(_abc_40319_new_n2188_));
INVX1 INVX1_339 ( .A(_abc_40319_new_n2192_), .Y(_abc_40319_new_n2193_));
INVX1 INVX1_34 ( .A(_abc_40319_new_n711_), .Y(_abc_40319_new_n712_));
INVX1 INVX1_340 ( .A(_abc_40319_new_n1175_), .Y(_abc_40319_new_n2196_));
INVX1 INVX1_341 ( .A(_abc_40319_new_n2202_), .Y(_abc_40319_new_n2203_));
INVX1 INVX1_342 ( .A(_abc_40319_new_n2205_), .Y(_abc_40319_new_n2206_));
INVX1 INVX1_343 ( .A(DATAI_22_), .Y(_abc_40319_new_n2213_));
INVX1 INVX1_344 ( .A(_abc_40319_new_n2217_), .Y(_abc_40319_new_n2218_));
INVX1 INVX1_345 ( .A(_abc_40319_new_n2222_), .Y(_abc_40319_new_n2223_));
INVX1 INVX1_346 ( .A(_abc_40319_new_n1325_), .Y(_abc_40319_new_n2228_));
INVX1 INVX1_347 ( .A(_abc_40319_new_n2230_), .Y(_abc_40319_new_n2231_));
INVX1 INVX1_348 ( .A(_abc_40319_new_n2233_), .Y(_abc_40319_new_n2234_));
INVX1 INVX1_349 ( .A(_abc_40319_new_n2239_), .Y(_abc_40319_new_n2240_));
INVX1 INVX1_35 ( .A(REG3_REG_6_), .Y(_abc_40319_new_n728_));
INVX1 INVX1_350 ( .A(_abc_40319_new_n944_), .Y(_abc_40319_new_n2246_));
INVX1 INVX1_351 ( .A(DATAI_27_), .Y(_abc_40319_new_n2258_));
INVX1 INVX1_352 ( .A(_abc_40319_new_n2088_), .Y(_abc_40319_new_n2262_));
INVX1 INVX1_353 ( .A(_abc_40319_new_n2266_), .Y(_abc_40319_new_n2267_));
INVX1 INVX1_354 ( .A(_abc_40319_new_n1956_), .Y(_abc_40319_new_n2284_));
INVX1 INVX1_355 ( .A(_abc_40319_new_n2026_), .Y(_abc_40319_new_n2294_));
INVX1 INVX1_356 ( .A(_abc_40319_new_n2039_), .Y(_abc_40319_new_n2296_));
INVX1 INVX1_357 ( .A(_abc_40319_new_n2049_), .Y(_abc_40319_new_n2298_));
INVX1 INVX1_358 ( .A(_abc_40319_new_n2093_), .Y(_abc_40319_new_n2303_));
INVX1 INVX1_359 ( .A(_abc_40319_new_n2113_), .Y(_abc_40319_new_n2305_));
INVX1 INVX1_36 ( .A(REG3_REG_3_), .Y(_abc_40319_new_n729_));
INVX1 INVX1_360 ( .A(_abc_40319_new_n2259_), .Y(_abc_40319_new_n2308_));
INVX1 INVX1_361 ( .A(_abc_40319_new_n2310_), .Y(_abc_40319_new_n2311_));
INVX1 INVX1_362 ( .A(_abc_40319_new_n2317_), .Y(_abc_40319_new_n2318_));
INVX1 INVX1_363 ( .A(_abc_40319_new_n2319_), .Y(_abc_40319_new_n2320_));
INVX1 INVX1_364 ( .A(_abc_40319_new_n2221_), .Y(_abc_40319_new_n2330_));
INVX1 INVX1_365 ( .A(_abc_40319_new_n2331_), .Y(_abc_40319_new_n2332_));
INVX1 INVX1_366 ( .A(_abc_40319_new_n2339_), .Y(_abc_40319_new_n2340_));
INVX1 INVX1_367 ( .A(_abc_40319_new_n2123_), .Y(_abc_40319_new_n2346_));
INVX1 INVX1_368 ( .A(_abc_40319_new_n2349_), .Y(_abc_40319_new_n2350_));
INVX1 INVX1_369 ( .A(_abc_40319_new_n2351_), .Y(_abc_40319_new_n2352_));
INVX1 INVX1_37 ( .A(REG3_REG_4_), .Y(_abc_40319_new_n730_));
INVX1 INVX1_370 ( .A(_abc_40319_new_n2312_), .Y(_abc_40319_new_n2353_));
INVX1 INVX1_371 ( .A(_abc_40319_new_n2359_), .Y(_abc_40319_new_n2360_));
INVX1 INVX1_372 ( .A(_abc_40319_new_n2355_), .Y(_abc_40319_new_n2370_));
INVX1 INVX1_373 ( .A(_abc_40319_new_n2334_), .Y(_abc_40319_new_n2373_));
INVX1 INVX1_374 ( .A(_abc_40319_new_n2219_), .Y(_abc_40319_new_n2380_));
INVX1 INVX1_375 ( .A(_abc_40319_new_n698_), .Y(_abc_40319_new_n2388_));
INVX1 INVX1_376 ( .A(_abc_40319_new_n2389_), .Y(_abc_40319_new_n2390_));
INVX1 INVX1_377 ( .A(_abc_40319_new_n2148_), .Y(_abc_40319_new_n2402_));
INVX1 INVX1_378 ( .A(_abc_40319_new_n2307_), .Y(_abc_40319_new_n2403_));
INVX1 INVX1_379 ( .A(_abc_40319_new_n2321_), .Y(_abc_40319_new_n2407_));
INVX1 INVX1_38 ( .A(REG3_REG_7_), .Y(_abc_40319_new_n735_));
INVX1 INVX1_380 ( .A(_abc_40319_new_n2144_), .Y(_abc_40319_new_n2426_));
INVX1 INVX1_381 ( .A(_abc_40319_new_n1276_), .Y(_abc_40319_new_n2427_));
INVX1 INVX1_382 ( .A(_abc_40319_new_n2438_), .Y(_abc_40319_new_n2444_));
INVX1 INVX1_383 ( .A(_abc_40319_new_n2446_), .Y(_abc_40319_new_n2447_));
INVX1 INVX1_384 ( .A(_abc_40319_new_n2124_), .Y(_abc_40319_new_n2454_));
INVX1 INVX1_385 ( .A(_abc_40319_new_n2127_), .Y(_abc_40319_new_n2455_));
INVX1 INVX1_386 ( .A(_abc_40319_new_n2133_), .Y(_abc_40319_new_n2456_));
INVX1 INVX1_387 ( .A(_abc_40319_new_n2473_), .Y(_abc_40319_new_n2474_));
INVX1 INVX1_388 ( .A(_abc_40319_new_n2377_), .Y(_abc_40319_new_n2484_));
INVX1 INVX1_389 ( .A(_abc_40319_new_n2486_), .Y(_abc_40319_new_n2487_));
INVX1 INVX1_39 ( .A(_abc_40319_new_n737_), .Y(_abc_40319_new_n738_));
INVX1 INVX1_390 ( .A(_abc_40319_new_n2490_), .Y(_abc_40319_new_n2491_));
INVX1 INVX1_391 ( .A(_abc_40319_new_n2494_), .Y(_abc_40319_new_n2495_));
INVX1 INVX1_392 ( .A(_abc_40319_new_n2406_), .Y(_abc_40319_new_n2499_));
INVX1 INVX1_393 ( .A(_abc_40319_new_n2404_), .Y(_abc_40319_new_n2506_));
INVX1 INVX1_394 ( .A(_abc_40319_new_n2512_), .Y(_abc_40319_new_n2513_));
INVX1 INVX1_395 ( .A(_abc_40319_new_n2519_), .Y(_abc_40319_new_n2520_));
INVX1 INVX1_396 ( .A(_abc_40319_new_n694_), .Y(_abc_40319_new_n2523_));
INVX1 INVX1_397 ( .A(_abc_40319_new_n2524_), .Y(_abc_40319_new_n2525_));
INVX1 INVX1_398 ( .A(_abc_40319_new_n2546_), .Y(_abc_40319_new_n2547_));
INVX1 INVX1_399 ( .A(_abc_40319_new_n2567_), .Y(_abc_40319_new_n2568_));
INVX1 INVX1_4 ( .A(IR_REG_17_), .Y(_abc_40319_new_n534_));
INVX1 INVX1_40 ( .A(_abc_40319_new_n614_), .Y(_abc_40319_new_n742_));
INVX1 INVX1_400 ( .A(_abc_40319_new_n2550_), .Y(_abc_40319_new_n2571_));
INVX1 INVX1_401 ( .A(_abc_40319_new_n2582_), .Y(_abc_40319_new_n2583_));
INVX1 INVX1_402 ( .A(_abc_40319_new_n2614_), .Y(_abc_40319_new_n2615_));
INVX1 INVX1_403 ( .A(_abc_40319_new_n2538_), .Y(_abc_40319_new_n2623_));
INVX1 INVX1_404 ( .A(_abc_40319_new_n2630_), .Y(_abc_40319_new_n2631_));
INVX1 INVX1_405 ( .A(REG2_REG_7_), .Y(_abc_40319_new_n2639_));
INVX1 INVX1_406 ( .A(_abc_40319_new_n2640_), .Y(_abc_40319_new_n2641_));
INVX1 INVX1_407 ( .A(_abc_40319_new_n942_), .Y(_abc_40319_new_n2642_));
INVX1 INVX1_408 ( .A(REG1_REG_7_), .Y(_abc_40319_new_n2653_));
INVX1 INVX1_409 ( .A(REG2_REG_8_), .Y(_abc_40319_new_n2663_));
INVX1 INVX1_41 ( .A(_abc_40319_new_n667_), .Y(_abc_40319_new_n749_));
INVX1 INVX1_410 ( .A(_abc_40319_new_n2665_), .Y(_abc_40319_new_n2667_));
INVX1 INVX1_411 ( .A(REG1_REG_8_), .Y(_abc_40319_new_n2672_));
INVX1 INVX1_412 ( .A(_abc_40319_new_n2683_), .Y(_abc_40319_new_n2684_));
INVX1 INVX1_413 ( .A(_abc_40319_new_n2542_), .Y(_abc_40319_new_n2686_));
INVX1 INVX1_414 ( .A(_abc_40319_new_n2688_), .Y(_abc_40319_new_n2689_));
INVX1 INVX1_415 ( .A(_abc_40319_new_n2664_), .Y(_abc_40319_new_n2697_));
INVX1 INVX1_416 ( .A(_abc_40319_new_n2700_), .Y(_abc_40319_new_n2701_));
INVX1 INVX1_417 ( .A(_abc_40319_new_n2543_), .Y(_abc_40319_new_n2711_));
INVX1 INVX1_418 ( .A(_abc_40319_new_n2725_), .Y(_abc_40319_new_n2726_));
INVX1 INVX1_419 ( .A(_abc_40319_new_n2695_), .Y(_abc_40319_new_n2727_));
INVX1 INVX1_42 ( .A(_abc_40319_new_n725_), .Y(_abc_40319_new_n753_));
INVX1 INVX1_420 ( .A(_abc_40319_new_n2728_), .Y(_abc_40319_new_n2731_));
INVX1 INVX1_421 ( .A(_abc_40319_new_n2732_), .Y(_abc_40319_new_n2733_));
INVX1 INVX1_422 ( .A(_abc_40319_new_n1369_), .Y(_abc_40319_new_n2738_));
INVX1 INVX1_423 ( .A(_abc_40319_new_n2739_), .Y(_abc_40319_new_n2740_));
INVX1 INVX1_424 ( .A(_abc_40319_new_n2741_), .Y(_abc_40319_new_n2742_));
INVX1 INVX1_425 ( .A(_abc_40319_new_n2748_), .Y(_abc_40319_new_n2749_));
INVX1 INVX1_426 ( .A(_abc_40319_new_n2750_), .Y(_abc_40319_new_n2751_));
INVX1 INVX1_427 ( .A(_abc_40319_new_n1348_), .Y(_abc_40319_new_n2761_));
INVX1 INVX1_428 ( .A(_abc_40319_new_n2763_), .Y(_abc_40319_new_n2764_));
INVX1 INVX1_429 ( .A(_abc_40319_new_n2785_), .Y(_abc_40319_new_n2786_));
INVX1 INVX1_43 ( .A(_abc_40319_new_n739_), .Y(_abc_40319_new_n754_));
INVX1 INVX1_430 ( .A(_abc_40319_new_n2771_), .Y(_abc_40319_new_n2792_));
INVX1 INVX1_431 ( .A(_abc_40319_new_n2770_), .Y(_abc_40319_new_n2815_));
INVX1 INVX1_432 ( .A(_abc_40319_new_n2789_), .Y(_abc_40319_new_n2816_));
INVX1 INVX1_433 ( .A(_abc_40319_new_n2834_), .Y(_abc_40319_new_n2835_));
INVX1 INVX1_434 ( .A(_abc_40319_new_n1221_), .Y(_abc_40319_new_n2836_));
INVX1 INVX1_435 ( .A(_abc_40319_new_n2837_), .Y(_abc_40319_new_n2838_));
INVX1 INVX1_436 ( .A(_abc_40319_new_n2790_), .Y(_abc_40319_new_n2840_));
INVX1 INVX1_437 ( .A(_abc_40319_new_n2813_), .Y(_abc_40319_new_n2841_));
INVX1 INVX1_438 ( .A(_abc_40319_new_n2853_), .Y(_abc_40319_new_n2854_));
INVX1 INVX1_439 ( .A(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2855_));
INVX1 INVX1_44 ( .A(_abc_40319_new_n740_), .Y(_abc_40319_new_n759_));
INVX1 INVX1_440 ( .A(_abc_40319_new_n2856_), .Y(_abc_40319_new_n2857_));
INVX1 INVX1_441 ( .A(_abc_40319_new_n1680_), .Y(_abc_40319_new_n2862_));
INVX1 INVX1_442 ( .A(_abc_40319_new_n2864_), .Y(_abc_40319_new_n2865_));
INVX1 INVX1_443 ( .A(_abc_40319_new_n2812_), .Y(_abc_40319_new_n2867_));
INVX1 INVX1_444 ( .A(_abc_40319_new_n1196_), .Y(_abc_40319_new_n2879_));
INVX1 INVX1_445 ( .A(_abc_40319_new_n1146_), .Y(_abc_40319_new_n2899_));
INVX1 INVX1_446 ( .A(_abc_40319_new_n2880_), .Y(_abc_40319_new_n2902_));
INVX1 INVX1_447 ( .A(_abc_40319_new_n2900_), .Y(_abc_40319_new_n2908_));
INVX1 INVX1_448 ( .A(_abc_40319_new_n2901_), .Y(_abc_40319_new_n2909_));
INVX1 INVX1_449 ( .A(_abc_40319_new_n2878_), .Y(_abc_40319_new_n2910_));
INVX1 INVX1_45 ( .A(REG2_REG_5_), .Y(_abc_40319_new_n770_));
INVX1 INVX1_450 ( .A(_abc_40319_new_n2915_), .Y(_abc_40319_new_n2916_));
INVX1 INVX1_451 ( .A(REG2_REG_18_), .Y(_abc_40319_new_n2917_));
INVX1 INVX1_452 ( .A(_abc_40319_new_n2918_), .Y(_abc_40319_new_n2919_));
INVX1 INVX1_453 ( .A(_abc_40319_new_n2932_), .Y(_abc_40319_new_n2935_));
INVX1 INVX1_454 ( .A(REG2_REG_19_), .Y(_abc_40319_new_n2939_));
INVX1 INVX1_455 ( .A(_abc_40319_new_n2960_), .Y(_abc_40319_new_n2990_));
INVX1 INVX1_456 ( .A(_abc_40319_new_n2991_), .Y(_abc_40319_new_n2992_));
INVX1 INVX1_457 ( .A(_abc_40319_new_n2961_), .Y(_abc_40319_new_n2996_));
INVX1 INVX1_458 ( .A(_abc_40319_new_n3006_), .Y(_abc_40319_new_n3007_));
INVX1 INVX1_459 ( .A(_abc_40319_new_n3018_), .Y(_abc_40319_new_n3019_));
INVX1 INVX1_46 ( .A(REG0_REG_5_), .Y(_abc_40319_new_n776_));
INVX1 INVX1_460 ( .A(_abc_40319_new_n2198_), .Y(_abc_40319_new_n3020_));
INVX1 INVX1_461 ( .A(_abc_40319_new_n3022_), .Y(_abc_40319_new_n3023_));
INVX1 INVX1_462 ( .A(_abc_40319_new_n3026_), .Y(_abc_40319_new_n3027_));
INVX1 INVX1_463 ( .A(_abc_40319_new_n2238_), .Y(_abc_40319_new_n3030_));
INVX1 INVX1_464 ( .A(_abc_40319_new_n3031_), .Y(_abc_40319_new_n3032_));
INVX1 INVX1_465 ( .A(_abc_40319_new_n3053_), .Y(_abc_40319_new_n3054_));
INVX1 INVX1_466 ( .A(_abc_40319_new_n3058_), .Y(_abc_40319_new_n3059_));
INVX1 INVX1_467 ( .A(_abc_40319_new_n3062_), .Y(_abc_40319_new_n3063_));
INVX1 INVX1_468 ( .A(_abc_40319_new_n3072_), .Y(_abc_40319_new_n3073_));
INVX1 INVX1_469 ( .A(_abc_40319_new_n3079_), .Y(_abc_40319_new_n3080_));
INVX1 INVX1_47 ( .A(_abc_40319_new_n727_), .Y(_abc_40319_new_n778_));
INVX1 INVX1_470 ( .A(_abc_40319_new_n3093_), .Y(_abc_40319_new_n3094_));
INVX1 INVX1_471 ( .A(_abc_40319_new_n3098_), .Y(_abc_40319_new_n3099_));
INVX1 INVX1_472 ( .A(_abc_40319_new_n3100_), .Y(_abc_40319_new_n3101_));
INVX1 INVX1_473 ( .A(_abc_40319_new_n3103_), .Y(_abc_40319_new_n3104_));
INVX1 INVX1_474 ( .A(_abc_40319_new_n2261_), .Y(_abc_40319_new_n3119_));
INVX1 INVX1_475 ( .A(_abc_40319_new_n3092_), .Y(_abc_40319_new_n3121_));
INVX1 INVX1_476 ( .A(_abc_40319_new_n3110_), .Y(_abc_40319_new_n3133_));
INVX1 INVX1_477 ( .A(_abc_40319_new_n2125_), .Y(_abc_40319_new_n3144_));
INVX1 INVX1_478 ( .A(_abc_40319_new_n3090_), .Y(_abc_40319_new_n3146_));
INVX1 INVX1_479 ( .A(DATAI_24_), .Y(_abc_40319_new_n3147_));
INVX1 INVX1_48 ( .A(REG3_REG_5_), .Y(_abc_40319_new_n779_));
INVX1 INVX1_480 ( .A(_abc_40319_new_n3005_), .Y(_abc_40319_new_n3155_));
INVX1 INVX1_481 ( .A(_abc_40319_new_n3160_), .Y(_abc_40319_new_n3161_));
INVX1 INVX1_482 ( .A(_abc_40319_new_n3108_), .Y(_abc_40319_new_n3164_));
INVX1 INVX1_483 ( .A(_abc_40319_new_n3171_), .Y(_abc_40319_new_n3172_));
INVX1 INVX1_484 ( .A(_abc_40319_new_n2457_), .Y(_abc_40319_new_n3178_));
INVX1 INVX1_485 ( .A(_abc_40319_new_n1072_), .Y(_abc_40319_new_n3192_));
INVX1 INVX1_486 ( .A(_abc_40319_new_n3200_), .Y(_abc_40319_new_n3201_));
INVX1 INVX1_487 ( .A(_abc_40319_new_n2134_), .Y(_abc_40319_new_n3203_));
INVX1 INVX1_488 ( .A(_abc_40319_new_n3220_), .Y(_abc_40319_new_n3221_));
INVX1 INVX1_489 ( .A(_abc_40319_new_n2975_), .Y(_abc_40319_new_n3224_));
INVX1 INVX1_49 ( .A(_abc_40319_new_n791_), .Y(_abc_40319_new_n792_));
INVX1 INVX1_490 ( .A(DATAI_20_), .Y(_abc_40319_new_n3247_));
INVX1 INVX1_491 ( .A(_abc_40319_new_n2974_), .Y(_abc_40319_new_n3248_));
INVX1 INVX1_492 ( .A(_abc_40319_new_n2143_), .Y(_abc_40319_new_n3265_));
INVX1 INVX1_493 ( .A(_abc_40319_new_n3283_), .Y(_abc_40319_new_n3284_));
INVX1 INVX1_494 ( .A(_abc_40319_new_n2498_), .Y(_abc_40319_new_n3290_));
INVX1 INVX1_495 ( .A(_abc_40319_new_n3316_), .Y(_abc_40319_new_n3317_));
INVX1 INVX1_496 ( .A(_abc_40319_new_n3331_), .Y(_abc_40319_new_n3332_));
INVX1 INVX1_497 ( .A(_abc_40319_new_n3340_), .Y(_abc_40319_new_n3341_));
INVX1 INVX1_498 ( .A(_abc_40319_new_n2327_), .Y(_abc_40319_new_n3346_));
INVX1 INVX1_499 ( .A(_abc_40319_new_n3348_), .Y(_abc_40319_new_n3349_));
INVX1 INVX1_5 ( .A(IR_REG_19_), .Y(_abc_40319_new_n537_));
INVX1 INVX1_50 ( .A(_abc_40319_new_n796_), .Y(_abc_40319_new_n797_));
INVX1 INVX1_500 ( .A(_abc_40319_new_n3352_), .Y(_abc_40319_new_n3353_));
INVX1 INVX1_501 ( .A(_abc_40319_new_n2985_), .Y(_abc_40319_new_n3368_));
INVX1 INVX1_502 ( .A(_abc_40319_new_n3382_), .Y(_abc_40319_new_n3386_));
INVX1 INVX1_503 ( .A(_abc_40319_new_n3409_), .Y(_abc_40319_new_n3410_));
INVX1 INVX1_504 ( .A(_abc_40319_new_n3412_), .Y(_abc_40319_new_n3413_));
INVX1 INVX1_505 ( .A(_abc_40319_new_n3414_), .Y(_abc_40319_new_n3415_));
INVX1 INVX1_506 ( .A(_abc_40319_new_n3424_), .Y(_abc_40319_new_n3425_));
INVX1 INVX1_507 ( .A(_abc_40319_new_n3433_), .Y(_abc_40319_new_n3434_));
INVX1 INVX1_508 ( .A(_abc_40319_new_n3448_), .Y(_abc_40319_new_n3449_));
INVX1 INVX1_509 ( .A(_abc_40319_new_n3454_), .Y(_abc_40319_new_n3455_));
INVX1 INVX1_51 ( .A(REG1_REG_4_), .Y(_abc_40319_new_n800_));
INVX1 INVX1_510 ( .A(_abc_40319_new_n2969_), .Y(_abc_40319_new_n3459_));
INVX1 INVX1_511 ( .A(_abc_40319_new_n3466_), .Y(_abc_40319_new_n3467_));
INVX1 INVX1_512 ( .A(_abc_40319_new_n3478_), .Y(_abc_40319_new_n3479_));
INVX1 INVX1_513 ( .A(_abc_40319_new_n3483_), .Y(_abc_40319_new_n3484_));
INVX1 INVX1_514 ( .A(_abc_40319_new_n3490_), .Y(_abc_40319_new_n3491_));
INVX1 INVX1_515 ( .A(_abc_40319_new_n3497_), .Y(_abc_40319_new_n3498_));
INVX1 INVX1_516 ( .A(_abc_40319_new_n3500_), .Y(_abc_40319_new_n3501_));
INVX1 INVX1_517 ( .A(_abc_40319_new_n3531_), .Y(_abc_40319_new_n3532_));
INVX1 INVX1_518 ( .A(_abc_40319_new_n3534_), .Y(_abc_40319_new_n3535_));
INVX1 INVX1_519 ( .A(_abc_40319_new_n3550_), .Y(_abc_40319_new_n3553_));
INVX1 INVX1_52 ( .A(REG2_REG_4_), .Y(_abc_40319_new_n801_));
INVX1 INVX1_520 ( .A(_abc_40319_new_n3047_), .Y(_abc_40319_new_n3564_));
INVX1 INVX1_521 ( .A(_abc_40319_new_n3569_), .Y(_abc_40319_new_n3570_));
INVX1 INVX1_522 ( .A(_abc_40319_new_n3043_), .Y(_abc_40319_new_n3598_));
INVX1 INVX1_523 ( .A(_abc_40319_new_n2468_), .Y(_abc_40319_new_n3613_));
INVX1 INVX1_524 ( .A(_abc_40319_new_n3622_), .Y(_abc_40319_new_n3623_));
INVX1 INVX1_525 ( .A(_abc_40319_new_n2225_), .Y(_abc_40319_new_n3631_));
INVX1 INVX1_526 ( .A(_abc_40319_new_n3653_), .Y(_abc_40319_new_n3654_));
INVX1 INVX1_527 ( .A(_abc_40319_new_n3657_), .Y(_abc_40319_new_n3658_));
INVX1 INVX1_528 ( .A(_abc_40319_new_n3659_), .Y(n493));
INVX1 INVX1_529 ( .A(_abc_40319_new_n3661_), .Y(n488));
INVX1 INVX1_53 ( .A(REG0_REG_4_), .Y(_abc_40319_new_n804_));
INVX1 INVX1_530 ( .A(_abc_40319_new_n3663_), .Y(n483));
INVX1 INVX1_531 ( .A(_abc_40319_new_n3665_), .Y(n478));
INVX1 INVX1_532 ( .A(_abc_40319_new_n3667_), .Y(n473));
INVX1 INVX1_533 ( .A(_abc_40319_new_n3669_), .Y(n468));
INVX1 INVX1_534 ( .A(_abc_40319_new_n3671_), .Y(n463));
INVX1 INVX1_535 ( .A(_abc_40319_new_n3673_), .Y(n458));
INVX1 INVX1_536 ( .A(_abc_40319_new_n3675_), .Y(n453));
INVX1 INVX1_537 ( .A(_abc_40319_new_n3677_), .Y(n448));
INVX1 INVX1_538 ( .A(_abc_40319_new_n3679_), .Y(n443));
INVX1 INVX1_539 ( .A(_abc_40319_new_n3681_), .Y(n438));
INVX1 INVX1_54 ( .A(_abc_40319_new_n810_), .Y(_abc_40319_new_n811_));
INVX1 INVX1_540 ( .A(_abc_40319_new_n3683_), .Y(n433));
INVX1 INVX1_541 ( .A(_abc_40319_new_n3685_), .Y(n428));
INVX1 INVX1_542 ( .A(_abc_40319_new_n3687_), .Y(n423));
INVX1 INVX1_543 ( .A(_abc_40319_new_n3689_), .Y(n418));
INVX1 INVX1_544 ( .A(_abc_40319_new_n3691_), .Y(n413));
INVX1 INVX1_545 ( .A(_abc_40319_new_n3693_), .Y(n408));
INVX1 INVX1_546 ( .A(_abc_40319_new_n3695_), .Y(n403));
INVX1 INVX1_547 ( .A(_abc_40319_new_n3697_), .Y(n398));
INVX1 INVX1_548 ( .A(_abc_40319_new_n3699_), .Y(n393));
INVX1 INVX1_549 ( .A(_abc_40319_new_n3701_), .Y(n388));
INVX1 INVX1_55 ( .A(_abc_40319_new_n821_), .Y(_abc_40319_new_n822_));
INVX1 INVX1_550 ( .A(_abc_40319_new_n3703_), .Y(n383));
INVX1 INVX1_551 ( .A(_abc_40319_new_n3705_), .Y(n378));
INVX1 INVX1_552 ( .A(_abc_40319_new_n3707_), .Y(n373));
INVX1 INVX1_553 ( .A(_abc_40319_new_n3709_), .Y(n368));
INVX1 INVX1_554 ( .A(_abc_40319_new_n3711_), .Y(n363));
INVX1 INVX1_555 ( .A(_abc_40319_new_n3713_), .Y(n358));
INVX1 INVX1_556 ( .A(_abc_40319_new_n3715_), .Y(n353));
INVX1 INVX1_557 ( .A(_abc_40319_new_n3717_), .Y(n348));
INVX1 INVX1_558 ( .A(DATAI_28_), .Y(_abc_40319_new_n3726_));
INVX1 INVX1_559 ( .A(_abc_40319_new_n3735_), .Y(_abc_40319_new_n3736_));
INVX1 INVX1_56 ( .A(DATAI_3_), .Y(_abc_40319_new_n823_));
INVX1 INVX1_560 ( .A(_abc_40319_new_n3739_), .Y(_abc_40319_new_n3740_));
INVX1 INVX1_561 ( .A(_abc_40319_new_n3744_), .Y(_abc_40319_new_n3745_));
INVX1 INVX1_562 ( .A(_abc_40319_new_n3750_), .Y(_abc_40319_new_n3751_));
INVX1 INVX1_563 ( .A(_abc_40319_new_n3757_), .Y(_abc_40319_new_n3758_));
INVX1 INVX1_564 ( .A(_abc_40319_new_n3812_), .Y(_abc_40319_new_n3813_));
INVX1 INVX1_565 ( .A(_abc_40319_new_n3823_), .Y(_abc_40319_new_n3824_));
INVX1 INVX1_566 ( .A(_abc_40319_new_n2118_), .Y(_abc_40319_new_n3827_));
INVX1 INVX1_567 ( .A(_abc_40319_new_n3848_), .Y(_abc_40319_new_n3849_));
INVX1 INVX1_568 ( .A(_abc_40319_new_n2982_), .Y(_abc_40319_new_n3855_));
INVX1 INVX1_569 ( .A(_abc_40319_new_n3877_), .Y(_abc_40319_new_n3878_));
INVX1 INVX1_57 ( .A(_abc_40319_new_n825_), .Y(_abc_40319_new_n826_));
INVX1 INVX1_570 ( .A(D_REG_1_), .Y(_abc_40319_new_n3882_));
INVX1 INVX1_571 ( .A(_abc_40319_new_n3887_), .Y(_abc_40319_new_n3888_));
INVX1 INVX1_572 ( .A(_abc_40319_new_n3889_), .Y(_abc_40319_new_n3890_));
INVX1 INVX1_573 ( .A(_abc_40319_new_n3620_), .Y(_abc_40319_new_n3891_));
INVX1 INVX1_574 ( .A(_abc_40319_new_n1005_), .Y(_abc_40319_new_n3893_));
INVX1 INVX1_575 ( .A(REG0_REG_3_), .Y(_abc_40319_new_n3914_));
INVX1 INVX1_576 ( .A(_abc_40319_new_n3927_), .Y(_abc_40319_new_n3928_));
INVX1 INVX1_577 ( .A(REG0_REG_7_), .Y(_abc_40319_new_n3936_));
INVX1 INVX1_578 ( .A(REG0_REG_8_), .Y(_abc_40319_new_n3943_));
INVX1 INVX1_579 ( .A(_abc_40319_new_n3505_), .Y(_abc_40319_new_n3949_));
INVX1 INVX1_58 ( .A(REG2_REG_3_), .Y(_abc_40319_new_n827_));
INVX1 INVX1_580 ( .A(_abc_40319_new_n3962_), .Y(_abc_40319_new_n3963_));
INVX1 INVX1_581 ( .A(_abc_40319_new_n4003_), .Y(_abc_40319_new_n4004_));
INVX1 INVX1_582 ( .A(_abc_40319_new_n3279_), .Y(_abc_40319_new_n4013_));
INVX1 INVX1_583 ( .A(_abc_40319_new_n4024_), .Y(_abc_40319_new_n4025_));
INVX1 INVX1_584 ( .A(_abc_40319_new_n4030_), .Y(_abc_40319_new_n4031_));
INVX1 INVX1_585 ( .A(_abc_40319_new_n4036_), .Y(_abc_40319_new_n4037_));
INVX1 INVX1_586 ( .A(_abc_40319_new_n4042_), .Y(_abc_40319_new_n4043_));
INVX1 INVX1_587 ( .A(_abc_40319_new_n4048_), .Y(_abc_40319_new_n4049_));
INVX1 INVX1_588 ( .A(_abc_40319_new_n4057_), .Y(_abc_40319_new_n4058_));
INVX1 INVX1_589 ( .A(_abc_40319_new_n4064_), .Y(_abc_40319_new_n4065_));
INVX1 INVX1_59 ( .A(REG1_REG_3_), .Y(_abc_40319_new_n828_));
INVX1 INVX1_590 ( .A(_abc_40319_new_n4084_), .Y(_abc_40319_new_n4085_));
INVX1 INVX1_591 ( .A(REG1_REG_2_), .Y(_abc_40319_new_n4091_));
INVX1 INVX1_592 ( .A(n1345), .Y(_abc_40319_new_n4158_));
INVX1 INVX1_6 ( .A(IR_REG_22_), .Y(_abc_40319_new_n543_));
INVX1 INVX1_60 ( .A(_abc_40319_new_n829_), .Y(_abc_40319_new_n830_));
INVX1 INVX1_61 ( .A(_abc_40319_new_n833_), .Y(_abc_40319_new_n834_));
INVX1 INVX1_62 ( .A(_abc_40319_new_n836_), .Y(_abc_40319_new_n837_));
INVX1 INVX1_63 ( .A(_abc_40319_new_n843_), .Y(_abc_40319_new_n844_));
INVX1 INVX1_64 ( .A(_abc_40319_new_n840_), .Y(_abc_40319_new_n846_));
INVX1 INVX1_65 ( .A(REG2_REG_2_), .Y(_abc_40319_new_n847_));
INVX1 INVX1_66 ( .A(REG0_REG_2_), .Y(_abc_40319_new_n848_));
INVX1 INVX1_67 ( .A(_abc_40319_new_n839_), .Y(_abc_40319_new_n853_));
INVX1 INVX1_68 ( .A(_abc_40319_new_n842_), .Y(_abc_40319_new_n855_));
INVX1 INVX1_69 ( .A(_abc_40319_new_n858_), .Y(_abc_40319_new_n859_));
INVX1 INVX1_7 ( .A(IR_REG_1_), .Y(_abc_40319_new_n544_));
INVX1 INVX1_70 ( .A(_abc_40319_new_n831_), .Y(_abc_40319_new_n861_));
INVX1 INVX1_71 ( .A(IR_REG_0_), .Y(_abc_40319_new_n871_));
INVX1 INVX1_72 ( .A(_abc_40319_new_n835_), .Y(_abc_40319_new_n872_));
INVX1 INVX1_73 ( .A(REG1_REG_1_), .Y(_abc_40319_new_n883_));
INVX1 INVX1_74 ( .A(REG0_REG_1_), .Y(_abc_40319_new_n884_));
INVX1 INVX1_75 ( .A(DATAI_1_), .Y(_abc_40319_new_n893_));
INVX1 INVX1_76 ( .A(_abc_40319_new_n880_), .Y(_abc_40319_new_n897_));
INVX1 INVX1_77 ( .A(_abc_40319_new_n881_), .Y(_abc_40319_new_n902_));
INVX1 INVX1_78 ( .A(REG0_REG_0_), .Y(_abc_40319_new_n906_));
INVX1 INVX1_79 ( .A(REG2_REG_0_), .Y(_abc_40319_new_n907_));
INVX1 INVX1_8 ( .A(IR_REG_5_), .Y(_abc_40319_new_n547_));
INVX1 INVX1_80 ( .A(REG1_REG_0_), .Y(_abc_40319_new_n909_));
INVX1 INVX1_81 ( .A(DATAI_0_), .Y(_abc_40319_new_n920_));
INVX1 INVX1_82 ( .A(REG1_REG_6_), .Y(_abc_40319_new_n945_));
INVX1 INVX1_83 ( .A(_abc_40319_new_n733_), .Y(_abc_40319_new_n946_));
INVX1 INVX1_84 ( .A(_abc_40319_new_n948_), .Y(_abc_40319_new_n949_));
INVX1 INVX1_85 ( .A(REG2_REG_6_), .Y(_abc_40319_new_n951_));
INVX1 INVX1_86 ( .A(REG0_REG_6_), .Y(_abc_40319_new_n952_));
INVX1 INVX1_87 ( .A(_abc_40319_new_n954_), .Y(_abc_40319_new_n959_));
INVX1 INVX1_88 ( .A(_abc_40319_new_n965_), .Y(_abc_40319_new_n966_));
INVX1 INVX1_89 ( .A(_abc_40319_new_n964_), .Y(_abc_40319_new_n968_));
INVX1 INVX1_9 ( .A(IR_REG_4_), .Y(_abc_40319_new_n548_));
INVX1 INVX1_90 ( .A(_abc_40319_new_n674_), .Y(_abc_40319_new_n972_));
INVX1 INVX1_91 ( .A(_abc_40319_new_n668_), .Y(_abc_40319_new_n973_));
INVX1 INVX1_92 ( .A(_abc_40319_new_n974_), .Y(_abc_40319_new_n975_));
INVX1 INVX1_93 ( .A(_abc_40319_new_n696_), .Y(_abc_40319_new_n977_));
INVX1 INVX1_94 ( .A(_abc_40319_new_n978_), .Y(_abc_40319_new_n979_));
INVX1 INVX1_95 ( .A(REG3_REG_8_), .Y(_abc_40319_new_n980_));
INVX1 INVX1_96 ( .A(_abc_40319_new_n982_), .Y(_abc_40319_new_n983_));
INVX1 INVX1_97 ( .A(_abc_40319_new_n987_), .Y(_abc_40319_new_n988_));
INVX1 INVX1_98 ( .A(_abc_40319_new_n976_), .Y(_abc_40319_new_n991_));
INVX1 INVX1_99 ( .A(_abc_40319_new_n663_), .Y(_abc_40319_new_n992_));
MUX2X1 MUX2X1_1 ( .A(_abc_40319_new_n744_), .B(REG1_REG_0_), .S(_abc_40319_new_n574_), .Y(_abc_40319_new_n928_));
MUX2X1 MUX2X1_2 ( .A(_abc_40319_new_n1369_), .B(DATAI_11_), .S(_abc_40319_new_n1341_), .Y(_abc_40319_new_n1370_));
MUX2X1 MUX2X1_3 ( .A(_abc_40319_new_n3455_), .B(_abc_40319_new_n1354_), .S(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3456_));
MUX2X1 MUX2X1_4 ( .A(_abc_40319_new_n3472_), .B(_abc_40319_new_n1373_), .S(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3473_));
NAND2X1 NAND2X1_1 ( .A(_abc_40319_new_n544_), .B(_abc_40319_new_n545_), .Y(_abc_40319_new_n546_));
NAND2X1 NAND2X1_10 ( .A(_abc_40319_new_n588_), .B(_abc_40319_new_n561_), .Y(_abc_40319_new_n589_));
NAND2X1 NAND2X1_100 ( .A(REG0_REG_16_), .B(_abc_40319_new_n724_), .Y(_abc_40319_new_n1177_));
NAND2X1 NAND2X1_101 ( .A(REG3_REG_14_), .B(REG3_REG_15_), .Y(_abc_40319_new_n1181_));
NAND2X1 NAND2X1_102 ( .A(IR_REG_31_), .B(_abc_40319_new_n1194_), .Y(_abc_40319_new_n1195_));
NAND2X1 NAND2X1_103 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n1214_), .Y(_abc_40319_new_n1215_));
NAND2X1 NAND2X1_104 ( .A(_abc_40319_new_n1218_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n1219_));
NAND2X1 NAND2X1_105 ( .A(IR_REG_31_), .B(_abc_40319_new_n1219_), .Y(_abc_40319_new_n1220_));
NAND2X1 NAND2X1_106 ( .A(REG3_REG_14_), .B(_abc_40319_new_n1028_), .Y(_abc_40319_new_n1229_));
NAND2X1 NAND2X1_107 ( .A(_abc_40319_new_n727_), .B(_abc_40319_new_n1230_), .Y(_abc_40319_new_n1231_));
NAND2X1 NAND2X1_108 ( .A(_abc_40319_new_n1234_), .B(_abc_40319_new_n1237_), .Y(_abc_40319_new_n1238_));
NAND2X1 NAND2X1_109 ( .A(IR_REG_14_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n1244_));
NAND2X1 NAND2X1_11 ( .A(IR_REG_28_), .B(_abc_40319_new_n591_), .Y(_abc_40319_new_n601_));
NAND2X1 NAND2X1_110 ( .A(_abc_40319_new_n727_), .B(_abc_40319_new_n1255_), .Y(_abc_40319_new_n1256_));
NAND2X1 NAND2X1_111 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n1264_), .Y(_abc_40319_new_n1266_));
NAND2X1 NAND2X1_112 ( .A(IR_REG_8_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n1272_));
NAND2X1 NAND2X1_113 ( .A(_abc_40319_new_n1277_), .B(_abc_40319_new_n1279_), .Y(_abc_40319_new_n1283_));
NAND2X1 NAND2X1_114 ( .A(_abc_40319_new_n1283_), .B(_abc_40319_new_n1287_), .Y(_abc_40319_new_n1288_));
NAND2X1 NAND2X1_115 ( .A(_abc_40319_new_n1289_), .B(_abc_40319_new_n1267_), .Y(_abc_40319_new_n1290_));
NAND2X1 NAND2X1_116 ( .A(IR_REG_31_), .B(_abc_40319_new_n1292_), .Y(_abc_40319_new_n1293_));
NAND2X1 NAND2X1_117 ( .A(REG3_REG_9_), .B(_abc_40319_new_n982_), .Y(_abc_40319_new_n1299_));
NAND2X1 NAND2X1_118 ( .A(_abc_40319_new_n1302_), .B(_abc_40319_new_n727_), .Y(_abc_40319_new_n1303_));
NAND2X1 NAND2X1_119 ( .A(IR_REG_13_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n1321_));
NAND2X1 NAND2X1_12 ( .A(_abc_40319_new_n605_), .B(_abc_40319_new_n557_), .Y(_abc_40319_new_n606_));
NAND2X1 NAND2X1_120 ( .A(_abc_40319_new_n1337_), .B(_abc_40319_new_n1339_), .Y(_abc_40319_new_n1340_));
NAND2X1 NAND2X1_121 ( .A(IR_REG_12_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n1347_));
NAND2X1 NAND2X1_122 ( .A(_abc_40319_new_n1341_), .B(_abc_40319_new_n1348_), .Y(_abc_40319_new_n1349_));
NAND2X1 NAND2X1_123 ( .A(_abc_40319_new_n727_), .B(_abc_40319_new_n1357_), .Y(_abc_40319_new_n1358_));
NAND2X1 NAND2X1_124 ( .A(_abc_40319_new_n1361_), .B(_abc_40319_new_n1363_), .Y(_abc_40319_new_n1364_));
NAND2X1 NAND2X1_125 ( .A(IR_REG_11_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n1368_));
NAND2X1 NAND2X1_126 ( .A(REG0_REG_11_), .B(_abc_40319_new_n724_), .Y(_abc_40319_new_n1375_));
NAND2X1 NAND2X1_127 ( .A(_abc_40319_new_n1026_), .B(_abc_40319_new_n1376_), .Y(_abc_40319_new_n1377_));
NAND2X1 NAND2X1_128 ( .A(_abc_40319_new_n1387_), .B(_abc_40319_new_n1344_), .Y(_abc_40319_new_n1388_));
NAND2X1 NAND2X1_129 ( .A(IR_REG_10_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n1389_));
NAND2X1 NAND2X1_13 ( .A(IR_REG_22_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n607_));
NAND2X1 NAND2X1_130 ( .A(REG2_REG_10_), .B(_abc_40319_new_n715_), .Y(_abc_40319_new_n1395_));
NAND2X1 NAND2X1_131 ( .A(_abc_40319_new_n1404_), .B(_abc_40319_new_n1406_), .Y(_abc_40319_new_n1408_));
NAND2X1 NAND2X1_132 ( .A(_abc_40319_new_n1382_), .B(_abc_40319_new_n1384_), .Y(_abc_40319_new_n1410_));
NAND2X1 NAND2X1_133 ( .A(_abc_40319_new_n1411_), .B(_abc_40319_new_n1365_), .Y(_abc_40319_new_n1412_));
NAND2X1 NAND2X1_134 ( .A(_abc_40319_new_n1266_), .B(_abc_40319_new_n1419_), .Y(_abc_40319_new_n1420_));
NAND2X1 NAND2X1_135 ( .A(_abc_40319_new_n1191_), .B(_abc_40319_new_n1193_), .Y(_abc_40319_new_n1423_));
NAND2X1 NAND2X1_136 ( .A(_abc_40319_new_n727_), .B(_abc_40319_new_n1432_), .Y(_abc_40319_new_n1433_));
NAND2X1 NAND2X1_137 ( .A(REG2_REG_19_), .B(_abc_40319_new_n715_), .Y(_abc_40319_new_n1434_));
NAND2X1 NAND2X1_138 ( .A(REG0_REG_19_), .B(_abc_40319_new_n724_), .Y(_abc_40319_new_n1435_));
NAND2X1 NAND2X1_139 ( .A(_abc_40319_new_n1445_), .B(_abc_40319_new_n1126_), .Y(_abc_40319_new_n1446_));
NAND2X1 NAND2X1_14 ( .A(_abc_40319_new_n554_), .B(_abc_40319_new_n553_), .Y(_abc_40319_new_n611_));
NAND2X1 NAND2X1_140 ( .A(REG2_REG_20_), .B(_abc_40319_new_n715_), .Y(_abc_40319_new_n1448_));
NAND2X1 NAND2X1_141 ( .A(REG0_REG_20_), .B(_abc_40319_new_n724_), .Y(_abc_40319_new_n1449_));
NAND2X1 NAND2X1_142 ( .A(REG1_REG_20_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n1450_));
NAND2X1 NAND2X1_143 ( .A(REG3_REG_21_), .B(_abc_40319_new_n1034_), .Y(_abc_40319_new_n1461_));
NAND2X1 NAND2X1_144 ( .A(_abc_40319_new_n1124_), .B(_abc_40319_new_n1126_), .Y(_abc_40319_new_n1462_));
NAND2X1 NAND2X1_145 ( .A(_abc_40319_new_n1462_), .B(_abc_40319_new_n1461_), .Y(_abc_40319_new_n1463_));
NAND2X1 NAND2X1_146 ( .A(REG0_REG_21_), .B(_abc_40319_new_n724_), .Y(_abc_40319_new_n1465_));
NAND2X1 NAND2X1_147 ( .A(REG1_REG_21_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n1466_));
NAND2X1 NAND2X1_148 ( .A(REG2_REG_21_), .B(_abc_40319_new_n715_), .Y(_abc_40319_new_n1467_));
NAND2X1 NAND2X1_149 ( .A(_abc_40319_new_n1439_), .B(_abc_40319_new_n1441_), .Y(_abc_40319_new_n1480_));
NAND2X1 NAND2X1_15 ( .A(B_REG), .B(_abc_40319_new_n623_), .Y(_abc_40319_new_n624_));
NAND2X1 NAND2X1_150 ( .A(_abc_40319_new_n1454_), .B(_abc_40319_new_n1456_), .Y(_abc_40319_new_n1482_));
NAND2X1 NAND2X1_151 ( .A(_abc_40319_new_n1095_), .B(_abc_40319_new_n1099_), .Y(_abc_40319_new_n1489_));
NAND2X1 NAND2X1_152 ( .A(REG1_REG_28_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n1501_));
NAND2X1 NAND2X1_153 ( .A(_abc_40319_new_n1266_), .B(_abc_40319_new_n1265_), .Y(_abc_40319_new_n1512_));
NAND2X1 NAND2X1_154 ( .A(_abc_40319_new_n1141_), .B(_abc_40319_new_n1487_), .Y(_abc_40319_new_n1525_));
NAND2X1 NAND2X1_155 ( .A(_abc_40319_new_n1121_), .B(_abc_40319_new_n1120_), .Y(_abc_40319_new_n1526_));
NAND2X1 NAND2X1_156 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1529_), .Y(_abc_40319_new_n1530_));
NAND2X1 NAND2X1_157 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1539_), .Y(_abc_40319_new_n1540_));
NAND2X1 NAND2X1_158 ( .A(_abc_40319_new_n917_), .B(_abc_40319_new_n930_), .Y(_abc_40319_new_n1549_));
NAND2X1 NAND2X1_159 ( .A(REG1_REG_29_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n1593_));
NAND2X1 NAND2X1_16 ( .A(_abc_40319_new_n567_), .B(_abc_40319_new_n572_), .Y(_abc_40319_new_n629_));
NAND2X1 NAND2X1_160 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1599_), .Y(_abc_40319_new_n1600_));
NAND2X1 NAND2X1_161 ( .A(_abc_40319_new_n1497_), .B(_abc_40319_new_n1498_), .Y(_abc_40319_new_n1601_));
NAND2X1 NAND2X1_162 ( .A(_abc_40319_new_n1283_), .B(_abc_40319_new_n1284_), .Y(_abc_40319_new_n1607_));
NAND2X1 NAND2X1_163 ( .A(_abc_40319_new_n1613_), .B(_abc_40319_new_n1619_), .Y(n1291));
NAND2X1 NAND2X1_164 ( .A(_abc_40319_new_n903_), .B(_abc_40319_new_n901_), .Y(_abc_40319_new_n1621_));
NAND2X1 NAND2X1_165 ( .A(_abc_40319_new_n1480_), .B(_abc_40319_new_n1633_), .Y(_abc_40319_new_n1634_));
NAND2X1 NAND2X1_166 ( .A(_abc_40319_new_n1364_), .B(_abc_40319_new_n1414_), .Y(_abc_40319_new_n1645_));
NAND2X1 NAND2X1_167 ( .A(_abc_40319_new_n676_), .B(_abc_40319_new_n1665_), .Y(_abc_40319_new_n1666_));
NAND2X1 NAND2X1_168 ( .A(_abc_40319_new_n1238_), .B(_abc_40319_new_n1421_), .Y(_abc_40319_new_n1673_));
NAND2X1 NAND2X1_169 ( .A(_abc_40319_new_n793_), .B(_abc_40319_new_n792_), .Y(_abc_40319_new_n1685_));
NAND2X1 NAND2X1_17 ( .A(_abc_40319_new_n654_), .B(_abc_40319_new_n656_), .Y(_abc_40319_new_n657_));
NAND2X1 NAND2X1_170 ( .A(_abc_40319_new_n1687_), .B(_abc_40319_new_n1692_), .Y(n1261));
NAND2X1 NAND2X1_171 ( .A(_abc_40319_new_n1489_), .B(_abc_40319_new_n1101_), .Y(_abc_40319_new_n1707_));
NAND2X1 NAND2X1_172 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1711_), .Y(_abc_40319_new_n1712_));
NAND2X1 NAND2X1_173 ( .A(_abc_40319_new_n1087_), .B(_abc_40319_new_n1058_), .Y(_abc_40319_new_n1713_));
NAND2X1 NAND2X1_174 ( .A(_abc_40319_new_n817_), .B(_abc_40319_new_n816_), .Y(_abc_40319_new_n1720_));
NAND2X1 NAND2X1_175 ( .A(_abc_40319_new_n925_), .B(_abc_40319_new_n929_), .Y(_abc_40319_new_n1746_));
NAND2X1 NAND2X1_176 ( .A(_abc_40319_new_n919_), .B(_abc_40319_new_n917_), .Y(_abc_40319_new_n1747_));
NAND2X1 NAND2X1_177 ( .A(_abc_40319_new_n1482_), .B(_abc_40319_new_n1458_), .Y(_abc_40319_new_n1757_));
NAND2X1 NAND2X1_178 ( .A(_abc_40319_new_n1364_), .B(_abc_40319_new_n1767_), .Y(_abc_40319_new_n1769_));
NAND2X1 NAND2X1_179 ( .A(_abc_40319_new_n1770_), .B(_abc_40319_new_n1769_), .Y(_abc_40319_new_n1771_));
NAND2X1 NAND2X1_18 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n614_), .Y(_abc_40319_new_n660_));
NAND2X1 NAND2X1_180 ( .A(_abc_40319_new_n1486_), .B(_abc_40319_new_n1479_), .Y(_abc_40319_new_n1781_));
NAND2X1 NAND2X1_181 ( .A(_abc_40319_new_n1141_), .B(_abc_40319_new_n1143_), .Y(_abc_40319_new_n1782_));
NAND2X1 NAND2X1_182 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1786_), .Y(_abc_40319_new_n1787_));
NAND2X1 NAND2X1_183 ( .A(_abc_40319_new_n1410_), .B(_abc_40319_new_n1646_), .Y(_abc_40319_new_n1793_));
NAND2X1 NAND2X1_184 ( .A(_abc_40319_new_n1163_), .B(_abc_40319_new_n1165_), .Y(_abc_40319_new_n1819_));
NAND2X1 NAND2X1_185 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1822_), .Y(_abc_40319_new_n1823_));
NAND2X1 NAND2X1_186 ( .A(_abc_40319_new_n1847_), .B(_abc_40319_new_n1845_), .Y(_abc_40319_new_n1848_));
NAND2X1 NAND2X1_187 ( .A(_abc_40319_new_n1844_), .B(_abc_40319_new_n1848_), .Y(_abc_40319_new_n1849_));
NAND2X1 NAND2X1_188 ( .A(_abc_40319_new_n976_), .B(_abc_40319_new_n1850_), .Y(_abc_40319_new_n1851_));
NAND2X1 NAND2X1_189 ( .A(_abc_40319_new_n1238_), .B(_abc_40319_new_n1240_), .Y(_abc_40319_new_n1859_));
NAND2X1 NAND2X1_19 ( .A(IR_REG_20_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n662_));
NAND2X1 NAND2X1_190 ( .A(REG1_REG_31_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n1880_));
NAND2X1 NAND2X1_191 ( .A(_abc_40319_new_n1886_), .B(_abc_40319_new_n1885_), .Y(_abc_40319_new_n1887_));
NAND2X1 NAND2X1_192 ( .A(_abc_40319_new_n836_), .B(_abc_40319_new_n1341_), .Y(_abc_40319_new_n1889_));
NAND2X1 NAND2X1_193 ( .A(_abc_40319_new_n1902_), .B(_abc_40319_new_n1905_), .Y(_abc_40319_new_n1906_));
NAND2X1 NAND2X1_194 ( .A(_abc_40319_new_n1934_), .B(_abc_40319_new_n1930_), .Y(_abc_40319_new_n1956_));
NAND2X1 NAND2X1_195 ( .A(_abc_40319_new_n1971_), .B(_abc_40319_new_n1953_), .Y(_abc_40319_new_n1972_));
NAND2X1 NAND2X1_196 ( .A(_abc_40319_new_n1951_), .B(_abc_40319_new_n1973_), .Y(_abc_40319_new_n1974_));
NAND2X1 NAND2X1_197 ( .A(_abc_40319_new_n1984_), .B(_abc_40319_new_n1979_), .Y(_abc_40319_new_n1994_));
NAND2X1 NAND2X1_198 ( .A(_abc_40319_new_n1983_), .B(_abc_40319_new_n1978_), .Y(_abc_40319_new_n1997_));
NAND2X1 NAND2X1_199 ( .A(_abc_40319_new_n2013_), .B(_abc_40319_new_n2012_), .Y(_abc_40319_new_n2014_));
NAND2X1 NAND2X1_2 ( .A(_abc_40319_new_n538_), .B(_abc_40319_new_n554_), .Y(_abc_40319_new_n555_));
NAND2X1 NAND2X1_20 ( .A(_abc_40319_new_n611_), .B(_abc_40319_new_n664_), .Y(_abc_40319_new_n665_));
NAND2X1 NAND2X1_200 ( .A(_abc_40319_new_n2018_), .B(_abc_40319_new_n2019_), .Y(_abc_40319_new_n2022_));
NAND2X1 NAND2X1_201 ( .A(_abc_40319_new_n2041_), .B(_abc_40319_new_n2042_), .Y(_abc_40319_new_n2045_));
NAND2X1 NAND2X1_202 ( .A(_abc_40319_new_n2057_), .B(_abc_40319_new_n2059_), .Y(_abc_40319_new_n2060_));
NAND2X1 NAND2X1_203 ( .A(_abc_40319_new_n2086_), .B(_abc_40319_new_n2079_), .Y(_abc_40319_new_n2087_));
NAND2X1 NAND2X1_204 ( .A(REG1_REG_30_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n2100_));
NAND2X1 NAND2X1_205 ( .A(_abc_40319_new_n1582_), .B(_abc_40319_new_n1505_), .Y(_abc_40319_new_n2119_));
NAND2X1 NAND2X1_206 ( .A(_abc_40319_new_n2118_), .B(_abc_40319_new_n2119_), .Y(_abc_40319_new_n2120_));
NAND2X1 NAND2X1_207 ( .A(_abc_40319_new_n1055_), .B(_abc_40319_new_n1496_), .Y(_abc_40319_new_n2124_));
NAND2X1 NAND2X1_208 ( .A(_abc_40319_new_n2123_), .B(_abc_40319_new_n2124_), .Y(_abc_40319_new_n2125_));
NAND2X1 NAND2X1_209 ( .A(_abc_40319_new_n1080_), .B(_abc_40319_new_n1078_), .Y(_abc_40319_new_n2128_));
NAND2X1 NAND2X1_21 ( .A(IR_REG_19_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n666_));
NAND2X1 NAND2X1_210 ( .A(_abc_40319_new_n2127_), .B(_abc_40319_new_n2128_), .Y(_abc_40319_new_n2129_));
NAND2X1 NAND2X1_211 ( .A(_abc_40319_new_n1085_), .B(_abc_40319_new_n1093_), .Y(_abc_40319_new_n2131_));
NAND2X1 NAND2X1_212 ( .A(_abc_40319_new_n1109_), .B(_abc_40319_new_n1710_), .Y(_abc_40319_new_n2135_));
NAND2X1 NAND2X1_213 ( .A(_abc_40319_new_n2137_), .B(_abc_40319_new_n2135_), .Y(_abc_40319_new_n2138_));
NAND2X1 NAND2X1_214 ( .A(_abc_40319_new_n2154_), .B(_abc_40319_new_n2153_), .Y(_abc_40319_new_n2155_));
NAND2X1 NAND2X1_215 ( .A(_abc_40319_new_n1198_), .B(_abc_40319_new_n1208_), .Y(_abc_40319_new_n2157_));
NAND2X1 NAND2X1_216 ( .A(_abc_40319_new_n2156_), .B(_abc_40319_new_n2157_), .Y(_abc_40319_new_n2158_));
NAND2X1 NAND2X1_217 ( .A(_abc_40319_new_n2161_), .B(_abc_40319_new_n2163_), .Y(_abc_40319_new_n2164_));
NAND2X1 NAND2X1_218 ( .A(_abc_40319_new_n2166_), .B(_abc_40319_new_n2168_), .Y(_abc_40319_new_n2169_));
NAND2X1 NAND2X1_219 ( .A(_abc_40319_new_n2165_), .B(_abc_40319_new_n2170_), .Y(_abc_40319_new_n2171_));
NAND2X1 NAND2X1_22 ( .A(_abc_40319_new_n670_), .B(_abc_40319_new_n674_), .Y(_abc_40319_new_n675_));
NAND2X1 NAND2X1_220 ( .A(_abc_40319_new_n799_), .B(_abc_40319_new_n1556_), .Y(_abc_40319_new_n2175_));
NAND2X1 NAND2X1_221 ( .A(_abc_40319_new_n2175_), .B(_abc_40319_new_n2174_), .Y(_abc_40319_new_n2176_));
NAND2X1 NAND2X1_222 ( .A(_abc_40319_new_n2177_), .B(_abc_40319_new_n2179_), .Y(_abc_40319_new_n2180_));
NAND2X1 NAND2X1_223 ( .A(_abc_40319_new_n2189_), .B(_abc_40319_new_n2188_), .Y(_abc_40319_new_n2190_));
NAND2X1 NAND2X1_224 ( .A(_abc_40319_new_n2196_), .B(_abc_40319_new_n1700_), .Y(_abc_40319_new_n2197_));
NAND2X1 NAND2X1_225 ( .A(_abc_40319_new_n2201_), .B(_abc_40319_new_n2203_), .Y(_abc_40319_new_n2204_));
NAND2X1 NAND2X1_226 ( .A(_abc_40319_new_n1401_), .B(_abc_40319_new_n1541_), .Y(_abc_40319_new_n2205_));
NAND2X1 NAND2X1_227 ( .A(_abc_40319_new_n2209_), .B(_abc_40319_new_n2200_), .Y(_abc_40319_new_n2210_));
NAND2X1 NAND2X1_228 ( .A(_abc_40319_new_n2215_), .B(_abc_40319_new_n2214_), .Y(_abc_40319_new_n2216_));
NAND2X1 NAND2X1_229 ( .A(_abc_40319_new_n2221_), .B(_abc_40319_new_n2223_), .Y(_abc_40319_new_n2224_));
NAND2X1 NAND2X1_23 ( .A(_abc_40319_new_n667_), .B(_abc_40319_new_n614_), .Y(_abc_40319_new_n682_));
NAND2X1 NAND2X1_230 ( .A(_abc_40319_new_n1902_), .B(_abc_40319_new_n1898_), .Y(_abc_40319_new_n2225_));
NAND2X1 NAND2X1_231 ( .A(_abc_40319_new_n769_), .B(_abc_40319_new_n788_), .Y(_abc_40319_new_n2233_));
NAND2X1 NAND2X1_232 ( .A(_abc_40319_new_n1905_), .B(_abc_40319_new_n1899_), .Y(_abc_40319_new_n2237_));
NAND2X1 NAND2X1_233 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n855_), .Y(_abc_40319_new_n2244_));
NAND2X1 NAND2X1_234 ( .A(_abc_40319_new_n2243_), .B(_abc_40319_new_n2244_), .Y(_abc_40319_new_n2245_));
NAND2X1 NAND2X1_235 ( .A(_abc_40319_new_n944_), .B(_abc_40319_new_n959_), .Y(_abc_40319_new_n2248_));
NAND2X1 NAND2X1_236 ( .A(_abc_40319_new_n2247_), .B(_abc_40319_new_n2248_), .Y(_abc_40319_new_n2249_));
NAND2X1 NAND2X1_237 ( .A(_abc_40319_new_n2250_), .B(_abc_40319_new_n2242_), .Y(_abc_40319_new_n2251_));
NAND2X1 NAND2X1_238 ( .A(_abc_40319_new_n1018_), .B(_abc_40319_new_n1592_), .Y(_abc_40319_new_n2260_));
NAND2X1 NAND2X1_239 ( .A(_abc_40319_new_n2259_), .B(_abc_40319_new_n2260_), .Y(_abc_40319_new_n2261_));
NAND2X1 NAND2X1_24 ( .A(IR_REG_31_), .B(_abc_40319_new_n688_), .Y(_abc_40319_new_n689_));
NAND2X1 NAND2X1_240 ( .A(_abc_40319_new_n1593_), .B(_abc_40319_new_n1597_), .Y(_abc_40319_new_n2264_));
NAND2X1 NAND2X1_241 ( .A(IR_REG_23_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n2274_));
NAND2X1 NAND2X1_242 ( .A(_abc_40319_new_n1898_), .B(_abc_40319_new_n1899_), .Y(_abc_40319_new_n2275_));
NAND2X1 NAND2X1_243 ( .A(_abc_40319_new_n2275_), .B(_abc_40319_new_n2276_), .Y(_abc_40319_new_n2277_));
NAND2X1 NAND2X1_244 ( .A(_abc_40319_new_n1928_), .B(_abc_40319_new_n1927_), .Y(_abc_40319_new_n2285_));
NAND2X1 NAND2X1_245 ( .A(_abc_40319_new_n1963_), .B(_abc_40319_new_n1962_), .Y(_abc_40319_new_n2286_));
NAND2X1 NAND2X1_246 ( .A(_abc_40319_new_n2285_), .B(_abc_40319_new_n2286_), .Y(_abc_40319_new_n2287_));
NAND2X1 NAND2X1_247 ( .A(_abc_40319_new_n2320_), .B(_abc_40319_new_n2325_), .Y(_abc_40319_new_n2326_));
NAND2X1 NAND2X1_248 ( .A(_abc_40319_new_n2333_), .B(_abc_40319_new_n2329_), .Y(_abc_40319_new_n2334_));
NAND2X1 NAND2X1_249 ( .A(_abc_40319_new_n2342_), .B(_abc_40319_new_n2335_), .Y(_abc_40319_new_n2343_));
NAND2X1 NAND2X1_25 ( .A(IR_REG_27_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n693_));
NAND2X1 NAND2X1_250 ( .A(_abc_40319_new_n2318_), .B(_abc_40319_new_n2344_), .Y(_abc_40319_new_n2345_));
NAND2X1 NAND2X1_251 ( .A(_abc_40319_new_n2350_), .B(_abc_40319_new_n2348_), .Y(_abc_40319_new_n2351_));
NAND2X1 NAND2X1_252 ( .A(_abc_40319_new_n2362_), .B(_abc_40319_new_n1905_), .Y(_abc_40319_new_n2363_));
NAND2X1 NAND2X1_253 ( .A(_abc_40319_new_n2373_), .B(_abc_40319_new_n2375_), .Y(_abc_40319_new_n2376_));
NAND2X1 NAND2X1_254 ( .A(_abc_40319_new_n2408_), .B(_abc_40319_new_n2407_), .Y(_abc_40319_new_n2409_));
NAND2X1 NAND2X1_255 ( .A(_abc_40319_new_n2307_), .B(_abc_40319_new_n2309_), .Y(_abc_40319_new_n2421_));
NAND2X1 NAND2X1_256 ( .A(_abc_40319_new_n2371_), .B(_abc_40319_new_n2370_), .Y(_abc_40319_new_n2425_));
NAND2X1 NAND2X1_257 ( .A(_abc_40319_new_n2234_), .B(_abc_40319_new_n2350_), .Y(_abc_40319_new_n2433_));
NAND2X1 NAND2X1_258 ( .A(_abc_40319_new_n2311_), .B(_abc_40319_new_n2401_), .Y(_abc_40319_new_n2443_));
NAND2X1 NAND2X1_259 ( .A(_abc_40319_new_n667_), .B(_abc_40319_new_n742_), .Y(_abc_40319_new_n2445_));
NAND2X1 NAND2X1_26 ( .A(_abc_40319_new_n693_), .B(_abc_40319_new_n692_), .Y(_abc_40319_new_n694_));
NAND2X1 NAND2X1_260 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n2450_), .Y(_abc_40319_new_n2451_));
NAND2X1 NAND2X1_261 ( .A(_abc_40319_new_n1877_), .B(_abc_40319_new_n2150_), .Y(_abc_40319_new_n2452_));
NAND2X1 NAND2X1_262 ( .A(_abc_40319_new_n2458_), .B(_abc_40319_new_n2406_), .Y(_abc_40319_new_n2459_));
NAND2X1 NAND2X1_263 ( .A(_abc_40319_new_n2332_), .B(_abc_40319_new_n2485_), .Y(_abc_40319_new_n2492_));
NAND2X1 NAND2X1_264 ( .A(_abc_40319_new_n2526_), .B(_abc_40319_new_n2527_), .Y(_abc_40319_new_n2528_));
NAND2X1 NAND2X1_265 ( .A(REG2_REG_1_), .B(_abc_40319_new_n2544_), .Y(_abc_40319_new_n2546_));
NAND2X1 NAND2X1_266 ( .A(REG1_REG_1_), .B(_abc_40319_new_n2532_), .Y(_abc_40319_new_n2550_));
NAND2X1 NAND2X1_267 ( .A(_abc_40319_new_n2551_), .B(_abc_40319_new_n2550_), .Y(_abc_40319_new_n2552_));
NAND2X1 NAND2X1_268 ( .A(_abc_40319_new_n2557_), .B(_abc_40319_new_n2556_), .Y(n1050));
NAND2X1 NAND2X1_269 ( .A(REG1_REG_2_), .B(_abc_40319_new_n836_), .Y(_abc_40319_new_n2569_));
NAND2X1 NAND2X1_27 ( .A(_abc_40319_new_n600_), .B(_abc_40319_new_n601_), .Y(_abc_40319_new_n695_));
NAND2X1 NAND2X1_270 ( .A(_abc_40319_new_n2569_), .B(_abc_40319_new_n2568_), .Y(_abc_40319_new_n2570_));
NAND2X1 NAND2X1_271 ( .A(REG1_REG_3_), .B(_abc_40319_new_n2581_), .Y(_abc_40319_new_n2584_));
NAND2X1 NAND2X1_272 ( .A(_abc_40319_new_n2584_), .B(_abc_40319_new_n2583_), .Y(_abc_40319_new_n2586_));
NAND2X1 NAND2X1_273 ( .A(REG2_REG_4_), .B(_abc_40319_new_n796_), .Y(_abc_40319_new_n2593_));
NAND2X1 NAND2X1_274 ( .A(_abc_40319_new_n801_), .B(_abc_40319_new_n797_), .Y(_abc_40319_new_n2594_));
NAND2X1 NAND2X1_275 ( .A(_abc_40319_new_n2593_), .B(_abc_40319_new_n2594_), .Y(_abc_40319_new_n2595_));
NAND2X1 NAND2X1_276 ( .A(REG1_REG_5_), .B(_abc_40319_new_n2612_), .Y(_abc_40319_new_n2613_));
NAND2X1 NAND2X1_277 ( .A(_abc_40319_new_n2613_), .B(_abc_40319_new_n2615_), .Y(_abc_40319_new_n2616_));
NAND2X1 NAND2X1_278 ( .A(_abc_40319_new_n770_), .B(_abc_40319_new_n767_), .Y(_abc_40319_new_n2628_));
NAND2X1 NAND2X1_279 ( .A(_abc_40319_new_n2637_), .B(_abc_40319_new_n2636_), .Y(n1030));
NAND2X1 NAND2X1_28 ( .A(IR_REG_30_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n708_));
NAND2X1 NAND2X1_280 ( .A(_abc_40319_new_n2639_), .B(_abc_40319_new_n691_), .Y(_abc_40319_new_n2645_));
NAND2X1 NAND2X1_281 ( .A(REG1_REG_7_), .B(_abc_40319_new_n690_), .Y(_abc_40319_new_n2652_));
NAND2X1 NAND2X1_282 ( .A(_abc_40319_new_n2653_), .B(_abc_40319_new_n691_), .Y(_abc_40319_new_n2654_));
NAND2X1 NAND2X1_283 ( .A(_abc_40319_new_n2652_), .B(_abc_40319_new_n2654_), .Y(_abc_40319_new_n2655_));
NAND2X1 NAND2X1_284 ( .A(_abc_40319_new_n2661_), .B(_abc_40319_new_n2660_), .Y(n1026));
NAND2X1 NAND2X1_285 ( .A(REG1_REG_6_), .B(_abc_40319_new_n2642_), .Y(_abc_40319_new_n2673_));
NAND2X1 NAND2X1_286 ( .A(_abc_40319_new_n2672_), .B(_abc_40319_new_n2675_), .Y(_abc_40319_new_n2676_));
NAND2X1 NAND2X1_287 ( .A(_abc_40319_new_n2677_), .B(_abc_40319_new_n2676_), .Y(_abc_40319_new_n2678_));
NAND2X1 NAND2X1_288 ( .A(ADDR_REG_8_), .B(_abc_40319_new_n2539_), .Y(_abc_40319_new_n2690_));
NAND2X1 NAND2X1_289 ( .A(REG2_REG_9_), .B(_abc_40319_new_n1294_), .Y(_abc_40319_new_n2694_));
NAND2X1 NAND2X1_29 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n699_), .Y(_abc_40319_new_n716_));
NAND2X1 NAND2X1_290 ( .A(_abc_40319_new_n1305_), .B(_abc_40319_new_n1295_), .Y(_abc_40319_new_n2695_));
NAND2X1 NAND2X1_291 ( .A(_abc_40319_new_n2694_), .B(_abc_40319_new_n2695_), .Y(_abc_40319_new_n2696_));
NAND2X1 NAND2X1_292 ( .A(_abc_40319_new_n1298_), .B(_abc_40319_new_n1295_), .Y(_abc_40319_new_n2702_));
NAND2X1 NAND2X1_293 ( .A(_abc_40319_new_n2702_), .B(_abc_40319_new_n2701_), .Y(_abc_40319_new_n2703_));
NAND2X1 NAND2X1_294 ( .A(_abc_40319_new_n1274_), .B(_abc_40319_new_n2677_), .Y(_abc_40319_new_n2704_));
NAND2X1 NAND2X1_295 ( .A(_abc_40319_new_n2676_), .B(_abc_40319_new_n2704_), .Y(_abc_40319_new_n2705_));
NAND2X1 NAND2X1_296 ( .A(ADDR_REG_9_), .B(_abc_40319_new_n2539_), .Y(_abc_40319_new_n2708_));
NAND2X1 NAND2X1_297 ( .A(REG1_REG_10_), .B(_abc_40319_new_n2716_), .Y(_abc_40319_new_n2717_));
NAND2X1 NAND2X1_298 ( .A(_abc_40319_new_n2718_), .B(_abc_40319_new_n2717_), .Y(_abc_40319_new_n2719_));
NAND2X1 NAND2X1_299 ( .A(REG2_REG_10_), .B(_abc_40319_new_n1390_), .Y(_abc_40319_new_n2724_));
NAND2X1 NAND2X1_3 ( .A(_abc_40319_new_n541_), .B(_abc_40319_new_n532_), .Y(_abc_40319_new_n563_));
NAND2X1 NAND2X1_30 ( .A(IR_REG_29_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n722_));
NAND2X1 NAND2X1_300 ( .A(_abc_40319_new_n2724_), .B(_abc_40319_new_n2726_), .Y(_abc_40319_new_n2730_));
NAND2X1 NAND2X1_301 ( .A(_abc_40319_new_n2742_), .B(_abc_40319_new_n2740_), .Y(_abc_40319_new_n2743_));
NAND2X1 NAND2X1_302 ( .A(_abc_40319_new_n1391_), .B(_abc_40319_new_n2717_), .Y(_abc_40319_new_n2744_));
NAND2X1 NAND2X1_303 ( .A(_abc_40319_new_n2751_), .B(_abc_40319_new_n2749_), .Y(_abc_40319_new_n2752_));
NAND2X1 NAND2X1_304 ( .A(ADDR_REG_11_), .B(_abc_40319_new_n2539_), .Y(_abc_40319_new_n2755_));
NAND2X1 NAND2X1_305 ( .A(REG1_REG_12_), .B(_abc_40319_new_n2761_), .Y(_abc_40319_new_n2762_));
NAND2X1 NAND2X1_306 ( .A(_abc_40319_new_n2762_), .B(_abc_40319_new_n2764_), .Y(_abc_40319_new_n2765_));
NAND2X1 NAND2X1_307 ( .A(ADDR_REG_12_), .B(_abc_40319_new_n2539_), .Y(_abc_40319_new_n2777_));
NAND2X1 NAND2X1_308 ( .A(_abc_40319_new_n2784_), .B(_abc_40319_new_n2786_), .Y(_abc_40319_new_n2787_));
NAND2X1 NAND2X1_309 ( .A(_abc_40319_new_n1252_), .B(_abc_40319_new_n2803_), .Y(_abc_40319_new_n2804_));
NAND2X1 NAND2X1_31 ( .A(_abc_40319_new_n722_), .B(_abc_40319_new_n721_), .Y(_abc_40319_new_n723_));
NAND2X1 NAND2X1_310 ( .A(_abc_40319_new_n2688_), .B(_abc_40319_new_n2819_), .Y(_abc_40319_new_n2820_));
NAND2X1 NAND2X1_311 ( .A(_abc_40319_new_n2822_), .B(_abc_40319_new_n2820_), .Y(_abc_40319_new_n2823_));
NAND2X1 NAND2X1_312 ( .A(_abc_40319_new_n2524_), .B(_abc_40319_new_n2819_), .Y(_abc_40319_new_n2824_));
NAND2X1 NAND2X1_313 ( .A(_abc_40319_new_n2804_), .B(_abc_40319_new_n2809_), .Y(_abc_40319_new_n2828_));
NAND2X1 NAND2X1_314 ( .A(_abc_40319_new_n1224_), .B(_abc_40319_new_n2828_), .Y(_abc_40319_new_n2829_));
NAND2X1 NAND2X1_315 ( .A(REG1_REG_15_), .B(_abc_40319_new_n2830_), .Y(_abc_40319_new_n2831_));
NAND2X1 NAND2X1_316 ( .A(_abc_40319_new_n2829_), .B(_abc_40319_new_n2831_), .Y(_abc_40319_new_n2832_));
NAND2X1 NAND2X1_317 ( .A(_abc_40319_new_n2835_), .B(_abc_40319_new_n2838_), .Y(_abc_40319_new_n2839_));
NAND2X1 NAND2X1_318 ( .A(_abc_40319_new_n2524_), .B(_abc_40319_new_n2844_), .Y(_abc_40319_new_n2845_));
NAND2X1 NAND2X1_319 ( .A(_abc_40319_new_n2688_), .B(_abc_40319_new_n2844_), .Y(_abc_40319_new_n2847_));
NAND2X1 NAND2X1_32 ( .A(REG3_REG_5_), .B(_abc_40319_new_n731_), .Y(_abc_40319_new_n732_));
NAND2X1 NAND2X1_320 ( .A(_abc_40319_new_n2849_), .B(_abc_40319_new_n2847_), .Y(_abc_40319_new_n2850_));
NAND2X1 NAND2X1_321 ( .A(_abc_40319_new_n2854_), .B(_abc_40319_new_n2857_), .Y(_abc_40319_new_n2858_));
NAND2X1 NAND2X1_322 ( .A(REG2_REG_16_), .B(_abc_40319_new_n2855_), .Y(_abc_40319_new_n2863_));
NAND2X1 NAND2X1_323 ( .A(_abc_40319_new_n2863_), .B(_abc_40319_new_n2865_), .Y(_abc_40319_new_n2866_));
NAND2X1 NAND2X1_324 ( .A(_abc_40319_new_n2688_), .B(_abc_40319_new_n2870_), .Y(_abc_40319_new_n2871_));
NAND2X1 NAND2X1_325 ( .A(_abc_40319_new_n2524_), .B(_abc_40319_new_n2870_), .Y(_abc_40319_new_n2874_));
NAND2X1 NAND2X1_326 ( .A(REG2_REG_17_), .B(_abc_40319_new_n2879_), .Y(_abc_40319_new_n2885_));
NAND2X1 NAND2X1_327 ( .A(_abc_40319_new_n1202_), .B(_abc_40319_new_n1196_), .Y(_abc_40319_new_n2886_));
NAND2X1 NAND2X1_328 ( .A(_abc_40319_new_n2886_), .B(_abc_40319_new_n2885_), .Y(_abc_40319_new_n2887_));
NAND2X1 NAND2X1_329 ( .A(_abc_40319_new_n2524_), .B(_abc_40319_new_n2890_), .Y(_abc_40319_new_n2891_));
NAND2X1 NAND2X1_33 ( .A(REG3_REG_7_), .B(_abc_40319_new_n733_), .Y(_abc_40319_new_n734_));
NAND2X1 NAND2X1_330 ( .A(_abc_40319_new_n2543_), .B(_abc_40319_new_n2892_), .Y(_abc_40319_new_n2893_));
NAND2X1 NAND2X1_331 ( .A(_abc_40319_new_n2919_), .B(_abc_40319_new_n2916_), .Y(_abc_40319_new_n2920_));
NAND2X1 NAND2X1_332 ( .A(_abc_40319_new_n2524_), .B(_abc_40319_new_n2945_), .Y(_abc_40319_new_n2946_));
NAND2X1 NAND2X1_333 ( .A(ADDR_REG_19_), .B(_abc_40319_new_n2539_), .Y(_abc_40319_new_n2951_));
NAND2X1 NAND2X1_334 ( .A(_abc_40319_new_n2958_), .B(_abc_40319_new_n2956_), .Y(_abc_40319_new_n2959_));
NAND2X1 NAND2X1_335 ( .A(_abc_40319_new_n2955_), .B(_abc_40319_new_n2960_), .Y(_abc_40319_new_n2961_));
NAND2X1 NAND2X1_336 ( .A(_abc_40319_new_n895_), .B(_abc_40319_new_n922_), .Y(_abc_40319_new_n2962_));
NAND2X1 NAND2X1_337 ( .A(_abc_40319_new_n825_), .B(_abc_40319_new_n2963_), .Y(_abc_40319_new_n2964_));
NAND2X1 NAND2X1_338 ( .A(_abc_40319_new_n1938_), .B(_abc_40319_new_n2965_), .Y(_abc_40319_new_n2966_));
NAND2X1 NAND2X1_339 ( .A(_abc_40319_new_n2388_), .B(_abc_40319_new_n2967_), .Y(_abc_40319_new_n2968_));
NAND2X1 NAND2X1_34 ( .A(_abc_40319_new_n736_), .B(_abc_40319_new_n734_), .Y(_abc_40319_new_n737_));
NAND2X1 NAND2X1_340 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n2980_), .Y(_abc_40319_new_n2981_));
NAND2X1 NAND2X1_341 ( .A(_abc_40319_new_n2987_), .B(_abc_40319_new_n2960_), .Y(_abc_40319_new_n2988_));
NAND2X1 NAND2X1_342 ( .A(_abc_40319_new_n2996_), .B(_abc_40319_new_n2997_), .Y(_abc_40319_new_n2998_));
NAND2X1 NAND2X1_343 ( .A(_abc_40319_new_n3001_), .B(_abc_40319_new_n2998_), .Y(n968));
NAND2X1 NAND2X1_344 ( .A(_abc_40319_new_n3045_), .B(_abc_40319_new_n3052_), .Y(_abc_40319_new_n3053_));
NAND2X1 NAND2X1_345 ( .A(_abc_40319_new_n3065_), .B(_abc_40319_new_n3063_), .Y(_abc_40319_new_n3066_));
NAND2X1 NAND2X1_346 ( .A(_abc_40319_new_n3073_), .B(_abc_40319_new_n3018_), .Y(_abc_40319_new_n3074_));
NAND2X1 NAND2X1_347 ( .A(_abc_40319_new_n3075_), .B(_abc_40319_new_n3071_), .Y(_abc_40319_new_n3076_));
NAND2X1 NAND2X1_348 ( .A(_abc_40319_new_n1080_), .B(_abc_40319_new_n1077_), .Y(_abc_40319_new_n3087_));
NAND2X1 NAND2X1_349 ( .A(_abc_40319_new_n3090_), .B(_abc_40319_new_n3081_), .Y(_abc_40319_new_n3091_));
NAND2X1 NAND2X1_35 ( .A(_abc_40319_new_n739_), .B(_abc_40319_new_n725_), .Y(_abc_40319_new_n740_));
NAND2X1 NAND2X1_350 ( .A(_abc_40319_new_n3091_), .B(_abc_40319_new_n3089_), .Y(_abc_40319_new_n3092_));
NAND2X1 NAND2X1_351 ( .A(_abc_40319_new_n2121_), .B(_abc_40319_new_n3096_), .Y(_abc_40319_new_n3097_));
NAND2X1 NAND2X1_352 ( .A(_abc_40319_new_n3095_), .B(_abc_40319_new_n3097_), .Y(_abc_40319_new_n3109_));
NAND2X1 NAND2X1_353 ( .A(_abc_40319_new_n2446_), .B(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3110_));
NAND2X1 NAND2X1_354 ( .A(REG2_REG_28_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3117_));
NAND2X1 NAND2X1_355 ( .A(_abc_40319_new_n3124_), .B(_abc_40319_new_n3123_), .Y(_abc_40319_new_n3125_));
NAND2X1 NAND2X1_356 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3125_), .Y(_abc_40319_new_n3134_));
NAND2X1 NAND2X1_357 ( .A(_abc_40319_new_n2996_), .B(_abc_40319_new_n3136_), .Y(_abc_40319_new_n3137_));
NAND2X1 NAND2X1_358 ( .A(REG2_REG_27_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3142_));
NAND2X1 NAND2X1_359 ( .A(_abc_40319_new_n2125_), .B(_abc_40319_new_n3152_), .Y(_abc_40319_new_n3153_));
NAND2X1 NAND2X1_36 ( .A(_abc_40319_new_n663_), .B(_abc_40319_new_n742_), .Y(_abc_40319_new_n743_));
NAND2X1 NAND2X1_360 ( .A(_abc_40319_new_n3151_), .B(_abc_40319_new_n3153_), .Y(_abc_40319_new_n3154_));
NAND2X1 NAND2X1_361 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3154_), .Y(_abc_40319_new_n3159_));
NAND2X1 NAND2X1_362 ( .A(nRESET_G), .B(_abc_40319_new_n3166_), .Y(_abc_40319_new_n3167_));
NAND2X1 NAND2X1_363 ( .A(_abc_40319_new_n3159_), .B(_abc_40319_new_n3170_), .Y(_abc_40319_new_n3171_));
NAND2X1 NAND2X1_364 ( .A(_abc_40319_new_n2130_), .B(_abc_40319_new_n3174_), .Y(_abc_40319_new_n3175_));
NAND2X1 NAND2X1_365 ( .A(_abc_40319_new_n3175_), .B(_abc_40319_new_n3176_), .Y(_abc_40319_new_n3177_));
NAND2X1 NAND2X1_366 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3177_), .Y(_abc_40319_new_n3189_));
NAND2X1 NAND2X1_367 ( .A(_abc_40319_new_n3189_), .B(_abc_40319_new_n3199_), .Y(_abc_40319_new_n3200_));
NAND2X1 NAND2X1_368 ( .A(_abc_40319_new_n3101_), .B(_abc_40319_new_n3204_), .Y(_abc_40319_new_n3205_));
NAND2X1 NAND2X1_369 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3204_), .Y(_abc_40319_new_n3210_));
NAND2X1 NAND2X1_37 ( .A(IR_REG_31_), .B(_abc_40319_new_n747_), .Y(_abc_40319_new_n748_));
NAND2X1 NAND2X1_370 ( .A(nRESET_G), .B(_abc_40319_new_n3215_), .Y(_abc_40319_new_n3216_));
NAND2X1 NAND2X1_371 ( .A(_abc_40319_new_n3210_), .B(_abc_40319_new_n3219_), .Y(_abc_40319_new_n3220_));
NAND2X1 NAND2X1_372 ( .A(_abc_40319_new_n3076_), .B(_abc_40319_new_n3027_), .Y(_abc_40319_new_n3228_));
NAND2X1 NAND2X1_373 ( .A(_abc_40319_new_n3101_), .B(_abc_40319_new_n3229_), .Y(_abc_40319_new_n3238_));
NAND2X1 NAND2X1_374 ( .A(_abc_40319_new_n3101_), .B(_abc_40319_new_n3255_), .Y(_abc_40319_new_n3258_));
NAND2X1 NAND2X1_375 ( .A(_abc_40319_new_n2960_), .B(_abc_40319_new_n3260_), .Y(_abc_40319_new_n3261_));
NAND2X1 NAND2X1_376 ( .A(_abc_40319_new_n2960_), .B(_abc_40319_new_n3273_), .Y(_abc_40319_new_n3274_));
NAND2X1 NAND2X1_377 ( .A(REG2_REG_21_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3275_));
NAND2X1 NAND2X1_378 ( .A(_abc_40319_new_n3101_), .B(_abc_40319_new_n3287_), .Y(_abc_40319_new_n3288_));
NAND2X1 NAND2X1_379 ( .A(_abc_40319_new_n2960_), .B(_abc_40319_new_n3294_), .Y(_abc_40319_new_n3295_));
NAND2X1 NAND2X1_38 ( .A(_abc_40319_new_n574_), .B(_abc_40319_new_n744_), .Y(_abc_40319_new_n757_));
NAND2X1 NAND2X1_380 ( .A(REG2_REG_20_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3296_));
NAND2X1 NAND2X1_381 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3287_), .Y(_abc_40319_new_n3297_));
NAND2X1 NAND2X1_382 ( .A(_abc_40319_new_n1159_), .B(_abc_40319_new_n2973_), .Y(_abc_40319_new_n3298_));
NAND2X1 NAND2X1_383 ( .A(_abc_40319_new_n3299_), .B(_abc_40319_new_n3249_), .Y(_abc_40319_new_n3300_));
NAND2X1 NAND2X1_384 ( .A(_abc_40319_new_n2960_), .B(_abc_40319_new_n3312_), .Y(_abc_40319_new_n3313_));
NAND2X1 NAND2X1_385 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3308_), .Y(_abc_40319_new_n3314_));
NAND2X1 NAND2X1_386 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3324_), .Y(_abc_40319_new_n3330_));
NAND2X1 NAND2X1_387 ( .A(_abc_40319_new_n3339_), .B(_abc_40319_new_n3330_), .Y(_abc_40319_new_n3340_));
NAND2X1 NAND2X1_388 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3344_), .Y(_abc_40319_new_n3365_));
NAND2X1 NAND2X1_389 ( .A(_abc_40319_new_n1261_), .B(_abc_40319_new_n2971_), .Y(_abc_40319_new_n3377_));
NAND2X1 NAND2X1_39 ( .A(_abc_40319_new_n678_), .B(_abc_40319_new_n574_), .Y(_abc_40319_new_n758_));
NAND2X1 NAND2X1_390 ( .A(_abc_40319_new_n2996_), .B(_abc_40319_new_n3379_), .Y(_abc_40319_new_n3380_));
NAND2X1 NAND2X1_391 ( .A(_abc_40319_new_n1176_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3389_));
NAND2X1 NAND2X1_392 ( .A(_abc_40319_new_n2996_), .B(_abc_40319_new_n3395_), .Y(_abc_40319_new_n3396_));
NAND2X1 NAND2X1_393 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3398_), .Y(_abc_40319_new_n3399_));
NAND2X1 NAND2X1_394 ( .A(_abc_40319_new_n1225_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3403_));
NAND2X1 NAND2X1_395 ( .A(_abc_40319_new_n3399_), .B(_abc_40319_new_n3404_), .Y(_abc_40319_new_n3405_));
NAND2X1 NAND2X1_396 ( .A(_abc_40319_new_n2996_), .B(_abc_40319_new_n3436_), .Y(_abc_40319_new_n3437_));
NAND2X1 NAND2X1_397 ( .A(_abc_40319_new_n3101_), .B(_abc_40319_new_n3463_), .Y(_abc_40319_new_n3470_));
NAND2X1 NAND2X1_398 ( .A(_abc_40319_new_n2996_), .B(_abc_40319_new_n3485_), .Y(_abc_40319_new_n3486_));
NAND2X1 NAND2X1_399 ( .A(_abc_40319_new_n3502_), .B(_abc_40319_new_n3459_), .Y(_abc_40319_new_n3503_));
NAND2X1 NAND2X1_4 ( .A(_abc_40319_new_n562_), .B(_abc_40319_new_n564_), .Y(_abc_40319_new_n565_));
NAND2X1 NAND2X1_40 ( .A(_abc_40319_new_n757_), .B(_abc_40319_new_n760_), .Y(_abc_40319_new_n761_));
NAND2X1 NAND2X1_400 ( .A(_abc_40319_new_n3101_), .B(_abc_40319_new_n3514_), .Y(_abc_40319_new_n3515_));
NAND2X1 NAND2X1_401 ( .A(_abc_40319_new_n3518_), .B(_abc_40319_new_n2996_), .Y(_abc_40319_new_n3519_));
NAND2X1 NAND2X1_402 ( .A(_abc_40319_new_n3537_), .B(_abc_40319_new_n2996_), .Y(_abc_40319_new_n3538_));
NAND2X1 NAND2X1_403 ( .A(_abc_40319_new_n3539_), .B(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3540_));
NAND2X1 NAND2X1_404 ( .A(_abc_40319_new_n3554_), .B(_abc_40319_new_n2996_), .Y(_abc_40319_new_n3555_));
NAND2X1 NAND2X1_405 ( .A(_abc_40319_new_n951_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3556_));
NAND2X1 NAND2X1_406 ( .A(_abc_40319_new_n3571_), .B(_abc_40319_new_n2996_), .Y(_abc_40319_new_n3572_));
NAND2X1 NAND2X1_407 ( .A(_abc_40319_new_n3572_), .B(_abc_40319_new_n3576_), .Y(_abc_40319_new_n3577_));
NAND2X1 NAND2X1_408 ( .A(_abc_40319_new_n3597_), .B(_abc_40319_new_n3601_), .Y(_abc_40319_new_n3602_));
NAND2X1 NAND2X1_409 ( .A(_abc_40319_new_n3605_), .B(_abc_40319_new_n2964_), .Y(_abc_40319_new_n3606_));
NAND2X1 NAND2X1_41 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n526_), .Y(_abc_40319_new_n763_));
NAND2X1 NAND2X1_410 ( .A(_abc_40319_new_n3604_), .B(_abc_40319_new_n3610_), .Y(n833));
NAND2X1 NAND2X1_411 ( .A(_abc_40319_new_n3647_), .B(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3648_));
NAND2X1 NAND2X1_412 ( .A(_abc_40319_new_n3649_), .B(_abc_40319_new_n3651_), .Y(n818));
NAND2X1 NAND2X1_413 ( .A(D_REG_31_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3659_));
NAND2X1 NAND2X1_414 ( .A(D_REG_30_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3661_));
NAND2X1 NAND2X1_415 ( .A(D_REG_29_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3663_));
NAND2X1 NAND2X1_416 ( .A(D_REG_28_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3665_));
NAND2X1 NAND2X1_417 ( .A(D_REG_27_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3667_));
NAND2X1 NAND2X1_418 ( .A(D_REG_26_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3669_));
NAND2X1 NAND2X1_419 ( .A(D_REG_25_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3671_));
NAND2X1 NAND2X1_42 ( .A(IR_REG_31_), .B(_abc_40319_new_n765_), .Y(_abc_40319_new_n766_));
NAND2X1 NAND2X1_420 ( .A(D_REG_24_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3673_));
NAND2X1 NAND2X1_421 ( .A(D_REG_23_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3675_));
NAND2X1 NAND2X1_422 ( .A(D_REG_22_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3677_));
NAND2X1 NAND2X1_423 ( .A(D_REG_21_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3679_));
NAND2X1 NAND2X1_424 ( .A(D_REG_20_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3681_));
NAND2X1 NAND2X1_425 ( .A(D_REG_19_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3683_));
NAND2X1 NAND2X1_426 ( .A(D_REG_18_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3685_));
NAND2X1 NAND2X1_427 ( .A(D_REG_17_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3687_));
NAND2X1 NAND2X1_428 ( .A(D_REG_16_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3689_));
NAND2X1 NAND2X1_429 ( .A(D_REG_15_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3691_));
NAND2X1 NAND2X1_43 ( .A(REG1_REG_5_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n771_));
NAND2X1 NAND2X1_430 ( .A(D_REG_14_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3693_));
NAND2X1 NAND2X1_431 ( .A(D_REG_13_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3695_));
NAND2X1 NAND2X1_432 ( .A(D_REG_12_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3697_));
NAND2X1 NAND2X1_433 ( .A(D_REG_11_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3699_));
NAND2X1 NAND2X1_434 ( .A(D_REG_10_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3701_));
NAND2X1 NAND2X1_435 ( .A(D_REG_9_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3703_));
NAND2X1 NAND2X1_436 ( .A(D_REG_8_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3705_));
NAND2X1 NAND2X1_437 ( .A(D_REG_7_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3707_));
NAND2X1 NAND2X1_438 ( .A(D_REG_6_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3709_));
NAND2X1 NAND2X1_439 ( .A(D_REG_5_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3711_));
NAND2X1 NAND2X1_44 ( .A(_abc_40319_new_n780_), .B(_abc_40319_new_n732_), .Y(_abc_40319_new_n781_));
NAND2X1 NAND2X1_440 ( .A(D_REG_4_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3713_));
NAND2X1 NAND2X1_441 ( .A(D_REG_3_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3715_));
NAND2X1 NAND2X1_442 ( .A(D_REG_2_), .B(_abc_40319_new_n3658_), .Y(_abc_40319_new_n3717_));
NAND2X1 NAND2X1_443 ( .A(_abc_40319_new_n3723_), .B(_abc_40319_new_n3724_), .Y(n323));
NAND2X1 NAND2X1_444 ( .A(IR_REG_28_), .B(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3727_));
NAND2X1 NAND2X1_445 ( .A(_abc_40319_new_n542_), .B(_abc_40319_new_n558_), .Y(_abc_40319_new_n3742_));
NAND2X1 NAND2X1_446 ( .A(_abc_40319_new_n3753_), .B(_abc_40319_new_n3754_), .Y(n283));
NAND2X1 NAND2X1_447 ( .A(_abc_40319_new_n3763_), .B(_abc_40319_new_n3764_), .Y(n268));
NAND2X1 NAND2X1_448 ( .A(_abc_40319_new_n3769_), .B(_abc_40319_new_n3771_), .Y(n258));
NAND2X1 NAND2X1_449 ( .A(_abc_40319_new_n3776_), .B(_abc_40319_new_n3777_), .Y(n248));
NAND2X1 NAND2X1_45 ( .A(_abc_40319_new_n757_), .B(_abc_40319_new_n789_), .Y(_abc_40319_new_n790_));
NAND2X1 NAND2X1_450 ( .A(IR_REG_12_), .B(_abc_40319_new_n3720_), .Y(_abc_40319_new_n3782_));
NAND2X1 NAND2X1_451 ( .A(_abc_40319_new_n3793_), .B(_abc_40319_new_n3794_), .Y(n223));
NAND2X1 NAND2X1_452 ( .A(_abc_40319_new_n3796_), .B(_abc_40319_new_n3797_), .Y(n218));
NAND2X1 NAND2X1_453 ( .A(_abc_40319_new_n3799_), .B(_abc_40319_new_n3800_), .Y(n213));
NAND2X1 NAND2X1_454 ( .A(_abc_40319_new_n3802_), .B(_abc_40319_new_n3803_), .Y(n208));
NAND2X1 NAND2X1_455 ( .A(_abc_40319_new_n3808_), .B(_abc_40319_new_n3809_), .Y(n198));
NAND2X1 NAND2X1_456 ( .A(_abc_40319_new_n3829_), .B(_abc_40319_new_n3835_), .Y(_abc_40319_new_n3836_));
NAND2X1 NAND2X1_457 ( .A(_abc_40319_new_n2266_), .B(_abc_40319_new_n3842_), .Y(_abc_40319_new_n3843_));
NAND2X1 NAND2X1_458 ( .A(_abc_40319_new_n3841_), .B(_abc_40319_new_n3843_), .Y(_abc_40319_new_n3844_));
NAND2X1 NAND2X1_459 ( .A(_abc_40319_new_n3849_), .B(_abc_40319_new_n3846_), .Y(_abc_40319_new_n3850_));
NAND2X1 NAND2X1_46 ( .A(IR_REG_31_), .B(_abc_40319_new_n794_), .Y(_abc_40319_new_n795_));
NAND2X1 NAND2X1_460 ( .A(_abc_40319_new_n3837_), .B(_abc_40319_new_n3851_), .Y(_abc_40319_new_n3852_));
NAND2X1 NAND2X1_461 ( .A(_abc_40319_new_n2960_), .B(_abc_40319_new_n3852_), .Y(_abc_40319_new_n3853_));
NAND2X1 NAND2X1_462 ( .A(_abc_40319_new_n3133_), .B(_abc_40319_new_n3844_), .Y(_abc_40319_new_n3854_));
NAND2X1 NAND2X1_463 ( .A(REG3_REG_17_), .B(_abc_40319_new_n3861_), .Y(_abc_40319_new_n3862_));
NAND2X1 NAND2X1_464 ( .A(_abc_40319_new_n3893_), .B(_abc_40319_new_n2237_), .Y(_abc_40319_new_n3900_));
NAND2X1 NAND2X1_465 ( .A(_abc_40319_new_n3893_), .B(_abc_40319_new_n3567_), .Y(_abc_40319_new_n3920_));
NAND2X1 NAND2X1_466 ( .A(_abc_40319_new_n3893_), .B(_abc_40319_new_n3553_), .Y(_abc_40319_new_n3932_));
NAND2X1 NAND2X1_467 ( .A(_abc_40319_new_n3536_), .B(_abc_40319_new_n2968_), .Y(_abc_40319_new_n3937_));
NAND2X1 NAND2X1_468 ( .A(_abc_40319_new_n3939_), .B(_abc_40319_new_n3535_), .Y(_abc_40319_new_n3940_));
NAND2X1 NAND2X1_469 ( .A(_abc_40319_new_n3951_), .B(_abc_40319_new_n3501_), .Y(_abc_40319_new_n3952_));
NAND2X1 NAND2X1_47 ( .A(_abc_40319_new_n806_), .B(_abc_40319_new_n727_), .Y(_abc_40319_new_n807_));
NAND2X1 NAND2X1_470 ( .A(_abc_40319_new_n3961_), .B(_abc_40319_new_n3960_), .Y(_abc_40319_new_n3962_));
NAND2X1 NAND2X1_471 ( .A(_abc_40319_new_n3620_), .B(_abc_40319_new_n3417_), .Y(_abc_40319_new_n3977_));
NAND2X1 NAND2X1_472 ( .A(_abc_40319_new_n3982_), .B(_abc_40319_new_n3983_), .Y(_abc_40319_new_n3984_));
NAND2X1 NAND2X1_473 ( .A(_abc_40319_new_n3893_), .B(_abc_40319_new_n3344_), .Y(_abc_40319_new_n3997_));
NAND2X1 NAND2X1_474 ( .A(_abc_40319_new_n4007_), .B(_abc_40319_new_n4008_), .Y(_abc_40319_new_n4009_));
NAND2X1 NAND2X1_475 ( .A(_abc_40319_new_n3620_), .B(_abc_40319_new_n3251_), .Y(_abc_40319_new_n4020_));
NAND2X1 NAND2X1_476 ( .A(_abc_40319_new_n3893_), .B(_abc_40319_new_n3255_), .Y(_abc_40319_new_n4021_));
NAND2X1 NAND2X1_477 ( .A(_abc_40319_new_n3620_), .B(_abc_40319_new_n3136_), .Y(_abc_40319_new_n4052_));
NAND2X1 NAND2X1_478 ( .A(_abc_40319_new_n3893_), .B(_abc_40319_new_n3844_), .Y(_abc_40319_new_n4068_));
NAND2X1 NAND2X1_479 ( .A(_abc_40319_new_n4073_), .B(_abc_40319_new_n4072_), .Y(n643));
NAND2X1 NAND2X1_48 ( .A(_abc_40319_new_n750_), .B(_abc_40319_new_n574_), .Y(_abc_40319_new_n812_));
NAND2X1 NAND2X1_480 ( .A(_abc_40319_new_n4082_), .B(_abc_40319_new_n4081_), .Y(n653));
NAND2X1 NAND2X1_481 ( .A(_abc_40319_new_n656_), .B(_abc_40319_new_n3887_), .Y(_abc_40319_new_n4084_));
NAND2X1 NAND2X1_482 ( .A(_abc_40319_new_n4134_), .B(_abc_40319_new_n4133_), .Y(n763));
NAND2X1 NAND2X1_483 ( .A(_abc_40319_new_n4151_), .B(_abc_40319_new_n4150_), .Y(n803));
NAND2X1 NAND2X1_484 ( .A(_abc_40319_new_n4156_), .B(_abc_40319_new_n4155_), .Y(n813));
NAND2X1 NAND2X1_49 ( .A(_abc_40319_new_n811_), .B(_abc_40319_new_n815_), .Y(_abc_40319_new_n817_));
NAND2X1 NAND2X1_5 ( .A(IR_REG_31_), .B(_abc_40319_new_n565_), .Y(_abc_40319_new_n566_));
NAND2X1 NAND2X1_50 ( .A(IR_REG_3_), .B(_abc_40319_new_n546_), .Y(_abc_40319_new_n818_));
NAND2X1 NAND2X1_51 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n818_), .Y(_abc_40319_new_n819_));
NAND2X1 NAND2X1_52 ( .A(IR_REG_31_), .B(_abc_40319_new_n819_), .Y(_abc_40319_new_n820_));
NAND2X1 NAND2X1_53 ( .A(_abc_40319_new_n831_), .B(_abc_40319_new_n830_), .Y(_abc_40319_new_n832_));
NAND2X1 NAND2X1_54 ( .A(_abc_40319_new_n840_), .B(_abc_40319_new_n841_), .Y(_abc_40319_new_n842_));
NAND2X1 NAND2X1_55 ( .A(_abc_40319_new_n867_), .B(_abc_40319_new_n863_), .Y(_abc_40319_new_n868_));
NAND2X1 NAND2X1_56 ( .A(IR_REG_1_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n874_));
NAND2X1 NAND2X1_57 ( .A(_abc_40319_new_n879_), .B(_abc_40319_new_n878_), .Y(_abc_40319_new_n880_));
NAND2X1 NAND2X1_58 ( .A(REG3_REG_1_), .B(_abc_40319_new_n727_), .Y(_abc_40319_new_n888_));
NAND2X1 NAND2X1_59 ( .A(_abc_40319_new_n887_), .B(_abc_40319_new_n888_), .Y(_abc_40319_new_n889_));
NAND2X1 NAND2X1_6 ( .A(IR_REG_26_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n570_));
NAND2X1 NAND2X1_60 ( .A(_abc_40319_new_n899_), .B(_abc_40319_new_n891_), .Y(_abc_40319_new_n900_));
NAND2X1 NAND2X1_61 ( .A(_abc_40319_new_n881_), .B(_abc_40319_new_n900_), .Y(_abc_40319_new_n901_));
NAND2X1 NAND2X1_62 ( .A(_abc_40319_new_n574_), .B(_abc_40319_new_n904_), .Y(_abc_40319_new_n905_));
NAND2X1 NAND2X1_63 ( .A(REG3_REG_0_), .B(_abc_40319_new_n727_), .Y(_abc_40319_new_n910_));
NAND2X1 NAND2X1_64 ( .A(_abc_40319_new_n745_), .B(_abc_40319_new_n916_), .Y(_abc_40319_new_n917_));
NAND2X1 NAND2X1_65 ( .A(_abc_40319_new_n857_), .B(_abc_40319_new_n851_), .Y(_abc_40319_new_n932_));
NAND2X1 NAND2X1_66 ( .A(_abc_40319_new_n792_), .B(_abc_40319_new_n936_), .Y(_abc_40319_new_n937_));
NAND2X1 NAND2X1_67 ( .A(_abc_40319_new_n685_), .B(_abc_40319_new_n550_), .Y(_abc_40319_new_n938_));
NAND2X1 NAND2X1_68 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n685_), .Y(_abc_40319_new_n941_));
NAND2X1 NAND2X1_69 ( .A(_abc_40319_new_n728_), .B(_abc_40319_new_n732_), .Y(_abc_40319_new_n947_));
NAND2X1 NAND2X1_7 ( .A(_abc_40319_new_n560_), .B(_abc_40319_new_n573_), .Y(_abc_40319_new_n574_));
NAND2X1 NAND2X1_70 ( .A(_abc_40319_new_n757_), .B(_abc_40319_new_n960_), .Y(_abc_40319_new_n961_));
NAND2X1 NAND2X1_71 ( .A(_abc_40319_new_n963_), .B(_abc_40319_new_n964_), .Y(_abc_40319_new_n965_));
NAND2X1 NAND2X1_72 ( .A(_abc_40319_new_n985_), .B(_abc_40319_new_n986_), .Y(_abc_40319_new_n987_));
NAND2X1 NAND2X1_73 ( .A(_abc_40319_new_n992_), .B(_abc_40319_new_n1004_), .Y(_abc_40319_new_n1005_));
NAND2X1 NAND2X1_74 ( .A(REG3_REG_12_), .B(REG3_REG_13_), .Y(_abc_40319_new_n1027_));
NAND2X1 NAND2X1_75 ( .A(REG3_REG_16_), .B(REG3_REG_17_), .Y(_abc_40319_new_n1030_));
NAND2X1 NAND2X1_76 ( .A(REG3_REG_18_), .B(_abc_40319_new_n1031_), .Y(_abc_40319_new_n1032_));
NAND2X1 NAND2X1_77 ( .A(REG3_REG_27_), .B(_abc_40319_new_n1039_), .Y(_abc_40319_new_n1040_));
NAND2X1 NAND2X1_78 ( .A(_abc_40319_new_n1038_), .B(_abc_40319_new_n1040_), .Y(_abc_40319_new_n1041_));
NAND2X1 NAND2X1_79 ( .A(REG1_REG_27_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n1043_));
NAND2X1 NAND2X1_8 ( .A(_abc_40319_new_n556_), .B(_abc_40319_new_n553_), .Y(_abc_40319_new_n576_));
NAND2X1 NAND2X1_80 ( .A(_abc_40319_new_n1047_), .B(_abc_40319_new_n1049_), .Y(_abc_40319_new_n1051_));
NAND2X1 NAND2X1_81 ( .A(REG3_REG_24_), .B(_abc_40319_new_n1036_), .Y(_abc_40319_new_n1058_));
NAND2X1 NAND2X1_82 ( .A(REG1_REG_26_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n1062_));
NAND2X1 NAND2X1_83 ( .A(_abc_40319_new_n1064_), .B(_abc_40319_new_n1060_), .Y(_abc_40319_new_n1065_));
NAND2X1 NAND2X1_84 ( .A(_abc_40319_new_n1066_), .B(_abc_40319_new_n1068_), .Y(_abc_40319_new_n1069_));
NAND2X1 NAND2X1_85 ( .A(_abc_40319_new_n1057_), .B(_abc_40319_new_n1058_), .Y(_abc_40319_new_n1071_));
NAND2X1 NAND2X1_86 ( .A(_abc_40319_new_n1037_), .B(_abc_40319_new_n1071_), .Y(_abc_40319_new_n1072_));
NAND2X1 NAND2X1_87 ( .A(REG2_REG_25_), .B(_abc_40319_new_n715_), .Y(_abc_40319_new_n1074_));
NAND2X1 NAND2X1_88 ( .A(REG2_REG_24_), .B(_abc_40319_new_n715_), .Y(_abc_40319_new_n1090_));
NAND2X1 NAND2X1_89 ( .A(_abc_40319_new_n1079_), .B(_abc_40319_new_n1082_), .Y(_abc_40319_new_n1103_));
NAND2X1 NAND2X1_9 ( .A(_abc_40319_new_n578_), .B(_abc_40319_new_n577_), .Y(_abc_40319_new_n579_));
NAND2X1 NAND2X1_90 ( .A(REG1_REG_23_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n1112_));
NAND2X1 NAND2X1_91 ( .A(_abc_40319_new_n1116_), .B(_abc_40319_new_n1119_), .Y(_abc_40319_new_n1121_));
NAND2X1 NAND2X1_92 ( .A(REG3_REG_20_), .B(_abc_40319_new_n1033_), .Y(_abc_40319_new_n1126_));
NAND2X1 NAND2X1_93 ( .A(_abc_40319_new_n1127_), .B(_abc_40319_new_n1035_), .Y(_abc_40319_new_n1128_));
NAND2X1 NAND2X1_94 ( .A(REG1_REG_22_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n1131_));
NAND2X1 NAND2X1_95 ( .A(REG2_REG_22_), .B(_abc_40319_new_n715_), .Y(_abc_40319_new_n1132_));
NAND2X1 NAND2X1_96 ( .A(_abc_40319_new_n1136_), .B(_abc_40319_new_n1140_), .Y(_abc_40319_new_n1141_));
NAND2X1 NAND2X1_97 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n594_), .Y(_abc_40319_new_n1145_));
NAND2X1 NAND2X1_98 ( .A(_abc_40319_new_n1152_), .B(_abc_40319_new_n1032_), .Y(_abc_40319_new_n1153_));
NAND2X1 NAND2X1_99 ( .A(_abc_40319_new_n1158_), .B(_abc_40319_new_n1162_), .Y(_abc_40319_new_n1163_));
NAND3X1 NAND3X1_1 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n525_), .C(_abc_40319_new_n526_), .Y(_abc_40319_new_n527_));
NAND3X1 NAND3X1_10 ( .A(_abc_40319_new_n561_), .B(_abc_40319_new_n541_), .C(_abc_40319_new_n532_), .Y(_abc_40319_new_n562_));
NAND3X1 NAND3X1_100 ( .A(_abc_40319_new_n2190_), .B(_abc_40319_new_n2186_), .C(_abc_40319_new_n2181_), .Y(_abc_40319_new_n2191_));
NAND3X1 NAND3X1_101 ( .A(_abc_40319_new_n2143_), .B(_abc_40319_new_n2211_), .C(_abc_40319_new_n2172_), .Y(_abc_40319_new_n2212_));
NAND3X1 NAND3X1_102 ( .A(_abc_40319_new_n2231_), .B(_abc_40319_new_n2235_), .C(_abc_40319_new_n2226_), .Y(_abc_40319_new_n2236_));
NAND3X1 NAND3X1_103 ( .A(_abc_40319_new_n2216_), .B(_abc_40319_new_n2220_), .C(_abc_40319_new_n2252_), .Y(_abc_40319_new_n2253_));
NAND3X1 NAND3X1_104 ( .A(_abc_40319_new_n2130_), .B(_abc_40319_new_n2134_), .C(_abc_40319_new_n2255_), .Y(_abc_40319_new_n2256_));
NAND3X1 NAND3X1_105 ( .A(_abc_40319_new_n2121_), .B(_abc_40319_new_n2268_), .C(_abc_40319_new_n2257_), .Y(_abc_40319_new_n2269_));
NAND3X1 NAND3X1_106 ( .A(_abc_40319_new_n1967_), .B(_abc_40319_new_n1935_), .C(_abc_40319_new_n1929_), .Y(_abc_40319_new_n2289_));
NAND3X1 NAND3X1_107 ( .A(_abc_40319_new_n1953_), .B(_abc_40319_new_n2289_), .C(_abc_40319_new_n2288_), .Y(_abc_40319_new_n2290_));
NAND3X1 NAND3X1_108 ( .A(_abc_40319_new_n2118_), .B(_abc_40319_new_n2307_), .C(_abc_40319_new_n2309_), .Y(_abc_40319_new_n2310_));
NAND3X1 NAND3X1_109 ( .A(_abc_40319_new_n2135_), .B(_abc_40319_new_n2312_), .C(_abc_40319_new_n2131_), .Y(_abc_40319_new_n2313_));
NAND3X1 NAND3X1_11 ( .A(_abc_40319_new_n590_), .B(_abc_40319_new_n541_), .C(_abc_40319_new_n532_), .Y(_abc_40319_new_n591_));
NAND3X1 NAND3X1_110 ( .A(_abc_40319_new_n2313_), .B(_abc_40319_new_n2314_), .C(_abc_40319_new_n2316_), .Y(_abc_40319_new_n2317_));
NAND3X1 NAND3X1_111 ( .A(_abc_40319_new_n2359_), .B(_abc_40319_new_n2363_), .C(_abc_40319_new_n2364_), .Y(_abc_40319_new_n2365_));
NAND3X1 NAND3X1_112 ( .A(_abc_40319_new_n2369_), .B(_abc_40319_new_n2371_), .C(_abc_40319_new_n2370_), .Y(_abc_40319_new_n2372_));
NAND3X1 NAND3X1_113 ( .A(_abc_40319_new_n2377_), .B(_abc_40319_new_n2373_), .C(_abc_40319_new_n2318_), .Y(_abc_40319_new_n2378_));
NAND3X1 NAND3X1_114 ( .A(_abc_40319_new_n2378_), .B(_abc_40319_new_n2372_), .C(_abc_40319_new_n2376_), .Y(_abc_40319_new_n2379_));
NAND3X1 NAND3X1_115 ( .A(_abc_40319_new_n2371_), .B(_abc_40319_new_n2391_), .C(_abc_40319_new_n2370_), .Y(_abc_40319_new_n2392_));
NAND3X1 NAND3X1_116 ( .A(_abc_40319_new_n2178_), .B(_abc_40319_new_n2348_), .C(_abc_40319_new_n2370_), .Y(_abc_40319_new_n2398_));
NAND3X1 NAND3X1_117 ( .A(_abc_40319_new_n2392_), .B(_abc_40319_new_n2398_), .C(_abc_40319_new_n2397_), .Y(_abc_40319_new_n2399_));
NAND3X1 NAND3X1_118 ( .A(_abc_40319_new_n2345_), .B(_abc_40319_new_n2368_), .C(_abc_40319_new_n2400_), .Y(_abc_40319_new_n2401_));
NAND3X1 NAND3X1_119 ( .A(_abc_40319_new_n2154_), .B(_abc_40319_new_n2307_), .C(_abc_40319_new_n2309_), .Y(_abc_40319_new_n2418_));
NAND3X1 NAND3X1_12 ( .A(_abc_40319_new_n534_), .B(_abc_40319_new_n594_), .C(_abc_40319_new_n595_), .Y(_abc_40319_new_n596_));
NAND3X1 NAND3X1_120 ( .A(_abc_40319_new_n2152_), .B(_abc_40319_new_n2174_), .C(_abc_40319_new_n2118_), .Y(_abc_40319_new_n2422_));
NAND3X1 NAND3X1_121 ( .A(_abc_40319_new_n2338_), .B(_abc_40319_new_n2428_), .C(_abc_40319_new_n2426_), .Y(_abc_40319_new_n2429_));
NAND3X1 NAND3X1_122 ( .A(_abc_40319_new_n2118_), .B(_abc_40319_new_n2307_), .C(_abc_40319_new_n2430_), .Y(_abc_40319_new_n2431_));
NAND3X1 NAND3X1_123 ( .A(_abc_40319_new_n2420_), .B(_abc_40319_new_n2437_), .C(_abc_40319_new_n2415_), .Y(_abc_40319_new_n2438_));
NAND3X1 NAND3X1_124 ( .A(_abc_40319_new_n2270_), .B(_abc_40319_new_n2441_), .C(_abc_40319_new_n2115_), .Y(_abc_40319_new_n2442_));
NAND3X1 NAND3X1_125 ( .A(_abc_40319_new_n2448_), .B(_abc_40319_new_n2443_), .C(_abc_40319_new_n2444_), .Y(_abc_40319_new_n2449_));
NAND3X1 NAND3X1_126 ( .A(_abc_40319_new_n2457_), .B(_abc_40319_new_n2460_), .C(_abc_40319_new_n2459_), .Y(_abc_40319_new_n2461_));
NAND3X1 NAND3X1_127 ( .A(_abc_40319_new_n2484_), .B(_abc_40319_new_n2374_), .C(_abc_40319_new_n2487_), .Y(_abc_40319_new_n2488_));
NAND3X1 NAND3X1_128 ( .A(_abc_40319_new_n2128_), .B(_abc_40319_new_n2503_), .C(_abc_40319_new_n2498_), .Y(_abc_40319_new_n2504_));
NAND3X1 NAND3X1_129 ( .A(_abc_40319_new_n2452_), .B(_abc_40319_new_n2513_), .C(_abc_40319_new_n2510_), .Y(_abc_40319_new_n2514_));
NAND3X1 NAND3X1_13 ( .A(_abc_40319_new_n543_), .B(_abc_40319_new_n575_), .C(_abc_40319_new_n597_), .Y(_abc_40319_new_n598_));
NAND3X1 NAND3X1_130 ( .A(_abc_40319_new_n2449_), .B(_abc_40319_new_n2518_), .C(_abc_40319_new_n2515_), .Y(_abc_40319_new_n2519_));
NAND3X1 NAND3X1_131 ( .A(_abc_40319_new_n2562_), .B(_abc_40319_new_n2575_), .C(_abc_40319_new_n2561_), .Y(n1046));
NAND3X1 NAND3X1_132 ( .A(_abc_40319_new_n2604_), .B(_abc_40319_new_n2605_), .C(_abc_40319_new_n2561_), .Y(n1038));
NAND3X1 NAND3X1_133 ( .A(_abc_40319_new_n2673_), .B(_abc_40319_new_n2652_), .C(_abc_40319_new_n2650_), .Y(_abc_40319_new_n2674_));
NAND3X1 NAND3X1_134 ( .A(REG1_REG_8_), .B(_abc_40319_new_n2654_), .C(_abc_40319_new_n2674_), .Y(_abc_40319_new_n2677_));
NAND3X1 NAND3X1_135 ( .A(_abc_40319_new_n2685_), .B(_abc_40319_new_n2692_), .C(_abc_40319_new_n2682_), .Y(n1022));
NAND3X1 NAND3X1_136 ( .A(_abc_40319_new_n2702_), .B(_abc_40319_new_n2676_), .C(_abc_40319_new_n2704_), .Y(_abc_40319_new_n2715_));
NAND3X1 NAND3X1_137 ( .A(_abc_40319_new_n1394_), .B(_abc_40319_new_n2701_), .C(_abc_40319_new_n2715_), .Y(_abc_40319_new_n2718_));
NAND3X1 NAND3X1_138 ( .A(_abc_40319_new_n1800_), .B(_abc_40319_new_n2755_), .C(_abc_40319_new_n2757_), .Y(_abc_40319_new_n2758_));
NAND3X1 NAND3X1_139 ( .A(_abc_40319_new_n2717_), .B(_abc_40319_new_n2740_), .C(_abc_40319_new_n2766_), .Y(_abc_40319_new_n2767_));
NAND3X1 NAND3X1_14 ( .A(_abc_40319_new_n532_), .B(_abc_40319_new_n590_), .C(_abc_40319_new_n599_), .Y(_abc_40319_new_n600_));
NAND3X1 NAND3X1_140 ( .A(_abc_40319_new_n2724_), .B(_abc_40319_new_n2749_), .C(_abc_40319_new_n2773_), .Y(_abc_40319_new_n2774_));
NAND3X1 NAND3X1_141 ( .A(_abc_40319_new_n1655_), .B(_abc_40319_new_n2777_), .C(_abc_40319_new_n2779_), .Y(_abc_40319_new_n2780_));
NAND3X1 NAND3X1_142 ( .A(_abc_40319_new_n2742_), .B(_abc_40319_new_n2764_), .C(_abc_40319_new_n2767_), .Y(_abc_40319_new_n2783_));
NAND3X1 NAND3X1_143 ( .A(_abc_40319_new_n1326_), .B(_abc_40319_new_n2762_), .C(_abc_40319_new_n2783_), .Y(_abc_40319_new_n2784_));
NAND3X1 NAND3X1_144 ( .A(_abc_40319_new_n2751_), .B(_abc_40319_new_n2792_), .C(_abc_40319_new_n2774_), .Y(_abc_40319_new_n2793_));
NAND3X1 NAND3X1_145 ( .A(_abc_40319_new_n2815_), .B(_abc_40319_new_n2816_), .C(_abc_40319_new_n2793_), .Y(_abc_40319_new_n2817_));
NAND3X1 NAND3X1_146 ( .A(_abc_40319_new_n2840_), .B(_abc_40319_new_n2841_), .C(_abc_40319_new_n2817_), .Y(_abc_40319_new_n2842_));
NAND3X1 NAND3X1_147 ( .A(_abc_40319_new_n2867_), .B(_abc_40319_new_n2835_), .C(_abc_40319_new_n2842_), .Y(_abc_40319_new_n2868_));
NAND3X1 NAND3X1_148 ( .A(_abc_40319_new_n2862_), .B(_abc_40319_new_n2872_), .C(_abc_40319_new_n2871_), .Y(_abc_40319_new_n2873_));
NAND3X1 NAND3X1_149 ( .A(_abc_40319_new_n2829_), .B(_abc_40319_new_n2857_), .C(_abc_40319_new_n2859_), .Y(_abc_40319_new_n2882_));
NAND3X1 NAND3X1_15 ( .A(_abc_40319_new_n534_), .B(_abc_40319_new_n595_), .C(_abc_40319_new_n532_), .Y(_abc_40319_new_n604_));
NAND3X1 NAND3X1_150 ( .A(_abc_40319_new_n2838_), .B(_abc_40319_new_n2865_), .C(_abc_40319_new_n2868_), .Y(_abc_40319_new_n2888_));
NAND3X1 NAND3X1_151 ( .A(_abc_40319_new_n2831_), .B(_abc_40319_new_n2854_), .C(_abc_40319_new_n2903_), .Y(_abc_40319_new_n2904_));
NAND3X1 NAND3X1_152 ( .A(_abc_40319_new_n2857_), .B(_abc_40319_new_n2902_), .C(_abc_40319_new_n2904_), .Y(_abc_40319_new_n2905_));
NAND3X1 NAND3X1_153 ( .A(_abc_40319_new_n2854_), .B(_abc_40319_new_n2910_), .C(_abc_40319_new_n2882_), .Y(_abc_40319_new_n2911_));
NAND3X1 NAND3X1_154 ( .A(_abc_40319_new_n2908_), .B(_abc_40319_new_n2909_), .C(_abc_40319_new_n2912_), .Y(_abc_40319_new_n2913_));
NAND3X1 NAND3X1_155 ( .A(_abc_40319_new_n2863_), .B(_abc_40319_new_n2885_), .C(_abc_40319_new_n2888_), .Y(_abc_40319_new_n2921_));
NAND3X1 NAND3X1_156 ( .A(_abc_40319_new_n2927_), .B(_abc_40319_new_n2928_), .C(_abc_40319_new_n2925_), .Y(n982));
NAND3X1 NAND3X1_157 ( .A(_abc_40319_new_n2910_), .B(_abc_40319_new_n2909_), .C(_abc_40319_new_n2905_), .Y(_abc_40319_new_n2933_));
NAND3X1 NAND3X1_158 ( .A(_abc_40319_new_n2908_), .B(_abc_40319_new_n2932_), .C(_abc_40319_new_n2933_), .Y(_abc_40319_new_n2934_));
NAND3X1 NAND3X1_159 ( .A(_abc_40319_new_n2902_), .B(_abc_40319_new_n2908_), .C(_abc_40319_new_n2911_), .Y(_abc_40319_new_n2936_));
NAND3X1 NAND3X1_16 ( .A(_abc_40319_new_n632_), .B(_abc_40319_new_n633_), .C(_abc_40319_new_n634_), .Y(_abc_40319_new_n635_));
NAND3X1 NAND3X1_160 ( .A(_abc_40319_new_n2909_), .B(_abc_40319_new_n2935_), .C(_abc_40319_new_n2936_), .Y(_abc_40319_new_n2937_));
NAND3X1 NAND3X1_161 ( .A(_abc_40319_new_n2953_), .B(_abc_40319_new_n2948_), .C(_abc_40319_new_n2950_), .Y(n978));
NAND3X1 NAND3X1_162 ( .A(_abc_40319_new_n1370_), .B(_abc_40319_new_n1541_), .C(_abc_40319_new_n2969_), .Y(_abc_40319_new_n2970_));
NAND3X1 NAND3X1_163 ( .A(_abc_40319_new_n1865_), .B(_abc_40319_new_n1261_), .C(_abc_40319_new_n2971_), .Y(_abc_40319_new_n2972_));
NAND3X1 NAND3X1_164 ( .A(_abc_40319_new_n1159_), .B(_abc_40319_new_n1570_), .C(_abc_40319_new_n2973_), .Y(_abc_40319_new_n2974_));
NAND3X1 NAND3X1_165 ( .A(_abc_40319_new_n1108_), .B(_abc_40319_new_n1122_), .C(_abc_40319_new_n2975_), .Y(_abc_40319_new_n2976_));
NAND3X1 NAND3X1_166 ( .A(_abc_40319_new_n1017_), .B(_abc_40319_new_n1054_), .C(_abc_40319_new_n2977_), .Y(_abc_40319_new_n2978_));
NAND3X1 NAND3X1_167 ( .A(_abc_40319_new_n2088_), .B(_abc_40319_new_n2096_), .C(_abc_40319_new_n2979_), .Y(_abc_40319_new_n2980_));
NAND3X1 NAND3X1_168 ( .A(_abc_40319_new_n1877_), .B(_abc_40319_new_n2096_), .C(_abc_40319_new_n2982_), .Y(_abc_40319_new_n2983_));
NAND3X1 NAND3X1_169 ( .A(_abc_40319_new_n3044_), .B(_abc_40319_new_n3041_), .C(_abc_40319_new_n3039_), .Y(_abc_40319_new_n3045_));
NAND3X1 NAND3X1_17 ( .A(_abc_40319_new_n636_), .B(_abc_40319_new_n637_), .C(_abc_40319_new_n638_), .Y(_abc_40319_new_n639_));
NAND3X1 NAND3X1_170 ( .A(_abc_40319_new_n3007_), .B(_abc_40319_new_n3076_), .C(_abc_40319_new_n3027_), .Y(_abc_40319_new_n3077_));
NAND3X1 NAND3X1_171 ( .A(_abc_40319_new_n3101_), .B(_abc_40319_new_n3095_), .C(_abc_40319_new_n3097_), .Y(_abc_40319_new_n3102_));
NAND3X1 NAND3X1_172 ( .A(_abc_40319_new_n3107_), .B(_abc_40319_new_n3117_), .C(_abc_40319_new_n3116_), .Y(n958));
NAND3X1 NAND3X1_173 ( .A(_abc_40319_new_n3134_), .B(_abc_40319_new_n3139_), .C(_abc_40319_new_n3137_), .Y(_abc_40319_new_n3140_));
NAND3X1 NAND3X1_174 ( .A(_abc_40319_new_n3132_), .B(_abc_40319_new_n3142_), .C(_abc_40319_new_n3141_), .Y(n953));
NAND3X1 NAND3X1_175 ( .A(_abc_40319_new_n3148_), .B(_abc_40319_new_n3078_), .C(_abc_40319_new_n3077_), .Y(_abc_40319_new_n3149_));
NAND3X1 NAND3X1_176 ( .A(_abc_40319_new_n3087_), .B(_abc_40319_new_n3146_), .C(_abc_40319_new_n3149_), .Y(_abc_40319_new_n3150_));
NAND3X1 NAND3X1_177 ( .A(_abc_40319_new_n3144_), .B(_abc_40319_new_n3145_), .C(_abc_40319_new_n3150_), .Y(_abc_40319_new_n3151_));
NAND3X1 NAND3X1_178 ( .A(_abc_40319_new_n2353_), .B(_abc_40319_new_n2460_), .C(_abc_40319_new_n2138_), .Y(_abc_40319_new_n3235_));
NAND3X1 NAND3X1_179 ( .A(nRESET_G), .B(_abc_40319_new_n3227_), .C(_abc_40319_new_n3243_), .Y(_abc_40319_new_n3244_));
NAND3X1 NAND3X1_18 ( .A(_abc_40319_new_n644_), .B(_abc_40319_new_n645_), .C(_abc_40319_new_n646_), .Y(_abc_40319_new_n647_));
NAND3X1 NAND3X1_180 ( .A(nRESET_G), .B(_abc_40319_new_n3252_), .C(_abc_40319_new_n3262_), .Y(_abc_40319_new_n3263_));
NAND3X1 NAND3X1_181 ( .A(_abc_40319_new_n3275_), .B(_abc_40319_new_n3284_), .C(_abc_40319_new_n3274_), .Y(n923));
NAND3X1 NAND3X1_182 ( .A(_abc_40319_new_n3289_), .B(_abc_40319_new_n3293_), .C(_abc_40319_new_n3288_), .Y(_abc_40319_new_n3294_));
NAND3X1 NAND3X1_183 ( .A(_abc_40319_new_n3301_), .B(_abc_40319_new_n3304_), .C(_abc_40319_new_n3297_), .Y(_abc_40319_new_n3305_));
NAND3X1 NAND3X1_184 ( .A(_abc_40319_new_n3295_), .B(_abc_40319_new_n3296_), .C(_abc_40319_new_n3306_), .Y(n918));
NAND3X1 NAND3X1_185 ( .A(_abc_40319_new_n3314_), .B(_abc_40319_new_n3322_), .C(_abc_40319_new_n3313_), .Y(n913));
NAND3X1 NAND3X1_186 ( .A(_abc_40319_new_n1739_), .B(_abc_40319_new_n1309_), .C(_abc_40319_new_n3347_), .Y(_abc_40319_new_n3348_));
NAND3X1 NAND3X1_187 ( .A(_abc_40319_new_n3365_), .B(_abc_40319_new_n3374_), .C(_abc_40319_new_n3364_), .Y(n903));
NAND3X1 NAND3X1_188 ( .A(nRESET_G), .B(_abc_40319_new_n3376_), .C(_abc_40319_new_n3392_), .Y(n898));
NAND3X1 NAND3X1_189 ( .A(nRESET_G), .B(_abc_40319_new_n3394_), .C(_abc_40319_new_n3406_), .Y(n893));
NAND3X1 NAND3X1_19 ( .A(_abc_40319_new_n648_), .B(_abc_40319_new_n649_), .C(_abc_40319_new_n650_), .Y(_abc_40319_new_n651_));
NAND3X1 NAND3X1_190 ( .A(_abc_40319_new_n3441_), .B(_abc_40319_new_n3442_), .C(_abc_40319_new_n3437_), .Y(_abc_40319_new_n3443_));
NAND3X1 NAND3X1_191 ( .A(nRESET_G), .B(_abc_40319_new_n3447_), .C(_abc_40319_new_n3457_), .Y(n878));
NAND3X1 NAND3X1_192 ( .A(nRESET_G), .B(_abc_40319_new_n3462_), .C(_abc_40319_new_n3474_), .Y(n873));
NAND3X1 NAND3X1_193 ( .A(_abc_40319_new_n3488_), .B(_abc_40319_new_n3492_), .C(_abc_40319_new_n3486_), .Y(_abc_40319_new_n3493_));
NAND3X1 NAND3X1_194 ( .A(_abc_40319_new_n3522_), .B(_abc_40319_new_n3524_), .C(_abc_40319_new_n3519_), .Y(_abc_40319_new_n3525_));
NAND3X1 NAND3X1_195 ( .A(_abc_40319_new_n3541_), .B(_abc_40319_new_n3542_), .C(_abc_40319_new_n3538_), .Y(_abc_40319_new_n3543_));
NAND3X1 NAND3X1_196 ( .A(_abc_40319_new_n3559_), .B(_abc_40319_new_n3555_), .C(_abc_40319_new_n3558_), .Y(_abc_40319_new_n3560_));
NAND3X1 NAND3X1_197 ( .A(_abc_40319_new_n706_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n704_), .Y(_abc_40319_new_n3719_));
NAND3X1 NAND3X1_198 ( .A(nRESET_G), .B(_abc_40319_new_n3721_), .C(_abc_40319_new_n3719_), .Y(n328));
NAND3X1 NAND3X1_199 ( .A(_abc_40319_new_n591_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n587_), .Y(_abc_40319_new_n3731_));
NAND3X1 NAND3X1_2 ( .A(_abc_40319_new_n529_), .B(_abc_40319_new_n528_), .C(_abc_40319_new_n530_), .Y(_abc_40319_new_n531_));
NAND3X1 NAND3X1_20 ( .A(_abc_40319_new_n643_), .B(_abc_40319_new_n640_), .C(_abc_40319_new_n652_), .Y(_abc_40319_new_n653_));
NAND3X1 NAND3X1_200 ( .A(nRESET_G), .B(_abc_40319_new_n3732_), .C(_abc_40319_new_n3731_), .Y(n313));
NAND3X1 NAND3X1_201 ( .A(nRESET_G), .B(_abc_40319_new_n3761_), .C(_abc_40319_new_n3760_), .Y(n273));
NAND3X1 NAND3X1_202 ( .A(nRESET_G), .B(_abc_40319_new_n3767_), .C(_abc_40319_new_n3766_), .Y(n263));
NAND3X1 NAND3X1_203 ( .A(nRESET_G), .B(_abc_40319_new_n3774_), .C(_abc_40319_new_n3773_), .Y(n253));
NAND3X1 NAND3X1_204 ( .A(nRESET_G), .B(_abc_40319_new_n3780_), .C(_abc_40319_new_n3779_), .Y(n243));
NAND3X1 NAND3X1_205 ( .A(nRESET_G), .B(_abc_40319_new_n3788_), .C(_abc_40319_new_n3787_), .Y(n233));
NAND3X1 NAND3X1_206 ( .A(nRESET_G), .B(_abc_40319_new_n3791_), .C(_abc_40319_new_n3790_), .Y(n228));
NAND3X1 NAND3X1_207 ( .A(nRESET_G), .B(_abc_40319_new_n3806_), .C(_abc_40319_new_n3805_), .Y(n203));
NAND3X1 NAND3X1_208 ( .A(_abc_40319_new_n3815_), .B(_abc_40319_new_n3653_), .C(_abc_40319_new_n546_), .Y(_abc_40319_new_n3816_));
NAND3X1 NAND3X1_209 ( .A(nRESET_G), .B(_abc_40319_new_n3817_), .C(_abc_40319_new_n3816_), .Y(n188));
NAND3X1 NAND3X1_21 ( .A(_abc_40319_new_n684_), .B(_abc_40319_new_n685_), .C(_abc_40319_new_n550_), .Y(_abc_40319_new_n686_));
NAND3X1 NAND3X1_210 ( .A(_abc_40319_new_n608_), .B(_abc_40319_new_n667_), .C(_abc_40319_new_n663_), .Y(_abc_40319_new_n3823_));
NAND3X1 NAND3X1_211 ( .A(_abc_40319_new_n3838_), .B(_abc_40319_new_n2267_), .C(_abc_40319_new_n3840_), .Y(_abc_40319_new_n3841_));
NAND3X1 NAND3X1_212 ( .A(REG3_REG_14_), .B(REG3_REG_15_), .C(_abc_40319_new_n3859_), .Y(_abc_40319_new_n3860_));
NAND3X1 NAND3X1_213 ( .A(REG3_REG_19_), .B(REG3_REG_20_), .C(_abc_40319_new_n3863_), .Y(_abc_40319_new_n3864_));
NAND3X1 NAND3X1_214 ( .A(REG3_REG_24_), .B(REG3_REG_23_), .C(_abc_40319_new_n3866_), .Y(_abc_40319_new_n3867_));
NAND3X1 NAND3X1_215 ( .A(REG3_REG_27_), .B(REG3_REG_28_), .C(_abc_40319_new_n3869_), .Y(_abc_40319_new_n3870_));
NAND3X1 NAND3X1_216 ( .A(_abc_40319_new_n3854_), .B(_abc_40319_new_n3875_), .C(_abc_40319_new_n3853_), .Y(n963));
NAND3X1 NAND3X1_217 ( .A(_abc_40319_new_n654_), .B(_abc_40319_new_n3885_), .C(_abc_40319_new_n630_), .Y(_abc_40319_new_n3886_));
NAND3X1 NAND3X1_218 ( .A(_abc_40319_new_n3623_), .B(_abc_40319_new_n3910_), .C(_abc_40319_new_n3619_), .Y(_abc_40319_new_n3911_));
NAND3X1 NAND3X1_219 ( .A(_abc_40319_new_n3573_), .B(_abc_40319_new_n3920_), .C(_abc_40319_new_n3921_), .Y(_abc_40319_new_n3922_));
NAND3X1 NAND3X1_22 ( .A(IR_REG_31_), .B(_abc_40319_new_n591_), .C(_abc_40319_new_n587_), .Y(_abc_40319_new_n692_));
NAND3X1 NAND3X1_220 ( .A(_abc_40319_new_n3925_), .B(_abc_40319_new_n3926_), .C(_abc_40319_new_n3585_), .Y(_abc_40319_new_n3927_));
NAND3X1 NAND3X1_221 ( .A(_abc_40319_new_n3931_), .B(_abc_40319_new_n3932_), .C(_abc_40319_new_n3552_), .Y(_abc_40319_new_n3933_));
NAND3X1 NAND3X1_222 ( .A(_abc_40319_new_n3944_), .B(_abc_40319_new_n3945_), .C(_abc_40319_new_n3517_), .Y(_abc_40319_new_n3946_));
NAND3X1 NAND3X1_223 ( .A(_abc_40319_new_n3955_), .B(_abc_40319_new_n3956_), .C(_abc_40319_new_n3484_), .Y(_abc_40319_new_n3957_));
NAND3X1 NAND3X1_224 ( .A(_abc_40319_new_n3967_), .B(_abc_40319_new_n3968_), .C(_abc_40319_new_n3455_), .Y(_abc_40319_new_n3969_));
NAND3X1 NAND3X1_225 ( .A(_abc_40319_new_n3972_), .B(_abc_40319_new_n3973_), .C(_abc_40319_new_n3434_), .Y(_abc_40319_new_n3974_));
NAND3X1 NAND3X1_226 ( .A(_abc_40319_new_n3418_), .B(_abc_40319_new_n3977_), .C(_abc_40319_new_n3978_), .Y(_abc_40319_new_n3979_));
NAND3X1 NAND3X1_227 ( .A(nRESET_G), .B(_abc_40319_new_n3992_), .C(_abc_40319_new_n3991_), .Y(n578));
NAND3X1 NAND3X1_228 ( .A(_abc_40319_new_n3996_), .B(_abc_40319_new_n3997_), .C(_abc_40319_new_n3994_), .Y(_abc_40319_new_n3998_));
NAND3X1 NAND3X1_229 ( .A(_abc_40319_new_n4001_), .B(_abc_40319_new_n4002_), .C(_abc_40319_new_n3329_), .Y(_abc_40319_new_n4003_));
NAND3X1 NAND3X1_23 ( .A(_abc_40319_new_n543_), .B(_abc_40319_new_n701_), .C(_abc_40319_new_n700_), .Y(_abc_40319_new_n702_));
NAND3X1 NAND3X1_230 ( .A(nRESET_G), .B(_abc_40319_new_n4011_), .C(_abc_40319_new_n4010_), .Y(n593));
NAND3X1 NAND3X1_231 ( .A(nRESET_G), .B(_abc_40319_new_n4018_), .C(_abc_40319_new_n4017_), .Y(n603));
NAND3X1 NAND3X1_232 ( .A(_abc_40319_new_n4020_), .B(_abc_40319_new_n3260_), .C(_abc_40319_new_n4023_), .Y(_abc_40319_new_n4024_));
NAND3X1 NAND3X1_233 ( .A(_abc_40319_new_n4028_), .B(_abc_40319_new_n4029_), .C(_abc_40319_new_n3240_), .Y(_abc_40319_new_n4030_));
NAND3X1 NAND3X1_234 ( .A(_abc_40319_new_n4034_), .B(_abc_40319_new_n4035_), .C(_abc_40319_new_n3209_), .Y(_abc_40319_new_n4036_));
NAND3X1 NAND3X1_235 ( .A(_abc_40319_new_n4040_), .B(_abc_40319_new_n4041_), .C(_abc_40319_new_n3188_), .Y(_abc_40319_new_n4042_));
NAND3X1 NAND3X1_236 ( .A(_abc_40319_new_n4047_), .B(_abc_40319_new_n3158_), .C(_abc_40319_new_n4046_), .Y(_abc_40319_new_n4048_));
NAND3X1 NAND3X1_237 ( .A(_abc_40319_new_n3131_), .B(_abc_40319_new_n4052_), .C(_abc_40319_new_n4056_), .Y(_abc_40319_new_n4057_));
NAND3X1 NAND3X1_238 ( .A(_abc_40319_new_n4063_), .B(_abc_40319_new_n3106_), .C(_abc_40319_new_n4061_), .Y(_abc_40319_new_n4064_));
NAND3X1 NAND3X1_239 ( .A(_abc_40319_new_n3620_), .B(_abc_40319_new_n3856_), .C(_abc_40319_new_n3855_), .Y(_abc_40319_new_n4070_));
NAND3X1 NAND3X1_24 ( .A(_abc_40319_new_n699_), .B(_abc_40319_new_n590_), .C(_abc_40319_new_n703_), .Y(_abc_40319_new_n704_));
NAND3X1 NAND3X1_240 ( .A(_abc_40319_new_n3837_), .B(_abc_40319_new_n4070_), .C(_abc_40319_new_n3851_), .Y(_abc_40319_new_n4071_));
NAND3X1 NAND3X1_25 ( .A(IR_REG_31_), .B(_abc_40319_new_n706_), .C(_abc_40319_new_n704_), .Y(_abc_40319_new_n707_));
NAND3X1 NAND3X1_26 ( .A(_abc_40319_new_n532_), .B(_abc_40319_new_n590_), .C(_abc_40319_new_n710_), .Y(_abc_40319_new_n711_));
NAND3X1 NAND3X1_27 ( .A(IR_REG_31_), .B(_abc_40319_new_n711_), .C(_abc_40319_new_n720_), .Y(_abc_40319_new_n721_));
NAND3X1 NAND3X1_28 ( .A(_abc_40319_new_n682_), .B(_abc_40319_new_n660_), .C(_abc_40319_new_n743_), .Y(_abc_40319_new_n744_));
NAND3X1 NAND3X1_29 ( .A(_abc_40319_new_n755_), .B(_abc_40319_new_n752_), .C(_abc_40319_new_n745_), .Y(_abc_40319_new_n756_));
NAND3X1 NAND3X1_3 ( .A(_abc_40319_new_n533_), .B(_abc_40319_new_n534_), .C(_abc_40319_new_n535_), .Y(_abc_40319_new_n536_));
NAND3X1 NAND3X1_30 ( .A(_abc_40319_new_n716_), .B(_abc_40319_new_n719_), .C(_abc_40319_new_n773_), .Y(_abc_40319_new_n774_));
NAND3X1 NAND3X1_31 ( .A(_abc_40319_new_n707_), .B(_abc_40319_new_n708_), .C(_abc_40319_new_n773_), .Y(_abc_40319_new_n777_));
NAND3X1 NAND3X1_32 ( .A(_abc_40319_new_n786_), .B(_abc_40319_new_n785_), .C(_abc_40319_new_n745_), .Y(_abc_40319_new_n787_));
NAND3X1 NAND3X1_33 ( .A(_abc_40319_new_n784_), .B(_abc_40319_new_n787_), .C(_abc_40319_new_n790_), .Y(_abc_40319_new_n793_));
NAND3X1 NAND3X1_34 ( .A(_abc_40319_new_n707_), .B(_abc_40319_new_n708_), .C(_abc_40319_new_n723_), .Y(_abc_40319_new_n802_));
NAND3X1 NAND3X1_35 ( .A(_abc_40319_new_n757_), .B(_abc_40319_new_n850_), .C(_abc_40319_new_n845_), .Y(_abc_40319_new_n851_));
NAND3X1 NAND3X1_36 ( .A(_abc_40319_new_n844_), .B(_abc_40319_new_n857_), .C(_abc_40319_new_n851_), .Y(_abc_40319_new_n858_));
NAND3X1 NAND3X1_37 ( .A(_abc_40319_new_n757_), .B(_abc_40319_new_n862_), .C(_abc_40319_new_n860_), .Y(_abc_40319_new_n863_));
NAND3X1 NAND3X1_38 ( .A(REG2_REG_1_), .B(_abc_40319_new_n773_), .C(_abc_40319_new_n886_), .Y(_abc_40319_new_n887_));
NAND3X1 NAND3X1_39 ( .A(_abc_40319_new_n757_), .B(_abc_40319_new_n890_), .C(_abc_40319_new_n882_), .Y(_abc_40319_new_n891_));
NAND3X1 NAND3X1_4 ( .A(_abc_40319_new_n537_), .B(_abc_40319_new_n538_), .C(_abc_40319_new_n539_), .Y(_abc_40319_new_n540_));
NAND3X1 NAND3X1_40 ( .A(_abc_40319_new_n902_), .B(_abc_40319_new_n899_), .C(_abc_40319_new_n891_), .Y(_abc_40319_new_n903_));
NAND3X1 NAND3X1_41 ( .A(_abc_40319_new_n757_), .B(_abc_40319_new_n915_), .C(_abc_40319_new_n918_), .Y(_abc_40319_new_n919_));
NAND3X1 NAND3X1_42 ( .A(_abc_40319_new_n927_), .B(_abc_40319_new_n926_), .C(_abc_40319_new_n928_), .Y(_abc_40319_new_n929_));
NAND3X1 NAND3X1_43 ( .A(_abc_40319_new_n919_), .B(_abc_40319_new_n925_), .C(_abc_40319_new_n929_), .Y(_abc_40319_new_n930_));
NAND3X1 NAND3X1_44 ( .A(_abc_40319_new_n917_), .B(_abc_40319_new_n903_), .C(_abc_40319_new_n930_), .Y(_abc_40319_new_n931_));
NAND3X1 NAND3X1_45 ( .A(_abc_40319_new_n901_), .B(_abc_40319_new_n931_), .C(_abc_40319_new_n933_), .Y(_abc_40319_new_n934_));
NAND3X1 NAND3X1_46 ( .A(_abc_40319_new_n817_), .B(_abc_40319_new_n934_), .C(_abc_40319_new_n870_), .Y(_abc_40319_new_n935_));
NAND3X1 NAND3X1_47 ( .A(_abc_40319_new_n793_), .B(_abc_40319_new_n816_), .C(_abc_40319_new_n935_), .Y(_abc_40319_new_n936_));
NAND3X1 NAND3X1_48 ( .A(_abc_40319_new_n957_), .B(_abc_40319_new_n956_), .C(_abc_40319_new_n745_), .Y(_abc_40319_new_n958_));
NAND3X1 NAND3X1_49 ( .A(_abc_40319_new_n955_), .B(_abc_40319_new_n958_), .C(_abc_40319_new_n961_), .Y(_abc_40319_new_n963_));
NAND3X1 NAND3X1_5 ( .A(_abc_40319_new_n523_), .B(_abc_40319_new_n541_), .C(_abc_40319_new_n532_), .Y(_abc_40319_new_n542_));
NAND3X1 NAND3X1_50 ( .A(_abc_40319_new_n741_), .B(_abc_40319_new_n756_), .C(_abc_40319_new_n761_), .Y(_abc_40319_new_n964_));
NAND3X1 NAND3X1_51 ( .A(REG3_REG_9_), .B(_abc_40319_new_n1025_), .C(_abc_40319_new_n982_), .Y(_abc_40319_new_n1026_));
NAND3X1 NAND3X1_52 ( .A(REG3_REG_14_), .B(REG3_REG_15_), .C(_abc_40319_new_n1028_), .Y(_abc_40319_new_n1029_));
NAND3X1 NAND3X1_53 ( .A(REG3_REG_21_), .B(REG3_REG_22_), .C(_abc_40319_new_n1034_), .Y(_abc_40319_new_n1035_));
NAND3X1 NAND3X1_54 ( .A(REG3_REG_25_), .B(REG3_REG_24_), .C(_abc_40319_new_n1036_), .Y(_abc_40319_new_n1037_));
NAND3X1 NAND3X1_55 ( .A(_abc_40319_new_n727_), .B(_abc_40319_new_n1059_), .C(_abc_40319_new_n1056_), .Y(_abc_40319_new_n1060_));
NAND3X1 NAND3X1_56 ( .A(_abc_40319_new_n727_), .B(_abc_40319_new_n1087_), .C(_abc_40319_new_n1058_), .Y(_abc_40319_new_n1088_));
NAND3X1 NAND3X1_57 ( .A(_abc_40319_new_n963_), .B(_abc_40319_new_n793_), .C(_abc_40319_new_n964_), .Y(_abc_40319_new_n1280_));
NAND3X1 NAND3X1_58 ( .A(_abc_40319_new_n816_), .B(_abc_40319_new_n1281_), .C(_abc_40319_new_n935_), .Y(_abc_40319_new_n1282_));
NAND3X1 NAND3X1_59 ( .A(_abc_40319_new_n963_), .B(_abc_40319_new_n964_), .C(_abc_40319_new_n791_), .Y(_abc_40319_new_n1285_));
NAND3X1 NAND3X1_6 ( .A(_abc_40319_new_n547_), .B(_abc_40319_new_n524_), .C(_abc_40319_new_n548_), .Y(_abc_40319_new_n549_));
NAND3X1 NAND3X1_60 ( .A(_abc_40319_new_n1284_), .B(_abc_40319_new_n1285_), .C(_abc_40319_new_n1286_), .Y(_abc_40319_new_n1287_));
NAND3X1 NAND3X1_61 ( .A(_abc_40319_new_n1312_), .B(_abc_40319_new_n1288_), .C(_abc_40319_new_n1282_), .Y(_abc_40319_new_n1314_));
NAND3X1 NAND3X1_62 ( .A(IR_REG_31_), .B(_abc_40319_new_n1342_), .C(_abc_40319_new_n1345_), .Y(_abc_40319_new_n1346_));
NAND3X1 NAND3X1_63 ( .A(_abc_40319_new_n1414_), .B(_abc_40319_new_n1416_), .C(_abc_40319_new_n1412_), .Y(_abc_40319_new_n1417_));
NAND3X1 NAND3X1_64 ( .A(_abc_40319_new_n1240_), .B(_abc_40319_new_n1265_), .C(_abc_40319_new_n1420_), .Y(_abc_40319_new_n1421_));
NAND3X1 NAND3X1_65 ( .A(_abc_40319_new_n1217_), .B(_abc_40319_new_n1238_), .C(_abc_40319_new_n1421_), .Y(_abc_40319_new_n1422_));
NAND3X1 NAND3X1_66 ( .A(_abc_40319_new_n1165_), .B(_abc_40319_new_n1426_), .C(_abc_40319_new_n1422_), .Y(_abc_40319_new_n1427_));
NAND3X1 NAND3X1_67 ( .A(_abc_40319_new_n1434_), .B(_abc_40319_new_n1435_), .C(_abc_40319_new_n1433_), .Y(_abc_40319_new_n1436_));
NAND3X1 NAND3X1_68 ( .A(_abc_40319_new_n1448_), .B(_abc_40319_new_n1450_), .C(_abc_40319_new_n1449_), .Y(_abc_40319_new_n1451_));
NAND3X1 NAND3X1_69 ( .A(_abc_40319_new_n1466_), .B(_abc_40319_new_n1467_), .C(_abc_40319_new_n1465_), .Y(_abc_40319_new_n1468_));
NAND3X1 NAND3X1_7 ( .A(_abc_40319_new_n528_), .B(_abc_40319_new_n551_), .C(_abc_40319_new_n550_), .Y(_abc_40319_new_n552_));
NAND3X1 NAND3X1_70 ( .A(_abc_40319_new_n1163_), .B(_abc_40319_new_n1478_), .C(_abc_40319_new_n1427_), .Y(_abc_40319_new_n1479_));
NAND3X1 NAND3X1_71 ( .A(_abc_40319_new_n1143_), .B(_abc_40319_new_n1486_), .C(_abc_40319_new_n1479_), .Y(_abc_40319_new_n1487_));
NAND3X1 NAND3X1_72 ( .A(_abc_40319_new_n1121_), .B(_abc_40319_new_n1141_), .C(_abc_40319_new_n1487_), .Y(_abc_40319_new_n1488_));
NAND3X1 NAND3X1_73 ( .A(_abc_40319_new_n1530_), .B(_abc_40319_new_n1534_), .C(_abc_40319_new_n1528_), .Y(n1316));
NAND3X1 NAND3X1_74 ( .A(REG3_REG_27_), .B(REG3_REG_28_), .C(_abc_40319_new_n1039_), .Y(_abc_40319_new_n1595_));
NAND3X1 NAND3X1_75 ( .A(_abc_40319_new_n1101_), .B(_abc_40319_new_n1120_), .C(_abc_40319_new_n1488_), .Y(_abc_40319_new_n1662_));
NAND3X1 NAND3X1_76 ( .A(_abc_40319_new_n1712_), .B(_abc_40319_new_n1717_), .C(_abc_40319_new_n1709_), .Y(n1251));
NAND3X1 NAND3X1_77 ( .A(_abc_40319_new_n1722_), .B(_abc_40319_new_n1725_), .C(_abc_40319_new_n1730_), .Y(n1246));
NAND3X1 NAND3X1_78 ( .A(_abc_40319_new_n1787_), .B(_abc_40319_new_n1791_), .C(_abc_40319_new_n1785_), .Y(n1221));
NAND3X1 NAND3X1_79 ( .A(_abc_40319_new_n1811_), .B(_abc_40319_new_n1808_), .C(_abc_40319_new_n1816_), .Y(n1211));
NAND3X1 NAND3X1_8 ( .A(_abc_40319_new_n543_), .B(_abc_40319_new_n556_), .C(_abc_40319_new_n553_), .Y(_abc_40319_new_n557_));
NAND3X1 NAND3X1_80 ( .A(_abc_40319_new_n1823_), .B(_abc_40319_new_n1828_), .C(_abc_40319_new_n1821_), .Y(n1206));
NAND3X1 NAND3X1_81 ( .A(_abc_40319_new_n1660_), .B(_abc_40319_new_n1489_), .C(_abc_40319_new_n1662_), .Y(_abc_40319_new_n1845_));
NAND3X1 NAND3X1_82 ( .A(_abc_40319_new_n1864_), .B(_abc_40319_new_n1868_), .C(_abc_40319_new_n1861_), .Y(n1191));
NAND3X1 NAND3X1_83 ( .A(_abc_40319_new_n580_), .B(_abc_40319_new_n608_), .C(_abc_40319_new_n992_), .Y(_abc_40319_new_n1888_));
NAND3X1 NAND3X1_84 ( .A(_abc_40319_new_n877_), .B(_abc_40319_new_n879_), .C(_abc_40319_new_n878_), .Y(_abc_40319_new_n1902_));
NAND3X1 NAND3X1_85 ( .A(_abc_40319_new_n1904_), .B(_abc_40319_new_n914_), .C(_abc_40319_new_n1903_), .Y(_abc_40319_new_n1905_));
NAND3X1 NAND3X1_86 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1898_), .C(_abc_40319_new_n1906_), .Y(_abc_40319_new_n1907_));
NAND3X1 NAND3X1_87 ( .A(_abc_40319_new_n1925_), .B(_abc_40319_new_n1926_), .C(_abc_40319_new_n1924_), .Y(_abc_40319_new_n1927_));
NAND3X1 NAND3X1_88 ( .A(_abc_40319_new_n1932_), .B(_abc_40319_new_n1933_), .C(_abc_40319_new_n1931_), .Y(_abc_40319_new_n1934_));
NAND3X1 NAND3X1_89 ( .A(_abc_40319_new_n1936_), .B(_abc_40319_new_n1937_), .C(_abc_40319_new_n1939_), .Y(_abc_40319_new_n1940_));
NAND3X1 NAND3X1_9 ( .A(IR_REG_31_), .B(_abc_40319_new_n542_), .C(_abc_40319_new_n558_), .Y(_abc_40319_new_n559_));
NAND3X1 NAND3X1_90 ( .A(_abc_40319_new_n1940_), .B(_abc_40319_new_n1935_), .C(_abc_40319_new_n1929_), .Y(_abc_40319_new_n1941_));
NAND3X1 NAND3X1_91 ( .A(_abc_40319_new_n1923_), .B(_abc_40319_new_n1942_), .C(_abc_40319_new_n1922_), .Y(_abc_40319_new_n1943_));
NAND3X1 NAND3X1_92 ( .A(_abc_40319_new_n1946_), .B(_abc_40319_new_n1944_), .C(_abc_40319_new_n1945_), .Y(_abc_40319_new_n1947_));
NAND3X1 NAND3X1_93 ( .A(_abc_40319_new_n1960_), .B(_abc_40319_new_n1961_), .C(_abc_40319_new_n1959_), .Y(_abc_40319_new_n1962_));
NAND3X1 NAND3X1_94 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1351_), .C(_abc_40319_new_n1349_), .Y(_abc_40319_new_n1981_));
NAND3X1 NAND3X1_95 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n1982_), .C(_abc_40319_new_n1981_), .Y(_abc_40319_new_n1983_));
NAND3X1 NAND3X1_96 ( .A(_abc_40319_new_n1972_), .B(_abc_40319_new_n1974_), .C(_abc_40319_new_n1991_), .Y(_abc_40319_new_n1992_));
NAND3X1 NAND3X1_97 ( .A(_abc_40319_new_n2027_), .B(_abc_40319_new_n2028_), .C(_abc_40319_new_n2029_), .Y(_abc_40319_new_n2030_));
NAND3X1 NAND3X1_98 ( .A(_abc_40319_new_n615_), .B(_abc_40319_new_n663_), .C(_abc_40319_new_n2114_), .Y(_abc_40319_new_n2115_));
NAND3X1 NAND3X1_99 ( .A(_abc_40319_new_n2147_), .B(_abc_40319_new_n2151_), .C(_abc_40319_new_n2159_), .Y(_abc_40319_new_n2160_));
NOR2X1 NOR2X1_1 ( .A(IR_REG_5_), .B(IR_REG_4_), .Y(_abc_40319_new_n525_));
NOR2X1 NOR2X1_10 ( .A(IR_REG_19_), .B(IR_REG_18_), .Y(_abc_40319_new_n554_));
NOR2X1 NOR2X1_100 ( .A(_abc_40319_new_n1307_), .B(_abc_40319_new_n1304_), .Y(_abc_40319_new_n1308_));
NOR2X1 NOR2X1_101 ( .A(IR_REG_10_), .B(_abc_40319_new_n1290_), .Y(_abc_40319_new_n1343_));
NOR2X1 NOR2X1_102 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n1378_), .Y(_abc_40319_new_n1379_));
NOR2X1 NOR2X1_103 ( .A(_abc_40319_new_n1400_), .B(_abc_40319_new_n1396_), .Y(_abc_40319_new_n1401_));
NOR2X1 NOR2X1_104 ( .A(_abc_40319_new_n1361_), .B(_abc_40319_new_n1363_), .Y(_abc_40319_new_n1413_));
NOR2X1 NOR2X1_105 ( .A(_abc_40319_new_n1337_), .B(_abc_40319_new_n1339_), .Y(_abc_40319_new_n1415_));
NOR2X1 NOR2X1_106 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n1214_), .Y(_abc_40319_new_n1425_));
NOR2X1 NOR2X1_107 ( .A(_abc_40319_new_n1430_), .B(_abc_40319_new_n802_), .Y(_abc_40319_new_n1431_));
NOR2X1 NOR2X1_108 ( .A(_abc_40319_new_n778_), .B(_abc_40319_new_n1446_), .Y(_abc_40319_new_n1447_));
NOR2X1 NOR2X1_109 ( .A(_abc_40319_new_n1454_), .B(_abc_40319_new_n1456_), .Y(_abc_40319_new_n1457_));
NOR2X1 NOR2X1_11 ( .A(IR_REG_24_), .B(IR_REG_25_), .Y(_abc_40319_new_n561_));
NOR2X1 NOR2X1_110 ( .A(_abc_40319_new_n778_), .B(_abc_40319_new_n1463_), .Y(_abc_40319_new_n1464_));
NOR2X1 NOR2X1_111 ( .A(_abc_40319_new_n1470_), .B(_abc_40319_new_n1473_), .Y(_abc_40319_new_n1481_));
NOR2X1 NOR2X1_112 ( .A(_abc_40319_new_n1483_), .B(_abc_40319_new_n1481_), .Y(_abc_40319_new_n1484_));
NOR2X1 NOR2X1_113 ( .A(_abc_40319_new_n1107_), .B(_abc_40319_new_n1492_), .Y(_abc_40319_new_n1493_));
NOR2X1 NOR2X1_114 ( .A(_abc_40319_new_n1504_), .B(_abc_40319_new_n1499_), .Y(_abc_40319_new_n1505_));
NOR2X1 NOR2X1_115 ( .A(_abc_40319_new_n1335_), .B(_abc_40319_new_n1332_), .Y(_abc_40319_new_n1514_));
NOR2X1 NOR2X1_116 ( .A(_abc_40319_new_n1514_), .B(_abc_40319_new_n979_), .Y(_abc_40319_new_n1515_));
NOR2X1 NOR2X1_117 ( .A(_abc_40319_new_n1516_), .B(_abc_40319_new_n989_), .Y(_abc_40319_new_n1517_));
NOR2X1 NOR2X1_118 ( .A(_abc_40319_new_n1110_), .B(_abc_40319_new_n1003_), .Y(_abc_40319_new_n1531_));
NOR2X1 NOR2X1_119 ( .A(_abc_40319_new_n1533_), .B(_abc_40319_new_n1531_), .Y(_abc_40319_new_n1534_));
NOR2X1 NOR2X1_12 ( .A(_abc_40319_new_n567_), .B(_abc_40319_new_n572_), .Y(_abc_40319_new_n573_));
NOR2X1 NOR2X1_120 ( .A(_abc_40319_new_n1404_), .B(_abc_40319_new_n1406_), .Y(_abc_40319_new_n1536_));
NOR2X1 NOR2X1_121 ( .A(_abc_40319_new_n1536_), .B(_abc_40319_new_n1409_), .Y(_abc_40319_new_n1537_));
NOR2X1 NOR2X1_122 ( .A(_abc_40319_new_n1156_), .B(_abc_40319_new_n979_), .Y(_abc_40319_new_n1566_));
NOR2X1 NOR2X1_123 ( .A(_abc_40319_new_n1567_), .B(_abc_40319_new_n989_), .Y(_abc_40319_new_n1568_));
NOR2X1 NOR2X1_124 ( .A(_abc_40319_new_n1050_), .B(_abc_40319_new_n1107_), .Y(_abc_40319_new_n1578_));
NOR2X1 NOR2X1_125 ( .A(_abc_40319_new_n1052_), .B(_abc_40319_new_n1586_), .Y(_abc_40319_new_n1587_));
NOR2X1 NOR2X1_126 ( .A(_abc_40319_new_n1050_), .B(_abc_40319_new_n1589_), .Y(_abc_40319_new_n1590_));
NOR2X1 NOR2X1_127 ( .A(_abc_40319_new_n1471_), .B(_abc_40319_new_n1474_), .Y(_abc_40319_new_n1632_));
NOR2X1 NOR2X1_128 ( .A(_abc_40319_new_n1481_), .B(_abc_40319_new_n1475_), .Y(_abc_40319_new_n1637_));
NOR2X1 NOR2X1_129 ( .A(_abc_40319_new_n1379_), .B(_abc_40319_new_n979_), .Y(_abc_40319_new_n1651_));
NOR2X1 NOR2X1_13 ( .A(_abc_40319_new_n580_), .B(_abc_40319_new_n574_), .Y(_abc_40319_new_n581_));
NOR2X1 NOR2X1_130 ( .A(_abc_40319_new_n1514_), .B(_abc_40319_new_n989_), .Y(_abc_40319_new_n1652_));
NOR2X1 NOR2X1_131 ( .A(_abc_40319_new_n1191_), .B(_abc_40319_new_n1193_), .Y(_abc_40319_new_n1675_));
NOR2X1 NOR2X1_132 ( .A(_abc_40319_new_n1675_), .B(_abc_40319_new_n1424_), .Y(_abc_40319_new_n1676_));
NOR2X1 NOR2X1_133 ( .A(_abc_40319_new_n1425_), .B(_abc_40319_new_n1216_), .Y(_abc_40319_new_n1694_));
NOR2X1 NOR2X1_134 ( .A(_abc_40319_new_n865_), .B(_abc_40319_new_n979_), .Y(_abc_40319_new_n1723_));
NOR2X1 NOR2X1_135 ( .A(_abc_40319_new_n788_), .B(_abc_40319_new_n989_), .Y(_abc_40319_new_n1724_));
NOR2X1 NOR2X1_136 ( .A(_abc_40319_new_n988_), .B(_abc_40319_new_n979_), .Y(_abc_40319_new_n1736_));
NOR2X1 NOR2X1_137 ( .A(_abc_40319_new_n1401_), .B(_abc_40319_new_n989_), .Y(_abc_40319_new_n1737_));
NOR2X1 NOR2X1_138 ( .A(_abc_40319_new_n1468_), .B(_abc_40319_new_n1464_), .Y(_abc_40319_new_n1760_));
NOR2X1 NOR2X1_139 ( .A(_abc_40319_new_n991_), .B(_abc_40319_new_n1774_), .Y(_abc_40319_new_n1775_));
NOR2X1 NOR2X1_14 ( .A(RESET_G), .B(_abc_40319_new_n583_), .Y(n1345));
NOR2X1 NOR2X1_140 ( .A(_abc_40319_new_n1775_), .B(_abc_40319_new_n1778_), .Y(_abc_40319_new_n1779_));
NOR2X1 NOR2X1_141 ( .A(_abc_40319_new_n1128_), .B(_abc_40319_new_n1003_), .Y(_abc_40319_new_n1788_));
NOR2X1 NOR2X1_142 ( .A(_abc_40319_new_n1790_), .B(_abc_40319_new_n1788_), .Y(_abc_40319_new_n1791_));
NOR2X1 NOR2X1_143 ( .A(_abc_40319_new_n1401_), .B(_abc_40319_new_n979_), .Y(_abc_40319_new_n1795_));
NOR2X1 NOR2X1_144 ( .A(_abc_40319_new_n1796_), .B(_abc_40319_new_n989_), .Y(_abc_40319_new_n1797_));
NOR2X1 NOR2X1_145 ( .A(_abc_40319_new_n844_), .B(_abc_40319_new_n1552_), .Y(_abc_40319_new_n1805_));
NOR2X1 NOR2X1_146 ( .A(_abc_40319_new_n859_), .B(_abc_40319_new_n1805_), .Y(_abc_40319_new_n1806_));
NOR2X1 NOR2X1_147 ( .A(_abc_40319_new_n897_), .B(_abc_40319_new_n979_), .Y(_abc_40319_new_n1809_));
NOR2X1 NOR2X1_148 ( .A(_abc_40319_new_n865_), .B(_abc_40319_new_n989_), .Y(_abc_40319_new_n1810_));
NOR2X1 NOR2X1_149 ( .A(_abc_40319_new_n962_), .B(_abc_40319_new_n1830_), .Y(_abc_40319_new_n1831_));
NOR2X1 NOR2X1_15 ( .A(STATE_REG), .B(RESET_G), .Y(n1336));
NOR2X1 NOR2X1_150 ( .A(_abc_40319_new_n788_), .B(_abc_40319_new_n979_), .Y(_abc_40319_new_n1834_));
NOR2X1 NOR2X1_151 ( .A(_abc_40319_new_n759_), .B(_abc_40319_new_n989_), .Y(_abc_40319_new_n1835_));
NOR2X1 NOR2X1_152 ( .A(_abc_40319_new_n1102_), .B(_abc_40319_new_n1083_), .Y(_abc_40319_new_n1843_));
NOR2X1 NOR2X1_153 ( .A(_abc_40319_new_n1258_), .B(_abc_40319_new_n979_), .Y(_abc_40319_new_n1862_));
NOR2X1 NOR2X1_154 ( .A(_abc_40319_new_n1700_), .B(_abc_40319_new_n989_), .Y(_abc_40319_new_n1863_));
NOR2X1 NOR2X1_155 ( .A(_abc_40319_new_n618_), .B(_abc_40319_new_n1870_), .Y(_abc_40319_new_n1871_));
NOR2X1 NOR2X1_156 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n663_), .Y(_abc_40319_new_n1873_));
NOR2X1 NOR2X1_157 ( .A(_abc_40319_new_n1878_), .B(_abc_40319_new_n1881_), .Y(_abc_40319_new_n1882_));
NOR2X1 NOR2X1_158 ( .A(_abc_40319_new_n1890_), .B(_abc_40319_new_n1891_), .Y(_abc_40319_new_n1892_));
NOR2X1 NOR2X1_159 ( .A(_abc_40319_new_n825_), .B(_abc_40319_new_n1873_), .Y(_abc_40319_new_n1910_));
NOR2X1 NOR2X1_16 ( .A(IR_REG_31_), .B(IR_REG_27_), .Y(_abc_40319_new_n586_));
NOR2X1 NOR2X1_160 ( .A(_abc_40319_new_n1910_), .B(_abc_40319_new_n1911_), .Y(_abc_40319_new_n1912_));
NOR2X1 NOR2X1_161 ( .A(_abc_40319_new_n1928_), .B(_abc_40319_new_n1927_), .Y(_abc_40319_new_n1955_));
NOR2X1 NOR2X1_162 ( .A(_abc_40319_new_n1966_), .B(_abc_40319_new_n1968_), .Y(_abc_40319_new_n1969_));
NOR2X1 NOR2X1_163 ( .A(_abc_40319_new_n1963_), .B(_abc_40319_new_n1962_), .Y(_abc_40319_new_n1971_));
NOR2X1 NOR2X1_164 ( .A(_abc_40319_new_n1873_), .B(_abc_40319_new_n1370_), .Y(_abc_40319_new_n1985_));
NOR2X1 NOR2X1_165 ( .A(_abc_40319_new_n1977_), .B(_abc_40319_new_n1976_), .Y(_abc_40319_new_n1996_));
NOR2X1 NOR2X1_166 ( .A(_abc_40319_new_n2000_), .B(_abc_40319_new_n1999_), .Y(_abc_40319_new_n2005_));
NOR2X1 NOR2X1_167 ( .A(_abc_40319_new_n2088_), .B(_abc_40319_new_n1873_), .Y(_abc_40319_new_n2089_));
NOR2X1 NOR2X1_168 ( .A(_abc_40319_new_n2089_), .B(_abc_40319_new_n2090_), .Y(_abc_40319_new_n2091_));
NOR2X1 NOR2X1_169 ( .A(_abc_40319_new_n2098_), .B(_abc_40319_new_n2101_), .Y(_abc_40319_new_n2102_));
NOR2X1 NOR2X1_17 ( .A(IR_REG_27_), .B(_abc_40319_new_n589_), .Y(_abc_40319_new_n590_));
NOR2X1 NOR2X1_170 ( .A(_abc_40319_new_n992_), .B(_abc_40319_new_n742_), .Y(_abc_40319_new_n2116_));
NOR2X1 NOR2X1_171 ( .A(_abc_40319_new_n1085_), .B(_abc_40319_new_n1093_), .Y(_abc_40319_new_n2133_));
NOR2X1 NOR2X1_172 ( .A(_abc_40319_new_n2133_), .B(_abc_40319_new_n2132_), .Y(_abc_40319_new_n2134_));
NOR2X1 NOR2X1_173 ( .A(_abc_40319_new_n1459_), .B(_abc_40319_new_n1469_), .Y(_abc_40319_new_n2142_));
NOR2X1 NOR2X1_174 ( .A(_abc_40319_new_n2141_), .B(_abc_40319_new_n2142_), .Y(_abc_40319_new_n2143_));
NOR2X1 NOR2X1_175 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n1883_), .Y(_abc_40319_new_n2144_));
NOR2X1 NOR2X1_176 ( .A(_abc_40319_new_n2146_), .B(_abc_40319_new_n2144_), .Y(_abc_40319_new_n2147_));
NOR2X1 NOR2X1_177 ( .A(_abc_40319_new_n2096_), .B(_abc_40319_new_n2103_), .Y(_abc_40319_new_n2148_));
NOR2X1 NOR2X1_178 ( .A(_abc_40319_new_n2150_), .B(_abc_40319_new_n2148_), .Y(_abc_40319_new_n2151_));
NOR2X1 NOR2X1_179 ( .A(_abc_40319_new_n825_), .B(_abc_40319_new_n832_), .Y(_abc_40319_new_n2152_));
NOR2X1 NOR2X1_18 ( .A(IR_REG_31_), .B(IR_REG_28_), .Y(_abc_40319_new_n593_));
NOR2X1 NOR2X1_180 ( .A(_abc_40319_new_n2155_), .B(_abc_40319_new_n2158_), .Y(_abc_40319_new_n2159_));
NOR2X1 NOR2X1_181 ( .A(_abc_40319_new_n1159_), .B(_abc_40319_new_n1157_), .Y(_abc_40319_new_n2162_));
NOR2X1 NOR2X1_182 ( .A(_abc_40319_new_n1570_), .B(_abc_40319_new_n1437_), .Y(_abc_40319_new_n2167_));
NOR2X1 NOR2X1_183 ( .A(_abc_40319_new_n2160_), .B(_abc_40319_new_n2171_), .Y(_abc_40319_new_n2172_));
NOR2X1 NOR2X1_184 ( .A(_abc_40319_new_n799_), .B(_abc_40319_new_n1556_), .Y(_abc_40319_new_n2173_));
NOR2X1 NOR2X1_185 ( .A(_abc_40319_new_n1370_), .B(_abc_40319_new_n1380_), .Y(_abc_40319_new_n2178_));
NOR2X1 NOR2X1_186 ( .A(_abc_40319_new_n2176_), .B(_abc_40319_new_n2180_), .Y(_abc_40319_new_n2181_));
NOR2X1 NOR2X1_187 ( .A(_abc_40319_new_n1297_), .B(_abc_40319_new_n1309_), .Y(_abc_40319_new_n2182_));
NOR2X1 NOR2X1_188 ( .A(_abc_40319_new_n2184_), .B(_abc_40319_new_n2182_), .Y(_abc_40319_new_n2185_));
NOR2X1 NOR2X1_189 ( .A(_abc_40319_new_n698_), .B(_abc_40319_new_n740_), .Y(_abc_40319_new_n2187_));
NOR2X1 NOR2X1_19 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n614_), .Y(_abc_40319_new_n615_));
NOR2X1 NOR2X1_190 ( .A(_abc_40319_new_n1276_), .B(_abc_40319_new_n987_), .Y(_abc_40319_new_n2194_));
NOR2X1 NOR2X1_191 ( .A(_abc_40319_new_n2194_), .B(_abc_40319_new_n2193_), .Y(_abc_40319_new_n2195_));
NOR2X1 NOR2X1_192 ( .A(_abc_40319_new_n2195_), .B(_abc_40319_new_n2199_), .Y(_abc_40319_new_n2200_));
NOR2X1 NOR2X1_193 ( .A(_abc_40319_new_n1360_), .B(_abc_40319_new_n1654_), .Y(_abc_40319_new_n2202_));
NOR2X1 NOR2X1_194 ( .A(_abc_40319_new_n1401_), .B(_abc_40319_new_n1541_), .Y(_abc_40319_new_n2207_));
NOR2X1 NOR2X1_195 ( .A(_abc_40319_new_n2207_), .B(_abc_40319_new_n2206_), .Y(_abc_40319_new_n2208_));
NOR2X1 NOR2X1_196 ( .A(_abc_40319_new_n2208_), .B(_abc_40319_new_n2204_), .Y(_abc_40319_new_n2209_));
NOR2X1 NOR2X1_197 ( .A(_abc_40319_new_n2191_), .B(_abc_40319_new_n2210_), .Y(_abc_40319_new_n2211_));
NOR2X1 NOR2X1_198 ( .A(_abc_40319_new_n1442_), .B(_abc_40319_new_n1452_), .Y(_abc_40319_new_n2219_));
NOR2X1 NOR2X1_199 ( .A(_abc_40319_new_n2218_), .B(_abc_40319_new_n2219_), .Y(_abc_40319_new_n2220_));
NOR2X1 NOR2X1_2 ( .A(IR_REG_13_), .B(IR_REG_6_), .Y(_abc_40319_new_n529_));
NOR2X1 NOR2X1_20 ( .A(_abc_40319_new_n618_), .B(_abc_40319_new_n619_), .Y(_abc_40319_new_n620_));
NOR2X1 NOR2X1_200 ( .A(_abc_40319_new_n1865_), .B(_abc_40319_new_n1233_), .Y(_abc_40319_new_n2222_));
NOR2X1 NOR2X1_201 ( .A(_abc_40319_new_n2225_), .B(_abc_40319_new_n2224_), .Y(_abc_40319_new_n2226_));
NOR2X1 NOR2X1_202 ( .A(_abc_40319_new_n1325_), .B(_abc_40319_new_n1336_), .Y(_abc_40319_new_n2227_));
NOR2X1 NOR2X1_203 ( .A(_abc_40319_new_n2228_), .B(_abc_40319_new_n1514_), .Y(_abc_40319_new_n2229_));
NOR2X1 NOR2X1_204 ( .A(_abc_40319_new_n2229_), .B(_abc_40319_new_n2227_), .Y(_abc_40319_new_n2230_));
NOR2X1 NOR2X1_205 ( .A(_abc_40319_new_n769_), .B(_abc_40319_new_n788_), .Y(_abc_40319_new_n2232_));
NOR2X1 NOR2X1_206 ( .A(_abc_40319_new_n2232_), .B(_abc_40319_new_n2234_), .Y(_abc_40319_new_n2235_));
NOR2X1 NOR2X1_207 ( .A(_abc_40319_new_n1248_), .B(_abc_40319_new_n1259_), .Y(_abc_40319_new_n2238_));
NOR2X1 NOR2X1_208 ( .A(_abc_40319_new_n2240_), .B(_abc_40319_new_n2238_), .Y(_abc_40319_new_n2241_));
NOR2X1 NOR2X1_209 ( .A(_abc_40319_new_n2237_), .B(_abc_40319_new_n2241_), .Y(_abc_40319_new_n2242_));
NOR2X1 NOR2X1_21 ( .A(_abc_40319_new_n622_), .B(_abc_40319_new_n624_), .Y(_abc_40319_new_n625_));
NOR2X1 NOR2X1_210 ( .A(_abc_40319_new_n2245_), .B(_abc_40319_new_n2249_), .Y(_abc_40319_new_n2250_));
NOR2X1 NOR2X1_211 ( .A(_abc_40319_new_n2251_), .B(_abc_40319_new_n2236_), .Y(_abc_40319_new_n2252_));
NOR2X1 NOR2X1_212 ( .A(_abc_40319_new_n2253_), .B(_abc_40319_new_n2212_), .Y(_abc_40319_new_n2254_));
NOR2X1 NOR2X1_213 ( .A(_abc_40319_new_n2125_), .B(_abc_40319_new_n2256_), .Y(_abc_40319_new_n2257_));
NOR2X1 NOR2X1_214 ( .A(_abc_40319_new_n2262_), .B(_abc_40319_new_n1598_), .Y(_abc_40319_new_n2263_));
NOR2X1 NOR2X1_215 ( .A(_abc_40319_new_n2088_), .B(_abc_40319_new_n2264_), .Y(_abc_40319_new_n2265_));
NOR2X1 NOR2X1_216 ( .A(_abc_40319_new_n2265_), .B(_abc_40319_new_n2263_), .Y(_abc_40319_new_n2266_));
NOR2X1 NOR2X1_217 ( .A(_abc_40319_new_n2261_), .B(_abc_40319_new_n2267_), .Y(_abc_40319_new_n2268_));
NOR2X1 NOR2X1_218 ( .A(_abc_40319_new_n1896_), .B(_abc_40319_new_n2272_), .Y(_abc_40319_new_n2273_));
NOR2X1 NOR2X1_219 ( .A(_abc_40319_new_n2144_), .B(_abc_40319_new_n2308_), .Y(_abc_40319_new_n2309_));
NOR2X1 NOR2X1_22 ( .A(_abc_40319_new_n626_), .B(_abc_40319_new_n625_), .Y(_abc_40319_new_n627_));
NOR2X1 NOR2X1_220 ( .A(_abc_40319_new_n1123_), .B(_abc_40319_new_n1137_), .Y(_abc_40319_new_n2312_));
NOR2X1 NOR2X1_221 ( .A(_abc_40319_new_n2319_), .B(_abc_40319_new_n2324_), .Y(_abc_40319_new_n2329_));
NOR2X1 NOR2X1_222 ( .A(_abc_40319_new_n2332_), .B(_abc_40319_new_n2330_), .Y(_abc_40319_new_n2333_));
NOR2X1 NOR2X1_223 ( .A(_abc_40319_new_n2328_), .B(_abc_40319_new_n2334_), .Y(_abc_40319_new_n2335_));
NOR2X1 NOR2X1_224 ( .A(_abc_40319_new_n2341_), .B(_abc_40319_new_n2337_), .Y(_abc_40319_new_n2342_));
NOR2X1 NOR2X1_225 ( .A(_abc_40319_new_n2346_), .B(_abc_40319_new_n2347_), .Y(_abc_40319_new_n2348_));
NOR2X1 NOR2X1_226 ( .A(_abc_40319_new_n2358_), .B(_abc_40319_new_n2173_), .Y(_abc_40319_new_n2359_));
NOR2X1 NOR2X1_227 ( .A(_abc_40319_new_n1902_), .B(_abc_40319_new_n2360_), .Y(_abc_40319_new_n2361_));
NOR2X1 NOR2X1_228 ( .A(_abc_40319_new_n1004_), .B(_abc_40319_new_n742_), .Y(_abc_40319_new_n2362_));
NOR2X1 NOR2X1_229 ( .A(_abc_40319_new_n2275_), .B(_abc_40319_new_n2356_), .Y(_abc_40319_new_n2364_));
NOR2X1 NOR2X1_23 ( .A(D_REG_12_), .B(D_REG_15_), .Y(_abc_40319_new_n632_));
NOR2X1 NOR2X1_230 ( .A(_abc_40319_new_n2365_), .B(_abc_40319_new_n2366_), .Y(_abc_40319_new_n2367_));
NOR2X1 NOR2X1_231 ( .A(_abc_40319_new_n1739_), .B(_abc_40319_new_n1309_), .Y(_abc_40319_new_n2369_));
NOR2X1 NOR2X1_232 ( .A(_abc_40319_new_n2374_), .B(_abc_40319_new_n2317_), .Y(_abc_40319_new_n2375_));
NOR2X1 NOR2X1_233 ( .A(_abc_40319_new_n2228_), .B(_abc_40319_new_n1336_), .Y(_abc_40319_new_n2377_));
NOR2X1 NOR2X1_234 ( .A(_abc_40319_new_n2196_), .B(_abc_40319_new_n1189_), .Y(_abc_40319_new_n2381_));
NOR2X1 NOR2X1_235 ( .A(_abc_40319_new_n1261_), .B(_abc_40319_new_n1259_), .Y(_abc_40319_new_n2384_));
NOR2X1 NOR2X1_236 ( .A(_abc_40319_new_n2386_), .B(_abc_40319_new_n2317_), .Y(_abc_40319_new_n2387_));
NOR2X1 NOR2X1_237 ( .A(_abc_40319_new_n2388_), .B(_abc_40319_new_n740_), .Y(_abc_40319_new_n2389_));
NOR2X1 NOR2X1_238 ( .A(_abc_40319_new_n2390_), .B(_abc_40319_new_n2339_), .Y(_abc_40319_new_n2391_));
NOR2X1 NOR2X1_239 ( .A(_abc_40319_new_n1541_), .B(_abc_40319_new_n1402_), .Y(_abc_40319_new_n2394_));
NOR2X1 NOR2X1_24 ( .A(D_REG_14_), .B(D_REG_17_), .Y(_abc_40319_new_n633_));
NOR2X1 NOR2X1_240 ( .A(_abc_40319_new_n2395_), .B(_abc_40319_new_n2355_), .Y(_abc_40319_new_n2396_));
NOR2X1 NOR2X1_241 ( .A(_abc_40319_new_n1122_), .B(_abc_40319_new_n1135_), .Y(_abc_40319_new_n2405_));
NOR2X1 NOR2X1_242 ( .A(_abc_40319_new_n2142_), .B(_abc_40319_new_n2405_), .Y(_abc_40319_new_n2406_));
NOR2X1 NOR2X1_243 ( .A(_abc_40319_new_n2175_), .B(_abc_40319_new_n2310_), .Y(_abc_40319_new_n2416_));
NOR2X1 NOR2X1_244 ( .A(_abc_40319_new_n2422_), .B(_abc_40319_new_n2421_), .Y(_abc_40319_new_n2423_));
NOR2X1 NOR2X1_245 ( .A(_abc_40319_new_n987_), .B(_abc_40319_new_n2427_), .Y(_abc_40319_new_n2428_));
NOR2X1 NOR2X1_246 ( .A(_abc_40319_new_n2429_), .B(_abc_40319_new_n2308_), .Y(_abc_40319_new_n2430_));
NOR2X1 NOR2X1_247 ( .A(_abc_40319_new_n2425_), .B(_abc_40319_new_n2431_), .Y(_abc_40319_new_n2432_));
NOR2X1 NOR2X1_248 ( .A(_abc_40319_new_n2433_), .B(_abc_40319_new_n2355_), .Y(_abc_40319_new_n2434_));
NOR2X1 NOR2X1_249 ( .A(_abc_40319_new_n663_), .B(_abc_40319_new_n2445_), .Y(_abc_40319_new_n2446_));
NOR2X1 NOR2X1_25 ( .A(D_REG_5_), .B(D_REG_13_), .Y(_abc_40319_new_n634_));
NOR2X1 NOR2X1_250 ( .A(_abc_40319_new_n667_), .B(_abc_40319_new_n743_), .Y(_abc_40319_new_n2450_));
NOR2X1 NOR2X1_251 ( .A(_abc_40319_new_n2465_), .B(_abc_40319_new_n2466_), .Y(_abc_40319_new_n2467_));
NOR2X1 NOR2X1_252 ( .A(_abc_40319_new_n2480_), .B(_abc_40319_new_n2328_), .Y(_abc_40319_new_n2481_));
NOR2X1 NOR2X1_253 ( .A(_abc_40319_new_n2179_), .B(_abc_40319_new_n2328_), .Y(_abc_40319_new_n2483_));
NOR2X1 NOR2X1_254 ( .A(_abc_40319_new_n2222_), .B(_abc_40319_new_n2381_), .Y(_abc_40319_new_n2485_));
NOR2X1 NOR2X1_255 ( .A(_abc_40319_new_n2483_), .B(_abc_40319_new_n2488_), .Y(_abc_40319_new_n2489_));
NOR2X1 NOR2X1_256 ( .A(_abc_40319_new_n2496_), .B(_abc_40319_new_n2491_), .Y(_abc_40319_new_n2497_));
NOR2X1 NOR2X1_257 ( .A(_abc_40319_new_n2167_), .B(_abc_40319_new_n2219_), .Y(_abc_40319_new_n2500_));
NOR2X1 NOR2X1_258 ( .A(_abc_40319_new_n2499_), .B(_abc_40319_new_n2501_), .Y(_abc_40319_new_n2502_));
NOR2X1 NOR2X1_259 ( .A(_abc_40319_new_n2508_), .B(_abc_40319_new_n2506_), .Y(_abc_40319_new_n2509_));
NOR2X1 NOR2X1_26 ( .A(D_REG_19_), .B(D_REG_18_), .Y(_abc_40319_new_n636_));
NOR2X1 NOR2X1_260 ( .A(_abc_40319_new_n749_), .B(_abc_40319_new_n743_), .Y(_abc_40319_new_n2517_));
NOR2X1 NOR2X1_261 ( .A(_abc_40319_new_n977_), .B(_abc_40319_new_n2523_), .Y(_abc_40319_new_n2524_));
NOR2X1 NOR2X1_262 ( .A(IR_REG_0_), .B(REG1_REG_0_), .Y(_abc_40319_new_n2531_));
NOR2X1 NOR2X1_263 ( .A(_abc_40319_new_n871_), .B(_abc_40319_new_n909_), .Y(_abc_40319_new_n2532_));
NOR2X1 NOR2X1_264 ( .A(_abc_40319_new_n2531_), .B(_abc_40319_new_n2532_), .Y(_abc_40319_new_n2533_));
NOR2X1 NOR2X1_265 ( .A(_abc_40319_new_n581_), .B(n1341), .Y(_abc_40319_new_n2539_));
NOR2X1 NOR2X1_266 ( .A(_abc_40319_new_n1872_), .B(_abc_40319_new_n2539_), .Y(_abc_40319_new_n2542_));
NOR2X1 NOR2X1_267 ( .A(_abc_40319_new_n972_), .B(_abc_40319_new_n2539_), .Y(_abc_40319_new_n2543_));
NOR2X1 NOR2X1_268 ( .A(_abc_40319_new_n871_), .B(_abc_40319_new_n907_), .Y(_abc_40319_new_n2544_));
NOR2X1 NOR2X1_269 ( .A(REG2_REG_1_), .B(_abc_40319_new_n2544_), .Y(_abc_40319_new_n2545_));
NOR2X1 NOR2X1_27 ( .A(D_REG_21_), .B(D_REG_20_), .Y(_abc_40319_new_n637_));
NOR2X1 NOR2X1_270 ( .A(_abc_40319_new_n2545_), .B(_abc_40319_new_n2547_), .Y(_abc_40319_new_n2548_));
NOR2X1 NOR2X1_271 ( .A(_abc_40319_new_n2559_), .B(_abc_40319_new_n1749_), .Y(_abc_40319_new_n2560_));
NOR2X1 NOR2X1_272 ( .A(_abc_40319_new_n2565_), .B(_abc_40319_new_n2525_), .Y(_abc_40319_new_n2566_));
NOR2X1 NOR2X1_273 ( .A(REG1_REG_2_), .B(_abc_40319_new_n836_), .Y(_abc_40319_new_n2567_));
NOR2X1 NOR2X1_274 ( .A(REG1_REG_3_), .B(_abc_40319_new_n2581_), .Y(_abc_40319_new_n2582_));
NOR2X1 NOR2X1_275 ( .A(_abc_40319_new_n822_), .B(_abc_40319_new_n2586_), .Y(_abc_40319_new_n2587_));
NOR2X1 NOR2X1_276 ( .A(REG1_REG_5_), .B(_abc_40319_new_n2612_), .Y(_abc_40319_new_n2614_));
NOR2X1 NOR2X1_277 ( .A(_abc_40319_new_n2639_), .B(_abc_40319_new_n691_), .Y(_abc_40319_new_n2640_));
NOR2X1 NOR2X1_278 ( .A(_abc_40319_new_n2646_), .B(_abc_40319_new_n2648_), .Y(_abc_40319_new_n2649_));
NOR2X1 NOR2X1_279 ( .A(_abc_40319_new_n2655_), .B(_abc_40319_new_n2651_), .Y(_abc_40319_new_n2657_));
NOR2X1 NOR2X1_28 ( .A(D_REG_16_), .B(D_REG_22_), .Y(_abc_40319_new_n638_));
NOR2X1 NOR2X1_280 ( .A(_abc_40319_new_n2663_), .B(_abc_40319_new_n1274_), .Y(_abc_40319_new_n2664_));
NOR2X1 NOR2X1_281 ( .A(REG2_REG_8_), .B(_abc_40319_new_n1273_), .Y(_abc_40319_new_n2668_));
NOR2X1 NOR2X1_282 ( .A(_abc_40319_new_n2525_), .B(_abc_40319_new_n2670_), .Y(_abc_40319_new_n2671_));
NOR2X1 NOR2X1_283 ( .A(_abc_40319_new_n694_), .B(_abc_40319_new_n2686_), .Y(_abc_40319_new_n2687_));
NOR2X1 NOR2X1_284 ( .A(_abc_40319_new_n2525_), .B(_abc_40319_new_n2686_), .Y(_abc_40319_new_n2688_));
NOR2X1 NOR2X1_285 ( .A(_abc_40319_new_n1298_), .B(_abc_40319_new_n1295_), .Y(_abc_40319_new_n2700_));
NOR2X1 NOR2X1_286 ( .A(_abc_40319_new_n2712_), .B(_abc_40319_new_n2710_), .Y(_abc_40319_new_n2713_));
NOR2X1 NOR2X1_287 ( .A(REG2_REG_10_), .B(_abc_40319_new_n1390_), .Y(_abc_40319_new_n2725_));
NOR2X1 NOR2X1_288 ( .A(_abc_40319_new_n1372_), .B(_abc_40319_new_n2738_), .Y(_abc_40319_new_n2739_));
NOR2X1 NOR2X1_289 ( .A(REG1_REG_11_), .B(_abc_40319_new_n1369_), .Y(_abc_40319_new_n2741_));
NOR2X1 NOR2X1_29 ( .A(_abc_40319_new_n635_), .B(_abc_40319_new_n639_), .Y(_abc_40319_new_n640_));
NOR2X1 NOR2X1_290 ( .A(_abc_40319_new_n1373_), .B(_abc_40319_new_n2738_), .Y(_abc_40319_new_n2748_));
NOR2X1 NOR2X1_291 ( .A(REG2_REG_11_), .B(_abc_40319_new_n1369_), .Y(_abc_40319_new_n2750_));
NOR2X1 NOR2X1_292 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n2738_), .Y(_abc_40319_new_n2756_));
NOR2X1 NOR2X1_293 ( .A(REG1_REG_12_), .B(_abc_40319_new_n2761_), .Y(_abc_40319_new_n2763_));
NOR2X1 NOR2X1_294 ( .A(_abc_40319_new_n1354_), .B(_abc_40319_new_n1348_), .Y(_abc_40319_new_n2770_));
NOR2X1 NOR2X1_295 ( .A(REG2_REG_12_), .B(_abc_40319_new_n2761_), .Y(_abc_40319_new_n2771_));
NOR2X1 NOR2X1_296 ( .A(_abc_40319_new_n2770_), .B(_abc_40319_new_n2771_), .Y(_abc_40319_new_n2772_));
NOR2X1 NOR2X1_297 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n1348_), .Y(_abc_40319_new_n2778_));
NOR2X1 NOR2X1_298 ( .A(_abc_40319_new_n1333_), .B(_abc_40319_new_n1323_), .Y(_abc_40319_new_n2789_));
NOR2X1 NOR2X1_299 ( .A(REG2_REG_13_), .B(_abc_40319_new_n1322_), .Y(_abc_40319_new_n2790_));
NOR2X1 NOR2X1_3 ( .A(_abc_40319_new_n527_), .B(_abc_40319_new_n531_), .Y(_abc_40319_new_n532_));
NOR2X1 NOR2X1_30 ( .A(D_REG_24_), .B(D_REG_23_), .Y(_abc_40319_new_n641_));
NOR2X1 NOR2X1_300 ( .A(_abc_40319_new_n2790_), .B(_abc_40319_new_n2789_), .Y(_abc_40319_new_n2791_));
NOR2X1 NOR2X1_301 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n1323_), .Y(_abc_40319_new_n2797_));
NOR2X1 NOR2X1_302 ( .A(_abc_40319_new_n2808_), .B(_abc_40319_new_n2809_), .Y(_abc_40319_new_n2810_));
NOR2X1 NOR2X1_303 ( .A(_abc_40319_new_n2810_), .B(_abc_40319_new_n2807_), .Y(_abc_40319_new_n2811_));
NOR2X1 NOR2X1_304 ( .A(_abc_40319_new_n1249_), .B(_abc_40319_new_n1246_), .Y(_abc_40319_new_n2812_));
NOR2X1 NOR2X1_305 ( .A(REG2_REG_14_), .B(_abc_40319_new_n1245_), .Y(_abc_40319_new_n2813_));
NOR2X1 NOR2X1_306 ( .A(_abc_40319_new_n2813_), .B(_abc_40319_new_n2812_), .Y(_abc_40319_new_n2814_));
NOR2X1 NOR2X1_307 ( .A(_abc_40319_new_n1225_), .B(_abc_40319_new_n1221_), .Y(_abc_40319_new_n2834_));
NOR2X1 NOR2X1_308 ( .A(REG2_REG_15_), .B(_abc_40319_new_n2836_), .Y(_abc_40319_new_n2837_));
NOR2X1 NOR2X1_309 ( .A(_abc_40319_new_n1179_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2853_));
NOR2X1 NOR2X1_31 ( .A(D_REG_11_), .B(D_REG_10_), .Y(_abc_40319_new_n642_));
NOR2X1 NOR2X1_310 ( .A(REG1_REG_16_), .B(_abc_40319_new_n2855_), .Y(_abc_40319_new_n2856_));
NOR2X1 NOR2X1_311 ( .A(REG2_REG_16_), .B(_abc_40319_new_n2855_), .Y(_abc_40319_new_n2864_));
NOR2X1 NOR2X1_312 ( .A(_abc_40319_new_n1199_), .B(_abc_40319_new_n1196_), .Y(_abc_40319_new_n2878_));
NOR2X1 NOR2X1_313 ( .A(REG1_REG_17_), .B(_abc_40319_new_n2879_), .Y(_abc_40319_new_n2880_));
NOR2X1 NOR2X1_314 ( .A(_abc_40319_new_n2878_), .B(_abc_40319_new_n2880_), .Y(_abc_40319_new_n2881_));
NOR2X1 NOR2X1_315 ( .A(REG1_REG_18_), .B(_abc_40319_new_n2899_), .Y(_abc_40319_new_n2900_));
NOR2X1 NOR2X1_316 ( .A(_abc_40319_new_n1149_), .B(_abc_40319_new_n1146_), .Y(_abc_40319_new_n2901_));
NOR2X1 NOR2X1_317 ( .A(REG2_REG_18_), .B(_abc_40319_new_n2899_), .Y(_abc_40319_new_n2915_));
NOR2X1 NOR2X1_318 ( .A(_abc_40319_new_n2917_), .B(_abc_40319_new_n1146_), .Y(_abc_40319_new_n2918_));
NOR2X1 NOR2X1_319 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n1146_), .Y(_abc_40319_new_n2926_));
NOR2X1 NOR2X1_32 ( .A(D_REG_26_), .B(D_REG_25_), .Y(_abc_40319_new_n644_));
NOR2X1 NOR2X1_320 ( .A(_abc_40319_new_n1430_), .B(_abc_40319_new_n667_), .Y(_abc_40319_new_n2930_));
NOR2X1 NOR2X1_321 ( .A(REG1_REG_19_), .B(_abc_40319_new_n749_), .Y(_abc_40319_new_n2931_));
NOR2X1 NOR2X1_322 ( .A(_abc_40319_new_n2930_), .B(_abc_40319_new_n2931_), .Y(_abc_40319_new_n2932_));
NOR2X1 NOR2X1_323 ( .A(_abc_40319_new_n2942_), .B(_abc_40319_new_n2946_), .Y(_abc_40319_new_n2949_));
NOR2X1 NOR2X1_324 ( .A(_abc_40319_new_n660_), .B(_abc_40319_new_n973_), .Y(_abc_40319_new_n2955_));
NOR2X1 NOR2X1_325 ( .A(_abc_40319_new_n656_), .B(_abc_40319_new_n630_), .Y(_abc_40319_new_n2956_));
NOR2X1 NOR2X1_326 ( .A(_abc_40319_new_n972_), .B(_abc_40319_new_n2957_), .Y(_abc_40319_new_n2958_));
NOR2X1 NOR2X1_327 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n2962_), .Y(_abc_40319_new_n2963_));
NOR2X1 NOR2X1_328 ( .A(_abc_40319_new_n799_), .B(_abc_40319_new_n2964_), .Y(_abc_40319_new_n2965_));
NOR2X1 NOR2X1_329 ( .A(_abc_40319_new_n944_), .B(_abc_40319_new_n2966_), .Y(_abc_40319_new_n2967_));
NOR2X1 NOR2X1_33 ( .A(D_REG_2_), .B(D_REG_29_), .Y(_abc_40319_new_n645_));
NOR2X1 NOR2X1_330 ( .A(_abc_40319_new_n1582_), .B(_abc_40319_new_n2978_), .Y(_abc_40319_new_n2979_));
NOR2X1 NOR2X1_331 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n2991_));
NOR2X1 NOR2X1_332 ( .A(_abc_40319_new_n619_), .B(_abc_40319_new_n2993_), .Y(_abc_40319_new_n2994_));
NOR2X1 NOR2X1_333 ( .A(_abc_40319_new_n619_), .B(_abc_40319_new_n3000_), .Y(_abc_40319_new_n3001_));
NOR2X1 NOR2X1_334 ( .A(_abc_40319_new_n1108_), .B(_abc_40319_new_n1710_), .Y(_abc_40319_new_n3006_));
NOR2X1 NOR2X1_335 ( .A(_abc_40319_new_n1443_), .B(_abc_40319_new_n1452_), .Y(_abc_40319_new_n3009_));
NOR2X1 NOR2X1_336 ( .A(_abc_40319_new_n3008_), .B(_abc_40319_new_n3011_), .Y(_abc_40319_new_n3012_));
NOR2X1 NOR2X1_337 ( .A(_abc_40319_new_n1148_), .B(_abc_40319_new_n1157_), .Y(_abc_40319_new_n3017_));
NOR2X1 NOR2X1_338 ( .A(_abc_40319_new_n3017_), .B(_abc_40319_new_n3011_), .Y(_abc_40319_new_n3018_));
NOR2X1 NOR2X1_339 ( .A(_abc_40319_new_n1223_), .B(_abc_40319_new_n1233_), .Y(_abc_40319_new_n3028_));
NOR2X1 NOR2X1_34 ( .A(D_REG_28_), .B(D_REG_27_), .Y(_abc_40319_new_n646_));
NOR2X1 NOR2X1_340 ( .A(_abc_40319_new_n922_), .B(_abc_40319_new_n912_), .Y(_abc_40319_new_n3037_));
NOR2X1 NOR2X1_341 ( .A(_abc_40319_new_n769_), .B(_abc_40319_new_n783_), .Y(_abc_40319_new_n3040_));
NOR2X1 NOR2X1_342 ( .A(_abc_40319_new_n826_), .B(_abc_40319_new_n832_), .Y(_abc_40319_new_n3042_));
NOR2X1 NOR2X1_343 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n842_), .Y(_abc_40319_new_n3043_));
NOR2X1 NOR2X1_344 ( .A(_abc_40319_new_n3043_), .B(_abc_40319_new_n3042_), .Y(_abc_40319_new_n3044_));
NOR2X1 NOR2X1_345 ( .A(_abc_40319_new_n2184_), .B(_abc_40319_new_n2207_), .Y(_abc_40319_new_n3056_));
NOR2X1 NOR2X1_346 ( .A(_abc_40319_new_n3082_), .B(_abc_40319_new_n3080_), .Y(_abc_40319_new_n3083_));
NOR2X1 NOR2X1_347 ( .A(_abc_40319_new_n1017_), .B(_abc_40319_new_n1592_), .Y(_abc_40319_new_n3086_));
NOR2X1 NOR2X1_348 ( .A(_abc_40319_new_n1084_), .B(_abc_40319_new_n1093_), .Y(_abc_40319_new_n3090_));
NOR2X1 NOR2X1_349 ( .A(_abc_40319_new_n3094_), .B(_abc_40319_new_n3085_), .Y(_abc_40319_new_n3096_));
NOR2X1 NOR2X1_35 ( .A(D_REG_7_), .B(D_REG_4_), .Y(_abc_40319_new_n648_));
NOR2X1 NOR2X1_350 ( .A(_abc_40319_new_n977_), .B(_abc_40319_new_n616_), .Y(_abc_40319_new_n3103_));
NOR2X1 NOR2X1_351 ( .A(_abc_40319_new_n2985_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3108_));
NOR2X1 NOR2X1_352 ( .A(_abc_40319_new_n1085_), .B(_abc_40319_new_n2976_), .Y(_abc_40319_new_n3160_));
NOR2X1 NOR2X1_353 ( .A(_abc_40319_new_n3178_), .B(_abc_40319_new_n3181_), .Y(_abc_40319_new_n3182_));
NOR2X1 NOR2X1_354 ( .A(_abc_40319_new_n2354_), .B(_abc_40319_new_n3182_), .Y(_abc_40319_new_n3183_));
NOR2X1 NOR2X1_355 ( .A(_abc_40319_new_n2133_), .B(_abc_40319_new_n3183_), .Y(_abc_40319_new_n3184_));
NOR2X1 NOR2X1_356 ( .A(_abc_40319_new_n1070_), .B(_abc_40319_new_n3160_), .Y(_abc_40319_new_n3190_));
NOR2X1 NOR2X1_357 ( .A(_abc_40319_new_n2977_), .B(_abc_40319_new_n3190_), .Y(_abc_40319_new_n3191_));
NOR2X1 NOR2X1_358 ( .A(REG2_REG_25_), .B(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3193_));
NOR2X1 NOR2X1_359 ( .A(_abc_40319_new_n1070_), .B(_abc_40319_new_n994_), .Y(_abc_40319_new_n3194_));
NOR2X1 NOR2X1_36 ( .A(D_REG_3_), .B(D_REG_6_), .Y(_abc_40319_new_n649_));
NOR2X1 NOR2X1_360 ( .A(_abc_40319_new_n3194_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3195_));
NOR2X1 NOR2X1_361 ( .A(_abc_40319_new_n2499_), .B(_abc_40319_new_n3230_), .Y(_abc_40319_new_n3233_));
NOR2X1 NOR2X1_362 ( .A(REG2_REG_23_), .B(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3241_));
NOR2X1 NOR2X1_363 ( .A(_abc_40319_new_n1459_), .B(_abc_40319_new_n994_), .Y(_abc_40319_new_n3279_));
NOR2X1 NOR2X1_364 ( .A(_abc_40319_new_n1442_), .B(_abc_40319_new_n994_), .Y(_abc_40319_new_n3302_));
NOR2X1 NOR2X1_365 ( .A(_abc_40319_new_n1570_), .B(_abc_40319_new_n994_), .Y(_abc_40319_new_n3316_));
NOR2X1 NOR2X1_366 ( .A(_abc_40319_new_n1175_), .B(_abc_40319_new_n2972_), .Y(_abc_40319_new_n3331_));
NOR2X1 NOR2X1_367 ( .A(_abc_40319_new_n2394_), .B(_abc_40319_new_n2178_), .Y(_abc_40319_new_n3347_));
NOR2X1 NOR2X1_368 ( .A(_abc_40319_new_n1211_), .B(_abc_40319_new_n3331_), .Y(_abc_40319_new_n3366_));
NOR2X1 NOR2X1_369 ( .A(_abc_40319_new_n2973_), .B(_abc_40319_new_n3366_), .Y(_abc_40319_new_n3367_));
NOR2X1 NOR2X1_37 ( .A(D_REG_31_), .B(D_REG_8_), .Y(_abc_40319_new_n650_));
NOR2X1 NOR2X1_370 ( .A(_abc_40319_new_n3381_), .B(_abc_40319_new_n3391_), .Y(_abc_40319_new_n3392_));
NOR2X1 NOR2X1_371 ( .A(_abc_40319_new_n3397_), .B(_abc_40319_new_n3405_), .Y(_abc_40319_new_n3406_));
NOR2X1 NOR2X1_372 ( .A(_abc_40319_new_n1352_), .B(_abc_40319_new_n2970_), .Y(_abc_40319_new_n3414_));
NOR2X1 NOR2X1_373 ( .A(_abc_40319_new_n3418_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3419_));
NOR2X1 NOR2X1_374 ( .A(_abc_40319_new_n2228_), .B(_abc_40319_new_n3414_), .Y(_abc_40319_new_n3435_));
NOR2X1 NOR2X1_375 ( .A(_abc_40319_new_n2971_), .B(_abc_40319_new_n3435_), .Y(_abc_40319_new_n3436_));
NOR2X1 NOR2X1_376 ( .A(_abc_40319_new_n2228_), .B(_abc_40319_new_n994_), .Y(_abc_40319_new_n3438_));
NOR2X1 NOR2X1_377 ( .A(_abc_40319_new_n3438_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3439_));
NOR2X1 NOR2X1_378 ( .A(_abc_40319_new_n3451_), .B(_abc_40319_new_n3456_), .Y(_abc_40319_new_n3457_));
NOR2X1 NOR2X1_379 ( .A(_abc_40319_new_n3465_), .B(_abc_40319_new_n3473_), .Y(_abc_40319_new_n3474_));
NOR2X1 NOR2X1_38 ( .A(_abc_40319_new_n647_), .B(_abc_40319_new_n651_), .Y(_abc_40319_new_n652_));
NOR2X1 NOR2X1_380 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n1541_), .Y(_abc_40319_new_n3489_));
NOR2X1 NOR2X1_381 ( .A(_abc_40319_new_n2427_), .B(_abc_40319_new_n994_), .Y(_abc_40319_new_n3520_));
NOR2X1 NOR2X1_382 ( .A(_abc_40319_new_n1308_), .B(_abc_40319_new_n2985_), .Y(_abc_40319_new_n3521_));
NOR2X1 NOR2X1_383 ( .A(_abc_40319_new_n663_), .B(_abc_40319_new_n660_), .Y(_abc_40319_new_n3620_));
NOR2X1 NOR2X1_384 ( .A(_abc_40319_new_n912_), .B(_abc_40319_new_n3104_), .Y(_abc_40319_new_n3630_));
NOR2X1 NOR2X1_385 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n618_), .Y(_abc_40319_new_n3653_));
NOR2X1 NOR2X1_386 ( .A(IR_REG_31_), .B(_abc_40319_new_n618_), .Y(_abc_40319_new_n3720_));
NOR2X1 NOR2X1_387 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1170_), .Y(_abc_40319_new_n3770_));
NOR2X1 NOR2X1_388 ( .A(_abc_40319_new_n3825_), .B(_abc_40319_new_n3003_), .Y(_abc_40319_new_n3826_));
NOR2X1 NOR2X1_389 ( .A(_abc_40319_new_n1581_), .B(_abc_40319_new_n2267_), .Y(_abc_40319_new_n3828_));
NOR2X1 NOR2X1_39 ( .A(_abc_40319_new_n630_), .B(_abc_40319_new_n657_), .Y(_abc_40319_new_n658_));
NOR2X1 NOR2X1_390 ( .A(_abc_40319_new_n3827_), .B(_abc_40319_new_n3832_), .Y(_abc_40319_new_n3833_));
NOR2X1 NOR2X1_391 ( .A(_abc_40319_new_n1327_), .B(_abc_40319_new_n1026_), .Y(_abc_40319_new_n3858_));
NOR2X1 NOR2X1_392 ( .A(_abc_40319_new_n1184_), .B(_abc_40319_new_n3860_), .Y(_abc_40319_new_n3861_));
NOR2X1 NOR2X1_393 ( .A(_abc_40319_new_n1151_), .B(_abc_40319_new_n3862_), .Y(_abc_40319_new_n3863_));
NOR2X1 NOR2X1_394 ( .A(_abc_40319_new_n1124_), .B(_abc_40319_new_n3864_), .Y(_abc_40319_new_n3865_));
NOR2X1 NOR2X1_395 ( .A(_abc_40319_new_n1057_), .B(_abc_40319_new_n3867_), .Y(_abc_40319_new_n3868_));
NOR2X1 NOR2X1_396 ( .A(_abc_40319_new_n2088_), .B(_abc_40319_new_n994_), .Y(_abc_40319_new_n3871_));
NOR2X1 NOR2X1_397 ( .A(_abc_40319_new_n972_), .B(_abc_40319_new_n3886_), .Y(_abc_40319_new_n3887_));
NOR2X1 NOR2X1_398 ( .A(_abc_40319_new_n656_), .B(_abc_40319_new_n3888_), .Y(_abc_40319_new_n3889_));
NOR2X1 NOR2X1_399 ( .A(_abc_40319_new_n3891_), .B(_abc_40319_new_n3300_), .Y(_abc_40319_new_n3892_));
NOR2X1 NOR2X1_4 ( .A(IR_REG_15_), .B(IR_REG_14_), .Y(_abc_40319_new_n535_));
NOR2X1 NOR2X1_40 ( .A(_abc_40319_new_n667_), .B(_abc_40319_new_n663_), .Y(_abc_40319_new_n668_));
NOR2X1 NOR2X1_400 ( .A(_abc_40319_new_n3294_), .B(_abc_40319_new_n3896_), .Y(_abc_40319_new_n3897_));
NOR2X1 NOR2X1_401 ( .A(_abc_40319_new_n3345_), .B(_abc_40319_new_n3363_), .Y(_abc_40319_new_n3994_));
NOR2X1 NOR2X1_402 ( .A(_abc_40319_new_n1017_), .B(_abc_40319_new_n994_), .Y(_abc_40319_new_n4053_));
NOR2X1 NOR2X1_403 ( .A(_abc_40319_new_n2985_), .B(_abc_40319_new_n1505_), .Y(_abc_40319_new_n4055_));
NOR2X1 NOR2X1_404 ( .A(_abc_40319_new_n1005_), .B(_abc_40319_new_n3109_), .Y(_abc_40319_new_n4062_));
NOR2X1 NOR2X1_41 ( .A(_abc_40319_new_n580_), .B(_abc_40319_new_n671_), .Y(_abc_40319_new_n672_));
NOR2X1 NOR2X1_42 ( .A(_abc_40319_new_n618_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n674_));
NOR2X1 NOR2X1_43 ( .A(_abc_40319_new_n675_), .B(_abc_40319_new_n659_), .Y(_abc_40319_new_n676_));
NOR2X1 NOR2X1_44 ( .A(_abc_40319_new_n663_), .B(_abc_40319_new_n614_), .Y(_abc_40319_new_n678_));
NOR2X1 NOR2X1_45 ( .A(_abc_40319_new_n667_), .B(_abc_40319_new_n609_), .Y(_abc_40319_new_n680_));
NOR2X1 NOR2X1_46 ( .A(_abc_40319_new_n663_), .B(_abc_40319_new_n680_), .Y(_abc_40319_new_n681_));
NOR2X1 NOR2X1_47 ( .A(_abc_40319_new_n536_), .B(_abc_40319_new_n540_), .Y(_abc_40319_new_n700_));
NOR2X1 NOR2X1_48 ( .A(IR_REG_28_), .B(IR_REG_29_), .Y(_abc_40319_new_n701_));
NOR2X1 NOR2X1_49 ( .A(_abc_40319_new_n552_), .B(_abc_40319_new_n702_), .Y(_abc_40319_new_n703_));
NOR2X1 NOR2X1_5 ( .A(IR_REG_20_), .B(IR_REG_21_), .Y(_abc_40319_new_n538_));
NOR2X1 NOR2X1_50 ( .A(IR_REG_30_), .B(_abc_40319_new_n711_), .Y(_abc_40319_new_n717_));
NOR2X1 NOR2X1_51 ( .A(_abc_40319_new_n729_), .B(_abc_40319_new_n730_), .Y(_abc_40319_new_n731_));
NOR2X1 NOR2X1_52 ( .A(_abc_40319_new_n728_), .B(_abc_40319_new_n732_), .Y(_abc_40319_new_n733_));
NOR2X1 NOR2X1_53 ( .A(_abc_40319_new_n782_), .B(_abc_40319_new_n775_), .Y(_abc_40319_new_n788_));
NOR2X1 NOR2X1_54 ( .A(REG3_REG_3_), .B(REG3_REG_4_), .Y(_abc_40319_new_n805_));
NOR2X1 NOR2X1_55 ( .A(_abc_40319_new_n805_), .B(_abc_40319_new_n731_), .Y(_abc_40319_new_n806_));
NOR2X1 NOR2X1_56 ( .A(_abc_40319_new_n758_), .B(_abc_40319_new_n855_), .Y(_abc_40319_new_n856_));
NOR2X1 NOR2X1_57 ( .A(_abc_40319_new_n829_), .B(_abc_40319_new_n861_), .Y(_abc_40319_new_n865_));
NOR2X1 NOR2X1_58 ( .A(_abc_40319_new_n758_), .B(_abc_40319_new_n865_), .Y(_abc_40319_new_n866_));
NOR2X1 NOR2X1_59 ( .A(_abc_40319_new_n758_), .B(_abc_40319_new_n897_), .Y(_abc_40319_new_n898_));
NOR2X1 NOR2X1_6 ( .A(IR_REG_23_), .B(IR_REG_18_), .Y(_abc_40319_new_n539_));
NOR2X1 NOR2X1_60 ( .A(_abc_40319_new_n908_), .B(_abc_40319_new_n911_), .Y(_abc_40319_new_n912_));
NOR2X1 NOR2X1_61 ( .A(_abc_40319_new_n912_), .B(_abc_40319_new_n758_), .Y(_abc_40319_new_n924_));
NOR2X1 NOR2X1_62 ( .A(_abc_40319_new_n973_), .B(_abc_40319_new_n616_), .Y(_abc_40319_new_n974_));
NOR2X1 NOR2X1_63 ( .A(_abc_40319_new_n975_), .B(_abc_40319_new_n972_), .Y(_abc_40319_new_n976_));
NOR2X1 NOR2X1_64 ( .A(_abc_40319_new_n977_), .B(_abc_40319_new_n659_), .Y(_abc_40319_new_n978_));
NOR2X1 NOR2X1_65 ( .A(_abc_40319_new_n980_), .B(_abc_40319_new_n734_), .Y(_abc_40319_new_n982_));
NOR2X1 NOR2X1_66 ( .A(_abc_40319_new_n992_), .B(_abc_40319_new_n660_), .Y(_abc_40319_new_n993_));
NOR2X1 NOR2X1_67 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n972_), .Y(_abc_40319_new_n995_));
NOR2X1 NOR2X1_68 ( .A(_abc_40319_new_n668_), .B(_abc_40319_new_n616_), .Y(_abc_40319_new_n997_));
NOR2X1 NOR2X1_69 ( .A(_abc_40319_new_n608_), .B(_abc_40319_new_n749_), .Y(_abc_40319_new_n1004_));
NOR2X1 NOR2X1_7 ( .A(IR_REG_2_), .B(IR_REG_0_), .Y(_abc_40319_new_n545_));
NOR2X1 NOR2X1_70 ( .A(_abc_40319_new_n742_), .B(_abc_40319_new_n1005_), .Y(_abc_40319_new_n1006_));
NOR2X1 NOR2X1_71 ( .A(_abc_40319_new_n1007_), .B(_abc_40319_new_n972_), .Y(_abc_40319_new_n1008_));
NOR2X1 NOR2X1_72 ( .A(_abc_40319_new_n1023_), .B(_abc_40319_new_n1024_), .Y(_abc_40319_new_n1025_));
NOR2X1 NOR2X1_73 ( .A(_abc_40319_new_n1027_), .B(_abc_40319_new_n1026_), .Y(_abc_40319_new_n1028_));
NOR2X1 NOR2X1_74 ( .A(_abc_40319_new_n1030_), .B(_abc_40319_new_n1029_), .Y(_abc_40319_new_n1031_));
NOR2X1 NOR2X1_75 ( .A(_abc_40319_new_n1022_), .B(_abc_40319_new_n1032_), .Y(_abc_40319_new_n1033_));
NOR2X1 NOR2X1_76 ( .A(_abc_40319_new_n1021_), .B(_abc_40319_new_n1035_), .Y(_abc_40319_new_n1036_));
NOR2X1 NOR2X1_77 ( .A(_abc_40319_new_n1019_), .B(_abc_40319_new_n1037_), .Y(_abc_40319_new_n1039_));
NOR2X1 NOR2X1_78 ( .A(_abc_40319_new_n1047_), .B(_abc_40319_new_n1049_), .Y(_abc_40319_new_n1050_));
NOR2X1 NOR2X1_79 ( .A(_abc_40319_new_n1095_), .B(_abc_40319_new_n1099_), .Y(_abc_40319_new_n1100_));
NOR2X1 NOR2X1_8 ( .A(_abc_40319_new_n549_), .B(_abc_40319_new_n546_), .Y(_abc_40319_new_n550_));
NOR2X1 NOR2X1_80 ( .A(_abc_40319_new_n1066_), .B(_abc_40319_new_n1068_), .Y(_abc_40319_new_n1102_));
NOR2X1 NOR2X1_81 ( .A(_abc_40319_new_n1102_), .B(_abc_40319_new_n1104_), .Y(_abc_40319_new_n1105_));
NOR2X1 NOR2X1_82 ( .A(_abc_40319_new_n778_), .B(_abc_40319_new_n1128_), .Y(_abc_40319_new_n1129_));
NOR2X1 NOR2X1_83 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1129_), .Y(_abc_40319_new_n1137_));
NOR2X1 NOR2X1_84 ( .A(_abc_40319_new_n1136_), .B(_abc_40319_new_n1140_), .Y(_abc_40319_new_n1142_));
NOR2X1 NOR2X1_85 ( .A(_abc_40319_new_n1149_), .B(_abc_40319_new_n802_), .Y(_abc_40319_new_n1150_));
NOR2X1 NOR2X1_86 ( .A(_abc_40319_new_n1150_), .B(_abc_40319_new_n1155_), .Y(_abc_40319_new_n1156_));
NOR2X1 NOR2X1_87 ( .A(_abc_40319_new_n1158_), .B(_abc_40319_new_n1162_), .Y(_abc_40319_new_n1164_));
NOR2X1 NOR2X1_88 ( .A(IR_REG_14_), .B(_abc_40319_new_n552_), .Y(_abc_40319_new_n1166_));
NOR2X1 NOR2X1_89 ( .A(IR_REG_15_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n1168_));
NOR2X1 NOR2X1_9 ( .A(_abc_40319_new_n536_), .B(_abc_40319_new_n552_), .Y(_abc_40319_new_n553_));
NOR2X1 NOR2X1_90 ( .A(IR_REG_16_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n1170_));
NOR2X1 NOR2X1_91 ( .A(_abc_40319_new_n533_), .B(_abc_40319_new_n1168_), .Y(_abc_40319_new_n1171_));
NOR2X1 NOR2X1_92 ( .A(_abc_40319_new_n1181_), .B(_abc_40319_new_n1180_), .Y(_abc_40319_new_n1182_));
NOR2X1 NOR2X1_93 ( .A(REG3_REG_16_), .B(_abc_40319_new_n1182_), .Y(_abc_40319_new_n1183_));
NOR2X1 NOR2X1_94 ( .A(_abc_40319_new_n1184_), .B(_abc_40319_new_n1029_), .Y(_abc_40319_new_n1185_));
NOR2X1 NOR2X1_95 ( .A(_abc_40319_new_n1185_), .B(_abc_40319_new_n1183_), .Y(_abc_40319_new_n1186_));
NOR2X1 NOR2X1_96 ( .A(_abc_40319_new_n1201_), .B(_abc_40319_new_n1207_), .Y(_abc_40319_new_n1208_));
NOR2X1 NOR2X1_97 ( .A(_abc_40319_new_n1234_), .B(_abc_40319_new_n1237_), .Y(_abc_40319_new_n1239_));
NOR2X1 NOR2X1_98 ( .A(_abc_40319_new_n1251_), .B(_abc_40319_new_n1257_), .Y(_abc_40319_new_n1258_));
NOR2X1 NOR2X1_99 ( .A(IR_REG_8_), .B(_abc_40319_new_n686_), .Y(_abc_40319_new_n1267_));
NOR3X1 NOR3X1_1 ( .A(IR_REG_2_), .B(IR_REG_0_), .C(IR_REG_1_), .Y(_abc_40319_new_n526_));
NOR3X1 NOR3X1_10 ( .A(_abc_40319_new_n1965_), .B(_abc_40319_new_n1954_), .C(_abc_40319_new_n1969_), .Y(_abc_40319_new_n1970_));
NOR3X1 NOR3X1_11 ( .A(_abc_40319_new_n1890_), .B(_abc_40319_new_n1891_), .C(_abc_40319_new_n2271_), .Y(_abc_40319_new_n2272_));
NOR3X1 NOR3X1_12 ( .A(_abc_40319_new_n1910_), .B(_abc_40319_new_n1911_), .C(_abc_40319_new_n2279_), .Y(_abc_40319_new_n2280_));
NOR3X1 NOR3X1_13 ( .A(_abc_40319_new_n2355_), .B(_abc_40319_new_n2356_), .C(_abc_40319_new_n2351_), .Y(_abc_40319_new_n2357_));
NOR3X1 NOR3X1_14 ( .A(_abc_40319_new_n2337_), .B(_abc_40319_new_n2346_), .C(_abc_40319_new_n2347_), .Y(_abc_40319_new_n2371_));
NOR3X1 NOR3X1_15 ( .A(_abc_40319_new_n2387_), .B(_abc_40319_new_n2399_), .C(_abc_40319_new_n2379_), .Y(_abc_40319_new_n2400_));
NOR3X1 NOR3X1_16 ( .A(_abc_40319_new_n2244_), .B(_abc_40319_new_n2417_), .C(_abc_40319_new_n2418_), .Y(_abc_40319_new_n2419_));
NOR3X1 NOR3X1_17 ( .A(_abc_40319_new_n1276_), .B(_abc_40319_new_n1297_), .C(_abc_40319_new_n2968_), .Y(_abc_40319_new_n2969_));
NOR3X1 NOR3X1_18 ( .A(_abc_40319_new_n1325_), .B(_abc_40319_new_n1352_), .C(_abc_40319_new_n2970_), .Y(_abc_40319_new_n2971_));
NOR3X1 NOR3X1_19 ( .A(_abc_40319_new_n1175_), .B(_abc_40319_new_n1198_), .C(_abc_40319_new_n2972_), .Y(_abc_40319_new_n2973_));
NOR3X1 NOR3X1_2 ( .A(IR_REG_9_), .B(IR_REG_8_), .C(IR_REG_7_), .Y(_abc_40319_new_n528_));
NOR3X1 NOR3X1_20 ( .A(_abc_40319_new_n1443_), .B(_abc_40319_new_n1460_), .C(_abc_40319_new_n2974_), .Y(_abc_40319_new_n2975_));
NOR3X1 NOR3X1_21 ( .A(_abc_40319_new_n1080_), .B(_abc_40319_new_n1085_), .C(_abc_40319_new_n2976_), .Y(_abc_40319_new_n2977_));
NOR3X1 NOR3X1_22 ( .A(_abc_40319_new_n1582_), .B(_abc_40319_new_n2262_), .C(_abc_40319_new_n2978_), .Y(_abc_40319_new_n2982_));
NOR3X1 NOR3X1_23 ( .A(_abc_40319_new_n4053_), .B(_abc_40319_new_n4055_), .C(_abc_40319_new_n4054_), .Y(_abc_40319_new_n4056_));
NOR3X1 NOR3X1_3 ( .A(IR_REG_12_), .B(IR_REG_10_), .C(IR_REG_11_), .Y(_abc_40319_new_n530_));
NOR3X1 NOR3X1_4 ( .A(IR_REG_22_), .B(_abc_40319_new_n536_), .C(_abc_40319_new_n540_), .Y(_abc_40319_new_n541_));
NOR3X1 NOR3X1_5 ( .A(IR_REG_15_), .B(IR_REG_14_), .C(IR_REG_16_), .Y(_abc_40319_new_n595_));
NOR3X1 NOR3X1_6 ( .A(IR_REG_20_), .B(IR_REG_19_), .C(IR_REG_21_), .Y(_abc_40319_new_n597_));
NOR3X1 NOR3X1_7 ( .A(IR_REG_28_), .B(_abc_40319_new_n596_), .C(_abc_40319_new_n598_), .Y(_abc_40319_new_n599_));
NOR3X1 NOR3X1_8 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n596_), .C(_abc_40319_new_n598_), .Y(_abc_40319_new_n710_));
NOR3X1 NOR3X1_9 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n663_), .C(_abc_40319_new_n1870_), .Y(_abc_40319_new_n1875_));
OAI21X1 OAI21X1_1 ( .A(IR_REG_23_), .B(_abc_40319_new_n557_), .C(IR_REG_24_), .Y(_abc_40319_new_n558_));
OAI21X1 OAI21X1_10 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n606_), .C(_abc_40319_new_n607_), .Y(_abc_40319_new_n608_));
OAI21X1 OAI21X1_100 ( .A(_abc_40319_new_n658_), .B(_abc_40319_new_n991_), .C(_abc_40319_new_n1001_), .Y(_abc_40319_new_n1002_));
OAI21X1 OAI21X1_101 ( .A(_abc_40319_new_n996_), .B(_abc_40319_new_n659_), .C(_abc_40319_new_n1009_), .Y(_abc_40319_new_n1010_));
OAI21X1 OAI21X1_102 ( .A(_abc_40319_new_n735_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1012_));
OAI21X1 OAI21X1_103 ( .A(_abc_40319_new_n737_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1013_), .Y(_abc_40319_new_n1014_));
OAI21X1 OAI21X1_104 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n971_), .C(_abc_40319_new_n1015_), .Y(n1331));
OAI21X1 OAI21X1_105 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_27_), .Y(_abc_40319_new_n1017_));
OAI21X1 OAI21X1_106 ( .A(_abc_40319_new_n1019_), .B(_abc_40319_new_n1037_), .C(_abc_40319_new_n1020_), .Y(_abc_40319_new_n1038_));
OAI21X1 OAI21X1_107 ( .A(_abc_40319_new_n1042_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n1043_), .Y(_abc_40319_new_n1044_));
OAI21X1 OAI21X1_108 ( .A(_abc_40319_new_n778_), .B(_abc_40319_new_n1041_), .C(_abc_40319_new_n1045_), .Y(_abc_40319_new_n1046_));
OAI21X1 OAI21X1_109 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_26_), .Y(_abc_40319_new_n1054_));
OAI21X1 OAI21X1_11 ( .A(IR_REG_20_), .B(_abc_40319_new_n611_), .C(IR_REG_21_), .Y(_abc_40319_new_n612_));
OAI21X1 OAI21X1_110 ( .A(_abc_40319_new_n1057_), .B(_abc_40319_new_n1058_), .C(_abc_40319_new_n1019_), .Y(_abc_40319_new_n1059_));
OAI21X1 OAI21X1_111 ( .A(_abc_40319_new_n1061_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n1062_), .Y(_abc_40319_new_n1063_));
OAI21X1 OAI21X1_112 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_25_), .Y(_abc_40319_new_n1070_));
OAI21X1 OAI21X1_113 ( .A(_abc_40319_new_n1073_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n1074_), .Y(_abc_40319_new_n1075_));
OAI21X1 OAI21X1_114 ( .A(_abc_40319_new_n778_), .B(_abc_40319_new_n1072_), .C(_abc_40319_new_n1076_), .Y(_abc_40319_new_n1077_));
OAI21X1 OAI21X1_115 ( .A(_abc_40319_new_n1079_), .B(_abc_40319_new_n1082_), .C(_abc_40319_new_n1069_), .Y(_abc_40319_new_n1083_));
OAI21X1 OAI21X1_116 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_24_), .Y(_abc_40319_new_n1084_));
OAI21X1 OAI21X1_117 ( .A(_abc_40319_new_n1021_), .B(_abc_40319_new_n1035_), .C(_abc_40319_new_n1086_), .Y(_abc_40319_new_n1087_));
OAI21X1 OAI21X1_118 ( .A(_abc_40319_new_n1089_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n1090_), .Y(_abc_40319_new_n1091_));
OAI21X1 OAI21X1_119 ( .A(_abc_40319_new_n1083_), .B(_abc_40319_new_n1101_), .C(_abc_40319_new_n1105_), .Y(_abc_40319_new_n1106_));
OAI21X1 OAI21X1_12 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n613_), .C(_abc_40319_new_n610_), .Y(_abc_40319_new_n614_));
OAI21X1 OAI21X1_120 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_23_), .Y(_abc_40319_new_n1108_));
OAI21X1 OAI21X1_121 ( .A(_abc_40319_new_n1111_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n1112_), .Y(_abc_40319_new_n1113_));
OAI21X1 OAI21X1_122 ( .A(_abc_40319_new_n778_), .B(_abc_40319_new_n1110_), .C(_abc_40319_new_n1114_), .Y(_abc_40319_new_n1115_));
OAI21X1 OAI21X1_123 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_22_), .Y(_abc_40319_new_n1122_));
OAI21X1 OAI21X1_124 ( .A(_abc_40319_new_n1124_), .B(_abc_40319_new_n1126_), .C(_abc_40319_new_n1125_), .Y(_abc_40319_new_n1127_));
OAI21X1 OAI21X1_125 ( .A(_abc_40319_new_n1130_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n1133_), .Y(_abc_40319_new_n1134_));
OAI21X1 OAI21X1_126 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n1144_), .C(_abc_40319_new_n1145_), .Y(_abc_40319_new_n1146_));
OAI21X1 OAI21X1_127 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_18_), .Y(_abc_40319_new_n1147_));
OAI21X1 OAI21X1_128 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n1146_), .C(_abc_40319_new_n1147_), .Y(_abc_40319_new_n1148_));
OAI21X1 OAI21X1_129 ( .A(_abc_40319_new_n1030_), .B(_abc_40319_new_n1029_), .C(_abc_40319_new_n1151_), .Y(_abc_40319_new_n1152_));
OAI21X1 OAI21X1_13 ( .A(_abc_40319_new_n580_), .B(_abc_40319_new_n616_), .C(_abc_40319_new_n603_), .Y(_abc_40319_new_n617_));
OAI21X1 OAI21X1_130 ( .A(_abc_40319_new_n778_), .B(_abc_40319_new_n1153_), .C(_abc_40319_new_n1154_), .Y(_abc_40319_new_n1155_));
OAI21X1 OAI21X1_131 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1170_), .C(IR_REG_31_), .Y(_abc_40319_new_n1172_));
OAI21X1 OAI21X1_132 ( .A(IR_REG_31_), .B(IR_REG_16_), .C(_abc_40319_new_n1172_), .Y(_abc_40319_new_n1173_));
OAI21X1 OAI21X1_133 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_16_), .Y(_abc_40319_new_n1174_));
OAI21X1 OAI21X1_134 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n1173_), .C(_abc_40319_new_n1174_), .Y(_abc_40319_new_n1175_));
OAI21X1 OAI21X1_135 ( .A(_abc_40319_new_n1176_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n1177_), .Y(_abc_40319_new_n1178_));
OAI21X1 OAI21X1_136 ( .A(_abc_40319_new_n534_), .B(_abc_40319_new_n1170_), .C(_abc_40319_new_n604_), .Y(_abc_40319_new_n1194_));
OAI21X1 OAI21X1_137 ( .A(IR_REG_31_), .B(IR_REG_17_), .C(_abc_40319_new_n1195_), .Y(_abc_40319_new_n1196_));
OAI21X1 OAI21X1_138 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_17_), .Y(_abc_40319_new_n1197_));
OAI21X1 OAI21X1_139 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n1196_), .C(_abc_40319_new_n1197_), .Y(_abc_40319_new_n1198_));
OAI21X1 OAI21X1_14 ( .A(_abc_40319_new_n581_), .B(_abc_40319_new_n617_), .C(_abc_40319_new_n620_), .Y(n1341));
OAI21X1 OAI21X1_140 ( .A(_abc_40319_new_n1191_), .B(_abc_40319_new_n1193_), .C(_abc_40319_new_n1215_), .Y(_abc_40319_new_n1216_));
OAI21X1 OAI21X1_141 ( .A(IR_REG_14_), .B(_abc_40319_new_n552_), .C(IR_REG_15_), .Y(_abc_40319_new_n1218_));
OAI21X1 OAI21X1_142 ( .A(IR_REG_31_), .B(IR_REG_15_), .C(_abc_40319_new_n1220_), .Y(_abc_40319_new_n1221_));
OAI21X1 OAI21X1_143 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_15_), .Y(_abc_40319_new_n1222_));
OAI21X1 OAI21X1_144 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n1221_), .C(_abc_40319_new_n1222_), .Y(_abc_40319_new_n1223_));
OAI21X1 OAI21X1_145 ( .A(_abc_40319_new_n1227_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n1231_), .Y(_abc_40319_new_n1232_));
OAI21X1 OAI21X1_146 ( .A(_abc_40319_new_n527_), .B(_abc_40319_new_n531_), .C(IR_REG_14_), .Y(_abc_40319_new_n1241_));
OAI21X1 OAI21X1_147 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n1243_), .C(_abc_40319_new_n1244_), .Y(_abc_40319_new_n1245_));
OAI21X1 OAI21X1_148 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_14_), .Y(_abc_40319_new_n1247_));
OAI21X1 OAI21X1_149 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n1246_), .C(_abc_40319_new_n1247_), .Y(_abc_40319_new_n1248_));
OAI21X1 OAI21X1_15 ( .A(B_REG), .B(_abc_40319_new_n623_), .C(_abc_40319_new_n571_), .Y(_abc_40319_new_n626_));
OAI21X1 OAI21X1_150 ( .A(_abc_40319_new_n1027_), .B(_abc_40319_new_n1026_), .C(_abc_40319_new_n1253_), .Y(_abc_40319_new_n1254_));
OAI21X1 OAI21X1_151 ( .A(_abc_40319_new_n1252_), .B(_abc_40319_new_n802_), .C(_abc_40319_new_n1256_), .Y(_abc_40319_new_n1257_));
OAI21X1 OAI21X1_152 ( .A(IR_REG_7_), .B(_abc_40319_new_n938_), .C(IR_REG_8_), .Y(_abc_40319_new_n1269_));
OAI21X1 OAI21X1_153 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n1271_), .C(_abc_40319_new_n1272_), .Y(_abc_40319_new_n1273_));
OAI21X1 OAI21X1_154 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_8_), .Y(_abc_40319_new_n1275_));
OAI21X1 OAI21X1_155 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n1274_), .C(_abc_40319_new_n1275_), .Y(_abc_40319_new_n1276_));
OAI21X1 OAI21X1_156 ( .A(_abc_40319_new_n962_), .B(_abc_40319_new_n762_), .C(_abc_40319_new_n964_), .Y(_abc_40319_new_n1286_));
OAI21X1 OAI21X1_157 ( .A(IR_REG_8_), .B(_abc_40319_new_n686_), .C(IR_REG_9_), .Y(_abc_40319_new_n1291_));
OAI21X1 OAI21X1_158 ( .A(IR_REG_31_), .B(_abc_40319_new_n1289_), .C(_abc_40319_new_n1293_), .Y(_abc_40319_new_n1294_));
OAI21X1 OAI21X1_159 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_9_), .Y(_abc_40319_new_n1296_));
OAI21X1 OAI21X1_16 ( .A(D_REG_1_), .B(_abc_40319_new_n628_), .C(_abc_40319_new_n629_), .Y(_abc_40319_new_n630_));
OAI21X1 OAI21X1_160 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n1295_), .C(_abc_40319_new_n1296_), .Y(_abc_40319_new_n1297_));
OAI21X1 OAI21X1_161 ( .A(_abc_40319_new_n980_), .B(_abc_40319_new_n734_), .C(_abc_40319_new_n1300_), .Y(_abc_40319_new_n1301_));
OAI21X1 OAI21X1_162 ( .A(_abc_40319_new_n1298_), .B(_abc_40319_new_n802_), .C(_abc_40319_new_n1303_), .Y(_abc_40319_new_n1304_));
OAI21X1 OAI21X1_163 ( .A(_abc_40319_new_n1318_), .B(_abc_40319_new_n1290_), .C(IR_REG_13_), .Y(_abc_40319_new_n1319_));
OAI21X1 OAI21X1_164 ( .A(_abc_40319_new_n527_), .B(_abc_40319_new_n531_), .C(_abc_40319_new_n1319_), .Y(_abc_40319_new_n1320_));
OAI21X1 OAI21X1_165 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n1320_), .C(_abc_40319_new_n1321_), .Y(_abc_40319_new_n1322_));
OAI21X1 OAI21X1_166 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_13_), .Y(_abc_40319_new_n1324_));
OAI21X1 OAI21X1_167 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n1323_), .C(_abc_40319_new_n1324_), .Y(_abc_40319_new_n1325_));
OAI21X1 OAI21X1_168 ( .A(_abc_40319_new_n1327_), .B(_abc_40319_new_n1026_), .C(_abc_40319_new_n1328_), .Y(_abc_40319_new_n1329_));
OAI21X1 OAI21X1_169 ( .A(IR_REG_11_), .B(_abc_40319_new_n1344_), .C(IR_REG_12_), .Y(_abc_40319_new_n1345_));
OAI21X1 OAI21X1_17 ( .A(_abc_40319_new_n631_), .B(_abc_40319_new_n653_), .C(_abc_40319_new_n627_), .Y(_abc_40319_new_n654_));
OAI21X1 OAI21X1_170 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(_abc_40319_new_n1350_), .Y(_abc_40319_new_n1351_));
OAI21X1 OAI21X1_171 ( .A(_abc_40319_new_n1356_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n1358_), .Y(_abc_40319_new_n1359_));
OAI21X1 OAI21X1_172 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n1367_), .C(_abc_40319_new_n1368_), .Y(_abc_40319_new_n1369_));
OAI21X1 OAI21X1_173 ( .A(_abc_40319_new_n1023_), .B(_abc_40319_new_n1299_), .C(_abc_40319_new_n1024_), .Y(_abc_40319_new_n1376_));
OAI21X1 OAI21X1_174 ( .A(_abc_40319_new_n778_), .B(_abc_40319_new_n1377_), .C(_abc_40319_new_n1375_), .Y(_abc_40319_new_n1378_));
OAI21X1 OAI21X1_175 ( .A(_abc_40319_new_n1382_), .B(_abc_40319_new_n1384_), .C(_abc_40319_new_n1365_), .Y(_abc_40319_new_n1385_));
OAI21X1 OAI21X1_176 ( .A(IR_REG_9_), .B(_abc_40319_new_n1268_), .C(IR_REG_10_), .Y(_abc_40319_new_n1387_));
OAI21X1 OAI21X1_177 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n1388_), .C(_abc_40319_new_n1389_), .Y(_abc_40319_new_n1390_));
OAI21X1 OAI21X1_178 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_10_), .Y(_abc_40319_new_n1392_));
OAI21X1 OAI21X1_179 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n1391_), .C(_abc_40319_new_n1392_), .Y(_abc_40319_new_n1393_));
OAI21X1 OAI21X1_18 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n661_), .C(_abc_40319_new_n662_), .Y(_abc_40319_new_n663_));
OAI21X1 OAI21X1_180 ( .A(_abc_40319_new_n1394_), .B(_abc_40319_new_n802_), .C(_abc_40319_new_n1395_), .Y(_abc_40319_new_n1396_));
OAI21X1 OAI21X1_181 ( .A(_abc_40319_new_n1404_), .B(_abc_40319_new_n1406_), .C(_abc_40319_new_n1386_), .Y(_abc_40319_new_n1407_));
OAI21X1 OAI21X1_182 ( .A(_abc_40319_new_n1407_), .B(_abc_40319_new_n1317_), .C(_abc_40319_new_n1418_), .Y(_abc_40319_new_n1419_));
OAI21X1 OAI21X1_183 ( .A(_abc_40319_new_n1424_), .B(_abc_40319_new_n1425_), .C(_abc_40319_new_n1215_), .Y(_abc_40319_new_n1426_));
OAI21X1 OAI21X1_184 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_19_), .Y(_abc_40319_new_n1428_));
OAI21X1 OAI21X1_185 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n749_), .C(_abc_40319_new_n1428_), .Y(_abc_40319_new_n1429_));
OAI21X1 OAI21X1_186 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_20_), .Y(_abc_40319_new_n1442_));
OAI21X1 OAI21X1_187 ( .A(_abc_40319_new_n1022_), .B(_abc_40319_new_n1032_), .C(_abc_40319_new_n1444_), .Y(_abc_40319_new_n1445_));
OAI21X1 OAI21X1_188 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_21_), .Y(_abc_40319_new_n1459_));
OAI21X1 OAI21X1_189 ( .A(_abc_40319_new_n1471_), .B(_abc_40319_new_n1474_), .C(_abc_40319_new_n1458_), .Y(_abc_40319_new_n1475_));
OAI21X1 OAI21X1_19 ( .A(IR_REG_18_), .B(_abc_40319_new_n604_), .C(IR_REG_19_), .Y(_abc_40319_new_n664_));
OAI21X1 OAI21X1_190 ( .A(_abc_40319_new_n1439_), .B(_abc_40319_new_n1441_), .C(_abc_40319_new_n1476_), .Y(_abc_40319_new_n1477_));
OAI21X1 OAI21X1_191 ( .A(_abc_40319_new_n1480_), .B(_abc_40319_new_n1475_), .C(_abc_40319_new_n1484_), .Y(_abc_40319_new_n1485_));
OAI21X1 OAI21X1_192 ( .A(_abc_40319_new_n1471_), .B(_abc_40319_new_n1474_), .C(_abc_40319_new_n1485_), .Y(_abc_40319_new_n1486_));
OAI21X1 OAI21X1_193 ( .A(_abc_40319_new_n1053_), .B(_abc_40319_new_n1493_), .C(_abc_40319_new_n676_), .Y(_abc_40319_new_n1495_));
OAI21X1 OAI21X1_194 ( .A(_abc_40319_new_n1020_), .B(_abc_40319_new_n1056_), .C(REG3_REG_28_), .Y(_abc_40319_new_n1497_));
OAI21X1 OAI21X1_195 ( .A(_abc_40319_new_n1500_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n1501_), .Y(_abc_40319_new_n1502_));
OAI21X1 OAI21X1_196 ( .A(_abc_40319_new_n1020_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1507_));
OAI21X1 OAI21X1_197 ( .A(_abc_40319_new_n1041_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1508_), .Y(_abc_40319_new_n1509_));
OAI21X1 OAI21X1_198 ( .A(_abc_40319_new_n1494_), .B(_abc_40319_new_n1495_), .C(_abc_40319_new_n1510_), .Y(n1326));
OAI21X1 OAI21X1_199 ( .A(_abc_40319_new_n1517_), .B(_abc_40319_new_n1515_), .C(_abc_40319_new_n976_), .Y(_abc_40319_new_n1518_));
OAI21X1 OAI21X1_2 ( .A(_abc_40319_new_n523_), .B(IR_REG_31_), .C(_abc_40319_new_n559_), .Y(_abc_40319_new_n560_));
OAI21X1 OAI21X1_20 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n665_), .C(_abc_40319_new_n666_), .Y(_abc_40319_new_n667_));
OAI21X1 OAI21X1_200 ( .A(_abc_40319_new_n1261_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1520_), .Y(_abc_40319_new_n1521_));
OAI21X1 OAI21X1_201 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1513_), .C(_abc_40319_new_n1523_), .Y(n1321));
OAI21X1 OAI21X1_202 ( .A(_abc_40319_new_n1525_), .B(_abc_40319_new_n1526_), .C(_abc_40319_new_n1527_), .Y(_abc_40319_new_n1528_));
OAI21X1 OAI21X1_203 ( .A(_abc_40319_new_n1108_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1532_), .Y(_abc_40319_new_n1533_));
OAI21X1 OAI21X1_204 ( .A(_abc_40319_new_n1541_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1542_), .Y(_abc_40319_new_n1543_));
OAI21X1 OAI21X1_205 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1538_), .C(_abc_40319_new_n1545_), .Y(n1311));
OAI21X1 OAI21X1_206 ( .A(_abc_40319_new_n1548_), .B(_abc_40319_new_n1550_), .C(_abc_40319_new_n903_), .Y(_abc_40319_new_n1551_));
OAI21X1 OAI21X1_207 ( .A(_abc_40319_new_n844_), .B(_abc_40319_new_n1552_), .C(_abc_40319_new_n1551_), .Y(_abc_40319_new_n1553_));
OAI21X1 OAI21X1_208 ( .A(_abc_40319_new_n843_), .B(_abc_40319_new_n932_), .C(_abc_40319_new_n1553_), .Y(_abc_40319_new_n1554_));
OAI21X1 OAI21X1_209 ( .A(_abc_40319_new_n729_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1558_));
OAI21X1 OAI21X1_21 ( .A(_abc_40319_new_n660_), .B(_abc_40319_new_n668_), .C(_abc_40319_new_n616_), .Y(_abc_40319_new_n669_));
OAI21X1 OAI21X1_210 ( .A(REG3_REG_3_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1559_), .Y(_abc_40319_new_n1560_));
OAI21X1 OAI21X1_211 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1555_), .C(_abc_40319_new_n1561_), .Y(n1306));
OAI21X1 OAI21X1_212 ( .A(_abc_40319_new_n1568_), .B(_abc_40319_new_n1566_), .C(_abc_40319_new_n976_), .Y(_abc_40319_new_n1569_));
OAI21X1 OAI21X1_213 ( .A(_abc_40319_new_n1022_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1571_));
OAI21X1 OAI21X1_214 ( .A(_abc_40319_new_n1570_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1572_), .Y(_abc_40319_new_n1573_));
OAI21X1 OAI21X1_215 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1565_), .C(_abc_40319_new_n1575_), .Y(n1301));
OAI21X1 OAI21X1_216 ( .A(_abc_40319_new_n1491_), .B(_abc_40319_new_n1577_), .C(_abc_40319_new_n1578_), .Y(_abc_40319_new_n1579_));
OAI21X1 OAI21X1_217 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_28_), .Y(_abc_40319_new_n1581_));
OAI21X1 OAI21X1_218 ( .A(_abc_40319_new_n1107_), .B(_abc_40319_new_n1492_), .C(_abc_40319_new_n1051_), .Y(_abc_40319_new_n1588_));
OAI21X1 OAI21X1_219 ( .A(_abc_40319_new_n1581_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1602_), .Y(_abc_40319_new_n1603_));
OAI21X1 OAI21X1_22 ( .A(IR_REG_6_), .B(_abc_40319_new_n527_), .C(IR_REG_7_), .Y(_abc_40319_new_n687_));
OAI21X1 OAI21X1_220 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1591_), .C(_abc_40319_new_n1605_), .Y(n1296));
OAI21X1 OAI21X1_221 ( .A(_abc_40319_new_n811_), .B(_abc_40319_new_n815_), .C(_abc_40319_new_n935_), .Y(_abc_40319_new_n1609_));
OAI21X1 OAI21X1_222 ( .A(_abc_40319_new_n1280_), .B(_abc_40319_new_n1609_), .C(_abc_40319_new_n1610_), .Y(_abc_40319_new_n1611_));
OAI21X1 OAI21X1_223 ( .A(_abc_40319_new_n1608_), .B(_abc_40319_new_n1611_), .C(_abc_40319_new_n1612_), .Y(_abc_40319_new_n1613_));
OAI21X1 OAI21X1_224 ( .A(_abc_40319_new_n980_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1616_));
OAI21X1 OAI21X1_225 ( .A(_abc_40319_new_n1615_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1617_), .Y(_abc_40319_new_n1618_));
OAI21X1 OAI21X1_226 ( .A(_abc_40319_new_n1624_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1625_));
OAI21X1 OAI21X1_227 ( .A(_abc_40319_new_n1624_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1626_), .Y(_abc_40319_new_n1627_));
OAI21X1 OAI21X1_228 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1622_), .C(_abc_40319_new_n1628_), .Y(n1286));
OAI21X1 OAI21X1_229 ( .A(_abc_40319_new_n1439_), .B(_abc_40319_new_n1441_), .C(_abc_40319_new_n1563_), .Y(_abc_40319_new_n1633_));
OAI21X1 OAI21X1_23 ( .A(IR_REG_31_), .B(_abc_40319_new_n684_), .C(_abc_40319_new_n689_), .Y(_abc_40319_new_n690_));
OAI21X1 OAI21X1_230 ( .A(_abc_40319_new_n1632_), .B(_abc_40319_new_n1481_), .C(_abc_40319_new_n1635_), .Y(_abc_40319_new_n1636_));
OAI21X1 OAI21X1_231 ( .A(_abc_40319_new_n1483_), .B(_abc_40319_new_n1634_), .C(_abc_40319_new_n1637_), .Y(_abc_40319_new_n1638_));
OAI21X1 OAI21X1_232 ( .A(_abc_40319_new_n1124_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1640_));
OAI21X1 OAI21X1_233 ( .A(_abc_40319_new_n1463_), .B(_abc_40319_new_n1001_), .C(_abc_40319_new_n1641_), .Y(_abc_40319_new_n1642_));
OAI21X1 OAI21X1_234 ( .A(_abc_40319_new_n991_), .B(_abc_40319_new_n1631_), .C(_abc_40319_new_n1643_), .Y(n1281));
OAI21X1 OAI21X1_235 ( .A(_abc_40319_new_n1536_), .B(_abc_40319_new_n1317_), .C(_abc_40319_new_n1408_), .Y(_abc_40319_new_n1647_));
OAI21X1 OAI21X1_236 ( .A(_abc_40319_new_n1645_), .B(_abc_40319_new_n1648_), .C(_abc_40319_new_n676_), .Y(_abc_40319_new_n1650_));
OAI21X1 OAI21X1_237 ( .A(_abc_40319_new_n1652_), .B(_abc_40319_new_n1651_), .C(_abc_40319_new_n976_), .Y(_abc_40319_new_n1653_));
OAI21X1 OAI21X1_238 ( .A(_abc_40319_new_n1654_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1655_), .Y(_abc_40319_new_n1656_));
OAI21X1 OAI21X1_239 ( .A(_abc_40319_new_n1649_), .B(_abc_40319_new_n1650_), .C(_abc_40319_new_n1658_), .Y(n1276));
OAI21X1 OAI21X1_24 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_7_), .Y(_abc_40319_new_n697_));
OAI21X1 OAI21X1_240 ( .A(_abc_40319_new_n1100_), .B(_abc_40319_new_n1664_), .C(_abc_40319_new_n1661_), .Y(_abc_40319_new_n1665_));
OAI21X1 OAI21X1_241 ( .A(_abc_40319_new_n1057_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1668_));
OAI21X1 OAI21X1_242 ( .A(_abc_40319_new_n1072_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1669_), .Y(_abc_40319_new_n1670_));
OAI21X1 OAI21X1_243 ( .A(_abc_40319_new_n1663_), .B(_abc_40319_new_n1666_), .C(_abc_40319_new_n1671_), .Y(n1271));
OAI21X1 OAI21X1_244 ( .A(_abc_40319_new_n1676_), .B(_abc_40319_new_n1674_), .C(_abc_40319_new_n676_), .Y(_abc_40319_new_n1678_));
OAI21X1 OAI21X1_245 ( .A(_abc_40319_new_n1184_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1680_));
OAI21X1 OAI21X1_246 ( .A(_abc_40319_new_n1187_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1681_), .Y(_abc_40319_new_n1682_));
OAI21X1 OAI21X1_247 ( .A(_abc_40319_new_n1677_), .B(_abc_40319_new_n1678_), .C(_abc_40319_new_n1683_), .Y(n1266));
OAI21X1 OAI21X1_248 ( .A(_abc_40319_new_n1609_), .B(_abc_40319_new_n1685_), .C(_abc_40319_new_n1686_), .Y(_abc_40319_new_n1687_));
OAI21X1 OAI21X1_249 ( .A(_abc_40319_new_n779_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1689_));
OAI21X1 OAI21X1_25 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n691_), .C(_abc_40319_new_n697_), .Y(_abc_40319_new_n698_));
OAI21X1 OAI21X1_250 ( .A(_abc_40319_new_n781_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1690_), .Y(_abc_40319_new_n1691_));
OAI21X1 OAI21X1_251 ( .A(_abc_40319_new_n1424_), .B(_abc_40319_new_n1674_), .C(_abc_40319_new_n1694_), .Y(_abc_40319_new_n1695_));
OAI21X1 OAI21X1_252 ( .A(_abc_40319_new_n1675_), .B(_abc_40319_new_n1673_), .C(_abc_40319_new_n1423_), .Y(_abc_40319_new_n1698_));
OAI21X1 OAI21X1_253 ( .A(_abc_40319_new_n1697_), .B(_abc_40319_new_n1698_), .C(_abc_40319_new_n1695_), .Y(_abc_40319_new_n1699_));
OAI21X1 OAI21X1_254 ( .A(_abc_40319_new_n1203_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1702_));
OAI21X1 OAI21X1_255 ( .A(_abc_40319_new_n1206_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1703_), .Y(_abc_40319_new_n1704_));
OAI21X1 OAI21X1_256 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1699_), .C(_abc_40319_new_n1705_), .Y(n1256));
OAI21X1 OAI21X1_257 ( .A(_abc_40319_new_n1577_), .B(_abc_40319_new_n1707_), .C(_abc_40319_new_n1708_), .Y(_abc_40319_new_n1709_));
OAI21X1 OAI21X1_258 ( .A(_abc_40319_new_n1084_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1715_), .Y(_abc_40319_new_n1716_));
OAI21X1 OAI21X1_259 ( .A(_abc_40319_new_n1719_), .B(_abc_40319_new_n1720_), .C(_abc_40319_new_n1721_), .Y(_abc_40319_new_n1722_));
OAI21X1 OAI21X1_26 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n591_), .C(IR_REG_30_), .Y(_abc_40319_new_n706_));
OAI21X1 OAI21X1_260 ( .A(_abc_40319_new_n1724_), .B(_abc_40319_new_n1723_), .C(_abc_40319_new_n976_), .Y(_abc_40319_new_n1725_));
OAI21X1 OAI21X1_261 ( .A(_abc_40319_new_n730_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1727_));
OAI21X1 OAI21X1_262 ( .A(_abc_40319_new_n1726_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1728_), .Y(_abc_40319_new_n1729_));
OAI21X1 OAI21X1_263 ( .A(_abc_40319_new_n1316_), .B(_abc_40319_new_n1733_), .C(_abc_40319_new_n676_), .Y(_abc_40319_new_n1735_));
OAI21X1 OAI21X1_264 ( .A(_abc_40319_new_n1737_), .B(_abc_40319_new_n1736_), .C(_abc_40319_new_n976_), .Y(_abc_40319_new_n1738_));
OAI21X1 OAI21X1_265 ( .A(_abc_40319_new_n1300_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1740_));
OAI21X1 OAI21X1_266 ( .A(_abc_40319_new_n1739_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1741_), .Y(_abc_40319_new_n1742_));
OAI21X1 OAI21X1_267 ( .A(_abc_40319_new_n1734_), .B(_abc_40319_new_n1735_), .C(_abc_40319_new_n1744_), .Y(n1241));
OAI21X1 OAI21X1_268 ( .A(_abc_40319_new_n1750_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1752_));
OAI21X1 OAI21X1_269 ( .A(_abc_40319_new_n1750_), .B(_abc_40319_new_n1001_), .C(_abc_40319_new_n1753_), .Y(_abc_40319_new_n1754_));
OAI21X1 OAI21X1_27 ( .A(_abc_40319_new_n712_), .B(_abc_40319_new_n713_), .C(IR_REG_31_), .Y(_abc_40319_new_n714_));
OAI21X1 OAI21X1_270 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1749_), .C(_abc_40319_new_n1755_), .Y(n1236));
OAI21X1 OAI21X1_271 ( .A(_abc_40319_new_n1444_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1762_));
OAI21X1 OAI21X1_272 ( .A(_abc_40319_new_n1446_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1763_), .Y(_abc_40319_new_n1764_));
OAI21X1 OAI21X1_273 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1758_), .C(_abc_40319_new_n1765_), .Y(n1231));
OAI21X1 OAI21X1_274 ( .A(_abc_40319_new_n1413_), .B(_abc_40319_new_n1767_), .C(_abc_40319_new_n1365_), .Y(_abc_40319_new_n1768_));
OAI21X1 OAI21X1_275 ( .A(_abc_40319_new_n1415_), .B(_abc_40319_new_n1768_), .C(_abc_40319_new_n1771_), .Y(_abc_40319_new_n1772_));
OAI21X1 OAI21X1_276 ( .A(_abc_40319_new_n1328_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1776_));
OAI21X1 OAI21X1_277 ( .A(_abc_40319_new_n1331_), .B(_abc_40319_new_n1001_), .C(_abc_40319_new_n1777_), .Y(_abc_40319_new_n1778_));
OAI21X1 OAI21X1_278 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1772_), .C(_abc_40319_new_n1779_), .Y(n1226));
OAI21X1 OAI21X1_279 ( .A(_abc_40319_new_n1781_), .B(_abc_40319_new_n1783_), .C(_abc_40319_new_n1784_), .Y(_abc_40319_new_n1785_));
OAI21X1 OAI21X1_28 ( .A(_abc_40319_new_n717_), .B(_abc_40319_new_n718_), .C(IR_REG_31_), .Y(_abc_40319_new_n719_));
OAI21X1 OAI21X1_280 ( .A(_abc_40319_new_n1122_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1789_), .Y(_abc_40319_new_n1790_));
OAI21X1 OAI21X1_281 ( .A(_abc_40319_new_n1797_), .B(_abc_40319_new_n1795_), .C(_abc_40319_new_n976_), .Y(_abc_40319_new_n1798_));
OAI21X1 OAI21X1_282 ( .A(_abc_40319_new_n1370_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1800_), .Y(_abc_40319_new_n1801_));
OAI21X1 OAI21X1_283 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1794_), .C(_abc_40319_new_n1803_), .Y(n1216));
OAI21X1 OAI21X1_284 ( .A(_abc_40319_new_n1551_), .B(_abc_40319_new_n1806_), .C(_abc_40319_new_n1807_), .Y(_abc_40319_new_n1808_));
OAI21X1 OAI21X1_285 ( .A(_abc_40319_new_n1810_), .B(_abc_40319_new_n1809_), .C(_abc_40319_new_n976_), .Y(_abc_40319_new_n1811_));
OAI21X1 OAI21X1_286 ( .A(_abc_40319_new_n1812_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1813_));
OAI21X1 OAI21X1_287 ( .A(_abc_40319_new_n853_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1814_), .Y(_abc_40319_new_n1815_));
OAI21X1 OAI21X1_288 ( .A(_abc_40319_new_n1818_), .B(_abc_40319_new_n1819_), .C(_abc_40319_new_n1820_), .Y(_abc_40319_new_n1821_));
OAI21X1 OAI21X1_289 ( .A(_abc_40319_new_n1151_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1825_));
OAI21X1 OAI21X1_29 ( .A(IR_REG_28_), .B(_abc_40319_new_n591_), .C(IR_REG_29_), .Y(_abc_40319_new_n720_));
OAI21X1 OAI21X1_290 ( .A(_abc_40319_new_n1159_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1826_), .Y(_abc_40319_new_n1827_));
OAI21X1 OAI21X1_291 ( .A(_abc_40319_new_n1831_), .B(_abc_40319_new_n937_), .C(_abc_40319_new_n676_), .Y(_abc_40319_new_n1833_));
OAI21X1 OAI21X1_292 ( .A(_abc_40319_new_n728_), .B(_abc_40319_new_n1011_), .C(nRESET_G), .Y(_abc_40319_new_n1837_));
OAI21X1 OAI21X1_293 ( .A(_abc_40319_new_n949_), .B(_abc_40319_new_n1003_), .C(_abc_40319_new_n1838_), .Y(_abc_40319_new_n1839_));
OAI21X1 OAI21X1_294 ( .A(_abc_40319_new_n1833_), .B(_abc_40319_new_n1832_), .C(_abc_40319_new_n1840_), .Y(n1201));
OAI21X1 OAI21X1_295 ( .A(_abc_40319_new_n1095_), .B(_abc_40319_new_n1099_), .C(_abc_40319_new_n1103_), .Y(_abc_40319_new_n1842_));
OAI21X1 OAI21X1_296 ( .A(_abc_40319_new_n1842_), .B(_abc_40319_new_n1664_), .C(_abc_40319_new_n1843_), .Y(_abc_40319_new_n1844_));
OAI21X1 OAI21X1_297 ( .A(_abc_40319_new_n1054_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1853_), .Y(_abc_40319_new_n1854_));
OAI21X1 OAI21X1_298 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n1849_), .C(_abc_40319_new_n1856_), .Y(n1196));
OAI21X1 OAI21X1_299 ( .A(_abc_40319_new_n1858_), .B(_abc_40319_new_n1859_), .C(_abc_40319_new_n1860_), .Y(_abc_40319_new_n1861_));
OAI21X1 OAI21X1_3 ( .A(IR_REG_24_), .B(_abc_40319_new_n563_), .C(IR_REG_25_), .Y(_abc_40319_new_n564_));
OAI21X1 OAI21X1_30 ( .A(_abc_40319_new_n728_), .B(_abc_40319_new_n732_), .C(_abc_40319_new_n735_), .Y(_abc_40319_new_n736_));
OAI21X1 OAI21X1_300 ( .A(_abc_40319_new_n1863_), .B(_abc_40319_new_n1862_), .C(_abc_40319_new_n976_), .Y(_abc_40319_new_n1864_));
OAI21X1 OAI21X1_301 ( .A(_abc_40319_new_n1865_), .B(_abc_40319_new_n1519_), .C(_abc_40319_new_n1866_), .Y(_abc_40319_new_n1867_));
OAI21X1 OAI21X1_302 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_31_), .Y(_abc_40319_new_n1876_));
OAI21X1 OAI21X1_303 ( .A(_abc_40319_new_n1879_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n1880_), .Y(_abc_40319_new_n1881_));
OAI21X1 OAI21X1_304 ( .A(_abc_40319_new_n855_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1892_), .Y(_abc_40319_new_n1893_));
OAI21X1 OAI21X1_305 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n663_), .C(_abc_40319_new_n580_), .Y(_abc_40319_new_n1894_));
OAI21X1 OAI21X1_306 ( .A(_abc_40319_new_n885_), .B(_abc_40319_new_n889_), .C(_abc_40319_new_n895_), .Y(_abc_40319_new_n1898_));
OAI21X1 OAI21X1_307 ( .A(_abc_40319_new_n908_), .B(_abc_40319_new_n911_), .C(_abc_40319_new_n922_), .Y(_abc_40319_new_n1899_));
OAI21X1 OAI21X1_308 ( .A(_abc_40319_new_n895_), .B(_abc_40319_new_n880_), .C(_abc_40319_new_n1875_), .Y(_abc_40319_new_n1901_));
OAI21X1 OAI21X1_309 ( .A(_abc_40319_new_n1900_), .B(_abc_40319_new_n1901_), .C(_abc_40319_new_n1907_), .Y(_abc_40319_new_n1908_));
OAI21X1 OAI21X1_31 ( .A(_abc_40319_new_n604_), .B(_abc_40319_new_n555_), .C(_abc_40319_new_n612_), .Y(_abc_40319_new_n747_));
OAI21X1 OAI21X1_310 ( .A(_abc_40319_new_n865_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1912_), .Y(_abc_40319_new_n1913_));
OAI21X1 OAI21X1_311 ( .A(_abc_40319_new_n1726_), .B(_abc_40319_new_n1874_), .C(_abc_40319_new_n580_), .Y(_abc_40319_new_n1917_));
OAI21X1 OAI21X1_312 ( .A(_abc_40319_new_n1556_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1919_), .Y(_abc_40319_new_n1920_));
OAI21X1 OAI21X1_313 ( .A(_abc_40319_new_n1916_), .B(_abc_40319_new_n1909_), .C(_abc_40319_new_n1921_), .Y(_abc_40319_new_n1922_));
OAI21X1 OAI21X1_314 ( .A(_abc_40319_new_n754_), .B(_abc_40319_new_n753_), .C(_abc_40319_new_n1875_), .Y(_abc_40319_new_n1924_));
OAI21X1 OAI21X1_315 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n663_), .C(_abc_40319_new_n698_), .Y(_abc_40319_new_n1925_));
OAI21X1 OAI21X1_316 ( .A(_abc_40319_new_n953_), .B(_abc_40319_new_n950_), .C(_abc_40319_new_n1870_), .Y(_abc_40319_new_n1926_));
OAI21X1 OAI21X1_317 ( .A(_abc_40319_new_n950_), .B(_abc_40319_new_n953_), .C(_abc_40319_new_n1875_), .Y(_abc_40319_new_n1931_));
OAI21X1 OAI21X1_318 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n663_), .C(_abc_40319_new_n944_), .Y(_abc_40319_new_n1932_));
OAI21X1 OAI21X1_319 ( .A(_abc_40319_new_n782_), .B(_abc_40319_new_n775_), .C(_abc_40319_new_n1870_), .Y(_abc_40319_new_n1933_));
OAI21X1 OAI21X1_32 ( .A(_abc_40319_new_n751_), .B(_abc_40319_new_n746_), .C(_abc_40319_new_n698_), .Y(_abc_40319_new_n752_));
OAI21X1 OAI21X1_320 ( .A(_abc_40319_new_n775_), .B(_abc_40319_new_n782_), .C(_abc_40319_new_n1875_), .Y(_abc_40319_new_n1936_));
OAI21X1 OAI21X1_321 ( .A(_abc_40319_new_n1396_), .B(_abc_40319_new_n1400_), .C(_abc_40319_new_n1875_), .Y(_abc_40319_new_n1944_));
OAI21X1 OAI21X1_322 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n663_), .C(_abc_40319_new_n1393_), .Y(_abc_40319_new_n1945_));
OAI21X1 OAI21X1_323 ( .A(_abc_40319_new_n1307_), .B(_abc_40319_new_n1304_), .C(_abc_40319_new_n1870_), .Y(_abc_40319_new_n1946_));
OAI21X1 OAI21X1_324 ( .A(_abc_40319_new_n1308_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1949_), .Y(_abc_40319_new_n1950_));
OAI21X1 OAI21X1_325 ( .A(_abc_40319_new_n1957_), .B(_abc_40319_new_n1958_), .C(_abc_40319_new_n1875_), .Y(_abc_40319_new_n1959_));
OAI21X1 OAI21X1_326 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n663_), .C(_abc_40319_new_n1276_), .Y(_abc_40319_new_n1960_));
OAI21X1 OAI21X1_327 ( .A(_abc_40319_new_n754_), .B(_abc_40319_new_n753_), .C(_abc_40319_new_n1870_), .Y(_abc_40319_new_n1961_));
OAI21X1 OAI21X1_328 ( .A(_abc_40319_new_n1956_), .B(_abc_40319_new_n1955_), .C(_abc_40319_new_n1964_), .Y(_abc_40319_new_n1965_));
OAI21X1 OAI21X1_329 ( .A(_abc_40319_new_n1514_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1975_), .Y(_abc_40319_new_n1976_));
OAI21X1 OAI21X1_33 ( .A(_abc_40319_new_n753_), .B(_abc_40319_new_n754_), .C(_abc_40319_new_n679_), .Y(_abc_40319_new_n755_));
OAI21X1 OAI21X1_330 ( .A(_abc_40319_new_n1977_), .B(_abc_40319_new_n1976_), .C(_abc_40319_new_n1978_), .Y(_abc_40319_new_n1979_));
OAI21X1 OAI21X1_331 ( .A(_abc_40319_new_n1355_), .B(_abc_40319_new_n1359_), .C(_abc_40319_new_n1875_), .Y(_abc_40319_new_n1980_));
OAI21X1 OAI21X1_332 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n1378_), .C(_abc_40319_new_n1870_), .Y(_abc_40319_new_n1982_));
OAI21X1 OAI21X1_333 ( .A(_abc_40319_new_n1977_), .B(_abc_40319_new_n1976_), .C(_abc_40319_new_n1983_), .Y(_abc_40319_new_n1984_));
OAI21X1 OAI21X1_334 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n1378_), .C(_abc_40319_new_n1875_), .Y(_abc_40319_new_n1986_));
OAI21X1 OAI21X1_335 ( .A(_abc_40319_new_n580_), .B(_abc_40319_new_n1401_), .C(_abc_40319_new_n1986_), .Y(_abc_40319_new_n1987_));
OAI21X1 OAI21X1_336 ( .A(_abc_40319_new_n1258_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1998_), .Y(_abc_40319_new_n1999_));
OAI21X1 OAI21X1_337 ( .A(_abc_40319_new_n1996_), .B(_abc_40319_new_n1997_), .C(_abc_40319_new_n2001_), .Y(_abc_40319_new_n2002_));
OAI21X1 OAI21X1_338 ( .A(_abc_40319_new_n2004_), .B(_abc_40319_new_n1993_), .C(_abc_40319_new_n2009_), .Y(_abc_40319_new_n2010_));
OAI21X1 OAI21X1_339 ( .A(_abc_40319_new_n580_), .B(_abc_40319_new_n1516_), .C(_abc_40319_new_n2011_), .Y(_abc_40319_new_n2012_));
OAI21X1 OAI21X1_34 ( .A(_abc_40319_new_n758_), .B(_abc_40319_new_n759_), .C(_abc_40319_new_n752_), .Y(_abc_40319_new_n760_));
OAI21X1 OAI21X1_340 ( .A(_abc_40319_new_n2007_), .B(_abc_40319_new_n2008_), .C(_abc_40319_new_n2014_), .Y(_abc_40319_new_n2015_));
OAI21X1 OAI21X1_341 ( .A(_abc_40319_new_n1888_), .B(_abc_40319_new_n1208_), .C(_abc_40319_new_n2017_), .Y(_abc_40319_new_n2018_));
OAI21X1 OAI21X1_342 ( .A(_abc_40319_new_n2025_), .B(_abc_40319_new_n2024_), .C(_abc_40319_new_n2022_), .Y(_abc_40319_new_n2026_));
OAI21X1 OAI21X1_343 ( .A(_abc_40319_new_n1150_), .B(_abc_40319_new_n1155_), .C(_abc_40319_new_n1870_), .Y(_abc_40319_new_n2027_));
OAI21X1 OAI21X1_344 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n663_), .C(_abc_40319_new_n1429_), .Y(_abc_40319_new_n2028_));
OAI21X1 OAI21X1_345 ( .A(_abc_40319_new_n1431_), .B(_abc_40319_new_n1436_), .C(_abc_40319_new_n1875_), .Y(_abc_40319_new_n2029_));
OAI21X1 OAI21X1_346 ( .A(_abc_40319_new_n2026_), .B(_abc_40319_new_n2021_), .C(_abc_40319_new_n2033_), .Y(_abc_40319_new_n2034_));
OAI21X1 OAI21X1_347 ( .A(_abc_40319_new_n1567_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n2036_), .Y(_abc_40319_new_n2037_));
OAI21X1 OAI21X1_348 ( .A(_abc_40319_new_n1888_), .B(_abc_40319_new_n1760_), .C(_abc_40319_new_n2040_), .Y(_abc_40319_new_n2041_));
OAI21X1 OAI21X1_349 ( .A(_abc_40319_new_n2048_), .B(_abc_40319_new_n2047_), .C(_abc_40319_new_n2045_), .Y(_abc_40319_new_n2049_));
OAI21X1 OAI21X1_35 ( .A(IR_REG_4_), .B(_abc_40319_new_n763_), .C(IR_REG_5_), .Y(_abc_40319_new_n764_));
OAI21X1 OAI21X1_350 ( .A(_abc_40319_new_n1888_), .B(_abc_40319_new_n1710_), .C(_abc_40319_new_n2050_), .Y(_abc_40319_new_n2051_));
OAI21X1 OAI21X1_351 ( .A(_abc_40319_new_n2049_), .B(_abc_40319_new_n2044_), .C(_abc_40319_new_n2054_), .Y(_abc_40319_new_n2055_));
OAI21X1 OAI21X1_352 ( .A(_abc_40319_new_n1888_), .B(_abc_40319_new_n1093_), .C(_abc_40319_new_n2056_), .Y(_abc_40319_new_n2057_));
OAI21X1 OAI21X1_353 ( .A(_abc_40319_new_n2052_), .B(_abc_40319_new_n2053_), .C(_abc_40319_new_n2060_), .Y(_abc_40319_new_n2061_));
OAI21X1 OAI21X1_354 ( .A(_abc_40319_new_n1888_), .B(_abc_40319_new_n1078_), .C(_abc_40319_new_n2063_), .Y(_abc_40319_new_n2064_));
OAI21X1 OAI21X1_355 ( .A(_abc_40319_new_n1888_), .B(_abc_40319_new_n1496_), .C(_abc_40319_new_n2068_), .Y(_abc_40319_new_n2069_));
OAI21X1 OAI21X1_356 ( .A(_abc_40319_new_n2073_), .B(_abc_40319_new_n2067_), .C(_abc_40319_new_n2078_), .Y(_abc_40319_new_n2079_));
OAI21X1 OAI21X1_357 ( .A(_abc_40319_new_n1888_), .B(_abc_40319_new_n1505_), .C(_abc_40319_new_n2080_), .Y(_abc_40319_new_n2081_));
OAI21X1 OAI21X1_358 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_29_), .Y(_abc_40319_new_n2088_));
OAI21X1 OAI21X1_359 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_30_), .Y(_abc_40319_new_n2096_));
OAI21X1 OAI21X1_36 ( .A(_abc_40319_new_n546_), .B(_abc_40319_new_n549_), .C(_abc_40319_new_n764_), .Y(_abc_40319_new_n765_));
OAI21X1 OAI21X1_360 ( .A(_abc_40319_new_n2099_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n2100_), .Y(_abc_40319_new_n2101_));
OAI21X1 OAI21X1_361 ( .A(_abc_40319_new_n2098_), .B(_abc_40319_new_n2101_), .C(_abc_40319_new_n1883_), .Y(_abc_40319_new_n2106_));
OAI21X1 OAI21X1_362 ( .A(_abc_40319_new_n992_), .B(_abc_40319_new_n2106_), .C(_abc_40319_new_n2107_), .Y(_abc_40319_new_n2108_));
OAI21X1 OAI21X1_363 ( .A(_abc_40319_new_n2113_), .B(_abc_40319_new_n2112_), .C(_abc_40319_new_n1887_), .Y(_abc_40319_new_n2114_));
OAI21X1 OAI21X1_364 ( .A(_abc_40319_new_n1504_), .B(_abc_40319_new_n1499_), .C(_abc_40319_new_n1581_), .Y(_abc_40319_new_n2118_));
OAI21X1 OAI21X1_365 ( .A(_abc_40319_new_n2122_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n1065_), .Y(_abc_40319_new_n2123_));
OAI21X1 OAI21X1_366 ( .A(_abc_40319_new_n2126_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n1077_), .Y(_abc_40319_new_n2127_));
OAI21X1 OAI21X1_367 ( .A(_abc_40319_new_n2136_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n1115_), .Y(_abc_40319_new_n2137_));
OAI21X1 OAI21X1_368 ( .A(_abc_40319_new_n1468_), .B(_abc_40319_new_n1464_), .C(_abc_40319_new_n1459_), .Y(_abc_40319_new_n2140_));
OAI21X1 OAI21X1_369 ( .A(_abc_40319_new_n1878_), .B(_abc_40319_new_n1881_), .C(_abc_40319_new_n1876_), .Y(_abc_40319_new_n2145_));
OAI21X1 OAI21X1_37 ( .A(IR_REG_31_), .B(IR_REG_5_), .C(_abc_40319_new_n766_), .Y(_abc_40319_new_n767_));
OAI21X1 OAI21X1_370 ( .A(_abc_40319_new_n2098_), .B(_abc_40319_new_n2101_), .C(_abc_40319_new_n2096_), .Y(_abc_40319_new_n2149_));
OAI21X1 OAI21X1_371 ( .A(_abc_40319_new_n829_), .B(_abc_40319_new_n861_), .C(_abc_40319_new_n825_), .Y(_abc_40319_new_n2154_));
OAI21X1 OAI21X1_372 ( .A(_abc_40319_new_n1201_), .B(_abc_40319_new_n1207_), .C(_abc_40319_new_n1211_), .Y(_abc_40319_new_n2156_));
OAI21X1 OAI21X1_373 ( .A(_abc_40319_new_n1150_), .B(_abc_40319_new_n1155_), .C(_abc_40319_new_n1159_), .Y(_abc_40319_new_n2161_));
OAI21X1 OAI21X1_374 ( .A(_abc_40319_new_n1431_), .B(_abc_40319_new_n1436_), .C(_abc_40319_new_n1570_), .Y(_abc_40319_new_n2166_));
OAI21X1 OAI21X1_375 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n1378_), .C(_abc_40319_new_n1370_), .Y(_abc_40319_new_n2177_));
OAI21X1 OAI21X1_376 ( .A(_abc_40319_new_n1304_), .B(_abc_40319_new_n1307_), .C(_abc_40319_new_n1297_), .Y(_abc_40319_new_n2183_));
OAI21X1 OAI21X1_377 ( .A(_abc_40319_new_n754_), .B(_abc_40319_new_n753_), .C(_abc_40319_new_n698_), .Y(_abc_40319_new_n2189_));
OAI21X1 OAI21X1_378 ( .A(_abc_40319_new_n1957_), .B(_abc_40319_new_n1958_), .C(_abc_40319_new_n1276_), .Y(_abc_40319_new_n2192_));
OAI21X1 OAI21X1_379 ( .A(_abc_40319_new_n1178_), .B(_abc_40319_new_n1188_), .C(_abc_40319_new_n1175_), .Y(_abc_40319_new_n2198_));
OAI21X1 OAI21X1_38 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_5_), .Y(_abc_40319_new_n768_));
OAI21X1 OAI21X1_380 ( .A(_abc_40319_new_n1355_), .B(_abc_40319_new_n1359_), .C(_abc_40319_new_n1654_), .Y(_abc_40319_new_n2201_));
OAI21X1 OAI21X1_381 ( .A(_abc_40319_new_n2213_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n1137_), .Y(_abc_40319_new_n2214_));
OAI21X1 OAI21X1_382 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1129_), .C(_abc_40319_new_n1123_), .Y(_abc_40319_new_n2215_));
OAI21X1 OAI21X1_383 ( .A(_abc_40319_new_n1451_), .B(_abc_40319_new_n1447_), .C(_abc_40319_new_n1442_), .Y(_abc_40319_new_n2217_));
OAI21X1 OAI21X1_384 ( .A(_abc_40319_new_n1226_), .B(_abc_40319_new_n1232_), .C(_abc_40319_new_n1865_), .Y(_abc_40319_new_n2221_));
OAI21X1 OAI21X1_385 ( .A(_abc_40319_new_n1251_), .B(_abc_40319_new_n1257_), .C(_abc_40319_new_n1248_), .Y(_abc_40319_new_n2239_));
OAI21X1 OAI21X1_386 ( .A(_abc_40319_new_n849_), .B(_abc_40319_new_n846_), .C(_abc_40319_new_n853_), .Y(_abc_40319_new_n2243_));
OAI21X1 OAI21X1_387 ( .A(_abc_40319_new_n953_), .B(_abc_40319_new_n950_), .C(_abc_40319_new_n2246_), .Y(_abc_40319_new_n2247_));
OAI21X1 OAI21X1_388 ( .A(_abc_40319_new_n2258_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n1046_), .Y(_abc_40319_new_n2259_));
OAI21X1 OAI21X1_389 ( .A(_abc_40319_new_n2273_), .B(_abc_40319_new_n2278_), .C(_abc_40319_new_n2281_), .Y(_abc_40319_new_n2282_));
OAI21X1 OAI21X1_39 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n767_), .C(_abc_40319_new_n768_), .Y(_abc_40319_new_n769_));
OAI21X1 OAI21X1_390 ( .A(_abc_40319_new_n1992_), .B(_abc_40319_new_n2291_), .C(_abc_40319_new_n2003_), .Y(_abc_40319_new_n2292_));
OAI21X1 OAI21X1_391 ( .A(_abc_40319_new_n2020_), .B(_abc_40319_new_n2293_), .C(_abc_40319_new_n2294_), .Y(_abc_40319_new_n2295_));
OAI21X1 OAI21X1_392 ( .A(_abc_40319_new_n2043_), .B(_abc_40319_new_n2297_), .C(_abc_40319_new_n2298_), .Y(_abc_40319_new_n2299_));
OAI21X1 OAI21X1_393 ( .A(_abc_40319_new_n2066_), .B(_abc_40319_new_n2300_), .C(_abc_40319_new_n2072_), .Y(_abc_40319_new_n2301_));
OAI21X1 OAI21X1_394 ( .A(_abc_40319_new_n2303_), .B(_abc_40319_new_n2302_), .C(_abc_40319_new_n2110_), .Y(_abc_40319_new_n2304_));
OAI21X1 OAI21X1_395 ( .A(_abc_40319_new_n1443_), .B(_abc_40319_new_n1567_), .C(_abc_40319_new_n2140_), .Y(_abc_40319_new_n2319_));
OAI21X1 OAI21X1_396 ( .A(_abc_40319_new_n1148_), .B(_abc_40319_new_n1156_), .C(_abc_40319_new_n2166_), .Y(_abc_40319_new_n2321_));
OAI21X1 OAI21X1_397 ( .A(_abc_40319_new_n1178_), .B(_abc_40319_new_n1188_), .C(_abc_40319_new_n2196_), .Y(_abc_40319_new_n2322_));
OAI21X1 OAI21X1_398 ( .A(_abc_40319_new_n2156_), .B(_abc_40319_new_n2162_), .C(_abc_40319_new_n2322_), .Y(_abc_40319_new_n2323_));
OAI21X1 OAI21X1_399 ( .A(_abc_40319_new_n2223_), .B(_abc_40319_new_n2324_), .C(_abc_40319_new_n2168_), .Y(_abc_40319_new_n2325_));
OAI21X1 OAI21X1_4 ( .A(IR_REG_31_), .B(IR_REG_25_), .C(_abc_40319_new_n566_), .Y(_abc_40319_new_n567_));
OAI21X1 OAI21X1_40 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n772_), .C(_abc_40319_new_n709_), .Y(_abc_40319_new_n773_));
OAI21X1 OAI21X1_400 ( .A(_abc_40319_new_n1332_), .B(_abc_40319_new_n1335_), .C(_abc_40319_new_n2228_), .Y(_abc_40319_new_n2327_));
OAI21X1 OAI21X1_401 ( .A(_abc_40319_new_n1796_), .B(_abc_40319_new_n1352_), .C(_abc_40319_new_n2327_), .Y(_abc_40319_new_n2328_));
OAI21X1 OAI21X1_402 ( .A(_abc_40319_new_n1251_), .B(_abc_40319_new_n1257_), .C(_abc_40319_new_n1261_), .Y(_abc_40319_new_n2331_));
OAI21X1 OAI21X1_403 ( .A(_abc_40319_new_n1396_), .B(_abc_40319_new_n1400_), .C(_abc_40319_new_n1541_), .Y(_abc_40319_new_n2336_));
OAI21X1 OAI21X1_404 ( .A(_abc_40319_new_n2177_), .B(_abc_40319_new_n2202_), .C(_abc_40319_new_n2336_), .Y(_abc_40319_new_n2337_));
OAI21X1 OAI21X1_405 ( .A(_abc_40319_new_n1304_), .B(_abc_40319_new_n1307_), .C(_abc_40319_new_n1739_), .Y(_abc_40319_new_n2338_));
OAI21X1 OAI21X1_406 ( .A(_abc_40319_new_n988_), .B(_abc_40319_new_n1276_), .C(_abc_40319_new_n2338_), .Y(_abc_40319_new_n2339_));
OAI21X1 OAI21X1_407 ( .A(_abc_40319_new_n698_), .B(_abc_40319_new_n759_), .C(_abc_40319_new_n2340_), .Y(_abc_40319_new_n2341_));
OAI21X1 OAI21X1_408 ( .A(_abc_40319_new_n2248_), .B(_abc_40319_new_n2343_), .C(_abc_40319_new_n2326_), .Y(_abc_40319_new_n2344_));
OAI21X1 OAI21X1_409 ( .A(_abc_40319_new_n2132_), .B(_abc_40319_new_n2137_), .C(_abc_40319_new_n2315_), .Y(_abc_40319_new_n2347_));
OAI21X1 OAI21X1_41 ( .A(_abc_40319_new_n770_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n771_), .Y(_abc_40319_new_n775_));
OAI21X1 OAI21X1_410 ( .A(_abc_40319_new_n944_), .B(_abc_40319_new_n959_), .C(_abc_40319_new_n2342_), .Y(_abc_40319_new_n2349_));
OAI21X1 OAI21X1_411 ( .A(_abc_40319_new_n1108_), .B(_abc_40319_new_n1115_), .C(_abc_40319_new_n2131_), .Y(_abc_40319_new_n2354_));
OAI21X1 OAI21X1_412 ( .A(_abc_40319_new_n2353_), .B(_abc_40319_new_n2354_), .C(_abc_40319_new_n2335_), .Y(_abc_40319_new_n2355_));
OAI21X1 OAI21X1_413 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n855_), .C(_abc_40319_new_n2154_), .Y(_abc_40319_new_n2358_));
OAI21X1 OAI21X1_414 ( .A(_abc_40319_new_n1123_), .B(_abc_40319_new_n1137_), .C(_abc_40319_new_n2335_), .Y(_abc_40319_new_n2366_));
OAI21X1 OAI21X1_415 ( .A(_abc_40319_new_n1325_), .B(_abc_40319_new_n1514_), .C(_abc_40319_new_n2202_), .Y(_abc_40319_new_n2374_));
OAI21X1 OAI21X1_416 ( .A(_abc_40319_new_n2156_), .B(_abc_40319_new_n2162_), .C(_abc_40319_new_n2381_), .Y(_abc_40319_new_n2382_));
OAI21X1 OAI21X1_417 ( .A(_abc_40319_new_n2321_), .B(_abc_40319_new_n2382_), .C(_abc_40319_new_n2380_), .Y(_abc_40319_new_n2383_));
OAI21X1 OAI21X1_418 ( .A(_abc_40319_new_n1054_), .B(_abc_40319_new_n1065_), .C(_abc_40319_new_n2128_), .Y(_abc_40319_new_n2393_));
OAI21X1 OAI21X1_419 ( .A(_abc_40319_new_n2177_), .B(_abc_40319_new_n2202_), .C(_abc_40319_new_n2394_), .Y(_abc_40319_new_n2395_));
OAI21X1 OAI21X1_42 ( .A(_abc_40319_new_n729_), .B(_abc_40319_new_n730_), .C(_abc_40319_new_n779_), .Y(_abc_40319_new_n780_));
OAI21X1 OAI21X1_420 ( .A(_abc_40319_new_n1159_), .B(_abc_40319_new_n1157_), .C(_abc_40319_new_n2157_), .Y(_abc_40319_new_n2408_));
OAI21X1 OAI21X1_421 ( .A(_abc_40319_new_n2319_), .B(_abc_40319_new_n2409_), .C(_abc_40319_new_n2406_), .Y(_abc_40319_new_n2410_));
OAI21X1 OAI21X1_422 ( .A(_abc_40319_new_n2354_), .B(_abc_40319_new_n2410_), .C(_abc_40319_new_n2259_), .Y(_abc_40319_new_n2411_));
OAI21X1 OAI21X1_423 ( .A(_abc_40319_new_n2411_), .B(_abc_40319_new_n2317_), .C(_abc_40319_new_n2404_), .Y(_abc_40319_new_n2412_));
OAI21X1 OAI21X1_424 ( .A(_abc_40319_new_n2403_), .B(_abc_40319_new_n2413_), .C(_abc_40319_new_n2402_), .Y(_abc_40319_new_n2414_));
OAI21X1 OAI21X1_425 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n1883_), .C(_abc_40319_new_n2414_), .Y(_abc_40319_new_n2415_));
OAI21X1 OAI21X1_426 ( .A(_abc_40319_new_n799_), .B(_abc_40319_new_n1556_), .C(_abc_40319_new_n2118_), .Y(_abc_40319_new_n2417_));
OAI21X1 OAI21X1_427 ( .A(_abc_40319_new_n2416_), .B(_abc_40319_new_n2419_), .C(_abc_40319_new_n2357_), .Y(_abc_40319_new_n2420_));
OAI21X1 OAI21X1_428 ( .A(_abc_40319_new_n616_), .B(_abc_40319_new_n2306_), .C(_abc_40319_new_n2440_), .Y(_abc_40319_new_n2441_));
OAI21X1 OAI21X1_429 ( .A(_abc_40319_new_n749_), .B(_abc_40319_new_n1874_), .C(_abc_40319_new_n2447_), .Y(_abc_40319_new_n2448_));
OAI21X1 OAI21X1_43 ( .A(_abc_40319_new_n751_), .B(_abc_40319_new_n746_), .C(_abc_40319_new_n769_), .Y(_abc_40319_new_n785_));
OAI21X1 OAI21X1_430 ( .A(_abc_40319_new_n1055_), .B(_abc_40319_new_n1496_), .C(_abc_40319_new_n2259_), .Y(_abc_40319_new_n2453_));
OAI21X1 OAI21X1_431 ( .A(_abc_40319_new_n2166_), .B(_abc_40319_new_n2219_), .C(_abc_40319_new_n2217_), .Y(_abc_40319_new_n2458_));
OAI21X1 OAI21X1_432 ( .A(_abc_40319_new_n1122_), .B(_abc_40319_new_n1135_), .C(_abc_40319_new_n2141_), .Y(_abc_40319_new_n2460_));
OAI21X1 OAI21X1_433 ( .A(_abc_40319_new_n1108_), .B(_abc_40319_new_n1115_), .C(_abc_40319_new_n2461_), .Y(_abc_40319_new_n2462_));
OAI21X1 OAI21X1_434 ( .A(_abc_40319_new_n2132_), .B(_abc_40319_new_n2462_), .C(_abc_40319_new_n2456_), .Y(_abc_40319_new_n2463_));
OAI21X1 OAI21X1_435 ( .A(_abc_40319_new_n987_), .B(_abc_40319_new_n2427_), .C(_abc_40319_new_n2390_), .Y(_abc_40319_new_n2465_));
OAI21X1 OAI21X1_436 ( .A(_abc_40319_new_n877_), .B(_abc_40319_new_n897_), .C(_abc_40319_new_n1906_), .Y(_abc_40319_new_n2468_));
OAI21X1 OAI21X1_437 ( .A(_abc_40319_new_n853_), .B(_abc_40319_new_n842_), .C(_abc_40319_new_n2468_), .Y(_abc_40319_new_n2469_));
OAI21X1 OAI21X1_438 ( .A(_abc_40319_new_n2152_), .B(_abc_40319_new_n2470_), .C(_abc_40319_new_n2154_), .Y(_abc_40319_new_n2471_));
OAI21X1 OAI21X1_439 ( .A(_abc_40319_new_n1726_), .B(_abc_40319_new_n809_), .C(_abc_40319_new_n2472_), .Y(_abc_40319_new_n2473_));
OAI21X1 OAI21X1_44 ( .A(_abc_40319_new_n775_), .B(_abc_40319_new_n782_), .C(_abc_40319_new_n679_), .Y(_abc_40319_new_n786_));
OAI21X1 OAI21X1_440 ( .A(_abc_40319_new_n2173_), .B(_abc_40319_new_n2232_), .C(_abc_40319_new_n2472_), .Y(_abc_40319_new_n2475_));
OAI21X1 OAI21X1_441 ( .A(_abc_40319_new_n944_), .B(_abc_40319_new_n959_), .C(_abc_40319_new_n2475_), .Y(_abc_40319_new_n2476_));
OAI21X1 OAI21X1_442 ( .A(_abc_40319_new_n698_), .B(_abc_40319_new_n759_), .C(_abc_40319_new_n2477_), .Y(_abc_40319_new_n2478_));
OAI21X1 OAI21X1_443 ( .A(_abc_40319_new_n1393_), .B(_abc_40319_new_n1401_), .C(_abc_40319_new_n2177_), .Y(_abc_40319_new_n2480_));
OAI21X1 OAI21X1_444 ( .A(_abc_40319_new_n2340_), .B(_abc_40319_new_n2466_), .C(_abc_40319_new_n2481_), .Y(_abc_40319_new_n2482_));
OAI21X1 OAI21X1_445 ( .A(_abc_40319_new_n1261_), .B(_abc_40319_new_n1259_), .C(_abc_40319_new_n2485_), .Y(_abc_40319_new_n2486_));
OAI21X1 OAI21X1_446 ( .A(_abc_40319_new_n2479_), .B(_abc_40319_new_n2482_), .C(_abc_40319_new_n2489_), .Y(_abc_40319_new_n2490_));
OAI21X1 OAI21X1_447 ( .A(_abc_40319_new_n2381_), .B(_abc_40319_new_n2493_), .C(_abc_40319_new_n2492_), .Y(_abc_40319_new_n2494_));
OAI21X1 OAI21X1_448 ( .A(_abc_40319_new_n1198_), .B(_abc_40319_new_n1208_), .C(_abc_40319_new_n2495_), .Y(_abc_40319_new_n2496_));
OAI21X1 OAI21X1_449 ( .A(_abc_40319_new_n2408_), .B(_abc_40319_new_n2497_), .C(_abc_40319_new_n2161_), .Y(_abc_40319_new_n2498_));
OAI21X1 OAI21X1_45 ( .A(_abc_40319_new_n758_), .B(_abc_40319_new_n788_), .C(_abc_40319_new_n785_), .Y(_abc_40319_new_n789_));
OAI21X1 OAI21X1_450 ( .A(_abc_40319_new_n1108_), .B(_abc_40319_new_n1115_), .C(_abc_40319_new_n2500_), .Y(_abc_40319_new_n2501_));
OAI21X1 OAI21X1_451 ( .A(_abc_40319_new_n2088_), .B(_abc_40319_new_n2264_), .C(_abc_40319_new_n2507_), .Y(_abc_40319_new_n2508_));
OAI21X1 OAI21X1_452 ( .A(_abc_40319_new_n2453_), .B(_abc_40319_new_n2505_), .C(_abc_40319_new_n2509_), .Y(_abc_40319_new_n2510_));
OAI21X1 OAI21X1_453 ( .A(_abc_40319_new_n2118_), .B(_abc_40319_new_n2508_), .C(_abc_40319_new_n2511_), .Y(_abc_40319_new_n2512_));
OAI21X1 OAI21X1_454 ( .A(_abc_40319_new_n1007_), .B(_abc_40319_new_n2114_), .C(_abc_40319_new_n2520_), .Y(_abc_40319_new_n2521_));
OAI21X1 OAI21X1_455 ( .A(_abc_40319_new_n2525_), .B(_abc_40319_new_n975_), .C(_abc_40319_new_n1870_), .Y(_abc_40319_new_n2526_));
OAI21X1 OAI21X1_456 ( .A(_abc_40319_new_n1872_), .B(_abc_40319_new_n2522_), .C(_abc_40319_new_n2529_), .Y(n1186));
OAI21X1 OAI21X1_457 ( .A(_abc_40319_new_n593_), .B(_abc_40319_new_n602_), .C(IR_REG_0_), .Y(_abc_40319_new_n2534_));
OAI21X1 OAI21X1_458 ( .A(_abc_40319_new_n871_), .B(_abc_40319_new_n907_), .C(_abc_40319_new_n2524_), .Y(_abc_40319_new_n2535_));
OAI21X1 OAI21X1_459 ( .A(_abc_40319_new_n1871_), .B(_abc_40319_new_n674_), .C(n1341), .Y(_abc_40319_new_n2538_));
OAI21X1 OAI21X1_46 ( .A(IR_REG_31_), .B(_abc_40319_new_n548_), .C(_abc_40319_new_n795_), .Y(_abc_40319_new_n796_));
OAI21X1 OAI21X1_460 ( .A(_abc_40319_new_n2537_), .B(_abc_40319_new_n2538_), .C(_abc_40319_new_n2540_), .Y(n1054));
OAI21X1 OAI21X1_461 ( .A(_abc_40319_new_n871_), .B(_abc_40319_new_n909_), .C(_abc_40319_new_n883_), .Y(_abc_40319_new_n2551_));
OAI21X1 OAI21X1_462 ( .A(_abc_40319_new_n2549_), .B(_abc_40319_new_n2525_), .C(_abc_40319_new_n2554_), .Y(_abc_40319_new_n2555_));
OAI21X1 OAI21X1_463 ( .A(_abc_40319_new_n2542_), .B(_abc_40319_new_n2543_), .C(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2556_));
OAI21X1 OAI21X1_464 ( .A(_abc_40319_new_n586_), .B(_abc_40319_new_n592_), .C(_abc_40319_new_n696_), .Y(_abc_40319_new_n2559_));
OAI21X1 OAI21X1_465 ( .A(_abc_40319_new_n2536_), .B(_abc_40319_new_n2560_), .C(n1345), .Y(_abc_40319_new_n2561_));
OAI21X1 OAI21X1_466 ( .A(REG2_REG_2_), .B(_abc_40319_new_n836_), .C(_abc_40319_new_n2564_), .Y(_abc_40319_new_n2577_));
OAI21X1 OAI21X1_467 ( .A(_abc_40319_new_n847_), .B(_abc_40319_new_n837_), .C(_abc_40319_new_n2577_), .Y(_abc_40319_new_n2578_));
OAI21X1 OAI21X1_468 ( .A(_abc_40319_new_n2567_), .B(_abc_40319_new_n2572_), .C(_abc_40319_new_n2569_), .Y(_abc_40319_new_n2581_));
OAI21X1 OAI21X1_469 ( .A(_abc_40319_new_n2585_), .B(_abc_40319_new_n2587_), .C(_abc_40319_new_n2523_), .Y(_abc_40319_new_n2588_));
OAI21X1 OAI21X1_47 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_4_), .Y(_abc_40319_new_n798_));
OAI21X1 OAI21X1_470 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n821_), .C(_abc_40319_new_n2588_), .Y(_abc_40319_new_n2589_));
OAI21X1 OAI21X1_471 ( .A(_abc_40319_new_n2590_), .B(_abc_40319_new_n2538_), .C(_abc_40319_new_n2591_), .Y(n1042));
OAI21X1 OAI21X1_472 ( .A(REG2_REG_3_), .B(_abc_40319_new_n822_), .C(_abc_40319_new_n2578_), .Y(_abc_40319_new_n2596_));
OAI21X1 OAI21X1_473 ( .A(_abc_40319_new_n827_), .B(_abc_40319_new_n821_), .C(_abc_40319_new_n2596_), .Y(_abc_40319_new_n2597_));
OAI21X1 OAI21X1_474 ( .A(_abc_40319_new_n821_), .B(_abc_40319_new_n2582_), .C(_abc_40319_new_n2584_), .Y(_abc_40319_new_n2599_));
OAI21X1 OAI21X1_475 ( .A(_abc_40319_new_n2525_), .B(_abc_40319_new_n2598_), .C(_abc_40319_new_n2602_), .Y(_abc_40319_new_n2603_));
OAI21X1 OAI21X1_476 ( .A(REG2_REG_4_), .B(_abc_40319_new_n796_), .C(_abc_40319_new_n2597_), .Y(_abc_40319_new_n2607_));
OAI21X1 OAI21X1_477 ( .A(REG1_REG_4_), .B(_abc_40319_new_n796_), .C(_abc_40319_new_n2599_), .Y(_abc_40319_new_n2611_));
OAI21X1 OAI21X1_478 ( .A(_abc_40319_new_n800_), .B(_abc_40319_new_n797_), .C(_abc_40319_new_n2611_), .Y(_abc_40319_new_n2612_));
OAI21X1 OAI21X1_479 ( .A(_abc_40319_new_n767_), .B(_abc_40319_new_n2616_), .C(_abc_40319_new_n2617_), .Y(_abc_40319_new_n2618_));
OAI21X1 OAI21X1_48 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n797_), .C(_abc_40319_new_n798_), .Y(_abc_40319_new_n799_));
OAI21X1 OAI21X1_480 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n767_), .C(_abc_40319_new_n2618_), .Y(_abc_40319_new_n2619_));
OAI21X1 OAI21X1_481 ( .A(_abc_40319_new_n2538_), .B(_abc_40319_new_n2620_), .C(_abc_40319_new_n2621_), .Y(n1034));
OAI21X1 OAI21X1_482 ( .A(_abc_40319_new_n767_), .B(_abc_40319_new_n2614_), .C(_abc_40319_new_n2613_), .Y(_abc_40319_new_n2624_));
OAI21X1 OAI21X1_483 ( .A(_abc_40319_new_n2625_), .B(_abc_40319_new_n2624_), .C(_abc_40319_new_n2523_), .Y(_abc_40319_new_n2626_));
OAI21X1 OAI21X1_484 ( .A(_abc_40319_new_n770_), .B(_abc_40319_new_n767_), .C(_abc_40319_new_n2608_), .Y(_abc_40319_new_n2629_));
OAI21X1 OAI21X1_485 ( .A(_abc_40319_new_n2631_), .B(_abc_40319_new_n2632_), .C(_abc_40319_new_n2633_), .Y(_abc_40319_new_n2634_));
OAI21X1 OAI21X1_486 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n942_), .C(_abc_40319_new_n2634_), .Y(_abc_40319_new_n2635_));
OAI21X1 OAI21X1_487 ( .A(_abc_40319_new_n2627_), .B(_abc_40319_new_n2635_), .C(_abc_40319_new_n2623_), .Y(_abc_40319_new_n2636_));
OAI21X1 OAI21X1_488 ( .A(REG2_REG_6_), .B(_abc_40319_new_n2642_), .C(_abc_40319_new_n2630_), .Y(_abc_40319_new_n2643_));
OAI21X1 OAI21X1_489 ( .A(_abc_40319_new_n951_), .B(_abc_40319_new_n942_), .C(_abc_40319_new_n2643_), .Y(_abc_40319_new_n2644_));
OAI21X1 OAI21X1_49 ( .A(_abc_40319_new_n804_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n807_), .Y(_abc_40319_new_n808_));
OAI21X1 OAI21X1_490 ( .A(REG2_REG_7_), .B(_abc_40319_new_n690_), .C(_abc_40319_new_n2644_), .Y(_abc_40319_new_n2647_));
OAI21X1 OAI21X1_491 ( .A(_abc_40319_new_n2640_), .B(_abc_40319_new_n2647_), .C(_abc_40319_new_n2524_), .Y(_abc_40319_new_n2648_));
OAI21X1 OAI21X1_492 ( .A(REG1_REG_6_), .B(_abc_40319_new_n2642_), .C(_abc_40319_new_n2624_), .Y(_abc_40319_new_n2650_));
OAI21X1 OAI21X1_493 ( .A(_abc_40319_new_n945_), .B(_abc_40319_new_n942_), .C(_abc_40319_new_n2650_), .Y(_abc_40319_new_n2651_));
OAI21X1 OAI21X1_494 ( .A(_abc_40319_new_n2657_), .B(_abc_40319_new_n2656_), .C(_abc_40319_new_n2523_), .Y(_abc_40319_new_n2658_));
OAI21X1 OAI21X1_495 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n691_), .C(_abc_40319_new_n2658_), .Y(_abc_40319_new_n2659_));
OAI21X1 OAI21X1_496 ( .A(_abc_40319_new_n2659_), .B(_abc_40319_new_n2649_), .C(_abc_40319_new_n2623_), .Y(_abc_40319_new_n2660_));
OAI21X1 OAI21X1_497 ( .A(_abc_40319_new_n2639_), .B(_abc_40319_new_n691_), .C(_abc_40319_new_n2647_), .Y(_abc_40319_new_n2665_));
OAI21X1 OAI21X1_498 ( .A(REG2_REG_8_), .B(_abc_40319_new_n1273_), .C(_abc_40319_new_n2665_), .Y(_abc_40319_new_n2666_));
OAI21X1 OAI21X1_499 ( .A(_abc_40319_new_n2664_), .B(_abc_40319_new_n2668_), .C(_abc_40319_new_n2667_), .Y(_abc_40319_new_n2669_));
OAI21X1 OAI21X1_5 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n569_), .C(_abc_40319_new_n570_), .Y(_abc_40319_new_n571_));
OAI21X1 OAI21X1_50 ( .A(_abc_40319_new_n671_), .B(_abc_40319_new_n681_), .C(_abc_40319_new_n812_), .Y(_abc_40319_new_n813_));
OAI21X1 OAI21X1_500 ( .A(_abc_40319_new_n2664_), .B(_abc_40319_new_n2666_), .C(_abc_40319_new_n2669_), .Y(_abc_40319_new_n2670_));
OAI21X1 OAI21X1_501 ( .A(REG1_REG_7_), .B(_abc_40319_new_n690_), .C(_abc_40319_new_n2674_), .Y(_abc_40319_new_n2675_));
OAI21X1 OAI21X1_502 ( .A(_abc_40319_new_n586_), .B(_abc_40319_new_n592_), .C(_abc_40319_new_n2679_), .Y(_abc_40319_new_n2680_));
OAI21X1 OAI21X1_503 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n1274_), .C(_abc_40319_new_n2680_), .Y(_abc_40319_new_n2681_));
OAI21X1 OAI21X1_504 ( .A(_abc_40319_new_n2671_), .B(_abc_40319_new_n2681_), .C(_abc_40319_new_n2543_), .Y(_abc_40319_new_n2682_));
OAI21X1 OAI21X1_505 ( .A(_abc_40319_new_n593_), .B(_abc_40319_new_n602_), .C(_abc_40319_new_n2542_), .Y(_abc_40319_new_n2683_));
OAI21X1 OAI21X1_506 ( .A(_abc_40319_new_n2689_), .B(_abc_40319_new_n2670_), .C(_abc_40319_new_n2690_), .Y(_abc_40319_new_n2691_));
OAI21X1 OAI21X1_507 ( .A(_abc_40319_new_n593_), .B(_abc_40319_new_n602_), .C(_abc_40319_new_n1294_), .Y(_abc_40319_new_n2709_));
OAI21X1 OAI21X1_508 ( .A(_abc_40319_new_n2709_), .B(_abc_40319_new_n2686_), .C(_abc_40319_new_n2708_), .Y(_abc_40319_new_n2710_));
OAI21X1 OAI21X1_509 ( .A(_abc_40319_new_n2709_), .B(_abc_40319_new_n2711_), .C(_abc_40319_new_n1741_), .Y(_abc_40319_new_n2712_));
OAI21X1 OAI21X1_51 ( .A(IR_REG_31_), .B(IR_REG_3_), .C(_abc_40319_new_n820_), .Y(_abc_40319_new_n821_));
OAI21X1 OAI21X1_510 ( .A(_abc_40319_new_n2538_), .B(_abc_40319_new_n2707_), .C(_abc_40319_new_n2713_), .Y(n1018));
OAI21X1 OAI21X1_511 ( .A(_abc_40319_new_n1298_), .B(_abc_40319_new_n1295_), .C(_abc_40319_new_n2715_), .Y(_abc_40319_new_n2716_));
OAI21X1 OAI21X1_512 ( .A(_abc_40319_new_n1391_), .B(_abc_40319_new_n2683_), .C(_abc_40319_new_n1542_), .Y(_abc_40319_new_n2722_));
OAI21X1 OAI21X1_513 ( .A(_abc_40319_new_n2727_), .B(_abc_40319_new_n2698_), .C(_abc_40319_new_n2694_), .Y(_abc_40319_new_n2728_));
OAI21X1 OAI21X1_514 ( .A(_abc_40319_new_n2542_), .B(_abc_40319_new_n2543_), .C(_abc_40319_new_n2524_), .Y(_abc_40319_new_n2732_));
OAI21X1 OAI21X1_515 ( .A(_abc_40319_new_n2730_), .B(_abc_40319_new_n2731_), .C(_abc_40319_new_n2733_), .Y(_abc_40319_new_n2734_));
OAI21X1 OAI21X1_516 ( .A(_abc_40319_new_n2729_), .B(_abc_40319_new_n2734_), .C(_abc_40319_new_n2723_), .Y(_abc_40319_new_n2735_));
OAI21X1 OAI21X1_517 ( .A(_abc_40319_new_n2711_), .B(_abc_40319_new_n2721_), .C(_abc_40319_new_n2736_), .Y(n1014));
OAI21X1 OAI21X1_518 ( .A(REG1_REG_10_), .B(_abc_40319_new_n2716_), .C(_abc_40319_new_n2744_), .Y(_abc_40319_new_n2745_));
OAI21X1 OAI21X1_519 ( .A(_abc_40319_new_n2542_), .B(_abc_40319_new_n2543_), .C(_abc_40319_new_n2523_), .Y(_abc_40319_new_n2747_));
OAI21X1 OAI21X1_52 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(_abc_40319_new_n823_), .Y(_abc_40319_new_n824_));
OAI21X1 OAI21X1_520 ( .A(_abc_40319_new_n2725_), .B(_abc_40319_new_n2731_), .C(_abc_40319_new_n2724_), .Y(_abc_40319_new_n2753_));
OAI21X1 OAI21X1_521 ( .A(_abc_40319_new_n2542_), .B(_abc_40319_new_n2543_), .C(_abc_40319_new_n2756_), .Y(_abc_40319_new_n2757_));
OAI21X1 OAI21X1_522 ( .A(_abc_40319_new_n2746_), .B(_abc_40319_new_n2747_), .C(_abc_40319_new_n2759_), .Y(n1010));
OAI21X1 OAI21X1_523 ( .A(REG1_REG_10_), .B(_abc_40319_new_n2716_), .C(_abc_40319_new_n1390_), .Y(_abc_40319_new_n2766_));
OAI21X1 OAI21X1_524 ( .A(REG1_REG_11_), .B(_abc_40319_new_n1369_), .C(_abc_40319_new_n2767_), .Y(_abc_40319_new_n2768_));
OAI21X1 OAI21X1_525 ( .A(REG2_REG_10_), .B(_abc_40319_new_n1390_), .C(_abc_40319_new_n2728_), .Y(_abc_40319_new_n2773_));
OAI21X1 OAI21X1_526 ( .A(REG2_REG_11_), .B(_abc_40319_new_n1369_), .C(_abc_40319_new_n2774_), .Y(_abc_40319_new_n2775_));
OAI21X1 OAI21X1_527 ( .A(_abc_40319_new_n2542_), .B(_abc_40319_new_n2543_), .C(_abc_40319_new_n2778_), .Y(_abc_40319_new_n2779_));
OAI21X1 OAI21X1_528 ( .A(_abc_40319_new_n2747_), .B(_abc_40319_new_n2769_), .C(_abc_40319_new_n2781_), .Y(n1006));
OAI21X1 OAI21X1_529 ( .A(_abc_40319_new_n1354_), .B(_abc_40319_new_n1348_), .C(_abc_40319_new_n2793_), .Y(_abc_40319_new_n2794_));
OAI21X1 OAI21X1_53 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n822_), .C(_abc_40319_new_n824_), .Y(_abc_40319_new_n825_));
OAI21X1 OAI21X1_530 ( .A(_abc_40319_new_n2791_), .B(_abc_40319_new_n2794_), .C(_abc_40319_new_n2795_), .Y(_abc_40319_new_n2796_));
OAI21X1 OAI21X1_531 ( .A(_abc_40319_new_n2747_), .B(_abc_40319_new_n2788_), .C(_abc_40319_new_n2801_), .Y(n1002));
OAI21X1 OAI21X1_532 ( .A(_abc_40319_new_n2785_), .B(_abc_40319_new_n2805_), .C(REG1_REG_14_), .Y(_abc_40319_new_n2806_));
OAI21X1 OAI21X1_533 ( .A(_abc_40319_new_n1252_), .B(_abc_40319_new_n2803_), .C(_abc_40319_new_n1246_), .Y(_abc_40319_new_n2809_));
OAI21X1 OAI21X1_534 ( .A(REG2_REG_13_), .B(_abc_40319_new_n1322_), .C(_abc_40319_new_n2817_), .Y(_abc_40319_new_n2818_));
OAI21X1 OAI21X1_535 ( .A(_abc_40319_new_n1246_), .B(_abc_40319_new_n2683_), .C(_abc_40319_new_n1520_), .Y(_abc_40319_new_n2821_));
OAI21X1 OAI21X1_536 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n1246_), .C(_abc_40319_new_n2824_), .Y(_abc_40319_new_n2825_));
OAI21X1 OAI21X1_537 ( .A(_abc_40319_new_n2747_), .B(_abc_40319_new_n2811_), .C(_abc_40319_new_n2826_), .Y(n998));
OAI21X1 OAI21X1_538 ( .A(_abc_40319_new_n1249_), .B(_abc_40319_new_n1246_), .C(_abc_40319_new_n2842_), .Y(_abc_40319_new_n2843_));
OAI21X1 OAI21X1_539 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n1221_), .C(_abc_40319_new_n2845_), .Y(_abc_40319_new_n2846_));
OAI21X1 OAI21X1_54 ( .A(IR_REG_0_), .B(IR_REG_1_), .C(IR_REG_31_), .Y(_abc_40319_new_n835_));
OAI21X1 OAI21X1_540 ( .A(_abc_40319_new_n1221_), .B(_abc_40319_new_n2683_), .C(_abc_40319_new_n1866_), .Y(_abc_40319_new_n2848_));
OAI21X1 OAI21X1_541 ( .A(_abc_40319_new_n2747_), .B(_abc_40319_new_n2833_), .C(_abc_40319_new_n2851_), .Y(n994));
OAI21X1 OAI21X1_542 ( .A(_abc_40319_new_n1224_), .B(_abc_40319_new_n2828_), .C(_abc_40319_new_n1221_), .Y(_abc_40319_new_n2859_));
OAI21X1 OAI21X1_543 ( .A(REG1_REG_15_), .B(_abc_40319_new_n2830_), .C(_abc_40319_new_n2859_), .Y(_abc_40319_new_n2860_));
OAI21X1 OAI21X1_544 ( .A(REG2_REG_15_), .B(_abc_40319_new_n2836_), .C(_abc_40319_new_n2868_), .Y(_abc_40319_new_n2869_));
OAI21X1 OAI21X1_545 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n1173_), .C(_abc_40319_new_n2874_), .Y(_abc_40319_new_n2875_));
OAI21X1 OAI21X1_546 ( .A(_abc_40319_new_n2747_), .B(_abc_40319_new_n2861_), .C(_abc_40319_new_n2876_), .Y(n990));
OAI21X1 OAI21X1_547 ( .A(_abc_40319_new_n1179_), .B(_abc_40319_new_n1173_), .C(_abc_40319_new_n2882_), .Y(_abc_40319_new_n2883_));
OAI21X1 OAI21X1_548 ( .A(_abc_40319_new_n1176_), .B(_abc_40319_new_n1173_), .C(_abc_40319_new_n2888_), .Y(_abc_40319_new_n2889_));
OAI21X1 OAI21X1_549 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n1196_), .C(_abc_40319_new_n2891_), .Y(_abc_40319_new_n2892_));
OAI21X1 OAI21X1_55 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_2_), .Y(_abc_40319_new_n838_));
OAI21X1 OAI21X1_550 ( .A(_abc_40319_new_n1196_), .B(_abc_40319_new_n2683_), .C(_abc_40319_new_n2894_), .Y(_abc_40319_new_n2895_));
OAI21X1 OAI21X1_551 ( .A(_abc_40319_new_n2747_), .B(_abc_40319_new_n2884_), .C(_abc_40319_new_n2897_), .Y(n986));
OAI21X1 OAI21X1_552 ( .A(REG1_REG_15_), .B(_abc_40319_new_n2830_), .C(_abc_40319_new_n2836_), .Y(_abc_40319_new_n2903_));
OAI21X1 OAI21X1_553 ( .A(_abc_40319_new_n1199_), .B(_abc_40319_new_n1196_), .C(_abc_40319_new_n2905_), .Y(_abc_40319_new_n2906_));
OAI21X1 OAI21X1_554 ( .A(_abc_40319_new_n2900_), .B(_abc_40319_new_n2901_), .C(_abc_40319_new_n2906_), .Y(_abc_40319_new_n2907_));
OAI21X1 OAI21X1_555 ( .A(REG1_REG_17_), .B(_abc_40319_new_n2879_), .C(_abc_40319_new_n2911_), .Y(_abc_40319_new_n2912_));
OAI21X1 OAI21X1_556 ( .A(REG2_REG_17_), .B(_abc_40319_new_n2879_), .C(_abc_40319_new_n2921_), .Y(_abc_40319_new_n2922_));
OAI21X1 OAI21X1_557 ( .A(_abc_40319_new_n2920_), .B(_abc_40319_new_n2922_), .C(_abc_40319_new_n2524_), .Y(_abc_40319_new_n2923_));
OAI21X1 OAI21X1_558 ( .A(_abc_40319_new_n2924_), .B(_abc_40319_new_n2914_), .C(_abc_40319_new_n2623_), .Y(_abc_40319_new_n2925_));
OAI21X1 OAI21X1_559 ( .A(REG2_REG_18_), .B(_abc_40319_new_n2899_), .C(_abc_40319_new_n2940_), .Y(_abc_40319_new_n2941_));
OAI21X1 OAI21X1_56 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n837_), .C(_abc_40319_new_n838_), .Y(_abc_40319_new_n839_));
OAI21X1 OAI21X1_560 ( .A(_abc_40319_new_n2939_), .B(_abc_40319_new_n667_), .C(_abc_40319_new_n2919_), .Y(_abc_40319_new_n2943_));
OAI21X1 OAI21X1_561 ( .A(_abc_40319_new_n2915_), .B(_abc_40319_new_n2922_), .C(_abc_40319_new_n2944_), .Y(_abc_40319_new_n2945_));
OAI21X1 OAI21X1_562 ( .A(_abc_40319_new_n2947_), .B(_abc_40319_new_n2938_), .C(_abc_40319_new_n2543_), .Y(_abc_40319_new_n2948_));
OAI21X1 OAI21X1_563 ( .A(_abc_40319_new_n2949_), .B(_abc_40319_new_n2938_), .C(_abc_40319_new_n2542_), .Y(_abc_40319_new_n2950_));
OAI21X1 OAI21X1_564 ( .A(_abc_40319_new_n616_), .B(_abc_40319_new_n668_), .C(_abc_40319_new_n654_), .Y(_abc_40319_new_n2957_));
OAI21X1 OAI21X1_565 ( .A(_abc_40319_new_n972_), .B(_abc_40319_new_n1007_), .C(_abc_40319_new_n2959_), .Y(_abc_40319_new_n2960_));
OAI21X1 OAI21X1_566 ( .A(_abc_40319_new_n593_), .B(_abc_40319_new_n602_), .C(_abc_40319_new_n615_), .Y(_abc_40319_new_n2985_));
OAI21X1 OAI21X1_567 ( .A(_abc_40319_new_n1878_), .B(_abc_40319_new_n1881_), .C(_abc_40319_new_n2986_), .Y(_abc_40319_new_n2987_));
OAI21X1 OAI21X1_568 ( .A(REG2_REG_31_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n2988_), .Y(_abc_40319_new_n2989_));
OAI21X1 OAI21X1_569 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n2992_), .C(_abc_40319_new_n2989_), .Y(_abc_40319_new_n2993_));
OAI21X1 OAI21X1_57 ( .A(_abc_40319_new_n751_), .B(_abc_40319_new_n746_), .C(_abc_40319_new_n839_), .Y(_abc_40319_new_n845_));
OAI21X1 OAI21X1_570 ( .A(_abc_40319_new_n2961_), .B(_abc_40319_new_n2984_), .C(_abc_40319_new_n2994_), .Y(n973));
OAI21X1 OAI21X1_571 ( .A(REG2_REG_30_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n2988_), .Y(_abc_40319_new_n2999_));
OAI21X1 OAI21X1_572 ( .A(_abc_40319_new_n2096_), .B(_abc_40319_new_n2992_), .C(_abc_40319_new_n2999_), .Y(_abc_40319_new_n3000_));
OAI21X1 OAI21X1_573 ( .A(_abc_40319_new_n2453_), .B(_abc_40319_new_n2505_), .C(_abc_40319_new_n2260_), .Y(_abc_40319_new_n3003_));
OAI21X1 OAI21X1_574 ( .A(_abc_40319_new_n609_), .B(_abc_40319_new_n749_), .C(_abc_40319_new_n743_), .Y(_abc_40319_new_n3005_));
OAI21X1 OAI21X1_575 ( .A(_abc_40319_new_n1150_), .B(_abc_40319_new_n1155_), .C(_abc_40319_new_n1148_), .Y(_abc_40319_new_n3008_));
OAI21X1 OAI21X1_576 ( .A(_abc_40319_new_n1460_), .B(_abc_40319_new_n1469_), .C(_abc_40319_new_n3010_), .Y(_abc_40319_new_n3011_));
OAI21X1 OAI21X1_577 ( .A(_abc_40319_new_n1443_), .B(_abc_40319_new_n1452_), .C(_abc_40319_new_n3013_), .Y(_abc_40319_new_n3014_));
OAI21X1 OAI21X1_578 ( .A(_abc_40319_new_n1459_), .B(_abc_40319_new_n1760_), .C(_abc_40319_new_n3014_), .Y(_abc_40319_new_n3015_));
OAI21X1 OAI21X1_579 ( .A(_abc_40319_new_n1198_), .B(_abc_40319_new_n3020_), .C(_abc_40319_new_n1209_), .Y(_abc_40319_new_n3021_));
OAI21X1 OAI21X1_58 ( .A(_abc_40319_new_n846_), .B(_abc_40319_new_n849_), .C(_abc_40319_new_n679_), .Y(_abc_40319_new_n850_));
OAI21X1 OAI21X1_580 ( .A(_abc_40319_new_n1211_), .B(_abc_40319_new_n2198_), .C(_abc_40319_new_n3021_), .Y(_abc_40319_new_n3022_));
OAI21X1 OAI21X1_581 ( .A(_abc_40319_new_n3019_), .B(_abc_40319_new_n3023_), .C(_abc_40319_new_n3016_), .Y(_abc_40319_new_n3024_));
OAI21X1 OAI21X1_582 ( .A(_abc_40319_new_n1123_), .B(_abc_40319_new_n1135_), .C(_abc_40319_new_n3024_), .Y(_abc_40319_new_n3025_));
OAI21X1 OAI21X1_583 ( .A(_abc_40319_new_n1122_), .B(_abc_40319_new_n1137_), .C(_abc_40319_new_n3025_), .Y(_abc_40319_new_n3026_));
OAI21X1 OAI21X1_584 ( .A(_abc_40319_new_n1226_), .B(_abc_40319_new_n1232_), .C(_abc_40319_new_n1223_), .Y(_abc_40319_new_n3029_));
OAI21X1 OAI21X1_585 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n1378_), .C(_abc_40319_new_n1371_), .Y(_abc_40319_new_n3033_));
OAI21X1 OAI21X1_586 ( .A(_abc_40319_new_n3033_), .B(_abc_40319_new_n3032_), .C(_abc_40319_new_n3034_), .Y(_abc_40319_new_n3035_));
OAI21X1 OAI21X1_587 ( .A(_abc_40319_new_n1325_), .B(_abc_40319_new_n1336_), .C(_abc_40319_new_n3035_), .Y(_abc_40319_new_n3036_));
OAI21X1 OAI21X1_588 ( .A(_abc_40319_new_n877_), .B(_abc_40319_new_n880_), .C(_abc_40319_new_n3037_), .Y(_abc_40319_new_n3038_));
OAI21X1 OAI21X1_589 ( .A(_abc_40319_new_n895_), .B(_abc_40319_new_n897_), .C(_abc_40319_new_n3038_), .Y(_abc_40319_new_n3039_));
OAI21X1 OAI21X1_59 ( .A(_abc_40319_new_n663_), .B(_abc_40319_new_n680_), .C(_abc_40319_new_n574_), .Y(_abc_40319_new_n852_));
OAI21X1 OAI21X1_590 ( .A(_abc_40319_new_n829_), .B(_abc_40319_new_n861_), .C(_abc_40319_new_n826_), .Y(_abc_40319_new_n3046_));
OAI21X1 OAI21X1_591 ( .A(_abc_40319_new_n849_), .B(_abc_40319_new_n846_), .C(_abc_40319_new_n839_), .Y(_abc_40319_new_n3047_));
OAI21X1 OAI21X1_592 ( .A(_abc_40319_new_n3047_), .B(_abc_40319_new_n3042_), .C(_abc_40319_new_n3046_), .Y(_abc_40319_new_n3048_));
OAI21X1 OAI21X1_593 ( .A(_abc_40319_new_n803_), .B(_abc_40319_new_n808_), .C(_abc_40319_new_n799_), .Y(_abc_40319_new_n3049_));
OAI21X1 OAI21X1_594 ( .A(_abc_40319_new_n782_), .B(_abc_40319_new_n775_), .C(_abc_40319_new_n769_), .Y(_abc_40319_new_n3050_));
OAI21X1 OAI21X1_595 ( .A(_abc_40319_new_n3049_), .B(_abc_40319_new_n3040_), .C(_abc_40319_new_n3050_), .Y(_abc_40319_new_n3051_));
OAI21X1 OAI21X1_596 ( .A(_abc_40319_new_n1297_), .B(_abc_40319_new_n1309_), .C(_abc_40319_new_n2205_), .Y(_abc_40319_new_n3055_));
OAI21X1 OAI21X1_597 ( .A(_abc_40319_new_n2192_), .B(_abc_40319_new_n3055_), .C(_abc_40319_new_n3056_), .Y(_abc_40319_new_n3057_));
OAI21X1 OAI21X1_598 ( .A(_abc_40319_new_n953_), .B(_abc_40319_new_n950_), .C(_abc_40319_new_n944_), .Y(_abc_40319_new_n3058_));
OAI21X1 OAI21X1_599 ( .A(_abc_40319_new_n698_), .B(_abc_40319_new_n3059_), .C(_abc_40319_new_n740_), .Y(_abc_40319_new_n3060_));
OAI21X1 OAI21X1_6 ( .A(IR_REG_22_), .B(_abc_40319_new_n576_), .C(IR_REG_23_), .Y(_abc_40319_new_n577_));
OAI21X1 OAI21X1_60 ( .A(_abc_40319_new_n856_), .B(_abc_40319_new_n854_), .C(_abc_40319_new_n745_), .Y(_abc_40319_new_n857_));
OAI21X1 OAI21X1_600 ( .A(_abc_40319_new_n2388_), .B(_abc_40319_new_n3058_), .C(_abc_40319_new_n3060_), .Y(_abc_40319_new_n3061_));
OAI21X1 OAI21X1_601 ( .A(_abc_40319_new_n3054_), .B(_abc_40319_new_n3066_), .C(_abc_40319_new_n3064_), .Y(_abc_40319_new_n3067_));
OAI21X1 OAI21X1_602 ( .A(_abc_40319_new_n1371_), .B(_abc_40319_new_n1380_), .C(_abc_40319_new_n3067_), .Y(_abc_40319_new_n3068_));
OAI21X1 OAI21X1_603 ( .A(_abc_40319_new_n3032_), .B(_abc_40319_new_n3068_), .C(_abc_40319_new_n3036_), .Y(_abc_40319_new_n3069_));
OAI21X1 OAI21X1_604 ( .A(_abc_40319_new_n3028_), .B(_abc_40319_new_n3070_), .C(_abc_40319_new_n3029_), .Y(_abc_40319_new_n3071_));
OAI21X1 OAI21X1_605 ( .A(_abc_40319_new_n1198_), .B(_abc_40319_new_n1209_), .C(_abc_40319_new_n2197_), .Y(_abc_40319_new_n3072_));
OAI21X1 OAI21X1_606 ( .A(_abc_40319_new_n2136_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n1710_), .Y(_abc_40319_new_n3078_));
OAI21X1 OAI21X1_607 ( .A(_abc_40319_new_n2258_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n1592_), .Y(_abc_40319_new_n3079_));
OAI21X1 OAI21X1_608 ( .A(_abc_40319_new_n1085_), .B(_abc_40319_new_n1094_), .C(_abc_40319_new_n3081_), .Y(_abc_40319_new_n3082_));
OAI21X1 OAI21X1_609 ( .A(_abc_40319_new_n1054_), .B(_abc_40319_new_n1496_), .C(_abc_40319_new_n3087_), .Y(_abc_40319_new_n3088_));
OAI21X1 OAI21X1_61 ( .A(_abc_40319_new_n751_), .B(_abc_40319_new_n746_), .C(_abc_40319_new_n826_), .Y(_abc_40319_new_n860_));
OAI21X1 OAI21X1_610 ( .A(_abc_40319_new_n1055_), .B(_abc_40319_new_n1065_), .C(_abc_40319_new_n3088_), .Y(_abc_40319_new_n3089_));
OAI21X1 OAI21X1_611 ( .A(_abc_40319_new_n3094_), .B(_abc_40319_new_n3085_), .C(_abc_40319_new_n2120_), .Y(_abc_40319_new_n3095_));
OAI21X1 OAI21X1_612 ( .A(_abc_40319_new_n614_), .B(_abc_40319_new_n1874_), .C(_abc_40319_new_n749_), .Y(_abc_40319_new_n3098_));
OAI21X1 OAI21X1_613 ( .A(_abc_40319_new_n608_), .B(_abc_40319_new_n678_), .C(_abc_40319_new_n3099_), .Y(_abc_40319_new_n3100_));
OAI21X1 OAI21X1_614 ( .A(_abc_40319_new_n1592_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3102_), .Y(_abc_40319_new_n3105_));
OAI21X1 OAI21X1_615 ( .A(_abc_40319_new_n1581_), .B(_abc_40319_new_n2992_), .C(_abc_40319_new_n3112_), .Y(_abc_40319_new_n3113_));
OAI21X1 OAI21X1_616 ( .A(_abc_40319_new_n3109_), .B(_abc_40319_new_n3110_), .C(_abc_40319_new_n3114_), .Y(_abc_40319_new_n3115_));
OAI21X1 OAI21X1_617 ( .A(_abc_40319_new_n1109_), .B(_abc_40319_new_n1115_), .C(_abc_40319_new_n3077_), .Y(_abc_40319_new_n3120_));
OAI21X1 OAI21X1_618 ( .A(_abc_40319_new_n3082_), .B(_abc_40319_new_n3120_), .C(_abc_40319_new_n3121_), .Y(_abc_40319_new_n3122_));
OAI21X1 OAI21X1_619 ( .A(_abc_40319_new_n3080_), .B(_abc_40319_new_n3086_), .C(_abc_40319_new_n3122_), .Y(_abc_40319_new_n3124_));
OAI21X1 OAI21X1_62 ( .A(_abc_40319_new_n829_), .B(_abc_40319_new_n861_), .C(_abc_40319_new_n679_), .Y(_abc_40319_new_n862_));
OAI21X1 OAI21X1_620 ( .A(_abc_40319_new_n2454_), .B(_abc_40319_new_n3126_), .C(_abc_40319_new_n2123_), .Y(_abc_40319_new_n3127_));
OAI21X1 OAI21X1_621 ( .A(_abc_40319_new_n3119_), .B(_abc_40319_new_n3127_), .C(_abc_40319_new_n3005_), .Y(_abc_40319_new_n3129_));
OAI21X1 OAI21X1_622 ( .A(_abc_40319_new_n2122_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n2977_), .Y(_abc_40319_new_n3135_));
OAI21X1 OAI21X1_623 ( .A(_abc_40319_new_n1009_), .B(_abc_40319_new_n1041_), .C(nRESET_G), .Y(_abc_40319_new_n3138_));
OAI21X1 OAI21X1_624 ( .A(_abc_40319_new_n2126_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n1078_), .Y(_abc_40319_new_n3145_));
OAI21X1 OAI21X1_625 ( .A(_abc_40319_new_n3147_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n1093_), .Y(_abc_40319_new_n3148_));
OAI21X1 OAI21X1_626 ( .A(_abc_40319_new_n1080_), .B(_abc_40319_new_n1077_), .C(_abc_40319_new_n3150_), .Y(_abc_40319_new_n3152_));
OAI21X1 OAI21X1_627 ( .A(_abc_40319_new_n1080_), .B(_abc_40319_new_n3161_), .C(_abc_40319_new_n1055_), .Y(_abc_40319_new_n3162_));
OAI21X1 OAI21X1_628 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n1054_), .C(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3165_));
OAI21X1 OAI21X1_629 ( .A(REG2_REG_26_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3165_), .Y(_abc_40319_new_n3166_));
OAI21X1 OAI21X1_63 ( .A(_abc_40319_new_n866_), .B(_abc_40319_new_n864_), .C(_abc_40319_new_n745_), .Y(_abc_40319_new_n867_));
OAI21X1 OAI21X1_630 ( .A(_abc_40319_new_n1592_), .B(_abc_40319_new_n3164_), .C(_abc_40319_new_n3168_), .Y(_abc_40319_new_n3169_));
OAI21X1 OAI21X1_631 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3158_), .C(_abc_40319_new_n3172_), .Y(n948));
OAI21X1 OAI21X1_632 ( .A(_abc_40319_new_n1084_), .B(_abc_40319_new_n1093_), .C(_abc_40319_new_n3149_), .Y(_abc_40319_new_n3174_));
OAI21X1 OAI21X1_633 ( .A(_abc_40319_new_n3179_), .B(_abc_40319_new_n2491_), .C(_abc_40319_new_n2500_), .Y(_abc_40319_new_n3180_));
OAI21X1 OAI21X1_634 ( .A(_abc_40319_new_n2129_), .B(_abc_40319_new_n3184_), .C(_abc_40319_new_n3005_), .Y(_abc_40319_new_n3186_));
OAI21X1 OAI21X1_635 ( .A(_abc_40319_new_n3193_), .B(_abc_40319_new_n3195_), .C(nRESET_G), .Y(_abc_40319_new_n3196_));
OAI21X1 OAI21X1_636 ( .A(_abc_40319_new_n1496_), .B(_abc_40319_new_n3164_), .C(_abc_40319_new_n3197_), .Y(_abc_40319_new_n3198_));
OAI21X1 OAI21X1_637 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3188_), .C(_abc_40319_new_n3201_), .Y(n943));
OAI21X1 OAI21X1_638 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3207_), .C(_abc_40319_new_n3205_), .Y(_abc_40319_new_n3208_));
OAI21X1 OAI21X1_639 ( .A(_abc_40319_new_n2213_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n2975_), .Y(_abc_40319_new_n3211_));
OAI21X1 OAI21X1_64 ( .A(_abc_40319_new_n871_), .B(_abc_40319_new_n544_), .C(_abc_40319_new_n872_), .Y(_abc_40319_new_n873_));
OAI21X1 OAI21X1_640 ( .A(_abc_40319_new_n1109_), .B(_abc_40319_new_n3211_), .C(_abc_40319_new_n1085_), .Y(_abc_40319_new_n3212_));
OAI21X1 OAI21X1_641 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n1084_), .C(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3214_));
OAI21X1 OAI21X1_642 ( .A(REG2_REG_24_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3214_), .Y(_abc_40319_new_n3215_));
OAI21X1 OAI21X1_643 ( .A(_abc_40319_new_n1078_), .B(_abc_40319_new_n3164_), .C(_abc_40319_new_n3217_), .Y(_abc_40319_new_n3218_));
OAI21X1 OAI21X1_644 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3209_), .C(_abc_40319_new_n3221_), .Y(n938));
OAI21X1 OAI21X1_645 ( .A(_abc_40319_new_n1123_), .B(_abc_40319_new_n3224_), .C(_abc_40319_new_n1109_), .Y(_abc_40319_new_n3225_));
OAI21X1 OAI21X1_646 ( .A(_abc_40319_new_n1108_), .B(_abc_40319_new_n1115_), .C(_abc_40319_new_n2457_), .Y(_abc_40319_new_n3232_));
OAI21X1 OAI21X1_647 ( .A(_abc_40319_new_n1122_), .B(_abc_40319_new_n1135_), .C(_abc_40319_new_n2139_), .Y(_abc_40319_new_n3234_));
OAI21X1 OAI21X1_648 ( .A(_abc_40319_new_n3231_), .B(_abc_40319_new_n3232_), .C(_abc_40319_new_n3236_), .Y(_abc_40319_new_n3237_));
OAI21X1 OAI21X1_649 ( .A(_abc_40319_new_n1137_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3238_), .Y(_abc_40319_new_n3239_));
OAI21X1 OAI21X1_65 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_1_), .Y(_abc_40319_new_n876_));
OAI21X1 OAI21X1_650 ( .A(_abc_40319_new_n3247_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n3248_), .Y(_abc_40319_new_n3249_));
OAI21X1 OAI21X1_651 ( .A(_abc_40319_new_n1460_), .B(_abc_40319_new_n3249_), .C(_abc_40319_new_n1123_), .Y(_abc_40319_new_n3250_));
OAI21X1 OAI21X1_652 ( .A(_abc_40319_new_n3019_), .B(_abc_40319_new_n3253_), .C(_abc_40319_new_n3016_), .Y(_abc_40319_new_n3254_));
OAI21X1 OAI21X1_653 ( .A(_abc_40319_new_n1760_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3258_), .Y(_abc_40319_new_n3259_));
OAI21X1 OAI21X1_654 ( .A(_abc_40319_new_n3017_), .B(_abc_40319_new_n3253_), .C(_abc_40319_new_n3008_), .Y(_abc_40319_new_n3266_));
OAI21X1 OAI21X1_655 ( .A(_abc_40319_new_n1429_), .B(_abc_40319_new_n1437_), .C(_abc_40319_new_n3266_), .Y(_abc_40319_new_n3267_));
OAI21X1 OAI21X1_656 ( .A(_abc_40319_new_n3009_), .B(_abc_40319_new_n3267_), .C(_abc_40319_new_n3014_), .Y(_abc_40319_new_n3268_));
OAI21X1 OAI21X1_657 ( .A(_abc_40319_new_n3265_), .B(_abc_40319_new_n3230_), .C(_abc_40319_new_n3005_), .Y(_abc_40319_new_n3270_));
OAI21X1 OAI21X1_658 ( .A(_abc_40319_new_n3100_), .B(_abc_40319_new_n3269_), .C(_abc_40319_new_n3272_), .Y(_abc_40319_new_n3273_));
OAI21X1 OAI21X1_659 ( .A(_abc_40319_new_n1443_), .B(_abc_40319_new_n2974_), .C(_abc_40319_new_n1460_), .Y(_abc_40319_new_n3276_));
OAI21X1 OAI21X1_66 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n875_), .C(_abc_40319_new_n876_), .Y(_abc_40319_new_n877_));
OAI21X1 OAI21X1_660 ( .A(_abc_40319_new_n1463_), .B(_abc_40319_new_n1009_), .C(nRESET_G), .Y(_abc_40319_new_n3278_));
OAI21X1 OAI21X1_661 ( .A(_abc_40319_new_n1137_), .B(_abc_40319_new_n3164_), .C(_abc_40319_new_n3280_), .Y(_abc_40319_new_n3281_));
OAI21X1 OAI21X1_662 ( .A(_abc_40319_new_n3110_), .B(_abc_40319_new_n3269_), .C(_abc_40319_new_n3282_), .Y(_abc_40319_new_n3283_));
OAI21X1 OAI21X1_663 ( .A(_abc_40319_new_n1570_), .B(_abc_40319_new_n1759_), .C(_abc_40319_new_n3267_), .Y(_abc_40319_new_n3286_));
OAI21X1 OAI21X1_664 ( .A(_abc_40319_new_n1431_), .B(_abc_40319_new_n1436_), .C(_abc_40319_new_n3103_), .Y(_abc_40319_new_n3289_));
OAI21X1 OAI21X1_665 ( .A(_abc_40319_new_n2167_), .B(_abc_40319_new_n3290_), .C(_abc_40319_new_n2166_), .Y(_abc_40319_new_n3291_));
OAI21X1 OAI21X1_666 ( .A(_abc_40319_new_n2220_), .B(_abc_40319_new_n3291_), .C(_abc_40319_new_n3292_), .Y(_abc_40319_new_n3293_));
OAI21X1 OAI21X1_667 ( .A(_abc_40319_new_n1429_), .B(_abc_40319_new_n3298_), .C(_abc_40319_new_n1443_), .Y(_abc_40319_new_n3299_));
OAI21X1 OAI21X1_668 ( .A(_abc_40319_new_n1446_), .B(_abc_40319_new_n1009_), .C(nRESET_G), .Y(_abc_40319_new_n3303_));
OAI21X1 OAI21X1_669 ( .A(_abc_40319_new_n2170_), .B(_abc_40319_new_n2498_), .C(_abc_40319_new_n3005_), .Y(_abc_40319_new_n3309_));
OAI21X1 OAI21X1_67 ( .A(_abc_40319_new_n751_), .B(_abc_40319_new_n746_), .C(_abc_40319_new_n877_), .Y(_abc_40319_new_n882_));
OAI21X1 OAI21X1_670 ( .A(_abc_40319_new_n1156_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3311_), .Y(_abc_40319_new_n3312_));
OAI21X1 OAI21X1_671 ( .A(_abc_40319_new_n3317_), .B(_abc_40319_new_n2990_), .C(_abc_40319_new_n3318_), .Y(_abc_40319_new_n3319_));
OAI21X1 OAI21X1_672 ( .A(_abc_40319_new_n1567_), .B(_abc_40319_new_n3164_), .C(_abc_40319_new_n3320_), .Y(_abc_40319_new_n3321_));
OAI21X1 OAI21X1_673 ( .A(_abc_40319_new_n2496_), .B(_abc_40319_new_n2491_), .C(_abc_40319_new_n2157_), .Y(_abc_40319_new_n3325_));
OAI21X1 OAI21X1_674 ( .A(_abc_40319_new_n2164_), .B(_abc_40319_new_n3325_), .C(_abc_40319_new_n3326_), .Y(_abc_40319_new_n3327_));
OAI21X1 OAI21X1_675 ( .A(_abc_40319_new_n1208_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3327_), .Y(_abc_40319_new_n3328_));
OAI21X1 OAI21X1_676 ( .A(_abc_40319_new_n1198_), .B(_abc_40319_new_n3332_), .C(_abc_40319_new_n1148_), .Y(_abc_40319_new_n3333_));
OAI21X1 OAI21X1_677 ( .A(_abc_40319_new_n1159_), .B(_abc_40319_new_n2992_), .C(_abc_40319_new_n3335_), .Y(_abc_40319_new_n3336_));
OAI21X1 OAI21X1_678 ( .A(_abc_40319_new_n1759_), .B(_abc_40319_new_n3164_), .C(_abc_40319_new_n3337_), .Y(_abc_40319_new_n3338_));
OAI21X1 OAI21X1_679 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3329_), .C(_abc_40319_new_n3341_), .Y(n908));
OAI21X1 OAI21X1_68 ( .A(IR_REG_31_), .B(_abc_40319_new_n699_), .C(_abc_40319_new_n707_), .Y(_abc_40319_new_n886_));
OAI21X1 OAI21X1_680 ( .A(_abc_40319_new_n2480_), .B(_abc_40319_new_n3349_), .C(_abc_40319_new_n2179_), .Y(_abc_40319_new_n3350_));
OAI21X1 OAI21X1_681 ( .A(_abc_40319_new_n754_), .B(_abc_40319_new_n753_), .C(_abc_40319_new_n2388_), .Y(_abc_40319_new_n3351_));
OAI21X1 OAI21X1_682 ( .A(_abc_40319_new_n1276_), .B(_abc_40319_new_n988_), .C(_abc_40319_new_n3351_), .Y(_abc_40319_new_n3352_));
OAI21X1 OAI21X1_683 ( .A(_abc_40319_new_n2389_), .B(_abc_40319_new_n2477_), .C(_abc_40319_new_n3353_), .Y(_abc_40319_new_n3354_));
OAI21X1 OAI21X1_684 ( .A(_abc_40319_new_n987_), .B(_abc_40319_new_n2427_), .C(_abc_40319_new_n3354_), .Y(_abc_40319_new_n3355_));
OAI21X1 OAI21X1_685 ( .A(_abc_40319_new_n1739_), .B(_abc_40319_new_n1309_), .C(_abc_40319_new_n3347_), .Y(_abc_40319_new_n3356_));
OAI21X1 OAI21X1_686 ( .A(_abc_40319_new_n3356_), .B(_abc_40319_new_n3355_), .C(_abc_40319_new_n3350_), .Y(_abc_40319_new_n3357_));
OAI21X1 OAI21X1_687 ( .A(_abc_40319_new_n1654_), .B(_abc_40319_new_n1360_), .C(_abc_40319_new_n3357_), .Y(_abc_40319_new_n3358_));
OAI21X1 OAI21X1_688 ( .A(_abc_40319_new_n1352_), .B(_abc_40319_new_n1796_), .C(_abc_40319_new_n3358_), .Y(_abc_40319_new_n3359_));
OAI21X1 OAI21X1_689 ( .A(_abc_40319_new_n2486_), .B(_abc_40319_new_n3360_), .C(_abc_40319_new_n2495_), .Y(_abc_40319_new_n3361_));
OAI21X1 OAI21X1_69 ( .A(_abc_40319_new_n885_), .B(_abc_40319_new_n889_), .C(_abc_40319_new_n679_), .Y(_abc_40319_new_n890_));
OAI21X1 OAI21X1_690 ( .A(_abc_40319_new_n3345_), .B(_abc_40319_new_n3363_), .C(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3364_));
OAI21X1 OAI21X1_691 ( .A(_abc_40319_new_n1150_), .B(_abc_40319_new_n1155_), .C(_abc_40319_new_n3368_), .Y(_abc_40319_new_n3369_));
OAI21X1 OAI21X1_692 ( .A(_abc_40319_new_n1202_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3370_), .Y(_abc_40319_new_n3371_));
OAI21X1 OAI21X1_693 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3369_), .C(_abc_40319_new_n3372_), .Y(_abc_40319_new_n3373_));
OAI21X1 OAI21X1_694 ( .A(_abc_40319_new_n1223_), .B(_abc_40319_new_n3377_), .C(_abc_40319_new_n1175_), .Y(_abc_40319_new_n3378_));
OAI21X1 OAI21X1_695 ( .A(_abc_40319_new_n2196_), .B(_abc_40319_new_n2992_), .C(_abc_40319_new_n3380_), .Y(_abc_40319_new_n3381_));
OAI21X1 OAI21X1_696 ( .A(_abc_40319_new_n2384_), .B(_abc_40319_new_n3360_), .C(_abc_40319_new_n2331_), .Y(_abc_40319_new_n3383_));
OAI21X1 OAI21X1_697 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3385_), .C(_abc_40319_new_n3387_), .Y(_abc_40319_new_n3388_));
OAI21X1 OAI21X1_698 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3388_), .C(_abc_40319_new_n3389_), .Y(_abc_40319_new_n3390_));
OAI21X1 OAI21X1_699 ( .A(_abc_40319_new_n3110_), .B(_abc_40319_new_n3382_), .C(_abc_40319_new_n3390_), .Y(_abc_40319_new_n3391_));
OAI21X1 OAI21X1_7 ( .A(IR_REG_31_), .B(_abc_40319_new_n575_), .C(_abc_40319_new_n579_), .Y(_abc_40319_new_n580_));
OAI21X1 OAI21X1_70 ( .A(IR_REG_31_), .B(_abc_40319_new_n544_), .C(_abc_40319_new_n873_), .Y(_abc_40319_new_n892_));
OAI21X1 OAI21X1_700 ( .A(_abc_40319_new_n1865_), .B(_abc_40319_new_n2992_), .C(_abc_40319_new_n3396_), .Y(_abc_40319_new_n3397_));
OAI21X1 OAI21X1_701 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3400_), .C(_abc_40319_new_n3401_), .Y(_abc_40319_new_n3402_));
OAI21X1 OAI21X1_702 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3402_), .C(_abc_40319_new_n3403_), .Y(_abc_40319_new_n3404_));
OAI21X1 OAI21X1_703 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3408_), .C(_abc_40319_new_n3411_), .Y(_abc_40319_new_n3412_));
OAI21X1 OAI21X1_704 ( .A(_abc_40319_new_n1325_), .B(_abc_40319_new_n3415_), .C(_abc_40319_new_n1248_), .Y(_abc_40319_new_n3416_));
OAI21X1 OAI21X1_705 ( .A(_abc_40319_new_n1249_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3420_), .Y(_abc_40319_new_n3421_));
OAI21X1 OAI21X1_706 ( .A(_abc_40319_new_n3110_), .B(_abc_40319_new_n3409_), .C(_abc_40319_new_n3423_), .Y(_abc_40319_new_n3424_));
OAI21X1 OAI21X1_707 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3413_), .C(_abc_40319_new_n3425_), .Y(n888));
OAI21X1 OAI21X1_708 ( .A(_abc_40319_new_n1370_), .B(_abc_40319_new_n1379_), .C(_abc_40319_new_n3068_), .Y(_abc_40319_new_n3428_));
OAI21X1 OAI21X1_709 ( .A(_abc_40319_new_n1352_), .B(_abc_40319_new_n1360_), .C(_abc_40319_new_n3428_), .Y(_abc_40319_new_n3429_));
OAI21X1 OAI21X1_71 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(_abc_40319_new_n893_), .Y(_abc_40319_new_n894_));
OAI21X1 OAI21X1_710 ( .A(_abc_40319_new_n1654_), .B(_abc_40319_new_n1796_), .C(_abc_40319_new_n3429_), .Y(_abc_40319_new_n3430_));
OAI21X1 OAI21X1_711 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3427_), .C(_abc_40319_new_n3432_), .Y(_abc_40319_new_n3433_));
OAI21X1 OAI21X1_712 ( .A(_abc_40319_new_n1258_), .B(_abc_40319_new_n2985_), .C(_abc_40319_new_n3439_), .Y(_abc_40319_new_n3440_));
OAI21X1 OAI21X1_713 ( .A(REG2_REG_13_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3440_), .Y(_abc_40319_new_n3441_));
OAI21X1 OAI21X1_714 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3434_), .C(_abc_40319_new_n3444_), .Y(n883));
OAI21X1 OAI21X1_715 ( .A(_abc_40319_new_n1514_), .B(_abc_40319_new_n3164_), .C(_abc_40319_new_n3450_), .Y(_abc_40319_new_n3451_));
OAI21X1 OAI21X1_716 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3452_), .C(_abc_40319_new_n3453_), .Y(_abc_40319_new_n3454_));
OAI21X1 OAI21X1_717 ( .A(_abc_40319_new_n1393_), .B(_abc_40319_new_n3459_), .C(_abc_40319_new_n1371_), .Y(_abc_40319_new_n3460_));
OAI21X1 OAI21X1_718 ( .A(_abc_40319_new_n1796_), .B(_abc_40319_new_n3164_), .C(_abc_40319_new_n3464_), .Y(_abc_40319_new_n3465_));
OAI21X1 OAI21X1_719 ( .A(_abc_40319_new_n2369_), .B(_abc_40319_new_n3355_), .C(_abc_40319_new_n2338_), .Y(_abc_40319_new_n3466_));
OAI21X1 OAI21X1_72 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n892_), .C(_abc_40319_new_n894_), .Y(_abc_40319_new_n895_));
OAI21X1 OAI21X1_720 ( .A(_abc_40319_new_n2394_), .B(_abc_40319_new_n3467_), .C(_abc_40319_new_n2336_), .Y(_abc_40319_new_n3468_));
OAI21X1 OAI21X1_721 ( .A(_abc_40319_new_n1401_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3470_), .Y(_abc_40319_new_n3471_));
OAI21X1 OAI21X1_722 ( .A(_abc_40319_new_n2194_), .B(_abc_40319_new_n3477_), .C(_abc_40319_new_n2192_), .Y(_abc_40319_new_n3478_));
OAI21X1 OAI21X1_723 ( .A(_abc_40319_new_n2182_), .B(_abc_40319_new_n3479_), .C(_abc_40319_new_n2183_), .Y(_abc_40319_new_n3480_));
OAI21X1 OAI21X1_724 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3476_), .C(_abc_40319_new_n3482_), .Y(_abc_40319_new_n3483_));
OAI21X1 OAI21X1_725 ( .A(_abc_40319_new_n1399_), .B(_abc_40319_new_n1009_), .C(nRESET_G), .Y(_abc_40319_new_n3487_));
OAI21X1 OAI21X1_726 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n1378_), .C(_abc_40319_new_n3368_), .Y(_abc_40319_new_n3490_));
OAI21X1 OAI21X1_727 ( .A(_abc_40319_new_n3489_), .B(_abc_40319_new_n3491_), .C(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3492_));
OAI21X1 OAI21X1_728 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3484_), .C(_abc_40319_new_n3494_), .Y(n868));
OAI21X1 OAI21X1_729 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3496_), .C(_abc_40319_new_n3499_), .Y(_abc_40319_new_n3500_));
OAI21X1 OAI21X1_73 ( .A(_abc_40319_new_n898_), .B(_abc_40319_new_n896_), .C(_abc_40319_new_n745_), .Y(_abc_40319_new_n899_));
OAI21X1 OAI21X1_730 ( .A(_abc_40319_new_n1276_), .B(_abc_40319_new_n2968_), .C(_abc_40319_new_n1297_), .Y(_abc_40319_new_n3502_));
OAI21X1 OAI21X1_731 ( .A(_abc_40319_new_n1396_), .B(_abc_40319_new_n1400_), .C(_abc_40319_new_n3368_), .Y(_abc_40319_new_n3504_));
OAI21X1 OAI21X1_732 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n1739_), .C(_abc_40319_new_n3504_), .Y(_abc_40319_new_n3505_));
OAI21X1 OAI21X1_733 ( .A(_abc_40319_new_n1305_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3506_), .Y(_abc_40319_new_n3507_));
OAI21X1 OAI21X1_734 ( .A(_abc_40319_new_n2961_), .B(_abc_40319_new_n3503_), .C(_abc_40319_new_n3508_), .Y(_abc_40319_new_n3509_));
OAI21X1 OAI21X1_735 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3501_), .C(_abc_40319_new_n3510_), .Y(n863));
OAI21X1 OAI21X1_736 ( .A(_abc_40319_new_n2389_), .B(_abc_40319_new_n2477_), .C(_abc_40319_new_n3351_), .Y(_abc_40319_new_n3512_));
OAI21X1 OAI21X1_737 ( .A(_abc_40319_new_n759_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3515_), .Y(_abc_40319_new_n3516_));
OAI21X1 OAI21X1_738 ( .A(_abc_40319_new_n3520_), .B(_abc_40319_new_n3521_), .C(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3522_));
OAI21X1 OAI21X1_739 ( .A(_abc_40319_new_n1615_), .B(_abc_40319_new_n1009_), .C(nRESET_G), .Y(_abc_40319_new_n3523_));
OAI21X1 OAI21X1_74 ( .A(_abc_40319_new_n749_), .B(_abc_40319_new_n742_), .C(_abc_40319_new_n681_), .Y(_abc_40319_new_n904_));
OAI21X1 OAI21X1_740 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3517_), .C(_abc_40319_new_n3526_), .Y(n858));
OAI21X1 OAI21X1_741 ( .A(_abc_40319_new_n944_), .B(_abc_40319_new_n954_), .C(_abc_40319_new_n3053_), .Y(_abc_40319_new_n3529_));
OAI21X1 OAI21X1_742 ( .A(_abc_40319_new_n2246_), .B(_abc_40319_new_n959_), .C(_abc_40319_new_n3529_), .Y(_abc_40319_new_n3530_));
OAI21X1 OAI21X1_743 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3528_), .C(_abc_40319_new_n3533_), .Y(_abc_40319_new_n3534_));
OAI21X1 OAI21X1_744 ( .A(_abc_40319_new_n944_), .B(_abc_40319_new_n2966_), .C(_abc_40319_new_n698_), .Y(_abc_40319_new_n3536_));
OAI21X1 OAI21X1_745 ( .A(REG2_REG_7_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3540_), .Y(_abc_40319_new_n3541_));
OAI21X1 OAI21X1_746 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3535_), .C(_abc_40319_new_n3544_), .Y(n853));
OAI21X1 OAI21X1_747 ( .A(_abc_40319_new_n1726_), .B(_abc_40319_new_n809_), .C(_abc_40319_new_n2471_), .Y(_abc_40319_new_n3546_));
OAI21X1 OAI21X1_748 ( .A(_abc_40319_new_n799_), .B(_abc_40319_new_n1556_), .C(_abc_40319_new_n3546_), .Y(_abc_40319_new_n3547_));
OAI21X1 OAI21X1_749 ( .A(_abc_40319_new_n2232_), .B(_abc_40319_new_n3547_), .C(_abc_40319_new_n2233_), .Y(_abc_40319_new_n3548_));
OAI21X1 OAI21X1_75 ( .A(_abc_40319_new_n909_), .B(_abc_40319_new_n802_), .C(_abc_40319_new_n910_), .Y(_abc_40319_new_n911_));
OAI21X1 OAI21X1_750 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3557_), .C(_abc_40319_new_n3556_), .Y(_abc_40319_new_n3558_));
OAI21X1 OAI21X1_751 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3552_), .C(_abc_40319_new_n3561_), .Y(n848));
OAI21X1 OAI21X1_752 ( .A(_abc_40319_new_n3564_), .B(_abc_40319_new_n3039_), .C(_abc_40319_new_n3044_), .Y(_abc_40319_new_n3565_));
OAI21X1 OAI21X1_753 ( .A(_abc_40319_new_n825_), .B(_abc_40319_new_n865_), .C(_abc_40319_new_n3565_), .Y(_abc_40319_new_n3566_));
OAI21X1 OAI21X1_754 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3563_), .C(_abc_40319_new_n3568_), .Y(_abc_40319_new_n3569_));
OAI21X1 OAI21X1_755 ( .A(_abc_40319_new_n3573_), .B(_abc_40319_new_n2990_), .C(_abc_40319_new_n3574_), .Y(_abc_40319_new_n3575_));
OAI21X1 OAI21X1_756 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3570_), .C(_abc_40319_new_n3578_), .Y(n838));
OAI21X1 OAI21X1_757 ( .A(_abc_40319_new_n799_), .B(_abc_40319_new_n809_), .C(_abc_40319_new_n3566_), .Y(_abc_40319_new_n3581_));
OAI21X1 OAI21X1_758 ( .A(_abc_40319_new_n1726_), .B(_abc_40319_new_n1556_), .C(_abc_40319_new_n3581_), .Y(_abc_40319_new_n3582_));
OAI21X1 OAI21X1_759 ( .A(_abc_40319_new_n799_), .B(_abc_40319_new_n2964_), .C(_abc_40319_new_n769_), .Y(_abc_40319_new_n3586_));
OAI21X1 OAI21X1_76 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_0_), .Y(_abc_40319_new_n913_));
OAI21X1 OAI21X1_760 ( .A(_abc_40319_new_n781_), .B(_abc_40319_new_n1009_), .C(nRESET_G), .Y(_abc_40319_new_n3590_));
OAI21X1 OAI21X1_761 ( .A(_abc_40319_new_n3110_), .B(_abc_40319_new_n3583_), .C(_abc_40319_new_n3591_), .Y(_abc_40319_new_n3592_));
OAI21X1 OAI21X1_762 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n3585_), .C(_abc_40319_new_n3594_), .Y(n843));
OAI21X1 OAI21X1_763 ( .A(_abc_40319_new_n2155_), .B(_abc_40319_new_n2470_), .C(_abc_40319_new_n3596_), .Y(_abc_40319_new_n3597_));
OAI21X1 OAI21X1_764 ( .A(_abc_40319_new_n3564_), .B(_abc_40319_new_n3039_), .C(_abc_40319_new_n3598_), .Y(_abc_40319_new_n3599_));
OAI21X1 OAI21X1_765 ( .A(_abc_40319_new_n3603_), .B(_abc_40319_new_n3602_), .C(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3604_));
OAI21X1 OAI21X1_766 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n2962_), .C(_abc_40319_new_n826_), .Y(_abc_40319_new_n3605_));
OAI21X1 OAI21X1_767 ( .A(REG3_REG_3_), .B(_abc_40319_new_n1009_), .C(nRESET_G), .Y(_abc_40319_new_n3607_));
OAI21X1 OAI21X1_768 ( .A(_abc_40319_new_n2961_), .B(_abc_40319_new_n3606_), .C(_abc_40319_new_n3608_), .Y(_abc_40319_new_n3609_));
OAI21X1 OAI21X1_769 ( .A(_abc_40319_new_n3613_), .B(_abc_40319_new_n2245_), .C(_abc_40319_new_n3614_), .Y(_abc_40319_new_n3615_));
OAI21X1 OAI21X1_77 ( .A(_abc_40319_new_n871_), .B(_abc_40319_new_n603_), .C(_abc_40319_new_n913_), .Y(_abc_40319_new_n914_));
OAI21X1 OAI21X1_770 ( .A(_abc_40319_new_n3100_), .B(_abc_40319_new_n3612_), .C(_abc_40319_new_n3615_), .Y(_abc_40319_new_n3616_));
OAI21X1 OAI21X1_771 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n2962_), .C(_abc_40319_new_n3620_), .Y(_abc_40319_new_n3621_));
OAI21X1 OAI21X1_772 ( .A(_abc_40319_new_n667_), .B(_abc_40319_new_n3623_), .C(_abc_40319_new_n3619_), .Y(_abc_40319_new_n3624_));
OAI21X1 OAI21X1_773 ( .A(_abc_40319_new_n847_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3625_), .Y(_abc_40319_new_n3626_));
OAI21X1 OAI21X1_774 ( .A(_abc_40319_new_n3110_), .B(_abc_40319_new_n3612_), .C(_abc_40319_new_n3627_), .Y(n828));
OAI21X1 OAI21X1_775 ( .A(_abc_40319_new_n1905_), .B(_abc_40319_new_n3631_), .C(_abc_40319_new_n3632_), .Y(_abc_40319_new_n3633_));
OAI21X1 OAI21X1_776 ( .A(_abc_40319_new_n3100_), .B(_abc_40319_new_n3629_), .C(_abc_40319_new_n3633_), .Y(_abc_40319_new_n3634_));
OAI21X1 OAI21X1_777 ( .A(_abc_40319_new_n895_), .B(_abc_40319_new_n922_), .C(_abc_40319_new_n3636_), .Y(_abc_40319_new_n3637_));
OAI21X1 OAI21X1_778 ( .A(_abc_40319_new_n667_), .B(_abc_40319_new_n3637_), .C(_abc_40319_new_n3638_), .Y(_abc_40319_new_n3639_));
OAI21X1 OAI21X1_779 ( .A(_abc_40319_new_n3639_), .B(_abc_40319_new_n3635_), .C(_abc_40319_new_n2960_), .Y(_abc_40319_new_n3640_));
OAI21X1 OAI21X1_78 ( .A(_abc_40319_new_n912_), .B(_abc_40319_new_n905_), .C(_abc_40319_new_n915_), .Y(_abc_40319_new_n916_));
OAI21X1 OAI21X1_780 ( .A(_abc_40319_new_n1624_), .B(_abc_40319_new_n1009_), .C(nRESET_G), .Y(_abc_40319_new_n3641_));
OAI21X1 OAI21X1_781 ( .A(_abc_40319_new_n3110_), .B(_abc_40319_new_n3629_), .C(_abc_40319_new_n3643_), .Y(n823));
OAI21X1 OAI21X1_782 ( .A(_abc_40319_new_n3005_), .B(_abc_40319_new_n3101_), .C(_abc_40319_new_n2237_), .Y(_abc_40319_new_n3645_));
OAI21X1 OAI21X1_783 ( .A(_abc_40319_new_n897_), .B(_abc_40319_new_n2985_), .C(_abc_40319_new_n3645_), .Y(_abc_40319_new_n3646_));
OAI21X1 OAI21X1_784 ( .A(_abc_40319_new_n993_), .B(_abc_40319_new_n2955_), .C(_abc_40319_new_n914_), .Y(_abc_40319_new_n3647_));
OAI21X1 OAI21X1_785 ( .A(_abc_40319_new_n1750_), .B(_abc_40319_new_n1009_), .C(nRESET_G), .Y(_abc_40319_new_n3650_));
OAI21X1 OAI21X1_786 ( .A(_abc_40319_new_n3654_), .B(_abc_40319_new_n704_), .C(_abc_40319_new_n3655_), .Y(n333));
OAI21X1 OAI21X1_787 ( .A(_abc_40319_new_n627_), .B(_abc_40319_new_n972_), .C(nRESET_G), .Y(_abc_40319_new_n3657_));
OAI21X1 OAI21X1_788 ( .A(_abc_40319_new_n3726_), .B(_abc_40319_new_n1011_), .C(_abc_40319_new_n3727_), .Y(_abc_40319_new_n3728_));
OAI21X1 OAI21X1_789 ( .A(_abc_40319_new_n3654_), .B(_abc_40319_new_n695_), .C(nRESET_G), .Y(_abc_40319_new_n3729_));
OAI21X1 OAI21X1_79 ( .A(_abc_40319_new_n908_), .B(_abc_40319_new_n911_), .C(_abc_40319_new_n683_), .Y(_abc_40319_new_n918_));
OAI21X1 OAI21X1_790 ( .A(_abc_40319_new_n2122_), .B(_abc_40319_new_n1011_), .C(_abc_40319_new_n3734_), .Y(_abc_40319_new_n3735_));
OAI21X1 OAI21X1_791 ( .A(_abc_40319_new_n3654_), .B(_abc_40319_new_n569_), .C(_abc_40319_new_n3736_), .Y(n308));
OAI21X1 OAI21X1_792 ( .A(_abc_40319_new_n2126_), .B(_abc_40319_new_n1011_), .C(_abc_40319_new_n3738_), .Y(_abc_40319_new_n3739_));
OAI21X1 OAI21X1_793 ( .A(_abc_40319_new_n3654_), .B(_abc_40319_new_n565_), .C(_abc_40319_new_n3740_), .Y(n303));
OAI21X1 OAI21X1_794 ( .A(_abc_40319_new_n3147_), .B(_abc_40319_new_n1011_), .C(_abc_40319_new_n3743_), .Y(_abc_40319_new_n3744_));
OAI21X1 OAI21X1_795 ( .A(_abc_40319_new_n3654_), .B(_abc_40319_new_n3742_), .C(_abc_40319_new_n3745_), .Y(n298));
OAI21X1 OAI21X1_796 ( .A(_abc_40319_new_n618_), .B(_abc_40319_new_n1870_), .C(_abc_40319_new_n3747_), .Y(n293));
OAI21X1 OAI21X1_797 ( .A(_abc_40319_new_n2213_), .B(_abc_40319_new_n1011_), .C(_abc_40319_new_n3749_), .Y(_abc_40319_new_n3750_));
OAI21X1 OAI21X1_798 ( .A(_abc_40319_new_n3654_), .B(_abc_40319_new_n606_), .C(_abc_40319_new_n3751_), .Y(n288));
OAI21X1 OAI21X1_799 ( .A(_abc_40319_new_n3247_), .B(_abc_40319_new_n1011_), .C(_abc_40319_new_n3756_), .Y(_abc_40319_new_n3757_));
OAI21X1 OAI21X1_8 ( .A(IR_REG_26_), .B(_abc_40319_new_n562_), .C(IR_REG_27_), .Y(_abc_40319_new_n587_));
OAI21X1 OAI21X1_80 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(_abc_40319_new_n920_), .Y(_abc_40319_new_n921_));
OAI21X1 OAI21X1_800 ( .A(_abc_40319_new_n3654_), .B(_abc_40319_new_n661_), .C(_abc_40319_new_n3758_), .Y(n278));
OAI21X1 OAI21X1_801 ( .A(_abc_40319_new_n1350_), .B(_abc_40319_new_n1011_), .C(_abc_40319_new_n3782_), .Y(_abc_40319_new_n3783_));
OAI21X1 OAI21X1_802 ( .A(_abc_40319_new_n1318_), .B(_abc_40319_new_n1290_), .C(_abc_40319_new_n1345_), .Y(_abc_40319_new_n3784_));
OAI21X1 OAI21X1_803 ( .A(_abc_40319_new_n3654_), .B(_abc_40319_new_n3784_), .C(nRESET_G), .Y(_abc_40319_new_n3785_));
OAI21X1 OAI21X1_804 ( .A(_abc_40319_new_n823_), .B(_abc_40319_new_n1011_), .C(_abc_40319_new_n3811_), .Y(_abc_40319_new_n3812_));
OAI21X1 OAI21X1_805 ( .A(_abc_40319_new_n819_), .B(_abc_40319_new_n3654_), .C(_abc_40319_new_n3813_), .Y(n193));
OAI21X1 OAI21X1_806 ( .A(IR_REG_0_), .B(IR_REG_1_), .C(IR_REG_2_), .Y(_abc_40319_new_n3815_));
OAI21X1 OAI21X1_807 ( .A(_abc_40319_new_n618_), .B(_abc_40319_new_n875_), .C(_abc_40319_new_n3819_), .Y(n183));
OAI21X1 OAI21X1_808 ( .A(_abc_40319_new_n920_), .B(_abc_40319_new_n1011_), .C(_abc_40319_new_n3821_), .Y(n178));
OAI21X1 OAI21X1_809 ( .A(_abc_40319_new_n2265_), .B(_abc_40319_new_n2263_), .C(_abc_40319_new_n2119_), .Y(_abc_40319_new_n3825_));
OAI21X1 OAI21X1_81 ( .A(IR_REG_0_), .B(_abc_40319_new_n603_), .C(_abc_40319_new_n921_), .Y(_abc_40319_new_n922_));
OAI21X1 OAI21X1_810 ( .A(_abc_40319_new_n1017_), .B(_abc_40319_new_n1046_), .C(_abc_40319_new_n2124_), .Y(_abc_40319_new_n3830_));
OAI21X1 OAI21X1_811 ( .A(_abc_40319_new_n1046_), .B(_abc_40319_new_n2346_), .C(_abc_40319_new_n1017_), .Y(_abc_40319_new_n3831_));
OAI21X1 OAI21X1_812 ( .A(_abc_40319_new_n1592_), .B(_abc_40319_new_n2123_), .C(_abc_40319_new_n2266_), .Y(_abc_40319_new_n3832_));
OAI21X1 OAI21X1_813 ( .A(_abc_40319_new_n3830_), .B(_abc_40319_new_n3126_), .C(_abc_40319_new_n3834_), .Y(_abc_40319_new_n3835_));
OAI21X1 OAI21X1_814 ( .A(_abc_40319_new_n3836_), .B(_abc_40319_new_n3826_), .C(_abc_40319_new_n3824_), .Y(_abc_40319_new_n3837_));
OAI21X1 OAI21X1_815 ( .A(_abc_40319_new_n1504_), .B(_abc_40319_new_n1499_), .C(_abc_40319_new_n1582_), .Y(_abc_40319_new_n3838_));
OAI21X1 OAI21X1_816 ( .A(_abc_40319_new_n3726_), .B(_abc_40319_new_n1341_), .C(_abc_40319_new_n1505_), .Y(_abc_40319_new_n3839_));
OAI21X1 OAI21X1_817 ( .A(_abc_40319_new_n3094_), .B(_abc_40319_new_n3085_), .C(_abc_40319_new_n3839_), .Y(_abc_40319_new_n3840_));
OAI21X1 OAI21X1_818 ( .A(_abc_40319_new_n1505_), .B(_abc_40319_new_n1581_), .C(_abc_40319_new_n3840_), .Y(_abc_40319_new_n3842_));
OAI21X1 OAI21X1_819 ( .A(_abc_40319_new_n749_), .B(_abc_40319_new_n1874_), .C(_abc_40319_new_n743_), .Y(_abc_40319_new_n3845_));
OAI21X1 OAI21X1_82 ( .A(_abc_40319_new_n924_), .B(_abc_40319_new_n923_), .C(_abc_40319_new_n745_), .Y(_abc_40319_new_n925_));
OAI21X1 OAI21X1_820 ( .A(_abc_40319_new_n3836_), .B(_abc_40319_new_n3826_), .C(_abc_40319_new_n3845_), .Y(_abc_40319_new_n3846_));
OAI21X1 OAI21X1_821 ( .A(_abc_40319_new_n2098_), .B(_abc_40319_new_n2101_), .C(_abc_40319_new_n2986_), .Y(_abc_40319_new_n3847_));
OAI21X1 OAI21X1_822 ( .A(_abc_40319_new_n3104_), .B(_abc_40319_new_n1505_), .C(_abc_40319_new_n3847_), .Y(_abc_40319_new_n3848_));
OAI21X1 OAI21X1_823 ( .A(_abc_40319_new_n1582_), .B(_abc_40319_new_n2978_), .C(_abc_40319_new_n2262_), .Y(_abc_40319_new_n3856_));
OAI21X1 OAI21X1_824 ( .A(_abc_40319_new_n1594_), .B(_abc_40319_new_n2960_), .C(nRESET_G), .Y(_abc_40319_new_n3872_));
OAI21X1 OAI21X1_825 ( .A(_abc_40319_new_n1009_), .B(_abc_40319_new_n3870_), .C(_abc_40319_new_n3873_), .Y(_abc_40319_new_n3874_));
OAI21X1 OAI21X1_826 ( .A(_abc_40319_new_n625_), .B(_abc_40319_new_n626_), .C(_abc_40319_new_n674_), .Y(_abc_40319_new_n3877_));
OAI21X1 OAI21X1_827 ( .A(_abc_40319_new_n622_), .B(_abc_40319_new_n572_), .C(_abc_40319_new_n623_), .Y(_abc_40319_new_n3879_));
OAI21X1 OAI21X1_828 ( .A(_abc_40319_new_n619_), .B(_abc_40319_new_n3879_), .C(_abc_40319_new_n3657_), .Y(_abc_40319_new_n3880_));
OAI21X1 OAI21X1_829 ( .A(_abc_40319_new_n655_), .B(_abc_40319_new_n3878_), .C(_abc_40319_new_n3880_), .Y(n338));
OAI21X1 OAI21X1_83 ( .A(_abc_40319_new_n751_), .B(_abc_40319_new_n746_), .C(_abc_40319_new_n914_), .Y(_abc_40319_new_n926_));
OAI21X1 OAI21X1_830 ( .A(_abc_40319_new_n3882_), .B(_abc_40319_new_n3878_), .C(_abc_40319_new_n3883_), .Y(n343));
OAI21X1 OAI21X1_831 ( .A(_abc_40319_new_n615_), .B(_abc_40319_new_n3620_), .C(_abc_40319_new_n973_), .Y(_abc_40319_new_n3885_));
OAI21X1 OAI21X1_832 ( .A(_abc_40319_new_n1760_), .B(_abc_40319_new_n2985_), .C(_abc_40319_new_n3894_), .Y(_abc_40319_new_n3895_));
OAI21X1 OAI21X1_833 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n3897_), .C(_abc_40319_new_n3898_), .Y(n598));
OAI21X1 OAI21X1_834 ( .A(_abc_40319_new_n660_), .B(_abc_40319_new_n922_), .C(_abc_40319_new_n3900_), .Y(_abc_40319_new_n3901_));
OAI21X1 OAI21X1_835 ( .A(_abc_40319_new_n3646_), .B(_abc_40319_new_n3901_), .C(_abc_40319_new_n3889_), .Y(_abc_40319_new_n3902_));
OAI21X1 OAI21X1_836 ( .A(_abc_40319_new_n906_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3903_), .Y(n498));
OAI21X1 OAI21X1_837 ( .A(_abc_40319_new_n1005_), .B(_abc_40319_new_n3629_), .C(_abc_40319_new_n3905_), .Y(_abc_40319_new_n3906_));
OAI21X1 OAI21X1_838 ( .A(_abc_40319_new_n884_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3908_), .Y(n503));
OAI21X1 OAI21X1_839 ( .A(_abc_40319_new_n848_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3912_), .Y(n508));
OAI21X1 OAI21X1_84 ( .A(_abc_40319_new_n908_), .B(_abc_40319_new_n911_), .C(_abc_40319_new_n679_), .Y(_abc_40319_new_n927_));
OAI21X1 OAI21X1_840 ( .A(_abc_40319_new_n3891_), .B(_abc_40319_new_n3606_), .C(_abc_40319_new_n3915_), .Y(_abc_40319_new_n3916_));
OAI21X1 OAI21X1_841 ( .A(_abc_40319_new_n3914_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3918_), .Y(n513));
OAI21X1 OAI21X1_842 ( .A(_abc_40319_new_n804_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3923_), .Y(n518));
OAI21X1 OAI21X1_843 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n3928_), .C(_abc_40319_new_n3929_), .Y(n523));
OAI21X1 OAI21X1_844 ( .A(_abc_40319_new_n952_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3934_), .Y(n528));
OAI21X1 OAI21X1_845 ( .A(_abc_40319_new_n3891_), .B(_abc_40319_new_n3937_), .C(_abc_40319_new_n3539_), .Y(_abc_40319_new_n3938_));
OAI21X1 OAI21X1_846 ( .A(_abc_40319_new_n3936_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3941_), .Y(n533));
OAI21X1 OAI21X1_847 ( .A(_abc_40319_new_n3943_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3947_), .Y(n538));
OAI21X1 OAI21X1_848 ( .A(_abc_40319_new_n3891_), .B(_abc_40319_new_n3503_), .C(_abc_40319_new_n3949_), .Y(_abc_40319_new_n3950_));
OAI21X1 OAI21X1_849 ( .A(_abc_40319_new_n1306_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3953_), .Y(n543));
OAI21X1 OAI21X1_85 ( .A(_abc_40319_new_n549_), .B(_abc_40319_new_n546_), .C(IR_REG_6_), .Y(_abc_40319_new_n939_));
OAI21X1 OAI21X1_850 ( .A(_abc_40319_new_n1397_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3958_), .Y(n548));
OAI21X1 OAI21X1_851 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n3964_), .C(_abc_40319_new_n3965_), .Y(n553));
OAI21X1 OAI21X1_852 ( .A(_abc_40319_new_n1356_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3970_), .Y(n558));
OAI21X1 OAI21X1_853 ( .A(_abc_40319_new_n1334_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3975_), .Y(n563));
OAI21X1 OAI21X1_854 ( .A(_abc_40319_new_n1250_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3980_), .Y(n568));
OAI21X1 OAI21X1_855 ( .A(_abc_40319_new_n3984_), .B(_abc_40319_new_n3402_), .C(_abc_40319_new_n3889_), .Y(_abc_40319_new_n3985_));
OAI21X1 OAI21X1_856 ( .A(_abc_40319_new_n1227_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3986_), .Y(n573));
OAI21X1 OAI21X1_857 ( .A(_abc_40319_new_n1005_), .B(_abc_40319_new_n3382_), .C(_abc_40319_new_n3989_), .Y(_abc_40319_new_n3990_));
OAI21X1 OAI21X1_858 ( .A(_abc_40319_new_n3990_), .B(_abc_40319_new_n3388_), .C(_abc_40319_new_n3889_), .Y(_abc_40319_new_n3991_));
OAI21X1 OAI21X1_859 ( .A(_abc_40319_new_n656_), .B(_abc_40319_new_n3888_), .C(REG0_REG_16_), .Y(_abc_40319_new_n3992_));
OAI21X1 OAI21X1_86 ( .A(_abc_40319_new_n568_), .B(_abc_40319_new_n940_), .C(_abc_40319_new_n941_), .Y(_abc_40319_new_n942_));
OAI21X1 OAI21X1_860 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n1211_), .C(_abc_40319_new_n3369_), .Y(_abc_40319_new_n3995_));
OAI21X1 OAI21X1_861 ( .A(_abc_40319_new_n1200_), .B(_abc_40319_new_n3889_), .C(_abc_40319_new_n3999_), .Y(n583));
OAI21X1 OAI21X1_862 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n4004_), .C(_abc_40319_new_n4005_), .Y(n588));
OAI21X1 OAI21X1_863 ( .A(_abc_40319_new_n4009_), .B(_abc_40319_new_n3312_), .C(_abc_40319_new_n3889_), .Y(_abc_40319_new_n4010_));
OAI21X1 OAI21X1_864 ( .A(_abc_40319_new_n656_), .B(_abc_40319_new_n3888_), .C(REG0_REG_19_), .Y(_abc_40319_new_n4011_));
OAI21X1 OAI21X1_865 ( .A(_abc_40319_new_n2985_), .B(_abc_40319_new_n1137_), .C(_abc_40319_new_n4013_), .Y(_abc_40319_new_n4014_));
OAI21X1 OAI21X1_866 ( .A(_abc_40319_new_n1005_), .B(_abc_40319_new_n3269_), .C(_abc_40319_new_n4015_), .Y(_abc_40319_new_n4016_));
OAI21X1 OAI21X1_867 ( .A(_abc_40319_new_n3273_), .B(_abc_40319_new_n4016_), .C(_abc_40319_new_n3889_), .Y(_abc_40319_new_n4017_));
OAI21X1 OAI21X1_868 ( .A(_abc_40319_new_n656_), .B(_abc_40319_new_n3888_), .C(REG0_REG_21_), .Y(_abc_40319_new_n4018_));
OAI21X1 OAI21X1_869 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n1122_), .C(_abc_40319_new_n4021_), .Y(_abc_40319_new_n4022_));
OAI21X1 OAI21X1_87 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n694_), .C(DATAI_6_), .Y(_abc_40319_new_n943_));
OAI21X1 OAI21X1_870 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n4025_), .C(_abc_40319_new_n4026_), .Y(n608));
OAI21X1 OAI21X1_871 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n4031_), .C(_abc_40319_new_n4032_), .Y(n613));
OAI21X1 OAI21X1_872 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n4037_), .C(_abc_40319_new_n4038_), .Y(n618));
OAI21X1 OAI21X1_873 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n4043_), .C(_abc_40319_new_n4044_), .Y(n623));
OAI21X1 OAI21X1_874 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n4049_), .C(_abc_40319_new_n4050_), .Y(n628));
OAI21X1 OAI21X1_875 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n4058_), .C(_abc_40319_new_n4059_), .Y(n633));
OAI21X1 OAI21X1_876 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n4065_), .C(_abc_40319_new_n4066_), .Y(n638));
OAI21X1 OAI21X1_877 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n2088_), .C(_abc_40319_new_n4068_), .Y(_abc_40319_new_n4069_));
OAI21X1 OAI21X1_878 ( .A(_abc_40319_new_n4069_), .B(_abc_40319_new_n4071_), .C(_abc_40319_new_n3889_), .Y(_abc_40319_new_n4072_));
OAI21X1 OAI21X1_879 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n2096_), .C(_abc_40319_new_n2987_), .Y(_abc_40319_new_n4075_));
OAI21X1 OAI21X1_88 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n942_), .C(_abc_40319_new_n943_), .Y(_abc_40319_new_n944_));
OAI21X1 OAI21X1_880 ( .A(_abc_40319_new_n3890_), .B(_abc_40319_new_n4076_), .C(_abc_40319_new_n4077_), .Y(n648));
OAI21X1 OAI21X1_881 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n1876_), .C(_abc_40319_new_n2987_), .Y(_abc_40319_new_n4080_));
OAI21X1 OAI21X1_882 ( .A(_abc_40319_new_n4080_), .B(_abc_40319_new_n4079_), .C(_abc_40319_new_n3889_), .Y(_abc_40319_new_n4081_));
OAI21X1 OAI21X1_883 ( .A(_abc_40319_new_n3646_), .B(_abc_40319_new_n3901_), .C(_abc_40319_new_n4085_), .Y(_abc_40319_new_n4086_));
OAI21X1 OAI21X1_884 ( .A(_abc_40319_new_n909_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4087_), .Y(n658));
OAI21X1 OAI21X1_885 ( .A(_abc_40319_new_n883_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4089_), .Y(n663));
OAI21X1 OAI21X1_886 ( .A(_abc_40319_new_n4091_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4092_), .Y(n668));
OAI21X1 OAI21X1_887 ( .A(_abc_40319_new_n828_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4094_), .Y(n673));
OAI21X1 OAI21X1_888 ( .A(_abc_40319_new_n800_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4096_), .Y(n678));
OAI21X1 OAI21X1_889 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n3928_), .C(_abc_40319_new_n4098_), .Y(n683));
OAI21X1 OAI21X1_89 ( .A(_abc_40319_new_n751_), .B(_abc_40319_new_n746_), .C(_abc_40319_new_n944_), .Y(_abc_40319_new_n956_));
OAI21X1 OAI21X1_890 ( .A(_abc_40319_new_n945_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4100_), .Y(n688));
OAI21X1 OAI21X1_891 ( .A(_abc_40319_new_n2653_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4102_), .Y(n693));
OAI21X1 OAI21X1_892 ( .A(_abc_40319_new_n2672_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4104_), .Y(n698));
OAI21X1 OAI21X1_893 ( .A(_abc_40319_new_n1298_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4106_), .Y(n703));
OAI21X1 OAI21X1_894 ( .A(_abc_40319_new_n1394_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4108_), .Y(n708));
OAI21X1 OAI21X1_895 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n3964_), .C(_abc_40319_new_n4110_), .Y(n713));
OAI21X1 OAI21X1_896 ( .A(_abc_40319_new_n1353_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4112_), .Y(n718));
OAI21X1 OAI21X1_897 ( .A(_abc_40319_new_n1326_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4114_), .Y(n723));
OAI21X1 OAI21X1_898 ( .A(_abc_40319_new_n1252_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4116_), .Y(n728));
OAI21X1 OAI21X1_899 ( .A(_abc_40319_new_n3984_), .B(_abc_40319_new_n3402_), .C(_abc_40319_new_n4085_), .Y(_abc_40319_new_n4118_));
OAI21X1 OAI21X1_9 ( .A(_abc_40319_new_n555_), .B(_abc_40319_new_n604_), .C(IR_REG_22_), .Y(_abc_40319_new_n605_));
OAI21X1 OAI21X1_90 ( .A(_abc_40319_new_n950_), .B(_abc_40319_new_n953_), .C(_abc_40319_new_n679_), .Y(_abc_40319_new_n957_));
OAI21X1 OAI21X1_900 ( .A(_abc_40319_new_n1224_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4119_), .Y(n733));
OAI21X1 OAI21X1_901 ( .A(_abc_40319_new_n3990_), .B(_abc_40319_new_n3388_), .C(_abc_40319_new_n4085_), .Y(_abc_40319_new_n4121_));
OAI21X1 OAI21X1_902 ( .A(_abc_40319_new_n1179_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4122_), .Y(n738));
OAI21X1 OAI21X1_903 ( .A(_abc_40319_new_n1199_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4124_), .Y(n743));
OAI21X1 OAI21X1_904 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n4004_), .C(_abc_40319_new_n4126_), .Y(n748));
OAI21X1 OAI21X1_905 ( .A(_abc_40319_new_n4009_), .B(_abc_40319_new_n3312_), .C(_abc_40319_new_n4085_), .Y(_abc_40319_new_n4128_));
OAI21X1 OAI21X1_906 ( .A(_abc_40319_new_n1430_), .B(_abc_40319_new_n4085_), .C(_abc_40319_new_n4129_), .Y(n753));
OAI21X1 OAI21X1_907 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n3897_), .C(_abc_40319_new_n4131_), .Y(n758));
OAI21X1 OAI21X1_908 ( .A(_abc_40319_new_n3273_), .B(_abc_40319_new_n4016_), .C(_abc_40319_new_n4085_), .Y(_abc_40319_new_n4133_));
OAI21X1 OAI21X1_909 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n4025_), .C(_abc_40319_new_n4136_), .Y(n768));
OAI21X1 OAI21X1_91 ( .A(_abc_40319_new_n758_), .B(_abc_40319_new_n959_), .C(_abc_40319_new_n956_), .Y(_abc_40319_new_n960_));
OAI21X1 OAI21X1_910 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n4031_), .C(_abc_40319_new_n4138_), .Y(n773));
OAI21X1 OAI21X1_911 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n4037_), .C(_abc_40319_new_n4140_), .Y(n778));
OAI21X1 OAI21X1_912 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n4043_), .C(_abc_40319_new_n4142_), .Y(n783));
OAI21X1 OAI21X1_913 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n4049_), .C(_abc_40319_new_n4144_), .Y(n788));
OAI21X1 OAI21X1_914 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n4058_), .C(_abc_40319_new_n4146_), .Y(n793));
OAI21X1 OAI21X1_915 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n4065_), .C(_abc_40319_new_n4148_), .Y(n798));
OAI21X1 OAI21X1_916 ( .A(_abc_40319_new_n4069_), .B(_abc_40319_new_n4071_), .C(_abc_40319_new_n4085_), .Y(_abc_40319_new_n4150_));
OAI21X1 OAI21X1_917 ( .A(_abc_40319_new_n4084_), .B(_abc_40319_new_n4076_), .C(_abc_40319_new_n4153_), .Y(n808));
OAI21X1 OAI21X1_918 ( .A(_abc_40319_new_n4080_), .B(_abc_40319_new_n4079_), .C(_abc_40319_new_n4085_), .Y(_abc_40319_new_n4155_));
OAI21X1 OAI21X1_919 ( .A(_abc_40319_new_n912_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4159_), .Y(n1058));
OAI21X1 OAI21X1_92 ( .A(_abc_40319_new_n962_), .B(_abc_40319_new_n937_), .C(_abc_40319_new_n966_), .Y(_abc_40319_new_n967_));
OAI21X1 OAI21X1_920 ( .A(_abc_40319_new_n897_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4161_), .Y(n1062));
OAI21X1 OAI21X1_921 ( .A(_abc_40319_new_n855_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4163_), .Y(n1066));
OAI21X1 OAI21X1_922 ( .A(_abc_40319_new_n865_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4165_), .Y(n1070));
OAI21X1 OAI21X1_923 ( .A(_abc_40319_new_n1556_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4167_), .Y(n1074));
OAI21X1 OAI21X1_924 ( .A(_abc_40319_new_n788_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4169_), .Y(n1078));
OAI21X1 OAI21X1_925 ( .A(_abc_40319_new_n959_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4171_), .Y(n1082));
OAI21X1 OAI21X1_926 ( .A(_abc_40319_new_n759_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4173_), .Y(n1086));
OAI21X1 OAI21X1_927 ( .A(_abc_40319_new_n988_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4175_), .Y(n1090));
OAI21X1 OAI21X1_928 ( .A(_abc_40319_new_n1308_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4177_), .Y(n1094));
OAI21X1 OAI21X1_929 ( .A(_abc_40319_new_n1401_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4179_), .Y(n1098));
OAI21X1 OAI21X1_93 ( .A(_abc_40319_new_n762_), .B(_abc_40319_new_n968_), .C(_abc_40319_new_n969_), .Y(_abc_40319_new_n970_));
OAI21X1 OAI21X1_930 ( .A(_abc_40319_new_n1379_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4181_), .Y(n1102));
OAI21X1 OAI21X1_931 ( .A(_abc_40319_new_n1796_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4183_), .Y(n1106));
OAI21X1 OAI21X1_932 ( .A(_abc_40319_new_n1514_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4185_), .Y(n1110));
OAI21X1 OAI21X1_933 ( .A(_abc_40319_new_n1258_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4187_), .Y(n1114));
OAI21X1 OAI21X1_934 ( .A(_abc_40319_new_n1516_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4189_), .Y(n1118));
OAI21X1 OAI21X1_935 ( .A(_abc_40319_new_n1700_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4191_), .Y(n1122));
OAI21X1 OAI21X1_936 ( .A(_abc_40319_new_n1208_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4193_), .Y(n1126));
OAI21X1 OAI21X1_937 ( .A(_abc_40319_new_n1156_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4195_), .Y(n1130));
OAI21X1 OAI21X1_938 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1759_), .C(_abc_40319_new_n4197_), .Y(n1134));
OAI21X1 OAI21X1_939 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1567_), .C(_abc_40319_new_n4199_), .Y(n1138));
OAI21X1 OAI21X1_94 ( .A(_abc_40319_new_n762_), .B(_abc_40319_new_n967_), .C(_abc_40319_new_n970_), .Y(_abc_40319_new_n971_));
OAI21X1 OAI21X1_940 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1760_), .C(_abc_40319_new_n4201_), .Y(n1142));
OAI21X1 OAI21X1_941 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1137_), .C(_abc_40319_new_n4203_), .Y(n1146));
OAI21X1 OAI21X1_942 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1710_), .C(_abc_40319_new_n4205_), .Y(n1150));
OAI21X1 OAI21X1_943 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1093_), .C(_abc_40319_new_n4207_), .Y(n1154));
OAI21X1 OAI21X1_944 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1078_), .C(_abc_40319_new_n4209_), .Y(n1158));
OAI21X1 OAI21X1_945 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1496_), .C(_abc_40319_new_n4211_), .Y(n1162));
OAI21X1 OAI21X1_946 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1592_), .C(_abc_40319_new_n4213_), .Y(n1166));
OAI21X1 OAI21X1_947 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1505_), .C(_abc_40319_new_n4215_), .Y(n1170));
OAI21X1 OAI21X1_948 ( .A(_abc_40319_new_n4158_), .B(_abc_40319_new_n1598_), .C(_abc_40319_new_n4217_), .Y(n1174));
OAI21X1 OAI21X1_949 ( .A(_abc_40319_new_n2102_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4219_), .Y(n1178));
OAI21X1 OAI21X1_95 ( .A(_abc_40319_new_n735_), .B(_abc_40319_new_n946_), .C(_abc_40319_new_n980_), .Y(_abc_40319_new_n981_));
OAI21X1 OAI21X1_950 ( .A(_abc_40319_new_n1882_), .B(_abc_40319_new_n4158_), .C(_abc_40319_new_n4221_), .Y(n1182));
OAI21X1 OAI21X1_96 ( .A(_abc_40319_new_n593_), .B(_abc_40319_new_n602_), .C(_abc_40319_new_n658_), .Y(_abc_40319_new_n989_));
OAI21X1 OAI21X1_97 ( .A(_abc_40319_new_n669_), .B(_abc_40319_new_n658_), .C(_abc_40319_new_n672_), .Y(_abc_40319_new_n998_));
OAI21X1 OAI21X1_98 ( .A(_abc_40319_new_n997_), .B(_abc_40319_new_n998_), .C(STATE_REG), .Y(_abc_40319_new_n999_));
OAI21X1 OAI21X1_99 ( .A(_abc_40319_new_n658_), .B(_abc_40319_new_n996_), .C(_abc_40319_new_n999_), .Y(_abc_40319_new_n1000_));
OAI22X1 OAI22X1_1 ( .A(_abc_40319_new_n593_), .B(_abc_40319_new_n602_), .C(_abc_40319_new_n586_), .D(_abc_40319_new_n592_), .Y(_abc_40319_new_n603_));
OAI22X1 OAI22X1_10 ( .A(_abc_40319_new_n988_), .B(_abc_40319_new_n989_), .C(_abc_40319_new_n959_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n990_));
OAI22X1 OAI22X1_11 ( .A(_abc_40319_new_n758_), .B(_abc_40319_new_n1070_), .C(_abc_40319_new_n905_), .D(_abc_40319_new_n1078_), .Y(_abc_40319_new_n1079_));
OAI22X1 OAI22X1_12 ( .A(_abc_40319_new_n1096_), .B(_abc_40319_new_n1084_), .C(_abc_40319_new_n758_), .D(_abc_40319_new_n1093_), .Y(_abc_40319_new_n1097_));
OAI22X1 OAI22X1_13 ( .A(_abc_40319_new_n1096_), .B(_abc_40319_new_n1122_), .C(_abc_40319_new_n758_), .D(_abc_40319_new_n1137_), .Y(_abc_40319_new_n1138_));
OAI22X1 OAI22X1_14 ( .A(_abc_40319_new_n1096_), .B(_abc_40319_new_n1159_), .C(_abc_40319_new_n758_), .D(_abc_40319_new_n1156_), .Y(_abc_40319_new_n1160_));
OAI22X1 OAI22X1_15 ( .A(_abc_40319_new_n1179_), .B(_abc_40319_new_n802_), .C(_abc_40319_new_n778_), .D(_abc_40319_new_n1187_), .Y(_abc_40319_new_n1188_));
OAI22X1 OAI22X1_16 ( .A(_abc_40319_new_n1200_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n1199_), .D(_abc_40319_new_n802_), .Y(_abc_40319_new_n1201_));
OAI22X1 OAI22X1_17 ( .A(_abc_40319_new_n1202_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n778_), .D(_abc_40319_new_n1206_), .Y(_abc_40319_new_n1207_));
OAI22X1 OAI22X1_18 ( .A(_abc_40319_new_n1096_), .B(_abc_40319_new_n1211_), .C(_abc_40319_new_n758_), .D(_abc_40319_new_n1208_), .Y(_abc_40319_new_n1212_));
OAI22X1 OAI22X1_19 ( .A(_abc_40319_new_n1225_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n1224_), .D(_abc_40319_new_n802_), .Y(_abc_40319_new_n1226_));
OAI22X1 OAI22X1_2 ( .A(_abc_40319_new_n776_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n781_), .D(_abc_40319_new_n778_), .Y(_abc_40319_new_n782_));
OAI22X1 OAI22X1_20 ( .A(_abc_40319_new_n1249_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n1250_), .D(_abc_40319_new_n777_), .Y(_abc_40319_new_n1251_));
OAI22X1 OAI22X1_21 ( .A(_abc_40319_new_n758_), .B(_abc_40319_new_n1258_), .C(_abc_40319_new_n1261_), .D(_abc_40319_new_n1096_), .Y(_abc_40319_new_n1262_));
OAI22X1 OAI22X1_22 ( .A(_abc_40319_new_n1305_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n1306_), .D(_abc_40319_new_n777_), .Y(_abc_40319_new_n1307_));
OAI22X1 OAI22X1_23 ( .A(_abc_40319_new_n1326_), .B(_abc_40319_new_n802_), .C(_abc_40319_new_n778_), .D(_abc_40319_new_n1331_), .Y(_abc_40319_new_n1332_));
OAI22X1 OAI22X1_24 ( .A(_abc_40319_new_n1333_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n1334_), .D(_abc_40319_new_n777_), .Y(_abc_40319_new_n1335_));
OAI22X1 OAI22X1_25 ( .A(_abc_40319_new_n1354_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n1353_), .D(_abc_40319_new_n802_), .Y(_abc_40319_new_n1355_));
OAI22X1 OAI22X1_26 ( .A(_abc_40319_new_n1373_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n1372_), .D(_abc_40319_new_n802_), .Y(_abc_40319_new_n1374_));
OAI22X1 OAI22X1_27 ( .A(_abc_40319_new_n758_), .B(_abc_40319_new_n1379_), .C(_abc_40319_new_n1370_), .D(_abc_40319_new_n1096_), .Y(_abc_40319_new_n1383_));
OAI22X1 OAI22X1_28 ( .A(_abc_40319_new_n1397_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n1399_), .D(_abc_40319_new_n778_), .Y(_abc_40319_new_n1400_));
OAI22X1 OAI22X1_29 ( .A(_abc_40319_new_n979_), .B(_abc_40319_new_n1496_), .C(_abc_40319_new_n989_), .D(_abc_40319_new_n1505_), .Y(_abc_40319_new_n1506_));
OAI22X1 OAI22X1_3 ( .A(_abc_40319_new_n801_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n800_), .D(_abc_40319_new_n802_), .Y(_abc_40319_new_n803_));
OAI22X1 OAI22X1_30 ( .A(_abc_40319_new_n989_), .B(_abc_40319_new_n1093_), .C(_abc_40319_new_n1137_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1529_));
OAI22X1 OAI22X1_31 ( .A(_abc_40319_new_n989_), .B(_abc_40319_new_n1379_), .C(_abc_40319_new_n1308_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1539_));
OAI22X1 OAI22X1_32 ( .A(_abc_40319_new_n1556_), .B(_abc_40319_new_n989_), .C(_abc_40319_new_n855_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1557_));
OAI22X1 OAI22X1_33 ( .A(_abc_40319_new_n1096_), .B(_abc_40319_new_n1581_), .C(_abc_40319_new_n758_), .D(_abc_40319_new_n1505_), .Y(_abc_40319_new_n1584_));
OAI22X1 OAI22X1_34 ( .A(_abc_40319_new_n1594_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n778_), .D(_abc_40319_new_n1595_), .Y(_abc_40319_new_n1596_));
OAI22X1 OAI22X1_35 ( .A(_abc_40319_new_n979_), .B(_abc_40319_new_n1592_), .C(_abc_40319_new_n989_), .D(_abc_40319_new_n1598_), .Y(_abc_40319_new_n1599_));
OAI22X1 OAI22X1_36 ( .A(_abc_40319_new_n989_), .B(_abc_40319_new_n1308_), .C(_abc_40319_new_n759_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1614_));
OAI22X1 OAI22X1_37 ( .A(_abc_40319_new_n855_), .B(_abc_40319_new_n989_), .C(_abc_40319_new_n912_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1623_));
OAI22X1 OAI22X1_38 ( .A(_abc_40319_new_n658_), .B(_abc_40319_new_n1463_), .C(_abc_40319_new_n1137_), .D(_abc_40319_new_n989_), .Y(_abc_40319_new_n1630_));
OAI22X1 OAI22X1_39 ( .A(_abc_40319_new_n979_), .B(_abc_40319_new_n1093_), .C(_abc_40319_new_n989_), .D(_abc_40319_new_n1496_), .Y(_abc_40319_new_n1667_));
OAI22X1 OAI22X1_4 ( .A(_abc_40319_new_n827_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n828_), .D(_abc_40319_new_n802_), .Y(_abc_40319_new_n829_));
OAI22X1 OAI22X1_40 ( .A(_abc_40319_new_n989_), .B(_abc_40319_new_n1208_), .C(_abc_40319_new_n1516_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1679_));
OAI22X1 OAI22X1_41 ( .A(_abc_40319_new_n959_), .B(_abc_40319_new_n989_), .C(_abc_40319_new_n1556_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1688_));
OAI22X1 OAI22X1_42 ( .A(_abc_40319_new_n989_), .B(_abc_40319_new_n1156_), .C(_abc_40319_new_n1700_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1701_));
OAI22X1 OAI22X1_43 ( .A(_abc_40319_new_n979_), .B(_abc_40319_new_n1710_), .C(_abc_40319_new_n989_), .D(_abc_40319_new_n1078_), .Y(_abc_40319_new_n1711_));
OAI22X1 OAI22X1_44 ( .A(_abc_40319_new_n1750_), .B(_abc_40319_new_n658_), .C(_abc_40319_new_n897_), .D(_abc_40319_new_n989_), .Y(_abc_40319_new_n1751_));
OAI22X1 OAI22X1_45 ( .A(_abc_40319_new_n989_), .B(_abc_40319_new_n1760_), .C(_abc_40319_new_n1759_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1761_));
OAI22X1 OAI22X1_46 ( .A(_abc_40319_new_n658_), .B(_abc_40319_new_n1331_), .C(_abc_40319_new_n1258_), .D(_abc_40319_new_n989_), .Y(_abc_40319_new_n1773_));
OAI22X1 OAI22X1_47 ( .A(_abc_40319_new_n989_), .B(_abc_40319_new_n1710_), .C(_abc_40319_new_n1760_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1786_));
OAI22X1 OAI22X1_48 ( .A(_abc_40319_new_n989_), .B(_abc_40319_new_n1759_), .C(_abc_40319_new_n1208_), .D(_abc_40319_new_n979_), .Y(_abc_40319_new_n1822_));
OAI22X1 OAI22X1_49 ( .A(_abc_40319_new_n979_), .B(_abc_40319_new_n1078_), .C(_abc_40319_new_n989_), .D(_abc_40319_new_n1592_), .Y(_abc_40319_new_n1850_));
OAI22X1 OAI22X1_5 ( .A(_abc_40319_new_n847_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n848_), .D(_abc_40319_new_n777_), .Y(_abc_40319_new_n849_));
OAI22X1 OAI22X1_50 ( .A(_abc_40319_new_n1897_), .B(_abc_40319_new_n1893_), .C(_abc_40319_new_n1913_), .D(_abc_40319_new_n1915_), .Y(_abc_40319_new_n1916_));
OAI22X1 OAI22X1_51 ( .A(_abc_40319_new_n698_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n740_), .Y(_abc_40319_new_n1928_));
OAI22X1 OAI22X1_52 ( .A(_abc_40319_new_n944_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n954_), .Y(_abc_40319_new_n1930_));
OAI22X1 OAI22X1_53 ( .A(_abc_40319_new_n1393_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n1402_), .Y(_abc_40319_new_n1948_));
OAI22X1 OAI22X1_54 ( .A(_abc_40319_new_n1276_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n987_), .Y(_abc_40319_new_n1963_));
OAI22X1 OAI22X1_55 ( .A(_abc_40319_new_n1934_), .B(_abc_40319_new_n1930_), .C(_abc_40319_new_n1928_), .D(_abc_40319_new_n1927_), .Y(_abc_40319_new_n1966_));
OAI22X1 OAI22X1_56 ( .A(_abc_40319_new_n1325_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n1336_), .Y(_abc_40319_new_n1977_));
OAI22X1 OAI22X1_57 ( .A(_abc_40319_new_n1360_), .B(_abc_40319_new_n1894_), .C(_abc_40319_new_n1888_), .D(_abc_40319_new_n1352_), .Y(_abc_40319_new_n1978_));
OAI22X1 OAI22X1_58 ( .A(_abc_40319_new_n1371_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n1380_), .Y(_abc_40319_new_n1989_));
OAI22X1 OAI22X1_59 ( .A(_abc_40319_new_n1947_), .B(_abc_40319_new_n1948_), .C(_abc_40319_new_n1989_), .D(_abc_40319_new_n1988_), .Y(_abc_40319_new_n1990_));
OAI22X1 OAI22X1_6 ( .A(_abc_40319_new_n884_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n883_), .D(_abc_40319_new_n802_), .Y(_abc_40319_new_n885_));
OAI22X1 OAI22X1_60 ( .A(_abc_40319_new_n1248_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n1259_), .Y(_abc_40319_new_n2000_));
OAI22X1 OAI22X1_61 ( .A(_abc_40319_new_n1873_), .B(_abc_40319_new_n1865_), .C(_abc_40319_new_n580_), .D(_abc_40319_new_n1258_), .Y(_abc_40319_new_n2006_));
OAI22X1 OAI22X1_62 ( .A(_abc_40319_new_n1175_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n1189_), .Y(_abc_40319_new_n2013_));
OAI22X1 OAI22X1_63 ( .A(_abc_40319_new_n1198_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n1209_), .Y(_abc_40319_new_n2019_));
OAI22X1 OAI22X1_64 ( .A(_abc_40319_new_n2012_), .B(_abc_40319_new_n2013_), .C(_abc_40319_new_n2018_), .D(_abc_40319_new_n2019_), .Y(_abc_40319_new_n2020_));
OAI22X1 OAI22X1_65 ( .A(_abc_40319_new_n1873_), .B(_abc_40319_new_n1159_), .C(_abc_40319_new_n580_), .D(_abc_40319_new_n1208_), .Y(_abc_40319_new_n2023_));
OAI22X1 OAI22X1_66 ( .A(_abc_40319_new_n1443_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n1452_), .Y(_abc_40319_new_n2038_));
OAI22X1 OAI22X1_67 ( .A(_abc_40319_new_n1460_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n1469_), .Y(_abc_40319_new_n2042_));
OAI22X1 OAI22X1_68 ( .A(_abc_40319_new_n2037_), .B(_abc_40319_new_n2038_), .C(_abc_40319_new_n2041_), .D(_abc_40319_new_n2042_), .Y(_abc_40319_new_n2043_));
OAI22X1 OAI22X1_69 ( .A(_abc_40319_new_n1873_), .B(_abc_40319_new_n1122_), .C(_abc_40319_new_n580_), .D(_abc_40319_new_n1760_), .Y(_abc_40319_new_n2046_));
OAI22X1 OAI22X1_7 ( .A(_abc_40319_new_n906_), .B(_abc_40319_new_n777_), .C(_abc_40319_new_n907_), .D(_abc_40319_new_n774_), .Y(_abc_40319_new_n908_));
OAI22X1 OAI22X1_70 ( .A(_abc_40319_new_n1080_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n1077_), .Y(_abc_40319_new_n2065_));
OAI22X1 OAI22X1_71 ( .A(_abc_40319_new_n2057_), .B(_abc_40319_new_n2059_), .C(_abc_40319_new_n2065_), .D(_abc_40319_new_n2064_), .Y(_abc_40319_new_n2066_));
OAI22X1 OAI22X1_72 ( .A(_abc_40319_new_n580_), .B(_abc_40319_new_n1496_), .C(_abc_40319_new_n1888_), .D(_abc_40319_new_n1592_), .Y(_abc_40319_new_n2075_));
OAI22X1 OAI22X1_73 ( .A(_abc_40319_new_n1582_), .B(_abc_40319_new_n1888_), .C(_abc_40319_new_n1894_), .D(_abc_40319_new_n1580_), .Y(_abc_40319_new_n2083_));
OAI22X1 OAI22X1_74 ( .A(_abc_40319_new_n2076_), .B(_abc_40319_new_n2077_), .C(_abc_40319_new_n2082_), .D(_abc_40319_new_n2084_), .Y(_abc_40319_new_n2085_));
OAI22X1 OAI22X1_75 ( .A(_abc_40319_new_n1888_), .B(_abc_40319_new_n1598_), .C(_abc_40319_new_n580_), .D(_abc_40319_new_n1505_), .Y(_abc_40319_new_n2090_));
OAI22X1 OAI22X1_76 ( .A(_abc_40319_new_n1885_), .B(_abc_40319_new_n1886_), .C(_abc_40319_new_n2105_), .D(_abc_40319_new_n2109_), .Y(_abc_40319_new_n2113_));
OAI22X1 OAI22X1_77 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n837_), .C(_abc_40319_new_n2573_), .D(_abc_40319_new_n694_), .Y(_abc_40319_new_n2574_));
OAI22X1 OAI22X1_78 ( .A(_abc_40319_new_n2566_), .B(_abc_40319_new_n2574_), .C(_abc_40319_new_n2542_), .D(_abc_40319_new_n2543_), .Y(_abc_40319_new_n2575_));
OAI22X1 OAI22X1_79 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n749_), .C(_abc_40319_new_n2942_), .D(_abc_40319_new_n2946_), .Y(_abc_40319_new_n2947_));
OAI22X1 OAI22X1_8 ( .A(_abc_40319_new_n945_), .B(_abc_40319_new_n802_), .C(_abc_40319_new_n949_), .D(_abc_40319_new_n778_), .Y(_abc_40319_new_n950_));
OAI22X1 OAI22X1_80 ( .A(_abc_40319_new_n1570_), .B(_abc_40319_new_n1759_), .C(_abc_40319_new_n1442_), .D(_abc_40319_new_n1567_), .Y(_abc_40319_new_n3013_));
OAI22X1 OAI22X1_81 ( .A(_abc_40319_new_n1460_), .B(_abc_40319_new_n1469_), .C(_abc_40319_new_n3015_), .D(_abc_40319_new_n3012_), .Y(_abc_40319_new_n3016_));
OAI22X1 OAI22X1_82 ( .A(_abc_40319_new_n1496_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3128_), .D(_abc_40319_new_n3129_), .Y(_abc_40319_new_n3130_));
OAI22X1 OAI22X1_83 ( .A(_abc_40319_new_n1078_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3155_), .D(_abc_40319_new_n3156_), .Y(_abc_40319_new_n3157_));
OAI22X1 OAI22X1_84 ( .A(_abc_40319_new_n1093_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3185_), .D(_abc_40319_new_n3186_), .Y(_abc_40319_new_n3187_));
OAI22X1 OAI22X1_85 ( .A(_abc_40319_new_n1009_), .B(_abc_40319_new_n1110_), .C(_abc_40319_new_n1093_), .D(_abc_40319_new_n3164_), .Y(_abc_40319_new_n3223_));
OAI22X1 OAI22X1_86 ( .A(_abc_40319_new_n1009_), .B(_abc_40319_new_n1128_), .C(_abc_40319_new_n1710_), .D(_abc_40319_new_n3164_), .Y(_abc_40319_new_n3246_));
OAI22X1 OAI22X1_87 ( .A(_abc_40319_new_n1700_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3155_), .D(_abc_40319_new_n3362_), .Y(_abc_40319_new_n3363_));
OAI22X1 OAI22X1_88 ( .A(_abc_40319_new_n788_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3100_), .D(_abc_40319_new_n3550_), .Y(_abc_40319_new_n3551_));
OAI22X1 OAI22X1_89 ( .A(_abc_40319_new_n759_), .B(_abc_40319_new_n2985_), .C(_abc_40319_new_n2246_), .D(_abc_40319_new_n994_), .Y(_abc_40319_new_n3557_));
OAI22X1 OAI22X1_9 ( .A(_abc_40319_new_n951_), .B(_abc_40319_new_n774_), .C(_abc_40319_new_n952_), .D(_abc_40319_new_n777_), .Y(_abc_40319_new_n953_));
OAI22X1 OAI22X1_90 ( .A(_abc_40319_new_n1556_), .B(_abc_40319_new_n3104_), .C(_abc_40319_new_n3100_), .D(_abc_40319_new_n3583_), .Y(_abc_40319_new_n3584_));
OAI22X1 OAI22X1_91 ( .A(_abc_40319_new_n1938_), .B(_abc_40319_new_n994_), .C(_abc_40319_new_n2985_), .D(_abc_40319_new_n959_), .Y(_abc_40319_new_n3589_));
OAI22X1 OAI22X1_92 ( .A(_abc_40319_new_n825_), .B(_abc_40319_new_n994_), .C(_abc_40319_new_n2985_), .D(_abc_40319_new_n1556_), .Y(_abc_40319_new_n3603_));
OAI22X1 OAI22X1_93 ( .A(REG2_REG_0_), .B(_abc_40319_new_n2960_), .C(_abc_40319_new_n3646_), .D(_abc_40319_new_n3648_), .Y(_abc_40319_new_n3649_));
OAI22X1 OAI22X1_94 ( .A(_abc_40319_new_n994_), .B(_abc_40319_new_n2196_), .C(_abc_40319_new_n2985_), .D(_abc_40319_new_n1208_), .Y(_abc_40319_new_n3988_));
OR2X2 OR2X2_1 ( .A(IR_REG_31_), .B(IR_REG_21_), .Y(_abc_40319_new_n610_));
OR2X2 OR2X2_10 ( .A(_abc_40319_new_n1119_), .B(_abc_40319_new_n1116_), .Y(_abc_40319_new_n1120_));
OR2X2 OR2X2_11 ( .A(_abc_40319_new_n1129_), .B(_abc_40319_new_n1134_), .Y(_abc_40319_new_n1135_));
OR2X2 OR2X2_12 ( .A(_abc_40319_new_n1026_), .B(_abc_40319_new_n1027_), .Y(_abc_40319_new_n1180_));
OR2X2 OR2X2_13 ( .A(_abc_40319_new_n1188_), .B(_abc_40319_new_n1178_), .Y(_abc_40319_new_n1189_));
OR2X2 OR2X2_14 ( .A(_abc_40319_new_n1232_), .B(_abc_40319_new_n1226_), .Y(_abc_40319_new_n1233_));
OR2X2 OR2X2_15 ( .A(_abc_40319_new_n1264_), .B(_abc_40319_new_n1260_), .Y(_abc_40319_new_n1265_));
OR2X2 OR2X2_16 ( .A(_abc_40319_new_n1279_), .B(_abc_40319_new_n1277_), .Y(_abc_40319_new_n1284_));
OR2X2 OR2X2_17 ( .A(_abc_40319_new_n1332_), .B(_abc_40319_new_n1335_), .Y(_abc_40319_new_n1336_));
OR2X2 OR2X2_18 ( .A(_abc_40319_new_n1290_), .B(_abc_40319_new_n1318_), .Y(_abc_40319_new_n1342_));
OR2X2 OR2X2_19 ( .A(_abc_40319_new_n1359_), .B(_abc_40319_new_n1355_), .Y(_abc_40319_new_n1360_));
OR2X2 OR2X2_2 ( .A(D_REG_30_), .B(D_REG_9_), .Y(_abc_40319_new_n631_));
OR2X2 OR2X2_20 ( .A(_abc_40319_new_n1436_), .B(_abc_40319_new_n1431_), .Y(_abc_40319_new_n1437_));
OR2X2 OR2X2_21 ( .A(_abc_40319_new_n1447_), .B(_abc_40319_new_n1451_), .Y(_abc_40319_new_n1452_));
OR2X2 OR2X2_22 ( .A(_abc_40319_new_n1464_), .B(_abc_40319_new_n1468_), .Y(_abc_40319_new_n1469_));
OR2X2 OR2X2_23 ( .A(_abc_40319_new_n1083_), .B(_abc_40319_new_n1490_), .Y(_abc_40319_new_n1491_));
OR2X2 OR2X2_24 ( .A(_abc_40319_new_n1040_), .B(REG3_REG_28_), .Y(_abc_40319_new_n1498_));
OR2X2 OR2X2_25 ( .A(_abc_40319_new_n1384_), .B(_abc_40319_new_n1382_), .Y(_abc_40319_new_n1646_));
OR2X2 OR2X2_26 ( .A(_abc_40319_new_n1082_), .B(_abc_40319_new_n1079_), .Y(_abc_40319_new_n1660_));
OR2X2 OR2X2_27 ( .A(_abc_40319_new_n1834_), .B(_abc_40319_new_n1835_), .Y(_abc_40319_new_n1836_));
OR2X2 OR2X2_28 ( .A(_abc_40319_new_n1920_), .B(_abc_40319_new_n1918_), .Y(_abc_40319_new_n1923_));
OR2X2 OR2X2_29 ( .A(_abc_40319_new_n1927_), .B(_abc_40319_new_n1928_), .Y(_abc_40319_new_n1929_));
OR2X2 OR2X2_3 ( .A(IR_REG_31_), .B(IR_REG_29_), .Y(_abc_40319_new_n709_));
OR2X2 OR2X2_30 ( .A(_abc_40319_new_n1930_), .B(_abc_40319_new_n1934_), .Y(_abc_40319_new_n1935_));
OR2X2 OR2X2_31 ( .A(_abc_40319_new_n1987_), .B(_abc_40319_new_n1985_), .Y(_abc_40319_new_n1988_));
OR2X2 OR2X2_32 ( .A(_abc_40319_new_n2269_), .B(_abc_40319_new_n2117_), .Y(_abc_40319_new_n2270_));
OR2X2 OR2X2_33 ( .A(_abc_40319_new_n2132_), .B(_abc_40319_new_n2137_), .Y(_abc_40319_new_n2314_));
OR2X2 OR2X2_34 ( .A(_abc_40319_new_n2323_), .B(_abc_40319_new_n2321_), .Y(_abc_40319_new_n2324_));
OR2X2 OR2X2_35 ( .A(_abc_40319_new_n2369_), .B(_abc_40319_new_n2394_), .Y(_abc_40319_new_n2466_));
OR2X2 OR2X2_36 ( .A(_abc_40319_new_n2514_), .B(_abc_40319_new_n2451_), .Y(_abc_40319_new_n2515_));
OR2X2 OR2X2_37 ( .A(_abc_40319_new_n3055_), .B(_abc_40319_new_n2194_), .Y(_abc_40319_new_n3062_));
OR2X2 OR2X2_38 ( .A(_abc_40319_new_n3106_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3107_));
OR2X2 OR2X2_39 ( .A(_abc_40319_new_n3122_), .B(_abc_40319_new_n3119_), .Y(_abc_40319_new_n3123_));
OR2X2 OR2X2_4 ( .A(_abc_40319_new_n775_), .B(_abc_40319_new_n782_), .Y(_abc_40319_new_n783_));
OR2X2 OR2X2_40 ( .A(_abc_40319_new_n3131_), .B(_abc_40319_new_n2990_), .Y(_abc_40319_new_n3132_));
OR2X2 OR2X2_41 ( .A(_abc_40319_new_n3174_), .B(_abc_40319_new_n2130_), .Y(_abc_40319_new_n3176_));
OR2X2 OR2X2_42 ( .A(_abc_40319_new_n2496_), .B(_abc_40319_new_n2321_), .Y(_abc_40319_new_n3179_));
OR2X2 OR2X2_43 ( .A(_abc_40319_new_n3244_), .B(_abc_40319_new_n3223_), .Y(n933));
OR2X2 OR2X2_44 ( .A(_abc_40319_new_n2960_), .B(REG2_REG_22_), .Y(_abc_40319_new_n3256_));
OR2X2 OR2X2_45 ( .A(_abc_40319_new_n3263_), .B(_abc_40319_new_n3246_), .Y(n928));
OR2X2 OR2X2_46 ( .A(_abc_40319_new_n3300_), .B(_abc_40319_new_n2961_), .Y(_abc_40319_new_n3301_));
OR2X2 OR2X2_47 ( .A(_abc_40319_new_n3419_), .B(_abc_40319_new_n3421_), .Y(_abc_40319_new_n3422_));
OR2X2 OR2X2_48 ( .A(_abc_40319_new_n3592_), .B(_abc_40319_new_n3588_), .Y(_abc_40319_new_n3593_));
OR2X2 OR2X2_49 ( .A(_abc_40319_new_n3634_), .B(_abc_40319_new_n3630_), .Y(_abc_40319_new_n3635_));
OR2X2 OR2X2_5 ( .A(_abc_40319_new_n808_), .B(_abc_40319_new_n803_), .Y(_abc_40319_new_n809_));
OR2X2 OR2X2_50 ( .A(_abc_40319_new_n3729_), .B(_abc_40319_new_n3728_), .Y(n318));
OR2X2 OR2X2_51 ( .A(_abc_40319_new_n665_), .B(_abc_40319_new_n3654_), .Y(_abc_40319_new_n3760_));
OR2X2 OR2X2_52 ( .A(_abc_40319_new_n1194_), .B(_abc_40319_new_n3654_), .Y(_abc_40319_new_n3766_));
OR2X2 OR2X2_53 ( .A(_abc_40319_new_n1219_), .B(_abc_40319_new_n3654_), .Y(_abc_40319_new_n3773_));
OR2X2 OR2X2_54 ( .A(_abc_40319_new_n1320_), .B(_abc_40319_new_n3654_), .Y(_abc_40319_new_n3779_));
OR2X2 OR2X2_55 ( .A(_abc_40319_new_n3785_), .B(_abc_40319_new_n3783_), .Y(n238));
OR2X2 OR2X2_56 ( .A(_abc_40319_new_n1367_), .B(_abc_40319_new_n3654_), .Y(_abc_40319_new_n3787_));
OR2X2 OR2X2_57 ( .A(_abc_40319_new_n1388_), .B(_abc_40319_new_n3654_), .Y(_abc_40319_new_n3790_));
OR2X2 OR2X2_58 ( .A(_abc_40319_new_n765_), .B(_abc_40319_new_n3654_), .Y(_abc_40319_new_n3805_));
OR2X2 OR2X2_59 ( .A(_abc_40319_new_n3895_), .B(_abc_40319_new_n3892_), .Y(_abc_40319_new_n3896_));
OR2X2 OR2X2_6 ( .A(_abc_40319_new_n815_), .B(_abc_40319_new_n811_), .Y(_abc_40319_new_n816_));
OR2X2 OR2X2_60 ( .A(_abc_40319_new_n3635_), .B(_abc_40319_new_n3906_), .Y(_abc_40319_new_n3907_));
OR2X2 OR2X2_61 ( .A(_abc_40319_new_n3612_), .B(_abc_40319_new_n1005_), .Y(_abc_40319_new_n3910_));
OR2X2 OR2X2_62 ( .A(_abc_40319_new_n3916_), .B(_abc_40319_new_n3602_), .Y(_abc_40319_new_n3917_));
OR2X2 OR2X2_63 ( .A(_abc_40319_new_n3583_), .B(_abc_40319_new_n1005_), .Y(_abc_40319_new_n3925_));
OR2X2 OR2X2_7 ( .A(_abc_40319_new_n950_), .B(_abc_40319_new_n953_), .Y(_abc_40319_new_n954_));
OR2X2 OR2X2_8 ( .A(_abc_40319_new_n1052_), .B(_abc_40319_new_n1050_), .Y(_abc_40319_new_n1053_));
OR2X2 OR2X2_9 ( .A(_abc_40319_new_n1037_), .B(_abc_40319_new_n1019_), .Y(_abc_40319_new_n1056_));
XNOR2X1 XNOR2X1_1 ( .A(_abc_40319_new_n562_), .B(IR_REG_26_), .Y(_abc_40319_new_n569_));
XNOR2X1 XNOR2X1_10 ( .A(_abc_40319_new_n1117_), .B(_abc_40319_new_n745_), .Y(_abc_40319_new_n1118_));
XNOR2X1 XNOR2X1_11 ( .A(_abc_40319_new_n1138_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1139_));
XNOR2X1 XNOR2X1_12 ( .A(_abc_40319_new_n604_), .B(_abc_40319_new_n594_), .Y(_abc_40319_new_n1144_));
XNOR2X1 XNOR2X1_13 ( .A(_abc_40319_new_n1160_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1161_));
XNOR2X1 XNOR2X1_14 ( .A(_abc_40319_new_n1192_), .B(_abc_40319_new_n745_), .Y(_abc_40319_new_n1193_));
XNOR2X1 XNOR2X1_15 ( .A(_abc_40319_new_n1212_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1213_));
XNOR2X1 XNOR2X1_16 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n745_), .Y(_abc_40319_new_n1236_));
XNOR2X1 XNOR2X1_17 ( .A(_abc_40319_new_n1262_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1263_));
XNOR2X1 XNOR2X1_18 ( .A(_abc_40319_new_n1278_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1279_));
XNOR2X1 XNOR2X1_19 ( .A(_abc_40319_new_n1338_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1339_));
XNOR2X1 XNOR2X1_2 ( .A(_abc_40319_new_n611_), .B(IR_REG_20_), .Y(_abc_40319_new_n661_));
XNOR2X1 XNOR2X1_20 ( .A(_abc_40319_new_n1026_), .B(REG3_REG_12_), .Y(_abc_40319_new_n1357_));
XNOR2X1 XNOR2X1_21 ( .A(_abc_40319_new_n1362_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1363_));
XNOR2X1 XNOR2X1_22 ( .A(_abc_40319_new_n1343_), .B(_abc_40319_new_n1366_), .Y(_abc_40319_new_n1367_));
XNOR2X1 XNOR2X1_23 ( .A(_abc_40319_new_n1383_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1384_));
XNOR2X1 XNOR2X1_24 ( .A(_abc_40319_new_n1299_), .B(REG3_REG_10_), .Y(_abc_40319_new_n1398_));
XNOR2X1 XNOR2X1_25 ( .A(_abc_40319_new_n1032_), .B(REG3_REG_19_), .Y(_abc_40319_new_n1432_));
XNOR2X1 XNOR2X1_26 ( .A(_abc_40319_new_n1440_), .B(_abc_40319_new_n745_), .Y(_abc_40319_new_n1441_));
XNOR2X1 XNOR2X1_27 ( .A(_abc_40319_new_n1455_), .B(_abc_40319_new_n745_), .Y(_abc_40319_new_n1456_));
XNOR2X1 XNOR2X1_28 ( .A(_abc_40319_new_n1472_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1473_));
XNOR2X1 XNOR2X1_29 ( .A(_abc_40319_new_n868_), .B(_abc_40319_new_n834_), .Y(_abc_40319_new_n1547_));
XNOR2X1 XNOR2X1_3 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n548_), .Y(_abc_40319_new_n794_));
XNOR2X1 XNOR2X1_30 ( .A(_abc_40319_new_n1554_), .B(_abc_40319_new_n1547_), .Y(_abc_40319_new_n1555_));
XNOR2X1 XNOR2X1_31 ( .A(_abc_40319_new_n1441_), .B(_abc_40319_new_n1438_), .Y(_abc_40319_new_n1564_));
XNOR2X1 XNOR2X1_32 ( .A(_abc_40319_new_n1563_), .B(_abc_40319_new_n1564_), .Y(_abc_40319_new_n1565_));
XNOR2X1 XNOR2X1_33 ( .A(_abc_40319_new_n1584_), .B(_abc_40319_new_n745_), .Y(_abc_40319_new_n1585_));
XNOR2X1 XNOR2X1_34 ( .A(_abc_40319_new_n2548_), .B(_abc_40319_new_n892_), .Y(_abc_40319_new_n2549_));
XNOR2X1 XNOR2X1_35 ( .A(_abc_40319_new_n892_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2553_));
XNOR2X1 XNOR2X1_36 ( .A(_abc_40319_new_n836_), .B(REG2_REG_2_), .Y(_abc_40319_new_n2563_));
XNOR2X1 XNOR2X1_37 ( .A(_abc_40319_new_n2570_), .B(_abc_40319_new_n2572_), .Y(_abc_40319_new_n2573_));
XNOR2X1 XNOR2X1_38 ( .A(_abc_40319_new_n821_), .B(REG2_REG_3_), .Y(_abc_40319_new_n2579_));
XNOR2X1 XNOR2X1_39 ( .A(_abc_40319_new_n796_), .B(REG1_REG_4_), .Y(_abc_40319_new_n2600_));
XNOR2X1 XNOR2X1_4 ( .A(_abc_40319_new_n835_), .B(IR_REG_2_), .Y(_abc_40319_new_n836_));
XNOR2X1 XNOR2X1_40 ( .A(_abc_40319_new_n2599_), .B(_abc_40319_new_n2600_), .Y(_abc_40319_new_n2601_));
XNOR2X1 XNOR2X1_41 ( .A(_abc_40319_new_n767_), .B(REG2_REG_5_), .Y(_abc_40319_new_n2609_));
XNOR2X1 XNOR2X1_42 ( .A(_abc_40319_new_n2608_), .B(_abc_40319_new_n2609_), .Y(_abc_40319_new_n2610_));
XNOR2X1 XNOR2X1_43 ( .A(_abc_40319_new_n942_), .B(REG1_REG_6_), .Y(_abc_40319_new_n2625_));
XNOR2X1 XNOR2X1_44 ( .A(_abc_40319_new_n942_), .B(_abc_40319_new_n951_), .Y(_abc_40319_new_n2632_));
XNOR2X1 XNOR2X1_45 ( .A(_abc_40319_new_n2678_), .B(_abc_40319_new_n1273_), .Y(_abc_40319_new_n2679_));
XNOR2X1 XNOR2X1_46 ( .A(_abc_40319_new_n2719_), .B(_abc_40319_new_n1390_), .Y(_abc_40319_new_n2720_));
XNOR2X1 XNOR2X1_47 ( .A(_abc_40319_new_n2745_), .B(_abc_40319_new_n2743_), .Y(_abc_40319_new_n2746_));
XNOR2X1 XNOR2X1_48 ( .A(_abc_40319_new_n2753_), .B(_abc_40319_new_n2752_), .Y(_abc_40319_new_n2754_));
XNOR2X1 XNOR2X1_49 ( .A(_abc_40319_new_n2768_), .B(_abc_40319_new_n2765_), .Y(_abc_40319_new_n2769_));
XNOR2X1 XNOR2X1_5 ( .A(_abc_40319_new_n1048_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1049_));
XNOR2X1 XNOR2X1_50 ( .A(_abc_40319_new_n2775_), .B(_abc_40319_new_n2772_), .Y(_abc_40319_new_n2776_));
XNOR2X1 XNOR2X1_51 ( .A(_abc_40319_new_n2787_), .B(_abc_40319_new_n1323_), .Y(_abc_40319_new_n2788_));
XNOR2X1 XNOR2X1_52 ( .A(_abc_40319_new_n2818_), .B(_abc_40319_new_n2814_), .Y(_abc_40319_new_n2819_));
XNOR2X1 XNOR2X1_53 ( .A(_abc_40319_new_n2832_), .B(_abc_40319_new_n1221_), .Y(_abc_40319_new_n2833_));
XNOR2X1 XNOR2X1_54 ( .A(_abc_40319_new_n2843_), .B(_abc_40319_new_n2839_), .Y(_abc_40319_new_n2844_));
XNOR2X1 XNOR2X1_55 ( .A(_abc_40319_new_n2860_), .B(_abc_40319_new_n2858_), .Y(_abc_40319_new_n2861_));
XNOR2X1 XNOR2X1_56 ( .A(_abc_40319_new_n2883_), .B(_abc_40319_new_n2881_), .Y(_abc_40319_new_n2884_));
XNOR2X1 XNOR2X1_57 ( .A(_abc_40319_new_n2889_), .B(_abc_40319_new_n2887_), .Y(_abc_40319_new_n2890_));
XNOR2X1 XNOR2X1_58 ( .A(_abc_40319_new_n667_), .B(_abc_40319_new_n2939_), .Y(_abc_40319_new_n2940_));
XNOR2X1 XNOR2X1_59 ( .A(_abc_40319_new_n2982_), .B(_abc_40319_new_n2097_), .Y(_abc_40319_new_n2997_));
XNOR2X1 XNOR2X1_6 ( .A(_abc_40319_new_n1067_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1068_));
XNOR2X1 XNOR2X1_60 ( .A(_abc_40319_new_n3003_), .B(_abc_40319_new_n2121_), .Y(_abc_40319_new_n3004_));
XNOR2X1 XNOR2X1_61 ( .A(_abc_40319_new_n2978_), .B(_abc_40319_new_n1581_), .Y(_abc_40319_new_n3111_));
XNOR2X1 XNOR2X1_62 ( .A(_abc_40319_new_n3135_), .B(_abc_40319_new_n1017_), .Y(_abc_40319_new_n3136_));
XNOR2X1 XNOR2X1_63 ( .A(_abc_40319_new_n3126_), .B(_abc_40319_new_n2125_), .Y(_abc_40319_new_n3156_));
XNOR2X1 XNOR2X1_64 ( .A(_abc_40319_new_n3120_), .B(_abc_40319_new_n3203_), .Y(_abc_40319_new_n3204_));
XNOR2X1 XNOR2X1_65 ( .A(_abc_40319_new_n3206_), .B(_abc_40319_new_n3203_), .Y(_abc_40319_new_n3207_));
XNOR2X1 XNOR2X1_66 ( .A(_abc_40319_new_n3228_), .B(_abc_40319_new_n2139_), .Y(_abc_40319_new_n3229_));
XNOR2X1 XNOR2X1_67 ( .A(_abc_40319_new_n3254_), .B(_abc_40319_new_n2216_), .Y(_abc_40319_new_n3255_));
XNOR2X1 XNOR2X1_68 ( .A(_abc_40319_new_n3268_), .B(_abc_40319_new_n3265_), .Y(_abc_40319_new_n3269_));
XNOR2X1 XNOR2X1_69 ( .A(_abc_40319_new_n3286_), .B(_abc_40319_new_n2220_), .Y(_abc_40319_new_n3287_));
XNOR2X1 XNOR2X1_7 ( .A(_abc_40319_new_n1081_), .B(_abc_40319_new_n745_), .Y(_abc_40319_new_n1082_));
XNOR2X1 XNOR2X1_70 ( .A(_abc_40319_new_n3266_), .B(_abc_40319_new_n2170_), .Y(_abc_40319_new_n3308_));
XNOR2X1 XNOR2X1_71 ( .A(_abc_40319_new_n3298_), .B(_abc_40319_new_n1570_), .Y(_abc_40319_new_n3315_));
XNOR2X1 XNOR2X1_72 ( .A(_abc_40319_new_n3253_), .B(_abc_40319_new_n2164_), .Y(_abc_40319_new_n3324_));
XNOR2X1 XNOR2X1_73 ( .A(_abc_40319_new_n3343_), .B(_abc_40319_new_n2158_), .Y(_abc_40319_new_n3344_));
XNOR2X1 XNOR2X1_74 ( .A(_abc_40319_new_n3071_), .B(_abc_40319_new_n2199_), .Y(_abc_40319_new_n3382_));
XNOR2X1 XNOR2X1_75 ( .A(_abc_40319_new_n3384_), .B(_abc_40319_new_n2199_), .Y(_abc_40319_new_n3385_));
XNOR2X1 XNOR2X1_76 ( .A(_abc_40319_new_n3377_), .B(_abc_40319_new_n1865_), .Y(_abc_40319_new_n3395_));
XNOR2X1 XNOR2X1_77 ( .A(_abc_40319_new_n3070_), .B(_abc_40319_new_n2224_), .Y(_abc_40319_new_n3398_));
XNOR2X1 XNOR2X1_78 ( .A(_abc_40319_new_n3360_), .B(_abc_40319_new_n2241_), .Y(_abc_40319_new_n3408_));
XNOR2X1 XNOR2X1_79 ( .A(_abc_40319_new_n3069_), .B(_abc_40319_new_n2241_), .Y(_abc_40319_new_n3409_));
XNOR2X1 XNOR2X1_8 ( .A(_abc_40319_new_n1097_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1098_));
XNOR2X1 XNOR2X1_80 ( .A(_abc_40319_new_n3359_), .B(_abc_40319_new_n2231_), .Y(_abc_40319_new_n3427_));
XNOR2X1 XNOR2X1_81 ( .A(_abc_40319_new_n3430_), .B(_abc_40319_new_n2231_), .Y(_abc_40319_new_n3431_));
XNOR2X1 XNOR2X1_82 ( .A(_abc_40319_new_n2970_), .B(_abc_40319_new_n1654_), .Y(_abc_40319_new_n3446_));
XNOR2X1 XNOR2X1_83 ( .A(_abc_40319_new_n3428_), .B(_abc_40319_new_n2204_), .Y(_abc_40319_new_n3448_));
XNOR2X1 XNOR2X1_84 ( .A(_abc_40319_new_n3468_), .B(_abc_40319_new_n2180_), .Y(_abc_40319_new_n3469_));
XNOR2X1 XNOR2X1_85 ( .A(_abc_40319_new_n2969_), .B(_abc_40319_new_n1393_), .Y(_abc_40319_new_n3485_));
XNOR2X1 XNOR2X1_86 ( .A(_abc_40319_new_n3355_), .B(_abc_40319_new_n2185_), .Y(_abc_40319_new_n3496_));
XNOR2X1 XNOR2X1_87 ( .A(_abc_40319_new_n3478_), .B(_abc_40319_new_n2185_), .Y(_abc_40319_new_n3497_));
XNOR2X1 XNOR2X1_88 ( .A(_abc_40319_new_n3512_), .B(_abc_40319_new_n2195_), .Y(_abc_40319_new_n3513_));
XNOR2X1 XNOR2X1_89 ( .A(_abc_40319_new_n3477_), .B(_abc_40319_new_n2195_), .Y(_abc_40319_new_n3514_));
XNOR2X1 XNOR2X1_9 ( .A(_abc_40319_new_n1035_), .B(_abc_40319_new_n1021_), .Y(_abc_40319_new_n1110_));
XNOR2X1 XNOR2X1_90 ( .A(_abc_40319_new_n2968_), .B(_abc_40319_new_n2427_), .Y(_abc_40319_new_n3518_));
XNOR2X1 XNOR2X1_91 ( .A(_abc_40319_new_n3053_), .B(_abc_40319_new_n2249_), .Y(_abc_40319_new_n3550_));
XNOR2X1 XNOR2X1_92 ( .A(_abc_40319_new_n2966_), .B(_abc_40319_new_n2246_), .Y(_abc_40319_new_n3554_));
XNOR2X1 XNOR2X1_93 ( .A(_abc_40319_new_n2964_), .B(_abc_40319_new_n1726_), .Y(_abc_40319_new_n3571_));
XNOR2X1 XNOR2X1_94 ( .A(_abc_40319_new_n3599_), .B(_abc_40319_new_n2155_), .Y(_abc_40319_new_n3600_));
XNOR2X1 XNOR2X1_95 ( .A(_abc_40319_new_n3039_), .B(_abc_40319_new_n2245_), .Y(_abc_40319_new_n3612_));
XNOR2X1 XNOR2X1_96 ( .A(_abc_40319_new_n3037_), .B(_abc_40319_new_n2225_), .Y(_abc_40319_new_n3629_));
XOR2X1 XOR2X1_1 ( .A(_abc_40319_new_n814_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n815_));
XOR2X1 XOR2X1_10 ( .A(_abc_40319_new_n1647_), .B(_abc_40319_new_n1793_), .Y(_abc_40319_new_n1794_));
XOR2X1 XOR2X1_11 ( .A(_abc_40319_new_n2564_), .B(_abc_40319_new_n2563_), .Y(_abc_40319_new_n2565_));
XOR2X1 XOR2X1_12 ( .A(_abc_40319_new_n2579_), .B(_abc_40319_new_n2578_), .Y(_abc_40319_new_n2580_));
XOR2X1 XOR2X1_13 ( .A(_abc_40319_new_n2597_), .B(_abc_40319_new_n2595_), .Y(_abc_40319_new_n2598_));
XOR2X1 XOR2X1_14 ( .A(_abc_40319_new_n2698_), .B(_abc_40319_new_n2696_), .Y(_abc_40319_new_n2699_));
XOR2X1 XOR2X1_15 ( .A(_abc_40319_new_n2705_), .B(_abc_40319_new_n2703_), .Y(_abc_40319_new_n2706_));
XOR2X1 XOR2X1_16 ( .A(_abc_40319_new_n2869_), .B(_abc_40319_new_n2866_), .Y(_abc_40319_new_n2870_));
XOR2X1 XOR2X1_17 ( .A(_abc_40319_new_n3231_), .B(_abc_40319_new_n2216_), .Y(_abc_40319_new_n3257_));
XOR2X1 XOR2X1_18 ( .A(_abc_40319_new_n3361_), .B(_abc_40319_new_n2158_), .Y(_abc_40319_new_n3362_));
XOR2X1 XOR2X1_19 ( .A(_abc_40319_new_n3383_), .B(_abc_40319_new_n2224_), .Y(_abc_40319_new_n3400_));
XOR2X1 XOR2X1_2 ( .A(_abc_40319_new_n1310_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1311_));
XOR2X1 XOR2X1_20 ( .A(_abc_40319_new_n3357_), .B(_abc_40319_new_n2204_), .Y(_abc_40319_new_n3452_));
XOR2X1 XOR2X1_21 ( .A(_abc_40319_new_n3067_), .B(_abc_40319_new_n2180_), .Y(_abc_40319_new_n3463_));
XOR2X1 XOR2X1_22 ( .A(_abc_40319_new_n3466_), .B(_abc_40319_new_n2208_), .Y(_abc_40319_new_n3476_));
XOR2X1 XOR2X1_23 ( .A(_abc_40319_new_n3480_), .B(_abc_40319_new_n2208_), .Y(_abc_40319_new_n3481_));
XOR2X1 XOR2X1_24 ( .A(_abc_40319_new_n2477_), .B(_abc_40319_new_n2190_), .Y(_abc_40319_new_n3528_));
XOR2X1 XOR2X1_25 ( .A(_abc_40319_new_n3530_), .B(_abc_40319_new_n2190_), .Y(_abc_40319_new_n3531_));
XOR2X1 XOR2X1_26 ( .A(_abc_40319_new_n3548_), .B(_abc_40319_new_n2249_), .Y(_abc_40319_new_n3549_));
XOR2X1 XOR2X1_27 ( .A(_abc_40319_new_n2471_), .B(_abc_40319_new_n2176_), .Y(_abc_40319_new_n3563_));
XOR2X1 XOR2X1_28 ( .A(_abc_40319_new_n3566_), .B(_abc_40319_new_n2176_), .Y(_abc_40319_new_n3567_));
XOR2X1 XOR2X1_29 ( .A(_abc_40319_new_n3547_), .B(_abc_40319_new_n2235_), .Y(_abc_40319_new_n3580_));
XOR2X1 XOR2X1_3 ( .A(_abc_40319_new_n1405_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1406_));
XOR2X1 XOR2X1_30 ( .A(_abc_40319_new_n3582_), .B(_abc_40319_new_n2235_), .Y(_abc_40319_new_n3583_));
XOR2X1 XOR2X1_4 ( .A(_abc_40319_new_n1419_), .B(_abc_40319_new_n1512_), .Y(_abc_40319_new_n1513_));
XOR2X1 XOR2X1_5 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n1537_), .Y(_abc_40319_new_n1538_));
XOR2X1 XOR2X1_6 ( .A(_abc_40319_new_n1585_), .B(_abc_40319_new_n1583_), .Y(_abc_40319_new_n1586_));
XOR2X1 XOR2X1_7 ( .A(_abc_40319_new_n1621_), .B(_abc_40319_new_n1549_), .Y(_abc_40319_new_n1622_));
XOR2X1 XOR2X1_8 ( .A(_abc_40319_new_n1747_), .B(_abc_40319_new_n1746_), .Y(_abc_40319_new_n1748_));
XOR2X1 XOR2X1_9 ( .A(_abc_40319_new_n1634_), .B(_abc_40319_new_n1757_), .Y(_abc_40319_new_n1758_));


endmodule