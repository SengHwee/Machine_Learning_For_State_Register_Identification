module fpSqrt(rst, clk, ce, ld, \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] , \o[8] , \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] , \o[16] , \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] , \o[24] , \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] , \o[32] , \o[33] , \o[34] , \o[35] , \o[36] , \o[37] , \o[38] , \o[39] , \o[40] , \o[41] , \o[42] , \o[43] , \o[44] , \o[45] , \o[46] , \o[47] , \o[48] , \o[49] , \o[50] , \o[51] , \o[52] , \o[53] , \o[54] , \o[55] , \o[56] , \o[57] , \o[58] , \o[59] , \o[60] , \o[61] , \o[62] , \o[63] , \o[64] , \o[65] , \o[66] , \o[67] , \o[68] , \o[69] , \o[70] , \o[71] , \o[72] , \o[73] , \o[74] , \o[75] , \o[76] , \o[77] , \o[78] , \o[79] , \o[80] , \o[81] , \o[82] , \o[83] , \o[84] , \o[85] , \o[86] , \o[87] , \o[88] , \o[89] , \o[90] , \o[91] , \o[92] , \o[93] , \o[94] , \o[95] , \o[96] , \o[97] , \o[98] , \o[99] , \o[100] , \o[101] , \o[102] , \o[103] , \o[104] , \o[105] , \o[106] , \o[107] , \o[108] , \o[109] , \o[110] , \o[111] , \o[112] , \o[113] , \o[114] , \o[115] , \o[116] , \o[117] , \o[118] , \o[119] , \o[120] , \o[121] , \o[122] , \o[123] , \o[124] , \o[125] , \o[126] , \o[127] , \o[128] , \o[129] , \o[130] , \o[131] , \o[132] , \o[133] , \o[134] , \o[135] , \o[136] , \o[137] , \o[138] , \o[139] , \o[140] , \o[141] , \o[142] , \o[143] , \o[144] , \o[145] , \o[146] , \o[147] , \o[148] , \o[149] , \o[150] , \o[151] , \o[152] , \o[153] , \o[154] , \o[155] , \o[156] , \o[157] , \o[158] , \o[159] , \o[160] , \o[161] , \o[162] , \o[163] , \o[164] , \o[165] , \o[166] , \o[167] , \o[168] , \o[169] , \o[170] , \o[171] , \o[172] , \o[173] , \o[174] , \o[175] , \o[176] , \o[177] , \o[178] , \o[179] , \o[180] , \o[181] , \o[182] , \o[183] , \o[184] , \o[185] , \o[186] , \o[187] , \o[188] , \o[189] , \o[190] , \o[191] , \o[192] , \o[193] , \o[194] , \o[195] , \o[196] , \o[197] , \o[198] , \o[199] , \o[200] , \o[201] , \o[202] , \o[203] , \o[204] , \o[205] , \o[206] , \o[207] , \o[208] , \o[209] , \o[210] , \o[211] , \o[212] , \o[213] , \o[214] , \o[215] , \o[216] , \o[217] , \o[218] , \o[219] , \o[220] , \o[221] , \o[222] , \o[223] , \o[224] , \o[225] , \o[226] , \o[227] , \o[228] , \o[229] , \o[230] , \o[231] , \o[232] , \o[233] , \o[234] , \o[235] , \o[236] , \o[237] , \o[238] , \o[239] , \o[240] , \o[241] , done);

wire _abc_73687_new_n1001_; 
wire _abc_73687_new_n1002_; 
wire _abc_73687_new_n1004_; 
wire _abc_73687_new_n1005_; 
wire _abc_73687_new_n1007_; 
wire _abc_73687_new_n1008_; 
wire _abc_73687_new_n1010_; 
wire _abc_73687_new_n1011_; 
wire _abc_73687_new_n1013_; 
wire _abc_73687_new_n1014_; 
wire _abc_73687_new_n1016_; 
wire _abc_73687_new_n1017_; 
wire _abc_73687_new_n1019_; 
wire _abc_73687_new_n1020_; 
wire _abc_73687_new_n1022_; 
wire _abc_73687_new_n1023_; 
wire _abc_73687_new_n1025_; 
wire _abc_73687_new_n1026_; 
wire _abc_73687_new_n1028_; 
wire _abc_73687_new_n1029_; 
wire _abc_73687_new_n1031_; 
wire _abc_73687_new_n1032_; 
wire _abc_73687_new_n1034_; 
wire _abc_73687_new_n1035_; 
wire _abc_73687_new_n1037_; 
wire _abc_73687_new_n1038_; 
wire _abc_73687_new_n1040_; 
wire _abc_73687_new_n1041_; 
wire _abc_73687_new_n1043_; 
wire _abc_73687_new_n1044_; 
wire _abc_73687_new_n1046_; 
wire _abc_73687_new_n1047_; 
wire _abc_73687_new_n1049_; 
wire _abc_73687_new_n1050_; 
wire _abc_73687_new_n1052_; 
wire _abc_73687_new_n1053_; 
wire _abc_73687_new_n1055_; 
wire _abc_73687_new_n1056_; 
wire _abc_73687_new_n1058_; 
wire _abc_73687_new_n1059_; 
wire _abc_73687_new_n1061_; 
wire _abc_73687_new_n1062_; 
wire _abc_73687_new_n1064_; 
wire _abc_73687_new_n1065_; 
wire _abc_73687_new_n1067_; 
wire _abc_73687_new_n1068_; 
wire _abc_73687_new_n1070_; 
wire _abc_73687_new_n1071_; 
wire _abc_73687_new_n1073_; 
wire _abc_73687_new_n1074_; 
wire _abc_73687_new_n1076_; 
wire _abc_73687_new_n1077_; 
wire _abc_73687_new_n1079_; 
wire _abc_73687_new_n1080_; 
wire _abc_73687_new_n1082_; 
wire _abc_73687_new_n1083_; 
wire _abc_73687_new_n1085_; 
wire _abc_73687_new_n1086_; 
wire _abc_73687_new_n1088_; 
wire _abc_73687_new_n1089_; 
wire _abc_73687_new_n1091_; 
wire _abc_73687_new_n1092_; 
wire _abc_73687_new_n1094_; 
wire _abc_73687_new_n1095_; 
wire _abc_73687_new_n1097_; 
wire _abc_73687_new_n1098_; 
wire _abc_73687_new_n1100_; 
wire _abc_73687_new_n1101_; 
wire _abc_73687_new_n1103_; 
wire _abc_73687_new_n1104_; 
wire _abc_73687_new_n1106_; 
wire _abc_73687_new_n1107_; 
wire _abc_73687_new_n1109_; 
wire _abc_73687_new_n1110_; 
wire _abc_73687_new_n1112_; 
wire _abc_73687_new_n1113_; 
wire _abc_73687_new_n1115_; 
wire _abc_73687_new_n1116_; 
wire _abc_73687_new_n1118_; 
wire _abc_73687_new_n1119_; 
wire _abc_73687_new_n1121_; 
wire _abc_73687_new_n1122_; 
wire _abc_73687_new_n1124_; 
wire _abc_73687_new_n1125_; 
wire _abc_73687_new_n1127_; 
wire _abc_73687_new_n1128_; 
wire _abc_73687_new_n1130_; 
wire _abc_73687_new_n1131_; 
wire _abc_73687_new_n1133_; 
wire _abc_73687_new_n1134_; 
wire _abc_73687_new_n1136_; 
wire _abc_73687_new_n1137_; 
wire _abc_73687_new_n1139_; 
wire _abc_73687_new_n1140_; 
wire _abc_73687_new_n1142_; 
wire _abc_73687_new_n1143_; 
wire _abc_73687_new_n1145_; 
wire _abc_73687_new_n1146_; 
wire _abc_73687_new_n1148_; 
wire _abc_73687_new_n1149_; 
wire _abc_73687_new_n1151_; 
wire _abc_73687_new_n1152_; 
wire _abc_73687_new_n1154_; 
wire _abc_73687_new_n1155_; 
wire _abc_73687_new_n1157_; 
wire _abc_73687_new_n1158_; 
wire _abc_73687_new_n1160_; 
wire _abc_73687_new_n1161_; 
wire _abc_73687_new_n1163_; 
wire _abc_73687_new_n1164_; 
wire _abc_73687_new_n1169_; 
wire _abc_73687_new_n1170_; 
wire _abc_73687_new_n1171_; 
wire _abc_73687_new_n1173_; 
wire _abc_73687_new_n1174_; 
wire _abc_73687_new_n1176_; 
wire _abc_73687_new_n1177_; 
wire _abc_73687_new_n1179_; 
wire _abc_73687_new_n1180_; 
wire _abc_73687_new_n1182_; 
wire _abc_73687_new_n1183_; 
wire _abc_73687_new_n1185_; 
wire _abc_73687_new_n1186_; 
wire _abc_73687_new_n1188_; 
wire _abc_73687_new_n1189_; 
wire _abc_73687_new_n1191_; 
wire _abc_73687_new_n1192_; 
wire _abc_73687_new_n1194_; 
wire _abc_73687_new_n1195_; 
wire _abc_73687_new_n1197_; 
wire _abc_73687_new_n1198_; 
wire _abc_73687_new_n1200_; 
wire _abc_73687_new_n1201_; 
wire _abc_73687_new_n1203_; 
wire _abc_73687_new_n1204_; 
wire _abc_73687_new_n1206_; 
wire _abc_73687_new_n1207_; 
wire _abc_73687_new_n1209_; 
wire _abc_73687_new_n1210_; 
wire _abc_73687_new_n1212_; 
wire _abc_73687_new_n1213_; 
wire _abc_73687_new_n1215_; 
wire _abc_73687_new_n1216_; 
wire _abc_73687_new_n1218_; 
wire _abc_73687_new_n1219_; 
wire _abc_73687_new_n1221_; 
wire _abc_73687_new_n1222_; 
wire _abc_73687_new_n1224_; 
wire _abc_73687_new_n1225_; 
wire _abc_73687_new_n1227_; 
wire _abc_73687_new_n1228_; 
wire _abc_73687_new_n1230_; 
wire _abc_73687_new_n1231_; 
wire _abc_73687_new_n1233_; 
wire _abc_73687_new_n1234_; 
wire _abc_73687_new_n1236_; 
wire _abc_73687_new_n1237_; 
wire _abc_73687_new_n1239_; 
wire _abc_73687_new_n1240_; 
wire _abc_73687_new_n1242_; 
wire _abc_73687_new_n1243_; 
wire _abc_73687_new_n1245_; 
wire _abc_73687_new_n1246_; 
wire _abc_73687_new_n1248_; 
wire _abc_73687_new_n1249_; 
wire _abc_73687_new_n1251_; 
wire _abc_73687_new_n1252_; 
wire _abc_73687_new_n1254_; 
wire _abc_73687_new_n1255_; 
wire _abc_73687_new_n1257_; 
wire _abc_73687_new_n1258_; 
wire _abc_73687_new_n1260_; 
wire _abc_73687_new_n1261_; 
wire _abc_73687_new_n1263_; 
wire _abc_73687_new_n1264_; 
wire _abc_73687_new_n1266_; 
wire _abc_73687_new_n1267_; 
wire _abc_73687_new_n1269_; 
wire _abc_73687_new_n1270_; 
wire _abc_73687_new_n1272_; 
wire _abc_73687_new_n1273_; 
wire _abc_73687_new_n1275_; 
wire _abc_73687_new_n1276_; 
wire _abc_73687_new_n1278_; 
wire _abc_73687_new_n1279_; 
wire _abc_73687_new_n1281_; 
wire _abc_73687_new_n1282_; 
wire _abc_73687_new_n1284_; 
wire _abc_73687_new_n1285_; 
wire _abc_73687_new_n1287_; 
wire _abc_73687_new_n1288_; 
wire _abc_73687_new_n1290_; 
wire _abc_73687_new_n1291_; 
wire _abc_73687_new_n1293_; 
wire _abc_73687_new_n1294_; 
wire _abc_73687_new_n1296_; 
wire _abc_73687_new_n1297_; 
wire _abc_73687_new_n1299_; 
wire _abc_73687_new_n1300_; 
wire _abc_73687_new_n1302_; 
wire _abc_73687_new_n1303_; 
wire _abc_73687_new_n1305_; 
wire _abc_73687_new_n1306_; 
wire _abc_73687_new_n1308_; 
wire _abc_73687_new_n1309_; 
wire _abc_73687_new_n1311_; 
wire _abc_73687_new_n1312_; 
wire _abc_73687_new_n1314_; 
wire _abc_73687_new_n1315_; 
wire _abc_73687_new_n1317_; 
wire _abc_73687_new_n1318_; 
wire _abc_73687_new_n1320_; 
wire _abc_73687_new_n1321_; 
wire _abc_73687_new_n1323_; 
wire _abc_73687_new_n1324_; 
wire _abc_73687_new_n1326_; 
wire _abc_73687_new_n1327_; 
wire _abc_73687_new_n1329_; 
wire _abc_73687_new_n1330_; 
wire _abc_73687_new_n1332_; 
wire _abc_73687_new_n1333_; 
wire _abc_73687_new_n1335_; 
wire _abc_73687_new_n1336_; 
wire _abc_73687_new_n1338_; 
wire _abc_73687_new_n1339_; 
wire _abc_73687_new_n1341_; 
wire _abc_73687_new_n1342_; 
wire _abc_73687_new_n1344_; 
wire _abc_73687_new_n1345_; 
wire _abc_73687_new_n1347_; 
wire _abc_73687_new_n1348_; 
wire _abc_73687_new_n1350_; 
wire _abc_73687_new_n1351_; 
wire _abc_73687_new_n1353_; 
wire _abc_73687_new_n1354_; 
wire _abc_73687_new_n1356_; 
wire _abc_73687_new_n1357_; 
wire _abc_73687_new_n1359_; 
wire _abc_73687_new_n1360_; 
wire _abc_73687_new_n1362_; 
wire _abc_73687_new_n1363_; 
wire _abc_73687_new_n1365_; 
wire _abc_73687_new_n1366_; 
wire _abc_73687_new_n1368_; 
wire _abc_73687_new_n1369_; 
wire _abc_73687_new_n1371_; 
wire _abc_73687_new_n1372_; 
wire _abc_73687_new_n1374_; 
wire _abc_73687_new_n1375_; 
wire _abc_73687_new_n1377_; 
wire _abc_73687_new_n1378_; 
wire _abc_73687_new_n1380_; 
wire _abc_73687_new_n1381_; 
wire _abc_73687_new_n1383_; 
wire _abc_73687_new_n1384_; 
wire _abc_73687_new_n1386_; 
wire _abc_73687_new_n1387_; 
wire _abc_73687_new_n1389_; 
wire _abc_73687_new_n1390_; 
wire _abc_73687_new_n1392_; 
wire _abc_73687_new_n1393_; 
wire _abc_73687_new_n1395_; 
wire _abc_73687_new_n1396_; 
wire _abc_73687_new_n1398_; 
wire _abc_73687_new_n1399_; 
wire _abc_73687_new_n1401_; 
wire _abc_73687_new_n1402_; 
wire _abc_73687_new_n1404_; 
wire _abc_73687_new_n1405_; 
wire _abc_73687_new_n1407_; 
wire _abc_73687_new_n1408_; 
wire _abc_73687_new_n1410_; 
wire _abc_73687_new_n1411_; 
wire _abc_73687_new_n1413_; 
wire _abc_73687_new_n1414_; 
wire _abc_73687_new_n1416_; 
wire _abc_73687_new_n1417_; 
wire _abc_73687_new_n1419_; 
wire _abc_73687_new_n1420_; 
wire _abc_73687_new_n1422_; 
wire _abc_73687_new_n1423_; 
wire _abc_73687_new_n1425_; 
wire _abc_73687_new_n1426_; 
wire _abc_73687_new_n1428_; 
wire _abc_73687_new_n1429_; 
wire _abc_73687_new_n1431_; 
wire _abc_73687_new_n1432_; 
wire _abc_73687_new_n1434_; 
wire _abc_73687_new_n1435_; 
wire _abc_73687_new_n1437_; 
wire _abc_73687_new_n1438_; 
wire _abc_73687_new_n1440_; 
wire _abc_73687_new_n1441_; 
wire _abc_73687_new_n1443_; 
wire _abc_73687_new_n1444_; 
wire _abc_73687_new_n1446_; 
wire _abc_73687_new_n1447_; 
wire _abc_73687_new_n1449_; 
wire _abc_73687_new_n1450_; 
wire _abc_73687_new_n1452_; 
wire _abc_73687_new_n1453_; 
wire _abc_73687_new_n1455_; 
wire _abc_73687_new_n1456_; 
wire _abc_73687_new_n1458_; 
wire _abc_73687_new_n1459_; 
wire _abc_73687_new_n1461_; 
wire _abc_73687_new_n1462_; 
wire _abc_73687_new_n1464_; 
wire _abc_73687_new_n1465_; 
wire _abc_73687_new_n1467_; 
wire _abc_73687_new_n1468_; 
wire _abc_73687_new_n1470_; 
wire _abc_73687_new_n1471_; 
wire _abc_73687_new_n1473_; 
wire _abc_73687_new_n1474_; 
wire _abc_73687_new_n1476_; 
wire _abc_73687_new_n1477_; 
wire _abc_73687_new_n1479_; 
wire _abc_73687_new_n1480_; 
wire _abc_73687_new_n1482_; 
wire _abc_73687_new_n1483_; 
wire _abc_73687_new_n1485_; 
wire _abc_73687_new_n1486_; 
wire _abc_73687_new_n1488_; 
wire _abc_73687_new_n1489_; 
wire _abc_73687_new_n1491_; 
wire _abc_73687_new_n1492_; 
wire _abc_73687_new_n1494_; 
wire _abc_73687_new_n1495_; 
wire _abc_73687_new_n1497_; 
wire _abc_73687_new_n1498_; 
wire _abc_73687_new_n1500_; 
wire _abc_73687_new_n1501_; 
wire _abc_73687_new_n1503_; 
wire _abc_73687_new_n1504_; 
wire _abc_73687_new_n1507_; 
wire _abc_73687_new_n1508_; 
wire _abc_73687_new_n1509_; 
wire _abc_73687_new_n1510_; 
wire _abc_73687_new_n1511_; 
wire _abc_73687_new_n1512_; 
wire _abc_73687_new_n1514_; 
wire _abc_73687_new_n1515_; 
wire _abc_73687_new_n1516_; 
wire _abc_73687_new_n1517_; 
wire _abc_73687_new_n1518_; 
wire _abc_73687_new_n1519_; 
wire _abc_73687_new_n1521_; 
wire _abc_73687_new_n1522_; 
wire _abc_73687_new_n1523_; 
wire _abc_73687_new_n1524_; 
wire _abc_73687_new_n1525_; 
wire _abc_73687_new_n1526_; 
wire _abc_73687_new_n1527_; 
wire _abc_73687_new_n1528_; 
wire _abc_73687_new_n1529_; 
wire _abc_73687_new_n1531_; 
wire _abc_73687_new_n1532_; 
wire _abc_73687_new_n1533_; 
wire _abc_73687_new_n1534_; 
wire _abc_73687_new_n1535_; 
wire _abc_73687_new_n1536_; 
wire _abc_73687_new_n1537_; 
wire _abc_73687_new_n1538_; 
wire _abc_73687_new_n1539_; 
wire _abc_73687_new_n1540_; 
wire _abc_73687_new_n1541_; 
wire _abc_73687_new_n1542_; 
wire _abc_73687_new_n1543_; 
wire _abc_73687_new_n1544_; 
wire _abc_73687_new_n1545_; 
wire _abc_73687_new_n1546_; 
wire _abc_73687_new_n1548_; 
wire _abc_73687_new_n1549_; 
wire _abc_73687_new_n1550_; 
wire _abc_73687_new_n1551_; 
wire _abc_73687_new_n1552_; 
wire _abc_73687_new_n1553_; 
wire _abc_73687_new_n1554_; 
wire _abc_73687_new_n1555_; 
wire _abc_73687_new_n1556_; 
wire _abc_73687_new_n1557_; 
wire _abc_73687_new_n1558_; 
wire _abc_73687_new_n1559_; 
wire _abc_73687_new_n1561_; 
wire _abc_73687_new_n1562_; 
wire _abc_73687_new_n1563_; 
wire _abc_73687_new_n1564_; 
wire _abc_73687_new_n1565_; 
wire _abc_73687_new_n1566_; 
wire _abc_73687_new_n1567_; 
wire _abc_73687_new_n1568_; 
wire _abc_73687_new_n1569_; 
wire _abc_73687_new_n1570_; 
wire _abc_73687_new_n1571_; 
wire _abc_73687_new_n1572_; 
wire _abc_73687_new_n1574_; 
wire _abc_73687_new_n1575_; 
wire _abc_73687_new_n1576_; 
wire _abc_73687_new_n1577_; 
wire _abc_73687_new_n1578_; 
wire _abc_73687_new_n1579_; 
wire _abc_73687_new_n1580_; 
wire _abc_73687_new_n1581_; 
wire _abc_73687_new_n1582_; 
wire _abc_73687_new_n1583_; 
wire _abc_73687_new_n1584_; 
wire _abc_73687_new_n1585_; 
wire _abc_73687_new_n1587_; 
wire _abc_73687_new_n1588_; 
wire _abc_73687_new_n1589_; 
wire _abc_73687_new_n1590_; 
wire _abc_73687_new_n1591_; 
wire _abc_73687_new_n1592_; 
wire _abc_73687_new_n1593_; 
wire _abc_73687_new_n1594_; 
wire _abc_73687_new_n1595_; 
wire _abc_73687_new_n1596_; 
wire _abc_73687_new_n1597_; 
wire _abc_73687_new_n1598_; 
wire _abc_73687_new_n1600_; 
wire _abc_73687_new_n1601_; 
wire _abc_73687_new_n1602_; 
wire _abc_73687_new_n1603_; 
wire _abc_73687_new_n1604_; 
wire _abc_73687_new_n1605_; 
wire _abc_73687_new_n1606_; 
wire _abc_73687_new_n1607_; 
wire _abc_73687_new_n1608_; 
wire _abc_73687_new_n1609_; 
wire _abc_73687_new_n1610_; 
wire _abc_73687_new_n1611_; 
wire _abc_73687_new_n1613_; 
wire _abc_73687_new_n1614_; 
wire _abc_73687_new_n1615_; 
wire _abc_73687_new_n1616_; 
wire _abc_73687_new_n1617_; 
wire _abc_73687_new_n1618_; 
wire _abc_73687_new_n1619_; 
wire _abc_73687_new_n1620_; 
wire _abc_73687_new_n1621_; 
wire _abc_73687_new_n1622_; 
wire _abc_73687_new_n1623_; 
wire _abc_73687_new_n1624_; 
wire _abc_73687_new_n1626_; 
wire _abc_73687_new_n1627_; 
wire _abc_73687_new_n1628_; 
wire _abc_73687_new_n1629_; 
wire _abc_73687_new_n1630_; 
wire _abc_73687_new_n1631_; 
wire _abc_73687_new_n1632_; 
wire _abc_73687_new_n1633_; 
wire _abc_73687_new_n1634_; 
wire _abc_73687_new_n1635_; 
wire _abc_73687_new_n1636_; 
wire _abc_73687_new_n1637_; 
wire _abc_73687_new_n1638_; 
wire _abc_73687_new_n1639_; 
wire _abc_73687_new_n1640_; 
wire _abc_73687_new_n1642_; 
wire _abc_73687_new_n1643_; 
wire _abc_73687_new_n1644_; 
wire _abc_73687_new_n1645_; 
wire _abc_73687_new_n1646_; 
wire _abc_73687_new_n1647_; 
wire _abc_73687_new_n1648_; 
wire _abc_73687_new_n1649_; 
wire _abc_73687_new_n1650_; 
wire _abc_73687_new_n1651_; 
wire _abc_73687_new_n1652_; 
wire _abc_73687_new_n1653_; 
wire _abc_73687_new_n1655_; 
wire _abc_73687_new_n1656_; 
wire _abc_73687_new_n1657_; 
wire _abc_73687_new_n1658_; 
wire _abc_73687_new_n1659_; 
wire _abc_73687_new_n1660_; 
wire _abc_73687_new_n1661_; 
wire _abc_73687_new_n1662_; 
wire _abc_73687_new_n1663_; 
wire _abc_73687_new_n1664_; 
wire _abc_73687_new_n1665_; 
wire _abc_73687_new_n1666_; 
wire _abc_73687_new_n1667_; 
wire _abc_73687_new_n1669_; 
wire _abc_73687_new_n1670_; 
wire _abc_73687_new_n1671_; 
wire _abc_73687_new_n1672_; 
wire _abc_73687_new_n1673_; 
wire _abc_73687_new_n1674_; 
wire _abc_73687_new_n1675_; 
wire _abc_73687_new_n1676_; 
wire _abc_73687_new_n1677_; 
wire _abc_73687_new_n1678_; 
wire _abc_73687_new_n1679_; 
wire _abc_73687_new_n1681_; 
wire _abc_73687_new_n1682_; 
wire _abc_73687_new_n1683_; 
wire _abc_73687_new_n1684_; 
wire _abc_73687_new_n1685_; 
wire _abc_73687_new_n1686_; 
wire _abc_73687_new_n1687_; 
wire _abc_73687_new_n753_; 
wire _abc_73687_new_n830_; 
wire _abc_73687_new_n831_; 
wire _abc_73687_new_n833_; 
wire _abc_73687_new_n834_; 
wire _abc_73687_new_n836_; 
wire _abc_73687_new_n837_; 
wire _abc_73687_new_n839_; 
wire _abc_73687_new_n840_; 
wire _abc_73687_new_n842_; 
wire _abc_73687_new_n843_; 
wire _abc_73687_new_n845_; 
wire _abc_73687_new_n846_; 
wire _abc_73687_new_n848_; 
wire _abc_73687_new_n849_; 
wire _abc_73687_new_n851_; 
wire _abc_73687_new_n852_; 
wire _abc_73687_new_n854_; 
wire _abc_73687_new_n855_; 
wire _abc_73687_new_n857_; 
wire _abc_73687_new_n858_; 
wire _abc_73687_new_n860_; 
wire _abc_73687_new_n861_; 
wire _abc_73687_new_n863_; 
wire _abc_73687_new_n864_; 
wire _abc_73687_new_n866_; 
wire _abc_73687_new_n867_; 
wire _abc_73687_new_n869_; 
wire _abc_73687_new_n870_; 
wire _abc_73687_new_n872_; 
wire _abc_73687_new_n873_; 
wire _abc_73687_new_n875_; 
wire _abc_73687_new_n876_; 
wire _abc_73687_new_n878_; 
wire _abc_73687_new_n879_; 
wire _abc_73687_new_n881_; 
wire _abc_73687_new_n882_; 
wire _abc_73687_new_n884_; 
wire _abc_73687_new_n885_; 
wire _abc_73687_new_n887_; 
wire _abc_73687_new_n888_; 
wire _abc_73687_new_n890_; 
wire _abc_73687_new_n891_; 
wire _abc_73687_new_n893_; 
wire _abc_73687_new_n894_; 
wire _abc_73687_new_n896_; 
wire _abc_73687_new_n897_; 
wire _abc_73687_new_n899_; 
wire _abc_73687_new_n900_; 
wire _abc_73687_new_n902_; 
wire _abc_73687_new_n903_; 
wire _abc_73687_new_n905_; 
wire _abc_73687_new_n906_; 
wire _abc_73687_new_n908_; 
wire _abc_73687_new_n909_; 
wire _abc_73687_new_n911_; 
wire _abc_73687_new_n912_; 
wire _abc_73687_new_n914_; 
wire _abc_73687_new_n915_; 
wire _abc_73687_new_n917_; 
wire _abc_73687_new_n918_; 
wire _abc_73687_new_n920_; 
wire _abc_73687_new_n921_; 
wire _abc_73687_new_n923_; 
wire _abc_73687_new_n924_; 
wire _abc_73687_new_n926_; 
wire _abc_73687_new_n927_; 
wire _abc_73687_new_n929_; 
wire _abc_73687_new_n930_; 
wire _abc_73687_new_n932_; 
wire _abc_73687_new_n933_; 
wire _abc_73687_new_n935_; 
wire _abc_73687_new_n936_; 
wire _abc_73687_new_n938_; 
wire _abc_73687_new_n939_; 
wire _abc_73687_new_n941_; 
wire _abc_73687_new_n942_; 
wire _abc_73687_new_n944_; 
wire _abc_73687_new_n945_; 
wire _abc_73687_new_n947_; 
wire _abc_73687_new_n948_; 
wire _abc_73687_new_n950_; 
wire _abc_73687_new_n951_; 
wire _abc_73687_new_n953_; 
wire _abc_73687_new_n954_; 
wire _abc_73687_new_n956_; 
wire _abc_73687_new_n957_; 
wire _abc_73687_new_n959_; 
wire _abc_73687_new_n960_; 
wire _abc_73687_new_n962_; 
wire _abc_73687_new_n963_; 
wire _abc_73687_new_n965_; 
wire _abc_73687_new_n966_; 
wire _abc_73687_new_n968_; 
wire _abc_73687_new_n969_; 
wire _abc_73687_new_n971_; 
wire _abc_73687_new_n972_; 
wire _abc_73687_new_n974_; 
wire _abc_73687_new_n975_; 
wire _abc_73687_new_n977_; 
wire _abc_73687_new_n978_; 
wire _abc_73687_new_n980_; 
wire _abc_73687_new_n981_; 
wire _abc_73687_new_n983_; 
wire _abc_73687_new_n984_; 
wire _abc_73687_new_n986_; 
wire _abc_73687_new_n987_; 
wire _abc_73687_new_n989_; 
wire _abc_73687_new_n990_; 
wire _abc_73687_new_n992_; 
wire _abc_73687_new_n993_; 
wire _abc_73687_new_n995_; 
wire _abc_73687_new_n996_; 
wire _abc_73687_new_n998_; 
wire _abc_73687_new_n999_; 
wire aNan; 
input \a[0] ;
input \a[100] ;
input \a[101] ;
input \a[102] ;
input \a[103] ;
input \a[104] ;
input \a[105] ;
input \a[106] ;
input \a[107] ;
input \a[108] ;
input \a[109] ;
input \a[10] ;
input \a[110] ;
input \a[111] ;
input \a[112] ;
input \a[113] ;
input \a[114] ;
input \a[115] ;
input \a[116] ;
input \a[117] ;
input \a[118] ;
input \a[119] ;
input \a[11] ;
input \a[120] ;
input \a[121] ;
input \a[122] ;
input \a[123] ;
input \a[124] ;
input \a[125] ;
input \a[126] ;
input \a[127] ;
input \a[12] ;
input \a[13] ;
input \a[14] ;
input \a[15] ;
input \a[16] ;
input \a[17] ;
input \a[18] ;
input \a[19] ;
input \a[1] ;
input \a[20] ;
input \a[21] ;
input \a[22] ;
input \a[23] ;
input \a[24] ;
input \a[25] ;
input \a[26] ;
input \a[27] ;
input \a[28] ;
input \a[29] ;
input \a[2] ;
input \a[30] ;
input \a[31] ;
input \a[32] ;
input \a[33] ;
input \a[34] ;
input \a[35] ;
input \a[36] ;
input \a[37] ;
input \a[38] ;
input \a[39] ;
input \a[3] ;
input \a[40] ;
input \a[41] ;
input \a[42] ;
input \a[43] ;
input \a[44] ;
input \a[45] ;
input \a[46] ;
input \a[47] ;
input \a[48] ;
input \a[49] ;
input \a[4] ;
input \a[50] ;
input \a[51] ;
input \a[52] ;
input \a[53] ;
input \a[54] ;
input \a[55] ;
input \a[56] ;
input \a[57] ;
input \a[58] ;
input \a[59] ;
input \a[5] ;
input \a[60] ;
input \a[61] ;
input \a[62] ;
input \a[63] ;
input \a[64] ;
input \a[65] ;
input \a[66] ;
input \a[67] ;
input \a[68] ;
input \a[69] ;
input \a[6] ;
input \a[70] ;
input \a[71] ;
input \a[72] ;
input \a[73] ;
input \a[74] ;
input \a[75] ;
input \a[76] ;
input \a[77] ;
input \a[78] ;
input \a[79] ;
input \a[7] ;
input \a[80] ;
input \a[81] ;
input \a[82] ;
input \a[83] ;
input \a[84] ;
input \a[85] ;
input \a[86] ;
input \a[87] ;
input \a[88] ;
input \a[89] ;
input \a[8] ;
input \a[90] ;
input \a[91] ;
input \a[92] ;
input \a[93] ;
input \a[94] ;
input \a[95] ;
input \a[96] ;
input \a[97] ;
input \a[98] ;
input \a[99] ;
input \a[9] ;
input ce;
input clk;
output done;
wire fracta1_0_; 
wire fracta1_100_; 
wire fracta1_101_; 
wire fracta1_102_; 
wire fracta1_103_; 
wire fracta1_104_; 
wire fracta1_105_; 
wire fracta1_106_; 
wire fracta1_107_; 
wire fracta1_108_; 
wire fracta1_109_; 
wire fracta1_10_; 
wire fracta1_110_; 
wire fracta1_111_; 
wire fracta1_112_; 
wire fracta1_113_; 
wire fracta1_11_; 
wire fracta1_12_; 
wire fracta1_13_; 
wire fracta1_14_; 
wire fracta1_15_; 
wire fracta1_16_; 
wire fracta1_17_; 
wire fracta1_18_; 
wire fracta1_19_; 
wire fracta1_1_; 
wire fracta1_20_; 
wire fracta1_21_; 
wire fracta1_22_; 
wire fracta1_23_; 
wire fracta1_24_; 
wire fracta1_25_; 
wire fracta1_26_; 
wire fracta1_27_; 
wire fracta1_28_; 
wire fracta1_29_; 
wire fracta1_2_; 
wire fracta1_30_; 
wire fracta1_31_; 
wire fracta1_32_; 
wire fracta1_33_; 
wire fracta1_34_; 
wire fracta1_35_; 
wire fracta1_36_; 
wire fracta1_37_; 
wire fracta1_38_; 
wire fracta1_39_; 
wire fracta1_3_; 
wire fracta1_40_; 
wire fracta1_41_; 
wire fracta1_42_; 
wire fracta1_43_; 
wire fracta1_44_; 
wire fracta1_45_; 
wire fracta1_46_; 
wire fracta1_47_; 
wire fracta1_48_; 
wire fracta1_49_; 
wire fracta1_4_; 
wire fracta1_50_; 
wire fracta1_51_; 
wire fracta1_52_; 
wire fracta1_53_; 
wire fracta1_54_; 
wire fracta1_55_; 
wire fracta1_56_; 
wire fracta1_57_; 
wire fracta1_58_; 
wire fracta1_59_; 
wire fracta1_5_; 
wire fracta1_60_; 
wire fracta1_61_; 
wire fracta1_62_; 
wire fracta1_63_; 
wire fracta1_64_; 
wire fracta1_65_; 
wire fracta1_66_; 
wire fracta1_67_; 
wire fracta1_68_; 
wire fracta1_69_; 
wire fracta1_6_; 
wire fracta1_70_; 
wire fracta1_71_; 
wire fracta1_72_; 
wire fracta1_73_; 
wire fracta1_74_; 
wire fracta1_75_; 
wire fracta1_76_; 
wire fracta1_77_; 
wire fracta1_78_; 
wire fracta1_79_; 
wire fracta1_7_; 
wire fracta1_80_; 
wire fracta1_81_; 
wire fracta1_82_; 
wire fracta1_83_; 
wire fracta1_84_; 
wire fracta1_85_; 
wire fracta1_86_; 
wire fracta1_87_; 
wire fracta1_88_; 
wire fracta1_89_; 
wire fracta1_8_; 
wire fracta1_90_; 
wire fracta1_91_; 
wire fracta1_92_; 
wire fracta1_93_; 
wire fracta1_94_; 
wire fracta1_95_; 
wire fracta1_96_; 
wire fracta1_97_; 
wire fracta1_98_; 
wire fracta1_99_; 
wire fracta1_9_; 
wire fracta_112_; 
input ld;
output \o[0] ;
output \o[100] ;
output \o[101] ;
output \o[102] ;
output \o[103] ;
output \o[104] ;
output \o[105] ;
output \o[106] ;
output \o[107] ;
output \o[108] ;
output \o[109] ;
output \o[10] ;
output \o[110] ;
output \o[111] ;
output \o[112] ;
output \o[113] ;
output \o[114] ;
output \o[115] ;
output \o[116] ;
output \o[117] ;
output \o[118] ;
output \o[119] ;
output \o[11] ;
output \o[120] ;
output \o[121] ;
output \o[122] ;
output \o[123] ;
output \o[124] ;
output \o[125] ;
output \o[126] ;
output \o[127] ;
output \o[128] ;
output \o[129] ;
output \o[12] ;
output \o[130] ;
output \o[131] ;
output \o[132] ;
output \o[133] ;
output \o[134] ;
output \o[135] ;
output \o[136] ;
output \o[137] ;
output \o[138] ;
output \o[139] ;
output \o[13] ;
output \o[140] ;
output \o[141] ;
output \o[142] ;
output \o[143] ;
output \o[144] ;
output \o[145] ;
output \o[146] ;
output \o[147] ;
output \o[148] ;
output \o[149] ;
output \o[14] ;
output \o[150] ;
output \o[151] ;
output \o[152] ;
output \o[153] ;
output \o[154] ;
output \o[155] ;
output \o[156] ;
output \o[157] ;
output \o[158] ;
output \o[159] ;
output \o[15] ;
output \o[160] ;
output \o[161] ;
output \o[162] ;
output \o[163] ;
output \o[164] ;
output \o[165] ;
output \o[166] ;
output \o[167] ;
output \o[168] ;
output \o[169] ;
output \o[16] ;
output \o[170] ;
output \o[171] ;
output \o[172] ;
output \o[173] ;
output \o[174] ;
output \o[175] ;
output \o[176] ;
output \o[177] ;
output \o[178] ;
output \o[179] ;
output \o[17] ;
output \o[180] ;
output \o[181] ;
output \o[182] ;
output \o[183] ;
output \o[184] ;
output \o[185] ;
output \o[186] ;
output \o[187] ;
output \o[188] ;
output \o[189] ;
output \o[18] ;
output \o[190] ;
output \o[191] ;
output \o[192] ;
output \o[193] ;
output \o[194] ;
output \o[195] ;
output \o[196] ;
output \o[197] ;
output \o[198] ;
output \o[199] ;
output \o[19] ;
output \o[1] ;
output \o[200] ;
output \o[201] ;
output \o[202] ;
output \o[203] ;
output \o[204] ;
output \o[205] ;
output \o[206] ;
output \o[207] ;
output \o[208] ;
output \o[209] ;
output \o[20] ;
output \o[210] ;
output \o[211] ;
output \o[212] ;
output \o[213] ;
output \o[214] ;
output \o[215] ;
output \o[216] ;
output \o[217] ;
output \o[218] ;
output \o[219] ;
output \o[21] ;
output \o[220] ;
output \o[221] ;
output \o[222] ;
output \o[223] ;
output \o[224] ;
output \o[225] ;
output \o[226] ;
output \o[227] ;
output \o[228] ;
output \o[229] ;
output \o[22] ;
output \o[230] ;
output \o[231] ;
output \o[232] ;
output \o[233] ;
output \o[234] ;
output \o[235] ;
output \o[236] ;
output \o[237] ;
output \o[238] ;
output \o[239] ;
output \o[23] ;
output \o[240] ;
output \o[241] ;
output \o[24] ;
output \o[25] ;
output \o[26] ;
output \o[27] ;
output \o[28] ;
output \o[29] ;
output \o[2] ;
output \o[30] ;
output \o[31] ;
output \o[32] ;
output \o[33] ;
output \o[34] ;
output \o[35] ;
output \o[36] ;
output \o[37] ;
output \o[38] ;
output \o[39] ;
output \o[3] ;
output \o[40] ;
output \o[41] ;
output \o[42] ;
output \o[43] ;
output \o[44] ;
output \o[45] ;
output \o[46] ;
output \o[47] ;
output \o[48] ;
output \o[49] ;
output \o[4] ;
output \o[50] ;
output \o[51] ;
output \o[52] ;
output \o[53] ;
output \o[54] ;
output \o[55] ;
output \o[56] ;
output \o[57] ;
output \o[58] ;
output \o[59] ;
output \o[5] ;
output \o[60] ;
output \o[61] ;
output \o[62] ;
output \o[63] ;
output \o[64] ;
output \o[65] ;
output \o[66] ;
output \o[67] ;
output \o[68] ;
output \o[69] ;
output \o[6] ;
output \o[70] ;
output \o[71] ;
output \o[72] ;
output \o[73] ;
output \o[74] ;
output \o[75] ;
output \o[76] ;
output \o[77] ;
output \o[78] ;
output \o[79] ;
output \o[7] ;
output \o[80] ;
output \o[81] ;
output \o[82] ;
output \o[83] ;
output \o[84] ;
output \o[85] ;
output \o[86] ;
output \o[87] ;
output \o[88] ;
output \o[89] ;
output \o[8] ;
output \o[90] ;
output \o[91] ;
output \o[92] ;
output \o[93] ;
output \o[94] ;
output \o[95] ;
output \o[96] ;
output \o[97] ;
output \o[98] ;
output \o[99] ;
output \o[9] ;
input rst;
wire sqrto_0_; 
wire sqrto_100_; 
wire sqrto_101_; 
wire sqrto_102_; 
wire sqrto_103_; 
wire sqrto_104_; 
wire sqrto_105_; 
wire sqrto_106_; 
wire sqrto_107_; 
wire sqrto_108_; 
wire sqrto_109_; 
wire sqrto_10_; 
wire sqrto_110_; 
wire sqrto_111_; 
wire sqrto_112_; 
wire sqrto_113_; 
wire sqrto_114_; 
wire sqrto_115_; 
wire sqrto_116_; 
wire sqrto_117_; 
wire sqrto_118_; 
wire sqrto_119_; 
wire sqrto_11_; 
wire sqrto_120_; 
wire sqrto_121_; 
wire sqrto_122_; 
wire sqrto_123_; 
wire sqrto_124_; 
wire sqrto_125_; 
wire sqrto_126_; 
wire sqrto_127_; 
wire sqrto_128_; 
wire sqrto_129_; 
wire sqrto_12_; 
wire sqrto_130_; 
wire sqrto_131_; 
wire sqrto_132_; 
wire sqrto_133_; 
wire sqrto_134_; 
wire sqrto_135_; 
wire sqrto_136_; 
wire sqrto_137_; 
wire sqrto_138_; 
wire sqrto_139_; 
wire sqrto_13_; 
wire sqrto_140_; 
wire sqrto_141_; 
wire sqrto_142_; 
wire sqrto_143_; 
wire sqrto_144_; 
wire sqrto_145_; 
wire sqrto_146_; 
wire sqrto_147_; 
wire sqrto_148_; 
wire sqrto_149_; 
wire sqrto_14_; 
wire sqrto_150_; 
wire sqrto_151_; 
wire sqrto_152_; 
wire sqrto_153_; 
wire sqrto_154_; 
wire sqrto_155_; 
wire sqrto_156_; 
wire sqrto_157_; 
wire sqrto_158_; 
wire sqrto_159_; 
wire sqrto_15_; 
wire sqrto_160_; 
wire sqrto_161_; 
wire sqrto_162_; 
wire sqrto_163_; 
wire sqrto_164_; 
wire sqrto_165_; 
wire sqrto_166_; 
wire sqrto_167_; 
wire sqrto_168_; 
wire sqrto_169_; 
wire sqrto_16_; 
wire sqrto_170_; 
wire sqrto_171_; 
wire sqrto_172_; 
wire sqrto_173_; 
wire sqrto_174_; 
wire sqrto_175_; 
wire sqrto_176_; 
wire sqrto_177_; 
wire sqrto_178_; 
wire sqrto_179_; 
wire sqrto_17_; 
wire sqrto_180_; 
wire sqrto_181_; 
wire sqrto_182_; 
wire sqrto_183_; 
wire sqrto_184_; 
wire sqrto_185_; 
wire sqrto_186_; 
wire sqrto_187_; 
wire sqrto_188_; 
wire sqrto_189_; 
wire sqrto_18_; 
wire sqrto_190_; 
wire sqrto_191_; 
wire sqrto_192_; 
wire sqrto_193_; 
wire sqrto_194_; 
wire sqrto_195_; 
wire sqrto_196_; 
wire sqrto_197_; 
wire sqrto_198_; 
wire sqrto_199_; 
wire sqrto_19_; 
wire sqrto_1_; 
wire sqrto_200_; 
wire sqrto_201_; 
wire sqrto_202_; 
wire sqrto_203_; 
wire sqrto_204_; 
wire sqrto_205_; 
wire sqrto_206_; 
wire sqrto_207_; 
wire sqrto_208_; 
wire sqrto_209_; 
wire sqrto_20_; 
wire sqrto_210_; 
wire sqrto_211_; 
wire sqrto_212_; 
wire sqrto_213_; 
wire sqrto_214_; 
wire sqrto_215_; 
wire sqrto_216_; 
wire sqrto_217_; 
wire sqrto_218_; 
wire sqrto_219_; 
wire sqrto_21_; 
wire sqrto_220_; 
wire sqrto_221_; 
wire sqrto_222_; 
wire sqrto_223_; 
wire sqrto_224_; 
wire sqrto_225_; 
wire sqrto_22_; 
wire sqrto_23_; 
wire sqrto_24_; 
wire sqrto_25_; 
wire sqrto_26_; 
wire sqrto_27_; 
wire sqrto_28_; 
wire sqrto_29_; 
wire sqrto_2_; 
wire sqrto_30_; 
wire sqrto_31_; 
wire sqrto_32_; 
wire sqrto_33_; 
wire sqrto_34_; 
wire sqrto_35_; 
wire sqrto_36_; 
wire sqrto_37_; 
wire sqrto_38_; 
wire sqrto_39_; 
wire sqrto_3_; 
wire sqrto_40_; 
wire sqrto_41_; 
wire sqrto_42_; 
wire sqrto_43_; 
wire sqrto_44_; 
wire sqrto_45_; 
wire sqrto_46_; 
wire sqrto_47_; 
wire sqrto_48_; 
wire sqrto_49_; 
wire sqrto_4_; 
wire sqrto_50_; 
wire sqrto_51_; 
wire sqrto_52_; 
wire sqrto_53_; 
wire sqrto_54_; 
wire sqrto_55_; 
wire sqrto_56_; 
wire sqrto_57_; 
wire sqrto_58_; 
wire sqrto_59_; 
wire sqrto_5_; 
wire sqrto_60_; 
wire sqrto_61_; 
wire sqrto_62_; 
wire sqrto_63_; 
wire sqrto_64_; 
wire sqrto_65_; 
wire sqrto_66_; 
wire sqrto_67_; 
wire sqrto_68_; 
wire sqrto_69_; 
wire sqrto_6_; 
wire sqrto_70_; 
wire sqrto_71_; 
wire sqrto_72_; 
wire sqrto_73_; 
wire sqrto_74_; 
wire sqrto_75_; 
wire sqrto_76_; 
wire sqrto_77_; 
wire sqrto_78_; 
wire sqrto_79_; 
wire sqrto_7_; 
wire sqrto_80_; 
wire sqrto_81_; 
wire sqrto_82_; 
wire sqrto_83_; 
wire sqrto_84_; 
wire sqrto_85_; 
wire sqrto_86_; 
wire sqrto_87_; 
wire sqrto_88_; 
wire sqrto_89_; 
wire sqrto_8_; 
wire sqrto_90_; 
wire sqrto_91_; 
wire sqrto_92_; 
wire sqrto_93_; 
wire sqrto_94_; 
wire sqrto_95_; 
wire sqrto_96_; 
wire sqrto_97_; 
wire sqrto_98_; 
wire sqrto_99_; 
wire sqrto_9_; 
wire u1__abc_51895_new_n137_; 
wire u1__abc_51895_new_n138_; 
wire u1__abc_51895_new_n139_; 
wire u1__abc_51895_new_n140_; 
wire u1__abc_51895_new_n141_; 
wire u1__abc_51895_new_n142_; 
wire u1__abc_51895_new_n143_; 
wire u1__abc_51895_new_n144_; 
wire u1__abc_51895_new_n145_; 
wire u1__abc_51895_new_n146_; 
wire u1__abc_51895_new_n147_; 
wire u1__abc_51895_new_n148_; 
wire u1__abc_51895_new_n149_; 
wire u1__abc_51895_new_n152_; 
wire u1__abc_51895_new_n153_; 
wire u1__abc_51895_new_n154_; 
wire u1__abc_51895_new_n155_; 
wire u1__abc_51895_new_n156_; 
wire u1__abc_51895_new_n157_; 
wire u1__abc_51895_new_n158_; 
wire u1__abc_51895_new_n159_; 
wire u1__abc_51895_new_n160_; 
wire u1__abc_51895_new_n161_; 
wire u1__abc_51895_new_n162_; 
wire u1__abc_51895_new_n163_; 
wire u1__abc_51895_new_n164_; 
wire u1__abc_51895_new_n166_; 
wire u1__abc_51895_new_n167_; 
wire u1__abc_51895_new_n168_; 
wire u1__abc_51895_new_n169_; 
wire u1__abc_51895_new_n170_; 
wire u1__abc_51895_new_n171_; 
wire u1__abc_51895_new_n172_; 
wire u1__abc_51895_new_n173_; 
wire u1__abc_51895_new_n174_; 
wire u1__abc_51895_new_n175_; 
wire u1__abc_51895_new_n176_; 
wire u1__abc_51895_new_n177_; 
wire u1__abc_51895_new_n178_; 
wire u1__abc_51895_new_n179_; 
wire u1__abc_51895_new_n180_; 
wire u1__abc_51895_new_n181_; 
wire u1__abc_51895_new_n182_; 
wire u1__abc_51895_new_n183_; 
wire u1__abc_51895_new_n184_; 
wire u1__abc_51895_new_n185_; 
wire u1__abc_51895_new_n186_; 
wire u1__abc_51895_new_n187_; 
wire u1__abc_51895_new_n188_; 
wire u1__abc_51895_new_n189_; 
wire u1__abc_51895_new_n190_; 
wire u1__abc_51895_new_n191_; 
wire u1__abc_51895_new_n192_; 
wire u1__abc_51895_new_n193_; 
wire u1__abc_51895_new_n194_; 
wire u1__abc_51895_new_n195_; 
wire u1__abc_51895_new_n196_; 
wire u1__abc_51895_new_n197_; 
wire u1__abc_51895_new_n198_; 
wire u1__abc_51895_new_n199_; 
wire u1__abc_51895_new_n200_; 
wire u1__abc_51895_new_n201_; 
wire u1__abc_51895_new_n202_; 
wire u1__abc_51895_new_n203_; 
wire u1__abc_51895_new_n204_; 
wire u1__abc_51895_new_n205_; 
wire u1__abc_51895_new_n206_; 
wire u1__abc_51895_new_n207_; 
wire u1__abc_51895_new_n208_; 
wire u1__abc_51895_new_n209_; 
wire u1__abc_51895_new_n210_; 
wire u1__abc_51895_new_n211_; 
wire u1__abc_51895_new_n212_; 
wire u1__abc_51895_new_n213_; 
wire u1__abc_51895_new_n214_; 
wire u1__abc_51895_new_n215_; 
wire u1__abc_51895_new_n216_; 
wire u1__abc_51895_new_n217_; 
wire u1__abc_51895_new_n218_; 
wire u1__abc_51895_new_n219_; 
wire u1__abc_51895_new_n220_; 
wire u1__abc_51895_new_n221_; 
wire u1__abc_51895_new_n222_; 
wire u1__abc_51895_new_n223_; 
wire u1__abc_51895_new_n224_; 
wire u1__abc_51895_new_n225_; 
wire u1__abc_51895_new_n226_; 
wire u1__abc_51895_new_n227_; 
wire u1__abc_51895_new_n228_; 
wire u1__abc_51895_new_n229_; 
wire u1__abc_51895_new_n230_; 
wire u1__abc_51895_new_n231_; 
wire u1__abc_51895_new_n232_; 
wire u1__abc_51895_new_n233_; 
wire u1__abc_51895_new_n234_; 
wire u1__abc_51895_new_n235_; 
wire u1__abc_51895_new_n236_; 
wire u1__abc_51895_new_n237_; 
wire u1__abc_51895_new_n238_; 
wire u1__abc_51895_new_n239_; 
wire u1__abc_51895_new_n240_; 
wire u1__abc_51895_new_n241_; 
wire u1__abc_51895_new_n242_; 
wire u1__abc_51895_new_n243_; 
wire u1__abc_51895_new_n244_; 
wire u1__abc_51895_new_n245_; 
wire u1__abc_51895_new_n246_; 
wire u1__abc_51895_new_n247_; 
wire u1__abc_51895_new_n248_; 
wire u1__abc_51895_new_n249_; 
wire u1__abc_51895_new_n250_; 
wire u1__abc_51895_new_n251_; 
wire u1__abc_51895_new_n252_; 
wire u1__abc_51895_new_n253_; 
wire u1__abc_51895_new_n254_; 
wire u1__abc_51895_new_n255_; 
wire u1__abc_51895_new_n256_; 
wire u1__abc_51895_new_n257_; 
wire u1__abc_51895_new_n258_; 
wire u1__abc_51895_new_n259_; 
wire u1__abc_51895_new_n260_; 
wire u1__abc_51895_new_n261_; 
wire u1__abc_51895_new_n262_; 
wire u1__abc_51895_new_n263_; 
wire u1__abc_51895_new_n264_; 
wire u1__abc_51895_new_n265_; 
wire u1__abc_51895_new_n266_; 
wire u1__abc_51895_new_n267_; 
wire u1__abc_51895_new_n268_; 
wire u1__abc_51895_new_n269_; 
wire u1__abc_51895_new_n270_; 
wire u1__abc_51895_new_n271_; 
wire u1__abc_51895_new_n272_; 
wire u1__abc_51895_new_n273_; 
wire u1__abc_51895_new_n274_; 
wire u1__abc_51895_new_n275_; 
wire u1__abc_51895_new_n276_; 
wire u1__abc_51895_new_n277_; 
wire u1__abc_51895_new_n278_; 
wire u1__abc_51895_new_n279_; 
wire u1__abc_51895_new_n280_; 
wire u1__abc_51895_new_n281_; 
wire u1__abc_51895_new_n282_; 
wire u1__abc_51895_new_n283_; 
wire u1__abc_51895_new_n284_; 
wire u1__abc_51895_new_n285_; 
wire u1__abc_51895_new_n286_; 
wire u1__abc_51895_new_n287_; 
wire u1__abc_51895_new_n288_; 
wire u1__abc_51895_new_n289_; 
wire u1__abc_51895_new_n290_; 
wire u1__abc_51895_new_n291_; 
wire u1__abc_51895_new_n292_; 
wire u1__abc_51895_new_n293_; 
wire u1__abc_51895_new_n294_; 
wire u1__abc_51895_new_n295_; 
wire u1__abc_51895_new_n296_; 
wire u1__abc_51895_new_n297_; 
wire u1__abc_51895_new_n298_; 
wire u1__abc_51895_new_n299_; 
wire u1__abc_51895_new_n300_; 
wire u1__abc_51895_new_n301_; 
wire u1__abc_51895_new_n302_; 
wire u1__abc_51895_new_n303_; 
wire u1__abc_51895_new_n304_; 
wire u1__abc_51895_new_n305_; 
wire u1__abc_51895_new_n306_; 
wire u1__abc_51895_new_n307_; 
wire u1__abc_51895_new_n308_; 
wire u1__abc_51895_new_n309_; 
wire u1__abc_51895_new_n310_; 
wire u1__abc_51895_new_n311_; 
wire u1__abc_51895_new_n312_; 
wire u1__abc_51895_new_n313_; 
wire u1__abc_51895_new_n314_; 
wire u1__abc_51895_new_n315_; 
wire u1__abc_51895_new_n316_; 
wire u1__abc_51895_new_n317_; 
wire u1__abc_51895_new_n318_; 
wire u1__abc_51895_new_n319_; 
wire u1__abc_51895_new_n320_; 
wire u1__abc_51895_new_n321_; 
wire u1__abc_51895_new_n322_; 
wire u1__abc_51895_new_n323_; 
wire u1__abc_51895_new_n324_; 
wire u1__abc_51895_new_n325_; 
wire u1__abc_51895_new_n326_; 
wire u1__abc_51895_new_n327_; 
wire u1__abc_51895_new_n328_; 
wire u1__abc_51895_new_n329_; 
wire u1__abc_51895_new_n330_; 
wire u1__abc_51895_new_n331_; 
wire u1__abc_51895_new_n332_; 
wire u1__abc_51895_new_n333_; 
wire u1__abc_51895_new_n334_; 
wire u1__abc_51895_new_n335_; 
wire u1__abc_51895_new_n336_; 
wire u1__abc_51895_new_n337_; 
wire u1__abc_51895_new_n338_; 
wire u1__abc_51895_new_n339_; 
wire u1__abc_51895_new_n340_; 
wire u1__abc_51895_new_n341_; 
wire u1__abc_51895_new_n342_; 
wire u1__abc_51895_new_n343_; 
wire u1__abc_51895_new_n344_; 
wire u1__abc_51895_new_n345_; 
wire u1__abc_51895_new_n346_; 
wire u1__abc_51895_new_n347_; 
wire u1__abc_51895_new_n348_; 
wire u1__abc_51895_new_n349_; 
wire u1__abc_51895_new_n350_; 
wire u1__abc_51895_new_n351_; 
wire u1__abc_51895_new_n352_; 
wire u1__abc_51895_new_n353_; 
wire u1__abc_51895_new_n354_; 
wire u1__abc_51895_new_n355_; 
wire u1__abc_51895_new_n356_; 
wire u1__abc_51895_new_n357_; 
wire u1__abc_51895_new_n358_; 
wire u1__abc_51895_new_n359_; 
wire u1__abc_51895_new_n360_; 
wire u1__abc_51895_new_n361_; 
wire u1__abc_51895_new_n362_; 
wire u1__abc_51895_new_n363_; 
wire u1__abc_51895_new_n364_; 
wire u1__abc_51895_new_n365_; 
wire u1__abc_51895_new_n366_; 
wire u1__abc_51895_new_n367_; 
wire u1__abc_51895_new_n368_; 
wire u1__abc_51895_new_n369_; 
wire u1__abc_51895_new_n370_; 
wire u1__abc_51895_new_n371_; 
wire u1__abc_51895_new_n372_; 
wire u1__abc_51895_new_n373_; 
wire u1__abc_51895_new_n374_; 
wire u1__abc_51895_new_n375_; 
wire u1__abc_51895_new_n376_; 
wire u1__abc_51895_new_n377_; 
wire u1__abc_51895_new_n378_; 
wire u1__abc_51895_new_n379_; 
wire u1__abc_51895_new_n380_; 
wire u1__abc_51895_new_n381_; 
wire u1__abc_51895_new_n382_; 
wire u1__abc_51895_new_n383_; 
wire u1__abc_51895_new_n384_; 
wire u1__abc_51895_new_n385_; 
wire u1__abc_51895_new_n386_; 
wire u1__abc_51895_new_n387_; 
wire u1__abc_51895_new_n392_; 
wire u1_mz; 
wire u1_xinf; 
wire u2__0cnt_7_0__0_; 
wire u2__0cnt_7_0__1_; 
wire u2__0cnt_7_0__2_; 
wire u2__0cnt_7_0__3_; 
wire u2__0cnt_7_0__4_; 
wire u2__0cnt_7_0__5_; 
wire u2__0cnt_7_0__6_; 
wire u2__0cnt_7_0__7_; 
wire u2__0remHi_451_0__0_; 
wire u2__0remHi_451_0__100_; 
wire u2__0remHi_451_0__101_; 
wire u2__0remHi_451_0__102_; 
wire u2__0remHi_451_0__103_; 
wire u2__0remHi_451_0__104_; 
wire u2__0remHi_451_0__105_; 
wire u2__0remHi_451_0__106_; 
wire u2__0remHi_451_0__107_; 
wire u2__0remHi_451_0__108_; 
wire u2__0remHi_451_0__109_; 
wire u2__0remHi_451_0__10_; 
wire u2__0remHi_451_0__110_; 
wire u2__0remHi_451_0__111_; 
wire u2__0remHi_451_0__112_; 
wire u2__0remHi_451_0__113_; 
wire u2__0remHi_451_0__114_; 
wire u2__0remHi_451_0__115_; 
wire u2__0remHi_451_0__116_; 
wire u2__0remHi_451_0__117_; 
wire u2__0remHi_451_0__118_; 
wire u2__0remHi_451_0__119_; 
wire u2__0remHi_451_0__11_; 
wire u2__0remHi_451_0__120_; 
wire u2__0remHi_451_0__121_; 
wire u2__0remHi_451_0__122_; 
wire u2__0remHi_451_0__123_; 
wire u2__0remHi_451_0__124_; 
wire u2__0remHi_451_0__125_; 
wire u2__0remHi_451_0__126_; 
wire u2__0remHi_451_0__127_; 
wire u2__0remHi_451_0__128_; 
wire u2__0remHi_451_0__129_; 
wire u2__0remHi_451_0__12_; 
wire u2__0remHi_451_0__130_; 
wire u2__0remHi_451_0__131_; 
wire u2__0remHi_451_0__132_; 
wire u2__0remHi_451_0__133_; 
wire u2__0remHi_451_0__134_; 
wire u2__0remHi_451_0__135_; 
wire u2__0remHi_451_0__136_; 
wire u2__0remHi_451_0__137_; 
wire u2__0remHi_451_0__138_; 
wire u2__0remHi_451_0__139_; 
wire u2__0remHi_451_0__13_; 
wire u2__0remHi_451_0__140_; 
wire u2__0remHi_451_0__141_; 
wire u2__0remHi_451_0__142_; 
wire u2__0remHi_451_0__143_; 
wire u2__0remHi_451_0__144_; 
wire u2__0remHi_451_0__145_; 
wire u2__0remHi_451_0__146_; 
wire u2__0remHi_451_0__147_; 
wire u2__0remHi_451_0__148_; 
wire u2__0remHi_451_0__149_; 
wire u2__0remHi_451_0__14_; 
wire u2__0remHi_451_0__150_; 
wire u2__0remHi_451_0__151_; 
wire u2__0remHi_451_0__152_; 
wire u2__0remHi_451_0__153_; 
wire u2__0remHi_451_0__154_; 
wire u2__0remHi_451_0__155_; 
wire u2__0remHi_451_0__156_; 
wire u2__0remHi_451_0__157_; 
wire u2__0remHi_451_0__158_; 
wire u2__0remHi_451_0__159_; 
wire u2__0remHi_451_0__15_; 
wire u2__0remHi_451_0__160_; 
wire u2__0remHi_451_0__161_; 
wire u2__0remHi_451_0__162_; 
wire u2__0remHi_451_0__163_; 
wire u2__0remHi_451_0__164_; 
wire u2__0remHi_451_0__165_; 
wire u2__0remHi_451_0__166_; 
wire u2__0remHi_451_0__167_; 
wire u2__0remHi_451_0__168_; 
wire u2__0remHi_451_0__169_; 
wire u2__0remHi_451_0__16_; 
wire u2__0remHi_451_0__170_; 
wire u2__0remHi_451_0__171_; 
wire u2__0remHi_451_0__172_; 
wire u2__0remHi_451_0__173_; 
wire u2__0remHi_451_0__174_; 
wire u2__0remHi_451_0__175_; 
wire u2__0remHi_451_0__176_; 
wire u2__0remHi_451_0__177_; 
wire u2__0remHi_451_0__178_; 
wire u2__0remHi_451_0__179_; 
wire u2__0remHi_451_0__17_; 
wire u2__0remHi_451_0__180_; 
wire u2__0remHi_451_0__181_; 
wire u2__0remHi_451_0__182_; 
wire u2__0remHi_451_0__183_; 
wire u2__0remHi_451_0__184_; 
wire u2__0remHi_451_0__185_; 
wire u2__0remHi_451_0__186_; 
wire u2__0remHi_451_0__187_; 
wire u2__0remHi_451_0__188_; 
wire u2__0remHi_451_0__189_; 
wire u2__0remHi_451_0__18_; 
wire u2__0remHi_451_0__190_; 
wire u2__0remHi_451_0__191_; 
wire u2__0remHi_451_0__192_; 
wire u2__0remHi_451_0__193_; 
wire u2__0remHi_451_0__194_; 
wire u2__0remHi_451_0__195_; 
wire u2__0remHi_451_0__196_; 
wire u2__0remHi_451_0__197_; 
wire u2__0remHi_451_0__198_; 
wire u2__0remHi_451_0__199_; 
wire u2__0remHi_451_0__19_; 
wire u2__0remHi_451_0__1_; 
wire u2__0remHi_451_0__200_; 
wire u2__0remHi_451_0__201_; 
wire u2__0remHi_451_0__202_; 
wire u2__0remHi_451_0__203_; 
wire u2__0remHi_451_0__204_; 
wire u2__0remHi_451_0__205_; 
wire u2__0remHi_451_0__206_; 
wire u2__0remHi_451_0__207_; 
wire u2__0remHi_451_0__208_; 
wire u2__0remHi_451_0__209_; 
wire u2__0remHi_451_0__20_; 
wire u2__0remHi_451_0__210_; 
wire u2__0remHi_451_0__211_; 
wire u2__0remHi_451_0__212_; 
wire u2__0remHi_451_0__213_; 
wire u2__0remHi_451_0__214_; 
wire u2__0remHi_451_0__215_; 
wire u2__0remHi_451_0__216_; 
wire u2__0remHi_451_0__217_; 
wire u2__0remHi_451_0__218_; 
wire u2__0remHi_451_0__219_; 
wire u2__0remHi_451_0__21_; 
wire u2__0remHi_451_0__220_; 
wire u2__0remHi_451_0__221_; 
wire u2__0remHi_451_0__222_; 
wire u2__0remHi_451_0__223_; 
wire u2__0remHi_451_0__224_; 
wire u2__0remHi_451_0__225_; 
wire u2__0remHi_451_0__226_; 
wire u2__0remHi_451_0__227_; 
wire u2__0remHi_451_0__228_; 
wire u2__0remHi_451_0__229_; 
wire u2__0remHi_451_0__22_; 
wire u2__0remHi_451_0__230_; 
wire u2__0remHi_451_0__231_; 
wire u2__0remHi_451_0__232_; 
wire u2__0remHi_451_0__233_; 
wire u2__0remHi_451_0__234_; 
wire u2__0remHi_451_0__235_; 
wire u2__0remHi_451_0__236_; 
wire u2__0remHi_451_0__237_; 
wire u2__0remHi_451_0__238_; 
wire u2__0remHi_451_0__239_; 
wire u2__0remHi_451_0__23_; 
wire u2__0remHi_451_0__240_; 
wire u2__0remHi_451_0__241_; 
wire u2__0remHi_451_0__242_; 
wire u2__0remHi_451_0__243_; 
wire u2__0remHi_451_0__244_; 
wire u2__0remHi_451_0__245_; 
wire u2__0remHi_451_0__246_; 
wire u2__0remHi_451_0__247_; 
wire u2__0remHi_451_0__248_; 
wire u2__0remHi_451_0__249_; 
wire u2__0remHi_451_0__24_; 
wire u2__0remHi_451_0__250_; 
wire u2__0remHi_451_0__251_; 
wire u2__0remHi_451_0__252_; 
wire u2__0remHi_451_0__253_; 
wire u2__0remHi_451_0__254_; 
wire u2__0remHi_451_0__255_; 
wire u2__0remHi_451_0__256_; 
wire u2__0remHi_451_0__257_; 
wire u2__0remHi_451_0__258_; 
wire u2__0remHi_451_0__259_; 
wire u2__0remHi_451_0__25_; 
wire u2__0remHi_451_0__260_; 
wire u2__0remHi_451_0__261_; 
wire u2__0remHi_451_0__262_; 
wire u2__0remHi_451_0__263_; 
wire u2__0remHi_451_0__264_; 
wire u2__0remHi_451_0__265_; 
wire u2__0remHi_451_0__266_; 
wire u2__0remHi_451_0__267_; 
wire u2__0remHi_451_0__268_; 
wire u2__0remHi_451_0__269_; 
wire u2__0remHi_451_0__26_; 
wire u2__0remHi_451_0__270_; 
wire u2__0remHi_451_0__271_; 
wire u2__0remHi_451_0__272_; 
wire u2__0remHi_451_0__273_; 
wire u2__0remHi_451_0__274_; 
wire u2__0remHi_451_0__275_; 
wire u2__0remHi_451_0__276_; 
wire u2__0remHi_451_0__277_; 
wire u2__0remHi_451_0__278_; 
wire u2__0remHi_451_0__279_; 
wire u2__0remHi_451_0__27_; 
wire u2__0remHi_451_0__280_; 
wire u2__0remHi_451_0__281_; 
wire u2__0remHi_451_0__282_; 
wire u2__0remHi_451_0__283_; 
wire u2__0remHi_451_0__284_; 
wire u2__0remHi_451_0__285_; 
wire u2__0remHi_451_0__286_; 
wire u2__0remHi_451_0__287_; 
wire u2__0remHi_451_0__288_; 
wire u2__0remHi_451_0__289_; 
wire u2__0remHi_451_0__28_; 
wire u2__0remHi_451_0__290_; 
wire u2__0remHi_451_0__291_; 
wire u2__0remHi_451_0__292_; 
wire u2__0remHi_451_0__293_; 
wire u2__0remHi_451_0__294_; 
wire u2__0remHi_451_0__295_; 
wire u2__0remHi_451_0__296_; 
wire u2__0remHi_451_0__297_; 
wire u2__0remHi_451_0__298_; 
wire u2__0remHi_451_0__299_; 
wire u2__0remHi_451_0__29_; 
wire u2__0remHi_451_0__2_; 
wire u2__0remHi_451_0__300_; 
wire u2__0remHi_451_0__301_; 
wire u2__0remHi_451_0__302_; 
wire u2__0remHi_451_0__303_; 
wire u2__0remHi_451_0__304_; 
wire u2__0remHi_451_0__305_; 
wire u2__0remHi_451_0__306_; 
wire u2__0remHi_451_0__307_; 
wire u2__0remHi_451_0__308_; 
wire u2__0remHi_451_0__309_; 
wire u2__0remHi_451_0__30_; 
wire u2__0remHi_451_0__310_; 
wire u2__0remHi_451_0__311_; 
wire u2__0remHi_451_0__312_; 
wire u2__0remHi_451_0__313_; 
wire u2__0remHi_451_0__314_; 
wire u2__0remHi_451_0__315_; 
wire u2__0remHi_451_0__316_; 
wire u2__0remHi_451_0__317_; 
wire u2__0remHi_451_0__318_; 
wire u2__0remHi_451_0__319_; 
wire u2__0remHi_451_0__31_; 
wire u2__0remHi_451_0__320_; 
wire u2__0remHi_451_0__321_; 
wire u2__0remHi_451_0__322_; 
wire u2__0remHi_451_0__323_; 
wire u2__0remHi_451_0__324_; 
wire u2__0remHi_451_0__325_; 
wire u2__0remHi_451_0__326_; 
wire u2__0remHi_451_0__327_; 
wire u2__0remHi_451_0__328_; 
wire u2__0remHi_451_0__329_; 
wire u2__0remHi_451_0__32_; 
wire u2__0remHi_451_0__330_; 
wire u2__0remHi_451_0__331_; 
wire u2__0remHi_451_0__332_; 
wire u2__0remHi_451_0__333_; 
wire u2__0remHi_451_0__334_; 
wire u2__0remHi_451_0__335_; 
wire u2__0remHi_451_0__336_; 
wire u2__0remHi_451_0__337_; 
wire u2__0remHi_451_0__338_; 
wire u2__0remHi_451_0__339_; 
wire u2__0remHi_451_0__33_; 
wire u2__0remHi_451_0__340_; 
wire u2__0remHi_451_0__341_; 
wire u2__0remHi_451_0__342_; 
wire u2__0remHi_451_0__343_; 
wire u2__0remHi_451_0__344_; 
wire u2__0remHi_451_0__345_; 
wire u2__0remHi_451_0__346_; 
wire u2__0remHi_451_0__347_; 
wire u2__0remHi_451_0__348_; 
wire u2__0remHi_451_0__349_; 
wire u2__0remHi_451_0__34_; 
wire u2__0remHi_451_0__350_; 
wire u2__0remHi_451_0__351_; 
wire u2__0remHi_451_0__352_; 
wire u2__0remHi_451_0__353_; 
wire u2__0remHi_451_0__354_; 
wire u2__0remHi_451_0__355_; 
wire u2__0remHi_451_0__356_; 
wire u2__0remHi_451_0__357_; 
wire u2__0remHi_451_0__358_; 
wire u2__0remHi_451_0__359_; 
wire u2__0remHi_451_0__35_; 
wire u2__0remHi_451_0__360_; 
wire u2__0remHi_451_0__361_; 
wire u2__0remHi_451_0__362_; 
wire u2__0remHi_451_0__363_; 
wire u2__0remHi_451_0__364_; 
wire u2__0remHi_451_0__365_; 
wire u2__0remHi_451_0__366_; 
wire u2__0remHi_451_0__367_; 
wire u2__0remHi_451_0__368_; 
wire u2__0remHi_451_0__369_; 
wire u2__0remHi_451_0__36_; 
wire u2__0remHi_451_0__370_; 
wire u2__0remHi_451_0__371_; 
wire u2__0remHi_451_0__372_; 
wire u2__0remHi_451_0__373_; 
wire u2__0remHi_451_0__374_; 
wire u2__0remHi_451_0__375_; 
wire u2__0remHi_451_0__376_; 
wire u2__0remHi_451_0__377_; 
wire u2__0remHi_451_0__378_; 
wire u2__0remHi_451_0__379_; 
wire u2__0remHi_451_0__37_; 
wire u2__0remHi_451_0__380_; 
wire u2__0remHi_451_0__381_; 
wire u2__0remHi_451_0__382_; 
wire u2__0remHi_451_0__383_; 
wire u2__0remHi_451_0__384_; 
wire u2__0remHi_451_0__385_; 
wire u2__0remHi_451_0__386_; 
wire u2__0remHi_451_0__387_; 
wire u2__0remHi_451_0__388_; 
wire u2__0remHi_451_0__389_; 
wire u2__0remHi_451_0__38_; 
wire u2__0remHi_451_0__390_; 
wire u2__0remHi_451_0__391_; 
wire u2__0remHi_451_0__392_; 
wire u2__0remHi_451_0__393_; 
wire u2__0remHi_451_0__394_; 
wire u2__0remHi_451_0__395_; 
wire u2__0remHi_451_0__396_; 
wire u2__0remHi_451_0__397_; 
wire u2__0remHi_451_0__398_; 
wire u2__0remHi_451_0__399_; 
wire u2__0remHi_451_0__39_; 
wire u2__0remHi_451_0__3_; 
wire u2__0remHi_451_0__400_; 
wire u2__0remHi_451_0__401_; 
wire u2__0remHi_451_0__402_; 
wire u2__0remHi_451_0__403_; 
wire u2__0remHi_451_0__404_; 
wire u2__0remHi_451_0__405_; 
wire u2__0remHi_451_0__406_; 
wire u2__0remHi_451_0__407_; 
wire u2__0remHi_451_0__408_; 
wire u2__0remHi_451_0__409_; 
wire u2__0remHi_451_0__40_; 
wire u2__0remHi_451_0__410_; 
wire u2__0remHi_451_0__411_; 
wire u2__0remHi_451_0__412_; 
wire u2__0remHi_451_0__413_; 
wire u2__0remHi_451_0__414_; 
wire u2__0remHi_451_0__415_; 
wire u2__0remHi_451_0__416_; 
wire u2__0remHi_451_0__417_; 
wire u2__0remHi_451_0__418_; 
wire u2__0remHi_451_0__419_; 
wire u2__0remHi_451_0__41_; 
wire u2__0remHi_451_0__420_; 
wire u2__0remHi_451_0__421_; 
wire u2__0remHi_451_0__422_; 
wire u2__0remHi_451_0__423_; 
wire u2__0remHi_451_0__424_; 
wire u2__0remHi_451_0__425_; 
wire u2__0remHi_451_0__426_; 
wire u2__0remHi_451_0__427_; 
wire u2__0remHi_451_0__428_; 
wire u2__0remHi_451_0__429_; 
wire u2__0remHi_451_0__42_; 
wire u2__0remHi_451_0__430_; 
wire u2__0remHi_451_0__431_; 
wire u2__0remHi_451_0__432_; 
wire u2__0remHi_451_0__433_; 
wire u2__0remHi_451_0__434_; 
wire u2__0remHi_451_0__435_; 
wire u2__0remHi_451_0__436_; 
wire u2__0remHi_451_0__437_; 
wire u2__0remHi_451_0__438_; 
wire u2__0remHi_451_0__439_; 
wire u2__0remHi_451_0__43_; 
wire u2__0remHi_451_0__440_; 
wire u2__0remHi_451_0__441_; 
wire u2__0remHi_451_0__442_; 
wire u2__0remHi_451_0__443_; 
wire u2__0remHi_451_0__444_; 
wire u2__0remHi_451_0__445_; 
wire u2__0remHi_451_0__446_; 
wire u2__0remHi_451_0__447_; 
wire u2__0remHi_451_0__448_; 
wire u2__0remHi_451_0__449_; 
wire u2__0remHi_451_0__44_; 
wire u2__0remHi_451_0__45_; 
wire u2__0remHi_451_0__46_; 
wire u2__0remHi_451_0__47_; 
wire u2__0remHi_451_0__48_; 
wire u2__0remHi_451_0__49_; 
wire u2__0remHi_451_0__4_; 
wire u2__0remHi_451_0__50_; 
wire u2__0remHi_451_0__51_; 
wire u2__0remHi_451_0__52_; 
wire u2__0remHi_451_0__53_; 
wire u2__0remHi_451_0__54_; 
wire u2__0remHi_451_0__55_; 
wire u2__0remHi_451_0__56_; 
wire u2__0remHi_451_0__57_; 
wire u2__0remHi_451_0__58_; 
wire u2__0remHi_451_0__59_; 
wire u2__0remHi_451_0__5_; 
wire u2__0remHi_451_0__60_; 
wire u2__0remHi_451_0__61_; 
wire u2__0remHi_451_0__62_; 
wire u2__0remHi_451_0__63_; 
wire u2__0remHi_451_0__64_; 
wire u2__0remHi_451_0__65_; 
wire u2__0remHi_451_0__66_; 
wire u2__0remHi_451_0__67_; 
wire u2__0remHi_451_0__68_; 
wire u2__0remHi_451_0__69_; 
wire u2__0remHi_451_0__6_; 
wire u2__0remHi_451_0__70_; 
wire u2__0remHi_451_0__71_; 
wire u2__0remHi_451_0__72_; 
wire u2__0remHi_451_0__73_; 
wire u2__0remHi_451_0__74_; 
wire u2__0remHi_451_0__75_; 
wire u2__0remHi_451_0__76_; 
wire u2__0remHi_451_0__77_; 
wire u2__0remHi_451_0__78_; 
wire u2__0remHi_451_0__79_; 
wire u2__0remHi_451_0__7_; 
wire u2__0remHi_451_0__80_; 
wire u2__0remHi_451_0__81_; 
wire u2__0remHi_451_0__82_; 
wire u2__0remHi_451_0__83_; 
wire u2__0remHi_451_0__84_; 
wire u2__0remHi_451_0__85_; 
wire u2__0remHi_451_0__86_; 
wire u2__0remHi_451_0__87_; 
wire u2__0remHi_451_0__88_; 
wire u2__0remHi_451_0__89_; 
wire u2__0remHi_451_0__8_; 
wire u2__0remHi_451_0__90_; 
wire u2__0remHi_451_0__91_; 
wire u2__0remHi_451_0__92_; 
wire u2__0remHi_451_0__93_; 
wire u2__0remHi_451_0__94_; 
wire u2__0remHi_451_0__95_; 
wire u2__0remHi_451_0__96_; 
wire u2__0remHi_451_0__97_; 
wire u2__0remHi_451_0__98_; 
wire u2__0remHi_451_0__99_; 
wire u2__0remHi_451_0__9_; 
wire u2__0remLo_451_0__0_; 
wire u2__0remLo_451_0__100_; 
wire u2__0remLo_451_0__101_; 
wire u2__0remLo_451_0__102_; 
wire u2__0remLo_451_0__103_; 
wire u2__0remLo_451_0__104_; 
wire u2__0remLo_451_0__105_; 
wire u2__0remLo_451_0__106_; 
wire u2__0remLo_451_0__107_; 
wire u2__0remLo_451_0__108_; 
wire u2__0remLo_451_0__109_; 
wire u2__0remLo_451_0__10_; 
wire u2__0remLo_451_0__110_; 
wire u2__0remLo_451_0__111_; 
wire u2__0remLo_451_0__112_; 
wire u2__0remLo_451_0__113_; 
wire u2__0remLo_451_0__114_; 
wire u2__0remLo_451_0__115_; 
wire u2__0remLo_451_0__116_; 
wire u2__0remLo_451_0__117_; 
wire u2__0remLo_451_0__118_; 
wire u2__0remLo_451_0__119_; 
wire u2__0remLo_451_0__11_; 
wire u2__0remLo_451_0__120_; 
wire u2__0remLo_451_0__121_; 
wire u2__0remLo_451_0__122_; 
wire u2__0remLo_451_0__123_; 
wire u2__0remLo_451_0__124_; 
wire u2__0remLo_451_0__125_; 
wire u2__0remLo_451_0__126_; 
wire u2__0remLo_451_0__127_; 
wire u2__0remLo_451_0__128_; 
wire u2__0remLo_451_0__129_; 
wire u2__0remLo_451_0__12_; 
wire u2__0remLo_451_0__130_; 
wire u2__0remLo_451_0__131_; 
wire u2__0remLo_451_0__132_; 
wire u2__0remLo_451_0__133_; 
wire u2__0remLo_451_0__134_; 
wire u2__0remLo_451_0__135_; 
wire u2__0remLo_451_0__136_; 
wire u2__0remLo_451_0__137_; 
wire u2__0remLo_451_0__138_; 
wire u2__0remLo_451_0__139_; 
wire u2__0remLo_451_0__13_; 
wire u2__0remLo_451_0__140_; 
wire u2__0remLo_451_0__141_; 
wire u2__0remLo_451_0__142_; 
wire u2__0remLo_451_0__143_; 
wire u2__0remLo_451_0__144_; 
wire u2__0remLo_451_0__145_; 
wire u2__0remLo_451_0__146_; 
wire u2__0remLo_451_0__147_; 
wire u2__0remLo_451_0__148_; 
wire u2__0remLo_451_0__149_; 
wire u2__0remLo_451_0__14_; 
wire u2__0remLo_451_0__150_; 
wire u2__0remLo_451_0__151_; 
wire u2__0remLo_451_0__152_; 
wire u2__0remLo_451_0__153_; 
wire u2__0remLo_451_0__154_; 
wire u2__0remLo_451_0__155_; 
wire u2__0remLo_451_0__156_; 
wire u2__0remLo_451_0__157_; 
wire u2__0remLo_451_0__158_; 
wire u2__0remLo_451_0__159_; 
wire u2__0remLo_451_0__15_; 
wire u2__0remLo_451_0__160_; 
wire u2__0remLo_451_0__161_; 
wire u2__0remLo_451_0__162_; 
wire u2__0remLo_451_0__163_; 
wire u2__0remLo_451_0__164_; 
wire u2__0remLo_451_0__165_; 
wire u2__0remLo_451_0__166_; 
wire u2__0remLo_451_0__167_; 
wire u2__0remLo_451_0__168_; 
wire u2__0remLo_451_0__169_; 
wire u2__0remLo_451_0__16_; 
wire u2__0remLo_451_0__170_; 
wire u2__0remLo_451_0__171_; 
wire u2__0remLo_451_0__172_; 
wire u2__0remLo_451_0__173_; 
wire u2__0remLo_451_0__174_; 
wire u2__0remLo_451_0__175_; 
wire u2__0remLo_451_0__176_; 
wire u2__0remLo_451_0__177_; 
wire u2__0remLo_451_0__178_; 
wire u2__0remLo_451_0__179_; 
wire u2__0remLo_451_0__17_; 
wire u2__0remLo_451_0__180_; 
wire u2__0remLo_451_0__181_; 
wire u2__0remLo_451_0__182_; 
wire u2__0remLo_451_0__183_; 
wire u2__0remLo_451_0__184_; 
wire u2__0remLo_451_0__185_; 
wire u2__0remLo_451_0__186_; 
wire u2__0remLo_451_0__187_; 
wire u2__0remLo_451_0__188_; 
wire u2__0remLo_451_0__189_; 
wire u2__0remLo_451_0__18_; 
wire u2__0remLo_451_0__190_; 
wire u2__0remLo_451_0__191_; 
wire u2__0remLo_451_0__192_; 
wire u2__0remLo_451_0__193_; 
wire u2__0remLo_451_0__194_; 
wire u2__0remLo_451_0__195_; 
wire u2__0remLo_451_0__196_; 
wire u2__0remLo_451_0__197_; 
wire u2__0remLo_451_0__198_; 
wire u2__0remLo_451_0__199_; 
wire u2__0remLo_451_0__19_; 
wire u2__0remLo_451_0__1_; 
wire u2__0remLo_451_0__200_; 
wire u2__0remLo_451_0__201_; 
wire u2__0remLo_451_0__202_; 
wire u2__0remLo_451_0__203_; 
wire u2__0remLo_451_0__204_; 
wire u2__0remLo_451_0__205_; 
wire u2__0remLo_451_0__206_; 
wire u2__0remLo_451_0__207_; 
wire u2__0remLo_451_0__208_; 
wire u2__0remLo_451_0__209_; 
wire u2__0remLo_451_0__20_; 
wire u2__0remLo_451_0__210_; 
wire u2__0remLo_451_0__211_; 
wire u2__0remLo_451_0__212_; 
wire u2__0remLo_451_0__213_; 
wire u2__0remLo_451_0__214_; 
wire u2__0remLo_451_0__215_; 
wire u2__0remLo_451_0__216_; 
wire u2__0remLo_451_0__217_; 
wire u2__0remLo_451_0__218_; 
wire u2__0remLo_451_0__219_; 
wire u2__0remLo_451_0__21_; 
wire u2__0remLo_451_0__220_; 
wire u2__0remLo_451_0__221_; 
wire u2__0remLo_451_0__222_; 
wire u2__0remLo_451_0__223_; 
wire u2__0remLo_451_0__224_; 
wire u2__0remLo_451_0__225_; 
wire u2__0remLo_451_0__226_; 
wire u2__0remLo_451_0__227_; 
wire u2__0remLo_451_0__228_; 
wire u2__0remLo_451_0__229_; 
wire u2__0remLo_451_0__22_; 
wire u2__0remLo_451_0__230_; 
wire u2__0remLo_451_0__231_; 
wire u2__0remLo_451_0__232_; 
wire u2__0remLo_451_0__233_; 
wire u2__0remLo_451_0__234_; 
wire u2__0remLo_451_0__235_; 
wire u2__0remLo_451_0__236_; 
wire u2__0remLo_451_0__237_; 
wire u2__0remLo_451_0__238_; 
wire u2__0remLo_451_0__239_; 
wire u2__0remLo_451_0__23_; 
wire u2__0remLo_451_0__240_; 
wire u2__0remLo_451_0__241_; 
wire u2__0remLo_451_0__242_; 
wire u2__0remLo_451_0__243_; 
wire u2__0remLo_451_0__244_; 
wire u2__0remLo_451_0__245_; 
wire u2__0remLo_451_0__246_; 
wire u2__0remLo_451_0__247_; 
wire u2__0remLo_451_0__248_; 
wire u2__0remLo_451_0__249_; 
wire u2__0remLo_451_0__24_; 
wire u2__0remLo_451_0__250_; 
wire u2__0remLo_451_0__251_; 
wire u2__0remLo_451_0__252_; 
wire u2__0remLo_451_0__253_; 
wire u2__0remLo_451_0__254_; 
wire u2__0remLo_451_0__255_; 
wire u2__0remLo_451_0__256_; 
wire u2__0remLo_451_0__257_; 
wire u2__0remLo_451_0__258_; 
wire u2__0remLo_451_0__259_; 
wire u2__0remLo_451_0__25_; 
wire u2__0remLo_451_0__260_; 
wire u2__0remLo_451_0__261_; 
wire u2__0remLo_451_0__262_; 
wire u2__0remLo_451_0__263_; 
wire u2__0remLo_451_0__264_; 
wire u2__0remLo_451_0__265_; 
wire u2__0remLo_451_0__266_; 
wire u2__0remLo_451_0__267_; 
wire u2__0remLo_451_0__268_; 
wire u2__0remLo_451_0__269_; 
wire u2__0remLo_451_0__26_; 
wire u2__0remLo_451_0__270_; 
wire u2__0remLo_451_0__271_; 
wire u2__0remLo_451_0__272_; 
wire u2__0remLo_451_0__273_; 
wire u2__0remLo_451_0__274_; 
wire u2__0remLo_451_0__275_; 
wire u2__0remLo_451_0__276_; 
wire u2__0remLo_451_0__277_; 
wire u2__0remLo_451_0__278_; 
wire u2__0remLo_451_0__279_; 
wire u2__0remLo_451_0__27_; 
wire u2__0remLo_451_0__280_; 
wire u2__0remLo_451_0__281_; 
wire u2__0remLo_451_0__282_; 
wire u2__0remLo_451_0__283_; 
wire u2__0remLo_451_0__284_; 
wire u2__0remLo_451_0__285_; 
wire u2__0remLo_451_0__286_; 
wire u2__0remLo_451_0__287_; 
wire u2__0remLo_451_0__288_; 
wire u2__0remLo_451_0__289_; 
wire u2__0remLo_451_0__28_; 
wire u2__0remLo_451_0__290_; 
wire u2__0remLo_451_0__291_; 
wire u2__0remLo_451_0__292_; 
wire u2__0remLo_451_0__293_; 
wire u2__0remLo_451_0__294_; 
wire u2__0remLo_451_0__295_; 
wire u2__0remLo_451_0__296_; 
wire u2__0remLo_451_0__297_; 
wire u2__0remLo_451_0__298_; 
wire u2__0remLo_451_0__299_; 
wire u2__0remLo_451_0__29_; 
wire u2__0remLo_451_0__2_; 
wire u2__0remLo_451_0__300_; 
wire u2__0remLo_451_0__301_; 
wire u2__0remLo_451_0__302_; 
wire u2__0remLo_451_0__303_; 
wire u2__0remLo_451_0__304_; 
wire u2__0remLo_451_0__305_; 
wire u2__0remLo_451_0__306_; 
wire u2__0remLo_451_0__307_; 
wire u2__0remLo_451_0__308_; 
wire u2__0remLo_451_0__309_; 
wire u2__0remLo_451_0__30_; 
wire u2__0remLo_451_0__310_; 
wire u2__0remLo_451_0__311_; 
wire u2__0remLo_451_0__312_; 
wire u2__0remLo_451_0__313_; 
wire u2__0remLo_451_0__314_; 
wire u2__0remLo_451_0__315_; 
wire u2__0remLo_451_0__316_; 
wire u2__0remLo_451_0__317_; 
wire u2__0remLo_451_0__318_; 
wire u2__0remLo_451_0__319_; 
wire u2__0remLo_451_0__31_; 
wire u2__0remLo_451_0__320_; 
wire u2__0remLo_451_0__321_; 
wire u2__0remLo_451_0__322_; 
wire u2__0remLo_451_0__323_; 
wire u2__0remLo_451_0__324_; 
wire u2__0remLo_451_0__325_; 
wire u2__0remLo_451_0__326_; 
wire u2__0remLo_451_0__327_; 
wire u2__0remLo_451_0__328_; 
wire u2__0remLo_451_0__329_; 
wire u2__0remLo_451_0__32_; 
wire u2__0remLo_451_0__330_; 
wire u2__0remLo_451_0__331_; 
wire u2__0remLo_451_0__332_; 
wire u2__0remLo_451_0__333_; 
wire u2__0remLo_451_0__334_; 
wire u2__0remLo_451_0__335_; 
wire u2__0remLo_451_0__336_; 
wire u2__0remLo_451_0__337_; 
wire u2__0remLo_451_0__338_; 
wire u2__0remLo_451_0__339_; 
wire u2__0remLo_451_0__33_; 
wire u2__0remLo_451_0__340_; 
wire u2__0remLo_451_0__341_; 
wire u2__0remLo_451_0__342_; 
wire u2__0remLo_451_0__343_; 
wire u2__0remLo_451_0__344_; 
wire u2__0remLo_451_0__345_; 
wire u2__0remLo_451_0__346_; 
wire u2__0remLo_451_0__347_; 
wire u2__0remLo_451_0__348_; 
wire u2__0remLo_451_0__349_; 
wire u2__0remLo_451_0__34_; 
wire u2__0remLo_451_0__350_; 
wire u2__0remLo_451_0__351_; 
wire u2__0remLo_451_0__352_; 
wire u2__0remLo_451_0__353_; 
wire u2__0remLo_451_0__354_; 
wire u2__0remLo_451_0__355_; 
wire u2__0remLo_451_0__356_; 
wire u2__0remLo_451_0__357_; 
wire u2__0remLo_451_0__358_; 
wire u2__0remLo_451_0__359_; 
wire u2__0remLo_451_0__35_; 
wire u2__0remLo_451_0__360_; 
wire u2__0remLo_451_0__361_; 
wire u2__0remLo_451_0__362_; 
wire u2__0remLo_451_0__363_; 
wire u2__0remLo_451_0__364_; 
wire u2__0remLo_451_0__365_; 
wire u2__0remLo_451_0__366_; 
wire u2__0remLo_451_0__367_; 
wire u2__0remLo_451_0__368_; 
wire u2__0remLo_451_0__369_; 
wire u2__0remLo_451_0__36_; 
wire u2__0remLo_451_0__370_; 
wire u2__0remLo_451_0__371_; 
wire u2__0remLo_451_0__372_; 
wire u2__0remLo_451_0__373_; 
wire u2__0remLo_451_0__374_; 
wire u2__0remLo_451_0__375_; 
wire u2__0remLo_451_0__376_; 
wire u2__0remLo_451_0__377_; 
wire u2__0remLo_451_0__378_; 
wire u2__0remLo_451_0__379_; 
wire u2__0remLo_451_0__37_; 
wire u2__0remLo_451_0__380_; 
wire u2__0remLo_451_0__381_; 
wire u2__0remLo_451_0__382_; 
wire u2__0remLo_451_0__383_; 
wire u2__0remLo_451_0__384_; 
wire u2__0remLo_451_0__385_; 
wire u2__0remLo_451_0__386_; 
wire u2__0remLo_451_0__387_; 
wire u2__0remLo_451_0__388_; 
wire u2__0remLo_451_0__389_; 
wire u2__0remLo_451_0__38_; 
wire u2__0remLo_451_0__390_; 
wire u2__0remLo_451_0__391_; 
wire u2__0remLo_451_0__392_; 
wire u2__0remLo_451_0__393_; 
wire u2__0remLo_451_0__394_; 
wire u2__0remLo_451_0__395_; 
wire u2__0remLo_451_0__396_; 
wire u2__0remLo_451_0__397_; 
wire u2__0remLo_451_0__398_; 
wire u2__0remLo_451_0__399_; 
wire u2__0remLo_451_0__39_; 
wire u2__0remLo_451_0__3_; 
wire u2__0remLo_451_0__400_; 
wire u2__0remLo_451_0__401_; 
wire u2__0remLo_451_0__402_; 
wire u2__0remLo_451_0__403_; 
wire u2__0remLo_451_0__404_; 
wire u2__0remLo_451_0__405_; 
wire u2__0remLo_451_0__406_; 
wire u2__0remLo_451_0__407_; 
wire u2__0remLo_451_0__408_; 
wire u2__0remLo_451_0__409_; 
wire u2__0remLo_451_0__40_; 
wire u2__0remLo_451_0__410_; 
wire u2__0remLo_451_0__411_; 
wire u2__0remLo_451_0__412_; 
wire u2__0remLo_451_0__413_; 
wire u2__0remLo_451_0__414_; 
wire u2__0remLo_451_0__415_; 
wire u2__0remLo_451_0__416_; 
wire u2__0remLo_451_0__417_; 
wire u2__0remLo_451_0__418_; 
wire u2__0remLo_451_0__419_; 
wire u2__0remLo_451_0__41_; 
wire u2__0remLo_451_0__420_; 
wire u2__0remLo_451_0__421_; 
wire u2__0remLo_451_0__422_; 
wire u2__0remLo_451_0__423_; 
wire u2__0remLo_451_0__424_; 
wire u2__0remLo_451_0__425_; 
wire u2__0remLo_451_0__426_; 
wire u2__0remLo_451_0__427_; 
wire u2__0remLo_451_0__428_; 
wire u2__0remLo_451_0__429_; 
wire u2__0remLo_451_0__42_; 
wire u2__0remLo_451_0__430_; 
wire u2__0remLo_451_0__431_; 
wire u2__0remLo_451_0__432_; 
wire u2__0remLo_451_0__433_; 
wire u2__0remLo_451_0__434_; 
wire u2__0remLo_451_0__435_; 
wire u2__0remLo_451_0__436_; 
wire u2__0remLo_451_0__437_; 
wire u2__0remLo_451_0__438_; 
wire u2__0remLo_451_0__439_; 
wire u2__0remLo_451_0__43_; 
wire u2__0remLo_451_0__440_; 
wire u2__0remLo_451_0__441_; 
wire u2__0remLo_451_0__442_; 
wire u2__0remLo_451_0__443_; 
wire u2__0remLo_451_0__444_; 
wire u2__0remLo_451_0__445_; 
wire u2__0remLo_451_0__446_; 
wire u2__0remLo_451_0__447_; 
wire u2__0remLo_451_0__448_; 
wire u2__0remLo_451_0__449_; 
wire u2__0remLo_451_0__44_; 
wire u2__0remLo_451_0__450_; 
wire u2__0remLo_451_0__451_; 
wire u2__0remLo_451_0__45_; 
wire u2__0remLo_451_0__46_; 
wire u2__0remLo_451_0__47_; 
wire u2__0remLo_451_0__48_; 
wire u2__0remLo_451_0__49_; 
wire u2__0remLo_451_0__4_; 
wire u2__0remLo_451_0__50_; 
wire u2__0remLo_451_0__51_; 
wire u2__0remLo_451_0__52_; 
wire u2__0remLo_451_0__53_; 
wire u2__0remLo_451_0__54_; 
wire u2__0remLo_451_0__55_; 
wire u2__0remLo_451_0__56_; 
wire u2__0remLo_451_0__57_; 
wire u2__0remLo_451_0__58_; 
wire u2__0remLo_451_0__59_; 
wire u2__0remLo_451_0__5_; 
wire u2__0remLo_451_0__60_; 
wire u2__0remLo_451_0__61_; 
wire u2__0remLo_451_0__62_; 
wire u2__0remLo_451_0__63_; 
wire u2__0remLo_451_0__64_; 
wire u2__0remLo_451_0__65_; 
wire u2__0remLo_451_0__66_; 
wire u2__0remLo_451_0__67_; 
wire u2__0remLo_451_0__68_; 
wire u2__0remLo_451_0__69_; 
wire u2__0remLo_451_0__6_; 
wire u2__0remLo_451_0__70_; 
wire u2__0remLo_451_0__71_; 
wire u2__0remLo_451_0__72_; 
wire u2__0remLo_451_0__73_; 
wire u2__0remLo_451_0__74_; 
wire u2__0remLo_451_0__75_; 
wire u2__0remLo_451_0__76_; 
wire u2__0remLo_451_0__77_; 
wire u2__0remLo_451_0__78_; 
wire u2__0remLo_451_0__79_; 
wire u2__0remLo_451_0__7_; 
wire u2__0remLo_451_0__80_; 
wire u2__0remLo_451_0__81_; 
wire u2__0remLo_451_0__82_; 
wire u2__0remLo_451_0__83_; 
wire u2__0remLo_451_0__84_; 
wire u2__0remLo_451_0__85_; 
wire u2__0remLo_451_0__86_; 
wire u2__0remLo_451_0__87_; 
wire u2__0remLo_451_0__88_; 
wire u2__0remLo_451_0__89_; 
wire u2__0remLo_451_0__8_; 
wire u2__0remLo_451_0__90_; 
wire u2__0remLo_451_0__91_; 
wire u2__0remLo_451_0__92_; 
wire u2__0remLo_451_0__93_; 
wire u2__0remLo_451_0__94_; 
wire u2__0remLo_451_0__95_; 
wire u2__0remLo_451_0__96_; 
wire u2__0remLo_451_0__97_; 
wire u2__0remLo_451_0__98_; 
wire u2__0remLo_451_0__99_; 
wire u2__0remLo_451_0__9_; 
wire u2__0root_452_0__0_; 
wire u2__0root_452_0__100_; 
wire u2__0root_452_0__101_; 
wire u2__0root_452_0__102_; 
wire u2__0root_452_0__103_; 
wire u2__0root_452_0__104_; 
wire u2__0root_452_0__105_; 
wire u2__0root_452_0__106_; 
wire u2__0root_452_0__107_; 
wire u2__0root_452_0__108_; 
wire u2__0root_452_0__109_; 
wire u2__0root_452_0__10_; 
wire u2__0root_452_0__110_; 
wire u2__0root_452_0__111_; 
wire u2__0root_452_0__112_; 
wire u2__0root_452_0__113_; 
wire u2__0root_452_0__114_; 
wire u2__0root_452_0__115_; 
wire u2__0root_452_0__116_; 
wire u2__0root_452_0__117_; 
wire u2__0root_452_0__118_; 
wire u2__0root_452_0__119_; 
wire u2__0root_452_0__11_; 
wire u2__0root_452_0__120_; 
wire u2__0root_452_0__121_; 
wire u2__0root_452_0__122_; 
wire u2__0root_452_0__123_; 
wire u2__0root_452_0__124_; 
wire u2__0root_452_0__125_; 
wire u2__0root_452_0__126_; 
wire u2__0root_452_0__127_; 
wire u2__0root_452_0__128_; 
wire u2__0root_452_0__129_; 
wire u2__0root_452_0__12_; 
wire u2__0root_452_0__130_; 
wire u2__0root_452_0__131_; 
wire u2__0root_452_0__132_; 
wire u2__0root_452_0__133_; 
wire u2__0root_452_0__134_; 
wire u2__0root_452_0__135_; 
wire u2__0root_452_0__136_; 
wire u2__0root_452_0__137_; 
wire u2__0root_452_0__138_; 
wire u2__0root_452_0__139_; 
wire u2__0root_452_0__13_; 
wire u2__0root_452_0__140_; 
wire u2__0root_452_0__141_; 
wire u2__0root_452_0__142_; 
wire u2__0root_452_0__143_; 
wire u2__0root_452_0__144_; 
wire u2__0root_452_0__145_; 
wire u2__0root_452_0__146_; 
wire u2__0root_452_0__147_; 
wire u2__0root_452_0__148_; 
wire u2__0root_452_0__149_; 
wire u2__0root_452_0__14_; 
wire u2__0root_452_0__150_; 
wire u2__0root_452_0__151_; 
wire u2__0root_452_0__152_; 
wire u2__0root_452_0__153_; 
wire u2__0root_452_0__154_; 
wire u2__0root_452_0__155_; 
wire u2__0root_452_0__156_; 
wire u2__0root_452_0__157_; 
wire u2__0root_452_0__158_; 
wire u2__0root_452_0__159_; 
wire u2__0root_452_0__15_; 
wire u2__0root_452_0__160_; 
wire u2__0root_452_0__161_; 
wire u2__0root_452_0__162_; 
wire u2__0root_452_0__163_; 
wire u2__0root_452_0__164_; 
wire u2__0root_452_0__165_; 
wire u2__0root_452_0__166_; 
wire u2__0root_452_0__167_; 
wire u2__0root_452_0__168_; 
wire u2__0root_452_0__169_; 
wire u2__0root_452_0__16_; 
wire u2__0root_452_0__170_; 
wire u2__0root_452_0__171_; 
wire u2__0root_452_0__172_; 
wire u2__0root_452_0__173_; 
wire u2__0root_452_0__174_; 
wire u2__0root_452_0__175_; 
wire u2__0root_452_0__176_; 
wire u2__0root_452_0__177_; 
wire u2__0root_452_0__178_; 
wire u2__0root_452_0__179_; 
wire u2__0root_452_0__17_; 
wire u2__0root_452_0__180_; 
wire u2__0root_452_0__181_; 
wire u2__0root_452_0__182_; 
wire u2__0root_452_0__183_; 
wire u2__0root_452_0__184_; 
wire u2__0root_452_0__185_; 
wire u2__0root_452_0__186_; 
wire u2__0root_452_0__187_; 
wire u2__0root_452_0__188_; 
wire u2__0root_452_0__189_; 
wire u2__0root_452_0__18_; 
wire u2__0root_452_0__190_; 
wire u2__0root_452_0__191_; 
wire u2__0root_452_0__192_; 
wire u2__0root_452_0__193_; 
wire u2__0root_452_0__194_; 
wire u2__0root_452_0__195_; 
wire u2__0root_452_0__196_; 
wire u2__0root_452_0__197_; 
wire u2__0root_452_0__198_; 
wire u2__0root_452_0__199_; 
wire u2__0root_452_0__19_; 
wire u2__0root_452_0__1_; 
wire u2__0root_452_0__200_; 
wire u2__0root_452_0__201_; 
wire u2__0root_452_0__202_; 
wire u2__0root_452_0__203_; 
wire u2__0root_452_0__204_; 
wire u2__0root_452_0__205_; 
wire u2__0root_452_0__206_; 
wire u2__0root_452_0__207_; 
wire u2__0root_452_0__208_; 
wire u2__0root_452_0__209_; 
wire u2__0root_452_0__20_; 
wire u2__0root_452_0__210_; 
wire u2__0root_452_0__211_; 
wire u2__0root_452_0__212_; 
wire u2__0root_452_0__213_; 
wire u2__0root_452_0__214_; 
wire u2__0root_452_0__215_; 
wire u2__0root_452_0__216_; 
wire u2__0root_452_0__217_; 
wire u2__0root_452_0__218_; 
wire u2__0root_452_0__219_; 
wire u2__0root_452_0__21_; 
wire u2__0root_452_0__220_; 
wire u2__0root_452_0__221_; 
wire u2__0root_452_0__222_; 
wire u2__0root_452_0__223_; 
wire u2__0root_452_0__224_; 
wire u2__0root_452_0__225_; 
wire u2__0root_452_0__226_; 
wire u2__0root_452_0__227_; 
wire u2__0root_452_0__228_; 
wire u2__0root_452_0__229_; 
wire u2__0root_452_0__22_; 
wire u2__0root_452_0__230_; 
wire u2__0root_452_0__231_; 
wire u2__0root_452_0__232_; 
wire u2__0root_452_0__233_; 
wire u2__0root_452_0__234_; 
wire u2__0root_452_0__235_; 
wire u2__0root_452_0__236_; 
wire u2__0root_452_0__237_; 
wire u2__0root_452_0__238_; 
wire u2__0root_452_0__239_; 
wire u2__0root_452_0__23_; 
wire u2__0root_452_0__240_; 
wire u2__0root_452_0__241_; 
wire u2__0root_452_0__242_; 
wire u2__0root_452_0__243_; 
wire u2__0root_452_0__244_; 
wire u2__0root_452_0__245_; 
wire u2__0root_452_0__246_; 
wire u2__0root_452_0__247_; 
wire u2__0root_452_0__248_; 
wire u2__0root_452_0__249_; 
wire u2__0root_452_0__24_; 
wire u2__0root_452_0__250_; 
wire u2__0root_452_0__251_; 
wire u2__0root_452_0__252_; 
wire u2__0root_452_0__253_; 
wire u2__0root_452_0__254_; 
wire u2__0root_452_0__255_; 
wire u2__0root_452_0__256_; 
wire u2__0root_452_0__257_; 
wire u2__0root_452_0__258_; 
wire u2__0root_452_0__259_; 
wire u2__0root_452_0__25_; 
wire u2__0root_452_0__260_; 
wire u2__0root_452_0__261_; 
wire u2__0root_452_0__262_; 
wire u2__0root_452_0__263_; 
wire u2__0root_452_0__264_; 
wire u2__0root_452_0__265_; 
wire u2__0root_452_0__266_; 
wire u2__0root_452_0__267_; 
wire u2__0root_452_0__268_; 
wire u2__0root_452_0__269_; 
wire u2__0root_452_0__26_; 
wire u2__0root_452_0__270_; 
wire u2__0root_452_0__271_; 
wire u2__0root_452_0__272_; 
wire u2__0root_452_0__273_; 
wire u2__0root_452_0__274_; 
wire u2__0root_452_0__275_; 
wire u2__0root_452_0__276_; 
wire u2__0root_452_0__277_; 
wire u2__0root_452_0__278_; 
wire u2__0root_452_0__279_; 
wire u2__0root_452_0__27_; 
wire u2__0root_452_0__280_; 
wire u2__0root_452_0__281_; 
wire u2__0root_452_0__282_; 
wire u2__0root_452_0__283_; 
wire u2__0root_452_0__284_; 
wire u2__0root_452_0__285_; 
wire u2__0root_452_0__286_; 
wire u2__0root_452_0__287_; 
wire u2__0root_452_0__288_; 
wire u2__0root_452_0__289_; 
wire u2__0root_452_0__28_; 
wire u2__0root_452_0__290_; 
wire u2__0root_452_0__291_; 
wire u2__0root_452_0__292_; 
wire u2__0root_452_0__293_; 
wire u2__0root_452_0__294_; 
wire u2__0root_452_0__295_; 
wire u2__0root_452_0__296_; 
wire u2__0root_452_0__297_; 
wire u2__0root_452_0__298_; 
wire u2__0root_452_0__299_; 
wire u2__0root_452_0__29_; 
wire u2__0root_452_0__2_; 
wire u2__0root_452_0__300_; 
wire u2__0root_452_0__301_; 
wire u2__0root_452_0__302_; 
wire u2__0root_452_0__303_; 
wire u2__0root_452_0__304_; 
wire u2__0root_452_0__305_; 
wire u2__0root_452_0__306_; 
wire u2__0root_452_0__307_; 
wire u2__0root_452_0__308_; 
wire u2__0root_452_0__309_; 
wire u2__0root_452_0__30_; 
wire u2__0root_452_0__310_; 
wire u2__0root_452_0__311_; 
wire u2__0root_452_0__312_; 
wire u2__0root_452_0__313_; 
wire u2__0root_452_0__314_; 
wire u2__0root_452_0__315_; 
wire u2__0root_452_0__316_; 
wire u2__0root_452_0__317_; 
wire u2__0root_452_0__318_; 
wire u2__0root_452_0__319_; 
wire u2__0root_452_0__31_; 
wire u2__0root_452_0__320_; 
wire u2__0root_452_0__321_; 
wire u2__0root_452_0__322_; 
wire u2__0root_452_0__323_; 
wire u2__0root_452_0__324_; 
wire u2__0root_452_0__325_; 
wire u2__0root_452_0__326_; 
wire u2__0root_452_0__327_; 
wire u2__0root_452_0__328_; 
wire u2__0root_452_0__329_; 
wire u2__0root_452_0__32_; 
wire u2__0root_452_0__330_; 
wire u2__0root_452_0__331_; 
wire u2__0root_452_0__332_; 
wire u2__0root_452_0__333_; 
wire u2__0root_452_0__334_; 
wire u2__0root_452_0__335_; 
wire u2__0root_452_0__336_; 
wire u2__0root_452_0__337_; 
wire u2__0root_452_0__338_; 
wire u2__0root_452_0__339_; 
wire u2__0root_452_0__33_; 
wire u2__0root_452_0__340_; 
wire u2__0root_452_0__341_; 
wire u2__0root_452_0__342_; 
wire u2__0root_452_0__343_; 
wire u2__0root_452_0__344_; 
wire u2__0root_452_0__345_; 
wire u2__0root_452_0__346_; 
wire u2__0root_452_0__347_; 
wire u2__0root_452_0__348_; 
wire u2__0root_452_0__349_; 
wire u2__0root_452_0__34_; 
wire u2__0root_452_0__350_; 
wire u2__0root_452_0__351_; 
wire u2__0root_452_0__352_; 
wire u2__0root_452_0__353_; 
wire u2__0root_452_0__354_; 
wire u2__0root_452_0__355_; 
wire u2__0root_452_0__356_; 
wire u2__0root_452_0__357_; 
wire u2__0root_452_0__358_; 
wire u2__0root_452_0__359_; 
wire u2__0root_452_0__35_; 
wire u2__0root_452_0__360_; 
wire u2__0root_452_0__361_; 
wire u2__0root_452_0__362_; 
wire u2__0root_452_0__363_; 
wire u2__0root_452_0__364_; 
wire u2__0root_452_0__365_; 
wire u2__0root_452_0__366_; 
wire u2__0root_452_0__367_; 
wire u2__0root_452_0__368_; 
wire u2__0root_452_0__369_; 
wire u2__0root_452_0__36_; 
wire u2__0root_452_0__370_; 
wire u2__0root_452_0__371_; 
wire u2__0root_452_0__372_; 
wire u2__0root_452_0__373_; 
wire u2__0root_452_0__374_; 
wire u2__0root_452_0__375_; 
wire u2__0root_452_0__376_; 
wire u2__0root_452_0__377_; 
wire u2__0root_452_0__378_; 
wire u2__0root_452_0__379_; 
wire u2__0root_452_0__37_; 
wire u2__0root_452_0__380_; 
wire u2__0root_452_0__381_; 
wire u2__0root_452_0__382_; 
wire u2__0root_452_0__383_; 
wire u2__0root_452_0__384_; 
wire u2__0root_452_0__385_; 
wire u2__0root_452_0__386_; 
wire u2__0root_452_0__387_; 
wire u2__0root_452_0__388_; 
wire u2__0root_452_0__389_; 
wire u2__0root_452_0__38_; 
wire u2__0root_452_0__390_; 
wire u2__0root_452_0__391_; 
wire u2__0root_452_0__392_; 
wire u2__0root_452_0__393_; 
wire u2__0root_452_0__394_; 
wire u2__0root_452_0__395_; 
wire u2__0root_452_0__396_; 
wire u2__0root_452_0__397_; 
wire u2__0root_452_0__398_; 
wire u2__0root_452_0__399_; 
wire u2__0root_452_0__39_; 
wire u2__0root_452_0__3_; 
wire u2__0root_452_0__400_; 
wire u2__0root_452_0__401_; 
wire u2__0root_452_0__402_; 
wire u2__0root_452_0__403_; 
wire u2__0root_452_0__404_; 
wire u2__0root_452_0__405_; 
wire u2__0root_452_0__406_; 
wire u2__0root_452_0__407_; 
wire u2__0root_452_0__408_; 
wire u2__0root_452_0__409_; 
wire u2__0root_452_0__40_; 
wire u2__0root_452_0__410_; 
wire u2__0root_452_0__411_; 
wire u2__0root_452_0__412_; 
wire u2__0root_452_0__413_; 
wire u2__0root_452_0__414_; 
wire u2__0root_452_0__415_; 
wire u2__0root_452_0__416_; 
wire u2__0root_452_0__417_; 
wire u2__0root_452_0__418_; 
wire u2__0root_452_0__419_; 
wire u2__0root_452_0__41_; 
wire u2__0root_452_0__420_; 
wire u2__0root_452_0__421_; 
wire u2__0root_452_0__422_; 
wire u2__0root_452_0__423_; 
wire u2__0root_452_0__424_; 
wire u2__0root_452_0__425_; 
wire u2__0root_452_0__426_; 
wire u2__0root_452_0__427_; 
wire u2__0root_452_0__428_; 
wire u2__0root_452_0__429_; 
wire u2__0root_452_0__42_; 
wire u2__0root_452_0__430_; 
wire u2__0root_452_0__431_; 
wire u2__0root_452_0__432_; 
wire u2__0root_452_0__433_; 
wire u2__0root_452_0__434_; 
wire u2__0root_452_0__435_; 
wire u2__0root_452_0__436_; 
wire u2__0root_452_0__437_; 
wire u2__0root_452_0__438_; 
wire u2__0root_452_0__439_; 
wire u2__0root_452_0__43_; 
wire u2__0root_452_0__440_; 
wire u2__0root_452_0__441_; 
wire u2__0root_452_0__442_; 
wire u2__0root_452_0__443_; 
wire u2__0root_452_0__444_; 
wire u2__0root_452_0__445_; 
wire u2__0root_452_0__446_; 
wire u2__0root_452_0__447_; 
wire u2__0root_452_0__448_; 
wire u2__0root_452_0__449_; 
wire u2__0root_452_0__44_; 
wire u2__0root_452_0__450_; 
wire u2__0root_452_0__45_; 
wire u2__0root_452_0__46_; 
wire u2__0root_452_0__47_; 
wire u2__0root_452_0__48_; 
wire u2__0root_452_0__49_; 
wire u2__0root_452_0__4_; 
wire u2__0root_452_0__50_; 
wire u2__0root_452_0__51_; 
wire u2__0root_452_0__52_; 
wire u2__0root_452_0__53_; 
wire u2__0root_452_0__54_; 
wire u2__0root_452_0__55_; 
wire u2__0root_452_0__56_; 
wire u2__0root_452_0__57_; 
wire u2__0root_452_0__58_; 
wire u2__0root_452_0__59_; 
wire u2__0root_452_0__5_; 
wire u2__0root_452_0__60_; 
wire u2__0root_452_0__61_; 
wire u2__0root_452_0__62_; 
wire u2__0root_452_0__63_; 
wire u2__0root_452_0__64_; 
wire u2__0root_452_0__65_; 
wire u2__0root_452_0__66_; 
wire u2__0root_452_0__67_; 
wire u2__0root_452_0__68_; 
wire u2__0root_452_0__69_; 
wire u2__0root_452_0__6_; 
wire u2__0root_452_0__70_; 
wire u2__0root_452_0__71_; 
wire u2__0root_452_0__72_; 
wire u2__0root_452_0__73_; 
wire u2__0root_452_0__74_; 
wire u2__0root_452_0__75_; 
wire u2__0root_452_0__76_; 
wire u2__0root_452_0__77_; 
wire u2__0root_452_0__78_; 
wire u2__0root_452_0__79_; 
wire u2__0root_452_0__7_; 
wire u2__0root_452_0__80_; 
wire u2__0root_452_0__81_; 
wire u2__0root_452_0__82_; 
wire u2__0root_452_0__83_; 
wire u2__0root_452_0__84_; 
wire u2__0root_452_0__85_; 
wire u2__0root_452_0__86_; 
wire u2__0root_452_0__87_; 
wire u2__0root_452_0__88_; 
wire u2__0root_452_0__89_; 
wire u2__0root_452_0__8_; 
wire u2__0root_452_0__90_; 
wire u2__0root_452_0__91_; 
wire u2__0root_452_0__92_; 
wire u2__0root_452_0__93_; 
wire u2__0root_452_0__94_; 
wire u2__0root_452_0__95_; 
wire u2__0root_452_0__96_; 
wire u2__0root_452_0__97_; 
wire u2__0root_452_0__98_; 
wire u2__0root_452_0__99_; 
wire u2__0root_452_0__9_; 
wire u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_0_; 
wire u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_1_; 
wire u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_2_; 
wire u2__abc_52155_new_n10000_; 
wire u2__abc_52155_new_n10001_; 
wire u2__abc_52155_new_n10002_; 
wire u2__abc_52155_new_n10003_; 
wire u2__abc_52155_new_n10004_; 
wire u2__abc_52155_new_n10005_; 
wire u2__abc_52155_new_n10006_; 
wire u2__abc_52155_new_n10007_; 
wire u2__abc_52155_new_n10008_; 
wire u2__abc_52155_new_n10009_; 
wire u2__abc_52155_new_n10010_; 
wire u2__abc_52155_new_n10011_; 
wire u2__abc_52155_new_n10012_; 
wire u2__abc_52155_new_n10013_; 
wire u2__abc_52155_new_n10015_; 
wire u2__abc_52155_new_n10016_; 
wire u2__abc_52155_new_n10017_; 
wire u2__abc_52155_new_n10018_; 
wire u2__abc_52155_new_n10019_; 
wire u2__abc_52155_new_n10020_; 
wire u2__abc_52155_new_n10021_; 
wire u2__abc_52155_new_n10022_; 
wire u2__abc_52155_new_n10023_; 
wire u2__abc_52155_new_n10024_; 
wire u2__abc_52155_new_n10025_; 
wire u2__abc_52155_new_n10026_; 
wire u2__abc_52155_new_n10027_; 
wire u2__abc_52155_new_n10028_; 
wire u2__abc_52155_new_n10029_; 
wire u2__abc_52155_new_n10030_; 
wire u2__abc_52155_new_n10031_; 
wire u2__abc_52155_new_n10032_; 
wire u2__abc_52155_new_n10033_; 
wire u2__abc_52155_new_n10035_; 
wire u2__abc_52155_new_n10036_; 
wire u2__abc_52155_new_n10037_; 
wire u2__abc_52155_new_n10038_; 
wire u2__abc_52155_new_n10039_; 
wire u2__abc_52155_new_n10040_; 
wire u2__abc_52155_new_n10041_; 
wire u2__abc_52155_new_n10042_; 
wire u2__abc_52155_new_n10043_; 
wire u2__abc_52155_new_n10044_; 
wire u2__abc_52155_new_n10045_; 
wire u2__abc_52155_new_n10046_; 
wire u2__abc_52155_new_n10047_; 
wire u2__abc_52155_new_n10048_; 
wire u2__abc_52155_new_n10049_; 
wire u2__abc_52155_new_n10050_; 
wire u2__abc_52155_new_n10052_; 
wire u2__abc_52155_new_n10053_; 
wire u2__abc_52155_new_n10054_; 
wire u2__abc_52155_new_n10055_; 
wire u2__abc_52155_new_n10056_; 
wire u2__abc_52155_new_n10057_; 
wire u2__abc_52155_new_n10058_; 
wire u2__abc_52155_new_n10059_; 
wire u2__abc_52155_new_n10060_; 
wire u2__abc_52155_new_n10061_; 
wire u2__abc_52155_new_n10062_; 
wire u2__abc_52155_new_n10063_; 
wire u2__abc_52155_new_n10064_; 
wire u2__abc_52155_new_n10065_; 
wire u2__abc_52155_new_n10066_; 
wire u2__abc_52155_new_n10067_; 
wire u2__abc_52155_new_n10068_; 
wire u2__abc_52155_new_n10069_; 
wire u2__abc_52155_new_n10070_; 
wire u2__abc_52155_new_n10071_; 
wire u2__abc_52155_new_n10073_; 
wire u2__abc_52155_new_n10074_; 
wire u2__abc_52155_new_n10075_; 
wire u2__abc_52155_new_n10076_; 
wire u2__abc_52155_new_n10077_; 
wire u2__abc_52155_new_n10078_; 
wire u2__abc_52155_new_n10079_; 
wire u2__abc_52155_new_n10080_; 
wire u2__abc_52155_new_n10081_; 
wire u2__abc_52155_new_n10082_; 
wire u2__abc_52155_new_n10083_; 
wire u2__abc_52155_new_n10084_; 
wire u2__abc_52155_new_n10085_; 
wire u2__abc_52155_new_n10086_; 
wire u2__abc_52155_new_n10087_; 
wire u2__abc_52155_new_n10088_; 
wire u2__abc_52155_new_n10090_; 
wire u2__abc_52155_new_n10091_; 
wire u2__abc_52155_new_n10092_; 
wire u2__abc_52155_new_n10093_; 
wire u2__abc_52155_new_n10094_; 
wire u2__abc_52155_new_n10095_; 
wire u2__abc_52155_new_n10096_; 
wire u2__abc_52155_new_n10097_; 
wire u2__abc_52155_new_n10098_; 
wire u2__abc_52155_new_n10099_; 
wire u2__abc_52155_new_n10100_; 
wire u2__abc_52155_new_n10101_; 
wire u2__abc_52155_new_n10102_; 
wire u2__abc_52155_new_n10103_; 
wire u2__abc_52155_new_n10104_; 
wire u2__abc_52155_new_n10105_; 
wire u2__abc_52155_new_n10106_; 
wire u2__abc_52155_new_n10107_; 
wire u2__abc_52155_new_n10108_; 
wire u2__abc_52155_new_n10110_; 
wire u2__abc_52155_new_n10111_; 
wire u2__abc_52155_new_n10112_; 
wire u2__abc_52155_new_n10113_; 
wire u2__abc_52155_new_n10114_; 
wire u2__abc_52155_new_n10115_; 
wire u2__abc_52155_new_n10116_; 
wire u2__abc_52155_new_n10117_; 
wire u2__abc_52155_new_n10118_; 
wire u2__abc_52155_new_n10119_; 
wire u2__abc_52155_new_n10120_; 
wire u2__abc_52155_new_n10121_; 
wire u2__abc_52155_new_n10122_; 
wire u2__abc_52155_new_n10123_; 
wire u2__abc_52155_new_n10124_; 
wire u2__abc_52155_new_n10125_; 
wire u2__abc_52155_new_n10127_; 
wire u2__abc_52155_new_n10128_; 
wire u2__abc_52155_new_n10129_; 
wire u2__abc_52155_new_n10130_; 
wire u2__abc_52155_new_n10131_; 
wire u2__abc_52155_new_n10132_; 
wire u2__abc_52155_new_n10133_; 
wire u2__abc_52155_new_n10134_; 
wire u2__abc_52155_new_n10135_; 
wire u2__abc_52155_new_n10136_; 
wire u2__abc_52155_new_n10137_; 
wire u2__abc_52155_new_n10138_; 
wire u2__abc_52155_new_n10139_; 
wire u2__abc_52155_new_n10140_; 
wire u2__abc_52155_new_n10141_; 
wire u2__abc_52155_new_n10142_; 
wire u2__abc_52155_new_n10143_; 
wire u2__abc_52155_new_n10144_; 
wire u2__abc_52155_new_n10145_; 
wire u2__abc_52155_new_n10146_; 
wire u2__abc_52155_new_n10147_; 
wire u2__abc_52155_new_n10148_; 
wire u2__abc_52155_new_n10149_; 
wire u2__abc_52155_new_n10150_; 
wire u2__abc_52155_new_n10151_; 
wire u2__abc_52155_new_n10152_; 
wire u2__abc_52155_new_n10153_; 
wire u2__abc_52155_new_n10154_; 
wire u2__abc_52155_new_n10155_; 
wire u2__abc_52155_new_n10156_; 
wire u2__abc_52155_new_n10157_; 
wire u2__abc_52155_new_n10158_; 
wire u2__abc_52155_new_n10159_; 
wire u2__abc_52155_new_n10160_; 
wire u2__abc_52155_new_n10161_; 
wire u2__abc_52155_new_n10162_; 
wire u2__abc_52155_new_n10163_; 
wire u2__abc_52155_new_n10165_; 
wire u2__abc_52155_new_n10166_; 
wire u2__abc_52155_new_n10167_; 
wire u2__abc_52155_new_n10168_; 
wire u2__abc_52155_new_n10169_; 
wire u2__abc_52155_new_n10170_; 
wire u2__abc_52155_new_n10171_; 
wire u2__abc_52155_new_n10172_; 
wire u2__abc_52155_new_n10173_; 
wire u2__abc_52155_new_n10174_; 
wire u2__abc_52155_new_n10175_; 
wire u2__abc_52155_new_n10176_; 
wire u2__abc_52155_new_n10177_; 
wire u2__abc_52155_new_n10178_; 
wire u2__abc_52155_new_n10179_; 
wire u2__abc_52155_new_n10180_; 
wire u2__abc_52155_new_n10182_; 
wire u2__abc_52155_new_n10183_; 
wire u2__abc_52155_new_n10184_; 
wire u2__abc_52155_new_n10185_; 
wire u2__abc_52155_new_n10186_; 
wire u2__abc_52155_new_n10187_; 
wire u2__abc_52155_new_n10188_; 
wire u2__abc_52155_new_n10189_; 
wire u2__abc_52155_new_n10190_; 
wire u2__abc_52155_new_n10191_; 
wire u2__abc_52155_new_n10192_; 
wire u2__abc_52155_new_n10193_; 
wire u2__abc_52155_new_n10194_; 
wire u2__abc_52155_new_n10195_; 
wire u2__abc_52155_new_n10196_; 
wire u2__abc_52155_new_n10197_; 
wire u2__abc_52155_new_n10198_; 
wire u2__abc_52155_new_n10199_; 
wire u2__abc_52155_new_n10200_; 
wire u2__abc_52155_new_n10201_; 
wire u2__abc_52155_new_n10203_; 
wire u2__abc_52155_new_n10204_; 
wire u2__abc_52155_new_n10205_; 
wire u2__abc_52155_new_n10206_; 
wire u2__abc_52155_new_n10207_; 
wire u2__abc_52155_new_n10208_; 
wire u2__abc_52155_new_n10209_; 
wire u2__abc_52155_new_n10210_; 
wire u2__abc_52155_new_n10211_; 
wire u2__abc_52155_new_n10212_; 
wire u2__abc_52155_new_n10213_; 
wire u2__abc_52155_new_n10214_; 
wire u2__abc_52155_new_n10215_; 
wire u2__abc_52155_new_n10216_; 
wire u2__abc_52155_new_n10217_; 
wire u2__abc_52155_new_n10218_; 
wire u2__abc_52155_new_n10219_; 
wire u2__abc_52155_new_n10221_; 
wire u2__abc_52155_new_n10222_; 
wire u2__abc_52155_new_n10223_; 
wire u2__abc_52155_new_n10224_; 
wire u2__abc_52155_new_n10225_; 
wire u2__abc_52155_new_n10226_; 
wire u2__abc_52155_new_n10227_; 
wire u2__abc_52155_new_n10228_; 
wire u2__abc_52155_new_n10229_; 
wire u2__abc_52155_new_n10230_; 
wire u2__abc_52155_new_n10231_; 
wire u2__abc_52155_new_n10232_; 
wire u2__abc_52155_new_n10233_; 
wire u2__abc_52155_new_n10234_; 
wire u2__abc_52155_new_n10235_; 
wire u2__abc_52155_new_n10236_; 
wire u2__abc_52155_new_n10237_; 
wire u2__abc_52155_new_n10238_; 
wire u2__abc_52155_new_n10239_; 
wire u2__abc_52155_new_n10240_; 
wire u2__abc_52155_new_n10241_; 
wire u2__abc_52155_new_n10243_; 
wire u2__abc_52155_new_n10244_; 
wire u2__abc_52155_new_n10245_; 
wire u2__abc_52155_new_n10246_; 
wire u2__abc_52155_new_n10247_; 
wire u2__abc_52155_new_n10248_; 
wire u2__abc_52155_new_n10249_; 
wire u2__abc_52155_new_n10250_; 
wire u2__abc_52155_new_n10251_; 
wire u2__abc_52155_new_n10252_; 
wire u2__abc_52155_new_n10253_; 
wire u2__abc_52155_new_n10254_; 
wire u2__abc_52155_new_n10255_; 
wire u2__abc_52155_new_n10256_; 
wire u2__abc_52155_new_n10257_; 
wire u2__abc_52155_new_n10258_; 
wire u2__abc_52155_new_n10259_; 
wire u2__abc_52155_new_n10261_; 
wire u2__abc_52155_new_n10262_; 
wire u2__abc_52155_new_n10263_; 
wire u2__abc_52155_new_n10264_; 
wire u2__abc_52155_new_n10265_; 
wire u2__abc_52155_new_n10266_; 
wire u2__abc_52155_new_n10267_; 
wire u2__abc_52155_new_n10268_; 
wire u2__abc_52155_new_n10269_; 
wire u2__abc_52155_new_n10270_; 
wire u2__abc_52155_new_n10271_; 
wire u2__abc_52155_new_n10272_; 
wire u2__abc_52155_new_n10273_; 
wire u2__abc_52155_new_n10274_; 
wire u2__abc_52155_new_n10275_; 
wire u2__abc_52155_new_n10276_; 
wire u2__abc_52155_new_n10277_; 
wire u2__abc_52155_new_n10278_; 
wire u2__abc_52155_new_n10279_; 
wire u2__abc_52155_new_n10280_; 
wire u2__abc_52155_new_n10282_; 
wire u2__abc_52155_new_n10283_; 
wire u2__abc_52155_new_n10284_; 
wire u2__abc_52155_new_n10285_; 
wire u2__abc_52155_new_n10286_; 
wire u2__abc_52155_new_n10287_; 
wire u2__abc_52155_new_n10288_; 
wire u2__abc_52155_new_n10289_; 
wire u2__abc_52155_new_n10290_; 
wire u2__abc_52155_new_n10291_; 
wire u2__abc_52155_new_n10292_; 
wire u2__abc_52155_new_n10293_; 
wire u2__abc_52155_new_n10294_; 
wire u2__abc_52155_new_n10295_; 
wire u2__abc_52155_new_n10296_; 
wire u2__abc_52155_new_n10297_; 
wire u2__abc_52155_new_n10298_; 
wire u2__abc_52155_new_n10300_; 
wire u2__abc_52155_new_n10301_; 
wire u2__abc_52155_new_n10302_; 
wire u2__abc_52155_new_n10303_; 
wire u2__abc_52155_new_n10304_; 
wire u2__abc_52155_new_n10305_; 
wire u2__abc_52155_new_n10306_; 
wire u2__abc_52155_new_n10307_; 
wire u2__abc_52155_new_n10308_; 
wire u2__abc_52155_new_n10309_; 
wire u2__abc_52155_new_n10310_; 
wire u2__abc_52155_new_n10311_; 
wire u2__abc_52155_new_n10312_; 
wire u2__abc_52155_new_n10313_; 
wire u2__abc_52155_new_n10314_; 
wire u2__abc_52155_new_n10315_; 
wire u2__abc_52155_new_n10316_; 
wire u2__abc_52155_new_n10317_; 
wire u2__abc_52155_new_n10318_; 
wire u2__abc_52155_new_n10319_; 
wire u2__abc_52155_new_n10320_; 
wire u2__abc_52155_new_n10321_; 
wire u2__abc_52155_new_n10322_; 
wire u2__abc_52155_new_n10323_; 
wire u2__abc_52155_new_n10324_; 
wire u2__abc_52155_new_n10326_; 
wire u2__abc_52155_new_n10327_; 
wire u2__abc_52155_new_n10328_; 
wire u2__abc_52155_new_n10329_; 
wire u2__abc_52155_new_n10330_; 
wire u2__abc_52155_new_n10331_; 
wire u2__abc_52155_new_n10332_; 
wire u2__abc_52155_new_n10333_; 
wire u2__abc_52155_new_n10334_; 
wire u2__abc_52155_new_n10335_; 
wire u2__abc_52155_new_n10336_; 
wire u2__abc_52155_new_n10337_; 
wire u2__abc_52155_new_n10338_; 
wire u2__abc_52155_new_n10339_; 
wire u2__abc_52155_new_n10340_; 
wire u2__abc_52155_new_n10341_; 
wire u2__abc_52155_new_n10343_; 
wire u2__abc_52155_new_n10344_; 
wire u2__abc_52155_new_n10345_; 
wire u2__abc_52155_new_n10346_; 
wire u2__abc_52155_new_n10347_; 
wire u2__abc_52155_new_n10348_; 
wire u2__abc_52155_new_n10349_; 
wire u2__abc_52155_new_n10350_; 
wire u2__abc_52155_new_n10351_; 
wire u2__abc_52155_new_n10352_; 
wire u2__abc_52155_new_n10353_; 
wire u2__abc_52155_new_n10354_; 
wire u2__abc_52155_new_n10355_; 
wire u2__abc_52155_new_n10356_; 
wire u2__abc_52155_new_n10357_; 
wire u2__abc_52155_new_n10358_; 
wire u2__abc_52155_new_n10359_; 
wire u2__abc_52155_new_n10361_; 
wire u2__abc_52155_new_n10362_; 
wire u2__abc_52155_new_n10363_; 
wire u2__abc_52155_new_n10364_; 
wire u2__abc_52155_new_n10365_; 
wire u2__abc_52155_new_n10366_; 
wire u2__abc_52155_new_n10367_; 
wire u2__abc_52155_new_n10368_; 
wire u2__abc_52155_new_n10369_; 
wire u2__abc_52155_new_n10370_; 
wire u2__abc_52155_new_n10371_; 
wire u2__abc_52155_new_n10372_; 
wire u2__abc_52155_new_n10373_; 
wire u2__abc_52155_new_n10374_; 
wire u2__abc_52155_new_n10375_; 
wire u2__abc_52155_new_n10376_; 
wire u2__abc_52155_new_n10377_; 
wire u2__abc_52155_new_n10379_; 
wire u2__abc_52155_new_n10380_; 
wire u2__abc_52155_new_n10381_; 
wire u2__abc_52155_new_n10382_; 
wire u2__abc_52155_new_n10383_; 
wire u2__abc_52155_new_n10384_; 
wire u2__abc_52155_new_n10385_; 
wire u2__abc_52155_new_n10386_; 
wire u2__abc_52155_new_n10387_; 
wire u2__abc_52155_new_n10388_; 
wire u2__abc_52155_new_n10389_; 
wire u2__abc_52155_new_n10390_; 
wire u2__abc_52155_new_n10391_; 
wire u2__abc_52155_new_n10392_; 
wire u2__abc_52155_new_n10393_; 
wire u2__abc_52155_new_n10394_; 
wire u2__abc_52155_new_n10395_; 
wire u2__abc_52155_new_n10396_; 
wire u2__abc_52155_new_n10397_; 
wire u2__abc_52155_new_n10398_; 
wire u2__abc_52155_new_n10399_; 
wire u2__abc_52155_new_n10400_; 
wire u2__abc_52155_new_n10401_; 
wire u2__abc_52155_new_n10403_; 
wire u2__abc_52155_new_n10404_; 
wire u2__abc_52155_new_n10405_; 
wire u2__abc_52155_new_n10406_; 
wire u2__abc_52155_new_n10407_; 
wire u2__abc_52155_new_n10408_; 
wire u2__abc_52155_new_n10409_; 
wire u2__abc_52155_new_n10410_; 
wire u2__abc_52155_new_n10411_; 
wire u2__abc_52155_new_n10412_; 
wire u2__abc_52155_new_n10413_; 
wire u2__abc_52155_new_n10414_; 
wire u2__abc_52155_new_n10415_; 
wire u2__abc_52155_new_n10416_; 
wire u2__abc_52155_new_n10417_; 
wire u2__abc_52155_new_n10418_; 
wire u2__abc_52155_new_n10420_; 
wire u2__abc_52155_new_n10421_; 
wire u2__abc_52155_new_n10422_; 
wire u2__abc_52155_new_n10423_; 
wire u2__abc_52155_new_n10424_; 
wire u2__abc_52155_new_n10425_; 
wire u2__abc_52155_new_n10426_; 
wire u2__abc_52155_new_n10427_; 
wire u2__abc_52155_new_n10428_; 
wire u2__abc_52155_new_n10429_; 
wire u2__abc_52155_new_n10430_; 
wire u2__abc_52155_new_n10431_; 
wire u2__abc_52155_new_n10432_; 
wire u2__abc_52155_new_n10433_; 
wire u2__abc_52155_new_n10434_; 
wire u2__abc_52155_new_n10435_; 
wire u2__abc_52155_new_n10436_; 
wire u2__abc_52155_new_n10437_; 
wire u2__abc_52155_new_n10439_; 
wire u2__abc_52155_new_n10440_; 
wire u2__abc_52155_new_n10441_; 
wire u2__abc_52155_new_n10442_; 
wire u2__abc_52155_new_n10443_; 
wire u2__abc_52155_new_n10444_; 
wire u2__abc_52155_new_n10445_; 
wire u2__abc_52155_new_n10446_; 
wire u2__abc_52155_new_n10447_; 
wire u2__abc_52155_new_n10448_; 
wire u2__abc_52155_new_n10449_; 
wire u2__abc_52155_new_n10450_; 
wire u2__abc_52155_new_n10451_; 
wire u2__abc_52155_new_n10452_; 
wire u2__abc_52155_new_n10453_; 
wire u2__abc_52155_new_n10454_; 
wire u2__abc_52155_new_n10456_; 
wire u2__abc_52155_new_n10457_; 
wire u2__abc_52155_new_n10458_; 
wire u2__abc_52155_new_n10459_; 
wire u2__abc_52155_new_n10460_; 
wire u2__abc_52155_new_n10461_; 
wire u2__abc_52155_new_n10462_; 
wire u2__abc_52155_new_n10463_; 
wire u2__abc_52155_new_n10464_; 
wire u2__abc_52155_new_n10465_; 
wire u2__abc_52155_new_n10466_; 
wire u2__abc_52155_new_n10467_; 
wire u2__abc_52155_new_n10468_; 
wire u2__abc_52155_new_n10469_; 
wire u2__abc_52155_new_n10470_; 
wire u2__abc_52155_new_n10471_; 
wire u2__abc_52155_new_n10472_; 
wire u2__abc_52155_new_n10473_; 
wire u2__abc_52155_new_n10474_; 
wire u2__abc_52155_new_n10475_; 
wire u2__abc_52155_new_n10476_; 
wire u2__abc_52155_new_n10477_; 
wire u2__abc_52155_new_n10478_; 
wire u2__abc_52155_new_n10479_; 
wire u2__abc_52155_new_n10480_; 
wire u2__abc_52155_new_n10481_; 
wire u2__abc_52155_new_n10483_; 
wire u2__abc_52155_new_n10484_; 
wire u2__abc_52155_new_n10485_; 
wire u2__abc_52155_new_n10486_; 
wire u2__abc_52155_new_n10487_; 
wire u2__abc_52155_new_n10488_; 
wire u2__abc_52155_new_n10489_; 
wire u2__abc_52155_new_n10490_; 
wire u2__abc_52155_new_n10491_; 
wire u2__abc_52155_new_n10492_; 
wire u2__abc_52155_new_n10493_; 
wire u2__abc_52155_new_n10494_; 
wire u2__abc_52155_new_n10495_; 
wire u2__abc_52155_new_n10496_; 
wire u2__abc_52155_new_n10497_; 
wire u2__abc_52155_new_n10498_; 
wire u2__abc_52155_new_n10500_; 
wire u2__abc_52155_new_n10501_; 
wire u2__abc_52155_new_n10502_; 
wire u2__abc_52155_new_n10503_; 
wire u2__abc_52155_new_n10504_; 
wire u2__abc_52155_new_n10505_; 
wire u2__abc_52155_new_n10506_; 
wire u2__abc_52155_new_n10507_; 
wire u2__abc_52155_new_n10508_; 
wire u2__abc_52155_new_n10509_; 
wire u2__abc_52155_new_n10510_; 
wire u2__abc_52155_new_n10511_; 
wire u2__abc_52155_new_n10512_; 
wire u2__abc_52155_new_n10513_; 
wire u2__abc_52155_new_n10514_; 
wire u2__abc_52155_new_n10515_; 
wire u2__abc_52155_new_n10516_; 
wire u2__abc_52155_new_n10518_; 
wire u2__abc_52155_new_n10519_; 
wire u2__abc_52155_new_n10520_; 
wire u2__abc_52155_new_n10521_; 
wire u2__abc_52155_new_n10522_; 
wire u2__abc_52155_new_n10523_; 
wire u2__abc_52155_new_n10524_; 
wire u2__abc_52155_new_n10525_; 
wire u2__abc_52155_new_n10526_; 
wire u2__abc_52155_new_n10527_; 
wire u2__abc_52155_new_n10528_; 
wire u2__abc_52155_new_n10529_; 
wire u2__abc_52155_new_n10530_; 
wire u2__abc_52155_new_n10531_; 
wire u2__abc_52155_new_n10532_; 
wire u2__abc_52155_new_n10533_; 
wire u2__abc_52155_new_n10534_; 
wire u2__abc_52155_new_n10536_; 
wire u2__abc_52155_new_n10537_; 
wire u2__abc_52155_new_n10538_; 
wire u2__abc_52155_new_n10539_; 
wire u2__abc_52155_new_n10540_; 
wire u2__abc_52155_new_n10541_; 
wire u2__abc_52155_new_n10542_; 
wire u2__abc_52155_new_n10543_; 
wire u2__abc_52155_new_n10544_; 
wire u2__abc_52155_new_n10545_; 
wire u2__abc_52155_new_n10546_; 
wire u2__abc_52155_new_n10547_; 
wire u2__abc_52155_new_n10548_; 
wire u2__abc_52155_new_n10549_; 
wire u2__abc_52155_new_n10550_; 
wire u2__abc_52155_new_n10551_; 
wire u2__abc_52155_new_n10552_; 
wire u2__abc_52155_new_n10553_; 
wire u2__abc_52155_new_n10555_; 
wire u2__abc_52155_new_n10556_; 
wire u2__abc_52155_new_n10557_; 
wire u2__abc_52155_new_n10558_; 
wire u2__abc_52155_new_n10559_; 
wire u2__abc_52155_new_n10560_; 
wire u2__abc_52155_new_n10561_; 
wire u2__abc_52155_new_n10562_; 
wire u2__abc_52155_new_n10563_; 
wire u2__abc_52155_new_n10564_; 
wire u2__abc_52155_new_n10565_; 
wire u2__abc_52155_new_n10566_; 
wire u2__abc_52155_new_n10567_; 
wire u2__abc_52155_new_n10568_; 
wire u2__abc_52155_new_n10569_; 
wire u2__abc_52155_new_n10570_; 
wire u2__abc_52155_new_n10572_; 
wire u2__abc_52155_new_n10573_; 
wire u2__abc_52155_new_n10574_; 
wire u2__abc_52155_new_n10575_; 
wire u2__abc_52155_new_n10576_; 
wire u2__abc_52155_new_n10577_; 
wire u2__abc_52155_new_n10578_; 
wire u2__abc_52155_new_n10579_; 
wire u2__abc_52155_new_n10580_; 
wire u2__abc_52155_new_n10581_; 
wire u2__abc_52155_new_n10582_; 
wire u2__abc_52155_new_n10583_; 
wire u2__abc_52155_new_n10584_; 
wire u2__abc_52155_new_n10585_; 
wire u2__abc_52155_new_n10586_; 
wire u2__abc_52155_new_n10587_; 
wire u2__abc_52155_new_n10589_; 
wire u2__abc_52155_new_n10590_; 
wire u2__abc_52155_new_n10591_; 
wire u2__abc_52155_new_n10592_; 
wire u2__abc_52155_new_n10593_; 
wire u2__abc_52155_new_n10594_; 
wire u2__abc_52155_new_n10595_; 
wire u2__abc_52155_new_n10596_; 
wire u2__abc_52155_new_n10597_; 
wire u2__abc_52155_new_n10598_; 
wire u2__abc_52155_new_n10599_; 
wire u2__abc_52155_new_n10600_; 
wire u2__abc_52155_new_n10601_; 
wire u2__abc_52155_new_n10602_; 
wire u2__abc_52155_new_n10603_; 
wire u2__abc_52155_new_n10604_; 
wire u2__abc_52155_new_n10606_; 
wire u2__abc_52155_new_n10607_; 
wire u2__abc_52155_new_n10608_; 
wire u2__abc_52155_new_n10609_; 
wire u2__abc_52155_new_n10610_; 
wire u2__abc_52155_new_n10611_; 
wire u2__abc_52155_new_n10612_; 
wire u2__abc_52155_new_n10613_; 
wire u2__abc_52155_new_n10614_; 
wire u2__abc_52155_new_n10615_; 
wire u2__abc_52155_new_n10616_; 
wire u2__abc_52155_new_n10617_; 
wire u2__abc_52155_new_n10618_; 
wire u2__abc_52155_new_n10619_; 
wire u2__abc_52155_new_n10620_; 
wire u2__abc_52155_new_n10621_; 
wire u2__abc_52155_new_n10622_; 
wire u2__abc_52155_new_n10623_; 
wire u2__abc_52155_new_n10624_; 
wire u2__abc_52155_new_n10625_; 
wire u2__abc_52155_new_n10626_; 
wire u2__abc_52155_new_n10627_; 
wire u2__abc_52155_new_n10628_; 
wire u2__abc_52155_new_n10629_; 
wire u2__abc_52155_new_n10630_; 
wire u2__abc_52155_new_n10631_; 
wire u2__abc_52155_new_n10632_; 
wire u2__abc_52155_new_n10633_; 
wire u2__abc_52155_new_n10634_; 
wire u2__abc_52155_new_n10635_; 
wire u2__abc_52155_new_n10637_; 
wire u2__abc_52155_new_n10638_; 
wire u2__abc_52155_new_n10639_; 
wire u2__abc_52155_new_n10640_; 
wire u2__abc_52155_new_n10641_; 
wire u2__abc_52155_new_n10642_; 
wire u2__abc_52155_new_n10643_; 
wire u2__abc_52155_new_n10644_; 
wire u2__abc_52155_new_n10645_; 
wire u2__abc_52155_new_n10646_; 
wire u2__abc_52155_new_n10647_; 
wire u2__abc_52155_new_n10648_; 
wire u2__abc_52155_new_n10649_; 
wire u2__abc_52155_new_n10650_; 
wire u2__abc_52155_new_n10651_; 
wire u2__abc_52155_new_n10652_; 
wire u2__abc_52155_new_n10654_; 
wire u2__abc_52155_new_n10655_; 
wire u2__abc_52155_new_n10656_; 
wire u2__abc_52155_new_n10657_; 
wire u2__abc_52155_new_n10658_; 
wire u2__abc_52155_new_n10659_; 
wire u2__abc_52155_new_n10660_; 
wire u2__abc_52155_new_n10661_; 
wire u2__abc_52155_new_n10662_; 
wire u2__abc_52155_new_n10663_; 
wire u2__abc_52155_new_n10664_; 
wire u2__abc_52155_new_n10665_; 
wire u2__abc_52155_new_n10666_; 
wire u2__abc_52155_new_n10667_; 
wire u2__abc_52155_new_n10668_; 
wire u2__abc_52155_new_n10669_; 
wire u2__abc_52155_new_n10670_; 
wire u2__abc_52155_new_n10671_; 
wire u2__abc_52155_new_n10673_; 
wire u2__abc_52155_new_n10674_; 
wire u2__abc_52155_new_n10675_; 
wire u2__abc_52155_new_n10676_; 
wire u2__abc_52155_new_n10677_; 
wire u2__abc_52155_new_n10678_; 
wire u2__abc_52155_new_n10679_; 
wire u2__abc_52155_new_n10680_; 
wire u2__abc_52155_new_n10681_; 
wire u2__abc_52155_new_n10682_; 
wire u2__abc_52155_new_n10683_; 
wire u2__abc_52155_new_n10684_; 
wire u2__abc_52155_new_n10685_; 
wire u2__abc_52155_new_n10686_; 
wire u2__abc_52155_new_n10687_; 
wire u2__abc_52155_new_n10688_; 
wire u2__abc_52155_new_n10690_; 
wire u2__abc_52155_new_n10691_; 
wire u2__abc_52155_new_n10692_; 
wire u2__abc_52155_new_n10693_; 
wire u2__abc_52155_new_n10694_; 
wire u2__abc_52155_new_n10695_; 
wire u2__abc_52155_new_n10696_; 
wire u2__abc_52155_new_n10697_; 
wire u2__abc_52155_new_n10698_; 
wire u2__abc_52155_new_n10699_; 
wire u2__abc_52155_new_n10700_; 
wire u2__abc_52155_new_n10701_; 
wire u2__abc_52155_new_n10702_; 
wire u2__abc_52155_new_n10703_; 
wire u2__abc_52155_new_n10704_; 
wire u2__abc_52155_new_n10705_; 
wire u2__abc_52155_new_n10706_; 
wire u2__abc_52155_new_n10707_; 
wire u2__abc_52155_new_n10708_; 
wire u2__abc_52155_new_n10709_; 
wire u2__abc_52155_new_n10710_; 
wire u2__abc_52155_new_n10711_; 
wire u2__abc_52155_new_n10713_; 
wire u2__abc_52155_new_n10714_; 
wire u2__abc_52155_new_n10715_; 
wire u2__abc_52155_new_n10716_; 
wire u2__abc_52155_new_n10717_; 
wire u2__abc_52155_new_n10718_; 
wire u2__abc_52155_new_n10719_; 
wire u2__abc_52155_new_n10720_; 
wire u2__abc_52155_new_n10721_; 
wire u2__abc_52155_new_n10722_; 
wire u2__abc_52155_new_n10723_; 
wire u2__abc_52155_new_n10724_; 
wire u2__abc_52155_new_n10725_; 
wire u2__abc_52155_new_n10726_; 
wire u2__abc_52155_new_n10727_; 
wire u2__abc_52155_new_n10728_; 
wire u2__abc_52155_new_n10730_; 
wire u2__abc_52155_new_n10731_; 
wire u2__abc_52155_new_n10732_; 
wire u2__abc_52155_new_n10733_; 
wire u2__abc_52155_new_n10734_; 
wire u2__abc_52155_new_n10735_; 
wire u2__abc_52155_new_n10736_; 
wire u2__abc_52155_new_n10737_; 
wire u2__abc_52155_new_n10738_; 
wire u2__abc_52155_new_n10739_; 
wire u2__abc_52155_new_n10740_; 
wire u2__abc_52155_new_n10741_; 
wire u2__abc_52155_new_n10742_; 
wire u2__abc_52155_new_n10743_; 
wire u2__abc_52155_new_n10744_; 
wire u2__abc_52155_new_n10745_; 
wire u2__abc_52155_new_n10746_; 
wire u2__abc_52155_new_n10747_; 
wire u2__abc_52155_new_n10749_; 
wire u2__abc_52155_new_n10750_; 
wire u2__abc_52155_new_n10751_; 
wire u2__abc_52155_new_n10752_; 
wire u2__abc_52155_new_n10753_; 
wire u2__abc_52155_new_n10754_; 
wire u2__abc_52155_new_n10755_; 
wire u2__abc_52155_new_n10756_; 
wire u2__abc_52155_new_n10757_; 
wire u2__abc_52155_new_n10758_; 
wire u2__abc_52155_new_n10759_; 
wire u2__abc_52155_new_n10760_; 
wire u2__abc_52155_new_n10761_; 
wire u2__abc_52155_new_n10762_; 
wire u2__abc_52155_new_n10763_; 
wire u2__abc_52155_new_n10764_; 
wire u2__abc_52155_new_n10766_; 
wire u2__abc_52155_new_n10767_; 
wire u2__abc_52155_new_n10768_; 
wire u2__abc_52155_new_n10769_; 
wire u2__abc_52155_new_n10770_; 
wire u2__abc_52155_new_n10771_; 
wire u2__abc_52155_new_n10772_; 
wire u2__abc_52155_new_n10773_; 
wire u2__abc_52155_new_n10774_; 
wire u2__abc_52155_new_n10775_; 
wire u2__abc_52155_new_n10776_; 
wire u2__abc_52155_new_n10777_; 
wire u2__abc_52155_new_n10778_; 
wire u2__abc_52155_new_n10779_; 
wire u2__abc_52155_new_n10780_; 
wire u2__abc_52155_new_n10781_; 
wire u2__abc_52155_new_n10782_; 
wire u2__abc_52155_new_n10783_; 
wire u2__abc_52155_new_n10784_; 
wire u2__abc_52155_new_n10785_; 
wire u2__abc_52155_new_n10786_; 
wire u2__abc_52155_new_n10787_; 
wire u2__abc_52155_new_n10788_; 
wire u2__abc_52155_new_n10789_; 
wire u2__abc_52155_new_n10790_; 
wire u2__abc_52155_new_n10791_; 
wire u2__abc_52155_new_n10792_; 
wire u2__abc_52155_new_n10793_; 
wire u2__abc_52155_new_n10795_; 
wire u2__abc_52155_new_n10796_; 
wire u2__abc_52155_new_n10797_; 
wire u2__abc_52155_new_n10798_; 
wire u2__abc_52155_new_n10799_; 
wire u2__abc_52155_new_n10800_; 
wire u2__abc_52155_new_n10801_; 
wire u2__abc_52155_new_n10802_; 
wire u2__abc_52155_new_n10803_; 
wire u2__abc_52155_new_n10804_; 
wire u2__abc_52155_new_n10805_; 
wire u2__abc_52155_new_n10806_; 
wire u2__abc_52155_new_n10807_; 
wire u2__abc_52155_new_n10808_; 
wire u2__abc_52155_new_n10809_; 
wire u2__abc_52155_new_n10810_; 
wire u2__abc_52155_new_n10812_; 
wire u2__abc_52155_new_n10813_; 
wire u2__abc_52155_new_n10814_; 
wire u2__abc_52155_new_n10815_; 
wire u2__abc_52155_new_n10816_; 
wire u2__abc_52155_new_n10817_; 
wire u2__abc_52155_new_n10818_; 
wire u2__abc_52155_new_n10819_; 
wire u2__abc_52155_new_n10820_; 
wire u2__abc_52155_new_n10821_; 
wire u2__abc_52155_new_n10822_; 
wire u2__abc_52155_new_n10823_; 
wire u2__abc_52155_new_n10824_; 
wire u2__abc_52155_new_n10825_; 
wire u2__abc_52155_new_n10826_; 
wire u2__abc_52155_new_n10827_; 
wire u2__abc_52155_new_n10828_; 
wire u2__abc_52155_new_n10829_; 
wire u2__abc_52155_new_n10830_; 
wire u2__abc_52155_new_n10832_; 
wire u2__abc_52155_new_n10833_; 
wire u2__abc_52155_new_n10834_; 
wire u2__abc_52155_new_n10835_; 
wire u2__abc_52155_new_n10836_; 
wire u2__abc_52155_new_n10837_; 
wire u2__abc_52155_new_n10838_; 
wire u2__abc_52155_new_n10839_; 
wire u2__abc_52155_new_n10840_; 
wire u2__abc_52155_new_n10841_; 
wire u2__abc_52155_new_n10842_; 
wire u2__abc_52155_new_n10843_; 
wire u2__abc_52155_new_n10844_; 
wire u2__abc_52155_new_n10845_; 
wire u2__abc_52155_new_n10846_; 
wire u2__abc_52155_new_n10847_; 
wire u2__abc_52155_new_n10848_; 
wire u2__abc_52155_new_n10850_; 
wire u2__abc_52155_new_n10851_; 
wire u2__abc_52155_new_n10852_; 
wire u2__abc_52155_new_n10853_; 
wire u2__abc_52155_new_n10854_; 
wire u2__abc_52155_new_n10855_; 
wire u2__abc_52155_new_n10856_; 
wire u2__abc_52155_new_n10857_; 
wire u2__abc_52155_new_n10858_; 
wire u2__abc_52155_new_n10859_; 
wire u2__abc_52155_new_n10860_; 
wire u2__abc_52155_new_n10861_; 
wire u2__abc_52155_new_n10862_; 
wire u2__abc_52155_new_n10863_; 
wire u2__abc_52155_new_n10864_; 
wire u2__abc_52155_new_n10865_; 
wire u2__abc_52155_new_n10866_; 
wire u2__abc_52155_new_n10867_; 
wire u2__abc_52155_new_n10868_; 
wire u2__abc_52155_new_n10869_; 
wire u2__abc_52155_new_n10870_; 
wire u2__abc_52155_new_n10871_; 
wire u2__abc_52155_new_n10873_; 
wire u2__abc_52155_new_n10874_; 
wire u2__abc_52155_new_n10875_; 
wire u2__abc_52155_new_n10876_; 
wire u2__abc_52155_new_n10877_; 
wire u2__abc_52155_new_n10878_; 
wire u2__abc_52155_new_n10879_; 
wire u2__abc_52155_new_n10880_; 
wire u2__abc_52155_new_n10881_; 
wire u2__abc_52155_new_n10882_; 
wire u2__abc_52155_new_n10883_; 
wire u2__abc_52155_new_n10884_; 
wire u2__abc_52155_new_n10885_; 
wire u2__abc_52155_new_n10886_; 
wire u2__abc_52155_new_n10887_; 
wire u2__abc_52155_new_n10888_; 
wire u2__abc_52155_new_n10890_; 
wire u2__abc_52155_new_n10891_; 
wire u2__abc_52155_new_n10892_; 
wire u2__abc_52155_new_n10893_; 
wire u2__abc_52155_new_n10894_; 
wire u2__abc_52155_new_n10895_; 
wire u2__abc_52155_new_n10896_; 
wire u2__abc_52155_new_n10897_; 
wire u2__abc_52155_new_n10898_; 
wire u2__abc_52155_new_n10899_; 
wire u2__abc_52155_new_n10900_; 
wire u2__abc_52155_new_n10901_; 
wire u2__abc_52155_new_n10902_; 
wire u2__abc_52155_new_n10903_; 
wire u2__abc_52155_new_n10904_; 
wire u2__abc_52155_new_n10905_; 
wire u2__abc_52155_new_n10907_; 
wire u2__abc_52155_new_n10908_; 
wire u2__abc_52155_new_n10909_; 
wire u2__abc_52155_new_n10910_; 
wire u2__abc_52155_new_n10911_; 
wire u2__abc_52155_new_n10912_; 
wire u2__abc_52155_new_n10913_; 
wire u2__abc_52155_new_n10914_; 
wire u2__abc_52155_new_n10915_; 
wire u2__abc_52155_new_n10916_; 
wire u2__abc_52155_new_n10917_; 
wire u2__abc_52155_new_n10918_; 
wire u2__abc_52155_new_n10919_; 
wire u2__abc_52155_new_n10920_; 
wire u2__abc_52155_new_n10921_; 
wire u2__abc_52155_new_n10922_; 
wire u2__abc_52155_new_n10924_; 
wire u2__abc_52155_new_n10925_; 
wire u2__abc_52155_new_n10926_; 
wire u2__abc_52155_new_n10927_; 
wire u2__abc_52155_new_n10928_; 
wire u2__abc_52155_new_n10929_; 
wire u2__abc_52155_new_n10930_; 
wire u2__abc_52155_new_n10931_; 
wire u2__abc_52155_new_n10932_; 
wire u2__abc_52155_new_n10933_; 
wire u2__abc_52155_new_n10934_; 
wire u2__abc_52155_new_n10935_; 
wire u2__abc_52155_new_n10936_; 
wire u2__abc_52155_new_n10937_; 
wire u2__abc_52155_new_n10938_; 
wire u2__abc_52155_new_n10939_; 
wire u2__abc_52155_new_n10940_; 
wire u2__abc_52155_new_n10941_; 
wire u2__abc_52155_new_n10942_; 
wire u2__abc_52155_new_n10943_; 
wire u2__abc_52155_new_n10944_; 
wire u2__abc_52155_new_n10945_; 
wire u2__abc_52155_new_n10946_; 
wire u2__abc_52155_new_n10947_; 
wire u2__abc_52155_new_n10949_; 
wire u2__abc_52155_new_n10950_; 
wire u2__abc_52155_new_n10951_; 
wire u2__abc_52155_new_n10952_; 
wire u2__abc_52155_new_n10953_; 
wire u2__abc_52155_new_n10954_; 
wire u2__abc_52155_new_n10955_; 
wire u2__abc_52155_new_n10956_; 
wire u2__abc_52155_new_n10957_; 
wire u2__abc_52155_new_n10958_; 
wire u2__abc_52155_new_n10959_; 
wire u2__abc_52155_new_n10960_; 
wire u2__abc_52155_new_n10961_; 
wire u2__abc_52155_new_n10962_; 
wire u2__abc_52155_new_n10963_; 
wire u2__abc_52155_new_n10964_; 
wire u2__abc_52155_new_n10966_; 
wire u2__abc_52155_new_n10967_; 
wire u2__abc_52155_new_n10968_; 
wire u2__abc_52155_new_n10969_; 
wire u2__abc_52155_new_n10970_; 
wire u2__abc_52155_new_n10971_; 
wire u2__abc_52155_new_n10972_; 
wire u2__abc_52155_new_n10973_; 
wire u2__abc_52155_new_n10974_; 
wire u2__abc_52155_new_n10975_; 
wire u2__abc_52155_new_n10976_; 
wire u2__abc_52155_new_n10977_; 
wire u2__abc_52155_new_n10978_; 
wire u2__abc_52155_new_n10979_; 
wire u2__abc_52155_new_n10980_; 
wire u2__abc_52155_new_n10981_; 
wire u2__abc_52155_new_n10982_; 
wire u2__abc_52155_new_n10983_; 
wire u2__abc_52155_new_n10984_; 
wire u2__abc_52155_new_n10986_; 
wire u2__abc_52155_new_n10987_; 
wire u2__abc_52155_new_n10988_; 
wire u2__abc_52155_new_n10989_; 
wire u2__abc_52155_new_n10990_; 
wire u2__abc_52155_new_n10991_; 
wire u2__abc_52155_new_n10992_; 
wire u2__abc_52155_new_n10993_; 
wire u2__abc_52155_new_n10994_; 
wire u2__abc_52155_new_n10995_; 
wire u2__abc_52155_new_n10996_; 
wire u2__abc_52155_new_n10997_; 
wire u2__abc_52155_new_n10998_; 
wire u2__abc_52155_new_n10999_; 
wire u2__abc_52155_new_n11000_; 
wire u2__abc_52155_new_n11001_; 
wire u2__abc_52155_new_n11003_; 
wire u2__abc_52155_new_n11004_; 
wire u2__abc_52155_new_n11005_; 
wire u2__abc_52155_new_n11006_; 
wire u2__abc_52155_new_n11007_; 
wire u2__abc_52155_new_n11008_; 
wire u2__abc_52155_new_n11009_; 
wire u2__abc_52155_new_n11010_; 
wire u2__abc_52155_new_n11011_; 
wire u2__abc_52155_new_n11012_; 
wire u2__abc_52155_new_n11013_; 
wire u2__abc_52155_new_n11014_; 
wire u2__abc_52155_new_n11015_; 
wire u2__abc_52155_new_n11016_; 
wire u2__abc_52155_new_n11017_; 
wire u2__abc_52155_new_n11018_; 
wire u2__abc_52155_new_n11019_; 
wire u2__abc_52155_new_n11020_; 
wire u2__abc_52155_new_n11022_; 
wire u2__abc_52155_new_n11023_; 
wire u2__abc_52155_new_n11024_; 
wire u2__abc_52155_new_n11025_; 
wire u2__abc_52155_new_n11026_; 
wire u2__abc_52155_new_n11027_; 
wire u2__abc_52155_new_n11028_; 
wire u2__abc_52155_new_n11029_; 
wire u2__abc_52155_new_n11030_; 
wire u2__abc_52155_new_n11031_; 
wire u2__abc_52155_new_n11032_; 
wire u2__abc_52155_new_n11033_; 
wire u2__abc_52155_new_n11034_; 
wire u2__abc_52155_new_n11035_; 
wire u2__abc_52155_new_n11036_; 
wire u2__abc_52155_new_n11037_; 
wire u2__abc_52155_new_n11039_; 
wire u2__abc_52155_new_n11040_; 
wire u2__abc_52155_new_n11041_; 
wire u2__abc_52155_new_n11042_; 
wire u2__abc_52155_new_n11043_; 
wire u2__abc_52155_new_n11044_; 
wire u2__abc_52155_new_n11045_; 
wire u2__abc_52155_new_n11046_; 
wire u2__abc_52155_new_n11047_; 
wire u2__abc_52155_new_n11048_; 
wire u2__abc_52155_new_n11049_; 
wire u2__abc_52155_new_n11050_; 
wire u2__abc_52155_new_n11051_; 
wire u2__abc_52155_new_n11052_; 
wire u2__abc_52155_new_n11053_; 
wire u2__abc_52155_new_n11054_; 
wire u2__abc_52155_new_n11055_; 
wire u2__abc_52155_new_n11056_; 
wire u2__abc_52155_new_n11058_; 
wire u2__abc_52155_new_n11059_; 
wire u2__abc_52155_new_n11060_; 
wire u2__abc_52155_new_n11061_; 
wire u2__abc_52155_new_n11062_; 
wire u2__abc_52155_new_n11063_; 
wire u2__abc_52155_new_n11064_; 
wire u2__abc_52155_new_n11065_; 
wire u2__abc_52155_new_n11066_; 
wire u2__abc_52155_new_n11067_; 
wire u2__abc_52155_new_n11068_; 
wire u2__abc_52155_new_n11069_; 
wire u2__abc_52155_new_n11070_; 
wire u2__abc_52155_new_n11071_; 
wire u2__abc_52155_new_n11072_; 
wire u2__abc_52155_new_n11073_; 
wire u2__abc_52155_new_n11075_; 
wire u2__abc_52155_new_n11076_; 
wire u2__abc_52155_new_n11077_; 
wire u2__abc_52155_new_n11078_; 
wire u2__abc_52155_new_n11079_; 
wire u2__abc_52155_new_n11080_; 
wire u2__abc_52155_new_n11081_; 
wire u2__abc_52155_new_n11082_; 
wire u2__abc_52155_new_n11083_; 
wire u2__abc_52155_new_n11084_; 
wire u2__abc_52155_new_n11085_; 
wire u2__abc_52155_new_n11086_; 
wire u2__abc_52155_new_n11087_; 
wire u2__abc_52155_new_n11088_; 
wire u2__abc_52155_new_n11089_; 
wire u2__abc_52155_new_n11090_; 
wire u2__abc_52155_new_n11091_; 
wire u2__abc_52155_new_n11092_; 
wire u2__abc_52155_new_n11093_; 
wire u2__abc_52155_new_n11094_; 
wire u2__abc_52155_new_n11095_; 
wire u2__abc_52155_new_n11096_; 
wire u2__abc_52155_new_n11097_; 
wire u2__abc_52155_new_n11098_; 
wire u2__abc_52155_new_n11099_; 
wire u2__abc_52155_new_n11100_; 
wire u2__abc_52155_new_n11101_; 
wire u2__abc_52155_new_n11102_; 
wire u2__abc_52155_new_n11103_; 
wire u2__abc_52155_new_n11104_; 
wire u2__abc_52155_new_n11105_; 
wire u2__abc_52155_new_n11106_; 
wire u2__abc_52155_new_n11107_; 
wire u2__abc_52155_new_n11108_; 
wire u2__abc_52155_new_n11109_; 
wire u2__abc_52155_new_n11111_; 
wire u2__abc_52155_new_n11112_; 
wire u2__abc_52155_new_n11113_; 
wire u2__abc_52155_new_n11114_; 
wire u2__abc_52155_new_n11115_; 
wire u2__abc_52155_new_n11116_; 
wire u2__abc_52155_new_n11117_; 
wire u2__abc_52155_new_n11118_; 
wire u2__abc_52155_new_n11119_; 
wire u2__abc_52155_new_n11120_; 
wire u2__abc_52155_new_n11121_; 
wire u2__abc_52155_new_n11122_; 
wire u2__abc_52155_new_n11123_; 
wire u2__abc_52155_new_n11124_; 
wire u2__abc_52155_new_n11125_; 
wire u2__abc_52155_new_n11126_; 
wire u2__abc_52155_new_n11128_; 
wire u2__abc_52155_new_n11129_; 
wire u2__abc_52155_new_n11130_; 
wire u2__abc_52155_new_n11131_; 
wire u2__abc_52155_new_n11132_; 
wire u2__abc_52155_new_n11133_; 
wire u2__abc_52155_new_n11134_; 
wire u2__abc_52155_new_n11135_; 
wire u2__abc_52155_new_n11136_; 
wire u2__abc_52155_new_n11137_; 
wire u2__abc_52155_new_n11138_; 
wire u2__abc_52155_new_n11139_; 
wire u2__abc_52155_new_n11140_; 
wire u2__abc_52155_new_n11141_; 
wire u2__abc_52155_new_n11142_; 
wire u2__abc_52155_new_n11143_; 
wire u2__abc_52155_new_n11144_; 
wire u2__abc_52155_new_n11145_; 
wire u2__abc_52155_new_n11146_; 
wire u2__abc_52155_new_n11148_; 
wire u2__abc_52155_new_n11149_; 
wire u2__abc_52155_new_n11150_; 
wire u2__abc_52155_new_n11151_; 
wire u2__abc_52155_new_n11152_; 
wire u2__abc_52155_new_n11153_; 
wire u2__abc_52155_new_n11154_; 
wire u2__abc_52155_new_n11155_; 
wire u2__abc_52155_new_n11156_; 
wire u2__abc_52155_new_n11157_; 
wire u2__abc_52155_new_n11158_; 
wire u2__abc_52155_new_n11159_; 
wire u2__abc_52155_new_n11160_; 
wire u2__abc_52155_new_n11161_; 
wire u2__abc_52155_new_n11162_; 
wire u2__abc_52155_new_n11163_; 
wire u2__abc_52155_new_n11165_; 
wire u2__abc_52155_new_n11166_; 
wire u2__abc_52155_new_n11167_; 
wire u2__abc_52155_new_n11168_; 
wire u2__abc_52155_new_n11169_; 
wire u2__abc_52155_new_n11170_; 
wire u2__abc_52155_new_n11171_; 
wire u2__abc_52155_new_n11172_; 
wire u2__abc_52155_new_n11173_; 
wire u2__abc_52155_new_n11174_; 
wire u2__abc_52155_new_n11175_; 
wire u2__abc_52155_new_n11176_; 
wire u2__abc_52155_new_n11177_; 
wire u2__abc_52155_new_n11178_; 
wire u2__abc_52155_new_n11179_; 
wire u2__abc_52155_new_n11180_; 
wire u2__abc_52155_new_n11181_; 
wire u2__abc_52155_new_n11182_; 
wire u2__abc_52155_new_n11184_; 
wire u2__abc_52155_new_n11185_; 
wire u2__abc_52155_new_n11186_; 
wire u2__abc_52155_new_n11187_; 
wire u2__abc_52155_new_n11188_; 
wire u2__abc_52155_new_n11189_; 
wire u2__abc_52155_new_n11190_; 
wire u2__abc_52155_new_n11191_; 
wire u2__abc_52155_new_n11192_; 
wire u2__abc_52155_new_n11193_; 
wire u2__abc_52155_new_n11194_; 
wire u2__abc_52155_new_n11195_; 
wire u2__abc_52155_new_n11196_; 
wire u2__abc_52155_new_n11197_; 
wire u2__abc_52155_new_n11198_; 
wire u2__abc_52155_new_n11199_; 
wire u2__abc_52155_new_n11201_; 
wire u2__abc_52155_new_n11202_; 
wire u2__abc_52155_new_n11203_; 
wire u2__abc_52155_new_n11204_; 
wire u2__abc_52155_new_n11205_; 
wire u2__abc_52155_new_n11206_; 
wire u2__abc_52155_new_n11207_; 
wire u2__abc_52155_new_n11208_; 
wire u2__abc_52155_new_n11209_; 
wire u2__abc_52155_new_n11210_; 
wire u2__abc_52155_new_n11211_; 
wire u2__abc_52155_new_n11212_; 
wire u2__abc_52155_new_n11213_; 
wire u2__abc_52155_new_n11214_; 
wire u2__abc_52155_new_n11215_; 
wire u2__abc_52155_new_n11216_; 
wire u2__abc_52155_new_n11217_; 
wire u2__abc_52155_new_n11218_; 
wire u2__abc_52155_new_n11220_; 
wire u2__abc_52155_new_n11221_; 
wire u2__abc_52155_new_n11222_; 
wire u2__abc_52155_new_n11223_; 
wire u2__abc_52155_new_n11224_; 
wire u2__abc_52155_new_n11225_; 
wire u2__abc_52155_new_n11226_; 
wire u2__abc_52155_new_n11227_; 
wire u2__abc_52155_new_n11228_; 
wire u2__abc_52155_new_n11229_; 
wire u2__abc_52155_new_n11230_; 
wire u2__abc_52155_new_n11231_; 
wire u2__abc_52155_new_n11232_; 
wire u2__abc_52155_new_n11233_; 
wire u2__abc_52155_new_n11234_; 
wire u2__abc_52155_new_n11235_; 
wire u2__abc_52155_new_n11237_; 
wire u2__abc_52155_new_n11238_; 
wire u2__abc_52155_new_n11239_; 
wire u2__abc_52155_new_n11240_; 
wire u2__abc_52155_new_n11241_; 
wire u2__abc_52155_new_n11242_; 
wire u2__abc_52155_new_n11243_; 
wire u2__abc_52155_new_n11244_; 
wire u2__abc_52155_new_n11245_; 
wire u2__abc_52155_new_n11246_; 
wire u2__abc_52155_new_n11247_; 
wire u2__abc_52155_new_n11248_; 
wire u2__abc_52155_new_n11249_; 
wire u2__abc_52155_new_n11250_; 
wire u2__abc_52155_new_n11251_; 
wire u2__abc_52155_new_n11252_; 
wire u2__abc_52155_new_n11253_; 
wire u2__abc_52155_new_n11254_; 
wire u2__abc_52155_new_n11255_; 
wire u2__abc_52155_new_n11256_; 
wire u2__abc_52155_new_n11257_; 
wire u2__abc_52155_new_n11258_; 
wire u2__abc_52155_new_n11259_; 
wire u2__abc_52155_new_n11260_; 
wire u2__abc_52155_new_n11261_; 
wire u2__abc_52155_new_n11262_; 
wire u2__abc_52155_new_n11263_; 
wire u2__abc_52155_new_n11264_; 
wire u2__abc_52155_new_n11265_; 
wire u2__abc_52155_new_n11267_; 
wire u2__abc_52155_new_n11268_; 
wire u2__abc_52155_new_n11269_; 
wire u2__abc_52155_new_n11270_; 
wire u2__abc_52155_new_n11271_; 
wire u2__abc_52155_new_n11272_; 
wire u2__abc_52155_new_n11273_; 
wire u2__abc_52155_new_n11274_; 
wire u2__abc_52155_new_n11275_; 
wire u2__abc_52155_new_n11276_; 
wire u2__abc_52155_new_n11277_; 
wire u2__abc_52155_new_n11278_; 
wire u2__abc_52155_new_n11279_; 
wire u2__abc_52155_new_n11280_; 
wire u2__abc_52155_new_n11281_; 
wire u2__abc_52155_new_n11282_; 
wire u2__abc_52155_new_n11284_; 
wire u2__abc_52155_new_n11285_; 
wire u2__abc_52155_new_n11286_; 
wire u2__abc_52155_new_n11287_; 
wire u2__abc_52155_new_n11288_; 
wire u2__abc_52155_new_n11289_; 
wire u2__abc_52155_new_n11290_; 
wire u2__abc_52155_new_n11291_; 
wire u2__abc_52155_new_n11292_; 
wire u2__abc_52155_new_n11293_; 
wire u2__abc_52155_new_n11294_; 
wire u2__abc_52155_new_n11295_; 
wire u2__abc_52155_new_n11296_; 
wire u2__abc_52155_new_n11297_; 
wire u2__abc_52155_new_n11298_; 
wire u2__abc_52155_new_n11299_; 
wire u2__abc_52155_new_n11300_; 
wire u2__abc_52155_new_n11301_; 
wire u2__abc_52155_new_n11302_; 
wire u2__abc_52155_new_n11304_; 
wire u2__abc_52155_new_n11305_; 
wire u2__abc_52155_new_n11306_; 
wire u2__abc_52155_new_n11307_; 
wire u2__abc_52155_new_n11308_; 
wire u2__abc_52155_new_n11309_; 
wire u2__abc_52155_new_n11310_; 
wire u2__abc_52155_new_n11311_; 
wire u2__abc_52155_new_n11312_; 
wire u2__abc_52155_new_n11313_; 
wire u2__abc_52155_new_n11314_; 
wire u2__abc_52155_new_n11315_; 
wire u2__abc_52155_new_n11316_; 
wire u2__abc_52155_new_n11317_; 
wire u2__abc_52155_new_n11318_; 
wire u2__abc_52155_new_n11319_; 
wire u2__abc_52155_new_n11321_; 
wire u2__abc_52155_new_n11322_; 
wire u2__abc_52155_new_n11323_; 
wire u2__abc_52155_new_n11324_; 
wire u2__abc_52155_new_n11325_; 
wire u2__abc_52155_new_n11326_; 
wire u2__abc_52155_new_n11327_; 
wire u2__abc_52155_new_n11328_; 
wire u2__abc_52155_new_n11329_; 
wire u2__abc_52155_new_n11330_; 
wire u2__abc_52155_new_n11331_; 
wire u2__abc_52155_new_n11332_; 
wire u2__abc_52155_new_n11333_; 
wire u2__abc_52155_new_n11334_; 
wire u2__abc_52155_new_n11335_; 
wire u2__abc_52155_new_n11336_; 
wire u2__abc_52155_new_n11337_; 
wire u2__abc_52155_new_n11338_; 
wire u2__abc_52155_new_n11339_; 
wire u2__abc_52155_new_n11340_; 
wire u2__abc_52155_new_n11342_; 
wire u2__abc_52155_new_n11343_; 
wire u2__abc_52155_new_n11344_; 
wire u2__abc_52155_new_n11345_; 
wire u2__abc_52155_new_n11346_; 
wire u2__abc_52155_new_n11347_; 
wire u2__abc_52155_new_n11348_; 
wire u2__abc_52155_new_n11349_; 
wire u2__abc_52155_new_n11350_; 
wire u2__abc_52155_new_n11351_; 
wire u2__abc_52155_new_n11352_; 
wire u2__abc_52155_new_n11353_; 
wire u2__abc_52155_new_n11354_; 
wire u2__abc_52155_new_n11355_; 
wire u2__abc_52155_new_n11356_; 
wire u2__abc_52155_new_n11357_; 
wire u2__abc_52155_new_n11359_; 
wire u2__abc_52155_new_n11360_; 
wire u2__abc_52155_new_n11361_; 
wire u2__abc_52155_new_n11362_; 
wire u2__abc_52155_new_n11363_; 
wire u2__abc_52155_new_n11364_; 
wire u2__abc_52155_new_n11365_; 
wire u2__abc_52155_new_n11366_; 
wire u2__abc_52155_new_n11367_; 
wire u2__abc_52155_new_n11368_; 
wire u2__abc_52155_new_n11369_; 
wire u2__abc_52155_new_n11370_; 
wire u2__abc_52155_new_n11371_; 
wire u2__abc_52155_new_n11372_; 
wire u2__abc_52155_new_n11373_; 
wire u2__abc_52155_new_n11374_; 
wire u2__abc_52155_new_n11375_; 
wire u2__abc_52155_new_n11376_; 
wire u2__abc_52155_new_n11378_; 
wire u2__abc_52155_new_n11379_; 
wire u2__abc_52155_new_n11380_; 
wire u2__abc_52155_new_n11381_; 
wire u2__abc_52155_new_n11382_; 
wire u2__abc_52155_new_n11383_; 
wire u2__abc_52155_new_n11384_; 
wire u2__abc_52155_new_n11385_; 
wire u2__abc_52155_new_n11386_; 
wire u2__abc_52155_new_n11387_; 
wire u2__abc_52155_new_n11388_; 
wire u2__abc_52155_new_n11389_; 
wire u2__abc_52155_new_n11390_; 
wire u2__abc_52155_new_n11391_; 
wire u2__abc_52155_new_n11392_; 
wire u2__abc_52155_new_n11393_; 
wire u2__abc_52155_new_n11395_; 
wire u2__abc_52155_new_n11396_; 
wire u2__abc_52155_new_n11397_; 
wire u2__abc_52155_new_n11398_; 
wire u2__abc_52155_new_n11399_; 
wire u2__abc_52155_new_n11400_; 
wire u2__abc_52155_new_n11401_; 
wire u2__abc_52155_new_n11402_; 
wire u2__abc_52155_new_n11403_; 
wire u2__abc_52155_new_n11404_; 
wire u2__abc_52155_new_n11405_; 
wire u2__abc_52155_new_n11406_; 
wire u2__abc_52155_new_n11407_; 
wire u2__abc_52155_new_n11408_; 
wire u2__abc_52155_new_n11409_; 
wire u2__abc_52155_new_n11410_; 
wire u2__abc_52155_new_n11411_; 
wire u2__abc_52155_new_n11412_; 
wire u2__abc_52155_new_n11413_; 
wire u2__abc_52155_new_n11414_; 
wire u2__abc_52155_new_n11415_; 
wire u2__abc_52155_new_n11416_; 
wire u2__abc_52155_new_n11417_; 
wire u2__abc_52155_new_n11418_; 
wire u2__abc_52155_new_n11419_; 
wire u2__abc_52155_new_n11420_; 
wire u2__abc_52155_new_n11421_; 
wire u2__abc_52155_new_n11422_; 
wire u2__abc_52155_new_n11423_; 
wire u2__abc_52155_new_n11424_; 
wire u2__abc_52155_new_n11426_; 
wire u2__abc_52155_new_n11427_; 
wire u2__abc_52155_new_n11428_; 
wire u2__abc_52155_new_n11429_; 
wire u2__abc_52155_new_n11430_; 
wire u2__abc_52155_new_n11431_; 
wire u2__abc_52155_new_n11432_; 
wire u2__abc_52155_new_n11433_; 
wire u2__abc_52155_new_n11434_; 
wire u2__abc_52155_new_n11435_; 
wire u2__abc_52155_new_n11436_; 
wire u2__abc_52155_new_n11437_; 
wire u2__abc_52155_new_n11438_; 
wire u2__abc_52155_new_n11439_; 
wire u2__abc_52155_new_n11440_; 
wire u2__abc_52155_new_n11441_; 
wire u2__abc_52155_new_n11443_; 
wire u2__abc_52155_new_n11444_; 
wire u2__abc_52155_new_n11445_; 
wire u2__abc_52155_new_n11446_; 
wire u2__abc_52155_new_n11447_; 
wire u2__abc_52155_new_n11448_; 
wire u2__abc_52155_new_n11449_; 
wire u2__abc_52155_new_n11450_; 
wire u2__abc_52155_new_n11451_; 
wire u2__abc_52155_new_n11452_; 
wire u2__abc_52155_new_n11453_; 
wire u2__abc_52155_new_n11454_; 
wire u2__abc_52155_new_n11455_; 
wire u2__abc_52155_new_n11456_; 
wire u2__abc_52155_new_n11457_; 
wire u2__abc_52155_new_n11458_; 
wire u2__abc_52155_new_n11459_; 
wire u2__abc_52155_new_n11461_; 
wire u2__abc_52155_new_n11462_; 
wire u2__abc_52155_new_n11463_; 
wire u2__abc_52155_new_n11464_; 
wire u2__abc_52155_new_n11465_; 
wire u2__abc_52155_new_n11466_; 
wire u2__abc_52155_new_n11467_; 
wire u2__abc_52155_new_n11468_; 
wire u2__abc_52155_new_n11469_; 
wire u2__abc_52155_new_n11470_; 
wire u2__abc_52155_new_n11471_; 
wire u2__abc_52155_new_n11472_; 
wire u2__abc_52155_new_n11473_; 
wire u2__abc_52155_new_n11474_; 
wire u2__abc_52155_new_n11475_; 
wire u2__abc_52155_new_n11476_; 
wire u2__abc_52155_new_n11477_; 
wire u2__abc_52155_new_n11479_; 
wire u2__abc_52155_new_n11480_; 
wire u2__abc_52155_new_n11481_; 
wire u2__abc_52155_new_n11482_; 
wire u2__abc_52155_new_n11483_; 
wire u2__abc_52155_new_n11484_; 
wire u2__abc_52155_new_n11485_; 
wire u2__abc_52155_new_n11486_; 
wire u2__abc_52155_new_n11487_; 
wire u2__abc_52155_new_n11488_; 
wire u2__abc_52155_new_n11489_; 
wire u2__abc_52155_new_n11490_; 
wire u2__abc_52155_new_n11491_; 
wire u2__abc_52155_new_n11492_; 
wire u2__abc_52155_new_n11493_; 
wire u2__abc_52155_new_n11494_; 
wire u2__abc_52155_new_n11495_; 
wire u2__abc_52155_new_n11496_; 
wire u2__abc_52155_new_n11497_; 
wire u2__abc_52155_new_n11498_; 
wire u2__abc_52155_new_n11499_; 
wire u2__abc_52155_new_n11500_; 
wire u2__abc_52155_new_n11501_; 
wire u2__abc_52155_new_n11503_; 
wire u2__abc_52155_new_n11504_; 
wire u2__abc_52155_new_n11505_; 
wire u2__abc_52155_new_n11506_; 
wire u2__abc_52155_new_n11507_; 
wire u2__abc_52155_new_n11508_; 
wire u2__abc_52155_new_n11509_; 
wire u2__abc_52155_new_n11510_; 
wire u2__abc_52155_new_n11511_; 
wire u2__abc_52155_new_n11512_; 
wire u2__abc_52155_new_n11513_; 
wire u2__abc_52155_new_n11514_; 
wire u2__abc_52155_new_n11515_; 
wire u2__abc_52155_new_n11516_; 
wire u2__abc_52155_new_n11517_; 
wire u2__abc_52155_new_n11518_; 
wire u2__abc_52155_new_n11520_; 
wire u2__abc_52155_new_n11521_; 
wire u2__abc_52155_new_n11522_; 
wire u2__abc_52155_new_n11523_; 
wire u2__abc_52155_new_n11524_; 
wire u2__abc_52155_new_n11525_; 
wire u2__abc_52155_new_n11526_; 
wire u2__abc_52155_new_n11527_; 
wire u2__abc_52155_new_n11528_; 
wire u2__abc_52155_new_n11529_; 
wire u2__abc_52155_new_n11530_; 
wire u2__abc_52155_new_n11531_; 
wire u2__abc_52155_new_n11532_; 
wire u2__abc_52155_new_n11533_; 
wire u2__abc_52155_new_n11534_; 
wire u2__abc_52155_new_n11535_; 
wire u2__abc_52155_new_n11537_; 
wire u2__abc_52155_new_n11538_; 
wire u2__abc_52155_new_n11539_; 
wire u2__abc_52155_new_n11540_; 
wire u2__abc_52155_new_n11541_; 
wire u2__abc_52155_new_n11542_; 
wire u2__abc_52155_new_n11543_; 
wire u2__abc_52155_new_n11544_; 
wire u2__abc_52155_new_n11545_; 
wire u2__abc_52155_new_n11546_; 
wire u2__abc_52155_new_n11547_; 
wire u2__abc_52155_new_n11548_; 
wire u2__abc_52155_new_n11549_; 
wire u2__abc_52155_new_n11550_; 
wire u2__abc_52155_new_n11551_; 
wire u2__abc_52155_new_n11552_; 
wire u2__abc_52155_new_n11554_; 
wire u2__abc_52155_new_n11555_; 
wire u2__abc_52155_new_n11556_; 
wire u2__abc_52155_new_n11557_; 
wire u2__abc_52155_new_n11558_; 
wire u2__abc_52155_new_n11559_; 
wire u2__abc_52155_new_n11560_; 
wire u2__abc_52155_new_n11561_; 
wire u2__abc_52155_new_n11562_; 
wire u2__abc_52155_new_n11563_; 
wire u2__abc_52155_new_n11564_; 
wire u2__abc_52155_new_n11565_; 
wire u2__abc_52155_new_n11566_; 
wire u2__abc_52155_new_n11567_; 
wire u2__abc_52155_new_n11568_; 
wire u2__abc_52155_new_n11569_; 
wire u2__abc_52155_new_n11570_; 
wire u2__abc_52155_new_n11571_; 
wire u2__abc_52155_new_n11572_; 
wire u2__abc_52155_new_n11573_; 
wire u2__abc_52155_new_n11574_; 
wire u2__abc_52155_new_n11575_; 
wire u2__abc_52155_new_n11576_; 
wire u2__abc_52155_new_n11577_; 
wire u2__abc_52155_new_n11579_; 
wire u2__abc_52155_new_n11580_; 
wire u2__abc_52155_new_n11581_; 
wire u2__abc_52155_new_n11582_; 
wire u2__abc_52155_new_n11583_; 
wire u2__abc_52155_new_n11584_; 
wire u2__abc_52155_new_n11585_; 
wire u2__abc_52155_new_n11586_; 
wire u2__abc_52155_new_n11587_; 
wire u2__abc_52155_new_n11588_; 
wire u2__abc_52155_new_n11589_; 
wire u2__abc_52155_new_n11590_; 
wire u2__abc_52155_new_n11591_; 
wire u2__abc_52155_new_n11592_; 
wire u2__abc_52155_new_n11593_; 
wire u2__abc_52155_new_n11594_; 
wire u2__abc_52155_new_n11596_; 
wire u2__abc_52155_new_n11597_; 
wire u2__abc_52155_new_n11598_; 
wire u2__abc_52155_new_n11599_; 
wire u2__abc_52155_new_n11600_; 
wire u2__abc_52155_new_n11601_; 
wire u2__abc_52155_new_n11602_; 
wire u2__abc_52155_new_n11603_; 
wire u2__abc_52155_new_n11604_; 
wire u2__abc_52155_new_n11605_; 
wire u2__abc_52155_new_n11606_; 
wire u2__abc_52155_new_n11607_; 
wire u2__abc_52155_new_n11608_; 
wire u2__abc_52155_new_n11609_; 
wire u2__abc_52155_new_n11610_; 
wire u2__abc_52155_new_n11611_; 
wire u2__abc_52155_new_n11612_; 
wire u2__abc_52155_new_n11613_; 
wire u2__abc_52155_new_n11615_; 
wire u2__abc_52155_new_n11616_; 
wire u2__abc_52155_new_n11617_; 
wire u2__abc_52155_new_n11618_; 
wire u2__abc_52155_new_n11619_; 
wire u2__abc_52155_new_n11620_; 
wire u2__abc_52155_new_n11621_; 
wire u2__abc_52155_new_n11622_; 
wire u2__abc_52155_new_n11623_; 
wire u2__abc_52155_new_n11624_; 
wire u2__abc_52155_new_n11625_; 
wire u2__abc_52155_new_n11626_; 
wire u2__abc_52155_new_n11627_; 
wire u2__abc_52155_new_n11628_; 
wire u2__abc_52155_new_n11629_; 
wire u2__abc_52155_new_n11630_; 
wire u2__abc_52155_new_n11632_; 
wire u2__abc_52155_new_n11633_; 
wire u2__abc_52155_new_n11634_; 
wire u2__abc_52155_new_n11635_; 
wire u2__abc_52155_new_n11636_; 
wire u2__abc_52155_new_n11637_; 
wire u2__abc_52155_new_n11638_; 
wire u2__abc_52155_new_n11639_; 
wire u2__abc_52155_new_n11640_; 
wire u2__abc_52155_new_n11641_; 
wire u2__abc_52155_new_n11642_; 
wire u2__abc_52155_new_n11643_; 
wire u2__abc_52155_new_n11644_; 
wire u2__abc_52155_new_n11645_; 
wire u2__abc_52155_new_n11646_; 
wire u2__abc_52155_new_n11647_; 
wire u2__abc_52155_new_n11648_; 
wire u2__abc_52155_new_n11649_; 
wire u2__abc_52155_new_n11650_; 
wire u2__abc_52155_new_n11651_; 
wire u2__abc_52155_new_n11652_; 
wire u2__abc_52155_new_n11653_; 
wire u2__abc_52155_new_n11655_; 
wire u2__abc_52155_new_n11656_; 
wire u2__abc_52155_new_n11657_; 
wire u2__abc_52155_new_n11658_; 
wire u2__abc_52155_new_n11659_; 
wire u2__abc_52155_new_n11660_; 
wire u2__abc_52155_new_n11661_; 
wire u2__abc_52155_new_n11662_; 
wire u2__abc_52155_new_n11663_; 
wire u2__abc_52155_new_n11664_; 
wire u2__abc_52155_new_n11665_; 
wire u2__abc_52155_new_n11666_; 
wire u2__abc_52155_new_n11667_; 
wire u2__abc_52155_new_n11668_; 
wire u2__abc_52155_new_n11669_; 
wire u2__abc_52155_new_n11670_; 
wire u2__abc_52155_new_n11672_; 
wire u2__abc_52155_new_n11673_; 
wire u2__abc_52155_new_n11674_; 
wire u2__abc_52155_new_n11675_; 
wire u2__abc_52155_new_n11676_; 
wire u2__abc_52155_new_n11677_; 
wire u2__abc_52155_new_n11678_; 
wire u2__abc_52155_new_n11679_; 
wire u2__abc_52155_new_n11680_; 
wire u2__abc_52155_new_n11681_; 
wire u2__abc_52155_new_n11682_; 
wire u2__abc_52155_new_n11683_; 
wire u2__abc_52155_new_n11684_; 
wire u2__abc_52155_new_n11685_; 
wire u2__abc_52155_new_n11686_; 
wire u2__abc_52155_new_n11687_; 
wire u2__abc_52155_new_n11688_; 
wire u2__abc_52155_new_n11689_; 
wire u2__abc_52155_new_n11691_; 
wire u2__abc_52155_new_n11692_; 
wire u2__abc_52155_new_n11693_; 
wire u2__abc_52155_new_n11694_; 
wire u2__abc_52155_new_n11695_; 
wire u2__abc_52155_new_n11696_; 
wire u2__abc_52155_new_n11697_; 
wire u2__abc_52155_new_n11698_; 
wire u2__abc_52155_new_n11699_; 
wire u2__abc_52155_new_n11700_; 
wire u2__abc_52155_new_n11701_; 
wire u2__abc_52155_new_n11702_; 
wire u2__abc_52155_new_n11703_; 
wire u2__abc_52155_new_n11704_; 
wire u2__abc_52155_new_n11705_; 
wire u2__abc_52155_new_n11706_; 
wire u2__abc_52155_new_n11708_; 
wire u2__abc_52155_new_n11709_; 
wire u2__abc_52155_new_n11710_; 
wire u2__abc_52155_new_n11711_; 
wire u2__abc_52155_new_n11712_; 
wire u2__abc_52155_new_n11713_; 
wire u2__abc_52155_new_n11714_; 
wire u2__abc_52155_new_n11715_; 
wire u2__abc_52155_new_n11716_; 
wire u2__abc_52155_new_n11717_; 
wire u2__abc_52155_new_n11718_; 
wire u2__abc_52155_new_n11719_; 
wire u2__abc_52155_new_n11720_; 
wire u2__abc_52155_new_n11721_; 
wire u2__abc_52155_new_n11722_; 
wire u2__abc_52155_new_n11723_; 
wire u2__abc_52155_new_n11724_; 
wire u2__abc_52155_new_n11725_; 
wire u2__abc_52155_new_n11726_; 
wire u2__abc_52155_new_n11727_; 
wire u2__abc_52155_new_n11728_; 
wire u2__abc_52155_new_n11729_; 
wire u2__abc_52155_new_n11730_; 
wire u2__abc_52155_new_n11731_; 
wire u2__abc_52155_new_n11732_; 
wire u2__abc_52155_new_n11733_; 
wire u2__abc_52155_new_n11735_; 
wire u2__abc_52155_new_n11736_; 
wire u2__abc_52155_new_n11737_; 
wire u2__abc_52155_new_n11738_; 
wire u2__abc_52155_new_n11739_; 
wire u2__abc_52155_new_n11740_; 
wire u2__abc_52155_new_n11741_; 
wire u2__abc_52155_new_n11742_; 
wire u2__abc_52155_new_n11743_; 
wire u2__abc_52155_new_n11744_; 
wire u2__abc_52155_new_n11745_; 
wire u2__abc_52155_new_n11746_; 
wire u2__abc_52155_new_n11747_; 
wire u2__abc_52155_new_n11748_; 
wire u2__abc_52155_new_n11749_; 
wire u2__abc_52155_new_n11750_; 
wire u2__abc_52155_new_n11752_; 
wire u2__abc_52155_new_n11753_; 
wire u2__abc_52155_new_n11754_; 
wire u2__abc_52155_new_n11755_; 
wire u2__abc_52155_new_n11756_; 
wire u2__abc_52155_new_n11757_; 
wire u2__abc_52155_new_n11758_; 
wire u2__abc_52155_new_n11759_; 
wire u2__abc_52155_new_n11760_; 
wire u2__abc_52155_new_n11761_; 
wire u2__abc_52155_new_n11762_; 
wire u2__abc_52155_new_n11763_; 
wire u2__abc_52155_new_n11764_; 
wire u2__abc_52155_new_n11765_; 
wire u2__abc_52155_new_n11766_; 
wire u2__abc_52155_new_n11767_; 
wire u2__abc_52155_new_n11768_; 
wire u2__abc_52155_new_n11769_; 
wire u2__abc_52155_new_n11770_; 
wire u2__abc_52155_new_n11772_; 
wire u2__abc_52155_new_n11773_; 
wire u2__abc_52155_new_n11774_; 
wire u2__abc_52155_new_n11775_; 
wire u2__abc_52155_new_n11776_; 
wire u2__abc_52155_new_n11777_; 
wire u2__abc_52155_new_n11778_; 
wire u2__abc_52155_new_n11779_; 
wire u2__abc_52155_new_n11780_; 
wire u2__abc_52155_new_n11781_; 
wire u2__abc_52155_new_n11782_; 
wire u2__abc_52155_new_n11783_; 
wire u2__abc_52155_new_n11784_; 
wire u2__abc_52155_new_n11785_; 
wire u2__abc_52155_new_n11786_; 
wire u2__abc_52155_new_n11787_; 
wire u2__abc_52155_new_n11789_; 
wire u2__abc_52155_new_n11790_; 
wire u2__abc_52155_new_n11791_; 
wire u2__abc_52155_new_n11792_; 
wire u2__abc_52155_new_n11793_; 
wire u2__abc_52155_new_n11794_; 
wire u2__abc_52155_new_n11795_; 
wire u2__abc_52155_new_n11796_; 
wire u2__abc_52155_new_n11797_; 
wire u2__abc_52155_new_n11798_; 
wire u2__abc_52155_new_n11799_; 
wire u2__abc_52155_new_n11800_; 
wire u2__abc_52155_new_n11801_; 
wire u2__abc_52155_new_n11802_; 
wire u2__abc_52155_new_n11803_; 
wire u2__abc_52155_new_n11804_; 
wire u2__abc_52155_new_n11805_; 
wire u2__abc_52155_new_n11806_; 
wire u2__abc_52155_new_n11807_; 
wire u2__abc_52155_new_n11808_; 
wire u2__abc_52155_new_n11810_; 
wire u2__abc_52155_new_n11811_; 
wire u2__abc_52155_new_n11812_; 
wire u2__abc_52155_new_n11813_; 
wire u2__abc_52155_new_n11814_; 
wire u2__abc_52155_new_n11815_; 
wire u2__abc_52155_new_n11816_; 
wire u2__abc_52155_new_n11817_; 
wire u2__abc_52155_new_n11818_; 
wire u2__abc_52155_new_n11819_; 
wire u2__abc_52155_new_n11820_; 
wire u2__abc_52155_new_n11821_; 
wire u2__abc_52155_new_n11822_; 
wire u2__abc_52155_new_n11823_; 
wire u2__abc_52155_new_n11824_; 
wire u2__abc_52155_new_n11825_; 
wire u2__abc_52155_new_n11827_; 
wire u2__abc_52155_new_n11828_; 
wire u2__abc_52155_new_n11829_; 
wire u2__abc_52155_new_n11830_; 
wire u2__abc_52155_new_n11831_; 
wire u2__abc_52155_new_n11832_; 
wire u2__abc_52155_new_n11833_; 
wire u2__abc_52155_new_n11834_; 
wire u2__abc_52155_new_n11835_; 
wire u2__abc_52155_new_n11836_; 
wire u2__abc_52155_new_n11837_; 
wire u2__abc_52155_new_n11838_; 
wire u2__abc_52155_new_n11839_; 
wire u2__abc_52155_new_n11840_; 
wire u2__abc_52155_new_n11841_; 
wire u2__abc_52155_new_n11842_; 
wire u2__abc_52155_new_n11844_; 
wire u2__abc_52155_new_n11845_; 
wire u2__abc_52155_new_n11846_; 
wire u2__abc_52155_new_n11847_; 
wire u2__abc_52155_new_n11848_; 
wire u2__abc_52155_new_n11849_; 
wire u2__abc_52155_new_n11850_; 
wire u2__abc_52155_new_n11851_; 
wire u2__abc_52155_new_n11852_; 
wire u2__abc_52155_new_n11853_; 
wire u2__abc_52155_new_n11854_; 
wire u2__abc_52155_new_n11855_; 
wire u2__abc_52155_new_n11856_; 
wire u2__abc_52155_new_n11857_; 
wire u2__abc_52155_new_n11858_; 
wire u2__abc_52155_new_n11859_; 
wire u2__abc_52155_new_n11861_; 
wire u2__abc_52155_new_n11862_; 
wire u2__abc_52155_new_n11863_; 
wire u2__abc_52155_new_n11864_; 
wire u2__abc_52155_new_n11865_; 
wire u2__abc_52155_new_n11866_; 
wire u2__abc_52155_new_n11867_; 
wire u2__abc_52155_new_n11868_; 
wire u2__abc_52155_new_n11869_; 
wire u2__abc_52155_new_n11870_; 
wire u2__abc_52155_new_n11871_; 
wire u2__abc_52155_new_n11872_; 
wire u2__abc_52155_new_n11873_; 
wire u2__abc_52155_new_n11874_; 
wire u2__abc_52155_new_n11875_; 
wire u2__abc_52155_new_n11876_; 
wire u2__abc_52155_new_n11877_; 
wire u2__abc_52155_new_n11878_; 
wire u2__abc_52155_new_n11879_; 
wire u2__abc_52155_new_n11880_; 
wire u2__abc_52155_new_n11881_; 
wire u2__abc_52155_new_n11882_; 
wire u2__abc_52155_new_n11883_; 
wire u2__abc_52155_new_n11884_; 
wire u2__abc_52155_new_n11886_; 
wire u2__abc_52155_new_n11887_; 
wire u2__abc_52155_new_n11888_; 
wire u2__abc_52155_new_n11889_; 
wire u2__abc_52155_new_n11890_; 
wire u2__abc_52155_new_n11891_; 
wire u2__abc_52155_new_n11892_; 
wire u2__abc_52155_new_n11893_; 
wire u2__abc_52155_new_n11894_; 
wire u2__abc_52155_new_n11895_; 
wire u2__abc_52155_new_n11896_; 
wire u2__abc_52155_new_n11897_; 
wire u2__abc_52155_new_n11898_; 
wire u2__abc_52155_new_n11899_; 
wire u2__abc_52155_new_n11900_; 
wire u2__abc_52155_new_n11901_; 
wire u2__abc_52155_new_n11903_; 
wire u2__abc_52155_new_n11904_; 
wire u2__abc_52155_new_n11905_; 
wire u2__abc_52155_new_n11906_; 
wire u2__abc_52155_new_n11907_; 
wire u2__abc_52155_new_n11908_; 
wire u2__abc_52155_new_n11909_; 
wire u2__abc_52155_new_n11910_; 
wire u2__abc_52155_new_n11911_; 
wire u2__abc_52155_new_n11912_; 
wire u2__abc_52155_new_n11913_; 
wire u2__abc_52155_new_n11914_; 
wire u2__abc_52155_new_n11915_; 
wire u2__abc_52155_new_n11916_; 
wire u2__abc_52155_new_n11917_; 
wire u2__abc_52155_new_n11918_; 
wire u2__abc_52155_new_n11919_; 
wire u2__abc_52155_new_n11920_; 
wire u2__abc_52155_new_n11921_; 
wire u2__abc_52155_new_n11923_; 
wire u2__abc_52155_new_n11924_; 
wire u2__abc_52155_new_n11925_; 
wire u2__abc_52155_new_n11926_; 
wire u2__abc_52155_new_n11927_; 
wire u2__abc_52155_new_n11928_; 
wire u2__abc_52155_new_n11929_; 
wire u2__abc_52155_new_n11930_; 
wire u2__abc_52155_new_n11931_; 
wire u2__abc_52155_new_n11932_; 
wire u2__abc_52155_new_n11933_; 
wire u2__abc_52155_new_n11934_; 
wire u2__abc_52155_new_n11935_; 
wire u2__abc_52155_new_n11936_; 
wire u2__abc_52155_new_n11937_; 
wire u2__abc_52155_new_n11938_; 
wire u2__abc_52155_new_n11940_; 
wire u2__abc_52155_new_n11941_; 
wire u2__abc_52155_new_n11942_; 
wire u2__abc_52155_new_n11943_; 
wire u2__abc_52155_new_n11944_; 
wire u2__abc_52155_new_n11945_; 
wire u2__abc_52155_new_n11946_; 
wire u2__abc_52155_new_n11947_; 
wire u2__abc_52155_new_n11948_; 
wire u2__abc_52155_new_n11949_; 
wire u2__abc_52155_new_n11950_; 
wire u2__abc_52155_new_n11951_; 
wire u2__abc_52155_new_n11952_; 
wire u2__abc_52155_new_n11953_; 
wire u2__abc_52155_new_n11954_; 
wire u2__abc_52155_new_n11955_; 
wire u2__abc_52155_new_n11956_; 
wire u2__abc_52155_new_n11957_; 
wire u2__abc_52155_new_n11958_; 
wire u2__abc_52155_new_n11959_; 
wire u2__abc_52155_new_n11961_; 
wire u2__abc_52155_new_n11962_; 
wire u2__abc_52155_new_n11963_; 
wire u2__abc_52155_new_n11964_; 
wire u2__abc_52155_new_n11965_; 
wire u2__abc_52155_new_n11966_; 
wire u2__abc_52155_new_n11967_; 
wire u2__abc_52155_new_n11968_; 
wire u2__abc_52155_new_n11969_; 
wire u2__abc_52155_new_n11970_; 
wire u2__abc_52155_new_n11971_; 
wire u2__abc_52155_new_n11972_; 
wire u2__abc_52155_new_n11973_; 
wire u2__abc_52155_new_n11974_; 
wire u2__abc_52155_new_n11975_; 
wire u2__abc_52155_new_n11976_; 
wire u2__abc_52155_new_n11978_; 
wire u2__abc_52155_new_n11979_; 
wire u2__abc_52155_new_n11980_; 
wire u2__abc_52155_new_n11981_; 
wire u2__abc_52155_new_n11982_; 
wire u2__abc_52155_new_n11983_; 
wire u2__abc_52155_new_n11984_; 
wire u2__abc_52155_new_n11985_; 
wire u2__abc_52155_new_n11986_; 
wire u2__abc_52155_new_n11987_; 
wire u2__abc_52155_new_n11988_; 
wire u2__abc_52155_new_n11989_; 
wire u2__abc_52155_new_n11990_; 
wire u2__abc_52155_new_n11991_; 
wire u2__abc_52155_new_n11992_; 
wire u2__abc_52155_new_n11993_; 
wire u2__abc_52155_new_n11994_; 
wire u2__abc_52155_new_n11995_; 
wire u2__abc_52155_new_n11997_; 
wire u2__abc_52155_new_n11998_; 
wire u2__abc_52155_new_n11999_; 
wire u2__abc_52155_new_n12000_; 
wire u2__abc_52155_new_n12001_; 
wire u2__abc_52155_new_n12002_; 
wire u2__abc_52155_new_n12003_; 
wire u2__abc_52155_new_n12004_; 
wire u2__abc_52155_new_n12005_; 
wire u2__abc_52155_new_n12006_; 
wire u2__abc_52155_new_n12007_; 
wire u2__abc_52155_new_n12008_; 
wire u2__abc_52155_new_n12009_; 
wire u2__abc_52155_new_n12010_; 
wire u2__abc_52155_new_n12011_; 
wire u2__abc_52155_new_n12012_; 
wire u2__abc_52155_new_n12014_; 
wire u2__abc_52155_new_n12015_; 
wire u2__abc_52155_new_n12016_; 
wire u2__abc_52155_new_n12017_; 
wire u2__abc_52155_new_n12018_; 
wire u2__abc_52155_new_n12019_; 
wire u2__abc_52155_new_n12020_; 
wire u2__abc_52155_new_n12021_; 
wire u2__abc_52155_new_n12022_; 
wire u2__abc_52155_new_n12023_; 
wire u2__abc_52155_new_n12024_; 
wire u2__abc_52155_new_n12025_; 
wire u2__abc_52155_new_n12026_; 
wire u2__abc_52155_new_n12027_; 
wire u2__abc_52155_new_n12028_; 
wire u2__abc_52155_new_n12029_; 
wire u2__abc_52155_new_n12030_; 
wire u2__abc_52155_new_n12031_; 
wire u2__abc_52155_new_n12032_; 
wire u2__abc_52155_new_n12033_; 
wire u2__abc_52155_new_n12034_; 
wire u2__abc_52155_new_n12035_; 
wire u2__abc_52155_new_n12036_; 
wire u2__abc_52155_new_n12037_; 
wire u2__abc_52155_new_n12038_; 
wire u2__abc_52155_new_n12039_; 
wire u2__abc_52155_new_n12040_; 
wire u2__abc_52155_new_n12041_; 
wire u2__abc_52155_new_n12042_; 
wire u2__abc_52155_new_n12043_; 
wire u2__abc_52155_new_n12044_; 
wire u2__abc_52155_new_n12045_; 
wire u2__abc_52155_new_n12046_; 
wire u2__abc_52155_new_n12048_; 
wire u2__abc_52155_new_n12049_; 
wire u2__abc_52155_new_n12050_; 
wire u2__abc_52155_new_n12051_; 
wire u2__abc_52155_new_n12052_; 
wire u2__abc_52155_new_n12053_; 
wire u2__abc_52155_new_n12054_; 
wire u2__abc_52155_new_n12055_; 
wire u2__abc_52155_new_n12056_; 
wire u2__abc_52155_new_n12057_; 
wire u2__abc_52155_new_n12058_; 
wire u2__abc_52155_new_n12059_; 
wire u2__abc_52155_new_n12060_; 
wire u2__abc_52155_new_n12061_; 
wire u2__abc_52155_new_n12062_; 
wire u2__abc_52155_new_n12063_; 
wire u2__abc_52155_new_n12065_; 
wire u2__abc_52155_new_n12066_; 
wire u2__abc_52155_new_n12067_; 
wire u2__abc_52155_new_n12068_; 
wire u2__abc_52155_new_n12069_; 
wire u2__abc_52155_new_n12070_; 
wire u2__abc_52155_new_n12071_; 
wire u2__abc_52155_new_n12072_; 
wire u2__abc_52155_new_n12073_; 
wire u2__abc_52155_new_n12074_; 
wire u2__abc_52155_new_n12075_; 
wire u2__abc_52155_new_n12076_; 
wire u2__abc_52155_new_n12077_; 
wire u2__abc_52155_new_n12078_; 
wire u2__abc_52155_new_n12079_; 
wire u2__abc_52155_new_n12080_; 
wire u2__abc_52155_new_n12081_; 
wire u2__abc_52155_new_n12082_; 
wire u2__abc_52155_new_n12084_; 
wire u2__abc_52155_new_n12085_; 
wire u2__abc_52155_new_n12086_; 
wire u2__abc_52155_new_n12087_; 
wire u2__abc_52155_new_n12088_; 
wire u2__abc_52155_new_n12089_; 
wire u2__abc_52155_new_n12090_; 
wire u2__abc_52155_new_n12091_; 
wire u2__abc_52155_new_n12092_; 
wire u2__abc_52155_new_n12093_; 
wire u2__abc_52155_new_n12094_; 
wire u2__abc_52155_new_n12095_; 
wire u2__abc_52155_new_n12096_; 
wire u2__abc_52155_new_n12097_; 
wire u2__abc_52155_new_n12098_; 
wire u2__abc_52155_new_n12099_; 
wire u2__abc_52155_new_n12101_; 
wire u2__abc_52155_new_n12102_; 
wire u2__abc_52155_new_n12103_; 
wire u2__abc_52155_new_n12104_; 
wire u2__abc_52155_new_n12105_; 
wire u2__abc_52155_new_n12106_; 
wire u2__abc_52155_new_n12107_; 
wire u2__abc_52155_new_n12108_; 
wire u2__abc_52155_new_n12109_; 
wire u2__abc_52155_new_n12110_; 
wire u2__abc_52155_new_n12111_; 
wire u2__abc_52155_new_n12112_; 
wire u2__abc_52155_new_n12113_; 
wire u2__abc_52155_new_n12114_; 
wire u2__abc_52155_new_n12115_; 
wire u2__abc_52155_new_n12116_; 
wire u2__abc_52155_new_n12117_; 
wire u2__abc_52155_new_n12118_; 
wire u2__abc_52155_new_n12119_; 
wire u2__abc_52155_new_n12120_; 
wire u2__abc_52155_new_n12121_; 
wire u2__abc_52155_new_n12122_; 
wire u2__abc_52155_new_n12123_; 
wire u2__abc_52155_new_n12124_; 
wire u2__abc_52155_new_n12126_; 
wire u2__abc_52155_new_n12127_; 
wire u2__abc_52155_new_n12128_; 
wire u2__abc_52155_new_n12129_; 
wire u2__abc_52155_new_n12130_; 
wire u2__abc_52155_new_n12131_; 
wire u2__abc_52155_new_n12132_; 
wire u2__abc_52155_new_n12133_; 
wire u2__abc_52155_new_n12134_; 
wire u2__abc_52155_new_n12135_; 
wire u2__abc_52155_new_n12136_; 
wire u2__abc_52155_new_n12137_; 
wire u2__abc_52155_new_n12138_; 
wire u2__abc_52155_new_n12139_; 
wire u2__abc_52155_new_n12140_; 
wire u2__abc_52155_new_n12141_; 
wire u2__abc_52155_new_n12143_; 
wire u2__abc_52155_new_n12144_; 
wire u2__abc_52155_new_n12145_; 
wire u2__abc_52155_new_n12146_; 
wire u2__abc_52155_new_n12147_; 
wire u2__abc_52155_new_n12148_; 
wire u2__abc_52155_new_n12149_; 
wire u2__abc_52155_new_n12150_; 
wire u2__abc_52155_new_n12151_; 
wire u2__abc_52155_new_n12152_; 
wire u2__abc_52155_new_n12153_; 
wire u2__abc_52155_new_n12154_; 
wire u2__abc_52155_new_n12155_; 
wire u2__abc_52155_new_n12156_; 
wire u2__abc_52155_new_n12157_; 
wire u2__abc_52155_new_n12158_; 
wire u2__abc_52155_new_n12159_; 
wire u2__abc_52155_new_n12160_; 
wire u2__abc_52155_new_n12162_; 
wire u2__abc_52155_new_n12163_; 
wire u2__abc_52155_new_n12164_; 
wire u2__abc_52155_new_n12165_; 
wire u2__abc_52155_new_n12166_; 
wire u2__abc_52155_new_n12167_; 
wire u2__abc_52155_new_n12168_; 
wire u2__abc_52155_new_n12169_; 
wire u2__abc_52155_new_n12170_; 
wire u2__abc_52155_new_n12171_; 
wire u2__abc_52155_new_n12172_; 
wire u2__abc_52155_new_n12173_; 
wire u2__abc_52155_new_n12174_; 
wire u2__abc_52155_new_n12175_; 
wire u2__abc_52155_new_n12176_; 
wire u2__abc_52155_new_n12177_; 
wire u2__abc_52155_new_n12179_; 
wire u2__abc_52155_new_n12180_; 
wire u2__abc_52155_new_n12181_; 
wire u2__abc_52155_new_n12182_; 
wire u2__abc_52155_new_n12183_; 
wire u2__abc_52155_new_n12184_; 
wire u2__abc_52155_new_n12185_; 
wire u2__abc_52155_new_n12186_; 
wire u2__abc_52155_new_n12187_; 
wire u2__abc_52155_new_n12188_; 
wire u2__abc_52155_new_n12189_; 
wire u2__abc_52155_new_n12190_; 
wire u2__abc_52155_new_n12191_; 
wire u2__abc_52155_new_n12192_; 
wire u2__abc_52155_new_n12193_; 
wire u2__abc_52155_new_n12194_; 
wire u2__abc_52155_new_n12195_; 
wire u2__abc_52155_new_n12196_; 
wire u2__abc_52155_new_n12197_; 
wire u2__abc_52155_new_n12198_; 
wire u2__abc_52155_new_n12199_; 
wire u2__abc_52155_new_n12200_; 
wire u2__abc_52155_new_n12201_; 
wire u2__abc_52155_new_n12202_; 
wire u2__abc_52155_new_n12204_; 
wire u2__abc_52155_new_n12205_; 
wire u2__abc_52155_new_n12206_; 
wire u2__abc_52155_new_n12207_; 
wire u2__abc_52155_new_n12208_; 
wire u2__abc_52155_new_n12209_; 
wire u2__abc_52155_new_n12210_; 
wire u2__abc_52155_new_n12211_; 
wire u2__abc_52155_new_n12212_; 
wire u2__abc_52155_new_n12213_; 
wire u2__abc_52155_new_n12214_; 
wire u2__abc_52155_new_n12215_; 
wire u2__abc_52155_new_n12216_; 
wire u2__abc_52155_new_n12217_; 
wire u2__abc_52155_new_n12218_; 
wire u2__abc_52155_new_n12219_; 
wire u2__abc_52155_new_n12221_; 
wire u2__abc_52155_new_n12222_; 
wire u2__abc_52155_new_n12223_; 
wire u2__abc_52155_new_n12224_; 
wire u2__abc_52155_new_n12225_; 
wire u2__abc_52155_new_n12226_; 
wire u2__abc_52155_new_n12227_; 
wire u2__abc_52155_new_n12228_; 
wire u2__abc_52155_new_n12229_; 
wire u2__abc_52155_new_n12230_; 
wire u2__abc_52155_new_n12231_; 
wire u2__abc_52155_new_n12232_; 
wire u2__abc_52155_new_n12233_; 
wire u2__abc_52155_new_n12234_; 
wire u2__abc_52155_new_n12235_; 
wire u2__abc_52155_new_n12236_; 
wire u2__abc_52155_new_n12237_; 
wire u2__abc_52155_new_n12238_; 
wire u2__abc_52155_new_n12239_; 
wire u2__abc_52155_new_n12241_; 
wire u2__abc_52155_new_n12242_; 
wire u2__abc_52155_new_n12243_; 
wire u2__abc_52155_new_n12244_; 
wire u2__abc_52155_new_n12245_; 
wire u2__abc_52155_new_n12246_; 
wire u2__abc_52155_new_n12247_; 
wire u2__abc_52155_new_n12248_; 
wire u2__abc_52155_new_n12249_; 
wire u2__abc_52155_new_n12250_; 
wire u2__abc_52155_new_n12251_; 
wire u2__abc_52155_new_n12252_; 
wire u2__abc_52155_new_n12253_; 
wire u2__abc_52155_new_n12254_; 
wire u2__abc_52155_new_n12255_; 
wire u2__abc_52155_new_n12256_; 
wire u2__abc_52155_new_n12258_; 
wire u2__abc_52155_new_n12259_; 
wire u2__abc_52155_new_n12260_; 
wire u2__abc_52155_new_n12261_; 
wire u2__abc_52155_new_n12262_; 
wire u2__abc_52155_new_n12263_; 
wire u2__abc_52155_new_n12264_; 
wire u2__abc_52155_new_n12265_; 
wire u2__abc_52155_new_n12266_; 
wire u2__abc_52155_new_n12267_; 
wire u2__abc_52155_new_n12268_; 
wire u2__abc_52155_new_n12269_; 
wire u2__abc_52155_new_n12270_; 
wire u2__abc_52155_new_n12271_; 
wire u2__abc_52155_new_n12272_; 
wire u2__abc_52155_new_n12273_; 
wire u2__abc_52155_new_n12274_; 
wire u2__abc_52155_new_n12275_; 
wire u2__abc_52155_new_n12277_; 
wire u2__abc_52155_new_n12278_; 
wire u2__abc_52155_new_n12279_; 
wire u2__abc_52155_new_n12280_; 
wire u2__abc_52155_new_n12281_; 
wire u2__abc_52155_new_n12282_; 
wire u2__abc_52155_new_n12283_; 
wire u2__abc_52155_new_n12284_; 
wire u2__abc_52155_new_n12285_; 
wire u2__abc_52155_new_n12286_; 
wire u2__abc_52155_new_n12287_; 
wire u2__abc_52155_new_n12288_; 
wire u2__abc_52155_new_n12289_; 
wire u2__abc_52155_new_n12290_; 
wire u2__abc_52155_new_n12291_; 
wire u2__abc_52155_new_n12292_; 
wire u2__abc_52155_new_n12294_; 
wire u2__abc_52155_new_n12295_; 
wire u2__abc_52155_new_n12296_; 
wire u2__abc_52155_new_n12297_; 
wire u2__abc_52155_new_n12298_; 
wire u2__abc_52155_new_n12299_; 
wire u2__abc_52155_new_n12300_; 
wire u2__abc_52155_new_n12301_; 
wire u2__abc_52155_new_n12302_; 
wire u2__abc_52155_new_n12303_; 
wire u2__abc_52155_new_n12304_; 
wire u2__abc_52155_new_n12305_; 
wire u2__abc_52155_new_n12306_; 
wire u2__abc_52155_new_n12307_; 
wire u2__abc_52155_new_n12308_; 
wire u2__abc_52155_new_n12309_; 
wire u2__abc_52155_new_n12310_; 
wire u2__abc_52155_new_n12311_; 
wire u2__abc_52155_new_n12313_; 
wire u2__abc_52155_new_n12314_; 
wire u2__abc_52155_new_n12315_; 
wire u2__abc_52155_new_n12316_; 
wire u2__abc_52155_new_n12317_; 
wire u2__abc_52155_new_n12318_; 
wire u2__abc_52155_new_n12319_; 
wire u2__abc_52155_new_n12320_; 
wire u2__abc_52155_new_n12321_; 
wire u2__abc_52155_new_n12322_; 
wire u2__abc_52155_new_n12323_; 
wire u2__abc_52155_new_n12324_; 
wire u2__abc_52155_new_n12325_; 
wire u2__abc_52155_new_n12326_; 
wire u2__abc_52155_new_n12327_; 
wire u2__abc_52155_new_n12328_; 
wire u2__abc_52155_new_n12330_; 
wire u2__abc_52155_new_n12331_; 
wire u2__abc_52155_new_n12332_; 
wire u2__abc_52155_new_n12333_; 
wire u2__abc_52155_new_n12334_; 
wire u2__abc_52155_new_n12335_; 
wire u2__abc_52155_new_n12336_; 
wire u2__abc_52155_new_n12337_; 
wire u2__abc_52155_new_n12338_; 
wire u2__abc_52155_new_n12339_; 
wire u2__abc_52155_new_n12340_; 
wire u2__abc_52155_new_n12341_; 
wire u2__abc_52155_new_n12342_; 
wire u2__abc_52155_new_n12343_; 
wire u2__abc_52155_new_n12344_; 
wire u2__abc_52155_new_n12345_; 
wire u2__abc_52155_new_n12346_; 
wire u2__abc_52155_new_n12347_; 
wire u2__abc_52155_new_n12348_; 
wire u2__abc_52155_new_n12349_; 
wire u2__abc_52155_new_n12350_; 
wire u2__abc_52155_new_n12351_; 
wire u2__abc_52155_new_n12352_; 
wire u2__abc_52155_new_n12353_; 
wire u2__abc_52155_new_n12354_; 
wire u2__abc_52155_new_n12355_; 
wire u2__abc_52155_new_n12356_; 
wire u2__abc_52155_new_n12357_; 
wire u2__abc_52155_new_n12358_; 
wire u2__abc_52155_new_n12359_; 
wire u2__abc_52155_new_n12360_; 
wire u2__abc_52155_new_n12361_; 
wire u2__abc_52155_new_n12362_; 
wire u2__abc_52155_new_n12363_; 
wire u2__abc_52155_new_n12364_; 
wire u2__abc_52155_new_n12366_; 
wire u2__abc_52155_new_n12367_; 
wire u2__abc_52155_new_n12368_; 
wire u2__abc_52155_new_n12369_; 
wire u2__abc_52155_new_n12370_; 
wire u2__abc_52155_new_n12371_; 
wire u2__abc_52155_new_n12372_; 
wire u2__abc_52155_new_n12373_; 
wire u2__abc_52155_new_n12374_; 
wire u2__abc_52155_new_n12375_; 
wire u2__abc_52155_new_n12376_; 
wire u2__abc_52155_new_n12377_; 
wire u2__abc_52155_new_n12378_; 
wire u2__abc_52155_new_n12379_; 
wire u2__abc_52155_new_n12380_; 
wire u2__abc_52155_new_n12381_; 
wire u2__abc_52155_new_n12383_; 
wire u2__abc_52155_new_n12384_; 
wire u2__abc_52155_new_n12385_; 
wire u2__abc_52155_new_n12386_; 
wire u2__abc_52155_new_n12387_; 
wire u2__abc_52155_new_n12388_; 
wire u2__abc_52155_new_n12389_; 
wire u2__abc_52155_new_n12390_; 
wire u2__abc_52155_new_n12391_; 
wire u2__abc_52155_new_n12392_; 
wire u2__abc_52155_new_n12393_; 
wire u2__abc_52155_new_n12394_; 
wire u2__abc_52155_new_n12395_; 
wire u2__abc_52155_new_n12396_; 
wire u2__abc_52155_new_n12397_; 
wire u2__abc_52155_new_n12398_; 
wire u2__abc_52155_new_n12399_; 
wire u2__abc_52155_new_n12400_; 
wire u2__abc_52155_new_n12401_; 
wire u2__abc_52155_new_n12403_; 
wire u2__abc_52155_new_n12404_; 
wire u2__abc_52155_new_n12405_; 
wire u2__abc_52155_new_n12406_; 
wire u2__abc_52155_new_n12407_; 
wire u2__abc_52155_new_n12408_; 
wire u2__abc_52155_new_n12409_; 
wire u2__abc_52155_new_n12410_; 
wire u2__abc_52155_new_n12411_; 
wire u2__abc_52155_new_n12412_; 
wire u2__abc_52155_new_n12413_; 
wire u2__abc_52155_new_n12414_; 
wire u2__abc_52155_new_n12415_; 
wire u2__abc_52155_new_n12416_; 
wire u2__abc_52155_new_n12417_; 
wire u2__abc_52155_new_n12418_; 
wire u2__abc_52155_new_n12420_; 
wire u2__abc_52155_new_n12421_; 
wire u2__abc_52155_new_n12422_; 
wire u2__abc_52155_new_n12423_; 
wire u2__abc_52155_new_n12424_; 
wire u2__abc_52155_new_n12425_; 
wire u2__abc_52155_new_n12426_; 
wire u2__abc_52155_new_n12427_; 
wire u2__abc_52155_new_n12428_; 
wire u2__abc_52155_new_n12429_; 
wire u2__abc_52155_new_n12430_; 
wire u2__abc_52155_new_n12431_; 
wire u2__abc_52155_new_n12432_; 
wire u2__abc_52155_new_n12433_; 
wire u2__abc_52155_new_n12434_; 
wire u2__abc_52155_new_n12435_; 
wire u2__abc_52155_new_n12436_; 
wire u2__abc_52155_new_n12437_; 
wire u2__abc_52155_new_n12438_; 
wire u2__abc_52155_new_n12439_; 
wire u2__abc_52155_new_n12441_; 
wire u2__abc_52155_new_n12442_; 
wire u2__abc_52155_new_n12443_; 
wire u2__abc_52155_new_n12444_; 
wire u2__abc_52155_new_n12445_; 
wire u2__abc_52155_new_n12446_; 
wire u2__abc_52155_new_n12447_; 
wire u2__abc_52155_new_n12448_; 
wire u2__abc_52155_new_n12449_; 
wire u2__abc_52155_new_n12450_; 
wire u2__abc_52155_new_n12451_; 
wire u2__abc_52155_new_n12452_; 
wire u2__abc_52155_new_n12453_; 
wire u2__abc_52155_new_n12454_; 
wire u2__abc_52155_new_n12455_; 
wire u2__abc_52155_new_n12456_; 
wire u2__abc_52155_new_n12458_; 
wire u2__abc_52155_new_n12459_; 
wire u2__abc_52155_new_n12460_; 
wire u2__abc_52155_new_n12461_; 
wire u2__abc_52155_new_n12462_; 
wire u2__abc_52155_new_n12463_; 
wire u2__abc_52155_new_n12464_; 
wire u2__abc_52155_new_n12465_; 
wire u2__abc_52155_new_n12466_; 
wire u2__abc_52155_new_n12467_; 
wire u2__abc_52155_new_n12468_; 
wire u2__abc_52155_new_n12469_; 
wire u2__abc_52155_new_n12470_; 
wire u2__abc_52155_new_n12471_; 
wire u2__abc_52155_new_n12472_; 
wire u2__abc_52155_new_n12473_; 
wire u2__abc_52155_new_n12475_; 
wire u2__abc_52155_new_n12476_; 
wire u2__abc_52155_new_n12477_; 
wire u2__abc_52155_new_n12478_; 
wire u2__abc_52155_new_n12479_; 
wire u2__abc_52155_new_n12480_; 
wire u2__abc_52155_new_n12481_; 
wire u2__abc_52155_new_n12482_; 
wire u2__abc_52155_new_n12483_; 
wire u2__abc_52155_new_n12484_; 
wire u2__abc_52155_new_n12485_; 
wire u2__abc_52155_new_n12486_; 
wire u2__abc_52155_new_n12487_; 
wire u2__abc_52155_new_n12488_; 
wire u2__abc_52155_new_n12489_; 
wire u2__abc_52155_new_n12490_; 
wire u2__abc_52155_new_n12492_; 
wire u2__abc_52155_new_n12493_; 
wire u2__abc_52155_new_n12494_; 
wire u2__abc_52155_new_n12495_; 
wire u2__abc_52155_new_n12496_; 
wire u2__abc_52155_new_n12497_; 
wire u2__abc_52155_new_n12498_; 
wire u2__abc_52155_new_n12499_; 
wire u2__abc_52155_new_n12500_; 
wire u2__abc_52155_new_n12501_; 
wire u2__abc_52155_new_n12502_; 
wire u2__abc_52155_new_n12503_; 
wire u2__abc_52155_new_n12504_; 
wire u2__abc_52155_new_n12505_; 
wire u2__abc_52155_new_n12506_; 
wire u2__abc_52155_new_n12507_; 
wire u2__abc_52155_new_n12508_; 
wire u2__abc_52155_new_n12509_; 
wire u2__abc_52155_new_n12510_; 
wire u2__abc_52155_new_n12511_; 
wire u2__abc_52155_new_n12512_; 
wire u2__abc_52155_new_n12513_; 
wire u2__abc_52155_new_n12514_; 
wire u2__abc_52155_new_n12515_; 
wire u2__abc_52155_new_n12517_; 
wire u2__abc_52155_new_n12518_; 
wire u2__abc_52155_new_n12519_; 
wire u2__abc_52155_new_n12520_; 
wire u2__abc_52155_new_n12521_; 
wire u2__abc_52155_new_n12522_; 
wire u2__abc_52155_new_n12523_; 
wire u2__abc_52155_new_n12524_; 
wire u2__abc_52155_new_n12525_; 
wire u2__abc_52155_new_n12526_; 
wire u2__abc_52155_new_n12527_; 
wire u2__abc_52155_new_n12528_; 
wire u2__abc_52155_new_n12529_; 
wire u2__abc_52155_new_n12530_; 
wire u2__abc_52155_new_n12531_; 
wire u2__abc_52155_new_n12532_; 
wire u2__abc_52155_new_n12534_; 
wire u2__abc_52155_new_n12535_; 
wire u2__abc_52155_new_n12536_; 
wire u2__abc_52155_new_n12537_; 
wire u2__abc_52155_new_n12538_; 
wire u2__abc_52155_new_n12539_; 
wire u2__abc_52155_new_n12540_; 
wire u2__abc_52155_new_n12541_; 
wire u2__abc_52155_new_n12542_; 
wire u2__abc_52155_new_n12543_; 
wire u2__abc_52155_new_n12544_; 
wire u2__abc_52155_new_n12545_; 
wire u2__abc_52155_new_n12546_; 
wire u2__abc_52155_new_n12547_; 
wire u2__abc_52155_new_n12548_; 
wire u2__abc_52155_new_n12549_; 
wire u2__abc_52155_new_n12550_; 
wire u2__abc_52155_new_n12551_; 
wire u2__abc_52155_new_n12552_; 
wire u2__abc_52155_new_n12554_; 
wire u2__abc_52155_new_n12555_; 
wire u2__abc_52155_new_n12556_; 
wire u2__abc_52155_new_n12557_; 
wire u2__abc_52155_new_n12558_; 
wire u2__abc_52155_new_n12559_; 
wire u2__abc_52155_new_n12560_; 
wire u2__abc_52155_new_n12561_; 
wire u2__abc_52155_new_n12562_; 
wire u2__abc_52155_new_n12563_; 
wire u2__abc_52155_new_n12564_; 
wire u2__abc_52155_new_n12565_; 
wire u2__abc_52155_new_n12566_; 
wire u2__abc_52155_new_n12567_; 
wire u2__abc_52155_new_n12568_; 
wire u2__abc_52155_new_n12569_; 
wire u2__abc_52155_new_n12571_; 
wire u2__abc_52155_new_n12572_; 
wire u2__abc_52155_new_n12573_; 
wire u2__abc_52155_new_n12574_; 
wire u2__abc_52155_new_n12575_; 
wire u2__abc_52155_new_n12576_; 
wire u2__abc_52155_new_n12577_; 
wire u2__abc_52155_new_n12578_; 
wire u2__abc_52155_new_n12579_; 
wire u2__abc_52155_new_n12580_; 
wire u2__abc_52155_new_n12581_; 
wire u2__abc_52155_new_n12582_; 
wire u2__abc_52155_new_n12583_; 
wire u2__abc_52155_new_n12584_; 
wire u2__abc_52155_new_n12585_; 
wire u2__abc_52155_new_n12586_; 
wire u2__abc_52155_new_n12587_; 
wire u2__abc_52155_new_n12588_; 
wire u2__abc_52155_new_n12589_; 
wire u2__abc_52155_new_n12590_; 
wire u2__abc_52155_new_n12592_; 
wire u2__abc_52155_new_n12593_; 
wire u2__abc_52155_new_n12594_; 
wire u2__abc_52155_new_n12595_; 
wire u2__abc_52155_new_n12596_; 
wire u2__abc_52155_new_n12597_; 
wire u2__abc_52155_new_n12598_; 
wire u2__abc_52155_new_n12599_; 
wire u2__abc_52155_new_n12600_; 
wire u2__abc_52155_new_n12601_; 
wire u2__abc_52155_new_n12602_; 
wire u2__abc_52155_new_n12603_; 
wire u2__abc_52155_new_n12604_; 
wire u2__abc_52155_new_n12605_; 
wire u2__abc_52155_new_n12606_; 
wire u2__abc_52155_new_n12607_; 
wire u2__abc_52155_new_n12609_; 
wire u2__abc_52155_new_n12610_; 
wire u2__abc_52155_new_n12611_; 
wire u2__abc_52155_new_n12612_; 
wire u2__abc_52155_new_n12613_; 
wire u2__abc_52155_new_n12614_; 
wire u2__abc_52155_new_n12615_; 
wire u2__abc_52155_new_n12616_; 
wire u2__abc_52155_new_n12617_; 
wire u2__abc_52155_new_n12618_; 
wire u2__abc_52155_new_n12619_; 
wire u2__abc_52155_new_n12620_; 
wire u2__abc_52155_new_n12621_; 
wire u2__abc_52155_new_n12622_; 
wire u2__abc_52155_new_n12623_; 
wire u2__abc_52155_new_n12624_; 
wire u2__abc_52155_new_n12625_; 
wire u2__abc_52155_new_n12626_; 
wire u2__abc_52155_new_n12628_; 
wire u2__abc_52155_new_n12629_; 
wire u2__abc_52155_new_n12630_; 
wire u2__abc_52155_new_n12631_; 
wire u2__abc_52155_new_n12632_; 
wire u2__abc_52155_new_n12633_; 
wire u2__abc_52155_new_n12634_; 
wire u2__abc_52155_new_n12635_; 
wire u2__abc_52155_new_n12636_; 
wire u2__abc_52155_new_n12637_; 
wire u2__abc_52155_new_n12638_; 
wire u2__abc_52155_new_n12639_; 
wire u2__abc_52155_new_n12640_; 
wire u2__abc_52155_new_n12641_; 
wire u2__abc_52155_new_n12642_; 
wire u2__abc_52155_new_n12643_; 
wire u2__abc_52155_new_n12645_; 
wire u2__abc_52155_new_n12646_; 
wire u2__abc_52155_new_n12647_; 
wire u2__abc_52155_new_n12648_; 
wire u2__abc_52155_new_n12649_; 
wire u2__abc_52155_new_n12650_; 
wire u2__abc_52155_new_n12651_; 
wire u2__abc_52155_new_n12652_; 
wire u2__abc_52155_new_n12653_; 
wire u2__abc_52155_new_n12654_; 
wire u2__abc_52155_new_n12655_; 
wire u2__abc_52155_new_n12656_; 
wire u2__abc_52155_new_n12657_; 
wire u2__abc_52155_new_n12658_; 
wire u2__abc_52155_new_n12659_; 
wire u2__abc_52155_new_n12660_; 
wire u2__abc_52155_new_n12661_; 
wire u2__abc_52155_new_n12662_; 
wire u2__abc_52155_new_n12663_; 
wire u2__abc_52155_new_n12664_; 
wire u2__abc_52155_new_n12665_; 
wire u2__abc_52155_new_n12666_; 
wire u2__abc_52155_new_n12667_; 
wire u2__abc_52155_new_n12668_; 
wire u2__abc_52155_new_n12669_; 
wire u2__abc_52155_new_n12670_; 
wire u2__abc_52155_new_n12671_; 
wire u2__abc_52155_new_n12672_; 
wire u2__abc_52155_new_n12673_; 
wire u2__abc_52155_new_n12674_; 
wire u2__abc_52155_new_n12675_; 
wire u2__abc_52155_new_n12676_; 
wire u2__abc_52155_new_n12678_; 
wire u2__abc_52155_new_n12679_; 
wire u2__abc_52155_new_n12680_; 
wire u2__abc_52155_new_n12681_; 
wire u2__abc_52155_new_n12682_; 
wire u2__abc_52155_new_n12683_; 
wire u2__abc_52155_new_n12684_; 
wire u2__abc_52155_new_n12685_; 
wire u2__abc_52155_new_n12686_; 
wire u2__abc_52155_new_n12687_; 
wire u2__abc_52155_new_n12688_; 
wire u2__abc_52155_new_n12689_; 
wire u2__abc_52155_new_n12690_; 
wire u2__abc_52155_new_n12691_; 
wire u2__abc_52155_new_n12692_; 
wire u2__abc_52155_new_n12693_; 
wire u2__abc_52155_new_n12695_; 
wire u2__abc_52155_new_n12696_; 
wire u2__abc_52155_new_n12697_; 
wire u2__abc_52155_new_n12698_; 
wire u2__abc_52155_new_n12699_; 
wire u2__abc_52155_new_n12700_; 
wire u2__abc_52155_new_n12701_; 
wire u2__abc_52155_new_n12702_; 
wire u2__abc_52155_new_n12703_; 
wire u2__abc_52155_new_n12704_; 
wire u2__abc_52155_new_n12705_; 
wire u2__abc_52155_new_n12706_; 
wire u2__abc_52155_new_n12707_; 
wire u2__abc_52155_new_n12708_; 
wire u2__abc_52155_new_n12709_; 
wire u2__abc_52155_new_n12710_; 
wire u2__abc_52155_new_n12711_; 
wire u2__abc_52155_new_n12712_; 
wire u2__abc_52155_new_n12713_; 
wire u2__abc_52155_new_n12715_; 
wire u2__abc_52155_new_n12716_; 
wire u2__abc_52155_new_n12717_; 
wire u2__abc_52155_new_n12718_; 
wire u2__abc_52155_new_n12719_; 
wire u2__abc_52155_new_n12720_; 
wire u2__abc_52155_new_n12721_; 
wire u2__abc_52155_new_n12722_; 
wire u2__abc_52155_new_n12723_; 
wire u2__abc_52155_new_n12724_; 
wire u2__abc_52155_new_n12725_; 
wire u2__abc_52155_new_n12726_; 
wire u2__abc_52155_new_n12727_; 
wire u2__abc_52155_new_n12728_; 
wire u2__abc_52155_new_n12729_; 
wire u2__abc_52155_new_n12730_; 
wire u2__abc_52155_new_n12732_; 
wire u2__abc_52155_new_n12733_; 
wire u2__abc_52155_new_n12734_; 
wire u2__abc_52155_new_n12735_; 
wire u2__abc_52155_new_n12736_; 
wire u2__abc_52155_new_n12737_; 
wire u2__abc_52155_new_n12738_; 
wire u2__abc_52155_new_n12739_; 
wire u2__abc_52155_new_n12740_; 
wire u2__abc_52155_new_n12741_; 
wire u2__abc_52155_new_n12742_; 
wire u2__abc_52155_new_n12743_; 
wire u2__abc_52155_new_n12744_; 
wire u2__abc_52155_new_n12745_; 
wire u2__abc_52155_new_n12746_; 
wire u2__abc_52155_new_n12747_; 
wire u2__abc_52155_new_n12748_; 
wire u2__abc_52155_new_n12749_; 
wire u2__abc_52155_new_n12750_; 
wire u2__abc_52155_new_n12751_; 
wire u2__abc_52155_new_n12753_; 
wire u2__abc_52155_new_n12754_; 
wire u2__abc_52155_new_n12755_; 
wire u2__abc_52155_new_n12756_; 
wire u2__abc_52155_new_n12757_; 
wire u2__abc_52155_new_n12758_; 
wire u2__abc_52155_new_n12759_; 
wire u2__abc_52155_new_n12760_; 
wire u2__abc_52155_new_n12761_; 
wire u2__abc_52155_new_n12762_; 
wire u2__abc_52155_new_n12763_; 
wire u2__abc_52155_new_n12764_; 
wire u2__abc_52155_new_n12765_; 
wire u2__abc_52155_new_n12766_; 
wire u2__abc_52155_new_n12767_; 
wire u2__abc_52155_new_n12768_; 
wire u2__abc_52155_new_n12770_; 
wire u2__abc_52155_new_n12771_; 
wire u2__abc_52155_new_n12772_; 
wire u2__abc_52155_new_n12773_; 
wire u2__abc_52155_new_n12774_; 
wire u2__abc_52155_new_n12775_; 
wire u2__abc_52155_new_n12776_; 
wire u2__abc_52155_new_n12777_; 
wire u2__abc_52155_new_n12778_; 
wire u2__abc_52155_new_n12779_; 
wire u2__abc_52155_new_n12780_; 
wire u2__abc_52155_new_n12781_; 
wire u2__abc_52155_new_n12782_; 
wire u2__abc_52155_new_n12783_; 
wire u2__abc_52155_new_n12784_; 
wire u2__abc_52155_new_n12785_; 
wire u2__abc_52155_new_n12786_; 
wire u2__abc_52155_new_n12787_; 
wire u2__abc_52155_new_n12789_; 
wire u2__abc_52155_new_n12790_; 
wire u2__abc_52155_new_n12791_; 
wire u2__abc_52155_new_n12792_; 
wire u2__abc_52155_new_n12793_; 
wire u2__abc_52155_new_n12794_; 
wire u2__abc_52155_new_n12795_; 
wire u2__abc_52155_new_n12796_; 
wire u2__abc_52155_new_n12797_; 
wire u2__abc_52155_new_n12798_; 
wire u2__abc_52155_new_n12799_; 
wire u2__abc_52155_new_n12800_; 
wire u2__abc_52155_new_n12801_; 
wire u2__abc_52155_new_n12802_; 
wire u2__abc_52155_new_n12803_; 
wire u2__abc_52155_new_n12804_; 
wire u2__abc_52155_new_n12806_; 
wire u2__abc_52155_new_n12807_; 
wire u2__abc_52155_new_n12808_; 
wire u2__abc_52155_new_n12809_; 
wire u2__abc_52155_new_n12810_; 
wire u2__abc_52155_new_n12811_; 
wire u2__abc_52155_new_n12812_; 
wire u2__abc_52155_new_n12813_; 
wire u2__abc_52155_new_n12814_; 
wire u2__abc_52155_new_n12815_; 
wire u2__abc_52155_new_n12816_; 
wire u2__abc_52155_new_n12817_; 
wire u2__abc_52155_new_n12818_; 
wire u2__abc_52155_new_n12819_; 
wire u2__abc_52155_new_n12820_; 
wire u2__abc_52155_new_n12821_; 
wire u2__abc_52155_new_n12822_; 
wire u2__abc_52155_new_n12823_; 
wire u2__abc_52155_new_n12824_; 
wire u2__abc_52155_new_n12825_; 
wire u2__abc_52155_new_n12826_; 
wire u2__abc_52155_new_n12827_; 
wire u2__abc_52155_new_n12828_; 
wire u2__abc_52155_new_n12829_; 
wire u2__abc_52155_new_n12830_; 
wire u2__abc_52155_new_n12831_; 
wire u2__abc_52155_new_n12833_; 
wire u2__abc_52155_new_n12834_; 
wire u2__abc_52155_new_n12835_; 
wire u2__abc_52155_new_n12836_; 
wire u2__abc_52155_new_n12837_; 
wire u2__abc_52155_new_n12838_; 
wire u2__abc_52155_new_n12839_; 
wire u2__abc_52155_new_n12840_; 
wire u2__abc_52155_new_n12841_; 
wire u2__abc_52155_new_n12842_; 
wire u2__abc_52155_new_n12843_; 
wire u2__abc_52155_new_n12844_; 
wire u2__abc_52155_new_n12845_; 
wire u2__abc_52155_new_n12846_; 
wire u2__abc_52155_new_n12847_; 
wire u2__abc_52155_new_n12848_; 
wire u2__abc_52155_new_n12850_; 
wire u2__abc_52155_new_n12851_; 
wire u2__abc_52155_new_n12852_; 
wire u2__abc_52155_new_n12853_; 
wire u2__abc_52155_new_n12854_; 
wire u2__abc_52155_new_n12855_; 
wire u2__abc_52155_new_n12856_; 
wire u2__abc_52155_new_n12857_; 
wire u2__abc_52155_new_n12858_; 
wire u2__abc_52155_new_n12859_; 
wire u2__abc_52155_new_n12860_; 
wire u2__abc_52155_new_n12861_; 
wire u2__abc_52155_new_n12862_; 
wire u2__abc_52155_new_n12863_; 
wire u2__abc_52155_new_n12864_; 
wire u2__abc_52155_new_n12865_; 
wire u2__abc_52155_new_n12866_; 
wire u2__abc_52155_new_n12867_; 
wire u2__abc_52155_new_n12868_; 
wire u2__abc_52155_new_n12870_; 
wire u2__abc_52155_new_n12871_; 
wire u2__abc_52155_new_n12872_; 
wire u2__abc_52155_new_n12873_; 
wire u2__abc_52155_new_n12874_; 
wire u2__abc_52155_new_n12875_; 
wire u2__abc_52155_new_n12876_; 
wire u2__abc_52155_new_n12877_; 
wire u2__abc_52155_new_n12878_; 
wire u2__abc_52155_new_n12879_; 
wire u2__abc_52155_new_n12880_; 
wire u2__abc_52155_new_n12881_; 
wire u2__abc_52155_new_n12882_; 
wire u2__abc_52155_new_n12883_; 
wire u2__abc_52155_new_n12884_; 
wire u2__abc_52155_new_n12885_; 
wire u2__abc_52155_new_n12887_; 
wire u2__abc_52155_new_n12888_; 
wire u2__abc_52155_new_n12889_; 
wire u2__abc_52155_new_n12890_; 
wire u2__abc_52155_new_n12891_; 
wire u2__abc_52155_new_n12892_; 
wire u2__abc_52155_new_n12893_; 
wire u2__abc_52155_new_n12894_; 
wire u2__abc_52155_new_n12895_; 
wire u2__abc_52155_new_n12896_; 
wire u2__abc_52155_new_n12897_; 
wire u2__abc_52155_new_n12898_; 
wire u2__abc_52155_new_n12899_; 
wire u2__abc_52155_new_n12900_; 
wire u2__abc_52155_new_n12901_; 
wire u2__abc_52155_new_n12902_; 
wire u2__abc_52155_new_n12903_; 
wire u2__abc_52155_new_n12904_; 
wire u2__abc_52155_new_n12906_; 
wire u2__abc_52155_new_n12907_; 
wire u2__abc_52155_new_n12908_; 
wire u2__abc_52155_new_n12909_; 
wire u2__abc_52155_new_n12910_; 
wire u2__abc_52155_new_n12911_; 
wire u2__abc_52155_new_n12912_; 
wire u2__abc_52155_new_n12913_; 
wire u2__abc_52155_new_n12914_; 
wire u2__abc_52155_new_n12915_; 
wire u2__abc_52155_new_n12916_; 
wire u2__abc_52155_new_n12917_; 
wire u2__abc_52155_new_n12918_; 
wire u2__abc_52155_new_n12919_; 
wire u2__abc_52155_new_n12920_; 
wire u2__abc_52155_new_n12921_; 
wire u2__abc_52155_new_n12923_; 
wire u2__abc_52155_new_n12924_; 
wire u2__abc_52155_new_n12925_; 
wire u2__abc_52155_new_n12926_; 
wire u2__abc_52155_new_n12927_; 
wire u2__abc_52155_new_n12928_; 
wire u2__abc_52155_new_n12929_; 
wire u2__abc_52155_new_n12930_; 
wire u2__abc_52155_new_n12931_; 
wire u2__abc_52155_new_n12932_; 
wire u2__abc_52155_new_n12933_; 
wire u2__abc_52155_new_n12934_; 
wire u2__abc_52155_new_n12935_; 
wire u2__abc_52155_new_n12936_; 
wire u2__abc_52155_new_n12937_; 
wire u2__abc_52155_new_n12938_; 
wire u2__abc_52155_new_n12939_; 
wire u2__abc_52155_new_n12940_; 
wire u2__abc_52155_new_n12942_; 
wire u2__abc_52155_new_n12943_; 
wire u2__abc_52155_new_n12944_; 
wire u2__abc_52155_new_n12945_; 
wire u2__abc_52155_new_n12946_; 
wire u2__abc_52155_new_n12947_; 
wire u2__abc_52155_new_n12948_; 
wire u2__abc_52155_new_n12949_; 
wire u2__abc_52155_new_n12950_; 
wire u2__abc_52155_new_n12951_; 
wire u2__abc_52155_new_n12952_; 
wire u2__abc_52155_new_n12953_; 
wire u2__abc_52155_new_n12954_; 
wire u2__abc_52155_new_n12955_; 
wire u2__abc_52155_new_n12956_; 
wire u2__abc_52155_new_n12957_; 
wire u2__abc_52155_new_n12959_; 
wire u2__abc_52155_new_n12960_; 
wire u2__abc_52155_new_n12961_; 
wire u2__abc_52155_new_n12962_; 
wire u2__abc_52155_new_n12963_; 
wire u2__abc_52155_new_n12964_; 
wire u2__abc_52155_new_n12965_; 
wire u2__abc_52155_new_n12966_; 
wire u2__abc_52155_new_n12967_; 
wire u2__abc_52155_new_n12968_; 
wire u2__abc_52155_new_n12969_; 
wire u2__abc_52155_new_n12970_; 
wire u2__abc_52155_new_n12971_; 
wire u2__abc_52155_new_n12972_; 
wire u2__abc_52155_new_n12973_; 
wire u2__abc_52155_new_n12974_; 
wire u2__abc_52155_new_n12975_; 
wire u2__abc_52155_new_n12976_; 
wire u2__abc_52155_new_n12977_; 
wire u2__abc_52155_new_n12978_; 
wire u2__abc_52155_new_n12979_; 
wire u2__abc_52155_new_n12980_; 
wire u2__abc_52155_new_n12981_; 
wire u2__abc_52155_new_n12982_; 
wire u2__abc_52155_new_n12983_; 
wire u2__abc_52155_new_n12984_; 
wire u2__abc_52155_new_n12985_; 
wire u2__abc_52155_new_n12986_; 
wire u2__abc_52155_new_n12987_; 
wire u2__abc_52155_new_n12988_; 
wire u2__abc_52155_new_n12989_; 
wire u2__abc_52155_new_n12991_; 
wire u2__abc_52155_new_n12992_; 
wire u2__abc_52155_new_n12993_; 
wire u2__abc_52155_new_n12994_; 
wire u2__abc_52155_new_n12995_; 
wire u2__abc_52155_new_n12996_; 
wire u2__abc_52155_new_n12997_; 
wire u2__abc_52155_new_n12998_; 
wire u2__abc_52155_new_n12999_; 
wire u2__abc_52155_new_n13000_; 
wire u2__abc_52155_new_n13001_; 
wire u2__abc_52155_new_n13002_; 
wire u2__abc_52155_new_n13003_; 
wire u2__abc_52155_new_n13004_; 
wire u2__abc_52155_new_n13005_; 
wire u2__abc_52155_new_n13006_; 
wire u2__abc_52155_new_n13008_; 
wire u2__abc_52155_new_n13009_; 
wire u2__abc_52155_new_n13010_; 
wire u2__abc_52155_new_n13011_; 
wire u2__abc_52155_new_n13012_; 
wire u2__abc_52155_new_n13013_; 
wire u2__abc_52155_new_n13014_; 
wire u2__abc_52155_new_n13015_; 
wire u2__abc_52155_new_n13016_; 
wire u2__abc_52155_new_n13017_; 
wire u2__abc_52155_new_n13018_; 
wire u2__abc_52155_new_n13019_; 
wire u2__abc_52155_new_n13020_; 
wire u2__abc_52155_new_n13021_; 
wire u2__abc_52155_new_n13022_; 
wire u2__abc_52155_new_n13023_; 
wire u2__abc_52155_new_n13024_; 
wire u2__abc_52155_new_n13025_; 
wire u2__abc_52155_new_n13027_; 
wire u2__abc_52155_new_n13028_; 
wire u2__abc_52155_new_n13029_; 
wire u2__abc_52155_new_n13030_; 
wire u2__abc_52155_new_n13031_; 
wire u2__abc_52155_new_n13032_; 
wire u2__abc_52155_new_n13033_; 
wire u2__abc_52155_new_n13034_; 
wire u2__abc_52155_new_n13035_; 
wire u2__abc_52155_new_n13036_; 
wire u2__abc_52155_new_n13037_; 
wire u2__abc_52155_new_n13038_; 
wire u2__abc_52155_new_n13039_; 
wire u2__abc_52155_new_n13040_; 
wire u2__abc_52155_new_n13041_; 
wire u2__abc_52155_new_n13042_; 
wire u2__abc_52155_new_n13044_; 
wire u2__abc_52155_new_n13045_; 
wire u2__abc_52155_new_n13046_; 
wire u2__abc_52155_new_n13047_; 
wire u2__abc_52155_new_n13048_; 
wire u2__abc_52155_new_n13049_; 
wire u2__abc_52155_new_n13050_; 
wire u2__abc_52155_new_n13051_; 
wire u2__abc_52155_new_n13052_; 
wire u2__abc_52155_new_n13053_; 
wire u2__abc_52155_new_n13054_; 
wire u2__abc_52155_new_n13055_; 
wire u2__abc_52155_new_n13056_; 
wire u2__abc_52155_new_n13057_; 
wire u2__abc_52155_new_n13058_; 
wire u2__abc_52155_new_n13059_; 
wire u2__abc_52155_new_n13060_; 
wire u2__abc_52155_new_n13061_; 
wire u2__abc_52155_new_n13062_; 
wire u2__abc_52155_new_n13063_; 
wire u2__abc_52155_new_n13064_; 
wire u2__abc_52155_new_n13065_; 
wire u2__abc_52155_new_n13066_; 
wire u2__abc_52155_new_n13068_; 
wire u2__abc_52155_new_n13069_; 
wire u2__abc_52155_new_n13070_; 
wire u2__abc_52155_new_n13071_; 
wire u2__abc_52155_new_n13072_; 
wire u2__abc_52155_new_n13073_; 
wire u2__abc_52155_new_n13074_; 
wire u2__abc_52155_new_n13075_; 
wire u2__abc_52155_new_n13076_; 
wire u2__abc_52155_new_n13077_; 
wire u2__abc_52155_new_n13078_; 
wire u2__abc_52155_new_n13079_; 
wire u2__abc_52155_new_n13080_; 
wire u2__abc_52155_new_n13081_; 
wire u2__abc_52155_new_n13082_; 
wire u2__abc_52155_new_n13083_; 
wire u2__abc_52155_new_n13085_; 
wire u2__abc_52155_new_n13086_; 
wire u2__abc_52155_new_n13087_; 
wire u2__abc_52155_new_n13088_; 
wire u2__abc_52155_new_n13089_; 
wire u2__abc_52155_new_n13090_; 
wire u2__abc_52155_new_n13091_; 
wire u2__abc_52155_new_n13092_; 
wire u2__abc_52155_new_n13093_; 
wire u2__abc_52155_new_n13094_; 
wire u2__abc_52155_new_n13095_; 
wire u2__abc_52155_new_n13096_; 
wire u2__abc_52155_new_n13097_; 
wire u2__abc_52155_new_n13098_; 
wire u2__abc_52155_new_n13099_; 
wire u2__abc_52155_new_n13100_; 
wire u2__abc_52155_new_n13101_; 
wire u2__abc_52155_new_n13102_; 
wire u2__abc_52155_new_n13104_; 
wire u2__abc_52155_new_n13105_; 
wire u2__abc_52155_new_n13106_; 
wire u2__abc_52155_new_n13107_; 
wire u2__abc_52155_new_n13108_; 
wire u2__abc_52155_new_n13109_; 
wire u2__abc_52155_new_n13110_; 
wire u2__abc_52155_new_n13111_; 
wire u2__abc_52155_new_n13112_; 
wire u2__abc_52155_new_n13113_; 
wire u2__abc_52155_new_n13114_; 
wire u2__abc_52155_new_n13115_; 
wire u2__abc_52155_new_n13116_; 
wire u2__abc_52155_new_n13117_; 
wire u2__abc_52155_new_n13118_; 
wire u2__abc_52155_new_n13119_; 
wire u2__abc_52155_new_n13121_; 
wire u2__abc_52155_new_n13122_; 
wire u2__abc_52155_new_n13123_; 
wire u2__abc_52155_new_n13124_; 
wire u2__abc_52155_new_n13125_; 
wire u2__abc_52155_new_n13126_; 
wire u2__abc_52155_new_n13127_; 
wire u2__abc_52155_new_n13128_; 
wire u2__abc_52155_new_n13129_; 
wire u2__abc_52155_new_n13130_; 
wire u2__abc_52155_new_n13131_; 
wire u2__abc_52155_new_n13132_; 
wire u2__abc_52155_new_n13133_; 
wire u2__abc_52155_new_n13134_; 
wire u2__abc_52155_new_n13135_; 
wire u2__abc_52155_new_n13136_; 
wire u2__abc_52155_new_n13137_; 
wire u2__abc_52155_new_n13138_; 
wire u2__abc_52155_new_n13139_; 
wire u2__abc_52155_new_n13140_; 
wire u2__abc_52155_new_n13141_; 
wire u2__abc_52155_new_n13142_; 
wire u2__abc_52155_new_n13143_; 
wire u2__abc_52155_new_n13144_; 
wire u2__abc_52155_new_n13145_; 
wire u2__abc_52155_new_n13147_; 
wire u2__abc_52155_new_n13148_; 
wire u2__abc_52155_new_n13149_; 
wire u2__abc_52155_new_n13150_; 
wire u2__abc_52155_new_n13151_; 
wire u2__abc_52155_new_n13152_; 
wire u2__abc_52155_new_n13153_; 
wire u2__abc_52155_new_n13154_; 
wire u2__abc_52155_new_n13155_; 
wire u2__abc_52155_new_n13156_; 
wire u2__abc_52155_new_n13157_; 
wire u2__abc_52155_new_n13158_; 
wire u2__abc_52155_new_n13159_; 
wire u2__abc_52155_new_n13160_; 
wire u2__abc_52155_new_n13161_; 
wire u2__abc_52155_new_n13162_; 
wire u2__abc_52155_new_n13164_; 
wire u2__abc_52155_new_n13165_; 
wire u2__abc_52155_new_n13166_; 
wire u2__abc_52155_new_n13167_; 
wire u2__abc_52155_new_n13168_; 
wire u2__abc_52155_new_n13169_; 
wire u2__abc_52155_new_n13170_; 
wire u2__abc_52155_new_n13171_; 
wire u2__abc_52155_new_n13172_; 
wire u2__abc_52155_new_n13173_; 
wire u2__abc_52155_new_n13174_; 
wire u2__abc_52155_new_n13175_; 
wire u2__abc_52155_new_n13176_; 
wire u2__abc_52155_new_n13177_; 
wire u2__abc_52155_new_n13178_; 
wire u2__abc_52155_new_n13179_; 
wire u2__abc_52155_new_n13180_; 
wire u2__abc_52155_new_n13181_; 
wire u2__abc_52155_new_n13183_; 
wire u2__abc_52155_new_n13184_; 
wire u2__abc_52155_new_n13185_; 
wire u2__abc_52155_new_n13186_; 
wire u2__abc_52155_new_n13187_; 
wire u2__abc_52155_new_n13188_; 
wire u2__abc_52155_new_n13189_; 
wire u2__abc_52155_new_n13190_; 
wire u2__abc_52155_new_n13191_; 
wire u2__abc_52155_new_n13192_; 
wire u2__abc_52155_new_n13193_; 
wire u2__abc_52155_new_n13194_; 
wire u2__abc_52155_new_n13195_; 
wire u2__abc_52155_new_n13196_; 
wire u2__abc_52155_new_n13197_; 
wire u2__abc_52155_new_n13198_; 
wire u2__abc_52155_new_n13200_; 
wire u2__abc_52155_new_n13201_; 
wire u2__abc_52155_new_n13202_; 
wire u2__abc_52155_new_n13203_; 
wire u2__abc_52155_new_n13204_; 
wire u2__abc_52155_new_n13205_; 
wire u2__abc_52155_new_n13206_; 
wire u2__abc_52155_new_n13207_; 
wire u2__abc_52155_new_n13208_; 
wire u2__abc_52155_new_n13209_; 
wire u2__abc_52155_new_n13210_; 
wire u2__abc_52155_new_n13211_; 
wire u2__abc_52155_new_n13212_; 
wire u2__abc_52155_new_n13213_; 
wire u2__abc_52155_new_n13214_; 
wire u2__abc_52155_new_n13215_; 
wire u2__abc_52155_new_n13216_; 
wire u2__abc_52155_new_n13217_; 
wire u2__abc_52155_new_n13218_; 
wire u2__abc_52155_new_n13219_; 
wire u2__abc_52155_new_n13220_; 
wire u2__abc_52155_new_n13221_; 
wire u2__abc_52155_new_n13222_; 
wire u2__abc_52155_new_n13224_; 
wire u2__abc_52155_new_n13225_; 
wire u2__abc_52155_new_n13226_; 
wire u2__abc_52155_new_n13227_; 
wire u2__abc_52155_new_n13228_; 
wire u2__abc_52155_new_n13229_; 
wire u2__abc_52155_new_n13230_; 
wire u2__abc_52155_new_n13231_; 
wire u2__abc_52155_new_n13232_; 
wire u2__abc_52155_new_n13233_; 
wire u2__abc_52155_new_n13234_; 
wire u2__abc_52155_new_n13235_; 
wire u2__abc_52155_new_n13236_; 
wire u2__abc_52155_new_n13237_; 
wire u2__abc_52155_new_n13238_; 
wire u2__abc_52155_new_n13239_; 
wire u2__abc_52155_new_n13241_; 
wire u2__abc_52155_new_n13242_; 
wire u2__abc_52155_new_n13243_; 
wire u2__abc_52155_new_n13244_; 
wire u2__abc_52155_new_n13245_; 
wire u2__abc_52155_new_n13246_; 
wire u2__abc_52155_new_n13247_; 
wire u2__abc_52155_new_n13248_; 
wire u2__abc_52155_new_n13249_; 
wire u2__abc_52155_new_n13250_; 
wire u2__abc_52155_new_n13251_; 
wire u2__abc_52155_new_n13252_; 
wire u2__abc_52155_new_n13253_; 
wire u2__abc_52155_new_n13254_; 
wire u2__abc_52155_new_n13255_; 
wire u2__abc_52155_new_n13256_; 
wire u2__abc_52155_new_n13257_; 
wire u2__abc_52155_new_n13258_; 
wire u2__abc_52155_new_n13260_; 
wire u2__abc_52155_new_n13261_; 
wire u2__abc_52155_new_n13262_; 
wire u2__abc_52155_new_n13263_; 
wire u2__abc_52155_new_n13264_; 
wire u2__abc_52155_new_n13265_; 
wire u2__abc_52155_new_n13266_; 
wire u2__abc_52155_new_n13267_; 
wire u2__abc_52155_new_n13268_; 
wire u2__abc_52155_new_n13269_; 
wire u2__abc_52155_new_n13270_; 
wire u2__abc_52155_new_n13271_; 
wire u2__abc_52155_new_n13272_; 
wire u2__abc_52155_new_n13273_; 
wire u2__abc_52155_new_n13274_; 
wire u2__abc_52155_new_n13275_; 
wire u2__abc_52155_new_n13277_; 
wire u2__abc_52155_new_n13278_; 
wire u2__abc_52155_new_n13279_; 
wire u2__abc_52155_new_n13280_; 
wire u2__abc_52155_new_n13281_; 
wire u2__abc_52155_new_n13282_; 
wire u2__abc_52155_new_n13283_; 
wire u2__abc_52155_new_n13284_; 
wire u2__abc_52155_new_n13285_; 
wire u2__abc_52155_new_n13286_; 
wire u2__abc_52155_new_n13287_; 
wire u2__abc_52155_new_n13288_; 
wire u2__abc_52155_new_n13289_; 
wire u2__abc_52155_new_n13290_; 
wire u2__abc_52155_new_n13291_; 
wire u2__abc_52155_new_n13292_; 
wire u2__abc_52155_new_n13293_; 
wire u2__abc_52155_new_n13294_; 
wire u2__abc_52155_new_n13295_; 
wire u2__abc_52155_new_n13296_; 
wire u2__abc_52155_new_n13297_; 
wire u2__abc_52155_new_n13298_; 
wire u2__abc_52155_new_n13299_; 
wire u2__abc_52155_new_n13300_; 
wire u2__abc_52155_new_n13301_; 
wire u2__abc_52155_new_n13302_; 
wire u2__abc_52155_new_n13303_; 
wire u2__abc_52155_new_n13304_; 
wire u2__abc_52155_new_n13305_; 
wire u2__abc_52155_new_n13306_; 
wire u2__abc_52155_new_n13307_; 
wire u2__abc_52155_new_n13308_; 
wire u2__abc_52155_new_n13310_; 
wire u2__abc_52155_new_n13311_; 
wire u2__abc_52155_new_n13312_; 
wire u2__abc_52155_new_n13313_; 
wire u2__abc_52155_new_n13314_; 
wire u2__abc_52155_new_n13315_; 
wire u2__abc_52155_new_n13316_; 
wire u2__abc_52155_new_n13317_; 
wire u2__abc_52155_new_n13318_; 
wire u2__abc_52155_new_n13319_; 
wire u2__abc_52155_new_n13320_; 
wire u2__abc_52155_new_n13321_; 
wire u2__abc_52155_new_n13322_; 
wire u2__abc_52155_new_n13323_; 
wire u2__abc_52155_new_n13324_; 
wire u2__abc_52155_new_n13325_; 
wire u2__abc_52155_new_n13327_; 
wire u2__abc_52155_new_n13328_; 
wire u2__abc_52155_new_n13329_; 
wire u2__abc_52155_new_n13330_; 
wire u2__abc_52155_new_n13331_; 
wire u2__abc_52155_new_n13332_; 
wire u2__abc_52155_new_n13333_; 
wire u2__abc_52155_new_n13334_; 
wire u2__abc_52155_new_n13335_; 
wire u2__abc_52155_new_n13336_; 
wire u2__abc_52155_new_n13337_; 
wire u2__abc_52155_new_n13338_; 
wire u2__abc_52155_new_n13339_; 
wire u2__abc_52155_new_n13340_; 
wire u2__abc_52155_new_n13341_; 
wire u2__abc_52155_new_n13342_; 
wire u2__abc_52155_new_n13343_; 
wire u2__abc_52155_new_n13344_; 
wire u2__abc_52155_new_n13346_; 
wire u2__abc_52155_new_n13347_; 
wire u2__abc_52155_new_n13348_; 
wire u2__abc_52155_new_n13349_; 
wire u2__abc_52155_new_n13350_; 
wire u2__abc_52155_new_n13351_; 
wire u2__abc_52155_new_n13352_; 
wire u2__abc_52155_new_n13353_; 
wire u2__abc_52155_new_n13354_; 
wire u2__abc_52155_new_n13355_; 
wire u2__abc_52155_new_n13356_; 
wire u2__abc_52155_new_n13357_; 
wire u2__abc_52155_new_n13358_; 
wire u2__abc_52155_new_n13359_; 
wire u2__abc_52155_new_n13360_; 
wire u2__abc_52155_new_n13361_; 
wire u2__abc_52155_new_n13363_; 
wire u2__abc_52155_new_n13364_; 
wire u2__abc_52155_new_n13365_; 
wire u2__abc_52155_new_n13366_; 
wire u2__abc_52155_new_n13367_; 
wire u2__abc_52155_new_n13368_; 
wire u2__abc_52155_new_n13369_; 
wire u2__abc_52155_new_n13370_; 
wire u2__abc_52155_new_n13371_; 
wire u2__abc_52155_new_n13372_; 
wire u2__abc_52155_new_n13373_; 
wire u2__abc_52155_new_n13374_; 
wire u2__abc_52155_new_n13375_; 
wire u2__abc_52155_new_n13376_; 
wire u2__abc_52155_new_n13377_; 
wire u2__abc_52155_new_n13378_; 
wire u2__abc_52155_new_n13379_; 
wire u2__abc_52155_new_n13380_; 
wire u2__abc_52155_new_n13381_; 
wire u2__abc_52155_new_n13382_; 
wire u2__abc_52155_new_n13383_; 
wire u2__abc_52155_new_n13384_; 
wire u2__abc_52155_new_n13385_; 
wire u2__abc_52155_new_n13387_; 
wire u2__abc_52155_new_n13388_; 
wire u2__abc_52155_new_n13389_; 
wire u2__abc_52155_new_n13390_; 
wire u2__abc_52155_new_n13391_; 
wire u2__abc_52155_new_n13392_; 
wire u2__abc_52155_new_n13393_; 
wire u2__abc_52155_new_n13394_; 
wire u2__abc_52155_new_n13395_; 
wire u2__abc_52155_new_n13396_; 
wire u2__abc_52155_new_n13397_; 
wire u2__abc_52155_new_n13398_; 
wire u2__abc_52155_new_n13399_; 
wire u2__abc_52155_new_n13400_; 
wire u2__abc_52155_new_n13401_; 
wire u2__abc_52155_new_n13402_; 
wire u2__abc_52155_new_n13404_; 
wire u2__abc_52155_new_n13405_; 
wire u2__abc_52155_new_n13406_; 
wire u2__abc_52155_new_n13407_; 
wire u2__abc_52155_new_n13408_; 
wire u2__abc_52155_new_n13409_; 
wire u2__abc_52155_new_n13410_; 
wire u2__abc_52155_new_n13411_; 
wire u2__abc_52155_new_n13412_; 
wire u2__abc_52155_new_n13413_; 
wire u2__abc_52155_new_n13414_; 
wire u2__abc_52155_new_n13415_; 
wire u2__abc_52155_new_n13416_; 
wire u2__abc_52155_new_n13417_; 
wire u2__abc_52155_new_n13418_; 
wire u2__abc_52155_new_n13419_; 
wire u2__abc_52155_new_n13420_; 
wire u2__abc_52155_new_n13421_; 
wire u2__abc_52155_new_n13423_; 
wire u2__abc_52155_new_n13424_; 
wire u2__abc_52155_new_n13425_; 
wire u2__abc_52155_new_n13426_; 
wire u2__abc_52155_new_n13427_; 
wire u2__abc_52155_new_n13428_; 
wire u2__abc_52155_new_n13429_; 
wire u2__abc_52155_new_n13430_; 
wire u2__abc_52155_new_n13431_; 
wire u2__abc_52155_new_n13432_; 
wire u2__abc_52155_new_n13433_; 
wire u2__abc_52155_new_n13434_; 
wire u2__abc_52155_new_n13435_; 
wire u2__abc_52155_new_n13436_; 
wire u2__abc_52155_new_n13437_; 
wire u2__abc_52155_new_n13438_; 
wire u2__abc_52155_new_n13440_; 
wire u2__abc_52155_new_n13441_; 
wire u2__abc_52155_new_n13442_; 
wire u2__abc_52155_new_n13443_; 
wire u2__abc_52155_new_n13444_; 
wire u2__abc_52155_new_n13445_; 
wire u2__abc_52155_new_n13446_; 
wire u2__abc_52155_new_n13447_; 
wire u2__abc_52155_new_n13448_; 
wire u2__abc_52155_new_n13449_; 
wire u2__abc_52155_new_n13450_; 
wire u2__abc_52155_new_n13451_; 
wire u2__abc_52155_new_n13452_; 
wire u2__abc_52155_new_n13453_; 
wire u2__abc_52155_new_n13454_; 
wire u2__abc_52155_new_n13455_; 
wire u2__abc_52155_new_n13456_; 
wire u2__abc_52155_new_n13457_; 
wire u2__abc_52155_new_n13458_; 
wire u2__abc_52155_new_n13459_; 
wire u2__abc_52155_new_n13460_; 
wire u2__abc_52155_new_n13461_; 
wire u2__abc_52155_new_n13462_; 
wire u2__abc_52155_new_n13463_; 
wire u2__abc_52155_new_n13464_; 
wire u2__abc_52155_new_n13466_; 
wire u2__abc_52155_new_n13467_; 
wire u2__abc_52155_new_n13468_; 
wire u2__abc_52155_new_n13469_; 
wire u2__abc_52155_new_n13470_; 
wire u2__abc_52155_new_n13471_; 
wire u2__abc_52155_new_n13472_; 
wire u2__abc_52155_new_n13473_; 
wire u2__abc_52155_new_n13474_; 
wire u2__abc_52155_new_n13475_; 
wire u2__abc_52155_new_n13476_; 
wire u2__abc_52155_new_n13477_; 
wire u2__abc_52155_new_n13478_; 
wire u2__abc_52155_new_n13479_; 
wire u2__abc_52155_new_n13480_; 
wire u2__abc_52155_new_n13481_; 
wire u2__abc_52155_new_n13483_; 
wire u2__abc_52155_new_n13484_; 
wire u2__abc_52155_new_n13485_; 
wire u2__abc_52155_new_n13486_; 
wire u2__abc_52155_new_n13487_; 
wire u2__abc_52155_new_n13488_; 
wire u2__abc_52155_new_n13489_; 
wire u2__abc_52155_new_n13490_; 
wire u2__abc_52155_new_n13491_; 
wire u2__abc_52155_new_n13492_; 
wire u2__abc_52155_new_n13493_; 
wire u2__abc_52155_new_n13494_; 
wire u2__abc_52155_new_n13495_; 
wire u2__abc_52155_new_n13496_; 
wire u2__abc_52155_new_n13497_; 
wire u2__abc_52155_new_n13498_; 
wire u2__abc_52155_new_n13499_; 
wire u2__abc_52155_new_n13500_; 
wire u2__abc_52155_new_n13501_; 
wire u2__abc_52155_new_n13503_; 
wire u2__abc_52155_new_n13504_; 
wire u2__abc_52155_new_n13505_; 
wire u2__abc_52155_new_n13506_; 
wire u2__abc_52155_new_n13507_; 
wire u2__abc_52155_new_n13508_; 
wire u2__abc_52155_new_n13509_; 
wire u2__abc_52155_new_n13510_; 
wire u2__abc_52155_new_n13511_; 
wire u2__abc_52155_new_n13512_; 
wire u2__abc_52155_new_n13513_; 
wire u2__abc_52155_new_n13514_; 
wire u2__abc_52155_new_n13515_; 
wire u2__abc_52155_new_n13516_; 
wire u2__abc_52155_new_n13517_; 
wire u2__abc_52155_new_n13518_; 
wire u2__abc_52155_new_n13520_; 
wire u2__abc_52155_new_n13521_; 
wire u2__abc_52155_new_n13522_; 
wire u2__abc_52155_new_n13523_; 
wire u2__abc_52155_new_n13524_; 
wire u2__abc_52155_new_n13525_; 
wire u2__abc_52155_new_n13526_; 
wire u2__abc_52155_new_n13527_; 
wire u2__abc_52155_new_n13528_; 
wire u2__abc_52155_new_n13529_; 
wire u2__abc_52155_new_n13530_; 
wire u2__abc_52155_new_n13531_; 
wire u2__abc_52155_new_n13532_; 
wire u2__abc_52155_new_n13533_; 
wire u2__abc_52155_new_n13534_; 
wire u2__abc_52155_new_n13535_; 
wire u2__abc_52155_new_n13536_; 
wire u2__abc_52155_new_n13537_; 
wire u2__abc_52155_new_n13538_; 
wire u2__abc_52155_new_n13539_; 
wire u2__abc_52155_new_n13541_; 
wire u2__abc_52155_new_n13542_; 
wire u2__abc_52155_new_n13543_; 
wire u2__abc_52155_new_n13544_; 
wire u2__abc_52155_new_n13545_; 
wire u2__abc_52155_new_n13546_; 
wire u2__abc_52155_new_n13547_; 
wire u2__abc_52155_new_n13548_; 
wire u2__abc_52155_new_n13549_; 
wire u2__abc_52155_new_n13550_; 
wire u2__abc_52155_new_n13551_; 
wire u2__abc_52155_new_n13552_; 
wire u2__abc_52155_new_n13553_; 
wire u2__abc_52155_new_n13554_; 
wire u2__abc_52155_new_n13555_; 
wire u2__abc_52155_new_n13556_; 
wire u2__abc_52155_new_n13558_; 
wire u2__abc_52155_new_n13559_; 
wire u2__abc_52155_new_n13560_; 
wire u2__abc_52155_new_n13561_; 
wire u2__abc_52155_new_n13562_; 
wire u2__abc_52155_new_n13563_; 
wire u2__abc_52155_new_n13564_; 
wire u2__abc_52155_new_n13565_; 
wire u2__abc_52155_new_n13566_; 
wire u2__abc_52155_new_n13567_; 
wire u2__abc_52155_new_n13568_; 
wire u2__abc_52155_new_n13569_; 
wire u2__abc_52155_new_n13570_; 
wire u2__abc_52155_new_n13571_; 
wire u2__abc_52155_new_n13572_; 
wire u2__abc_52155_new_n13573_; 
wire u2__abc_52155_new_n13574_; 
wire u2__abc_52155_new_n13575_; 
wire u2__abc_52155_new_n13577_; 
wire u2__abc_52155_new_n13578_; 
wire u2__abc_52155_new_n13579_; 
wire u2__abc_52155_new_n13580_; 
wire u2__abc_52155_new_n13581_; 
wire u2__abc_52155_new_n13582_; 
wire u2__abc_52155_new_n13583_; 
wire u2__abc_52155_new_n13584_; 
wire u2__abc_52155_new_n13585_; 
wire u2__abc_52155_new_n13586_; 
wire u2__abc_52155_new_n13587_; 
wire u2__abc_52155_new_n13588_; 
wire u2__abc_52155_new_n13589_; 
wire u2__abc_52155_new_n13590_; 
wire u2__abc_52155_new_n13591_; 
wire u2__abc_52155_new_n13592_; 
wire u2__abc_52155_new_n13594_; 
wire u2__abc_52155_new_n13595_; 
wire u2__abc_52155_new_n13596_; 
wire u2__abc_52155_new_n13597_; 
wire u2__abc_52155_new_n13598_; 
wire u2__abc_52155_new_n13599_; 
wire u2__abc_52155_new_n13600_; 
wire u2__abc_52155_new_n13601_; 
wire u2__abc_52155_new_n13602_; 
wire u2__abc_52155_new_n13603_; 
wire u2__abc_52155_new_n13604_; 
wire u2__abc_52155_new_n13605_; 
wire u2__abc_52155_new_n13606_; 
wire u2__abc_52155_new_n13607_; 
wire u2__abc_52155_new_n13608_; 
wire u2__abc_52155_new_n13609_; 
wire u2__abc_52155_new_n13610_; 
wire u2__abc_52155_new_n13611_; 
wire u2__abc_52155_new_n13612_; 
wire u2__abc_52155_new_n13613_; 
wire u2__abc_52155_new_n13614_; 
wire u2__abc_52155_new_n13615_; 
wire u2__abc_52155_new_n13616_; 
wire u2__abc_52155_new_n13617_; 
wire u2__abc_52155_new_n13618_; 
wire u2__abc_52155_new_n13619_; 
wire u2__abc_52155_new_n13620_; 
wire u2__abc_52155_new_n13621_; 
wire u2__abc_52155_new_n13622_; 
wire u2__abc_52155_new_n13624_; 
wire u2__abc_52155_new_n13625_; 
wire u2__abc_52155_new_n13626_; 
wire u2__abc_52155_new_n13627_; 
wire u2__abc_52155_new_n13628_; 
wire u2__abc_52155_new_n13629_; 
wire u2__abc_52155_new_n13630_; 
wire u2__abc_52155_new_n13631_; 
wire u2__abc_52155_new_n13632_; 
wire u2__abc_52155_new_n13633_; 
wire u2__abc_52155_new_n13634_; 
wire u2__abc_52155_new_n13635_; 
wire u2__abc_52155_new_n13636_; 
wire u2__abc_52155_new_n13637_; 
wire u2__abc_52155_new_n13638_; 
wire u2__abc_52155_new_n13639_; 
wire u2__abc_52155_new_n13641_; 
wire u2__abc_52155_new_n13642_; 
wire u2__abc_52155_new_n13643_; 
wire u2__abc_52155_new_n13644_; 
wire u2__abc_52155_new_n13645_; 
wire u2__abc_52155_new_n13646_; 
wire u2__abc_52155_new_n13647_; 
wire u2__abc_52155_new_n13648_; 
wire u2__abc_52155_new_n13649_; 
wire u2__abc_52155_new_n13650_; 
wire u2__abc_52155_new_n13651_; 
wire u2__abc_52155_new_n13652_; 
wire u2__abc_52155_new_n13653_; 
wire u2__abc_52155_new_n13654_; 
wire u2__abc_52155_new_n13655_; 
wire u2__abc_52155_new_n13656_; 
wire u2__abc_52155_new_n13657_; 
wire u2__abc_52155_new_n13658_; 
wire u2__abc_52155_new_n13659_; 
wire u2__abc_52155_new_n13661_; 
wire u2__abc_52155_new_n13662_; 
wire u2__abc_52155_new_n13663_; 
wire u2__abc_52155_new_n13664_; 
wire u2__abc_52155_new_n13665_; 
wire u2__abc_52155_new_n13666_; 
wire u2__abc_52155_new_n13667_; 
wire u2__abc_52155_new_n13668_; 
wire u2__abc_52155_new_n13669_; 
wire u2__abc_52155_new_n13670_; 
wire u2__abc_52155_new_n13671_; 
wire u2__abc_52155_new_n13672_; 
wire u2__abc_52155_new_n13673_; 
wire u2__abc_52155_new_n13674_; 
wire u2__abc_52155_new_n13675_; 
wire u2__abc_52155_new_n13676_; 
wire u2__abc_52155_new_n13678_; 
wire u2__abc_52155_new_n13679_; 
wire u2__abc_52155_new_n13680_; 
wire u2__abc_52155_new_n13681_; 
wire u2__abc_52155_new_n13682_; 
wire u2__abc_52155_new_n13683_; 
wire u2__abc_52155_new_n13684_; 
wire u2__abc_52155_new_n13685_; 
wire u2__abc_52155_new_n13686_; 
wire u2__abc_52155_new_n13687_; 
wire u2__abc_52155_new_n13688_; 
wire u2__abc_52155_new_n13689_; 
wire u2__abc_52155_new_n13690_; 
wire u2__abc_52155_new_n13691_; 
wire u2__abc_52155_new_n13692_; 
wire u2__abc_52155_new_n13693_; 
wire u2__abc_52155_new_n13694_; 
wire u2__abc_52155_new_n13695_; 
wire u2__abc_52155_new_n13696_; 
wire u2__abc_52155_new_n13697_; 
wire u2__abc_52155_new_n13699_; 
wire u2__abc_52155_new_n13700_; 
wire u2__abc_52155_new_n13701_; 
wire u2__abc_52155_new_n13702_; 
wire u2__abc_52155_new_n13703_; 
wire u2__abc_52155_new_n13704_; 
wire u2__abc_52155_new_n13705_; 
wire u2__abc_52155_new_n13706_; 
wire u2__abc_52155_new_n13707_; 
wire u2__abc_52155_new_n13708_; 
wire u2__abc_52155_new_n13709_; 
wire u2__abc_52155_new_n13710_; 
wire u2__abc_52155_new_n13711_; 
wire u2__abc_52155_new_n13712_; 
wire u2__abc_52155_new_n13713_; 
wire u2__abc_52155_new_n13714_; 
wire u2__abc_52155_new_n13716_; 
wire u2__abc_52155_new_n13717_; 
wire u2__abc_52155_new_n13718_; 
wire u2__abc_52155_new_n13719_; 
wire u2__abc_52155_new_n13720_; 
wire u2__abc_52155_new_n13721_; 
wire u2__abc_52155_new_n13722_; 
wire u2__abc_52155_new_n13723_; 
wire u2__abc_52155_new_n13724_; 
wire u2__abc_52155_new_n13725_; 
wire u2__abc_52155_new_n13726_; 
wire u2__abc_52155_new_n13727_; 
wire u2__abc_52155_new_n13728_; 
wire u2__abc_52155_new_n13729_; 
wire u2__abc_52155_new_n13730_; 
wire u2__abc_52155_new_n13731_; 
wire u2__abc_52155_new_n13733_; 
wire u2__abc_52155_new_n13734_; 
wire u2__abc_52155_new_n13735_; 
wire u2__abc_52155_new_n13736_; 
wire u2__abc_52155_new_n13737_; 
wire u2__abc_52155_new_n13738_; 
wire u2__abc_52155_new_n13739_; 
wire u2__abc_52155_new_n13740_; 
wire u2__abc_52155_new_n13741_; 
wire u2__abc_52155_new_n13742_; 
wire u2__abc_52155_new_n13743_; 
wire u2__abc_52155_new_n13744_; 
wire u2__abc_52155_new_n13745_; 
wire u2__abc_52155_new_n13746_; 
wire u2__abc_52155_new_n13747_; 
wire u2__abc_52155_new_n13748_; 
wire u2__abc_52155_new_n13750_; 
wire u2__abc_52155_new_n13751_; 
wire u2__abc_52155_new_n13752_; 
wire u2__abc_52155_new_n13753_; 
wire u2__abc_52155_new_n13754_; 
wire u2__abc_52155_new_n13755_; 
wire u2__abc_52155_new_n13756_; 
wire u2__abc_52155_new_n13757_; 
wire u2__abc_52155_new_n13758_; 
wire u2__abc_52155_new_n13759_; 
wire u2__abc_52155_new_n13760_; 
wire u2__abc_52155_new_n13761_; 
wire u2__abc_52155_new_n13762_; 
wire u2__abc_52155_new_n13763_; 
wire u2__abc_52155_new_n13764_; 
wire u2__abc_52155_new_n13765_; 
wire u2__abc_52155_new_n13766_; 
wire u2__abc_52155_new_n13767_; 
wire u2__abc_52155_new_n13768_; 
wire u2__abc_52155_new_n13769_; 
wire u2__abc_52155_new_n13770_; 
wire u2__abc_52155_new_n13771_; 
wire u2__abc_52155_new_n13772_; 
wire u2__abc_52155_new_n13773_; 
wire u2__abc_52155_new_n13775_; 
wire u2__abc_52155_new_n13776_; 
wire u2__abc_52155_new_n13777_; 
wire u2__abc_52155_new_n13778_; 
wire u2__abc_52155_new_n13779_; 
wire u2__abc_52155_new_n13780_; 
wire u2__abc_52155_new_n13781_; 
wire u2__abc_52155_new_n13782_; 
wire u2__abc_52155_new_n13783_; 
wire u2__abc_52155_new_n13784_; 
wire u2__abc_52155_new_n13785_; 
wire u2__abc_52155_new_n13786_; 
wire u2__abc_52155_new_n13787_; 
wire u2__abc_52155_new_n13788_; 
wire u2__abc_52155_new_n13789_; 
wire u2__abc_52155_new_n13790_; 
wire u2__abc_52155_new_n13792_; 
wire u2__abc_52155_new_n13793_; 
wire u2__abc_52155_new_n13794_; 
wire u2__abc_52155_new_n13795_; 
wire u2__abc_52155_new_n13796_; 
wire u2__abc_52155_new_n13797_; 
wire u2__abc_52155_new_n13798_; 
wire u2__abc_52155_new_n13799_; 
wire u2__abc_52155_new_n13800_; 
wire u2__abc_52155_new_n13801_; 
wire u2__abc_52155_new_n13802_; 
wire u2__abc_52155_new_n13803_; 
wire u2__abc_52155_new_n13804_; 
wire u2__abc_52155_new_n13805_; 
wire u2__abc_52155_new_n13806_; 
wire u2__abc_52155_new_n13807_; 
wire u2__abc_52155_new_n13808_; 
wire u2__abc_52155_new_n13809_; 
wire u2__abc_52155_new_n13811_; 
wire u2__abc_52155_new_n13812_; 
wire u2__abc_52155_new_n13813_; 
wire u2__abc_52155_new_n13814_; 
wire u2__abc_52155_new_n13815_; 
wire u2__abc_52155_new_n13816_; 
wire u2__abc_52155_new_n13817_; 
wire u2__abc_52155_new_n13818_; 
wire u2__abc_52155_new_n13819_; 
wire u2__abc_52155_new_n13820_; 
wire u2__abc_52155_new_n13821_; 
wire u2__abc_52155_new_n13822_; 
wire u2__abc_52155_new_n13823_; 
wire u2__abc_52155_new_n13824_; 
wire u2__abc_52155_new_n13825_; 
wire u2__abc_52155_new_n13826_; 
wire u2__abc_52155_new_n13828_; 
wire u2__abc_52155_new_n13829_; 
wire u2__abc_52155_new_n13830_; 
wire u2__abc_52155_new_n13831_; 
wire u2__abc_52155_new_n13832_; 
wire u2__abc_52155_new_n13833_; 
wire u2__abc_52155_new_n13834_; 
wire u2__abc_52155_new_n13835_; 
wire u2__abc_52155_new_n13836_; 
wire u2__abc_52155_new_n13837_; 
wire u2__abc_52155_new_n13838_; 
wire u2__abc_52155_new_n13839_; 
wire u2__abc_52155_new_n13840_; 
wire u2__abc_52155_new_n13841_; 
wire u2__abc_52155_new_n13842_; 
wire u2__abc_52155_new_n13843_; 
wire u2__abc_52155_new_n13844_; 
wire u2__abc_52155_new_n13845_; 
wire u2__abc_52155_new_n13846_; 
wire u2__abc_52155_new_n13847_; 
wire u2__abc_52155_new_n13848_; 
wire u2__abc_52155_new_n13849_; 
wire u2__abc_52155_new_n13850_; 
wire u2__abc_52155_new_n13851_; 
wire u2__abc_52155_new_n13853_; 
wire u2__abc_52155_new_n13854_; 
wire u2__abc_52155_new_n13855_; 
wire u2__abc_52155_new_n13856_; 
wire u2__abc_52155_new_n13857_; 
wire u2__abc_52155_new_n13858_; 
wire u2__abc_52155_new_n13859_; 
wire u2__abc_52155_new_n13860_; 
wire u2__abc_52155_new_n13861_; 
wire u2__abc_52155_new_n13862_; 
wire u2__abc_52155_new_n13863_; 
wire u2__abc_52155_new_n13864_; 
wire u2__abc_52155_new_n13865_; 
wire u2__abc_52155_new_n13866_; 
wire u2__abc_52155_new_n13867_; 
wire u2__abc_52155_new_n13868_; 
wire u2__abc_52155_new_n13870_; 
wire u2__abc_52155_new_n13871_; 
wire u2__abc_52155_new_n13872_; 
wire u2__abc_52155_new_n13873_; 
wire u2__abc_52155_new_n13874_; 
wire u2__abc_52155_new_n13875_; 
wire u2__abc_52155_new_n13876_; 
wire u2__abc_52155_new_n13877_; 
wire u2__abc_52155_new_n13878_; 
wire u2__abc_52155_new_n13879_; 
wire u2__abc_52155_new_n13880_; 
wire u2__abc_52155_new_n13881_; 
wire u2__abc_52155_new_n13882_; 
wire u2__abc_52155_new_n13883_; 
wire u2__abc_52155_new_n13884_; 
wire u2__abc_52155_new_n13885_; 
wire u2__abc_52155_new_n13886_; 
wire u2__abc_52155_new_n13887_; 
wire u2__abc_52155_new_n13889_; 
wire u2__abc_52155_new_n13890_; 
wire u2__abc_52155_new_n13891_; 
wire u2__abc_52155_new_n13892_; 
wire u2__abc_52155_new_n13893_; 
wire u2__abc_52155_new_n13894_; 
wire u2__abc_52155_new_n13895_; 
wire u2__abc_52155_new_n13896_; 
wire u2__abc_52155_new_n13897_; 
wire u2__abc_52155_new_n13898_; 
wire u2__abc_52155_new_n13899_; 
wire u2__abc_52155_new_n13900_; 
wire u2__abc_52155_new_n13901_; 
wire u2__abc_52155_new_n13902_; 
wire u2__abc_52155_new_n13903_; 
wire u2__abc_52155_new_n13904_; 
wire u2__abc_52155_new_n13906_; 
wire u2__abc_52155_new_n13907_; 
wire u2__abc_52155_new_n13908_; 
wire u2__abc_52155_new_n13909_; 
wire u2__abc_52155_new_n13910_; 
wire u2__abc_52155_new_n13911_; 
wire u2__abc_52155_new_n13912_; 
wire u2__abc_52155_new_n13913_; 
wire u2__abc_52155_new_n13914_; 
wire u2__abc_52155_new_n13915_; 
wire u2__abc_52155_new_n13916_; 
wire u2__abc_52155_new_n13917_; 
wire u2__abc_52155_new_n13918_; 
wire u2__abc_52155_new_n13919_; 
wire u2__abc_52155_new_n13920_; 
wire u2__abc_52155_new_n13921_; 
wire u2__abc_52155_new_n13922_; 
wire u2__abc_52155_new_n13923_; 
wire u2__abc_52155_new_n13924_; 
wire u2__abc_52155_new_n13925_; 
wire u2__abc_52155_new_n13926_; 
wire u2__abc_52155_new_n13927_; 
wire u2__abc_52155_new_n13928_; 
wire u2__abc_52155_new_n13929_; 
wire u2__abc_52155_new_n13930_; 
wire u2__abc_52155_new_n13931_; 
wire u2__abc_52155_new_n13932_; 
wire u2__abc_52155_new_n13933_; 
wire u2__abc_52155_new_n13934_; 
wire u2__abc_52155_new_n13935_; 
wire u2__abc_52155_new_n13936_; 
wire u2__abc_52155_new_n13937_; 
wire u2__abc_52155_new_n13938_; 
wire u2__abc_52155_new_n13939_; 
wire u2__abc_52155_new_n13940_; 
wire u2__abc_52155_new_n13941_; 
wire u2__abc_52155_new_n13943_; 
wire u2__abc_52155_new_n13944_; 
wire u2__abc_52155_new_n13945_; 
wire u2__abc_52155_new_n13946_; 
wire u2__abc_52155_new_n13947_; 
wire u2__abc_52155_new_n13948_; 
wire u2__abc_52155_new_n13949_; 
wire u2__abc_52155_new_n13950_; 
wire u2__abc_52155_new_n13951_; 
wire u2__abc_52155_new_n13952_; 
wire u2__abc_52155_new_n13953_; 
wire u2__abc_52155_new_n13954_; 
wire u2__abc_52155_new_n13955_; 
wire u2__abc_52155_new_n13956_; 
wire u2__abc_52155_new_n13957_; 
wire u2__abc_52155_new_n13958_; 
wire u2__abc_52155_new_n13960_; 
wire u2__abc_52155_new_n13961_; 
wire u2__abc_52155_new_n13962_; 
wire u2__abc_52155_new_n13963_; 
wire u2__abc_52155_new_n13964_; 
wire u2__abc_52155_new_n13965_; 
wire u2__abc_52155_new_n13966_; 
wire u2__abc_52155_new_n13967_; 
wire u2__abc_52155_new_n13968_; 
wire u2__abc_52155_new_n13969_; 
wire u2__abc_52155_new_n13970_; 
wire u2__abc_52155_new_n13971_; 
wire u2__abc_52155_new_n13972_; 
wire u2__abc_52155_new_n13973_; 
wire u2__abc_52155_new_n13974_; 
wire u2__abc_52155_new_n13975_; 
wire u2__abc_52155_new_n13976_; 
wire u2__abc_52155_new_n13977_; 
wire u2__abc_52155_new_n13978_; 
wire u2__abc_52155_new_n13980_; 
wire u2__abc_52155_new_n13981_; 
wire u2__abc_52155_new_n13982_; 
wire u2__abc_52155_new_n13983_; 
wire u2__abc_52155_new_n13984_; 
wire u2__abc_52155_new_n13985_; 
wire u2__abc_52155_new_n13986_; 
wire u2__abc_52155_new_n13987_; 
wire u2__abc_52155_new_n13988_; 
wire u2__abc_52155_new_n13989_; 
wire u2__abc_52155_new_n13990_; 
wire u2__abc_52155_new_n13991_; 
wire u2__abc_52155_new_n13992_; 
wire u2__abc_52155_new_n13993_; 
wire u2__abc_52155_new_n13994_; 
wire u2__abc_52155_new_n13995_; 
wire u2__abc_52155_new_n13997_; 
wire u2__abc_52155_new_n13998_; 
wire u2__abc_52155_new_n13999_; 
wire u2__abc_52155_new_n14000_; 
wire u2__abc_52155_new_n14001_; 
wire u2__abc_52155_new_n14002_; 
wire u2__abc_52155_new_n14003_; 
wire u2__abc_52155_new_n14004_; 
wire u2__abc_52155_new_n14005_; 
wire u2__abc_52155_new_n14006_; 
wire u2__abc_52155_new_n14007_; 
wire u2__abc_52155_new_n14008_; 
wire u2__abc_52155_new_n14009_; 
wire u2__abc_52155_new_n14010_; 
wire u2__abc_52155_new_n14011_; 
wire u2__abc_52155_new_n14012_; 
wire u2__abc_52155_new_n14013_; 
wire u2__abc_52155_new_n14014_; 
wire u2__abc_52155_new_n14015_; 
wire u2__abc_52155_new_n14016_; 
wire u2__abc_52155_new_n14018_; 
wire u2__abc_52155_new_n14019_; 
wire u2__abc_52155_new_n14020_; 
wire u2__abc_52155_new_n14021_; 
wire u2__abc_52155_new_n14022_; 
wire u2__abc_52155_new_n14023_; 
wire u2__abc_52155_new_n14024_; 
wire u2__abc_52155_new_n14025_; 
wire u2__abc_52155_new_n14026_; 
wire u2__abc_52155_new_n14027_; 
wire u2__abc_52155_new_n14028_; 
wire u2__abc_52155_new_n14029_; 
wire u2__abc_52155_new_n14030_; 
wire u2__abc_52155_new_n14031_; 
wire u2__abc_52155_new_n14032_; 
wire u2__abc_52155_new_n14033_; 
wire u2__abc_52155_new_n14035_; 
wire u2__abc_52155_new_n14036_; 
wire u2__abc_52155_new_n14037_; 
wire u2__abc_52155_new_n14038_; 
wire u2__abc_52155_new_n14039_; 
wire u2__abc_52155_new_n14040_; 
wire u2__abc_52155_new_n14041_; 
wire u2__abc_52155_new_n14042_; 
wire u2__abc_52155_new_n14043_; 
wire u2__abc_52155_new_n14044_; 
wire u2__abc_52155_new_n14045_; 
wire u2__abc_52155_new_n14046_; 
wire u2__abc_52155_new_n14047_; 
wire u2__abc_52155_new_n14048_; 
wire u2__abc_52155_new_n14049_; 
wire u2__abc_52155_new_n14050_; 
wire u2__abc_52155_new_n14051_; 
wire u2__abc_52155_new_n14052_; 
wire u2__abc_52155_new_n14054_; 
wire u2__abc_52155_new_n14055_; 
wire u2__abc_52155_new_n14056_; 
wire u2__abc_52155_new_n14057_; 
wire u2__abc_52155_new_n14058_; 
wire u2__abc_52155_new_n14059_; 
wire u2__abc_52155_new_n14060_; 
wire u2__abc_52155_new_n14061_; 
wire u2__abc_52155_new_n14062_; 
wire u2__abc_52155_new_n14063_; 
wire u2__abc_52155_new_n14064_; 
wire u2__abc_52155_new_n14065_; 
wire u2__abc_52155_new_n14066_; 
wire u2__abc_52155_new_n14067_; 
wire u2__abc_52155_new_n14068_; 
wire u2__abc_52155_new_n14069_; 
wire u2__abc_52155_new_n14071_; 
wire u2__abc_52155_new_n14072_; 
wire u2__abc_52155_new_n14073_; 
wire u2__abc_52155_new_n14074_; 
wire u2__abc_52155_new_n14075_; 
wire u2__abc_52155_new_n14076_; 
wire u2__abc_52155_new_n14077_; 
wire u2__abc_52155_new_n14078_; 
wire u2__abc_52155_new_n14079_; 
wire u2__abc_52155_new_n14080_; 
wire u2__abc_52155_new_n14081_; 
wire u2__abc_52155_new_n14082_; 
wire u2__abc_52155_new_n14083_; 
wire u2__abc_52155_new_n14084_; 
wire u2__abc_52155_new_n14085_; 
wire u2__abc_52155_new_n14086_; 
wire u2__abc_52155_new_n14087_; 
wire u2__abc_52155_new_n14088_; 
wire u2__abc_52155_new_n14089_; 
wire u2__abc_52155_new_n14090_; 
wire u2__abc_52155_new_n14091_; 
wire u2__abc_52155_new_n14092_; 
wire u2__abc_52155_new_n14093_; 
wire u2__abc_52155_new_n14094_; 
wire u2__abc_52155_new_n14095_; 
wire u2__abc_52155_new_n14097_; 
wire u2__abc_52155_new_n14098_; 
wire u2__abc_52155_new_n14099_; 
wire u2__abc_52155_new_n14100_; 
wire u2__abc_52155_new_n14101_; 
wire u2__abc_52155_new_n14102_; 
wire u2__abc_52155_new_n14103_; 
wire u2__abc_52155_new_n14104_; 
wire u2__abc_52155_new_n14105_; 
wire u2__abc_52155_new_n14106_; 
wire u2__abc_52155_new_n14107_; 
wire u2__abc_52155_new_n14108_; 
wire u2__abc_52155_new_n14109_; 
wire u2__abc_52155_new_n14110_; 
wire u2__abc_52155_new_n14111_; 
wire u2__abc_52155_new_n14112_; 
wire u2__abc_52155_new_n14114_; 
wire u2__abc_52155_new_n14115_; 
wire u2__abc_52155_new_n14116_; 
wire u2__abc_52155_new_n14117_; 
wire u2__abc_52155_new_n14118_; 
wire u2__abc_52155_new_n14119_; 
wire u2__abc_52155_new_n14120_; 
wire u2__abc_52155_new_n14121_; 
wire u2__abc_52155_new_n14122_; 
wire u2__abc_52155_new_n14123_; 
wire u2__abc_52155_new_n14124_; 
wire u2__abc_52155_new_n14125_; 
wire u2__abc_52155_new_n14126_; 
wire u2__abc_52155_new_n14127_; 
wire u2__abc_52155_new_n14128_; 
wire u2__abc_52155_new_n14129_; 
wire u2__abc_52155_new_n14130_; 
wire u2__abc_52155_new_n14131_; 
wire u2__abc_52155_new_n14132_; 
wire u2__abc_52155_new_n14134_; 
wire u2__abc_52155_new_n14135_; 
wire u2__abc_52155_new_n14136_; 
wire u2__abc_52155_new_n14137_; 
wire u2__abc_52155_new_n14138_; 
wire u2__abc_52155_new_n14139_; 
wire u2__abc_52155_new_n14140_; 
wire u2__abc_52155_new_n14141_; 
wire u2__abc_52155_new_n14142_; 
wire u2__abc_52155_new_n14143_; 
wire u2__abc_52155_new_n14144_; 
wire u2__abc_52155_new_n14145_; 
wire u2__abc_52155_new_n14146_; 
wire u2__abc_52155_new_n14147_; 
wire u2__abc_52155_new_n14148_; 
wire u2__abc_52155_new_n14149_; 
wire u2__abc_52155_new_n14151_; 
wire u2__abc_52155_new_n14152_; 
wire u2__abc_52155_new_n14153_; 
wire u2__abc_52155_new_n14154_; 
wire u2__abc_52155_new_n14155_; 
wire u2__abc_52155_new_n14156_; 
wire u2__abc_52155_new_n14157_; 
wire u2__abc_52155_new_n14158_; 
wire u2__abc_52155_new_n14159_; 
wire u2__abc_52155_new_n14160_; 
wire u2__abc_52155_new_n14161_; 
wire u2__abc_52155_new_n14162_; 
wire u2__abc_52155_new_n14163_; 
wire u2__abc_52155_new_n14164_; 
wire u2__abc_52155_new_n14165_; 
wire u2__abc_52155_new_n14166_; 
wire u2__abc_52155_new_n14167_; 
wire u2__abc_52155_new_n14168_; 
wire u2__abc_52155_new_n14169_; 
wire u2__abc_52155_new_n14170_; 
wire u2__abc_52155_new_n14172_; 
wire u2__abc_52155_new_n14173_; 
wire u2__abc_52155_new_n14174_; 
wire u2__abc_52155_new_n14175_; 
wire u2__abc_52155_new_n14176_; 
wire u2__abc_52155_new_n14177_; 
wire u2__abc_52155_new_n14178_; 
wire u2__abc_52155_new_n14179_; 
wire u2__abc_52155_new_n14180_; 
wire u2__abc_52155_new_n14181_; 
wire u2__abc_52155_new_n14182_; 
wire u2__abc_52155_new_n14183_; 
wire u2__abc_52155_new_n14184_; 
wire u2__abc_52155_new_n14185_; 
wire u2__abc_52155_new_n14186_; 
wire u2__abc_52155_new_n14187_; 
wire u2__abc_52155_new_n14189_; 
wire u2__abc_52155_new_n14190_; 
wire u2__abc_52155_new_n14191_; 
wire u2__abc_52155_new_n14192_; 
wire u2__abc_52155_new_n14193_; 
wire u2__abc_52155_new_n14194_; 
wire u2__abc_52155_new_n14195_; 
wire u2__abc_52155_new_n14196_; 
wire u2__abc_52155_new_n14197_; 
wire u2__abc_52155_new_n14198_; 
wire u2__abc_52155_new_n14199_; 
wire u2__abc_52155_new_n14200_; 
wire u2__abc_52155_new_n14201_; 
wire u2__abc_52155_new_n14202_; 
wire u2__abc_52155_new_n14203_; 
wire u2__abc_52155_new_n14204_; 
wire u2__abc_52155_new_n14205_; 
wire u2__abc_52155_new_n14206_; 
wire u2__abc_52155_new_n14208_; 
wire u2__abc_52155_new_n14209_; 
wire u2__abc_52155_new_n14210_; 
wire u2__abc_52155_new_n14211_; 
wire u2__abc_52155_new_n14212_; 
wire u2__abc_52155_new_n14213_; 
wire u2__abc_52155_new_n14214_; 
wire u2__abc_52155_new_n14215_; 
wire u2__abc_52155_new_n14216_; 
wire u2__abc_52155_new_n14217_; 
wire u2__abc_52155_new_n14218_; 
wire u2__abc_52155_new_n14219_; 
wire u2__abc_52155_new_n14220_; 
wire u2__abc_52155_new_n14221_; 
wire u2__abc_52155_new_n14222_; 
wire u2__abc_52155_new_n14223_; 
wire u2__abc_52155_new_n14225_; 
wire u2__abc_52155_new_n14226_; 
wire u2__abc_52155_new_n14227_; 
wire u2__abc_52155_new_n14228_; 
wire u2__abc_52155_new_n14229_; 
wire u2__abc_52155_new_n14230_; 
wire u2__abc_52155_new_n14231_; 
wire u2__abc_52155_new_n14232_; 
wire u2__abc_52155_new_n14233_; 
wire u2__abc_52155_new_n14234_; 
wire u2__abc_52155_new_n14235_; 
wire u2__abc_52155_new_n14236_; 
wire u2__abc_52155_new_n14237_; 
wire u2__abc_52155_new_n14238_; 
wire u2__abc_52155_new_n14239_; 
wire u2__abc_52155_new_n14240_; 
wire u2__abc_52155_new_n14241_; 
wire u2__abc_52155_new_n14242_; 
wire u2__abc_52155_new_n14243_; 
wire u2__abc_52155_new_n14244_; 
wire u2__abc_52155_new_n14245_; 
wire u2__abc_52155_new_n14246_; 
wire u2__abc_52155_new_n14247_; 
wire u2__abc_52155_new_n14248_; 
wire u2__abc_52155_new_n14249_; 
wire u2__abc_52155_new_n14250_; 
wire u2__abc_52155_new_n14251_; 
wire u2__abc_52155_new_n14252_; 
wire u2__abc_52155_new_n14253_; 
wire u2__abc_52155_new_n14255_; 
wire u2__abc_52155_new_n14256_; 
wire u2__abc_52155_new_n14257_; 
wire u2__abc_52155_new_n14258_; 
wire u2__abc_52155_new_n14259_; 
wire u2__abc_52155_new_n14260_; 
wire u2__abc_52155_new_n14261_; 
wire u2__abc_52155_new_n14262_; 
wire u2__abc_52155_new_n14263_; 
wire u2__abc_52155_new_n14264_; 
wire u2__abc_52155_new_n14265_; 
wire u2__abc_52155_new_n14266_; 
wire u2__abc_52155_new_n14267_; 
wire u2__abc_52155_new_n14268_; 
wire u2__abc_52155_new_n14269_; 
wire u2__abc_52155_new_n14270_; 
wire u2__abc_52155_new_n14272_; 
wire u2__abc_52155_new_n14273_; 
wire u2__abc_52155_new_n14274_; 
wire u2__abc_52155_new_n14275_; 
wire u2__abc_52155_new_n14276_; 
wire u2__abc_52155_new_n14277_; 
wire u2__abc_52155_new_n14278_; 
wire u2__abc_52155_new_n14279_; 
wire u2__abc_52155_new_n14280_; 
wire u2__abc_52155_new_n14281_; 
wire u2__abc_52155_new_n14282_; 
wire u2__abc_52155_new_n14283_; 
wire u2__abc_52155_new_n14284_; 
wire u2__abc_52155_new_n14285_; 
wire u2__abc_52155_new_n14286_; 
wire u2__abc_52155_new_n14287_; 
wire u2__abc_52155_new_n14288_; 
wire u2__abc_52155_new_n14289_; 
wire u2__abc_52155_new_n14291_; 
wire u2__abc_52155_new_n14292_; 
wire u2__abc_52155_new_n14293_; 
wire u2__abc_52155_new_n14294_; 
wire u2__abc_52155_new_n14295_; 
wire u2__abc_52155_new_n14296_; 
wire u2__abc_52155_new_n14297_; 
wire u2__abc_52155_new_n14298_; 
wire u2__abc_52155_new_n14299_; 
wire u2__abc_52155_new_n14300_; 
wire u2__abc_52155_new_n14301_; 
wire u2__abc_52155_new_n14302_; 
wire u2__abc_52155_new_n14303_; 
wire u2__abc_52155_new_n14304_; 
wire u2__abc_52155_new_n14305_; 
wire u2__abc_52155_new_n14306_; 
wire u2__abc_52155_new_n14308_; 
wire u2__abc_52155_new_n14309_; 
wire u2__abc_52155_new_n14310_; 
wire u2__abc_52155_new_n14311_; 
wire u2__abc_52155_new_n14312_; 
wire u2__abc_52155_new_n14313_; 
wire u2__abc_52155_new_n14314_; 
wire u2__abc_52155_new_n14315_; 
wire u2__abc_52155_new_n14316_; 
wire u2__abc_52155_new_n14317_; 
wire u2__abc_52155_new_n14318_; 
wire u2__abc_52155_new_n14319_; 
wire u2__abc_52155_new_n14320_; 
wire u2__abc_52155_new_n14321_; 
wire u2__abc_52155_new_n14322_; 
wire u2__abc_52155_new_n14323_; 
wire u2__abc_52155_new_n14324_; 
wire u2__abc_52155_new_n14325_; 
wire u2__abc_52155_new_n14326_; 
wire u2__abc_52155_new_n14327_; 
wire u2__abc_52155_new_n14328_; 
wire u2__abc_52155_new_n14329_; 
wire u2__abc_52155_new_n14330_; 
wire u2__abc_52155_new_n14332_; 
wire u2__abc_52155_new_n14333_; 
wire u2__abc_52155_new_n14334_; 
wire u2__abc_52155_new_n14335_; 
wire u2__abc_52155_new_n14336_; 
wire u2__abc_52155_new_n14337_; 
wire u2__abc_52155_new_n14338_; 
wire u2__abc_52155_new_n14339_; 
wire u2__abc_52155_new_n14340_; 
wire u2__abc_52155_new_n14341_; 
wire u2__abc_52155_new_n14342_; 
wire u2__abc_52155_new_n14343_; 
wire u2__abc_52155_new_n14344_; 
wire u2__abc_52155_new_n14345_; 
wire u2__abc_52155_new_n14346_; 
wire u2__abc_52155_new_n14347_; 
wire u2__abc_52155_new_n14349_; 
wire u2__abc_52155_new_n14350_; 
wire u2__abc_52155_new_n14351_; 
wire u2__abc_52155_new_n14352_; 
wire u2__abc_52155_new_n14353_; 
wire u2__abc_52155_new_n14354_; 
wire u2__abc_52155_new_n14355_; 
wire u2__abc_52155_new_n14356_; 
wire u2__abc_52155_new_n14357_; 
wire u2__abc_52155_new_n14358_; 
wire u2__abc_52155_new_n14359_; 
wire u2__abc_52155_new_n14360_; 
wire u2__abc_52155_new_n14361_; 
wire u2__abc_52155_new_n14362_; 
wire u2__abc_52155_new_n14363_; 
wire u2__abc_52155_new_n14364_; 
wire u2__abc_52155_new_n14365_; 
wire u2__abc_52155_new_n14366_; 
wire u2__abc_52155_new_n14368_; 
wire u2__abc_52155_new_n14369_; 
wire u2__abc_52155_new_n14370_; 
wire u2__abc_52155_new_n14371_; 
wire u2__abc_52155_new_n14372_; 
wire u2__abc_52155_new_n14373_; 
wire u2__abc_52155_new_n14374_; 
wire u2__abc_52155_new_n14375_; 
wire u2__abc_52155_new_n14376_; 
wire u2__abc_52155_new_n14377_; 
wire u2__abc_52155_new_n14378_; 
wire u2__abc_52155_new_n14379_; 
wire u2__abc_52155_new_n14380_; 
wire u2__abc_52155_new_n14381_; 
wire u2__abc_52155_new_n14382_; 
wire u2__abc_52155_new_n14383_; 
wire u2__abc_52155_new_n14385_; 
wire u2__abc_52155_new_n14386_; 
wire u2__abc_52155_new_n14387_; 
wire u2__abc_52155_new_n14388_; 
wire u2__abc_52155_new_n14389_; 
wire u2__abc_52155_new_n14390_; 
wire u2__abc_52155_new_n14391_; 
wire u2__abc_52155_new_n14392_; 
wire u2__abc_52155_new_n14393_; 
wire u2__abc_52155_new_n14394_; 
wire u2__abc_52155_new_n14395_; 
wire u2__abc_52155_new_n14396_; 
wire u2__abc_52155_new_n14397_; 
wire u2__abc_52155_new_n14398_; 
wire u2__abc_52155_new_n14399_; 
wire u2__abc_52155_new_n14400_; 
wire u2__abc_52155_new_n14401_; 
wire u2__abc_52155_new_n14402_; 
wire u2__abc_52155_new_n14403_; 
wire u2__abc_52155_new_n14404_; 
wire u2__abc_52155_new_n14405_; 
wire u2__abc_52155_new_n14406_; 
wire u2__abc_52155_new_n14407_; 
wire u2__abc_52155_new_n14408_; 
wire u2__abc_52155_new_n14409_; 
wire u2__abc_52155_new_n14410_; 
wire u2__abc_52155_new_n14412_; 
wire u2__abc_52155_new_n14413_; 
wire u2__abc_52155_new_n14414_; 
wire u2__abc_52155_new_n14415_; 
wire u2__abc_52155_new_n14416_; 
wire u2__abc_52155_new_n14417_; 
wire u2__abc_52155_new_n14418_; 
wire u2__abc_52155_new_n14419_; 
wire u2__abc_52155_new_n14420_; 
wire u2__abc_52155_new_n14421_; 
wire u2__abc_52155_new_n14422_; 
wire u2__abc_52155_new_n14423_; 
wire u2__abc_52155_new_n14424_; 
wire u2__abc_52155_new_n14425_; 
wire u2__abc_52155_new_n14426_; 
wire u2__abc_52155_new_n14427_; 
wire u2__abc_52155_new_n14429_; 
wire u2__abc_52155_new_n14430_; 
wire u2__abc_52155_new_n14431_; 
wire u2__abc_52155_new_n14432_; 
wire u2__abc_52155_new_n14433_; 
wire u2__abc_52155_new_n14434_; 
wire u2__abc_52155_new_n14435_; 
wire u2__abc_52155_new_n14436_; 
wire u2__abc_52155_new_n14437_; 
wire u2__abc_52155_new_n14438_; 
wire u2__abc_52155_new_n14439_; 
wire u2__abc_52155_new_n14440_; 
wire u2__abc_52155_new_n14441_; 
wire u2__abc_52155_new_n14442_; 
wire u2__abc_52155_new_n14443_; 
wire u2__abc_52155_new_n14444_; 
wire u2__abc_52155_new_n14445_; 
wire u2__abc_52155_new_n14446_; 
wire u2__abc_52155_new_n14448_; 
wire u2__abc_52155_new_n14449_; 
wire u2__abc_52155_new_n14450_; 
wire u2__abc_52155_new_n14451_; 
wire u2__abc_52155_new_n14452_; 
wire u2__abc_52155_new_n14453_; 
wire u2__abc_52155_new_n14454_; 
wire u2__abc_52155_new_n14455_; 
wire u2__abc_52155_new_n14456_; 
wire u2__abc_52155_new_n14457_; 
wire u2__abc_52155_new_n14458_; 
wire u2__abc_52155_new_n14459_; 
wire u2__abc_52155_new_n14460_; 
wire u2__abc_52155_new_n14461_; 
wire u2__abc_52155_new_n14462_; 
wire u2__abc_52155_new_n14463_; 
wire u2__abc_52155_new_n14465_; 
wire u2__abc_52155_new_n14466_; 
wire u2__abc_52155_new_n14467_; 
wire u2__abc_52155_new_n14468_; 
wire u2__abc_52155_new_n14469_; 
wire u2__abc_52155_new_n14470_; 
wire u2__abc_52155_new_n14471_; 
wire u2__abc_52155_new_n14472_; 
wire u2__abc_52155_new_n14473_; 
wire u2__abc_52155_new_n14474_; 
wire u2__abc_52155_new_n14475_; 
wire u2__abc_52155_new_n14476_; 
wire u2__abc_52155_new_n14477_; 
wire u2__abc_52155_new_n14478_; 
wire u2__abc_52155_new_n14479_; 
wire u2__abc_52155_new_n14480_; 
wire u2__abc_52155_new_n14481_; 
wire u2__abc_52155_new_n14482_; 
wire u2__abc_52155_new_n14483_; 
wire u2__abc_52155_new_n14484_; 
wire u2__abc_52155_new_n14485_; 
wire u2__abc_52155_new_n14486_; 
wire u2__abc_52155_new_n14487_; 
wire u2__abc_52155_new_n14489_; 
wire u2__abc_52155_new_n14490_; 
wire u2__abc_52155_new_n14491_; 
wire u2__abc_52155_new_n14492_; 
wire u2__abc_52155_new_n14493_; 
wire u2__abc_52155_new_n14494_; 
wire u2__abc_52155_new_n14495_; 
wire u2__abc_52155_new_n14496_; 
wire u2__abc_52155_new_n14497_; 
wire u2__abc_52155_new_n14498_; 
wire u2__abc_52155_new_n14499_; 
wire u2__abc_52155_new_n14500_; 
wire u2__abc_52155_new_n14501_; 
wire u2__abc_52155_new_n14502_; 
wire u2__abc_52155_new_n14503_; 
wire u2__abc_52155_new_n14504_; 
wire u2__abc_52155_new_n14506_; 
wire u2__abc_52155_new_n14507_; 
wire u2__abc_52155_new_n14508_; 
wire u2__abc_52155_new_n14509_; 
wire u2__abc_52155_new_n14510_; 
wire u2__abc_52155_new_n14511_; 
wire u2__abc_52155_new_n14512_; 
wire u2__abc_52155_new_n14513_; 
wire u2__abc_52155_new_n14514_; 
wire u2__abc_52155_new_n14515_; 
wire u2__abc_52155_new_n14516_; 
wire u2__abc_52155_new_n14517_; 
wire u2__abc_52155_new_n14518_; 
wire u2__abc_52155_new_n14519_; 
wire u2__abc_52155_new_n14520_; 
wire u2__abc_52155_new_n14521_; 
wire u2__abc_52155_new_n14522_; 
wire u2__abc_52155_new_n14523_; 
wire u2__abc_52155_new_n14525_; 
wire u2__abc_52155_new_n14526_; 
wire u2__abc_52155_new_n14527_; 
wire u2__abc_52155_new_n14528_; 
wire u2__abc_52155_new_n14529_; 
wire u2__abc_52155_new_n14530_; 
wire u2__abc_52155_new_n14531_; 
wire u2__abc_52155_new_n14532_; 
wire u2__abc_52155_new_n14533_; 
wire u2__abc_52155_new_n14534_; 
wire u2__abc_52155_new_n14535_; 
wire u2__abc_52155_new_n14536_; 
wire u2__abc_52155_new_n14537_; 
wire u2__abc_52155_new_n14538_; 
wire u2__abc_52155_new_n14539_; 
wire u2__abc_52155_new_n14540_; 
wire u2__abc_52155_new_n14542_; 
wire u2__abc_52155_new_n14543_; 
wire u2__abc_52155_new_n14544_; 
wire u2__abc_52155_new_n14545_; 
wire u2__abc_52155_new_n14546_; 
wire u2__abc_52155_new_n14547_; 
wire u2__abc_52155_new_n14548_; 
wire u2__abc_52155_new_n14549_; 
wire u2__abc_52155_new_n14550_; 
wire u2__abc_52155_new_n14551_; 
wire u2__abc_52155_new_n14552_; 
wire u2__abc_52155_new_n14553_; 
wire u2__abc_52155_new_n14554_; 
wire u2__abc_52155_new_n14555_; 
wire u2__abc_52155_new_n14556_; 
wire u2__abc_52155_new_n14557_; 
wire u2__abc_52155_new_n14558_; 
wire u2__abc_52155_new_n14559_; 
wire u2__abc_52155_new_n14560_; 
wire u2__abc_52155_new_n14561_; 
wire u2__abc_52155_new_n14562_; 
wire u2__abc_52155_new_n14563_; 
wire u2__abc_52155_new_n14564_; 
wire u2__abc_52155_new_n14565_; 
wire u2__abc_52155_new_n14566_; 
wire u2__abc_52155_new_n14567_; 
wire u2__abc_52155_new_n14568_; 
wire u2__abc_52155_new_n14569_; 
wire u2__abc_52155_new_n14570_; 
wire u2__abc_52155_new_n14571_; 
wire u2__abc_52155_new_n14572_; 
wire u2__abc_52155_new_n14573_; 
wire u2__abc_52155_new_n14575_; 
wire u2__abc_52155_new_n14576_; 
wire u2__abc_52155_new_n14577_; 
wire u2__abc_52155_new_n14578_; 
wire u2__abc_52155_new_n14579_; 
wire u2__abc_52155_new_n14580_; 
wire u2__abc_52155_new_n14581_; 
wire u2__abc_52155_new_n14582_; 
wire u2__abc_52155_new_n14583_; 
wire u2__abc_52155_new_n14584_; 
wire u2__abc_52155_new_n14585_; 
wire u2__abc_52155_new_n14586_; 
wire u2__abc_52155_new_n14587_; 
wire u2__abc_52155_new_n14588_; 
wire u2__abc_52155_new_n14589_; 
wire u2__abc_52155_new_n14590_; 
wire u2__abc_52155_new_n14592_; 
wire u2__abc_52155_new_n14593_; 
wire u2__abc_52155_new_n14594_; 
wire u2__abc_52155_new_n14595_; 
wire u2__abc_52155_new_n14596_; 
wire u2__abc_52155_new_n14597_; 
wire u2__abc_52155_new_n14598_; 
wire u2__abc_52155_new_n14599_; 
wire u2__abc_52155_new_n14600_; 
wire u2__abc_52155_new_n14601_; 
wire u2__abc_52155_new_n14602_; 
wire u2__abc_52155_new_n14603_; 
wire u2__abc_52155_new_n14604_; 
wire u2__abc_52155_new_n14605_; 
wire u2__abc_52155_new_n14606_; 
wire u2__abc_52155_new_n14607_; 
wire u2__abc_52155_new_n14608_; 
wire u2__abc_52155_new_n14609_; 
wire u2__abc_52155_new_n14611_; 
wire u2__abc_52155_new_n14612_; 
wire u2__abc_52155_new_n14613_; 
wire u2__abc_52155_new_n14614_; 
wire u2__abc_52155_new_n14615_; 
wire u2__abc_52155_new_n14616_; 
wire u2__abc_52155_new_n14617_; 
wire u2__abc_52155_new_n14618_; 
wire u2__abc_52155_new_n14619_; 
wire u2__abc_52155_new_n14620_; 
wire u2__abc_52155_new_n14621_; 
wire u2__abc_52155_new_n14622_; 
wire u2__abc_52155_new_n14623_; 
wire u2__abc_52155_new_n14624_; 
wire u2__abc_52155_new_n14625_; 
wire u2__abc_52155_new_n14626_; 
wire u2__abc_52155_new_n14628_; 
wire u2__abc_52155_new_n14629_; 
wire u2__abc_52155_new_n14630_; 
wire u2__abc_52155_new_n14631_; 
wire u2__abc_52155_new_n14632_; 
wire u2__abc_52155_new_n14633_; 
wire u2__abc_52155_new_n14634_; 
wire u2__abc_52155_new_n14635_; 
wire u2__abc_52155_new_n14636_; 
wire u2__abc_52155_new_n14637_; 
wire u2__abc_52155_new_n14638_; 
wire u2__abc_52155_new_n14639_; 
wire u2__abc_52155_new_n14640_; 
wire u2__abc_52155_new_n14641_; 
wire u2__abc_52155_new_n14642_; 
wire u2__abc_52155_new_n14643_; 
wire u2__abc_52155_new_n14644_; 
wire u2__abc_52155_new_n14645_; 
wire u2__abc_52155_new_n14646_; 
wire u2__abc_52155_new_n14647_; 
wire u2__abc_52155_new_n14648_; 
wire u2__abc_52155_new_n14649_; 
wire u2__abc_52155_new_n14650_; 
wire u2__abc_52155_new_n14652_; 
wire u2__abc_52155_new_n14653_; 
wire u2__abc_52155_new_n14654_; 
wire u2__abc_52155_new_n14655_; 
wire u2__abc_52155_new_n14656_; 
wire u2__abc_52155_new_n14657_; 
wire u2__abc_52155_new_n14658_; 
wire u2__abc_52155_new_n14659_; 
wire u2__abc_52155_new_n14660_; 
wire u2__abc_52155_new_n14661_; 
wire u2__abc_52155_new_n14662_; 
wire u2__abc_52155_new_n14663_; 
wire u2__abc_52155_new_n14664_; 
wire u2__abc_52155_new_n14665_; 
wire u2__abc_52155_new_n14666_; 
wire u2__abc_52155_new_n14667_; 
wire u2__abc_52155_new_n14669_; 
wire u2__abc_52155_new_n14670_; 
wire u2__abc_52155_new_n14671_; 
wire u2__abc_52155_new_n14672_; 
wire u2__abc_52155_new_n14673_; 
wire u2__abc_52155_new_n14674_; 
wire u2__abc_52155_new_n14675_; 
wire u2__abc_52155_new_n14676_; 
wire u2__abc_52155_new_n14677_; 
wire u2__abc_52155_new_n14678_; 
wire u2__abc_52155_new_n14679_; 
wire u2__abc_52155_new_n14680_; 
wire u2__abc_52155_new_n14681_; 
wire u2__abc_52155_new_n14682_; 
wire u2__abc_52155_new_n14683_; 
wire u2__abc_52155_new_n14684_; 
wire u2__abc_52155_new_n14685_; 
wire u2__abc_52155_new_n14686_; 
wire u2__abc_52155_new_n14688_; 
wire u2__abc_52155_new_n14689_; 
wire u2__abc_52155_new_n14690_; 
wire u2__abc_52155_new_n14691_; 
wire u2__abc_52155_new_n14692_; 
wire u2__abc_52155_new_n14693_; 
wire u2__abc_52155_new_n14694_; 
wire u2__abc_52155_new_n14695_; 
wire u2__abc_52155_new_n14696_; 
wire u2__abc_52155_new_n14697_; 
wire u2__abc_52155_new_n14698_; 
wire u2__abc_52155_new_n14699_; 
wire u2__abc_52155_new_n14700_; 
wire u2__abc_52155_new_n14701_; 
wire u2__abc_52155_new_n14702_; 
wire u2__abc_52155_new_n14703_; 
wire u2__abc_52155_new_n14705_; 
wire u2__abc_52155_new_n14706_; 
wire u2__abc_52155_new_n14707_; 
wire u2__abc_52155_new_n14708_; 
wire u2__abc_52155_new_n14709_; 
wire u2__abc_52155_new_n14710_; 
wire u2__abc_52155_new_n14711_; 
wire u2__abc_52155_new_n14712_; 
wire u2__abc_52155_new_n14713_; 
wire u2__abc_52155_new_n14714_; 
wire u2__abc_52155_new_n14715_; 
wire u2__abc_52155_new_n14716_; 
wire u2__abc_52155_new_n14717_; 
wire u2__abc_52155_new_n14718_; 
wire u2__abc_52155_new_n14719_; 
wire u2__abc_52155_new_n14720_; 
wire u2__abc_52155_new_n14721_; 
wire u2__abc_52155_new_n14722_; 
wire u2__abc_52155_new_n14723_; 
wire u2__abc_52155_new_n14724_; 
wire u2__abc_52155_new_n14725_; 
wire u2__abc_52155_new_n14726_; 
wire u2__abc_52155_new_n14727_; 
wire u2__abc_52155_new_n14728_; 
wire u2__abc_52155_new_n14729_; 
wire u2__abc_52155_new_n14730_; 
wire u2__abc_52155_new_n14732_; 
wire u2__abc_52155_new_n14733_; 
wire u2__abc_52155_new_n14734_; 
wire u2__abc_52155_new_n14735_; 
wire u2__abc_52155_new_n14736_; 
wire u2__abc_52155_new_n14737_; 
wire u2__abc_52155_new_n14738_; 
wire u2__abc_52155_new_n14739_; 
wire u2__abc_52155_new_n14740_; 
wire u2__abc_52155_new_n14741_; 
wire u2__abc_52155_new_n14742_; 
wire u2__abc_52155_new_n14743_; 
wire u2__abc_52155_new_n14744_; 
wire u2__abc_52155_new_n14745_; 
wire u2__abc_52155_new_n14746_; 
wire u2__abc_52155_new_n14747_; 
wire u2__abc_52155_new_n14749_; 
wire u2__abc_52155_new_n14750_; 
wire u2__abc_52155_new_n14751_; 
wire u2__abc_52155_new_n14752_; 
wire u2__abc_52155_new_n14753_; 
wire u2__abc_52155_new_n14754_; 
wire u2__abc_52155_new_n14755_; 
wire u2__abc_52155_new_n14756_; 
wire u2__abc_52155_new_n14757_; 
wire u2__abc_52155_new_n14758_; 
wire u2__abc_52155_new_n14759_; 
wire u2__abc_52155_new_n14760_; 
wire u2__abc_52155_new_n14761_; 
wire u2__abc_52155_new_n14762_; 
wire u2__abc_52155_new_n14763_; 
wire u2__abc_52155_new_n14764_; 
wire u2__abc_52155_new_n14765_; 
wire u2__abc_52155_new_n14766_; 
wire u2__abc_52155_new_n14767_; 
wire u2__abc_52155_new_n14769_; 
wire u2__abc_52155_new_n14770_; 
wire u2__abc_52155_new_n14771_; 
wire u2__abc_52155_new_n14772_; 
wire u2__abc_52155_new_n14773_; 
wire u2__abc_52155_new_n14774_; 
wire u2__abc_52155_new_n14775_; 
wire u2__abc_52155_new_n14776_; 
wire u2__abc_52155_new_n14777_; 
wire u2__abc_52155_new_n14778_; 
wire u2__abc_52155_new_n14779_; 
wire u2__abc_52155_new_n14780_; 
wire u2__abc_52155_new_n14781_; 
wire u2__abc_52155_new_n14782_; 
wire u2__abc_52155_new_n14783_; 
wire u2__abc_52155_new_n14784_; 
wire u2__abc_52155_new_n14786_; 
wire u2__abc_52155_new_n14787_; 
wire u2__abc_52155_new_n14788_; 
wire u2__abc_52155_new_n14789_; 
wire u2__abc_52155_new_n14790_; 
wire u2__abc_52155_new_n14791_; 
wire u2__abc_52155_new_n14792_; 
wire u2__abc_52155_new_n14793_; 
wire u2__abc_52155_new_n14794_; 
wire u2__abc_52155_new_n14795_; 
wire u2__abc_52155_new_n14796_; 
wire u2__abc_52155_new_n14797_; 
wire u2__abc_52155_new_n14798_; 
wire u2__abc_52155_new_n14799_; 
wire u2__abc_52155_new_n14800_; 
wire u2__abc_52155_new_n14801_; 
wire u2__abc_52155_new_n14802_; 
wire u2__abc_52155_new_n14803_; 
wire u2__abc_52155_new_n14804_; 
wire u2__abc_52155_new_n14805_; 
wire u2__abc_52155_new_n14807_; 
wire u2__abc_52155_new_n14808_; 
wire u2__abc_52155_new_n14809_; 
wire u2__abc_52155_new_n14810_; 
wire u2__abc_52155_new_n14811_; 
wire u2__abc_52155_new_n14812_; 
wire u2__abc_52155_new_n14813_; 
wire u2__abc_52155_new_n14814_; 
wire u2__abc_52155_new_n14815_; 
wire u2__abc_52155_new_n14816_; 
wire u2__abc_52155_new_n14817_; 
wire u2__abc_52155_new_n14818_; 
wire u2__abc_52155_new_n14819_; 
wire u2__abc_52155_new_n14820_; 
wire u2__abc_52155_new_n14821_; 
wire u2__abc_52155_new_n14822_; 
wire u2__abc_52155_new_n14824_; 
wire u2__abc_52155_new_n14825_; 
wire u2__abc_52155_new_n14826_; 
wire u2__abc_52155_new_n14827_; 
wire u2__abc_52155_new_n14828_; 
wire u2__abc_52155_new_n14829_; 
wire u2__abc_52155_new_n14830_; 
wire u2__abc_52155_new_n14831_; 
wire u2__abc_52155_new_n14832_; 
wire u2__abc_52155_new_n14833_; 
wire u2__abc_52155_new_n14834_; 
wire u2__abc_52155_new_n14835_; 
wire u2__abc_52155_new_n14836_; 
wire u2__abc_52155_new_n14837_; 
wire u2__abc_52155_new_n14838_; 
wire u2__abc_52155_new_n14839_; 
wire u2__abc_52155_new_n14840_; 
wire u2__abc_52155_new_n14841_; 
wire u2__abc_52155_new_n14843_; 
wire u2__abc_52155_new_n14844_; 
wire u2__abc_52155_new_n14845_; 
wire u2__abc_52155_new_n14846_; 
wire u2__abc_52155_new_n14847_; 
wire u2__abc_52155_new_n14848_; 
wire u2__abc_52155_new_n14849_; 
wire u2__abc_52155_new_n14850_; 
wire u2__abc_52155_new_n14851_; 
wire u2__abc_52155_new_n14852_; 
wire u2__abc_52155_new_n14853_; 
wire u2__abc_52155_new_n14854_; 
wire u2__abc_52155_new_n14855_; 
wire u2__abc_52155_new_n14856_; 
wire u2__abc_52155_new_n14857_; 
wire u2__abc_52155_new_n14858_; 
wire u2__abc_52155_new_n14860_; 
wire u2__abc_52155_new_n14861_; 
wire u2__abc_52155_new_n14862_; 
wire u2__abc_52155_new_n14863_; 
wire u2__abc_52155_new_n14864_; 
wire u2__abc_52155_new_n14865_; 
wire u2__abc_52155_new_n14866_; 
wire u2__abc_52155_new_n14867_; 
wire u2__abc_52155_new_n14868_; 
wire u2__abc_52155_new_n14869_; 
wire u2__abc_52155_new_n14870_; 
wire u2__abc_52155_new_n14871_; 
wire u2__abc_52155_new_n14872_; 
wire u2__abc_52155_new_n14873_; 
wire u2__abc_52155_new_n14874_; 
wire u2__abc_52155_new_n14875_; 
wire u2__abc_52155_new_n14876_; 
wire u2__abc_52155_new_n14877_; 
wire u2__abc_52155_new_n14878_; 
wire u2__abc_52155_new_n14879_; 
wire u2__abc_52155_new_n14880_; 
wire u2__abc_52155_new_n14881_; 
wire u2__abc_52155_new_n14882_; 
wire u2__abc_52155_new_n14883_; 
wire u2__abc_52155_new_n14884_; 
wire u2__abc_52155_new_n14885_; 
wire u2__abc_52155_new_n14886_; 
wire u2__abc_52155_new_n14887_; 
wire u2__abc_52155_new_n14888_; 
wire u2__abc_52155_new_n14889_; 
wire u2__abc_52155_new_n14891_; 
wire u2__abc_52155_new_n14892_; 
wire u2__abc_52155_new_n14893_; 
wire u2__abc_52155_new_n14894_; 
wire u2__abc_52155_new_n14895_; 
wire u2__abc_52155_new_n14896_; 
wire u2__abc_52155_new_n14897_; 
wire u2__abc_52155_new_n14898_; 
wire u2__abc_52155_new_n14899_; 
wire u2__abc_52155_new_n14900_; 
wire u2__abc_52155_new_n14901_; 
wire u2__abc_52155_new_n14902_; 
wire u2__abc_52155_new_n14903_; 
wire u2__abc_52155_new_n14904_; 
wire u2__abc_52155_new_n14905_; 
wire u2__abc_52155_new_n14906_; 
wire u2__abc_52155_new_n14908_; 
wire u2__abc_52155_new_n14909_; 
wire u2__abc_52155_new_n14910_; 
wire u2__abc_52155_new_n14911_; 
wire u2__abc_52155_new_n14912_; 
wire u2__abc_52155_new_n14913_; 
wire u2__abc_52155_new_n14914_; 
wire u2__abc_52155_new_n14915_; 
wire u2__abc_52155_new_n14916_; 
wire u2__abc_52155_new_n14917_; 
wire u2__abc_52155_new_n14918_; 
wire u2__abc_52155_new_n14919_; 
wire u2__abc_52155_new_n14920_; 
wire u2__abc_52155_new_n14921_; 
wire u2__abc_52155_new_n14922_; 
wire u2__abc_52155_new_n14923_; 
wire u2__abc_52155_new_n14924_; 
wire u2__abc_52155_new_n14925_; 
wire u2__abc_52155_new_n14927_; 
wire u2__abc_52155_new_n14928_; 
wire u2__abc_52155_new_n14929_; 
wire u2__abc_52155_new_n14930_; 
wire u2__abc_52155_new_n14931_; 
wire u2__abc_52155_new_n14932_; 
wire u2__abc_52155_new_n14933_; 
wire u2__abc_52155_new_n14934_; 
wire u2__abc_52155_new_n14935_; 
wire u2__abc_52155_new_n14936_; 
wire u2__abc_52155_new_n14937_; 
wire u2__abc_52155_new_n14938_; 
wire u2__abc_52155_new_n14939_; 
wire u2__abc_52155_new_n14940_; 
wire u2__abc_52155_new_n14941_; 
wire u2__abc_52155_new_n14942_; 
wire u2__abc_52155_new_n14944_; 
wire u2__abc_52155_new_n14945_; 
wire u2__abc_52155_new_n14946_; 
wire u2__abc_52155_new_n14947_; 
wire u2__abc_52155_new_n14948_; 
wire u2__abc_52155_new_n14949_; 
wire u2__abc_52155_new_n14950_; 
wire u2__abc_52155_new_n14951_; 
wire u2__abc_52155_new_n14952_; 
wire u2__abc_52155_new_n14953_; 
wire u2__abc_52155_new_n14954_; 
wire u2__abc_52155_new_n14955_; 
wire u2__abc_52155_new_n14956_; 
wire u2__abc_52155_new_n14957_; 
wire u2__abc_52155_new_n14958_; 
wire u2__abc_52155_new_n14959_; 
wire u2__abc_52155_new_n14960_; 
wire u2__abc_52155_new_n14961_; 
wire u2__abc_52155_new_n14962_; 
wire u2__abc_52155_new_n14963_; 
wire u2__abc_52155_new_n14964_; 
wire u2__abc_52155_new_n14965_; 
wire u2__abc_52155_new_n14966_; 
wire u2__abc_52155_new_n14968_; 
wire u2__abc_52155_new_n14969_; 
wire u2__abc_52155_new_n14970_; 
wire u2__abc_52155_new_n14971_; 
wire u2__abc_52155_new_n14972_; 
wire u2__abc_52155_new_n14973_; 
wire u2__abc_52155_new_n14974_; 
wire u2__abc_52155_new_n14975_; 
wire u2__abc_52155_new_n14976_; 
wire u2__abc_52155_new_n14977_; 
wire u2__abc_52155_new_n14978_; 
wire u2__abc_52155_new_n14979_; 
wire u2__abc_52155_new_n14980_; 
wire u2__abc_52155_new_n14981_; 
wire u2__abc_52155_new_n14982_; 
wire u2__abc_52155_new_n14983_; 
wire u2__abc_52155_new_n14985_; 
wire u2__abc_52155_new_n14986_; 
wire u2__abc_52155_new_n14987_; 
wire u2__abc_52155_new_n14988_; 
wire u2__abc_52155_new_n14989_; 
wire u2__abc_52155_new_n14990_; 
wire u2__abc_52155_new_n14991_; 
wire u2__abc_52155_new_n14992_; 
wire u2__abc_52155_new_n14993_; 
wire u2__abc_52155_new_n14994_; 
wire u2__abc_52155_new_n14995_; 
wire u2__abc_52155_new_n14996_; 
wire u2__abc_52155_new_n14997_; 
wire u2__abc_52155_new_n14998_; 
wire u2__abc_52155_new_n14999_; 
wire u2__abc_52155_new_n15000_; 
wire u2__abc_52155_new_n15002_; 
wire u2__abc_52155_new_n15003_; 
wire u2__abc_52155_new_n15004_; 
wire u2__abc_52155_new_n15005_; 
wire u2__abc_52155_new_n15006_; 
wire u2__abc_52155_new_n15007_; 
wire u2__abc_52155_new_n15008_; 
wire u2__abc_52155_new_n15009_; 
wire u2__abc_52155_new_n15010_; 
wire u2__abc_52155_new_n15011_; 
wire u2__abc_52155_new_n15012_; 
wire u2__abc_52155_new_n15013_; 
wire u2__abc_52155_new_n15014_; 
wire u2__abc_52155_new_n15015_; 
wire u2__abc_52155_new_n15016_; 
wire u2__abc_52155_new_n15017_; 
wire u2__abc_52155_new_n15019_; 
wire u2__abc_52155_new_n15020_; 
wire u2__abc_52155_new_n15021_; 
wire u2__abc_52155_new_n15022_; 
wire u2__abc_52155_new_n15023_; 
wire u2__abc_52155_new_n15024_; 
wire u2__abc_52155_new_n15025_; 
wire u2__abc_52155_new_n15026_; 
wire u2__abc_52155_new_n15027_; 
wire u2__abc_52155_new_n15028_; 
wire u2__abc_52155_new_n15029_; 
wire u2__abc_52155_new_n15030_; 
wire u2__abc_52155_new_n15031_; 
wire u2__abc_52155_new_n15032_; 
wire u2__abc_52155_new_n15033_; 
wire u2__abc_52155_new_n15034_; 
wire u2__abc_52155_new_n15035_; 
wire u2__abc_52155_new_n15036_; 
wire u2__abc_52155_new_n15037_; 
wire u2__abc_52155_new_n15038_; 
wire u2__abc_52155_new_n15039_; 
wire u2__abc_52155_new_n15040_; 
wire u2__abc_52155_new_n15041_; 
wire u2__abc_52155_new_n15042_; 
wire u2__abc_52155_new_n15044_; 
wire u2__abc_52155_new_n15045_; 
wire u2__abc_52155_new_n15046_; 
wire u2__abc_52155_new_n15047_; 
wire u2__abc_52155_new_n15048_; 
wire u2__abc_52155_new_n15049_; 
wire u2__abc_52155_new_n15050_; 
wire u2__abc_52155_new_n15051_; 
wire u2__abc_52155_new_n15052_; 
wire u2__abc_52155_new_n15053_; 
wire u2__abc_52155_new_n15054_; 
wire u2__abc_52155_new_n15055_; 
wire u2__abc_52155_new_n15056_; 
wire u2__abc_52155_new_n15057_; 
wire u2__abc_52155_new_n15058_; 
wire u2__abc_52155_new_n15059_; 
wire u2__abc_52155_new_n15061_; 
wire u2__abc_52155_new_n15062_; 
wire u2__abc_52155_new_n15063_; 
wire u2__abc_52155_new_n15064_; 
wire u2__abc_52155_new_n15065_; 
wire u2__abc_52155_new_n15066_; 
wire u2__abc_52155_new_n15067_; 
wire u2__abc_52155_new_n15068_; 
wire u2__abc_52155_new_n15069_; 
wire u2__abc_52155_new_n15070_; 
wire u2__abc_52155_new_n15071_; 
wire u2__abc_52155_new_n15072_; 
wire u2__abc_52155_new_n15073_; 
wire u2__abc_52155_new_n15074_; 
wire u2__abc_52155_new_n15075_; 
wire u2__abc_52155_new_n15076_; 
wire u2__abc_52155_new_n15077_; 
wire u2__abc_52155_new_n15078_; 
wire u2__abc_52155_new_n15079_; 
wire u2__abc_52155_new_n15081_; 
wire u2__abc_52155_new_n15082_; 
wire u2__abc_52155_new_n15083_; 
wire u2__abc_52155_new_n15084_; 
wire u2__abc_52155_new_n15085_; 
wire u2__abc_52155_new_n15086_; 
wire u2__abc_52155_new_n15087_; 
wire u2__abc_52155_new_n15088_; 
wire u2__abc_52155_new_n15089_; 
wire u2__abc_52155_new_n15090_; 
wire u2__abc_52155_new_n15091_; 
wire u2__abc_52155_new_n15092_; 
wire u2__abc_52155_new_n15093_; 
wire u2__abc_52155_new_n15094_; 
wire u2__abc_52155_new_n15095_; 
wire u2__abc_52155_new_n15096_; 
wire u2__abc_52155_new_n15098_; 
wire u2__abc_52155_new_n15099_; 
wire u2__abc_52155_new_n15100_; 
wire u2__abc_52155_new_n15101_; 
wire u2__abc_52155_new_n15102_; 
wire u2__abc_52155_new_n15103_; 
wire u2__abc_52155_new_n15104_; 
wire u2__abc_52155_new_n15105_; 
wire u2__abc_52155_new_n15106_; 
wire u2__abc_52155_new_n15107_; 
wire u2__abc_52155_new_n15108_; 
wire u2__abc_52155_new_n15109_; 
wire u2__abc_52155_new_n15110_; 
wire u2__abc_52155_new_n15111_; 
wire u2__abc_52155_new_n15112_; 
wire u2__abc_52155_new_n15113_; 
wire u2__abc_52155_new_n15114_; 
wire u2__abc_52155_new_n15115_; 
wire u2__abc_52155_new_n15117_; 
wire u2__abc_52155_new_n15118_; 
wire u2__abc_52155_new_n15119_; 
wire u2__abc_52155_new_n15120_; 
wire u2__abc_52155_new_n15121_; 
wire u2__abc_52155_new_n15122_; 
wire u2__abc_52155_new_n15123_; 
wire u2__abc_52155_new_n15124_; 
wire u2__abc_52155_new_n15125_; 
wire u2__abc_52155_new_n15126_; 
wire u2__abc_52155_new_n15127_; 
wire u2__abc_52155_new_n15128_; 
wire u2__abc_52155_new_n15129_; 
wire u2__abc_52155_new_n15130_; 
wire u2__abc_52155_new_n15131_; 
wire u2__abc_52155_new_n15132_; 
wire u2__abc_52155_new_n15134_; 
wire u2__abc_52155_new_n15135_; 
wire u2__abc_52155_new_n15136_; 
wire u2__abc_52155_new_n15137_; 
wire u2__abc_52155_new_n15138_; 
wire u2__abc_52155_new_n15139_; 
wire u2__abc_52155_new_n15140_; 
wire u2__abc_52155_new_n15141_; 
wire u2__abc_52155_new_n15142_; 
wire u2__abc_52155_new_n15143_; 
wire u2__abc_52155_new_n15144_; 
wire u2__abc_52155_new_n15145_; 
wire u2__abc_52155_new_n15146_; 
wire u2__abc_52155_new_n15147_; 
wire u2__abc_52155_new_n15148_; 
wire u2__abc_52155_new_n15149_; 
wire u2__abc_52155_new_n15150_; 
wire u2__abc_52155_new_n15151_; 
wire u2__abc_52155_new_n15153_; 
wire u2__abc_52155_new_n15154_; 
wire u2__abc_52155_new_n15155_; 
wire u2__abc_52155_new_n15156_; 
wire u2__abc_52155_new_n15157_; 
wire u2__abc_52155_new_n15158_; 
wire u2__abc_52155_new_n15159_; 
wire u2__abc_52155_new_n15160_; 
wire u2__abc_52155_new_n15161_; 
wire u2__abc_52155_new_n15162_; 
wire u2__abc_52155_new_n15163_; 
wire u2__abc_52155_new_n15164_; 
wire u2__abc_52155_new_n15165_; 
wire u2__abc_52155_new_n15166_; 
wire u2__abc_52155_new_n15167_; 
wire u2__abc_52155_new_n15168_; 
wire u2__abc_52155_new_n15170_; 
wire u2__abc_52155_new_n15171_; 
wire u2__abc_52155_new_n15172_; 
wire u2__abc_52155_new_n15173_; 
wire u2__abc_52155_new_n15174_; 
wire u2__abc_52155_new_n15175_; 
wire u2__abc_52155_new_n15176_; 
wire u2__abc_52155_new_n15177_; 
wire u2__abc_52155_new_n15178_; 
wire u2__abc_52155_new_n15179_; 
wire u2__abc_52155_new_n15180_; 
wire u2__abc_52155_new_n15181_; 
wire u2__abc_52155_new_n15182_; 
wire u2__abc_52155_new_n15183_; 
wire u2__abc_52155_new_n15184_; 
wire u2__abc_52155_new_n15185_; 
wire u2__abc_52155_new_n15186_; 
wire u2__abc_52155_new_n15187_; 
wire u2__abc_52155_new_n15188_; 
wire u2__abc_52155_new_n15189_; 
wire u2__abc_52155_new_n15190_; 
wire u2__abc_52155_new_n15191_; 
wire u2__abc_52155_new_n15192_; 
wire u2__abc_52155_new_n15193_; 
wire u2__abc_52155_new_n15194_; 
wire u2__abc_52155_new_n15195_; 
wire u2__abc_52155_new_n15196_; 
wire u2__abc_52155_new_n15197_; 
wire u2__abc_52155_new_n15198_; 
wire u2__abc_52155_new_n15199_; 
wire u2__abc_52155_new_n15200_; 
wire u2__abc_52155_new_n15201_; 
wire u2__abc_52155_new_n15202_; 
wire u2__abc_52155_new_n15203_; 
wire u2__abc_52155_new_n15204_; 
wire u2__abc_52155_new_n15205_; 
wire u2__abc_52155_new_n15206_; 
wire u2__abc_52155_new_n15207_; 
wire u2__abc_52155_new_n15208_; 
wire u2__abc_52155_new_n15209_; 
wire u2__abc_52155_new_n15210_; 
wire u2__abc_52155_new_n15212_; 
wire u2__abc_52155_new_n15213_; 
wire u2__abc_52155_new_n15214_; 
wire u2__abc_52155_new_n15215_; 
wire u2__abc_52155_new_n15216_; 
wire u2__abc_52155_new_n15217_; 
wire u2__abc_52155_new_n15218_; 
wire u2__abc_52155_new_n15219_; 
wire u2__abc_52155_new_n15220_; 
wire u2__abc_52155_new_n15221_; 
wire u2__abc_52155_new_n15222_; 
wire u2__abc_52155_new_n15223_; 
wire u2__abc_52155_new_n15224_; 
wire u2__abc_52155_new_n15225_; 
wire u2__abc_52155_new_n15226_; 
wire u2__abc_52155_new_n15227_; 
wire u2__abc_52155_new_n15229_; 
wire u2__abc_52155_new_n15230_; 
wire u2__abc_52155_new_n15231_; 
wire u2__abc_52155_new_n15232_; 
wire u2__abc_52155_new_n15233_; 
wire u2__abc_52155_new_n15234_; 
wire u2__abc_52155_new_n15235_; 
wire u2__abc_52155_new_n15236_; 
wire u2__abc_52155_new_n15237_; 
wire u2__abc_52155_new_n15238_; 
wire u2__abc_52155_new_n15239_; 
wire u2__abc_52155_new_n15240_; 
wire u2__abc_52155_new_n15241_; 
wire u2__abc_52155_new_n15242_; 
wire u2__abc_52155_new_n15243_; 
wire u2__abc_52155_new_n15244_; 
wire u2__abc_52155_new_n15245_; 
wire u2__abc_52155_new_n15246_; 
wire u2__abc_52155_new_n15248_; 
wire u2__abc_52155_new_n15249_; 
wire u2__abc_52155_new_n15250_; 
wire u2__abc_52155_new_n15251_; 
wire u2__abc_52155_new_n15252_; 
wire u2__abc_52155_new_n15253_; 
wire u2__abc_52155_new_n15254_; 
wire u2__abc_52155_new_n15255_; 
wire u2__abc_52155_new_n15256_; 
wire u2__abc_52155_new_n15257_; 
wire u2__abc_52155_new_n15258_; 
wire u2__abc_52155_new_n15259_; 
wire u2__abc_52155_new_n15260_; 
wire u2__abc_52155_new_n15261_; 
wire u2__abc_52155_new_n15262_; 
wire u2__abc_52155_new_n15263_; 
wire u2__abc_52155_new_n15265_; 
wire u2__abc_52155_new_n15266_; 
wire u2__abc_52155_new_n15267_; 
wire u2__abc_52155_new_n15268_; 
wire u2__abc_52155_new_n15269_; 
wire u2__abc_52155_new_n15270_; 
wire u2__abc_52155_new_n15271_; 
wire u2__abc_52155_new_n15272_; 
wire u2__abc_52155_new_n15273_; 
wire u2__abc_52155_new_n15274_; 
wire u2__abc_52155_new_n15275_; 
wire u2__abc_52155_new_n15276_; 
wire u2__abc_52155_new_n15277_; 
wire u2__abc_52155_new_n15278_; 
wire u2__abc_52155_new_n15279_; 
wire u2__abc_52155_new_n15280_; 
wire u2__abc_52155_new_n15281_; 
wire u2__abc_52155_new_n15282_; 
wire u2__abc_52155_new_n15283_; 
wire u2__abc_52155_new_n15284_; 
wire u2__abc_52155_new_n15285_; 
wire u2__abc_52155_new_n15286_; 
wire u2__abc_52155_new_n15288_; 
wire u2__abc_52155_new_n15289_; 
wire u2__abc_52155_new_n15290_; 
wire u2__abc_52155_new_n15291_; 
wire u2__abc_52155_new_n15292_; 
wire u2__abc_52155_new_n15293_; 
wire u2__abc_52155_new_n15294_; 
wire u2__abc_52155_new_n15295_; 
wire u2__abc_52155_new_n15296_; 
wire u2__abc_52155_new_n15297_; 
wire u2__abc_52155_new_n15298_; 
wire u2__abc_52155_new_n15299_; 
wire u2__abc_52155_new_n15300_; 
wire u2__abc_52155_new_n15301_; 
wire u2__abc_52155_new_n15302_; 
wire u2__abc_52155_new_n15303_; 
wire u2__abc_52155_new_n15305_; 
wire u2__abc_52155_new_n15306_; 
wire u2__abc_52155_new_n15307_; 
wire u2__abc_52155_new_n15308_; 
wire u2__abc_52155_new_n15309_; 
wire u2__abc_52155_new_n15310_; 
wire u2__abc_52155_new_n15311_; 
wire u2__abc_52155_new_n15312_; 
wire u2__abc_52155_new_n15313_; 
wire u2__abc_52155_new_n15314_; 
wire u2__abc_52155_new_n15315_; 
wire u2__abc_52155_new_n15316_; 
wire u2__abc_52155_new_n15317_; 
wire u2__abc_52155_new_n15318_; 
wire u2__abc_52155_new_n15319_; 
wire u2__abc_52155_new_n15320_; 
wire u2__abc_52155_new_n15321_; 
wire u2__abc_52155_new_n15322_; 
wire u2__abc_52155_new_n15324_; 
wire u2__abc_52155_new_n15325_; 
wire u2__abc_52155_new_n15326_; 
wire u2__abc_52155_new_n15327_; 
wire u2__abc_52155_new_n15328_; 
wire u2__abc_52155_new_n15329_; 
wire u2__abc_52155_new_n15330_; 
wire u2__abc_52155_new_n15331_; 
wire u2__abc_52155_new_n15332_; 
wire u2__abc_52155_new_n15333_; 
wire u2__abc_52155_new_n15334_; 
wire u2__abc_52155_new_n15335_; 
wire u2__abc_52155_new_n15336_; 
wire u2__abc_52155_new_n15337_; 
wire u2__abc_52155_new_n15338_; 
wire u2__abc_52155_new_n15339_; 
wire u2__abc_52155_new_n15341_; 
wire u2__abc_52155_new_n15342_; 
wire u2__abc_52155_new_n15343_; 
wire u2__abc_52155_new_n15344_; 
wire u2__abc_52155_new_n15345_; 
wire u2__abc_52155_new_n15346_; 
wire u2__abc_52155_new_n15347_; 
wire u2__abc_52155_new_n15348_; 
wire u2__abc_52155_new_n15349_; 
wire u2__abc_52155_new_n15350_; 
wire u2__abc_52155_new_n15351_; 
wire u2__abc_52155_new_n15352_; 
wire u2__abc_52155_new_n15353_; 
wire u2__abc_52155_new_n15354_; 
wire u2__abc_52155_new_n15355_; 
wire u2__abc_52155_new_n15356_; 
wire u2__abc_52155_new_n15357_; 
wire u2__abc_52155_new_n15358_; 
wire u2__abc_52155_new_n15359_; 
wire u2__abc_52155_new_n15360_; 
wire u2__abc_52155_new_n15361_; 
wire u2__abc_52155_new_n15362_; 
wire u2__abc_52155_new_n15363_; 
wire u2__abc_52155_new_n15364_; 
wire u2__abc_52155_new_n15366_; 
wire u2__abc_52155_new_n15367_; 
wire u2__abc_52155_new_n15368_; 
wire u2__abc_52155_new_n15369_; 
wire u2__abc_52155_new_n15370_; 
wire u2__abc_52155_new_n15371_; 
wire u2__abc_52155_new_n15372_; 
wire u2__abc_52155_new_n15373_; 
wire u2__abc_52155_new_n15374_; 
wire u2__abc_52155_new_n15375_; 
wire u2__abc_52155_new_n15376_; 
wire u2__abc_52155_new_n15377_; 
wire u2__abc_52155_new_n15378_; 
wire u2__abc_52155_new_n15379_; 
wire u2__abc_52155_new_n15380_; 
wire u2__abc_52155_new_n15381_; 
wire u2__abc_52155_new_n15383_; 
wire u2__abc_52155_new_n15384_; 
wire u2__abc_52155_new_n15385_; 
wire u2__abc_52155_new_n15386_; 
wire u2__abc_52155_new_n15387_; 
wire u2__abc_52155_new_n15388_; 
wire u2__abc_52155_new_n15389_; 
wire u2__abc_52155_new_n15390_; 
wire u2__abc_52155_new_n15391_; 
wire u2__abc_52155_new_n15392_; 
wire u2__abc_52155_new_n15393_; 
wire u2__abc_52155_new_n15394_; 
wire u2__abc_52155_new_n15395_; 
wire u2__abc_52155_new_n15396_; 
wire u2__abc_52155_new_n15397_; 
wire u2__abc_52155_new_n15398_; 
wire u2__abc_52155_new_n15400_; 
wire u2__abc_52155_new_n15401_; 
wire u2__abc_52155_new_n15402_; 
wire u2__abc_52155_new_n15403_; 
wire u2__abc_52155_new_n15404_; 
wire u2__abc_52155_new_n15405_; 
wire u2__abc_52155_new_n15406_; 
wire u2__abc_52155_new_n15407_; 
wire u2__abc_52155_new_n15408_; 
wire u2__abc_52155_new_n15409_; 
wire u2__abc_52155_new_n15410_; 
wire u2__abc_52155_new_n15411_; 
wire u2__abc_52155_new_n15412_; 
wire u2__abc_52155_new_n15413_; 
wire u2__abc_52155_new_n15414_; 
wire u2__abc_52155_new_n15415_; 
wire u2__abc_52155_new_n15417_; 
wire u2__abc_52155_new_n15418_; 
wire u2__abc_52155_new_n15419_; 
wire u2__abc_52155_new_n15420_; 
wire u2__abc_52155_new_n15421_; 
wire u2__abc_52155_new_n15422_; 
wire u2__abc_52155_new_n15423_; 
wire u2__abc_52155_new_n15424_; 
wire u2__abc_52155_new_n15425_; 
wire u2__abc_52155_new_n15426_; 
wire u2__abc_52155_new_n15427_; 
wire u2__abc_52155_new_n15428_; 
wire u2__abc_52155_new_n15429_; 
wire u2__abc_52155_new_n15430_; 
wire u2__abc_52155_new_n15431_; 
wire u2__abc_52155_new_n15432_; 
wire u2__abc_52155_new_n15433_; 
wire u2__abc_52155_new_n15434_; 
wire u2__abc_52155_new_n15435_; 
wire u2__abc_52155_new_n15436_; 
wire u2__abc_52155_new_n15437_; 
wire u2__abc_52155_new_n15438_; 
wire u2__abc_52155_new_n15439_; 
wire u2__abc_52155_new_n15441_; 
wire u2__abc_52155_new_n15442_; 
wire u2__abc_52155_new_n15443_; 
wire u2__abc_52155_new_n15444_; 
wire u2__abc_52155_new_n15445_; 
wire u2__abc_52155_new_n15446_; 
wire u2__abc_52155_new_n15447_; 
wire u2__abc_52155_new_n15448_; 
wire u2__abc_52155_new_n15449_; 
wire u2__abc_52155_new_n15450_; 
wire u2__abc_52155_new_n15451_; 
wire u2__abc_52155_new_n15452_; 
wire u2__abc_52155_new_n15453_; 
wire u2__abc_52155_new_n15454_; 
wire u2__abc_52155_new_n15455_; 
wire u2__abc_52155_new_n15456_; 
wire u2__abc_52155_new_n15458_; 
wire u2__abc_52155_new_n15459_; 
wire u2__abc_52155_new_n15460_; 
wire u2__abc_52155_new_n15461_; 
wire u2__abc_52155_new_n15462_; 
wire u2__abc_52155_new_n15463_; 
wire u2__abc_52155_new_n15464_; 
wire u2__abc_52155_new_n15465_; 
wire u2__abc_52155_new_n15466_; 
wire u2__abc_52155_new_n15467_; 
wire u2__abc_52155_new_n15468_; 
wire u2__abc_52155_new_n15469_; 
wire u2__abc_52155_new_n15470_; 
wire u2__abc_52155_new_n15471_; 
wire u2__abc_52155_new_n15472_; 
wire u2__abc_52155_new_n15473_; 
wire u2__abc_52155_new_n15474_; 
wire u2__abc_52155_new_n15475_; 
wire u2__abc_52155_new_n15477_; 
wire u2__abc_52155_new_n15478_; 
wire u2__abc_52155_new_n15479_; 
wire u2__abc_52155_new_n15480_; 
wire u2__abc_52155_new_n15481_; 
wire u2__abc_52155_new_n15482_; 
wire u2__abc_52155_new_n15483_; 
wire u2__abc_52155_new_n15484_; 
wire u2__abc_52155_new_n15485_; 
wire u2__abc_52155_new_n15486_; 
wire u2__abc_52155_new_n15487_; 
wire u2__abc_52155_new_n15488_; 
wire u2__abc_52155_new_n15489_; 
wire u2__abc_52155_new_n15490_; 
wire u2__abc_52155_new_n15491_; 
wire u2__abc_52155_new_n15492_; 
wire u2__abc_52155_new_n15494_; 
wire u2__abc_52155_new_n15495_; 
wire u2__abc_52155_new_n15496_; 
wire u2__abc_52155_new_n15497_; 
wire u2__abc_52155_new_n15498_; 
wire u2__abc_52155_new_n15499_; 
wire u2__abc_52155_new_n15500_; 
wire u2__abc_52155_new_n15501_; 
wire u2__abc_52155_new_n15502_; 
wire u2__abc_52155_new_n15503_; 
wire u2__abc_52155_new_n15504_; 
wire u2__abc_52155_new_n15505_; 
wire u2__abc_52155_new_n15506_; 
wire u2__abc_52155_new_n15507_; 
wire u2__abc_52155_new_n15508_; 
wire u2__abc_52155_new_n15509_; 
wire u2__abc_52155_new_n15510_; 
wire u2__abc_52155_new_n15511_; 
wire u2__abc_52155_new_n15512_; 
wire u2__abc_52155_new_n15513_; 
wire u2__abc_52155_new_n15514_; 
wire u2__abc_52155_new_n15515_; 
wire u2__abc_52155_new_n15516_; 
wire u2__abc_52155_new_n15517_; 
wire u2__abc_52155_new_n15519_; 
wire u2__abc_52155_new_n15520_; 
wire u2__abc_52155_new_n15521_; 
wire u2__abc_52155_new_n15522_; 
wire u2__abc_52155_new_n15523_; 
wire u2__abc_52155_new_n15524_; 
wire u2__abc_52155_new_n15525_; 
wire u2__abc_52155_new_n15526_; 
wire u2__abc_52155_new_n15527_; 
wire u2__abc_52155_new_n15528_; 
wire u2__abc_52155_new_n15529_; 
wire u2__abc_52155_new_n15530_; 
wire u2__abc_52155_new_n15531_; 
wire u2__abc_52155_new_n15532_; 
wire u2__abc_52155_new_n15533_; 
wire u2__abc_52155_new_n15534_; 
wire u2__abc_52155_new_n15536_; 
wire u2__abc_52155_new_n15537_; 
wire u2__abc_52155_new_n15538_; 
wire u2__abc_52155_new_n15539_; 
wire u2__abc_52155_new_n15540_; 
wire u2__abc_52155_new_n15541_; 
wire u2__abc_52155_new_n15542_; 
wire u2__abc_52155_new_n15543_; 
wire u2__abc_52155_new_n15544_; 
wire u2__abc_52155_new_n15545_; 
wire u2__abc_52155_new_n15546_; 
wire u2__abc_52155_new_n15547_; 
wire u2__abc_52155_new_n15548_; 
wire u2__abc_52155_new_n15549_; 
wire u2__abc_52155_new_n15550_; 
wire u2__abc_52155_new_n15551_; 
wire u2__abc_52155_new_n15552_; 
wire u2__abc_52155_new_n15553_; 
wire u2__abc_52155_new_n15554_; 
wire u2__abc_52155_new_n15556_; 
wire u2__abc_52155_new_n15557_; 
wire u2__abc_52155_new_n15558_; 
wire u2__abc_52155_new_n15559_; 
wire u2__abc_52155_new_n15560_; 
wire u2__abc_52155_new_n15561_; 
wire u2__abc_52155_new_n15562_; 
wire u2__abc_52155_new_n15563_; 
wire u2__abc_52155_new_n15564_; 
wire u2__abc_52155_new_n15565_; 
wire u2__abc_52155_new_n15566_; 
wire u2__abc_52155_new_n15567_; 
wire u2__abc_52155_new_n15568_; 
wire u2__abc_52155_new_n15569_; 
wire u2__abc_52155_new_n15570_; 
wire u2__abc_52155_new_n15571_; 
wire u2__abc_52155_new_n15573_; 
wire u2__abc_52155_new_n15574_; 
wire u2__abc_52155_new_n15575_; 
wire u2__abc_52155_new_n15576_; 
wire u2__abc_52155_new_n15577_; 
wire u2__abc_52155_new_n15578_; 
wire u2__abc_52155_new_n15579_; 
wire u2__abc_52155_new_n15580_; 
wire u2__abc_52155_new_n15581_; 
wire u2__abc_52155_new_n15582_; 
wire u2__abc_52155_new_n15583_; 
wire u2__abc_52155_new_n15584_; 
wire u2__abc_52155_new_n15585_; 
wire u2__abc_52155_new_n15586_; 
wire u2__abc_52155_new_n15587_; 
wire u2__abc_52155_new_n15588_; 
wire u2__abc_52155_new_n15589_; 
wire u2__abc_52155_new_n15590_; 
wire u2__abc_52155_new_n15591_; 
wire u2__abc_52155_new_n15592_; 
wire u2__abc_52155_new_n15594_; 
wire u2__abc_52155_new_n15595_; 
wire u2__abc_52155_new_n15596_; 
wire u2__abc_52155_new_n15597_; 
wire u2__abc_52155_new_n15598_; 
wire u2__abc_52155_new_n15599_; 
wire u2__abc_52155_new_n15600_; 
wire u2__abc_52155_new_n15601_; 
wire u2__abc_52155_new_n15602_; 
wire u2__abc_52155_new_n15603_; 
wire u2__abc_52155_new_n15604_; 
wire u2__abc_52155_new_n15605_; 
wire u2__abc_52155_new_n15606_; 
wire u2__abc_52155_new_n15607_; 
wire u2__abc_52155_new_n15608_; 
wire u2__abc_52155_new_n15609_; 
wire u2__abc_52155_new_n15611_; 
wire u2__abc_52155_new_n15612_; 
wire u2__abc_52155_new_n15613_; 
wire u2__abc_52155_new_n15614_; 
wire u2__abc_52155_new_n15615_; 
wire u2__abc_52155_new_n15616_; 
wire u2__abc_52155_new_n15617_; 
wire u2__abc_52155_new_n15618_; 
wire u2__abc_52155_new_n15619_; 
wire u2__abc_52155_new_n15620_; 
wire u2__abc_52155_new_n15621_; 
wire u2__abc_52155_new_n15622_; 
wire u2__abc_52155_new_n15623_; 
wire u2__abc_52155_new_n15624_; 
wire u2__abc_52155_new_n15625_; 
wire u2__abc_52155_new_n15626_; 
wire u2__abc_52155_new_n15627_; 
wire u2__abc_52155_new_n15628_; 
wire u2__abc_52155_new_n15630_; 
wire u2__abc_52155_new_n15631_; 
wire u2__abc_52155_new_n15632_; 
wire u2__abc_52155_new_n15633_; 
wire u2__abc_52155_new_n15634_; 
wire u2__abc_52155_new_n15635_; 
wire u2__abc_52155_new_n15636_; 
wire u2__abc_52155_new_n15637_; 
wire u2__abc_52155_new_n15638_; 
wire u2__abc_52155_new_n15639_; 
wire u2__abc_52155_new_n15640_; 
wire u2__abc_52155_new_n15641_; 
wire u2__abc_52155_new_n15642_; 
wire u2__abc_52155_new_n15643_; 
wire u2__abc_52155_new_n15644_; 
wire u2__abc_52155_new_n15645_; 
wire u2__abc_52155_new_n15647_; 
wire u2__abc_52155_new_n15648_; 
wire u2__abc_52155_new_n15649_; 
wire u2__abc_52155_new_n15650_; 
wire u2__abc_52155_new_n15651_; 
wire u2__abc_52155_new_n15652_; 
wire u2__abc_52155_new_n15653_; 
wire u2__abc_52155_new_n15654_; 
wire u2__abc_52155_new_n15655_; 
wire u2__abc_52155_new_n15656_; 
wire u2__abc_52155_new_n15657_; 
wire u2__abc_52155_new_n15658_; 
wire u2__abc_52155_new_n15659_; 
wire u2__abc_52155_new_n15660_; 
wire u2__abc_52155_new_n15661_; 
wire u2__abc_52155_new_n15662_; 
wire u2__abc_52155_new_n15663_; 
wire u2__abc_52155_new_n15664_; 
wire u2__abc_52155_new_n15665_; 
wire u2__abc_52155_new_n15666_; 
wire u2__abc_52155_new_n15667_; 
wire u2__abc_52155_new_n15668_; 
wire u2__abc_52155_new_n15669_; 
wire u2__abc_52155_new_n15670_; 
wire u2__abc_52155_new_n15672_; 
wire u2__abc_52155_new_n15673_; 
wire u2__abc_52155_new_n15674_; 
wire u2__abc_52155_new_n15675_; 
wire u2__abc_52155_new_n15676_; 
wire u2__abc_52155_new_n15677_; 
wire u2__abc_52155_new_n15678_; 
wire u2__abc_52155_new_n15679_; 
wire u2__abc_52155_new_n15680_; 
wire u2__abc_52155_new_n15681_; 
wire u2__abc_52155_new_n15682_; 
wire u2__abc_52155_new_n15683_; 
wire u2__abc_52155_new_n15684_; 
wire u2__abc_52155_new_n15685_; 
wire u2__abc_52155_new_n15686_; 
wire u2__abc_52155_new_n15687_; 
wire u2__abc_52155_new_n15689_; 
wire u2__abc_52155_new_n15690_; 
wire u2__abc_52155_new_n15691_; 
wire u2__abc_52155_new_n15692_; 
wire u2__abc_52155_new_n15693_; 
wire u2__abc_52155_new_n15694_; 
wire u2__abc_52155_new_n15695_; 
wire u2__abc_52155_new_n15696_; 
wire u2__abc_52155_new_n15697_; 
wire u2__abc_52155_new_n15698_; 
wire u2__abc_52155_new_n15699_; 
wire u2__abc_52155_new_n15700_; 
wire u2__abc_52155_new_n15701_; 
wire u2__abc_52155_new_n15702_; 
wire u2__abc_52155_new_n15703_; 
wire u2__abc_52155_new_n15704_; 
wire u2__abc_52155_new_n15705_; 
wire u2__abc_52155_new_n15706_; 
wire u2__abc_52155_new_n15708_; 
wire u2__abc_52155_new_n15709_; 
wire u2__abc_52155_new_n15710_; 
wire u2__abc_52155_new_n15711_; 
wire u2__abc_52155_new_n15712_; 
wire u2__abc_52155_new_n15713_; 
wire u2__abc_52155_new_n15714_; 
wire u2__abc_52155_new_n15715_; 
wire u2__abc_52155_new_n15716_; 
wire u2__abc_52155_new_n15717_; 
wire u2__abc_52155_new_n15718_; 
wire u2__abc_52155_new_n15719_; 
wire u2__abc_52155_new_n15720_; 
wire u2__abc_52155_new_n15721_; 
wire u2__abc_52155_new_n15722_; 
wire u2__abc_52155_new_n15723_; 
wire u2__abc_52155_new_n15725_; 
wire u2__abc_52155_new_n15726_; 
wire u2__abc_52155_new_n15727_; 
wire u2__abc_52155_new_n15728_; 
wire u2__abc_52155_new_n15729_; 
wire u2__abc_52155_new_n15730_; 
wire u2__abc_52155_new_n15731_; 
wire u2__abc_52155_new_n15732_; 
wire u2__abc_52155_new_n15733_; 
wire u2__abc_52155_new_n15734_; 
wire u2__abc_52155_new_n15735_; 
wire u2__abc_52155_new_n15736_; 
wire u2__abc_52155_new_n15737_; 
wire u2__abc_52155_new_n15738_; 
wire u2__abc_52155_new_n15739_; 
wire u2__abc_52155_new_n15740_; 
wire u2__abc_52155_new_n15741_; 
wire u2__abc_52155_new_n15742_; 
wire u2__abc_52155_new_n15743_; 
wire u2__abc_52155_new_n15744_; 
wire u2__abc_52155_new_n15745_; 
wire u2__abc_52155_new_n15746_; 
wire u2__abc_52155_new_n15748_; 
wire u2__abc_52155_new_n15749_; 
wire u2__abc_52155_new_n15750_; 
wire u2__abc_52155_new_n15751_; 
wire u2__abc_52155_new_n15752_; 
wire u2__abc_52155_new_n15753_; 
wire u2__abc_52155_new_n15754_; 
wire u2__abc_52155_new_n15755_; 
wire u2__abc_52155_new_n15756_; 
wire u2__abc_52155_new_n15757_; 
wire u2__abc_52155_new_n15758_; 
wire u2__abc_52155_new_n15759_; 
wire u2__abc_52155_new_n15760_; 
wire u2__abc_52155_new_n15761_; 
wire u2__abc_52155_new_n15762_; 
wire u2__abc_52155_new_n15763_; 
wire u2__abc_52155_new_n15765_; 
wire u2__abc_52155_new_n15766_; 
wire u2__abc_52155_new_n15767_; 
wire u2__abc_52155_new_n15768_; 
wire u2__abc_52155_new_n15769_; 
wire u2__abc_52155_new_n15770_; 
wire u2__abc_52155_new_n15771_; 
wire u2__abc_52155_new_n15772_; 
wire u2__abc_52155_new_n15773_; 
wire u2__abc_52155_new_n15774_; 
wire u2__abc_52155_new_n15775_; 
wire u2__abc_52155_new_n15776_; 
wire u2__abc_52155_new_n15777_; 
wire u2__abc_52155_new_n15778_; 
wire u2__abc_52155_new_n15779_; 
wire u2__abc_52155_new_n15780_; 
wire u2__abc_52155_new_n15781_; 
wire u2__abc_52155_new_n15782_; 
wire u2__abc_52155_new_n15784_; 
wire u2__abc_52155_new_n15785_; 
wire u2__abc_52155_new_n15786_; 
wire u2__abc_52155_new_n15787_; 
wire u2__abc_52155_new_n15788_; 
wire u2__abc_52155_new_n15789_; 
wire u2__abc_52155_new_n15790_; 
wire u2__abc_52155_new_n15791_; 
wire u2__abc_52155_new_n15792_; 
wire u2__abc_52155_new_n15793_; 
wire u2__abc_52155_new_n15794_; 
wire u2__abc_52155_new_n15795_; 
wire u2__abc_52155_new_n15796_; 
wire u2__abc_52155_new_n15797_; 
wire u2__abc_52155_new_n15798_; 
wire u2__abc_52155_new_n15799_; 
wire u2__abc_52155_new_n15801_; 
wire u2__abc_52155_new_n15802_; 
wire u2__abc_52155_new_n15803_; 
wire u2__abc_52155_new_n15804_; 
wire u2__abc_52155_new_n15805_; 
wire u2__abc_52155_new_n15806_; 
wire u2__abc_52155_new_n15807_; 
wire u2__abc_52155_new_n15808_; 
wire u2__abc_52155_new_n15809_; 
wire u2__abc_52155_new_n15810_; 
wire u2__abc_52155_new_n15811_; 
wire u2__abc_52155_new_n15812_; 
wire u2__abc_52155_new_n15813_; 
wire u2__abc_52155_new_n15814_; 
wire u2__abc_52155_new_n15815_; 
wire u2__abc_52155_new_n15816_; 
wire u2__abc_52155_new_n15817_; 
wire u2__abc_52155_new_n15818_; 
wire u2__abc_52155_new_n15819_; 
wire u2__abc_52155_new_n15820_; 
wire u2__abc_52155_new_n15821_; 
wire u2__abc_52155_new_n15822_; 
wire u2__abc_52155_new_n15823_; 
wire u2__abc_52155_new_n15824_; 
wire u2__abc_52155_new_n15825_; 
wire u2__abc_52155_new_n15826_; 
wire u2__abc_52155_new_n15827_; 
wire u2__abc_52155_new_n15828_; 
wire u2__abc_52155_new_n15829_; 
wire u2__abc_52155_new_n15830_; 
wire u2__abc_52155_new_n15832_; 
wire u2__abc_52155_new_n15833_; 
wire u2__abc_52155_new_n15834_; 
wire u2__abc_52155_new_n15835_; 
wire u2__abc_52155_new_n15836_; 
wire u2__abc_52155_new_n15837_; 
wire u2__abc_52155_new_n15838_; 
wire u2__abc_52155_new_n15839_; 
wire u2__abc_52155_new_n15840_; 
wire u2__abc_52155_new_n15841_; 
wire u2__abc_52155_new_n15842_; 
wire u2__abc_52155_new_n15843_; 
wire u2__abc_52155_new_n15844_; 
wire u2__abc_52155_new_n15845_; 
wire u2__abc_52155_new_n15846_; 
wire u2__abc_52155_new_n15847_; 
wire u2__abc_52155_new_n15849_; 
wire u2__abc_52155_new_n15850_; 
wire u2__abc_52155_new_n15851_; 
wire u2__abc_52155_new_n15852_; 
wire u2__abc_52155_new_n15853_; 
wire u2__abc_52155_new_n15854_; 
wire u2__abc_52155_new_n15855_; 
wire u2__abc_52155_new_n15856_; 
wire u2__abc_52155_new_n15857_; 
wire u2__abc_52155_new_n15858_; 
wire u2__abc_52155_new_n15859_; 
wire u2__abc_52155_new_n15860_; 
wire u2__abc_52155_new_n15861_; 
wire u2__abc_52155_new_n15862_; 
wire u2__abc_52155_new_n15863_; 
wire u2__abc_52155_new_n15864_; 
wire u2__abc_52155_new_n15865_; 
wire u2__abc_52155_new_n15866_; 
wire u2__abc_52155_new_n15868_; 
wire u2__abc_52155_new_n15869_; 
wire u2__abc_52155_new_n15870_; 
wire u2__abc_52155_new_n15871_; 
wire u2__abc_52155_new_n15872_; 
wire u2__abc_52155_new_n15873_; 
wire u2__abc_52155_new_n15874_; 
wire u2__abc_52155_new_n15875_; 
wire u2__abc_52155_new_n15876_; 
wire u2__abc_52155_new_n15877_; 
wire u2__abc_52155_new_n15878_; 
wire u2__abc_52155_new_n15879_; 
wire u2__abc_52155_new_n15880_; 
wire u2__abc_52155_new_n15881_; 
wire u2__abc_52155_new_n15882_; 
wire u2__abc_52155_new_n15883_; 
wire u2__abc_52155_new_n15885_; 
wire u2__abc_52155_new_n15886_; 
wire u2__abc_52155_new_n15887_; 
wire u2__abc_52155_new_n15888_; 
wire u2__abc_52155_new_n15889_; 
wire u2__abc_52155_new_n15890_; 
wire u2__abc_52155_new_n15891_; 
wire u2__abc_52155_new_n15892_; 
wire u2__abc_52155_new_n15893_; 
wire u2__abc_52155_new_n15894_; 
wire u2__abc_52155_new_n15895_; 
wire u2__abc_52155_new_n15896_; 
wire u2__abc_52155_new_n15897_; 
wire u2__abc_52155_new_n15898_; 
wire u2__abc_52155_new_n15899_; 
wire u2__abc_52155_new_n15900_; 
wire u2__abc_52155_new_n15901_; 
wire u2__abc_52155_new_n15902_; 
wire u2__abc_52155_new_n15903_; 
wire u2__abc_52155_new_n15904_; 
wire u2__abc_52155_new_n15905_; 
wire u2__abc_52155_new_n15906_; 
wire u2__abc_52155_new_n15908_; 
wire u2__abc_52155_new_n15909_; 
wire u2__abc_52155_new_n15910_; 
wire u2__abc_52155_new_n15911_; 
wire u2__abc_52155_new_n15912_; 
wire u2__abc_52155_new_n15913_; 
wire u2__abc_52155_new_n15914_; 
wire u2__abc_52155_new_n15915_; 
wire u2__abc_52155_new_n15916_; 
wire u2__abc_52155_new_n15917_; 
wire u2__abc_52155_new_n15918_; 
wire u2__abc_52155_new_n15919_; 
wire u2__abc_52155_new_n15920_; 
wire u2__abc_52155_new_n15921_; 
wire u2__abc_52155_new_n15922_; 
wire u2__abc_52155_new_n15923_; 
wire u2__abc_52155_new_n15925_; 
wire u2__abc_52155_new_n15926_; 
wire u2__abc_52155_new_n15927_; 
wire u2__abc_52155_new_n15928_; 
wire u2__abc_52155_new_n15929_; 
wire u2__abc_52155_new_n15930_; 
wire u2__abc_52155_new_n15931_; 
wire u2__abc_52155_new_n15932_; 
wire u2__abc_52155_new_n15933_; 
wire u2__abc_52155_new_n15934_; 
wire u2__abc_52155_new_n15935_; 
wire u2__abc_52155_new_n15936_; 
wire u2__abc_52155_new_n15937_; 
wire u2__abc_52155_new_n15938_; 
wire u2__abc_52155_new_n15939_; 
wire u2__abc_52155_new_n15940_; 
wire u2__abc_52155_new_n15941_; 
wire u2__abc_52155_new_n15942_; 
wire u2__abc_52155_new_n15944_; 
wire u2__abc_52155_new_n15945_; 
wire u2__abc_52155_new_n15946_; 
wire u2__abc_52155_new_n15947_; 
wire u2__abc_52155_new_n15948_; 
wire u2__abc_52155_new_n15949_; 
wire u2__abc_52155_new_n15950_; 
wire u2__abc_52155_new_n15951_; 
wire u2__abc_52155_new_n15952_; 
wire u2__abc_52155_new_n15953_; 
wire u2__abc_52155_new_n15954_; 
wire u2__abc_52155_new_n15955_; 
wire u2__abc_52155_new_n15956_; 
wire u2__abc_52155_new_n15957_; 
wire u2__abc_52155_new_n15958_; 
wire u2__abc_52155_new_n15959_; 
wire u2__abc_52155_new_n15961_; 
wire u2__abc_52155_new_n15962_; 
wire u2__abc_52155_new_n15963_; 
wire u2__abc_52155_new_n15964_; 
wire u2__abc_52155_new_n15965_; 
wire u2__abc_52155_new_n15966_; 
wire u2__abc_52155_new_n15967_; 
wire u2__abc_52155_new_n15968_; 
wire u2__abc_52155_new_n15969_; 
wire u2__abc_52155_new_n15970_; 
wire u2__abc_52155_new_n15971_; 
wire u2__abc_52155_new_n15972_; 
wire u2__abc_52155_new_n15973_; 
wire u2__abc_52155_new_n15974_; 
wire u2__abc_52155_new_n15975_; 
wire u2__abc_52155_new_n15976_; 
wire u2__abc_52155_new_n15977_; 
wire u2__abc_52155_new_n15978_; 
wire u2__abc_52155_new_n15979_; 
wire u2__abc_52155_new_n15980_; 
wire u2__abc_52155_new_n15981_; 
wire u2__abc_52155_new_n15982_; 
wire u2__abc_52155_new_n15983_; 
wire u2__abc_52155_new_n15984_; 
wire u2__abc_52155_new_n15986_; 
wire u2__abc_52155_new_n15987_; 
wire u2__abc_52155_new_n15988_; 
wire u2__abc_52155_new_n15989_; 
wire u2__abc_52155_new_n15990_; 
wire u2__abc_52155_new_n15991_; 
wire u2__abc_52155_new_n15992_; 
wire u2__abc_52155_new_n15993_; 
wire u2__abc_52155_new_n15994_; 
wire u2__abc_52155_new_n15995_; 
wire u2__abc_52155_new_n15996_; 
wire u2__abc_52155_new_n15997_; 
wire u2__abc_52155_new_n15998_; 
wire u2__abc_52155_new_n15999_; 
wire u2__abc_52155_new_n16000_; 
wire u2__abc_52155_new_n16001_; 
wire u2__abc_52155_new_n16003_; 
wire u2__abc_52155_new_n16004_; 
wire u2__abc_52155_new_n16005_; 
wire u2__abc_52155_new_n16006_; 
wire u2__abc_52155_new_n16007_; 
wire u2__abc_52155_new_n16008_; 
wire u2__abc_52155_new_n16009_; 
wire u2__abc_52155_new_n16010_; 
wire u2__abc_52155_new_n16011_; 
wire u2__abc_52155_new_n16012_; 
wire u2__abc_52155_new_n16013_; 
wire u2__abc_52155_new_n16014_; 
wire u2__abc_52155_new_n16015_; 
wire u2__abc_52155_new_n16016_; 
wire u2__abc_52155_new_n16017_; 
wire u2__abc_52155_new_n16018_; 
wire u2__abc_52155_new_n16020_; 
wire u2__abc_52155_new_n16021_; 
wire u2__abc_52155_new_n16022_; 
wire u2__abc_52155_new_n16023_; 
wire u2__abc_52155_new_n16024_; 
wire u2__abc_52155_new_n16025_; 
wire u2__abc_52155_new_n16026_; 
wire u2__abc_52155_new_n16027_; 
wire u2__abc_52155_new_n16028_; 
wire u2__abc_52155_new_n16029_; 
wire u2__abc_52155_new_n16030_; 
wire u2__abc_52155_new_n16031_; 
wire u2__abc_52155_new_n16032_; 
wire u2__abc_52155_new_n16033_; 
wire u2__abc_52155_new_n16034_; 
wire u2__abc_52155_new_n16035_; 
wire u2__abc_52155_new_n16037_; 
wire u2__abc_52155_new_n16038_; 
wire u2__abc_52155_new_n16039_; 
wire u2__abc_52155_new_n16040_; 
wire u2__abc_52155_new_n16041_; 
wire u2__abc_52155_new_n16042_; 
wire u2__abc_52155_new_n16043_; 
wire u2__abc_52155_new_n16044_; 
wire u2__abc_52155_new_n16045_; 
wire u2__abc_52155_new_n16046_; 
wire u2__abc_52155_new_n16047_; 
wire u2__abc_52155_new_n16048_; 
wire u2__abc_52155_new_n16049_; 
wire u2__abc_52155_new_n16050_; 
wire u2__abc_52155_new_n16051_; 
wire u2__abc_52155_new_n16052_; 
wire u2__abc_52155_new_n16053_; 
wire u2__abc_52155_new_n16054_; 
wire u2__abc_52155_new_n16055_; 
wire u2__abc_52155_new_n16056_; 
wire u2__abc_52155_new_n16057_; 
wire u2__abc_52155_new_n16058_; 
wire u2__abc_52155_new_n16059_; 
wire u2__abc_52155_new_n16061_; 
wire u2__abc_52155_new_n16062_; 
wire u2__abc_52155_new_n16063_; 
wire u2__abc_52155_new_n16064_; 
wire u2__abc_52155_new_n16065_; 
wire u2__abc_52155_new_n16066_; 
wire u2__abc_52155_new_n16067_; 
wire u2__abc_52155_new_n16068_; 
wire u2__abc_52155_new_n16069_; 
wire u2__abc_52155_new_n16070_; 
wire u2__abc_52155_new_n16071_; 
wire u2__abc_52155_new_n16072_; 
wire u2__abc_52155_new_n16073_; 
wire u2__abc_52155_new_n16074_; 
wire u2__abc_52155_new_n16075_; 
wire u2__abc_52155_new_n16076_; 
wire u2__abc_52155_new_n16078_; 
wire u2__abc_52155_new_n16079_; 
wire u2__abc_52155_new_n16080_; 
wire u2__abc_52155_new_n16081_; 
wire u2__abc_52155_new_n16082_; 
wire u2__abc_52155_new_n16083_; 
wire u2__abc_52155_new_n16084_; 
wire u2__abc_52155_new_n16085_; 
wire u2__abc_52155_new_n16086_; 
wire u2__abc_52155_new_n16087_; 
wire u2__abc_52155_new_n16088_; 
wire u2__abc_52155_new_n16089_; 
wire u2__abc_52155_new_n16090_; 
wire u2__abc_52155_new_n16091_; 
wire u2__abc_52155_new_n16092_; 
wire u2__abc_52155_new_n16093_; 
wire u2__abc_52155_new_n16094_; 
wire u2__abc_52155_new_n16095_; 
wire u2__abc_52155_new_n16097_; 
wire u2__abc_52155_new_n16098_; 
wire u2__abc_52155_new_n16099_; 
wire u2__abc_52155_new_n16100_; 
wire u2__abc_52155_new_n16101_; 
wire u2__abc_52155_new_n16102_; 
wire u2__abc_52155_new_n16103_; 
wire u2__abc_52155_new_n16104_; 
wire u2__abc_52155_new_n16105_; 
wire u2__abc_52155_new_n16106_; 
wire u2__abc_52155_new_n16107_; 
wire u2__abc_52155_new_n16108_; 
wire u2__abc_52155_new_n16109_; 
wire u2__abc_52155_new_n16110_; 
wire u2__abc_52155_new_n16111_; 
wire u2__abc_52155_new_n16112_; 
wire u2__abc_52155_new_n16114_; 
wire u2__abc_52155_new_n16115_; 
wire u2__abc_52155_new_n16116_; 
wire u2__abc_52155_new_n16117_; 
wire u2__abc_52155_new_n16118_; 
wire u2__abc_52155_new_n16119_; 
wire u2__abc_52155_new_n16120_; 
wire u2__abc_52155_new_n16121_; 
wire u2__abc_52155_new_n16122_; 
wire u2__abc_52155_new_n16123_; 
wire u2__abc_52155_new_n16124_; 
wire u2__abc_52155_new_n16125_; 
wire u2__abc_52155_new_n16126_; 
wire u2__abc_52155_new_n16127_; 
wire u2__abc_52155_new_n16128_; 
wire u2__abc_52155_new_n16129_; 
wire u2__abc_52155_new_n16130_; 
wire u2__abc_52155_new_n16131_; 
wire u2__abc_52155_new_n16132_; 
wire u2__abc_52155_new_n16133_; 
wire u2__abc_52155_new_n16134_; 
wire u2__abc_52155_new_n16135_; 
wire u2__abc_52155_new_n16136_; 
wire u2__abc_52155_new_n16137_; 
wire u2__abc_52155_new_n16138_; 
wire u2__abc_52155_new_n16139_; 
wire u2__abc_52155_new_n16141_; 
wire u2__abc_52155_new_n16142_; 
wire u2__abc_52155_new_n16143_; 
wire u2__abc_52155_new_n16144_; 
wire u2__abc_52155_new_n16145_; 
wire u2__abc_52155_new_n16146_; 
wire u2__abc_52155_new_n16147_; 
wire u2__abc_52155_new_n16148_; 
wire u2__abc_52155_new_n16149_; 
wire u2__abc_52155_new_n16150_; 
wire u2__abc_52155_new_n16151_; 
wire u2__abc_52155_new_n16152_; 
wire u2__abc_52155_new_n16153_; 
wire u2__abc_52155_new_n16154_; 
wire u2__abc_52155_new_n16155_; 
wire u2__abc_52155_new_n16156_; 
wire u2__abc_52155_new_n16158_; 
wire u2__abc_52155_new_n16159_; 
wire u2__abc_52155_new_n16160_; 
wire u2__abc_52155_new_n16161_; 
wire u2__abc_52155_new_n16162_; 
wire u2__abc_52155_new_n16163_; 
wire u2__abc_52155_new_n16164_; 
wire u2__abc_52155_new_n16165_; 
wire u2__abc_52155_new_n16166_; 
wire u2__abc_52155_new_n16167_; 
wire u2__abc_52155_new_n16168_; 
wire u2__abc_52155_new_n16169_; 
wire u2__abc_52155_new_n16170_; 
wire u2__abc_52155_new_n16171_; 
wire u2__abc_52155_new_n16172_; 
wire u2__abc_52155_new_n16173_; 
wire u2__abc_52155_new_n16174_; 
wire u2__abc_52155_new_n16175_; 
wire u2__abc_52155_new_n16176_; 
wire u2__abc_52155_new_n16178_; 
wire u2__abc_52155_new_n16179_; 
wire u2__abc_52155_new_n16180_; 
wire u2__abc_52155_new_n16181_; 
wire u2__abc_52155_new_n16182_; 
wire u2__abc_52155_new_n16183_; 
wire u2__abc_52155_new_n16184_; 
wire u2__abc_52155_new_n16185_; 
wire u2__abc_52155_new_n16186_; 
wire u2__abc_52155_new_n16187_; 
wire u2__abc_52155_new_n16188_; 
wire u2__abc_52155_new_n16189_; 
wire u2__abc_52155_new_n16190_; 
wire u2__abc_52155_new_n16191_; 
wire u2__abc_52155_new_n16192_; 
wire u2__abc_52155_new_n16193_; 
wire u2__abc_52155_new_n16195_; 
wire u2__abc_52155_new_n16196_; 
wire u2__abc_52155_new_n16197_; 
wire u2__abc_52155_new_n16198_; 
wire u2__abc_52155_new_n16199_; 
wire u2__abc_52155_new_n16200_; 
wire u2__abc_52155_new_n16201_; 
wire u2__abc_52155_new_n16202_; 
wire u2__abc_52155_new_n16203_; 
wire u2__abc_52155_new_n16204_; 
wire u2__abc_52155_new_n16205_; 
wire u2__abc_52155_new_n16206_; 
wire u2__abc_52155_new_n16207_; 
wire u2__abc_52155_new_n16208_; 
wire u2__abc_52155_new_n16209_; 
wire u2__abc_52155_new_n16210_; 
wire u2__abc_52155_new_n16211_; 
wire u2__abc_52155_new_n16212_; 
wire u2__abc_52155_new_n16214_; 
wire u2__abc_52155_new_n16215_; 
wire u2__abc_52155_new_n16216_; 
wire u2__abc_52155_new_n16217_; 
wire u2__abc_52155_new_n16218_; 
wire u2__abc_52155_new_n16219_; 
wire u2__abc_52155_new_n16220_; 
wire u2__abc_52155_new_n16221_; 
wire u2__abc_52155_new_n16222_; 
wire u2__abc_52155_new_n16223_; 
wire u2__abc_52155_new_n16224_; 
wire u2__abc_52155_new_n16225_; 
wire u2__abc_52155_new_n16226_; 
wire u2__abc_52155_new_n16227_; 
wire u2__abc_52155_new_n16228_; 
wire u2__abc_52155_new_n16229_; 
wire u2__abc_52155_new_n16231_; 
wire u2__abc_52155_new_n16232_; 
wire u2__abc_52155_new_n16233_; 
wire u2__abc_52155_new_n16234_; 
wire u2__abc_52155_new_n16235_; 
wire u2__abc_52155_new_n16236_; 
wire u2__abc_52155_new_n16237_; 
wire u2__abc_52155_new_n16238_; 
wire u2__abc_52155_new_n16239_; 
wire u2__abc_52155_new_n16240_; 
wire u2__abc_52155_new_n16241_; 
wire u2__abc_52155_new_n16242_; 
wire u2__abc_52155_new_n16243_; 
wire u2__abc_52155_new_n16244_; 
wire u2__abc_52155_new_n16245_; 
wire u2__abc_52155_new_n16246_; 
wire u2__abc_52155_new_n16248_; 
wire u2__abc_52155_new_n16249_; 
wire u2__abc_52155_new_n16250_; 
wire u2__abc_52155_new_n16251_; 
wire u2__abc_52155_new_n16252_; 
wire u2__abc_52155_new_n16253_; 
wire u2__abc_52155_new_n16254_; 
wire u2__abc_52155_new_n16255_; 
wire u2__abc_52155_new_n16256_; 
wire u2__abc_52155_new_n16257_; 
wire u2__abc_52155_new_n16258_; 
wire u2__abc_52155_new_n16259_; 
wire u2__abc_52155_new_n16260_; 
wire u2__abc_52155_new_n16261_; 
wire u2__abc_52155_new_n16262_; 
wire u2__abc_52155_new_n16263_; 
wire u2__abc_52155_new_n16265_; 
wire u2__abc_52155_new_n16266_; 
wire u2__abc_52155_new_n16267_; 
wire u2__abc_52155_new_n16268_; 
wire u2__abc_52155_new_n16269_; 
wire u2__abc_52155_new_n16270_; 
wire u2__abc_52155_new_n16271_; 
wire u2__abc_52155_new_n16272_; 
wire u2__abc_52155_new_n16273_; 
wire u2__abc_52155_new_n16274_; 
wire u2__abc_52155_new_n16275_; 
wire u2__abc_52155_new_n16276_; 
wire u2__abc_52155_new_n16277_; 
wire u2__abc_52155_new_n16278_; 
wire u2__abc_52155_new_n16279_; 
wire u2__abc_52155_new_n16280_; 
wire u2__abc_52155_new_n16281_; 
wire u2__abc_52155_new_n16282_; 
wire u2__abc_52155_new_n16283_; 
wire u2__abc_52155_new_n16284_; 
wire u2__abc_52155_new_n16285_; 
wire u2__abc_52155_new_n16286_; 
wire u2__abc_52155_new_n16287_; 
wire u2__abc_52155_new_n16288_; 
wire u2__abc_52155_new_n16289_; 
wire u2__abc_52155_new_n16290_; 
wire u2__abc_52155_new_n16291_; 
wire u2__abc_52155_new_n16292_; 
wire u2__abc_52155_new_n16293_; 
wire u2__abc_52155_new_n16294_; 
wire u2__abc_52155_new_n16296_; 
wire u2__abc_52155_new_n16297_; 
wire u2__abc_52155_new_n16298_; 
wire u2__abc_52155_new_n16299_; 
wire u2__abc_52155_new_n16300_; 
wire u2__abc_52155_new_n16301_; 
wire u2__abc_52155_new_n16302_; 
wire u2__abc_52155_new_n16303_; 
wire u2__abc_52155_new_n16304_; 
wire u2__abc_52155_new_n16305_; 
wire u2__abc_52155_new_n16306_; 
wire u2__abc_52155_new_n16307_; 
wire u2__abc_52155_new_n16308_; 
wire u2__abc_52155_new_n16309_; 
wire u2__abc_52155_new_n16310_; 
wire u2__abc_52155_new_n16311_; 
wire u2__abc_52155_new_n16313_; 
wire u2__abc_52155_new_n16314_; 
wire u2__abc_52155_new_n16315_; 
wire u2__abc_52155_new_n16316_; 
wire u2__abc_52155_new_n16317_; 
wire u2__abc_52155_new_n16318_; 
wire u2__abc_52155_new_n16319_; 
wire u2__abc_52155_new_n16320_; 
wire u2__abc_52155_new_n16321_; 
wire u2__abc_52155_new_n16322_; 
wire u2__abc_52155_new_n16323_; 
wire u2__abc_52155_new_n16324_; 
wire u2__abc_52155_new_n16325_; 
wire u2__abc_52155_new_n16326_; 
wire u2__abc_52155_new_n16327_; 
wire u2__abc_52155_new_n16328_; 
wire u2__abc_52155_new_n16329_; 
wire u2__abc_52155_new_n16330_; 
wire u2__abc_52155_new_n16331_; 
wire u2__abc_52155_new_n16333_; 
wire u2__abc_52155_new_n16334_; 
wire u2__abc_52155_new_n16335_; 
wire u2__abc_52155_new_n16336_; 
wire u2__abc_52155_new_n16337_; 
wire u2__abc_52155_new_n16338_; 
wire u2__abc_52155_new_n16339_; 
wire u2__abc_52155_new_n16340_; 
wire u2__abc_52155_new_n16341_; 
wire u2__abc_52155_new_n16342_; 
wire u2__abc_52155_new_n16343_; 
wire u2__abc_52155_new_n16344_; 
wire u2__abc_52155_new_n16345_; 
wire u2__abc_52155_new_n16346_; 
wire u2__abc_52155_new_n16347_; 
wire u2__abc_52155_new_n16348_; 
wire u2__abc_52155_new_n16350_; 
wire u2__abc_52155_new_n16351_; 
wire u2__abc_52155_new_n16352_; 
wire u2__abc_52155_new_n16353_; 
wire u2__abc_52155_new_n16354_; 
wire u2__abc_52155_new_n16355_; 
wire u2__abc_52155_new_n16356_; 
wire u2__abc_52155_new_n16357_; 
wire u2__abc_52155_new_n16358_; 
wire u2__abc_52155_new_n16359_; 
wire u2__abc_52155_new_n16360_; 
wire u2__abc_52155_new_n16361_; 
wire u2__abc_52155_new_n16362_; 
wire u2__abc_52155_new_n16363_; 
wire u2__abc_52155_new_n16364_; 
wire u2__abc_52155_new_n16365_; 
wire u2__abc_52155_new_n16366_; 
wire u2__abc_52155_new_n16367_; 
wire u2__abc_52155_new_n16368_; 
wire u2__abc_52155_new_n16369_; 
wire u2__abc_52155_new_n16371_; 
wire u2__abc_52155_new_n16372_; 
wire u2__abc_52155_new_n16373_; 
wire u2__abc_52155_new_n16374_; 
wire u2__abc_52155_new_n16375_; 
wire u2__abc_52155_new_n16376_; 
wire u2__abc_52155_new_n16377_; 
wire u2__abc_52155_new_n16378_; 
wire u2__abc_52155_new_n16379_; 
wire u2__abc_52155_new_n16380_; 
wire u2__abc_52155_new_n16381_; 
wire u2__abc_52155_new_n16382_; 
wire u2__abc_52155_new_n16383_; 
wire u2__abc_52155_new_n16384_; 
wire u2__abc_52155_new_n16385_; 
wire u2__abc_52155_new_n16386_; 
wire u2__abc_52155_new_n16388_; 
wire u2__abc_52155_new_n16389_; 
wire u2__abc_52155_new_n16390_; 
wire u2__abc_52155_new_n16391_; 
wire u2__abc_52155_new_n16392_; 
wire u2__abc_52155_new_n16393_; 
wire u2__abc_52155_new_n16394_; 
wire u2__abc_52155_new_n16395_; 
wire u2__abc_52155_new_n16396_; 
wire u2__abc_52155_new_n16397_; 
wire u2__abc_52155_new_n16398_; 
wire u2__abc_52155_new_n16399_; 
wire u2__abc_52155_new_n16400_; 
wire u2__abc_52155_new_n16401_; 
wire u2__abc_52155_new_n16402_; 
wire u2__abc_52155_new_n16403_; 
wire u2__abc_52155_new_n16404_; 
wire u2__abc_52155_new_n16405_; 
wire u2__abc_52155_new_n16407_; 
wire u2__abc_52155_new_n16408_; 
wire u2__abc_52155_new_n16409_; 
wire u2__abc_52155_new_n16410_; 
wire u2__abc_52155_new_n16411_; 
wire u2__abc_52155_new_n16412_; 
wire u2__abc_52155_new_n16413_; 
wire u2__abc_52155_new_n16414_; 
wire u2__abc_52155_new_n16415_; 
wire u2__abc_52155_new_n16416_; 
wire u2__abc_52155_new_n16417_; 
wire u2__abc_52155_new_n16418_; 
wire u2__abc_52155_new_n16419_; 
wire u2__abc_52155_new_n16420_; 
wire u2__abc_52155_new_n16421_; 
wire u2__abc_52155_new_n16422_; 
wire u2__abc_52155_new_n16424_; 
wire u2__abc_52155_new_n16425_; 
wire u2__abc_52155_new_n16426_; 
wire u2__abc_52155_new_n16427_; 
wire u2__abc_52155_new_n16428_; 
wire u2__abc_52155_new_n16429_; 
wire u2__abc_52155_new_n16430_; 
wire u2__abc_52155_new_n16431_; 
wire u2__abc_52155_new_n16432_; 
wire u2__abc_52155_new_n16433_; 
wire u2__abc_52155_new_n16434_; 
wire u2__abc_52155_new_n16435_; 
wire u2__abc_52155_new_n16436_; 
wire u2__abc_52155_new_n16437_; 
wire u2__abc_52155_new_n16438_; 
wire u2__abc_52155_new_n16439_; 
wire u2__abc_52155_new_n16440_; 
wire u2__abc_52155_new_n16441_; 
wire u2__abc_52155_new_n16442_; 
wire u2__abc_52155_new_n16443_; 
wire u2__abc_52155_new_n16444_; 
wire u2__abc_52155_new_n16445_; 
wire u2__abc_52155_new_n16446_; 
wire u2__abc_52155_new_n16447_; 
wire u2__abc_52155_new_n16448_; 
wire u2__abc_52155_new_n16449_; 
wire u2__abc_52155_new_n16450_; 
wire u2__abc_52155_new_n16451_; 
wire u2__abc_52155_new_n16453_; 
wire u2__abc_52155_new_n16454_; 
wire u2__abc_52155_new_n16455_; 
wire u2__abc_52155_new_n16456_; 
wire u2__abc_52155_new_n16457_; 
wire u2__abc_52155_new_n16458_; 
wire u2__abc_52155_new_n16459_; 
wire u2__abc_52155_new_n16460_; 
wire u2__abc_52155_new_n16461_; 
wire u2__abc_52155_new_n16462_; 
wire u2__abc_52155_new_n16463_; 
wire u2__abc_52155_new_n16464_; 
wire u2__abc_52155_new_n16465_; 
wire u2__abc_52155_new_n16466_; 
wire u2__abc_52155_new_n16467_; 
wire u2__abc_52155_new_n16468_; 
wire u2__abc_52155_new_n16470_; 
wire u2__abc_52155_new_n16471_; 
wire u2__abc_52155_new_n16472_; 
wire u2__abc_52155_new_n16473_; 
wire u2__abc_52155_new_n16474_; 
wire u2__abc_52155_new_n16475_; 
wire u2__abc_52155_new_n16477_; 
wire u2__abc_52155_new_n16478_; 
wire u2__abc_52155_new_n16479_; 
wire u2__abc_52155_new_n16480_; 
wire u2__abc_52155_new_n16481_; 
wire u2__abc_52155_new_n16483_; 
wire u2__abc_52155_new_n16484_; 
wire u2__abc_52155_new_n16485_; 
wire u2__abc_52155_new_n16486_; 
wire u2__abc_52155_new_n16487_; 
wire u2__abc_52155_new_n16488_; 
wire u2__abc_52155_new_n16489_; 
wire u2__abc_52155_new_n16490_; 
wire u2__abc_52155_new_n16492_; 
wire u2__abc_52155_new_n16493_; 
wire u2__abc_52155_new_n16494_; 
wire u2__abc_52155_new_n16495_; 
wire u2__abc_52155_new_n16496_; 
wire u2__abc_52155_new_n16497_; 
wire u2__abc_52155_new_n16498_; 
wire u2__abc_52155_new_n16500_; 
wire u2__abc_52155_new_n16501_; 
wire u2__abc_52155_new_n16502_; 
wire u2__abc_52155_new_n16503_; 
wire u2__abc_52155_new_n16505_; 
wire u2__abc_52155_new_n16506_; 
wire u2__abc_52155_new_n16507_; 
wire u2__abc_52155_new_n16508_; 
wire u2__abc_52155_new_n16510_; 
wire u2__abc_52155_new_n16511_; 
wire u2__abc_52155_new_n16512_; 
wire u2__abc_52155_new_n16513_; 
wire u2__abc_52155_new_n16514_; 
wire u2__abc_52155_new_n16516_; 
wire u2__abc_52155_new_n16517_; 
wire u2__abc_52155_new_n16518_; 
wire u2__abc_52155_new_n16519_; 
wire u2__abc_52155_new_n16520_; 
wire u2__abc_52155_new_n16522_; 
wire u2__abc_52155_new_n16523_; 
wire u2__abc_52155_new_n16525_; 
wire u2__abc_52155_new_n16527_; 
wire u2__abc_52155_new_n16528_; 
wire u2__abc_52155_new_n16529_; 
wire u2__abc_52155_new_n16530_; 
wire u2__abc_52155_new_n16532_; 
wire u2__abc_52155_new_n16533_; 
wire u2__abc_52155_new_n16534_; 
wire u2__abc_52155_new_n16535_; 
wire u2__abc_52155_new_n16537_; 
wire u2__abc_52155_new_n16538_; 
wire u2__abc_52155_new_n16539_; 
wire u2__abc_52155_new_n16540_; 
wire u2__abc_52155_new_n16542_; 
wire u2__abc_52155_new_n16543_; 
wire u2__abc_52155_new_n16544_; 
wire u2__abc_52155_new_n16545_; 
wire u2__abc_52155_new_n16547_; 
wire u2__abc_52155_new_n16548_; 
wire u2__abc_52155_new_n16549_; 
wire u2__abc_52155_new_n16550_; 
wire u2__abc_52155_new_n16552_; 
wire u2__abc_52155_new_n16553_; 
wire u2__abc_52155_new_n16554_; 
wire u2__abc_52155_new_n16555_; 
wire u2__abc_52155_new_n16557_; 
wire u2__abc_52155_new_n16558_; 
wire u2__abc_52155_new_n16559_; 
wire u2__abc_52155_new_n16560_; 
wire u2__abc_52155_new_n16562_; 
wire u2__abc_52155_new_n16563_; 
wire u2__abc_52155_new_n16564_; 
wire u2__abc_52155_new_n16565_; 
wire u2__abc_52155_new_n16567_; 
wire u2__abc_52155_new_n16568_; 
wire u2__abc_52155_new_n16569_; 
wire u2__abc_52155_new_n16570_; 
wire u2__abc_52155_new_n16572_; 
wire u2__abc_52155_new_n16573_; 
wire u2__abc_52155_new_n16574_; 
wire u2__abc_52155_new_n16575_; 
wire u2__abc_52155_new_n16577_; 
wire u2__abc_52155_new_n16578_; 
wire u2__abc_52155_new_n16579_; 
wire u2__abc_52155_new_n16580_; 
wire u2__abc_52155_new_n16582_; 
wire u2__abc_52155_new_n16583_; 
wire u2__abc_52155_new_n16584_; 
wire u2__abc_52155_new_n16585_; 
wire u2__abc_52155_new_n16587_; 
wire u2__abc_52155_new_n16588_; 
wire u2__abc_52155_new_n16589_; 
wire u2__abc_52155_new_n16590_; 
wire u2__abc_52155_new_n16592_; 
wire u2__abc_52155_new_n16593_; 
wire u2__abc_52155_new_n16594_; 
wire u2__abc_52155_new_n16595_; 
wire u2__abc_52155_new_n16597_; 
wire u2__abc_52155_new_n16598_; 
wire u2__abc_52155_new_n16599_; 
wire u2__abc_52155_new_n16600_; 
wire u2__abc_52155_new_n16602_; 
wire u2__abc_52155_new_n16603_; 
wire u2__abc_52155_new_n16604_; 
wire u2__abc_52155_new_n16605_; 
wire u2__abc_52155_new_n16607_; 
wire u2__abc_52155_new_n16608_; 
wire u2__abc_52155_new_n16609_; 
wire u2__abc_52155_new_n16610_; 
wire u2__abc_52155_new_n16612_; 
wire u2__abc_52155_new_n16613_; 
wire u2__abc_52155_new_n16614_; 
wire u2__abc_52155_new_n16615_; 
wire u2__abc_52155_new_n16617_; 
wire u2__abc_52155_new_n16618_; 
wire u2__abc_52155_new_n16619_; 
wire u2__abc_52155_new_n16620_; 
wire u2__abc_52155_new_n16622_; 
wire u2__abc_52155_new_n16623_; 
wire u2__abc_52155_new_n16624_; 
wire u2__abc_52155_new_n16625_; 
wire u2__abc_52155_new_n16627_; 
wire u2__abc_52155_new_n16628_; 
wire u2__abc_52155_new_n16629_; 
wire u2__abc_52155_new_n16630_; 
wire u2__abc_52155_new_n16632_; 
wire u2__abc_52155_new_n16633_; 
wire u2__abc_52155_new_n16634_; 
wire u2__abc_52155_new_n16635_; 
wire u2__abc_52155_new_n16637_; 
wire u2__abc_52155_new_n16638_; 
wire u2__abc_52155_new_n16639_; 
wire u2__abc_52155_new_n16640_; 
wire u2__abc_52155_new_n16642_; 
wire u2__abc_52155_new_n16643_; 
wire u2__abc_52155_new_n16644_; 
wire u2__abc_52155_new_n16645_; 
wire u2__abc_52155_new_n16647_; 
wire u2__abc_52155_new_n16648_; 
wire u2__abc_52155_new_n16649_; 
wire u2__abc_52155_new_n16650_; 
wire u2__abc_52155_new_n16652_; 
wire u2__abc_52155_new_n16653_; 
wire u2__abc_52155_new_n16654_; 
wire u2__abc_52155_new_n16655_; 
wire u2__abc_52155_new_n16657_; 
wire u2__abc_52155_new_n16658_; 
wire u2__abc_52155_new_n16659_; 
wire u2__abc_52155_new_n16660_; 
wire u2__abc_52155_new_n16662_; 
wire u2__abc_52155_new_n16663_; 
wire u2__abc_52155_new_n16664_; 
wire u2__abc_52155_new_n16665_; 
wire u2__abc_52155_new_n16667_; 
wire u2__abc_52155_new_n16668_; 
wire u2__abc_52155_new_n16669_; 
wire u2__abc_52155_new_n16670_; 
wire u2__abc_52155_new_n16672_; 
wire u2__abc_52155_new_n16673_; 
wire u2__abc_52155_new_n16674_; 
wire u2__abc_52155_new_n16675_; 
wire u2__abc_52155_new_n16677_; 
wire u2__abc_52155_new_n16678_; 
wire u2__abc_52155_new_n16679_; 
wire u2__abc_52155_new_n16680_; 
wire u2__abc_52155_new_n16681_; 
wire u2__abc_52155_new_n16682_; 
wire u2__abc_52155_new_n16683_; 
wire u2__abc_52155_new_n16684_; 
wire u2__abc_52155_new_n16685_; 
wire u2__abc_52155_new_n16686_; 
wire u2__abc_52155_new_n16688_; 
wire u2__abc_52155_new_n16689_; 
wire u2__abc_52155_new_n16690_; 
wire u2__abc_52155_new_n16691_; 
wire u2__abc_52155_new_n16692_; 
wire u2__abc_52155_new_n16694_; 
wire u2__abc_52155_new_n16695_; 
wire u2__abc_52155_new_n16696_; 
wire u2__abc_52155_new_n16697_; 
wire u2__abc_52155_new_n16698_; 
wire u2__abc_52155_new_n16699_; 
wire u2__abc_52155_new_n16700_; 
wire u2__abc_52155_new_n16701_; 
wire u2__abc_52155_new_n16703_; 
wire u2__abc_52155_new_n16704_; 
wire u2__abc_52155_new_n16705_; 
wire u2__abc_52155_new_n16706_; 
wire u2__abc_52155_new_n16707_; 
wire u2__abc_52155_new_n16709_; 
wire u2__abc_52155_new_n16710_; 
wire u2__abc_52155_new_n16711_; 
wire u2__abc_52155_new_n16712_; 
wire u2__abc_52155_new_n16713_; 
wire u2__abc_52155_new_n16715_; 
wire u2__abc_52155_new_n16716_; 
wire u2__abc_52155_new_n16717_; 
wire u2__abc_52155_new_n16718_; 
wire u2__abc_52155_new_n16719_; 
wire u2__abc_52155_new_n16721_; 
wire u2__abc_52155_new_n16722_; 
wire u2__abc_52155_new_n16723_; 
wire u2__abc_52155_new_n16724_; 
wire u2__abc_52155_new_n16725_; 
wire u2__abc_52155_new_n16727_; 
wire u2__abc_52155_new_n16728_; 
wire u2__abc_52155_new_n16729_; 
wire u2__abc_52155_new_n16730_; 
wire u2__abc_52155_new_n16731_; 
wire u2__abc_52155_new_n16733_; 
wire u2__abc_52155_new_n16734_; 
wire u2__abc_52155_new_n16735_; 
wire u2__abc_52155_new_n16736_; 
wire u2__abc_52155_new_n16737_; 
wire u2__abc_52155_new_n16739_; 
wire u2__abc_52155_new_n16740_; 
wire u2__abc_52155_new_n16741_; 
wire u2__abc_52155_new_n16742_; 
wire u2__abc_52155_new_n16743_; 
wire u2__abc_52155_new_n16745_; 
wire u2__abc_52155_new_n16746_; 
wire u2__abc_52155_new_n16747_; 
wire u2__abc_52155_new_n16748_; 
wire u2__abc_52155_new_n16749_; 
wire u2__abc_52155_new_n16751_; 
wire u2__abc_52155_new_n16752_; 
wire u2__abc_52155_new_n16753_; 
wire u2__abc_52155_new_n16754_; 
wire u2__abc_52155_new_n16755_; 
wire u2__abc_52155_new_n16757_; 
wire u2__abc_52155_new_n16758_; 
wire u2__abc_52155_new_n16759_; 
wire u2__abc_52155_new_n16760_; 
wire u2__abc_52155_new_n16761_; 
wire u2__abc_52155_new_n16763_; 
wire u2__abc_52155_new_n16764_; 
wire u2__abc_52155_new_n16765_; 
wire u2__abc_52155_new_n16766_; 
wire u2__abc_52155_new_n16767_; 
wire u2__abc_52155_new_n16769_; 
wire u2__abc_52155_new_n16770_; 
wire u2__abc_52155_new_n16771_; 
wire u2__abc_52155_new_n16772_; 
wire u2__abc_52155_new_n16773_; 
wire u2__abc_52155_new_n16774_; 
wire u2__abc_52155_new_n16775_; 
wire u2__abc_52155_new_n16776_; 
wire u2__abc_52155_new_n16778_; 
wire u2__abc_52155_new_n16779_; 
wire u2__abc_52155_new_n16780_; 
wire u2__abc_52155_new_n16781_; 
wire u2__abc_52155_new_n16782_; 
wire u2__abc_52155_new_n16784_; 
wire u2__abc_52155_new_n16785_; 
wire u2__abc_52155_new_n16786_; 
wire u2__abc_52155_new_n16787_; 
wire u2__abc_52155_new_n16788_; 
wire u2__abc_52155_new_n16790_; 
wire u2__abc_52155_new_n16791_; 
wire u2__abc_52155_new_n16792_; 
wire u2__abc_52155_new_n16793_; 
wire u2__abc_52155_new_n16794_; 
wire u2__abc_52155_new_n16796_; 
wire u2__abc_52155_new_n16797_; 
wire u2__abc_52155_new_n16798_; 
wire u2__abc_52155_new_n16799_; 
wire u2__abc_52155_new_n16800_; 
wire u2__abc_52155_new_n16802_; 
wire u2__abc_52155_new_n16803_; 
wire u2__abc_52155_new_n16804_; 
wire u2__abc_52155_new_n16805_; 
wire u2__abc_52155_new_n16806_; 
wire u2__abc_52155_new_n16808_; 
wire u2__abc_52155_new_n16809_; 
wire u2__abc_52155_new_n16810_; 
wire u2__abc_52155_new_n16811_; 
wire u2__abc_52155_new_n16812_; 
wire u2__abc_52155_new_n16814_; 
wire u2__abc_52155_new_n16815_; 
wire u2__abc_52155_new_n16816_; 
wire u2__abc_52155_new_n16817_; 
wire u2__abc_52155_new_n16818_; 
wire u2__abc_52155_new_n16820_; 
wire u2__abc_52155_new_n16821_; 
wire u2__abc_52155_new_n16822_; 
wire u2__abc_52155_new_n16823_; 
wire u2__abc_52155_new_n16824_; 
wire u2__abc_52155_new_n16826_; 
wire u2__abc_52155_new_n16827_; 
wire u2__abc_52155_new_n16828_; 
wire u2__abc_52155_new_n16829_; 
wire u2__abc_52155_new_n16830_; 
wire u2__abc_52155_new_n16832_; 
wire u2__abc_52155_new_n16833_; 
wire u2__abc_52155_new_n16834_; 
wire u2__abc_52155_new_n16835_; 
wire u2__abc_52155_new_n16836_; 
wire u2__abc_52155_new_n16838_; 
wire u2__abc_52155_new_n16839_; 
wire u2__abc_52155_new_n16840_; 
wire u2__abc_52155_new_n16841_; 
wire u2__abc_52155_new_n16842_; 
wire u2__abc_52155_new_n16844_; 
wire u2__abc_52155_new_n16845_; 
wire u2__abc_52155_new_n16846_; 
wire u2__abc_52155_new_n16847_; 
wire u2__abc_52155_new_n16848_; 
wire u2__abc_52155_new_n16850_; 
wire u2__abc_52155_new_n16851_; 
wire u2__abc_52155_new_n16852_; 
wire u2__abc_52155_new_n16853_; 
wire u2__abc_52155_new_n16854_; 
wire u2__abc_52155_new_n16856_; 
wire u2__abc_52155_new_n16857_; 
wire u2__abc_52155_new_n16858_; 
wire u2__abc_52155_new_n16859_; 
wire u2__abc_52155_new_n16860_; 
wire u2__abc_52155_new_n16862_; 
wire u2__abc_52155_new_n16863_; 
wire u2__abc_52155_new_n16864_; 
wire u2__abc_52155_new_n16865_; 
wire u2__abc_52155_new_n16866_; 
wire u2__abc_52155_new_n16867_; 
wire u2__abc_52155_new_n16868_; 
wire u2__abc_52155_new_n16869_; 
wire u2__abc_52155_new_n16871_; 
wire u2__abc_52155_new_n16872_; 
wire u2__abc_52155_new_n16873_; 
wire u2__abc_52155_new_n16874_; 
wire u2__abc_52155_new_n16875_; 
wire u2__abc_52155_new_n16877_; 
wire u2__abc_52155_new_n16878_; 
wire u2__abc_52155_new_n16879_; 
wire u2__abc_52155_new_n16880_; 
wire u2__abc_52155_new_n16881_; 
wire u2__abc_52155_new_n16883_; 
wire u2__abc_52155_new_n16884_; 
wire u2__abc_52155_new_n16885_; 
wire u2__abc_52155_new_n16886_; 
wire u2__abc_52155_new_n16887_; 
wire u2__abc_52155_new_n16889_; 
wire u2__abc_52155_new_n16890_; 
wire u2__abc_52155_new_n16891_; 
wire u2__abc_52155_new_n16892_; 
wire u2__abc_52155_new_n16893_; 
wire u2__abc_52155_new_n16894_; 
wire u2__abc_52155_new_n16895_; 
wire u2__abc_52155_new_n16896_; 
wire u2__abc_52155_new_n16898_; 
wire u2__abc_52155_new_n16899_; 
wire u2__abc_52155_new_n16900_; 
wire u2__abc_52155_new_n16901_; 
wire u2__abc_52155_new_n16902_; 
wire u2__abc_52155_new_n16904_; 
wire u2__abc_52155_new_n16905_; 
wire u2__abc_52155_new_n16906_; 
wire u2__abc_52155_new_n16907_; 
wire u2__abc_52155_new_n16908_; 
wire u2__abc_52155_new_n16910_; 
wire u2__abc_52155_new_n16911_; 
wire u2__abc_52155_new_n16912_; 
wire u2__abc_52155_new_n16913_; 
wire u2__abc_52155_new_n16914_; 
wire u2__abc_52155_new_n16916_; 
wire u2__abc_52155_new_n16917_; 
wire u2__abc_52155_new_n16918_; 
wire u2__abc_52155_new_n16919_; 
wire u2__abc_52155_new_n16920_; 
wire u2__abc_52155_new_n16922_; 
wire u2__abc_52155_new_n16923_; 
wire u2__abc_52155_new_n16924_; 
wire u2__abc_52155_new_n16925_; 
wire u2__abc_52155_new_n16926_; 
wire u2__abc_52155_new_n16928_; 
wire u2__abc_52155_new_n16929_; 
wire u2__abc_52155_new_n16930_; 
wire u2__abc_52155_new_n16931_; 
wire u2__abc_52155_new_n16932_; 
wire u2__abc_52155_new_n16934_; 
wire u2__abc_52155_new_n16935_; 
wire u2__abc_52155_new_n16936_; 
wire u2__abc_52155_new_n16937_; 
wire u2__abc_52155_new_n16938_; 
wire u2__abc_52155_new_n16940_; 
wire u2__abc_52155_new_n16941_; 
wire u2__abc_52155_new_n16942_; 
wire u2__abc_52155_new_n16943_; 
wire u2__abc_52155_new_n16944_; 
wire u2__abc_52155_new_n16946_; 
wire u2__abc_52155_new_n16947_; 
wire u2__abc_52155_new_n16948_; 
wire u2__abc_52155_new_n16949_; 
wire u2__abc_52155_new_n16950_; 
wire u2__abc_52155_new_n16951_; 
wire u2__abc_52155_new_n16952_; 
wire u2__abc_52155_new_n16953_; 
wire u2__abc_52155_new_n16955_; 
wire u2__abc_52155_new_n16956_; 
wire u2__abc_52155_new_n16957_; 
wire u2__abc_52155_new_n16958_; 
wire u2__abc_52155_new_n16959_; 
wire u2__abc_52155_new_n16961_; 
wire u2__abc_52155_new_n16962_; 
wire u2__abc_52155_new_n16963_; 
wire u2__abc_52155_new_n16964_; 
wire u2__abc_52155_new_n16965_; 
wire u2__abc_52155_new_n16967_; 
wire u2__abc_52155_new_n16968_; 
wire u2__abc_52155_new_n16969_; 
wire u2__abc_52155_new_n16970_; 
wire u2__abc_52155_new_n16971_; 
wire u2__abc_52155_new_n16973_; 
wire u2__abc_52155_new_n16974_; 
wire u2__abc_52155_new_n16975_; 
wire u2__abc_52155_new_n16976_; 
wire u2__abc_52155_new_n16977_; 
wire u2__abc_52155_new_n16979_; 
wire u2__abc_52155_new_n16980_; 
wire u2__abc_52155_new_n16981_; 
wire u2__abc_52155_new_n16982_; 
wire u2__abc_52155_new_n16983_; 
wire u2__abc_52155_new_n16985_; 
wire u2__abc_52155_new_n16986_; 
wire u2__abc_52155_new_n16987_; 
wire u2__abc_52155_new_n16988_; 
wire u2__abc_52155_new_n16989_; 
wire u2__abc_52155_new_n16990_; 
wire u2__abc_52155_new_n16991_; 
wire u2__abc_52155_new_n16992_; 
wire u2__abc_52155_new_n16994_; 
wire u2__abc_52155_new_n16995_; 
wire u2__abc_52155_new_n16996_; 
wire u2__abc_52155_new_n16997_; 
wire u2__abc_52155_new_n16998_; 
wire u2__abc_52155_new_n17000_; 
wire u2__abc_52155_new_n17001_; 
wire u2__abc_52155_new_n17002_; 
wire u2__abc_52155_new_n17003_; 
wire u2__abc_52155_new_n17004_; 
wire u2__abc_52155_new_n17006_; 
wire u2__abc_52155_new_n17007_; 
wire u2__abc_52155_new_n17008_; 
wire u2__abc_52155_new_n17009_; 
wire u2__abc_52155_new_n17010_; 
wire u2__abc_52155_new_n17012_; 
wire u2__abc_52155_new_n17013_; 
wire u2__abc_52155_new_n17014_; 
wire u2__abc_52155_new_n17015_; 
wire u2__abc_52155_new_n17016_; 
wire u2__abc_52155_new_n17018_; 
wire u2__abc_52155_new_n17019_; 
wire u2__abc_52155_new_n17020_; 
wire u2__abc_52155_new_n17021_; 
wire u2__abc_52155_new_n17022_; 
wire u2__abc_52155_new_n17024_; 
wire u2__abc_52155_new_n17025_; 
wire u2__abc_52155_new_n17026_; 
wire u2__abc_52155_new_n17027_; 
wire u2__abc_52155_new_n17028_; 
wire u2__abc_52155_new_n17030_; 
wire u2__abc_52155_new_n17031_; 
wire u2__abc_52155_new_n17032_; 
wire u2__abc_52155_new_n17033_; 
wire u2__abc_52155_new_n17034_; 
wire u2__abc_52155_new_n17036_; 
wire u2__abc_52155_new_n17037_; 
wire u2__abc_52155_new_n17038_; 
wire u2__abc_52155_new_n17039_; 
wire u2__abc_52155_new_n17040_; 
wire u2__abc_52155_new_n17042_; 
wire u2__abc_52155_new_n17043_; 
wire u2__abc_52155_new_n17044_; 
wire u2__abc_52155_new_n17045_; 
wire u2__abc_52155_new_n17046_; 
wire u2__abc_52155_new_n17048_; 
wire u2__abc_52155_new_n17049_; 
wire u2__abc_52155_new_n17050_; 
wire u2__abc_52155_new_n17051_; 
wire u2__abc_52155_new_n17052_; 
wire u2__abc_52155_new_n17054_; 
wire u2__abc_52155_new_n17055_; 
wire u2__abc_52155_new_n17056_; 
wire u2__abc_52155_new_n17057_; 
wire u2__abc_52155_new_n17058_; 
wire u2__abc_52155_new_n17060_; 
wire u2__abc_52155_new_n17061_; 
wire u2__abc_52155_new_n17062_; 
wire u2__abc_52155_new_n17063_; 
wire u2__abc_52155_new_n17064_; 
wire u2__abc_52155_new_n17066_; 
wire u2__abc_52155_new_n17067_; 
wire u2__abc_52155_new_n17068_; 
wire u2__abc_52155_new_n17069_; 
wire u2__abc_52155_new_n17070_; 
wire u2__abc_52155_new_n17072_; 
wire u2__abc_52155_new_n17073_; 
wire u2__abc_52155_new_n17074_; 
wire u2__abc_52155_new_n17075_; 
wire u2__abc_52155_new_n17076_; 
wire u2__abc_52155_new_n17078_; 
wire u2__abc_52155_new_n17079_; 
wire u2__abc_52155_new_n17080_; 
wire u2__abc_52155_new_n17081_; 
wire u2__abc_52155_new_n17082_; 
wire u2__abc_52155_new_n17084_; 
wire u2__abc_52155_new_n17085_; 
wire u2__abc_52155_new_n17086_; 
wire u2__abc_52155_new_n17087_; 
wire u2__abc_52155_new_n17088_; 
wire u2__abc_52155_new_n17089_; 
wire u2__abc_52155_new_n17091_; 
wire u2__abc_52155_new_n17092_; 
wire u2__abc_52155_new_n17093_; 
wire u2__abc_52155_new_n17094_; 
wire u2__abc_52155_new_n17095_; 
wire u2__abc_52155_new_n17096_; 
wire u2__abc_52155_new_n17097_; 
wire u2__abc_52155_new_n17098_; 
wire u2__abc_52155_new_n17100_; 
wire u2__abc_52155_new_n17101_; 
wire u2__abc_52155_new_n17102_; 
wire u2__abc_52155_new_n17103_; 
wire u2__abc_52155_new_n17104_; 
wire u2__abc_52155_new_n17106_; 
wire u2__abc_52155_new_n17107_; 
wire u2__abc_52155_new_n17108_; 
wire u2__abc_52155_new_n17109_; 
wire u2__abc_52155_new_n17110_; 
wire u2__abc_52155_new_n17112_; 
wire u2__abc_52155_new_n17113_; 
wire u2__abc_52155_new_n17114_; 
wire u2__abc_52155_new_n17115_; 
wire u2__abc_52155_new_n17116_; 
wire u2__abc_52155_new_n17118_; 
wire u2__abc_52155_new_n17119_; 
wire u2__abc_52155_new_n17120_; 
wire u2__abc_52155_new_n17121_; 
wire u2__abc_52155_new_n17122_; 
wire u2__abc_52155_new_n17124_; 
wire u2__abc_52155_new_n17125_; 
wire u2__abc_52155_new_n17126_; 
wire u2__abc_52155_new_n17127_; 
wire u2__abc_52155_new_n17128_; 
wire u2__abc_52155_new_n17130_; 
wire u2__abc_52155_new_n17131_; 
wire u2__abc_52155_new_n17132_; 
wire u2__abc_52155_new_n17133_; 
wire u2__abc_52155_new_n17134_; 
wire u2__abc_52155_new_n17136_; 
wire u2__abc_52155_new_n17137_; 
wire u2__abc_52155_new_n17138_; 
wire u2__abc_52155_new_n17139_; 
wire u2__abc_52155_new_n17140_; 
wire u2__abc_52155_new_n17142_; 
wire u2__abc_52155_new_n17143_; 
wire u2__abc_52155_new_n17144_; 
wire u2__abc_52155_new_n17145_; 
wire u2__abc_52155_new_n17146_; 
wire u2__abc_52155_new_n17148_; 
wire u2__abc_52155_new_n17149_; 
wire u2__abc_52155_new_n17150_; 
wire u2__abc_52155_new_n17151_; 
wire u2__abc_52155_new_n17152_; 
wire u2__abc_52155_new_n17154_; 
wire u2__abc_52155_new_n17155_; 
wire u2__abc_52155_new_n17156_; 
wire u2__abc_52155_new_n17157_; 
wire u2__abc_52155_new_n17158_; 
wire u2__abc_52155_new_n17160_; 
wire u2__abc_52155_new_n17161_; 
wire u2__abc_52155_new_n17162_; 
wire u2__abc_52155_new_n17163_; 
wire u2__abc_52155_new_n17164_; 
wire u2__abc_52155_new_n17166_; 
wire u2__abc_52155_new_n17167_; 
wire u2__abc_52155_new_n17168_; 
wire u2__abc_52155_new_n17169_; 
wire u2__abc_52155_new_n17170_; 
wire u2__abc_52155_new_n17172_; 
wire u2__abc_52155_new_n17173_; 
wire u2__abc_52155_new_n17174_; 
wire u2__abc_52155_new_n17175_; 
wire u2__abc_52155_new_n17176_; 
wire u2__abc_52155_new_n17177_; 
wire u2__abc_52155_new_n17178_; 
wire u2__abc_52155_new_n17179_; 
wire u2__abc_52155_new_n17181_; 
wire u2__abc_52155_new_n17182_; 
wire u2__abc_52155_new_n17183_; 
wire u2__abc_52155_new_n17184_; 
wire u2__abc_52155_new_n17185_; 
wire u2__abc_52155_new_n17187_; 
wire u2__abc_52155_new_n17188_; 
wire u2__abc_52155_new_n17189_; 
wire u2__abc_52155_new_n17190_; 
wire u2__abc_52155_new_n17191_; 
wire u2__abc_52155_new_n17193_; 
wire u2__abc_52155_new_n17194_; 
wire u2__abc_52155_new_n17195_; 
wire u2__abc_52155_new_n17196_; 
wire u2__abc_52155_new_n17197_; 
wire u2__abc_52155_new_n17199_; 
wire u2__abc_52155_new_n17200_; 
wire u2__abc_52155_new_n17201_; 
wire u2__abc_52155_new_n17202_; 
wire u2__abc_52155_new_n17203_; 
wire u2__abc_52155_new_n17204_; 
wire u2__abc_52155_new_n17205_; 
wire u2__abc_52155_new_n17206_; 
wire u2__abc_52155_new_n17208_; 
wire u2__abc_52155_new_n17209_; 
wire u2__abc_52155_new_n17210_; 
wire u2__abc_52155_new_n17211_; 
wire u2__abc_52155_new_n17212_; 
wire u2__abc_52155_new_n17214_; 
wire u2__abc_52155_new_n17215_; 
wire u2__abc_52155_new_n17216_; 
wire u2__abc_52155_new_n17217_; 
wire u2__abc_52155_new_n17218_; 
wire u2__abc_52155_new_n17220_; 
wire u2__abc_52155_new_n17221_; 
wire u2__abc_52155_new_n17222_; 
wire u2__abc_52155_new_n17223_; 
wire u2__abc_52155_new_n17224_; 
wire u2__abc_52155_new_n17226_; 
wire u2__abc_52155_new_n17227_; 
wire u2__abc_52155_new_n17228_; 
wire u2__abc_52155_new_n17229_; 
wire u2__abc_52155_new_n17230_; 
wire u2__abc_52155_new_n17232_; 
wire u2__abc_52155_new_n17233_; 
wire u2__abc_52155_new_n17234_; 
wire u2__abc_52155_new_n17235_; 
wire u2__abc_52155_new_n17236_; 
wire u2__abc_52155_new_n17238_; 
wire u2__abc_52155_new_n17239_; 
wire u2__abc_52155_new_n17240_; 
wire u2__abc_52155_new_n17241_; 
wire u2__abc_52155_new_n17242_; 
wire u2__abc_52155_new_n17244_; 
wire u2__abc_52155_new_n17245_; 
wire u2__abc_52155_new_n17246_; 
wire u2__abc_52155_new_n17247_; 
wire u2__abc_52155_new_n17248_; 
wire u2__abc_52155_new_n17250_; 
wire u2__abc_52155_new_n17251_; 
wire u2__abc_52155_new_n17252_; 
wire u2__abc_52155_new_n17253_; 
wire u2__abc_52155_new_n17254_; 
wire u2__abc_52155_new_n17256_; 
wire u2__abc_52155_new_n17257_; 
wire u2__abc_52155_new_n17258_; 
wire u2__abc_52155_new_n17259_; 
wire u2__abc_52155_new_n17260_; 
wire u2__abc_52155_new_n17262_; 
wire u2__abc_52155_new_n17263_; 
wire u2__abc_52155_new_n17264_; 
wire u2__abc_52155_new_n17265_; 
wire u2__abc_52155_new_n17266_; 
wire u2__abc_52155_new_n17268_; 
wire u2__abc_52155_new_n17269_; 
wire u2__abc_52155_new_n17270_; 
wire u2__abc_52155_new_n17271_; 
wire u2__abc_52155_new_n17272_; 
wire u2__abc_52155_new_n17274_; 
wire u2__abc_52155_new_n17275_; 
wire u2__abc_52155_new_n17276_; 
wire u2__abc_52155_new_n17277_; 
wire u2__abc_52155_new_n17278_; 
wire u2__abc_52155_new_n17280_; 
wire u2__abc_52155_new_n17281_; 
wire u2__abc_52155_new_n17282_; 
wire u2__abc_52155_new_n17283_; 
wire u2__abc_52155_new_n17284_; 
wire u2__abc_52155_new_n17286_; 
wire u2__abc_52155_new_n17287_; 
wire u2__abc_52155_new_n17288_; 
wire u2__abc_52155_new_n17289_; 
wire u2__abc_52155_new_n17290_; 
wire u2__abc_52155_new_n17292_; 
wire u2__abc_52155_new_n17293_; 
wire u2__abc_52155_new_n17294_; 
wire u2__abc_52155_new_n17295_; 
wire u2__abc_52155_new_n17296_; 
wire u2__abc_52155_new_n17297_; 
wire u2__abc_52155_new_n17298_; 
wire u2__abc_52155_new_n17299_; 
wire u2__abc_52155_new_n17301_; 
wire u2__abc_52155_new_n17302_; 
wire u2__abc_52155_new_n17303_; 
wire u2__abc_52155_new_n17304_; 
wire u2__abc_52155_new_n17305_; 
wire u2__abc_52155_new_n17307_; 
wire u2__abc_52155_new_n17308_; 
wire u2__abc_52155_new_n17309_; 
wire u2__abc_52155_new_n17310_; 
wire u2__abc_52155_new_n17311_; 
wire u2__abc_52155_new_n17313_; 
wire u2__abc_52155_new_n17314_; 
wire u2__abc_52155_new_n17315_; 
wire u2__abc_52155_new_n17316_; 
wire u2__abc_52155_new_n17317_; 
wire u2__abc_52155_new_n17319_; 
wire u2__abc_52155_new_n17320_; 
wire u2__abc_52155_new_n17321_; 
wire u2__abc_52155_new_n17322_; 
wire u2__abc_52155_new_n17323_; 
wire u2__abc_52155_new_n17325_; 
wire u2__abc_52155_new_n17326_; 
wire u2__abc_52155_new_n17327_; 
wire u2__abc_52155_new_n17328_; 
wire u2__abc_52155_new_n17329_; 
wire u2__abc_52155_new_n17331_; 
wire u2__abc_52155_new_n17332_; 
wire u2__abc_52155_new_n17333_; 
wire u2__abc_52155_new_n17334_; 
wire u2__abc_52155_new_n17335_; 
wire u2__abc_52155_new_n17337_; 
wire u2__abc_52155_new_n17338_; 
wire u2__abc_52155_new_n17339_; 
wire u2__abc_52155_new_n17340_; 
wire u2__abc_52155_new_n17341_; 
wire u2__abc_52155_new_n17343_; 
wire u2__abc_52155_new_n17344_; 
wire u2__abc_52155_new_n17345_; 
wire u2__abc_52155_new_n17346_; 
wire u2__abc_52155_new_n17347_; 
wire u2__abc_52155_new_n17349_; 
wire u2__abc_52155_new_n17350_; 
wire u2__abc_52155_new_n17351_; 
wire u2__abc_52155_new_n17352_; 
wire u2__abc_52155_new_n17353_; 
wire u2__abc_52155_new_n17355_; 
wire u2__abc_52155_new_n17356_; 
wire u2__abc_52155_new_n17357_; 
wire u2__abc_52155_new_n17358_; 
wire u2__abc_52155_new_n17359_; 
wire u2__abc_52155_new_n17361_; 
wire u2__abc_52155_new_n17362_; 
wire u2__abc_52155_new_n17363_; 
wire u2__abc_52155_new_n17364_; 
wire u2__abc_52155_new_n17365_; 
wire u2__abc_52155_new_n17367_; 
wire u2__abc_52155_new_n17368_; 
wire u2__abc_52155_new_n17369_; 
wire u2__abc_52155_new_n17370_; 
wire u2__abc_52155_new_n17371_; 
wire u2__abc_52155_new_n17373_; 
wire u2__abc_52155_new_n17374_; 
wire u2__abc_52155_new_n17375_; 
wire u2__abc_52155_new_n17376_; 
wire u2__abc_52155_new_n17377_; 
wire u2__abc_52155_new_n17378_; 
wire u2__abc_52155_new_n17379_; 
wire u2__abc_52155_new_n17380_; 
wire u2__abc_52155_new_n17382_; 
wire u2__abc_52155_new_n17383_; 
wire u2__abc_52155_new_n17384_; 
wire u2__abc_52155_new_n17385_; 
wire u2__abc_52155_new_n17386_; 
wire u2__abc_52155_new_n17388_; 
wire u2__abc_52155_new_n17389_; 
wire u2__abc_52155_new_n17390_; 
wire u2__abc_52155_new_n17391_; 
wire u2__abc_52155_new_n17392_; 
wire u2__abc_52155_new_n17394_; 
wire u2__abc_52155_new_n17395_; 
wire u2__abc_52155_new_n17396_; 
wire u2__abc_52155_new_n17397_; 
wire u2__abc_52155_new_n17398_; 
wire u2__abc_52155_new_n17400_; 
wire u2__abc_52155_new_n17401_; 
wire u2__abc_52155_new_n17402_; 
wire u2__abc_52155_new_n17403_; 
wire u2__abc_52155_new_n17404_; 
wire u2__abc_52155_new_n17406_; 
wire u2__abc_52155_new_n17407_; 
wire u2__abc_52155_new_n17408_; 
wire u2__abc_52155_new_n17409_; 
wire u2__abc_52155_new_n17410_; 
wire u2__abc_52155_new_n17412_; 
wire u2__abc_52155_new_n17413_; 
wire u2__abc_52155_new_n17414_; 
wire u2__abc_52155_new_n17415_; 
wire u2__abc_52155_new_n17416_; 
wire u2__abc_52155_new_n17418_; 
wire u2__abc_52155_new_n17419_; 
wire u2__abc_52155_new_n17420_; 
wire u2__abc_52155_new_n17421_; 
wire u2__abc_52155_new_n17422_; 
wire u2__abc_52155_new_n17424_; 
wire u2__abc_52155_new_n17425_; 
wire u2__abc_52155_new_n17426_; 
wire u2__abc_52155_new_n17427_; 
wire u2__abc_52155_new_n17428_; 
wire u2__abc_52155_new_n17430_; 
wire u2__abc_52155_new_n17431_; 
wire u2__abc_52155_new_n17432_; 
wire u2__abc_52155_new_n17433_; 
wire u2__abc_52155_new_n17434_; 
wire u2__abc_52155_new_n17436_; 
wire u2__abc_52155_new_n17437_; 
wire u2__abc_52155_new_n17438_; 
wire u2__abc_52155_new_n17439_; 
wire u2__abc_52155_new_n17440_; 
wire u2__abc_52155_new_n17442_; 
wire u2__abc_52155_new_n17443_; 
wire u2__abc_52155_new_n17444_; 
wire u2__abc_52155_new_n17445_; 
wire u2__abc_52155_new_n17446_; 
wire u2__abc_52155_new_n17448_; 
wire u2__abc_52155_new_n17449_; 
wire u2__abc_52155_new_n17450_; 
wire u2__abc_52155_new_n17451_; 
wire u2__abc_52155_new_n17452_; 
wire u2__abc_52155_new_n17454_; 
wire u2__abc_52155_new_n17455_; 
wire u2__abc_52155_new_n17456_; 
wire u2__abc_52155_new_n17457_; 
wire u2__abc_52155_new_n17458_; 
wire u2__abc_52155_new_n17460_; 
wire u2__abc_52155_new_n17461_; 
wire u2__abc_52155_new_n17462_; 
wire u2__abc_52155_new_n17463_; 
wire u2__abc_52155_new_n17464_; 
wire u2__abc_52155_new_n17466_; 
wire u2__abc_52155_new_n17467_; 
wire u2__abc_52155_new_n17468_; 
wire u2__abc_52155_new_n17469_; 
wire u2__abc_52155_new_n17470_; 
wire u2__abc_52155_new_n17472_; 
wire u2__abc_52155_new_n17473_; 
wire u2__abc_52155_new_n17474_; 
wire u2__abc_52155_new_n17475_; 
wire u2__abc_52155_new_n17476_; 
wire u2__abc_52155_new_n17478_; 
wire u2__abc_52155_new_n17479_; 
wire u2__abc_52155_new_n17480_; 
wire u2__abc_52155_new_n17481_; 
wire u2__abc_52155_new_n17482_; 
wire u2__abc_52155_new_n17484_; 
wire u2__abc_52155_new_n17485_; 
wire u2__abc_52155_new_n17486_; 
wire u2__abc_52155_new_n17487_; 
wire u2__abc_52155_new_n17488_; 
wire u2__abc_52155_new_n17489_; 
wire u2__abc_52155_new_n17490_; 
wire u2__abc_52155_new_n17491_; 
wire u2__abc_52155_new_n17493_; 
wire u2__abc_52155_new_n17494_; 
wire u2__abc_52155_new_n17495_; 
wire u2__abc_52155_new_n17496_; 
wire u2__abc_52155_new_n17497_; 
wire u2__abc_52155_new_n17498_; 
wire u2__abc_52155_new_n17499_; 
wire u2__abc_52155_new_n17500_; 
wire u2__abc_52155_new_n17502_; 
wire u2__abc_52155_new_n17503_; 
wire u2__abc_52155_new_n17504_; 
wire u2__abc_52155_new_n17505_; 
wire u2__abc_52155_new_n17506_; 
wire u2__abc_52155_new_n17508_; 
wire u2__abc_52155_new_n17509_; 
wire u2__abc_52155_new_n17510_; 
wire u2__abc_52155_new_n17511_; 
wire u2__abc_52155_new_n17512_; 
wire u2__abc_52155_new_n17514_; 
wire u2__abc_52155_new_n17515_; 
wire u2__abc_52155_new_n17516_; 
wire u2__abc_52155_new_n17517_; 
wire u2__abc_52155_new_n17518_; 
wire u2__abc_52155_new_n17520_; 
wire u2__abc_52155_new_n17521_; 
wire u2__abc_52155_new_n17522_; 
wire u2__abc_52155_new_n17523_; 
wire u2__abc_52155_new_n17524_; 
wire u2__abc_52155_new_n17526_; 
wire u2__abc_52155_new_n17527_; 
wire u2__abc_52155_new_n17528_; 
wire u2__abc_52155_new_n17529_; 
wire u2__abc_52155_new_n17530_; 
wire u2__abc_52155_new_n17532_; 
wire u2__abc_52155_new_n17533_; 
wire u2__abc_52155_new_n17534_; 
wire u2__abc_52155_new_n17535_; 
wire u2__abc_52155_new_n17536_; 
wire u2__abc_52155_new_n17538_; 
wire u2__abc_52155_new_n17539_; 
wire u2__abc_52155_new_n17540_; 
wire u2__abc_52155_new_n17541_; 
wire u2__abc_52155_new_n17542_; 
wire u2__abc_52155_new_n17544_; 
wire u2__abc_52155_new_n17545_; 
wire u2__abc_52155_new_n17546_; 
wire u2__abc_52155_new_n17547_; 
wire u2__abc_52155_new_n17548_; 
wire u2__abc_52155_new_n17550_; 
wire u2__abc_52155_new_n17551_; 
wire u2__abc_52155_new_n17552_; 
wire u2__abc_52155_new_n17553_; 
wire u2__abc_52155_new_n17554_; 
wire u2__abc_52155_new_n17556_; 
wire u2__abc_52155_new_n17557_; 
wire u2__abc_52155_new_n17558_; 
wire u2__abc_52155_new_n17559_; 
wire u2__abc_52155_new_n17560_; 
wire u2__abc_52155_new_n17562_; 
wire u2__abc_52155_new_n17563_; 
wire u2__abc_52155_new_n17564_; 
wire u2__abc_52155_new_n17565_; 
wire u2__abc_52155_new_n17566_; 
wire u2__abc_52155_new_n17568_; 
wire u2__abc_52155_new_n17569_; 
wire u2__abc_52155_new_n17570_; 
wire u2__abc_52155_new_n17571_; 
wire u2__abc_52155_new_n17572_; 
wire u2__abc_52155_new_n17574_; 
wire u2__abc_52155_new_n17575_; 
wire u2__abc_52155_new_n17576_; 
wire u2__abc_52155_new_n17577_; 
wire u2__abc_52155_new_n17578_; 
wire u2__abc_52155_new_n17580_; 
wire u2__abc_52155_new_n17581_; 
wire u2__abc_52155_new_n17582_; 
wire u2__abc_52155_new_n17583_; 
wire u2__abc_52155_new_n17584_; 
wire u2__abc_52155_new_n17586_; 
wire u2__abc_52155_new_n17587_; 
wire u2__abc_52155_new_n17588_; 
wire u2__abc_52155_new_n17589_; 
wire u2__abc_52155_new_n17590_; 
wire u2__abc_52155_new_n17592_; 
wire u2__abc_52155_new_n17593_; 
wire u2__abc_52155_new_n17594_; 
wire u2__abc_52155_new_n17595_; 
wire u2__abc_52155_new_n17596_; 
wire u2__abc_52155_new_n17598_; 
wire u2__abc_52155_new_n17599_; 
wire u2__abc_52155_new_n17600_; 
wire u2__abc_52155_new_n17601_; 
wire u2__abc_52155_new_n17602_; 
wire u2__abc_52155_new_n17604_; 
wire u2__abc_52155_new_n17605_; 
wire u2__abc_52155_new_n17606_; 
wire u2__abc_52155_new_n17607_; 
wire u2__abc_52155_new_n17608_; 
wire u2__abc_52155_new_n17610_; 
wire u2__abc_52155_new_n17611_; 
wire u2__abc_52155_new_n17612_; 
wire u2__abc_52155_new_n17613_; 
wire u2__abc_52155_new_n17614_; 
wire u2__abc_52155_new_n17616_; 
wire u2__abc_52155_new_n17617_; 
wire u2__abc_52155_new_n17618_; 
wire u2__abc_52155_new_n17619_; 
wire u2__abc_52155_new_n17620_; 
wire u2__abc_52155_new_n17622_; 
wire u2__abc_52155_new_n17623_; 
wire u2__abc_52155_new_n17624_; 
wire u2__abc_52155_new_n17625_; 
wire u2__abc_52155_new_n17626_; 
wire u2__abc_52155_new_n17628_; 
wire u2__abc_52155_new_n17629_; 
wire u2__abc_52155_new_n17630_; 
wire u2__abc_52155_new_n17631_; 
wire u2__abc_52155_new_n17632_; 
wire u2__abc_52155_new_n17634_; 
wire u2__abc_52155_new_n17635_; 
wire u2__abc_52155_new_n17636_; 
wire u2__abc_52155_new_n17637_; 
wire u2__abc_52155_new_n17638_; 
wire u2__abc_52155_new_n17640_; 
wire u2__abc_52155_new_n17641_; 
wire u2__abc_52155_new_n17642_; 
wire u2__abc_52155_new_n17643_; 
wire u2__abc_52155_new_n17644_; 
wire u2__abc_52155_new_n17646_; 
wire u2__abc_52155_new_n17647_; 
wire u2__abc_52155_new_n17648_; 
wire u2__abc_52155_new_n17649_; 
wire u2__abc_52155_new_n17650_; 
wire u2__abc_52155_new_n17652_; 
wire u2__abc_52155_new_n17653_; 
wire u2__abc_52155_new_n17654_; 
wire u2__abc_52155_new_n17655_; 
wire u2__abc_52155_new_n17656_; 
wire u2__abc_52155_new_n17658_; 
wire u2__abc_52155_new_n17659_; 
wire u2__abc_52155_new_n17660_; 
wire u2__abc_52155_new_n17661_; 
wire u2__abc_52155_new_n17662_; 
wire u2__abc_52155_new_n17664_; 
wire u2__abc_52155_new_n17665_; 
wire u2__abc_52155_new_n17666_; 
wire u2__abc_52155_new_n17667_; 
wire u2__abc_52155_new_n17668_; 
wire u2__abc_52155_new_n17670_; 
wire u2__abc_52155_new_n17671_; 
wire u2__abc_52155_new_n17672_; 
wire u2__abc_52155_new_n17673_; 
wire u2__abc_52155_new_n17674_; 
wire u2__abc_52155_new_n17676_; 
wire u2__abc_52155_new_n17677_; 
wire u2__abc_52155_new_n17678_; 
wire u2__abc_52155_new_n17679_; 
wire u2__abc_52155_new_n17680_; 
wire u2__abc_52155_new_n17682_; 
wire u2__abc_52155_new_n17683_; 
wire u2__abc_52155_new_n17684_; 
wire u2__abc_52155_new_n17685_; 
wire u2__abc_52155_new_n17686_; 
wire u2__abc_52155_new_n17688_; 
wire u2__abc_52155_new_n17689_; 
wire u2__abc_52155_new_n17690_; 
wire u2__abc_52155_new_n17691_; 
wire u2__abc_52155_new_n17692_; 
wire u2__abc_52155_new_n17693_; 
wire u2__abc_52155_new_n17694_; 
wire u2__abc_52155_new_n17695_; 
wire u2__abc_52155_new_n17697_; 
wire u2__abc_52155_new_n17698_; 
wire u2__abc_52155_new_n17699_; 
wire u2__abc_52155_new_n17700_; 
wire u2__abc_52155_new_n17701_; 
wire u2__abc_52155_new_n17703_; 
wire u2__abc_52155_new_n17704_; 
wire u2__abc_52155_new_n17705_; 
wire u2__abc_52155_new_n17706_; 
wire u2__abc_52155_new_n17707_; 
wire u2__abc_52155_new_n17709_; 
wire u2__abc_52155_new_n17710_; 
wire u2__abc_52155_new_n17711_; 
wire u2__abc_52155_new_n17712_; 
wire u2__abc_52155_new_n17713_; 
wire u2__abc_52155_new_n17715_; 
wire u2__abc_52155_new_n17716_; 
wire u2__abc_52155_new_n17717_; 
wire u2__abc_52155_new_n17718_; 
wire u2__abc_52155_new_n17719_; 
wire u2__abc_52155_new_n17721_; 
wire u2__abc_52155_new_n17722_; 
wire u2__abc_52155_new_n17723_; 
wire u2__abc_52155_new_n17724_; 
wire u2__abc_52155_new_n17725_; 
wire u2__abc_52155_new_n17727_; 
wire u2__abc_52155_new_n17728_; 
wire u2__abc_52155_new_n17729_; 
wire u2__abc_52155_new_n17730_; 
wire u2__abc_52155_new_n17731_; 
wire u2__abc_52155_new_n17733_; 
wire u2__abc_52155_new_n17734_; 
wire u2__abc_52155_new_n17735_; 
wire u2__abc_52155_new_n17736_; 
wire u2__abc_52155_new_n17737_; 
wire u2__abc_52155_new_n17739_; 
wire u2__abc_52155_new_n17740_; 
wire u2__abc_52155_new_n17741_; 
wire u2__abc_52155_new_n17742_; 
wire u2__abc_52155_new_n17743_; 
wire u2__abc_52155_new_n17745_; 
wire u2__abc_52155_new_n17746_; 
wire u2__abc_52155_new_n17747_; 
wire u2__abc_52155_new_n17748_; 
wire u2__abc_52155_new_n17749_; 
wire u2__abc_52155_new_n17750_; 
wire u2__abc_52155_new_n17751_; 
wire u2__abc_52155_new_n17752_; 
wire u2__abc_52155_new_n17754_; 
wire u2__abc_52155_new_n17755_; 
wire u2__abc_52155_new_n17756_; 
wire u2__abc_52155_new_n17757_; 
wire u2__abc_52155_new_n17758_; 
wire u2__abc_52155_new_n17760_; 
wire u2__abc_52155_new_n17761_; 
wire u2__abc_52155_new_n17762_; 
wire u2__abc_52155_new_n17763_; 
wire u2__abc_52155_new_n17764_; 
wire u2__abc_52155_new_n17766_; 
wire u2__abc_52155_new_n17767_; 
wire u2__abc_52155_new_n17768_; 
wire u2__abc_52155_new_n17769_; 
wire u2__abc_52155_new_n17770_; 
wire u2__abc_52155_new_n17772_; 
wire u2__abc_52155_new_n17773_; 
wire u2__abc_52155_new_n17774_; 
wire u2__abc_52155_new_n17775_; 
wire u2__abc_52155_new_n17776_; 
wire u2__abc_52155_new_n17778_; 
wire u2__abc_52155_new_n17779_; 
wire u2__abc_52155_new_n17780_; 
wire u2__abc_52155_new_n17781_; 
wire u2__abc_52155_new_n17782_; 
wire u2__abc_52155_new_n17784_; 
wire u2__abc_52155_new_n17785_; 
wire u2__abc_52155_new_n17786_; 
wire u2__abc_52155_new_n17787_; 
wire u2__abc_52155_new_n17788_; 
wire u2__abc_52155_new_n17790_; 
wire u2__abc_52155_new_n17791_; 
wire u2__abc_52155_new_n17792_; 
wire u2__abc_52155_new_n17793_; 
wire u2__abc_52155_new_n17794_; 
wire u2__abc_52155_new_n17796_; 
wire u2__abc_52155_new_n17797_; 
wire u2__abc_52155_new_n17798_; 
wire u2__abc_52155_new_n17799_; 
wire u2__abc_52155_new_n17800_; 
wire u2__abc_52155_new_n17802_; 
wire u2__abc_52155_new_n17803_; 
wire u2__abc_52155_new_n17804_; 
wire u2__abc_52155_new_n17805_; 
wire u2__abc_52155_new_n17806_; 
wire u2__abc_52155_new_n17808_; 
wire u2__abc_52155_new_n17809_; 
wire u2__abc_52155_new_n17810_; 
wire u2__abc_52155_new_n17811_; 
wire u2__abc_52155_new_n17812_; 
wire u2__abc_52155_new_n17814_; 
wire u2__abc_52155_new_n17815_; 
wire u2__abc_52155_new_n17816_; 
wire u2__abc_52155_new_n17817_; 
wire u2__abc_52155_new_n17818_; 
wire u2__abc_52155_new_n17820_; 
wire u2__abc_52155_new_n17821_; 
wire u2__abc_52155_new_n17822_; 
wire u2__abc_52155_new_n17823_; 
wire u2__abc_52155_new_n17824_; 
wire u2__abc_52155_new_n17826_; 
wire u2__abc_52155_new_n17827_; 
wire u2__abc_52155_new_n17828_; 
wire u2__abc_52155_new_n17829_; 
wire u2__abc_52155_new_n17830_; 
wire u2__abc_52155_new_n17832_; 
wire u2__abc_52155_new_n17833_; 
wire u2__abc_52155_new_n17834_; 
wire u2__abc_52155_new_n17835_; 
wire u2__abc_52155_new_n17836_; 
wire u2__abc_52155_new_n17838_; 
wire u2__abc_52155_new_n17839_; 
wire u2__abc_52155_new_n17840_; 
wire u2__abc_52155_new_n17841_; 
wire u2__abc_52155_new_n17842_; 
wire u2__abc_52155_new_n17844_; 
wire u2__abc_52155_new_n17845_; 
wire u2__abc_52155_new_n17846_; 
wire u2__abc_52155_new_n17847_; 
wire u2__abc_52155_new_n17848_; 
wire u2__abc_52155_new_n17850_; 
wire u2__abc_52155_new_n17851_; 
wire u2__abc_52155_new_n17852_; 
wire u2__abc_52155_new_n17853_; 
wire u2__abc_52155_new_n17854_; 
wire u2__abc_52155_new_n17856_; 
wire u2__abc_52155_new_n17857_; 
wire u2__abc_52155_new_n17858_; 
wire u2__abc_52155_new_n17859_; 
wire u2__abc_52155_new_n17860_; 
wire u2__abc_52155_new_n17862_; 
wire u2__abc_52155_new_n17863_; 
wire u2__abc_52155_new_n17864_; 
wire u2__abc_52155_new_n17865_; 
wire u2__abc_52155_new_n17866_; 
wire u2__abc_52155_new_n17868_; 
wire u2__abc_52155_new_n17869_; 
wire u2__abc_52155_new_n17870_; 
wire u2__abc_52155_new_n17871_; 
wire u2__abc_52155_new_n17872_; 
wire u2__abc_52155_new_n17874_; 
wire u2__abc_52155_new_n17875_; 
wire u2__abc_52155_new_n17876_; 
wire u2__abc_52155_new_n17877_; 
wire u2__abc_52155_new_n17878_; 
wire u2__abc_52155_new_n17880_; 
wire u2__abc_52155_new_n17881_; 
wire u2__abc_52155_new_n17882_; 
wire u2__abc_52155_new_n17883_; 
wire u2__abc_52155_new_n17884_; 
wire u2__abc_52155_new_n17886_; 
wire u2__abc_52155_new_n17887_; 
wire u2__abc_52155_new_n17888_; 
wire u2__abc_52155_new_n17889_; 
wire u2__abc_52155_new_n17890_; 
wire u2__abc_52155_new_n17891_; 
wire u2__abc_52155_new_n17892_; 
wire u2__abc_52155_new_n17893_; 
wire u2__abc_52155_new_n17895_; 
wire u2__abc_52155_new_n17896_; 
wire u2__abc_52155_new_n17897_; 
wire u2__abc_52155_new_n17898_; 
wire u2__abc_52155_new_n17899_; 
wire u2__abc_52155_new_n17900_; 
wire u2__abc_52155_new_n17901_; 
wire u2__abc_52155_new_n17902_; 
wire u2__abc_52155_new_n17904_; 
wire u2__abc_52155_new_n17905_; 
wire u2__abc_52155_new_n17906_; 
wire u2__abc_52155_new_n17907_; 
wire u2__abc_52155_new_n17908_; 
wire u2__abc_52155_new_n17910_; 
wire u2__abc_52155_new_n17911_; 
wire u2__abc_52155_new_n17912_; 
wire u2__abc_52155_new_n17913_; 
wire u2__abc_52155_new_n17914_; 
wire u2__abc_52155_new_n17916_; 
wire u2__abc_52155_new_n17917_; 
wire u2__abc_52155_new_n17918_; 
wire u2__abc_52155_new_n17919_; 
wire u2__abc_52155_new_n17920_; 
wire u2__abc_52155_new_n17922_; 
wire u2__abc_52155_new_n17923_; 
wire u2__abc_52155_new_n17924_; 
wire u2__abc_52155_new_n17925_; 
wire u2__abc_52155_new_n17926_; 
wire u2__abc_52155_new_n17928_; 
wire u2__abc_52155_new_n17929_; 
wire u2__abc_52155_new_n17930_; 
wire u2__abc_52155_new_n17931_; 
wire u2__abc_52155_new_n17932_; 
wire u2__abc_52155_new_n17934_; 
wire u2__abc_52155_new_n17935_; 
wire u2__abc_52155_new_n17936_; 
wire u2__abc_52155_new_n17937_; 
wire u2__abc_52155_new_n17938_; 
wire u2__abc_52155_new_n17940_; 
wire u2__abc_52155_new_n17941_; 
wire u2__abc_52155_new_n17942_; 
wire u2__abc_52155_new_n17943_; 
wire u2__abc_52155_new_n17944_; 
wire u2__abc_52155_new_n17946_; 
wire u2__abc_52155_new_n17947_; 
wire u2__abc_52155_new_n17948_; 
wire u2__abc_52155_new_n17949_; 
wire u2__abc_52155_new_n17950_; 
wire u2__abc_52155_new_n17952_; 
wire u2__abc_52155_new_n17953_; 
wire u2__abc_52155_new_n17954_; 
wire u2__abc_52155_new_n17955_; 
wire u2__abc_52155_new_n17956_; 
wire u2__abc_52155_new_n17958_; 
wire u2__abc_52155_new_n17959_; 
wire u2__abc_52155_new_n17960_; 
wire u2__abc_52155_new_n17961_; 
wire u2__abc_52155_new_n17962_; 
wire u2__abc_52155_new_n17964_; 
wire u2__abc_52155_new_n17965_; 
wire u2__abc_52155_new_n17966_; 
wire u2__abc_52155_new_n17967_; 
wire u2__abc_52155_new_n17968_; 
wire u2__abc_52155_new_n17970_; 
wire u2__abc_52155_new_n17971_; 
wire u2__abc_52155_new_n17972_; 
wire u2__abc_52155_new_n17973_; 
wire u2__abc_52155_new_n17974_; 
wire u2__abc_52155_new_n17976_; 
wire u2__abc_52155_new_n17977_; 
wire u2__abc_52155_new_n17978_; 
wire u2__abc_52155_new_n17979_; 
wire u2__abc_52155_new_n17980_; 
wire u2__abc_52155_new_n17982_; 
wire u2__abc_52155_new_n17983_; 
wire u2__abc_52155_new_n17984_; 
wire u2__abc_52155_new_n17985_; 
wire u2__abc_52155_new_n17986_; 
wire u2__abc_52155_new_n17987_; 
wire u2__abc_52155_new_n17988_; 
wire u2__abc_52155_new_n17989_; 
wire u2__abc_52155_new_n17991_; 
wire u2__abc_52155_new_n17992_; 
wire u2__abc_52155_new_n17993_; 
wire u2__abc_52155_new_n17994_; 
wire u2__abc_52155_new_n17995_; 
wire u2__abc_52155_new_n17997_; 
wire u2__abc_52155_new_n17998_; 
wire u2__abc_52155_new_n17999_; 
wire u2__abc_52155_new_n18000_; 
wire u2__abc_52155_new_n18001_; 
wire u2__abc_52155_new_n18003_; 
wire u2__abc_52155_new_n18004_; 
wire u2__abc_52155_new_n18005_; 
wire u2__abc_52155_new_n18006_; 
wire u2__abc_52155_new_n18007_; 
wire u2__abc_52155_new_n18009_; 
wire u2__abc_52155_new_n18010_; 
wire u2__abc_52155_new_n18011_; 
wire u2__abc_52155_new_n18012_; 
wire u2__abc_52155_new_n18013_; 
wire u2__abc_52155_new_n18015_; 
wire u2__abc_52155_new_n18016_; 
wire u2__abc_52155_new_n18017_; 
wire u2__abc_52155_new_n18018_; 
wire u2__abc_52155_new_n18019_; 
wire u2__abc_52155_new_n18021_; 
wire u2__abc_52155_new_n18022_; 
wire u2__abc_52155_new_n18023_; 
wire u2__abc_52155_new_n18024_; 
wire u2__abc_52155_new_n18025_; 
wire u2__abc_52155_new_n18027_; 
wire u2__abc_52155_new_n18028_; 
wire u2__abc_52155_new_n18029_; 
wire u2__abc_52155_new_n18030_; 
wire u2__abc_52155_new_n18031_; 
wire u2__abc_52155_new_n18033_; 
wire u2__abc_52155_new_n18034_; 
wire u2__abc_52155_new_n18035_; 
wire u2__abc_52155_new_n18036_; 
wire u2__abc_52155_new_n18037_; 
wire u2__abc_52155_new_n18039_; 
wire u2__abc_52155_new_n18040_; 
wire u2__abc_52155_new_n18041_; 
wire u2__abc_52155_new_n18042_; 
wire u2__abc_52155_new_n18043_; 
wire u2__abc_52155_new_n18045_; 
wire u2__abc_52155_new_n18046_; 
wire u2__abc_52155_new_n18047_; 
wire u2__abc_52155_new_n18048_; 
wire u2__abc_52155_new_n18049_; 
wire u2__abc_52155_new_n18051_; 
wire u2__abc_52155_new_n18052_; 
wire u2__abc_52155_new_n18053_; 
wire u2__abc_52155_new_n18054_; 
wire u2__abc_52155_new_n18055_; 
wire u2__abc_52155_new_n18057_; 
wire u2__abc_52155_new_n18058_; 
wire u2__abc_52155_new_n18059_; 
wire u2__abc_52155_new_n18060_; 
wire u2__abc_52155_new_n18061_; 
wire u2__abc_52155_new_n18063_; 
wire u2__abc_52155_new_n18064_; 
wire u2__abc_52155_new_n18065_; 
wire u2__abc_52155_new_n18066_; 
wire u2__abc_52155_new_n18067_; 
wire u2__abc_52155_new_n18069_; 
wire u2__abc_52155_new_n18070_; 
wire u2__abc_52155_new_n18071_; 
wire u2__abc_52155_new_n18072_; 
wire u2__abc_52155_new_n18073_; 
wire u2__abc_52155_new_n18075_; 
wire u2__abc_52155_new_n18076_; 
wire u2__abc_52155_new_n18077_; 
wire u2__abc_52155_new_n18078_; 
wire u2__abc_52155_new_n18079_; 
wire u2__abc_52155_new_n18081_; 
wire u2__abc_52155_new_n18082_; 
wire u2__abc_52155_new_n18083_; 
wire u2__abc_52155_new_n18084_; 
wire u2__abc_52155_new_n18085_; 
wire u2__abc_52155_new_n18087_; 
wire u2__abc_52155_new_n18088_; 
wire u2__abc_52155_new_n18089_; 
wire u2__abc_52155_new_n18090_; 
wire u2__abc_52155_new_n18091_; 
wire u2__abc_52155_new_n18092_; 
wire u2__abc_52155_new_n18093_; 
wire u2__abc_52155_new_n18094_; 
wire u2__abc_52155_new_n18096_; 
wire u2__abc_52155_new_n18097_; 
wire u2__abc_52155_new_n18098_; 
wire u2__abc_52155_new_n18099_; 
wire u2__abc_52155_new_n18101_; 
wire u2__abc_52155_new_n18102_; 
wire u2__abc_52155_new_n18103_; 
wire u2__abc_52155_new_n18104_; 
wire u2__abc_52155_new_n18106_; 
wire u2__abc_52155_new_n18107_; 
wire u2__abc_52155_new_n18108_; 
wire u2__abc_52155_new_n18109_; 
wire u2__abc_52155_new_n18111_; 
wire u2__abc_52155_new_n18112_; 
wire u2__abc_52155_new_n18113_; 
wire u2__abc_52155_new_n18114_; 
wire u2__abc_52155_new_n18116_; 
wire u2__abc_52155_new_n18117_; 
wire u2__abc_52155_new_n18118_; 
wire u2__abc_52155_new_n18119_; 
wire u2__abc_52155_new_n18121_; 
wire u2__abc_52155_new_n18122_; 
wire u2__abc_52155_new_n18123_; 
wire u2__abc_52155_new_n18124_; 
wire u2__abc_52155_new_n18126_; 
wire u2__abc_52155_new_n18127_; 
wire u2__abc_52155_new_n18128_; 
wire u2__abc_52155_new_n18129_; 
wire u2__abc_52155_new_n18131_; 
wire u2__abc_52155_new_n18132_; 
wire u2__abc_52155_new_n18133_; 
wire u2__abc_52155_new_n18134_; 
wire u2__abc_52155_new_n18136_; 
wire u2__abc_52155_new_n18137_; 
wire u2__abc_52155_new_n18138_; 
wire u2__abc_52155_new_n18139_; 
wire u2__abc_52155_new_n18141_; 
wire u2__abc_52155_new_n18142_; 
wire u2__abc_52155_new_n18143_; 
wire u2__abc_52155_new_n18144_; 
wire u2__abc_52155_new_n18146_; 
wire u2__abc_52155_new_n18147_; 
wire u2__abc_52155_new_n18148_; 
wire u2__abc_52155_new_n18149_; 
wire u2__abc_52155_new_n18151_; 
wire u2__abc_52155_new_n18152_; 
wire u2__abc_52155_new_n18153_; 
wire u2__abc_52155_new_n18154_; 
wire u2__abc_52155_new_n18156_; 
wire u2__abc_52155_new_n18157_; 
wire u2__abc_52155_new_n18158_; 
wire u2__abc_52155_new_n18159_; 
wire u2__abc_52155_new_n18161_; 
wire u2__abc_52155_new_n18162_; 
wire u2__abc_52155_new_n18163_; 
wire u2__abc_52155_new_n18164_; 
wire u2__abc_52155_new_n18166_; 
wire u2__abc_52155_new_n18167_; 
wire u2__abc_52155_new_n18168_; 
wire u2__abc_52155_new_n18169_; 
wire u2__abc_52155_new_n18171_; 
wire u2__abc_52155_new_n18172_; 
wire u2__abc_52155_new_n18173_; 
wire u2__abc_52155_new_n18174_; 
wire u2__abc_52155_new_n18176_; 
wire u2__abc_52155_new_n18177_; 
wire u2__abc_52155_new_n18178_; 
wire u2__abc_52155_new_n18179_; 
wire u2__abc_52155_new_n18181_; 
wire u2__abc_52155_new_n18182_; 
wire u2__abc_52155_new_n18183_; 
wire u2__abc_52155_new_n18184_; 
wire u2__abc_52155_new_n18186_; 
wire u2__abc_52155_new_n18187_; 
wire u2__abc_52155_new_n18188_; 
wire u2__abc_52155_new_n18189_; 
wire u2__abc_52155_new_n18191_; 
wire u2__abc_52155_new_n18192_; 
wire u2__abc_52155_new_n18193_; 
wire u2__abc_52155_new_n18194_; 
wire u2__abc_52155_new_n18196_; 
wire u2__abc_52155_new_n18197_; 
wire u2__abc_52155_new_n18198_; 
wire u2__abc_52155_new_n18199_; 
wire u2__abc_52155_new_n18201_; 
wire u2__abc_52155_new_n18202_; 
wire u2__abc_52155_new_n18203_; 
wire u2__abc_52155_new_n18204_; 
wire u2__abc_52155_new_n18206_; 
wire u2__abc_52155_new_n18207_; 
wire u2__abc_52155_new_n18208_; 
wire u2__abc_52155_new_n18209_; 
wire u2__abc_52155_new_n18211_; 
wire u2__abc_52155_new_n18212_; 
wire u2__abc_52155_new_n18213_; 
wire u2__abc_52155_new_n18214_; 
wire u2__abc_52155_new_n18216_; 
wire u2__abc_52155_new_n18217_; 
wire u2__abc_52155_new_n18218_; 
wire u2__abc_52155_new_n18219_; 
wire u2__abc_52155_new_n18221_; 
wire u2__abc_52155_new_n18222_; 
wire u2__abc_52155_new_n18223_; 
wire u2__abc_52155_new_n18224_; 
wire u2__abc_52155_new_n18226_; 
wire u2__abc_52155_new_n18227_; 
wire u2__abc_52155_new_n18228_; 
wire u2__abc_52155_new_n18229_; 
wire u2__abc_52155_new_n18231_; 
wire u2__abc_52155_new_n18232_; 
wire u2__abc_52155_new_n18233_; 
wire u2__abc_52155_new_n18234_; 
wire u2__abc_52155_new_n18236_; 
wire u2__abc_52155_new_n18237_; 
wire u2__abc_52155_new_n18238_; 
wire u2__abc_52155_new_n18239_; 
wire u2__abc_52155_new_n18241_; 
wire u2__abc_52155_new_n18242_; 
wire u2__abc_52155_new_n18243_; 
wire u2__abc_52155_new_n18244_; 
wire u2__abc_52155_new_n18246_; 
wire u2__abc_52155_new_n18247_; 
wire u2__abc_52155_new_n18248_; 
wire u2__abc_52155_new_n18249_; 
wire u2__abc_52155_new_n18251_; 
wire u2__abc_52155_new_n18252_; 
wire u2__abc_52155_new_n18253_; 
wire u2__abc_52155_new_n18254_; 
wire u2__abc_52155_new_n18256_; 
wire u2__abc_52155_new_n18257_; 
wire u2__abc_52155_new_n18258_; 
wire u2__abc_52155_new_n18259_; 
wire u2__abc_52155_new_n18261_; 
wire u2__abc_52155_new_n18262_; 
wire u2__abc_52155_new_n18263_; 
wire u2__abc_52155_new_n18264_; 
wire u2__abc_52155_new_n18266_; 
wire u2__abc_52155_new_n18267_; 
wire u2__abc_52155_new_n18268_; 
wire u2__abc_52155_new_n18269_; 
wire u2__abc_52155_new_n18271_; 
wire u2__abc_52155_new_n18272_; 
wire u2__abc_52155_new_n18273_; 
wire u2__abc_52155_new_n18274_; 
wire u2__abc_52155_new_n18276_; 
wire u2__abc_52155_new_n18277_; 
wire u2__abc_52155_new_n18278_; 
wire u2__abc_52155_new_n18279_; 
wire u2__abc_52155_new_n18281_; 
wire u2__abc_52155_new_n18282_; 
wire u2__abc_52155_new_n18283_; 
wire u2__abc_52155_new_n18284_; 
wire u2__abc_52155_new_n18286_; 
wire u2__abc_52155_new_n18287_; 
wire u2__abc_52155_new_n18288_; 
wire u2__abc_52155_new_n18289_; 
wire u2__abc_52155_new_n18291_; 
wire u2__abc_52155_new_n18292_; 
wire u2__abc_52155_new_n18293_; 
wire u2__abc_52155_new_n18294_; 
wire u2__abc_52155_new_n18296_; 
wire u2__abc_52155_new_n18297_; 
wire u2__abc_52155_new_n18298_; 
wire u2__abc_52155_new_n18299_; 
wire u2__abc_52155_new_n18301_; 
wire u2__abc_52155_new_n18302_; 
wire u2__abc_52155_new_n18303_; 
wire u2__abc_52155_new_n18304_; 
wire u2__abc_52155_new_n18306_; 
wire u2__abc_52155_new_n18307_; 
wire u2__abc_52155_new_n18308_; 
wire u2__abc_52155_new_n18309_; 
wire u2__abc_52155_new_n18311_; 
wire u2__abc_52155_new_n18312_; 
wire u2__abc_52155_new_n18313_; 
wire u2__abc_52155_new_n18314_; 
wire u2__abc_52155_new_n18316_; 
wire u2__abc_52155_new_n18317_; 
wire u2__abc_52155_new_n18318_; 
wire u2__abc_52155_new_n18319_; 
wire u2__abc_52155_new_n18321_; 
wire u2__abc_52155_new_n18322_; 
wire u2__abc_52155_new_n18323_; 
wire u2__abc_52155_new_n18324_; 
wire u2__abc_52155_new_n18326_; 
wire u2__abc_52155_new_n18327_; 
wire u2__abc_52155_new_n18328_; 
wire u2__abc_52155_new_n18329_; 
wire u2__abc_52155_new_n18331_; 
wire u2__abc_52155_new_n18332_; 
wire u2__abc_52155_new_n18333_; 
wire u2__abc_52155_new_n18334_; 
wire u2__abc_52155_new_n18336_; 
wire u2__abc_52155_new_n18337_; 
wire u2__abc_52155_new_n18338_; 
wire u2__abc_52155_new_n18339_; 
wire u2__abc_52155_new_n18341_; 
wire u2__abc_52155_new_n18342_; 
wire u2__abc_52155_new_n18343_; 
wire u2__abc_52155_new_n18344_; 
wire u2__abc_52155_new_n18346_; 
wire u2__abc_52155_new_n18347_; 
wire u2__abc_52155_new_n18348_; 
wire u2__abc_52155_new_n18349_; 
wire u2__abc_52155_new_n18351_; 
wire u2__abc_52155_new_n18352_; 
wire u2__abc_52155_new_n18353_; 
wire u2__abc_52155_new_n18354_; 
wire u2__abc_52155_new_n18356_; 
wire u2__abc_52155_new_n18357_; 
wire u2__abc_52155_new_n18358_; 
wire u2__abc_52155_new_n18359_; 
wire u2__abc_52155_new_n18361_; 
wire u2__abc_52155_new_n18362_; 
wire u2__abc_52155_new_n18363_; 
wire u2__abc_52155_new_n18364_; 
wire u2__abc_52155_new_n18366_; 
wire u2__abc_52155_new_n18367_; 
wire u2__abc_52155_new_n18368_; 
wire u2__abc_52155_new_n18369_; 
wire u2__abc_52155_new_n18371_; 
wire u2__abc_52155_new_n18372_; 
wire u2__abc_52155_new_n18373_; 
wire u2__abc_52155_new_n18374_; 
wire u2__abc_52155_new_n18376_; 
wire u2__abc_52155_new_n18377_; 
wire u2__abc_52155_new_n18378_; 
wire u2__abc_52155_new_n18379_; 
wire u2__abc_52155_new_n18381_; 
wire u2__abc_52155_new_n18382_; 
wire u2__abc_52155_new_n18383_; 
wire u2__abc_52155_new_n18384_; 
wire u2__abc_52155_new_n18386_; 
wire u2__abc_52155_new_n18387_; 
wire u2__abc_52155_new_n18388_; 
wire u2__abc_52155_new_n18389_; 
wire u2__abc_52155_new_n18391_; 
wire u2__abc_52155_new_n18392_; 
wire u2__abc_52155_new_n18393_; 
wire u2__abc_52155_new_n18394_; 
wire u2__abc_52155_new_n18396_; 
wire u2__abc_52155_new_n18397_; 
wire u2__abc_52155_new_n18398_; 
wire u2__abc_52155_new_n18399_; 
wire u2__abc_52155_new_n18401_; 
wire u2__abc_52155_new_n18402_; 
wire u2__abc_52155_new_n18403_; 
wire u2__abc_52155_new_n18404_; 
wire u2__abc_52155_new_n18406_; 
wire u2__abc_52155_new_n18407_; 
wire u2__abc_52155_new_n18408_; 
wire u2__abc_52155_new_n18409_; 
wire u2__abc_52155_new_n18411_; 
wire u2__abc_52155_new_n18412_; 
wire u2__abc_52155_new_n18413_; 
wire u2__abc_52155_new_n18414_; 
wire u2__abc_52155_new_n18416_; 
wire u2__abc_52155_new_n18417_; 
wire u2__abc_52155_new_n18418_; 
wire u2__abc_52155_new_n18419_; 
wire u2__abc_52155_new_n18421_; 
wire u2__abc_52155_new_n18422_; 
wire u2__abc_52155_new_n18423_; 
wire u2__abc_52155_new_n18424_; 
wire u2__abc_52155_new_n18426_; 
wire u2__abc_52155_new_n18427_; 
wire u2__abc_52155_new_n18428_; 
wire u2__abc_52155_new_n18429_; 
wire u2__abc_52155_new_n18431_; 
wire u2__abc_52155_new_n18432_; 
wire u2__abc_52155_new_n18433_; 
wire u2__abc_52155_new_n18434_; 
wire u2__abc_52155_new_n18436_; 
wire u2__abc_52155_new_n18437_; 
wire u2__abc_52155_new_n18438_; 
wire u2__abc_52155_new_n18439_; 
wire u2__abc_52155_new_n18441_; 
wire u2__abc_52155_new_n18442_; 
wire u2__abc_52155_new_n18443_; 
wire u2__abc_52155_new_n18444_; 
wire u2__abc_52155_new_n18446_; 
wire u2__abc_52155_new_n18447_; 
wire u2__abc_52155_new_n18448_; 
wire u2__abc_52155_new_n18449_; 
wire u2__abc_52155_new_n18451_; 
wire u2__abc_52155_new_n18452_; 
wire u2__abc_52155_new_n18453_; 
wire u2__abc_52155_new_n18454_; 
wire u2__abc_52155_new_n18456_; 
wire u2__abc_52155_new_n18457_; 
wire u2__abc_52155_new_n18458_; 
wire u2__abc_52155_new_n18459_; 
wire u2__abc_52155_new_n18461_; 
wire u2__abc_52155_new_n18462_; 
wire u2__abc_52155_new_n18463_; 
wire u2__abc_52155_new_n18464_; 
wire u2__abc_52155_new_n18466_; 
wire u2__abc_52155_new_n18467_; 
wire u2__abc_52155_new_n18468_; 
wire u2__abc_52155_new_n18469_; 
wire u2__abc_52155_new_n18471_; 
wire u2__abc_52155_new_n18472_; 
wire u2__abc_52155_new_n18473_; 
wire u2__abc_52155_new_n18474_; 
wire u2__abc_52155_new_n18476_; 
wire u2__abc_52155_new_n18477_; 
wire u2__abc_52155_new_n18478_; 
wire u2__abc_52155_new_n18479_; 
wire u2__abc_52155_new_n18481_; 
wire u2__abc_52155_new_n18482_; 
wire u2__abc_52155_new_n18483_; 
wire u2__abc_52155_new_n18484_; 
wire u2__abc_52155_new_n18486_; 
wire u2__abc_52155_new_n18487_; 
wire u2__abc_52155_new_n18488_; 
wire u2__abc_52155_new_n18489_; 
wire u2__abc_52155_new_n18491_; 
wire u2__abc_52155_new_n18492_; 
wire u2__abc_52155_new_n18493_; 
wire u2__abc_52155_new_n18494_; 
wire u2__abc_52155_new_n18496_; 
wire u2__abc_52155_new_n18497_; 
wire u2__abc_52155_new_n18498_; 
wire u2__abc_52155_new_n18499_; 
wire u2__abc_52155_new_n18501_; 
wire u2__abc_52155_new_n18502_; 
wire u2__abc_52155_new_n18503_; 
wire u2__abc_52155_new_n18504_; 
wire u2__abc_52155_new_n18506_; 
wire u2__abc_52155_new_n18507_; 
wire u2__abc_52155_new_n18508_; 
wire u2__abc_52155_new_n18509_; 
wire u2__abc_52155_new_n18511_; 
wire u2__abc_52155_new_n18512_; 
wire u2__abc_52155_new_n18513_; 
wire u2__abc_52155_new_n18514_; 
wire u2__abc_52155_new_n18516_; 
wire u2__abc_52155_new_n18517_; 
wire u2__abc_52155_new_n18518_; 
wire u2__abc_52155_new_n18519_; 
wire u2__abc_52155_new_n18521_; 
wire u2__abc_52155_new_n18522_; 
wire u2__abc_52155_new_n18523_; 
wire u2__abc_52155_new_n18524_; 
wire u2__abc_52155_new_n18526_; 
wire u2__abc_52155_new_n18527_; 
wire u2__abc_52155_new_n18528_; 
wire u2__abc_52155_new_n18529_; 
wire u2__abc_52155_new_n18531_; 
wire u2__abc_52155_new_n18532_; 
wire u2__abc_52155_new_n18533_; 
wire u2__abc_52155_new_n18534_; 
wire u2__abc_52155_new_n18536_; 
wire u2__abc_52155_new_n18537_; 
wire u2__abc_52155_new_n18538_; 
wire u2__abc_52155_new_n18539_; 
wire u2__abc_52155_new_n18541_; 
wire u2__abc_52155_new_n18542_; 
wire u2__abc_52155_new_n18543_; 
wire u2__abc_52155_new_n18544_; 
wire u2__abc_52155_new_n18546_; 
wire u2__abc_52155_new_n18547_; 
wire u2__abc_52155_new_n18548_; 
wire u2__abc_52155_new_n18549_; 
wire u2__abc_52155_new_n18551_; 
wire u2__abc_52155_new_n18552_; 
wire u2__abc_52155_new_n18553_; 
wire u2__abc_52155_new_n18554_; 
wire u2__abc_52155_new_n18556_; 
wire u2__abc_52155_new_n18557_; 
wire u2__abc_52155_new_n18558_; 
wire u2__abc_52155_new_n18559_; 
wire u2__abc_52155_new_n18561_; 
wire u2__abc_52155_new_n18562_; 
wire u2__abc_52155_new_n18563_; 
wire u2__abc_52155_new_n18564_; 
wire u2__abc_52155_new_n18566_; 
wire u2__abc_52155_new_n18567_; 
wire u2__abc_52155_new_n18568_; 
wire u2__abc_52155_new_n18569_; 
wire u2__abc_52155_new_n18571_; 
wire u2__abc_52155_new_n18572_; 
wire u2__abc_52155_new_n18573_; 
wire u2__abc_52155_new_n18574_; 
wire u2__abc_52155_new_n18576_; 
wire u2__abc_52155_new_n18577_; 
wire u2__abc_52155_new_n18578_; 
wire u2__abc_52155_new_n18579_; 
wire u2__abc_52155_new_n18581_; 
wire u2__abc_52155_new_n18582_; 
wire u2__abc_52155_new_n18583_; 
wire u2__abc_52155_new_n18584_; 
wire u2__abc_52155_new_n18586_; 
wire u2__abc_52155_new_n18587_; 
wire u2__abc_52155_new_n18588_; 
wire u2__abc_52155_new_n18589_; 
wire u2__abc_52155_new_n18591_; 
wire u2__abc_52155_new_n18592_; 
wire u2__abc_52155_new_n18593_; 
wire u2__abc_52155_new_n18594_; 
wire u2__abc_52155_new_n18596_; 
wire u2__abc_52155_new_n18597_; 
wire u2__abc_52155_new_n18598_; 
wire u2__abc_52155_new_n18599_; 
wire u2__abc_52155_new_n18601_; 
wire u2__abc_52155_new_n18602_; 
wire u2__abc_52155_new_n18603_; 
wire u2__abc_52155_new_n18604_; 
wire u2__abc_52155_new_n18606_; 
wire u2__abc_52155_new_n18607_; 
wire u2__abc_52155_new_n18608_; 
wire u2__abc_52155_new_n18609_; 
wire u2__abc_52155_new_n18611_; 
wire u2__abc_52155_new_n18612_; 
wire u2__abc_52155_new_n18613_; 
wire u2__abc_52155_new_n18614_; 
wire u2__abc_52155_new_n18616_; 
wire u2__abc_52155_new_n18617_; 
wire u2__abc_52155_new_n18618_; 
wire u2__abc_52155_new_n18619_; 
wire u2__abc_52155_new_n18621_; 
wire u2__abc_52155_new_n18622_; 
wire u2__abc_52155_new_n18623_; 
wire u2__abc_52155_new_n18624_; 
wire u2__abc_52155_new_n18626_; 
wire u2__abc_52155_new_n18627_; 
wire u2__abc_52155_new_n18628_; 
wire u2__abc_52155_new_n18629_; 
wire u2__abc_52155_new_n18631_; 
wire u2__abc_52155_new_n18632_; 
wire u2__abc_52155_new_n18633_; 
wire u2__abc_52155_new_n18634_; 
wire u2__abc_52155_new_n18636_; 
wire u2__abc_52155_new_n18637_; 
wire u2__abc_52155_new_n18638_; 
wire u2__abc_52155_new_n18639_; 
wire u2__abc_52155_new_n18641_; 
wire u2__abc_52155_new_n18642_; 
wire u2__abc_52155_new_n18643_; 
wire u2__abc_52155_new_n18644_; 
wire u2__abc_52155_new_n18646_; 
wire u2__abc_52155_new_n18647_; 
wire u2__abc_52155_new_n18648_; 
wire u2__abc_52155_new_n18649_; 
wire u2__abc_52155_new_n18651_; 
wire u2__abc_52155_new_n18652_; 
wire u2__abc_52155_new_n18653_; 
wire u2__abc_52155_new_n18654_; 
wire u2__abc_52155_new_n18656_; 
wire u2__abc_52155_new_n18657_; 
wire u2__abc_52155_new_n18658_; 
wire u2__abc_52155_new_n18659_; 
wire u2__abc_52155_new_n18661_; 
wire u2__abc_52155_new_n18662_; 
wire u2__abc_52155_new_n18663_; 
wire u2__abc_52155_new_n18664_; 
wire u2__abc_52155_new_n18666_; 
wire u2__abc_52155_new_n18667_; 
wire u2__abc_52155_new_n18668_; 
wire u2__abc_52155_new_n18669_; 
wire u2__abc_52155_new_n18671_; 
wire u2__abc_52155_new_n18672_; 
wire u2__abc_52155_new_n18673_; 
wire u2__abc_52155_new_n18674_; 
wire u2__abc_52155_new_n18676_; 
wire u2__abc_52155_new_n18677_; 
wire u2__abc_52155_new_n18678_; 
wire u2__abc_52155_new_n18679_; 
wire u2__abc_52155_new_n18681_; 
wire u2__abc_52155_new_n18682_; 
wire u2__abc_52155_new_n18683_; 
wire u2__abc_52155_new_n18684_; 
wire u2__abc_52155_new_n18686_; 
wire u2__abc_52155_new_n18687_; 
wire u2__abc_52155_new_n18688_; 
wire u2__abc_52155_new_n18689_; 
wire u2__abc_52155_new_n18691_; 
wire u2__abc_52155_new_n18692_; 
wire u2__abc_52155_new_n18693_; 
wire u2__abc_52155_new_n18694_; 
wire u2__abc_52155_new_n18696_; 
wire u2__abc_52155_new_n18697_; 
wire u2__abc_52155_new_n18698_; 
wire u2__abc_52155_new_n18699_; 
wire u2__abc_52155_new_n18701_; 
wire u2__abc_52155_new_n18702_; 
wire u2__abc_52155_new_n18703_; 
wire u2__abc_52155_new_n18704_; 
wire u2__abc_52155_new_n18706_; 
wire u2__abc_52155_new_n18707_; 
wire u2__abc_52155_new_n18708_; 
wire u2__abc_52155_new_n18709_; 
wire u2__abc_52155_new_n18711_; 
wire u2__abc_52155_new_n18712_; 
wire u2__abc_52155_new_n18713_; 
wire u2__abc_52155_new_n18714_; 
wire u2__abc_52155_new_n18716_; 
wire u2__abc_52155_new_n18717_; 
wire u2__abc_52155_new_n18718_; 
wire u2__abc_52155_new_n18719_; 
wire u2__abc_52155_new_n18721_; 
wire u2__abc_52155_new_n18722_; 
wire u2__abc_52155_new_n18723_; 
wire u2__abc_52155_new_n18724_; 
wire u2__abc_52155_new_n18726_; 
wire u2__abc_52155_new_n18727_; 
wire u2__abc_52155_new_n18728_; 
wire u2__abc_52155_new_n18729_; 
wire u2__abc_52155_new_n18731_; 
wire u2__abc_52155_new_n18732_; 
wire u2__abc_52155_new_n18733_; 
wire u2__abc_52155_new_n18734_; 
wire u2__abc_52155_new_n18736_; 
wire u2__abc_52155_new_n18737_; 
wire u2__abc_52155_new_n18738_; 
wire u2__abc_52155_new_n18739_; 
wire u2__abc_52155_new_n18741_; 
wire u2__abc_52155_new_n18742_; 
wire u2__abc_52155_new_n18743_; 
wire u2__abc_52155_new_n18744_; 
wire u2__abc_52155_new_n18746_; 
wire u2__abc_52155_new_n18747_; 
wire u2__abc_52155_new_n18748_; 
wire u2__abc_52155_new_n18749_; 
wire u2__abc_52155_new_n18751_; 
wire u2__abc_52155_new_n18752_; 
wire u2__abc_52155_new_n18753_; 
wire u2__abc_52155_new_n18754_; 
wire u2__abc_52155_new_n18756_; 
wire u2__abc_52155_new_n18757_; 
wire u2__abc_52155_new_n18758_; 
wire u2__abc_52155_new_n18759_; 
wire u2__abc_52155_new_n18761_; 
wire u2__abc_52155_new_n18762_; 
wire u2__abc_52155_new_n18763_; 
wire u2__abc_52155_new_n18764_; 
wire u2__abc_52155_new_n18766_; 
wire u2__abc_52155_new_n18767_; 
wire u2__abc_52155_new_n18768_; 
wire u2__abc_52155_new_n18769_; 
wire u2__abc_52155_new_n18771_; 
wire u2__abc_52155_new_n18772_; 
wire u2__abc_52155_new_n18773_; 
wire u2__abc_52155_new_n18774_; 
wire u2__abc_52155_new_n18776_; 
wire u2__abc_52155_new_n18777_; 
wire u2__abc_52155_new_n18778_; 
wire u2__abc_52155_new_n18779_; 
wire u2__abc_52155_new_n18781_; 
wire u2__abc_52155_new_n18782_; 
wire u2__abc_52155_new_n18783_; 
wire u2__abc_52155_new_n18784_; 
wire u2__abc_52155_new_n18786_; 
wire u2__abc_52155_new_n18787_; 
wire u2__abc_52155_new_n18788_; 
wire u2__abc_52155_new_n18789_; 
wire u2__abc_52155_new_n18791_; 
wire u2__abc_52155_new_n18792_; 
wire u2__abc_52155_new_n18793_; 
wire u2__abc_52155_new_n18794_; 
wire u2__abc_52155_new_n18796_; 
wire u2__abc_52155_new_n18797_; 
wire u2__abc_52155_new_n18798_; 
wire u2__abc_52155_new_n18799_; 
wire u2__abc_52155_new_n18801_; 
wire u2__abc_52155_new_n18802_; 
wire u2__abc_52155_new_n18803_; 
wire u2__abc_52155_new_n18804_; 
wire u2__abc_52155_new_n18806_; 
wire u2__abc_52155_new_n18807_; 
wire u2__abc_52155_new_n18808_; 
wire u2__abc_52155_new_n18809_; 
wire u2__abc_52155_new_n18811_; 
wire u2__abc_52155_new_n18812_; 
wire u2__abc_52155_new_n18813_; 
wire u2__abc_52155_new_n18814_; 
wire u2__abc_52155_new_n18816_; 
wire u2__abc_52155_new_n18817_; 
wire u2__abc_52155_new_n18818_; 
wire u2__abc_52155_new_n18819_; 
wire u2__abc_52155_new_n18821_; 
wire u2__abc_52155_new_n18822_; 
wire u2__abc_52155_new_n18823_; 
wire u2__abc_52155_new_n18824_; 
wire u2__abc_52155_new_n18826_; 
wire u2__abc_52155_new_n18827_; 
wire u2__abc_52155_new_n18828_; 
wire u2__abc_52155_new_n18829_; 
wire u2__abc_52155_new_n18831_; 
wire u2__abc_52155_new_n18832_; 
wire u2__abc_52155_new_n18833_; 
wire u2__abc_52155_new_n18834_; 
wire u2__abc_52155_new_n18836_; 
wire u2__abc_52155_new_n18837_; 
wire u2__abc_52155_new_n18838_; 
wire u2__abc_52155_new_n18839_; 
wire u2__abc_52155_new_n18841_; 
wire u2__abc_52155_new_n18842_; 
wire u2__abc_52155_new_n18843_; 
wire u2__abc_52155_new_n18844_; 
wire u2__abc_52155_new_n18846_; 
wire u2__abc_52155_new_n18847_; 
wire u2__abc_52155_new_n18848_; 
wire u2__abc_52155_new_n18849_; 
wire u2__abc_52155_new_n18851_; 
wire u2__abc_52155_new_n18852_; 
wire u2__abc_52155_new_n18853_; 
wire u2__abc_52155_new_n18854_; 
wire u2__abc_52155_new_n18856_; 
wire u2__abc_52155_new_n18857_; 
wire u2__abc_52155_new_n18858_; 
wire u2__abc_52155_new_n18859_; 
wire u2__abc_52155_new_n18861_; 
wire u2__abc_52155_new_n18862_; 
wire u2__abc_52155_new_n18863_; 
wire u2__abc_52155_new_n18864_; 
wire u2__abc_52155_new_n18866_; 
wire u2__abc_52155_new_n18867_; 
wire u2__abc_52155_new_n18868_; 
wire u2__abc_52155_new_n18869_; 
wire u2__abc_52155_new_n18871_; 
wire u2__abc_52155_new_n18872_; 
wire u2__abc_52155_new_n18873_; 
wire u2__abc_52155_new_n18874_; 
wire u2__abc_52155_new_n18876_; 
wire u2__abc_52155_new_n18877_; 
wire u2__abc_52155_new_n18878_; 
wire u2__abc_52155_new_n18879_; 
wire u2__abc_52155_new_n18881_; 
wire u2__abc_52155_new_n18882_; 
wire u2__abc_52155_new_n18883_; 
wire u2__abc_52155_new_n18884_; 
wire u2__abc_52155_new_n18886_; 
wire u2__abc_52155_new_n18887_; 
wire u2__abc_52155_new_n18888_; 
wire u2__abc_52155_new_n18889_; 
wire u2__abc_52155_new_n18891_; 
wire u2__abc_52155_new_n18892_; 
wire u2__abc_52155_new_n18893_; 
wire u2__abc_52155_new_n18894_; 
wire u2__abc_52155_new_n18896_; 
wire u2__abc_52155_new_n18897_; 
wire u2__abc_52155_new_n18898_; 
wire u2__abc_52155_new_n18899_; 
wire u2__abc_52155_new_n18901_; 
wire u2__abc_52155_new_n18902_; 
wire u2__abc_52155_new_n18903_; 
wire u2__abc_52155_new_n18904_; 
wire u2__abc_52155_new_n18906_; 
wire u2__abc_52155_new_n18907_; 
wire u2__abc_52155_new_n18908_; 
wire u2__abc_52155_new_n18909_; 
wire u2__abc_52155_new_n18911_; 
wire u2__abc_52155_new_n18912_; 
wire u2__abc_52155_new_n18913_; 
wire u2__abc_52155_new_n18914_; 
wire u2__abc_52155_new_n18916_; 
wire u2__abc_52155_new_n18917_; 
wire u2__abc_52155_new_n18918_; 
wire u2__abc_52155_new_n18919_; 
wire u2__abc_52155_new_n18921_; 
wire u2__abc_52155_new_n18922_; 
wire u2__abc_52155_new_n18923_; 
wire u2__abc_52155_new_n18924_; 
wire u2__abc_52155_new_n18926_; 
wire u2__abc_52155_new_n18927_; 
wire u2__abc_52155_new_n18928_; 
wire u2__abc_52155_new_n18929_; 
wire u2__abc_52155_new_n18931_; 
wire u2__abc_52155_new_n18932_; 
wire u2__abc_52155_new_n18933_; 
wire u2__abc_52155_new_n18934_; 
wire u2__abc_52155_new_n18936_; 
wire u2__abc_52155_new_n18937_; 
wire u2__abc_52155_new_n18938_; 
wire u2__abc_52155_new_n18939_; 
wire u2__abc_52155_new_n18941_; 
wire u2__abc_52155_new_n18942_; 
wire u2__abc_52155_new_n18943_; 
wire u2__abc_52155_new_n18944_; 
wire u2__abc_52155_new_n18946_; 
wire u2__abc_52155_new_n18947_; 
wire u2__abc_52155_new_n18948_; 
wire u2__abc_52155_new_n18949_; 
wire u2__abc_52155_new_n18951_; 
wire u2__abc_52155_new_n18952_; 
wire u2__abc_52155_new_n18953_; 
wire u2__abc_52155_new_n18954_; 
wire u2__abc_52155_new_n18956_; 
wire u2__abc_52155_new_n18957_; 
wire u2__abc_52155_new_n18958_; 
wire u2__abc_52155_new_n18959_; 
wire u2__abc_52155_new_n18961_; 
wire u2__abc_52155_new_n18962_; 
wire u2__abc_52155_new_n18963_; 
wire u2__abc_52155_new_n18964_; 
wire u2__abc_52155_new_n18966_; 
wire u2__abc_52155_new_n18967_; 
wire u2__abc_52155_new_n18968_; 
wire u2__abc_52155_new_n18969_; 
wire u2__abc_52155_new_n18971_; 
wire u2__abc_52155_new_n18972_; 
wire u2__abc_52155_new_n18973_; 
wire u2__abc_52155_new_n18974_; 
wire u2__abc_52155_new_n18976_; 
wire u2__abc_52155_new_n18977_; 
wire u2__abc_52155_new_n18978_; 
wire u2__abc_52155_new_n18979_; 
wire u2__abc_52155_new_n18981_; 
wire u2__abc_52155_new_n18982_; 
wire u2__abc_52155_new_n18983_; 
wire u2__abc_52155_new_n18984_; 
wire u2__abc_52155_new_n18986_; 
wire u2__abc_52155_new_n18987_; 
wire u2__abc_52155_new_n18988_; 
wire u2__abc_52155_new_n18989_; 
wire u2__abc_52155_new_n18991_; 
wire u2__abc_52155_new_n18992_; 
wire u2__abc_52155_new_n18993_; 
wire u2__abc_52155_new_n18994_; 
wire u2__abc_52155_new_n18996_; 
wire u2__abc_52155_new_n18997_; 
wire u2__abc_52155_new_n18998_; 
wire u2__abc_52155_new_n18999_; 
wire u2__abc_52155_new_n19001_; 
wire u2__abc_52155_new_n19002_; 
wire u2__abc_52155_new_n19003_; 
wire u2__abc_52155_new_n19004_; 
wire u2__abc_52155_new_n19006_; 
wire u2__abc_52155_new_n19007_; 
wire u2__abc_52155_new_n19008_; 
wire u2__abc_52155_new_n19009_; 
wire u2__abc_52155_new_n19011_; 
wire u2__abc_52155_new_n19012_; 
wire u2__abc_52155_new_n19013_; 
wire u2__abc_52155_new_n19014_; 
wire u2__abc_52155_new_n19016_; 
wire u2__abc_52155_new_n19017_; 
wire u2__abc_52155_new_n19018_; 
wire u2__abc_52155_new_n19019_; 
wire u2__abc_52155_new_n19021_; 
wire u2__abc_52155_new_n19022_; 
wire u2__abc_52155_new_n19023_; 
wire u2__abc_52155_new_n19024_; 
wire u2__abc_52155_new_n19026_; 
wire u2__abc_52155_new_n19027_; 
wire u2__abc_52155_new_n19028_; 
wire u2__abc_52155_new_n19029_; 
wire u2__abc_52155_new_n19031_; 
wire u2__abc_52155_new_n19032_; 
wire u2__abc_52155_new_n19033_; 
wire u2__abc_52155_new_n19034_; 
wire u2__abc_52155_new_n19036_; 
wire u2__abc_52155_new_n19037_; 
wire u2__abc_52155_new_n19038_; 
wire u2__abc_52155_new_n19039_; 
wire u2__abc_52155_new_n19041_; 
wire u2__abc_52155_new_n19042_; 
wire u2__abc_52155_new_n19043_; 
wire u2__abc_52155_new_n19044_; 
wire u2__abc_52155_new_n19046_; 
wire u2__abc_52155_new_n19047_; 
wire u2__abc_52155_new_n19048_; 
wire u2__abc_52155_new_n19049_; 
wire u2__abc_52155_new_n19051_; 
wire u2__abc_52155_new_n19052_; 
wire u2__abc_52155_new_n19053_; 
wire u2__abc_52155_new_n19054_; 
wire u2__abc_52155_new_n19056_; 
wire u2__abc_52155_new_n19057_; 
wire u2__abc_52155_new_n19058_; 
wire u2__abc_52155_new_n19059_; 
wire u2__abc_52155_new_n19061_; 
wire u2__abc_52155_new_n19062_; 
wire u2__abc_52155_new_n19063_; 
wire u2__abc_52155_new_n19064_; 
wire u2__abc_52155_new_n19066_; 
wire u2__abc_52155_new_n19068_; 
wire u2__abc_52155_new_n19069_; 
wire u2__abc_52155_new_n19070_; 
wire u2__abc_52155_new_n19071_; 
wire u2__abc_52155_new_n19072_; 
wire u2__abc_52155_new_n19073_; 
wire u2__abc_52155_new_n19074_; 
wire u2__abc_52155_new_n19075_; 
wire u2__abc_52155_new_n19076_; 
wire u2__abc_52155_new_n19077_; 
wire u2__abc_52155_new_n19078_; 
wire u2__abc_52155_new_n19080_; 
wire u2__abc_52155_new_n19081_; 
wire u2__abc_52155_new_n19082_; 
wire u2__abc_52155_new_n19083_; 
wire u2__abc_52155_new_n19084_; 
wire u2__abc_52155_new_n19085_; 
wire u2__abc_52155_new_n19086_; 
wire u2__abc_52155_new_n19087_; 
wire u2__abc_52155_new_n19088_; 
wire u2__abc_52155_new_n19089_; 
wire u2__abc_52155_new_n19090_; 
wire u2__abc_52155_new_n19092_; 
wire u2__abc_52155_new_n19093_; 
wire u2__abc_52155_new_n19094_; 
wire u2__abc_52155_new_n19095_; 
wire u2__abc_52155_new_n19096_; 
wire u2__abc_52155_new_n19097_; 
wire u2__abc_52155_new_n19098_; 
wire u2__abc_52155_new_n19099_; 
wire u2__abc_52155_new_n19100_; 
wire u2__abc_52155_new_n19101_; 
wire u2__abc_52155_new_n19102_; 
wire u2__abc_52155_new_n19104_; 
wire u2__abc_52155_new_n19105_; 
wire u2__abc_52155_new_n19106_; 
wire u2__abc_52155_new_n19107_; 
wire u2__abc_52155_new_n19108_; 
wire u2__abc_52155_new_n19109_; 
wire u2__abc_52155_new_n19110_; 
wire u2__abc_52155_new_n19111_; 
wire u2__abc_52155_new_n19112_; 
wire u2__abc_52155_new_n19113_; 
wire u2__abc_52155_new_n19114_; 
wire u2__abc_52155_new_n19116_; 
wire u2__abc_52155_new_n19117_; 
wire u2__abc_52155_new_n19118_; 
wire u2__abc_52155_new_n19119_; 
wire u2__abc_52155_new_n19120_; 
wire u2__abc_52155_new_n19121_; 
wire u2__abc_52155_new_n19122_; 
wire u2__abc_52155_new_n19123_; 
wire u2__abc_52155_new_n19124_; 
wire u2__abc_52155_new_n19125_; 
wire u2__abc_52155_new_n19126_; 
wire u2__abc_52155_new_n19128_; 
wire u2__abc_52155_new_n19129_; 
wire u2__abc_52155_new_n19130_; 
wire u2__abc_52155_new_n19131_; 
wire u2__abc_52155_new_n19132_; 
wire u2__abc_52155_new_n19133_; 
wire u2__abc_52155_new_n19134_; 
wire u2__abc_52155_new_n19135_; 
wire u2__abc_52155_new_n19136_; 
wire u2__abc_52155_new_n19137_; 
wire u2__abc_52155_new_n19138_; 
wire u2__abc_52155_new_n19140_; 
wire u2__abc_52155_new_n19141_; 
wire u2__abc_52155_new_n19142_; 
wire u2__abc_52155_new_n19143_; 
wire u2__abc_52155_new_n19144_; 
wire u2__abc_52155_new_n19145_; 
wire u2__abc_52155_new_n19146_; 
wire u2__abc_52155_new_n19147_; 
wire u2__abc_52155_new_n19148_; 
wire u2__abc_52155_new_n19149_; 
wire u2__abc_52155_new_n19150_; 
wire u2__abc_52155_new_n19152_; 
wire u2__abc_52155_new_n19153_; 
wire u2__abc_52155_new_n19154_; 
wire u2__abc_52155_new_n19155_; 
wire u2__abc_52155_new_n19156_; 
wire u2__abc_52155_new_n19157_; 
wire u2__abc_52155_new_n19158_; 
wire u2__abc_52155_new_n19159_; 
wire u2__abc_52155_new_n19160_; 
wire u2__abc_52155_new_n19161_; 
wire u2__abc_52155_new_n19162_; 
wire u2__abc_52155_new_n19164_; 
wire u2__abc_52155_new_n19165_; 
wire u2__abc_52155_new_n19166_; 
wire u2__abc_52155_new_n19167_; 
wire u2__abc_52155_new_n19168_; 
wire u2__abc_52155_new_n19169_; 
wire u2__abc_52155_new_n19170_; 
wire u2__abc_52155_new_n19171_; 
wire u2__abc_52155_new_n19172_; 
wire u2__abc_52155_new_n19173_; 
wire u2__abc_52155_new_n19174_; 
wire u2__abc_52155_new_n19176_; 
wire u2__abc_52155_new_n19177_; 
wire u2__abc_52155_new_n19178_; 
wire u2__abc_52155_new_n19179_; 
wire u2__abc_52155_new_n19180_; 
wire u2__abc_52155_new_n19181_; 
wire u2__abc_52155_new_n19182_; 
wire u2__abc_52155_new_n19183_; 
wire u2__abc_52155_new_n19184_; 
wire u2__abc_52155_new_n19185_; 
wire u2__abc_52155_new_n19186_; 
wire u2__abc_52155_new_n19188_; 
wire u2__abc_52155_new_n19189_; 
wire u2__abc_52155_new_n19190_; 
wire u2__abc_52155_new_n19191_; 
wire u2__abc_52155_new_n19192_; 
wire u2__abc_52155_new_n19193_; 
wire u2__abc_52155_new_n19194_; 
wire u2__abc_52155_new_n19195_; 
wire u2__abc_52155_new_n19196_; 
wire u2__abc_52155_new_n19197_; 
wire u2__abc_52155_new_n19198_; 
wire u2__abc_52155_new_n19200_; 
wire u2__abc_52155_new_n19201_; 
wire u2__abc_52155_new_n19202_; 
wire u2__abc_52155_new_n19203_; 
wire u2__abc_52155_new_n19204_; 
wire u2__abc_52155_new_n19205_; 
wire u2__abc_52155_new_n19206_; 
wire u2__abc_52155_new_n19207_; 
wire u2__abc_52155_new_n19208_; 
wire u2__abc_52155_new_n19209_; 
wire u2__abc_52155_new_n19210_; 
wire u2__abc_52155_new_n19212_; 
wire u2__abc_52155_new_n19213_; 
wire u2__abc_52155_new_n19214_; 
wire u2__abc_52155_new_n19215_; 
wire u2__abc_52155_new_n19216_; 
wire u2__abc_52155_new_n19217_; 
wire u2__abc_52155_new_n19218_; 
wire u2__abc_52155_new_n19219_; 
wire u2__abc_52155_new_n19220_; 
wire u2__abc_52155_new_n19221_; 
wire u2__abc_52155_new_n19222_; 
wire u2__abc_52155_new_n19224_; 
wire u2__abc_52155_new_n19225_; 
wire u2__abc_52155_new_n19226_; 
wire u2__abc_52155_new_n19227_; 
wire u2__abc_52155_new_n19228_; 
wire u2__abc_52155_new_n19229_; 
wire u2__abc_52155_new_n19230_; 
wire u2__abc_52155_new_n19231_; 
wire u2__abc_52155_new_n19232_; 
wire u2__abc_52155_new_n19233_; 
wire u2__abc_52155_new_n19234_; 
wire u2__abc_52155_new_n19236_; 
wire u2__abc_52155_new_n19237_; 
wire u2__abc_52155_new_n19238_; 
wire u2__abc_52155_new_n19239_; 
wire u2__abc_52155_new_n19240_; 
wire u2__abc_52155_new_n19241_; 
wire u2__abc_52155_new_n19242_; 
wire u2__abc_52155_new_n19243_; 
wire u2__abc_52155_new_n19244_; 
wire u2__abc_52155_new_n19245_; 
wire u2__abc_52155_new_n19246_; 
wire u2__abc_52155_new_n19248_; 
wire u2__abc_52155_new_n19249_; 
wire u2__abc_52155_new_n19250_; 
wire u2__abc_52155_new_n19251_; 
wire u2__abc_52155_new_n19252_; 
wire u2__abc_52155_new_n19253_; 
wire u2__abc_52155_new_n19254_; 
wire u2__abc_52155_new_n19255_; 
wire u2__abc_52155_new_n19256_; 
wire u2__abc_52155_new_n19257_; 
wire u2__abc_52155_new_n19258_; 
wire u2__abc_52155_new_n19260_; 
wire u2__abc_52155_new_n19261_; 
wire u2__abc_52155_new_n19262_; 
wire u2__abc_52155_new_n19263_; 
wire u2__abc_52155_new_n19264_; 
wire u2__abc_52155_new_n19265_; 
wire u2__abc_52155_new_n19266_; 
wire u2__abc_52155_new_n19267_; 
wire u2__abc_52155_new_n19268_; 
wire u2__abc_52155_new_n19269_; 
wire u2__abc_52155_new_n19270_; 
wire u2__abc_52155_new_n19272_; 
wire u2__abc_52155_new_n19273_; 
wire u2__abc_52155_new_n19274_; 
wire u2__abc_52155_new_n19275_; 
wire u2__abc_52155_new_n19276_; 
wire u2__abc_52155_new_n19277_; 
wire u2__abc_52155_new_n19278_; 
wire u2__abc_52155_new_n19279_; 
wire u2__abc_52155_new_n19280_; 
wire u2__abc_52155_new_n19281_; 
wire u2__abc_52155_new_n19282_; 
wire u2__abc_52155_new_n19284_; 
wire u2__abc_52155_new_n19285_; 
wire u2__abc_52155_new_n19286_; 
wire u2__abc_52155_new_n19287_; 
wire u2__abc_52155_new_n19288_; 
wire u2__abc_52155_new_n19289_; 
wire u2__abc_52155_new_n19290_; 
wire u2__abc_52155_new_n19291_; 
wire u2__abc_52155_new_n19292_; 
wire u2__abc_52155_new_n19293_; 
wire u2__abc_52155_new_n19294_; 
wire u2__abc_52155_new_n19296_; 
wire u2__abc_52155_new_n19297_; 
wire u2__abc_52155_new_n19298_; 
wire u2__abc_52155_new_n19299_; 
wire u2__abc_52155_new_n19300_; 
wire u2__abc_52155_new_n19301_; 
wire u2__abc_52155_new_n19302_; 
wire u2__abc_52155_new_n19303_; 
wire u2__abc_52155_new_n19304_; 
wire u2__abc_52155_new_n19305_; 
wire u2__abc_52155_new_n19306_; 
wire u2__abc_52155_new_n19308_; 
wire u2__abc_52155_new_n19309_; 
wire u2__abc_52155_new_n19310_; 
wire u2__abc_52155_new_n19311_; 
wire u2__abc_52155_new_n19312_; 
wire u2__abc_52155_new_n19313_; 
wire u2__abc_52155_new_n19314_; 
wire u2__abc_52155_new_n19315_; 
wire u2__abc_52155_new_n19316_; 
wire u2__abc_52155_new_n19317_; 
wire u2__abc_52155_new_n19318_; 
wire u2__abc_52155_new_n19320_; 
wire u2__abc_52155_new_n19321_; 
wire u2__abc_52155_new_n19322_; 
wire u2__abc_52155_new_n19323_; 
wire u2__abc_52155_new_n19324_; 
wire u2__abc_52155_new_n19325_; 
wire u2__abc_52155_new_n19326_; 
wire u2__abc_52155_new_n19327_; 
wire u2__abc_52155_new_n19328_; 
wire u2__abc_52155_new_n19329_; 
wire u2__abc_52155_new_n19330_; 
wire u2__abc_52155_new_n19332_; 
wire u2__abc_52155_new_n19333_; 
wire u2__abc_52155_new_n19334_; 
wire u2__abc_52155_new_n19335_; 
wire u2__abc_52155_new_n19336_; 
wire u2__abc_52155_new_n19337_; 
wire u2__abc_52155_new_n19338_; 
wire u2__abc_52155_new_n19339_; 
wire u2__abc_52155_new_n19340_; 
wire u2__abc_52155_new_n19341_; 
wire u2__abc_52155_new_n19342_; 
wire u2__abc_52155_new_n19344_; 
wire u2__abc_52155_new_n19345_; 
wire u2__abc_52155_new_n19346_; 
wire u2__abc_52155_new_n19347_; 
wire u2__abc_52155_new_n19348_; 
wire u2__abc_52155_new_n19349_; 
wire u2__abc_52155_new_n19350_; 
wire u2__abc_52155_new_n19351_; 
wire u2__abc_52155_new_n19352_; 
wire u2__abc_52155_new_n19353_; 
wire u2__abc_52155_new_n19354_; 
wire u2__abc_52155_new_n19356_; 
wire u2__abc_52155_new_n19357_; 
wire u2__abc_52155_new_n19358_; 
wire u2__abc_52155_new_n19359_; 
wire u2__abc_52155_new_n19360_; 
wire u2__abc_52155_new_n19361_; 
wire u2__abc_52155_new_n19362_; 
wire u2__abc_52155_new_n19363_; 
wire u2__abc_52155_new_n19364_; 
wire u2__abc_52155_new_n19365_; 
wire u2__abc_52155_new_n19366_; 
wire u2__abc_52155_new_n19368_; 
wire u2__abc_52155_new_n19369_; 
wire u2__abc_52155_new_n19370_; 
wire u2__abc_52155_new_n19371_; 
wire u2__abc_52155_new_n19372_; 
wire u2__abc_52155_new_n19373_; 
wire u2__abc_52155_new_n19374_; 
wire u2__abc_52155_new_n19375_; 
wire u2__abc_52155_new_n19376_; 
wire u2__abc_52155_new_n19377_; 
wire u2__abc_52155_new_n19378_; 
wire u2__abc_52155_new_n19380_; 
wire u2__abc_52155_new_n19381_; 
wire u2__abc_52155_new_n19382_; 
wire u2__abc_52155_new_n19383_; 
wire u2__abc_52155_new_n19384_; 
wire u2__abc_52155_new_n19385_; 
wire u2__abc_52155_new_n19386_; 
wire u2__abc_52155_new_n19387_; 
wire u2__abc_52155_new_n19388_; 
wire u2__abc_52155_new_n19389_; 
wire u2__abc_52155_new_n19390_; 
wire u2__abc_52155_new_n19392_; 
wire u2__abc_52155_new_n19393_; 
wire u2__abc_52155_new_n19394_; 
wire u2__abc_52155_new_n19395_; 
wire u2__abc_52155_new_n19396_; 
wire u2__abc_52155_new_n19397_; 
wire u2__abc_52155_new_n19398_; 
wire u2__abc_52155_new_n19399_; 
wire u2__abc_52155_new_n19400_; 
wire u2__abc_52155_new_n19401_; 
wire u2__abc_52155_new_n19402_; 
wire u2__abc_52155_new_n19404_; 
wire u2__abc_52155_new_n19405_; 
wire u2__abc_52155_new_n19406_; 
wire u2__abc_52155_new_n19407_; 
wire u2__abc_52155_new_n19408_; 
wire u2__abc_52155_new_n19409_; 
wire u2__abc_52155_new_n19410_; 
wire u2__abc_52155_new_n19411_; 
wire u2__abc_52155_new_n19412_; 
wire u2__abc_52155_new_n19413_; 
wire u2__abc_52155_new_n19414_; 
wire u2__abc_52155_new_n19416_; 
wire u2__abc_52155_new_n19417_; 
wire u2__abc_52155_new_n19418_; 
wire u2__abc_52155_new_n19419_; 
wire u2__abc_52155_new_n19420_; 
wire u2__abc_52155_new_n19421_; 
wire u2__abc_52155_new_n19422_; 
wire u2__abc_52155_new_n19423_; 
wire u2__abc_52155_new_n19424_; 
wire u2__abc_52155_new_n19425_; 
wire u2__abc_52155_new_n19426_; 
wire u2__abc_52155_new_n19428_; 
wire u2__abc_52155_new_n19429_; 
wire u2__abc_52155_new_n19430_; 
wire u2__abc_52155_new_n19431_; 
wire u2__abc_52155_new_n19432_; 
wire u2__abc_52155_new_n19433_; 
wire u2__abc_52155_new_n19434_; 
wire u2__abc_52155_new_n19435_; 
wire u2__abc_52155_new_n19436_; 
wire u2__abc_52155_new_n19437_; 
wire u2__abc_52155_new_n19438_; 
wire u2__abc_52155_new_n19440_; 
wire u2__abc_52155_new_n19441_; 
wire u2__abc_52155_new_n19442_; 
wire u2__abc_52155_new_n19443_; 
wire u2__abc_52155_new_n19444_; 
wire u2__abc_52155_new_n19445_; 
wire u2__abc_52155_new_n19446_; 
wire u2__abc_52155_new_n19447_; 
wire u2__abc_52155_new_n19448_; 
wire u2__abc_52155_new_n19449_; 
wire u2__abc_52155_new_n19450_; 
wire u2__abc_52155_new_n19452_; 
wire u2__abc_52155_new_n19453_; 
wire u2__abc_52155_new_n19454_; 
wire u2__abc_52155_new_n19455_; 
wire u2__abc_52155_new_n19456_; 
wire u2__abc_52155_new_n19457_; 
wire u2__abc_52155_new_n19458_; 
wire u2__abc_52155_new_n19459_; 
wire u2__abc_52155_new_n19460_; 
wire u2__abc_52155_new_n19461_; 
wire u2__abc_52155_new_n19462_; 
wire u2__abc_52155_new_n19464_; 
wire u2__abc_52155_new_n19465_; 
wire u2__abc_52155_new_n19466_; 
wire u2__abc_52155_new_n19467_; 
wire u2__abc_52155_new_n19468_; 
wire u2__abc_52155_new_n19469_; 
wire u2__abc_52155_new_n19470_; 
wire u2__abc_52155_new_n19471_; 
wire u2__abc_52155_new_n19472_; 
wire u2__abc_52155_new_n19473_; 
wire u2__abc_52155_new_n19474_; 
wire u2__abc_52155_new_n19476_; 
wire u2__abc_52155_new_n19477_; 
wire u2__abc_52155_new_n19478_; 
wire u2__abc_52155_new_n19479_; 
wire u2__abc_52155_new_n19480_; 
wire u2__abc_52155_new_n19481_; 
wire u2__abc_52155_new_n19482_; 
wire u2__abc_52155_new_n19483_; 
wire u2__abc_52155_new_n19484_; 
wire u2__abc_52155_new_n19485_; 
wire u2__abc_52155_new_n19486_; 
wire u2__abc_52155_new_n19488_; 
wire u2__abc_52155_new_n19489_; 
wire u2__abc_52155_new_n19490_; 
wire u2__abc_52155_new_n19491_; 
wire u2__abc_52155_new_n19492_; 
wire u2__abc_52155_new_n19493_; 
wire u2__abc_52155_new_n19494_; 
wire u2__abc_52155_new_n19495_; 
wire u2__abc_52155_new_n19496_; 
wire u2__abc_52155_new_n19497_; 
wire u2__abc_52155_new_n19498_; 
wire u2__abc_52155_new_n19500_; 
wire u2__abc_52155_new_n19501_; 
wire u2__abc_52155_new_n19502_; 
wire u2__abc_52155_new_n19503_; 
wire u2__abc_52155_new_n19504_; 
wire u2__abc_52155_new_n19505_; 
wire u2__abc_52155_new_n19506_; 
wire u2__abc_52155_new_n19507_; 
wire u2__abc_52155_new_n19508_; 
wire u2__abc_52155_new_n19509_; 
wire u2__abc_52155_new_n19510_; 
wire u2__abc_52155_new_n19512_; 
wire u2__abc_52155_new_n19513_; 
wire u2__abc_52155_new_n19514_; 
wire u2__abc_52155_new_n19515_; 
wire u2__abc_52155_new_n19516_; 
wire u2__abc_52155_new_n19517_; 
wire u2__abc_52155_new_n19518_; 
wire u2__abc_52155_new_n19519_; 
wire u2__abc_52155_new_n19520_; 
wire u2__abc_52155_new_n19521_; 
wire u2__abc_52155_new_n19522_; 
wire u2__abc_52155_new_n19524_; 
wire u2__abc_52155_new_n19525_; 
wire u2__abc_52155_new_n19526_; 
wire u2__abc_52155_new_n19527_; 
wire u2__abc_52155_new_n19528_; 
wire u2__abc_52155_new_n19529_; 
wire u2__abc_52155_new_n19530_; 
wire u2__abc_52155_new_n19531_; 
wire u2__abc_52155_new_n19532_; 
wire u2__abc_52155_new_n19533_; 
wire u2__abc_52155_new_n19534_; 
wire u2__abc_52155_new_n19536_; 
wire u2__abc_52155_new_n19537_; 
wire u2__abc_52155_new_n19538_; 
wire u2__abc_52155_new_n19539_; 
wire u2__abc_52155_new_n19540_; 
wire u2__abc_52155_new_n19541_; 
wire u2__abc_52155_new_n19542_; 
wire u2__abc_52155_new_n19543_; 
wire u2__abc_52155_new_n19544_; 
wire u2__abc_52155_new_n19545_; 
wire u2__abc_52155_new_n19546_; 
wire u2__abc_52155_new_n19548_; 
wire u2__abc_52155_new_n19549_; 
wire u2__abc_52155_new_n19550_; 
wire u2__abc_52155_new_n19551_; 
wire u2__abc_52155_new_n19552_; 
wire u2__abc_52155_new_n19553_; 
wire u2__abc_52155_new_n19554_; 
wire u2__abc_52155_new_n19555_; 
wire u2__abc_52155_new_n19556_; 
wire u2__abc_52155_new_n19557_; 
wire u2__abc_52155_new_n19558_; 
wire u2__abc_52155_new_n19560_; 
wire u2__abc_52155_new_n19561_; 
wire u2__abc_52155_new_n19562_; 
wire u2__abc_52155_new_n19563_; 
wire u2__abc_52155_new_n19564_; 
wire u2__abc_52155_new_n19565_; 
wire u2__abc_52155_new_n19566_; 
wire u2__abc_52155_new_n19567_; 
wire u2__abc_52155_new_n19568_; 
wire u2__abc_52155_new_n19569_; 
wire u2__abc_52155_new_n19570_; 
wire u2__abc_52155_new_n19572_; 
wire u2__abc_52155_new_n19573_; 
wire u2__abc_52155_new_n19574_; 
wire u2__abc_52155_new_n19575_; 
wire u2__abc_52155_new_n19576_; 
wire u2__abc_52155_new_n19577_; 
wire u2__abc_52155_new_n19578_; 
wire u2__abc_52155_new_n19579_; 
wire u2__abc_52155_new_n19580_; 
wire u2__abc_52155_new_n19581_; 
wire u2__abc_52155_new_n19582_; 
wire u2__abc_52155_new_n19584_; 
wire u2__abc_52155_new_n19585_; 
wire u2__abc_52155_new_n19586_; 
wire u2__abc_52155_new_n19587_; 
wire u2__abc_52155_new_n19588_; 
wire u2__abc_52155_new_n19589_; 
wire u2__abc_52155_new_n19590_; 
wire u2__abc_52155_new_n19591_; 
wire u2__abc_52155_new_n19592_; 
wire u2__abc_52155_new_n19593_; 
wire u2__abc_52155_new_n19594_; 
wire u2__abc_52155_new_n19596_; 
wire u2__abc_52155_new_n19597_; 
wire u2__abc_52155_new_n19598_; 
wire u2__abc_52155_new_n19599_; 
wire u2__abc_52155_new_n19600_; 
wire u2__abc_52155_new_n19601_; 
wire u2__abc_52155_new_n19602_; 
wire u2__abc_52155_new_n19603_; 
wire u2__abc_52155_new_n19604_; 
wire u2__abc_52155_new_n19605_; 
wire u2__abc_52155_new_n19606_; 
wire u2__abc_52155_new_n19608_; 
wire u2__abc_52155_new_n19609_; 
wire u2__abc_52155_new_n19610_; 
wire u2__abc_52155_new_n19611_; 
wire u2__abc_52155_new_n19612_; 
wire u2__abc_52155_new_n19613_; 
wire u2__abc_52155_new_n19614_; 
wire u2__abc_52155_new_n19615_; 
wire u2__abc_52155_new_n19616_; 
wire u2__abc_52155_new_n19617_; 
wire u2__abc_52155_new_n19618_; 
wire u2__abc_52155_new_n19620_; 
wire u2__abc_52155_new_n19621_; 
wire u2__abc_52155_new_n19622_; 
wire u2__abc_52155_new_n19623_; 
wire u2__abc_52155_new_n19624_; 
wire u2__abc_52155_new_n19625_; 
wire u2__abc_52155_new_n19626_; 
wire u2__abc_52155_new_n19627_; 
wire u2__abc_52155_new_n19628_; 
wire u2__abc_52155_new_n19629_; 
wire u2__abc_52155_new_n19630_; 
wire u2__abc_52155_new_n19632_; 
wire u2__abc_52155_new_n19633_; 
wire u2__abc_52155_new_n19634_; 
wire u2__abc_52155_new_n19635_; 
wire u2__abc_52155_new_n19636_; 
wire u2__abc_52155_new_n19637_; 
wire u2__abc_52155_new_n19638_; 
wire u2__abc_52155_new_n19639_; 
wire u2__abc_52155_new_n19640_; 
wire u2__abc_52155_new_n19641_; 
wire u2__abc_52155_new_n19642_; 
wire u2__abc_52155_new_n19644_; 
wire u2__abc_52155_new_n19645_; 
wire u2__abc_52155_new_n19646_; 
wire u2__abc_52155_new_n19647_; 
wire u2__abc_52155_new_n19648_; 
wire u2__abc_52155_new_n19649_; 
wire u2__abc_52155_new_n19650_; 
wire u2__abc_52155_new_n19651_; 
wire u2__abc_52155_new_n19652_; 
wire u2__abc_52155_new_n19653_; 
wire u2__abc_52155_new_n19654_; 
wire u2__abc_52155_new_n19656_; 
wire u2__abc_52155_new_n19657_; 
wire u2__abc_52155_new_n19658_; 
wire u2__abc_52155_new_n19659_; 
wire u2__abc_52155_new_n19660_; 
wire u2__abc_52155_new_n19661_; 
wire u2__abc_52155_new_n19662_; 
wire u2__abc_52155_new_n19663_; 
wire u2__abc_52155_new_n19664_; 
wire u2__abc_52155_new_n19665_; 
wire u2__abc_52155_new_n19666_; 
wire u2__abc_52155_new_n19668_; 
wire u2__abc_52155_new_n19669_; 
wire u2__abc_52155_new_n19670_; 
wire u2__abc_52155_new_n19671_; 
wire u2__abc_52155_new_n19672_; 
wire u2__abc_52155_new_n19673_; 
wire u2__abc_52155_new_n19674_; 
wire u2__abc_52155_new_n19675_; 
wire u2__abc_52155_new_n19676_; 
wire u2__abc_52155_new_n19677_; 
wire u2__abc_52155_new_n19678_; 
wire u2__abc_52155_new_n19680_; 
wire u2__abc_52155_new_n19681_; 
wire u2__abc_52155_new_n19682_; 
wire u2__abc_52155_new_n19683_; 
wire u2__abc_52155_new_n19684_; 
wire u2__abc_52155_new_n19685_; 
wire u2__abc_52155_new_n19686_; 
wire u2__abc_52155_new_n19687_; 
wire u2__abc_52155_new_n19688_; 
wire u2__abc_52155_new_n19689_; 
wire u2__abc_52155_new_n19690_; 
wire u2__abc_52155_new_n19692_; 
wire u2__abc_52155_new_n19693_; 
wire u2__abc_52155_new_n19694_; 
wire u2__abc_52155_new_n19695_; 
wire u2__abc_52155_new_n19696_; 
wire u2__abc_52155_new_n19697_; 
wire u2__abc_52155_new_n19698_; 
wire u2__abc_52155_new_n19699_; 
wire u2__abc_52155_new_n19700_; 
wire u2__abc_52155_new_n19701_; 
wire u2__abc_52155_new_n19702_; 
wire u2__abc_52155_new_n19704_; 
wire u2__abc_52155_new_n19705_; 
wire u2__abc_52155_new_n19706_; 
wire u2__abc_52155_new_n19707_; 
wire u2__abc_52155_new_n19708_; 
wire u2__abc_52155_new_n19709_; 
wire u2__abc_52155_new_n19710_; 
wire u2__abc_52155_new_n19711_; 
wire u2__abc_52155_new_n19712_; 
wire u2__abc_52155_new_n19713_; 
wire u2__abc_52155_new_n19714_; 
wire u2__abc_52155_new_n19716_; 
wire u2__abc_52155_new_n19717_; 
wire u2__abc_52155_new_n19718_; 
wire u2__abc_52155_new_n19719_; 
wire u2__abc_52155_new_n19720_; 
wire u2__abc_52155_new_n19721_; 
wire u2__abc_52155_new_n19722_; 
wire u2__abc_52155_new_n19723_; 
wire u2__abc_52155_new_n19724_; 
wire u2__abc_52155_new_n19725_; 
wire u2__abc_52155_new_n19726_; 
wire u2__abc_52155_new_n19728_; 
wire u2__abc_52155_new_n19729_; 
wire u2__abc_52155_new_n19730_; 
wire u2__abc_52155_new_n19731_; 
wire u2__abc_52155_new_n19732_; 
wire u2__abc_52155_new_n19733_; 
wire u2__abc_52155_new_n19734_; 
wire u2__abc_52155_new_n19735_; 
wire u2__abc_52155_new_n19736_; 
wire u2__abc_52155_new_n19737_; 
wire u2__abc_52155_new_n19738_; 
wire u2__abc_52155_new_n19740_; 
wire u2__abc_52155_new_n19741_; 
wire u2__abc_52155_new_n19742_; 
wire u2__abc_52155_new_n19743_; 
wire u2__abc_52155_new_n19744_; 
wire u2__abc_52155_new_n19745_; 
wire u2__abc_52155_new_n19746_; 
wire u2__abc_52155_new_n19747_; 
wire u2__abc_52155_new_n19748_; 
wire u2__abc_52155_new_n19749_; 
wire u2__abc_52155_new_n19750_; 
wire u2__abc_52155_new_n19752_; 
wire u2__abc_52155_new_n19753_; 
wire u2__abc_52155_new_n19754_; 
wire u2__abc_52155_new_n19755_; 
wire u2__abc_52155_new_n19756_; 
wire u2__abc_52155_new_n19757_; 
wire u2__abc_52155_new_n19758_; 
wire u2__abc_52155_new_n19759_; 
wire u2__abc_52155_new_n19760_; 
wire u2__abc_52155_new_n19761_; 
wire u2__abc_52155_new_n19762_; 
wire u2__abc_52155_new_n19764_; 
wire u2__abc_52155_new_n19765_; 
wire u2__abc_52155_new_n19766_; 
wire u2__abc_52155_new_n19767_; 
wire u2__abc_52155_new_n19768_; 
wire u2__abc_52155_new_n19769_; 
wire u2__abc_52155_new_n19770_; 
wire u2__abc_52155_new_n19771_; 
wire u2__abc_52155_new_n19772_; 
wire u2__abc_52155_new_n19773_; 
wire u2__abc_52155_new_n19774_; 
wire u2__abc_52155_new_n19776_; 
wire u2__abc_52155_new_n19777_; 
wire u2__abc_52155_new_n19778_; 
wire u2__abc_52155_new_n19779_; 
wire u2__abc_52155_new_n19780_; 
wire u2__abc_52155_new_n19781_; 
wire u2__abc_52155_new_n19782_; 
wire u2__abc_52155_new_n19783_; 
wire u2__abc_52155_new_n19784_; 
wire u2__abc_52155_new_n19785_; 
wire u2__abc_52155_new_n19786_; 
wire u2__abc_52155_new_n19788_; 
wire u2__abc_52155_new_n19789_; 
wire u2__abc_52155_new_n19790_; 
wire u2__abc_52155_new_n19791_; 
wire u2__abc_52155_new_n19792_; 
wire u2__abc_52155_new_n19793_; 
wire u2__abc_52155_new_n19794_; 
wire u2__abc_52155_new_n19795_; 
wire u2__abc_52155_new_n19796_; 
wire u2__abc_52155_new_n19797_; 
wire u2__abc_52155_new_n19798_; 
wire u2__abc_52155_new_n19800_; 
wire u2__abc_52155_new_n19801_; 
wire u2__abc_52155_new_n19802_; 
wire u2__abc_52155_new_n19803_; 
wire u2__abc_52155_new_n19804_; 
wire u2__abc_52155_new_n19805_; 
wire u2__abc_52155_new_n19806_; 
wire u2__abc_52155_new_n19807_; 
wire u2__abc_52155_new_n19808_; 
wire u2__abc_52155_new_n19809_; 
wire u2__abc_52155_new_n19810_; 
wire u2__abc_52155_new_n19812_; 
wire u2__abc_52155_new_n19813_; 
wire u2__abc_52155_new_n19814_; 
wire u2__abc_52155_new_n19815_; 
wire u2__abc_52155_new_n19816_; 
wire u2__abc_52155_new_n19817_; 
wire u2__abc_52155_new_n19818_; 
wire u2__abc_52155_new_n19819_; 
wire u2__abc_52155_new_n19820_; 
wire u2__abc_52155_new_n19821_; 
wire u2__abc_52155_new_n19822_; 
wire u2__abc_52155_new_n19824_; 
wire u2__abc_52155_new_n19825_; 
wire u2__abc_52155_new_n19826_; 
wire u2__abc_52155_new_n19827_; 
wire u2__abc_52155_new_n19828_; 
wire u2__abc_52155_new_n19829_; 
wire u2__abc_52155_new_n19830_; 
wire u2__abc_52155_new_n19831_; 
wire u2__abc_52155_new_n19832_; 
wire u2__abc_52155_new_n19833_; 
wire u2__abc_52155_new_n19834_; 
wire u2__abc_52155_new_n19836_; 
wire u2__abc_52155_new_n19837_; 
wire u2__abc_52155_new_n19838_; 
wire u2__abc_52155_new_n19839_; 
wire u2__abc_52155_new_n19840_; 
wire u2__abc_52155_new_n19841_; 
wire u2__abc_52155_new_n19842_; 
wire u2__abc_52155_new_n19843_; 
wire u2__abc_52155_new_n19844_; 
wire u2__abc_52155_new_n19845_; 
wire u2__abc_52155_new_n19846_; 
wire u2__abc_52155_new_n19848_; 
wire u2__abc_52155_new_n19849_; 
wire u2__abc_52155_new_n19850_; 
wire u2__abc_52155_new_n19851_; 
wire u2__abc_52155_new_n19852_; 
wire u2__abc_52155_new_n19853_; 
wire u2__abc_52155_new_n19854_; 
wire u2__abc_52155_new_n19855_; 
wire u2__abc_52155_new_n19856_; 
wire u2__abc_52155_new_n19857_; 
wire u2__abc_52155_new_n19858_; 
wire u2__abc_52155_new_n19860_; 
wire u2__abc_52155_new_n19861_; 
wire u2__abc_52155_new_n19862_; 
wire u2__abc_52155_new_n19863_; 
wire u2__abc_52155_new_n19864_; 
wire u2__abc_52155_new_n19865_; 
wire u2__abc_52155_new_n19866_; 
wire u2__abc_52155_new_n19867_; 
wire u2__abc_52155_new_n19868_; 
wire u2__abc_52155_new_n19869_; 
wire u2__abc_52155_new_n19870_; 
wire u2__abc_52155_new_n19872_; 
wire u2__abc_52155_new_n19873_; 
wire u2__abc_52155_new_n19874_; 
wire u2__abc_52155_new_n19875_; 
wire u2__abc_52155_new_n19876_; 
wire u2__abc_52155_new_n19877_; 
wire u2__abc_52155_new_n19878_; 
wire u2__abc_52155_new_n19879_; 
wire u2__abc_52155_new_n19880_; 
wire u2__abc_52155_new_n19881_; 
wire u2__abc_52155_new_n19882_; 
wire u2__abc_52155_new_n19884_; 
wire u2__abc_52155_new_n19885_; 
wire u2__abc_52155_new_n19886_; 
wire u2__abc_52155_new_n19887_; 
wire u2__abc_52155_new_n19888_; 
wire u2__abc_52155_new_n19889_; 
wire u2__abc_52155_new_n19890_; 
wire u2__abc_52155_new_n19891_; 
wire u2__abc_52155_new_n19892_; 
wire u2__abc_52155_new_n19893_; 
wire u2__abc_52155_new_n19894_; 
wire u2__abc_52155_new_n19896_; 
wire u2__abc_52155_new_n19897_; 
wire u2__abc_52155_new_n19898_; 
wire u2__abc_52155_new_n19899_; 
wire u2__abc_52155_new_n19900_; 
wire u2__abc_52155_new_n19901_; 
wire u2__abc_52155_new_n19902_; 
wire u2__abc_52155_new_n19903_; 
wire u2__abc_52155_new_n19904_; 
wire u2__abc_52155_new_n19905_; 
wire u2__abc_52155_new_n19906_; 
wire u2__abc_52155_new_n19908_; 
wire u2__abc_52155_new_n19909_; 
wire u2__abc_52155_new_n19910_; 
wire u2__abc_52155_new_n19911_; 
wire u2__abc_52155_new_n19912_; 
wire u2__abc_52155_new_n19913_; 
wire u2__abc_52155_new_n19914_; 
wire u2__abc_52155_new_n19915_; 
wire u2__abc_52155_new_n19916_; 
wire u2__abc_52155_new_n19917_; 
wire u2__abc_52155_new_n19918_; 
wire u2__abc_52155_new_n19920_; 
wire u2__abc_52155_new_n19921_; 
wire u2__abc_52155_new_n19922_; 
wire u2__abc_52155_new_n19923_; 
wire u2__abc_52155_new_n19924_; 
wire u2__abc_52155_new_n19925_; 
wire u2__abc_52155_new_n19926_; 
wire u2__abc_52155_new_n19927_; 
wire u2__abc_52155_new_n19928_; 
wire u2__abc_52155_new_n19929_; 
wire u2__abc_52155_new_n19930_; 
wire u2__abc_52155_new_n19932_; 
wire u2__abc_52155_new_n19933_; 
wire u2__abc_52155_new_n19934_; 
wire u2__abc_52155_new_n19935_; 
wire u2__abc_52155_new_n19936_; 
wire u2__abc_52155_new_n19937_; 
wire u2__abc_52155_new_n19938_; 
wire u2__abc_52155_new_n19939_; 
wire u2__abc_52155_new_n19940_; 
wire u2__abc_52155_new_n19941_; 
wire u2__abc_52155_new_n19942_; 
wire u2__abc_52155_new_n19944_; 
wire u2__abc_52155_new_n19945_; 
wire u2__abc_52155_new_n19946_; 
wire u2__abc_52155_new_n19947_; 
wire u2__abc_52155_new_n19948_; 
wire u2__abc_52155_new_n19949_; 
wire u2__abc_52155_new_n19950_; 
wire u2__abc_52155_new_n19951_; 
wire u2__abc_52155_new_n19952_; 
wire u2__abc_52155_new_n19953_; 
wire u2__abc_52155_new_n19954_; 
wire u2__abc_52155_new_n19956_; 
wire u2__abc_52155_new_n19957_; 
wire u2__abc_52155_new_n19958_; 
wire u2__abc_52155_new_n19959_; 
wire u2__abc_52155_new_n19960_; 
wire u2__abc_52155_new_n19961_; 
wire u2__abc_52155_new_n19962_; 
wire u2__abc_52155_new_n19963_; 
wire u2__abc_52155_new_n19964_; 
wire u2__abc_52155_new_n19965_; 
wire u2__abc_52155_new_n19966_; 
wire u2__abc_52155_new_n19968_; 
wire u2__abc_52155_new_n19969_; 
wire u2__abc_52155_new_n19970_; 
wire u2__abc_52155_new_n19971_; 
wire u2__abc_52155_new_n19972_; 
wire u2__abc_52155_new_n19973_; 
wire u2__abc_52155_new_n19974_; 
wire u2__abc_52155_new_n19975_; 
wire u2__abc_52155_new_n19976_; 
wire u2__abc_52155_new_n19977_; 
wire u2__abc_52155_new_n19978_; 
wire u2__abc_52155_new_n19980_; 
wire u2__abc_52155_new_n19981_; 
wire u2__abc_52155_new_n19982_; 
wire u2__abc_52155_new_n19983_; 
wire u2__abc_52155_new_n19984_; 
wire u2__abc_52155_new_n19985_; 
wire u2__abc_52155_new_n19986_; 
wire u2__abc_52155_new_n19987_; 
wire u2__abc_52155_new_n19988_; 
wire u2__abc_52155_new_n19989_; 
wire u2__abc_52155_new_n19990_; 
wire u2__abc_52155_new_n19992_; 
wire u2__abc_52155_new_n19993_; 
wire u2__abc_52155_new_n19994_; 
wire u2__abc_52155_new_n19995_; 
wire u2__abc_52155_new_n19996_; 
wire u2__abc_52155_new_n19997_; 
wire u2__abc_52155_new_n19998_; 
wire u2__abc_52155_new_n19999_; 
wire u2__abc_52155_new_n20000_; 
wire u2__abc_52155_new_n20001_; 
wire u2__abc_52155_new_n20002_; 
wire u2__abc_52155_new_n20004_; 
wire u2__abc_52155_new_n20005_; 
wire u2__abc_52155_new_n20006_; 
wire u2__abc_52155_new_n20007_; 
wire u2__abc_52155_new_n20008_; 
wire u2__abc_52155_new_n20009_; 
wire u2__abc_52155_new_n20010_; 
wire u2__abc_52155_new_n20011_; 
wire u2__abc_52155_new_n20012_; 
wire u2__abc_52155_new_n20013_; 
wire u2__abc_52155_new_n20014_; 
wire u2__abc_52155_new_n20016_; 
wire u2__abc_52155_new_n20017_; 
wire u2__abc_52155_new_n20018_; 
wire u2__abc_52155_new_n20019_; 
wire u2__abc_52155_new_n20020_; 
wire u2__abc_52155_new_n20021_; 
wire u2__abc_52155_new_n20022_; 
wire u2__abc_52155_new_n20023_; 
wire u2__abc_52155_new_n20024_; 
wire u2__abc_52155_new_n20025_; 
wire u2__abc_52155_new_n20026_; 
wire u2__abc_52155_new_n20028_; 
wire u2__abc_52155_new_n20029_; 
wire u2__abc_52155_new_n20030_; 
wire u2__abc_52155_new_n20031_; 
wire u2__abc_52155_new_n20032_; 
wire u2__abc_52155_new_n20033_; 
wire u2__abc_52155_new_n20034_; 
wire u2__abc_52155_new_n20035_; 
wire u2__abc_52155_new_n20036_; 
wire u2__abc_52155_new_n20037_; 
wire u2__abc_52155_new_n20038_; 
wire u2__abc_52155_new_n20040_; 
wire u2__abc_52155_new_n20041_; 
wire u2__abc_52155_new_n20042_; 
wire u2__abc_52155_new_n20043_; 
wire u2__abc_52155_new_n20044_; 
wire u2__abc_52155_new_n20045_; 
wire u2__abc_52155_new_n20046_; 
wire u2__abc_52155_new_n20047_; 
wire u2__abc_52155_new_n20048_; 
wire u2__abc_52155_new_n20049_; 
wire u2__abc_52155_new_n20050_; 
wire u2__abc_52155_new_n20052_; 
wire u2__abc_52155_new_n20053_; 
wire u2__abc_52155_new_n20054_; 
wire u2__abc_52155_new_n20055_; 
wire u2__abc_52155_new_n20056_; 
wire u2__abc_52155_new_n20057_; 
wire u2__abc_52155_new_n20058_; 
wire u2__abc_52155_new_n20059_; 
wire u2__abc_52155_new_n20060_; 
wire u2__abc_52155_new_n20061_; 
wire u2__abc_52155_new_n20062_; 
wire u2__abc_52155_new_n20064_; 
wire u2__abc_52155_new_n20065_; 
wire u2__abc_52155_new_n20066_; 
wire u2__abc_52155_new_n20067_; 
wire u2__abc_52155_new_n20068_; 
wire u2__abc_52155_new_n20069_; 
wire u2__abc_52155_new_n20070_; 
wire u2__abc_52155_new_n20071_; 
wire u2__abc_52155_new_n20072_; 
wire u2__abc_52155_new_n20073_; 
wire u2__abc_52155_new_n20074_; 
wire u2__abc_52155_new_n20076_; 
wire u2__abc_52155_new_n20077_; 
wire u2__abc_52155_new_n20078_; 
wire u2__abc_52155_new_n20079_; 
wire u2__abc_52155_new_n20080_; 
wire u2__abc_52155_new_n20081_; 
wire u2__abc_52155_new_n20082_; 
wire u2__abc_52155_new_n20083_; 
wire u2__abc_52155_new_n20084_; 
wire u2__abc_52155_new_n20085_; 
wire u2__abc_52155_new_n20086_; 
wire u2__abc_52155_new_n20088_; 
wire u2__abc_52155_new_n20089_; 
wire u2__abc_52155_new_n20090_; 
wire u2__abc_52155_new_n20091_; 
wire u2__abc_52155_new_n20092_; 
wire u2__abc_52155_new_n20093_; 
wire u2__abc_52155_new_n20094_; 
wire u2__abc_52155_new_n20095_; 
wire u2__abc_52155_new_n20096_; 
wire u2__abc_52155_new_n20097_; 
wire u2__abc_52155_new_n20098_; 
wire u2__abc_52155_new_n20100_; 
wire u2__abc_52155_new_n20101_; 
wire u2__abc_52155_new_n20102_; 
wire u2__abc_52155_new_n20103_; 
wire u2__abc_52155_new_n20104_; 
wire u2__abc_52155_new_n20105_; 
wire u2__abc_52155_new_n20106_; 
wire u2__abc_52155_new_n20107_; 
wire u2__abc_52155_new_n20108_; 
wire u2__abc_52155_new_n20109_; 
wire u2__abc_52155_new_n20110_; 
wire u2__abc_52155_new_n20112_; 
wire u2__abc_52155_new_n20113_; 
wire u2__abc_52155_new_n20114_; 
wire u2__abc_52155_new_n20115_; 
wire u2__abc_52155_new_n20116_; 
wire u2__abc_52155_new_n20117_; 
wire u2__abc_52155_new_n20118_; 
wire u2__abc_52155_new_n20119_; 
wire u2__abc_52155_new_n20120_; 
wire u2__abc_52155_new_n20121_; 
wire u2__abc_52155_new_n20122_; 
wire u2__abc_52155_new_n20124_; 
wire u2__abc_52155_new_n20125_; 
wire u2__abc_52155_new_n20126_; 
wire u2__abc_52155_new_n20127_; 
wire u2__abc_52155_new_n20128_; 
wire u2__abc_52155_new_n20129_; 
wire u2__abc_52155_new_n20130_; 
wire u2__abc_52155_new_n20131_; 
wire u2__abc_52155_new_n20132_; 
wire u2__abc_52155_new_n20133_; 
wire u2__abc_52155_new_n20134_; 
wire u2__abc_52155_new_n20136_; 
wire u2__abc_52155_new_n20137_; 
wire u2__abc_52155_new_n20138_; 
wire u2__abc_52155_new_n20139_; 
wire u2__abc_52155_new_n20140_; 
wire u2__abc_52155_new_n20141_; 
wire u2__abc_52155_new_n20142_; 
wire u2__abc_52155_new_n20143_; 
wire u2__abc_52155_new_n20144_; 
wire u2__abc_52155_new_n20145_; 
wire u2__abc_52155_new_n20146_; 
wire u2__abc_52155_new_n20148_; 
wire u2__abc_52155_new_n20149_; 
wire u2__abc_52155_new_n20150_; 
wire u2__abc_52155_new_n20151_; 
wire u2__abc_52155_new_n20152_; 
wire u2__abc_52155_new_n20153_; 
wire u2__abc_52155_new_n20154_; 
wire u2__abc_52155_new_n20155_; 
wire u2__abc_52155_new_n20156_; 
wire u2__abc_52155_new_n20157_; 
wire u2__abc_52155_new_n20158_; 
wire u2__abc_52155_new_n20160_; 
wire u2__abc_52155_new_n20161_; 
wire u2__abc_52155_new_n20162_; 
wire u2__abc_52155_new_n20163_; 
wire u2__abc_52155_new_n20164_; 
wire u2__abc_52155_new_n20165_; 
wire u2__abc_52155_new_n20166_; 
wire u2__abc_52155_new_n20167_; 
wire u2__abc_52155_new_n20168_; 
wire u2__abc_52155_new_n20169_; 
wire u2__abc_52155_new_n20170_; 
wire u2__abc_52155_new_n20172_; 
wire u2__abc_52155_new_n20173_; 
wire u2__abc_52155_new_n20174_; 
wire u2__abc_52155_new_n20175_; 
wire u2__abc_52155_new_n20176_; 
wire u2__abc_52155_new_n20177_; 
wire u2__abc_52155_new_n20178_; 
wire u2__abc_52155_new_n20179_; 
wire u2__abc_52155_new_n20180_; 
wire u2__abc_52155_new_n20181_; 
wire u2__abc_52155_new_n20182_; 
wire u2__abc_52155_new_n20184_; 
wire u2__abc_52155_new_n20185_; 
wire u2__abc_52155_new_n20186_; 
wire u2__abc_52155_new_n20187_; 
wire u2__abc_52155_new_n20188_; 
wire u2__abc_52155_new_n20189_; 
wire u2__abc_52155_new_n20190_; 
wire u2__abc_52155_new_n20191_; 
wire u2__abc_52155_new_n20192_; 
wire u2__abc_52155_new_n20193_; 
wire u2__abc_52155_new_n20194_; 
wire u2__abc_52155_new_n20196_; 
wire u2__abc_52155_new_n20197_; 
wire u2__abc_52155_new_n20198_; 
wire u2__abc_52155_new_n20199_; 
wire u2__abc_52155_new_n20200_; 
wire u2__abc_52155_new_n20201_; 
wire u2__abc_52155_new_n20202_; 
wire u2__abc_52155_new_n20203_; 
wire u2__abc_52155_new_n20204_; 
wire u2__abc_52155_new_n20205_; 
wire u2__abc_52155_new_n20206_; 
wire u2__abc_52155_new_n20208_; 
wire u2__abc_52155_new_n20209_; 
wire u2__abc_52155_new_n20210_; 
wire u2__abc_52155_new_n20211_; 
wire u2__abc_52155_new_n20212_; 
wire u2__abc_52155_new_n20213_; 
wire u2__abc_52155_new_n20214_; 
wire u2__abc_52155_new_n20215_; 
wire u2__abc_52155_new_n20216_; 
wire u2__abc_52155_new_n20217_; 
wire u2__abc_52155_new_n20218_; 
wire u2__abc_52155_new_n20220_; 
wire u2__abc_52155_new_n20221_; 
wire u2__abc_52155_new_n20222_; 
wire u2__abc_52155_new_n20223_; 
wire u2__abc_52155_new_n20224_; 
wire u2__abc_52155_new_n20225_; 
wire u2__abc_52155_new_n20226_; 
wire u2__abc_52155_new_n20227_; 
wire u2__abc_52155_new_n20228_; 
wire u2__abc_52155_new_n20229_; 
wire u2__abc_52155_new_n20230_; 
wire u2__abc_52155_new_n20232_; 
wire u2__abc_52155_new_n20233_; 
wire u2__abc_52155_new_n20234_; 
wire u2__abc_52155_new_n20235_; 
wire u2__abc_52155_new_n20236_; 
wire u2__abc_52155_new_n20237_; 
wire u2__abc_52155_new_n20238_; 
wire u2__abc_52155_new_n20239_; 
wire u2__abc_52155_new_n20240_; 
wire u2__abc_52155_new_n20241_; 
wire u2__abc_52155_new_n20242_; 
wire u2__abc_52155_new_n20244_; 
wire u2__abc_52155_new_n20245_; 
wire u2__abc_52155_new_n20246_; 
wire u2__abc_52155_new_n20247_; 
wire u2__abc_52155_new_n20248_; 
wire u2__abc_52155_new_n20249_; 
wire u2__abc_52155_new_n20250_; 
wire u2__abc_52155_new_n20251_; 
wire u2__abc_52155_new_n20252_; 
wire u2__abc_52155_new_n20253_; 
wire u2__abc_52155_new_n20254_; 
wire u2__abc_52155_new_n20256_; 
wire u2__abc_52155_new_n20257_; 
wire u2__abc_52155_new_n20258_; 
wire u2__abc_52155_new_n20259_; 
wire u2__abc_52155_new_n20260_; 
wire u2__abc_52155_new_n20261_; 
wire u2__abc_52155_new_n20262_; 
wire u2__abc_52155_new_n20263_; 
wire u2__abc_52155_new_n20264_; 
wire u2__abc_52155_new_n20265_; 
wire u2__abc_52155_new_n20266_; 
wire u2__abc_52155_new_n20268_; 
wire u2__abc_52155_new_n20269_; 
wire u2__abc_52155_new_n20270_; 
wire u2__abc_52155_new_n20271_; 
wire u2__abc_52155_new_n20272_; 
wire u2__abc_52155_new_n20273_; 
wire u2__abc_52155_new_n20274_; 
wire u2__abc_52155_new_n20275_; 
wire u2__abc_52155_new_n20276_; 
wire u2__abc_52155_new_n20277_; 
wire u2__abc_52155_new_n20278_; 
wire u2__abc_52155_new_n20280_; 
wire u2__abc_52155_new_n20281_; 
wire u2__abc_52155_new_n20282_; 
wire u2__abc_52155_new_n20283_; 
wire u2__abc_52155_new_n20284_; 
wire u2__abc_52155_new_n20285_; 
wire u2__abc_52155_new_n20286_; 
wire u2__abc_52155_new_n20287_; 
wire u2__abc_52155_new_n20288_; 
wire u2__abc_52155_new_n20289_; 
wire u2__abc_52155_new_n20290_; 
wire u2__abc_52155_new_n20292_; 
wire u2__abc_52155_new_n20293_; 
wire u2__abc_52155_new_n20294_; 
wire u2__abc_52155_new_n20295_; 
wire u2__abc_52155_new_n20296_; 
wire u2__abc_52155_new_n20297_; 
wire u2__abc_52155_new_n20298_; 
wire u2__abc_52155_new_n20299_; 
wire u2__abc_52155_new_n20300_; 
wire u2__abc_52155_new_n20301_; 
wire u2__abc_52155_new_n20302_; 
wire u2__abc_52155_new_n20304_; 
wire u2__abc_52155_new_n20305_; 
wire u2__abc_52155_new_n20306_; 
wire u2__abc_52155_new_n20307_; 
wire u2__abc_52155_new_n20308_; 
wire u2__abc_52155_new_n20309_; 
wire u2__abc_52155_new_n20310_; 
wire u2__abc_52155_new_n20311_; 
wire u2__abc_52155_new_n20312_; 
wire u2__abc_52155_new_n20313_; 
wire u2__abc_52155_new_n20314_; 
wire u2__abc_52155_new_n20316_; 
wire u2__abc_52155_new_n20317_; 
wire u2__abc_52155_new_n20318_; 
wire u2__abc_52155_new_n20319_; 
wire u2__abc_52155_new_n20320_; 
wire u2__abc_52155_new_n20321_; 
wire u2__abc_52155_new_n20322_; 
wire u2__abc_52155_new_n20323_; 
wire u2__abc_52155_new_n20324_; 
wire u2__abc_52155_new_n20325_; 
wire u2__abc_52155_new_n20326_; 
wire u2__abc_52155_new_n20328_; 
wire u2__abc_52155_new_n20329_; 
wire u2__abc_52155_new_n20330_; 
wire u2__abc_52155_new_n20331_; 
wire u2__abc_52155_new_n20332_; 
wire u2__abc_52155_new_n20333_; 
wire u2__abc_52155_new_n20334_; 
wire u2__abc_52155_new_n20335_; 
wire u2__abc_52155_new_n20336_; 
wire u2__abc_52155_new_n20337_; 
wire u2__abc_52155_new_n20338_; 
wire u2__abc_52155_new_n20340_; 
wire u2__abc_52155_new_n20341_; 
wire u2__abc_52155_new_n20342_; 
wire u2__abc_52155_new_n20343_; 
wire u2__abc_52155_new_n20344_; 
wire u2__abc_52155_new_n20345_; 
wire u2__abc_52155_new_n20346_; 
wire u2__abc_52155_new_n20347_; 
wire u2__abc_52155_new_n20348_; 
wire u2__abc_52155_new_n20349_; 
wire u2__abc_52155_new_n20350_; 
wire u2__abc_52155_new_n20352_; 
wire u2__abc_52155_new_n20353_; 
wire u2__abc_52155_new_n20354_; 
wire u2__abc_52155_new_n20355_; 
wire u2__abc_52155_new_n20356_; 
wire u2__abc_52155_new_n20357_; 
wire u2__abc_52155_new_n20358_; 
wire u2__abc_52155_new_n20359_; 
wire u2__abc_52155_new_n20360_; 
wire u2__abc_52155_new_n20361_; 
wire u2__abc_52155_new_n20362_; 
wire u2__abc_52155_new_n20364_; 
wire u2__abc_52155_new_n20365_; 
wire u2__abc_52155_new_n20366_; 
wire u2__abc_52155_new_n20367_; 
wire u2__abc_52155_new_n20368_; 
wire u2__abc_52155_new_n20369_; 
wire u2__abc_52155_new_n20370_; 
wire u2__abc_52155_new_n20371_; 
wire u2__abc_52155_new_n20372_; 
wire u2__abc_52155_new_n20373_; 
wire u2__abc_52155_new_n20374_; 
wire u2__abc_52155_new_n20376_; 
wire u2__abc_52155_new_n20377_; 
wire u2__abc_52155_new_n20378_; 
wire u2__abc_52155_new_n20379_; 
wire u2__abc_52155_new_n20380_; 
wire u2__abc_52155_new_n20381_; 
wire u2__abc_52155_new_n20382_; 
wire u2__abc_52155_new_n20383_; 
wire u2__abc_52155_new_n20384_; 
wire u2__abc_52155_new_n20385_; 
wire u2__abc_52155_new_n20386_; 
wire u2__abc_52155_new_n20388_; 
wire u2__abc_52155_new_n20389_; 
wire u2__abc_52155_new_n20390_; 
wire u2__abc_52155_new_n20391_; 
wire u2__abc_52155_new_n20392_; 
wire u2__abc_52155_new_n20393_; 
wire u2__abc_52155_new_n20394_; 
wire u2__abc_52155_new_n20395_; 
wire u2__abc_52155_new_n20396_; 
wire u2__abc_52155_new_n20397_; 
wire u2__abc_52155_new_n20398_; 
wire u2__abc_52155_new_n20400_; 
wire u2__abc_52155_new_n20401_; 
wire u2__abc_52155_new_n20402_; 
wire u2__abc_52155_new_n20403_; 
wire u2__abc_52155_new_n20404_; 
wire u2__abc_52155_new_n20405_; 
wire u2__abc_52155_new_n20406_; 
wire u2__abc_52155_new_n20407_; 
wire u2__abc_52155_new_n20408_; 
wire u2__abc_52155_new_n20409_; 
wire u2__abc_52155_new_n20410_; 
wire u2__abc_52155_new_n20412_; 
wire u2__abc_52155_new_n20413_; 
wire u2__abc_52155_new_n20414_; 
wire u2__abc_52155_new_n20415_; 
wire u2__abc_52155_new_n20416_; 
wire u2__abc_52155_new_n20417_; 
wire u2__abc_52155_new_n20418_; 
wire u2__abc_52155_new_n20419_; 
wire u2__abc_52155_new_n20420_; 
wire u2__abc_52155_new_n20421_; 
wire u2__abc_52155_new_n20422_; 
wire u2__abc_52155_new_n20424_; 
wire u2__abc_52155_new_n20425_; 
wire u2__abc_52155_new_n20426_; 
wire u2__abc_52155_new_n20427_; 
wire u2__abc_52155_new_n20428_; 
wire u2__abc_52155_new_n20429_; 
wire u2__abc_52155_new_n20430_; 
wire u2__abc_52155_new_n20431_; 
wire u2__abc_52155_new_n20432_; 
wire u2__abc_52155_new_n20433_; 
wire u2__abc_52155_new_n20434_; 
wire u2__abc_52155_new_n20436_; 
wire u2__abc_52155_new_n20437_; 
wire u2__abc_52155_new_n20438_; 
wire u2__abc_52155_new_n20439_; 
wire u2__abc_52155_new_n20440_; 
wire u2__abc_52155_new_n20441_; 
wire u2__abc_52155_new_n20442_; 
wire u2__abc_52155_new_n20443_; 
wire u2__abc_52155_new_n20444_; 
wire u2__abc_52155_new_n20445_; 
wire u2__abc_52155_new_n20446_; 
wire u2__abc_52155_new_n20448_; 
wire u2__abc_52155_new_n20449_; 
wire u2__abc_52155_new_n20450_; 
wire u2__abc_52155_new_n20451_; 
wire u2__abc_52155_new_n20452_; 
wire u2__abc_52155_new_n20453_; 
wire u2__abc_52155_new_n20454_; 
wire u2__abc_52155_new_n20455_; 
wire u2__abc_52155_new_n20456_; 
wire u2__abc_52155_new_n20457_; 
wire u2__abc_52155_new_n20458_; 
wire u2__abc_52155_new_n20460_; 
wire u2__abc_52155_new_n20461_; 
wire u2__abc_52155_new_n20462_; 
wire u2__abc_52155_new_n20463_; 
wire u2__abc_52155_new_n20464_; 
wire u2__abc_52155_new_n20465_; 
wire u2__abc_52155_new_n20466_; 
wire u2__abc_52155_new_n20467_; 
wire u2__abc_52155_new_n20468_; 
wire u2__abc_52155_new_n20469_; 
wire u2__abc_52155_new_n20470_; 
wire u2__abc_52155_new_n20472_; 
wire u2__abc_52155_new_n20473_; 
wire u2__abc_52155_new_n20474_; 
wire u2__abc_52155_new_n20475_; 
wire u2__abc_52155_new_n20476_; 
wire u2__abc_52155_new_n20477_; 
wire u2__abc_52155_new_n20478_; 
wire u2__abc_52155_new_n20479_; 
wire u2__abc_52155_new_n20480_; 
wire u2__abc_52155_new_n20481_; 
wire u2__abc_52155_new_n20482_; 
wire u2__abc_52155_new_n20484_; 
wire u2__abc_52155_new_n20485_; 
wire u2__abc_52155_new_n20486_; 
wire u2__abc_52155_new_n20487_; 
wire u2__abc_52155_new_n20488_; 
wire u2__abc_52155_new_n20489_; 
wire u2__abc_52155_new_n20490_; 
wire u2__abc_52155_new_n20491_; 
wire u2__abc_52155_new_n20492_; 
wire u2__abc_52155_new_n20493_; 
wire u2__abc_52155_new_n20494_; 
wire u2__abc_52155_new_n20496_; 
wire u2__abc_52155_new_n20497_; 
wire u2__abc_52155_new_n20498_; 
wire u2__abc_52155_new_n20499_; 
wire u2__abc_52155_new_n20500_; 
wire u2__abc_52155_new_n20501_; 
wire u2__abc_52155_new_n20502_; 
wire u2__abc_52155_new_n20503_; 
wire u2__abc_52155_new_n20504_; 
wire u2__abc_52155_new_n20505_; 
wire u2__abc_52155_new_n20506_; 
wire u2__abc_52155_new_n20508_; 
wire u2__abc_52155_new_n20509_; 
wire u2__abc_52155_new_n20510_; 
wire u2__abc_52155_new_n20511_; 
wire u2__abc_52155_new_n20512_; 
wire u2__abc_52155_new_n20513_; 
wire u2__abc_52155_new_n20514_; 
wire u2__abc_52155_new_n20515_; 
wire u2__abc_52155_new_n20516_; 
wire u2__abc_52155_new_n20517_; 
wire u2__abc_52155_new_n20518_; 
wire u2__abc_52155_new_n20520_; 
wire u2__abc_52155_new_n20521_; 
wire u2__abc_52155_new_n20522_; 
wire u2__abc_52155_new_n20523_; 
wire u2__abc_52155_new_n20524_; 
wire u2__abc_52155_new_n20525_; 
wire u2__abc_52155_new_n20526_; 
wire u2__abc_52155_new_n20527_; 
wire u2__abc_52155_new_n20528_; 
wire u2__abc_52155_new_n20529_; 
wire u2__abc_52155_new_n20530_; 
wire u2__abc_52155_new_n20532_; 
wire u2__abc_52155_new_n20533_; 
wire u2__abc_52155_new_n20534_; 
wire u2__abc_52155_new_n20535_; 
wire u2__abc_52155_new_n20536_; 
wire u2__abc_52155_new_n20537_; 
wire u2__abc_52155_new_n20538_; 
wire u2__abc_52155_new_n20539_; 
wire u2__abc_52155_new_n20540_; 
wire u2__abc_52155_new_n20541_; 
wire u2__abc_52155_new_n20542_; 
wire u2__abc_52155_new_n20544_; 
wire u2__abc_52155_new_n20545_; 
wire u2__abc_52155_new_n20546_; 
wire u2__abc_52155_new_n20547_; 
wire u2__abc_52155_new_n20548_; 
wire u2__abc_52155_new_n20549_; 
wire u2__abc_52155_new_n20550_; 
wire u2__abc_52155_new_n20551_; 
wire u2__abc_52155_new_n20552_; 
wire u2__abc_52155_new_n20553_; 
wire u2__abc_52155_new_n20554_; 
wire u2__abc_52155_new_n20556_; 
wire u2__abc_52155_new_n20557_; 
wire u2__abc_52155_new_n20558_; 
wire u2__abc_52155_new_n20559_; 
wire u2__abc_52155_new_n20560_; 
wire u2__abc_52155_new_n20561_; 
wire u2__abc_52155_new_n20562_; 
wire u2__abc_52155_new_n20563_; 
wire u2__abc_52155_new_n20564_; 
wire u2__abc_52155_new_n20565_; 
wire u2__abc_52155_new_n20566_; 
wire u2__abc_52155_new_n20568_; 
wire u2__abc_52155_new_n20569_; 
wire u2__abc_52155_new_n20570_; 
wire u2__abc_52155_new_n20571_; 
wire u2__abc_52155_new_n20572_; 
wire u2__abc_52155_new_n20573_; 
wire u2__abc_52155_new_n20574_; 
wire u2__abc_52155_new_n20575_; 
wire u2__abc_52155_new_n20576_; 
wire u2__abc_52155_new_n20577_; 
wire u2__abc_52155_new_n20578_; 
wire u2__abc_52155_new_n20580_; 
wire u2__abc_52155_new_n20581_; 
wire u2__abc_52155_new_n20582_; 
wire u2__abc_52155_new_n20583_; 
wire u2__abc_52155_new_n20584_; 
wire u2__abc_52155_new_n20585_; 
wire u2__abc_52155_new_n20586_; 
wire u2__abc_52155_new_n20587_; 
wire u2__abc_52155_new_n20588_; 
wire u2__abc_52155_new_n20589_; 
wire u2__abc_52155_new_n20590_; 
wire u2__abc_52155_new_n20592_; 
wire u2__abc_52155_new_n20593_; 
wire u2__abc_52155_new_n20594_; 
wire u2__abc_52155_new_n20595_; 
wire u2__abc_52155_new_n20596_; 
wire u2__abc_52155_new_n20597_; 
wire u2__abc_52155_new_n20598_; 
wire u2__abc_52155_new_n20599_; 
wire u2__abc_52155_new_n20600_; 
wire u2__abc_52155_new_n20601_; 
wire u2__abc_52155_new_n20602_; 
wire u2__abc_52155_new_n20604_; 
wire u2__abc_52155_new_n20605_; 
wire u2__abc_52155_new_n20606_; 
wire u2__abc_52155_new_n20607_; 
wire u2__abc_52155_new_n20608_; 
wire u2__abc_52155_new_n20609_; 
wire u2__abc_52155_new_n20610_; 
wire u2__abc_52155_new_n20611_; 
wire u2__abc_52155_new_n20612_; 
wire u2__abc_52155_new_n20613_; 
wire u2__abc_52155_new_n20614_; 
wire u2__abc_52155_new_n20616_; 
wire u2__abc_52155_new_n20617_; 
wire u2__abc_52155_new_n20618_; 
wire u2__abc_52155_new_n20619_; 
wire u2__abc_52155_new_n20620_; 
wire u2__abc_52155_new_n20621_; 
wire u2__abc_52155_new_n20622_; 
wire u2__abc_52155_new_n20623_; 
wire u2__abc_52155_new_n20624_; 
wire u2__abc_52155_new_n20625_; 
wire u2__abc_52155_new_n20626_; 
wire u2__abc_52155_new_n20628_; 
wire u2__abc_52155_new_n20629_; 
wire u2__abc_52155_new_n20630_; 
wire u2__abc_52155_new_n20631_; 
wire u2__abc_52155_new_n20632_; 
wire u2__abc_52155_new_n20633_; 
wire u2__abc_52155_new_n20634_; 
wire u2__abc_52155_new_n20635_; 
wire u2__abc_52155_new_n20636_; 
wire u2__abc_52155_new_n20637_; 
wire u2__abc_52155_new_n20638_; 
wire u2__abc_52155_new_n20640_; 
wire u2__abc_52155_new_n20641_; 
wire u2__abc_52155_new_n20642_; 
wire u2__abc_52155_new_n20643_; 
wire u2__abc_52155_new_n20644_; 
wire u2__abc_52155_new_n20645_; 
wire u2__abc_52155_new_n20646_; 
wire u2__abc_52155_new_n20647_; 
wire u2__abc_52155_new_n20648_; 
wire u2__abc_52155_new_n20649_; 
wire u2__abc_52155_new_n20650_; 
wire u2__abc_52155_new_n20652_; 
wire u2__abc_52155_new_n20653_; 
wire u2__abc_52155_new_n20654_; 
wire u2__abc_52155_new_n20655_; 
wire u2__abc_52155_new_n20656_; 
wire u2__abc_52155_new_n20657_; 
wire u2__abc_52155_new_n20658_; 
wire u2__abc_52155_new_n20659_; 
wire u2__abc_52155_new_n20660_; 
wire u2__abc_52155_new_n20661_; 
wire u2__abc_52155_new_n20662_; 
wire u2__abc_52155_new_n20664_; 
wire u2__abc_52155_new_n20665_; 
wire u2__abc_52155_new_n20666_; 
wire u2__abc_52155_new_n20667_; 
wire u2__abc_52155_new_n20668_; 
wire u2__abc_52155_new_n20669_; 
wire u2__abc_52155_new_n20670_; 
wire u2__abc_52155_new_n20671_; 
wire u2__abc_52155_new_n20672_; 
wire u2__abc_52155_new_n20673_; 
wire u2__abc_52155_new_n20674_; 
wire u2__abc_52155_new_n20676_; 
wire u2__abc_52155_new_n20677_; 
wire u2__abc_52155_new_n20678_; 
wire u2__abc_52155_new_n20679_; 
wire u2__abc_52155_new_n20680_; 
wire u2__abc_52155_new_n20681_; 
wire u2__abc_52155_new_n20682_; 
wire u2__abc_52155_new_n20683_; 
wire u2__abc_52155_new_n20684_; 
wire u2__abc_52155_new_n20685_; 
wire u2__abc_52155_new_n20686_; 
wire u2__abc_52155_new_n20688_; 
wire u2__abc_52155_new_n20689_; 
wire u2__abc_52155_new_n20690_; 
wire u2__abc_52155_new_n20691_; 
wire u2__abc_52155_new_n20692_; 
wire u2__abc_52155_new_n20693_; 
wire u2__abc_52155_new_n20694_; 
wire u2__abc_52155_new_n20695_; 
wire u2__abc_52155_new_n20696_; 
wire u2__abc_52155_new_n20697_; 
wire u2__abc_52155_new_n20698_; 
wire u2__abc_52155_new_n20700_; 
wire u2__abc_52155_new_n20701_; 
wire u2__abc_52155_new_n20702_; 
wire u2__abc_52155_new_n20703_; 
wire u2__abc_52155_new_n20704_; 
wire u2__abc_52155_new_n20705_; 
wire u2__abc_52155_new_n20706_; 
wire u2__abc_52155_new_n20707_; 
wire u2__abc_52155_new_n20708_; 
wire u2__abc_52155_new_n20709_; 
wire u2__abc_52155_new_n20710_; 
wire u2__abc_52155_new_n20712_; 
wire u2__abc_52155_new_n20713_; 
wire u2__abc_52155_new_n20714_; 
wire u2__abc_52155_new_n20715_; 
wire u2__abc_52155_new_n20716_; 
wire u2__abc_52155_new_n20717_; 
wire u2__abc_52155_new_n20718_; 
wire u2__abc_52155_new_n20719_; 
wire u2__abc_52155_new_n20720_; 
wire u2__abc_52155_new_n20721_; 
wire u2__abc_52155_new_n20722_; 
wire u2__abc_52155_new_n20724_; 
wire u2__abc_52155_new_n20725_; 
wire u2__abc_52155_new_n20726_; 
wire u2__abc_52155_new_n20727_; 
wire u2__abc_52155_new_n20728_; 
wire u2__abc_52155_new_n20729_; 
wire u2__abc_52155_new_n20730_; 
wire u2__abc_52155_new_n20731_; 
wire u2__abc_52155_new_n20732_; 
wire u2__abc_52155_new_n20733_; 
wire u2__abc_52155_new_n20734_; 
wire u2__abc_52155_new_n20736_; 
wire u2__abc_52155_new_n20737_; 
wire u2__abc_52155_new_n20738_; 
wire u2__abc_52155_new_n20739_; 
wire u2__abc_52155_new_n20740_; 
wire u2__abc_52155_new_n20741_; 
wire u2__abc_52155_new_n20742_; 
wire u2__abc_52155_new_n20743_; 
wire u2__abc_52155_new_n20744_; 
wire u2__abc_52155_new_n20745_; 
wire u2__abc_52155_new_n20746_; 
wire u2__abc_52155_new_n20748_; 
wire u2__abc_52155_new_n20749_; 
wire u2__abc_52155_new_n20750_; 
wire u2__abc_52155_new_n20751_; 
wire u2__abc_52155_new_n20752_; 
wire u2__abc_52155_new_n20753_; 
wire u2__abc_52155_new_n20754_; 
wire u2__abc_52155_new_n20755_; 
wire u2__abc_52155_new_n20756_; 
wire u2__abc_52155_new_n20757_; 
wire u2__abc_52155_new_n20758_; 
wire u2__abc_52155_new_n20760_; 
wire u2__abc_52155_new_n20761_; 
wire u2__abc_52155_new_n20762_; 
wire u2__abc_52155_new_n20763_; 
wire u2__abc_52155_new_n20764_; 
wire u2__abc_52155_new_n20765_; 
wire u2__abc_52155_new_n20766_; 
wire u2__abc_52155_new_n20767_; 
wire u2__abc_52155_new_n20768_; 
wire u2__abc_52155_new_n20769_; 
wire u2__abc_52155_new_n20770_; 
wire u2__abc_52155_new_n20772_; 
wire u2__abc_52155_new_n20773_; 
wire u2__abc_52155_new_n20774_; 
wire u2__abc_52155_new_n20775_; 
wire u2__abc_52155_new_n20776_; 
wire u2__abc_52155_new_n20777_; 
wire u2__abc_52155_new_n20778_; 
wire u2__abc_52155_new_n20779_; 
wire u2__abc_52155_new_n20780_; 
wire u2__abc_52155_new_n20781_; 
wire u2__abc_52155_new_n20782_; 
wire u2__abc_52155_new_n20784_; 
wire u2__abc_52155_new_n20785_; 
wire u2__abc_52155_new_n20786_; 
wire u2__abc_52155_new_n20787_; 
wire u2__abc_52155_new_n20788_; 
wire u2__abc_52155_new_n20789_; 
wire u2__abc_52155_new_n20790_; 
wire u2__abc_52155_new_n20791_; 
wire u2__abc_52155_new_n20792_; 
wire u2__abc_52155_new_n20793_; 
wire u2__abc_52155_new_n20794_; 
wire u2__abc_52155_new_n20796_; 
wire u2__abc_52155_new_n20797_; 
wire u2__abc_52155_new_n20798_; 
wire u2__abc_52155_new_n20799_; 
wire u2__abc_52155_new_n20800_; 
wire u2__abc_52155_new_n20801_; 
wire u2__abc_52155_new_n20802_; 
wire u2__abc_52155_new_n20803_; 
wire u2__abc_52155_new_n20804_; 
wire u2__abc_52155_new_n20805_; 
wire u2__abc_52155_new_n20806_; 
wire u2__abc_52155_new_n20808_; 
wire u2__abc_52155_new_n20809_; 
wire u2__abc_52155_new_n20810_; 
wire u2__abc_52155_new_n20811_; 
wire u2__abc_52155_new_n20812_; 
wire u2__abc_52155_new_n20813_; 
wire u2__abc_52155_new_n20814_; 
wire u2__abc_52155_new_n20815_; 
wire u2__abc_52155_new_n20816_; 
wire u2__abc_52155_new_n20817_; 
wire u2__abc_52155_new_n20818_; 
wire u2__abc_52155_new_n20820_; 
wire u2__abc_52155_new_n20821_; 
wire u2__abc_52155_new_n20822_; 
wire u2__abc_52155_new_n20823_; 
wire u2__abc_52155_new_n20824_; 
wire u2__abc_52155_new_n20825_; 
wire u2__abc_52155_new_n20826_; 
wire u2__abc_52155_new_n20827_; 
wire u2__abc_52155_new_n20828_; 
wire u2__abc_52155_new_n20829_; 
wire u2__abc_52155_new_n20830_; 
wire u2__abc_52155_new_n20832_; 
wire u2__abc_52155_new_n20833_; 
wire u2__abc_52155_new_n20834_; 
wire u2__abc_52155_new_n20835_; 
wire u2__abc_52155_new_n20836_; 
wire u2__abc_52155_new_n20837_; 
wire u2__abc_52155_new_n20838_; 
wire u2__abc_52155_new_n20839_; 
wire u2__abc_52155_new_n20840_; 
wire u2__abc_52155_new_n20841_; 
wire u2__abc_52155_new_n20842_; 
wire u2__abc_52155_new_n20844_; 
wire u2__abc_52155_new_n20845_; 
wire u2__abc_52155_new_n20846_; 
wire u2__abc_52155_new_n20847_; 
wire u2__abc_52155_new_n20848_; 
wire u2__abc_52155_new_n20849_; 
wire u2__abc_52155_new_n20850_; 
wire u2__abc_52155_new_n20851_; 
wire u2__abc_52155_new_n20852_; 
wire u2__abc_52155_new_n20853_; 
wire u2__abc_52155_new_n20854_; 
wire u2__abc_52155_new_n20856_; 
wire u2__abc_52155_new_n20857_; 
wire u2__abc_52155_new_n20858_; 
wire u2__abc_52155_new_n20859_; 
wire u2__abc_52155_new_n20860_; 
wire u2__abc_52155_new_n20861_; 
wire u2__abc_52155_new_n20862_; 
wire u2__abc_52155_new_n20863_; 
wire u2__abc_52155_new_n20864_; 
wire u2__abc_52155_new_n20865_; 
wire u2__abc_52155_new_n20866_; 
wire u2__abc_52155_new_n20868_; 
wire u2__abc_52155_new_n20869_; 
wire u2__abc_52155_new_n20870_; 
wire u2__abc_52155_new_n20871_; 
wire u2__abc_52155_new_n20872_; 
wire u2__abc_52155_new_n20873_; 
wire u2__abc_52155_new_n20874_; 
wire u2__abc_52155_new_n20875_; 
wire u2__abc_52155_new_n20876_; 
wire u2__abc_52155_new_n20877_; 
wire u2__abc_52155_new_n20878_; 
wire u2__abc_52155_new_n20880_; 
wire u2__abc_52155_new_n20881_; 
wire u2__abc_52155_new_n20882_; 
wire u2__abc_52155_new_n20883_; 
wire u2__abc_52155_new_n20884_; 
wire u2__abc_52155_new_n20885_; 
wire u2__abc_52155_new_n20886_; 
wire u2__abc_52155_new_n20887_; 
wire u2__abc_52155_new_n20888_; 
wire u2__abc_52155_new_n20889_; 
wire u2__abc_52155_new_n20890_; 
wire u2__abc_52155_new_n20892_; 
wire u2__abc_52155_new_n20893_; 
wire u2__abc_52155_new_n20894_; 
wire u2__abc_52155_new_n20895_; 
wire u2__abc_52155_new_n20896_; 
wire u2__abc_52155_new_n20897_; 
wire u2__abc_52155_new_n20898_; 
wire u2__abc_52155_new_n20899_; 
wire u2__abc_52155_new_n20900_; 
wire u2__abc_52155_new_n20901_; 
wire u2__abc_52155_new_n20902_; 
wire u2__abc_52155_new_n20904_; 
wire u2__abc_52155_new_n20905_; 
wire u2__abc_52155_new_n20906_; 
wire u2__abc_52155_new_n20907_; 
wire u2__abc_52155_new_n20908_; 
wire u2__abc_52155_new_n20909_; 
wire u2__abc_52155_new_n20910_; 
wire u2__abc_52155_new_n20911_; 
wire u2__abc_52155_new_n20912_; 
wire u2__abc_52155_new_n20913_; 
wire u2__abc_52155_new_n20914_; 
wire u2__abc_52155_new_n20916_; 
wire u2__abc_52155_new_n20917_; 
wire u2__abc_52155_new_n20918_; 
wire u2__abc_52155_new_n20919_; 
wire u2__abc_52155_new_n20920_; 
wire u2__abc_52155_new_n20921_; 
wire u2__abc_52155_new_n20922_; 
wire u2__abc_52155_new_n20923_; 
wire u2__abc_52155_new_n20924_; 
wire u2__abc_52155_new_n20925_; 
wire u2__abc_52155_new_n20926_; 
wire u2__abc_52155_new_n20928_; 
wire u2__abc_52155_new_n20929_; 
wire u2__abc_52155_new_n20930_; 
wire u2__abc_52155_new_n20931_; 
wire u2__abc_52155_new_n20932_; 
wire u2__abc_52155_new_n20933_; 
wire u2__abc_52155_new_n20934_; 
wire u2__abc_52155_new_n20935_; 
wire u2__abc_52155_new_n20936_; 
wire u2__abc_52155_new_n20937_; 
wire u2__abc_52155_new_n20938_; 
wire u2__abc_52155_new_n20940_; 
wire u2__abc_52155_new_n20941_; 
wire u2__abc_52155_new_n20942_; 
wire u2__abc_52155_new_n20943_; 
wire u2__abc_52155_new_n20944_; 
wire u2__abc_52155_new_n20945_; 
wire u2__abc_52155_new_n20946_; 
wire u2__abc_52155_new_n20947_; 
wire u2__abc_52155_new_n20948_; 
wire u2__abc_52155_new_n20949_; 
wire u2__abc_52155_new_n20950_; 
wire u2__abc_52155_new_n20952_; 
wire u2__abc_52155_new_n20953_; 
wire u2__abc_52155_new_n20954_; 
wire u2__abc_52155_new_n20955_; 
wire u2__abc_52155_new_n20956_; 
wire u2__abc_52155_new_n20957_; 
wire u2__abc_52155_new_n20958_; 
wire u2__abc_52155_new_n20959_; 
wire u2__abc_52155_new_n20960_; 
wire u2__abc_52155_new_n20961_; 
wire u2__abc_52155_new_n20962_; 
wire u2__abc_52155_new_n20964_; 
wire u2__abc_52155_new_n20965_; 
wire u2__abc_52155_new_n20966_; 
wire u2__abc_52155_new_n20967_; 
wire u2__abc_52155_new_n20968_; 
wire u2__abc_52155_new_n20969_; 
wire u2__abc_52155_new_n20970_; 
wire u2__abc_52155_new_n20971_; 
wire u2__abc_52155_new_n20972_; 
wire u2__abc_52155_new_n20973_; 
wire u2__abc_52155_new_n20974_; 
wire u2__abc_52155_new_n20976_; 
wire u2__abc_52155_new_n20977_; 
wire u2__abc_52155_new_n20978_; 
wire u2__abc_52155_new_n20979_; 
wire u2__abc_52155_new_n20980_; 
wire u2__abc_52155_new_n20981_; 
wire u2__abc_52155_new_n20982_; 
wire u2__abc_52155_new_n20983_; 
wire u2__abc_52155_new_n20984_; 
wire u2__abc_52155_new_n20985_; 
wire u2__abc_52155_new_n20986_; 
wire u2__abc_52155_new_n20988_; 
wire u2__abc_52155_new_n20989_; 
wire u2__abc_52155_new_n20990_; 
wire u2__abc_52155_new_n20991_; 
wire u2__abc_52155_new_n20992_; 
wire u2__abc_52155_new_n20993_; 
wire u2__abc_52155_new_n20994_; 
wire u2__abc_52155_new_n20995_; 
wire u2__abc_52155_new_n20996_; 
wire u2__abc_52155_new_n20997_; 
wire u2__abc_52155_new_n20998_; 
wire u2__abc_52155_new_n21000_; 
wire u2__abc_52155_new_n21001_; 
wire u2__abc_52155_new_n21002_; 
wire u2__abc_52155_new_n21003_; 
wire u2__abc_52155_new_n21004_; 
wire u2__abc_52155_new_n21005_; 
wire u2__abc_52155_new_n21006_; 
wire u2__abc_52155_new_n21007_; 
wire u2__abc_52155_new_n21008_; 
wire u2__abc_52155_new_n21009_; 
wire u2__abc_52155_new_n21010_; 
wire u2__abc_52155_new_n21012_; 
wire u2__abc_52155_new_n21013_; 
wire u2__abc_52155_new_n21014_; 
wire u2__abc_52155_new_n21015_; 
wire u2__abc_52155_new_n21016_; 
wire u2__abc_52155_new_n21017_; 
wire u2__abc_52155_new_n21018_; 
wire u2__abc_52155_new_n21019_; 
wire u2__abc_52155_new_n21020_; 
wire u2__abc_52155_new_n21021_; 
wire u2__abc_52155_new_n21022_; 
wire u2__abc_52155_new_n21024_; 
wire u2__abc_52155_new_n21025_; 
wire u2__abc_52155_new_n21026_; 
wire u2__abc_52155_new_n21027_; 
wire u2__abc_52155_new_n21028_; 
wire u2__abc_52155_new_n21029_; 
wire u2__abc_52155_new_n21030_; 
wire u2__abc_52155_new_n21031_; 
wire u2__abc_52155_new_n21032_; 
wire u2__abc_52155_new_n21033_; 
wire u2__abc_52155_new_n21034_; 
wire u2__abc_52155_new_n21036_; 
wire u2__abc_52155_new_n21037_; 
wire u2__abc_52155_new_n21038_; 
wire u2__abc_52155_new_n21039_; 
wire u2__abc_52155_new_n21040_; 
wire u2__abc_52155_new_n21041_; 
wire u2__abc_52155_new_n21042_; 
wire u2__abc_52155_new_n21043_; 
wire u2__abc_52155_new_n21044_; 
wire u2__abc_52155_new_n21045_; 
wire u2__abc_52155_new_n21046_; 
wire u2__abc_52155_new_n21048_; 
wire u2__abc_52155_new_n21049_; 
wire u2__abc_52155_new_n21050_; 
wire u2__abc_52155_new_n21051_; 
wire u2__abc_52155_new_n21052_; 
wire u2__abc_52155_new_n21053_; 
wire u2__abc_52155_new_n21054_; 
wire u2__abc_52155_new_n21055_; 
wire u2__abc_52155_new_n21056_; 
wire u2__abc_52155_new_n21057_; 
wire u2__abc_52155_new_n21058_; 
wire u2__abc_52155_new_n21060_; 
wire u2__abc_52155_new_n21061_; 
wire u2__abc_52155_new_n21062_; 
wire u2__abc_52155_new_n21063_; 
wire u2__abc_52155_new_n21064_; 
wire u2__abc_52155_new_n21065_; 
wire u2__abc_52155_new_n21066_; 
wire u2__abc_52155_new_n21067_; 
wire u2__abc_52155_new_n21068_; 
wire u2__abc_52155_new_n21069_; 
wire u2__abc_52155_new_n21070_; 
wire u2__abc_52155_new_n21072_; 
wire u2__abc_52155_new_n21073_; 
wire u2__abc_52155_new_n21074_; 
wire u2__abc_52155_new_n21075_; 
wire u2__abc_52155_new_n21076_; 
wire u2__abc_52155_new_n21077_; 
wire u2__abc_52155_new_n21078_; 
wire u2__abc_52155_new_n21079_; 
wire u2__abc_52155_new_n21080_; 
wire u2__abc_52155_new_n21081_; 
wire u2__abc_52155_new_n21082_; 
wire u2__abc_52155_new_n21084_; 
wire u2__abc_52155_new_n21085_; 
wire u2__abc_52155_new_n21086_; 
wire u2__abc_52155_new_n21087_; 
wire u2__abc_52155_new_n21088_; 
wire u2__abc_52155_new_n21089_; 
wire u2__abc_52155_new_n21090_; 
wire u2__abc_52155_new_n21091_; 
wire u2__abc_52155_new_n21092_; 
wire u2__abc_52155_new_n21093_; 
wire u2__abc_52155_new_n21094_; 
wire u2__abc_52155_new_n21096_; 
wire u2__abc_52155_new_n21097_; 
wire u2__abc_52155_new_n21098_; 
wire u2__abc_52155_new_n21099_; 
wire u2__abc_52155_new_n21100_; 
wire u2__abc_52155_new_n21101_; 
wire u2__abc_52155_new_n21102_; 
wire u2__abc_52155_new_n21103_; 
wire u2__abc_52155_new_n21104_; 
wire u2__abc_52155_new_n21105_; 
wire u2__abc_52155_new_n21106_; 
wire u2__abc_52155_new_n21108_; 
wire u2__abc_52155_new_n21109_; 
wire u2__abc_52155_new_n21110_; 
wire u2__abc_52155_new_n21111_; 
wire u2__abc_52155_new_n21112_; 
wire u2__abc_52155_new_n21113_; 
wire u2__abc_52155_new_n21114_; 
wire u2__abc_52155_new_n21115_; 
wire u2__abc_52155_new_n21116_; 
wire u2__abc_52155_new_n21117_; 
wire u2__abc_52155_new_n21118_; 
wire u2__abc_52155_new_n21120_; 
wire u2__abc_52155_new_n21121_; 
wire u2__abc_52155_new_n21122_; 
wire u2__abc_52155_new_n21123_; 
wire u2__abc_52155_new_n21124_; 
wire u2__abc_52155_new_n21125_; 
wire u2__abc_52155_new_n21126_; 
wire u2__abc_52155_new_n21127_; 
wire u2__abc_52155_new_n21128_; 
wire u2__abc_52155_new_n21129_; 
wire u2__abc_52155_new_n21130_; 
wire u2__abc_52155_new_n21132_; 
wire u2__abc_52155_new_n21133_; 
wire u2__abc_52155_new_n21134_; 
wire u2__abc_52155_new_n21135_; 
wire u2__abc_52155_new_n21136_; 
wire u2__abc_52155_new_n21137_; 
wire u2__abc_52155_new_n21138_; 
wire u2__abc_52155_new_n21139_; 
wire u2__abc_52155_new_n21140_; 
wire u2__abc_52155_new_n21141_; 
wire u2__abc_52155_new_n21142_; 
wire u2__abc_52155_new_n21144_; 
wire u2__abc_52155_new_n21145_; 
wire u2__abc_52155_new_n21146_; 
wire u2__abc_52155_new_n21147_; 
wire u2__abc_52155_new_n21148_; 
wire u2__abc_52155_new_n21149_; 
wire u2__abc_52155_new_n21150_; 
wire u2__abc_52155_new_n21151_; 
wire u2__abc_52155_new_n21152_; 
wire u2__abc_52155_new_n21153_; 
wire u2__abc_52155_new_n21154_; 
wire u2__abc_52155_new_n21156_; 
wire u2__abc_52155_new_n21157_; 
wire u2__abc_52155_new_n21158_; 
wire u2__abc_52155_new_n21159_; 
wire u2__abc_52155_new_n21160_; 
wire u2__abc_52155_new_n21161_; 
wire u2__abc_52155_new_n21162_; 
wire u2__abc_52155_new_n21163_; 
wire u2__abc_52155_new_n21164_; 
wire u2__abc_52155_new_n21165_; 
wire u2__abc_52155_new_n21166_; 
wire u2__abc_52155_new_n21168_; 
wire u2__abc_52155_new_n21169_; 
wire u2__abc_52155_new_n21170_; 
wire u2__abc_52155_new_n21171_; 
wire u2__abc_52155_new_n21172_; 
wire u2__abc_52155_new_n21173_; 
wire u2__abc_52155_new_n21174_; 
wire u2__abc_52155_new_n21175_; 
wire u2__abc_52155_new_n21176_; 
wire u2__abc_52155_new_n21177_; 
wire u2__abc_52155_new_n21178_; 
wire u2__abc_52155_new_n21180_; 
wire u2__abc_52155_new_n21181_; 
wire u2__abc_52155_new_n21182_; 
wire u2__abc_52155_new_n21183_; 
wire u2__abc_52155_new_n21184_; 
wire u2__abc_52155_new_n21185_; 
wire u2__abc_52155_new_n21186_; 
wire u2__abc_52155_new_n21187_; 
wire u2__abc_52155_new_n21188_; 
wire u2__abc_52155_new_n21189_; 
wire u2__abc_52155_new_n21190_; 
wire u2__abc_52155_new_n21192_; 
wire u2__abc_52155_new_n21193_; 
wire u2__abc_52155_new_n21194_; 
wire u2__abc_52155_new_n21195_; 
wire u2__abc_52155_new_n21196_; 
wire u2__abc_52155_new_n21197_; 
wire u2__abc_52155_new_n21198_; 
wire u2__abc_52155_new_n21199_; 
wire u2__abc_52155_new_n21200_; 
wire u2__abc_52155_new_n21201_; 
wire u2__abc_52155_new_n21202_; 
wire u2__abc_52155_new_n21204_; 
wire u2__abc_52155_new_n21205_; 
wire u2__abc_52155_new_n21206_; 
wire u2__abc_52155_new_n21207_; 
wire u2__abc_52155_new_n21208_; 
wire u2__abc_52155_new_n21209_; 
wire u2__abc_52155_new_n21210_; 
wire u2__abc_52155_new_n21211_; 
wire u2__abc_52155_new_n21212_; 
wire u2__abc_52155_new_n21213_; 
wire u2__abc_52155_new_n21214_; 
wire u2__abc_52155_new_n21216_; 
wire u2__abc_52155_new_n21217_; 
wire u2__abc_52155_new_n21218_; 
wire u2__abc_52155_new_n21219_; 
wire u2__abc_52155_new_n21220_; 
wire u2__abc_52155_new_n21221_; 
wire u2__abc_52155_new_n21222_; 
wire u2__abc_52155_new_n21223_; 
wire u2__abc_52155_new_n21224_; 
wire u2__abc_52155_new_n21225_; 
wire u2__abc_52155_new_n21226_; 
wire u2__abc_52155_new_n21228_; 
wire u2__abc_52155_new_n21229_; 
wire u2__abc_52155_new_n21230_; 
wire u2__abc_52155_new_n21231_; 
wire u2__abc_52155_new_n21232_; 
wire u2__abc_52155_new_n21233_; 
wire u2__abc_52155_new_n21234_; 
wire u2__abc_52155_new_n21235_; 
wire u2__abc_52155_new_n21236_; 
wire u2__abc_52155_new_n21237_; 
wire u2__abc_52155_new_n21238_; 
wire u2__abc_52155_new_n21240_; 
wire u2__abc_52155_new_n21241_; 
wire u2__abc_52155_new_n21242_; 
wire u2__abc_52155_new_n21243_; 
wire u2__abc_52155_new_n21244_; 
wire u2__abc_52155_new_n21245_; 
wire u2__abc_52155_new_n21246_; 
wire u2__abc_52155_new_n21247_; 
wire u2__abc_52155_new_n21248_; 
wire u2__abc_52155_new_n21249_; 
wire u2__abc_52155_new_n21250_; 
wire u2__abc_52155_new_n21252_; 
wire u2__abc_52155_new_n21253_; 
wire u2__abc_52155_new_n21254_; 
wire u2__abc_52155_new_n21255_; 
wire u2__abc_52155_new_n21256_; 
wire u2__abc_52155_new_n21257_; 
wire u2__abc_52155_new_n21258_; 
wire u2__abc_52155_new_n21259_; 
wire u2__abc_52155_new_n21260_; 
wire u2__abc_52155_new_n21261_; 
wire u2__abc_52155_new_n21262_; 
wire u2__abc_52155_new_n21264_; 
wire u2__abc_52155_new_n21265_; 
wire u2__abc_52155_new_n21266_; 
wire u2__abc_52155_new_n21267_; 
wire u2__abc_52155_new_n21268_; 
wire u2__abc_52155_new_n21269_; 
wire u2__abc_52155_new_n21270_; 
wire u2__abc_52155_new_n21271_; 
wire u2__abc_52155_new_n21272_; 
wire u2__abc_52155_new_n21273_; 
wire u2__abc_52155_new_n21274_; 
wire u2__abc_52155_new_n21276_; 
wire u2__abc_52155_new_n21277_; 
wire u2__abc_52155_new_n21278_; 
wire u2__abc_52155_new_n21279_; 
wire u2__abc_52155_new_n21280_; 
wire u2__abc_52155_new_n21281_; 
wire u2__abc_52155_new_n21282_; 
wire u2__abc_52155_new_n21283_; 
wire u2__abc_52155_new_n21284_; 
wire u2__abc_52155_new_n21285_; 
wire u2__abc_52155_new_n21286_; 
wire u2__abc_52155_new_n21288_; 
wire u2__abc_52155_new_n21289_; 
wire u2__abc_52155_new_n21290_; 
wire u2__abc_52155_new_n21291_; 
wire u2__abc_52155_new_n21292_; 
wire u2__abc_52155_new_n21293_; 
wire u2__abc_52155_new_n21294_; 
wire u2__abc_52155_new_n21295_; 
wire u2__abc_52155_new_n21296_; 
wire u2__abc_52155_new_n21297_; 
wire u2__abc_52155_new_n21298_; 
wire u2__abc_52155_new_n21300_; 
wire u2__abc_52155_new_n21301_; 
wire u2__abc_52155_new_n21302_; 
wire u2__abc_52155_new_n21303_; 
wire u2__abc_52155_new_n21304_; 
wire u2__abc_52155_new_n21305_; 
wire u2__abc_52155_new_n21306_; 
wire u2__abc_52155_new_n21307_; 
wire u2__abc_52155_new_n21308_; 
wire u2__abc_52155_new_n21309_; 
wire u2__abc_52155_new_n21310_; 
wire u2__abc_52155_new_n21312_; 
wire u2__abc_52155_new_n21313_; 
wire u2__abc_52155_new_n21314_; 
wire u2__abc_52155_new_n21315_; 
wire u2__abc_52155_new_n21316_; 
wire u2__abc_52155_new_n21317_; 
wire u2__abc_52155_new_n21318_; 
wire u2__abc_52155_new_n21319_; 
wire u2__abc_52155_new_n21320_; 
wire u2__abc_52155_new_n21321_; 
wire u2__abc_52155_new_n21322_; 
wire u2__abc_52155_new_n21324_; 
wire u2__abc_52155_new_n21325_; 
wire u2__abc_52155_new_n21326_; 
wire u2__abc_52155_new_n21327_; 
wire u2__abc_52155_new_n21328_; 
wire u2__abc_52155_new_n21329_; 
wire u2__abc_52155_new_n21330_; 
wire u2__abc_52155_new_n21331_; 
wire u2__abc_52155_new_n21332_; 
wire u2__abc_52155_new_n21333_; 
wire u2__abc_52155_new_n21334_; 
wire u2__abc_52155_new_n21336_; 
wire u2__abc_52155_new_n21337_; 
wire u2__abc_52155_new_n21338_; 
wire u2__abc_52155_new_n21339_; 
wire u2__abc_52155_new_n21340_; 
wire u2__abc_52155_new_n21341_; 
wire u2__abc_52155_new_n21342_; 
wire u2__abc_52155_new_n21343_; 
wire u2__abc_52155_new_n21344_; 
wire u2__abc_52155_new_n21345_; 
wire u2__abc_52155_new_n21346_; 
wire u2__abc_52155_new_n21348_; 
wire u2__abc_52155_new_n21349_; 
wire u2__abc_52155_new_n21350_; 
wire u2__abc_52155_new_n21351_; 
wire u2__abc_52155_new_n21352_; 
wire u2__abc_52155_new_n21353_; 
wire u2__abc_52155_new_n21354_; 
wire u2__abc_52155_new_n21355_; 
wire u2__abc_52155_new_n21356_; 
wire u2__abc_52155_new_n21357_; 
wire u2__abc_52155_new_n21358_; 
wire u2__abc_52155_new_n21360_; 
wire u2__abc_52155_new_n21361_; 
wire u2__abc_52155_new_n21362_; 
wire u2__abc_52155_new_n21363_; 
wire u2__abc_52155_new_n21364_; 
wire u2__abc_52155_new_n21365_; 
wire u2__abc_52155_new_n21366_; 
wire u2__abc_52155_new_n21367_; 
wire u2__abc_52155_new_n21368_; 
wire u2__abc_52155_new_n21369_; 
wire u2__abc_52155_new_n21370_; 
wire u2__abc_52155_new_n21372_; 
wire u2__abc_52155_new_n21373_; 
wire u2__abc_52155_new_n21374_; 
wire u2__abc_52155_new_n21375_; 
wire u2__abc_52155_new_n21376_; 
wire u2__abc_52155_new_n21377_; 
wire u2__abc_52155_new_n21378_; 
wire u2__abc_52155_new_n21379_; 
wire u2__abc_52155_new_n21380_; 
wire u2__abc_52155_new_n21381_; 
wire u2__abc_52155_new_n21382_; 
wire u2__abc_52155_new_n21384_; 
wire u2__abc_52155_new_n21385_; 
wire u2__abc_52155_new_n21386_; 
wire u2__abc_52155_new_n21387_; 
wire u2__abc_52155_new_n21388_; 
wire u2__abc_52155_new_n21389_; 
wire u2__abc_52155_new_n21390_; 
wire u2__abc_52155_new_n21391_; 
wire u2__abc_52155_new_n21392_; 
wire u2__abc_52155_new_n21393_; 
wire u2__abc_52155_new_n21394_; 
wire u2__abc_52155_new_n21396_; 
wire u2__abc_52155_new_n21397_; 
wire u2__abc_52155_new_n21398_; 
wire u2__abc_52155_new_n21399_; 
wire u2__abc_52155_new_n21400_; 
wire u2__abc_52155_new_n21401_; 
wire u2__abc_52155_new_n21402_; 
wire u2__abc_52155_new_n21403_; 
wire u2__abc_52155_new_n21404_; 
wire u2__abc_52155_new_n21405_; 
wire u2__abc_52155_new_n21406_; 
wire u2__abc_52155_new_n21408_; 
wire u2__abc_52155_new_n21409_; 
wire u2__abc_52155_new_n21410_; 
wire u2__abc_52155_new_n21411_; 
wire u2__abc_52155_new_n21412_; 
wire u2__abc_52155_new_n21413_; 
wire u2__abc_52155_new_n21414_; 
wire u2__abc_52155_new_n21415_; 
wire u2__abc_52155_new_n21416_; 
wire u2__abc_52155_new_n21417_; 
wire u2__abc_52155_new_n21418_; 
wire u2__abc_52155_new_n21420_; 
wire u2__abc_52155_new_n21421_; 
wire u2__abc_52155_new_n21422_; 
wire u2__abc_52155_new_n21423_; 
wire u2__abc_52155_new_n21424_; 
wire u2__abc_52155_new_n21425_; 
wire u2__abc_52155_new_n21426_; 
wire u2__abc_52155_new_n21427_; 
wire u2__abc_52155_new_n21428_; 
wire u2__abc_52155_new_n21429_; 
wire u2__abc_52155_new_n21430_; 
wire u2__abc_52155_new_n21432_; 
wire u2__abc_52155_new_n21433_; 
wire u2__abc_52155_new_n21434_; 
wire u2__abc_52155_new_n21435_; 
wire u2__abc_52155_new_n21436_; 
wire u2__abc_52155_new_n21437_; 
wire u2__abc_52155_new_n21438_; 
wire u2__abc_52155_new_n21439_; 
wire u2__abc_52155_new_n21440_; 
wire u2__abc_52155_new_n21441_; 
wire u2__abc_52155_new_n21442_; 
wire u2__abc_52155_new_n21444_; 
wire u2__abc_52155_new_n21445_; 
wire u2__abc_52155_new_n21446_; 
wire u2__abc_52155_new_n21447_; 
wire u2__abc_52155_new_n21448_; 
wire u2__abc_52155_new_n21449_; 
wire u2__abc_52155_new_n21450_; 
wire u2__abc_52155_new_n21451_; 
wire u2__abc_52155_new_n21452_; 
wire u2__abc_52155_new_n21453_; 
wire u2__abc_52155_new_n21454_; 
wire u2__abc_52155_new_n21456_; 
wire u2__abc_52155_new_n21457_; 
wire u2__abc_52155_new_n21458_; 
wire u2__abc_52155_new_n21459_; 
wire u2__abc_52155_new_n21460_; 
wire u2__abc_52155_new_n21461_; 
wire u2__abc_52155_new_n21462_; 
wire u2__abc_52155_new_n21463_; 
wire u2__abc_52155_new_n21464_; 
wire u2__abc_52155_new_n21465_; 
wire u2__abc_52155_new_n21466_; 
wire u2__abc_52155_new_n21468_; 
wire u2__abc_52155_new_n21469_; 
wire u2__abc_52155_new_n21470_; 
wire u2__abc_52155_new_n21471_; 
wire u2__abc_52155_new_n21472_; 
wire u2__abc_52155_new_n21473_; 
wire u2__abc_52155_new_n21474_; 
wire u2__abc_52155_new_n21475_; 
wire u2__abc_52155_new_n21476_; 
wire u2__abc_52155_new_n21477_; 
wire u2__abc_52155_new_n21478_; 
wire u2__abc_52155_new_n21480_; 
wire u2__abc_52155_new_n21481_; 
wire u2__abc_52155_new_n21482_; 
wire u2__abc_52155_new_n21483_; 
wire u2__abc_52155_new_n21484_; 
wire u2__abc_52155_new_n21485_; 
wire u2__abc_52155_new_n21486_; 
wire u2__abc_52155_new_n21487_; 
wire u2__abc_52155_new_n21488_; 
wire u2__abc_52155_new_n21489_; 
wire u2__abc_52155_new_n21490_; 
wire u2__abc_52155_new_n21492_; 
wire u2__abc_52155_new_n21493_; 
wire u2__abc_52155_new_n21494_; 
wire u2__abc_52155_new_n21495_; 
wire u2__abc_52155_new_n21496_; 
wire u2__abc_52155_new_n21497_; 
wire u2__abc_52155_new_n21498_; 
wire u2__abc_52155_new_n21499_; 
wire u2__abc_52155_new_n21500_; 
wire u2__abc_52155_new_n21501_; 
wire u2__abc_52155_new_n21502_; 
wire u2__abc_52155_new_n21504_; 
wire u2__abc_52155_new_n21505_; 
wire u2__abc_52155_new_n21506_; 
wire u2__abc_52155_new_n21507_; 
wire u2__abc_52155_new_n21508_; 
wire u2__abc_52155_new_n21509_; 
wire u2__abc_52155_new_n21510_; 
wire u2__abc_52155_new_n21511_; 
wire u2__abc_52155_new_n21512_; 
wire u2__abc_52155_new_n21513_; 
wire u2__abc_52155_new_n21514_; 
wire u2__abc_52155_new_n21516_; 
wire u2__abc_52155_new_n21517_; 
wire u2__abc_52155_new_n21518_; 
wire u2__abc_52155_new_n21519_; 
wire u2__abc_52155_new_n21520_; 
wire u2__abc_52155_new_n21521_; 
wire u2__abc_52155_new_n21522_; 
wire u2__abc_52155_new_n21523_; 
wire u2__abc_52155_new_n21524_; 
wire u2__abc_52155_new_n21525_; 
wire u2__abc_52155_new_n21526_; 
wire u2__abc_52155_new_n21528_; 
wire u2__abc_52155_new_n21529_; 
wire u2__abc_52155_new_n21530_; 
wire u2__abc_52155_new_n21531_; 
wire u2__abc_52155_new_n21532_; 
wire u2__abc_52155_new_n21533_; 
wire u2__abc_52155_new_n21534_; 
wire u2__abc_52155_new_n21535_; 
wire u2__abc_52155_new_n21536_; 
wire u2__abc_52155_new_n21537_; 
wire u2__abc_52155_new_n21538_; 
wire u2__abc_52155_new_n21540_; 
wire u2__abc_52155_new_n21541_; 
wire u2__abc_52155_new_n21542_; 
wire u2__abc_52155_new_n21543_; 
wire u2__abc_52155_new_n21544_; 
wire u2__abc_52155_new_n21545_; 
wire u2__abc_52155_new_n21546_; 
wire u2__abc_52155_new_n21547_; 
wire u2__abc_52155_new_n21548_; 
wire u2__abc_52155_new_n21549_; 
wire u2__abc_52155_new_n21550_; 
wire u2__abc_52155_new_n21552_; 
wire u2__abc_52155_new_n21553_; 
wire u2__abc_52155_new_n21554_; 
wire u2__abc_52155_new_n21555_; 
wire u2__abc_52155_new_n21556_; 
wire u2__abc_52155_new_n21557_; 
wire u2__abc_52155_new_n21558_; 
wire u2__abc_52155_new_n21559_; 
wire u2__abc_52155_new_n21560_; 
wire u2__abc_52155_new_n21561_; 
wire u2__abc_52155_new_n21562_; 
wire u2__abc_52155_new_n21564_; 
wire u2__abc_52155_new_n21565_; 
wire u2__abc_52155_new_n21566_; 
wire u2__abc_52155_new_n21567_; 
wire u2__abc_52155_new_n21568_; 
wire u2__abc_52155_new_n21569_; 
wire u2__abc_52155_new_n21570_; 
wire u2__abc_52155_new_n21571_; 
wire u2__abc_52155_new_n21572_; 
wire u2__abc_52155_new_n21573_; 
wire u2__abc_52155_new_n21574_; 
wire u2__abc_52155_new_n21576_; 
wire u2__abc_52155_new_n21577_; 
wire u2__abc_52155_new_n21578_; 
wire u2__abc_52155_new_n21579_; 
wire u2__abc_52155_new_n21580_; 
wire u2__abc_52155_new_n21581_; 
wire u2__abc_52155_new_n21582_; 
wire u2__abc_52155_new_n21583_; 
wire u2__abc_52155_new_n21584_; 
wire u2__abc_52155_new_n21585_; 
wire u2__abc_52155_new_n21586_; 
wire u2__abc_52155_new_n21588_; 
wire u2__abc_52155_new_n21589_; 
wire u2__abc_52155_new_n21590_; 
wire u2__abc_52155_new_n21591_; 
wire u2__abc_52155_new_n21592_; 
wire u2__abc_52155_new_n21593_; 
wire u2__abc_52155_new_n21594_; 
wire u2__abc_52155_new_n21595_; 
wire u2__abc_52155_new_n21596_; 
wire u2__abc_52155_new_n21597_; 
wire u2__abc_52155_new_n21598_; 
wire u2__abc_52155_new_n21600_; 
wire u2__abc_52155_new_n21601_; 
wire u2__abc_52155_new_n21602_; 
wire u2__abc_52155_new_n21603_; 
wire u2__abc_52155_new_n21604_; 
wire u2__abc_52155_new_n21605_; 
wire u2__abc_52155_new_n21606_; 
wire u2__abc_52155_new_n21607_; 
wire u2__abc_52155_new_n21608_; 
wire u2__abc_52155_new_n21609_; 
wire u2__abc_52155_new_n21610_; 
wire u2__abc_52155_new_n21612_; 
wire u2__abc_52155_new_n21613_; 
wire u2__abc_52155_new_n21614_; 
wire u2__abc_52155_new_n21615_; 
wire u2__abc_52155_new_n21616_; 
wire u2__abc_52155_new_n21617_; 
wire u2__abc_52155_new_n21618_; 
wire u2__abc_52155_new_n21619_; 
wire u2__abc_52155_new_n21620_; 
wire u2__abc_52155_new_n21621_; 
wire u2__abc_52155_new_n21622_; 
wire u2__abc_52155_new_n21624_; 
wire u2__abc_52155_new_n21625_; 
wire u2__abc_52155_new_n21626_; 
wire u2__abc_52155_new_n21627_; 
wire u2__abc_52155_new_n21628_; 
wire u2__abc_52155_new_n21629_; 
wire u2__abc_52155_new_n21630_; 
wire u2__abc_52155_new_n21631_; 
wire u2__abc_52155_new_n21632_; 
wire u2__abc_52155_new_n21633_; 
wire u2__abc_52155_new_n21634_; 
wire u2__abc_52155_new_n21636_; 
wire u2__abc_52155_new_n21637_; 
wire u2__abc_52155_new_n21638_; 
wire u2__abc_52155_new_n21639_; 
wire u2__abc_52155_new_n21640_; 
wire u2__abc_52155_new_n21641_; 
wire u2__abc_52155_new_n21642_; 
wire u2__abc_52155_new_n21643_; 
wire u2__abc_52155_new_n21644_; 
wire u2__abc_52155_new_n21645_; 
wire u2__abc_52155_new_n21646_; 
wire u2__abc_52155_new_n21648_; 
wire u2__abc_52155_new_n21649_; 
wire u2__abc_52155_new_n21650_; 
wire u2__abc_52155_new_n21651_; 
wire u2__abc_52155_new_n21652_; 
wire u2__abc_52155_new_n21653_; 
wire u2__abc_52155_new_n21654_; 
wire u2__abc_52155_new_n21655_; 
wire u2__abc_52155_new_n21656_; 
wire u2__abc_52155_new_n21657_; 
wire u2__abc_52155_new_n21658_; 
wire u2__abc_52155_new_n21660_; 
wire u2__abc_52155_new_n21661_; 
wire u2__abc_52155_new_n21662_; 
wire u2__abc_52155_new_n21663_; 
wire u2__abc_52155_new_n21664_; 
wire u2__abc_52155_new_n21665_; 
wire u2__abc_52155_new_n21666_; 
wire u2__abc_52155_new_n21667_; 
wire u2__abc_52155_new_n21668_; 
wire u2__abc_52155_new_n21669_; 
wire u2__abc_52155_new_n21670_; 
wire u2__abc_52155_new_n21672_; 
wire u2__abc_52155_new_n21673_; 
wire u2__abc_52155_new_n21674_; 
wire u2__abc_52155_new_n21675_; 
wire u2__abc_52155_new_n21676_; 
wire u2__abc_52155_new_n21677_; 
wire u2__abc_52155_new_n21678_; 
wire u2__abc_52155_new_n21679_; 
wire u2__abc_52155_new_n21680_; 
wire u2__abc_52155_new_n21681_; 
wire u2__abc_52155_new_n21682_; 
wire u2__abc_52155_new_n21684_; 
wire u2__abc_52155_new_n21685_; 
wire u2__abc_52155_new_n21686_; 
wire u2__abc_52155_new_n21687_; 
wire u2__abc_52155_new_n21688_; 
wire u2__abc_52155_new_n21689_; 
wire u2__abc_52155_new_n21690_; 
wire u2__abc_52155_new_n21691_; 
wire u2__abc_52155_new_n21692_; 
wire u2__abc_52155_new_n21693_; 
wire u2__abc_52155_new_n21694_; 
wire u2__abc_52155_new_n21696_; 
wire u2__abc_52155_new_n21697_; 
wire u2__abc_52155_new_n21698_; 
wire u2__abc_52155_new_n21699_; 
wire u2__abc_52155_new_n21700_; 
wire u2__abc_52155_new_n21701_; 
wire u2__abc_52155_new_n21702_; 
wire u2__abc_52155_new_n21703_; 
wire u2__abc_52155_new_n21704_; 
wire u2__abc_52155_new_n21705_; 
wire u2__abc_52155_new_n21706_; 
wire u2__abc_52155_new_n21708_; 
wire u2__abc_52155_new_n21709_; 
wire u2__abc_52155_new_n21710_; 
wire u2__abc_52155_new_n21711_; 
wire u2__abc_52155_new_n21712_; 
wire u2__abc_52155_new_n21713_; 
wire u2__abc_52155_new_n21714_; 
wire u2__abc_52155_new_n21715_; 
wire u2__abc_52155_new_n21716_; 
wire u2__abc_52155_new_n21717_; 
wire u2__abc_52155_new_n21718_; 
wire u2__abc_52155_new_n21720_; 
wire u2__abc_52155_new_n21721_; 
wire u2__abc_52155_new_n21722_; 
wire u2__abc_52155_new_n21723_; 
wire u2__abc_52155_new_n21724_; 
wire u2__abc_52155_new_n21725_; 
wire u2__abc_52155_new_n21726_; 
wire u2__abc_52155_new_n21727_; 
wire u2__abc_52155_new_n21728_; 
wire u2__abc_52155_new_n21729_; 
wire u2__abc_52155_new_n21730_; 
wire u2__abc_52155_new_n21732_; 
wire u2__abc_52155_new_n21733_; 
wire u2__abc_52155_new_n21734_; 
wire u2__abc_52155_new_n21735_; 
wire u2__abc_52155_new_n21736_; 
wire u2__abc_52155_new_n21737_; 
wire u2__abc_52155_new_n21738_; 
wire u2__abc_52155_new_n21739_; 
wire u2__abc_52155_new_n21740_; 
wire u2__abc_52155_new_n21741_; 
wire u2__abc_52155_new_n21742_; 
wire u2__abc_52155_new_n21744_; 
wire u2__abc_52155_new_n21745_; 
wire u2__abc_52155_new_n21746_; 
wire u2__abc_52155_new_n21747_; 
wire u2__abc_52155_new_n21748_; 
wire u2__abc_52155_new_n21749_; 
wire u2__abc_52155_new_n21750_; 
wire u2__abc_52155_new_n21751_; 
wire u2__abc_52155_new_n21752_; 
wire u2__abc_52155_new_n21753_; 
wire u2__abc_52155_new_n21754_; 
wire u2__abc_52155_new_n21756_; 
wire u2__abc_52155_new_n21757_; 
wire u2__abc_52155_new_n21758_; 
wire u2__abc_52155_new_n21759_; 
wire u2__abc_52155_new_n21760_; 
wire u2__abc_52155_new_n21761_; 
wire u2__abc_52155_new_n21762_; 
wire u2__abc_52155_new_n21763_; 
wire u2__abc_52155_new_n21764_; 
wire u2__abc_52155_new_n21765_; 
wire u2__abc_52155_new_n21766_; 
wire u2__abc_52155_new_n21768_; 
wire u2__abc_52155_new_n21769_; 
wire u2__abc_52155_new_n21770_; 
wire u2__abc_52155_new_n21771_; 
wire u2__abc_52155_new_n21772_; 
wire u2__abc_52155_new_n21773_; 
wire u2__abc_52155_new_n21774_; 
wire u2__abc_52155_new_n21775_; 
wire u2__abc_52155_new_n21776_; 
wire u2__abc_52155_new_n21777_; 
wire u2__abc_52155_new_n21778_; 
wire u2__abc_52155_new_n21780_; 
wire u2__abc_52155_new_n21781_; 
wire u2__abc_52155_new_n21782_; 
wire u2__abc_52155_new_n21783_; 
wire u2__abc_52155_new_n21784_; 
wire u2__abc_52155_new_n21785_; 
wire u2__abc_52155_new_n21786_; 
wire u2__abc_52155_new_n21787_; 
wire u2__abc_52155_new_n21788_; 
wire u2__abc_52155_new_n21789_; 
wire u2__abc_52155_new_n21790_; 
wire u2__abc_52155_new_n21792_; 
wire u2__abc_52155_new_n21793_; 
wire u2__abc_52155_new_n21794_; 
wire u2__abc_52155_new_n21795_; 
wire u2__abc_52155_new_n21796_; 
wire u2__abc_52155_new_n21797_; 
wire u2__abc_52155_new_n21798_; 
wire u2__abc_52155_new_n21799_; 
wire u2__abc_52155_new_n21800_; 
wire u2__abc_52155_new_n21801_; 
wire u2__abc_52155_new_n21802_; 
wire u2__abc_52155_new_n21804_; 
wire u2__abc_52155_new_n21805_; 
wire u2__abc_52155_new_n21806_; 
wire u2__abc_52155_new_n21807_; 
wire u2__abc_52155_new_n21808_; 
wire u2__abc_52155_new_n21809_; 
wire u2__abc_52155_new_n21810_; 
wire u2__abc_52155_new_n21811_; 
wire u2__abc_52155_new_n21812_; 
wire u2__abc_52155_new_n21813_; 
wire u2__abc_52155_new_n21814_; 
wire u2__abc_52155_new_n21816_; 
wire u2__abc_52155_new_n21817_; 
wire u2__abc_52155_new_n21818_; 
wire u2__abc_52155_new_n21819_; 
wire u2__abc_52155_new_n21820_; 
wire u2__abc_52155_new_n21821_; 
wire u2__abc_52155_new_n21822_; 
wire u2__abc_52155_new_n21823_; 
wire u2__abc_52155_new_n21824_; 
wire u2__abc_52155_new_n21825_; 
wire u2__abc_52155_new_n21826_; 
wire u2__abc_52155_new_n21828_; 
wire u2__abc_52155_new_n21829_; 
wire u2__abc_52155_new_n21830_; 
wire u2__abc_52155_new_n21831_; 
wire u2__abc_52155_new_n21832_; 
wire u2__abc_52155_new_n21833_; 
wire u2__abc_52155_new_n21834_; 
wire u2__abc_52155_new_n21835_; 
wire u2__abc_52155_new_n21836_; 
wire u2__abc_52155_new_n21837_; 
wire u2__abc_52155_new_n21838_; 
wire u2__abc_52155_new_n21840_; 
wire u2__abc_52155_new_n21841_; 
wire u2__abc_52155_new_n21842_; 
wire u2__abc_52155_new_n21843_; 
wire u2__abc_52155_new_n21844_; 
wire u2__abc_52155_new_n21845_; 
wire u2__abc_52155_new_n21846_; 
wire u2__abc_52155_new_n21847_; 
wire u2__abc_52155_new_n21848_; 
wire u2__abc_52155_new_n21849_; 
wire u2__abc_52155_new_n21850_; 
wire u2__abc_52155_new_n21852_; 
wire u2__abc_52155_new_n21853_; 
wire u2__abc_52155_new_n21854_; 
wire u2__abc_52155_new_n21855_; 
wire u2__abc_52155_new_n21856_; 
wire u2__abc_52155_new_n21857_; 
wire u2__abc_52155_new_n21858_; 
wire u2__abc_52155_new_n21859_; 
wire u2__abc_52155_new_n21860_; 
wire u2__abc_52155_new_n21861_; 
wire u2__abc_52155_new_n21862_; 
wire u2__abc_52155_new_n21864_; 
wire u2__abc_52155_new_n21865_; 
wire u2__abc_52155_new_n21866_; 
wire u2__abc_52155_new_n21867_; 
wire u2__abc_52155_new_n21868_; 
wire u2__abc_52155_new_n21869_; 
wire u2__abc_52155_new_n21870_; 
wire u2__abc_52155_new_n21871_; 
wire u2__abc_52155_new_n21872_; 
wire u2__abc_52155_new_n21873_; 
wire u2__abc_52155_new_n21874_; 
wire u2__abc_52155_new_n21876_; 
wire u2__abc_52155_new_n21877_; 
wire u2__abc_52155_new_n21878_; 
wire u2__abc_52155_new_n21879_; 
wire u2__abc_52155_new_n21880_; 
wire u2__abc_52155_new_n21881_; 
wire u2__abc_52155_new_n21882_; 
wire u2__abc_52155_new_n21883_; 
wire u2__abc_52155_new_n21884_; 
wire u2__abc_52155_new_n21885_; 
wire u2__abc_52155_new_n21886_; 
wire u2__abc_52155_new_n21888_; 
wire u2__abc_52155_new_n21889_; 
wire u2__abc_52155_new_n21890_; 
wire u2__abc_52155_new_n21891_; 
wire u2__abc_52155_new_n21892_; 
wire u2__abc_52155_new_n21893_; 
wire u2__abc_52155_new_n21894_; 
wire u2__abc_52155_new_n21895_; 
wire u2__abc_52155_new_n21896_; 
wire u2__abc_52155_new_n21897_; 
wire u2__abc_52155_new_n21898_; 
wire u2__abc_52155_new_n21900_; 
wire u2__abc_52155_new_n21901_; 
wire u2__abc_52155_new_n21902_; 
wire u2__abc_52155_new_n21903_; 
wire u2__abc_52155_new_n21904_; 
wire u2__abc_52155_new_n21905_; 
wire u2__abc_52155_new_n21906_; 
wire u2__abc_52155_new_n21907_; 
wire u2__abc_52155_new_n21908_; 
wire u2__abc_52155_new_n21909_; 
wire u2__abc_52155_new_n21910_; 
wire u2__abc_52155_new_n21912_; 
wire u2__abc_52155_new_n21913_; 
wire u2__abc_52155_new_n21914_; 
wire u2__abc_52155_new_n21915_; 
wire u2__abc_52155_new_n21916_; 
wire u2__abc_52155_new_n21917_; 
wire u2__abc_52155_new_n21918_; 
wire u2__abc_52155_new_n21919_; 
wire u2__abc_52155_new_n21920_; 
wire u2__abc_52155_new_n21921_; 
wire u2__abc_52155_new_n21922_; 
wire u2__abc_52155_new_n21924_; 
wire u2__abc_52155_new_n21925_; 
wire u2__abc_52155_new_n21926_; 
wire u2__abc_52155_new_n21927_; 
wire u2__abc_52155_new_n21928_; 
wire u2__abc_52155_new_n21929_; 
wire u2__abc_52155_new_n21930_; 
wire u2__abc_52155_new_n21931_; 
wire u2__abc_52155_new_n21932_; 
wire u2__abc_52155_new_n21933_; 
wire u2__abc_52155_new_n21934_; 
wire u2__abc_52155_new_n21936_; 
wire u2__abc_52155_new_n21937_; 
wire u2__abc_52155_new_n21938_; 
wire u2__abc_52155_new_n21939_; 
wire u2__abc_52155_new_n21940_; 
wire u2__abc_52155_new_n21941_; 
wire u2__abc_52155_new_n21942_; 
wire u2__abc_52155_new_n21943_; 
wire u2__abc_52155_new_n21944_; 
wire u2__abc_52155_new_n21945_; 
wire u2__abc_52155_new_n21946_; 
wire u2__abc_52155_new_n21948_; 
wire u2__abc_52155_new_n21949_; 
wire u2__abc_52155_new_n21950_; 
wire u2__abc_52155_new_n21951_; 
wire u2__abc_52155_new_n21952_; 
wire u2__abc_52155_new_n21953_; 
wire u2__abc_52155_new_n21954_; 
wire u2__abc_52155_new_n21955_; 
wire u2__abc_52155_new_n21956_; 
wire u2__abc_52155_new_n21957_; 
wire u2__abc_52155_new_n21958_; 
wire u2__abc_52155_new_n21960_; 
wire u2__abc_52155_new_n21961_; 
wire u2__abc_52155_new_n21962_; 
wire u2__abc_52155_new_n21963_; 
wire u2__abc_52155_new_n21964_; 
wire u2__abc_52155_new_n21965_; 
wire u2__abc_52155_new_n21966_; 
wire u2__abc_52155_new_n21967_; 
wire u2__abc_52155_new_n21968_; 
wire u2__abc_52155_new_n21969_; 
wire u2__abc_52155_new_n21970_; 
wire u2__abc_52155_new_n21972_; 
wire u2__abc_52155_new_n21973_; 
wire u2__abc_52155_new_n21974_; 
wire u2__abc_52155_new_n21975_; 
wire u2__abc_52155_new_n21976_; 
wire u2__abc_52155_new_n21977_; 
wire u2__abc_52155_new_n21978_; 
wire u2__abc_52155_new_n21979_; 
wire u2__abc_52155_new_n21980_; 
wire u2__abc_52155_new_n21981_; 
wire u2__abc_52155_new_n21982_; 
wire u2__abc_52155_new_n21984_; 
wire u2__abc_52155_new_n21985_; 
wire u2__abc_52155_new_n21986_; 
wire u2__abc_52155_new_n21987_; 
wire u2__abc_52155_new_n21988_; 
wire u2__abc_52155_new_n21989_; 
wire u2__abc_52155_new_n21990_; 
wire u2__abc_52155_new_n21991_; 
wire u2__abc_52155_new_n21992_; 
wire u2__abc_52155_new_n21993_; 
wire u2__abc_52155_new_n21994_; 
wire u2__abc_52155_new_n21996_; 
wire u2__abc_52155_new_n21997_; 
wire u2__abc_52155_new_n21998_; 
wire u2__abc_52155_new_n21999_; 
wire u2__abc_52155_new_n22000_; 
wire u2__abc_52155_new_n22001_; 
wire u2__abc_52155_new_n22002_; 
wire u2__abc_52155_new_n22003_; 
wire u2__abc_52155_new_n22004_; 
wire u2__abc_52155_new_n22005_; 
wire u2__abc_52155_new_n22006_; 
wire u2__abc_52155_new_n22008_; 
wire u2__abc_52155_new_n22009_; 
wire u2__abc_52155_new_n22010_; 
wire u2__abc_52155_new_n22011_; 
wire u2__abc_52155_new_n22012_; 
wire u2__abc_52155_new_n22013_; 
wire u2__abc_52155_new_n22014_; 
wire u2__abc_52155_new_n22015_; 
wire u2__abc_52155_new_n22016_; 
wire u2__abc_52155_new_n22017_; 
wire u2__abc_52155_new_n22018_; 
wire u2__abc_52155_new_n22020_; 
wire u2__abc_52155_new_n22021_; 
wire u2__abc_52155_new_n22022_; 
wire u2__abc_52155_new_n22023_; 
wire u2__abc_52155_new_n22024_; 
wire u2__abc_52155_new_n22025_; 
wire u2__abc_52155_new_n22026_; 
wire u2__abc_52155_new_n22027_; 
wire u2__abc_52155_new_n22028_; 
wire u2__abc_52155_new_n22029_; 
wire u2__abc_52155_new_n22030_; 
wire u2__abc_52155_new_n22032_; 
wire u2__abc_52155_new_n22033_; 
wire u2__abc_52155_new_n22034_; 
wire u2__abc_52155_new_n22035_; 
wire u2__abc_52155_new_n22036_; 
wire u2__abc_52155_new_n22037_; 
wire u2__abc_52155_new_n22038_; 
wire u2__abc_52155_new_n22039_; 
wire u2__abc_52155_new_n22040_; 
wire u2__abc_52155_new_n22041_; 
wire u2__abc_52155_new_n22042_; 
wire u2__abc_52155_new_n22044_; 
wire u2__abc_52155_new_n22045_; 
wire u2__abc_52155_new_n22046_; 
wire u2__abc_52155_new_n22047_; 
wire u2__abc_52155_new_n22048_; 
wire u2__abc_52155_new_n22049_; 
wire u2__abc_52155_new_n22050_; 
wire u2__abc_52155_new_n22051_; 
wire u2__abc_52155_new_n22052_; 
wire u2__abc_52155_new_n22053_; 
wire u2__abc_52155_new_n22054_; 
wire u2__abc_52155_new_n22056_; 
wire u2__abc_52155_new_n22057_; 
wire u2__abc_52155_new_n22058_; 
wire u2__abc_52155_new_n22059_; 
wire u2__abc_52155_new_n22060_; 
wire u2__abc_52155_new_n22061_; 
wire u2__abc_52155_new_n22062_; 
wire u2__abc_52155_new_n22063_; 
wire u2__abc_52155_new_n22064_; 
wire u2__abc_52155_new_n22065_; 
wire u2__abc_52155_new_n22066_; 
wire u2__abc_52155_new_n22068_; 
wire u2__abc_52155_new_n22069_; 
wire u2__abc_52155_new_n22070_; 
wire u2__abc_52155_new_n22071_; 
wire u2__abc_52155_new_n22072_; 
wire u2__abc_52155_new_n22073_; 
wire u2__abc_52155_new_n22074_; 
wire u2__abc_52155_new_n22075_; 
wire u2__abc_52155_new_n22076_; 
wire u2__abc_52155_new_n22077_; 
wire u2__abc_52155_new_n22078_; 
wire u2__abc_52155_new_n22080_; 
wire u2__abc_52155_new_n22081_; 
wire u2__abc_52155_new_n22082_; 
wire u2__abc_52155_new_n22083_; 
wire u2__abc_52155_new_n22084_; 
wire u2__abc_52155_new_n22085_; 
wire u2__abc_52155_new_n22086_; 
wire u2__abc_52155_new_n22087_; 
wire u2__abc_52155_new_n22088_; 
wire u2__abc_52155_new_n22089_; 
wire u2__abc_52155_new_n22090_; 
wire u2__abc_52155_new_n22092_; 
wire u2__abc_52155_new_n22093_; 
wire u2__abc_52155_new_n22094_; 
wire u2__abc_52155_new_n22095_; 
wire u2__abc_52155_new_n22096_; 
wire u2__abc_52155_new_n22097_; 
wire u2__abc_52155_new_n22098_; 
wire u2__abc_52155_new_n22099_; 
wire u2__abc_52155_new_n22100_; 
wire u2__abc_52155_new_n22101_; 
wire u2__abc_52155_new_n22102_; 
wire u2__abc_52155_new_n22104_; 
wire u2__abc_52155_new_n22105_; 
wire u2__abc_52155_new_n22106_; 
wire u2__abc_52155_new_n22107_; 
wire u2__abc_52155_new_n22108_; 
wire u2__abc_52155_new_n22109_; 
wire u2__abc_52155_new_n22110_; 
wire u2__abc_52155_new_n22111_; 
wire u2__abc_52155_new_n22112_; 
wire u2__abc_52155_new_n22113_; 
wire u2__abc_52155_new_n22114_; 
wire u2__abc_52155_new_n22116_; 
wire u2__abc_52155_new_n22117_; 
wire u2__abc_52155_new_n22118_; 
wire u2__abc_52155_new_n22119_; 
wire u2__abc_52155_new_n22120_; 
wire u2__abc_52155_new_n22121_; 
wire u2__abc_52155_new_n22122_; 
wire u2__abc_52155_new_n22123_; 
wire u2__abc_52155_new_n22124_; 
wire u2__abc_52155_new_n22125_; 
wire u2__abc_52155_new_n22126_; 
wire u2__abc_52155_new_n22128_; 
wire u2__abc_52155_new_n22129_; 
wire u2__abc_52155_new_n22130_; 
wire u2__abc_52155_new_n22131_; 
wire u2__abc_52155_new_n22132_; 
wire u2__abc_52155_new_n22133_; 
wire u2__abc_52155_new_n22134_; 
wire u2__abc_52155_new_n22135_; 
wire u2__abc_52155_new_n22136_; 
wire u2__abc_52155_new_n22137_; 
wire u2__abc_52155_new_n22138_; 
wire u2__abc_52155_new_n22140_; 
wire u2__abc_52155_new_n22141_; 
wire u2__abc_52155_new_n22142_; 
wire u2__abc_52155_new_n22143_; 
wire u2__abc_52155_new_n22144_; 
wire u2__abc_52155_new_n22145_; 
wire u2__abc_52155_new_n22146_; 
wire u2__abc_52155_new_n22147_; 
wire u2__abc_52155_new_n22148_; 
wire u2__abc_52155_new_n22149_; 
wire u2__abc_52155_new_n22150_; 
wire u2__abc_52155_new_n22152_; 
wire u2__abc_52155_new_n22153_; 
wire u2__abc_52155_new_n22154_; 
wire u2__abc_52155_new_n22155_; 
wire u2__abc_52155_new_n22156_; 
wire u2__abc_52155_new_n22157_; 
wire u2__abc_52155_new_n22158_; 
wire u2__abc_52155_new_n22159_; 
wire u2__abc_52155_new_n22160_; 
wire u2__abc_52155_new_n22161_; 
wire u2__abc_52155_new_n22162_; 
wire u2__abc_52155_new_n22164_; 
wire u2__abc_52155_new_n22165_; 
wire u2__abc_52155_new_n22166_; 
wire u2__abc_52155_new_n22167_; 
wire u2__abc_52155_new_n22168_; 
wire u2__abc_52155_new_n22169_; 
wire u2__abc_52155_new_n22170_; 
wire u2__abc_52155_new_n22171_; 
wire u2__abc_52155_new_n22172_; 
wire u2__abc_52155_new_n22173_; 
wire u2__abc_52155_new_n22174_; 
wire u2__abc_52155_new_n22176_; 
wire u2__abc_52155_new_n22177_; 
wire u2__abc_52155_new_n22178_; 
wire u2__abc_52155_new_n22179_; 
wire u2__abc_52155_new_n22180_; 
wire u2__abc_52155_new_n22181_; 
wire u2__abc_52155_new_n22182_; 
wire u2__abc_52155_new_n22183_; 
wire u2__abc_52155_new_n22184_; 
wire u2__abc_52155_new_n22185_; 
wire u2__abc_52155_new_n22186_; 
wire u2__abc_52155_new_n22188_; 
wire u2__abc_52155_new_n22189_; 
wire u2__abc_52155_new_n22190_; 
wire u2__abc_52155_new_n22191_; 
wire u2__abc_52155_new_n22192_; 
wire u2__abc_52155_new_n22193_; 
wire u2__abc_52155_new_n22194_; 
wire u2__abc_52155_new_n22195_; 
wire u2__abc_52155_new_n22196_; 
wire u2__abc_52155_new_n22197_; 
wire u2__abc_52155_new_n22198_; 
wire u2__abc_52155_new_n22200_; 
wire u2__abc_52155_new_n22201_; 
wire u2__abc_52155_new_n22202_; 
wire u2__abc_52155_new_n22203_; 
wire u2__abc_52155_new_n22204_; 
wire u2__abc_52155_new_n22205_; 
wire u2__abc_52155_new_n22206_; 
wire u2__abc_52155_new_n22207_; 
wire u2__abc_52155_new_n22208_; 
wire u2__abc_52155_new_n22209_; 
wire u2__abc_52155_new_n22210_; 
wire u2__abc_52155_new_n22212_; 
wire u2__abc_52155_new_n22213_; 
wire u2__abc_52155_new_n22214_; 
wire u2__abc_52155_new_n22215_; 
wire u2__abc_52155_new_n22216_; 
wire u2__abc_52155_new_n22217_; 
wire u2__abc_52155_new_n22218_; 
wire u2__abc_52155_new_n22219_; 
wire u2__abc_52155_new_n22220_; 
wire u2__abc_52155_new_n22221_; 
wire u2__abc_52155_new_n22222_; 
wire u2__abc_52155_new_n22224_; 
wire u2__abc_52155_new_n22225_; 
wire u2__abc_52155_new_n22226_; 
wire u2__abc_52155_new_n22227_; 
wire u2__abc_52155_new_n22228_; 
wire u2__abc_52155_new_n22229_; 
wire u2__abc_52155_new_n22230_; 
wire u2__abc_52155_new_n22231_; 
wire u2__abc_52155_new_n22232_; 
wire u2__abc_52155_new_n22233_; 
wire u2__abc_52155_new_n22234_; 
wire u2__abc_52155_new_n22236_; 
wire u2__abc_52155_new_n22237_; 
wire u2__abc_52155_new_n22238_; 
wire u2__abc_52155_new_n22239_; 
wire u2__abc_52155_new_n22240_; 
wire u2__abc_52155_new_n22241_; 
wire u2__abc_52155_new_n22242_; 
wire u2__abc_52155_new_n22243_; 
wire u2__abc_52155_new_n22244_; 
wire u2__abc_52155_new_n22245_; 
wire u2__abc_52155_new_n22246_; 
wire u2__abc_52155_new_n22248_; 
wire u2__abc_52155_new_n22249_; 
wire u2__abc_52155_new_n22250_; 
wire u2__abc_52155_new_n22251_; 
wire u2__abc_52155_new_n22252_; 
wire u2__abc_52155_new_n22253_; 
wire u2__abc_52155_new_n22254_; 
wire u2__abc_52155_new_n22255_; 
wire u2__abc_52155_new_n22256_; 
wire u2__abc_52155_new_n22257_; 
wire u2__abc_52155_new_n22258_; 
wire u2__abc_52155_new_n22260_; 
wire u2__abc_52155_new_n22261_; 
wire u2__abc_52155_new_n22262_; 
wire u2__abc_52155_new_n22263_; 
wire u2__abc_52155_new_n22264_; 
wire u2__abc_52155_new_n22265_; 
wire u2__abc_52155_new_n22266_; 
wire u2__abc_52155_new_n22267_; 
wire u2__abc_52155_new_n22268_; 
wire u2__abc_52155_new_n22269_; 
wire u2__abc_52155_new_n22270_; 
wire u2__abc_52155_new_n22272_; 
wire u2__abc_52155_new_n22273_; 
wire u2__abc_52155_new_n22274_; 
wire u2__abc_52155_new_n22275_; 
wire u2__abc_52155_new_n22276_; 
wire u2__abc_52155_new_n22277_; 
wire u2__abc_52155_new_n22278_; 
wire u2__abc_52155_new_n22279_; 
wire u2__abc_52155_new_n22280_; 
wire u2__abc_52155_new_n22281_; 
wire u2__abc_52155_new_n22282_; 
wire u2__abc_52155_new_n22284_; 
wire u2__abc_52155_new_n22285_; 
wire u2__abc_52155_new_n22286_; 
wire u2__abc_52155_new_n22287_; 
wire u2__abc_52155_new_n22288_; 
wire u2__abc_52155_new_n22289_; 
wire u2__abc_52155_new_n22290_; 
wire u2__abc_52155_new_n22291_; 
wire u2__abc_52155_new_n22292_; 
wire u2__abc_52155_new_n22293_; 
wire u2__abc_52155_new_n22294_; 
wire u2__abc_52155_new_n22296_; 
wire u2__abc_52155_new_n22297_; 
wire u2__abc_52155_new_n22298_; 
wire u2__abc_52155_new_n22299_; 
wire u2__abc_52155_new_n22300_; 
wire u2__abc_52155_new_n22301_; 
wire u2__abc_52155_new_n22302_; 
wire u2__abc_52155_new_n22303_; 
wire u2__abc_52155_new_n22304_; 
wire u2__abc_52155_new_n22305_; 
wire u2__abc_52155_new_n22306_; 
wire u2__abc_52155_new_n22308_; 
wire u2__abc_52155_new_n22309_; 
wire u2__abc_52155_new_n22310_; 
wire u2__abc_52155_new_n22311_; 
wire u2__abc_52155_new_n22312_; 
wire u2__abc_52155_new_n22313_; 
wire u2__abc_52155_new_n22314_; 
wire u2__abc_52155_new_n22315_; 
wire u2__abc_52155_new_n22316_; 
wire u2__abc_52155_new_n22317_; 
wire u2__abc_52155_new_n22318_; 
wire u2__abc_52155_new_n22320_; 
wire u2__abc_52155_new_n22321_; 
wire u2__abc_52155_new_n22322_; 
wire u2__abc_52155_new_n22323_; 
wire u2__abc_52155_new_n22324_; 
wire u2__abc_52155_new_n22325_; 
wire u2__abc_52155_new_n22326_; 
wire u2__abc_52155_new_n22327_; 
wire u2__abc_52155_new_n22328_; 
wire u2__abc_52155_new_n22329_; 
wire u2__abc_52155_new_n22330_; 
wire u2__abc_52155_new_n22332_; 
wire u2__abc_52155_new_n22333_; 
wire u2__abc_52155_new_n22334_; 
wire u2__abc_52155_new_n22335_; 
wire u2__abc_52155_new_n22336_; 
wire u2__abc_52155_new_n22337_; 
wire u2__abc_52155_new_n22338_; 
wire u2__abc_52155_new_n22339_; 
wire u2__abc_52155_new_n22340_; 
wire u2__abc_52155_new_n22341_; 
wire u2__abc_52155_new_n22342_; 
wire u2__abc_52155_new_n22344_; 
wire u2__abc_52155_new_n22345_; 
wire u2__abc_52155_new_n22346_; 
wire u2__abc_52155_new_n22347_; 
wire u2__abc_52155_new_n22348_; 
wire u2__abc_52155_new_n22349_; 
wire u2__abc_52155_new_n22350_; 
wire u2__abc_52155_new_n22351_; 
wire u2__abc_52155_new_n22352_; 
wire u2__abc_52155_new_n22353_; 
wire u2__abc_52155_new_n22354_; 
wire u2__abc_52155_new_n22356_; 
wire u2__abc_52155_new_n22357_; 
wire u2__abc_52155_new_n22358_; 
wire u2__abc_52155_new_n22359_; 
wire u2__abc_52155_new_n22360_; 
wire u2__abc_52155_new_n22361_; 
wire u2__abc_52155_new_n22362_; 
wire u2__abc_52155_new_n22363_; 
wire u2__abc_52155_new_n22364_; 
wire u2__abc_52155_new_n22365_; 
wire u2__abc_52155_new_n22366_; 
wire u2__abc_52155_new_n22368_; 
wire u2__abc_52155_new_n22369_; 
wire u2__abc_52155_new_n22370_; 
wire u2__abc_52155_new_n22371_; 
wire u2__abc_52155_new_n22372_; 
wire u2__abc_52155_new_n22373_; 
wire u2__abc_52155_new_n22374_; 
wire u2__abc_52155_new_n22375_; 
wire u2__abc_52155_new_n22376_; 
wire u2__abc_52155_new_n22377_; 
wire u2__abc_52155_new_n22378_; 
wire u2__abc_52155_new_n22380_; 
wire u2__abc_52155_new_n22381_; 
wire u2__abc_52155_new_n22382_; 
wire u2__abc_52155_new_n22383_; 
wire u2__abc_52155_new_n22384_; 
wire u2__abc_52155_new_n22385_; 
wire u2__abc_52155_new_n22386_; 
wire u2__abc_52155_new_n22387_; 
wire u2__abc_52155_new_n22388_; 
wire u2__abc_52155_new_n22389_; 
wire u2__abc_52155_new_n22390_; 
wire u2__abc_52155_new_n22392_; 
wire u2__abc_52155_new_n22393_; 
wire u2__abc_52155_new_n22394_; 
wire u2__abc_52155_new_n22395_; 
wire u2__abc_52155_new_n22396_; 
wire u2__abc_52155_new_n22397_; 
wire u2__abc_52155_new_n22398_; 
wire u2__abc_52155_new_n22399_; 
wire u2__abc_52155_new_n22400_; 
wire u2__abc_52155_new_n22401_; 
wire u2__abc_52155_new_n22402_; 
wire u2__abc_52155_new_n22404_; 
wire u2__abc_52155_new_n22405_; 
wire u2__abc_52155_new_n22406_; 
wire u2__abc_52155_new_n22407_; 
wire u2__abc_52155_new_n22408_; 
wire u2__abc_52155_new_n22409_; 
wire u2__abc_52155_new_n22410_; 
wire u2__abc_52155_new_n22411_; 
wire u2__abc_52155_new_n22412_; 
wire u2__abc_52155_new_n22413_; 
wire u2__abc_52155_new_n22414_; 
wire u2__abc_52155_new_n22416_; 
wire u2__abc_52155_new_n22417_; 
wire u2__abc_52155_new_n22418_; 
wire u2__abc_52155_new_n22419_; 
wire u2__abc_52155_new_n22420_; 
wire u2__abc_52155_new_n22421_; 
wire u2__abc_52155_new_n22422_; 
wire u2__abc_52155_new_n22423_; 
wire u2__abc_52155_new_n22424_; 
wire u2__abc_52155_new_n22425_; 
wire u2__abc_52155_new_n22426_; 
wire u2__abc_52155_new_n22428_; 
wire u2__abc_52155_new_n22429_; 
wire u2__abc_52155_new_n22430_; 
wire u2__abc_52155_new_n22431_; 
wire u2__abc_52155_new_n22432_; 
wire u2__abc_52155_new_n22433_; 
wire u2__abc_52155_new_n22434_; 
wire u2__abc_52155_new_n22435_; 
wire u2__abc_52155_new_n22436_; 
wire u2__abc_52155_new_n22437_; 
wire u2__abc_52155_new_n22438_; 
wire u2__abc_52155_new_n22440_; 
wire u2__abc_52155_new_n22441_; 
wire u2__abc_52155_new_n22442_; 
wire u2__abc_52155_new_n22443_; 
wire u2__abc_52155_new_n22444_; 
wire u2__abc_52155_new_n22445_; 
wire u2__abc_52155_new_n22446_; 
wire u2__abc_52155_new_n22447_; 
wire u2__abc_52155_new_n22448_; 
wire u2__abc_52155_new_n22449_; 
wire u2__abc_52155_new_n22450_; 
wire u2__abc_52155_new_n22452_; 
wire u2__abc_52155_new_n22453_; 
wire u2__abc_52155_new_n22454_; 
wire u2__abc_52155_new_n22455_; 
wire u2__abc_52155_new_n22456_; 
wire u2__abc_52155_new_n22457_; 
wire u2__abc_52155_new_n22458_; 
wire u2__abc_52155_new_n22459_; 
wire u2__abc_52155_new_n22460_; 
wire u2__abc_52155_new_n22461_; 
wire u2__abc_52155_new_n22462_; 
wire u2__abc_52155_new_n22464_; 
wire u2__abc_52155_new_n22465_; 
wire u2__abc_52155_new_n22466_; 
wire u2__abc_52155_new_n22467_; 
wire u2__abc_52155_new_n22468_; 
wire u2__abc_52155_new_n22469_; 
wire u2__abc_52155_new_n22470_; 
wire u2__abc_52155_new_n22471_; 
wire u2__abc_52155_new_n22472_; 
wire u2__abc_52155_new_n22473_; 
wire u2__abc_52155_new_n22474_; 
wire u2__abc_52155_new_n22476_; 
wire u2__abc_52155_new_n22477_; 
wire u2__abc_52155_new_n22478_; 
wire u2__abc_52155_new_n22479_; 
wire u2__abc_52155_new_n22480_; 
wire u2__abc_52155_new_n22481_; 
wire u2__abc_52155_new_n22482_; 
wire u2__abc_52155_new_n22483_; 
wire u2__abc_52155_new_n22484_; 
wire u2__abc_52155_new_n22485_; 
wire u2__abc_52155_new_n22486_; 
wire u2__abc_52155_new_n22488_; 
wire u2__abc_52155_new_n22489_; 
wire u2__abc_52155_new_n22490_; 
wire u2__abc_52155_new_n22491_; 
wire u2__abc_52155_new_n22492_; 
wire u2__abc_52155_new_n22493_; 
wire u2__abc_52155_new_n22494_; 
wire u2__abc_52155_new_n22495_; 
wire u2__abc_52155_new_n22496_; 
wire u2__abc_52155_new_n22497_; 
wire u2__abc_52155_new_n22498_; 
wire u2__abc_52155_new_n22500_; 
wire u2__abc_52155_new_n22501_; 
wire u2__abc_52155_new_n22502_; 
wire u2__abc_52155_new_n22503_; 
wire u2__abc_52155_new_n22504_; 
wire u2__abc_52155_new_n22505_; 
wire u2__abc_52155_new_n22506_; 
wire u2__abc_52155_new_n22507_; 
wire u2__abc_52155_new_n22508_; 
wire u2__abc_52155_new_n22509_; 
wire u2__abc_52155_new_n22510_; 
wire u2__abc_52155_new_n22512_; 
wire u2__abc_52155_new_n22513_; 
wire u2__abc_52155_new_n22514_; 
wire u2__abc_52155_new_n22515_; 
wire u2__abc_52155_new_n22516_; 
wire u2__abc_52155_new_n22517_; 
wire u2__abc_52155_new_n22518_; 
wire u2__abc_52155_new_n22519_; 
wire u2__abc_52155_new_n22520_; 
wire u2__abc_52155_new_n22521_; 
wire u2__abc_52155_new_n22522_; 
wire u2__abc_52155_new_n22524_; 
wire u2__abc_52155_new_n22525_; 
wire u2__abc_52155_new_n22526_; 
wire u2__abc_52155_new_n22527_; 
wire u2__abc_52155_new_n22528_; 
wire u2__abc_52155_new_n22529_; 
wire u2__abc_52155_new_n22530_; 
wire u2__abc_52155_new_n22531_; 
wire u2__abc_52155_new_n22532_; 
wire u2__abc_52155_new_n22533_; 
wire u2__abc_52155_new_n22534_; 
wire u2__abc_52155_new_n22536_; 
wire u2__abc_52155_new_n22537_; 
wire u2__abc_52155_new_n22538_; 
wire u2__abc_52155_new_n22539_; 
wire u2__abc_52155_new_n22540_; 
wire u2__abc_52155_new_n22541_; 
wire u2__abc_52155_new_n22542_; 
wire u2__abc_52155_new_n22543_; 
wire u2__abc_52155_new_n22544_; 
wire u2__abc_52155_new_n22545_; 
wire u2__abc_52155_new_n22546_; 
wire u2__abc_52155_new_n22548_; 
wire u2__abc_52155_new_n22549_; 
wire u2__abc_52155_new_n22550_; 
wire u2__abc_52155_new_n22551_; 
wire u2__abc_52155_new_n22552_; 
wire u2__abc_52155_new_n22553_; 
wire u2__abc_52155_new_n22554_; 
wire u2__abc_52155_new_n22555_; 
wire u2__abc_52155_new_n22556_; 
wire u2__abc_52155_new_n22557_; 
wire u2__abc_52155_new_n22558_; 
wire u2__abc_52155_new_n22560_; 
wire u2__abc_52155_new_n22561_; 
wire u2__abc_52155_new_n22562_; 
wire u2__abc_52155_new_n22563_; 
wire u2__abc_52155_new_n22564_; 
wire u2__abc_52155_new_n22565_; 
wire u2__abc_52155_new_n22566_; 
wire u2__abc_52155_new_n22567_; 
wire u2__abc_52155_new_n22568_; 
wire u2__abc_52155_new_n22569_; 
wire u2__abc_52155_new_n22570_; 
wire u2__abc_52155_new_n22572_; 
wire u2__abc_52155_new_n22573_; 
wire u2__abc_52155_new_n22574_; 
wire u2__abc_52155_new_n22575_; 
wire u2__abc_52155_new_n22576_; 
wire u2__abc_52155_new_n22577_; 
wire u2__abc_52155_new_n22578_; 
wire u2__abc_52155_new_n22579_; 
wire u2__abc_52155_new_n22580_; 
wire u2__abc_52155_new_n22581_; 
wire u2__abc_52155_new_n22582_; 
wire u2__abc_52155_new_n22584_; 
wire u2__abc_52155_new_n22585_; 
wire u2__abc_52155_new_n22586_; 
wire u2__abc_52155_new_n22587_; 
wire u2__abc_52155_new_n22588_; 
wire u2__abc_52155_new_n22589_; 
wire u2__abc_52155_new_n22590_; 
wire u2__abc_52155_new_n22591_; 
wire u2__abc_52155_new_n22592_; 
wire u2__abc_52155_new_n22593_; 
wire u2__abc_52155_new_n22594_; 
wire u2__abc_52155_new_n22596_; 
wire u2__abc_52155_new_n22597_; 
wire u2__abc_52155_new_n22598_; 
wire u2__abc_52155_new_n22599_; 
wire u2__abc_52155_new_n22600_; 
wire u2__abc_52155_new_n22601_; 
wire u2__abc_52155_new_n22602_; 
wire u2__abc_52155_new_n22603_; 
wire u2__abc_52155_new_n22604_; 
wire u2__abc_52155_new_n22605_; 
wire u2__abc_52155_new_n22606_; 
wire u2__abc_52155_new_n22608_; 
wire u2__abc_52155_new_n22609_; 
wire u2__abc_52155_new_n22610_; 
wire u2__abc_52155_new_n22611_; 
wire u2__abc_52155_new_n22612_; 
wire u2__abc_52155_new_n22613_; 
wire u2__abc_52155_new_n22614_; 
wire u2__abc_52155_new_n22615_; 
wire u2__abc_52155_new_n22616_; 
wire u2__abc_52155_new_n22617_; 
wire u2__abc_52155_new_n22618_; 
wire u2__abc_52155_new_n22620_; 
wire u2__abc_52155_new_n22621_; 
wire u2__abc_52155_new_n22622_; 
wire u2__abc_52155_new_n22623_; 
wire u2__abc_52155_new_n22624_; 
wire u2__abc_52155_new_n22625_; 
wire u2__abc_52155_new_n22626_; 
wire u2__abc_52155_new_n22627_; 
wire u2__abc_52155_new_n22628_; 
wire u2__abc_52155_new_n22629_; 
wire u2__abc_52155_new_n22630_; 
wire u2__abc_52155_new_n22632_; 
wire u2__abc_52155_new_n22633_; 
wire u2__abc_52155_new_n22634_; 
wire u2__abc_52155_new_n22635_; 
wire u2__abc_52155_new_n22636_; 
wire u2__abc_52155_new_n22637_; 
wire u2__abc_52155_new_n22638_; 
wire u2__abc_52155_new_n22639_; 
wire u2__abc_52155_new_n22640_; 
wire u2__abc_52155_new_n22641_; 
wire u2__abc_52155_new_n22642_; 
wire u2__abc_52155_new_n22644_; 
wire u2__abc_52155_new_n22645_; 
wire u2__abc_52155_new_n22646_; 
wire u2__abc_52155_new_n22647_; 
wire u2__abc_52155_new_n22648_; 
wire u2__abc_52155_new_n22649_; 
wire u2__abc_52155_new_n22650_; 
wire u2__abc_52155_new_n22651_; 
wire u2__abc_52155_new_n22652_; 
wire u2__abc_52155_new_n22653_; 
wire u2__abc_52155_new_n22654_; 
wire u2__abc_52155_new_n22656_; 
wire u2__abc_52155_new_n22657_; 
wire u2__abc_52155_new_n22658_; 
wire u2__abc_52155_new_n22659_; 
wire u2__abc_52155_new_n22660_; 
wire u2__abc_52155_new_n22661_; 
wire u2__abc_52155_new_n22662_; 
wire u2__abc_52155_new_n22663_; 
wire u2__abc_52155_new_n22664_; 
wire u2__abc_52155_new_n22665_; 
wire u2__abc_52155_new_n22666_; 
wire u2__abc_52155_new_n22668_; 
wire u2__abc_52155_new_n22669_; 
wire u2__abc_52155_new_n22670_; 
wire u2__abc_52155_new_n22671_; 
wire u2__abc_52155_new_n22672_; 
wire u2__abc_52155_new_n22673_; 
wire u2__abc_52155_new_n22674_; 
wire u2__abc_52155_new_n22675_; 
wire u2__abc_52155_new_n22676_; 
wire u2__abc_52155_new_n22677_; 
wire u2__abc_52155_new_n22678_; 
wire u2__abc_52155_new_n22680_; 
wire u2__abc_52155_new_n22681_; 
wire u2__abc_52155_new_n22682_; 
wire u2__abc_52155_new_n22683_; 
wire u2__abc_52155_new_n22684_; 
wire u2__abc_52155_new_n22685_; 
wire u2__abc_52155_new_n22686_; 
wire u2__abc_52155_new_n22687_; 
wire u2__abc_52155_new_n22688_; 
wire u2__abc_52155_new_n22689_; 
wire u2__abc_52155_new_n22690_; 
wire u2__abc_52155_new_n22692_; 
wire u2__abc_52155_new_n22693_; 
wire u2__abc_52155_new_n22694_; 
wire u2__abc_52155_new_n22695_; 
wire u2__abc_52155_new_n22696_; 
wire u2__abc_52155_new_n22697_; 
wire u2__abc_52155_new_n22698_; 
wire u2__abc_52155_new_n22699_; 
wire u2__abc_52155_new_n22700_; 
wire u2__abc_52155_new_n22701_; 
wire u2__abc_52155_new_n22702_; 
wire u2__abc_52155_new_n22704_; 
wire u2__abc_52155_new_n22705_; 
wire u2__abc_52155_new_n22706_; 
wire u2__abc_52155_new_n22707_; 
wire u2__abc_52155_new_n22708_; 
wire u2__abc_52155_new_n22709_; 
wire u2__abc_52155_new_n22710_; 
wire u2__abc_52155_new_n22711_; 
wire u2__abc_52155_new_n22712_; 
wire u2__abc_52155_new_n22713_; 
wire u2__abc_52155_new_n22714_; 
wire u2__abc_52155_new_n22716_; 
wire u2__abc_52155_new_n22717_; 
wire u2__abc_52155_new_n22718_; 
wire u2__abc_52155_new_n22719_; 
wire u2__abc_52155_new_n22720_; 
wire u2__abc_52155_new_n22721_; 
wire u2__abc_52155_new_n22722_; 
wire u2__abc_52155_new_n22723_; 
wire u2__abc_52155_new_n22724_; 
wire u2__abc_52155_new_n22725_; 
wire u2__abc_52155_new_n22726_; 
wire u2__abc_52155_new_n22728_; 
wire u2__abc_52155_new_n22729_; 
wire u2__abc_52155_new_n22730_; 
wire u2__abc_52155_new_n22731_; 
wire u2__abc_52155_new_n22732_; 
wire u2__abc_52155_new_n22733_; 
wire u2__abc_52155_new_n22734_; 
wire u2__abc_52155_new_n22735_; 
wire u2__abc_52155_new_n22736_; 
wire u2__abc_52155_new_n22737_; 
wire u2__abc_52155_new_n22738_; 
wire u2__abc_52155_new_n22740_; 
wire u2__abc_52155_new_n22741_; 
wire u2__abc_52155_new_n22742_; 
wire u2__abc_52155_new_n22743_; 
wire u2__abc_52155_new_n22744_; 
wire u2__abc_52155_new_n22745_; 
wire u2__abc_52155_new_n22746_; 
wire u2__abc_52155_new_n22747_; 
wire u2__abc_52155_new_n22748_; 
wire u2__abc_52155_new_n22749_; 
wire u2__abc_52155_new_n22750_; 
wire u2__abc_52155_new_n22752_; 
wire u2__abc_52155_new_n22753_; 
wire u2__abc_52155_new_n22754_; 
wire u2__abc_52155_new_n22755_; 
wire u2__abc_52155_new_n22756_; 
wire u2__abc_52155_new_n22757_; 
wire u2__abc_52155_new_n22758_; 
wire u2__abc_52155_new_n22759_; 
wire u2__abc_52155_new_n22760_; 
wire u2__abc_52155_new_n22761_; 
wire u2__abc_52155_new_n22762_; 
wire u2__abc_52155_new_n22764_; 
wire u2__abc_52155_new_n22765_; 
wire u2__abc_52155_new_n22766_; 
wire u2__abc_52155_new_n22767_; 
wire u2__abc_52155_new_n22768_; 
wire u2__abc_52155_new_n22769_; 
wire u2__abc_52155_new_n22770_; 
wire u2__abc_52155_new_n22771_; 
wire u2__abc_52155_new_n22772_; 
wire u2__abc_52155_new_n22773_; 
wire u2__abc_52155_new_n22774_; 
wire u2__abc_52155_new_n22776_; 
wire u2__abc_52155_new_n22777_; 
wire u2__abc_52155_new_n22778_; 
wire u2__abc_52155_new_n22779_; 
wire u2__abc_52155_new_n22780_; 
wire u2__abc_52155_new_n22781_; 
wire u2__abc_52155_new_n22782_; 
wire u2__abc_52155_new_n22783_; 
wire u2__abc_52155_new_n22784_; 
wire u2__abc_52155_new_n22785_; 
wire u2__abc_52155_new_n22786_; 
wire u2__abc_52155_new_n22788_; 
wire u2__abc_52155_new_n22789_; 
wire u2__abc_52155_new_n22790_; 
wire u2__abc_52155_new_n22791_; 
wire u2__abc_52155_new_n22792_; 
wire u2__abc_52155_new_n22793_; 
wire u2__abc_52155_new_n22794_; 
wire u2__abc_52155_new_n22795_; 
wire u2__abc_52155_new_n22796_; 
wire u2__abc_52155_new_n22797_; 
wire u2__abc_52155_new_n22798_; 
wire u2__abc_52155_new_n22800_; 
wire u2__abc_52155_new_n22801_; 
wire u2__abc_52155_new_n22802_; 
wire u2__abc_52155_new_n22803_; 
wire u2__abc_52155_new_n22804_; 
wire u2__abc_52155_new_n22805_; 
wire u2__abc_52155_new_n22806_; 
wire u2__abc_52155_new_n22807_; 
wire u2__abc_52155_new_n22808_; 
wire u2__abc_52155_new_n22809_; 
wire u2__abc_52155_new_n22810_; 
wire u2__abc_52155_new_n22812_; 
wire u2__abc_52155_new_n22813_; 
wire u2__abc_52155_new_n22814_; 
wire u2__abc_52155_new_n22815_; 
wire u2__abc_52155_new_n22816_; 
wire u2__abc_52155_new_n22817_; 
wire u2__abc_52155_new_n22818_; 
wire u2__abc_52155_new_n22819_; 
wire u2__abc_52155_new_n22820_; 
wire u2__abc_52155_new_n22821_; 
wire u2__abc_52155_new_n22822_; 
wire u2__abc_52155_new_n22824_; 
wire u2__abc_52155_new_n22825_; 
wire u2__abc_52155_new_n22826_; 
wire u2__abc_52155_new_n22827_; 
wire u2__abc_52155_new_n22828_; 
wire u2__abc_52155_new_n22829_; 
wire u2__abc_52155_new_n22830_; 
wire u2__abc_52155_new_n22831_; 
wire u2__abc_52155_new_n22832_; 
wire u2__abc_52155_new_n22833_; 
wire u2__abc_52155_new_n22834_; 
wire u2__abc_52155_new_n22836_; 
wire u2__abc_52155_new_n22837_; 
wire u2__abc_52155_new_n22838_; 
wire u2__abc_52155_new_n22839_; 
wire u2__abc_52155_new_n22840_; 
wire u2__abc_52155_new_n22841_; 
wire u2__abc_52155_new_n22842_; 
wire u2__abc_52155_new_n22843_; 
wire u2__abc_52155_new_n22844_; 
wire u2__abc_52155_new_n22845_; 
wire u2__abc_52155_new_n22846_; 
wire u2__abc_52155_new_n22848_; 
wire u2__abc_52155_new_n22849_; 
wire u2__abc_52155_new_n22850_; 
wire u2__abc_52155_new_n22851_; 
wire u2__abc_52155_new_n22852_; 
wire u2__abc_52155_new_n22853_; 
wire u2__abc_52155_new_n22854_; 
wire u2__abc_52155_new_n22855_; 
wire u2__abc_52155_new_n22856_; 
wire u2__abc_52155_new_n22857_; 
wire u2__abc_52155_new_n22858_; 
wire u2__abc_52155_new_n22860_; 
wire u2__abc_52155_new_n22861_; 
wire u2__abc_52155_new_n22862_; 
wire u2__abc_52155_new_n22863_; 
wire u2__abc_52155_new_n22864_; 
wire u2__abc_52155_new_n22865_; 
wire u2__abc_52155_new_n22866_; 
wire u2__abc_52155_new_n22867_; 
wire u2__abc_52155_new_n22868_; 
wire u2__abc_52155_new_n22869_; 
wire u2__abc_52155_new_n22870_; 
wire u2__abc_52155_new_n22872_; 
wire u2__abc_52155_new_n22873_; 
wire u2__abc_52155_new_n22874_; 
wire u2__abc_52155_new_n22875_; 
wire u2__abc_52155_new_n22876_; 
wire u2__abc_52155_new_n22877_; 
wire u2__abc_52155_new_n22878_; 
wire u2__abc_52155_new_n22879_; 
wire u2__abc_52155_new_n22880_; 
wire u2__abc_52155_new_n22881_; 
wire u2__abc_52155_new_n22882_; 
wire u2__abc_52155_new_n22884_; 
wire u2__abc_52155_new_n22885_; 
wire u2__abc_52155_new_n22886_; 
wire u2__abc_52155_new_n22887_; 
wire u2__abc_52155_new_n22888_; 
wire u2__abc_52155_new_n22889_; 
wire u2__abc_52155_new_n22890_; 
wire u2__abc_52155_new_n22891_; 
wire u2__abc_52155_new_n22892_; 
wire u2__abc_52155_new_n22893_; 
wire u2__abc_52155_new_n22894_; 
wire u2__abc_52155_new_n22896_; 
wire u2__abc_52155_new_n22897_; 
wire u2__abc_52155_new_n22898_; 
wire u2__abc_52155_new_n22899_; 
wire u2__abc_52155_new_n22900_; 
wire u2__abc_52155_new_n22901_; 
wire u2__abc_52155_new_n22902_; 
wire u2__abc_52155_new_n22903_; 
wire u2__abc_52155_new_n22904_; 
wire u2__abc_52155_new_n22905_; 
wire u2__abc_52155_new_n22906_; 
wire u2__abc_52155_new_n22908_; 
wire u2__abc_52155_new_n22909_; 
wire u2__abc_52155_new_n22910_; 
wire u2__abc_52155_new_n22911_; 
wire u2__abc_52155_new_n22912_; 
wire u2__abc_52155_new_n22913_; 
wire u2__abc_52155_new_n22914_; 
wire u2__abc_52155_new_n22915_; 
wire u2__abc_52155_new_n22916_; 
wire u2__abc_52155_new_n22917_; 
wire u2__abc_52155_new_n22918_; 
wire u2__abc_52155_new_n22920_; 
wire u2__abc_52155_new_n22921_; 
wire u2__abc_52155_new_n22922_; 
wire u2__abc_52155_new_n22923_; 
wire u2__abc_52155_new_n22924_; 
wire u2__abc_52155_new_n22925_; 
wire u2__abc_52155_new_n22926_; 
wire u2__abc_52155_new_n22927_; 
wire u2__abc_52155_new_n22928_; 
wire u2__abc_52155_new_n22929_; 
wire u2__abc_52155_new_n22930_; 
wire u2__abc_52155_new_n22932_; 
wire u2__abc_52155_new_n22933_; 
wire u2__abc_52155_new_n22934_; 
wire u2__abc_52155_new_n22935_; 
wire u2__abc_52155_new_n22936_; 
wire u2__abc_52155_new_n22937_; 
wire u2__abc_52155_new_n22938_; 
wire u2__abc_52155_new_n22939_; 
wire u2__abc_52155_new_n22940_; 
wire u2__abc_52155_new_n22941_; 
wire u2__abc_52155_new_n22942_; 
wire u2__abc_52155_new_n22944_; 
wire u2__abc_52155_new_n22945_; 
wire u2__abc_52155_new_n22946_; 
wire u2__abc_52155_new_n22947_; 
wire u2__abc_52155_new_n22948_; 
wire u2__abc_52155_new_n22949_; 
wire u2__abc_52155_new_n22950_; 
wire u2__abc_52155_new_n22951_; 
wire u2__abc_52155_new_n22952_; 
wire u2__abc_52155_new_n22953_; 
wire u2__abc_52155_new_n22954_; 
wire u2__abc_52155_new_n22956_; 
wire u2__abc_52155_new_n22957_; 
wire u2__abc_52155_new_n22958_; 
wire u2__abc_52155_new_n22959_; 
wire u2__abc_52155_new_n22960_; 
wire u2__abc_52155_new_n22961_; 
wire u2__abc_52155_new_n22962_; 
wire u2__abc_52155_new_n22963_; 
wire u2__abc_52155_new_n22964_; 
wire u2__abc_52155_new_n22965_; 
wire u2__abc_52155_new_n22966_; 
wire u2__abc_52155_new_n22968_; 
wire u2__abc_52155_new_n22969_; 
wire u2__abc_52155_new_n22970_; 
wire u2__abc_52155_new_n22971_; 
wire u2__abc_52155_new_n22972_; 
wire u2__abc_52155_new_n22973_; 
wire u2__abc_52155_new_n22974_; 
wire u2__abc_52155_new_n22975_; 
wire u2__abc_52155_new_n22976_; 
wire u2__abc_52155_new_n22977_; 
wire u2__abc_52155_new_n22978_; 
wire u2__abc_52155_new_n22980_; 
wire u2__abc_52155_new_n22981_; 
wire u2__abc_52155_new_n22982_; 
wire u2__abc_52155_new_n22983_; 
wire u2__abc_52155_new_n22984_; 
wire u2__abc_52155_new_n22985_; 
wire u2__abc_52155_new_n22986_; 
wire u2__abc_52155_new_n22987_; 
wire u2__abc_52155_new_n22988_; 
wire u2__abc_52155_new_n22989_; 
wire u2__abc_52155_new_n22990_; 
wire u2__abc_52155_new_n22992_; 
wire u2__abc_52155_new_n22993_; 
wire u2__abc_52155_new_n22994_; 
wire u2__abc_52155_new_n22995_; 
wire u2__abc_52155_new_n22996_; 
wire u2__abc_52155_new_n22997_; 
wire u2__abc_52155_new_n22998_; 
wire u2__abc_52155_new_n22999_; 
wire u2__abc_52155_new_n23000_; 
wire u2__abc_52155_new_n23001_; 
wire u2__abc_52155_new_n23002_; 
wire u2__abc_52155_new_n23004_; 
wire u2__abc_52155_new_n23005_; 
wire u2__abc_52155_new_n23006_; 
wire u2__abc_52155_new_n23007_; 
wire u2__abc_52155_new_n23008_; 
wire u2__abc_52155_new_n23009_; 
wire u2__abc_52155_new_n23010_; 
wire u2__abc_52155_new_n23011_; 
wire u2__abc_52155_new_n23012_; 
wire u2__abc_52155_new_n23013_; 
wire u2__abc_52155_new_n23014_; 
wire u2__abc_52155_new_n23016_; 
wire u2__abc_52155_new_n23017_; 
wire u2__abc_52155_new_n23018_; 
wire u2__abc_52155_new_n23019_; 
wire u2__abc_52155_new_n23020_; 
wire u2__abc_52155_new_n23021_; 
wire u2__abc_52155_new_n23022_; 
wire u2__abc_52155_new_n23023_; 
wire u2__abc_52155_new_n23024_; 
wire u2__abc_52155_new_n23025_; 
wire u2__abc_52155_new_n23026_; 
wire u2__abc_52155_new_n23028_; 
wire u2__abc_52155_new_n23029_; 
wire u2__abc_52155_new_n23030_; 
wire u2__abc_52155_new_n23031_; 
wire u2__abc_52155_new_n23032_; 
wire u2__abc_52155_new_n23033_; 
wire u2__abc_52155_new_n23034_; 
wire u2__abc_52155_new_n23035_; 
wire u2__abc_52155_new_n23036_; 
wire u2__abc_52155_new_n23037_; 
wire u2__abc_52155_new_n23038_; 
wire u2__abc_52155_new_n23040_; 
wire u2__abc_52155_new_n23041_; 
wire u2__abc_52155_new_n23042_; 
wire u2__abc_52155_new_n23043_; 
wire u2__abc_52155_new_n23044_; 
wire u2__abc_52155_new_n23045_; 
wire u2__abc_52155_new_n23046_; 
wire u2__abc_52155_new_n23047_; 
wire u2__abc_52155_new_n23048_; 
wire u2__abc_52155_new_n23049_; 
wire u2__abc_52155_new_n23050_; 
wire u2__abc_52155_new_n23052_; 
wire u2__abc_52155_new_n23053_; 
wire u2__abc_52155_new_n23054_; 
wire u2__abc_52155_new_n23055_; 
wire u2__abc_52155_new_n23056_; 
wire u2__abc_52155_new_n23057_; 
wire u2__abc_52155_new_n23058_; 
wire u2__abc_52155_new_n23059_; 
wire u2__abc_52155_new_n23060_; 
wire u2__abc_52155_new_n23061_; 
wire u2__abc_52155_new_n23062_; 
wire u2__abc_52155_new_n23064_; 
wire u2__abc_52155_new_n23065_; 
wire u2__abc_52155_new_n23066_; 
wire u2__abc_52155_new_n23067_; 
wire u2__abc_52155_new_n23068_; 
wire u2__abc_52155_new_n23069_; 
wire u2__abc_52155_new_n23070_; 
wire u2__abc_52155_new_n23071_; 
wire u2__abc_52155_new_n23072_; 
wire u2__abc_52155_new_n23073_; 
wire u2__abc_52155_new_n23074_; 
wire u2__abc_52155_new_n23076_; 
wire u2__abc_52155_new_n23077_; 
wire u2__abc_52155_new_n23078_; 
wire u2__abc_52155_new_n23079_; 
wire u2__abc_52155_new_n23080_; 
wire u2__abc_52155_new_n23081_; 
wire u2__abc_52155_new_n23082_; 
wire u2__abc_52155_new_n23083_; 
wire u2__abc_52155_new_n23084_; 
wire u2__abc_52155_new_n23085_; 
wire u2__abc_52155_new_n23086_; 
wire u2__abc_52155_new_n23088_; 
wire u2__abc_52155_new_n23089_; 
wire u2__abc_52155_new_n23090_; 
wire u2__abc_52155_new_n23091_; 
wire u2__abc_52155_new_n23092_; 
wire u2__abc_52155_new_n23093_; 
wire u2__abc_52155_new_n23094_; 
wire u2__abc_52155_new_n23095_; 
wire u2__abc_52155_new_n23096_; 
wire u2__abc_52155_new_n23097_; 
wire u2__abc_52155_new_n23098_; 
wire u2__abc_52155_new_n23100_; 
wire u2__abc_52155_new_n23101_; 
wire u2__abc_52155_new_n23102_; 
wire u2__abc_52155_new_n23103_; 
wire u2__abc_52155_new_n23104_; 
wire u2__abc_52155_new_n23105_; 
wire u2__abc_52155_new_n23106_; 
wire u2__abc_52155_new_n23107_; 
wire u2__abc_52155_new_n23108_; 
wire u2__abc_52155_new_n23109_; 
wire u2__abc_52155_new_n23110_; 
wire u2__abc_52155_new_n23112_; 
wire u2__abc_52155_new_n23113_; 
wire u2__abc_52155_new_n23114_; 
wire u2__abc_52155_new_n23115_; 
wire u2__abc_52155_new_n23116_; 
wire u2__abc_52155_new_n23117_; 
wire u2__abc_52155_new_n23118_; 
wire u2__abc_52155_new_n23119_; 
wire u2__abc_52155_new_n23120_; 
wire u2__abc_52155_new_n23121_; 
wire u2__abc_52155_new_n23122_; 
wire u2__abc_52155_new_n23124_; 
wire u2__abc_52155_new_n23125_; 
wire u2__abc_52155_new_n23126_; 
wire u2__abc_52155_new_n23127_; 
wire u2__abc_52155_new_n23128_; 
wire u2__abc_52155_new_n23129_; 
wire u2__abc_52155_new_n23130_; 
wire u2__abc_52155_new_n23131_; 
wire u2__abc_52155_new_n23132_; 
wire u2__abc_52155_new_n23133_; 
wire u2__abc_52155_new_n23134_; 
wire u2__abc_52155_new_n23136_; 
wire u2__abc_52155_new_n23137_; 
wire u2__abc_52155_new_n23138_; 
wire u2__abc_52155_new_n23139_; 
wire u2__abc_52155_new_n23140_; 
wire u2__abc_52155_new_n23141_; 
wire u2__abc_52155_new_n23142_; 
wire u2__abc_52155_new_n23143_; 
wire u2__abc_52155_new_n23144_; 
wire u2__abc_52155_new_n23145_; 
wire u2__abc_52155_new_n23146_; 
wire u2__abc_52155_new_n23148_; 
wire u2__abc_52155_new_n23149_; 
wire u2__abc_52155_new_n23150_; 
wire u2__abc_52155_new_n23151_; 
wire u2__abc_52155_new_n23152_; 
wire u2__abc_52155_new_n23153_; 
wire u2__abc_52155_new_n23154_; 
wire u2__abc_52155_new_n23155_; 
wire u2__abc_52155_new_n23156_; 
wire u2__abc_52155_new_n23157_; 
wire u2__abc_52155_new_n23158_; 
wire u2__abc_52155_new_n23160_; 
wire u2__abc_52155_new_n23161_; 
wire u2__abc_52155_new_n23162_; 
wire u2__abc_52155_new_n23163_; 
wire u2__abc_52155_new_n23164_; 
wire u2__abc_52155_new_n23165_; 
wire u2__abc_52155_new_n23166_; 
wire u2__abc_52155_new_n23167_; 
wire u2__abc_52155_new_n23168_; 
wire u2__abc_52155_new_n23169_; 
wire u2__abc_52155_new_n23170_; 
wire u2__abc_52155_new_n23172_; 
wire u2__abc_52155_new_n23173_; 
wire u2__abc_52155_new_n23174_; 
wire u2__abc_52155_new_n23175_; 
wire u2__abc_52155_new_n23176_; 
wire u2__abc_52155_new_n23177_; 
wire u2__abc_52155_new_n23178_; 
wire u2__abc_52155_new_n23179_; 
wire u2__abc_52155_new_n23180_; 
wire u2__abc_52155_new_n23181_; 
wire u2__abc_52155_new_n23182_; 
wire u2__abc_52155_new_n23184_; 
wire u2__abc_52155_new_n23185_; 
wire u2__abc_52155_new_n23186_; 
wire u2__abc_52155_new_n23187_; 
wire u2__abc_52155_new_n23188_; 
wire u2__abc_52155_new_n23189_; 
wire u2__abc_52155_new_n23190_; 
wire u2__abc_52155_new_n23191_; 
wire u2__abc_52155_new_n23192_; 
wire u2__abc_52155_new_n23193_; 
wire u2__abc_52155_new_n23194_; 
wire u2__abc_52155_new_n23196_; 
wire u2__abc_52155_new_n23197_; 
wire u2__abc_52155_new_n23198_; 
wire u2__abc_52155_new_n23199_; 
wire u2__abc_52155_new_n23200_; 
wire u2__abc_52155_new_n23201_; 
wire u2__abc_52155_new_n23202_; 
wire u2__abc_52155_new_n23203_; 
wire u2__abc_52155_new_n23204_; 
wire u2__abc_52155_new_n23205_; 
wire u2__abc_52155_new_n23206_; 
wire u2__abc_52155_new_n23208_; 
wire u2__abc_52155_new_n23209_; 
wire u2__abc_52155_new_n23210_; 
wire u2__abc_52155_new_n23211_; 
wire u2__abc_52155_new_n23212_; 
wire u2__abc_52155_new_n23213_; 
wire u2__abc_52155_new_n23214_; 
wire u2__abc_52155_new_n23215_; 
wire u2__abc_52155_new_n23216_; 
wire u2__abc_52155_new_n23217_; 
wire u2__abc_52155_new_n23218_; 
wire u2__abc_52155_new_n23220_; 
wire u2__abc_52155_new_n23221_; 
wire u2__abc_52155_new_n23222_; 
wire u2__abc_52155_new_n23223_; 
wire u2__abc_52155_new_n23224_; 
wire u2__abc_52155_new_n23225_; 
wire u2__abc_52155_new_n23226_; 
wire u2__abc_52155_new_n23227_; 
wire u2__abc_52155_new_n23228_; 
wire u2__abc_52155_new_n23229_; 
wire u2__abc_52155_new_n23230_; 
wire u2__abc_52155_new_n23232_; 
wire u2__abc_52155_new_n23233_; 
wire u2__abc_52155_new_n23234_; 
wire u2__abc_52155_new_n23235_; 
wire u2__abc_52155_new_n23236_; 
wire u2__abc_52155_new_n23237_; 
wire u2__abc_52155_new_n23238_; 
wire u2__abc_52155_new_n23239_; 
wire u2__abc_52155_new_n23240_; 
wire u2__abc_52155_new_n23241_; 
wire u2__abc_52155_new_n23242_; 
wire u2__abc_52155_new_n23244_; 
wire u2__abc_52155_new_n23245_; 
wire u2__abc_52155_new_n23246_; 
wire u2__abc_52155_new_n23247_; 
wire u2__abc_52155_new_n23248_; 
wire u2__abc_52155_new_n23249_; 
wire u2__abc_52155_new_n23250_; 
wire u2__abc_52155_new_n23251_; 
wire u2__abc_52155_new_n23252_; 
wire u2__abc_52155_new_n23253_; 
wire u2__abc_52155_new_n23254_; 
wire u2__abc_52155_new_n23256_; 
wire u2__abc_52155_new_n23257_; 
wire u2__abc_52155_new_n23258_; 
wire u2__abc_52155_new_n23259_; 
wire u2__abc_52155_new_n23260_; 
wire u2__abc_52155_new_n23261_; 
wire u2__abc_52155_new_n23262_; 
wire u2__abc_52155_new_n23263_; 
wire u2__abc_52155_new_n23264_; 
wire u2__abc_52155_new_n23265_; 
wire u2__abc_52155_new_n23266_; 
wire u2__abc_52155_new_n23268_; 
wire u2__abc_52155_new_n23269_; 
wire u2__abc_52155_new_n23270_; 
wire u2__abc_52155_new_n23271_; 
wire u2__abc_52155_new_n23272_; 
wire u2__abc_52155_new_n23273_; 
wire u2__abc_52155_new_n23274_; 
wire u2__abc_52155_new_n23275_; 
wire u2__abc_52155_new_n23276_; 
wire u2__abc_52155_new_n23277_; 
wire u2__abc_52155_new_n23278_; 
wire u2__abc_52155_new_n23280_; 
wire u2__abc_52155_new_n23281_; 
wire u2__abc_52155_new_n23282_; 
wire u2__abc_52155_new_n23283_; 
wire u2__abc_52155_new_n23284_; 
wire u2__abc_52155_new_n23285_; 
wire u2__abc_52155_new_n23286_; 
wire u2__abc_52155_new_n23287_; 
wire u2__abc_52155_new_n23288_; 
wire u2__abc_52155_new_n23289_; 
wire u2__abc_52155_new_n23290_; 
wire u2__abc_52155_new_n23292_; 
wire u2__abc_52155_new_n23293_; 
wire u2__abc_52155_new_n23294_; 
wire u2__abc_52155_new_n23295_; 
wire u2__abc_52155_new_n23296_; 
wire u2__abc_52155_new_n23297_; 
wire u2__abc_52155_new_n23298_; 
wire u2__abc_52155_new_n23299_; 
wire u2__abc_52155_new_n23300_; 
wire u2__abc_52155_new_n23301_; 
wire u2__abc_52155_new_n23302_; 
wire u2__abc_52155_new_n23304_; 
wire u2__abc_52155_new_n23305_; 
wire u2__abc_52155_new_n23306_; 
wire u2__abc_52155_new_n23307_; 
wire u2__abc_52155_new_n23308_; 
wire u2__abc_52155_new_n23309_; 
wire u2__abc_52155_new_n23310_; 
wire u2__abc_52155_new_n23311_; 
wire u2__abc_52155_new_n23312_; 
wire u2__abc_52155_new_n23313_; 
wire u2__abc_52155_new_n23314_; 
wire u2__abc_52155_new_n23316_; 
wire u2__abc_52155_new_n23317_; 
wire u2__abc_52155_new_n23318_; 
wire u2__abc_52155_new_n23319_; 
wire u2__abc_52155_new_n23320_; 
wire u2__abc_52155_new_n23321_; 
wire u2__abc_52155_new_n23322_; 
wire u2__abc_52155_new_n23323_; 
wire u2__abc_52155_new_n23324_; 
wire u2__abc_52155_new_n23325_; 
wire u2__abc_52155_new_n23326_; 
wire u2__abc_52155_new_n23328_; 
wire u2__abc_52155_new_n23329_; 
wire u2__abc_52155_new_n23330_; 
wire u2__abc_52155_new_n23331_; 
wire u2__abc_52155_new_n23332_; 
wire u2__abc_52155_new_n23333_; 
wire u2__abc_52155_new_n23334_; 
wire u2__abc_52155_new_n23335_; 
wire u2__abc_52155_new_n23336_; 
wire u2__abc_52155_new_n23337_; 
wire u2__abc_52155_new_n23338_; 
wire u2__abc_52155_new_n23340_; 
wire u2__abc_52155_new_n23341_; 
wire u2__abc_52155_new_n23342_; 
wire u2__abc_52155_new_n23343_; 
wire u2__abc_52155_new_n23344_; 
wire u2__abc_52155_new_n23345_; 
wire u2__abc_52155_new_n23346_; 
wire u2__abc_52155_new_n23347_; 
wire u2__abc_52155_new_n23348_; 
wire u2__abc_52155_new_n23349_; 
wire u2__abc_52155_new_n23350_; 
wire u2__abc_52155_new_n23352_; 
wire u2__abc_52155_new_n23353_; 
wire u2__abc_52155_new_n23354_; 
wire u2__abc_52155_new_n23355_; 
wire u2__abc_52155_new_n23356_; 
wire u2__abc_52155_new_n23357_; 
wire u2__abc_52155_new_n23358_; 
wire u2__abc_52155_new_n23359_; 
wire u2__abc_52155_new_n23360_; 
wire u2__abc_52155_new_n23361_; 
wire u2__abc_52155_new_n23362_; 
wire u2__abc_52155_new_n23364_; 
wire u2__abc_52155_new_n23365_; 
wire u2__abc_52155_new_n23366_; 
wire u2__abc_52155_new_n23367_; 
wire u2__abc_52155_new_n23368_; 
wire u2__abc_52155_new_n23369_; 
wire u2__abc_52155_new_n23370_; 
wire u2__abc_52155_new_n23371_; 
wire u2__abc_52155_new_n23372_; 
wire u2__abc_52155_new_n23373_; 
wire u2__abc_52155_new_n23374_; 
wire u2__abc_52155_new_n23376_; 
wire u2__abc_52155_new_n23377_; 
wire u2__abc_52155_new_n23378_; 
wire u2__abc_52155_new_n23379_; 
wire u2__abc_52155_new_n23380_; 
wire u2__abc_52155_new_n23381_; 
wire u2__abc_52155_new_n23382_; 
wire u2__abc_52155_new_n23383_; 
wire u2__abc_52155_new_n23384_; 
wire u2__abc_52155_new_n23385_; 
wire u2__abc_52155_new_n23386_; 
wire u2__abc_52155_new_n23388_; 
wire u2__abc_52155_new_n23389_; 
wire u2__abc_52155_new_n23390_; 
wire u2__abc_52155_new_n23391_; 
wire u2__abc_52155_new_n23392_; 
wire u2__abc_52155_new_n23393_; 
wire u2__abc_52155_new_n23394_; 
wire u2__abc_52155_new_n23395_; 
wire u2__abc_52155_new_n23396_; 
wire u2__abc_52155_new_n23397_; 
wire u2__abc_52155_new_n23398_; 
wire u2__abc_52155_new_n23400_; 
wire u2__abc_52155_new_n23401_; 
wire u2__abc_52155_new_n23402_; 
wire u2__abc_52155_new_n23403_; 
wire u2__abc_52155_new_n23404_; 
wire u2__abc_52155_new_n23405_; 
wire u2__abc_52155_new_n23406_; 
wire u2__abc_52155_new_n23407_; 
wire u2__abc_52155_new_n23408_; 
wire u2__abc_52155_new_n23409_; 
wire u2__abc_52155_new_n23410_; 
wire u2__abc_52155_new_n23412_; 
wire u2__abc_52155_new_n23413_; 
wire u2__abc_52155_new_n23414_; 
wire u2__abc_52155_new_n23415_; 
wire u2__abc_52155_new_n23416_; 
wire u2__abc_52155_new_n23417_; 
wire u2__abc_52155_new_n23418_; 
wire u2__abc_52155_new_n23419_; 
wire u2__abc_52155_new_n23420_; 
wire u2__abc_52155_new_n23421_; 
wire u2__abc_52155_new_n23422_; 
wire u2__abc_52155_new_n23424_; 
wire u2__abc_52155_new_n23425_; 
wire u2__abc_52155_new_n23426_; 
wire u2__abc_52155_new_n23427_; 
wire u2__abc_52155_new_n23428_; 
wire u2__abc_52155_new_n23429_; 
wire u2__abc_52155_new_n23430_; 
wire u2__abc_52155_new_n23431_; 
wire u2__abc_52155_new_n23432_; 
wire u2__abc_52155_new_n23433_; 
wire u2__abc_52155_new_n23434_; 
wire u2__abc_52155_new_n23436_; 
wire u2__abc_52155_new_n23437_; 
wire u2__abc_52155_new_n23438_; 
wire u2__abc_52155_new_n23439_; 
wire u2__abc_52155_new_n23440_; 
wire u2__abc_52155_new_n23441_; 
wire u2__abc_52155_new_n23442_; 
wire u2__abc_52155_new_n23443_; 
wire u2__abc_52155_new_n23444_; 
wire u2__abc_52155_new_n23445_; 
wire u2__abc_52155_new_n23446_; 
wire u2__abc_52155_new_n23448_; 
wire u2__abc_52155_new_n23449_; 
wire u2__abc_52155_new_n23450_; 
wire u2__abc_52155_new_n23451_; 
wire u2__abc_52155_new_n23452_; 
wire u2__abc_52155_new_n23453_; 
wire u2__abc_52155_new_n23454_; 
wire u2__abc_52155_new_n23455_; 
wire u2__abc_52155_new_n23456_; 
wire u2__abc_52155_new_n23457_; 
wire u2__abc_52155_new_n23458_; 
wire u2__abc_52155_new_n23460_; 
wire u2__abc_52155_new_n23461_; 
wire u2__abc_52155_new_n23462_; 
wire u2__abc_52155_new_n23463_; 
wire u2__abc_52155_new_n23464_; 
wire u2__abc_52155_new_n23465_; 
wire u2__abc_52155_new_n23466_; 
wire u2__abc_52155_new_n23467_; 
wire u2__abc_52155_new_n23468_; 
wire u2__abc_52155_new_n23469_; 
wire u2__abc_52155_new_n23470_; 
wire u2__abc_52155_new_n23472_; 
wire u2__abc_52155_new_n23473_; 
wire u2__abc_52155_new_n23474_; 
wire u2__abc_52155_new_n23475_; 
wire u2__abc_52155_new_n23476_; 
wire u2__abc_52155_new_n23477_; 
wire u2__abc_52155_new_n23478_; 
wire u2__abc_52155_new_n23479_; 
wire u2__abc_52155_new_n23480_; 
wire u2__abc_52155_new_n23481_; 
wire u2__abc_52155_new_n23482_; 
wire u2__abc_52155_new_n23484_; 
wire u2__abc_52155_new_n23485_; 
wire u2__abc_52155_new_n23486_; 
wire u2__abc_52155_new_n23487_; 
wire u2__abc_52155_new_n23488_; 
wire u2__abc_52155_new_n23489_; 
wire u2__abc_52155_new_n23490_; 
wire u2__abc_52155_new_n23491_; 
wire u2__abc_52155_new_n23492_; 
wire u2__abc_52155_new_n23493_; 
wire u2__abc_52155_new_n23494_; 
wire u2__abc_52155_new_n23496_; 
wire u2__abc_52155_new_n23497_; 
wire u2__abc_52155_new_n23498_; 
wire u2__abc_52155_new_n23499_; 
wire u2__abc_52155_new_n23500_; 
wire u2__abc_52155_new_n23501_; 
wire u2__abc_52155_new_n23502_; 
wire u2__abc_52155_new_n23503_; 
wire u2__abc_52155_new_n23504_; 
wire u2__abc_52155_new_n23505_; 
wire u2__abc_52155_new_n23506_; 
wire u2__abc_52155_new_n23508_; 
wire u2__abc_52155_new_n23509_; 
wire u2__abc_52155_new_n23510_; 
wire u2__abc_52155_new_n23511_; 
wire u2__abc_52155_new_n23512_; 
wire u2__abc_52155_new_n23513_; 
wire u2__abc_52155_new_n23514_; 
wire u2__abc_52155_new_n23515_; 
wire u2__abc_52155_new_n23516_; 
wire u2__abc_52155_new_n23517_; 
wire u2__abc_52155_new_n23518_; 
wire u2__abc_52155_new_n23520_; 
wire u2__abc_52155_new_n23521_; 
wire u2__abc_52155_new_n23522_; 
wire u2__abc_52155_new_n23523_; 
wire u2__abc_52155_new_n23524_; 
wire u2__abc_52155_new_n23525_; 
wire u2__abc_52155_new_n23526_; 
wire u2__abc_52155_new_n23527_; 
wire u2__abc_52155_new_n23528_; 
wire u2__abc_52155_new_n23529_; 
wire u2__abc_52155_new_n23530_; 
wire u2__abc_52155_new_n23532_; 
wire u2__abc_52155_new_n23533_; 
wire u2__abc_52155_new_n23534_; 
wire u2__abc_52155_new_n23535_; 
wire u2__abc_52155_new_n23536_; 
wire u2__abc_52155_new_n23537_; 
wire u2__abc_52155_new_n23538_; 
wire u2__abc_52155_new_n23539_; 
wire u2__abc_52155_new_n23540_; 
wire u2__abc_52155_new_n23541_; 
wire u2__abc_52155_new_n23542_; 
wire u2__abc_52155_new_n23544_; 
wire u2__abc_52155_new_n23545_; 
wire u2__abc_52155_new_n23546_; 
wire u2__abc_52155_new_n23547_; 
wire u2__abc_52155_new_n23548_; 
wire u2__abc_52155_new_n23549_; 
wire u2__abc_52155_new_n23550_; 
wire u2__abc_52155_new_n23551_; 
wire u2__abc_52155_new_n23552_; 
wire u2__abc_52155_new_n23553_; 
wire u2__abc_52155_new_n23554_; 
wire u2__abc_52155_new_n23556_; 
wire u2__abc_52155_new_n23557_; 
wire u2__abc_52155_new_n23558_; 
wire u2__abc_52155_new_n23559_; 
wire u2__abc_52155_new_n23560_; 
wire u2__abc_52155_new_n23561_; 
wire u2__abc_52155_new_n23562_; 
wire u2__abc_52155_new_n23563_; 
wire u2__abc_52155_new_n23564_; 
wire u2__abc_52155_new_n23565_; 
wire u2__abc_52155_new_n23566_; 
wire u2__abc_52155_new_n23568_; 
wire u2__abc_52155_new_n23569_; 
wire u2__abc_52155_new_n23570_; 
wire u2__abc_52155_new_n23571_; 
wire u2__abc_52155_new_n23572_; 
wire u2__abc_52155_new_n23573_; 
wire u2__abc_52155_new_n23574_; 
wire u2__abc_52155_new_n23575_; 
wire u2__abc_52155_new_n23576_; 
wire u2__abc_52155_new_n23577_; 
wire u2__abc_52155_new_n23578_; 
wire u2__abc_52155_new_n23580_; 
wire u2__abc_52155_new_n23581_; 
wire u2__abc_52155_new_n23582_; 
wire u2__abc_52155_new_n23583_; 
wire u2__abc_52155_new_n23584_; 
wire u2__abc_52155_new_n23585_; 
wire u2__abc_52155_new_n23586_; 
wire u2__abc_52155_new_n23587_; 
wire u2__abc_52155_new_n23588_; 
wire u2__abc_52155_new_n23589_; 
wire u2__abc_52155_new_n23590_; 
wire u2__abc_52155_new_n23592_; 
wire u2__abc_52155_new_n23593_; 
wire u2__abc_52155_new_n23594_; 
wire u2__abc_52155_new_n23595_; 
wire u2__abc_52155_new_n23596_; 
wire u2__abc_52155_new_n23597_; 
wire u2__abc_52155_new_n23598_; 
wire u2__abc_52155_new_n23599_; 
wire u2__abc_52155_new_n23600_; 
wire u2__abc_52155_new_n23601_; 
wire u2__abc_52155_new_n23602_; 
wire u2__abc_52155_new_n23604_; 
wire u2__abc_52155_new_n23605_; 
wire u2__abc_52155_new_n23606_; 
wire u2__abc_52155_new_n23607_; 
wire u2__abc_52155_new_n23608_; 
wire u2__abc_52155_new_n23609_; 
wire u2__abc_52155_new_n23610_; 
wire u2__abc_52155_new_n23611_; 
wire u2__abc_52155_new_n23612_; 
wire u2__abc_52155_new_n23613_; 
wire u2__abc_52155_new_n23614_; 
wire u2__abc_52155_new_n23616_; 
wire u2__abc_52155_new_n23617_; 
wire u2__abc_52155_new_n23618_; 
wire u2__abc_52155_new_n23619_; 
wire u2__abc_52155_new_n23620_; 
wire u2__abc_52155_new_n23621_; 
wire u2__abc_52155_new_n23622_; 
wire u2__abc_52155_new_n23623_; 
wire u2__abc_52155_new_n23624_; 
wire u2__abc_52155_new_n23625_; 
wire u2__abc_52155_new_n23626_; 
wire u2__abc_52155_new_n23628_; 
wire u2__abc_52155_new_n23629_; 
wire u2__abc_52155_new_n23630_; 
wire u2__abc_52155_new_n23631_; 
wire u2__abc_52155_new_n23632_; 
wire u2__abc_52155_new_n23633_; 
wire u2__abc_52155_new_n23634_; 
wire u2__abc_52155_new_n23635_; 
wire u2__abc_52155_new_n23636_; 
wire u2__abc_52155_new_n23637_; 
wire u2__abc_52155_new_n23638_; 
wire u2__abc_52155_new_n23640_; 
wire u2__abc_52155_new_n23641_; 
wire u2__abc_52155_new_n23642_; 
wire u2__abc_52155_new_n23643_; 
wire u2__abc_52155_new_n23644_; 
wire u2__abc_52155_new_n23645_; 
wire u2__abc_52155_new_n23646_; 
wire u2__abc_52155_new_n23647_; 
wire u2__abc_52155_new_n23648_; 
wire u2__abc_52155_new_n23649_; 
wire u2__abc_52155_new_n23650_; 
wire u2__abc_52155_new_n23652_; 
wire u2__abc_52155_new_n23653_; 
wire u2__abc_52155_new_n23654_; 
wire u2__abc_52155_new_n23655_; 
wire u2__abc_52155_new_n23656_; 
wire u2__abc_52155_new_n23657_; 
wire u2__abc_52155_new_n23658_; 
wire u2__abc_52155_new_n23659_; 
wire u2__abc_52155_new_n23660_; 
wire u2__abc_52155_new_n23661_; 
wire u2__abc_52155_new_n23662_; 
wire u2__abc_52155_new_n23664_; 
wire u2__abc_52155_new_n23665_; 
wire u2__abc_52155_new_n23666_; 
wire u2__abc_52155_new_n23667_; 
wire u2__abc_52155_new_n23668_; 
wire u2__abc_52155_new_n23669_; 
wire u2__abc_52155_new_n23670_; 
wire u2__abc_52155_new_n23671_; 
wire u2__abc_52155_new_n23672_; 
wire u2__abc_52155_new_n23673_; 
wire u2__abc_52155_new_n23674_; 
wire u2__abc_52155_new_n23676_; 
wire u2__abc_52155_new_n23677_; 
wire u2__abc_52155_new_n23678_; 
wire u2__abc_52155_new_n23679_; 
wire u2__abc_52155_new_n23680_; 
wire u2__abc_52155_new_n23681_; 
wire u2__abc_52155_new_n23682_; 
wire u2__abc_52155_new_n23683_; 
wire u2__abc_52155_new_n23684_; 
wire u2__abc_52155_new_n23685_; 
wire u2__abc_52155_new_n23686_; 
wire u2__abc_52155_new_n23688_; 
wire u2__abc_52155_new_n23689_; 
wire u2__abc_52155_new_n23690_; 
wire u2__abc_52155_new_n23691_; 
wire u2__abc_52155_new_n23692_; 
wire u2__abc_52155_new_n23693_; 
wire u2__abc_52155_new_n23694_; 
wire u2__abc_52155_new_n23695_; 
wire u2__abc_52155_new_n23696_; 
wire u2__abc_52155_new_n23697_; 
wire u2__abc_52155_new_n23698_; 
wire u2__abc_52155_new_n23700_; 
wire u2__abc_52155_new_n23701_; 
wire u2__abc_52155_new_n23702_; 
wire u2__abc_52155_new_n23703_; 
wire u2__abc_52155_new_n23704_; 
wire u2__abc_52155_new_n23705_; 
wire u2__abc_52155_new_n23706_; 
wire u2__abc_52155_new_n23707_; 
wire u2__abc_52155_new_n23708_; 
wire u2__abc_52155_new_n23709_; 
wire u2__abc_52155_new_n23710_; 
wire u2__abc_52155_new_n23712_; 
wire u2__abc_52155_new_n23713_; 
wire u2__abc_52155_new_n23714_; 
wire u2__abc_52155_new_n23715_; 
wire u2__abc_52155_new_n23716_; 
wire u2__abc_52155_new_n23717_; 
wire u2__abc_52155_new_n23718_; 
wire u2__abc_52155_new_n23719_; 
wire u2__abc_52155_new_n23720_; 
wire u2__abc_52155_new_n23721_; 
wire u2__abc_52155_new_n23722_; 
wire u2__abc_52155_new_n23724_; 
wire u2__abc_52155_new_n23725_; 
wire u2__abc_52155_new_n23726_; 
wire u2__abc_52155_new_n23727_; 
wire u2__abc_52155_new_n23728_; 
wire u2__abc_52155_new_n23729_; 
wire u2__abc_52155_new_n23730_; 
wire u2__abc_52155_new_n23731_; 
wire u2__abc_52155_new_n23732_; 
wire u2__abc_52155_new_n23733_; 
wire u2__abc_52155_new_n23734_; 
wire u2__abc_52155_new_n23736_; 
wire u2__abc_52155_new_n23737_; 
wire u2__abc_52155_new_n23738_; 
wire u2__abc_52155_new_n23739_; 
wire u2__abc_52155_new_n23740_; 
wire u2__abc_52155_new_n23741_; 
wire u2__abc_52155_new_n23742_; 
wire u2__abc_52155_new_n23743_; 
wire u2__abc_52155_new_n23744_; 
wire u2__abc_52155_new_n23745_; 
wire u2__abc_52155_new_n23746_; 
wire u2__abc_52155_new_n23748_; 
wire u2__abc_52155_new_n23749_; 
wire u2__abc_52155_new_n23750_; 
wire u2__abc_52155_new_n23751_; 
wire u2__abc_52155_new_n23752_; 
wire u2__abc_52155_new_n23753_; 
wire u2__abc_52155_new_n23754_; 
wire u2__abc_52155_new_n23755_; 
wire u2__abc_52155_new_n23756_; 
wire u2__abc_52155_new_n23757_; 
wire u2__abc_52155_new_n23758_; 
wire u2__abc_52155_new_n23760_; 
wire u2__abc_52155_new_n23761_; 
wire u2__abc_52155_new_n23762_; 
wire u2__abc_52155_new_n23763_; 
wire u2__abc_52155_new_n23764_; 
wire u2__abc_52155_new_n23765_; 
wire u2__abc_52155_new_n23766_; 
wire u2__abc_52155_new_n23767_; 
wire u2__abc_52155_new_n23768_; 
wire u2__abc_52155_new_n23769_; 
wire u2__abc_52155_new_n23770_; 
wire u2__abc_52155_new_n23772_; 
wire u2__abc_52155_new_n23773_; 
wire u2__abc_52155_new_n23774_; 
wire u2__abc_52155_new_n23775_; 
wire u2__abc_52155_new_n23776_; 
wire u2__abc_52155_new_n23777_; 
wire u2__abc_52155_new_n23778_; 
wire u2__abc_52155_new_n23779_; 
wire u2__abc_52155_new_n23780_; 
wire u2__abc_52155_new_n23781_; 
wire u2__abc_52155_new_n23782_; 
wire u2__abc_52155_new_n23784_; 
wire u2__abc_52155_new_n23785_; 
wire u2__abc_52155_new_n23786_; 
wire u2__abc_52155_new_n23787_; 
wire u2__abc_52155_new_n23788_; 
wire u2__abc_52155_new_n23789_; 
wire u2__abc_52155_new_n23790_; 
wire u2__abc_52155_new_n23791_; 
wire u2__abc_52155_new_n23792_; 
wire u2__abc_52155_new_n23793_; 
wire u2__abc_52155_new_n23794_; 
wire u2__abc_52155_new_n23796_; 
wire u2__abc_52155_new_n23797_; 
wire u2__abc_52155_new_n23798_; 
wire u2__abc_52155_new_n23799_; 
wire u2__abc_52155_new_n23800_; 
wire u2__abc_52155_new_n23801_; 
wire u2__abc_52155_new_n23802_; 
wire u2__abc_52155_new_n23803_; 
wire u2__abc_52155_new_n23804_; 
wire u2__abc_52155_new_n23805_; 
wire u2__abc_52155_new_n23806_; 
wire u2__abc_52155_new_n23808_; 
wire u2__abc_52155_new_n23809_; 
wire u2__abc_52155_new_n23810_; 
wire u2__abc_52155_new_n23811_; 
wire u2__abc_52155_new_n23812_; 
wire u2__abc_52155_new_n23813_; 
wire u2__abc_52155_new_n23814_; 
wire u2__abc_52155_new_n23815_; 
wire u2__abc_52155_new_n23816_; 
wire u2__abc_52155_new_n23817_; 
wire u2__abc_52155_new_n23818_; 
wire u2__abc_52155_new_n23820_; 
wire u2__abc_52155_new_n23821_; 
wire u2__abc_52155_new_n23822_; 
wire u2__abc_52155_new_n23823_; 
wire u2__abc_52155_new_n23824_; 
wire u2__abc_52155_new_n23825_; 
wire u2__abc_52155_new_n23826_; 
wire u2__abc_52155_new_n23827_; 
wire u2__abc_52155_new_n23828_; 
wire u2__abc_52155_new_n23829_; 
wire u2__abc_52155_new_n23830_; 
wire u2__abc_52155_new_n23832_; 
wire u2__abc_52155_new_n23833_; 
wire u2__abc_52155_new_n23834_; 
wire u2__abc_52155_new_n23835_; 
wire u2__abc_52155_new_n23836_; 
wire u2__abc_52155_new_n23837_; 
wire u2__abc_52155_new_n23838_; 
wire u2__abc_52155_new_n23839_; 
wire u2__abc_52155_new_n23840_; 
wire u2__abc_52155_new_n23841_; 
wire u2__abc_52155_new_n23842_; 
wire u2__abc_52155_new_n23844_; 
wire u2__abc_52155_new_n23845_; 
wire u2__abc_52155_new_n23846_; 
wire u2__abc_52155_new_n23847_; 
wire u2__abc_52155_new_n23848_; 
wire u2__abc_52155_new_n23849_; 
wire u2__abc_52155_new_n23850_; 
wire u2__abc_52155_new_n23851_; 
wire u2__abc_52155_new_n23852_; 
wire u2__abc_52155_new_n23853_; 
wire u2__abc_52155_new_n23854_; 
wire u2__abc_52155_new_n23856_; 
wire u2__abc_52155_new_n23857_; 
wire u2__abc_52155_new_n23858_; 
wire u2__abc_52155_new_n23859_; 
wire u2__abc_52155_new_n23860_; 
wire u2__abc_52155_new_n23861_; 
wire u2__abc_52155_new_n23862_; 
wire u2__abc_52155_new_n23863_; 
wire u2__abc_52155_new_n23864_; 
wire u2__abc_52155_new_n23865_; 
wire u2__abc_52155_new_n23866_; 
wire u2__abc_52155_new_n23868_; 
wire u2__abc_52155_new_n23869_; 
wire u2__abc_52155_new_n23870_; 
wire u2__abc_52155_new_n23871_; 
wire u2__abc_52155_new_n23872_; 
wire u2__abc_52155_new_n23873_; 
wire u2__abc_52155_new_n23874_; 
wire u2__abc_52155_new_n23875_; 
wire u2__abc_52155_new_n23876_; 
wire u2__abc_52155_new_n23877_; 
wire u2__abc_52155_new_n23878_; 
wire u2__abc_52155_new_n23880_; 
wire u2__abc_52155_new_n23881_; 
wire u2__abc_52155_new_n23882_; 
wire u2__abc_52155_new_n23883_; 
wire u2__abc_52155_new_n23884_; 
wire u2__abc_52155_new_n23885_; 
wire u2__abc_52155_new_n23886_; 
wire u2__abc_52155_new_n23887_; 
wire u2__abc_52155_new_n23888_; 
wire u2__abc_52155_new_n23889_; 
wire u2__abc_52155_new_n23890_; 
wire u2__abc_52155_new_n23892_; 
wire u2__abc_52155_new_n23893_; 
wire u2__abc_52155_new_n23894_; 
wire u2__abc_52155_new_n23895_; 
wire u2__abc_52155_new_n23896_; 
wire u2__abc_52155_new_n23897_; 
wire u2__abc_52155_new_n23898_; 
wire u2__abc_52155_new_n23899_; 
wire u2__abc_52155_new_n23900_; 
wire u2__abc_52155_new_n23901_; 
wire u2__abc_52155_new_n23902_; 
wire u2__abc_52155_new_n23904_; 
wire u2__abc_52155_new_n23905_; 
wire u2__abc_52155_new_n23906_; 
wire u2__abc_52155_new_n23907_; 
wire u2__abc_52155_new_n23908_; 
wire u2__abc_52155_new_n23909_; 
wire u2__abc_52155_new_n23910_; 
wire u2__abc_52155_new_n23911_; 
wire u2__abc_52155_new_n23912_; 
wire u2__abc_52155_new_n23913_; 
wire u2__abc_52155_new_n23914_; 
wire u2__abc_52155_new_n23916_; 
wire u2__abc_52155_new_n23917_; 
wire u2__abc_52155_new_n23918_; 
wire u2__abc_52155_new_n23919_; 
wire u2__abc_52155_new_n23920_; 
wire u2__abc_52155_new_n23921_; 
wire u2__abc_52155_new_n23922_; 
wire u2__abc_52155_new_n23923_; 
wire u2__abc_52155_new_n23924_; 
wire u2__abc_52155_new_n23925_; 
wire u2__abc_52155_new_n23926_; 
wire u2__abc_52155_new_n23928_; 
wire u2__abc_52155_new_n23929_; 
wire u2__abc_52155_new_n23930_; 
wire u2__abc_52155_new_n23931_; 
wire u2__abc_52155_new_n23932_; 
wire u2__abc_52155_new_n23933_; 
wire u2__abc_52155_new_n23934_; 
wire u2__abc_52155_new_n23935_; 
wire u2__abc_52155_new_n23936_; 
wire u2__abc_52155_new_n23937_; 
wire u2__abc_52155_new_n23938_; 
wire u2__abc_52155_new_n23940_; 
wire u2__abc_52155_new_n23941_; 
wire u2__abc_52155_new_n23942_; 
wire u2__abc_52155_new_n23943_; 
wire u2__abc_52155_new_n23944_; 
wire u2__abc_52155_new_n23945_; 
wire u2__abc_52155_new_n23946_; 
wire u2__abc_52155_new_n23947_; 
wire u2__abc_52155_new_n23948_; 
wire u2__abc_52155_new_n23949_; 
wire u2__abc_52155_new_n23950_; 
wire u2__abc_52155_new_n23952_; 
wire u2__abc_52155_new_n23953_; 
wire u2__abc_52155_new_n23954_; 
wire u2__abc_52155_new_n23955_; 
wire u2__abc_52155_new_n23956_; 
wire u2__abc_52155_new_n23957_; 
wire u2__abc_52155_new_n23958_; 
wire u2__abc_52155_new_n23959_; 
wire u2__abc_52155_new_n23960_; 
wire u2__abc_52155_new_n23961_; 
wire u2__abc_52155_new_n23962_; 
wire u2__abc_52155_new_n23964_; 
wire u2__abc_52155_new_n23965_; 
wire u2__abc_52155_new_n23966_; 
wire u2__abc_52155_new_n23967_; 
wire u2__abc_52155_new_n23968_; 
wire u2__abc_52155_new_n23969_; 
wire u2__abc_52155_new_n23970_; 
wire u2__abc_52155_new_n23971_; 
wire u2__abc_52155_new_n23972_; 
wire u2__abc_52155_new_n23973_; 
wire u2__abc_52155_new_n23974_; 
wire u2__abc_52155_new_n23976_; 
wire u2__abc_52155_new_n23977_; 
wire u2__abc_52155_new_n23978_; 
wire u2__abc_52155_new_n23979_; 
wire u2__abc_52155_new_n23980_; 
wire u2__abc_52155_new_n23981_; 
wire u2__abc_52155_new_n23982_; 
wire u2__abc_52155_new_n23983_; 
wire u2__abc_52155_new_n23984_; 
wire u2__abc_52155_new_n23985_; 
wire u2__abc_52155_new_n23986_; 
wire u2__abc_52155_new_n23988_; 
wire u2__abc_52155_new_n23989_; 
wire u2__abc_52155_new_n23990_; 
wire u2__abc_52155_new_n23991_; 
wire u2__abc_52155_new_n23992_; 
wire u2__abc_52155_new_n23993_; 
wire u2__abc_52155_new_n23994_; 
wire u2__abc_52155_new_n23995_; 
wire u2__abc_52155_new_n23996_; 
wire u2__abc_52155_new_n23997_; 
wire u2__abc_52155_new_n23998_; 
wire u2__abc_52155_new_n24000_; 
wire u2__abc_52155_new_n24001_; 
wire u2__abc_52155_new_n24002_; 
wire u2__abc_52155_new_n24003_; 
wire u2__abc_52155_new_n24004_; 
wire u2__abc_52155_new_n24005_; 
wire u2__abc_52155_new_n24006_; 
wire u2__abc_52155_new_n24007_; 
wire u2__abc_52155_new_n24008_; 
wire u2__abc_52155_new_n24009_; 
wire u2__abc_52155_new_n24010_; 
wire u2__abc_52155_new_n24012_; 
wire u2__abc_52155_new_n24013_; 
wire u2__abc_52155_new_n24014_; 
wire u2__abc_52155_new_n24015_; 
wire u2__abc_52155_new_n24016_; 
wire u2__abc_52155_new_n24017_; 
wire u2__abc_52155_new_n24018_; 
wire u2__abc_52155_new_n24019_; 
wire u2__abc_52155_new_n24020_; 
wire u2__abc_52155_new_n24021_; 
wire u2__abc_52155_new_n24022_; 
wire u2__abc_52155_new_n24024_; 
wire u2__abc_52155_new_n24025_; 
wire u2__abc_52155_new_n24026_; 
wire u2__abc_52155_new_n24027_; 
wire u2__abc_52155_new_n24028_; 
wire u2__abc_52155_new_n24029_; 
wire u2__abc_52155_new_n24030_; 
wire u2__abc_52155_new_n24031_; 
wire u2__abc_52155_new_n24032_; 
wire u2__abc_52155_new_n24033_; 
wire u2__abc_52155_new_n24034_; 
wire u2__abc_52155_new_n24036_; 
wire u2__abc_52155_new_n24037_; 
wire u2__abc_52155_new_n24038_; 
wire u2__abc_52155_new_n24039_; 
wire u2__abc_52155_new_n24040_; 
wire u2__abc_52155_new_n24041_; 
wire u2__abc_52155_new_n24042_; 
wire u2__abc_52155_new_n24043_; 
wire u2__abc_52155_new_n24044_; 
wire u2__abc_52155_new_n24045_; 
wire u2__abc_52155_new_n24046_; 
wire u2__abc_52155_new_n24048_; 
wire u2__abc_52155_new_n24049_; 
wire u2__abc_52155_new_n24050_; 
wire u2__abc_52155_new_n24051_; 
wire u2__abc_52155_new_n24052_; 
wire u2__abc_52155_new_n24053_; 
wire u2__abc_52155_new_n24054_; 
wire u2__abc_52155_new_n24055_; 
wire u2__abc_52155_new_n24056_; 
wire u2__abc_52155_new_n24057_; 
wire u2__abc_52155_new_n24058_; 
wire u2__abc_52155_new_n24060_; 
wire u2__abc_52155_new_n24061_; 
wire u2__abc_52155_new_n24062_; 
wire u2__abc_52155_new_n24063_; 
wire u2__abc_52155_new_n24064_; 
wire u2__abc_52155_new_n24065_; 
wire u2__abc_52155_new_n24066_; 
wire u2__abc_52155_new_n24067_; 
wire u2__abc_52155_new_n24068_; 
wire u2__abc_52155_new_n24069_; 
wire u2__abc_52155_new_n24070_; 
wire u2__abc_52155_new_n24072_; 
wire u2__abc_52155_new_n24073_; 
wire u2__abc_52155_new_n24074_; 
wire u2__abc_52155_new_n24075_; 
wire u2__abc_52155_new_n24076_; 
wire u2__abc_52155_new_n24077_; 
wire u2__abc_52155_new_n24078_; 
wire u2__abc_52155_new_n24079_; 
wire u2__abc_52155_new_n24080_; 
wire u2__abc_52155_new_n24081_; 
wire u2__abc_52155_new_n24082_; 
wire u2__abc_52155_new_n24084_; 
wire u2__abc_52155_new_n24085_; 
wire u2__abc_52155_new_n24086_; 
wire u2__abc_52155_new_n24087_; 
wire u2__abc_52155_new_n24088_; 
wire u2__abc_52155_new_n24089_; 
wire u2__abc_52155_new_n24090_; 
wire u2__abc_52155_new_n24091_; 
wire u2__abc_52155_new_n24092_; 
wire u2__abc_52155_new_n24093_; 
wire u2__abc_52155_new_n24094_; 
wire u2__abc_52155_new_n24096_; 
wire u2__abc_52155_new_n24097_; 
wire u2__abc_52155_new_n24098_; 
wire u2__abc_52155_new_n24099_; 
wire u2__abc_52155_new_n24100_; 
wire u2__abc_52155_new_n24101_; 
wire u2__abc_52155_new_n24102_; 
wire u2__abc_52155_new_n24103_; 
wire u2__abc_52155_new_n24104_; 
wire u2__abc_52155_new_n24105_; 
wire u2__abc_52155_new_n24106_; 
wire u2__abc_52155_new_n24108_; 
wire u2__abc_52155_new_n24109_; 
wire u2__abc_52155_new_n24110_; 
wire u2__abc_52155_new_n24111_; 
wire u2__abc_52155_new_n24112_; 
wire u2__abc_52155_new_n24113_; 
wire u2__abc_52155_new_n24114_; 
wire u2__abc_52155_new_n24115_; 
wire u2__abc_52155_new_n24116_; 
wire u2__abc_52155_new_n24117_; 
wire u2__abc_52155_new_n24118_; 
wire u2__abc_52155_new_n24120_; 
wire u2__abc_52155_new_n24121_; 
wire u2__abc_52155_new_n24122_; 
wire u2__abc_52155_new_n24123_; 
wire u2__abc_52155_new_n24124_; 
wire u2__abc_52155_new_n24125_; 
wire u2__abc_52155_new_n24126_; 
wire u2__abc_52155_new_n24127_; 
wire u2__abc_52155_new_n24128_; 
wire u2__abc_52155_new_n24129_; 
wire u2__abc_52155_new_n24130_; 
wire u2__abc_52155_new_n24132_; 
wire u2__abc_52155_new_n24133_; 
wire u2__abc_52155_new_n24134_; 
wire u2__abc_52155_new_n24135_; 
wire u2__abc_52155_new_n24136_; 
wire u2__abc_52155_new_n24137_; 
wire u2__abc_52155_new_n24138_; 
wire u2__abc_52155_new_n24139_; 
wire u2__abc_52155_new_n24140_; 
wire u2__abc_52155_new_n24141_; 
wire u2__abc_52155_new_n24142_; 
wire u2__abc_52155_new_n24144_; 
wire u2__abc_52155_new_n24145_; 
wire u2__abc_52155_new_n24146_; 
wire u2__abc_52155_new_n24147_; 
wire u2__abc_52155_new_n24148_; 
wire u2__abc_52155_new_n24149_; 
wire u2__abc_52155_new_n24150_; 
wire u2__abc_52155_new_n24151_; 
wire u2__abc_52155_new_n24152_; 
wire u2__abc_52155_new_n24153_; 
wire u2__abc_52155_new_n24154_; 
wire u2__abc_52155_new_n24156_; 
wire u2__abc_52155_new_n24157_; 
wire u2__abc_52155_new_n24158_; 
wire u2__abc_52155_new_n24159_; 
wire u2__abc_52155_new_n24160_; 
wire u2__abc_52155_new_n24161_; 
wire u2__abc_52155_new_n24162_; 
wire u2__abc_52155_new_n24163_; 
wire u2__abc_52155_new_n24164_; 
wire u2__abc_52155_new_n24165_; 
wire u2__abc_52155_new_n24166_; 
wire u2__abc_52155_new_n24168_; 
wire u2__abc_52155_new_n24169_; 
wire u2__abc_52155_new_n24170_; 
wire u2__abc_52155_new_n24171_; 
wire u2__abc_52155_new_n24172_; 
wire u2__abc_52155_new_n24173_; 
wire u2__abc_52155_new_n24174_; 
wire u2__abc_52155_new_n24175_; 
wire u2__abc_52155_new_n24176_; 
wire u2__abc_52155_new_n24177_; 
wire u2__abc_52155_new_n24178_; 
wire u2__abc_52155_new_n24180_; 
wire u2__abc_52155_new_n24181_; 
wire u2__abc_52155_new_n24182_; 
wire u2__abc_52155_new_n24183_; 
wire u2__abc_52155_new_n24184_; 
wire u2__abc_52155_new_n24185_; 
wire u2__abc_52155_new_n24186_; 
wire u2__abc_52155_new_n24187_; 
wire u2__abc_52155_new_n24188_; 
wire u2__abc_52155_new_n24189_; 
wire u2__abc_52155_new_n24190_; 
wire u2__abc_52155_new_n24192_; 
wire u2__abc_52155_new_n24193_; 
wire u2__abc_52155_new_n24194_; 
wire u2__abc_52155_new_n24195_; 
wire u2__abc_52155_new_n24196_; 
wire u2__abc_52155_new_n24197_; 
wire u2__abc_52155_new_n24198_; 
wire u2__abc_52155_new_n24199_; 
wire u2__abc_52155_new_n24200_; 
wire u2__abc_52155_new_n24201_; 
wire u2__abc_52155_new_n24202_; 
wire u2__abc_52155_new_n24204_; 
wire u2__abc_52155_new_n24205_; 
wire u2__abc_52155_new_n24206_; 
wire u2__abc_52155_new_n24207_; 
wire u2__abc_52155_new_n24208_; 
wire u2__abc_52155_new_n24209_; 
wire u2__abc_52155_new_n24210_; 
wire u2__abc_52155_new_n24211_; 
wire u2__abc_52155_new_n24212_; 
wire u2__abc_52155_new_n24213_; 
wire u2__abc_52155_new_n24214_; 
wire u2__abc_52155_new_n24216_; 
wire u2__abc_52155_new_n24217_; 
wire u2__abc_52155_new_n24218_; 
wire u2__abc_52155_new_n24219_; 
wire u2__abc_52155_new_n24220_; 
wire u2__abc_52155_new_n24221_; 
wire u2__abc_52155_new_n24222_; 
wire u2__abc_52155_new_n24223_; 
wire u2__abc_52155_new_n24224_; 
wire u2__abc_52155_new_n24225_; 
wire u2__abc_52155_new_n24226_; 
wire u2__abc_52155_new_n24228_; 
wire u2__abc_52155_new_n24229_; 
wire u2__abc_52155_new_n24230_; 
wire u2__abc_52155_new_n24231_; 
wire u2__abc_52155_new_n24232_; 
wire u2__abc_52155_new_n24233_; 
wire u2__abc_52155_new_n24234_; 
wire u2__abc_52155_new_n24235_; 
wire u2__abc_52155_new_n24236_; 
wire u2__abc_52155_new_n24237_; 
wire u2__abc_52155_new_n24238_; 
wire u2__abc_52155_new_n24240_; 
wire u2__abc_52155_new_n24241_; 
wire u2__abc_52155_new_n24242_; 
wire u2__abc_52155_new_n24243_; 
wire u2__abc_52155_new_n24244_; 
wire u2__abc_52155_new_n24245_; 
wire u2__abc_52155_new_n24246_; 
wire u2__abc_52155_new_n24247_; 
wire u2__abc_52155_new_n24248_; 
wire u2__abc_52155_new_n24249_; 
wire u2__abc_52155_new_n24250_; 
wire u2__abc_52155_new_n24252_; 
wire u2__abc_52155_new_n24253_; 
wire u2__abc_52155_new_n24254_; 
wire u2__abc_52155_new_n24255_; 
wire u2__abc_52155_new_n24256_; 
wire u2__abc_52155_new_n24257_; 
wire u2__abc_52155_new_n24258_; 
wire u2__abc_52155_new_n24259_; 
wire u2__abc_52155_new_n24260_; 
wire u2__abc_52155_new_n24261_; 
wire u2__abc_52155_new_n24262_; 
wire u2__abc_52155_new_n24264_; 
wire u2__abc_52155_new_n24265_; 
wire u2__abc_52155_new_n24266_; 
wire u2__abc_52155_new_n24267_; 
wire u2__abc_52155_new_n24268_; 
wire u2__abc_52155_new_n24269_; 
wire u2__abc_52155_new_n24270_; 
wire u2__abc_52155_new_n24271_; 
wire u2__abc_52155_new_n24272_; 
wire u2__abc_52155_new_n24273_; 
wire u2__abc_52155_new_n24274_; 
wire u2__abc_52155_new_n24276_; 
wire u2__abc_52155_new_n24277_; 
wire u2__abc_52155_new_n24278_; 
wire u2__abc_52155_new_n24279_; 
wire u2__abc_52155_new_n24280_; 
wire u2__abc_52155_new_n24281_; 
wire u2__abc_52155_new_n24282_; 
wire u2__abc_52155_new_n24283_; 
wire u2__abc_52155_new_n24284_; 
wire u2__abc_52155_new_n24285_; 
wire u2__abc_52155_new_n24286_; 
wire u2__abc_52155_new_n24288_; 
wire u2__abc_52155_new_n24289_; 
wire u2__abc_52155_new_n24290_; 
wire u2__abc_52155_new_n24291_; 
wire u2__abc_52155_new_n24292_; 
wire u2__abc_52155_new_n24293_; 
wire u2__abc_52155_new_n24294_; 
wire u2__abc_52155_new_n24295_; 
wire u2__abc_52155_new_n24296_; 
wire u2__abc_52155_new_n24297_; 
wire u2__abc_52155_new_n24298_; 
wire u2__abc_52155_new_n24300_; 
wire u2__abc_52155_new_n24301_; 
wire u2__abc_52155_new_n24302_; 
wire u2__abc_52155_new_n24303_; 
wire u2__abc_52155_new_n24304_; 
wire u2__abc_52155_new_n24305_; 
wire u2__abc_52155_new_n24306_; 
wire u2__abc_52155_new_n24307_; 
wire u2__abc_52155_new_n24308_; 
wire u2__abc_52155_new_n24309_; 
wire u2__abc_52155_new_n24310_; 
wire u2__abc_52155_new_n24312_; 
wire u2__abc_52155_new_n24313_; 
wire u2__abc_52155_new_n24314_; 
wire u2__abc_52155_new_n24315_; 
wire u2__abc_52155_new_n24316_; 
wire u2__abc_52155_new_n24317_; 
wire u2__abc_52155_new_n24318_; 
wire u2__abc_52155_new_n24319_; 
wire u2__abc_52155_new_n24320_; 
wire u2__abc_52155_new_n24321_; 
wire u2__abc_52155_new_n24322_; 
wire u2__abc_52155_new_n24324_; 
wire u2__abc_52155_new_n24325_; 
wire u2__abc_52155_new_n24326_; 
wire u2__abc_52155_new_n24327_; 
wire u2__abc_52155_new_n24328_; 
wire u2__abc_52155_new_n24329_; 
wire u2__abc_52155_new_n24330_; 
wire u2__abc_52155_new_n24331_; 
wire u2__abc_52155_new_n24332_; 
wire u2__abc_52155_new_n24333_; 
wire u2__abc_52155_new_n24334_; 
wire u2__abc_52155_new_n24336_; 
wire u2__abc_52155_new_n24337_; 
wire u2__abc_52155_new_n24338_; 
wire u2__abc_52155_new_n24339_; 
wire u2__abc_52155_new_n24340_; 
wire u2__abc_52155_new_n24341_; 
wire u2__abc_52155_new_n24342_; 
wire u2__abc_52155_new_n24343_; 
wire u2__abc_52155_new_n24344_; 
wire u2__abc_52155_new_n24345_; 
wire u2__abc_52155_new_n24346_; 
wire u2__abc_52155_new_n24348_; 
wire u2__abc_52155_new_n24349_; 
wire u2__abc_52155_new_n24350_; 
wire u2__abc_52155_new_n24351_; 
wire u2__abc_52155_new_n24352_; 
wire u2__abc_52155_new_n24353_; 
wire u2__abc_52155_new_n24354_; 
wire u2__abc_52155_new_n24355_; 
wire u2__abc_52155_new_n24356_; 
wire u2__abc_52155_new_n24357_; 
wire u2__abc_52155_new_n24358_; 
wire u2__abc_52155_new_n24360_; 
wire u2__abc_52155_new_n24361_; 
wire u2__abc_52155_new_n24362_; 
wire u2__abc_52155_new_n24363_; 
wire u2__abc_52155_new_n24364_; 
wire u2__abc_52155_new_n24365_; 
wire u2__abc_52155_new_n24366_; 
wire u2__abc_52155_new_n24367_; 
wire u2__abc_52155_new_n24368_; 
wire u2__abc_52155_new_n24369_; 
wire u2__abc_52155_new_n24370_; 
wire u2__abc_52155_new_n24372_; 
wire u2__abc_52155_new_n24373_; 
wire u2__abc_52155_new_n24374_; 
wire u2__abc_52155_new_n24375_; 
wire u2__abc_52155_new_n24376_; 
wire u2__abc_52155_new_n24377_; 
wire u2__abc_52155_new_n24378_; 
wire u2__abc_52155_new_n24379_; 
wire u2__abc_52155_new_n24380_; 
wire u2__abc_52155_new_n24381_; 
wire u2__abc_52155_new_n24382_; 
wire u2__abc_52155_new_n24384_; 
wire u2__abc_52155_new_n24385_; 
wire u2__abc_52155_new_n24386_; 
wire u2__abc_52155_new_n24387_; 
wire u2__abc_52155_new_n24388_; 
wire u2__abc_52155_new_n24389_; 
wire u2__abc_52155_new_n24390_; 
wire u2__abc_52155_new_n24391_; 
wire u2__abc_52155_new_n24392_; 
wire u2__abc_52155_new_n24393_; 
wire u2__abc_52155_new_n24394_; 
wire u2__abc_52155_new_n24396_; 
wire u2__abc_52155_new_n24397_; 
wire u2__abc_52155_new_n24398_; 
wire u2__abc_52155_new_n24399_; 
wire u2__abc_52155_new_n24400_; 
wire u2__abc_52155_new_n24401_; 
wire u2__abc_52155_new_n24402_; 
wire u2__abc_52155_new_n24403_; 
wire u2__abc_52155_new_n24404_; 
wire u2__abc_52155_new_n24405_; 
wire u2__abc_52155_new_n24406_; 
wire u2__abc_52155_new_n24408_; 
wire u2__abc_52155_new_n24409_; 
wire u2__abc_52155_new_n24410_; 
wire u2__abc_52155_new_n24411_; 
wire u2__abc_52155_new_n24412_; 
wire u2__abc_52155_new_n24413_; 
wire u2__abc_52155_new_n24414_; 
wire u2__abc_52155_new_n24415_; 
wire u2__abc_52155_new_n24416_; 
wire u2__abc_52155_new_n24417_; 
wire u2__abc_52155_new_n24418_; 
wire u2__abc_52155_new_n24420_; 
wire u2__abc_52155_new_n24421_; 
wire u2__abc_52155_new_n24422_; 
wire u2__abc_52155_new_n24423_; 
wire u2__abc_52155_new_n24424_; 
wire u2__abc_52155_new_n24425_; 
wire u2__abc_52155_new_n24426_; 
wire u2__abc_52155_new_n24427_; 
wire u2__abc_52155_new_n24428_; 
wire u2__abc_52155_new_n24429_; 
wire u2__abc_52155_new_n24430_; 
wire u2__abc_52155_new_n24432_; 
wire u2__abc_52155_new_n24433_; 
wire u2__abc_52155_new_n24434_; 
wire u2__abc_52155_new_n24435_; 
wire u2__abc_52155_new_n24436_; 
wire u2__abc_52155_new_n24437_; 
wire u2__abc_52155_new_n24438_; 
wire u2__abc_52155_new_n24439_; 
wire u2__abc_52155_new_n24440_; 
wire u2__abc_52155_new_n24441_; 
wire u2__abc_52155_new_n24442_; 
wire u2__abc_52155_new_n24444_; 
wire u2__abc_52155_new_n24445_; 
wire u2__abc_52155_new_n24446_; 
wire u2__abc_52155_new_n24447_; 
wire u2__abc_52155_new_n24448_; 
wire u2__abc_52155_new_n24449_; 
wire u2__abc_52155_new_n24450_; 
wire u2__abc_52155_new_n24451_; 
wire u2__abc_52155_new_n24452_; 
wire u2__abc_52155_new_n24453_; 
wire u2__abc_52155_new_n24454_; 
wire u2__abc_52155_new_n24456_; 
wire u2__abc_52155_new_n24457_; 
wire u2__abc_52155_new_n24458_; 
wire u2__abc_52155_new_n24459_; 
wire u2__abc_52155_new_n24460_; 
wire u2__abc_52155_new_n24461_; 
wire u2__abc_52155_new_n24462_; 
wire u2__abc_52155_new_n24463_; 
wire u2__abc_52155_new_n24464_; 
wire u2__abc_52155_new_n24465_; 
wire u2__abc_52155_new_n24466_; 
wire u2__abc_52155_new_n2962_; 
wire u2__abc_52155_new_n2963_; 
wire u2__abc_52155_new_n2964_; 
wire u2__abc_52155_new_n2965_; 
wire u2__abc_52155_new_n2966_; 
wire u2__abc_52155_new_n2967_; 
wire u2__abc_52155_new_n2968_; 
wire u2__abc_52155_new_n2969_; 
wire u2__abc_52155_new_n2970_; 
wire u2__abc_52155_new_n2971_; 
wire u2__abc_52155_new_n2972_; 
wire u2__abc_52155_new_n2973_; 
wire u2__abc_52155_new_n2974_; 
wire u2__abc_52155_new_n2975_; 
wire u2__abc_52155_new_n2976_; 
wire u2__abc_52155_new_n2977_; 
wire u2__abc_52155_new_n2978_; 
wire u2__abc_52155_new_n2980_; 
wire u2__abc_52155_new_n2981_; 
wire u2__abc_52155_new_n2982_; 
wire u2__abc_52155_new_n2983_; 
wire u2__abc_52155_new_n2984_; 
wire u2__abc_52155_new_n2985_; 
wire u2__abc_52155_new_n2986_; 
wire u2__abc_52155_new_n2987_; 
wire u2__abc_52155_new_n2989_; 
wire u2__abc_52155_new_n2990_; 
wire u2__abc_52155_new_n2991_; 
wire u2__abc_52155_new_n2992_; 
wire u2__abc_52155_new_n2993_; 
wire u2__abc_52155_new_n2994_; 
wire u2__abc_52155_new_n2995_; 
wire u2__abc_52155_new_n2997_; 
wire u2__abc_52155_new_n2998_; 
wire u2__abc_52155_new_n2999_; 
wire u2__abc_52155_new_n3000_; 
wire u2__abc_52155_new_n3001_; 
wire u2__abc_52155_new_n3002_; 
wire u2__abc_52155_new_n3003_; 
wire u2__abc_52155_new_n3004_; 
wire u2__abc_52155_new_n3005_; 
wire u2__abc_52155_new_n3006_; 
wire u2__abc_52155_new_n3007_; 
wire u2__abc_52155_new_n3008_; 
wire u2__abc_52155_new_n3009_; 
wire u2__abc_52155_new_n3010_; 
wire u2__abc_52155_new_n3011_; 
wire u2__abc_52155_new_n3012_; 
wire u2__abc_52155_new_n3013_; 
wire u2__abc_52155_new_n3014_; 
wire u2__abc_52155_new_n3015_; 
wire u2__abc_52155_new_n3016_; 
wire u2__abc_52155_new_n3017_; 
wire u2__abc_52155_new_n3018_; 
wire u2__abc_52155_new_n3019_; 
wire u2__abc_52155_new_n3020_; 
wire u2__abc_52155_new_n3021_; 
wire u2__abc_52155_new_n3022_; 
wire u2__abc_52155_new_n3023_; 
wire u2__abc_52155_new_n3024_; 
wire u2__abc_52155_new_n3025_; 
wire u2__abc_52155_new_n3026_; 
wire u2__abc_52155_new_n3027_; 
wire u2__abc_52155_new_n3028_; 
wire u2__abc_52155_new_n3029_; 
wire u2__abc_52155_new_n3030_; 
wire u2__abc_52155_new_n3031_; 
wire u2__abc_52155_new_n3032_; 
wire u2__abc_52155_new_n3033_; 
wire u2__abc_52155_new_n3034_; 
wire u2__abc_52155_new_n3035_; 
wire u2__abc_52155_new_n3036_; 
wire u2__abc_52155_new_n3037_; 
wire u2__abc_52155_new_n3038_; 
wire u2__abc_52155_new_n3039_; 
wire u2__abc_52155_new_n3040_; 
wire u2__abc_52155_new_n3041_; 
wire u2__abc_52155_new_n3042_; 
wire u2__abc_52155_new_n3043_; 
wire u2__abc_52155_new_n3044_; 
wire u2__abc_52155_new_n3045_; 
wire u2__abc_52155_new_n3046_; 
wire u2__abc_52155_new_n3047_; 
wire u2__abc_52155_new_n3048_; 
wire u2__abc_52155_new_n3049_; 
wire u2__abc_52155_new_n3050_; 
wire u2__abc_52155_new_n3051_; 
wire u2__abc_52155_new_n3052_; 
wire u2__abc_52155_new_n3053_; 
wire u2__abc_52155_new_n3054_; 
wire u2__abc_52155_new_n3055_; 
wire u2__abc_52155_new_n3056_; 
wire u2__abc_52155_new_n3057_; 
wire u2__abc_52155_new_n3058_; 
wire u2__abc_52155_new_n3059_; 
wire u2__abc_52155_new_n3060_; 
wire u2__abc_52155_new_n3061_; 
wire u2__abc_52155_new_n3062_; 
wire u2__abc_52155_new_n3063_; 
wire u2__abc_52155_new_n3064_; 
wire u2__abc_52155_new_n3065_; 
wire u2__abc_52155_new_n3066_; 
wire u2__abc_52155_new_n3067_; 
wire u2__abc_52155_new_n3068_; 
wire u2__abc_52155_new_n3069_; 
wire u2__abc_52155_new_n3070_; 
wire u2__abc_52155_new_n3071_; 
wire u2__abc_52155_new_n3072_; 
wire u2__abc_52155_new_n3073_; 
wire u2__abc_52155_new_n3074_; 
wire u2__abc_52155_new_n3075_; 
wire u2__abc_52155_new_n3076_; 
wire u2__abc_52155_new_n3077_; 
wire u2__abc_52155_new_n3078_; 
wire u2__abc_52155_new_n3079_; 
wire u2__abc_52155_new_n3080_; 
wire u2__abc_52155_new_n3081_; 
wire u2__abc_52155_new_n3082_; 
wire u2__abc_52155_new_n3083_; 
wire u2__abc_52155_new_n3084_; 
wire u2__abc_52155_new_n3085_; 
wire u2__abc_52155_new_n3086_; 
wire u2__abc_52155_new_n3087_; 
wire u2__abc_52155_new_n3088_; 
wire u2__abc_52155_new_n3089_; 
wire u2__abc_52155_new_n3090_; 
wire u2__abc_52155_new_n3091_; 
wire u2__abc_52155_new_n3092_; 
wire u2__abc_52155_new_n3093_; 
wire u2__abc_52155_new_n3094_; 
wire u2__abc_52155_new_n3095_; 
wire u2__abc_52155_new_n3096_; 
wire u2__abc_52155_new_n3097_; 
wire u2__abc_52155_new_n3098_; 
wire u2__abc_52155_new_n3099_; 
wire u2__abc_52155_new_n3100_; 
wire u2__abc_52155_new_n3101_; 
wire u2__abc_52155_new_n3102_; 
wire u2__abc_52155_new_n3103_; 
wire u2__abc_52155_new_n3104_; 
wire u2__abc_52155_new_n3105_; 
wire u2__abc_52155_new_n3106_; 
wire u2__abc_52155_new_n3107_; 
wire u2__abc_52155_new_n3108_; 
wire u2__abc_52155_new_n3109_; 
wire u2__abc_52155_new_n3110_; 
wire u2__abc_52155_new_n3111_; 
wire u2__abc_52155_new_n3112_; 
wire u2__abc_52155_new_n3113_; 
wire u2__abc_52155_new_n3114_; 
wire u2__abc_52155_new_n3115_; 
wire u2__abc_52155_new_n3116_; 
wire u2__abc_52155_new_n3117_; 
wire u2__abc_52155_new_n3118_; 
wire u2__abc_52155_new_n3119_; 
wire u2__abc_52155_new_n3120_; 
wire u2__abc_52155_new_n3121_; 
wire u2__abc_52155_new_n3122_; 
wire u2__abc_52155_new_n3123_; 
wire u2__abc_52155_new_n3124_; 
wire u2__abc_52155_new_n3125_; 
wire u2__abc_52155_new_n3126_; 
wire u2__abc_52155_new_n3127_; 
wire u2__abc_52155_new_n3128_; 
wire u2__abc_52155_new_n3129_; 
wire u2__abc_52155_new_n3130_; 
wire u2__abc_52155_new_n3131_; 
wire u2__abc_52155_new_n3132_; 
wire u2__abc_52155_new_n3133_; 
wire u2__abc_52155_new_n3134_; 
wire u2__abc_52155_new_n3135_; 
wire u2__abc_52155_new_n3136_; 
wire u2__abc_52155_new_n3137_; 
wire u2__abc_52155_new_n3138_; 
wire u2__abc_52155_new_n3139_; 
wire u2__abc_52155_new_n3140_; 
wire u2__abc_52155_new_n3141_; 
wire u2__abc_52155_new_n3142_; 
wire u2__abc_52155_new_n3143_; 
wire u2__abc_52155_new_n3144_; 
wire u2__abc_52155_new_n3145_; 
wire u2__abc_52155_new_n3146_; 
wire u2__abc_52155_new_n3147_; 
wire u2__abc_52155_new_n3148_; 
wire u2__abc_52155_new_n3149_; 
wire u2__abc_52155_new_n3150_; 
wire u2__abc_52155_new_n3151_; 
wire u2__abc_52155_new_n3152_; 
wire u2__abc_52155_new_n3153_; 
wire u2__abc_52155_new_n3154_; 
wire u2__abc_52155_new_n3155_; 
wire u2__abc_52155_new_n3156_; 
wire u2__abc_52155_new_n3157_; 
wire u2__abc_52155_new_n3158_; 
wire u2__abc_52155_new_n3159_; 
wire u2__abc_52155_new_n3160_; 
wire u2__abc_52155_new_n3161_; 
wire u2__abc_52155_new_n3162_; 
wire u2__abc_52155_new_n3163_; 
wire u2__abc_52155_new_n3164_; 
wire u2__abc_52155_new_n3165_; 
wire u2__abc_52155_new_n3166_; 
wire u2__abc_52155_new_n3167_; 
wire u2__abc_52155_new_n3168_; 
wire u2__abc_52155_new_n3169_; 
wire u2__abc_52155_new_n3170_; 
wire u2__abc_52155_new_n3171_; 
wire u2__abc_52155_new_n3172_; 
wire u2__abc_52155_new_n3173_; 
wire u2__abc_52155_new_n3174_; 
wire u2__abc_52155_new_n3175_; 
wire u2__abc_52155_new_n3176_; 
wire u2__abc_52155_new_n3177_; 
wire u2__abc_52155_new_n3178_; 
wire u2__abc_52155_new_n3179_; 
wire u2__abc_52155_new_n3180_; 
wire u2__abc_52155_new_n3181_; 
wire u2__abc_52155_new_n3182_; 
wire u2__abc_52155_new_n3183_; 
wire u2__abc_52155_new_n3184_; 
wire u2__abc_52155_new_n3185_; 
wire u2__abc_52155_new_n3186_; 
wire u2__abc_52155_new_n3187_; 
wire u2__abc_52155_new_n3188_; 
wire u2__abc_52155_new_n3189_; 
wire u2__abc_52155_new_n3190_; 
wire u2__abc_52155_new_n3191_; 
wire u2__abc_52155_new_n3192_; 
wire u2__abc_52155_new_n3193_; 
wire u2__abc_52155_new_n3194_; 
wire u2__abc_52155_new_n3195_; 
wire u2__abc_52155_new_n3196_; 
wire u2__abc_52155_new_n3197_; 
wire u2__abc_52155_new_n3198_; 
wire u2__abc_52155_new_n3199_; 
wire u2__abc_52155_new_n3200_; 
wire u2__abc_52155_new_n3201_; 
wire u2__abc_52155_new_n3202_; 
wire u2__abc_52155_new_n3203_; 
wire u2__abc_52155_new_n3204_; 
wire u2__abc_52155_new_n3205_; 
wire u2__abc_52155_new_n3206_; 
wire u2__abc_52155_new_n3207_; 
wire u2__abc_52155_new_n3208_; 
wire u2__abc_52155_new_n3209_; 
wire u2__abc_52155_new_n3210_; 
wire u2__abc_52155_new_n3211_; 
wire u2__abc_52155_new_n3212_; 
wire u2__abc_52155_new_n3213_; 
wire u2__abc_52155_new_n3214_; 
wire u2__abc_52155_new_n3215_; 
wire u2__abc_52155_new_n3216_; 
wire u2__abc_52155_new_n3217_; 
wire u2__abc_52155_new_n3218_; 
wire u2__abc_52155_new_n3219_; 
wire u2__abc_52155_new_n3220_; 
wire u2__abc_52155_new_n3221_; 
wire u2__abc_52155_new_n3222_; 
wire u2__abc_52155_new_n3223_; 
wire u2__abc_52155_new_n3224_; 
wire u2__abc_52155_new_n3225_; 
wire u2__abc_52155_new_n3226_; 
wire u2__abc_52155_new_n3227_; 
wire u2__abc_52155_new_n3228_; 
wire u2__abc_52155_new_n3229_; 
wire u2__abc_52155_new_n3230_; 
wire u2__abc_52155_new_n3231_; 
wire u2__abc_52155_new_n3232_; 
wire u2__abc_52155_new_n3233_; 
wire u2__abc_52155_new_n3234_; 
wire u2__abc_52155_new_n3235_; 
wire u2__abc_52155_new_n3236_; 
wire u2__abc_52155_new_n3237_; 
wire u2__abc_52155_new_n3238_; 
wire u2__abc_52155_new_n3239_; 
wire u2__abc_52155_new_n3240_; 
wire u2__abc_52155_new_n3241_; 
wire u2__abc_52155_new_n3242_; 
wire u2__abc_52155_new_n3243_; 
wire u2__abc_52155_new_n3244_; 
wire u2__abc_52155_new_n3245_; 
wire u2__abc_52155_new_n3246_; 
wire u2__abc_52155_new_n3247_; 
wire u2__abc_52155_new_n3248_; 
wire u2__abc_52155_new_n3249_; 
wire u2__abc_52155_new_n3250_; 
wire u2__abc_52155_new_n3251_; 
wire u2__abc_52155_new_n3252_; 
wire u2__abc_52155_new_n3253_; 
wire u2__abc_52155_new_n3254_; 
wire u2__abc_52155_new_n3255_; 
wire u2__abc_52155_new_n3256_; 
wire u2__abc_52155_new_n3257_; 
wire u2__abc_52155_new_n3258_; 
wire u2__abc_52155_new_n3259_; 
wire u2__abc_52155_new_n3260_; 
wire u2__abc_52155_new_n3261_; 
wire u2__abc_52155_new_n3262_; 
wire u2__abc_52155_new_n3263_; 
wire u2__abc_52155_new_n3264_; 
wire u2__abc_52155_new_n3265_; 
wire u2__abc_52155_new_n3266_; 
wire u2__abc_52155_new_n3267_; 
wire u2__abc_52155_new_n3268_; 
wire u2__abc_52155_new_n3269_; 
wire u2__abc_52155_new_n3270_; 
wire u2__abc_52155_new_n3271_; 
wire u2__abc_52155_new_n3272_; 
wire u2__abc_52155_new_n3273_; 
wire u2__abc_52155_new_n3274_; 
wire u2__abc_52155_new_n3275_; 
wire u2__abc_52155_new_n3276_; 
wire u2__abc_52155_new_n3277_; 
wire u2__abc_52155_new_n3278_; 
wire u2__abc_52155_new_n3279_; 
wire u2__abc_52155_new_n3280_; 
wire u2__abc_52155_new_n3281_; 
wire u2__abc_52155_new_n3282_; 
wire u2__abc_52155_new_n3283_; 
wire u2__abc_52155_new_n3284_; 
wire u2__abc_52155_new_n3285_; 
wire u2__abc_52155_new_n3286_; 
wire u2__abc_52155_new_n3287_; 
wire u2__abc_52155_new_n3288_; 
wire u2__abc_52155_new_n3289_; 
wire u2__abc_52155_new_n3290_; 
wire u2__abc_52155_new_n3291_; 
wire u2__abc_52155_new_n3292_; 
wire u2__abc_52155_new_n3293_; 
wire u2__abc_52155_new_n3294_; 
wire u2__abc_52155_new_n3295_; 
wire u2__abc_52155_new_n3296_; 
wire u2__abc_52155_new_n3297_; 
wire u2__abc_52155_new_n3298_; 
wire u2__abc_52155_new_n3299_; 
wire u2__abc_52155_new_n3300_; 
wire u2__abc_52155_new_n3301_; 
wire u2__abc_52155_new_n3302_; 
wire u2__abc_52155_new_n3303_; 
wire u2__abc_52155_new_n3304_; 
wire u2__abc_52155_new_n3305_; 
wire u2__abc_52155_new_n3306_; 
wire u2__abc_52155_new_n3307_; 
wire u2__abc_52155_new_n3308_; 
wire u2__abc_52155_new_n3309_; 
wire u2__abc_52155_new_n3310_; 
wire u2__abc_52155_new_n3311_; 
wire u2__abc_52155_new_n3312_; 
wire u2__abc_52155_new_n3313_; 
wire u2__abc_52155_new_n3314_; 
wire u2__abc_52155_new_n3315_; 
wire u2__abc_52155_new_n3316_; 
wire u2__abc_52155_new_n3317_; 
wire u2__abc_52155_new_n3318_; 
wire u2__abc_52155_new_n3319_; 
wire u2__abc_52155_new_n3320_; 
wire u2__abc_52155_new_n3321_; 
wire u2__abc_52155_new_n3322_; 
wire u2__abc_52155_new_n3323_; 
wire u2__abc_52155_new_n3324_; 
wire u2__abc_52155_new_n3325_; 
wire u2__abc_52155_new_n3326_; 
wire u2__abc_52155_new_n3327_; 
wire u2__abc_52155_new_n3328_; 
wire u2__abc_52155_new_n3329_; 
wire u2__abc_52155_new_n3330_; 
wire u2__abc_52155_new_n3331_; 
wire u2__abc_52155_new_n3332_; 
wire u2__abc_52155_new_n3333_; 
wire u2__abc_52155_new_n3334_; 
wire u2__abc_52155_new_n3335_; 
wire u2__abc_52155_new_n3336_; 
wire u2__abc_52155_new_n3337_; 
wire u2__abc_52155_new_n3338_; 
wire u2__abc_52155_new_n3339_; 
wire u2__abc_52155_new_n3340_; 
wire u2__abc_52155_new_n3341_; 
wire u2__abc_52155_new_n3342_; 
wire u2__abc_52155_new_n3343_; 
wire u2__abc_52155_new_n3344_; 
wire u2__abc_52155_new_n3345_; 
wire u2__abc_52155_new_n3346_; 
wire u2__abc_52155_new_n3347_; 
wire u2__abc_52155_new_n3348_; 
wire u2__abc_52155_new_n3349_; 
wire u2__abc_52155_new_n3350_; 
wire u2__abc_52155_new_n3351_; 
wire u2__abc_52155_new_n3352_; 
wire u2__abc_52155_new_n3353_; 
wire u2__abc_52155_new_n3354_; 
wire u2__abc_52155_new_n3355_; 
wire u2__abc_52155_new_n3356_; 
wire u2__abc_52155_new_n3357_; 
wire u2__abc_52155_new_n3358_; 
wire u2__abc_52155_new_n3359_; 
wire u2__abc_52155_new_n3360_; 
wire u2__abc_52155_new_n3361_; 
wire u2__abc_52155_new_n3362_; 
wire u2__abc_52155_new_n3363_; 
wire u2__abc_52155_new_n3364_; 
wire u2__abc_52155_new_n3365_; 
wire u2__abc_52155_new_n3366_; 
wire u2__abc_52155_new_n3367_; 
wire u2__abc_52155_new_n3368_; 
wire u2__abc_52155_new_n3369_; 
wire u2__abc_52155_new_n3370_; 
wire u2__abc_52155_new_n3371_; 
wire u2__abc_52155_new_n3372_; 
wire u2__abc_52155_new_n3373_; 
wire u2__abc_52155_new_n3374_; 
wire u2__abc_52155_new_n3375_; 
wire u2__abc_52155_new_n3376_; 
wire u2__abc_52155_new_n3377_; 
wire u2__abc_52155_new_n3378_; 
wire u2__abc_52155_new_n3379_; 
wire u2__abc_52155_new_n3380_; 
wire u2__abc_52155_new_n3381_; 
wire u2__abc_52155_new_n3382_; 
wire u2__abc_52155_new_n3383_; 
wire u2__abc_52155_new_n3384_; 
wire u2__abc_52155_new_n3385_; 
wire u2__abc_52155_new_n3386_; 
wire u2__abc_52155_new_n3387_; 
wire u2__abc_52155_new_n3388_; 
wire u2__abc_52155_new_n3389_; 
wire u2__abc_52155_new_n3390_; 
wire u2__abc_52155_new_n3391_; 
wire u2__abc_52155_new_n3392_; 
wire u2__abc_52155_new_n3393_; 
wire u2__abc_52155_new_n3394_; 
wire u2__abc_52155_new_n3395_; 
wire u2__abc_52155_new_n3396_; 
wire u2__abc_52155_new_n3397_; 
wire u2__abc_52155_new_n3398_; 
wire u2__abc_52155_new_n3399_; 
wire u2__abc_52155_new_n3400_; 
wire u2__abc_52155_new_n3401_; 
wire u2__abc_52155_new_n3402_; 
wire u2__abc_52155_new_n3403_; 
wire u2__abc_52155_new_n3404_; 
wire u2__abc_52155_new_n3405_; 
wire u2__abc_52155_new_n3406_; 
wire u2__abc_52155_new_n3407_; 
wire u2__abc_52155_new_n3408_; 
wire u2__abc_52155_new_n3409_; 
wire u2__abc_52155_new_n3410_; 
wire u2__abc_52155_new_n3411_; 
wire u2__abc_52155_new_n3412_; 
wire u2__abc_52155_new_n3413_; 
wire u2__abc_52155_new_n3414_; 
wire u2__abc_52155_new_n3415_; 
wire u2__abc_52155_new_n3416_; 
wire u2__abc_52155_new_n3417_; 
wire u2__abc_52155_new_n3418_; 
wire u2__abc_52155_new_n3419_; 
wire u2__abc_52155_new_n3420_; 
wire u2__abc_52155_new_n3421_; 
wire u2__abc_52155_new_n3422_; 
wire u2__abc_52155_new_n3423_; 
wire u2__abc_52155_new_n3424_; 
wire u2__abc_52155_new_n3425_; 
wire u2__abc_52155_new_n3426_; 
wire u2__abc_52155_new_n3427_; 
wire u2__abc_52155_new_n3428_; 
wire u2__abc_52155_new_n3429_; 
wire u2__abc_52155_new_n3430_; 
wire u2__abc_52155_new_n3431_; 
wire u2__abc_52155_new_n3432_; 
wire u2__abc_52155_new_n3433_; 
wire u2__abc_52155_new_n3434_; 
wire u2__abc_52155_new_n3435_; 
wire u2__abc_52155_new_n3436_; 
wire u2__abc_52155_new_n3437_; 
wire u2__abc_52155_new_n3438_; 
wire u2__abc_52155_new_n3439_; 
wire u2__abc_52155_new_n3440_; 
wire u2__abc_52155_new_n3441_; 
wire u2__abc_52155_new_n3442_; 
wire u2__abc_52155_new_n3443_; 
wire u2__abc_52155_new_n3444_; 
wire u2__abc_52155_new_n3445_; 
wire u2__abc_52155_new_n3446_; 
wire u2__abc_52155_new_n3447_; 
wire u2__abc_52155_new_n3448_; 
wire u2__abc_52155_new_n3449_; 
wire u2__abc_52155_new_n3450_; 
wire u2__abc_52155_new_n3451_; 
wire u2__abc_52155_new_n3452_; 
wire u2__abc_52155_new_n3453_; 
wire u2__abc_52155_new_n3454_; 
wire u2__abc_52155_new_n3455_; 
wire u2__abc_52155_new_n3456_; 
wire u2__abc_52155_new_n3457_; 
wire u2__abc_52155_new_n3458_; 
wire u2__abc_52155_new_n3459_; 
wire u2__abc_52155_new_n3460_; 
wire u2__abc_52155_new_n3461_; 
wire u2__abc_52155_new_n3462_; 
wire u2__abc_52155_new_n3463_; 
wire u2__abc_52155_new_n3464_; 
wire u2__abc_52155_new_n3465_; 
wire u2__abc_52155_new_n3466_; 
wire u2__abc_52155_new_n3467_; 
wire u2__abc_52155_new_n3468_; 
wire u2__abc_52155_new_n3469_; 
wire u2__abc_52155_new_n3470_; 
wire u2__abc_52155_new_n3471_; 
wire u2__abc_52155_new_n3472_; 
wire u2__abc_52155_new_n3473_; 
wire u2__abc_52155_new_n3474_; 
wire u2__abc_52155_new_n3475_; 
wire u2__abc_52155_new_n3476_; 
wire u2__abc_52155_new_n3477_; 
wire u2__abc_52155_new_n3478_; 
wire u2__abc_52155_new_n3479_; 
wire u2__abc_52155_new_n3480_; 
wire u2__abc_52155_new_n3481_; 
wire u2__abc_52155_new_n3482_; 
wire u2__abc_52155_new_n3483_; 
wire u2__abc_52155_new_n3484_; 
wire u2__abc_52155_new_n3485_; 
wire u2__abc_52155_new_n3486_; 
wire u2__abc_52155_new_n3487_; 
wire u2__abc_52155_new_n3488_; 
wire u2__abc_52155_new_n3489_; 
wire u2__abc_52155_new_n3490_; 
wire u2__abc_52155_new_n3491_; 
wire u2__abc_52155_new_n3492_; 
wire u2__abc_52155_new_n3493_; 
wire u2__abc_52155_new_n3494_; 
wire u2__abc_52155_new_n3495_; 
wire u2__abc_52155_new_n3496_; 
wire u2__abc_52155_new_n3497_; 
wire u2__abc_52155_new_n3498_; 
wire u2__abc_52155_new_n3499_; 
wire u2__abc_52155_new_n3500_; 
wire u2__abc_52155_new_n3501_; 
wire u2__abc_52155_new_n3502_; 
wire u2__abc_52155_new_n3503_; 
wire u2__abc_52155_new_n3504_; 
wire u2__abc_52155_new_n3505_; 
wire u2__abc_52155_new_n3506_; 
wire u2__abc_52155_new_n3507_; 
wire u2__abc_52155_new_n3508_; 
wire u2__abc_52155_new_n3509_; 
wire u2__abc_52155_new_n3510_; 
wire u2__abc_52155_new_n3511_; 
wire u2__abc_52155_new_n3512_; 
wire u2__abc_52155_new_n3513_; 
wire u2__abc_52155_new_n3514_; 
wire u2__abc_52155_new_n3515_; 
wire u2__abc_52155_new_n3516_; 
wire u2__abc_52155_new_n3517_; 
wire u2__abc_52155_new_n3518_; 
wire u2__abc_52155_new_n3519_; 
wire u2__abc_52155_new_n3520_; 
wire u2__abc_52155_new_n3521_; 
wire u2__abc_52155_new_n3522_; 
wire u2__abc_52155_new_n3523_; 
wire u2__abc_52155_new_n3524_; 
wire u2__abc_52155_new_n3525_; 
wire u2__abc_52155_new_n3526_; 
wire u2__abc_52155_new_n3527_; 
wire u2__abc_52155_new_n3528_; 
wire u2__abc_52155_new_n3529_; 
wire u2__abc_52155_new_n3530_; 
wire u2__abc_52155_new_n3531_; 
wire u2__abc_52155_new_n3532_; 
wire u2__abc_52155_new_n3533_; 
wire u2__abc_52155_new_n3534_; 
wire u2__abc_52155_new_n3535_; 
wire u2__abc_52155_new_n3536_; 
wire u2__abc_52155_new_n3537_; 
wire u2__abc_52155_new_n3538_; 
wire u2__abc_52155_new_n3539_; 
wire u2__abc_52155_new_n3540_; 
wire u2__abc_52155_new_n3541_; 
wire u2__abc_52155_new_n3542_; 
wire u2__abc_52155_new_n3543_; 
wire u2__abc_52155_new_n3544_; 
wire u2__abc_52155_new_n3545_; 
wire u2__abc_52155_new_n3546_; 
wire u2__abc_52155_new_n3547_; 
wire u2__abc_52155_new_n3548_; 
wire u2__abc_52155_new_n3549_; 
wire u2__abc_52155_new_n3550_; 
wire u2__abc_52155_new_n3551_; 
wire u2__abc_52155_new_n3552_; 
wire u2__abc_52155_new_n3553_; 
wire u2__abc_52155_new_n3554_; 
wire u2__abc_52155_new_n3555_; 
wire u2__abc_52155_new_n3556_; 
wire u2__abc_52155_new_n3557_; 
wire u2__abc_52155_new_n3558_; 
wire u2__abc_52155_new_n3559_; 
wire u2__abc_52155_new_n3560_; 
wire u2__abc_52155_new_n3561_; 
wire u2__abc_52155_new_n3562_; 
wire u2__abc_52155_new_n3563_; 
wire u2__abc_52155_new_n3564_; 
wire u2__abc_52155_new_n3565_; 
wire u2__abc_52155_new_n3566_; 
wire u2__abc_52155_new_n3567_; 
wire u2__abc_52155_new_n3568_; 
wire u2__abc_52155_new_n3569_; 
wire u2__abc_52155_new_n3570_; 
wire u2__abc_52155_new_n3571_; 
wire u2__abc_52155_new_n3572_; 
wire u2__abc_52155_new_n3573_; 
wire u2__abc_52155_new_n3574_; 
wire u2__abc_52155_new_n3575_; 
wire u2__abc_52155_new_n3576_; 
wire u2__abc_52155_new_n3577_; 
wire u2__abc_52155_new_n3578_; 
wire u2__abc_52155_new_n3579_; 
wire u2__abc_52155_new_n3580_; 
wire u2__abc_52155_new_n3581_; 
wire u2__abc_52155_new_n3582_; 
wire u2__abc_52155_new_n3583_; 
wire u2__abc_52155_new_n3584_; 
wire u2__abc_52155_new_n3585_; 
wire u2__abc_52155_new_n3586_; 
wire u2__abc_52155_new_n3587_; 
wire u2__abc_52155_new_n3588_; 
wire u2__abc_52155_new_n3589_; 
wire u2__abc_52155_new_n3590_; 
wire u2__abc_52155_new_n3591_; 
wire u2__abc_52155_new_n3592_; 
wire u2__abc_52155_new_n3593_; 
wire u2__abc_52155_new_n3594_; 
wire u2__abc_52155_new_n3595_; 
wire u2__abc_52155_new_n3596_; 
wire u2__abc_52155_new_n3597_; 
wire u2__abc_52155_new_n3598_; 
wire u2__abc_52155_new_n3599_; 
wire u2__abc_52155_new_n3600_; 
wire u2__abc_52155_new_n3601_; 
wire u2__abc_52155_new_n3602_; 
wire u2__abc_52155_new_n3603_; 
wire u2__abc_52155_new_n3604_; 
wire u2__abc_52155_new_n3605_; 
wire u2__abc_52155_new_n3606_; 
wire u2__abc_52155_new_n3607_; 
wire u2__abc_52155_new_n3608_; 
wire u2__abc_52155_new_n3609_; 
wire u2__abc_52155_new_n3610_; 
wire u2__abc_52155_new_n3611_; 
wire u2__abc_52155_new_n3612_; 
wire u2__abc_52155_new_n3613_; 
wire u2__abc_52155_new_n3614_; 
wire u2__abc_52155_new_n3615_; 
wire u2__abc_52155_new_n3616_; 
wire u2__abc_52155_new_n3617_; 
wire u2__abc_52155_new_n3618_; 
wire u2__abc_52155_new_n3619_; 
wire u2__abc_52155_new_n3620_; 
wire u2__abc_52155_new_n3621_; 
wire u2__abc_52155_new_n3622_; 
wire u2__abc_52155_new_n3623_; 
wire u2__abc_52155_new_n3624_; 
wire u2__abc_52155_new_n3625_; 
wire u2__abc_52155_new_n3626_; 
wire u2__abc_52155_new_n3627_; 
wire u2__abc_52155_new_n3628_; 
wire u2__abc_52155_new_n3629_; 
wire u2__abc_52155_new_n3630_; 
wire u2__abc_52155_new_n3631_; 
wire u2__abc_52155_new_n3632_; 
wire u2__abc_52155_new_n3633_; 
wire u2__abc_52155_new_n3634_; 
wire u2__abc_52155_new_n3635_; 
wire u2__abc_52155_new_n3636_; 
wire u2__abc_52155_new_n3637_; 
wire u2__abc_52155_new_n3638_; 
wire u2__abc_52155_new_n3639_; 
wire u2__abc_52155_new_n3640_; 
wire u2__abc_52155_new_n3641_; 
wire u2__abc_52155_new_n3642_; 
wire u2__abc_52155_new_n3643_; 
wire u2__abc_52155_new_n3644_; 
wire u2__abc_52155_new_n3645_; 
wire u2__abc_52155_new_n3646_; 
wire u2__abc_52155_new_n3647_; 
wire u2__abc_52155_new_n3648_; 
wire u2__abc_52155_new_n3649_; 
wire u2__abc_52155_new_n3650_; 
wire u2__abc_52155_new_n3651_; 
wire u2__abc_52155_new_n3652_; 
wire u2__abc_52155_new_n3653_; 
wire u2__abc_52155_new_n3654_; 
wire u2__abc_52155_new_n3655_; 
wire u2__abc_52155_new_n3656_; 
wire u2__abc_52155_new_n3657_; 
wire u2__abc_52155_new_n3658_; 
wire u2__abc_52155_new_n3659_; 
wire u2__abc_52155_new_n3660_; 
wire u2__abc_52155_new_n3661_; 
wire u2__abc_52155_new_n3662_; 
wire u2__abc_52155_new_n3663_; 
wire u2__abc_52155_new_n3664_; 
wire u2__abc_52155_new_n3665_; 
wire u2__abc_52155_new_n3666_; 
wire u2__abc_52155_new_n3667_; 
wire u2__abc_52155_new_n3668_; 
wire u2__abc_52155_new_n3669_; 
wire u2__abc_52155_new_n3670_; 
wire u2__abc_52155_new_n3671_; 
wire u2__abc_52155_new_n3672_; 
wire u2__abc_52155_new_n3673_; 
wire u2__abc_52155_new_n3674_; 
wire u2__abc_52155_new_n3675_; 
wire u2__abc_52155_new_n3676_; 
wire u2__abc_52155_new_n3677_; 
wire u2__abc_52155_new_n3678_; 
wire u2__abc_52155_new_n3679_; 
wire u2__abc_52155_new_n3680_; 
wire u2__abc_52155_new_n3681_; 
wire u2__abc_52155_new_n3682_; 
wire u2__abc_52155_new_n3683_; 
wire u2__abc_52155_new_n3684_; 
wire u2__abc_52155_new_n3685_; 
wire u2__abc_52155_new_n3686_; 
wire u2__abc_52155_new_n3687_; 
wire u2__abc_52155_new_n3688_; 
wire u2__abc_52155_new_n3689_; 
wire u2__abc_52155_new_n3690_; 
wire u2__abc_52155_new_n3691_; 
wire u2__abc_52155_new_n3692_; 
wire u2__abc_52155_new_n3693_; 
wire u2__abc_52155_new_n3694_; 
wire u2__abc_52155_new_n3695_; 
wire u2__abc_52155_new_n3696_; 
wire u2__abc_52155_new_n3697_; 
wire u2__abc_52155_new_n3698_; 
wire u2__abc_52155_new_n3699_; 
wire u2__abc_52155_new_n3700_; 
wire u2__abc_52155_new_n3701_; 
wire u2__abc_52155_new_n3702_; 
wire u2__abc_52155_new_n3703_; 
wire u2__abc_52155_new_n3704_; 
wire u2__abc_52155_new_n3705_; 
wire u2__abc_52155_new_n3706_; 
wire u2__abc_52155_new_n3707_; 
wire u2__abc_52155_new_n3708_; 
wire u2__abc_52155_new_n3709_; 
wire u2__abc_52155_new_n3710_; 
wire u2__abc_52155_new_n3711_; 
wire u2__abc_52155_new_n3712_; 
wire u2__abc_52155_new_n3713_; 
wire u2__abc_52155_new_n3714_; 
wire u2__abc_52155_new_n3715_; 
wire u2__abc_52155_new_n3716_; 
wire u2__abc_52155_new_n3717_; 
wire u2__abc_52155_new_n3718_; 
wire u2__abc_52155_new_n3719_; 
wire u2__abc_52155_new_n3720_; 
wire u2__abc_52155_new_n3721_; 
wire u2__abc_52155_new_n3722_; 
wire u2__abc_52155_new_n3723_; 
wire u2__abc_52155_new_n3724_; 
wire u2__abc_52155_new_n3725_; 
wire u2__abc_52155_new_n3726_; 
wire u2__abc_52155_new_n3727_; 
wire u2__abc_52155_new_n3728_; 
wire u2__abc_52155_new_n3729_; 
wire u2__abc_52155_new_n3730_; 
wire u2__abc_52155_new_n3731_; 
wire u2__abc_52155_new_n3732_; 
wire u2__abc_52155_new_n3733_; 
wire u2__abc_52155_new_n3734_; 
wire u2__abc_52155_new_n3735_; 
wire u2__abc_52155_new_n3736_; 
wire u2__abc_52155_new_n3737_; 
wire u2__abc_52155_new_n3738_; 
wire u2__abc_52155_new_n3739_; 
wire u2__abc_52155_new_n3740_; 
wire u2__abc_52155_new_n3741_; 
wire u2__abc_52155_new_n3742_; 
wire u2__abc_52155_new_n3743_; 
wire u2__abc_52155_new_n3744_; 
wire u2__abc_52155_new_n3745_; 
wire u2__abc_52155_new_n3746_; 
wire u2__abc_52155_new_n3747_; 
wire u2__abc_52155_new_n3748_; 
wire u2__abc_52155_new_n3749_; 
wire u2__abc_52155_new_n3750_; 
wire u2__abc_52155_new_n3751_; 
wire u2__abc_52155_new_n3752_; 
wire u2__abc_52155_new_n3753_; 
wire u2__abc_52155_new_n3754_; 
wire u2__abc_52155_new_n3755_; 
wire u2__abc_52155_new_n3756_; 
wire u2__abc_52155_new_n3757_; 
wire u2__abc_52155_new_n3758_; 
wire u2__abc_52155_new_n3759_; 
wire u2__abc_52155_new_n3760_; 
wire u2__abc_52155_new_n3761_; 
wire u2__abc_52155_new_n3762_; 
wire u2__abc_52155_new_n3763_; 
wire u2__abc_52155_new_n3764_; 
wire u2__abc_52155_new_n3765_; 
wire u2__abc_52155_new_n3766_; 
wire u2__abc_52155_new_n3767_; 
wire u2__abc_52155_new_n3768_; 
wire u2__abc_52155_new_n3769_; 
wire u2__abc_52155_new_n3770_; 
wire u2__abc_52155_new_n3771_; 
wire u2__abc_52155_new_n3772_; 
wire u2__abc_52155_new_n3773_; 
wire u2__abc_52155_new_n3774_; 
wire u2__abc_52155_new_n3775_; 
wire u2__abc_52155_new_n3776_; 
wire u2__abc_52155_new_n3777_; 
wire u2__abc_52155_new_n3778_; 
wire u2__abc_52155_new_n3779_; 
wire u2__abc_52155_new_n3780_; 
wire u2__abc_52155_new_n3781_; 
wire u2__abc_52155_new_n3782_; 
wire u2__abc_52155_new_n3783_; 
wire u2__abc_52155_new_n3784_; 
wire u2__abc_52155_new_n3785_; 
wire u2__abc_52155_new_n3786_; 
wire u2__abc_52155_new_n3787_; 
wire u2__abc_52155_new_n3788_; 
wire u2__abc_52155_new_n3789_; 
wire u2__abc_52155_new_n3790_; 
wire u2__abc_52155_new_n3791_; 
wire u2__abc_52155_new_n3792_; 
wire u2__abc_52155_new_n3793_; 
wire u2__abc_52155_new_n3794_; 
wire u2__abc_52155_new_n3795_; 
wire u2__abc_52155_new_n3796_; 
wire u2__abc_52155_new_n3797_; 
wire u2__abc_52155_new_n3798_; 
wire u2__abc_52155_new_n3799_; 
wire u2__abc_52155_new_n3800_; 
wire u2__abc_52155_new_n3801_; 
wire u2__abc_52155_new_n3802_; 
wire u2__abc_52155_new_n3803_; 
wire u2__abc_52155_new_n3804_; 
wire u2__abc_52155_new_n3805_; 
wire u2__abc_52155_new_n3806_; 
wire u2__abc_52155_new_n3807_; 
wire u2__abc_52155_new_n3808_; 
wire u2__abc_52155_new_n3809_; 
wire u2__abc_52155_new_n3810_; 
wire u2__abc_52155_new_n3811_; 
wire u2__abc_52155_new_n3812_; 
wire u2__abc_52155_new_n3813_; 
wire u2__abc_52155_new_n3814_; 
wire u2__abc_52155_new_n3815_; 
wire u2__abc_52155_new_n3816_; 
wire u2__abc_52155_new_n3817_; 
wire u2__abc_52155_new_n3818_; 
wire u2__abc_52155_new_n3819_; 
wire u2__abc_52155_new_n3820_; 
wire u2__abc_52155_new_n3821_; 
wire u2__abc_52155_new_n3822_; 
wire u2__abc_52155_new_n3823_; 
wire u2__abc_52155_new_n3824_; 
wire u2__abc_52155_new_n3825_; 
wire u2__abc_52155_new_n3826_; 
wire u2__abc_52155_new_n3827_; 
wire u2__abc_52155_new_n3828_; 
wire u2__abc_52155_new_n3829_; 
wire u2__abc_52155_new_n3830_; 
wire u2__abc_52155_new_n3831_; 
wire u2__abc_52155_new_n3832_; 
wire u2__abc_52155_new_n3833_; 
wire u2__abc_52155_new_n3834_; 
wire u2__abc_52155_new_n3835_; 
wire u2__abc_52155_new_n3836_; 
wire u2__abc_52155_new_n3837_; 
wire u2__abc_52155_new_n3838_; 
wire u2__abc_52155_new_n3839_; 
wire u2__abc_52155_new_n3840_; 
wire u2__abc_52155_new_n3841_; 
wire u2__abc_52155_new_n3842_; 
wire u2__abc_52155_new_n3843_; 
wire u2__abc_52155_new_n3844_; 
wire u2__abc_52155_new_n3845_; 
wire u2__abc_52155_new_n3846_; 
wire u2__abc_52155_new_n3847_; 
wire u2__abc_52155_new_n3848_; 
wire u2__abc_52155_new_n3849_; 
wire u2__abc_52155_new_n3850_; 
wire u2__abc_52155_new_n3851_; 
wire u2__abc_52155_new_n3852_; 
wire u2__abc_52155_new_n3853_; 
wire u2__abc_52155_new_n3854_; 
wire u2__abc_52155_new_n3855_; 
wire u2__abc_52155_new_n3856_; 
wire u2__abc_52155_new_n3857_; 
wire u2__abc_52155_new_n3858_; 
wire u2__abc_52155_new_n3859_; 
wire u2__abc_52155_new_n3860_; 
wire u2__abc_52155_new_n3861_; 
wire u2__abc_52155_new_n3862_; 
wire u2__abc_52155_new_n3863_; 
wire u2__abc_52155_new_n3864_; 
wire u2__abc_52155_new_n3865_; 
wire u2__abc_52155_new_n3866_; 
wire u2__abc_52155_new_n3867_; 
wire u2__abc_52155_new_n3868_; 
wire u2__abc_52155_new_n3869_; 
wire u2__abc_52155_new_n3870_; 
wire u2__abc_52155_new_n3871_; 
wire u2__abc_52155_new_n3872_; 
wire u2__abc_52155_new_n3873_; 
wire u2__abc_52155_new_n3874_; 
wire u2__abc_52155_new_n3875_; 
wire u2__abc_52155_new_n3876_; 
wire u2__abc_52155_new_n3877_; 
wire u2__abc_52155_new_n3878_; 
wire u2__abc_52155_new_n3879_; 
wire u2__abc_52155_new_n3880_; 
wire u2__abc_52155_new_n3881_; 
wire u2__abc_52155_new_n3882_; 
wire u2__abc_52155_new_n3883_; 
wire u2__abc_52155_new_n3884_; 
wire u2__abc_52155_new_n3885_; 
wire u2__abc_52155_new_n3886_; 
wire u2__abc_52155_new_n3887_; 
wire u2__abc_52155_new_n3888_; 
wire u2__abc_52155_new_n3889_; 
wire u2__abc_52155_new_n3890_; 
wire u2__abc_52155_new_n3891_; 
wire u2__abc_52155_new_n3892_; 
wire u2__abc_52155_new_n3893_; 
wire u2__abc_52155_new_n3894_; 
wire u2__abc_52155_new_n3895_; 
wire u2__abc_52155_new_n3896_; 
wire u2__abc_52155_new_n3897_; 
wire u2__abc_52155_new_n3898_; 
wire u2__abc_52155_new_n3899_; 
wire u2__abc_52155_new_n3900_; 
wire u2__abc_52155_new_n3901_; 
wire u2__abc_52155_new_n3902_; 
wire u2__abc_52155_new_n3903_; 
wire u2__abc_52155_new_n3904_; 
wire u2__abc_52155_new_n3905_; 
wire u2__abc_52155_new_n3906_; 
wire u2__abc_52155_new_n3907_; 
wire u2__abc_52155_new_n3908_; 
wire u2__abc_52155_new_n3909_; 
wire u2__abc_52155_new_n3910_; 
wire u2__abc_52155_new_n3911_; 
wire u2__abc_52155_new_n3912_; 
wire u2__abc_52155_new_n3913_; 
wire u2__abc_52155_new_n3914_; 
wire u2__abc_52155_new_n3915_; 
wire u2__abc_52155_new_n3916_; 
wire u2__abc_52155_new_n3917_; 
wire u2__abc_52155_new_n3918_; 
wire u2__abc_52155_new_n3919_; 
wire u2__abc_52155_new_n3920_; 
wire u2__abc_52155_new_n3921_; 
wire u2__abc_52155_new_n3922_; 
wire u2__abc_52155_new_n3923_; 
wire u2__abc_52155_new_n3924_; 
wire u2__abc_52155_new_n3925_; 
wire u2__abc_52155_new_n3926_; 
wire u2__abc_52155_new_n3927_; 
wire u2__abc_52155_new_n3928_; 
wire u2__abc_52155_new_n3929_; 
wire u2__abc_52155_new_n3930_; 
wire u2__abc_52155_new_n3931_; 
wire u2__abc_52155_new_n3932_; 
wire u2__abc_52155_new_n3933_; 
wire u2__abc_52155_new_n3934_; 
wire u2__abc_52155_new_n3935_; 
wire u2__abc_52155_new_n3936_; 
wire u2__abc_52155_new_n3937_; 
wire u2__abc_52155_new_n3938_; 
wire u2__abc_52155_new_n3939_; 
wire u2__abc_52155_new_n3940_; 
wire u2__abc_52155_new_n3941_; 
wire u2__abc_52155_new_n3942_; 
wire u2__abc_52155_new_n3943_; 
wire u2__abc_52155_new_n3944_; 
wire u2__abc_52155_new_n3945_; 
wire u2__abc_52155_new_n3946_; 
wire u2__abc_52155_new_n3947_; 
wire u2__abc_52155_new_n3948_; 
wire u2__abc_52155_new_n3949_; 
wire u2__abc_52155_new_n3950_; 
wire u2__abc_52155_new_n3951_; 
wire u2__abc_52155_new_n3952_; 
wire u2__abc_52155_new_n3953_; 
wire u2__abc_52155_new_n3954_; 
wire u2__abc_52155_new_n3955_; 
wire u2__abc_52155_new_n3956_; 
wire u2__abc_52155_new_n3957_; 
wire u2__abc_52155_new_n3958_; 
wire u2__abc_52155_new_n3959_; 
wire u2__abc_52155_new_n3960_; 
wire u2__abc_52155_new_n3961_; 
wire u2__abc_52155_new_n3962_; 
wire u2__abc_52155_new_n3963_; 
wire u2__abc_52155_new_n3964_; 
wire u2__abc_52155_new_n3965_; 
wire u2__abc_52155_new_n3966_; 
wire u2__abc_52155_new_n3967_; 
wire u2__abc_52155_new_n3968_; 
wire u2__abc_52155_new_n3969_; 
wire u2__abc_52155_new_n3970_; 
wire u2__abc_52155_new_n3971_; 
wire u2__abc_52155_new_n3972_; 
wire u2__abc_52155_new_n3973_; 
wire u2__abc_52155_new_n3974_; 
wire u2__abc_52155_new_n3975_; 
wire u2__abc_52155_new_n3976_; 
wire u2__abc_52155_new_n3977_; 
wire u2__abc_52155_new_n3978_; 
wire u2__abc_52155_new_n3979_; 
wire u2__abc_52155_new_n3980_; 
wire u2__abc_52155_new_n3981_; 
wire u2__abc_52155_new_n3982_; 
wire u2__abc_52155_new_n3983_; 
wire u2__abc_52155_new_n3984_; 
wire u2__abc_52155_new_n3985_; 
wire u2__abc_52155_new_n3986_; 
wire u2__abc_52155_new_n3987_; 
wire u2__abc_52155_new_n3988_; 
wire u2__abc_52155_new_n3989_; 
wire u2__abc_52155_new_n3990_; 
wire u2__abc_52155_new_n3991_; 
wire u2__abc_52155_new_n3992_; 
wire u2__abc_52155_new_n3993_; 
wire u2__abc_52155_new_n3994_; 
wire u2__abc_52155_new_n3995_; 
wire u2__abc_52155_new_n3996_; 
wire u2__abc_52155_new_n3997_; 
wire u2__abc_52155_new_n3998_; 
wire u2__abc_52155_new_n3999_; 
wire u2__abc_52155_new_n4000_; 
wire u2__abc_52155_new_n4001_; 
wire u2__abc_52155_new_n4002_; 
wire u2__abc_52155_new_n4003_; 
wire u2__abc_52155_new_n4004_; 
wire u2__abc_52155_new_n4005_; 
wire u2__abc_52155_new_n4006_; 
wire u2__abc_52155_new_n4007_; 
wire u2__abc_52155_new_n4008_; 
wire u2__abc_52155_new_n4009_; 
wire u2__abc_52155_new_n4010_; 
wire u2__abc_52155_new_n4011_; 
wire u2__abc_52155_new_n4012_; 
wire u2__abc_52155_new_n4013_; 
wire u2__abc_52155_new_n4014_; 
wire u2__abc_52155_new_n4015_; 
wire u2__abc_52155_new_n4016_; 
wire u2__abc_52155_new_n4017_; 
wire u2__abc_52155_new_n4018_; 
wire u2__abc_52155_new_n4019_; 
wire u2__abc_52155_new_n4020_; 
wire u2__abc_52155_new_n4021_; 
wire u2__abc_52155_new_n4022_; 
wire u2__abc_52155_new_n4023_; 
wire u2__abc_52155_new_n4024_; 
wire u2__abc_52155_new_n4025_; 
wire u2__abc_52155_new_n4026_; 
wire u2__abc_52155_new_n4027_; 
wire u2__abc_52155_new_n4028_; 
wire u2__abc_52155_new_n4029_; 
wire u2__abc_52155_new_n4030_; 
wire u2__abc_52155_new_n4031_; 
wire u2__abc_52155_new_n4032_; 
wire u2__abc_52155_new_n4033_; 
wire u2__abc_52155_new_n4034_; 
wire u2__abc_52155_new_n4035_; 
wire u2__abc_52155_new_n4036_; 
wire u2__abc_52155_new_n4037_; 
wire u2__abc_52155_new_n4038_; 
wire u2__abc_52155_new_n4039_; 
wire u2__abc_52155_new_n4040_; 
wire u2__abc_52155_new_n4041_; 
wire u2__abc_52155_new_n4042_; 
wire u2__abc_52155_new_n4043_; 
wire u2__abc_52155_new_n4044_; 
wire u2__abc_52155_new_n4045_; 
wire u2__abc_52155_new_n4046_; 
wire u2__abc_52155_new_n4047_; 
wire u2__abc_52155_new_n4048_; 
wire u2__abc_52155_new_n4049_; 
wire u2__abc_52155_new_n4050_; 
wire u2__abc_52155_new_n4051_; 
wire u2__abc_52155_new_n4052_; 
wire u2__abc_52155_new_n4053_; 
wire u2__abc_52155_new_n4054_; 
wire u2__abc_52155_new_n4055_; 
wire u2__abc_52155_new_n4056_; 
wire u2__abc_52155_new_n4057_; 
wire u2__abc_52155_new_n4058_; 
wire u2__abc_52155_new_n4059_; 
wire u2__abc_52155_new_n4060_; 
wire u2__abc_52155_new_n4061_; 
wire u2__abc_52155_new_n4062_; 
wire u2__abc_52155_new_n4063_; 
wire u2__abc_52155_new_n4064_; 
wire u2__abc_52155_new_n4065_; 
wire u2__abc_52155_new_n4066_; 
wire u2__abc_52155_new_n4067_; 
wire u2__abc_52155_new_n4068_; 
wire u2__abc_52155_new_n4069_; 
wire u2__abc_52155_new_n4070_; 
wire u2__abc_52155_new_n4071_; 
wire u2__abc_52155_new_n4072_; 
wire u2__abc_52155_new_n4073_; 
wire u2__abc_52155_new_n4074_; 
wire u2__abc_52155_new_n4075_; 
wire u2__abc_52155_new_n4076_; 
wire u2__abc_52155_new_n4077_; 
wire u2__abc_52155_new_n4078_; 
wire u2__abc_52155_new_n4079_; 
wire u2__abc_52155_new_n4080_; 
wire u2__abc_52155_new_n4081_; 
wire u2__abc_52155_new_n4082_; 
wire u2__abc_52155_new_n4083_; 
wire u2__abc_52155_new_n4084_; 
wire u2__abc_52155_new_n4085_; 
wire u2__abc_52155_new_n4086_; 
wire u2__abc_52155_new_n4087_; 
wire u2__abc_52155_new_n4088_; 
wire u2__abc_52155_new_n4089_; 
wire u2__abc_52155_new_n4090_; 
wire u2__abc_52155_new_n4091_; 
wire u2__abc_52155_new_n4092_; 
wire u2__abc_52155_new_n4093_; 
wire u2__abc_52155_new_n4094_; 
wire u2__abc_52155_new_n4095_; 
wire u2__abc_52155_new_n4096_; 
wire u2__abc_52155_new_n4097_; 
wire u2__abc_52155_new_n4098_; 
wire u2__abc_52155_new_n4099_; 
wire u2__abc_52155_new_n4100_; 
wire u2__abc_52155_new_n4101_; 
wire u2__abc_52155_new_n4102_; 
wire u2__abc_52155_new_n4103_; 
wire u2__abc_52155_new_n4104_; 
wire u2__abc_52155_new_n4105_; 
wire u2__abc_52155_new_n4106_; 
wire u2__abc_52155_new_n4107_; 
wire u2__abc_52155_new_n4108_; 
wire u2__abc_52155_new_n4109_; 
wire u2__abc_52155_new_n4110_; 
wire u2__abc_52155_new_n4111_; 
wire u2__abc_52155_new_n4112_; 
wire u2__abc_52155_new_n4113_; 
wire u2__abc_52155_new_n4114_; 
wire u2__abc_52155_new_n4115_; 
wire u2__abc_52155_new_n4116_; 
wire u2__abc_52155_new_n4117_; 
wire u2__abc_52155_new_n4118_; 
wire u2__abc_52155_new_n4119_; 
wire u2__abc_52155_new_n4120_; 
wire u2__abc_52155_new_n4121_; 
wire u2__abc_52155_new_n4122_; 
wire u2__abc_52155_new_n4123_; 
wire u2__abc_52155_new_n4124_; 
wire u2__abc_52155_new_n4125_; 
wire u2__abc_52155_new_n4126_; 
wire u2__abc_52155_new_n4127_; 
wire u2__abc_52155_new_n4128_; 
wire u2__abc_52155_new_n4129_; 
wire u2__abc_52155_new_n4130_; 
wire u2__abc_52155_new_n4131_; 
wire u2__abc_52155_new_n4132_; 
wire u2__abc_52155_new_n4133_; 
wire u2__abc_52155_new_n4134_; 
wire u2__abc_52155_new_n4135_; 
wire u2__abc_52155_new_n4136_; 
wire u2__abc_52155_new_n4137_; 
wire u2__abc_52155_new_n4138_; 
wire u2__abc_52155_new_n4139_; 
wire u2__abc_52155_new_n4140_; 
wire u2__abc_52155_new_n4141_; 
wire u2__abc_52155_new_n4142_; 
wire u2__abc_52155_new_n4143_; 
wire u2__abc_52155_new_n4144_; 
wire u2__abc_52155_new_n4145_; 
wire u2__abc_52155_new_n4146_; 
wire u2__abc_52155_new_n4147_; 
wire u2__abc_52155_new_n4148_; 
wire u2__abc_52155_new_n4149_; 
wire u2__abc_52155_new_n4150_; 
wire u2__abc_52155_new_n4151_; 
wire u2__abc_52155_new_n4152_; 
wire u2__abc_52155_new_n4153_; 
wire u2__abc_52155_new_n4154_; 
wire u2__abc_52155_new_n4155_; 
wire u2__abc_52155_new_n4156_; 
wire u2__abc_52155_new_n4157_; 
wire u2__abc_52155_new_n4158_; 
wire u2__abc_52155_new_n4159_; 
wire u2__abc_52155_new_n4160_; 
wire u2__abc_52155_new_n4161_; 
wire u2__abc_52155_new_n4162_; 
wire u2__abc_52155_new_n4163_; 
wire u2__abc_52155_new_n4164_; 
wire u2__abc_52155_new_n4165_; 
wire u2__abc_52155_new_n4166_; 
wire u2__abc_52155_new_n4167_; 
wire u2__abc_52155_new_n4168_; 
wire u2__abc_52155_new_n4169_; 
wire u2__abc_52155_new_n4170_; 
wire u2__abc_52155_new_n4171_; 
wire u2__abc_52155_new_n4172_; 
wire u2__abc_52155_new_n4173_; 
wire u2__abc_52155_new_n4174_; 
wire u2__abc_52155_new_n4175_; 
wire u2__abc_52155_new_n4176_; 
wire u2__abc_52155_new_n4177_; 
wire u2__abc_52155_new_n4178_; 
wire u2__abc_52155_new_n4179_; 
wire u2__abc_52155_new_n4180_; 
wire u2__abc_52155_new_n4181_; 
wire u2__abc_52155_new_n4182_; 
wire u2__abc_52155_new_n4183_; 
wire u2__abc_52155_new_n4184_; 
wire u2__abc_52155_new_n4185_; 
wire u2__abc_52155_new_n4186_; 
wire u2__abc_52155_new_n4187_; 
wire u2__abc_52155_new_n4188_; 
wire u2__abc_52155_new_n4189_; 
wire u2__abc_52155_new_n4190_; 
wire u2__abc_52155_new_n4191_; 
wire u2__abc_52155_new_n4192_; 
wire u2__abc_52155_new_n4193_; 
wire u2__abc_52155_new_n4194_; 
wire u2__abc_52155_new_n4195_; 
wire u2__abc_52155_new_n4196_; 
wire u2__abc_52155_new_n4197_; 
wire u2__abc_52155_new_n4198_; 
wire u2__abc_52155_new_n4199_; 
wire u2__abc_52155_new_n4200_; 
wire u2__abc_52155_new_n4201_; 
wire u2__abc_52155_new_n4202_; 
wire u2__abc_52155_new_n4203_; 
wire u2__abc_52155_new_n4204_; 
wire u2__abc_52155_new_n4205_; 
wire u2__abc_52155_new_n4206_; 
wire u2__abc_52155_new_n4207_; 
wire u2__abc_52155_new_n4208_; 
wire u2__abc_52155_new_n4209_; 
wire u2__abc_52155_new_n4210_; 
wire u2__abc_52155_new_n4211_; 
wire u2__abc_52155_new_n4212_; 
wire u2__abc_52155_new_n4213_; 
wire u2__abc_52155_new_n4214_; 
wire u2__abc_52155_new_n4215_; 
wire u2__abc_52155_new_n4216_; 
wire u2__abc_52155_new_n4217_; 
wire u2__abc_52155_new_n4218_; 
wire u2__abc_52155_new_n4219_; 
wire u2__abc_52155_new_n4220_; 
wire u2__abc_52155_new_n4221_; 
wire u2__abc_52155_new_n4222_; 
wire u2__abc_52155_new_n4223_; 
wire u2__abc_52155_new_n4224_; 
wire u2__abc_52155_new_n4225_; 
wire u2__abc_52155_new_n4226_; 
wire u2__abc_52155_new_n4227_; 
wire u2__abc_52155_new_n4228_; 
wire u2__abc_52155_new_n4229_; 
wire u2__abc_52155_new_n4230_; 
wire u2__abc_52155_new_n4231_; 
wire u2__abc_52155_new_n4232_; 
wire u2__abc_52155_new_n4233_; 
wire u2__abc_52155_new_n4234_; 
wire u2__abc_52155_new_n4235_; 
wire u2__abc_52155_new_n4236_; 
wire u2__abc_52155_new_n4237_; 
wire u2__abc_52155_new_n4238_; 
wire u2__abc_52155_new_n4239_; 
wire u2__abc_52155_new_n4240_; 
wire u2__abc_52155_new_n4241_; 
wire u2__abc_52155_new_n4242_; 
wire u2__abc_52155_new_n4243_; 
wire u2__abc_52155_new_n4244_; 
wire u2__abc_52155_new_n4245_; 
wire u2__abc_52155_new_n4246_; 
wire u2__abc_52155_new_n4247_; 
wire u2__abc_52155_new_n4248_; 
wire u2__abc_52155_new_n4249_; 
wire u2__abc_52155_new_n4250_; 
wire u2__abc_52155_new_n4251_; 
wire u2__abc_52155_new_n4252_; 
wire u2__abc_52155_new_n4253_; 
wire u2__abc_52155_new_n4254_; 
wire u2__abc_52155_new_n4255_; 
wire u2__abc_52155_new_n4256_; 
wire u2__abc_52155_new_n4257_; 
wire u2__abc_52155_new_n4258_; 
wire u2__abc_52155_new_n4259_; 
wire u2__abc_52155_new_n4260_; 
wire u2__abc_52155_new_n4261_; 
wire u2__abc_52155_new_n4262_; 
wire u2__abc_52155_new_n4263_; 
wire u2__abc_52155_new_n4264_; 
wire u2__abc_52155_new_n4265_; 
wire u2__abc_52155_new_n4266_; 
wire u2__abc_52155_new_n4267_; 
wire u2__abc_52155_new_n4268_; 
wire u2__abc_52155_new_n4269_; 
wire u2__abc_52155_new_n4270_; 
wire u2__abc_52155_new_n4271_; 
wire u2__abc_52155_new_n4272_; 
wire u2__abc_52155_new_n4273_; 
wire u2__abc_52155_new_n4274_; 
wire u2__abc_52155_new_n4275_; 
wire u2__abc_52155_new_n4276_; 
wire u2__abc_52155_new_n4277_; 
wire u2__abc_52155_new_n4278_; 
wire u2__abc_52155_new_n4279_; 
wire u2__abc_52155_new_n4280_; 
wire u2__abc_52155_new_n4281_; 
wire u2__abc_52155_new_n4282_; 
wire u2__abc_52155_new_n4283_; 
wire u2__abc_52155_new_n4284_; 
wire u2__abc_52155_new_n4285_; 
wire u2__abc_52155_new_n4286_; 
wire u2__abc_52155_new_n4287_; 
wire u2__abc_52155_new_n4288_; 
wire u2__abc_52155_new_n4289_; 
wire u2__abc_52155_new_n4290_; 
wire u2__abc_52155_new_n4291_; 
wire u2__abc_52155_new_n4292_; 
wire u2__abc_52155_new_n4293_; 
wire u2__abc_52155_new_n4294_; 
wire u2__abc_52155_new_n4295_; 
wire u2__abc_52155_new_n4296_; 
wire u2__abc_52155_new_n4297_; 
wire u2__abc_52155_new_n4298_; 
wire u2__abc_52155_new_n4299_; 
wire u2__abc_52155_new_n4300_; 
wire u2__abc_52155_new_n4301_; 
wire u2__abc_52155_new_n4302_; 
wire u2__abc_52155_new_n4303_; 
wire u2__abc_52155_new_n4304_; 
wire u2__abc_52155_new_n4305_; 
wire u2__abc_52155_new_n4306_; 
wire u2__abc_52155_new_n4307_; 
wire u2__abc_52155_new_n4308_; 
wire u2__abc_52155_new_n4309_; 
wire u2__abc_52155_new_n4310_; 
wire u2__abc_52155_new_n4311_; 
wire u2__abc_52155_new_n4312_; 
wire u2__abc_52155_new_n4313_; 
wire u2__abc_52155_new_n4314_; 
wire u2__abc_52155_new_n4315_; 
wire u2__abc_52155_new_n4316_; 
wire u2__abc_52155_new_n4317_; 
wire u2__abc_52155_new_n4318_; 
wire u2__abc_52155_new_n4319_; 
wire u2__abc_52155_new_n4320_; 
wire u2__abc_52155_new_n4321_; 
wire u2__abc_52155_new_n4322_; 
wire u2__abc_52155_new_n4323_; 
wire u2__abc_52155_new_n4324_; 
wire u2__abc_52155_new_n4325_; 
wire u2__abc_52155_new_n4326_; 
wire u2__abc_52155_new_n4327_; 
wire u2__abc_52155_new_n4328_; 
wire u2__abc_52155_new_n4329_; 
wire u2__abc_52155_new_n4330_; 
wire u2__abc_52155_new_n4331_; 
wire u2__abc_52155_new_n4332_; 
wire u2__abc_52155_new_n4333_; 
wire u2__abc_52155_new_n4334_; 
wire u2__abc_52155_new_n4335_; 
wire u2__abc_52155_new_n4336_; 
wire u2__abc_52155_new_n4337_; 
wire u2__abc_52155_new_n4338_; 
wire u2__abc_52155_new_n4339_; 
wire u2__abc_52155_new_n4340_; 
wire u2__abc_52155_new_n4341_; 
wire u2__abc_52155_new_n4342_; 
wire u2__abc_52155_new_n4343_; 
wire u2__abc_52155_new_n4344_; 
wire u2__abc_52155_new_n4345_; 
wire u2__abc_52155_new_n4346_; 
wire u2__abc_52155_new_n4347_; 
wire u2__abc_52155_new_n4348_; 
wire u2__abc_52155_new_n4349_; 
wire u2__abc_52155_new_n4350_; 
wire u2__abc_52155_new_n4351_; 
wire u2__abc_52155_new_n4352_; 
wire u2__abc_52155_new_n4353_; 
wire u2__abc_52155_new_n4354_; 
wire u2__abc_52155_new_n4355_; 
wire u2__abc_52155_new_n4356_; 
wire u2__abc_52155_new_n4357_; 
wire u2__abc_52155_new_n4358_; 
wire u2__abc_52155_new_n4359_; 
wire u2__abc_52155_new_n4360_; 
wire u2__abc_52155_new_n4361_; 
wire u2__abc_52155_new_n4362_; 
wire u2__abc_52155_new_n4363_; 
wire u2__abc_52155_new_n4364_; 
wire u2__abc_52155_new_n4365_; 
wire u2__abc_52155_new_n4366_; 
wire u2__abc_52155_new_n4367_; 
wire u2__abc_52155_new_n4368_; 
wire u2__abc_52155_new_n4369_; 
wire u2__abc_52155_new_n4370_; 
wire u2__abc_52155_new_n4371_; 
wire u2__abc_52155_new_n4372_; 
wire u2__abc_52155_new_n4373_; 
wire u2__abc_52155_new_n4374_; 
wire u2__abc_52155_new_n4375_; 
wire u2__abc_52155_new_n4376_; 
wire u2__abc_52155_new_n4377_; 
wire u2__abc_52155_new_n4378_; 
wire u2__abc_52155_new_n4379_; 
wire u2__abc_52155_new_n4380_; 
wire u2__abc_52155_new_n4381_; 
wire u2__abc_52155_new_n4382_; 
wire u2__abc_52155_new_n4383_; 
wire u2__abc_52155_new_n4384_; 
wire u2__abc_52155_new_n4385_; 
wire u2__abc_52155_new_n4386_; 
wire u2__abc_52155_new_n4387_; 
wire u2__abc_52155_new_n4388_; 
wire u2__abc_52155_new_n4389_; 
wire u2__abc_52155_new_n4390_; 
wire u2__abc_52155_new_n4391_; 
wire u2__abc_52155_new_n4392_; 
wire u2__abc_52155_new_n4393_; 
wire u2__abc_52155_new_n4394_; 
wire u2__abc_52155_new_n4395_; 
wire u2__abc_52155_new_n4396_; 
wire u2__abc_52155_new_n4397_; 
wire u2__abc_52155_new_n4398_; 
wire u2__abc_52155_new_n4399_; 
wire u2__abc_52155_new_n4400_; 
wire u2__abc_52155_new_n4401_; 
wire u2__abc_52155_new_n4402_; 
wire u2__abc_52155_new_n4403_; 
wire u2__abc_52155_new_n4404_; 
wire u2__abc_52155_new_n4405_; 
wire u2__abc_52155_new_n4406_; 
wire u2__abc_52155_new_n4407_; 
wire u2__abc_52155_new_n4408_; 
wire u2__abc_52155_new_n4409_; 
wire u2__abc_52155_new_n4410_; 
wire u2__abc_52155_new_n4411_; 
wire u2__abc_52155_new_n4412_; 
wire u2__abc_52155_new_n4413_; 
wire u2__abc_52155_new_n4414_; 
wire u2__abc_52155_new_n4415_; 
wire u2__abc_52155_new_n4416_; 
wire u2__abc_52155_new_n4417_; 
wire u2__abc_52155_new_n4418_; 
wire u2__abc_52155_new_n4419_; 
wire u2__abc_52155_new_n4420_; 
wire u2__abc_52155_new_n4421_; 
wire u2__abc_52155_new_n4422_; 
wire u2__abc_52155_new_n4423_; 
wire u2__abc_52155_new_n4424_; 
wire u2__abc_52155_new_n4425_; 
wire u2__abc_52155_new_n4426_; 
wire u2__abc_52155_new_n4427_; 
wire u2__abc_52155_new_n4428_; 
wire u2__abc_52155_new_n4429_; 
wire u2__abc_52155_new_n4430_; 
wire u2__abc_52155_new_n4431_; 
wire u2__abc_52155_new_n4432_; 
wire u2__abc_52155_new_n4433_; 
wire u2__abc_52155_new_n4434_; 
wire u2__abc_52155_new_n4435_; 
wire u2__abc_52155_new_n4436_; 
wire u2__abc_52155_new_n4437_; 
wire u2__abc_52155_new_n4438_; 
wire u2__abc_52155_new_n4439_; 
wire u2__abc_52155_new_n4440_; 
wire u2__abc_52155_new_n4441_; 
wire u2__abc_52155_new_n4442_; 
wire u2__abc_52155_new_n4443_; 
wire u2__abc_52155_new_n4444_; 
wire u2__abc_52155_new_n4445_; 
wire u2__abc_52155_new_n4446_; 
wire u2__abc_52155_new_n4447_; 
wire u2__abc_52155_new_n4448_; 
wire u2__abc_52155_new_n4449_; 
wire u2__abc_52155_new_n4450_; 
wire u2__abc_52155_new_n4451_; 
wire u2__abc_52155_new_n4452_; 
wire u2__abc_52155_new_n4453_; 
wire u2__abc_52155_new_n4454_; 
wire u2__abc_52155_new_n4455_; 
wire u2__abc_52155_new_n4456_; 
wire u2__abc_52155_new_n4457_; 
wire u2__abc_52155_new_n4458_; 
wire u2__abc_52155_new_n4459_; 
wire u2__abc_52155_new_n4460_; 
wire u2__abc_52155_new_n4461_; 
wire u2__abc_52155_new_n4462_; 
wire u2__abc_52155_new_n4463_; 
wire u2__abc_52155_new_n4464_; 
wire u2__abc_52155_new_n4465_; 
wire u2__abc_52155_new_n4466_; 
wire u2__abc_52155_new_n4467_; 
wire u2__abc_52155_new_n4468_; 
wire u2__abc_52155_new_n4469_; 
wire u2__abc_52155_new_n4470_; 
wire u2__abc_52155_new_n4471_; 
wire u2__abc_52155_new_n4472_; 
wire u2__abc_52155_new_n4473_; 
wire u2__abc_52155_new_n4474_; 
wire u2__abc_52155_new_n4475_; 
wire u2__abc_52155_new_n4476_; 
wire u2__abc_52155_new_n4477_; 
wire u2__abc_52155_new_n4478_; 
wire u2__abc_52155_new_n4479_; 
wire u2__abc_52155_new_n4480_; 
wire u2__abc_52155_new_n4481_; 
wire u2__abc_52155_new_n4482_; 
wire u2__abc_52155_new_n4483_; 
wire u2__abc_52155_new_n4484_; 
wire u2__abc_52155_new_n4485_; 
wire u2__abc_52155_new_n4486_; 
wire u2__abc_52155_new_n4487_; 
wire u2__abc_52155_new_n4488_; 
wire u2__abc_52155_new_n4489_; 
wire u2__abc_52155_new_n4490_; 
wire u2__abc_52155_new_n4491_; 
wire u2__abc_52155_new_n4492_; 
wire u2__abc_52155_new_n4493_; 
wire u2__abc_52155_new_n4494_; 
wire u2__abc_52155_new_n4495_; 
wire u2__abc_52155_new_n4496_; 
wire u2__abc_52155_new_n4497_; 
wire u2__abc_52155_new_n4498_; 
wire u2__abc_52155_new_n4499_; 
wire u2__abc_52155_new_n4500_; 
wire u2__abc_52155_new_n4501_; 
wire u2__abc_52155_new_n4502_; 
wire u2__abc_52155_new_n4503_; 
wire u2__abc_52155_new_n4504_; 
wire u2__abc_52155_new_n4505_; 
wire u2__abc_52155_new_n4506_; 
wire u2__abc_52155_new_n4507_; 
wire u2__abc_52155_new_n4508_; 
wire u2__abc_52155_new_n4509_; 
wire u2__abc_52155_new_n4510_; 
wire u2__abc_52155_new_n4511_; 
wire u2__abc_52155_new_n4512_; 
wire u2__abc_52155_new_n4513_; 
wire u2__abc_52155_new_n4514_; 
wire u2__abc_52155_new_n4515_; 
wire u2__abc_52155_new_n4516_; 
wire u2__abc_52155_new_n4517_; 
wire u2__abc_52155_new_n4518_; 
wire u2__abc_52155_new_n4519_; 
wire u2__abc_52155_new_n4520_; 
wire u2__abc_52155_new_n4521_; 
wire u2__abc_52155_new_n4522_; 
wire u2__abc_52155_new_n4523_; 
wire u2__abc_52155_new_n4524_; 
wire u2__abc_52155_new_n4525_; 
wire u2__abc_52155_new_n4526_; 
wire u2__abc_52155_new_n4527_; 
wire u2__abc_52155_new_n4528_; 
wire u2__abc_52155_new_n4529_; 
wire u2__abc_52155_new_n4530_; 
wire u2__abc_52155_new_n4531_; 
wire u2__abc_52155_new_n4532_; 
wire u2__abc_52155_new_n4533_; 
wire u2__abc_52155_new_n4534_; 
wire u2__abc_52155_new_n4535_; 
wire u2__abc_52155_new_n4536_; 
wire u2__abc_52155_new_n4537_; 
wire u2__abc_52155_new_n4538_; 
wire u2__abc_52155_new_n4539_; 
wire u2__abc_52155_new_n4540_; 
wire u2__abc_52155_new_n4541_; 
wire u2__abc_52155_new_n4542_; 
wire u2__abc_52155_new_n4543_; 
wire u2__abc_52155_new_n4544_; 
wire u2__abc_52155_new_n4545_; 
wire u2__abc_52155_new_n4546_; 
wire u2__abc_52155_new_n4547_; 
wire u2__abc_52155_new_n4548_; 
wire u2__abc_52155_new_n4549_; 
wire u2__abc_52155_new_n4550_; 
wire u2__abc_52155_new_n4551_; 
wire u2__abc_52155_new_n4552_; 
wire u2__abc_52155_new_n4553_; 
wire u2__abc_52155_new_n4554_; 
wire u2__abc_52155_new_n4555_; 
wire u2__abc_52155_new_n4556_; 
wire u2__abc_52155_new_n4557_; 
wire u2__abc_52155_new_n4558_; 
wire u2__abc_52155_new_n4559_; 
wire u2__abc_52155_new_n4560_; 
wire u2__abc_52155_new_n4561_; 
wire u2__abc_52155_new_n4562_; 
wire u2__abc_52155_new_n4563_; 
wire u2__abc_52155_new_n4564_; 
wire u2__abc_52155_new_n4565_; 
wire u2__abc_52155_new_n4566_; 
wire u2__abc_52155_new_n4567_; 
wire u2__abc_52155_new_n4568_; 
wire u2__abc_52155_new_n4569_; 
wire u2__abc_52155_new_n4570_; 
wire u2__abc_52155_new_n4571_; 
wire u2__abc_52155_new_n4572_; 
wire u2__abc_52155_new_n4573_; 
wire u2__abc_52155_new_n4574_; 
wire u2__abc_52155_new_n4575_; 
wire u2__abc_52155_new_n4576_; 
wire u2__abc_52155_new_n4577_; 
wire u2__abc_52155_new_n4578_; 
wire u2__abc_52155_new_n4579_; 
wire u2__abc_52155_new_n4580_; 
wire u2__abc_52155_new_n4581_; 
wire u2__abc_52155_new_n4582_; 
wire u2__abc_52155_new_n4583_; 
wire u2__abc_52155_new_n4584_; 
wire u2__abc_52155_new_n4585_; 
wire u2__abc_52155_new_n4586_; 
wire u2__abc_52155_new_n4587_; 
wire u2__abc_52155_new_n4588_; 
wire u2__abc_52155_new_n4589_; 
wire u2__abc_52155_new_n4590_; 
wire u2__abc_52155_new_n4591_; 
wire u2__abc_52155_new_n4592_; 
wire u2__abc_52155_new_n4593_; 
wire u2__abc_52155_new_n4594_; 
wire u2__abc_52155_new_n4595_; 
wire u2__abc_52155_new_n4596_; 
wire u2__abc_52155_new_n4597_; 
wire u2__abc_52155_new_n4598_; 
wire u2__abc_52155_new_n4599_; 
wire u2__abc_52155_new_n4600_; 
wire u2__abc_52155_new_n4601_; 
wire u2__abc_52155_new_n4602_; 
wire u2__abc_52155_new_n4603_; 
wire u2__abc_52155_new_n4604_; 
wire u2__abc_52155_new_n4605_; 
wire u2__abc_52155_new_n4606_; 
wire u2__abc_52155_new_n4607_; 
wire u2__abc_52155_new_n4608_; 
wire u2__abc_52155_new_n4609_; 
wire u2__abc_52155_new_n4610_; 
wire u2__abc_52155_new_n4611_; 
wire u2__abc_52155_new_n4612_; 
wire u2__abc_52155_new_n4613_; 
wire u2__abc_52155_new_n4614_; 
wire u2__abc_52155_new_n4615_; 
wire u2__abc_52155_new_n4616_; 
wire u2__abc_52155_new_n4617_; 
wire u2__abc_52155_new_n4618_; 
wire u2__abc_52155_new_n4619_; 
wire u2__abc_52155_new_n4620_; 
wire u2__abc_52155_new_n4621_; 
wire u2__abc_52155_new_n4622_; 
wire u2__abc_52155_new_n4623_; 
wire u2__abc_52155_new_n4624_; 
wire u2__abc_52155_new_n4625_; 
wire u2__abc_52155_new_n4626_; 
wire u2__abc_52155_new_n4627_; 
wire u2__abc_52155_new_n4628_; 
wire u2__abc_52155_new_n4629_; 
wire u2__abc_52155_new_n4630_; 
wire u2__abc_52155_new_n4631_; 
wire u2__abc_52155_new_n4632_; 
wire u2__abc_52155_new_n4633_; 
wire u2__abc_52155_new_n4634_; 
wire u2__abc_52155_new_n4635_; 
wire u2__abc_52155_new_n4636_; 
wire u2__abc_52155_new_n4637_; 
wire u2__abc_52155_new_n4638_; 
wire u2__abc_52155_new_n4639_; 
wire u2__abc_52155_new_n4640_; 
wire u2__abc_52155_new_n4641_; 
wire u2__abc_52155_new_n4642_; 
wire u2__abc_52155_new_n4643_; 
wire u2__abc_52155_new_n4644_; 
wire u2__abc_52155_new_n4645_; 
wire u2__abc_52155_new_n4646_; 
wire u2__abc_52155_new_n4647_; 
wire u2__abc_52155_new_n4648_; 
wire u2__abc_52155_new_n4649_; 
wire u2__abc_52155_new_n4650_; 
wire u2__abc_52155_new_n4651_; 
wire u2__abc_52155_new_n4652_; 
wire u2__abc_52155_new_n4653_; 
wire u2__abc_52155_new_n4654_; 
wire u2__abc_52155_new_n4655_; 
wire u2__abc_52155_new_n4656_; 
wire u2__abc_52155_new_n4657_; 
wire u2__abc_52155_new_n4658_; 
wire u2__abc_52155_new_n4659_; 
wire u2__abc_52155_new_n4660_; 
wire u2__abc_52155_new_n4661_; 
wire u2__abc_52155_new_n4662_; 
wire u2__abc_52155_new_n4663_; 
wire u2__abc_52155_new_n4664_; 
wire u2__abc_52155_new_n4665_; 
wire u2__abc_52155_new_n4666_; 
wire u2__abc_52155_new_n4667_; 
wire u2__abc_52155_new_n4668_; 
wire u2__abc_52155_new_n4669_; 
wire u2__abc_52155_new_n4670_; 
wire u2__abc_52155_new_n4671_; 
wire u2__abc_52155_new_n4672_; 
wire u2__abc_52155_new_n4673_; 
wire u2__abc_52155_new_n4674_; 
wire u2__abc_52155_new_n4675_; 
wire u2__abc_52155_new_n4676_; 
wire u2__abc_52155_new_n4677_; 
wire u2__abc_52155_new_n4678_; 
wire u2__abc_52155_new_n4679_; 
wire u2__abc_52155_new_n4680_; 
wire u2__abc_52155_new_n4681_; 
wire u2__abc_52155_new_n4682_; 
wire u2__abc_52155_new_n4683_; 
wire u2__abc_52155_new_n4684_; 
wire u2__abc_52155_new_n4685_; 
wire u2__abc_52155_new_n4686_; 
wire u2__abc_52155_new_n4687_; 
wire u2__abc_52155_new_n4688_; 
wire u2__abc_52155_new_n4689_; 
wire u2__abc_52155_new_n4690_; 
wire u2__abc_52155_new_n4691_; 
wire u2__abc_52155_new_n4692_; 
wire u2__abc_52155_new_n4693_; 
wire u2__abc_52155_new_n4694_; 
wire u2__abc_52155_new_n4695_; 
wire u2__abc_52155_new_n4696_; 
wire u2__abc_52155_new_n4697_; 
wire u2__abc_52155_new_n4698_; 
wire u2__abc_52155_new_n4699_; 
wire u2__abc_52155_new_n4700_; 
wire u2__abc_52155_new_n4701_; 
wire u2__abc_52155_new_n4702_; 
wire u2__abc_52155_new_n4703_; 
wire u2__abc_52155_new_n4704_; 
wire u2__abc_52155_new_n4705_; 
wire u2__abc_52155_new_n4706_; 
wire u2__abc_52155_new_n4707_; 
wire u2__abc_52155_new_n4708_; 
wire u2__abc_52155_new_n4709_; 
wire u2__abc_52155_new_n4710_; 
wire u2__abc_52155_new_n4711_; 
wire u2__abc_52155_new_n4712_; 
wire u2__abc_52155_new_n4713_; 
wire u2__abc_52155_new_n4714_; 
wire u2__abc_52155_new_n4715_; 
wire u2__abc_52155_new_n4716_; 
wire u2__abc_52155_new_n4717_; 
wire u2__abc_52155_new_n4718_; 
wire u2__abc_52155_new_n4719_; 
wire u2__abc_52155_new_n4720_; 
wire u2__abc_52155_new_n4721_; 
wire u2__abc_52155_new_n4722_; 
wire u2__abc_52155_new_n4723_; 
wire u2__abc_52155_new_n4724_; 
wire u2__abc_52155_new_n4725_; 
wire u2__abc_52155_new_n4726_; 
wire u2__abc_52155_new_n4727_; 
wire u2__abc_52155_new_n4728_; 
wire u2__abc_52155_new_n4729_; 
wire u2__abc_52155_new_n4730_; 
wire u2__abc_52155_new_n4731_; 
wire u2__abc_52155_new_n4732_; 
wire u2__abc_52155_new_n4733_; 
wire u2__abc_52155_new_n4734_; 
wire u2__abc_52155_new_n4735_; 
wire u2__abc_52155_new_n4736_; 
wire u2__abc_52155_new_n4737_; 
wire u2__abc_52155_new_n4738_; 
wire u2__abc_52155_new_n4739_; 
wire u2__abc_52155_new_n4740_; 
wire u2__abc_52155_new_n4741_; 
wire u2__abc_52155_new_n4742_; 
wire u2__abc_52155_new_n4743_; 
wire u2__abc_52155_new_n4744_; 
wire u2__abc_52155_new_n4745_; 
wire u2__abc_52155_new_n4746_; 
wire u2__abc_52155_new_n4747_; 
wire u2__abc_52155_new_n4748_; 
wire u2__abc_52155_new_n4749_; 
wire u2__abc_52155_new_n4750_; 
wire u2__abc_52155_new_n4751_; 
wire u2__abc_52155_new_n4752_; 
wire u2__abc_52155_new_n4753_; 
wire u2__abc_52155_new_n4754_; 
wire u2__abc_52155_new_n4755_; 
wire u2__abc_52155_new_n4756_; 
wire u2__abc_52155_new_n4757_; 
wire u2__abc_52155_new_n4758_; 
wire u2__abc_52155_new_n4759_; 
wire u2__abc_52155_new_n4760_; 
wire u2__abc_52155_new_n4761_; 
wire u2__abc_52155_new_n4762_; 
wire u2__abc_52155_new_n4763_; 
wire u2__abc_52155_new_n4764_; 
wire u2__abc_52155_new_n4765_; 
wire u2__abc_52155_new_n4766_; 
wire u2__abc_52155_new_n4767_; 
wire u2__abc_52155_new_n4768_; 
wire u2__abc_52155_new_n4769_; 
wire u2__abc_52155_new_n4770_; 
wire u2__abc_52155_new_n4771_; 
wire u2__abc_52155_new_n4772_; 
wire u2__abc_52155_new_n4773_; 
wire u2__abc_52155_new_n4774_; 
wire u2__abc_52155_new_n4775_; 
wire u2__abc_52155_new_n4776_; 
wire u2__abc_52155_new_n4777_; 
wire u2__abc_52155_new_n4778_; 
wire u2__abc_52155_new_n4779_; 
wire u2__abc_52155_new_n4780_; 
wire u2__abc_52155_new_n4781_; 
wire u2__abc_52155_new_n4782_; 
wire u2__abc_52155_new_n4783_; 
wire u2__abc_52155_new_n4784_; 
wire u2__abc_52155_new_n4785_; 
wire u2__abc_52155_new_n4786_; 
wire u2__abc_52155_new_n4787_; 
wire u2__abc_52155_new_n4788_; 
wire u2__abc_52155_new_n4789_; 
wire u2__abc_52155_new_n4790_; 
wire u2__abc_52155_new_n4791_; 
wire u2__abc_52155_new_n4792_; 
wire u2__abc_52155_new_n4793_; 
wire u2__abc_52155_new_n4794_; 
wire u2__abc_52155_new_n4795_; 
wire u2__abc_52155_new_n4796_; 
wire u2__abc_52155_new_n4797_; 
wire u2__abc_52155_new_n4798_; 
wire u2__abc_52155_new_n4799_; 
wire u2__abc_52155_new_n4800_; 
wire u2__abc_52155_new_n4801_; 
wire u2__abc_52155_new_n4802_; 
wire u2__abc_52155_new_n4803_; 
wire u2__abc_52155_new_n4804_; 
wire u2__abc_52155_new_n4805_; 
wire u2__abc_52155_new_n4806_; 
wire u2__abc_52155_new_n4807_; 
wire u2__abc_52155_new_n4808_; 
wire u2__abc_52155_new_n4809_; 
wire u2__abc_52155_new_n4810_; 
wire u2__abc_52155_new_n4811_; 
wire u2__abc_52155_new_n4812_; 
wire u2__abc_52155_new_n4813_; 
wire u2__abc_52155_new_n4814_; 
wire u2__abc_52155_new_n4815_; 
wire u2__abc_52155_new_n4816_; 
wire u2__abc_52155_new_n4817_; 
wire u2__abc_52155_new_n4818_; 
wire u2__abc_52155_new_n4819_; 
wire u2__abc_52155_new_n4820_; 
wire u2__abc_52155_new_n4821_; 
wire u2__abc_52155_new_n4822_; 
wire u2__abc_52155_new_n4823_; 
wire u2__abc_52155_new_n4824_; 
wire u2__abc_52155_new_n4825_; 
wire u2__abc_52155_new_n4826_; 
wire u2__abc_52155_new_n4827_; 
wire u2__abc_52155_new_n4828_; 
wire u2__abc_52155_new_n4829_; 
wire u2__abc_52155_new_n4830_; 
wire u2__abc_52155_new_n4831_; 
wire u2__abc_52155_new_n4832_; 
wire u2__abc_52155_new_n4833_; 
wire u2__abc_52155_new_n4834_; 
wire u2__abc_52155_new_n4835_; 
wire u2__abc_52155_new_n4836_; 
wire u2__abc_52155_new_n4837_; 
wire u2__abc_52155_new_n4838_; 
wire u2__abc_52155_new_n4839_; 
wire u2__abc_52155_new_n4840_; 
wire u2__abc_52155_new_n4841_; 
wire u2__abc_52155_new_n4842_; 
wire u2__abc_52155_new_n4843_; 
wire u2__abc_52155_new_n4844_; 
wire u2__abc_52155_new_n4845_; 
wire u2__abc_52155_new_n4846_; 
wire u2__abc_52155_new_n4847_; 
wire u2__abc_52155_new_n4848_; 
wire u2__abc_52155_new_n4849_; 
wire u2__abc_52155_new_n4850_; 
wire u2__abc_52155_new_n4851_; 
wire u2__abc_52155_new_n4852_; 
wire u2__abc_52155_new_n4853_; 
wire u2__abc_52155_new_n4854_; 
wire u2__abc_52155_new_n4855_; 
wire u2__abc_52155_new_n4856_; 
wire u2__abc_52155_new_n4857_; 
wire u2__abc_52155_new_n4858_; 
wire u2__abc_52155_new_n4859_; 
wire u2__abc_52155_new_n4860_; 
wire u2__abc_52155_new_n4861_; 
wire u2__abc_52155_new_n4862_; 
wire u2__abc_52155_new_n4863_; 
wire u2__abc_52155_new_n4864_; 
wire u2__abc_52155_new_n4865_; 
wire u2__abc_52155_new_n4866_; 
wire u2__abc_52155_new_n4867_; 
wire u2__abc_52155_new_n4868_; 
wire u2__abc_52155_new_n4869_; 
wire u2__abc_52155_new_n4870_; 
wire u2__abc_52155_new_n4871_; 
wire u2__abc_52155_new_n4872_; 
wire u2__abc_52155_new_n4873_; 
wire u2__abc_52155_new_n4874_; 
wire u2__abc_52155_new_n4875_; 
wire u2__abc_52155_new_n4876_; 
wire u2__abc_52155_new_n4877_; 
wire u2__abc_52155_new_n4878_; 
wire u2__abc_52155_new_n4879_; 
wire u2__abc_52155_new_n4880_; 
wire u2__abc_52155_new_n4881_; 
wire u2__abc_52155_new_n4882_; 
wire u2__abc_52155_new_n4883_; 
wire u2__abc_52155_new_n4884_; 
wire u2__abc_52155_new_n4885_; 
wire u2__abc_52155_new_n4886_; 
wire u2__abc_52155_new_n4887_; 
wire u2__abc_52155_new_n4888_; 
wire u2__abc_52155_new_n4889_; 
wire u2__abc_52155_new_n4890_; 
wire u2__abc_52155_new_n4891_; 
wire u2__abc_52155_new_n4892_; 
wire u2__abc_52155_new_n4893_; 
wire u2__abc_52155_new_n4894_; 
wire u2__abc_52155_new_n4895_; 
wire u2__abc_52155_new_n4896_; 
wire u2__abc_52155_new_n4897_; 
wire u2__abc_52155_new_n4898_; 
wire u2__abc_52155_new_n4899_; 
wire u2__abc_52155_new_n4900_; 
wire u2__abc_52155_new_n4901_; 
wire u2__abc_52155_new_n4902_; 
wire u2__abc_52155_new_n4903_; 
wire u2__abc_52155_new_n4904_; 
wire u2__abc_52155_new_n4905_; 
wire u2__abc_52155_new_n4906_; 
wire u2__abc_52155_new_n4907_; 
wire u2__abc_52155_new_n4908_; 
wire u2__abc_52155_new_n4909_; 
wire u2__abc_52155_new_n4910_; 
wire u2__abc_52155_new_n4911_; 
wire u2__abc_52155_new_n4912_; 
wire u2__abc_52155_new_n4913_; 
wire u2__abc_52155_new_n4914_; 
wire u2__abc_52155_new_n4915_; 
wire u2__abc_52155_new_n4916_; 
wire u2__abc_52155_new_n4917_; 
wire u2__abc_52155_new_n4918_; 
wire u2__abc_52155_new_n4919_; 
wire u2__abc_52155_new_n4920_; 
wire u2__abc_52155_new_n4921_; 
wire u2__abc_52155_new_n4922_; 
wire u2__abc_52155_new_n4923_; 
wire u2__abc_52155_new_n4924_; 
wire u2__abc_52155_new_n4925_; 
wire u2__abc_52155_new_n4926_; 
wire u2__abc_52155_new_n4927_; 
wire u2__abc_52155_new_n4928_; 
wire u2__abc_52155_new_n4929_; 
wire u2__abc_52155_new_n4930_; 
wire u2__abc_52155_new_n4931_; 
wire u2__abc_52155_new_n4932_; 
wire u2__abc_52155_new_n4933_; 
wire u2__abc_52155_new_n4934_; 
wire u2__abc_52155_new_n4935_; 
wire u2__abc_52155_new_n4936_; 
wire u2__abc_52155_new_n4937_; 
wire u2__abc_52155_new_n4938_; 
wire u2__abc_52155_new_n4939_; 
wire u2__abc_52155_new_n4940_; 
wire u2__abc_52155_new_n4941_; 
wire u2__abc_52155_new_n4942_; 
wire u2__abc_52155_new_n4943_; 
wire u2__abc_52155_new_n4944_; 
wire u2__abc_52155_new_n4945_; 
wire u2__abc_52155_new_n4946_; 
wire u2__abc_52155_new_n4947_; 
wire u2__abc_52155_new_n4948_; 
wire u2__abc_52155_new_n4949_; 
wire u2__abc_52155_new_n4950_; 
wire u2__abc_52155_new_n4951_; 
wire u2__abc_52155_new_n4952_; 
wire u2__abc_52155_new_n4953_; 
wire u2__abc_52155_new_n4954_; 
wire u2__abc_52155_new_n4955_; 
wire u2__abc_52155_new_n4956_; 
wire u2__abc_52155_new_n4957_; 
wire u2__abc_52155_new_n4958_; 
wire u2__abc_52155_new_n4959_; 
wire u2__abc_52155_new_n4960_; 
wire u2__abc_52155_new_n4961_; 
wire u2__abc_52155_new_n4962_; 
wire u2__abc_52155_new_n4963_; 
wire u2__abc_52155_new_n4964_; 
wire u2__abc_52155_new_n4965_; 
wire u2__abc_52155_new_n4966_; 
wire u2__abc_52155_new_n4967_; 
wire u2__abc_52155_new_n4968_; 
wire u2__abc_52155_new_n4969_; 
wire u2__abc_52155_new_n4970_; 
wire u2__abc_52155_new_n4971_; 
wire u2__abc_52155_new_n4972_; 
wire u2__abc_52155_new_n4973_; 
wire u2__abc_52155_new_n4974_; 
wire u2__abc_52155_new_n4975_; 
wire u2__abc_52155_new_n4976_; 
wire u2__abc_52155_new_n4977_; 
wire u2__abc_52155_new_n4978_; 
wire u2__abc_52155_new_n4979_; 
wire u2__abc_52155_new_n4980_; 
wire u2__abc_52155_new_n4981_; 
wire u2__abc_52155_new_n4982_; 
wire u2__abc_52155_new_n4983_; 
wire u2__abc_52155_new_n4984_; 
wire u2__abc_52155_new_n4985_; 
wire u2__abc_52155_new_n4986_; 
wire u2__abc_52155_new_n4987_; 
wire u2__abc_52155_new_n4988_; 
wire u2__abc_52155_new_n4989_; 
wire u2__abc_52155_new_n4990_; 
wire u2__abc_52155_new_n4991_; 
wire u2__abc_52155_new_n4992_; 
wire u2__abc_52155_new_n4993_; 
wire u2__abc_52155_new_n4994_; 
wire u2__abc_52155_new_n4995_; 
wire u2__abc_52155_new_n4996_; 
wire u2__abc_52155_new_n4997_; 
wire u2__abc_52155_new_n4998_; 
wire u2__abc_52155_new_n4999_; 
wire u2__abc_52155_new_n5000_; 
wire u2__abc_52155_new_n5001_; 
wire u2__abc_52155_new_n5002_; 
wire u2__abc_52155_new_n5003_; 
wire u2__abc_52155_new_n5004_; 
wire u2__abc_52155_new_n5005_; 
wire u2__abc_52155_new_n5006_; 
wire u2__abc_52155_new_n5007_; 
wire u2__abc_52155_new_n5008_; 
wire u2__abc_52155_new_n5009_; 
wire u2__abc_52155_new_n5010_; 
wire u2__abc_52155_new_n5011_; 
wire u2__abc_52155_new_n5012_; 
wire u2__abc_52155_new_n5013_; 
wire u2__abc_52155_new_n5014_; 
wire u2__abc_52155_new_n5015_; 
wire u2__abc_52155_new_n5016_; 
wire u2__abc_52155_new_n5017_; 
wire u2__abc_52155_new_n5018_; 
wire u2__abc_52155_new_n5019_; 
wire u2__abc_52155_new_n5020_; 
wire u2__abc_52155_new_n5021_; 
wire u2__abc_52155_new_n5022_; 
wire u2__abc_52155_new_n5023_; 
wire u2__abc_52155_new_n5024_; 
wire u2__abc_52155_new_n5025_; 
wire u2__abc_52155_new_n5026_; 
wire u2__abc_52155_new_n5027_; 
wire u2__abc_52155_new_n5028_; 
wire u2__abc_52155_new_n5029_; 
wire u2__abc_52155_new_n5030_; 
wire u2__abc_52155_new_n5031_; 
wire u2__abc_52155_new_n5032_; 
wire u2__abc_52155_new_n5033_; 
wire u2__abc_52155_new_n5034_; 
wire u2__abc_52155_new_n5035_; 
wire u2__abc_52155_new_n5036_; 
wire u2__abc_52155_new_n5037_; 
wire u2__abc_52155_new_n5038_; 
wire u2__abc_52155_new_n5039_; 
wire u2__abc_52155_new_n5040_; 
wire u2__abc_52155_new_n5041_; 
wire u2__abc_52155_new_n5042_; 
wire u2__abc_52155_new_n5043_; 
wire u2__abc_52155_new_n5044_; 
wire u2__abc_52155_new_n5045_; 
wire u2__abc_52155_new_n5046_; 
wire u2__abc_52155_new_n5047_; 
wire u2__abc_52155_new_n5048_; 
wire u2__abc_52155_new_n5049_; 
wire u2__abc_52155_new_n5050_; 
wire u2__abc_52155_new_n5051_; 
wire u2__abc_52155_new_n5052_; 
wire u2__abc_52155_new_n5053_; 
wire u2__abc_52155_new_n5054_; 
wire u2__abc_52155_new_n5055_; 
wire u2__abc_52155_new_n5056_; 
wire u2__abc_52155_new_n5057_; 
wire u2__abc_52155_new_n5058_; 
wire u2__abc_52155_new_n5059_; 
wire u2__abc_52155_new_n5060_; 
wire u2__abc_52155_new_n5061_; 
wire u2__abc_52155_new_n5062_; 
wire u2__abc_52155_new_n5063_; 
wire u2__abc_52155_new_n5064_; 
wire u2__abc_52155_new_n5065_; 
wire u2__abc_52155_new_n5066_; 
wire u2__abc_52155_new_n5067_; 
wire u2__abc_52155_new_n5068_; 
wire u2__abc_52155_new_n5069_; 
wire u2__abc_52155_new_n5070_; 
wire u2__abc_52155_new_n5071_; 
wire u2__abc_52155_new_n5072_; 
wire u2__abc_52155_new_n5073_; 
wire u2__abc_52155_new_n5074_; 
wire u2__abc_52155_new_n5075_; 
wire u2__abc_52155_new_n5076_; 
wire u2__abc_52155_new_n5077_; 
wire u2__abc_52155_new_n5078_; 
wire u2__abc_52155_new_n5079_; 
wire u2__abc_52155_new_n5080_; 
wire u2__abc_52155_new_n5081_; 
wire u2__abc_52155_new_n5082_; 
wire u2__abc_52155_new_n5083_; 
wire u2__abc_52155_new_n5084_; 
wire u2__abc_52155_new_n5085_; 
wire u2__abc_52155_new_n5086_; 
wire u2__abc_52155_new_n5087_; 
wire u2__abc_52155_new_n5088_; 
wire u2__abc_52155_new_n5089_; 
wire u2__abc_52155_new_n5090_; 
wire u2__abc_52155_new_n5091_; 
wire u2__abc_52155_new_n5092_; 
wire u2__abc_52155_new_n5093_; 
wire u2__abc_52155_new_n5094_; 
wire u2__abc_52155_new_n5095_; 
wire u2__abc_52155_new_n5096_; 
wire u2__abc_52155_new_n5097_; 
wire u2__abc_52155_new_n5098_; 
wire u2__abc_52155_new_n5099_; 
wire u2__abc_52155_new_n5100_; 
wire u2__abc_52155_new_n5101_; 
wire u2__abc_52155_new_n5102_; 
wire u2__abc_52155_new_n5103_; 
wire u2__abc_52155_new_n5104_; 
wire u2__abc_52155_new_n5105_; 
wire u2__abc_52155_new_n5106_; 
wire u2__abc_52155_new_n5107_; 
wire u2__abc_52155_new_n5108_; 
wire u2__abc_52155_new_n5109_; 
wire u2__abc_52155_new_n5110_; 
wire u2__abc_52155_new_n5111_; 
wire u2__abc_52155_new_n5112_; 
wire u2__abc_52155_new_n5113_; 
wire u2__abc_52155_new_n5114_; 
wire u2__abc_52155_new_n5115_; 
wire u2__abc_52155_new_n5116_; 
wire u2__abc_52155_new_n5117_; 
wire u2__abc_52155_new_n5118_; 
wire u2__abc_52155_new_n5119_; 
wire u2__abc_52155_new_n5120_; 
wire u2__abc_52155_new_n5121_; 
wire u2__abc_52155_new_n5122_; 
wire u2__abc_52155_new_n5123_; 
wire u2__abc_52155_new_n5124_; 
wire u2__abc_52155_new_n5125_; 
wire u2__abc_52155_new_n5126_; 
wire u2__abc_52155_new_n5127_; 
wire u2__abc_52155_new_n5128_; 
wire u2__abc_52155_new_n5129_; 
wire u2__abc_52155_new_n5130_; 
wire u2__abc_52155_new_n5131_; 
wire u2__abc_52155_new_n5132_; 
wire u2__abc_52155_new_n5133_; 
wire u2__abc_52155_new_n5134_; 
wire u2__abc_52155_new_n5135_; 
wire u2__abc_52155_new_n5136_; 
wire u2__abc_52155_new_n5137_; 
wire u2__abc_52155_new_n5138_; 
wire u2__abc_52155_new_n5139_; 
wire u2__abc_52155_new_n5140_; 
wire u2__abc_52155_new_n5141_; 
wire u2__abc_52155_new_n5142_; 
wire u2__abc_52155_new_n5143_; 
wire u2__abc_52155_new_n5144_; 
wire u2__abc_52155_new_n5145_; 
wire u2__abc_52155_new_n5146_; 
wire u2__abc_52155_new_n5147_; 
wire u2__abc_52155_new_n5148_; 
wire u2__abc_52155_new_n5149_; 
wire u2__abc_52155_new_n5150_; 
wire u2__abc_52155_new_n5151_; 
wire u2__abc_52155_new_n5152_; 
wire u2__abc_52155_new_n5153_; 
wire u2__abc_52155_new_n5154_; 
wire u2__abc_52155_new_n5155_; 
wire u2__abc_52155_new_n5156_; 
wire u2__abc_52155_new_n5157_; 
wire u2__abc_52155_new_n5158_; 
wire u2__abc_52155_new_n5159_; 
wire u2__abc_52155_new_n5160_; 
wire u2__abc_52155_new_n5161_; 
wire u2__abc_52155_new_n5162_; 
wire u2__abc_52155_new_n5163_; 
wire u2__abc_52155_new_n5164_; 
wire u2__abc_52155_new_n5165_; 
wire u2__abc_52155_new_n5166_; 
wire u2__abc_52155_new_n5167_; 
wire u2__abc_52155_new_n5168_; 
wire u2__abc_52155_new_n5169_; 
wire u2__abc_52155_new_n5170_; 
wire u2__abc_52155_new_n5171_; 
wire u2__abc_52155_new_n5172_; 
wire u2__abc_52155_new_n5173_; 
wire u2__abc_52155_new_n5174_; 
wire u2__abc_52155_new_n5175_; 
wire u2__abc_52155_new_n5176_; 
wire u2__abc_52155_new_n5177_; 
wire u2__abc_52155_new_n5178_; 
wire u2__abc_52155_new_n5179_; 
wire u2__abc_52155_new_n5180_; 
wire u2__abc_52155_new_n5181_; 
wire u2__abc_52155_new_n5182_; 
wire u2__abc_52155_new_n5183_; 
wire u2__abc_52155_new_n5184_; 
wire u2__abc_52155_new_n5185_; 
wire u2__abc_52155_new_n5186_; 
wire u2__abc_52155_new_n5187_; 
wire u2__abc_52155_new_n5188_; 
wire u2__abc_52155_new_n5189_; 
wire u2__abc_52155_new_n5190_; 
wire u2__abc_52155_new_n5191_; 
wire u2__abc_52155_new_n5192_; 
wire u2__abc_52155_new_n5193_; 
wire u2__abc_52155_new_n5194_; 
wire u2__abc_52155_new_n5195_; 
wire u2__abc_52155_new_n5196_; 
wire u2__abc_52155_new_n5197_; 
wire u2__abc_52155_new_n5198_; 
wire u2__abc_52155_new_n5199_; 
wire u2__abc_52155_new_n5200_; 
wire u2__abc_52155_new_n5201_; 
wire u2__abc_52155_new_n5202_; 
wire u2__abc_52155_new_n5203_; 
wire u2__abc_52155_new_n5204_; 
wire u2__abc_52155_new_n5205_; 
wire u2__abc_52155_new_n5206_; 
wire u2__abc_52155_new_n5207_; 
wire u2__abc_52155_new_n5208_; 
wire u2__abc_52155_new_n5209_; 
wire u2__abc_52155_new_n5210_; 
wire u2__abc_52155_new_n5211_; 
wire u2__abc_52155_new_n5212_; 
wire u2__abc_52155_new_n5213_; 
wire u2__abc_52155_new_n5214_; 
wire u2__abc_52155_new_n5215_; 
wire u2__abc_52155_new_n5216_; 
wire u2__abc_52155_new_n5217_; 
wire u2__abc_52155_new_n5218_; 
wire u2__abc_52155_new_n5219_; 
wire u2__abc_52155_new_n5220_; 
wire u2__abc_52155_new_n5221_; 
wire u2__abc_52155_new_n5222_; 
wire u2__abc_52155_new_n5223_; 
wire u2__abc_52155_new_n5224_; 
wire u2__abc_52155_new_n5225_; 
wire u2__abc_52155_new_n5226_; 
wire u2__abc_52155_new_n5227_; 
wire u2__abc_52155_new_n5228_; 
wire u2__abc_52155_new_n5229_; 
wire u2__abc_52155_new_n5230_; 
wire u2__abc_52155_new_n5231_; 
wire u2__abc_52155_new_n5232_; 
wire u2__abc_52155_new_n5233_; 
wire u2__abc_52155_new_n5234_; 
wire u2__abc_52155_new_n5235_; 
wire u2__abc_52155_new_n5236_; 
wire u2__abc_52155_new_n5237_; 
wire u2__abc_52155_new_n5238_; 
wire u2__abc_52155_new_n5239_; 
wire u2__abc_52155_new_n5240_; 
wire u2__abc_52155_new_n5241_; 
wire u2__abc_52155_new_n5242_; 
wire u2__abc_52155_new_n5243_; 
wire u2__abc_52155_new_n5244_; 
wire u2__abc_52155_new_n5245_; 
wire u2__abc_52155_new_n5246_; 
wire u2__abc_52155_new_n5247_; 
wire u2__abc_52155_new_n5248_; 
wire u2__abc_52155_new_n5249_; 
wire u2__abc_52155_new_n5250_; 
wire u2__abc_52155_new_n5251_; 
wire u2__abc_52155_new_n5252_; 
wire u2__abc_52155_new_n5253_; 
wire u2__abc_52155_new_n5254_; 
wire u2__abc_52155_new_n5255_; 
wire u2__abc_52155_new_n5256_; 
wire u2__abc_52155_new_n5257_; 
wire u2__abc_52155_new_n5258_; 
wire u2__abc_52155_new_n5259_; 
wire u2__abc_52155_new_n5260_; 
wire u2__abc_52155_new_n5261_; 
wire u2__abc_52155_new_n5262_; 
wire u2__abc_52155_new_n5263_; 
wire u2__abc_52155_new_n5264_; 
wire u2__abc_52155_new_n5265_; 
wire u2__abc_52155_new_n5266_; 
wire u2__abc_52155_new_n5267_; 
wire u2__abc_52155_new_n5268_; 
wire u2__abc_52155_new_n5269_; 
wire u2__abc_52155_new_n5270_; 
wire u2__abc_52155_new_n5271_; 
wire u2__abc_52155_new_n5272_; 
wire u2__abc_52155_new_n5273_; 
wire u2__abc_52155_new_n5274_; 
wire u2__abc_52155_new_n5275_; 
wire u2__abc_52155_new_n5276_; 
wire u2__abc_52155_new_n5277_; 
wire u2__abc_52155_new_n5278_; 
wire u2__abc_52155_new_n5279_; 
wire u2__abc_52155_new_n5280_; 
wire u2__abc_52155_new_n5281_; 
wire u2__abc_52155_new_n5282_; 
wire u2__abc_52155_new_n5283_; 
wire u2__abc_52155_new_n5284_; 
wire u2__abc_52155_new_n5285_; 
wire u2__abc_52155_new_n5286_; 
wire u2__abc_52155_new_n5287_; 
wire u2__abc_52155_new_n5288_; 
wire u2__abc_52155_new_n5289_; 
wire u2__abc_52155_new_n5290_; 
wire u2__abc_52155_new_n5291_; 
wire u2__abc_52155_new_n5292_; 
wire u2__abc_52155_new_n5293_; 
wire u2__abc_52155_new_n5294_; 
wire u2__abc_52155_new_n5295_; 
wire u2__abc_52155_new_n5296_; 
wire u2__abc_52155_new_n5297_; 
wire u2__abc_52155_new_n5298_; 
wire u2__abc_52155_new_n5299_; 
wire u2__abc_52155_new_n5300_; 
wire u2__abc_52155_new_n5301_; 
wire u2__abc_52155_new_n5302_; 
wire u2__abc_52155_new_n5303_; 
wire u2__abc_52155_new_n5304_; 
wire u2__abc_52155_new_n5305_; 
wire u2__abc_52155_new_n5306_; 
wire u2__abc_52155_new_n5307_; 
wire u2__abc_52155_new_n5308_; 
wire u2__abc_52155_new_n5309_; 
wire u2__abc_52155_new_n5310_; 
wire u2__abc_52155_new_n5311_; 
wire u2__abc_52155_new_n5312_; 
wire u2__abc_52155_new_n5313_; 
wire u2__abc_52155_new_n5314_; 
wire u2__abc_52155_new_n5315_; 
wire u2__abc_52155_new_n5316_; 
wire u2__abc_52155_new_n5317_; 
wire u2__abc_52155_new_n5318_; 
wire u2__abc_52155_new_n5319_; 
wire u2__abc_52155_new_n5320_; 
wire u2__abc_52155_new_n5321_; 
wire u2__abc_52155_new_n5322_; 
wire u2__abc_52155_new_n5323_; 
wire u2__abc_52155_new_n5324_; 
wire u2__abc_52155_new_n5325_; 
wire u2__abc_52155_new_n5326_; 
wire u2__abc_52155_new_n5327_; 
wire u2__abc_52155_new_n5328_; 
wire u2__abc_52155_new_n5329_; 
wire u2__abc_52155_new_n5330_; 
wire u2__abc_52155_new_n5331_; 
wire u2__abc_52155_new_n5332_; 
wire u2__abc_52155_new_n5333_; 
wire u2__abc_52155_new_n5334_; 
wire u2__abc_52155_new_n5335_; 
wire u2__abc_52155_new_n5336_; 
wire u2__abc_52155_new_n5337_; 
wire u2__abc_52155_new_n5338_; 
wire u2__abc_52155_new_n5339_; 
wire u2__abc_52155_new_n5340_; 
wire u2__abc_52155_new_n5341_; 
wire u2__abc_52155_new_n5342_; 
wire u2__abc_52155_new_n5343_; 
wire u2__abc_52155_new_n5344_; 
wire u2__abc_52155_new_n5345_; 
wire u2__abc_52155_new_n5346_; 
wire u2__abc_52155_new_n5347_; 
wire u2__abc_52155_new_n5348_; 
wire u2__abc_52155_new_n5349_; 
wire u2__abc_52155_new_n5350_; 
wire u2__abc_52155_new_n5351_; 
wire u2__abc_52155_new_n5352_; 
wire u2__abc_52155_new_n5353_; 
wire u2__abc_52155_new_n5354_; 
wire u2__abc_52155_new_n5355_; 
wire u2__abc_52155_new_n5356_; 
wire u2__abc_52155_new_n5357_; 
wire u2__abc_52155_new_n5358_; 
wire u2__abc_52155_new_n5359_; 
wire u2__abc_52155_new_n5360_; 
wire u2__abc_52155_new_n5361_; 
wire u2__abc_52155_new_n5362_; 
wire u2__abc_52155_new_n5363_; 
wire u2__abc_52155_new_n5364_; 
wire u2__abc_52155_new_n5365_; 
wire u2__abc_52155_new_n5366_; 
wire u2__abc_52155_new_n5367_; 
wire u2__abc_52155_new_n5368_; 
wire u2__abc_52155_new_n5369_; 
wire u2__abc_52155_new_n5370_; 
wire u2__abc_52155_new_n5371_; 
wire u2__abc_52155_new_n5372_; 
wire u2__abc_52155_new_n5373_; 
wire u2__abc_52155_new_n5374_; 
wire u2__abc_52155_new_n5375_; 
wire u2__abc_52155_new_n5376_; 
wire u2__abc_52155_new_n5377_; 
wire u2__abc_52155_new_n5378_; 
wire u2__abc_52155_new_n5379_; 
wire u2__abc_52155_new_n5380_; 
wire u2__abc_52155_new_n5381_; 
wire u2__abc_52155_new_n5382_; 
wire u2__abc_52155_new_n5383_; 
wire u2__abc_52155_new_n5384_; 
wire u2__abc_52155_new_n5385_; 
wire u2__abc_52155_new_n5386_; 
wire u2__abc_52155_new_n5387_; 
wire u2__abc_52155_new_n5388_; 
wire u2__abc_52155_new_n5389_; 
wire u2__abc_52155_new_n5390_; 
wire u2__abc_52155_new_n5391_; 
wire u2__abc_52155_new_n5392_; 
wire u2__abc_52155_new_n5393_; 
wire u2__abc_52155_new_n5394_; 
wire u2__abc_52155_new_n5395_; 
wire u2__abc_52155_new_n5396_; 
wire u2__abc_52155_new_n5397_; 
wire u2__abc_52155_new_n5398_; 
wire u2__abc_52155_new_n5399_; 
wire u2__abc_52155_new_n5400_; 
wire u2__abc_52155_new_n5401_; 
wire u2__abc_52155_new_n5402_; 
wire u2__abc_52155_new_n5403_; 
wire u2__abc_52155_new_n5404_; 
wire u2__abc_52155_new_n5405_; 
wire u2__abc_52155_new_n5406_; 
wire u2__abc_52155_new_n5407_; 
wire u2__abc_52155_new_n5408_; 
wire u2__abc_52155_new_n5409_; 
wire u2__abc_52155_new_n5410_; 
wire u2__abc_52155_new_n5411_; 
wire u2__abc_52155_new_n5412_; 
wire u2__abc_52155_new_n5413_; 
wire u2__abc_52155_new_n5414_; 
wire u2__abc_52155_new_n5415_; 
wire u2__abc_52155_new_n5416_; 
wire u2__abc_52155_new_n5417_; 
wire u2__abc_52155_new_n5418_; 
wire u2__abc_52155_new_n5419_; 
wire u2__abc_52155_new_n5420_; 
wire u2__abc_52155_new_n5421_; 
wire u2__abc_52155_new_n5422_; 
wire u2__abc_52155_new_n5423_; 
wire u2__abc_52155_new_n5424_; 
wire u2__abc_52155_new_n5425_; 
wire u2__abc_52155_new_n5426_; 
wire u2__abc_52155_new_n5427_; 
wire u2__abc_52155_new_n5428_; 
wire u2__abc_52155_new_n5429_; 
wire u2__abc_52155_new_n5430_; 
wire u2__abc_52155_new_n5431_; 
wire u2__abc_52155_new_n5432_; 
wire u2__abc_52155_new_n5433_; 
wire u2__abc_52155_new_n5434_; 
wire u2__abc_52155_new_n5435_; 
wire u2__abc_52155_new_n5436_; 
wire u2__abc_52155_new_n5437_; 
wire u2__abc_52155_new_n5438_; 
wire u2__abc_52155_new_n5439_; 
wire u2__abc_52155_new_n5440_; 
wire u2__abc_52155_new_n5441_; 
wire u2__abc_52155_new_n5442_; 
wire u2__abc_52155_new_n5443_; 
wire u2__abc_52155_new_n5444_; 
wire u2__abc_52155_new_n5445_; 
wire u2__abc_52155_new_n5446_; 
wire u2__abc_52155_new_n5447_; 
wire u2__abc_52155_new_n5448_; 
wire u2__abc_52155_new_n5449_; 
wire u2__abc_52155_new_n5450_; 
wire u2__abc_52155_new_n5451_; 
wire u2__abc_52155_new_n5452_; 
wire u2__abc_52155_new_n5453_; 
wire u2__abc_52155_new_n5454_; 
wire u2__abc_52155_new_n5455_; 
wire u2__abc_52155_new_n5456_; 
wire u2__abc_52155_new_n5457_; 
wire u2__abc_52155_new_n5458_; 
wire u2__abc_52155_new_n5459_; 
wire u2__abc_52155_new_n5460_; 
wire u2__abc_52155_new_n5461_; 
wire u2__abc_52155_new_n5462_; 
wire u2__abc_52155_new_n5463_; 
wire u2__abc_52155_new_n5464_; 
wire u2__abc_52155_new_n5465_; 
wire u2__abc_52155_new_n5466_; 
wire u2__abc_52155_new_n5467_; 
wire u2__abc_52155_new_n5468_; 
wire u2__abc_52155_new_n5469_; 
wire u2__abc_52155_new_n5470_; 
wire u2__abc_52155_new_n5471_; 
wire u2__abc_52155_new_n5472_; 
wire u2__abc_52155_new_n5473_; 
wire u2__abc_52155_new_n5474_; 
wire u2__abc_52155_new_n5475_; 
wire u2__abc_52155_new_n5476_; 
wire u2__abc_52155_new_n5477_; 
wire u2__abc_52155_new_n5478_; 
wire u2__abc_52155_new_n5479_; 
wire u2__abc_52155_new_n5480_; 
wire u2__abc_52155_new_n5481_; 
wire u2__abc_52155_new_n5482_; 
wire u2__abc_52155_new_n5483_; 
wire u2__abc_52155_new_n5484_; 
wire u2__abc_52155_new_n5485_; 
wire u2__abc_52155_new_n5486_; 
wire u2__abc_52155_new_n5487_; 
wire u2__abc_52155_new_n5488_; 
wire u2__abc_52155_new_n5489_; 
wire u2__abc_52155_new_n5490_; 
wire u2__abc_52155_new_n5491_; 
wire u2__abc_52155_new_n5492_; 
wire u2__abc_52155_new_n5493_; 
wire u2__abc_52155_new_n5494_; 
wire u2__abc_52155_new_n5495_; 
wire u2__abc_52155_new_n5496_; 
wire u2__abc_52155_new_n5497_; 
wire u2__abc_52155_new_n5498_; 
wire u2__abc_52155_new_n5499_; 
wire u2__abc_52155_new_n5500_; 
wire u2__abc_52155_new_n5501_; 
wire u2__abc_52155_new_n5502_; 
wire u2__abc_52155_new_n5503_; 
wire u2__abc_52155_new_n5504_; 
wire u2__abc_52155_new_n5505_; 
wire u2__abc_52155_new_n5506_; 
wire u2__abc_52155_new_n5507_; 
wire u2__abc_52155_new_n5508_; 
wire u2__abc_52155_new_n5509_; 
wire u2__abc_52155_new_n5510_; 
wire u2__abc_52155_new_n5511_; 
wire u2__abc_52155_new_n5512_; 
wire u2__abc_52155_new_n5513_; 
wire u2__abc_52155_new_n5514_; 
wire u2__abc_52155_new_n5515_; 
wire u2__abc_52155_new_n5516_; 
wire u2__abc_52155_new_n5517_; 
wire u2__abc_52155_new_n5518_; 
wire u2__abc_52155_new_n5519_; 
wire u2__abc_52155_new_n5520_; 
wire u2__abc_52155_new_n5521_; 
wire u2__abc_52155_new_n5522_; 
wire u2__abc_52155_new_n5523_; 
wire u2__abc_52155_new_n5524_; 
wire u2__abc_52155_new_n5525_; 
wire u2__abc_52155_new_n5526_; 
wire u2__abc_52155_new_n5527_; 
wire u2__abc_52155_new_n5528_; 
wire u2__abc_52155_new_n5529_; 
wire u2__abc_52155_new_n5530_; 
wire u2__abc_52155_new_n5531_; 
wire u2__abc_52155_new_n5532_; 
wire u2__abc_52155_new_n5533_; 
wire u2__abc_52155_new_n5534_; 
wire u2__abc_52155_new_n5535_; 
wire u2__abc_52155_new_n5536_; 
wire u2__abc_52155_new_n5537_; 
wire u2__abc_52155_new_n5538_; 
wire u2__abc_52155_new_n5539_; 
wire u2__abc_52155_new_n5540_; 
wire u2__abc_52155_new_n5541_; 
wire u2__abc_52155_new_n5542_; 
wire u2__abc_52155_new_n5543_; 
wire u2__abc_52155_new_n5544_; 
wire u2__abc_52155_new_n5545_; 
wire u2__abc_52155_new_n5546_; 
wire u2__abc_52155_new_n5547_; 
wire u2__abc_52155_new_n5548_; 
wire u2__abc_52155_new_n5549_; 
wire u2__abc_52155_new_n5550_; 
wire u2__abc_52155_new_n5551_; 
wire u2__abc_52155_new_n5552_; 
wire u2__abc_52155_new_n5553_; 
wire u2__abc_52155_new_n5554_; 
wire u2__abc_52155_new_n5555_; 
wire u2__abc_52155_new_n5556_; 
wire u2__abc_52155_new_n5557_; 
wire u2__abc_52155_new_n5558_; 
wire u2__abc_52155_new_n5559_; 
wire u2__abc_52155_new_n5560_; 
wire u2__abc_52155_new_n5561_; 
wire u2__abc_52155_new_n5562_; 
wire u2__abc_52155_new_n5563_; 
wire u2__abc_52155_new_n5564_; 
wire u2__abc_52155_new_n5565_; 
wire u2__abc_52155_new_n5566_; 
wire u2__abc_52155_new_n5567_; 
wire u2__abc_52155_new_n5568_; 
wire u2__abc_52155_new_n5569_; 
wire u2__abc_52155_new_n5570_; 
wire u2__abc_52155_new_n5571_; 
wire u2__abc_52155_new_n5572_; 
wire u2__abc_52155_new_n5573_; 
wire u2__abc_52155_new_n5574_; 
wire u2__abc_52155_new_n5575_; 
wire u2__abc_52155_new_n5576_; 
wire u2__abc_52155_new_n5577_; 
wire u2__abc_52155_new_n5578_; 
wire u2__abc_52155_new_n5579_; 
wire u2__abc_52155_new_n5580_; 
wire u2__abc_52155_new_n5581_; 
wire u2__abc_52155_new_n5582_; 
wire u2__abc_52155_new_n5583_; 
wire u2__abc_52155_new_n5584_; 
wire u2__abc_52155_new_n5585_; 
wire u2__abc_52155_new_n5586_; 
wire u2__abc_52155_new_n5587_; 
wire u2__abc_52155_new_n5588_; 
wire u2__abc_52155_new_n5589_; 
wire u2__abc_52155_new_n5590_; 
wire u2__abc_52155_new_n5591_; 
wire u2__abc_52155_new_n5592_; 
wire u2__abc_52155_new_n5593_; 
wire u2__abc_52155_new_n5594_; 
wire u2__abc_52155_new_n5595_; 
wire u2__abc_52155_new_n5596_; 
wire u2__abc_52155_new_n5597_; 
wire u2__abc_52155_new_n5598_; 
wire u2__abc_52155_new_n5599_; 
wire u2__abc_52155_new_n5600_; 
wire u2__abc_52155_new_n5601_; 
wire u2__abc_52155_new_n5602_; 
wire u2__abc_52155_new_n5603_; 
wire u2__abc_52155_new_n5604_; 
wire u2__abc_52155_new_n5605_; 
wire u2__abc_52155_new_n5606_; 
wire u2__abc_52155_new_n5607_; 
wire u2__abc_52155_new_n5608_; 
wire u2__abc_52155_new_n5609_; 
wire u2__abc_52155_new_n5610_; 
wire u2__abc_52155_new_n5611_; 
wire u2__abc_52155_new_n5612_; 
wire u2__abc_52155_new_n5613_; 
wire u2__abc_52155_new_n5614_; 
wire u2__abc_52155_new_n5615_; 
wire u2__abc_52155_new_n5616_; 
wire u2__abc_52155_new_n5617_; 
wire u2__abc_52155_new_n5618_; 
wire u2__abc_52155_new_n5619_; 
wire u2__abc_52155_new_n5620_; 
wire u2__abc_52155_new_n5621_; 
wire u2__abc_52155_new_n5622_; 
wire u2__abc_52155_new_n5623_; 
wire u2__abc_52155_new_n5624_; 
wire u2__abc_52155_new_n5625_; 
wire u2__abc_52155_new_n5626_; 
wire u2__abc_52155_new_n5627_; 
wire u2__abc_52155_new_n5628_; 
wire u2__abc_52155_new_n5629_; 
wire u2__abc_52155_new_n5630_; 
wire u2__abc_52155_new_n5631_; 
wire u2__abc_52155_new_n5632_; 
wire u2__abc_52155_new_n5633_; 
wire u2__abc_52155_new_n5634_; 
wire u2__abc_52155_new_n5635_; 
wire u2__abc_52155_new_n5636_; 
wire u2__abc_52155_new_n5637_; 
wire u2__abc_52155_new_n5638_; 
wire u2__abc_52155_new_n5639_; 
wire u2__abc_52155_new_n5640_; 
wire u2__abc_52155_new_n5641_; 
wire u2__abc_52155_new_n5642_; 
wire u2__abc_52155_new_n5643_; 
wire u2__abc_52155_new_n5644_; 
wire u2__abc_52155_new_n5645_; 
wire u2__abc_52155_new_n5646_; 
wire u2__abc_52155_new_n5647_; 
wire u2__abc_52155_new_n5648_; 
wire u2__abc_52155_new_n5649_; 
wire u2__abc_52155_new_n5650_; 
wire u2__abc_52155_new_n5651_; 
wire u2__abc_52155_new_n5652_; 
wire u2__abc_52155_new_n5653_; 
wire u2__abc_52155_new_n5654_; 
wire u2__abc_52155_new_n5655_; 
wire u2__abc_52155_new_n5656_; 
wire u2__abc_52155_new_n5657_; 
wire u2__abc_52155_new_n5658_; 
wire u2__abc_52155_new_n5659_; 
wire u2__abc_52155_new_n5660_; 
wire u2__abc_52155_new_n5661_; 
wire u2__abc_52155_new_n5662_; 
wire u2__abc_52155_new_n5663_; 
wire u2__abc_52155_new_n5664_; 
wire u2__abc_52155_new_n5665_; 
wire u2__abc_52155_new_n5666_; 
wire u2__abc_52155_new_n5667_; 
wire u2__abc_52155_new_n5668_; 
wire u2__abc_52155_new_n5669_; 
wire u2__abc_52155_new_n5670_; 
wire u2__abc_52155_new_n5671_; 
wire u2__abc_52155_new_n5672_; 
wire u2__abc_52155_new_n5673_; 
wire u2__abc_52155_new_n5674_; 
wire u2__abc_52155_new_n5675_; 
wire u2__abc_52155_new_n5676_; 
wire u2__abc_52155_new_n5677_; 
wire u2__abc_52155_new_n5678_; 
wire u2__abc_52155_new_n5679_; 
wire u2__abc_52155_new_n5680_; 
wire u2__abc_52155_new_n5681_; 
wire u2__abc_52155_new_n5682_; 
wire u2__abc_52155_new_n5683_; 
wire u2__abc_52155_new_n5684_; 
wire u2__abc_52155_new_n5685_; 
wire u2__abc_52155_new_n5686_; 
wire u2__abc_52155_new_n5687_; 
wire u2__abc_52155_new_n5688_; 
wire u2__abc_52155_new_n5689_; 
wire u2__abc_52155_new_n5690_; 
wire u2__abc_52155_new_n5691_; 
wire u2__abc_52155_new_n5692_; 
wire u2__abc_52155_new_n5693_; 
wire u2__abc_52155_new_n5694_; 
wire u2__abc_52155_new_n5695_; 
wire u2__abc_52155_new_n5696_; 
wire u2__abc_52155_new_n5697_; 
wire u2__abc_52155_new_n5698_; 
wire u2__abc_52155_new_n5699_; 
wire u2__abc_52155_new_n5700_; 
wire u2__abc_52155_new_n5701_; 
wire u2__abc_52155_new_n5702_; 
wire u2__abc_52155_new_n5703_; 
wire u2__abc_52155_new_n5704_; 
wire u2__abc_52155_new_n5705_; 
wire u2__abc_52155_new_n5706_; 
wire u2__abc_52155_new_n5707_; 
wire u2__abc_52155_new_n5708_; 
wire u2__abc_52155_new_n5709_; 
wire u2__abc_52155_new_n5710_; 
wire u2__abc_52155_new_n5711_; 
wire u2__abc_52155_new_n5712_; 
wire u2__abc_52155_new_n5713_; 
wire u2__abc_52155_new_n5714_; 
wire u2__abc_52155_new_n5715_; 
wire u2__abc_52155_new_n5716_; 
wire u2__abc_52155_new_n5717_; 
wire u2__abc_52155_new_n5718_; 
wire u2__abc_52155_new_n5719_; 
wire u2__abc_52155_new_n5720_; 
wire u2__abc_52155_new_n5721_; 
wire u2__abc_52155_new_n5722_; 
wire u2__abc_52155_new_n5723_; 
wire u2__abc_52155_new_n5724_; 
wire u2__abc_52155_new_n5725_; 
wire u2__abc_52155_new_n5726_; 
wire u2__abc_52155_new_n5727_; 
wire u2__abc_52155_new_n5728_; 
wire u2__abc_52155_new_n5729_; 
wire u2__abc_52155_new_n5730_; 
wire u2__abc_52155_new_n5731_; 
wire u2__abc_52155_new_n5732_; 
wire u2__abc_52155_new_n5733_; 
wire u2__abc_52155_new_n5734_; 
wire u2__abc_52155_new_n5735_; 
wire u2__abc_52155_new_n5736_; 
wire u2__abc_52155_new_n5737_; 
wire u2__abc_52155_new_n5738_; 
wire u2__abc_52155_new_n5739_; 
wire u2__abc_52155_new_n5740_; 
wire u2__abc_52155_new_n5741_; 
wire u2__abc_52155_new_n5742_; 
wire u2__abc_52155_new_n5743_; 
wire u2__abc_52155_new_n5744_; 
wire u2__abc_52155_new_n5745_; 
wire u2__abc_52155_new_n5746_; 
wire u2__abc_52155_new_n5747_; 
wire u2__abc_52155_new_n5748_; 
wire u2__abc_52155_new_n5749_; 
wire u2__abc_52155_new_n5750_; 
wire u2__abc_52155_new_n5751_; 
wire u2__abc_52155_new_n5752_; 
wire u2__abc_52155_new_n5753_; 
wire u2__abc_52155_new_n5754_; 
wire u2__abc_52155_new_n5755_; 
wire u2__abc_52155_new_n5756_; 
wire u2__abc_52155_new_n5757_; 
wire u2__abc_52155_new_n5758_; 
wire u2__abc_52155_new_n5759_; 
wire u2__abc_52155_new_n5760_; 
wire u2__abc_52155_new_n5761_; 
wire u2__abc_52155_new_n5762_; 
wire u2__abc_52155_new_n5763_; 
wire u2__abc_52155_new_n5764_; 
wire u2__abc_52155_new_n5765_; 
wire u2__abc_52155_new_n5766_; 
wire u2__abc_52155_new_n5767_; 
wire u2__abc_52155_new_n5768_; 
wire u2__abc_52155_new_n5769_; 
wire u2__abc_52155_new_n5770_; 
wire u2__abc_52155_new_n5771_; 
wire u2__abc_52155_new_n5772_; 
wire u2__abc_52155_new_n5773_; 
wire u2__abc_52155_new_n5774_; 
wire u2__abc_52155_new_n5775_; 
wire u2__abc_52155_new_n5776_; 
wire u2__abc_52155_new_n5777_; 
wire u2__abc_52155_new_n5778_; 
wire u2__abc_52155_new_n5779_; 
wire u2__abc_52155_new_n5780_; 
wire u2__abc_52155_new_n5781_; 
wire u2__abc_52155_new_n5782_; 
wire u2__abc_52155_new_n5783_; 
wire u2__abc_52155_new_n5784_; 
wire u2__abc_52155_new_n5785_; 
wire u2__abc_52155_new_n5786_; 
wire u2__abc_52155_new_n5787_; 
wire u2__abc_52155_new_n5788_; 
wire u2__abc_52155_new_n5789_; 
wire u2__abc_52155_new_n5790_; 
wire u2__abc_52155_new_n5791_; 
wire u2__abc_52155_new_n5792_; 
wire u2__abc_52155_new_n5793_; 
wire u2__abc_52155_new_n5794_; 
wire u2__abc_52155_new_n5795_; 
wire u2__abc_52155_new_n5796_; 
wire u2__abc_52155_new_n5797_; 
wire u2__abc_52155_new_n5798_; 
wire u2__abc_52155_new_n5799_; 
wire u2__abc_52155_new_n5800_; 
wire u2__abc_52155_new_n5801_; 
wire u2__abc_52155_new_n5802_; 
wire u2__abc_52155_new_n5803_; 
wire u2__abc_52155_new_n5804_; 
wire u2__abc_52155_new_n5805_; 
wire u2__abc_52155_new_n5806_; 
wire u2__abc_52155_new_n5807_; 
wire u2__abc_52155_new_n5808_; 
wire u2__abc_52155_new_n5809_; 
wire u2__abc_52155_new_n5810_; 
wire u2__abc_52155_new_n5811_; 
wire u2__abc_52155_new_n5812_; 
wire u2__abc_52155_new_n5813_; 
wire u2__abc_52155_new_n5814_; 
wire u2__abc_52155_new_n5815_; 
wire u2__abc_52155_new_n5816_; 
wire u2__abc_52155_new_n5817_; 
wire u2__abc_52155_new_n5818_; 
wire u2__abc_52155_new_n5819_; 
wire u2__abc_52155_new_n5820_; 
wire u2__abc_52155_new_n5821_; 
wire u2__abc_52155_new_n5822_; 
wire u2__abc_52155_new_n5823_; 
wire u2__abc_52155_new_n5824_; 
wire u2__abc_52155_new_n5825_; 
wire u2__abc_52155_new_n5826_; 
wire u2__abc_52155_new_n5827_; 
wire u2__abc_52155_new_n5828_; 
wire u2__abc_52155_new_n5829_; 
wire u2__abc_52155_new_n5830_; 
wire u2__abc_52155_new_n5831_; 
wire u2__abc_52155_new_n5832_; 
wire u2__abc_52155_new_n5833_; 
wire u2__abc_52155_new_n5834_; 
wire u2__abc_52155_new_n5835_; 
wire u2__abc_52155_new_n5836_; 
wire u2__abc_52155_new_n5837_; 
wire u2__abc_52155_new_n5838_; 
wire u2__abc_52155_new_n5839_; 
wire u2__abc_52155_new_n5840_; 
wire u2__abc_52155_new_n5841_; 
wire u2__abc_52155_new_n5842_; 
wire u2__abc_52155_new_n5843_; 
wire u2__abc_52155_new_n5844_; 
wire u2__abc_52155_new_n5845_; 
wire u2__abc_52155_new_n5846_; 
wire u2__abc_52155_new_n5847_; 
wire u2__abc_52155_new_n5848_; 
wire u2__abc_52155_new_n5849_; 
wire u2__abc_52155_new_n5850_; 
wire u2__abc_52155_new_n5851_; 
wire u2__abc_52155_new_n5852_; 
wire u2__abc_52155_new_n5853_; 
wire u2__abc_52155_new_n5854_; 
wire u2__abc_52155_new_n5855_; 
wire u2__abc_52155_new_n5856_; 
wire u2__abc_52155_new_n5857_; 
wire u2__abc_52155_new_n5858_; 
wire u2__abc_52155_new_n5859_; 
wire u2__abc_52155_new_n5860_; 
wire u2__abc_52155_new_n5861_; 
wire u2__abc_52155_new_n5862_; 
wire u2__abc_52155_new_n5863_; 
wire u2__abc_52155_new_n5864_; 
wire u2__abc_52155_new_n5865_; 
wire u2__abc_52155_new_n5866_; 
wire u2__abc_52155_new_n5867_; 
wire u2__abc_52155_new_n5868_; 
wire u2__abc_52155_new_n5869_; 
wire u2__abc_52155_new_n5870_; 
wire u2__abc_52155_new_n5871_; 
wire u2__abc_52155_new_n5872_; 
wire u2__abc_52155_new_n5873_; 
wire u2__abc_52155_new_n5874_; 
wire u2__abc_52155_new_n5875_; 
wire u2__abc_52155_new_n5876_; 
wire u2__abc_52155_new_n5877_; 
wire u2__abc_52155_new_n5878_; 
wire u2__abc_52155_new_n5879_; 
wire u2__abc_52155_new_n5880_; 
wire u2__abc_52155_new_n5881_; 
wire u2__abc_52155_new_n5882_; 
wire u2__abc_52155_new_n5883_; 
wire u2__abc_52155_new_n5884_; 
wire u2__abc_52155_new_n5885_; 
wire u2__abc_52155_new_n5886_; 
wire u2__abc_52155_new_n5887_; 
wire u2__abc_52155_new_n5888_; 
wire u2__abc_52155_new_n5889_; 
wire u2__abc_52155_new_n5890_; 
wire u2__abc_52155_new_n5891_; 
wire u2__abc_52155_new_n5892_; 
wire u2__abc_52155_new_n5893_; 
wire u2__abc_52155_new_n5894_; 
wire u2__abc_52155_new_n5895_; 
wire u2__abc_52155_new_n5896_; 
wire u2__abc_52155_new_n5897_; 
wire u2__abc_52155_new_n5898_; 
wire u2__abc_52155_new_n5899_; 
wire u2__abc_52155_new_n5900_; 
wire u2__abc_52155_new_n5901_; 
wire u2__abc_52155_new_n5902_; 
wire u2__abc_52155_new_n5903_; 
wire u2__abc_52155_new_n5904_; 
wire u2__abc_52155_new_n5905_; 
wire u2__abc_52155_new_n5906_; 
wire u2__abc_52155_new_n5907_; 
wire u2__abc_52155_new_n5908_; 
wire u2__abc_52155_new_n5909_; 
wire u2__abc_52155_new_n5910_; 
wire u2__abc_52155_new_n5911_; 
wire u2__abc_52155_new_n5912_; 
wire u2__abc_52155_new_n5913_; 
wire u2__abc_52155_new_n5914_; 
wire u2__abc_52155_new_n5915_; 
wire u2__abc_52155_new_n5916_; 
wire u2__abc_52155_new_n5917_; 
wire u2__abc_52155_new_n5918_; 
wire u2__abc_52155_new_n5919_; 
wire u2__abc_52155_new_n5920_; 
wire u2__abc_52155_new_n5921_; 
wire u2__abc_52155_new_n5922_; 
wire u2__abc_52155_new_n5923_; 
wire u2__abc_52155_new_n5924_; 
wire u2__abc_52155_new_n5925_; 
wire u2__abc_52155_new_n5926_; 
wire u2__abc_52155_new_n5927_; 
wire u2__abc_52155_new_n5928_; 
wire u2__abc_52155_new_n5929_; 
wire u2__abc_52155_new_n5930_; 
wire u2__abc_52155_new_n5931_; 
wire u2__abc_52155_new_n5932_; 
wire u2__abc_52155_new_n5933_; 
wire u2__abc_52155_new_n5934_; 
wire u2__abc_52155_new_n5935_; 
wire u2__abc_52155_new_n5936_; 
wire u2__abc_52155_new_n5937_; 
wire u2__abc_52155_new_n5938_; 
wire u2__abc_52155_new_n5939_; 
wire u2__abc_52155_new_n5940_; 
wire u2__abc_52155_new_n5941_; 
wire u2__abc_52155_new_n5942_; 
wire u2__abc_52155_new_n5943_; 
wire u2__abc_52155_new_n5944_; 
wire u2__abc_52155_new_n5945_; 
wire u2__abc_52155_new_n5946_; 
wire u2__abc_52155_new_n5947_; 
wire u2__abc_52155_new_n5948_; 
wire u2__abc_52155_new_n5949_; 
wire u2__abc_52155_new_n5950_; 
wire u2__abc_52155_new_n5951_; 
wire u2__abc_52155_new_n5952_; 
wire u2__abc_52155_new_n5953_; 
wire u2__abc_52155_new_n5954_; 
wire u2__abc_52155_new_n5955_; 
wire u2__abc_52155_new_n5956_; 
wire u2__abc_52155_new_n5957_; 
wire u2__abc_52155_new_n5958_; 
wire u2__abc_52155_new_n5959_; 
wire u2__abc_52155_new_n5960_; 
wire u2__abc_52155_new_n5961_; 
wire u2__abc_52155_new_n5962_; 
wire u2__abc_52155_new_n5963_; 
wire u2__abc_52155_new_n5964_; 
wire u2__abc_52155_new_n5965_; 
wire u2__abc_52155_new_n5966_; 
wire u2__abc_52155_new_n5967_; 
wire u2__abc_52155_new_n5968_; 
wire u2__abc_52155_new_n5969_; 
wire u2__abc_52155_new_n5970_; 
wire u2__abc_52155_new_n5971_; 
wire u2__abc_52155_new_n5972_; 
wire u2__abc_52155_new_n5973_; 
wire u2__abc_52155_new_n5974_; 
wire u2__abc_52155_new_n5975_; 
wire u2__abc_52155_new_n5976_; 
wire u2__abc_52155_new_n5977_; 
wire u2__abc_52155_new_n5978_; 
wire u2__abc_52155_new_n5979_; 
wire u2__abc_52155_new_n5980_; 
wire u2__abc_52155_new_n5981_; 
wire u2__abc_52155_new_n5982_; 
wire u2__abc_52155_new_n5983_; 
wire u2__abc_52155_new_n5984_; 
wire u2__abc_52155_new_n5985_; 
wire u2__abc_52155_new_n5986_; 
wire u2__abc_52155_new_n5987_; 
wire u2__abc_52155_new_n5988_; 
wire u2__abc_52155_new_n5989_; 
wire u2__abc_52155_new_n5990_; 
wire u2__abc_52155_new_n5991_; 
wire u2__abc_52155_new_n5992_; 
wire u2__abc_52155_new_n5993_; 
wire u2__abc_52155_new_n5994_; 
wire u2__abc_52155_new_n5995_; 
wire u2__abc_52155_new_n5996_; 
wire u2__abc_52155_new_n5997_; 
wire u2__abc_52155_new_n5998_; 
wire u2__abc_52155_new_n5999_; 
wire u2__abc_52155_new_n6000_; 
wire u2__abc_52155_new_n6001_; 
wire u2__abc_52155_new_n6002_; 
wire u2__abc_52155_new_n6003_; 
wire u2__abc_52155_new_n6004_; 
wire u2__abc_52155_new_n6005_; 
wire u2__abc_52155_new_n6006_; 
wire u2__abc_52155_new_n6007_; 
wire u2__abc_52155_new_n6008_; 
wire u2__abc_52155_new_n6009_; 
wire u2__abc_52155_new_n6010_; 
wire u2__abc_52155_new_n6011_; 
wire u2__abc_52155_new_n6012_; 
wire u2__abc_52155_new_n6013_; 
wire u2__abc_52155_new_n6014_; 
wire u2__abc_52155_new_n6015_; 
wire u2__abc_52155_new_n6016_; 
wire u2__abc_52155_new_n6017_; 
wire u2__abc_52155_new_n6018_; 
wire u2__abc_52155_new_n6019_; 
wire u2__abc_52155_new_n6020_; 
wire u2__abc_52155_new_n6021_; 
wire u2__abc_52155_new_n6022_; 
wire u2__abc_52155_new_n6023_; 
wire u2__abc_52155_new_n6024_; 
wire u2__abc_52155_new_n6025_; 
wire u2__abc_52155_new_n6026_; 
wire u2__abc_52155_new_n6027_; 
wire u2__abc_52155_new_n6028_; 
wire u2__abc_52155_new_n6029_; 
wire u2__abc_52155_new_n6030_; 
wire u2__abc_52155_new_n6031_; 
wire u2__abc_52155_new_n6032_; 
wire u2__abc_52155_new_n6033_; 
wire u2__abc_52155_new_n6034_; 
wire u2__abc_52155_new_n6035_; 
wire u2__abc_52155_new_n6036_; 
wire u2__abc_52155_new_n6037_; 
wire u2__abc_52155_new_n6038_; 
wire u2__abc_52155_new_n6039_; 
wire u2__abc_52155_new_n6040_; 
wire u2__abc_52155_new_n6041_; 
wire u2__abc_52155_new_n6042_; 
wire u2__abc_52155_new_n6043_; 
wire u2__abc_52155_new_n6044_; 
wire u2__abc_52155_new_n6045_; 
wire u2__abc_52155_new_n6046_; 
wire u2__abc_52155_new_n6047_; 
wire u2__abc_52155_new_n6048_; 
wire u2__abc_52155_new_n6049_; 
wire u2__abc_52155_new_n6050_; 
wire u2__abc_52155_new_n6051_; 
wire u2__abc_52155_new_n6052_; 
wire u2__abc_52155_new_n6053_; 
wire u2__abc_52155_new_n6054_; 
wire u2__abc_52155_new_n6055_; 
wire u2__abc_52155_new_n6056_; 
wire u2__abc_52155_new_n6057_; 
wire u2__abc_52155_new_n6058_; 
wire u2__abc_52155_new_n6059_; 
wire u2__abc_52155_new_n6060_; 
wire u2__abc_52155_new_n6061_; 
wire u2__abc_52155_new_n6062_; 
wire u2__abc_52155_new_n6063_; 
wire u2__abc_52155_new_n6064_; 
wire u2__abc_52155_new_n6065_; 
wire u2__abc_52155_new_n6066_; 
wire u2__abc_52155_new_n6067_; 
wire u2__abc_52155_new_n6068_; 
wire u2__abc_52155_new_n6069_; 
wire u2__abc_52155_new_n6070_; 
wire u2__abc_52155_new_n6071_; 
wire u2__abc_52155_new_n6072_; 
wire u2__abc_52155_new_n6073_; 
wire u2__abc_52155_new_n6074_; 
wire u2__abc_52155_new_n6075_; 
wire u2__abc_52155_new_n6076_; 
wire u2__abc_52155_new_n6077_; 
wire u2__abc_52155_new_n6078_; 
wire u2__abc_52155_new_n6079_; 
wire u2__abc_52155_new_n6080_; 
wire u2__abc_52155_new_n6081_; 
wire u2__abc_52155_new_n6082_; 
wire u2__abc_52155_new_n6083_; 
wire u2__abc_52155_new_n6084_; 
wire u2__abc_52155_new_n6085_; 
wire u2__abc_52155_new_n6086_; 
wire u2__abc_52155_new_n6087_; 
wire u2__abc_52155_new_n6088_; 
wire u2__abc_52155_new_n6089_; 
wire u2__abc_52155_new_n6090_; 
wire u2__abc_52155_new_n6091_; 
wire u2__abc_52155_new_n6092_; 
wire u2__abc_52155_new_n6093_; 
wire u2__abc_52155_new_n6094_; 
wire u2__abc_52155_new_n6095_; 
wire u2__abc_52155_new_n6096_; 
wire u2__abc_52155_new_n6097_; 
wire u2__abc_52155_new_n6098_; 
wire u2__abc_52155_new_n6099_; 
wire u2__abc_52155_new_n6100_; 
wire u2__abc_52155_new_n6101_; 
wire u2__abc_52155_new_n6102_; 
wire u2__abc_52155_new_n6103_; 
wire u2__abc_52155_new_n6104_; 
wire u2__abc_52155_new_n6105_; 
wire u2__abc_52155_new_n6106_; 
wire u2__abc_52155_new_n6107_; 
wire u2__abc_52155_new_n6108_; 
wire u2__abc_52155_new_n6109_; 
wire u2__abc_52155_new_n6110_; 
wire u2__abc_52155_new_n6111_; 
wire u2__abc_52155_new_n6112_; 
wire u2__abc_52155_new_n6113_; 
wire u2__abc_52155_new_n6114_; 
wire u2__abc_52155_new_n6115_; 
wire u2__abc_52155_new_n6116_; 
wire u2__abc_52155_new_n6117_; 
wire u2__abc_52155_new_n6118_; 
wire u2__abc_52155_new_n6119_; 
wire u2__abc_52155_new_n6120_; 
wire u2__abc_52155_new_n6121_; 
wire u2__abc_52155_new_n6122_; 
wire u2__abc_52155_new_n6123_; 
wire u2__abc_52155_new_n6124_; 
wire u2__abc_52155_new_n6125_; 
wire u2__abc_52155_new_n6126_; 
wire u2__abc_52155_new_n6127_; 
wire u2__abc_52155_new_n6128_; 
wire u2__abc_52155_new_n6129_; 
wire u2__abc_52155_new_n6130_; 
wire u2__abc_52155_new_n6131_; 
wire u2__abc_52155_new_n6132_; 
wire u2__abc_52155_new_n6133_; 
wire u2__abc_52155_new_n6134_; 
wire u2__abc_52155_new_n6135_; 
wire u2__abc_52155_new_n6136_; 
wire u2__abc_52155_new_n6137_; 
wire u2__abc_52155_new_n6138_; 
wire u2__abc_52155_new_n6139_; 
wire u2__abc_52155_new_n6140_; 
wire u2__abc_52155_new_n6141_; 
wire u2__abc_52155_new_n6142_; 
wire u2__abc_52155_new_n6143_; 
wire u2__abc_52155_new_n6144_; 
wire u2__abc_52155_new_n6145_; 
wire u2__abc_52155_new_n6146_; 
wire u2__abc_52155_new_n6147_; 
wire u2__abc_52155_new_n6148_; 
wire u2__abc_52155_new_n6149_; 
wire u2__abc_52155_new_n6150_; 
wire u2__abc_52155_new_n6151_; 
wire u2__abc_52155_new_n6152_; 
wire u2__abc_52155_new_n6153_; 
wire u2__abc_52155_new_n6154_; 
wire u2__abc_52155_new_n6155_; 
wire u2__abc_52155_new_n6156_; 
wire u2__abc_52155_new_n6157_; 
wire u2__abc_52155_new_n6158_; 
wire u2__abc_52155_new_n6159_; 
wire u2__abc_52155_new_n6160_; 
wire u2__abc_52155_new_n6161_; 
wire u2__abc_52155_new_n6162_; 
wire u2__abc_52155_new_n6163_; 
wire u2__abc_52155_new_n6164_; 
wire u2__abc_52155_new_n6165_; 
wire u2__abc_52155_new_n6166_; 
wire u2__abc_52155_new_n6167_; 
wire u2__abc_52155_new_n6168_; 
wire u2__abc_52155_new_n6169_; 
wire u2__abc_52155_new_n6170_; 
wire u2__abc_52155_new_n6171_; 
wire u2__abc_52155_new_n6172_; 
wire u2__abc_52155_new_n6173_; 
wire u2__abc_52155_new_n6174_; 
wire u2__abc_52155_new_n6175_; 
wire u2__abc_52155_new_n6176_; 
wire u2__abc_52155_new_n6177_; 
wire u2__abc_52155_new_n6178_; 
wire u2__abc_52155_new_n6179_; 
wire u2__abc_52155_new_n6180_; 
wire u2__abc_52155_new_n6181_; 
wire u2__abc_52155_new_n6182_; 
wire u2__abc_52155_new_n6183_; 
wire u2__abc_52155_new_n6184_; 
wire u2__abc_52155_new_n6185_; 
wire u2__abc_52155_new_n6186_; 
wire u2__abc_52155_new_n6187_; 
wire u2__abc_52155_new_n6188_; 
wire u2__abc_52155_new_n6189_; 
wire u2__abc_52155_new_n6190_; 
wire u2__abc_52155_new_n6191_; 
wire u2__abc_52155_new_n6192_; 
wire u2__abc_52155_new_n6193_; 
wire u2__abc_52155_new_n6194_; 
wire u2__abc_52155_new_n6195_; 
wire u2__abc_52155_new_n6196_; 
wire u2__abc_52155_new_n6197_; 
wire u2__abc_52155_new_n6198_; 
wire u2__abc_52155_new_n6199_; 
wire u2__abc_52155_new_n6200_; 
wire u2__abc_52155_new_n6201_; 
wire u2__abc_52155_new_n6202_; 
wire u2__abc_52155_new_n6203_; 
wire u2__abc_52155_new_n6204_; 
wire u2__abc_52155_new_n6205_; 
wire u2__abc_52155_new_n6206_; 
wire u2__abc_52155_new_n6207_; 
wire u2__abc_52155_new_n6208_; 
wire u2__abc_52155_new_n6209_; 
wire u2__abc_52155_new_n6210_; 
wire u2__abc_52155_new_n6211_; 
wire u2__abc_52155_new_n6212_; 
wire u2__abc_52155_new_n6213_; 
wire u2__abc_52155_new_n6214_; 
wire u2__abc_52155_new_n6215_; 
wire u2__abc_52155_new_n6216_; 
wire u2__abc_52155_new_n6217_; 
wire u2__abc_52155_new_n6218_; 
wire u2__abc_52155_new_n6219_; 
wire u2__abc_52155_new_n6220_; 
wire u2__abc_52155_new_n6221_; 
wire u2__abc_52155_new_n6222_; 
wire u2__abc_52155_new_n6223_; 
wire u2__abc_52155_new_n6224_; 
wire u2__abc_52155_new_n6225_; 
wire u2__abc_52155_new_n6226_; 
wire u2__abc_52155_new_n6227_; 
wire u2__abc_52155_new_n6228_; 
wire u2__abc_52155_new_n6229_; 
wire u2__abc_52155_new_n6230_; 
wire u2__abc_52155_new_n6231_; 
wire u2__abc_52155_new_n6232_; 
wire u2__abc_52155_new_n6233_; 
wire u2__abc_52155_new_n6234_; 
wire u2__abc_52155_new_n6235_; 
wire u2__abc_52155_new_n6236_; 
wire u2__abc_52155_new_n6237_; 
wire u2__abc_52155_new_n6238_; 
wire u2__abc_52155_new_n6239_; 
wire u2__abc_52155_new_n6240_; 
wire u2__abc_52155_new_n6241_; 
wire u2__abc_52155_new_n6242_; 
wire u2__abc_52155_new_n6243_; 
wire u2__abc_52155_new_n6244_; 
wire u2__abc_52155_new_n6245_; 
wire u2__abc_52155_new_n6246_; 
wire u2__abc_52155_new_n6247_; 
wire u2__abc_52155_new_n6248_; 
wire u2__abc_52155_new_n6249_; 
wire u2__abc_52155_new_n6250_; 
wire u2__abc_52155_new_n6251_; 
wire u2__abc_52155_new_n6252_; 
wire u2__abc_52155_new_n6253_; 
wire u2__abc_52155_new_n6254_; 
wire u2__abc_52155_new_n6255_; 
wire u2__abc_52155_new_n6256_; 
wire u2__abc_52155_new_n6257_; 
wire u2__abc_52155_new_n6258_; 
wire u2__abc_52155_new_n6259_; 
wire u2__abc_52155_new_n6260_; 
wire u2__abc_52155_new_n6261_; 
wire u2__abc_52155_new_n6262_; 
wire u2__abc_52155_new_n6263_; 
wire u2__abc_52155_new_n6264_; 
wire u2__abc_52155_new_n6265_; 
wire u2__abc_52155_new_n6266_; 
wire u2__abc_52155_new_n6267_; 
wire u2__abc_52155_new_n6268_; 
wire u2__abc_52155_new_n6269_; 
wire u2__abc_52155_new_n6270_; 
wire u2__abc_52155_new_n6271_; 
wire u2__abc_52155_new_n6272_; 
wire u2__abc_52155_new_n6273_; 
wire u2__abc_52155_new_n6274_; 
wire u2__abc_52155_new_n6275_; 
wire u2__abc_52155_new_n6276_; 
wire u2__abc_52155_new_n6277_; 
wire u2__abc_52155_new_n6278_; 
wire u2__abc_52155_new_n6279_; 
wire u2__abc_52155_new_n6280_; 
wire u2__abc_52155_new_n6281_; 
wire u2__abc_52155_new_n6282_; 
wire u2__abc_52155_new_n6283_; 
wire u2__abc_52155_new_n6284_; 
wire u2__abc_52155_new_n6285_; 
wire u2__abc_52155_new_n6286_; 
wire u2__abc_52155_new_n6287_; 
wire u2__abc_52155_new_n6288_; 
wire u2__abc_52155_new_n6289_; 
wire u2__abc_52155_new_n6290_; 
wire u2__abc_52155_new_n6291_; 
wire u2__abc_52155_new_n6292_; 
wire u2__abc_52155_new_n6293_; 
wire u2__abc_52155_new_n6294_; 
wire u2__abc_52155_new_n6295_; 
wire u2__abc_52155_new_n6296_; 
wire u2__abc_52155_new_n6297_; 
wire u2__abc_52155_new_n6298_; 
wire u2__abc_52155_new_n6299_; 
wire u2__abc_52155_new_n6300_; 
wire u2__abc_52155_new_n6301_; 
wire u2__abc_52155_new_n6302_; 
wire u2__abc_52155_new_n6303_; 
wire u2__abc_52155_new_n6304_; 
wire u2__abc_52155_new_n6305_; 
wire u2__abc_52155_new_n6306_; 
wire u2__abc_52155_new_n6307_; 
wire u2__abc_52155_new_n6308_; 
wire u2__abc_52155_new_n6309_; 
wire u2__abc_52155_new_n6310_; 
wire u2__abc_52155_new_n6311_; 
wire u2__abc_52155_new_n6312_; 
wire u2__abc_52155_new_n6313_; 
wire u2__abc_52155_new_n6314_; 
wire u2__abc_52155_new_n6315_; 
wire u2__abc_52155_new_n6316_; 
wire u2__abc_52155_new_n6317_; 
wire u2__abc_52155_new_n6318_; 
wire u2__abc_52155_new_n6319_; 
wire u2__abc_52155_new_n6320_; 
wire u2__abc_52155_new_n6321_; 
wire u2__abc_52155_new_n6322_; 
wire u2__abc_52155_new_n6323_; 
wire u2__abc_52155_new_n6324_; 
wire u2__abc_52155_new_n6325_; 
wire u2__abc_52155_new_n6326_; 
wire u2__abc_52155_new_n6327_; 
wire u2__abc_52155_new_n6328_; 
wire u2__abc_52155_new_n6329_; 
wire u2__abc_52155_new_n6330_; 
wire u2__abc_52155_new_n6331_; 
wire u2__abc_52155_new_n6332_; 
wire u2__abc_52155_new_n6333_; 
wire u2__abc_52155_new_n6334_; 
wire u2__abc_52155_new_n6335_; 
wire u2__abc_52155_new_n6336_; 
wire u2__abc_52155_new_n6337_; 
wire u2__abc_52155_new_n6338_; 
wire u2__abc_52155_new_n6339_; 
wire u2__abc_52155_new_n6340_; 
wire u2__abc_52155_new_n6341_; 
wire u2__abc_52155_new_n6342_; 
wire u2__abc_52155_new_n6343_; 
wire u2__abc_52155_new_n6344_; 
wire u2__abc_52155_new_n6345_; 
wire u2__abc_52155_new_n6346_; 
wire u2__abc_52155_new_n6347_; 
wire u2__abc_52155_new_n6348_; 
wire u2__abc_52155_new_n6349_; 
wire u2__abc_52155_new_n6350_; 
wire u2__abc_52155_new_n6351_; 
wire u2__abc_52155_new_n6352_; 
wire u2__abc_52155_new_n6353_; 
wire u2__abc_52155_new_n6354_; 
wire u2__abc_52155_new_n6355_; 
wire u2__abc_52155_new_n6356_; 
wire u2__abc_52155_new_n6357_; 
wire u2__abc_52155_new_n6358_; 
wire u2__abc_52155_new_n6359_; 
wire u2__abc_52155_new_n6360_; 
wire u2__abc_52155_new_n6361_; 
wire u2__abc_52155_new_n6362_; 
wire u2__abc_52155_new_n6363_; 
wire u2__abc_52155_new_n6364_; 
wire u2__abc_52155_new_n6365_; 
wire u2__abc_52155_new_n6366_; 
wire u2__abc_52155_new_n6367_; 
wire u2__abc_52155_new_n6368_; 
wire u2__abc_52155_new_n6369_; 
wire u2__abc_52155_new_n6370_; 
wire u2__abc_52155_new_n6371_; 
wire u2__abc_52155_new_n6372_; 
wire u2__abc_52155_new_n6373_; 
wire u2__abc_52155_new_n6374_; 
wire u2__abc_52155_new_n6375_; 
wire u2__abc_52155_new_n6376_; 
wire u2__abc_52155_new_n6377_; 
wire u2__abc_52155_new_n6378_; 
wire u2__abc_52155_new_n6379_; 
wire u2__abc_52155_new_n6380_; 
wire u2__abc_52155_new_n6381_; 
wire u2__abc_52155_new_n6382_; 
wire u2__abc_52155_new_n6383_; 
wire u2__abc_52155_new_n6384_; 
wire u2__abc_52155_new_n6385_; 
wire u2__abc_52155_new_n6386_; 
wire u2__abc_52155_new_n6387_; 
wire u2__abc_52155_new_n6388_; 
wire u2__abc_52155_new_n6389_; 
wire u2__abc_52155_new_n6390_; 
wire u2__abc_52155_new_n6391_; 
wire u2__abc_52155_new_n6392_; 
wire u2__abc_52155_new_n6393_; 
wire u2__abc_52155_new_n6394_; 
wire u2__abc_52155_new_n6395_; 
wire u2__abc_52155_new_n6396_; 
wire u2__abc_52155_new_n6397_; 
wire u2__abc_52155_new_n6398_; 
wire u2__abc_52155_new_n6399_; 
wire u2__abc_52155_new_n6400_; 
wire u2__abc_52155_new_n6401_; 
wire u2__abc_52155_new_n6402_; 
wire u2__abc_52155_new_n6403_; 
wire u2__abc_52155_new_n6404_; 
wire u2__abc_52155_new_n6405_; 
wire u2__abc_52155_new_n6406_; 
wire u2__abc_52155_new_n6407_; 
wire u2__abc_52155_new_n6408_; 
wire u2__abc_52155_new_n6409_; 
wire u2__abc_52155_new_n6410_; 
wire u2__abc_52155_new_n6411_; 
wire u2__abc_52155_new_n6412_; 
wire u2__abc_52155_new_n6413_; 
wire u2__abc_52155_new_n6414_; 
wire u2__abc_52155_new_n6415_; 
wire u2__abc_52155_new_n6416_; 
wire u2__abc_52155_new_n6417_; 
wire u2__abc_52155_new_n6418_; 
wire u2__abc_52155_new_n6419_; 
wire u2__abc_52155_new_n6420_; 
wire u2__abc_52155_new_n6421_; 
wire u2__abc_52155_new_n6422_; 
wire u2__abc_52155_new_n6423_; 
wire u2__abc_52155_new_n6424_; 
wire u2__abc_52155_new_n6425_; 
wire u2__abc_52155_new_n6426_; 
wire u2__abc_52155_new_n6427_; 
wire u2__abc_52155_new_n6428_; 
wire u2__abc_52155_new_n6429_; 
wire u2__abc_52155_new_n6430_; 
wire u2__abc_52155_new_n6431_; 
wire u2__abc_52155_new_n6432_; 
wire u2__abc_52155_new_n6433_; 
wire u2__abc_52155_new_n6434_; 
wire u2__abc_52155_new_n6435_; 
wire u2__abc_52155_new_n6436_; 
wire u2__abc_52155_new_n6437_; 
wire u2__abc_52155_new_n6438_; 
wire u2__abc_52155_new_n6439_; 
wire u2__abc_52155_new_n6440_; 
wire u2__abc_52155_new_n6441_; 
wire u2__abc_52155_new_n6442_; 
wire u2__abc_52155_new_n6443_; 
wire u2__abc_52155_new_n6444_; 
wire u2__abc_52155_new_n6445_; 
wire u2__abc_52155_new_n6446_; 
wire u2__abc_52155_new_n6447_; 
wire u2__abc_52155_new_n6448_; 
wire u2__abc_52155_new_n6449_; 
wire u2__abc_52155_new_n6450_; 
wire u2__abc_52155_new_n6451_; 
wire u2__abc_52155_new_n6452_; 
wire u2__abc_52155_new_n6453_; 
wire u2__abc_52155_new_n6454_; 
wire u2__abc_52155_new_n6455_; 
wire u2__abc_52155_new_n6456_; 
wire u2__abc_52155_new_n6457_; 
wire u2__abc_52155_new_n6458_; 
wire u2__abc_52155_new_n6459_; 
wire u2__abc_52155_new_n6460_; 
wire u2__abc_52155_new_n6461_; 
wire u2__abc_52155_new_n6462_; 
wire u2__abc_52155_new_n6463_; 
wire u2__abc_52155_new_n6464_; 
wire u2__abc_52155_new_n6465_; 
wire u2__abc_52155_new_n6466_; 
wire u2__abc_52155_new_n6467_; 
wire u2__abc_52155_new_n6468_; 
wire u2__abc_52155_new_n6469_; 
wire u2__abc_52155_new_n6470_; 
wire u2__abc_52155_new_n6471_; 
wire u2__abc_52155_new_n6472_; 
wire u2__abc_52155_new_n6473_; 
wire u2__abc_52155_new_n6474_; 
wire u2__abc_52155_new_n6475_; 
wire u2__abc_52155_new_n6476_; 
wire u2__abc_52155_new_n6477_; 
wire u2__abc_52155_new_n6478_; 
wire u2__abc_52155_new_n6479_; 
wire u2__abc_52155_new_n6480_; 
wire u2__abc_52155_new_n6481_; 
wire u2__abc_52155_new_n6482_; 
wire u2__abc_52155_new_n6483_; 
wire u2__abc_52155_new_n6484_; 
wire u2__abc_52155_new_n6485_; 
wire u2__abc_52155_new_n6486_; 
wire u2__abc_52155_new_n6487_; 
wire u2__abc_52155_new_n6488_; 
wire u2__abc_52155_new_n6489_; 
wire u2__abc_52155_new_n6490_; 
wire u2__abc_52155_new_n6491_; 
wire u2__abc_52155_new_n6492_; 
wire u2__abc_52155_new_n6493_; 
wire u2__abc_52155_new_n6494_; 
wire u2__abc_52155_new_n6495_; 
wire u2__abc_52155_new_n6496_; 
wire u2__abc_52155_new_n6497_; 
wire u2__abc_52155_new_n6498_; 
wire u2__abc_52155_new_n6499_; 
wire u2__abc_52155_new_n6500_; 
wire u2__abc_52155_new_n6501_; 
wire u2__abc_52155_new_n6502_; 
wire u2__abc_52155_new_n6503_; 
wire u2__abc_52155_new_n6504_; 
wire u2__abc_52155_new_n6505_; 
wire u2__abc_52155_new_n6506_; 
wire u2__abc_52155_new_n6507_; 
wire u2__abc_52155_new_n6508_; 
wire u2__abc_52155_new_n6509_; 
wire u2__abc_52155_new_n6510_; 
wire u2__abc_52155_new_n6511_; 
wire u2__abc_52155_new_n6512_; 
wire u2__abc_52155_new_n6513_; 
wire u2__abc_52155_new_n6514_; 
wire u2__abc_52155_new_n6515_; 
wire u2__abc_52155_new_n6516_; 
wire u2__abc_52155_new_n6517_; 
wire u2__abc_52155_new_n6518_; 
wire u2__abc_52155_new_n6519_; 
wire u2__abc_52155_new_n6520_; 
wire u2__abc_52155_new_n6521_; 
wire u2__abc_52155_new_n6522_; 
wire u2__abc_52155_new_n6523_; 
wire u2__abc_52155_new_n6524_; 
wire u2__abc_52155_new_n6525_; 
wire u2__abc_52155_new_n6526_; 
wire u2__abc_52155_new_n6527_; 
wire u2__abc_52155_new_n6528_; 
wire u2__abc_52155_new_n6529_; 
wire u2__abc_52155_new_n6530_; 
wire u2__abc_52155_new_n6531_; 
wire u2__abc_52155_new_n6532_; 
wire u2__abc_52155_new_n6533_; 
wire u2__abc_52155_new_n6534_; 
wire u2__abc_52155_new_n6535_; 
wire u2__abc_52155_new_n6536_; 
wire u2__abc_52155_new_n6537_; 
wire u2__abc_52155_new_n6538_; 
wire u2__abc_52155_new_n6539_; 
wire u2__abc_52155_new_n6540_; 
wire u2__abc_52155_new_n6541_; 
wire u2__abc_52155_new_n6542_; 
wire u2__abc_52155_new_n6543_; 
wire u2__abc_52155_new_n6544_; 
wire u2__abc_52155_new_n6545_; 
wire u2__abc_52155_new_n6546_; 
wire u2__abc_52155_new_n6547_; 
wire u2__abc_52155_new_n6548_; 
wire u2__abc_52155_new_n6549_; 
wire u2__abc_52155_new_n6550_; 
wire u2__abc_52155_new_n6551_; 
wire u2__abc_52155_new_n6552_; 
wire u2__abc_52155_new_n6553_; 
wire u2__abc_52155_new_n6554_; 
wire u2__abc_52155_new_n6555_; 
wire u2__abc_52155_new_n6556_; 
wire u2__abc_52155_new_n6557_; 
wire u2__abc_52155_new_n6558_; 
wire u2__abc_52155_new_n6559_; 
wire u2__abc_52155_new_n6560_; 
wire u2__abc_52155_new_n6561_; 
wire u2__abc_52155_new_n6562_; 
wire u2__abc_52155_new_n6563_; 
wire u2__abc_52155_new_n6564_; 
wire u2__abc_52155_new_n6565_; 
wire u2__abc_52155_new_n6566_; 
wire u2__abc_52155_new_n6567_; 
wire u2__abc_52155_new_n6568_; 
wire u2__abc_52155_new_n6569_; 
wire u2__abc_52155_new_n6570_; 
wire u2__abc_52155_new_n6571_; 
wire u2__abc_52155_new_n6572_; 
wire u2__abc_52155_new_n6573_; 
wire u2__abc_52155_new_n6574_; 
wire u2__abc_52155_new_n6575_; 
wire u2__abc_52155_new_n6576_; 
wire u2__abc_52155_new_n6577_; 
wire u2__abc_52155_new_n6578_; 
wire u2__abc_52155_new_n6579_; 
wire u2__abc_52155_new_n6580_; 
wire u2__abc_52155_new_n6581_; 
wire u2__abc_52155_new_n6582_; 
wire u2__abc_52155_new_n6583_; 
wire u2__abc_52155_new_n6584_; 
wire u2__abc_52155_new_n6585_; 
wire u2__abc_52155_new_n6586_; 
wire u2__abc_52155_new_n6587_; 
wire u2__abc_52155_new_n6588_; 
wire u2__abc_52155_new_n6589_; 
wire u2__abc_52155_new_n6590_; 
wire u2__abc_52155_new_n6591_; 
wire u2__abc_52155_new_n6592_; 
wire u2__abc_52155_new_n6593_; 
wire u2__abc_52155_new_n6594_; 
wire u2__abc_52155_new_n6595_; 
wire u2__abc_52155_new_n6596_; 
wire u2__abc_52155_new_n6597_; 
wire u2__abc_52155_new_n6598_; 
wire u2__abc_52155_new_n6599_; 
wire u2__abc_52155_new_n6600_; 
wire u2__abc_52155_new_n6601_; 
wire u2__abc_52155_new_n6602_; 
wire u2__abc_52155_new_n6603_; 
wire u2__abc_52155_new_n6604_; 
wire u2__abc_52155_new_n6605_; 
wire u2__abc_52155_new_n6606_; 
wire u2__abc_52155_new_n6607_; 
wire u2__abc_52155_new_n6608_; 
wire u2__abc_52155_new_n6609_; 
wire u2__abc_52155_new_n6610_; 
wire u2__abc_52155_new_n6611_; 
wire u2__abc_52155_new_n6612_; 
wire u2__abc_52155_new_n6613_; 
wire u2__abc_52155_new_n6614_; 
wire u2__abc_52155_new_n6615_; 
wire u2__abc_52155_new_n6616_; 
wire u2__abc_52155_new_n6617_; 
wire u2__abc_52155_new_n6618_; 
wire u2__abc_52155_new_n6619_; 
wire u2__abc_52155_new_n6620_; 
wire u2__abc_52155_new_n6621_; 
wire u2__abc_52155_new_n6622_; 
wire u2__abc_52155_new_n6623_; 
wire u2__abc_52155_new_n6624_; 
wire u2__abc_52155_new_n6625_; 
wire u2__abc_52155_new_n6626_; 
wire u2__abc_52155_new_n6627_; 
wire u2__abc_52155_new_n6628_; 
wire u2__abc_52155_new_n6629_; 
wire u2__abc_52155_new_n6630_; 
wire u2__abc_52155_new_n6631_; 
wire u2__abc_52155_new_n6632_; 
wire u2__abc_52155_new_n6633_; 
wire u2__abc_52155_new_n6634_; 
wire u2__abc_52155_new_n6635_; 
wire u2__abc_52155_new_n6636_; 
wire u2__abc_52155_new_n6637_; 
wire u2__abc_52155_new_n6638_; 
wire u2__abc_52155_new_n6639_; 
wire u2__abc_52155_new_n6640_; 
wire u2__abc_52155_new_n6641_; 
wire u2__abc_52155_new_n6642_; 
wire u2__abc_52155_new_n6643_; 
wire u2__abc_52155_new_n6644_; 
wire u2__abc_52155_new_n6645_; 
wire u2__abc_52155_new_n6646_; 
wire u2__abc_52155_new_n6647_; 
wire u2__abc_52155_new_n6648_; 
wire u2__abc_52155_new_n6649_; 
wire u2__abc_52155_new_n6650_; 
wire u2__abc_52155_new_n6651_; 
wire u2__abc_52155_new_n6652_; 
wire u2__abc_52155_new_n6653_; 
wire u2__abc_52155_new_n6654_; 
wire u2__abc_52155_new_n6655_; 
wire u2__abc_52155_new_n6656_; 
wire u2__abc_52155_new_n6657_; 
wire u2__abc_52155_new_n6658_; 
wire u2__abc_52155_new_n6659_; 
wire u2__abc_52155_new_n6660_; 
wire u2__abc_52155_new_n6661_; 
wire u2__abc_52155_new_n6662_; 
wire u2__abc_52155_new_n6663_; 
wire u2__abc_52155_new_n6664_; 
wire u2__abc_52155_new_n6665_; 
wire u2__abc_52155_new_n6666_; 
wire u2__abc_52155_new_n6667_; 
wire u2__abc_52155_new_n6668_; 
wire u2__abc_52155_new_n6669_; 
wire u2__abc_52155_new_n6670_; 
wire u2__abc_52155_new_n6671_; 
wire u2__abc_52155_new_n6672_; 
wire u2__abc_52155_new_n6673_; 
wire u2__abc_52155_new_n6674_; 
wire u2__abc_52155_new_n6675_; 
wire u2__abc_52155_new_n6676_; 
wire u2__abc_52155_new_n6677_; 
wire u2__abc_52155_new_n6678_; 
wire u2__abc_52155_new_n6679_; 
wire u2__abc_52155_new_n6680_; 
wire u2__abc_52155_new_n6681_; 
wire u2__abc_52155_new_n6682_; 
wire u2__abc_52155_new_n6683_; 
wire u2__abc_52155_new_n6684_; 
wire u2__abc_52155_new_n6685_; 
wire u2__abc_52155_new_n6686_; 
wire u2__abc_52155_new_n6687_; 
wire u2__abc_52155_new_n6688_; 
wire u2__abc_52155_new_n6689_; 
wire u2__abc_52155_new_n6690_; 
wire u2__abc_52155_new_n6691_; 
wire u2__abc_52155_new_n6692_; 
wire u2__abc_52155_new_n6693_; 
wire u2__abc_52155_new_n6694_; 
wire u2__abc_52155_new_n6695_; 
wire u2__abc_52155_new_n6696_; 
wire u2__abc_52155_new_n6697_; 
wire u2__abc_52155_new_n6698_; 
wire u2__abc_52155_new_n6699_; 
wire u2__abc_52155_new_n6700_; 
wire u2__abc_52155_new_n6701_; 
wire u2__abc_52155_new_n6702_; 
wire u2__abc_52155_new_n6703_; 
wire u2__abc_52155_new_n6704_; 
wire u2__abc_52155_new_n6705_; 
wire u2__abc_52155_new_n6706_; 
wire u2__abc_52155_new_n6707_; 
wire u2__abc_52155_new_n6708_; 
wire u2__abc_52155_new_n6709_; 
wire u2__abc_52155_new_n6710_; 
wire u2__abc_52155_new_n6711_; 
wire u2__abc_52155_new_n6712_; 
wire u2__abc_52155_new_n6713_; 
wire u2__abc_52155_new_n6714_; 
wire u2__abc_52155_new_n6715_; 
wire u2__abc_52155_new_n6716_; 
wire u2__abc_52155_new_n6717_; 
wire u2__abc_52155_new_n6718_; 
wire u2__abc_52155_new_n6719_; 
wire u2__abc_52155_new_n6720_; 
wire u2__abc_52155_new_n6721_; 
wire u2__abc_52155_new_n6722_; 
wire u2__abc_52155_new_n6723_; 
wire u2__abc_52155_new_n6724_; 
wire u2__abc_52155_new_n6725_; 
wire u2__abc_52155_new_n6726_; 
wire u2__abc_52155_new_n6727_; 
wire u2__abc_52155_new_n6728_; 
wire u2__abc_52155_new_n6729_; 
wire u2__abc_52155_new_n6730_; 
wire u2__abc_52155_new_n6731_; 
wire u2__abc_52155_new_n6732_; 
wire u2__abc_52155_new_n6733_; 
wire u2__abc_52155_new_n6734_; 
wire u2__abc_52155_new_n6735_; 
wire u2__abc_52155_new_n6736_; 
wire u2__abc_52155_new_n6737_; 
wire u2__abc_52155_new_n6738_; 
wire u2__abc_52155_new_n6739_; 
wire u2__abc_52155_new_n6740_; 
wire u2__abc_52155_new_n6741_; 
wire u2__abc_52155_new_n6742_; 
wire u2__abc_52155_new_n6743_; 
wire u2__abc_52155_new_n6744_; 
wire u2__abc_52155_new_n6745_; 
wire u2__abc_52155_new_n6746_; 
wire u2__abc_52155_new_n6747_; 
wire u2__abc_52155_new_n6748_; 
wire u2__abc_52155_new_n6749_; 
wire u2__abc_52155_new_n6750_; 
wire u2__abc_52155_new_n6751_; 
wire u2__abc_52155_new_n6752_; 
wire u2__abc_52155_new_n6753_; 
wire u2__abc_52155_new_n6754_; 
wire u2__abc_52155_new_n6755_; 
wire u2__abc_52155_new_n6756_; 
wire u2__abc_52155_new_n6757_; 
wire u2__abc_52155_new_n6758_; 
wire u2__abc_52155_new_n6759_; 
wire u2__abc_52155_new_n6760_; 
wire u2__abc_52155_new_n6761_; 
wire u2__abc_52155_new_n6762_; 
wire u2__abc_52155_new_n6763_; 
wire u2__abc_52155_new_n6764_; 
wire u2__abc_52155_new_n6765_; 
wire u2__abc_52155_new_n6766_; 
wire u2__abc_52155_new_n6767_; 
wire u2__abc_52155_new_n6768_; 
wire u2__abc_52155_new_n6769_; 
wire u2__abc_52155_new_n6770_; 
wire u2__abc_52155_new_n6771_; 
wire u2__abc_52155_new_n6772_; 
wire u2__abc_52155_new_n6773_; 
wire u2__abc_52155_new_n6774_; 
wire u2__abc_52155_new_n6775_; 
wire u2__abc_52155_new_n6776_; 
wire u2__abc_52155_new_n6777_; 
wire u2__abc_52155_new_n6778_; 
wire u2__abc_52155_new_n6779_; 
wire u2__abc_52155_new_n6780_; 
wire u2__abc_52155_new_n6781_; 
wire u2__abc_52155_new_n6782_; 
wire u2__abc_52155_new_n6783_; 
wire u2__abc_52155_new_n6784_; 
wire u2__abc_52155_new_n6785_; 
wire u2__abc_52155_new_n6786_; 
wire u2__abc_52155_new_n6787_; 
wire u2__abc_52155_new_n6788_; 
wire u2__abc_52155_new_n6789_; 
wire u2__abc_52155_new_n6790_; 
wire u2__abc_52155_new_n6791_; 
wire u2__abc_52155_new_n6792_; 
wire u2__abc_52155_new_n6793_; 
wire u2__abc_52155_new_n6794_; 
wire u2__abc_52155_new_n6795_; 
wire u2__abc_52155_new_n6796_; 
wire u2__abc_52155_new_n6797_; 
wire u2__abc_52155_new_n6798_; 
wire u2__abc_52155_new_n6799_; 
wire u2__abc_52155_new_n6800_; 
wire u2__abc_52155_new_n6801_; 
wire u2__abc_52155_new_n6802_; 
wire u2__abc_52155_new_n6803_; 
wire u2__abc_52155_new_n6804_; 
wire u2__abc_52155_new_n6805_; 
wire u2__abc_52155_new_n6806_; 
wire u2__abc_52155_new_n6807_; 
wire u2__abc_52155_new_n6808_; 
wire u2__abc_52155_new_n6809_; 
wire u2__abc_52155_new_n6810_; 
wire u2__abc_52155_new_n6811_; 
wire u2__abc_52155_new_n6812_; 
wire u2__abc_52155_new_n6813_; 
wire u2__abc_52155_new_n6814_; 
wire u2__abc_52155_new_n6815_; 
wire u2__abc_52155_new_n6816_; 
wire u2__abc_52155_new_n6817_; 
wire u2__abc_52155_new_n6818_; 
wire u2__abc_52155_new_n6819_; 
wire u2__abc_52155_new_n6820_; 
wire u2__abc_52155_new_n6821_; 
wire u2__abc_52155_new_n6822_; 
wire u2__abc_52155_new_n6823_; 
wire u2__abc_52155_new_n6824_; 
wire u2__abc_52155_new_n6825_; 
wire u2__abc_52155_new_n6826_; 
wire u2__abc_52155_new_n6827_; 
wire u2__abc_52155_new_n6828_; 
wire u2__abc_52155_new_n6829_; 
wire u2__abc_52155_new_n6830_; 
wire u2__abc_52155_new_n6831_; 
wire u2__abc_52155_new_n6832_; 
wire u2__abc_52155_new_n6833_; 
wire u2__abc_52155_new_n6834_; 
wire u2__abc_52155_new_n6835_; 
wire u2__abc_52155_new_n6836_; 
wire u2__abc_52155_new_n6837_; 
wire u2__abc_52155_new_n6838_; 
wire u2__abc_52155_new_n6839_; 
wire u2__abc_52155_new_n6840_; 
wire u2__abc_52155_new_n6841_; 
wire u2__abc_52155_new_n6842_; 
wire u2__abc_52155_new_n6843_; 
wire u2__abc_52155_new_n6844_; 
wire u2__abc_52155_new_n6845_; 
wire u2__abc_52155_new_n6846_; 
wire u2__abc_52155_new_n6847_; 
wire u2__abc_52155_new_n6848_; 
wire u2__abc_52155_new_n6849_; 
wire u2__abc_52155_new_n6850_; 
wire u2__abc_52155_new_n6851_; 
wire u2__abc_52155_new_n6852_; 
wire u2__abc_52155_new_n6853_; 
wire u2__abc_52155_new_n6854_; 
wire u2__abc_52155_new_n6855_; 
wire u2__abc_52155_new_n6856_; 
wire u2__abc_52155_new_n6857_; 
wire u2__abc_52155_new_n6858_; 
wire u2__abc_52155_new_n6859_; 
wire u2__abc_52155_new_n6860_; 
wire u2__abc_52155_new_n6861_; 
wire u2__abc_52155_new_n6862_; 
wire u2__abc_52155_new_n6863_; 
wire u2__abc_52155_new_n6864_; 
wire u2__abc_52155_new_n6865_; 
wire u2__abc_52155_new_n6866_; 
wire u2__abc_52155_new_n6867_; 
wire u2__abc_52155_new_n6868_; 
wire u2__abc_52155_new_n6869_; 
wire u2__abc_52155_new_n6870_; 
wire u2__abc_52155_new_n6871_; 
wire u2__abc_52155_new_n6872_; 
wire u2__abc_52155_new_n6873_; 
wire u2__abc_52155_new_n6874_; 
wire u2__abc_52155_new_n6875_; 
wire u2__abc_52155_new_n6876_; 
wire u2__abc_52155_new_n6877_; 
wire u2__abc_52155_new_n6878_; 
wire u2__abc_52155_new_n6879_; 
wire u2__abc_52155_new_n6880_; 
wire u2__abc_52155_new_n6881_; 
wire u2__abc_52155_new_n6882_; 
wire u2__abc_52155_new_n6883_; 
wire u2__abc_52155_new_n6884_; 
wire u2__abc_52155_new_n6885_; 
wire u2__abc_52155_new_n6886_; 
wire u2__abc_52155_new_n6887_; 
wire u2__abc_52155_new_n6888_; 
wire u2__abc_52155_new_n6889_; 
wire u2__abc_52155_new_n6890_; 
wire u2__abc_52155_new_n6891_; 
wire u2__abc_52155_new_n6892_; 
wire u2__abc_52155_new_n6893_; 
wire u2__abc_52155_new_n6894_; 
wire u2__abc_52155_new_n6895_; 
wire u2__abc_52155_new_n6896_; 
wire u2__abc_52155_new_n6897_; 
wire u2__abc_52155_new_n6898_; 
wire u2__abc_52155_new_n6899_; 
wire u2__abc_52155_new_n6900_; 
wire u2__abc_52155_new_n6901_; 
wire u2__abc_52155_new_n6902_; 
wire u2__abc_52155_new_n6903_; 
wire u2__abc_52155_new_n6904_; 
wire u2__abc_52155_new_n6905_; 
wire u2__abc_52155_new_n6906_; 
wire u2__abc_52155_new_n6907_; 
wire u2__abc_52155_new_n6908_; 
wire u2__abc_52155_new_n6909_; 
wire u2__abc_52155_new_n6910_; 
wire u2__abc_52155_new_n6911_; 
wire u2__abc_52155_new_n6912_; 
wire u2__abc_52155_new_n6913_; 
wire u2__abc_52155_new_n6914_; 
wire u2__abc_52155_new_n6915_; 
wire u2__abc_52155_new_n6916_; 
wire u2__abc_52155_new_n6917_; 
wire u2__abc_52155_new_n6918_; 
wire u2__abc_52155_new_n6919_; 
wire u2__abc_52155_new_n6920_; 
wire u2__abc_52155_new_n6921_; 
wire u2__abc_52155_new_n6922_; 
wire u2__abc_52155_new_n6923_; 
wire u2__abc_52155_new_n6924_; 
wire u2__abc_52155_new_n6925_; 
wire u2__abc_52155_new_n6926_; 
wire u2__abc_52155_new_n6927_; 
wire u2__abc_52155_new_n6928_; 
wire u2__abc_52155_new_n6929_; 
wire u2__abc_52155_new_n6930_; 
wire u2__abc_52155_new_n6931_; 
wire u2__abc_52155_new_n6932_; 
wire u2__abc_52155_new_n6933_; 
wire u2__abc_52155_new_n6934_; 
wire u2__abc_52155_new_n6935_; 
wire u2__abc_52155_new_n6936_; 
wire u2__abc_52155_new_n6937_; 
wire u2__abc_52155_new_n6938_; 
wire u2__abc_52155_new_n6939_; 
wire u2__abc_52155_new_n6940_; 
wire u2__abc_52155_new_n6941_; 
wire u2__abc_52155_new_n6942_; 
wire u2__abc_52155_new_n6943_; 
wire u2__abc_52155_new_n6944_; 
wire u2__abc_52155_new_n6945_; 
wire u2__abc_52155_new_n6946_; 
wire u2__abc_52155_new_n6947_; 
wire u2__abc_52155_new_n6948_; 
wire u2__abc_52155_new_n6949_; 
wire u2__abc_52155_new_n6950_; 
wire u2__abc_52155_new_n6951_; 
wire u2__abc_52155_new_n6952_; 
wire u2__abc_52155_new_n6953_; 
wire u2__abc_52155_new_n6954_; 
wire u2__abc_52155_new_n6955_; 
wire u2__abc_52155_new_n6956_; 
wire u2__abc_52155_new_n6957_; 
wire u2__abc_52155_new_n6958_; 
wire u2__abc_52155_new_n6959_; 
wire u2__abc_52155_new_n6960_; 
wire u2__abc_52155_new_n6961_; 
wire u2__abc_52155_new_n6962_; 
wire u2__abc_52155_new_n6963_; 
wire u2__abc_52155_new_n6964_; 
wire u2__abc_52155_new_n6965_; 
wire u2__abc_52155_new_n6966_; 
wire u2__abc_52155_new_n6967_; 
wire u2__abc_52155_new_n6968_; 
wire u2__abc_52155_new_n6969_; 
wire u2__abc_52155_new_n6970_; 
wire u2__abc_52155_new_n6971_; 
wire u2__abc_52155_new_n6972_; 
wire u2__abc_52155_new_n6973_; 
wire u2__abc_52155_new_n6974_; 
wire u2__abc_52155_new_n6975_; 
wire u2__abc_52155_new_n6976_; 
wire u2__abc_52155_new_n6977_; 
wire u2__abc_52155_new_n6978_; 
wire u2__abc_52155_new_n6979_; 
wire u2__abc_52155_new_n6980_; 
wire u2__abc_52155_new_n6981_; 
wire u2__abc_52155_new_n6982_; 
wire u2__abc_52155_new_n6983_; 
wire u2__abc_52155_new_n6984_; 
wire u2__abc_52155_new_n6985_; 
wire u2__abc_52155_new_n6986_; 
wire u2__abc_52155_new_n6987_; 
wire u2__abc_52155_new_n6988_; 
wire u2__abc_52155_new_n6989_; 
wire u2__abc_52155_new_n6990_; 
wire u2__abc_52155_new_n6991_; 
wire u2__abc_52155_new_n6992_; 
wire u2__abc_52155_new_n6993_; 
wire u2__abc_52155_new_n6994_; 
wire u2__abc_52155_new_n6995_; 
wire u2__abc_52155_new_n6996_; 
wire u2__abc_52155_new_n6997_; 
wire u2__abc_52155_new_n6998_; 
wire u2__abc_52155_new_n6999_; 
wire u2__abc_52155_new_n7000_; 
wire u2__abc_52155_new_n7001_; 
wire u2__abc_52155_new_n7002_; 
wire u2__abc_52155_new_n7003_; 
wire u2__abc_52155_new_n7004_; 
wire u2__abc_52155_new_n7005_; 
wire u2__abc_52155_new_n7006_; 
wire u2__abc_52155_new_n7007_; 
wire u2__abc_52155_new_n7008_; 
wire u2__abc_52155_new_n7009_; 
wire u2__abc_52155_new_n7010_; 
wire u2__abc_52155_new_n7011_; 
wire u2__abc_52155_new_n7012_; 
wire u2__abc_52155_new_n7013_; 
wire u2__abc_52155_new_n7014_; 
wire u2__abc_52155_new_n7015_; 
wire u2__abc_52155_new_n7016_; 
wire u2__abc_52155_new_n7017_; 
wire u2__abc_52155_new_n7018_; 
wire u2__abc_52155_new_n7019_; 
wire u2__abc_52155_new_n7020_; 
wire u2__abc_52155_new_n7021_; 
wire u2__abc_52155_new_n7022_; 
wire u2__abc_52155_new_n7023_; 
wire u2__abc_52155_new_n7024_; 
wire u2__abc_52155_new_n7025_; 
wire u2__abc_52155_new_n7026_; 
wire u2__abc_52155_new_n7027_; 
wire u2__abc_52155_new_n7028_; 
wire u2__abc_52155_new_n7029_; 
wire u2__abc_52155_new_n7030_; 
wire u2__abc_52155_new_n7031_; 
wire u2__abc_52155_new_n7032_; 
wire u2__abc_52155_new_n7033_; 
wire u2__abc_52155_new_n7034_; 
wire u2__abc_52155_new_n7035_; 
wire u2__abc_52155_new_n7036_; 
wire u2__abc_52155_new_n7037_; 
wire u2__abc_52155_new_n7038_; 
wire u2__abc_52155_new_n7039_; 
wire u2__abc_52155_new_n7040_; 
wire u2__abc_52155_new_n7041_; 
wire u2__abc_52155_new_n7042_; 
wire u2__abc_52155_new_n7043_; 
wire u2__abc_52155_new_n7044_; 
wire u2__abc_52155_new_n7045_; 
wire u2__abc_52155_new_n7046_; 
wire u2__abc_52155_new_n7047_; 
wire u2__abc_52155_new_n7048_; 
wire u2__abc_52155_new_n7049_; 
wire u2__abc_52155_new_n7050_; 
wire u2__abc_52155_new_n7051_; 
wire u2__abc_52155_new_n7052_; 
wire u2__abc_52155_new_n7053_; 
wire u2__abc_52155_new_n7054_; 
wire u2__abc_52155_new_n7055_; 
wire u2__abc_52155_new_n7056_; 
wire u2__abc_52155_new_n7057_; 
wire u2__abc_52155_new_n7058_; 
wire u2__abc_52155_new_n7059_; 
wire u2__abc_52155_new_n7060_; 
wire u2__abc_52155_new_n7061_; 
wire u2__abc_52155_new_n7062_; 
wire u2__abc_52155_new_n7063_; 
wire u2__abc_52155_new_n7064_; 
wire u2__abc_52155_new_n7065_; 
wire u2__abc_52155_new_n7066_; 
wire u2__abc_52155_new_n7067_; 
wire u2__abc_52155_new_n7068_; 
wire u2__abc_52155_new_n7069_; 
wire u2__abc_52155_new_n7070_; 
wire u2__abc_52155_new_n7071_; 
wire u2__abc_52155_new_n7072_; 
wire u2__abc_52155_new_n7073_; 
wire u2__abc_52155_new_n7074_; 
wire u2__abc_52155_new_n7075_; 
wire u2__abc_52155_new_n7076_; 
wire u2__abc_52155_new_n7077_; 
wire u2__abc_52155_new_n7078_; 
wire u2__abc_52155_new_n7079_; 
wire u2__abc_52155_new_n7080_; 
wire u2__abc_52155_new_n7081_; 
wire u2__abc_52155_new_n7082_; 
wire u2__abc_52155_new_n7083_; 
wire u2__abc_52155_new_n7084_; 
wire u2__abc_52155_new_n7085_; 
wire u2__abc_52155_new_n7086_; 
wire u2__abc_52155_new_n7087_; 
wire u2__abc_52155_new_n7088_; 
wire u2__abc_52155_new_n7089_; 
wire u2__abc_52155_new_n7090_; 
wire u2__abc_52155_new_n7091_; 
wire u2__abc_52155_new_n7092_; 
wire u2__abc_52155_new_n7093_; 
wire u2__abc_52155_new_n7094_; 
wire u2__abc_52155_new_n7095_; 
wire u2__abc_52155_new_n7096_; 
wire u2__abc_52155_new_n7097_; 
wire u2__abc_52155_new_n7098_; 
wire u2__abc_52155_new_n7099_; 
wire u2__abc_52155_new_n7100_; 
wire u2__abc_52155_new_n7101_; 
wire u2__abc_52155_new_n7102_; 
wire u2__abc_52155_new_n7103_; 
wire u2__abc_52155_new_n7104_; 
wire u2__abc_52155_new_n7105_; 
wire u2__abc_52155_new_n7106_; 
wire u2__abc_52155_new_n7107_; 
wire u2__abc_52155_new_n7108_; 
wire u2__abc_52155_new_n7109_; 
wire u2__abc_52155_new_n7110_; 
wire u2__abc_52155_new_n7111_; 
wire u2__abc_52155_new_n7112_; 
wire u2__abc_52155_new_n7113_; 
wire u2__abc_52155_new_n7114_; 
wire u2__abc_52155_new_n7115_; 
wire u2__abc_52155_new_n7116_; 
wire u2__abc_52155_new_n7117_; 
wire u2__abc_52155_new_n7118_; 
wire u2__abc_52155_new_n7119_; 
wire u2__abc_52155_new_n7120_; 
wire u2__abc_52155_new_n7121_; 
wire u2__abc_52155_new_n7122_; 
wire u2__abc_52155_new_n7123_; 
wire u2__abc_52155_new_n7124_; 
wire u2__abc_52155_new_n7125_; 
wire u2__abc_52155_new_n7126_; 
wire u2__abc_52155_new_n7127_; 
wire u2__abc_52155_new_n7128_; 
wire u2__abc_52155_new_n7129_; 
wire u2__abc_52155_new_n7130_; 
wire u2__abc_52155_new_n7131_; 
wire u2__abc_52155_new_n7132_; 
wire u2__abc_52155_new_n7133_; 
wire u2__abc_52155_new_n7134_; 
wire u2__abc_52155_new_n7135_; 
wire u2__abc_52155_new_n7136_; 
wire u2__abc_52155_new_n7137_; 
wire u2__abc_52155_new_n7138_; 
wire u2__abc_52155_new_n7139_; 
wire u2__abc_52155_new_n7140_; 
wire u2__abc_52155_new_n7141_; 
wire u2__abc_52155_new_n7142_; 
wire u2__abc_52155_new_n7143_; 
wire u2__abc_52155_new_n7144_; 
wire u2__abc_52155_new_n7145_; 
wire u2__abc_52155_new_n7146_; 
wire u2__abc_52155_new_n7147_; 
wire u2__abc_52155_new_n7148_; 
wire u2__abc_52155_new_n7149_; 
wire u2__abc_52155_new_n7150_; 
wire u2__abc_52155_new_n7151_; 
wire u2__abc_52155_new_n7152_; 
wire u2__abc_52155_new_n7153_; 
wire u2__abc_52155_new_n7154_; 
wire u2__abc_52155_new_n7155_; 
wire u2__abc_52155_new_n7156_; 
wire u2__abc_52155_new_n7157_; 
wire u2__abc_52155_new_n7158_; 
wire u2__abc_52155_new_n7159_; 
wire u2__abc_52155_new_n7160_; 
wire u2__abc_52155_new_n7161_; 
wire u2__abc_52155_new_n7162_; 
wire u2__abc_52155_new_n7163_; 
wire u2__abc_52155_new_n7164_; 
wire u2__abc_52155_new_n7165_; 
wire u2__abc_52155_new_n7166_; 
wire u2__abc_52155_new_n7167_; 
wire u2__abc_52155_new_n7168_; 
wire u2__abc_52155_new_n7169_; 
wire u2__abc_52155_new_n7170_; 
wire u2__abc_52155_new_n7171_; 
wire u2__abc_52155_new_n7172_; 
wire u2__abc_52155_new_n7173_; 
wire u2__abc_52155_new_n7174_; 
wire u2__abc_52155_new_n7175_; 
wire u2__abc_52155_new_n7176_; 
wire u2__abc_52155_new_n7177_; 
wire u2__abc_52155_new_n7178_; 
wire u2__abc_52155_new_n7179_; 
wire u2__abc_52155_new_n7180_; 
wire u2__abc_52155_new_n7181_; 
wire u2__abc_52155_new_n7182_; 
wire u2__abc_52155_new_n7183_; 
wire u2__abc_52155_new_n7184_; 
wire u2__abc_52155_new_n7185_; 
wire u2__abc_52155_new_n7186_; 
wire u2__abc_52155_new_n7187_; 
wire u2__abc_52155_new_n7188_; 
wire u2__abc_52155_new_n7189_; 
wire u2__abc_52155_new_n7190_; 
wire u2__abc_52155_new_n7191_; 
wire u2__abc_52155_new_n7192_; 
wire u2__abc_52155_new_n7193_; 
wire u2__abc_52155_new_n7194_; 
wire u2__abc_52155_new_n7195_; 
wire u2__abc_52155_new_n7196_; 
wire u2__abc_52155_new_n7197_; 
wire u2__abc_52155_new_n7198_; 
wire u2__abc_52155_new_n7199_; 
wire u2__abc_52155_new_n7200_; 
wire u2__abc_52155_new_n7201_; 
wire u2__abc_52155_new_n7202_; 
wire u2__abc_52155_new_n7203_; 
wire u2__abc_52155_new_n7204_; 
wire u2__abc_52155_new_n7205_; 
wire u2__abc_52155_new_n7206_; 
wire u2__abc_52155_new_n7207_; 
wire u2__abc_52155_new_n7208_; 
wire u2__abc_52155_new_n7209_; 
wire u2__abc_52155_new_n7210_; 
wire u2__abc_52155_new_n7211_; 
wire u2__abc_52155_new_n7212_; 
wire u2__abc_52155_new_n7213_; 
wire u2__abc_52155_new_n7214_; 
wire u2__abc_52155_new_n7215_; 
wire u2__abc_52155_new_n7216_; 
wire u2__abc_52155_new_n7217_; 
wire u2__abc_52155_new_n7218_; 
wire u2__abc_52155_new_n7219_; 
wire u2__abc_52155_new_n7220_; 
wire u2__abc_52155_new_n7221_; 
wire u2__abc_52155_new_n7222_; 
wire u2__abc_52155_new_n7223_; 
wire u2__abc_52155_new_n7224_; 
wire u2__abc_52155_new_n7225_; 
wire u2__abc_52155_new_n7226_; 
wire u2__abc_52155_new_n7227_; 
wire u2__abc_52155_new_n7228_; 
wire u2__abc_52155_new_n7229_; 
wire u2__abc_52155_new_n7230_; 
wire u2__abc_52155_new_n7231_; 
wire u2__abc_52155_new_n7232_; 
wire u2__abc_52155_new_n7233_; 
wire u2__abc_52155_new_n7234_; 
wire u2__abc_52155_new_n7235_; 
wire u2__abc_52155_new_n7236_; 
wire u2__abc_52155_new_n7237_; 
wire u2__abc_52155_new_n7238_; 
wire u2__abc_52155_new_n7239_; 
wire u2__abc_52155_new_n7240_; 
wire u2__abc_52155_new_n7241_; 
wire u2__abc_52155_new_n7242_; 
wire u2__abc_52155_new_n7243_; 
wire u2__abc_52155_new_n7244_; 
wire u2__abc_52155_new_n7245_; 
wire u2__abc_52155_new_n7246_; 
wire u2__abc_52155_new_n7247_; 
wire u2__abc_52155_new_n7248_; 
wire u2__abc_52155_new_n7249_; 
wire u2__abc_52155_new_n7250_; 
wire u2__abc_52155_new_n7251_; 
wire u2__abc_52155_new_n7252_; 
wire u2__abc_52155_new_n7253_; 
wire u2__abc_52155_new_n7254_; 
wire u2__abc_52155_new_n7255_; 
wire u2__abc_52155_new_n7256_; 
wire u2__abc_52155_new_n7257_; 
wire u2__abc_52155_new_n7258_; 
wire u2__abc_52155_new_n7259_; 
wire u2__abc_52155_new_n7260_; 
wire u2__abc_52155_new_n7261_; 
wire u2__abc_52155_new_n7262_; 
wire u2__abc_52155_new_n7263_; 
wire u2__abc_52155_new_n7264_; 
wire u2__abc_52155_new_n7265_; 
wire u2__abc_52155_new_n7266_; 
wire u2__abc_52155_new_n7267_; 
wire u2__abc_52155_new_n7268_; 
wire u2__abc_52155_new_n7269_; 
wire u2__abc_52155_new_n7270_; 
wire u2__abc_52155_new_n7271_; 
wire u2__abc_52155_new_n7272_; 
wire u2__abc_52155_new_n7273_; 
wire u2__abc_52155_new_n7274_; 
wire u2__abc_52155_new_n7275_; 
wire u2__abc_52155_new_n7276_; 
wire u2__abc_52155_new_n7277_; 
wire u2__abc_52155_new_n7278_; 
wire u2__abc_52155_new_n7279_; 
wire u2__abc_52155_new_n7280_; 
wire u2__abc_52155_new_n7281_; 
wire u2__abc_52155_new_n7282_; 
wire u2__abc_52155_new_n7283_; 
wire u2__abc_52155_new_n7284_; 
wire u2__abc_52155_new_n7285_; 
wire u2__abc_52155_new_n7286_; 
wire u2__abc_52155_new_n7287_; 
wire u2__abc_52155_new_n7288_; 
wire u2__abc_52155_new_n7289_; 
wire u2__abc_52155_new_n7290_; 
wire u2__abc_52155_new_n7291_; 
wire u2__abc_52155_new_n7292_; 
wire u2__abc_52155_new_n7293_; 
wire u2__abc_52155_new_n7294_; 
wire u2__abc_52155_new_n7295_; 
wire u2__abc_52155_new_n7296_; 
wire u2__abc_52155_new_n7297_; 
wire u2__abc_52155_new_n7298_; 
wire u2__abc_52155_new_n7299_; 
wire u2__abc_52155_new_n7300_; 
wire u2__abc_52155_new_n7301_; 
wire u2__abc_52155_new_n7302_; 
wire u2__abc_52155_new_n7303_; 
wire u2__abc_52155_new_n7304_; 
wire u2__abc_52155_new_n7305_; 
wire u2__abc_52155_new_n7306_; 
wire u2__abc_52155_new_n7307_; 
wire u2__abc_52155_new_n7308_; 
wire u2__abc_52155_new_n7309_; 
wire u2__abc_52155_new_n7310_; 
wire u2__abc_52155_new_n7311_; 
wire u2__abc_52155_new_n7312_; 
wire u2__abc_52155_new_n7313_; 
wire u2__abc_52155_new_n7314_; 
wire u2__abc_52155_new_n7315_; 
wire u2__abc_52155_new_n7316_; 
wire u2__abc_52155_new_n7317_; 
wire u2__abc_52155_new_n7318_; 
wire u2__abc_52155_new_n7319_; 
wire u2__abc_52155_new_n7320_; 
wire u2__abc_52155_new_n7321_; 
wire u2__abc_52155_new_n7322_; 
wire u2__abc_52155_new_n7323_; 
wire u2__abc_52155_new_n7324_; 
wire u2__abc_52155_new_n7325_; 
wire u2__abc_52155_new_n7326_; 
wire u2__abc_52155_new_n7327_; 
wire u2__abc_52155_new_n7328_; 
wire u2__abc_52155_new_n7329_; 
wire u2__abc_52155_new_n7330_; 
wire u2__abc_52155_new_n7331_; 
wire u2__abc_52155_new_n7332_; 
wire u2__abc_52155_new_n7333_; 
wire u2__abc_52155_new_n7334_; 
wire u2__abc_52155_new_n7335_; 
wire u2__abc_52155_new_n7336_; 
wire u2__abc_52155_new_n7337_; 
wire u2__abc_52155_new_n7338_; 
wire u2__abc_52155_new_n7339_; 
wire u2__abc_52155_new_n7340_; 
wire u2__abc_52155_new_n7341_; 
wire u2__abc_52155_new_n7342_; 
wire u2__abc_52155_new_n7343_; 
wire u2__abc_52155_new_n7344_; 
wire u2__abc_52155_new_n7345_; 
wire u2__abc_52155_new_n7346_; 
wire u2__abc_52155_new_n7347_; 
wire u2__abc_52155_new_n7348_; 
wire u2__abc_52155_new_n7349_; 
wire u2__abc_52155_new_n7350_; 
wire u2__abc_52155_new_n7351_; 
wire u2__abc_52155_new_n7352_; 
wire u2__abc_52155_new_n7353_; 
wire u2__abc_52155_new_n7354_; 
wire u2__abc_52155_new_n7355_; 
wire u2__abc_52155_new_n7356_; 
wire u2__abc_52155_new_n7357_; 
wire u2__abc_52155_new_n7358_; 
wire u2__abc_52155_new_n7359_; 
wire u2__abc_52155_new_n7360_; 
wire u2__abc_52155_new_n7361_; 
wire u2__abc_52155_new_n7362_; 
wire u2__abc_52155_new_n7363_; 
wire u2__abc_52155_new_n7364_; 
wire u2__abc_52155_new_n7365_; 
wire u2__abc_52155_new_n7366_; 
wire u2__abc_52155_new_n7367_; 
wire u2__abc_52155_new_n7368_; 
wire u2__abc_52155_new_n7369_; 
wire u2__abc_52155_new_n7370_; 
wire u2__abc_52155_new_n7371_; 
wire u2__abc_52155_new_n7372_; 
wire u2__abc_52155_new_n7373_; 
wire u2__abc_52155_new_n7374_; 
wire u2__abc_52155_new_n7375_; 
wire u2__abc_52155_new_n7376_; 
wire u2__abc_52155_new_n7377_; 
wire u2__abc_52155_new_n7378_; 
wire u2__abc_52155_new_n7379_; 
wire u2__abc_52155_new_n7380_; 
wire u2__abc_52155_new_n7381_; 
wire u2__abc_52155_new_n7382_; 
wire u2__abc_52155_new_n7383_; 
wire u2__abc_52155_new_n7384_; 
wire u2__abc_52155_new_n7385_; 
wire u2__abc_52155_new_n7386_; 
wire u2__abc_52155_new_n7387_; 
wire u2__abc_52155_new_n7388_; 
wire u2__abc_52155_new_n7389_; 
wire u2__abc_52155_new_n7390_; 
wire u2__abc_52155_new_n7391_; 
wire u2__abc_52155_new_n7392_; 
wire u2__abc_52155_new_n7393_; 
wire u2__abc_52155_new_n7394_; 
wire u2__abc_52155_new_n7395_; 
wire u2__abc_52155_new_n7396_; 
wire u2__abc_52155_new_n7397_; 
wire u2__abc_52155_new_n7398_; 
wire u2__abc_52155_new_n7399_; 
wire u2__abc_52155_new_n7400_; 
wire u2__abc_52155_new_n7401_; 
wire u2__abc_52155_new_n7402_; 
wire u2__abc_52155_new_n7403_; 
wire u2__abc_52155_new_n7404_; 
wire u2__abc_52155_new_n7405_; 
wire u2__abc_52155_new_n7406_; 
wire u2__abc_52155_new_n7407_; 
wire u2__abc_52155_new_n7408_; 
wire u2__abc_52155_new_n7409_; 
wire u2__abc_52155_new_n7410_; 
wire u2__abc_52155_new_n7411_; 
wire u2__abc_52155_new_n7412_; 
wire u2__abc_52155_new_n7413_; 
wire u2__abc_52155_new_n7414_; 
wire u2__abc_52155_new_n7415_; 
wire u2__abc_52155_new_n7416_; 
wire u2__abc_52155_new_n7417_; 
wire u2__abc_52155_new_n7418_; 
wire u2__abc_52155_new_n7419_; 
wire u2__abc_52155_new_n7420_; 
wire u2__abc_52155_new_n7421_; 
wire u2__abc_52155_new_n7422_; 
wire u2__abc_52155_new_n7423_; 
wire u2__abc_52155_new_n7424_; 
wire u2__abc_52155_new_n7425_; 
wire u2__abc_52155_new_n7426_; 
wire u2__abc_52155_new_n7427_; 
wire u2__abc_52155_new_n7428_; 
wire u2__abc_52155_new_n7429_; 
wire u2__abc_52155_new_n7430_; 
wire u2__abc_52155_new_n7431_; 
wire u2__abc_52155_new_n7432_; 
wire u2__abc_52155_new_n7433_; 
wire u2__abc_52155_new_n7434_; 
wire u2__abc_52155_new_n7435_; 
wire u2__abc_52155_new_n7436_; 
wire u2__abc_52155_new_n7437_; 
wire u2__abc_52155_new_n7438_; 
wire u2__abc_52155_new_n7439_; 
wire u2__abc_52155_new_n7440_; 
wire u2__abc_52155_new_n7441_; 
wire u2__abc_52155_new_n7442_; 
wire u2__abc_52155_new_n7443_; 
wire u2__abc_52155_new_n7444_; 
wire u2__abc_52155_new_n7445_; 
wire u2__abc_52155_new_n7446_; 
wire u2__abc_52155_new_n7447_; 
wire u2__abc_52155_new_n7448_; 
wire u2__abc_52155_new_n7449_; 
wire u2__abc_52155_new_n7450_; 
wire u2__abc_52155_new_n7451_; 
wire u2__abc_52155_new_n7452_; 
wire u2__abc_52155_new_n7453_; 
wire u2__abc_52155_new_n7454_; 
wire u2__abc_52155_new_n7455_; 
wire u2__abc_52155_new_n7456_; 
wire u2__abc_52155_new_n7457_; 
wire u2__abc_52155_new_n7458_; 
wire u2__abc_52155_new_n7459_; 
wire u2__abc_52155_new_n7460_; 
wire u2__abc_52155_new_n7461_; 
wire u2__abc_52155_new_n7462_; 
wire u2__abc_52155_new_n7463_; 
wire u2__abc_52155_new_n7464_; 
wire u2__abc_52155_new_n7465_; 
wire u2__abc_52155_new_n7466_; 
wire u2__abc_52155_new_n7467_; 
wire u2__abc_52155_new_n7468_; 
wire u2__abc_52155_new_n7469_; 
wire u2__abc_52155_new_n7470_; 
wire u2__abc_52155_new_n7471_; 
wire u2__abc_52155_new_n7472_; 
wire u2__abc_52155_new_n7473_; 
wire u2__abc_52155_new_n7474_; 
wire u2__abc_52155_new_n7475_; 
wire u2__abc_52155_new_n7476_; 
wire u2__abc_52155_new_n7477_; 
wire u2__abc_52155_new_n7478_; 
wire u2__abc_52155_new_n7479_; 
wire u2__abc_52155_new_n7480_; 
wire u2__abc_52155_new_n7481_; 
wire u2__abc_52155_new_n7482_; 
wire u2__abc_52155_new_n7483_; 
wire u2__abc_52155_new_n7484_; 
wire u2__abc_52155_new_n7485_; 
wire u2__abc_52155_new_n7486_; 
wire u2__abc_52155_new_n7487_; 
wire u2__abc_52155_new_n7488_; 
wire u2__abc_52155_new_n7489_; 
wire u2__abc_52155_new_n7490_; 
wire u2__abc_52155_new_n7491_; 
wire u2__abc_52155_new_n7492_; 
wire u2__abc_52155_new_n7493_; 
wire u2__abc_52155_new_n7494_; 
wire u2__abc_52155_new_n7495_; 
wire u2__abc_52155_new_n7496_; 
wire u2__abc_52155_new_n7497_; 
wire u2__abc_52155_new_n7498_; 
wire u2__abc_52155_new_n7499_; 
wire u2__abc_52155_new_n7500_; 
wire u2__abc_52155_new_n7501_; 
wire u2__abc_52155_new_n7502_; 
wire u2__abc_52155_new_n7503_; 
wire u2__abc_52155_new_n7504_; 
wire u2__abc_52155_new_n7505_; 
wire u2__abc_52155_new_n7506_; 
wire u2__abc_52155_new_n7507_; 
wire u2__abc_52155_new_n7508_; 
wire u2__abc_52155_new_n7509_; 
wire u2__abc_52155_new_n7510_; 
wire u2__abc_52155_new_n7511_; 
wire u2__abc_52155_new_n7512_; 
wire u2__abc_52155_new_n7513_; 
wire u2__abc_52155_new_n7514_; 
wire u2__abc_52155_new_n7515_; 
wire u2__abc_52155_new_n7516_; 
wire u2__abc_52155_new_n7517_; 
wire u2__abc_52155_new_n7518_; 
wire u2__abc_52155_new_n7519_; 
wire u2__abc_52155_new_n7520_; 
wire u2__abc_52155_new_n7521_; 
wire u2__abc_52155_new_n7522_; 
wire u2__abc_52155_new_n7523_; 
wire u2__abc_52155_new_n7524_; 
wire u2__abc_52155_new_n7525_; 
wire u2__abc_52155_new_n7526_; 
wire u2__abc_52155_new_n7527_; 
wire u2__abc_52155_new_n7528_; 
wire u2__abc_52155_new_n7529_; 
wire u2__abc_52155_new_n7530_; 
wire u2__abc_52155_new_n7531_; 
wire u2__abc_52155_new_n7532_; 
wire u2__abc_52155_new_n7533_; 
wire u2__abc_52155_new_n7534_; 
wire u2__abc_52155_new_n7535_; 
wire u2__abc_52155_new_n7536_; 
wire u2__abc_52155_new_n7537_; 
wire u2__abc_52155_new_n7538_; 
wire u2__abc_52155_new_n7539_; 
wire u2__abc_52155_new_n7540_; 
wire u2__abc_52155_new_n7541_; 
wire u2__abc_52155_new_n7542_; 
wire u2__abc_52155_new_n7543_; 
wire u2__abc_52155_new_n7544_; 
wire u2__abc_52155_new_n7545_; 
wire u2__abc_52155_new_n7546_; 
wire u2__abc_52155_new_n7547_; 
wire u2__abc_52155_new_n7548_; 
wire u2__abc_52155_new_n7549_; 
wire u2__abc_52155_new_n7550_; 
wire u2__abc_52155_new_n7551_; 
wire u2__abc_52155_new_n7552_; 
wire u2__abc_52155_new_n7553_; 
wire u2__abc_52155_new_n7554_; 
wire u2__abc_52155_new_n7555_; 
wire u2__abc_52155_new_n7556_; 
wire u2__abc_52155_new_n7557_; 
wire u2__abc_52155_new_n7558_; 
wire u2__abc_52155_new_n7559_; 
wire u2__abc_52155_new_n7560_; 
wire u2__abc_52155_new_n7561_; 
wire u2__abc_52155_new_n7562_; 
wire u2__abc_52155_new_n7563_; 
wire u2__abc_52155_new_n7564_; 
wire u2__abc_52155_new_n7565_; 
wire u2__abc_52155_new_n7566_; 
wire u2__abc_52155_new_n7567_; 
wire u2__abc_52155_new_n7568_; 
wire u2__abc_52155_new_n7569_; 
wire u2__abc_52155_new_n7570_; 
wire u2__abc_52155_new_n7571_; 
wire u2__abc_52155_new_n7572_; 
wire u2__abc_52155_new_n7573_; 
wire u2__abc_52155_new_n7574_; 
wire u2__abc_52155_new_n7575_; 
wire u2__abc_52155_new_n7576_; 
wire u2__abc_52155_new_n7577_; 
wire u2__abc_52155_new_n7578_; 
wire u2__abc_52155_new_n7579_; 
wire u2__abc_52155_new_n7580_; 
wire u2__abc_52155_new_n7581_; 
wire u2__abc_52155_new_n7582_; 
wire u2__abc_52155_new_n7583_; 
wire u2__abc_52155_new_n7584_; 
wire u2__abc_52155_new_n7585_; 
wire u2__abc_52155_new_n7586_; 
wire u2__abc_52155_new_n7587_; 
wire u2__abc_52155_new_n7588_; 
wire u2__abc_52155_new_n7589_; 
wire u2__abc_52155_new_n7590_; 
wire u2__abc_52155_new_n7591_; 
wire u2__abc_52155_new_n7592_; 
wire u2__abc_52155_new_n7593_; 
wire u2__abc_52155_new_n7594_; 
wire u2__abc_52155_new_n7595_; 
wire u2__abc_52155_new_n7596_; 
wire u2__abc_52155_new_n7597_; 
wire u2__abc_52155_new_n7598_; 
wire u2__abc_52155_new_n7599_; 
wire u2__abc_52155_new_n7600_; 
wire u2__abc_52155_new_n7601_; 
wire u2__abc_52155_new_n7602_; 
wire u2__abc_52155_new_n7603_; 
wire u2__abc_52155_new_n7604_; 
wire u2__abc_52155_new_n7605_; 
wire u2__abc_52155_new_n7606_; 
wire u2__abc_52155_new_n7607_; 
wire u2__abc_52155_new_n7608_; 
wire u2__abc_52155_new_n7609_; 
wire u2__abc_52155_new_n7610_; 
wire u2__abc_52155_new_n7611_; 
wire u2__abc_52155_new_n7612_; 
wire u2__abc_52155_new_n7613_; 
wire u2__abc_52155_new_n7614_; 
wire u2__abc_52155_new_n7615_; 
wire u2__abc_52155_new_n7616_; 
wire u2__abc_52155_new_n7617_; 
wire u2__abc_52155_new_n7618_; 
wire u2__abc_52155_new_n7619_; 
wire u2__abc_52155_new_n7620_; 
wire u2__abc_52155_new_n7621_; 
wire u2__abc_52155_new_n7622_; 
wire u2__abc_52155_new_n7623_; 
wire u2__abc_52155_new_n7624_; 
wire u2__abc_52155_new_n7625_; 
wire u2__abc_52155_new_n7626_; 
wire u2__abc_52155_new_n7627_; 
wire u2__abc_52155_new_n7628_; 
wire u2__abc_52155_new_n7629_; 
wire u2__abc_52155_new_n7630_; 
wire u2__abc_52155_new_n7631_; 
wire u2__abc_52155_new_n7632_; 
wire u2__abc_52155_new_n7633_; 
wire u2__abc_52155_new_n7635_; 
wire u2__abc_52155_new_n7636_; 
wire u2__abc_52155_new_n7637_; 
wire u2__abc_52155_new_n7638_; 
wire u2__abc_52155_new_n7639_; 
wire u2__abc_52155_new_n7640_; 
wire u2__abc_52155_new_n7641_; 
wire u2__abc_52155_new_n7642_; 
wire u2__abc_52155_new_n7643_; 
wire u2__abc_52155_new_n7644_; 
wire u2__abc_52155_new_n7645_; 
wire u2__abc_52155_new_n7646_; 
wire u2__abc_52155_new_n7647_; 
wire u2__abc_52155_new_n7649_; 
wire u2__abc_52155_new_n7650_; 
wire u2__abc_52155_new_n7651_; 
wire u2__abc_52155_new_n7652_; 
wire u2__abc_52155_new_n7653_; 
wire u2__abc_52155_new_n7654_; 
wire u2__abc_52155_new_n7655_; 
wire u2__abc_52155_new_n7656_; 
wire u2__abc_52155_new_n7657_; 
wire u2__abc_52155_new_n7658_; 
wire u2__abc_52155_new_n7659_; 
wire u2__abc_52155_new_n7660_; 
wire u2__abc_52155_new_n7661_; 
wire u2__abc_52155_new_n7662_; 
wire u2__abc_52155_new_n7663_; 
wire u2__abc_52155_new_n7664_; 
wire u2__abc_52155_new_n7665_; 
wire u2__abc_52155_new_n7667_; 
wire u2__abc_52155_new_n7668_; 
wire u2__abc_52155_new_n7669_; 
wire u2__abc_52155_new_n7670_; 
wire u2__abc_52155_new_n7671_; 
wire u2__abc_52155_new_n7672_; 
wire u2__abc_52155_new_n7673_; 
wire u2__abc_52155_new_n7674_; 
wire u2__abc_52155_new_n7675_; 
wire u2__abc_52155_new_n7676_; 
wire u2__abc_52155_new_n7677_; 
wire u2__abc_52155_new_n7678_; 
wire u2__abc_52155_new_n7679_; 
wire u2__abc_52155_new_n7680_; 
wire u2__abc_52155_new_n7681_; 
wire u2__abc_52155_new_n7682_; 
wire u2__abc_52155_new_n7683_; 
wire u2__abc_52155_new_n7684_; 
wire u2__abc_52155_new_n7686_; 
wire u2__abc_52155_new_n7687_; 
wire u2__abc_52155_new_n7688_; 
wire u2__abc_52155_new_n7689_; 
wire u2__abc_52155_new_n7690_; 
wire u2__abc_52155_new_n7691_; 
wire u2__abc_52155_new_n7692_; 
wire u2__abc_52155_new_n7693_; 
wire u2__abc_52155_new_n7694_; 
wire u2__abc_52155_new_n7695_; 
wire u2__abc_52155_new_n7696_; 
wire u2__abc_52155_new_n7697_; 
wire u2__abc_52155_new_n7698_; 
wire u2__abc_52155_new_n7699_; 
wire u2__abc_52155_new_n7700_; 
wire u2__abc_52155_new_n7701_; 
wire u2__abc_52155_new_n7703_; 
wire u2__abc_52155_new_n7704_; 
wire u2__abc_52155_new_n7705_; 
wire u2__abc_52155_new_n7706_; 
wire u2__abc_52155_new_n7707_; 
wire u2__abc_52155_new_n7708_; 
wire u2__abc_52155_new_n7709_; 
wire u2__abc_52155_new_n7710_; 
wire u2__abc_52155_new_n7711_; 
wire u2__abc_52155_new_n7712_; 
wire u2__abc_52155_new_n7713_; 
wire u2__abc_52155_new_n7714_; 
wire u2__abc_52155_new_n7715_; 
wire u2__abc_52155_new_n7716_; 
wire u2__abc_52155_new_n7717_; 
wire u2__abc_52155_new_n7718_; 
wire u2__abc_52155_new_n7719_; 
wire u2__abc_52155_new_n7721_; 
wire u2__abc_52155_new_n7722_; 
wire u2__abc_52155_new_n7723_; 
wire u2__abc_52155_new_n7724_; 
wire u2__abc_52155_new_n7725_; 
wire u2__abc_52155_new_n7726_; 
wire u2__abc_52155_new_n7727_; 
wire u2__abc_52155_new_n7728_; 
wire u2__abc_52155_new_n7729_; 
wire u2__abc_52155_new_n7730_; 
wire u2__abc_52155_new_n7731_; 
wire u2__abc_52155_new_n7732_; 
wire u2__abc_52155_new_n7733_; 
wire u2__abc_52155_new_n7734_; 
wire u2__abc_52155_new_n7735_; 
wire u2__abc_52155_new_n7736_; 
wire u2__abc_52155_new_n7737_; 
wire u2__abc_52155_new_n7738_; 
wire u2__abc_52155_new_n7739_; 
wire u2__abc_52155_new_n7741_; 
wire u2__abc_52155_new_n7742_; 
wire u2__abc_52155_new_n7743_; 
wire u2__abc_52155_new_n7744_; 
wire u2__abc_52155_new_n7745_; 
wire u2__abc_52155_new_n7746_; 
wire u2__abc_52155_new_n7747_; 
wire u2__abc_52155_new_n7748_; 
wire u2__abc_52155_new_n7749_; 
wire u2__abc_52155_new_n7750_; 
wire u2__abc_52155_new_n7751_; 
wire u2__abc_52155_new_n7752_; 
wire u2__abc_52155_new_n7753_; 
wire u2__abc_52155_new_n7754_; 
wire u2__abc_52155_new_n7755_; 
wire u2__abc_52155_new_n7756_; 
wire u2__abc_52155_new_n7757_; 
wire u2__abc_52155_new_n7758_; 
wire u2__abc_52155_new_n7760_; 
wire u2__abc_52155_new_n7761_; 
wire u2__abc_52155_new_n7762_; 
wire u2__abc_52155_new_n7763_; 
wire u2__abc_52155_new_n7764_; 
wire u2__abc_52155_new_n7765_; 
wire u2__abc_52155_new_n7766_; 
wire u2__abc_52155_new_n7767_; 
wire u2__abc_52155_new_n7768_; 
wire u2__abc_52155_new_n7769_; 
wire u2__abc_52155_new_n7770_; 
wire u2__abc_52155_new_n7771_; 
wire u2__abc_52155_new_n7772_; 
wire u2__abc_52155_new_n7773_; 
wire u2__abc_52155_new_n7774_; 
wire u2__abc_52155_new_n7775_; 
wire u2__abc_52155_new_n7776_; 
wire u2__abc_52155_new_n7777_; 
wire u2__abc_52155_new_n7778_; 
wire u2__abc_52155_new_n7779_; 
wire u2__abc_52155_new_n7780_; 
wire u2__abc_52155_new_n7782_; 
wire u2__abc_52155_new_n7783_; 
wire u2__abc_52155_new_n7784_; 
wire u2__abc_52155_new_n7785_; 
wire u2__abc_52155_new_n7786_; 
wire u2__abc_52155_new_n7787_; 
wire u2__abc_52155_new_n7788_; 
wire u2__abc_52155_new_n7789_; 
wire u2__abc_52155_new_n7790_; 
wire u2__abc_52155_new_n7791_; 
wire u2__abc_52155_new_n7792_; 
wire u2__abc_52155_new_n7793_; 
wire u2__abc_52155_new_n7794_; 
wire u2__abc_52155_new_n7795_; 
wire u2__abc_52155_new_n7796_; 
wire u2__abc_52155_new_n7797_; 
wire u2__abc_52155_new_n7799_; 
wire u2__abc_52155_new_n7800_; 
wire u2__abc_52155_new_n7801_; 
wire u2__abc_52155_new_n7802_; 
wire u2__abc_52155_new_n7803_; 
wire u2__abc_52155_new_n7804_; 
wire u2__abc_52155_new_n7805_; 
wire u2__abc_52155_new_n7806_; 
wire u2__abc_52155_new_n7807_; 
wire u2__abc_52155_new_n7808_; 
wire u2__abc_52155_new_n7809_; 
wire u2__abc_52155_new_n7810_; 
wire u2__abc_52155_new_n7811_; 
wire u2__abc_52155_new_n7812_; 
wire u2__abc_52155_new_n7813_; 
wire u2__abc_52155_new_n7814_; 
wire u2__abc_52155_new_n7815_; 
wire u2__abc_52155_new_n7816_; 
wire u2__abc_52155_new_n7817_; 
wire u2__abc_52155_new_n7819_; 
wire u2__abc_52155_new_n7820_; 
wire u2__abc_52155_new_n7821_; 
wire u2__abc_52155_new_n7822_; 
wire u2__abc_52155_new_n7823_; 
wire u2__abc_52155_new_n7824_; 
wire u2__abc_52155_new_n7825_; 
wire u2__abc_52155_new_n7826_; 
wire u2__abc_52155_new_n7827_; 
wire u2__abc_52155_new_n7828_; 
wire u2__abc_52155_new_n7829_; 
wire u2__abc_52155_new_n7830_; 
wire u2__abc_52155_new_n7831_; 
wire u2__abc_52155_new_n7832_; 
wire u2__abc_52155_new_n7833_; 
wire u2__abc_52155_new_n7834_; 
wire u2__abc_52155_new_n7835_; 
wire u2__abc_52155_new_n7837_; 
wire u2__abc_52155_new_n7838_; 
wire u2__abc_52155_new_n7839_; 
wire u2__abc_52155_new_n7840_; 
wire u2__abc_52155_new_n7841_; 
wire u2__abc_52155_new_n7842_; 
wire u2__abc_52155_new_n7843_; 
wire u2__abc_52155_new_n7844_; 
wire u2__abc_52155_new_n7845_; 
wire u2__abc_52155_new_n7846_; 
wire u2__abc_52155_new_n7847_; 
wire u2__abc_52155_new_n7848_; 
wire u2__abc_52155_new_n7849_; 
wire u2__abc_52155_new_n7850_; 
wire u2__abc_52155_new_n7851_; 
wire u2__abc_52155_new_n7852_; 
wire u2__abc_52155_new_n7853_; 
wire u2__abc_52155_new_n7854_; 
wire u2__abc_52155_new_n7856_; 
wire u2__abc_52155_new_n7857_; 
wire u2__abc_52155_new_n7858_; 
wire u2__abc_52155_new_n7859_; 
wire u2__abc_52155_new_n7860_; 
wire u2__abc_52155_new_n7861_; 
wire u2__abc_52155_new_n7862_; 
wire u2__abc_52155_new_n7863_; 
wire u2__abc_52155_new_n7864_; 
wire u2__abc_52155_new_n7865_; 
wire u2__abc_52155_new_n7866_; 
wire u2__abc_52155_new_n7867_; 
wire u2__abc_52155_new_n7868_; 
wire u2__abc_52155_new_n7869_; 
wire u2__abc_52155_new_n7870_; 
wire u2__abc_52155_new_n7871_; 
wire u2__abc_52155_new_n7872_; 
wire u2__abc_52155_new_n7874_; 
wire u2__abc_52155_new_n7875_; 
wire u2__abc_52155_new_n7876_; 
wire u2__abc_52155_new_n7877_; 
wire u2__abc_52155_new_n7878_; 
wire u2__abc_52155_new_n7879_; 
wire u2__abc_52155_new_n7880_; 
wire u2__abc_52155_new_n7881_; 
wire u2__abc_52155_new_n7882_; 
wire u2__abc_52155_new_n7883_; 
wire u2__abc_52155_new_n7884_; 
wire u2__abc_52155_new_n7885_; 
wire u2__abc_52155_new_n7886_; 
wire u2__abc_52155_new_n7887_; 
wire u2__abc_52155_new_n7888_; 
wire u2__abc_52155_new_n7889_; 
wire u2__abc_52155_new_n7890_; 
wire u2__abc_52155_new_n7891_; 
wire u2__abc_52155_new_n7892_; 
wire u2__abc_52155_new_n7893_; 
wire u2__abc_52155_new_n7894_; 
wire u2__abc_52155_new_n7895_; 
wire u2__abc_52155_new_n7897_; 
wire u2__abc_52155_new_n7898_; 
wire u2__abc_52155_new_n7899_; 
wire u2__abc_52155_new_n7900_; 
wire u2__abc_52155_new_n7901_; 
wire u2__abc_52155_new_n7902_; 
wire u2__abc_52155_new_n7903_; 
wire u2__abc_52155_new_n7904_; 
wire u2__abc_52155_new_n7905_; 
wire u2__abc_52155_new_n7906_; 
wire u2__abc_52155_new_n7907_; 
wire u2__abc_52155_new_n7908_; 
wire u2__abc_52155_new_n7909_; 
wire u2__abc_52155_new_n7910_; 
wire u2__abc_52155_new_n7911_; 
wire u2__abc_52155_new_n7912_; 
wire u2__abc_52155_new_n7914_; 
wire u2__abc_52155_new_n7915_; 
wire u2__abc_52155_new_n7916_; 
wire u2__abc_52155_new_n7917_; 
wire u2__abc_52155_new_n7918_; 
wire u2__abc_52155_new_n7919_; 
wire u2__abc_52155_new_n7920_; 
wire u2__abc_52155_new_n7921_; 
wire u2__abc_52155_new_n7922_; 
wire u2__abc_52155_new_n7923_; 
wire u2__abc_52155_new_n7924_; 
wire u2__abc_52155_new_n7925_; 
wire u2__abc_52155_new_n7926_; 
wire u2__abc_52155_new_n7927_; 
wire u2__abc_52155_new_n7928_; 
wire u2__abc_52155_new_n7929_; 
wire u2__abc_52155_new_n7930_; 
wire u2__abc_52155_new_n7931_; 
wire u2__abc_52155_new_n7932_; 
wire u2__abc_52155_new_n7933_; 
wire u2__abc_52155_new_n7934_; 
wire u2__abc_52155_new_n7935_; 
wire u2__abc_52155_new_n7936_; 
wire u2__abc_52155_new_n7937_; 
wire u2__abc_52155_new_n7938_; 
wire u2__abc_52155_new_n7939_; 
wire u2__abc_52155_new_n7940_; 
wire u2__abc_52155_new_n7941_; 
wire u2__abc_52155_new_n7942_; 
wire u2__abc_52155_new_n7944_; 
wire u2__abc_52155_new_n7945_; 
wire u2__abc_52155_new_n7946_; 
wire u2__abc_52155_new_n7947_; 
wire u2__abc_52155_new_n7948_; 
wire u2__abc_52155_new_n7949_; 
wire u2__abc_52155_new_n7950_; 
wire u2__abc_52155_new_n7951_; 
wire u2__abc_52155_new_n7952_; 
wire u2__abc_52155_new_n7953_; 
wire u2__abc_52155_new_n7954_; 
wire u2__abc_52155_new_n7955_; 
wire u2__abc_52155_new_n7956_; 
wire u2__abc_52155_new_n7957_; 
wire u2__abc_52155_new_n7958_; 
wire u2__abc_52155_new_n7959_; 
wire u2__abc_52155_new_n7961_; 
wire u2__abc_52155_new_n7962_; 
wire u2__abc_52155_new_n7963_; 
wire u2__abc_52155_new_n7964_; 
wire u2__abc_52155_new_n7965_; 
wire u2__abc_52155_new_n7966_; 
wire u2__abc_52155_new_n7967_; 
wire u2__abc_52155_new_n7968_; 
wire u2__abc_52155_new_n7969_; 
wire u2__abc_52155_new_n7970_; 
wire u2__abc_52155_new_n7971_; 
wire u2__abc_52155_new_n7972_; 
wire u2__abc_52155_new_n7973_; 
wire u2__abc_52155_new_n7974_; 
wire u2__abc_52155_new_n7975_; 
wire u2__abc_52155_new_n7976_; 
wire u2__abc_52155_new_n7977_; 
wire u2__abc_52155_new_n7979_; 
wire u2__abc_52155_new_n7980_; 
wire u2__abc_52155_new_n7981_; 
wire u2__abc_52155_new_n7982_; 
wire u2__abc_52155_new_n7983_; 
wire u2__abc_52155_new_n7984_; 
wire u2__abc_52155_new_n7985_; 
wire u2__abc_52155_new_n7986_; 
wire u2__abc_52155_new_n7987_; 
wire u2__abc_52155_new_n7988_; 
wire u2__abc_52155_new_n7989_; 
wire u2__abc_52155_new_n7990_; 
wire u2__abc_52155_new_n7991_; 
wire u2__abc_52155_new_n7992_; 
wire u2__abc_52155_new_n7993_; 
wire u2__abc_52155_new_n7994_; 
wire u2__abc_52155_new_n7995_; 
wire u2__abc_52155_new_n7997_; 
wire u2__abc_52155_new_n7998_; 
wire u2__abc_52155_new_n7999_; 
wire u2__abc_52155_new_n8000_; 
wire u2__abc_52155_new_n8001_; 
wire u2__abc_52155_new_n8002_; 
wire u2__abc_52155_new_n8003_; 
wire u2__abc_52155_new_n8004_; 
wire u2__abc_52155_new_n8005_; 
wire u2__abc_52155_new_n8006_; 
wire u2__abc_52155_new_n8007_; 
wire u2__abc_52155_new_n8008_; 
wire u2__abc_52155_new_n8009_; 
wire u2__abc_52155_new_n8010_; 
wire u2__abc_52155_new_n8011_; 
wire u2__abc_52155_new_n8012_; 
wire u2__abc_52155_new_n8013_; 
wire u2__abc_52155_new_n8014_; 
wire u2__abc_52155_new_n8015_; 
wire u2__abc_52155_new_n8016_; 
wire u2__abc_52155_new_n8017_; 
wire u2__abc_52155_new_n8018_; 
wire u2__abc_52155_new_n8019_; 
wire u2__abc_52155_new_n8020_; 
wire u2__abc_52155_new_n8021_; 
wire u2__abc_52155_new_n8023_; 
wire u2__abc_52155_new_n8024_; 
wire u2__abc_52155_new_n8025_; 
wire u2__abc_52155_new_n8026_; 
wire u2__abc_52155_new_n8027_; 
wire u2__abc_52155_new_n8028_; 
wire u2__abc_52155_new_n8029_; 
wire u2__abc_52155_new_n8030_; 
wire u2__abc_52155_new_n8031_; 
wire u2__abc_52155_new_n8032_; 
wire u2__abc_52155_new_n8033_; 
wire u2__abc_52155_new_n8034_; 
wire u2__abc_52155_new_n8035_; 
wire u2__abc_52155_new_n8036_; 
wire u2__abc_52155_new_n8037_; 
wire u2__abc_52155_new_n8038_; 
wire u2__abc_52155_new_n8039_; 
wire u2__abc_52155_new_n8041_; 
wire u2__abc_52155_new_n8042_; 
wire u2__abc_52155_new_n8043_; 
wire u2__abc_52155_new_n8044_; 
wire u2__abc_52155_new_n8045_; 
wire u2__abc_52155_new_n8046_; 
wire u2__abc_52155_new_n8047_; 
wire u2__abc_52155_new_n8048_; 
wire u2__abc_52155_new_n8049_; 
wire u2__abc_52155_new_n8050_; 
wire u2__abc_52155_new_n8051_; 
wire u2__abc_52155_new_n8052_; 
wire u2__abc_52155_new_n8053_; 
wire u2__abc_52155_new_n8054_; 
wire u2__abc_52155_new_n8055_; 
wire u2__abc_52155_new_n8056_; 
wire u2__abc_52155_new_n8057_; 
wire u2__abc_52155_new_n8058_; 
wire u2__abc_52155_new_n8059_; 
wire u2__abc_52155_new_n8060_; 
wire u2__abc_52155_new_n8062_; 
wire u2__abc_52155_new_n8063_; 
wire u2__abc_52155_new_n8064_; 
wire u2__abc_52155_new_n8065_; 
wire u2__abc_52155_new_n8066_; 
wire u2__abc_52155_new_n8067_; 
wire u2__abc_52155_new_n8068_; 
wire u2__abc_52155_new_n8069_; 
wire u2__abc_52155_new_n8070_; 
wire u2__abc_52155_new_n8071_; 
wire u2__abc_52155_new_n8072_; 
wire u2__abc_52155_new_n8073_; 
wire u2__abc_52155_new_n8074_; 
wire u2__abc_52155_new_n8075_; 
wire u2__abc_52155_new_n8076_; 
wire u2__abc_52155_new_n8077_; 
wire u2__abc_52155_new_n8078_; 
wire u2__abc_52155_new_n8080_; 
wire u2__abc_52155_new_n8081_; 
wire u2__abc_52155_new_n8082_; 
wire u2__abc_52155_new_n8083_; 
wire u2__abc_52155_new_n8084_; 
wire u2__abc_52155_new_n8085_; 
wire u2__abc_52155_new_n8086_; 
wire u2__abc_52155_new_n8087_; 
wire u2__abc_52155_new_n8088_; 
wire u2__abc_52155_new_n8089_; 
wire u2__abc_52155_new_n8090_; 
wire u2__abc_52155_new_n8091_; 
wire u2__abc_52155_new_n8092_; 
wire u2__abc_52155_new_n8093_; 
wire u2__abc_52155_new_n8094_; 
wire u2__abc_52155_new_n8095_; 
wire u2__abc_52155_new_n8096_; 
wire u2__abc_52155_new_n8097_; 
wire u2__abc_52155_new_n8098_; 
wire u2__abc_52155_new_n8099_; 
wire u2__abc_52155_new_n8100_; 
wire u2__abc_52155_new_n8101_; 
wire u2__abc_52155_new_n8102_; 
wire u2__abc_52155_new_n8103_; 
wire u2__abc_52155_new_n8104_; 
wire u2__abc_52155_new_n8105_; 
wire u2__abc_52155_new_n8107_; 
wire u2__abc_52155_new_n8108_; 
wire u2__abc_52155_new_n8109_; 
wire u2__abc_52155_new_n8110_; 
wire u2__abc_52155_new_n8111_; 
wire u2__abc_52155_new_n8112_; 
wire u2__abc_52155_new_n8113_; 
wire u2__abc_52155_new_n8114_; 
wire u2__abc_52155_new_n8115_; 
wire u2__abc_52155_new_n8116_; 
wire u2__abc_52155_new_n8117_; 
wire u2__abc_52155_new_n8118_; 
wire u2__abc_52155_new_n8119_; 
wire u2__abc_52155_new_n8120_; 
wire u2__abc_52155_new_n8121_; 
wire u2__abc_52155_new_n8122_; 
wire u2__abc_52155_new_n8124_; 
wire u2__abc_52155_new_n8125_; 
wire u2__abc_52155_new_n8126_; 
wire u2__abc_52155_new_n8127_; 
wire u2__abc_52155_new_n8128_; 
wire u2__abc_52155_new_n8129_; 
wire u2__abc_52155_new_n8130_; 
wire u2__abc_52155_new_n8131_; 
wire u2__abc_52155_new_n8132_; 
wire u2__abc_52155_new_n8133_; 
wire u2__abc_52155_new_n8134_; 
wire u2__abc_52155_new_n8135_; 
wire u2__abc_52155_new_n8136_; 
wire u2__abc_52155_new_n8137_; 
wire u2__abc_52155_new_n8138_; 
wire u2__abc_52155_new_n8139_; 
wire u2__abc_52155_new_n8140_; 
wire u2__abc_52155_new_n8141_; 
wire u2__abc_52155_new_n8142_; 
wire u2__abc_52155_new_n8144_; 
wire u2__abc_52155_new_n8145_; 
wire u2__abc_52155_new_n8146_; 
wire u2__abc_52155_new_n8147_; 
wire u2__abc_52155_new_n8148_; 
wire u2__abc_52155_new_n8149_; 
wire u2__abc_52155_new_n8150_; 
wire u2__abc_52155_new_n8151_; 
wire u2__abc_52155_new_n8152_; 
wire u2__abc_52155_new_n8153_; 
wire u2__abc_52155_new_n8154_; 
wire u2__abc_52155_new_n8155_; 
wire u2__abc_52155_new_n8156_; 
wire u2__abc_52155_new_n8157_; 
wire u2__abc_52155_new_n8158_; 
wire u2__abc_52155_new_n8159_; 
wire u2__abc_52155_new_n8160_; 
wire u2__abc_52155_new_n8162_; 
wire u2__abc_52155_new_n8163_; 
wire u2__abc_52155_new_n8164_; 
wire u2__abc_52155_new_n8165_; 
wire u2__abc_52155_new_n8166_; 
wire u2__abc_52155_new_n8167_; 
wire u2__abc_52155_new_n8168_; 
wire u2__abc_52155_new_n8169_; 
wire u2__abc_52155_new_n8170_; 
wire u2__abc_52155_new_n8171_; 
wire u2__abc_52155_new_n8172_; 
wire u2__abc_52155_new_n8173_; 
wire u2__abc_52155_new_n8174_; 
wire u2__abc_52155_new_n8175_; 
wire u2__abc_52155_new_n8176_; 
wire u2__abc_52155_new_n8177_; 
wire u2__abc_52155_new_n8178_; 
wire u2__abc_52155_new_n8179_; 
wire u2__abc_52155_new_n8180_; 
wire u2__abc_52155_new_n8181_; 
wire u2__abc_52155_new_n8182_; 
wire u2__abc_52155_new_n8183_; 
wire u2__abc_52155_new_n8184_; 
wire u2__abc_52155_new_n8186_; 
wire u2__abc_52155_new_n8187_; 
wire u2__abc_52155_new_n8188_; 
wire u2__abc_52155_new_n8189_; 
wire u2__abc_52155_new_n8190_; 
wire u2__abc_52155_new_n8191_; 
wire u2__abc_52155_new_n8192_; 
wire u2__abc_52155_new_n8193_; 
wire u2__abc_52155_new_n8194_; 
wire u2__abc_52155_new_n8195_; 
wire u2__abc_52155_new_n8196_; 
wire u2__abc_52155_new_n8197_; 
wire u2__abc_52155_new_n8198_; 
wire u2__abc_52155_new_n8199_; 
wire u2__abc_52155_new_n8200_; 
wire u2__abc_52155_new_n8201_; 
wire u2__abc_52155_new_n8203_; 
wire u2__abc_52155_new_n8204_; 
wire u2__abc_52155_new_n8205_; 
wire u2__abc_52155_new_n8206_; 
wire u2__abc_52155_new_n8207_; 
wire u2__abc_52155_new_n8208_; 
wire u2__abc_52155_new_n8209_; 
wire u2__abc_52155_new_n8210_; 
wire u2__abc_52155_new_n8211_; 
wire u2__abc_52155_new_n8212_; 
wire u2__abc_52155_new_n8213_; 
wire u2__abc_52155_new_n8214_; 
wire u2__abc_52155_new_n8215_; 
wire u2__abc_52155_new_n8216_; 
wire u2__abc_52155_new_n8217_; 
wire u2__abc_52155_new_n8218_; 
wire u2__abc_52155_new_n8219_; 
wire u2__abc_52155_new_n8220_; 
wire u2__abc_52155_new_n8221_; 
wire u2__abc_52155_new_n8223_; 
wire u2__abc_52155_new_n8224_; 
wire u2__abc_52155_new_n8225_; 
wire u2__abc_52155_new_n8226_; 
wire u2__abc_52155_new_n8227_; 
wire u2__abc_52155_new_n8228_; 
wire u2__abc_52155_new_n8229_; 
wire u2__abc_52155_new_n8230_; 
wire u2__abc_52155_new_n8231_; 
wire u2__abc_52155_new_n8232_; 
wire u2__abc_52155_new_n8233_; 
wire u2__abc_52155_new_n8234_; 
wire u2__abc_52155_new_n8235_; 
wire u2__abc_52155_new_n8236_; 
wire u2__abc_52155_new_n8237_; 
wire u2__abc_52155_new_n8238_; 
wire u2__abc_52155_new_n8240_; 
wire u2__abc_52155_new_n8241_; 
wire u2__abc_52155_new_n8242_; 
wire u2__abc_52155_new_n8243_; 
wire u2__abc_52155_new_n8244_; 
wire u2__abc_52155_new_n8245_; 
wire u2__abc_52155_new_n8246_; 
wire u2__abc_52155_new_n8247_; 
wire u2__abc_52155_new_n8248_; 
wire u2__abc_52155_new_n8249_; 
wire u2__abc_52155_new_n8250_; 
wire u2__abc_52155_new_n8251_; 
wire u2__abc_52155_new_n8252_; 
wire u2__abc_52155_new_n8253_; 
wire u2__abc_52155_new_n8254_; 
wire u2__abc_52155_new_n8255_; 
wire u2__abc_52155_new_n8256_; 
wire u2__abc_52155_new_n8257_; 
wire u2__abc_52155_new_n8258_; 
wire u2__abc_52155_new_n8259_; 
wire u2__abc_52155_new_n8260_; 
wire u2__abc_52155_new_n8261_; 
wire u2__abc_52155_new_n8263_; 
wire u2__abc_52155_new_n8264_; 
wire u2__abc_52155_new_n8265_; 
wire u2__abc_52155_new_n8266_; 
wire u2__abc_52155_new_n8267_; 
wire u2__abc_52155_new_n8268_; 
wire u2__abc_52155_new_n8269_; 
wire u2__abc_52155_new_n8270_; 
wire u2__abc_52155_new_n8271_; 
wire u2__abc_52155_new_n8272_; 
wire u2__abc_52155_new_n8273_; 
wire u2__abc_52155_new_n8274_; 
wire u2__abc_52155_new_n8275_; 
wire u2__abc_52155_new_n8276_; 
wire u2__abc_52155_new_n8277_; 
wire u2__abc_52155_new_n8278_; 
wire u2__abc_52155_new_n8280_; 
wire u2__abc_52155_new_n8281_; 
wire u2__abc_52155_new_n8282_; 
wire u2__abc_52155_new_n8283_; 
wire u2__abc_52155_new_n8284_; 
wire u2__abc_52155_new_n8285_; 
wire u2__abc_52155_new_n8286_; 
wire u2__abc_52155_new_n8287_; 
wire u2__abc_52155_new_n8288_; 
wire u2__abc_52155_new_n8289_; 
wire u2__abc_52155_new_n8290_; 
wire u2__abc_52155_new_n8291_; 
wire u2__abc_52155_new_n8292_; 
wire u2__abc_52155_new_n8293_; 
wire u2__abc_52155_new_n8294_; 
wire u2__abc_52155_new_n8295_; 
wire u2__abc_52155_new_n8296_; 
wire u2__abc_52155_new_n8298_; 
wire u2__abc_52155_new_n8299_; 
wire u2__abc_52155_new_n8300_; 
wire u2__abc_52155_new_n8301_; 
wire u2__abc_52155_new_n8302_; 
wire u2__abc_52155_new_n8303_; 
wire u2__abc_52155_new_n8304_; 
wire u2__abc_52155_new_n8305_; 
wire u2__abc_52155_new_n8306_; 
wire u2__abc_52155_new_n8307_; 
wire u2__abc_52155_new_n8308_; 
wire u2__abc_52155_new_n8309_; 
wire u2__abc_52155_new_n8310_; 
wire u2__abc_52155_new_n8311_; 
wire u2__abc_52155_new_n8312_; 
wire u2__abc_52155_new_n8313_; 
wire u2__abc_52155_new_n8314_; 
wire u2__abc_52155_new_n8316_; 
wire u2__abc_52155_new_n8317_; 
wire u2__abc_52155_new_n8318_; 
wire u2__abc_52155_new_n8319_; 
wire u2__abc_52155_new_n8320_; 
wire u2__abc_52155_new_n8321_; 
wire u2__abc_52155_new_n8322_; 
wire u2__abc_52155_new_n8323_; 
wire u2__abc_52155_new_n8324_; 
wire u2__abc_52155_new_n8325_; 
wire u2__abc_52155_new_n8326_; 
wire u2__abc_52155_new_n8327_; 
wire u2__abc_52155_new_n8328_; 
wire u2__abc_52155_new_n8329_; 
wire u2__abc_52155_new_n8330_; 
wire u2__abc_52155_new_n8331_; 
wire u2__abc_52155_new_n8332_; 
wire u2__abc_52155_new_n8333_; 
wire u2__abc_52155_new_n8334_; 
wire u2__abc_52155_new_n8335_; 
wire u2__abc_52155_new_n8336_; 
wire u2__abc_52155_new_n8337_; 
wire u2__abc_52155_new_n8338_; 
wire u2__abc_52155_new_n8339_; 
wire u2__abc_52155_new_n8340_; 
wire u2__abc_52155_new_n8342_; 
wire u2__abc_52155_new_n8343_; 
wire u2__abc_52155_new_n8344_; 
wire u2__abc_52155_new_n8345_; 
wire u2__abc_52155_new_n8346_; 
wire u2__abc_52155_new_n8347_; 
wire u2__abc_52155_new_n8348_; 
wire u2__abc_52155_new_n8349_; 
wire u2__abc_52155_new_n8350_; 
wire u2__abc_52155_new_n8351_; 
wire u2__abc_52155_new_n8352_; 
wire u2__abc_52155_new_n8353_; 
wire u2__abc_52155_new_n8354_; 
wire u2__abc_52155_new_n8355_; 
wire u2__abc_52155_new_n8356_; 
wire u2__abc_52155_new_n8357_; 
wire u2__abc_52155_new_n8358_; 
wire u2__abc_52155_new_n8360_; 
wire u2__abc_52155_new_n8361_; 
wire u2__abc_52155_new_n8362_; 
wire u2__abc_52155_new_n8363_; 
wire u2__abc_52155_new_n8364_; 
wire u2__abc_52155_new_n8365_; 
wire u2__abc_52155_new_n8366_; 
wire u2__abc_52155_new_n8367_; 
wire u2__abc_52155_new_n8368_; 
wire u2__abc_52155_new_n8369_; 
wire u2__abc_52155_new_n8370_; 
wire u2__abc_52155_new_n8371_; 
wire u2__abc_52155_new_n8372_; 
wire u2__abc_52155_new_n8373_; 
wire u2__abc_52155_new_n8374_; 
wire u2__abc_52155_new_n8375_; 
wire u2__abc_52155_new_n8376_; 
wire u2__abc_52155_new_n8377_; 
wire u2__abc_52155_new_n8378_; 
wire u2__abc_52155_new_n8379_; 
wire u2__abc_52155_new_n8381_; 
wire u2__abc_52155_new_n8382_; 
wire u2__abc_52155_new_n8383_; 
wire u2__abc_52155_new_n8384_; 
wire u2__abc_52155_new_n8385_; 
wire u2__abc_52155_new_n8386_; 
wire u2__abc_52155_new_n8387_; 
wire u2__abc_52155_new_n8388_; 
wire u2__abc_52155_new_n8389_; 
wire u2__abc_52155_new_n8390_; 
wire u2__abc_52155_new_n8391_; 
wire u2__abc_52155_new_n8392_; 
wire u2__abc_52155_new_n8393_; 
wire u2__abc_52155_new_n8394_; 
wire u2__abc_52155_new_n8395_; 
wire u2__abc_52155_new_n8396_; 
wire u2__abc_52155_new_n8397_; 
wire u2__abc_52155_new_n8399_; 
wire u2__abc_52155_new_n8400_; 
wire u2__abc_52155_new_n8401_; 
wire u2__abc_52155_new_n8402_; 
wire u2__abc_52155_new_n8403_; 
wire u2__abc_52155_new_n8404_; 
wire u2__abc_52155_new_n8405_; 
wire u2__abc_52155_new_n8406_; 
wire u2__abc_52155_new_n8407_; 
wire u2__abc_52155_new_n8408_; 
wire u2__abc_52155_new_n8409_; 
wire u2__abc_52155_new_n8410_; 
wire u2__abc_52155_new_n8411_; 
wire u2__abc_52155_new_n8412_; 
wire u2__abc_52155_new_n8413_; 
wire u2__abc_52155_new_n8414_; 
wire u2__abc_52155_new_n8415_; 
wire u2__abc_52155_new_n8416_; 
wire u2__abc_52155_new_n8417_; 
wire u2__abc_52155_new_n8418_; 
wire u2__abc_52155_new_n8419_; 
wire u2__abc_52155_new_n8420_; 
wire u2__abc_52155_new_n8421_; 
wire u2__abc_52155_new_n8422_; 
wire u2__abc_52155_new_n8423_; 
wire u2__abc_52155_new_n8425_; 
wire u2__abc_52155_new_n8426_; 
wire u2__abc_52155_new_n8427_; 
wire u2__abc_52155_new_n8428_; 
wire u2__abc_52155_new_n8429_; 
wire u2__abc_52155_new_n8430_; 
wire u2__abc_52155_new_n8431_; 
wire u2__abc_52155_new_n8432_; 
wire u2__abc_52155_new_n8433_; 
wire u2__abc_52155_new_n8434_; 
wire u2__abc_52155_new_n8435_; 
wire u2__abc_52155_new_n8436_; 
wire u2__abc_52155_new_n8437_; 
wire u2__abc_52155_new_n8438_; 
wire u2__abc_52155_new_n8439_; 
wire u2__abc_52155_new_n8440_; 
wire u2__abc_52155_new_n8442_; 
wire u2__abc_52155_new_n8443_; 
wire u2__abc_52155_new_n8444_; 
wire u2__abc_52155_new_n8445_; 
wire u2__abc_52155_new_n8446_; 
wire u2__abc_52155_new_n8447_; 
wire u2__abc_52155_new_n8448_; 
wire u2__abc_52155_new_n8449_; 
wire u2__abc_52155_new_n8450_; 
wire u2__abc_52155_new_n8451_; 
wire u2__abc_52155_new_n8452_; 
wire u2__abc_52155_new_n8453_; 
wire u2__abc_52155_new_n8454_; 
wire u2__abc_52155_new_n8455_; 
wire u2__abc_52155_new_n8456_; 
wire u2__abc_52155_new_n8457_; 
wire u2__abc_52155_new_n8458_; 
wire u2__abc_52155_new_n8460_; 
wire u2__abc_52155_new_n8461_; 
wire u2__abc_52155_new_n8462_; 
wire u2__abc_52155_new_n8463_; 
wire u2__abc_52155_new_n8464_; 
wire u2__abc_52155_new_n8465_; 
wire u2__abc_52155_new_n8466_; 
wire u2__abc_52155_new_n8467_; 
wire u2__abc_52155_new_n8468_; 
wire u2__abc_52155_new_n8469_; 
wire u2__abc_52155_new_n8470_; 
wire u2__abc_52155_new_n8471_; 
wire u2__abc_52155_new_n8472_; 
wire u2__abc_52155_new_n8473_; 
wire u2__abc_52155_new_n8474_; 
wire u2__abc_52155_new_n8475_; 
wire u2__abc_52155_new_n8476_; 
wire u2__abc_52155_new_n8478_; 
wire u2__abc_52155_new_n8479_; 
wire u2__abc_52155_new_n8480_; 
wire u2__abc_52155_new_n8481_; 
wire u2__abc_52155_new_n8482_; 
wire u2__abc_52155_new_n8483_; 
wire u2__abc_52155_new_n8484_; 
wire u2__abc_52155_new_n8485_; 
wire u2__abc_52155_new_n8486_; 
wire u2__abc_52155_new_n8487_; 
wire u2__abc_52155_new_n8488_; 
wire u2__abc_52155_new_n8489_; 
wire u2__abc_52155_new_n8490_; 
wire u2__abc_52155_new_n8491_; 
wire u2__abc_52155_new_n8492_; 
wire u2__abc_52155_new_n8493_; 
wire u2__abc_52155_new_n8494_; 
wire u2__abc_52155_new_n8495_; 
wire u2__abc_52155_new_n8496_; 
wire u2__abc_52155_new_n8497_; 
wire u2__abc_52155_new_n8498_; 
wire u2__abc_52155_new_n8499_; 
wire u2__abc_52155_new_n8500_; 
wire u2__abc_52155_new_n8502_; 
wire u2__abc_52155_new_n8503_; 
wire u2__abc_52155_new_n8504_; 
wire u2__abc_52155_new_n8505_; 
wire u2__abc_52155_new_n8506_; 
wire u2__abc_52155_new_n8507_; 
wire u2__abc_52155_new_n8508_; 
wire u2__abc_52155_new_n8509_; 
wire u2__abc_52155_new_n8510_; 
wire u2__abc_52155_new_n8511_; 
wire u2__abc_52155_new_n8512_; 
wire u2__abc_52155_new_n8513_; 
wire u2__abc_52155_new_n8514_; 
wire u2__abc_52155_new_n8515_; 
wire u2__abc_52155_new_n8516_; 
wire u2__abc_52155_new_n8517_; 
wire u2__abc_52155_new_n8519_; 
wire u2__abc_52155_new_n8520_; 
wire u2__abc_52155_new_n8521_; 
wire u2__abc_52155_new_n8522_; 
wire u2__abc_52155_new_n8523_; 
wire u2__abc_52155_new_n8524_; 
wire u2__abc_52155_new_n8525_; 
wire u2__abc_52155_new_n8526_; 
wire u2__abc_52155_new_n8527_; 
wire u2__abc_52155_new_n8528_; 
wire u2__abc_52155_new_n8529_; 
wire u2__abc_52155_new_n8530_; 
wire u2__abc_52155_new_n8531_; 
wire u2__abc_52155_new_n8532_; 
wire u2__abc_52155_new_n8533_; 
wire u2__abc_52155_new_n8534_; 
wire u2__abc_52155_new_n8535_; 
wire u2__abc_52155_new_n8536_; 
wire u2__abc_52155_new_n8538_; 
wire u2__abc_52155_new_n8539_; 
wire u2__abc_52155_new_n8540_; 
wire u2__abc_52155_new_n8541_; 
wire u2__abc_52155_new_n8542_; 
wire u2__abc_52155_new_n8543_; 
wire u2__abc_52155_new_n8544_; 
wire u2__abc_52155_new_n8545_; 
wire u2__abc_52155_new_n8546_; 
wire u2__abc_52155_new_n8547_; 
wire u2__abc_52155_new_n8548_; 
wire u2__abc_52155_new_n8549_; 
wire u2__abc_52155_new_n8550_; 
wire u2__abc_52155_new_n8551_; 
wire u2__abc_52155_new_n8552_; 
wire u2__abc_52155_new_n8553_; 
wire u2__abc_52155_new_n8555_; 
wire u2__abc_52155_new_n8556_; 
wire u2__abc_52155_new_n8557_; 
wire u2__abc_52155_new_n8558_; 
wire u2__abc_52155_new_n8559_; 
wire u2__abc_52155_new_n8560_; 
wire u2__abc_52155_new_n8561_; 
wire u2__abc_52155_new_n8562_; 
wire u2__abc_52155_new_n8563_; 
wire u2__abc_52155_new_n8564_; 
wire u2__abc_52155_new_n8565_; 
wire u2__abc_52155_new_n8566_; 
wire u2__abc_52155_new_n8567_; 
wire u2__abc_52155_new_n8568_; 
wire u2__abc_52155_new_n8569_; 
wire u2__abc_52155_new_n8570_; 
wire u2__abc_52155_new_n8571_; 
wire u2__abc_52155_new_n8572_; 
wire u2__abc_52155_new_n8573_; 
wire u2__abc_52155_new_n8574_; 
wire u2__abc_52155_new_n8575_; 
wire u2__abc_52155_new_n8576_; 
wire u2__abc_52155_new_n8577_; 
wire u2__abc_52155_new_n8578_; 
wire u2__abc_52155_new_n8579_; 
wire u2__abc_52155_new_n8580_; 
wire u2__abc_52155_new_n8582_; 
wire u2__abc_52155_new_n8583_; 
wire u2__abc_52155_new_n8584_; 
wire u2__abc_52155_new_n8585_; 
wire u2__abc_52155_new_n8586_; 
wire u2__abc_52155_new_n8587_; 
wire u2__abc_52155_new_n8588_; 
wire u2__abc_52155_new_n8589_; 
wire u2__abc_52155_new_n8590_; 
wire u2__abc_52155_new_n8591_; 
wire u2__abc_52155_new_n8592_; 
wire u2__abc_52155_new_n8593_; 
wire u2__abc_52155_new_n8594_; 
wire u2__abc_52155_new_n8595_; 
wire u2__abc_52155_new_n8596_; 
wire u2__abc_52155_new_n8597_; 
wire u2__abc_52155_new_n8599_; 
wire u2__abc_52155_new_n8600_; 
wire u2__abc_52155_new_n8601_; 
wire u2__abc_52155_new_n8602_; 
wire u2__abc_52155_new_n8603_; 
wire u2__abc_52155_new_n8604_; 
wire u2__abc_52155_new_n8605_; 
wire u2__abc_52155_new_n8606_; 
wire u2__abc_52155_new_n8607_; 
wire u2__abc_52155_new_n8608_; 
wire u2__abc_52155_new_n8609_; 
wire u2__abc_52155_new_n8610_; 
wire u2__abc_52155_new_n8611_; 
wire u2__abc_52155_new_n8612_; 
wire u2__abc_52155_new_n8613_; 
wire u2__abc_52155_new_n8614_; 
wire u2__abc_52155_new_n8615_; 
wire u2__abc_52155_new_n8616_; 
wire u2__abc_52155_new_n8617_; 
wire u2__abc_52155_new_n8619_; 
wire u2__abc_52155_new_n8620_; 
wire u2__abc_52155_new_n8621_; 
wire u2__abc_52155_new_n8622_; 
wire u2__abc_52155_new_n8623_; 
wire u2__abc_52155_new_n8624_; 
wire u2__abc_52155_new_n8625_; 
wire u2__abc_52155_new_n8626_; 
wire u2__abc_52155_new_n8627_; 
wire u2__abc_52155_new_n8628_; 
wire u2__abc_52155_new_n8629_; 
wire u2__abc_52155_new_n8630_; 
wire u2__abc_52155_new_n8631_; 
wire u2__abc_52155_new_n8632_; 
wire u2__abc_52155_new_n8633_; 
wire u2__abc_52155_new_n8634_; 
wire u2__abc_52155_new_n8635_; 
wire u2__abc_52155_new_n8637_; 
wire u2__abc_52155_new_n8638_; 
wire u2__abc_52155_new_n8639_; 
wire u2__abc_52155_new_n8640_; 
wire u2__abc_52155_new_n8641_; 
wire u2__abc_52155_new_n8642_; 
wire u2__abc_52155_new_n8643_; 
wire u2__abc_52155_new_n8644_; 
wire u2__abc_52155_new_n8645_; 
wire u2__abc_52155_new_n8646_; 
wire u2__abc_52155_new_n8647_; 
wire u2__abc_52155_new_n8648_; 
wire u2__abc_52155_new_n8649_; 
wire u2__abc_52155_new_n8650_; 
wire u2__abc_52155_new_n8651_; 
wire u2__abc_52155_new_n8652_; 
wire u2__abc_52155_new_n8653_; 
wire u2__abc_52155_new_n8654_; 
wire u2__abc_52155_new_n8655_; 
wire u2__abc_52155_new_n8656_; 
wire u2__abc_52155_new_n8657_; 
wire u2__abc_52155_new_n8658_; 
wire u2__abc_52155_new_n8660_; 
wire u2__abc_52155_new_n8661_; 
wire u2__abc_52155_new_n8662_; 
wire u2__abc_52155_new_n8663_; 
wire u2__abc_52155_new_n8664_; 
wire u2__abc_52155_new_n8665_; 
wire u2__abc_52155_new_n8666_; 
wire u2__abc_52155_new_n8667_; 
wire u2__abc_52155_new_n8668_; 
wire u2__abc_52155_new_n8669_; 
wire u2__abc_52155_new_n8670_; 
wire u2__abc_52155_new_n8671_; 
wire u2__abc_52155_new_n8672_; 
wire u2__abc_52155_new_n8673_; 
wire u2__abc_52155_new_n8674_; 
wire u2__abc_52155_new_n8675_; 
wire u2__abc_52155_new_n8677_; 
wire u2__abc_52155_new_n8678_; 
wire u2__abc_52155_new_n8679_; 
wire u2__abc_52155_new_n8680_; 
wire u2__abc_52155_new_n8681_; 
wire u2__abc_52155_new_n8682_; 
wire u2__abc_52155_new_n8683_; 
wire u2__abc_52155_new_n8684_; 
wire u2__abc_52155_new_n8685_; 
wire u2__abc_52155_new_n8686_; 
wire u2__abc_52155_new_n8687_; 
wire u2__abc_52155_new_n8688_; 
wire u2__abc_52155_new_n8689_; 
wire u2__abc_52155_new_n8690_; 
wire u2__abc_52155_new_n8691_; 
wire u2__abc_52155_new_n8692_; 
wire u2__abc_52155_new_n8693_; 
wire u2__abc_52155_new_n8694_; 
wire u2__abc_52155_new_n8696_; 
wire u2__abc_52155_new_n8697_; 
wire u2__abc_52155_new_n8698_; 
wire u2__abc_52155_new_n8699_; 
wire u2__abc_52155_new_n8700_; 
wire u2__abc_52155_new_n8701_; 
wire u2__abc_52155_new_n8702_; 
wire u2__abc_52155_new_n8703_; 
wire u2__abc_52155_new_n8704_; 
wire u2__abc_52155_new_n8705_; 
wire u2__abc_52155_new_n8706_; 
wire u2__abc_52155_new_n8707_; 
wire u2__abc_52155_new_n8708_; 
wire u2__abc_52155_new_n8709_; 
wire u2__abc_52155_new_n8710_; 
wire u2__abc_52155_new_n8711_; 
wire u2__abc_52155_new_n8713_; 
wire u2__abc_52155_new_n8714_; 
wire u2__abc_52155_new_n8715_; 
wire u2__abc_52155_new_n8716_; 
wire u2__abc_52155_new_n8717_; 
wire u2__abc_52155_new_n8718_; 
wire u2__abc_52155_new_n8719_; 
wire u2__abc_52155_new_n8720_; 
wire u2__abc_52155_new_n8721_; 
wire u2__abc_52155_new_n8722_; 
wire u2__abc_52155_new_n8723_; 
wire u2__abc_52155_new_n8724_; 
wire u2__abc_52155_new_n8725_; 
wire u2__abc_52155_new_n8726_; 
wire u2__abc_52155_new_n8727_; 
wire u2__abc_52155_new_n8728_; 
wire u2__abc_52155_new_n8729_; 
wire u2__abc_52155_new_n8730_; 
wire u2__abc_52155_new_n8731_; 
wire u2__abc_52155_new_n8732_; 
wire u2__abc_52155_new_n8733_; 
wire u2__abc_52155_new_n8734_; 
wire u2__abc_52155_new_n8735_; 
wire u2__abc_52155_new_n8736_; 
wire u2__abc_52155_new_n8738_; 
wire u2__abc_52155_new_n8739_; 
wire u2__abc_52155_new_n8740_; 
wire u2__abc_52155_new_n8741_; 
wire u2__abc_52155_new_n8742_; 
wire u2__abc_52155_new_n8743_; 
wire u2__abc_52155_new_n8744_; 
wire u2__abc_52155_new_n8745_; 
wire u2__abc_52155_new_n8746_; 
wire u2__abc_52155_new_n8747_; 
wire u2__abc_52155_new_n8748_; 
wire u2__abc_52155_new_n8749_; 
wire u2__abc_52155_new_n8750_; 
wire u2__abc_52155_new_n8751_; 
wire u2__abc_52155_new_n8752_; 
wire u2__abc_52155_new_n8753_; 
wire u2__abc_52155_new_n8755_; 
wire u2__abc_52155_new_n8756_; 
wire u2__abc_52155_new_n8757_; 
wire u2__abc_52155_new_n8758_; 
wire u2__abc_52155_new_n8759_; 
wire u2__abc_52155_new_n8760_; 
wire u2__abc_52155_new_n8761_; 
wire u2__abc_52155_new_n8762_; 
wire u2__abc_52155_new_n8763_; 
wire u2__abc_52155_new_n8764_; 
wire u2__abc_52155_new_n8765_; 
wire u2__abc_52155_new_n8766_; 
wire u2__abc_52155_new_n8767_; 
wire u2__abc_52155_new_n8768_; 
wire u2__abc_52155_new_n8769_; 
wire u2__abc_52155_new_n8770_; 
wire u2__abc_52155_new_n8771_; 
wire u2__abc_52155_new_n8772_; 
wire u2__abc_52155_new_n8773_; 
wire u2__abc_52155_new_n8775_; 
wire u2__abc_52155_new_n8776_; 
wire u2__abc_52155_new_n8777_; 
wire u2__abc_52155_new_n8778_; 
wire u2__abc_52155_new_n8779_; 
wire u2__abc_52155_new_n8780_; 
wire u2__abc_52155_new_n8781_; 
wire u2__abc_52155_new_n8782_; 
wire u2__abc_52155_new_n8783_; 
wire u2__abc_52155_new_n8784_; 
wire u2__abc_52155_new_n8785_; 
wire u2__abc_52155_new_n8786_; 
wire u2__abc_52155_new_n8787_; 
wire u2__abc_52155_new_n8788_; 
wire u2__abc_52155_new_n8789_; 
wire u2__abc_52155_new_n8790_; 
wire u2__abc_52155_new_n8792_; 
wire u2__abc_52155_new_n8793_; 
wire u2__abc_52155_new_n8794_; 
wire u2__abc_52155_new_n8795_; 
wire u2__abc_52155_new_n8796_; 
wire u2__abc_52155_new_n8797_; 
wire u2__abc_52155_new_n8798_; 
wire u2__abc_52155_new_n8799_; 
wire u2__abc_52155_new_n8800_; 
wire u2__abc_52155_new_n8801_; 
wire u2__abc_52155_new_n8802_; 
wire u2__abc_52155_new_n8803_; 
wire u2__abc_52155_new_n8804_; 
wire u2__abc_52155_new_n8805_; 
wire u2__abc_52155_new_n8806_; 
wire u2__abc_52155_new_n8807_; 
wire u2__abc_52155_new_n8808_; 
wire u2__abc_52155_new_n8809_; 
wire u2__abc_52155_new_n8810_; 
wire u2__abc_52155_new_n8811_; 
wire u2__abc_52155_new_n8813_; 
wire u2__abc_52155_new_n8814_; 
wire u2__abc_52155_new_n8815_; 
wire u2__abc_52155_new_n8816_; 
wire u2__abc_52155_new_n8817_; 
wire u2__abc_52155_new_n8818_; 
wire u2__abc_52155_new_n8819_; 
wire u2__abc_52155_new_n8820_; 
wire u2__abc_52155_new_n8821_; 
wire u2__abc_52155_new_n8822_; 
wire u2__abc_52155_new_n8823_; 
wire u2__abc_52155_new_n8824_; 
wire u2__abc_52155_new_n8825_; 
wire u2__abc_52155_new_n8826_; 
wire u2__abc_52155_new_n8827_; 
wire u2__abc_52155_new_n8828_; 
wire u2__abc_52155_new_n8830_; 
wire u2__abc_52155_new_n8831_; 
wire u2__abc_52155_new_n8832_; 
wire u2__abc_52155_new_n8833_; 
wire u2__abc_52155_new_n8834_; 
wire u2__abc_52155_new_n8835_; 
wire u2__abc_52155_new_n8836_; 
wire u2__abc_52155_new_n8837_; 
wire u2__abc_52155_new_n8838_; 
wire u2__abc_52155_new_n8839_; 
wire u2__abc_52155_new_n8840_; 
wire u2__abc_52155_new_n8841_; 
wire u2__abc_52155_new_n8842_; 
wire u2__abc_52155_new_n8843_; 
wire u2__abc_52155_new_n8844_; 
wire u2__abc_52155_new_n8845_; 
wire u2__abc_52155_new_n8846_; 
wire u2__abc_52155_new_n8848_; 
wire u2__abc_52155_new_n8849_; 
wire u2__abc_52155_new_n8850_; 
wire u2__abc_52155_new_n8851_; 
wire u2__abc_52155_new_n8852_; 
wire u2__abc_52155_new_n8853_; 
wire u2__abc_52155_new_n8854_; 
wire u2__abc_52155_new_n8855_; 
wire u2__abc_52155_new_n8856_; 
wire u2__abc_52155_new_n8857_; 
wire u2__abc_52155_new_n8858_; 
wire u2__abc_52155_new_n8859_; 
wire u2__abc_52155_new_n8860_; 
wire u2__abc_52155_new_n8861_; 
wire u2__abc_52155_new_n8862_; 
wire u2__abc_52155_new_n8863_; 
wire u2__abc_52155_new_n8865_; 
wire u2__abc_52155_new_n8866_; 
wire u2__abc_52155_new_n8867_; 
wire u2__abc_52155_new_n8868_; 
wire u2__abc_52155_new_n8869_; 
wire u2__abc_52155_new_n8870_; 
wire u2__abc_52155_new_n8871_; 
wire u2__abc_52155_new_n8872_; 
wire u2__abc_52155_new_n8873_; 
wire u2__abc_52155_new_n8874_; 
wire u2__abc_52155_new_n8875_; 
wire u2__abc_52155_new_n8876_; 
wire u2__abc_52155_new_n8877_; 
wire u2__abc_52155_new_n8878_; 
wire u2__abc_52155_new_n8879_; 
wire u2__abc_52155_new_n8880_; 
wire u2__abc_52155_new_n8881_; 
wire u2__abc_52155_new_n8882_; 
wire u2__abc_52155_new_n8883_; 
wire u2__abc_52155_new_n8884_; 
wire u2__abc_52155_new_n8885_; 
wire u2__abc_52155_new_n8886_; 
wire u2__abc_52155_new_n8887_; 
wire u2__abc_52155_new_n8888_; 
wire u2__abc_52155_new_n8889_; 
wire u2__abc_52155_new_n8890_; 
wire u2__abc_52155_new_n8892_; 
wire u2__abc_52155_new_n8893_; 
wire u2__abc_52155_new_n8894_; 
wire u2__abc_52155_new_n8895_; 
wire u2__abc_52155_new_n8896_; 
wire u2__abc_52155_new_n8897_; 
wire u2__abc_52155_new_n8898_; 
wire u2__abc_52155_new_n8899_; 
wire u2__abc_52155_new_n8900_; 
wire u2__abc_52155_new_n8901_; 
wire u2__abc_52155_new_n8902_; 
wire u2__abc_52155_new_n8903_; 
wire u2__abc_52155_new_n8904_; 
wire u2__abc_52155_new_n8905_; 
wire u2__abc_52155_new_n8906_; 
wire u2__abc_52155_new_n8907_; 
wire u2__abc_52155_new_n8909_; 
wire u2__abc_52155_new_n8910_; 
wire u2__abc_52155_new_n8911_; 
wire u2__abc_52155_new_n8912_; 
wire u2__abc_52155_new_n8913_; 
wire u2__abc_52155_new_n8914_; 
wire u2__abc_52155_new_n8915_; 
wire u2__abc_52155_new_n8916_; 
wire u2__abc_52155_new_n8917_; 
wire u2__abc_52155_new_n8918_; 
wire u2__abc_52155_new_n8919_; 
wire u2__abc_52155_new_n8920_; 
wire u2__abc_52155_new_n8921_; 
wire u2__abc_52155_new_n8922_; 
wire u2__abc_52155_new_n8923_; 
wire u2__abc_52155_new_n8924_; 
wire u2__abc_52155_new_n8925_; 
wire u2__abc_52155_new_n8926_; 
wire u2__abc_52155_new_n8927_; 
wire u2__abc_52155_new_n8928_; 
wire u2__abc_52155_new_n8930_; 
wire u2__abc_52155_new_n8931_; 
wire u2__abc_52155_new_n8932_; 
wire u2__abc_52155_new_n8933_; 
wire u2__abc_52155_new_n8934_; 
wire u2__abc_52155_new_n8935_; 
wire u2__abc_52155_new_n8936_; 
wire u2__abc_52155_new_n8937_; 
wire u2__abc_52155_new_n8938_; 
wire u2__abc_52155_new_n8939_; 
wire u2__abc_52155_new_n8940_; 
wire u2__abc_52155_new_n8941_; 
wire u2__abc_52155_new_n8942_; 
wire u2__abc_52155_new_n8943_; 
wire u2__abc_52155_new_n8944_; 
wire u2__abc_52155_new_n8945_; 
wire u2__abc_52155_new_n8946_; 
wire u2__abc_52155_new_n8948_; 
wire u2__abc_52155_new_n8949_; 
wire u2__abc_52155_new_n8950_; 
wire u2__abc_52155_new_n8951_; 
wire u2__abc_52155_new_n8952_; 
wire u2__abc_52155_new_n8953_; 
wire u2__abc_52155_new_n8954_; 
wire u2__abc_52155_new_n8955_; 
wire u2__abc_52155_new_n8956_; 
wire u2__abc_52155_new_n8957_; 
wire u2__abc_52155_new_n8958_; 
wire u2__abc_52155_new_n8959_; 
wire u2__abc_52155_new_n8960_; 
wire u2__abc_52155_new_n8961_; 
wire u2__abc_52155_new_n8962_; 
wire u2__abc_52155_new_n8963_; 
wire u2__abc_52155_new_n8964_; 
wire u2__abc_52155_new_n8965_; 
wire u2__abc_52155_new_n8966_; 
wire u2__abc_52155_new_n8967_; 
wire u2__abc_52155_new_n8968_; 
wire u2__abc_52155_new_n8970_; 
wire u2__abc_52155_new_n8971_; 
wire u2__abc_52155_new_n8972_; 
wire u2__abc_52155_new_n8973_; 
wire u2__abc_52155_new_n8974_; 
wire u2__abc_52155_new_n8975_; 
wire u2__abc_52155_new_n8976_; 
wire u2__abc_52155_new_n8977_; 
wire u2__abc_52155_new_n8978_; 
wire u2__abc_52155_new_n8979_; 
wire u2__abc_52155_new_n8980_; 
wire u2__abc_52155_new_n8981_; 
wire u2__abc_52155_new_n8982_; 
wire u2__abc_52155_new_n8983_; 
wire u2__abc_52155_new_n8984_; 
wire u2__abc_52155_new_n8985_; 
wire u2__abc_52155_new_n8986_; 
wire u2__abc_52155_new_n8987_; 
wire u2__abc_52155_new_n8989_; 
wire u2__abc_52155_new_n8990_; 
wire u2__abc_52155_new_n8991_; 
wire u2__abc_52155_new_n8992_; 
wire u2__abc_52155_new_n8993_; 
wire u2__abc_52155_new_n8994_; 
wire u2__abc_52155_new_n8995_; 
wire u2__abc_52155_new_n8996_; 
wire u2__abc_52155_new_n8997_; 
wire u2__abc_52155_new_n8998_; 
wire u2__abc_52155_new_n8999_; 
wire u2__abc_52155_new_n9000_; 
wire u2__abc_52155_new_n9001_; 
wire u2__abc_52155_new_n9002_; 
wire u2__abc_52155_new_n9003_; 
wire u2__abc_52155_new_n9004_; 
wire u2__abc_52155_new_n9006_; 
wire u2__abc_52155_new_n9007_; 
wire u2__abc_52155_new_n9008_; 
wire u2__abc_52155_new_n9009_; 
wire u2__abc_52155_new_n9010_; 
wire u2__abc_52155_new_n9011_; 
wire u2__abc_52155_new_n9012_; 
wire u2__abc_52155_new_n9013_; 
wire u2__abc_52155_new_n9014_; 
wire u2__abc_52155_new_n9015_; 
wire u2__abc_52155_new_n9016_; 
wire u2__abc_52155_new_n9017_; 
wire u2__abc_52155_new_n9018_; 
wire u2__abc_52155_new_n9019_; 
wire u2__abc_52155_new_n9020_; 
wire u2__abc_52155_new_n9021_; 
wire u2__abc_52155_new_n9022_; 
wire u2__abc_52155_new_n9024_; 
wire u2__abc_52155_new_n9025_; 
wire u2__abc_52155_new_n9026_; 
wire u2__abc_52155_new_n9027_; 
wire u2__abc_52155_new_n9028_; 
wire u2__abc_52155_new_n9029_; 
wire u2__abc_52155_new_n9030_; 
wire u2__abc_52155_new_n9031_; 
wire u2__abc_52155_new_n9032_; 
wire u2__abc_52155_new_n9033_; 
wire u2__abc_52155_new_n9034_; 
wire u2__abc_52155_new_n9035_; 
wire u2__abc_52155_new_n9036_; 
wire u2__abc_52155_new_n9037_; 
wire u2__abc_52155_new_n9038_; 
wire u2__abc_52155_new_n9039_; 
wire u2__abc_52155_new_n9040_; 
wire u2__abc_52155_new_n9041_; 
wire u2__abc_52155_new_n9042_; 
wire u2__abc_52155_new_n9043_; 
wire u2__abc_52155_new_n9044_; 
wire u2__abc_52155_new_n9045_; 
wire u2__abc_52155_new_n9046_; 
wire u2__abc_52155_new_n9047_; 
wire u2__abc_52155_new_n9048_; 
wire u2__abc_52155_new_n9049_; 
wire u2__abc_52155_new_n9050_; 
wire u2__abc_52155_new_n9051_; 
wire u2__abc_52155_new_n9053_; 
wire u2__abc_52155_new_n9054_; 
wire u2__abc_52155_new_n9055_; 
wire u2__abc_52155_new_n9056_; 
wire u2__abc_52155_new_n9057_; 
wire u2__abc_52155_new_n9058_; 
wire u2__abc_52155_new_n9059_; 
wire u2__abc_52155_new_n9060_; 
wire u2__abc_52155_new_n9061_; 
wire u2__abc_52155_new_n9062_; 
wire u2__abc_52155_new_n9063_; 
wire u2__abc_52155_new_n9064_; 
wire u2__abc_52155_new_n9065_; 
wire u2__abc_52155_new_n9066_; 
wire u2__abc_52155_new_n9067_; 
wire u2__abc_52155_new_n9068_; 
wire u2__abc_52155_new_n9070_; 
wire u2__abc_52155_new_n9071_; 
wire u2__abc_52155_new_n9072_; 
wire u2__abc_52155_new_n9073_; 
wire u2__abc_52155_new_n9074_; 
wire u2__abc_52155_new_n9075_; 
wire u2__abc_52155_new_n9076_; 
wire u2__abc_52155_new_n9077_; 
wire u2__abc_52155_new_n9078_; 
wire u2__abc_52155_new_n9079_; 
wire u2__abc_52155_new_n9080_; 
wire u2__abc_52155_new_n9081_; 
wire u2__abc_52155_new_n9082_; 
wire u2__abc_52155_new_n9083_; 
wire u2__abc_52155_new_n9084_; 
wire u2__abc_52155_new_n9085_; 
wire u2__abc_52155_new_n9086_; 
wire u2__abc_52155_new_n9087_; 
wire u2__abc_52155_new_n9088_; 
wire u2__abc_52155_new_n9089_; 
wire u2__abc_52155_new_n9091_; 
wire u2__abc_52155_new_n9092_; 
wire u2__abc_52155_new_n9093_; 
wire u2__abc_52155_new_n9094_; 
wire u2__abc_52155_new_n9095_; 
wire u2__abc_52155_new_n9096_; 
wire u2__abc_52155_new_n9097_; 
wire u2__abc_52155_new_n9098_; 
wire u2__abc_52155_new_n9099_; 
wire u2__abc_52155_new_n9100_; 
wire u2__abc_52155_new_n9101_; 
wire u2__abc_52155_new_n9102_; 
wire u2__abc_52155_new_n9103_; 
wire u2__abc_52155_new_n9104_; 
wire u2__abc_52155_new_n9105_; 
wire u2__abc_52155_new_n9106_; 
wire u2__abc_52155_new_n9107_; 
wire u2__abc_52155_new_n9109_; 
wire u2__abc_52155_new_n9110_; 
wire u2__abc_52155_new_n9111_; 
wire u2__abc_52155_new_n9112_; 
wire u2__abc_52155_new_n9113_; 
wire u2__abc_52155_new_n9114_; 
wire u2__abc_52155_new_n9115_; 
wire u2__abc_52155_new_n9116_; 
wire u2__abc_52155_new_n9117_; 
wire u2__abc_52155_new_n9118_; 
wire u2__abc_52155_new_n9119_; 
wire u2__abc_52155_new_n9120_; 
wire u2__abc_52155_new_n9121_; 
wire u2__abc_52155_new_n9122_; 
wire u2__abc_52155_new_n9123_; 
wire u2__abc_52155_new_n9124_; 
wire u2__abc_52155_new_n9125_; 
wire u2__abc_52155_new_n9126_; 
wire u2__abc_52155_new_n9127_; 
wire u2__abc_52155_new_n9128_; 
wire u2__abc_52155_new_n9129_; 
wire u2__abc_52155_new_n9130_; 
wire u2__abc_52155_new_n9132_; 
wire u2__abc_52155_new_n9133_; 
wire u2__abc_52155_new_n9134_; 
wire u2__abc_52155_new_n9135_; 
wire u2__abc_52155_new_n9136_; 
wire u2__abc_52155_new_n9137_; 
wire u2__abc_52155_new_n9138_; 
wire u2__abc_52155_new_n9139_; 
wire u2__abc_52155_new_n9140_; 
wire u2__abc_52155_new_n9141_; 
wire u2__abc_52155_new_n9142_; 
wire u2__abc_52155_new_n9143_; 
wire u2__abc_52155_new_n9144_; 
wire u2__abc_52155_new_n9145_; 
wire u2__abc_52155_new_n9146_; 
wire u2__abc_52155_new_n9147_; 
wire u2__abc_52155_new_n9149_; 
wire u2__abc_52155_new_n9150_; 
wire u2__abc_52155_new_n9151_; 
wire u2__abc_52155_new_n9152_; 
wire u2__abc_52155_new_n9153_; 
wire u2__abc_52155_new_n9154_; 
wire u2__abc_52155_new_n9155_; 
wire u2__abc_52155_new_n9156_; 
wire u2__abc_52155_new_n9157_; 
wire u2__abc_52155_new_n9158_; 
wire u2__abc_52155_new_n9159_; 
wire u2__abc_52155_new_n9160_; 
wire u2__abc_52155_new_n9161_; 
wire u2__abc_52155_new_n9162_; 
wire u2__abc_52155_new_n9163_; 
wire u2__abc_52155_new_n9164_; 
wire u2__abc_52155_new_n9166_; 
wire u2__abc_52155_new_n9167_; 
wire u2__abc_52155_new_n9168_; 
wire u2__abc_52155_new_n9169_; 
wire u2__abc_52155_new_n9170_; 
wire u2__abc_52155_new_n9171_; 
wire u2__abc_52155_new_n9172_; 
wire u2__abc_52155_new_n9173_; 
wire u2__abc_52155_new_n9174_; 
wire u2__abc_52155_new_n9175_; 
wire u2__abc_52155_new_n9176_; 
wire u2__abc_52155_new_n9177_; 
wire u2__abc_52155_new_n9178_; 
wire u2__abc_52155_new_n9179_; 
wire u2__abc_52155_new_n9180_; 
wire u2__abc_52155_new_n9181_; 
wire u2__abc_52155_new_n9183_; 
wire u2__abc_52155_new_n9184_; 
wire u2__abc_52155_new_n9185_; 
wire u2__abc_52155_new_n9186_; 
wire u2__abc_52155_new_n9187_; 
wire u2__abc_52155_new_n9188_; 
wire u2__abc_52155_new_n9189_; 
wire u2__abc_52155_new_n9190_; 
wire u2__abc_52155_new_n9191_; 
wire u2__abc_52155_new_n9192_; 
wire u2__abc_52155_new_n9193_; 
wire u2__abc_52155_new_n9194_; 
wire u2__abc_52155_new_n9195_; 
wire u2__abc_52155_new_n9196_; 
wire u2__abc_52155_new_n9197_; 
wire u2__abc_52155_new_n9198_; 
wire u2__abc_52155_new_n9199_; 
wire u2__abc_52155_new_n9200_; 
wire u2__abc_52155_new_n9201_; 
wire u2__abc_52155_new_n9202_; 
wire u2__abc_52155_new_n9203_; 
wire u2__abc_52155_new_n9204_; 
wire u2__abc_52155_new_n9205_; 
wire u2__abc_52155_new_n9206_; 
wire u2__abc_52155_new_n9207_; 
wire u2__abc_52155_new_n9208_; 
wire u2__abc_52155_new_n9210_; 
wire u2__abc_52155_new_n9211_; 
wire u2__abc_52155_new_n9212_; 
wire u2__abc_52155_new_n9213_; 
wire u2__abc_52155_new_n9214_; 
wire u2__abc_52155_new_n9215_; 
wire u2__abc_52155_new_n9216_; 
wire u2__abc_52155_new_n9217_; 
wire u2__abc_52155_new_n9218_; 
wire u2__abc_52155_new_n9219_; 
wire u2__abc_52155_new_n9220_; 
wire u2__abc_52155_new_n9221_; 
wire u2__abc_52155_new_n9222_; 
wire u2__abc_52155_new_n9223_; 
wire u2__abc_52155_new_n9224_; 
wire u2__abc_52155_new_n9225_; 
wire u2__abc_52155_new_n9227_; 
wire u2__abc_52155_new_n9228_; 
wire u2__abc_52155_new_n9229_; 
wire u2__abc_52155_new_n9230_; 
wire u2__abc_52155_new_n9231_; 
wire u2__abc_52155_new_n9232_; 
wire u2__abc_52155_new_n9233_; 
wire u2__abc_52155_new_n9234_; 
wire u2__abc_52155_new_n9235_; 
wire u2__abc_52155_new_n9236_; 
wire u2__abc_52155_new_n9237_; 
wire u2__abc_52155_new_n9238_; 
wire u2__abc_52155_new_n9239_; 
wire u2__abc_52155_new_n9240_; 
wire u2__abc_52155_new_n9241_; 
wire u2__abc_52155_new_n9242_; 
wire u2__abc_52155_new_n9243_; 
wire u2__abc_52155_new_n9244_; 
wire u2__abc_52155_new_n9245_; 
wire u2__abc_52155_new_n9246_; 
wire u2__abc_52155_new_n9248_; 
wire u2__abc_52155_new_n9249_; 
wire u2__abc_52155_new_n9250_; 
wire u2__abc_52155_new_n9251_; 
wire u2__abc_52155_new_n9252_; 
wire u2__abc_52155_new_n9253_; 
wire u2__abc_52155_new_n9254_; 
wire u2__abc_52155_new_n9255_; 
wire u2__abc_52155_new_n9256_; 
wire u2__abc_52155_new_n9257_; 
wire u2__abc_52155_new_n9258_; 
wire u2__abc_52155_new_n9259_; 
wire u2__abc_52155_new_n9260_; 
wire u2__abc_52155_new_n9261_; 
wire u2__abc_52155_new_n9262_; 
wire u2__abc_52155_new_n9263_; 
wire u2__abc_52155_new_n9264_; 
wire u2__abc_52155_new_n9266_; 
wire u2__abc_52155_new_n9267_; 
wire u2__abc_52155_new_n9268_; 
wire u2__abc_52155_new_n9269_; 
wire u2__abc_52155_new_n9270_; 
wire u2__abc_52155_new_n9271_; 
wire u2__abc_52155_new_n9272_; 
wire u2__abc_52155_new_n9273_; 
wire u2__abc_52155_new_n9274_; 
wire u2__abc_52155_new_n9275_; 
wire u2__abc_52155_new_n9276_; 
wire u2__abc_52155_new_n9277_; 
wire u2__abc_52155_new_n9278_; 
wire u2__abc_52155_new_n9279_; 
wire u2__abc_52155_new_n9280_; 
wire u2__abc_52155_new_n9281_; 
wire u2__abc_52155_new_n9282_; 
wire u2__abc_52155_new_n9283_; 
wire u2__abc_52155_new_n9284_; 
wire u2__abc_52155_new_n9285_; 
wire u2__abc_52155_new_n9286_; 
wire u2__abc_52155_new_n9287_; 
wire u2__abc_52155_new_n9289_; 
wire u2__abc_52155_new_n9290_; 
wire u2__abc_52155_new_n9291_; 
wire u2__abc_52155_new_n9292_; 
wire u2__abc_52155_new_n9293_; 
wire u2__abc_52155_new_n9294_; 
wire u2__abc_52155_new_n9295_; 
wire u2__abc_52155_new_n9296_; 
wire u2__abc_52155_new_n9297_; 
wire u2__abc_52155_new_n9298_; 
wire u2__abc_52155_new_n9299_; 
wire u2__abc_52155_new_n9300_; 
wire u2__abc_52155_new_n9301_; 
wire u2__abc_52155_new_n9302_; 
wire u2__abc_52155_new_n9303_; 
wire u2__abc_52155_new_n9304_; 
wire u2__abc_52155_new_n9306_; 
wire u2__abc_52155_new_n9307_; 
wire u2__abc_52155_new_n9308_; 
wire u2__abc_52155_new_n9309_; 
wire u2__abc_52155_new_n9310_; 
wire u2__abc_52155_new_n9311_; 
wire u2__abc_52155_new_n9312_; 
wire u2__abc_52155_new_n9313_; 
wire u2__abc_52155_new_n9314_; 
wire u2__abc_52155_new_n9315_; 
wire u2__abc_52155_new_n9316_; 
wire u2__abc_52155_new_n9317_; 
wire u2__abc_52155_new_n9318_; 
wire u2__abc_52155_new_n9319_; 
wire u2__abc_52155_new_n9320_; 
wire u2__abc_52155_new_n9321_; 
wire u2__abc_52155_new_n9322_; 
wire u2__abc_52155_new_n9323_; 
wire u2__abc_52155_new_n9325_; 
wire u2__abc_52155_new_n9326_; 
wire u2__abc_52155_new_n9327_; 
wire u2__abc_52155_new_n9328_; 
wire u2__abc_52155_new_n9329_; 
wire u2__abc_52155_new_n9330_; 
wire u2__abc_52155_new_n9331_; 
wire u2__abc_52155_new_n9332_; 
wire u2__abc_52155_new_n9333_; 
wire u2__abc_52155_new_n9334_; 
wire u2__abc_52155_new_n9335_; 
wire u2__abc_52155_new_n9336_; 
wire u2__abc_52155_new_n9337_; 
wire u2__abc_52155_new_n9338_; 
wire u2__abc_52155_new_n9339_; 
wire u2__abc_52155_new_n9340_; 
wire u2__abc_52155_new_n9342_; 
wire u2__abc_52155_new_n9343_; 
wire u2__abc_52155_new_n9344_; 
wire u2__abc_52155_new_n9345_; 
wire u2__abc_52155_new_n9346_; 
wire u2__abc_52155_new_n9347_; 
wire u2__abc_52155_new_n9348_; 
wire u2__abc_52155_new_n9349_; 
wire u2__abc_52155_new_n9350_; 
wire u2__abc_52155_new_n9351_; 
wire u2__abc_52155_new_n9352_; 
wire u2__abc_52155_new_n9353_; 
wire u2__abc_52155_new_n9354_; 
wire u2__abc_52155_new_n9355_; 
wire u2__abc_52155_new_n9356_; 
wire u2__abc_52155_new_n9357_; 
wire u2__abc_52155_new_n9358_; 
wire u2__abc_52155_new_n9359_; 
wire u2__abc_52155_new_n9360_; 
wire u2__abc_52155_new_n9361_; 
wire u2__abc_52155_new_n9362_; 
wire u2__abc_52155_new_n9363_; 
wire u2__abc_52155_new_n9364_; 
wire u2__abc_52155_new_n9365_; 
wire u2__abc_52155_new_n9366_; 
wire u2__abc_52155_new_n9367_; 
wire u2__abc_52155_new_n9368_; 
wire u2__abc_52155_new_n9370_; 
wire u2__abc_52155_new_n9371_; 
wire u2__abc_52155_new_n9372_; 
wire u2__abc_52155_new_n9373_; 
wire u2__abc_52155_new_n9374_; 
wire u2__abc_52155_new_n9375_; 
wire u2__abc_52155_new_n9376_; 
wire u2__abc_52155_new_n9377_; 
wire u2__abc_52155_new_n9378_; 
wire u2__abc_52155_new_n9379_; 
wire u2__abc_52155_new_n9380_; 
wire u2__abc_52155_new_n9381_; 
wire u2__abc_52155_new_n9382_; 
wire u2__abc_52155_new_n9383_; 
wire u2__abc_52155_new_n9384_; 
wire u2__abc_52155_new_n9385_; 
wire u2__abc_52155_new_n9387_; 
wire u2__abc_52155_new_n9388_; 
wire u2__abc_52155_new_n9389_; 
wire u2__abc_52155_new_n9390_; 
wire u2__abc_52155_new_n9391_; 
wire u2__abc_52155_new_n9392_; 
wire u2__abc_52155_new_n9393_; 
wire u2__abc_52155_new_n9394_; 
wire u2__abc_52155_new_n9395_; 
wire u2__abc_52155_new_n9396_; 
wire u2__abc_52155_new_n9397_; 
wire u2__abc_52155_new_n9398_; 
wire u2__abc_52155_new_n9399_; 
wire u2__abc_52155_new_n9400_; 
wire u2__abc_52155_new_n9401_; 
wire u2__abc_52155_new_n9402_; 
wire u2__abc_52155_new_n9403_; 
wire u2__abc_52155_new_n9404_; 
wire u2__abc_52155_new_n9405_; 
wire u2__abc_52155_new_n9407_; 
wire u2__abc_52155_new_n9408_; 
wire u2__abc_52155_new_n9409_; 
wire u2__abc_52155_new_n9410_; 
wire u2__abc_52155_new_n9411_; 
wire u2__abc_52155_new_n9412_; 
wire u2__abc_52155_new_n9413_; 
wire u2__abc_52155_new_n9414_; 
wire u2__abc_52155_new_n9415_; 
wire u2__abc_52155_new_n9416_; 
wire u2__abc_52155_new_n9417_; 
wire u2__abc_52155_new_n9418_; 
wire u2__abc_52155_new_n9419_; 
wire u2__abc_52155_new_n9420_; 
wire u2__abc_52155_new_n9421_; 
wire u2__abc_52155_new_n9422_; 
wire u2__abc_52155_new_n9424_; 
wire u2__abc_52155_new_n9425_; 
wire u2__abc_52155_new_n9426_; 
wire u2__abc_52155_new_n9427_; 
wire u2__abc_52155_new_n9428_; 
wire u2__abc_52155_new_n9429_; 
wire u2__abc_52155_new_n9430_; 
wire u2__abc_52155_new_n9431_; 
wire u2__abc_52155_new_n9432_; 
wire u2__abc_52155_new_n9433_; 
wire u2__abc_52155_new_n9434_; 
wire u2__abc_52155_new_n9435_; 
wire u2__abc_52155_new_n9436_; 
wire u2__abc_52155_new_n9437_; 
wire u2__abc_52155_new_n9438_; 
wire u2__abc_52155_new_n9439_; 
wire u2__abc_52155_new_n9440_; 
wire u2__abc_52155_new_n9441_; 
wire u2__abc_52155_new_n9443_; 
wire u2__abc_52155_new_n9444_; 
wire u2__abc_52155_new_n9445_; 
wire u2__abc_52155_new_n9446_; 
wire u2__abc_52155_new_n9447_; 
wire u2__abc_52155_new_n9448_; 
wire u2__abc_52155_new_n9449_; 
wire u2__abc_52155_new_n9450_; 
wire u2__abc_52155_new_n9451_; 
wire u2__abc_52155_new_n9452_; 
wire u2__abc_52155_new_n9453_; 
wire u2__abc_52155_new_n9454_; 
wire u2__abc_52155_new_n9455_; 
wire u2__abc_52155_new_n9456_; 
wire u2__abc_52155_new_n9457_; 
wire u2__abc_52155_new_n9458_; 
wire u2__abc_52155_new_n9460_; 
wire u2__abc_52155_new_n9461_; 
wire u2__abc_52155_new_n9462_; 
wire u2__abc_52155_new_n9463_; 
wire u2__abc_52155_new_n9464_; 
wire u2__abc_52155_new_n9465_; 
wire u2__abc_52155_new_n9466_; 
wire u2__abc_52155_new_n9467_; 
wire u2__abc_52155_new_n9468_; 
wire u2__abc_52155_new_n9469_; 
wire u2__abc_52155_new_n9470_; 
wire u2__abc_52155_new_n9471_; 
wire u2__abc_52155_new_n9472_; 
wire u2__abc_52155_new_n9473_; 
wire u2__abc_52155_new_n9474_; 
wire u2__abc_52155_new_n9475_; 
wire u2__abc_52155_new_n9476_; 
wire u2__abc_52155_new_n9477_; 
wire u2__abc_52155_new_n9479_; 
wire u2__abc_52155_new_n9480_; 
wire u2__abc_52155_new_n9481_; 
wire u2__abc_52155_new_n9482_; 
wire u2__abc_52155_new_n9483_; 
wire u2__abc_52155_new_n9484_; 
wire u2__abc_52155_new_n9485_; 
wire u2__abc_52155_new_n9486_; 
wire u2__abc_52155_new_n9487_; 
wire u2__abc_52155_new_n9488_; 
wire u2__abc_52155_new_n9489_; 
wire u2__abc_52155_new_n9490_; 
wire u2__abc_52155_new_n9491_; 
wire u2__abc_52155_new_n9492_; 
wire u2__abc_52155_new_n9493_; 
wire u2__abc_52155_new_n9494_; 
wire u2__abc_52155_new_n9496_; 
wire u2__abc_52155_new_n9497_; 
wire u2__abc_52155_new_n9498_; 
wire u2__abc_52155_new_n9499_; 
wire u2__abc_52155_new_n9500_; 
wire u2__abc_52155_new_n9501_; 
wire u2__abc_52155_new_n9502_; 
wire u2__abc_52155_new_n9503_; 
wire u2__abc_52155_new_n9504_; 
wire u2__abc_52155_new_n9505_; 
wire u2__abc_52155_new_n9506_; 
wire u2__abc_52155_new_n9507_; 
wire u2__abc_52155_new_n9508_; 
wire u2__abc_52155_new_n9509_; 
wire u2__abc_52155_new_n9510_; 
wire u2__abc_52155_new_n9511_; 
wire u2__abc_52155_new_n9512_; 
wire u2__abc_52155_new_n9513_; 
wire u2__abc_52155_new_n9514_; 
wire u2__abc_52155_new_n9515_; 
wire u2__abc_52155_new_n9516_; 
wire u2__abc_52155_new_n9517_; 
wire u2__abc_52155_new_n9518_; 
wire u2__abc_52155_new_n9519_; 
wire u2__abc_52155_new_n9520_; 
wire u2__abc_52155_new_n9521_; 
wire u2__abc_52155_new_n9522_; 
wire u2__abc_52155_new_n9523_; 
wire u2__abc_52155_new_n9524_; 
wire u2__abc_52155_new_n9525_; 
wire u2__abc_52155_new_n9526_; 
wire u2__abc_52155_new_n9527_; 
wire u2__abc_52155_new_n9528_; 
wire u2__abc_52155_new_n9529_; 
wire u2__abc_52155_new_n9530_; 
wire u2__abc_52155_new_n9531_; 
wire u2__abc_52155_new_n9532_; 
wire u2__abc_52155_new_n9533_; 
wire u2__abc_52155_new_n9535_; 
wire u2__abc_52155_new_n9536_; 
wire u2__abc_52155_new_n9537_; 
wire u2__abc_52155_new_n9538_; 
wire u2__abc_52155_new_n9539_; 
wire u2__abc_52155_new_n9540_; 
wire u2__abc_52155_new_n9541_; 
wire u2__abc_52155_new_n9542_; 
wire u2__abc_52155_new_n9543_; 
wire u2__abc_52155_new_n9544_; 
wire u2__abc_52155_new_n9545_; 
wire u2__abc_52155_new_n9546_; 
wire u2__abc_52155_new_n9547_; 
wire u2__abc_52155_new_n9548_; 
wire u2__abc_52155_new_n9549_; 
wire u2__abc_52155_new_n9550_; 
wire u2__abc_52155_new_n9552_; 
wire u2__abc_52155_new_n9553_; 
wire u2__abc_52155_new_n9554_; 
wire u2__abc_52155_new_n9555_; 
wire u2__abc_52155_new_n9556_; 
wire u2__abc_52155_new_n9557_; 
wire u2__abc_52155_new_n9558_; 
wire u2__abc_52155_new_n9559_; 
wire u2__abc_52155_new_n9560_; 
wire u2__abc_52155_new_n9561_; 
wire u2__abc_52155_new_n9562_; 
wire u2__abc_52155_new_n9563_; 
wire u2__abc_52155_new_n9564_; 
wire u2__abc_52155_new_n9565_; 
wire u2__abc_52155_new_n9566_; 
wire u2__abc_52155_new_n9567_; 
wire u2__abc_52155_new_n9568_; 
wire u2__abc_52155_new_n9569_; 
wire u2__abc_52155_new_n9570_; 
wire u2__abc_52155_new_n9572_; 
wire u2__abc_52155_new_n9573_; 
wire u2__abc_52155_new_n9574_; 
wire u2__abc_52155_new_n9575_; 
wire u2__abc_52155_new_n9576_; 
wire u2__abc_52155_new_n9577_; 
wire u2__abc_52155_new_n9578_; 
wire u2__abc_52155_new_n9579_; 
wire u2__abc_52155_new_n9580_; 
wire u2__abc_52155_new_n9581_; 
wire u2__abc_52155_new_n9582_; 
wire u2__abc_52155_new_n9583_; 
wire u2__abc_52155_new_n9584_; 
wire u2__abc_52155_new_n9585_; 
wire u2__abc_52155_new_n9586_; 
wire u2__abc_52155_new_n9587_; 
wire u2__abc_52155_new_n9588_; 
wire u2__abc_52155_new_n9590_; 
wire u2__abc_52155_new_n9591_; 
wire u2__abc_52155_new_n9592_; 
wire u2__abc_52155_new_n9593_; 
wire u2__abc_52155_new_n9594_; 
wire u2__abc_52155_new_n9595_; 
wire u2__abc_52155_new_n9596_; 
wire u2__abc_52155_new_n9597_; 
wire u2__abc_52155_new_n9598_; 
wire u2__abc_52155_new_n9599_; 
wire u2__abc_52155_new_n9600_; 
wire u2__abc_52155_new_n9601_; 
wire u2__abc_52155_new_n9602_; 
wire u2__abc_52155_new_n9603_; 
wire u2__abc_52155_new_n9604_; 
wire u2__abc_52155_new_n9605_; 
wire u2__abc_52155_new_n9606_; 
wire u2__abc_52155_new_n9607_; 
wire u2__abc_52155_new_n9608_; 
wire u2__abc_52155_new_n9609_; 
wire u2__abc_52155_new_n9610_; 
wire u2__abc_52155_new_n9611_; 
wire u2__abc_52155_new_n9613_; 
wire u2__abc_52155_new_n9614_; 
wire u2__abc_52155_new_n9615_; 
wire u2__abc_52155_new_n9616_; 
wire u2__abc_52155_new_n9617_; 
wire u2__abc_52155_new_n9618_; 
wire u2__abc_52155_new_n9619_; 
wire u2__abc_52155_new_n9620_; 
wire u2__abc_52155_new_n9621_; 
wire u2__abc_52155_new_n9622_; 
wire u2__abc_52155_new_n9623_; 
wire u2__abc_52155_new_n9624_; 
wire u2__abc_52155_new_n9625_; 
wire u2__abc_52155_new_n9626_; 
wire u2__abc_52155_new_n9627_; 
wire u2__abc_52155_new_n9628_; 
wire u2__abc_52155_new_n9630_; 
wire u2__abc_52155_new_n9631_; 
wire u2__abc_52155_new_n9632_; 
wire u2__abc_52155_new_n9633_; 
wire u2__abc_52155_new_n9634_; 
wire u2__abc_52155_new_n9635_; 
wire u2__abc_52155_new_n9636_; 
wire u2__abc_52155_new_n9637_; 
wire u2__abc_52155_new_n9638_; 
wire u2__abc_52155_new_n9639_; 
wire u2__abc_52155_new_n9640_; 
wire u2__abc_52155_new_n9641_; 
wire u2__abc_52155_new_n9642_; 
wire u2__abc_52155_new_n9643_; 
wire u2__abc_52155_new_n9644_; 
wire u2__abc_52155_new_n9645_; 
wire u2__abc_52155_new_n9646_; 
wire u2__abc_52155_new_n9647_; 
wire u2__abc_52155_new_n9649_; 
wire u2__abc_52155_new_n9650_; 
wire u2__abc_52155_new_n9651_; 
wire u2__abc_52155_new_n9652_; 
wire u2__abc_52155_new_n9653_; 
wire u2__abc_52155_new_n9654_; 
wire u2__abc_52155_new_n9655_; 
wire u2__abc_52155_new_n9656_; 
wire u2__abc_52155_new_n9657_; 
wire u2__abc_52155_new_n9658_; 
wire u2__abc_52155_new_n9659_; 
wire u2__abc_52155_new_n9660_; 
wire u2__abc_52155_new_n9661_; 
wire u2__abc_52155_new_n9662_; 
wire u2__abc_52155_new_n9663_; 
wire u2__abc_52155_new_n9664_; 
wire u2__abc_52155_new_n9666_; 
wire u2__abc_52155_new_n9667_; 
wire u2__abc_52155_new_n9668_; 
wire u2__abc_52155_new_n9669_; 
wire u2__abc_52155_new_n9670_; 
wire u2__abc_52155_new_n9671_; 
wire u2__abc_52155_new_n9672_; 
wire u2__abc_52155_new_n9673_; 
wire u2__abc_52155_new_n9674_; 
wire u2__abc_52155_new_n9675_; 
wire u2__abc_52155_new_n9676_; 
wire u2__abc_52155_new_n9677_; 
wire u2__abc_52155_new_n9678_; 
wire u2__abc_52155_new_n9679_; 
wire u2__abc_52155_new_n9680_; 
wire u2__abc_52155_new_n9681_; 
wire u2__abc_52155_new_n9682_; 
wire u2__abc_52155_new_n9683_; 
wire u2__abc_52155_new_n9684_; 
wire u2__abc_52155_new_n9685_; 
wire u2__abc_52155_new_n9686_; 
wire u2__abc_52155_new_n9687_; 
wire u2__abc_52155_new_n9688_; 
wire u2__abc_52155_new_n9689_; 
wire u2__abc_52155_new_n9691_; 
wire u2__abc_52155_new_n9692_; 
wire u2__abc_52155_new_n9693_; 
wire u2__abc_52155_new_n9694_; 
wire u2__abc_52155_new_n9695_; 
wire u2__abc_52155_new_n9696_; 
wire u2__abc_52155_new_n9697_; 
wire u2__abc_52155_new_n9698_; 
wire u2__abc_52155_new_n9699_; 
wire u2__abc_52155_new_n9700_; 
wire u2__abc_52155_new_n9701_; 
wire u2__abc_52155_new_n9702_; 
wire u2__abc_52155_new_n9703_; 
wire u2__abc_52155_new_n9704_; 
wire u2__abc_52155_new_n9705_; 
wire u2__abc_52155_new_n9706_; 
wire u2__abc_52155_new_n9708_; 
wire u2__abc_52155_new_n9709_; 
wire u2__abc_52155_new_n9710_; 
wire u2__abc_52155_new_n9711_; 
wire u2__abc_52155_new_n9712_; 
wire u2__abc_52155_new_n9713_; 
wire u2__abc_52155_new_n9714_; 
wire u2__abc_52155_new_n9715_; 
wire u2__abc_52155_new_n9716_; 
wire u2__abc_52155_new_n9717_; 
wire u2__abc_52155_new_n9718_; 
wire u2__abc_52155_new_n9719_; 
wire u2__abc_52155_new_n9720_; 
wire u2__abc_52155_new_n9721_; 
wire u2__abc_52155_new_n9722_; 
wire u2__abc_52155_new_n9723_; 
wire u2__abc_52155_new_n9724_; 
wire u2__abc_52155_new_n9725_; 
wire u2__abc_52155_new_n9727_; 
wire u2__abc_52155_new_n9728_; 
wire u2__abc_52155_new_n9729_; 
wire u2__abc_52155_new_n9730_; 
wire u2__abc_52155_new_n9731_; 
wire u2__abc_52155_new_n9732_; 
wire u2__abc_52155_new_n9733_; 
wire u2__abc_52155_new_n9734_; 
wire u2__abc_52155_new_n9735_; 
wire u2__abc_52155_new_n9736_; 
wire u2__abc_52155_new_n9737_; 
wire u2__abc_52155_new_n9738_; 
wire u2__abc_52155_new_n9739_; 
wire u2__abc_52155_new_n9740_; 
wire u2__abc_52155_new_n9741_; 
wire u2__abc_52155_new_n9742_; 
wire u2__abc_52155_new_n9744_; 
wire u2__abc_52155_new_n9745_; 
wire u2__abc_52155_new_n9746_; 
wire u2__abc_52155_new_n9747_; 
wire u2__abc_52155_new_n9748_; 
wire u2__abc_52155_new_n9749_; 
wire u2__abc_52155_new_n9750_; 
wire u2__abc_52155_new_n9751_; 
wire u2__abc_52155_new_n9752_; 
wire u2__abc_52155_new_n9753_; 
wire u2__abc_52155_new_n9754_; 
wire u2__abc_52155_new_n9755_; 
wire u2__abc_52155_new_n9756_; 
wire u2__abc_52155_new_n9757_; 
wire u2__abc_52155_new_n9758_; 
wire u2__abc_52155_new_n9759_; 
wire u2__abc_52155_new_n9760_; 
wire u2__abc_52155_new_n9761_; 
wire u2__abc_52155_new_n9762_; 
wire u2__abc_52155_new_n9763_; 
wire u2__abc_52155_new_n9764_; 
wire u2__abc_52155_new_n9765_; 
wire u2__abc_52155_new_n9767_; 
wire u2__abc_52155_new_n9768_; 
wire u2__abc_52155_new_n9769_; 
wire u2__abc_52155_new_n9770_; 
wire u2__abc_52155_new_n9771_; 
wire u2__abc_52155_new_n9772_; 
wire u2__abc_52155_new_n9773_; 
wire u2__abc_52155_new_n9774_; 
wire u2__abc_52155_new_n9775_; 
wire u2__abc_52155_new_n9776_; 
wire u2__abc_52155_new_n9777_; 
wire u2__abc_52155_new_n9778_; 
wire u2__abc_52155_new_n9779_; 
wire u2__abc_52155_new_n9780_; 
wire u2__abc_52155_new_n9781_; 
wire u2__abc_52155_new_n9782_; 
wire u2__abc_52155_new_n9784_; 
wire u2__abc_52155_new_n9785_; 
wire u2__abc_52155_new_n9786_; 
wire u2__abc_52155_new_n9787_; 
wire u2__abc_52155_new_n9788_; 
wire u2__abc_52155_new_n9789_; 
wire u2__abc_52155_new_n9790_; 
wire u2__abc_52155_new_n9791_; 
wire u2__abc_52155_new_n9792_; 
wire u2__abc_52155_new_n9793_; 
wire u2__abc_52155_new_n9794_; 
wire u2__abc_52155_new_n9795_; 
wire u2__abc_52155_new_n9796_; 
wire u2__abc_52155_new_n9797_; 
wire u2__abc_52155_new_n9798_; 
wire u2__abc_52155_new_n9799_; 
wire u2__abc_52155_new_n9800_; 
wire u2__abc_52155_new_n9801_; 
wire u2__abc_52155_new_n9803_; 
wire u2__abc_52155_new_n9804_; 
wire u2__abc_52155_new_n9805_; 
wire u2__abc_52155_new_n9806_; 
wire u2__abc_52155_new_n9807_; 
wire u2__abc_52155_new_n9808_; 
wire u2__abc_52155_new_n9809_; 
wire u2__abc_52155_new_n9810_; 
wire u2__abc_52155_new_n9811_; 
wire u2__abc_52155_new_n9812_; 
wire u2__abc_52155_new_n9813_; 
wire u2__abc_52155_new_n9814_; 
wire u2__abc_52155_new_n9815_; 
wire u2__abc_52155_new_n9816_; 
wire u2__abc_52155_new_n9817_; 
wire u2__abc_52155_new_n9818_; 
wire u2__abc_52155_new_n9820_; 
wire u2__abc_52155_new_n9821_; 
wire u2__abc_52155_new_n9822_; 
wire u2__abc_52155_new_n9823_; 
wire u2__abc_52155_new_n9824_; 
wire u2__abc_52155_new_n9825_; 
wire u2__abc_52155_new_n9826_; 
wire u2__abc_52155_new_n9827_; 
wire u2__abc_52155_new_n9828_; 
wire u2__abc_52155_new_n9829_; 
wire u2__abc_52155_new_n9830_; 
wire u2__abc_52155_new_n9831_; 
wire u2__abc_52155_new_n9832_; 
wire u2__abc_52155_new_n9833_; 
wire u2__abc_52155_new_n9834_; 
wire u2__abc_52155_new_n9835_; 
wire u2__abc_52155_new_n9836_; 
wire u2__abc_52155_new_n9837_; 
wire u2__abc_52155_new_n9838_; 
wire u2__abc_52155_new_n9839_; 
wire u2__abc_52155_new_n9840_; 
wire u2__abc_52155_new_n9841_; 
wire u2__abc_52155_new_n9842_; 
wire u2__abc_52155_new_n9843_; 
wire u2__abc_52155_new_n9844_; 
wire u2__abc_52155_new_n9845_; 
wire u2__abc_52155_new_n9847_; 
wire u2__abc_52155_new_n9848_; 
wire u2__abc_52155_new_n9849_; 
wire u2__abc_52155_new_n9850_; 
wire u2__abc_52155_new_n9851_; 
wire u2__abc_52155_new_n9852_; 
wire u2__abc_52155_new_n9853_; 
wire u2__abc_52155_new_n9854_; 
wire u2__abc_52155_new_n9855_; 
wire u2__abc_52155_new_n9856_; 
wire u2__abc_52155_new_n9857_; 
wire u2__abc_52155_new_n9858_; 
wire u2__abc_52155_new_n9859_; 
wire u2__abc_52155_new_n9860_; 
wire u2__abc_52155_new_n9861_; 
wire u2__abc_52155_new_n9862_; 
wire u2__abc_52155_new_n9864_; 
wire u2__abc_52155_new_n9865_; 
wire u2__abc_52155_new_n9866_; 
wire u2__abc_52155_new_n9867_; 
wire u2__abc_52155_new_n9868_; 
wire u2__abc_52155_new_n9869_; 
wire u2__abc_52155_new_n9870_; 
wire u2__abc_52155_new_n9871_; 
wire u2__abc_52155_new_n9872_; 
wire u2__abc_52155_new_n9873_; 
wire u2__abc_52155_new_n9874_; 
wire u2__abc_52155_new_n9875_; 
wire u2__abc_52155_new_n9876_; 
wire u2__abc_52155_new_n9877_; 
wire u2__abc_52155_new_n9878_; 
wire u2__abc_52155_new_n9879_; 
wire u2__abc_52155_new_n9880_; 
wire u2__abc_52155_new_n9881_; 
wire u2__abc_52155_new_n9882_; 
wire u2__abc_52155_new_n9884_; 
wire u2__abc_52155_new_n9885_; 
wire u2__abc_52155_new_n9886_; 
wire u2__abc_52155_new_n9887_; 
wire u2__abc_52155_new_n9888_; 
wire u2__abc_52155_new_n9889_; 
wire u2__abc_52155_new_n9890_; 
wire u2__abc_52155_new_n9891_; 
wire u2__abc_52155_new_n9892_; 
wire u2__abc_52155_new_n9893_; 
wire u2__abc_52155_new_n9894_; 
wire u2__abc_52155_new_n9895_; 
wire u2__abc_52155_new_n9896_; 
wire u2__abc_52155_new_n9897_; 
wire u2__abc_52155_new_n9898_; 
wire u2__abc_52155_new_n9899_; 
wire u2__abc_52155_new_n9901_; 
wire u2__abc_52155_new_n9902_; 
wire u2__abc_52155_new_n9903_; 
wire u2__abc_52155_new_n9904_; 
wire u2__abc_52155_new_n9905_; 
wire u2__abc_52155_new_n9906_; 
wire u2__abc_52155_new_n9907_; 
wire u2__abc_52155_new_n9908_; 
wire u2__abc_52155_new_n9909_; 
wire u2__abc_52155_new_n9910_; 
wire u2__abc_52155_new_n9911_; 
wire u2__abc_52155_new_n9912_; 
wire u2__abc_52155_new_n9913_; 
wire u2__abc_52155_new_n9914_; 
wire u2__abc_52155_new_n9915_; 
wire u2__abc_52155_new_n9916_; 
wire u2__abc_52155_new_n9917_; 
wire u2__abc_52155_new_n9918_; 
wire u2__abc_52155_new_n9919_; 
wire u2__abc_52155_new_n9920_; 
wire u2__abc_52155_new_n9922_; 
wire u2__abc_52155_new_n9923_; 
wire u2__abc_52155_new_n9924_; 
wire u2__abc_52155_new_n9925_; 
wire u2__abc_52155_new_n9926_; 
wire u2__abc_52155_new_n9927_; 
wire u2__abc_52155_new_n9928_; 
wire u2__abc_52155_new_n9929_; 
wire u2__abc_52155_new_n9930_; 
wire u2__abc_52155_new_n9931_; 
wire u2__abc_52155_new_n9932_; 
wire u2__abc_52155_new_n9933_; 
wire u2__abc_52155_new_n9934_; 
wire u2__abc_52155_new_n9935_; 
wire u2__abc_52155_new_n9936_; 
wire u2__abc_52155_new_n9937_; 
wire u2__abc_52155_new_n9939_; 
wire u2__abc_52155_new_n9940_; 
wire u2__abc_52155_new_n9941_; 
wire u2__abc_52155_new_n9942_; 
wire u2__abc_52155_new_n9943_; 
wire u2__abc_52155_new_n9944_; 
wire u2__abc_52155_new_n9945_; 
wire u2__abc_52155_new_n9946_; 
wire u2__abc_52155_new_n9947_; 
wire u2__abc_52155_new_n9948_; 
wire u2__abc_52155_new_n9949_; 
wire u2__abc_52155_new_n9950_; 
wire u2__abc_52155_new_n9951_; 
wire u2__abc_52155_new_n9952_; 
wire u2__abc_52155_new_n9953_; 
wire u2__abc_52155_new_n9954_; 
wire u2__abc_52155_new_n9956_; 
wire u2__abc_52155_new_n9957_; 
wire u2__abc_52155_new_n9958_; 
wire u2__abc_52155_new_n9959_; 
wire u2__abc_52155_new_n9960_; 
wire u2__abc_52155_new_n9961_; 
wire u2__abc_52155_new_n9962_; 
wire u2__abc_52155_new_n9963_; 
wire u2__abc_52155_new_n9964_; 
wire u2__abc_52155_new_n9965_; 
wire u2__abc_52155_new_n9966_; 
wire u2__abc_52155_new_n9967_; 
wire u2__abc_52155_new_n9968_; 
wire u2__abc_52155_new_n9969_; 
wire u2__abc_52155_new_n9970_; 
wire u2__abc_52155_new_n9971_; 
wire u2__abc_52155_new_n9973_; 
wire u2__abc_52155_new_n9974_; 
wire u2__abc_52155_new_n9975_; 
wire u2__abc_52155_new_n9976_; 
wire u2__abc_52155_new_n9977_; 
wire u2__abc_52155_new_n9978_; 
wire u2__abc_52155_new_n9979_; 
wire u2__abc_52155_new_n9980_; 
wire u2__abc_52155_new_n9981_; 
wire u2__abc_52155_new_n9982_; 
wire u2__abc_52155_new_n9983_; 
wire u2__abc_52155_new_n9984_; 
wire u2__abc_52155_new_n9985_; 
wire u2__abc_52155_new_n9986_; 
wire u2__abc_52155_new_n9987_; 
wire u2__abc_52155_new_n9988_; 
wire u2__abc_52155_new_n9989_; 
wire u2__abc_52155_new_n9990_; 
wire u2__abc_52155_new_n9991_; 
wire u2__abc_52155_new_n9992_; 
wire u2__abc_52155_new_n9993_; 
wire u2__abc_52155_new_n9994_; 
wire u2__abc_52155_new_n9995_; 
wire u2__abc_52155_new_n9996_; 
wire u2__abc_52155_new_n9998_; 
wire u2__abc_52155_new_n9999_; 
wire u2_cnt_0_; 
wire u2_cnt_1_; 
wire u2_cnt_2_; 
wire u2_cnt_3_; 
wire u2_cnt_4_; 
wire u2_cnt_5_; 
wire u2_cnt_6_; 
wire u2_cnt_7_; 
wire u2_o_226_; 
wire u2_o_227_; 
wire u2_o_228_; 
wire u2_o_229_; 
wire u2_o_230_; 
wire u2_o_231_; 
wire u2_o_232_; 
wire u2_o_233_; 
wire u2_o_234_; 
wire u2_o_235_; 
wire u2_o_236_; 
wire u2_o_237_; 
wire u2_o_238_; 
wire u2_o_239_; 
wire u2_o_240_; 
wire u2_o_241_; 
wire u2_o_242_; 
wire u2_o_243_; 
wire u2_o_244_; 
wire u2_o_245_; 
wire u2_o_246_; 
wire u2_o_247_; 
wire u2_o_248_; 
wire u2_o_249_; 
wire u2_o_250_; 
wire u2_o_251_; 
wire u2_o_252_; 
wire u2_o_253_; 
wire u2_o_254_; 
wire u2_o_255_; 
wire u2_o_256_; 
wire u2_o_257_; 
wire u2_o_258_; 
wire u2_o_259_; 
wire u2_o_260_; 
wire u2_o_261_; 
wire u2_o_262_; 
wire u2_o_263_; 
wire u2_o_264_; 
wire u2_o_265_; 
wire u2_o_266_; 
wire u2_o_267_; 
wire u2_o_268_; 
wire u2_o_269_; 
wire u2_o_270_; 
wire u2_o_271_; 
wire u2_o_272_; 
wire u2_o_273_; 
wire u2_o_274_; 
wire u2_o_275_; 
wire u2_o_276_; 
wire u2_o_277_; 
wire u2_o_278_; 
wire u2_o_279_; 
wire u2_o_280_; 
wire u2_o_281_; 
wire u2_o_282_; 
wire u2_o_283_; 
wire u2_o_284_; 
wire u2_o_285_; 
wire u2_o_286_; 
wire u2_o_287_; 
wire u2_o_288_; 
wire u2_o_289_; 
wire u2_o_290_; 
wire u2_o_291_; 
wire u2_o_292_; 
wire u2_o_293_; 
wire u2_o_294_; 
wire u2_o_295_; 
wire u2_o_296_; 
wire u2_o_297_; 
wire u2_o_298_; 
wire u2_o_299_; 
wire u2_o_300_; 
wire u2_o_301_; 
wire u2_o_302_; 
wire u2_o_303_; 
wire u2_o_304_; 
wire u2_o_305_; 
wire u2_o_306_; 
wire u2_o_307_; 
wire u2_o_308_; 
wire u2_o_309_; 
wire u2_o_310_; 
wire u2_o_311_; 
wire u2_o_312_; 
wire u2_o_313_; 
wire u2_o_314_; 
wire u2_o_315_; 
wire u2_o_316_; 
wire u2_o_317_; 
wire u2_o_318_; 
wire u2_o_319_; 
wire u2_o_320_; 
wire u2_o_321_; 
wire u2_o_322_; 
wire u2_o_323_; 
wire u2_o_324_; 
wire u2_o_325_; 
wire u2_o_326_; 
wire u2_o_327_; 
wire u2_o_328_; 
wire u2_o_329_; 
wire u2_o_330_; 
wire u2_o_331_; 
wire u2_o_332_; 
wire u2_o_333_; 
wire u2_o_334_; 
wire u2_o_335_; 
wire u2_o_336_; 
wire u2_o_337_; 
wire u2_o_338_; 
wire u2_o_339_; 
wire u2_o_340_; 
wire u2_o_341_; 
wire u2_o_342_; 
wire u2_o_343_; 
wire u2_o_344_; 
wire u2_o_345_; 
wire u2_o_346_; 
wire u2_o_347_; 
wire u2_o_348_; 
wire u2_o_349_; 
wire u2_o_350_; 
wire u2_o_351_; 
wire u2_o_352_; 
wire u2_o_353_; 
wire u2_o_354_; 
wire u2_o_355_; 
wire u2_o_356_; 
wire u2_o_357_; 
wire u2_o_358_; 
wire u2_o_359_; 
wire u2_o_360_; 
wire u2_o_361_; 
wire u2_o_362_; 
wire u2_o_363_; 
wire u2_o_364_; 
wire u2_o_365_; 
wire u2_o_366_; 
wire u2_o_367_; 
wire u2_o_368_; 
wire u2_o_369_; 
wire u2_o_370_; 
wire u2_o_371_; 
wire u2_o_372_; 
wire u2_o_373_; 
wire u2_o_374_; 
wire u2_o_375_; 
wire u2_o_376_; 
wire u2_o_377_; 
wire u2_o_378_; 
wire u2_o_379_; 
wire u2_o_380_; 
wire u2_o_381_; 
wire u2_o_382_; 
wire u2_o_383_; 
wire u2_o_384_; 
wire u2_o_385_; 
wire u2_o_386_; 
wire u2_o_387_; 
wire u2_o_388_; 
wire u2_o_389_; 
wire u2_o_390_; 
wire u2_o_391_; 
wire u2_o_392_; 
wire u2_o_393_; 
wire u2_o_394_; 
wire u2_o_395_; 
wire u2_o_396_; 
wire u2_o_397_; 
wire u2_o_398_; 
wire u2_o_399_; 
wire u2_o_400_; 
wire u2_o_401_; 
wire u2_o_402_; 
wire u2_o_403_; 
wire u2_o_404_; 
wire u2_o_405_; 
wire u2_o_406_; 
wire u2_o_407_; 
wire u2_o_408_; 
wire u2_o_409_; 
wire u2_o_410_; 
wire u2_o_411_; 
wire u2_o_412_; 
wire u2_o_413_; 
wire u2_o_414_; 
wire u2_o_415_; 
wire u2_o_416_; 
wire u2_o_417_; 
wire u2_o_418_; 
wire u2_o_419_; 
wire u2_o_420_; 
wire u2_o_421_; 
wire u2_o_422_; 
wire u2_o_423_; 
wire u2_o_424_; 
wire u2_o_425_; 
wire u2_o_426_; 
wire u2_o_427_; 
wire u2_o_428_; 
wire u2_o_429_; 
wire u2_o_430_; 
wire u2_o_431_; 
wire u2_o_432_; 
wire u2_o_433_; 
wire u2_o_434_; 
wire u2_o_435_; 
wire u2_o_436_; 
wire u2_o_437_; 
wire u2_o_438_; 
wire u2_o_439_; 
wire u2_o_440_; 
wire u2_o_441_; 
wire u2_o_442_; 
wire u2_o_443_; 
wire u2_o_444_; 
wire u2_o_445_; 
wire u2_o_446_; 
wire u2_o_447_; 
wire u2_o_448_; 
wire u2_o_449_; 
wire u2_remHiShift_0_; 
wire u2_remHiShift_1_; 
wire u2_remHi_0_; 
wire u2_remHi_100_; 
wire u2_remHi_101_; 
wire u2_remHi_102_; 
wire u2_remHi_103_; 
wire u2_remHi_104_; 
wire u2_remHi_105_; 
wire u2_remHi_106_; 
wire u2_remHi_107_; 
wire u2_remHi_108_; 
wire u2_remHi_109_; 
wire u2_remHi_10_; 
wire u2_remHi_110_; 
wire u2_remHi_111_; 
wire u2_remHi_112_; 
wire u2_remHi_113_; 
wire u2_remHi_114_; 
wire u2_remHi_115_; 
wire u2_remHi_116_; 
wire u2_remHi_117_; 
wire u2_remHi_118_; 
wire u2_remHi_119_; 
wire u2_remHi_11_; 
wire u2_remHi_120_; 
wire u2_remHi_121_; 
wire u2_remHi_122_; 
wire u2_remHi_123_; 
wire u2_remHi_124_; 
wire u2_remHi_125_; 
wire u2_remHi_126_; 
wire u2_remHi_127_; 
wire u2_remHi_128_; 
wire u2_remHi_129_; 
wire u2_remHi_12_; 
wire u2_remHi_130_; 
wire u2_remHi_131_; 
wire u2_remHi_132_; 
wire u2_remHi_133_; 
wire u2_remHi_134_; 
wire u2_remHi_135_; 
wire u2_remHi_136_; 
wire u2_remHi_137_; 
wire u2_remHi_138_; 
wire u2_remHi_139_; 
wire u2_remHi_13_; 
wire u2_remHi_140_; 
wire u2_remHi_141_; 
wire u2_remHi_142_; 
wire u2_remHi_143_; 
wire u2_remHi_144_; 
wire u2_remHi_145_; 
wire u2_remHi_146_; 
wire u2_remHi_147_; 
wire u2_remHi_148_; 
wire u2_remHi_149_; 
wire u2_remHi_14_; 
wire u2_remHi_150_; 
wire u2_remHi_151_; 
wire u2_remHi_152_; 
wire u2_remHi_153_; 
wire u2_remHi_154_; 
wire u2_remHi_155_; 
wire u2_remHi_156_; 
wire u2_remHi_157_; 
wire u2_remHi_158_; 
wire u2_remHi_159_; 
wire u2_remHi_15_; 
wire u2_remHi_160_; 
wire u2_remHi_161_; 
wire u2_remHi_162_; 
wire u2_remHi_163_; 
wire u2_remHi_164_; 
wire u2_remHi_165_; 
wire u2_remHi_166_; 
wire u2_remHi_167_; 
wire u2_remHi_168_; 
wire u2_remHi_169_; 
wire u2_remHi_16_; 
wire u2_remHi_170_; 
wire u2_remHi_171_; 
wire u2_remHi_172_; 
wire u2_remHi_173_; 
wire u2_remHi_174_; 
wire u2_remHi_175_; 
wire u2_remHi_176_; 
wire u2_remHi_177_; 
wire u2_remHi_178_; 
wire u2_remHi_179_; 
wire u2_remHi_17_; 
wire u2_remHi_180_; 
wire u2_remHi_181_; 
wire u2_remHi_182_; 
wire u2_remHi_183_; 
wire u2_remHi_184_; 
wire u2_remHi_185_; 
wire u2_remHi_186_; 
wire u2_remHi_187_; 
wire u2_remHi_188_; 
wire u2_remHi_189_; 
wire u2_remHi_18_; 
wire u2_remHi_190_; 
wire u2_remHi_191_; 
wire u2_remHi_192_; 
wire u2_remHi_193_; 
wire u2_remHi_194_; 
wire u2_remHi_195_; 
wire u2_remHi_196_; 
wire u2_remHi_197_; 
wire u2_remHi_198_; 
wire u2_remHi_199_; 
wire u2_remHi_19_; 
wire u2_remHi_1_; 
wire u2_remHi_200_; 
wire u2_remHi_201_; 
wire u2_remHi_202_; 
wire u2_remHi_203_; 
wire u2_remHi_204_; 
wire u2_remHi_205_; 
wire u2_remHi_206_; 
wire u2_remHi_207_; 
wire u2_remHi_208_; 
wire u2_remHi_209_; 
wire u2_remHi_20_; 
wire u2_remHi_210_; 
wire u2_remHi_211_; 
wire u2_remHi_212_; 
wire u2_remHi_213_; 
wire u2_remHi_214_; 
wire u2_remHi_215_; 
wire u2_remHi_216_; 
wire u2_remHi_217_; 
wire u2_remHi_218_; 
wire u2_remHi_219_; 
wire u2_remHi_21_; 
wire u2_remHi_220_; 
wire u2_remHi_221_; 
wire u2_remHi_222_; 
wire u2_remHi_223_; 
wire u2_remHi_224_; 
wire u2_remHi_225_; 
wire u2_remHi_226_; 
wire u2_remHi_227_; 
wire u2_remHi_228_; 
wire u2_remHi_229_; 
wire u2_remHi_22_; 
wire u2_remHi_230_; 
wire u2_remHi_231_; 
wire u2_remHi_232_; 
wire u2_remHi_233_; 
wire u2_remHi_234_; 
wire u2_remHi_235_; 
wire u2_remHi_236_; 
wire u2_remHi_237_; 
wire u2_remHi_238_; 
wire u2_remHi_239_; 
wire u2_remHi_23_; 
wire u2_remHi_240_; 
wire u2_remHi_241_; 
wire u2_remHi_242_; 
wire u2_remHi_243_; 
wire u2_remHi_244_; 
wire u2_remHi_245_; 
wire u2_remHi_246_; 
wire u2_remHi_247_; 
wire u2_remHi_248_; 
wire u2_remHi_249_; 
wire u2_remHi_24_; 
wire u2_remHi_250_; 
wire u2_remHi_251_; 
wire u2_remHi_252_; 
wire u2_remHi_253_; 
wire u2_remHi_254_; 
wire u2_remHi_255_; 
wire u2_remHi_256_; 
wire u2_remHi_257_; 
wire u2_remHi_258_; 
wire u2_remHi_259_; 
wire u2_remHi_25_; 
wire u2_remHi_260_; 
wire u2_remHi_261_; 
wire u2_remHi_262_; 
wire u2_remHi_263_; 
wire u2_remHi_264_; 
wire u2_remHi_265_; 
wire u2_remHi_266_; 
wire u2_remHi_267_; 
wire u2_remHi_268_; 
wire u2_remHi_269_; 
wire u2_remHi_26_; 
wire u2_remHi_270_; 
wire u2_remHi_271_; 
wire u2_remHi_272_; 
wire u2_remHi_273_; 
wire u2_remHi_274_; 
wire u2_remHi_275_; 
wire u2_remHi_276_; 
wire u2_remHi_277_; 
wire u2_remHi_278_; 
wire u2_remHi_279_; 
wire u2_remHi_27_; 
wire u2_remHi_280_; 
wire u2_remHi_281_; 
wire u2_remHi_282_; 
wire u2_remHi_283_; 
wire u2_remHi_284_; 
wire u2_remHi_285_; 
wire u2_remHi_286_; 
wire u2_remHi_287_; 
wire u2_remHi_288_; 
wire u2_remHi_289_; 
wire u2_remHi_28_; 
wire u2_remHi_290_; 
wire u2_remHi_291_; 
wire u2_remHi_292_; 
wire u2_remHi_293_; 
wire u2_remHi_294_; 
wire u2_remHi_295_; 
wire u2_remHi_296_; 
wire u2_remHi_297_; 
wire u2_remHi_298_; 
wire u2_remHi_299_; 
wire u2_remHi_29_; 
wire u2_remHi_2_; 
wire u2_remHi_300_; 
wire u2_remHi_301_; 
wire u2_remHi_302_; 
wire u2_remHi_303_; 
wire u2_remHi_304_; 
wire u2_remHi_305_; 
wire u2_remHi_306_; 
wire u2_remHi_307_; 
wire u2_remHi_308_; 
wire u2_remHi_309_; 
wire u2_remHi_30_; 
wire u2_remHi_310_; 
wire u2_remHi_311_; 
wire u2_remHi_312_; 
wire u2_remHi_313_; 
wire u2_remHi_314_; 
wire u2_remHi_315_; 
wire u2_remHi_316_; 
wire u2_remHi_317_; 
wire u2_remHi_318_; 
wire u2_remHi_319_; 
wire u2_remHi_31_; 
wire u2_remHi_320_; 
wire u2_remHi_321_; 
wire u2_remHi_322_; 
wire u2_remHi_323_; 
wire u2_remHi_324_; 
wire u2_remHi_325_; 
wire u2_remHi_326_; 
wire u2_remHi_327_; 
wire u2_remHi_328_; 
wire u2_remHi_329_; 
wire u2_remHi_32_; 
wire u2_remHi_330_; 
wire u2_remHi_331_; 
wire u2_remHi_332_; 
wire u2_remHi_333_; 
wire u2_remHi_334_; 
wire u2_remHi_335_; 
wire u2_remHi_336_; 
wire u2_remHi_337_; 
wire u2_remHi_338_; 
wire u2_remHi_339_; 
wire u2_remHi_33_; 
wire u2_remHi_340_; 
wire u2_remHi_341_; 
wire u2_remHi_342_; 
wire u2_remHi_343_; 
wire u2_remHi_344_; 
wire u2_remHi_345_; 
wire u2_remHi_346_; 
wire u2_remHi_347_; 
wire u2_remHi_348_; 
wire u2_remHi_349_; 
wire u2_remHi_34_; 
wire u2_remHi_350_; 
wire u2_remHi_351_; 
wire u2_remHi_352_; 
wire u2_remHi_353_; 
wire u2_remHi_354_; 
wire u2_remHi_355_; 
wire u2_remHi_356_; 
wire u2_remHi_357_; 
wire u2_remHi_358_; 
wire u2_remHi_359_; 
wire u2_remHi_35_; 
wire u2_remHi_360_; 
wire u2_remHi_361_; 
wire u2_remHi_362_; 
wire u2_remHi_363_; 
wire u2_remHi_364_; 
wire u2_remHi_365_; 
wire u2_remHi_366_; 
wire u2_remHi_367_; 
wire u2_remHi_368_; 
wire u2_remHi_369_; 
wire u2_remHi_36_; 
wire u2_remHi_370_; 
wire u2_remHi_371_; 
wire u2_remHi_372_; 
wire u2_remHi_373_; 
wire u2_remHi_374_; 
wire u2_remHi_375_; 
wire u2_remHi_376_; 
wire u2_remHi_377_; 
wire u2_remHi_378_; 
wire u2_remHi_379_; 
wire u2_remHi_37_; 
wire u2_remHi_380_; 
wire u2_remHi_381_; 
wire u2_remHi_382_; 
wire u2_remHi_383_; 
wire u2_remHi_384_; 
wire u2_remHi_385_; 
wire u2_remHi_386_; 
wire u2_remHi_387_; 
wire u2_remHi_388_; 
wire u2_remHi_389_; 
wire u2_remHi_38_; 
wire u2_remHi_390_; 
wire u2_remHi_391_; 
wire u2_remHi_392_; 
wire u2_remHi_393_; 
wire u2_remHi_394_; 
wire u2_remHi_395_; 
wire u2_remHi_396_; 
wire u2_remHi_397_; 
wire u2_remHi_398_; 
wire u2_remHi_399_; 
wire u2_remHi_39_; 
wire u2_remHi_3_; 
wire u2_remHi_400_; 
wire u2_remHi_401_; 
wire u2_remHi_402_; 
wire u2_remHi_403_; 
wire u2_remHi_404_; 
wire u2_remHi_405_; 
wire u2_remHi_406_; 
wire u2_remHi_407_; 
wire u2_remHi_408_; 
wire u2_remHi_409_; 
wire u2_remHi_40_; 
wire u2_remHi_410_; 
wire u2_remHi_411_; 
wire u2_remHi_412_; 
wire u2_remHi_413_; 
wire u2_remHi_414_; 
wire u2_remHi_415_; 
wire u2_remHi_416_; 
wire u2_remHi_417_; 
wire u2_remHi_418_; 
wire u2_remHi_419_; 
wire u2_remHi_41_; 
wire u2_remHi_420_; 
wire u2_remHi_421_; 
wire u2_remHi_422_; 
wire u2_remHi_423_; 
wire u2_remHi_424_; 
wire u2_remHi_425_; 
wire u2_remHi_426_; 
wire u2_remHi_427_; 
wire u2_remHi_428_; 
wire u2_remHi_429_; 
wire u2_remHi_42_; 
wire u2_remHi_430_; 
wire u2_remHi_431_; 
wire u2_remHi_432_; 
wire u2_remHi_433_; 
wire u2_remHi_434_; 
wire u2_remHi_435_; 
wire u2_remHi_436_; 
wire u2_remHi_437_; 
wire u2_remHi_438_; 
wire u2_remHi_439_; 
wire u2_remHi_43_; 
wire u2_remHi_440_; 
wire u2_remHi_441_; 
wire u2_remHi_442_; 
wire u2_remHi_443_; 
wire u2_remHi_444_; 
wire u2_remHi_445_; 
wire u2_remHi_446_; 
wire u2_remHi_447_; 
wire u2_remHi_448_; 
wire u2_remHi_449_; 
wire u2_remHi_44_; 
wire u2_remHi_45_; 
wire u2_remHi_46_; 
wire u2_remHi_47_; 
wire u2_remHi_48_; 
wire u2_remHi_49_; 
wire u2_remHi_4_; 
wire u2_remHi_50_; 
wire u2_remHi_51_; 
wire u2_remHi_52_; 
wire u2_remHi_53_; 
wire u2_remHi_54_; 
wire u2_remHi_55_; 
wire u2_remHi_56_; 
wire u2_remHi_57_; 
wire u2_remHi_58_; 
wire u2_remHi_59_; 
wire u2_remHi_5_; 
wire u2_remHi_60_; 
wire u2_remHi_61_; 
wire u2_remHi_62_; 
wire u2_remHi_63_; 
wire u2_remHi_64_; 
wire u2_remHi_65_; 
wire u2_remHi_66_; 
wire u2_remHi_67_; 
wire u2_remHi_68_; 
wire u2_remHi_69_; 
wire u2_remHi_6_; 
wire u2_remHi_70_; 
wire u2_remHi_71_; 
wire u2_remHi_72_; 
wire u2_remHi_73_; 
wire u2_remHi_74_; 
wire u2_remHi_75_; 
wire u2_remHi_76_; 
wire u2_remHi_77_; 
wire u2_remHi_78_; 
wire u2_remHi_79_; 
wire u2_remHi_7_; 
wire u2_remHi_80_; 
wire u2_remHi_81_; 
wire u2_remHi_82_; 
wire u2_remHi_83_; 
wire u2_remHi_84_; 
wire u2_remHi_85_; 
wire u2_remHi_86_; 
wire u2_remHi_87_; 
wire u2_remHi_88_; 
wire u2_remHi_89_; 
wire u2_remHi_8_; 
wire u2_remHi_90_; 
wire u2_remHi_91_; 
wire u2_remHi_92_; 
wire u2_remHi_93_; 
wire u2_remHi_94_; 
wire u2_remHi_95_; 
wire u2_remHi_96_; 
wire u2_remHi_97_; 
wire u2_remHi_98_; 
wire u2_remHi_99_; 
wire u2_remHi_9_; 
wire u2_remLo_0_; 
wire u2_remLo_100_; 
wire u2_remLo_101_; 
wire u2_remLo_102_; 
wire u2_remLo_103_; 
wire u2_remLo_104_; 
wire u2_remLo_105_; 
wire u2_remLo_106_; 
wire u2_remLo_107_; 
wire u2_remLo_108_; 
wire u2_remLo_109_; 
wire u2_remLo_10_; 
wire u2_remLo_110_; 
wire u2_remLo_111_; 
wire u2_remLo_112_; 
wire u2_remLo_113_; 
wire u2_remLo_114_; 
wire u2_remLo_115_; 
wire u2_remLo_116_; 
wire u2_remLo_117_; 
wire u2_remLo_118_; 
wire u2_remLo_119_; 
wire u2_remLo_11_; 
wire u2_remLo_120_; 
wire u2_remLo_121_; 
wire u2_remLo_122_; 
wire u2_remLo_123_; 
wire u2_remLo_124_; 
wire u2_remLo_125_; 
wire u2_remLo_126_; 
wire u2_remLo_127_; 
wire u2_remLo_128_; 
wire u2_remLo_129_; 
wire u2_remLo_12_; 
wire u2_remLo_130_; 
wire u2_remLo_131_; 
wire u2_remLo_132_; 
wire u2_remLo_133_; 
wire u2_remLo_134_; 
wire u2_remLo_135_; 
wire u2_remLo_136_; 
wire u2_remLo_137_; 
wire u2_remLo_138_; 
wire u2_remLo_139_; 
wire u2_remLo_13_; 
wire u2_remLo_140_; 
wire u2_remLo_141_; 
wire u2_remLo_142_; 
wire u2_remLo_143_; 
wire u2_remLo_144_; 
wire u2_remLo_145_; 
wire u2_remLo_146_; 
wire u2_remLo_147_; 
wire u2_remLo_148_; 
wire u2_remLo_149_; 
wire u2_remLo_14_; 
wire u2_remLo_150_; 
wire u2_remLo_151_; 
wire u2_remLo_152_; 
wire u2_remLo_153_; 
wire u2_remLo_154_; 
wire u2_remLo_155_; 
wire u2_remLo_156_; 
wire u2_remLo_157_; 
wire u2_remLo_158_; 
wire u2_remLo_159_; 
wire u2_remLo_15_; 
wire u2_remLo_160_; 
wire u2_remLo_161_; 
wire u2_remLo_162_; 
wire u2_remLo_163_; 
wire u2_remLo_164_; 
wire u2_remLo_165_; 
wire u2_remLo_166_; 
wire u2_remLo_167_; 
wire u2_remLo_168_; 
wire u2_remLo_169_; 
wire u2_remLo_16_; 
wire u2_remLo_170_; 
wire u2_remLo_171_; 
wire u2_remLo_172_; 
wire u2_remLo_173_; 
wire u2_remLo_174_; 
wire u2_remLo_175_; 
wire u2_remLo_176_; 
wire u2_remLo_177_; 
wire u2_remLo_178_; 
wire u2_remLo_179_; 
wire u2_remLo_17_; 
wire u2_remLo_180_; 
wire u2_remLo_181_; 
wire u2_remLo_182_; 
wire u2_remLo_183_; 
wire u2_remLo_184_; 
wire u2_remLo_185_; 
wire u2_remLo_186_; 
wire u2_remLo_187_; 
wire u2_remLo_188_; 
wire u2_remLo_189_; 
wire u2_remLo_18_; 
wire u2_remLo_190_; 
wire u2_remLo_191_; 
wire u2_remLo_192_; 
wire u2_remLo_193_; 
wire u2_remLo_194_; 
wire u2_remLo_195_; 
wire u2_remLo_196_; 
wire u2_remLo_197_; 
wire u2_remLo_198_; 
wire u2_remLo_199_; 
wire u2_remLo_19_; 
wire u2_remLo_1_; 
wire u2_remLo_200_; 
wire u2_remLo_201_; 
wire u2_remLo_202_; 
wire u2_remLo_203_; 
wire u2_remLo_204_; 
wire u2_remLo_205_; 
wire u2_remLo_206_; 
wire u2_remLo_207_; 
wire u2_remLo_208_; 
wire u2_remLo_209_; 
wire u2_remLo_20_; 
wire u2_remLo_210_; 
wire u2_remLo_211_; 
wire u2_remLo_212_; 
wire u2_remLo_213_; 
wire u2_remLo_214_; 
wire u2_remLo_215_; 
wire u2_remLo_216_; 
wire u2_remLo_217_; 
wire u2_remLo_218_; 
wire u2_remLo_219_; 
wire u2_remLo_21_; 
wire u2_remLo_220_; 
wire u2_remLo_221_; 
wire u2_remLo_222_; 
wire u2_remLo_223_; 
wire u2_remLo_224_; 
wire u2_remLo_225_; 
wire u2_remLo_226_; 
wire u2_remLo_227_; 
wire u2_remLo_228_; 
wire u2_remLo_229_; 
wire u2_remLo_22_; 
wire u2_remLo_230_; 
wire u2_remLo_231_; 
wire u2_remLo_232_; 
wire u2_remLo_233_; 
wire u2_remLo_234_; 
wire u2_remLo_235_; 
wire u2_remLo_236_; 
wire u2_remLo_237_; 
wire u2_remLo_238_; 
wire u2_remLo_239_; 
wire u2_remLo_23_; 
wire u2_remLo_240_; 
wire u2_remLo_241_; 
wire u2_remLo_242_; 
wire u2_remLo_243_; 
wire u2_remLo_244_; 
wire u2_remLo_245_; 
wire u2_remLo_246_; 
wire u2_remLo_247_; 
wire u2_remLo_248_; 
wire u2_remLo_249_; 
wire u2_remLo_24_; 
wire u2_remLo_250_; 
wire u2_remLo_251_; 
wire u2_remLo_252_; 
wire u2_remLo_253_; 
wire u2_remLo_254_; 
wire u2_remLo_255_; 
wire u2_remLo_256_; 
wire u2_remLo_257_; 
wire u2_remLo_258_; 
wire u2_remLo_259_; 
wire u2_remLo_25_; 
wire u2_remLo_260_; 
wire u2_remLo_261_; 
wire u2_remLo_262_; 
wire u2_remLo_263_; 
wire u2_remLo_264_; 
wire u2_remLo_265_; 
wire u2_remLo_266_; 
wire u2_remLo_267_; 
wire u2_remLo_268_; 
wire u2_remLo_269_; 
wire u2_remLo_26_; 
wire u2_remLo_270_; 
wire u2_remLo_271_; 
wire u2_remLo_272_; 
wire u2_remLo_273_; 
wire u2_remLo_274_; 
wire u2_remLo_275_; 
wire u2_remLo_276_; 
wire u2_remLo_277_; 
wire u2_remLo_278_; 
wire u2_remLo_279_; 
wire u2_remLo_27_; 
wire u2_remLo_280_; 
wire u2_remLo_281_; 
wire u2_remLo_282_; 
wire u2_remLo_283_; 
wire u2_remLo_284_; 
wire u2_remLo_285_; 
wire u2_remLo_286_; 
wire u2_remLo_287_; 
wire u2_remLo_288_; 
wire u2_remLo_289_; 
wire u2_remLo_28_; 
wire u2_remLo_290_; 
wire u2_remLo_291_; 
wire u2_remLo_292_; 
wire u2_remLo_293_; 
wire u2_remLo_294_; 
wire u2_remLo_295_; 
wire u2_remLo_296_; 
wire u2_remLo_297_; 
wire u2_remLo_298_; 
wire u2_remLo_299_; 
wire u2_remLo_29_; 
wire u2_remLo_2_; 
wire u2_remLo_300_; 
wire u2_remLo_301_; 
wire u2_remLo_302_; 
wire u2_remLo_303_; 
wire u2_remLo_304_; 
wire u2_remLo_305_; 
wire u2_remLo_306_; 
wire u2_remLo_307_; 
wire u2_remLo_308_; 
wire u2_remLo_309_; 
wire u2_remLo_30_; 
wire u2_remLo_310_; 
wire u2_remLo_311_; 
wire u2_remLo_312_; 
wire u2_remLo_313_; 
wire u2_remLo_314_; 
wire u2_remLo_315_; 
wire u2_remLo_316_; 
wire u2_remLo_317_; 
wire u2_remLo_318_; 
wire u2_remLo_319_; 
wire u2_remLo_31_; 
wire u2_remLo_320_; 
wire u2_remLo_321_; 
wire u2_remLo_322_; 
wire u2_remLo_323_; 
wire u2_remLo_324_; 
wire u2_remLo_325_; 
wire u2_remLo_326_; 
wire u2_remLo_327_; 
wire u2_remLo_328_; 
wire u2_remLo_329_; 
wire u2_remLo_32_; 
wire u2_remLo_330_; 
wire u2_remLo_331_; 
wire u2_remLo_332_; 
wire u2_remLo_333_; 
wire u2_remLo_334_; 
wire u2_remLo_335_; 
wire u2_remLo_336_; 
wire u2_remLo_337_; 
wire u2_remLo_338_; 
wire u2_remLo_339_; 
wire u2_remLo_33_; 
wire u2_remLo_340_; 
wire u2_remLo_341_; 
wire u2_remLo_342_; 
wire u2_remLo_343_; 
wire u2_remLo_344_; 
wire u2_remLo_345_; 
wire u2_remLo_346_; 
wire u2_remLo_347_; 
wire u2_remLo_348_; 
wire u2_remLo_349_; 
wire u2_remLo_34_; 
wire u2_remLo_350_; 
wire u2_remLo_351_; 
wire u2_remLo_352_; 
wire u2_remLo_353_; 
wire u2_remLo_354_; 
wire u2_remLo_355_; 
wire u2_remLo_356_; 
wire u2_remLo_357_; 
wire u2_remLo_358_; 
wire u2_remLo_359_; 
wire u2_remLo_35_; 
wire u2_remLo_360_; 
wire u2_remLo_361_; 
wire u2_remLo_362_; 
wire u2_remLo_363_; 
wire u2_remLo_364_; 
wire u2_remLo_365_; 
wire u2_remLo_366_; 
wire u2_remLo_367_; 
wire u2_remLo_368_; 
wire u2_remLo_369_; 
wire u2_remLo_36_; 
wire u2_remLo_370_; 
wire u2_remLo_371_; 
wire u2_remLo_372_; 
wire u2_remLo_373_; 
wire u2_remLo_374_; 
wire u2_remLo_375_; 
wire u2_remLo_376_; 
wire u2_remLo_377_; 
wire u2_remLo_378_; 
wire u2_remLo_379_; 
wire u2_remLo_37_; 
wire u2_remLo_380_; 
wire u2_remLo_381_; 
wire u2_remLo_382_; 
wire u2_remLo_383_; 
wire u2_remLo_384_; 
wire u2_remLo_385_; 
wire u2_remLo_386_; 
wire u2_remLo_387_; 
wire u2_remLo_388_; 
wire u2_remLo_389_; 
wire u2_remLo_38_; 
wire u2_remLo_390_; 
wire u2_remLo_391_; 
wire u2_remLo_392_; 
wire u2_remLo_393_; 
wire u2_remLo_394_; 
wire u2_remLo_395_; 
wire u2_remLo_396_; 
wire u2_remLo_397_; 
wire u2_remLo_398_; 
wire u2_remLo_399_; 
wire u2_remLo_39_; 
wire u2_remLo_3_; 
wire u2_remLo_400_; 
wire u2_remLo_401_; 
wire u2_remLo_402_; 
wire u2_remLo_403_; 
wire u2_remLo_404_; 
wire u2_remLo_405_; 
wire u2_remLo_406_; 
wire u2_remLo_407_; 
wire u2_remLo_408_; 
wire u2_remLo_409_; 
wire u2_remLo_40_; 
wire u2_remLo_410_; 
wire u2_remLo_411_; 
wire u2_remLo_412_; 
wire u2_remLo_413_; 
wire u2_remLo_414_; 
wire u2_remLo_415_; 
wire u2_remLo_416_; 
wire u2_remLo_417_; 
wire u2_remLo_418_; 
wire u2_remLo_419_; 
wire u2_remLo_41_; 
wire u2_remLo_420_; 
wire u2_remLo_421_; 
wire u2_remLo_422_; 
wire u2_remLo_423_; 
wire u2_remLo_424_; 
wire u2_remLo_425_; 
wire u2_remLo_426_; 
wire u2_remLo_427_; 
wire u2_remLo_428_; 
wire u2_remLo_429_; 
wire u2_remLo_42_; 
wire u2_remLo_430_; 
wire u2_remLo_431_; 
wire u2_remLo_432_; 
wire u2_remLo_433_; 
wire u2_remLo_434_; 
wire u2_remLo_435_; 
wire u2_remLo_436_; 
wire u2_remLo_437_; 
wire u2_remLo_438_; 
wire u2_remLo_439_; 
wire u2_remLo_43_; 
wire u2_remLo_440_; 
wire u2_remLo_441_; 
wire u2_remLo_442_; 
wire u2_remLo_443_; 
wire u2_remLo_444_; 
wire u2_remLo_445_; 
wire u2_remLo_446_; 
wire u2_remLo_447_; 
wire u2_remLo_448_; 
wire u2_remLo_449_; 
wire u2_remLo_44_; 
wire u2_remLo_45_; 
wire u2_remLo_46_; 
wire u2_remLo_47_; 
wire u2_remLo_48_; 
wire u2_remLo_49_; 
wire u2_remLo_4_; 
wire u2_remLo_50_; 
wire u2_remLo_51_; 
wire u2_remLo_52_; 
wire u2_remLo_53_; 
wire u2_remLo_54_; 
wire u2_remLo_55_; 
wire u2_remLo_56_; 
wire u2_remLo_57_; 
wire u2_remLo_58_; 
wire u2_remLo_59_; 
wire u2_remLo_5_; 
wire u2_remLo_60_; 
wire u2_remLo_61_; 
wire u2_remLo_62_; 
wire u2_remLo_63_; 
wire u2_remLo_64_; 
wire u2_remLo_65_; 
wire u2_remLo_66_; 
wire u2_remLo_67_; 
wire u2_remLo_68_; 
wire u2_remLo_69_; 
wire u2_remLo_6_; 
wire u2_remLo_70_; 
wire u2_remLo_71_; 
wire u2_remLo_72_; 
wire u2_remLo_73_; 
wire u2_remLo_74_; 
wire u2_remLo_75_; 
wire u2_remLo_76_; 
wire u2_remLo_77_; 
wire u2_remLo_78_; 
wire u2_remLo_79_; 
wire u2_remLo_7_; 
wire u2_remLo_80_; 
wire u2_remLo_81_; 
wire u2_remLo_82_; 
wire u2_remLo_83_; 
wire u2_remLo_84_; 
wire u2_remLo_85_; 
wire u2_remLo_86_; 
wire u2_remLo_87_; 
wire u2_remLo_88_; 
wire u2_remLo_89_; 
wire u2_remLo_8_; 
wire u2_remLo_90_; 
wire u2_remLo_91_; 
wire u2_remLo_92_; 
wire u2_remLo_93_; 
wire u2_remLo_94_; 
wire u2_remLo_95_; 
wire u2_remLo_96_; 
wire u2_remLo_97_; 
wire u2_remLo_98_; 
wire u2_remLo_99_; 
wire u2_remLo_9_; 
wire u2_root_0_; 
wire u2_state_0_; 
wire u2_state_2_; 
AND2X2 AND2X2_1 ( .A(_abc_73687_new_n753_), .B(sqrto_0_), .Y(\o[36] ));
AND2X2 AND2X2_10 ( .A(_abc_73687_new_n753_), .B(sqrto_9_), .Y(\o[45] ));
AND2X2 AND2X2_100 ( .A(_abc_73687_new_n900_), .B(_abc_73687_new_n899_), .Y(\o[135] ));
AND2X2 AND2X2_1000 ( .A(u2__abc_52155_new_n4022_), .B(sqrto_70_), .Y(u2__abc_52155_new_n4023_));
AND2X2 AND2X2_10000 ( .A(u2__abc_52155_new_n19954_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__74_));
AND2X2 AND2X2_10001 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_74_), .Y(u2__abc_52155_new_n19956_));
AND2X2 AND2X2_10002 ( .A(u2__abc_52155_new_n19946_), .B(sqrto_73_), .Y(u2__abc_52155_new_n19958_));
AND2X2 AND2X2_10003 ( .A(u2__abc_52155_new_n19959_), .B(u2__abc_52155_new_n19957_), .Y(u2__abc_52155_new_n19960_));
AND2X2 AND2X2_10004 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4069_), .Y(u2__abc_52155_new_n19962_));
AND2X2 AND2X2_10005 ( .A(u2__abc_52155_new_n19963_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19964_));
AND2X2 AND2X2_10006 ( .A(u2__abc_52155_new_n19961_), .B(u2__abc_52155_new_n19964_), .Y(u2__abc_52155_new_n19965_));
AND2X2 AND2X2_10007 ( .A(u2__abc_52155_new_n19966_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__75_));
AND2X2 AND2X2_10008 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_75_), .Y(u2__abc_52155_new_n19968_));
AND2X2 AND2X2_10009 ( .A(u2__abc_52155_new_n19958_), .B(sqrto_74_), .Y(u2__abc_52155_new_n19970_));
AND2X2 AND2X2_1001 ( .A(u2__abc_52155_new_n4021_), .B(u2__abc_52155_new_n4024_), .Y(u2__abc_52155_new_n4025_));
AND2X2 AND2X2_10010 ( .A(u2__abc_52155_new_n19971_), .B(u2__abc_52155_new_n19969_), .Y(u2__abc_52155_new_n19972_));
AND2X2 AND2X2_10011 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4062_), .Y(u2__abc_52155_new_n19974_));
AND2X2 AND2X2_10012 ( .A(u2__abc_52155_new_n19975_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19976_));
AND2X2 AND2X2_10013 ( .A(u2__abc_52155_new_n19973_), .B(u2__abc_52155_new_n19976_), .Y(u2__abc_52155_new_n19977_));
AND2X2 AND2X2_10014 ( .A(u2__abc_52155_new_n19978_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__76_));
AND2X2 AND2X2_10015 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_76_), .Y(u2__abc_52155_new_n19980_));
AND2X2 AND2X2_10016 ( .A(u2__abc_52155_new_n19970_), .B(sqrto_75_), .Y(u2__abc_52155_new_n19982_));
AND2X2 AND2X2_10017 ( .A(u2__abc_52155_new_n19983_), .B(u2__abc_52155_new_n19981_), .Y(u2__abc_52155_new_n19984_));
AND2X2 AND2X2_10018 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4047_), .Y(u2__abc_52155_new_n19986_));
AND2X2 AND2X2_10019 ( .A(u2__abc_52155_new_n19987_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19988_));
AND2X2 AND2X2_1002 ( .A(u2__abc_52155_new_n4026_), .B(u2_remHi_71_), .Y(u2__abc_52155_new_n4027_));
AND2X2 AND2X2_10020 ( .A(u2__abc_52155_new_n19985_), .B(u2__abc_52155_new_n19988_), .Y(u2__abc_52155_new_n19989_));
AND2X2 AND2X2_10021 ( .A(u2__abc_52155_new_n19990_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__77_));
AND2X2 AND2X2_10022 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_77_), .Y(u2__abc_52155_new_n19992_));
AND2X2 AND2X2_10023 ( .A(u2__abc_52155_new_n19982_), .B(sqrto_76_), .Y(u2__abc_52155_new_n19994_));
AND2X2 AND2X2_10024 ( .A(u2__abc_52155_new_n19995_), .B(u2__abc_52155_new_n19993_), .Y(u2__abc_52155_new_n19996_));
AND2X2 AND2X2_10025 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4054_), .Y(u2__abc_52155_new_n19998_));
AND2X2 AND2X2_10026 ( .A(u2__abc_52155_new_n19999_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20000_));
AND2X2 AND2X2_10027 ( .A(u2__abc_52155_new_n19997_), .B(u2__abc_52155_new_n20000_), .Y(u2__abc_52155_new_n20001_));
AND2X2 AND2X2_10028 ( .A(u2__abc_52155_new_n20002_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__78_));
AND2X2 AND2X2_10029 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_78_), .Y(u2__abc_52155_new_n20004_));
AND2X2 AND2X2_1003 ( .A(u2__abc_52155_new_n4029_), .B(sqrto_71_), .Y(u2__abc_52155_new_n4030_));
AND2X2 AND2X2_10030 ( .A(u2__abc_52155_new_n19994_), .B(sqrto_77_), .Y(u2__abc_52155_new_n20006_));
AND2X2 AND2X2_10031 ( .A(u2__abc_52155_new_n20007_), .B(u2__abc_52155_new_n20005_), .Y(u2__abc_52155_new_n20008_));
AND2X2 AND2X2_10032 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3958_), .Y(u2__abc_52155_new_n20010_));
AND2X2 AND2X2_10033 ( .A(u2__abc_52155_new_n20011_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20012_));
AND2X2 AND2X2_10034 ( .A(u2__abc_52155_new_n20009_), .B(u2__abc_52155_new_n20012_), .Y(u2__abc_52155_new_n20013_));
AND2X2 AND2X2_10035 ( .A(u2__abc_52155_new_n20014_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__79_));
AND2X2 AND2X2_10036 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_79_), .Y(u2__abc_52155_new_n20016_));
AND2X2 AND2X2_10037 ( .A(u2__abc_52155_new_n20006_), .B(sqrto_78_), .Y(u2__abc_52155_new_n20018_));
AND2X2 AND2X2_10038 ( .A(u2__abc_52155_new_n20019_), .B(u2__abc_52155_new_n20017_), .Y(u2__abc_52155_new_n20020_));
AND2X2 AND2X2_10039 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3965_), .Y(u2__abc_52155_new_n20022_));
AND2X2 AND2X2_1004 ( .A(u2__abc_52155_new_n4028_), .B(u2__abc_52155_new_n4031_), .Y(u2__abc_52155_new_n4032_));
AND2X2 AND2X2_10040 ( .A(u2__abc_52155_new_n20023_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20024_));
AND2X2 AND2X2_10041 ( .A(u2__abc_52155_new_n20021_), .B(u2__abc_52155_new_n20024_), .Y(u2__abc_52155_new_n20025_));
AND2X2 AND2X2_10042 ( .A(u2__abc_52155_new_n20026_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__80_));
AND2X2 AND2X2_10043 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_80_), .Y(u2__abc_52155_new_n20028_));
AND2X2 AND2X2_10044 ( .A(u2__abc_52155_new_n20018_), .B(sqrto_79_), .Y(u2__abc_52155_new_n20029_));
AND2X2 AND2X2_10045 ( .A(u2__abc_52155_new_n20030_), .B(u2__abc_52155_new_n20031_), .Y(u2__abc_52155_new_n20032_));
AND2X2 AND2X2_10046 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3973_), .Y(u2__abc_52155_new_n20034_));
AND2X2 AND2X2_10047 ( .A(u2__abc_52155_new_n20035_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20036_));
AND2X2 AND2X2_10048 ( .A(u2__abc_52155_new_n20033_), .B(u2__abc_52155_new_n20036_), .Y(u2__abc_52155_new_n20037_));
AND2X2 AND2X2_10049 ( .A(u2__abc_52155_new_n20038_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__81_));
AND2X2 AND2X2_1005 ( .A(u2__abc_52155_new_n4025_), .B(u2__abc_52155_new_n4032_), .Y(u2__abc_52155_new_n4033_));
AND2X2 AND2X2_10050 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_81_), .Y(u2__abc_52155_new_n20040_));
AND2X2 AND2X2_10051 ( .A(u2__abc_52155_new_n20029_), .B(sqrto_80_), .Y(u2__abc_52155_new_n20042_));
AND2X2 AND2X2_10052 ( .A(u2__abc_52155_new_n20043_), .B(u2__abc_52155_new_n20041_), .Y(u2__abc_52155_new_n20044_));
AND2X2 AND2X2_10053 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3978_), .Y(u2__abc_52155_new_n20046_));
AND2X2 AND2X2_10054 ( .A(u2__abc_52155_new_n20047_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20048_));
AND2X2 AND2X2_10055 ( .A(u2__abc_52155_new_n20045_), .B(u2__abc_52155_new_n20048_), .Y(u2__abc_52155_new_n20049_));
AND2X2 AND2X2_10056 ( .A(u2__abc_52155_new_n20050_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__82_));
AND2X2 AND2X2_10057 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_82_), .Y(u2__abc_52155_new_n20052_));
AND2X2 AND2X2_10058 ( .A(u2__abc_52155_new_n20042_), .B(sqrto_81_), .Y(u2__abc_52155_new_n20054_));
AND2X2 AND2X2_10059 ( .A(u2__abc_52155_new_n20055_), .B(u2__abc_52155_new_n20053_), .Y(u2__abc_52155_new_n20056_));
AND2X2 AND2X2_1006 ( .A(u2__abc_52155_new_n4034_), .B(u2_remHi_72_), .Y(u2__abc_52155_new_n4035_));
AND2X2 AND2X2_10060 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4008_), .Y(u2__abc_52155_new_n20058_));
AND2X2 AND2X2_10061 ( .A(u2__abc_52155_new_n20059_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20060_));
AND2X2 AND2X2_10062 ( .A(u2__abc_52155_new_n20057_), .B(u2__abc_52155_new_n20060_), .Y(u2__abc_52155_new_n20061_));
AND2X2 AND2X2_10063 ( .A(u2__abc_52155_new_n20062_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__83_));
AND2X2 AND2X2_10064 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_83_), .Y(u2__abc_52155_new_n20064_));
AND2X2 AND2X2_10065 ( .A(u2__abc_52155_new_n20054_), .B(sqrto_82_), .Y(u2__abc_52155_new_n20066_));
AND2X2 AND2X2_10066 ( .A(u2__abc_52155_new_n20067_), .B(u2__abc_52155_new_n20065_), .Y(u2__abc_52155_new_n20068_));
AND2X2 AND2X2_10067 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4001_), .Y(u2__abc_52155_new_n20070_));
AND2X2 AND2X2_10068 ( .A(u2__abc_52155_new_n20071_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20072_));
AND2X2 AND2X2_10069 ( .A(u2__abc_52155_new_n20069_), .B(u2__abc_52155_new_n20072_), .Y(u2__abc_52155_new_n20073_));
AND2X2 AND2X2_1007 ( .A(u2__abc_52155_new_n4036_), .B(sqrto_72_), .Y(u2__abc_52155_new_n4037_));
AND2X2 AND2X2_10070 ( .A(u2__abc_52155_new_n20074_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__84_));
AND2X2 AND2X2_10071 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_84_), .Y(u2__abc_52155_new_n20076_));
AND2X2 AND2X2_10072 ( .A(u2__abc_52155_new_n20066_), .B(sqrto_83_), .Y(u2__abc_52155_new_n20078_));
AND2X2 AND2X2_10073 ( .A(u2__abc_52155_new_n20079_), .B(u2__abc_52155_new_n20077_), .Y(u2__abc_52155_new_n20080_));
AND2X2 AND2X2_10074 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3986_), .Y(u2__abc_52155_new_n20082_));
AND2X2 AND2X2_10075 ( .A(u2__abc_52155_new_n20083_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20084_));
AND2X2 AND2X2_10076 ( .A(u2__abc_52155_new_n20081_), .B(u2__abc_52155_new_n20084_), .Y(u2__abc_52155_new_n20085_));
AND2X2 AND2X2_10077 ( .A(u2__abc_52155_new_n20086_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__85_));
AND2X2 AND2X2_10078 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_85_), .Y(u2__abc_52155_new_n20088_));
AND2X2 AND2X2_10079 ( .A(u2__abc_52155_new_n20078_), .B(sqrto_84_), .Y(u2__abc_52155_new_n20090_));
AND2X2 AND2X2_1008 ( .A(u2__abc_52155_new_n4039_), .B(u2_remHi_73_), .Y(u2__abc_52155_new_n4040_));
AND2X2 AND2X2_10080 ( .A(u2__abc_52155_new_n20091_), .B(u2__abc_52155_new_n20089_), .Y(u2__abc_52155_new_n20092_));
AND2X2 AND2X2_10081 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3993_), .Y(u2__abc_52155_new_n20094_));
AND2X2 AND2X2_10082 ( .A(u2__abc_52155_new_n20095_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20096_));
AND2X2 AND2X2_10083 ( .A(u2__abc_52155_new_n20093_), .B(u2__abc_52155_new_n20096_), .Y(u2__abc_52155_new_n20097_));
AND2X2 AND2X2_10084 ( .A(u2__abc_52155_new_n20098_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__86_));
AND2X2 AND2X2_10085 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_86_), .Y(u2__abc_52155_new_n20100_));
AND2X2 AND2X2_10086 ( .A(u2__abc_52155_new_n20090_), .B(sqrto_85_), .Y(u2__abc_52155_new_n20102_));
AND2X2 AND2X2_10087 ( .A(u2__abc_52155_new_n20103_), .B(u2__abc_52155_new_n20101_), .Y(u2__abc_52155_new_n20104_));
AND2X2 AND2X2_10088 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3948_), .Y(u2__abc_52155_new_n20106_));
AND2X2 AND2X2_10089 ( .A(u2__abc_52155_new_n20107_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20108_));
AND2X2 AND2X2_1009 ( .A(u2__abc_52155_new_n4041_), .B(sqrto_73_), .Y(u2__abc_52155_new_n4042_));
AND2X2 AND2X2_10090 ( .A(u2__abc_52155_new_n20105_), .B(u2__abc_52155_new_n20108_), .Y(u2__abc_52155_new_n20109_));
AND2X2 AND2X2_10091 ( .A(u2__abc_52155_new_n20110_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__87_));
AND2X2 AND2X2_10092 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_87_), .Y(u2__abc_52155_new_n20112_));
AND2X2 AND2X2_10093 ( .A(u2__abc_52155_new_n20102_), .B(sqrto_86_), .Y(u2__abc_52155_new_n20114_));
AND2X2 AND2X2_10094 ( .A(u2__abc_52155_new_n20115_), .B(u2__abc_52155_new_n20113_), .Y(u2__abc_52155_new_n20116_));
AND2X2 AND2X2_10095 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3941_), .Y(u2__abc_52155_new_n20118_));
AND2X2 AND2X2_10096 ( .A(u2__abc_52155_new_n20119_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20120_));
AND2X2 AND2X2_10097 ( .A(u2__abc_52155_new_n20117_), .B(u2__abc_52155_new_n20120_), .Y(u2__abc_52155_new_n20121_));
AND2X2 AND2X2_10098 ( .A(u2__abc_52155_new_n20122_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__88_));
AND2X2 AND2X2_10099 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_88_), .Y(u2__abc_52155_new_n20124_));
AND2X2 AND2X2_101 ( .A(_abc_73687_new_n903_), .B(_abc_73687_new_n902_), .Y(\o[136] ));
AND2X2 AND2X2_1010 ( .A(u2__abc_52155_new_n4045_), .B(u2__abc_52155_new_n4033_), .Y(u2__abc_52155_new_n4046_));
AND2X2 AND2X2_10100 ( .A(u2__abc_52155_new_n20114_), .B(sqrto_87_), .Y(u2__abc_52155_new_n20125_));
AND2X2 AND2X2_10101 ( .A(u2__abc_52155_new_n20126_), .B(u2__abc_52155_new_n20127_), .Y(u2__abc_52155_new_n20128_));
AND2X2 AND2X2_10102 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3926_), .Y(u2__abc_52155_new_n20130_));
AND2X2 AND2X2_10103 ( .A(u2__abc_52155_new_n20131_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20132_));
AND2X2 AND2X2_10104 ( .A(u2__abc_52155_new_n20129_), .B(u2__abc_52155_new_n20132_), .Y(u2__abc_52155_new_n20133_));
AND2X2 AND2X2_10105 ( .A(u2__abc_52155_new_n20134_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__89_));
AND2X2 AND2X2_10106 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_89_), .Y(u2__abc_52155_new_n20136_));
AND2X2 AND2X2_10107 ( .A(u2__abc_52155_new_n20125_), .B(sqrto_88_), .Y(u2__abc_52155_new_n20138_));
AND2X2 AND2X2_10108 ( .A(u2__abc_52155_new_n20139_), .B(u2__abc_52155_new_n20137_), .Y(u2__abc_52155_new_n20140_));
AND2X2 AND2X2_10109 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3933_), .Y(u2__abc_52155_new_n20142_));
AND2X2 AND2X2_1011 ( .A(u2__abc_52155_new_n4047_), .B(u2_remHi_76_), .Y(u2__abc_52155_new_n4048_));
AND2X2 AND2X2_10110 ( .A(u2__abc_52155_new_n20143_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20144_));
AND2X2 AND2X2_10111 ( .A(u2__abc_52155_new_n20141_), .B(u2__abc_52155_new_n20144_), .Y(u2__abc_52155_new_n20145_));
AND2X2 AND2X2_10112 ( .A(u2__abc_52155_new_n20146_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__90_));
AND2X2 AND2X2_10113 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_90_), .Y(u2__abc_52155_new_n20148_));
AND2X2 AND2X2_10114 ( .A(u2__abc_52155_new_n20138_), .B(sqrto_89_), .Y(u2__abc_52155_new_n20150_));
AND2X2 AND2X2_10115 ( .A(u2__abc_52155_new_n20151_), .B(u2__abc_52155_new_n20149_), .Y(u2__abc_52155_new_n20152_));
AND2X2 AND2X2_10116 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3917_), .Y(u2__abc_52155_new_n20154_));
AND2X2 AND2X2_10117 ( .A(u2__abc_52155_new_n20155_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20156_));
AND2X2 AND2X2_10118 ( .A(u2__abc_52155_new_n20153_), .B(u2__abc_52155_new_n20156_), .Y(u2__abc_52155_new_n20157_));
AND2X2 AND2X2_10119 ( .A(u2__abc_52155_new_n20158_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__91_));
AND2X2 AND2X2_1012 ( .A(u2__abc_52155_new_n4050_), .B(sqrto_76_), .Y(u2__abc_52155_new_n4051_));
AND2X2 AND2X2_10120 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_91_), .Y(u2__abc_52155_new_n20160_));
AND2X2 AND2X2_10121 ( .A(u2__abc_52155_new_n20150_), .B(sqrto_90_), .Y(u2__abc_52155_new_n20162_));
AND2X2 AND2X2_10122 ( .A(u2__abc_52155_new_n20163_), .B(u2__abc_52155_new_n20161_), .Y(u2__abc_52155_new_n20164_));
AND2X2 AND2X2_10123 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3910_), .Y(u2__abc_52155_new_n20166_));
AND2X2 AND2X2_10124 ( .A(u2__abc_52155_new_n20167_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20168_));
AND2X2 AND2X2_10125 ( .A(u2__abc_52155_new_n20165_), .B(u2__abc_52155_new_n20168_), .Y(u2__abc_52155_new_n20169_));
AND2X2 AND2X2_10126 ( .A(u2__abc_52155_new_n20170_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__92_));
AND2X2 AND2X2_10127 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_92_), .Y(u2__abc_52155_new_n20172_));
AND2X2 AND2X2_10128 ( .A(u2__abc_52155_new_n20162_), .B(sqrto_91_), .Y(u2__abc_52155_new_n20173_));
AND2X2 AND2X2_10129 ( .A(u2__abc_52155_new_n20174_), .B(u2__abc_52155_new_n20175_), .Y(u2__abc_52155_new_n20176_));
AND2X2 AND2X2_1013 ( .A(u2__abc_52155_new_n4049_), .B(u2__abc_52155_new_n4052_), .Y(u2__abc_52155_new_n4053_));
AND2X2 AND2X2_10130 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3895_), .Y(u2__abc_52155_new_n20178_));
AND2X2 AND2X2_10131 ( .A(u2__abc_52155_new_n20179_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20180_));
AND2X2 AND2X2_10132 ( .A(u2__abc_52155_new_n20177_), .B(u2__abc_52155_new_n20180_), .Y(u2__abc_52155_new_n20181_));
AND2X2 AND2X2_10133 ( .A(u2__abc_52155_new_n20182_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__93_));
AND2X2 AND2X2_10134 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_93_), .Y(u2__abc_52155_new_n20184_));
AND2X2 AND2X2_10135 ( .A(u2__abc_52155_new_n20173_), .B(sqrto_92_), .Y(u2__abc_52155_new_n20186_));
AND2X2 AND2X2_10136 ( .A(u2__abc_52155_new_n20187_), .B(u2__abc_52155_new_n20185_), .Y(u2__abc_52155_new_n20188_));
AND2X2 AND2X2_10137 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3902_), .Y(u2__abc_52155_new_n20190_));
AND2X2 AND2X2_10138 ( .A(u2__abc_52155_new_n20191_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20192_));
AND2X2 AND2X2_10139 ( .A(u2__abc_52155_new_n20189_), .B(u2__abc_52155_new_n20192_), .Y(u2__abc_52155_new_n20193_));
AND2X2 AND2X2_1014 ( .A(u2__abc_52155_new_n4054_), .B(u2_remHi_77_), .Y(u2__abc_52155_new_n4055_));
AND2X2 AND2X2_10140 ( .A(u2__abc_52155_new_n20194_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__94_));
AND2X2 AND2X2_10141 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_94_), .Y(u2__abc_52155_new_n20196_));
AND2X2 AND2X2_10142 ( .A(u2__abc_52155_new_n20186_), .B(sqrto_93_), .Y(u2__abc_52155_new_n20197_));
AND2X2 AND2X2_10143 ( .A(u2__abc_52155_new_n20198_), .B(u2__abc_52155_new_n20199_), .Y(u2__abc_52155_new_n20200_));
AND2X2 AND2X2_10144 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3852_), .Y(u2__abc_52155_new_n20202_));
AND2X2 AND2X2_10145 ( .A(u2__abc_52155_new_n20203_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20204_));
AND2X2 AND2X2_10146 ( .A(u2__abc_52155_new_n20201_), .B(u2__abc_52155_new_n20204_), .Y(u2__abc_52155_new_n20205_));
AND2X2 AND2X2_10147 ( .A(u2__abc_52155_new_n20206_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__95_));
AND2X2 AND2X2_10148 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_95_), .Y(u2__abc_52155_new_n20208_));
AND2X2 AND2X2_10149 ( .A(u2__abc_52155_new_n20197_), .B(sqrto_94_), .Y(u2__abc_52155_new_n20210_));
AND2X2 AND2X2_1015 ( .A(u2__abc_52155_new_n4057_), .B(sqrto_77_), .Y(u2__abc_52155_new_n4058_));
AND2X2 AND2X2_10150 ( .A(u2__abc_52155_new_n20211_), .B(u2__abc_52155_new_n20209_), .Y(u2__abc_52155_new_n20212_));
AND2X2 AND2X2_10151 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3845_), .Y(u2__abc_52155_new_n20214_));
AND2X2 AND2X2_10152 ( .A(u2__abc_52155_new_n20215_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20216_));
AND2X2 AND2X2_10153 ( .A(u2__abc_52155_new_n20213_), .B(u2__abc_52155_new_n20216_), .Y(u2__abc_52155_new_n20217_));
AND2X2 AND2X2_10154 ( .A(u2__abc_52155_new_n20218_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__96_));
AND2X2 AND2X2_10155 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_96_), .Y(u2__abc_52155_new_n20220_));
AND2X2 AND2X2_10156 ( .A(u2__abc_52155_new_n20210_), .B(sqrto_95_), .Y(u2__abc_52155_new_n20222_));
AND2X2 AND2X2_10157 ( .A(u2__abc_52155_new_n20223_), .B(u2__abc_52155_new_n20221_), .Y(u2__abc_52155_new_n20224_));
AND2X2 AND2X2_10158 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3833_), .Y(u2__abc_52155_new_n20226_));
AND2X2 AND2X2_10159 ( .A(u2__abc_52155_new_n20227_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20228_));
AND2X2 AND2X2_1016 ( .A(u2__abc_52155_new_n4056_), .B(u2__abc_52155_new_n4059_), .Y(u2__abc_52155_new_n4060_));
AND2X2 AND2X2_10160 ( .A(u2__abc_52155_new_n20225_), .B(u2__abc_52155_new_n20228_), .Y(u2__abc_52155_new_n20229_));
AND2X2 AND2X2_10161 ( .A(u2__abc_52155_new_n20230_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__97_));
AND2X2 AND2X2_10162 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_97_), .Y(u2__abc_52155_new_n20232_));
AND2X2 AND2X2_10163 ( .A(u2__abc_52155_new_n20222_), .B(sqrto_96_), .Y(u2__abc_52155_new_n20234_));
AND2X2 AND2X2_10164 ( .A(u2__abc_52155_new_n20235_), .B(u2__abc_52155_new_n20233_), .Y(u2__abc_52155_new_n20236_));
AND2X2 AND2X2_10165 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3838_), .Y(u2__abc_52155_new_n20238_));
AND2X2 AND2X2_10166 ( .A(u2__abc_52155_new_n20239_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20240_));
AND2X2 AND2X2_10167 ( .A(u2__abc_52155_new_n20237_), .B(u2__abc_52155_new_n20240_), .Y(u2__abc_52155_new_n20241_));
AND2X2 AND2X2_10168 ( .A(u2__abc_52155_new_n20242_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__98_));
AND2X2 AND2X2_10169 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_98_), .Y(u2__abc_52155_new_n20244_));
AND2X2 AND2X2_1017 ( .A(u2__abc_52155_new_n4053_), .B(u2__abc_52155_new_n4060_), .Y(u2__abc_52155_new_n4061_));
AND2X2 AND2X2_10170 ( .A(u2__abc_52155_new_n20234_), .B(sqrto_97_), .Y(u2__abc_52155_new_n20246_));
AND2X2 AND2X2_10171 ( .A(u2__abc_52155_new_n20247_), .B(u2__abc_52155_new_n20245_), .Y(u2__abc_52155_new_n20248_));
AND2X2 AND2X2_10172 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3883_), .Y(u2__abc_52155_new_n20250_));
AND2X2 AND2X2_10173 ( .A(u2__abc_52155_new_n20251_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20252_));
AND2X2 AND2X2_10174 ( .A(u2__abc_52155_new_n20249_), .B(u2__abc_52155_new_n20252_), .Y(u2__abc_52155_new_n20253_));
AND2X2 AND2X2_10175 ( .A(u2__abc_52155_new_n20254_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__99_));
AND2X2 AND2X2_10176 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_99_), .Y(u2__abc_52155_new_n20256_));
AND2X2 AND2X2_10177 ( .A(u2__abc_52155_new_n20246_), .B(sqrto_98_), .Y(u2__abc_52155_new_n20258_));
AND2X2 AND2X2_10178 ( .A(u2__abc_52155_new_n20259_), .B(u2__abc_52155_new_n20257_), .Y(u2__abc_52155_new_n20260_));
AND2X2 AND2X2_10179 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3876_), .Y(u2__abc_52155_new_n20262_));
AND2X2 AND2X2_1018 ( .A(u2__abc_52155_new_n4062_), .B(u2_remHi_75_), .Y(u2__abc_52155_new_n4063_));
AND2X2 AND2X2_10180 ( .A(u2__abc_52155_new_n20263_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20264_));
AND2X2 AND2X2_10181 ( .A(u2__abc_52155_new_n20261_), .B(u2__abc_52155_new_n20264_), .Y(u2__abc_52155_new_n20265_));
AND2X2 AND2X2_10182 ( .A(u2__abc_52155_new_n20266_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__100_));
AND2X2 AND2X2_10183 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_100_), .Y(u2__abc_52155_new_n20268_));
AND2X2 AND2X2_10184 ( .A(u2__abc_52155_new_n20258_), .B(sqrto_99_), .Y(u2__abc_52155_new_n20270_));
AND2X2 AND2X2_10185 ( .A(u2__abc_52155_new_n20271_), .B(u2__abc_52155_new_n20269_), .Y(u2__abc_52155_new_n20272_));
AND2X2 AND2X2_10186 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3861_), .Y(u2__abc_52155_new_n20274_));
AND2X2 AND2X2_10187 ( .A(u2__abc_52155_new_n20275_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20276_));
AND2X2 AND2X2_10188 ( .A(u2__abc_52155_new_n20273_), .B(u2__abc_52155_new_n20276_), .Y(u2__abc_52155_new_n20277_));
AND2X2 AND2X2_10189 ( .A(u2__abc_52155_new_n20278_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__101_));
AND2X2 AND2X2_1019 ( .A(u2__abc_52155_new_n4065_), .B(sqrto_75_), .Y(u2__abc_52155_new_n4066_));
AND2X2 AND2X2_10190 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_101_), .Y(u2__abc_52155_new_n20280_));
AND2X2 AND2X2_10191 ( .A(u2__abc_52155_new_n20270_), .B(sqrto_100_), .Y(u2__abc_52155_new_n20282_));
AND2X2 AND2X2_10192 ( .A(u2__abc_52155_new_n20283_), .B(u2__abc_52155_new_n20281_), .Y(u2__abc_52155_new_n20284_));
AND2X2 AND2X2_10193 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3868_), .Y(u2__abc_52155_new_n20286_));
AND2X2 AND2X2_10194 ( .A(u2__abc_52155_new_n20287_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20288_));
AND2X2 AND2X2_10195 ( .A(u2__abc_52155_new_n20285_), .B(u2__abc_52155_new_n20288_), .Y(u2__abc_52155_new_n20289_));
AND2X2 AND2X2_10196 ( .A(u2__abc_52155_new_n20290_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__102_));
AND2X2 AND2X2_10197 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_102_), .Y(u2__abc_52155_new_n20292_));
AND2X2 AND2X2_10198 ( .A(u2__abc_52155_new_n20282_), .B(sqrto_101_), .Y(u2__abc_52155_new_n20294_));
AND2X2 AND2X2_10199 ( .A(u2__abc_52155_new_n20295_), .B(u2__abc_52155_new_n20293_), .Y(u2__abc_52155_new_n20296_));
AND2X2 AND2X2_102 ( .A(_abc_73687_new_n906_), .B(_abc_73687_new_n905_), .Y(\o[137] ));
AND2X2 AND2X2_1020 ( .A(u2__abc_52155_new_n4064_), .B(u2__abc_52155_new_n4067_), .Y(u2__abc_52155_new_n4068_));
AND2X2 AND2X2_10200 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3792_), .Y(u2__abc_52155_new_n20298_));
AND2X2 AND2X2_10201 ( .A(u2__abc_52155_new_n20299_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20300_));
AND2X2 AND2X2_10202 ( .A(u2__abc_52155_new_n20297_), .B(u2__abc_52155_new_n20300_), .Y(u2__abc_52155_new_n20301_));
AND2X2 AND2X2_10203 ( .A(u2__abc_52155_new_n20302_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__103_));
AND2X2 AND2X2_10204 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_103_), .Y(u2__abc_52155_new_n20304_));
AND2X2 AND2X2_10205 ( .A(u2__abc_52155_new_n20294_), .B(sqrto_102_), .Y(u2__abc_52155_new_n20306_));
AND2X2 AND2X2_10206 ( .A(u2__abc_52155_new_n20307_), .B(u2__abc_52155_new_n20305_), .Y(u2__abc_52155_new_n20308_));
AND2X2 AND2X2_10207 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3785_), .Y(u2__abc_52155_new_n20310_));
AND2X2 AND2X2_10208 ( .A(u2__abc_52155_new_n20311_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20312_));
AND2X2 AND2X2_10209 ( .A(u2__abc_52155_new_n20309_), .B(u2__abc_52155_new_n20312_), .Y(u2__abc_52155_new_n20313_));
AND2X2 AND2X2_1021 ( .A(u2__abc_52155_new_n4069_), .B(u2_remHi_74_), .Y(u2__abc_52155_new_n4070_));
AND2X2 AND2X2_10210 ( .A(u2__abc_52155_new_n20314_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__104_));
AND2X2 AND2X2_10211 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_104_), .Y(u2__abc_52155_new_n20316_));
AND2X2 AND2X2_10212 ( .A(u2__abc_52155_new_n20306_), .B(sqrto_103_), .Y(u2__abc_52155_new_n20317_));
AND2X2 AND2X2_10213 ( .A(u2__abc_52155_new_n20318_), .B(u2__abc_52155_new_n20319_), .Y(u2__abc_52155_new_n20320_));
AND2X2 AND2X2_10214 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3770_), .Y(u2__abc_52155_new_n20322_));
AND2X2 AND2X2_10215 ( .A(u2__abc_52155_new_n20323_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20324_));
AND2X2 AND2X2_10216 ( .A(u2__abc_52155_new_n20321_), .B(u2__abc_52155_new_n20324_), .Y(u2__abc_52155_new_n20325_));
AND2X2 AND2X2_10217 ( .A(u2__abc_52155_new_n20326_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__105_));
AND2X2 AND2X2_10218 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_105_), .Y(u2__abc_52155_new_n20328_));
AND2X2 AND2X2_10219 ( .A(u2__abc_52155_new_n20317_), .B(sqrto_104_), .Y(u2__abc_52155_new_n20330_));
AND2X2 AND2X2_1022 ( .A(u2__abc_52155_new_n4072_), .B(sqrto_74_), .Y(u2__abc_52155_new_n4073_));
AND2X2 AND2X2_10220 ( .A(u2__abc_52155_new_n20331_), .B(u2__abc_52155_new_n20329_), .Y(u2__abc_52155_new_n20332_));
AND2X2 AND2X2_10221 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3777_), .Y(u2__abc_52155_new_n20334_));
AND2X2 AND2X2_10222 ( .A(u2__abc_52155_new_n20335_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20336_));
AND2X2 AND2X2_10223 ( .A(u2__abc_52155_new_n20333_), .B(u2__abc_52155_new_n20336_), .Y(u2__abc_52155_new_n20337_));
AND2X2 AND2X2_10224 ( .A(u2__abc_52155_new_n20338_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__106_));
AND2X2 AND2X2_10225 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_106_), .Y(u2__abc_52155_new_n20340_));
AND2X2 AND2X2_10226 ( .A(u2__abc_52155_new_n20330_), .B(sqrto_105_), .Y(u2__abc_52155_new_n20342_));
AND2X2 AND2X2_10227 ( .A(u2__abc_52155_new_n20343_), .B(u2__abc_52155_new_n20341_), .Y(u2__abc_52155_new_n20344_));
AND2X2 AND2X2_10228 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3823_), .Y(u2__abc_52155_new_n20346_));
AND2X2 AND2X2_10229 ( .A(u2__abc_52155_new_n20347_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20348_));
AND2X2 AND2X2_1023 ( .A(u2__abc_52155_new_n4071_), .B(u2__abc_52155_new_n4074_), .Y(u2__abc_52155_new_n4075_));
AND2X2 AND2X2_10230 ( .A(u2__abc_52155_new_n20345_), .B(u2__abc_52155_new_n20348_), .Y(u2__abc_52155_new_n20349_));
AND2X2 AND2X2_10231 ( .A(u2__abc_52155_new_n20350_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__107_));
AND2X2 AND2X2_10232 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_107_), .Y(u2__abc_52155_new_n20352_));
AND2X2 AND2X2_10233 ( .A(u2__abc_52155_new_n20342_), .B(sqrto_106_), .Y(u2__abc_52155_new_n20354_));
AND2X2 AND2X2_10234 ( .A(u2__abc_52155_new_n20355_), .B(u2__abc_52155_new_n20353_), .Y(u2__abc_52155_new_n20356_));
AND2X2 AND2X2_10235 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3816_), .Y(u2__abc_52155_new_n20358_));
AND2X2 AND2X2_10236 ( .A(u2__abc_52155_new_n20359_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20360_));
AND2X2 AND2X2_10237 ( .A(u2__abc_52155_new_n20357_), .B(u2__abc_52155_new_n20360_), .Y(u2__abc_52155_new_n20361_));
AND2X2 AND2X2_10238 ( .A(u2__abc_52155_new_n20362_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__108_));
AND2X2 AND2X2_10239 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_108_), .Y(u2__abc_52155_new_n20364_));
AND2X2 AND2X2_1024 ( .A(u2__abc_52155_new_n4068_), .B(u2__abc_52155_new_n4075_), .Y(u2__abc_52155_new_n4076_));
AND2X2 AND2X2_10240 ( .A(u2__abc_52155_new_n20354_), .B(sqrto_107_), .Y(u2__abc_52155_new_n20365_));
AND2X2 AND2X2_10241 ( .A(u2__abc_52155_new_n20366_), .B(u2__abc_52155_new_n20367_), .Y(u2__abc_52155_new_n20368_));
AND2X2 AND2X2_10242 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3801_), .Y(u2__abc_52155_new_n20370_));
AND2X2 AND2X2_10243 ( .A(u2__abc_52155_new_n20371_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20372_));
AND2X2 AND2X2_10244 ( .A(u2__abc_52155_new_n20369_), .B(u2__abc_52155_new_n20372_), .Y(u2__abc_52155_new_n20373_));
AND2X2 AND2X2_10245 ( .A(u2__abc_52155_new_n20374_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__109_));
AND2X2 AND2X2_10246 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_109_), .Y(u2__abc_52155_new_n20376_));
AND2X2 AND2X2_10247 ( .A(u2__abc_52155_new_n20365_), .B(sqrto_108_), .Y(u2__abc_52155_new_n20378_));
AND2X2 AND2X2_10248 ( .A(u2__abc_52155_new_n20379_), .B(u2__abc_52155_new_n20377_), .Y(u2__abc_52155_new_n20380_));
AND2X2 AND2X2_10249 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3808_), .Y(u2__abc_52155_new_n20382_));
AND2X2 AND2X2_1025 ( .A(u2__abc_52155_new_n4061_), .B(u2__abc_52155_new_n4076_), .Y(u2__abc_52155_new_n4077_));
AND2X2 AND2X2_10250 ( .A(u2__abc_52155_new_n20383_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20384_));
AND2X2 AND2X2_10251 ( .A(u2__abc_52155_new_n20381_), .B(u2__abc_52155_new_n20384_), .Y(u2__abc_52155_new_n20385_));
AND2X2 AND2X2_10252 ( .A(u2__abc_52155_new_n20386_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__110_));
AND2X2 AND2X2_10253 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_110_), .Y(u2__abc_52155_new_n20388_));
AND2X2 AND2X2_10254 ( .A(u2__abc_52155_new_n20378_), .B(sqrto_109_), .Y(u2__abc_52155_new_n20389_));
AND2X2 AND2X2_10255 ( .A(u2__abc_52155_new_n20390_), .B(u2__abc_52155_new_n20391_), .Y(u2__abc_52155_new_n20392_));
AND2X2 AND2X2_10256 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3706_), .Y(u2__abc_52155_new_n20394_));
AND2X2 AND2X2_10257 ( .A(u2__abc_52155_new_n20395_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20396_));
AND2X2 AND2X2_10258 ( .A(u2__abc_52155_new_n20393_), .B(u2__abc_52155_new_n20396_), .Y(u2__abc_52155_new_n20397_));
AND2X2 AND2X2_10259 ( .A(u2__abc_52155_new_n20398_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__111_));
AND2X2 AND2X2_1026 ( .A(u2__abc_52155_new_n4046_), .B(u2__abc_52155_new_n4077_), .Y(u2__abc_52155_new_n4078_));
AND2X2 AND2X2_10260 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_111_), .Y(u2__abc_52155_new_n20400_));
AND2X2 AND2X2_10261 ( .A(u2__abc_52155_new_n20389_), .B(sqrto_110_), .Y(u2__abc_52155_new_n20402_));
AND2X2 AND2X2_10262 ( .A(u2__abc_52155_new_n20403_), .B(u2__abc_52155_new_n20401_), .Y(u2__abc_52155_new_n20404_));
AND2X2 AND2X2_10263 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3713_), .Y(u2__abc_52155_new_n20406_));
AND2X2 AND2X2_10264 ( .A(u2__abc_52155_new_n20407_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20408_));
AND2X2 AND2X2_10265 ( .A(u2__abc_52155_new_n20405_), .B(u2__abc_52155_new_n20408_), .Y(u2__abc_52155_new_n20409_));
AND2X2 AND2X2_10266 ( .A(u2__abc_52155_new_n20410_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__112_));
AND2X2 AND2X2_10267 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_112_), .Y(u2__abc_52155_new_n20412_));
AND2X2 AND2X2_10268 ( .A(u2__abc_52155_new_n20402_), .B(sqrto_111_), .Y(u2__abc_52155_new_n20414_));
AND2X2 AND2X2_10269 ( .A(u2__abc_52155_new_n20415_), .B(u2__abc_52155_new_n20413_), .Y(u2__abc_52155_new_n20416_));
AND2X2 AND2X2_1027 ( .A(u2__abc_52155_new_n4079_), .B(u2_remHi_62_), .Y(u2__abc_52155_new_n4080_));
AND2X2 AND2X2_10270 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3721_), .Y(u2__abc_52155_new_n20418_));
AND2X2 AND2X2_10271 ( .A(u2__abc_52155_new_n20419_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20420_));
AND2X2 AND2X2_10272 ( .A(u2__abc_52155_new_n20417_), .B(u2__abc_52155_new_n20420_), .Y(u2__abc_52155_new_n20421_));
AND2X2 AND2X2_10273 ( .A(u2__abc_52155_new_n20422_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__113_));
AND2X2 AND2X2_10274 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_113_), .Y(u2__abc_52155_new_n20424_));
AND2X2 AND2X2_10275 ( .A(u2__abc_52155_new_n20414_), .B(sqrto_112_), .Y(u2__abc_52155_new_n20426_));
AND2X2 AND2X2_10276 ( .A(u2__abc_52155_new_n20427_), .B(u2__abc_52155_new_n20425_), .Y(u2__abc_52155_new_n20428_));
AND2X2 AND2X2_10277 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3728_), .Y(u2__abc_52155_new_n20430_));
AND2X2 AND2X2_10278 ( .A(u2__abc_52155_new_n20431_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20432_));
AND2X2 AND2X2_10279 ( .A(u2__abc_52155_new_n20429_), .B(u2__abc_52155_new_n20432_), .Y(u2__abc_52155_new_n20433_));
AND2X2 AND2X2_1028 ( .A(u2__abc_52155_new_n4081_), .B(u2__abc_52155_new_n4082_), .Y(u2__abc_52155_new_n4083_));
AND2X2 AND2X2_10280 ( .A(u2__abc_52155_new_n20434_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__114_));
AND2X2 AND2X2_10281 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_114_), .Y(u2__abc_52155_new_n20436_));
AND2X2 AND2X2_10282 ( .A(u2__abc_52155_new_n20426_), .B(sqrto_113_), .Y(u2__abc_52155_new_n20438_));
AND2X2 AND2X2_10283 ( .A(u2__abc_52155_new_n20439_), .B(u2__abc_52155_new_n20437_), .Y(u2__abc_52155_new_n20440_));
AND2X2 AND2X2_10284 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3759_), .Y(u2__abc_52155_new_n20442_));
AND2X2 AND2X2_10285 ( .A(u2__abc_52155_new_n20443_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20444_));
AND2X2 AND2X2_10286 ( .A(u2__abc_52155_new_n20441_), .B(u2__abc_52155_new_n20444_), .Y(u2__abc_52155_new_n20445_));
AND2X2 AND2X2_10287 ( .A(u2__abc_52155_new_n20446_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__115_));
AND2X2 AND2X2_10288 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_115_), .Y(u2__abc_52155_new_n20448_));
AND2X2 AND2X2_10289 ( .A(u2__abc_52155_new_n20438_), .B(sqrto_114_), .Y(u2__abc_52155_new_n20450_));
AND2X2 AND2X2_1029 ( .A(u2__abc_52155_new_n4084_), .B(u2_remHi_63_), .Y(u2__abc_52155_new_n4085_));
AND2X2 AND2X2_10290 ( .A(u2__abc_52155_new_n20451_), .B(u2__abc_52155_new_n20449_), .Y(u2__abc_52155_new_n20452_));
AND2X2 AND2X2_10291 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3752_), .Y(u2__abc_52155_new_n20454_));
AND2X2 AND2X2_10292 ( .A(u2__abc_52155_new_n20455_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20456_));
AND2X2 AND2X2_10293 ( .A(u2__abc_52155_new_n20453_), .B(u2__abc_52155_new_n20456_), .Y(u2__abc_52155_new_n20457_));
AND2X2 AND2X2_10294 ( .A(u2__abc_52155_new_n20458_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__116_));
AND2X2 AND2X2_10295 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_116_), .Y(u2__abc_52155_new_n20460_));
AND2X2 AND2X2_10296 ( .A(u2__abc_52155_new_n20450_), .B(sqrto_115_), .Y(u2__abc_52155_new_n20461_));
AND2X2 AND2X2_10297 ( .A(u2__abc_52155_new_n20462_), .B(u2__abc_52155_new_n20463_), .Y(u2__abc_52155_new_n20464_));
AND2X2 AND2X2_10298 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3737_), .Y(u2__abc_52155_new_n20466_));
AND2X2 AND2X2_10299 ( .A(u2__abc_52155_new_n20467_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20468_));
AND2X2 AND2X2_103 ( .A(_abc_73687_new_n909_), .B(_abc_73687_new_n908_), .Y(\o[138] ));
AND2X2 AND2X2_1030 ( .A(u2__abc_52155_new_n4087_), .B(sqrto_63_), .Y(u2__abc_52155_new_n4088_));
AND2X2 AND2X2_10300 ( .A(u2__abc_52155_new_n20465_), .B(u2__abc_52155_new_n20468_), .Y(u2__abc_52155_new_n20469_));
AND2X2 AND2X2_10301 ( .A(u2__abc_52155_new_n20470_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__117_));
AND2X2 AND2X2_10302 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_117_), .Y(u2__abc_52155_new_n20472_));
AND2X2 AND2X2_10303 ( .A(u2__abc_52155_new_n20461_), .B(sqrto_116_), .Y(u2__abc_52155_new_n20474_));
AND2X2 AND2X2_10304 ( .A(u2__abc_52155_new_n20475_), .B(u2__abc_52155_new_n20473_), .Y(u2__abc_52155_new_n20476_));
AND2X2 AND2X2_10305 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3744_), .Y(u2__abc_52155_new_n20478_));
AND2X2 AND2X2_10306 ( .A(u2__abc_52155_new_n20479_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20480_));
AND2X2 AND2X2_10307 ( .A(u2__abc_52155_new_n20477_), .B(u2__abc_52155_new_n20480_), .Y(u2__abc_52155_new_n20481_));
AND2X2 AND2X2_10308 ( .A(u2__abc_52155_new_n20482_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__118_));
AND2X2 AND2X2_10309 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_118_), .Y(u2__abc_52155_new_n20484_));
AND2X2 AND2X2_1031 ( .A(u2__abc_52155_new_n4086_), .B(u2__abc_52155_new_n4089_), .Y(u2__abc_52155_new_n4090_));
AND2X2 AND2X2_10310 ( .A(u2__abc_52155_new_n20474_), .B(sqrto_117_), .Y(u2__abc_52155_new_n20485_));
AND2X2 AND2X2_10311 ( .A(u2__abc_52155_new_n20486_), .B(u2__abc_52155_new_n20487_), .Y(u2__abc_52155_new_n20488_));
AND2X2 AND2X2_10312 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3643_), .Y(u2__abc_52155_new_n20490_));
AND2X2 AND2X2_10313 ( .A(u2__abc_52155_new_n20491_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20492_));
AND2X2 AND2X2_10314 ( .A(u2__abc_52155_new_n20489_), .B(u2__abc_52155_new_n20492_), .Y(u2__abc_52155_new_n20493_));
AND2X2 AND2X2_10315 ( .A(u2__abc_52155_new_n20494_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__119_));
AND2X2 AND2X2_10316 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_119_), .Y(u2__abc_52155_new_n20496_));
AND2X2 AND2X2_10317 ( .A(u2__abc_52155_new_n20485_), .B(sqrto_118_), .Y(u2__abc_52155_new_n20498_));
AND2X2 AND2X2_10318 ( .A(u2__abc_52155_new_n20499_), .B(u2__abc_52155_new_n20497_), .Y(u2__abc_52155_new_n20500_));
AND2X2 AND2X2_10319 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3650_), .Y(u2__abc_52155_new_n20502_));
AND2X2 AND2X2_1032 ( .A(u2__abc_52155_new_n4090_), .B(u2__abc_52155_new_n4083_), .Y(u2__abc_52155_new_n4091_));
AND2X2 AND2X2_10320 ( .A(u2__abc_52155_new_n20503_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20504_));
AND2X2 AND2X2_10321 ( .A(u2__abc_52155_new_n20501_), .B(u2__abc_52155_new_n20504_), .Y(u2__abc_52155_new_n20505_));
AND2X2 AND2X2_10322 ( .A(u2__abc_52155_new_n20506_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__120_));
AND2X2 AND2X2_10323 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_120_), .Y(u2__abc_52155_new_n20508_));
AND2X2 AND2X2_10324 ( .A(u2__abc_52155_new_n20498_), .B(sqrto_119_), .Y(u2__abc_52155_new_n20510_));
AND2X2 AND2X2_10325 ( .A(u2__abc_52155_new_n20511_), .B(u2__abc_52155_new_n20509_), .Y(u2__abc_52155_new_n20512_));
AND2X2 AND2X2_10326 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3658_), .Y(u2__abc_52155_new_n20514_));
AND2X2 AND2X2_10327 ( .A(u2__abc_52155_new_n20515_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20516_));
AND2X2 AND2X2_10328 ( .A(u2__abc_52155_new_n20513_), .B(u2__abc_52155_new_n20516_), .Y(u2__abc_52155_new_n20517_));
AND2X2 AND2X2_10329 ( .A(u2__abc_52155_new_n20518_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__121_));
AND2X2 AND2X2_1033 ( .A(u2__abc_52155_new_n4092_), .B(u2_remHi_64_), .Y(u2__abc_52155_new_n4093_));
AND2X2 AND2X2_10330 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_121_), .Y(u2__abc_52155_new_n20520_));
AND2X2 AND2X2_10331 ( .A(u2__abc_52155_new_n20510_), .B(sqrto_120_), .Y(u2__abc_52155_new_n20522_));
AND2X2 AND2X2_10332 ( .A(u2__abc_52155_new_n20523_), .B(u2__abc_52155_new_n20521_), .Y(u2__abc_52155_new_n20524_));
AND2X2 AND2X2_10333 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3665_), .Y(u2__abc_52155_new_n20526_));
AND2X2 AND2X2_10334 ( .A(u2__abc_52155_new_n20527_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20528_));
AND2X2 AND2X2_10335 ( .A(u2__abc_52155_new_n20525_), .B(u2__abc_52155_new_n20528_), .Y(u2__abc_52155_new_n20529_));
AND2X2 AND2X2_10336 ( .A(u2__abc_52155_new_n20530_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__122_));
AND2X2 AND2X2_10337 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_122_), .Y(u2__abc_52155_new_n20532_));
AND2X2 AND2X2_10338 ( .A(u2__abc_52155_new_n20522_), .B(sqrto_121_), .Y(u2__abc_52155_new_n20533_));
AND2X2 AND2X2_10339 ( .A(u2__abc_52155_new_n20534_), .B(u2__abc_52155_new_n20535_), .Y(u2__abc_52155_new_n20536_));
AND2X2 AND2X2_1034 ( .A(u2__abc_52155_new_n4094_), .B(sqrto_64_), .Y(u2__abc_52155_new_n4095_));
AND2X2 AND2X2_10340 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3696_), .Y(u2__abc_52155_new_n20538_));
AND2X2 AND2X2_10341 ( .A(u2__abc_52155_new_n20539_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20540_));
AND2X2 AND2X2_10342 ( .A(u2__abc_52155_new_n20537_), .B(u2__abc_52155_new_n20540_), .Y(u2__abc_52155_new_n20541_));
AND2X2 AND2X2_10343 ( .A(u2__abc_52155_new_n20542_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__123_));
AND2X2 AND2X2_10344 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_123_), .Y(u2__abc_52155_new_n20544_));
AND2X2 AND2X2_10345 ( .A(u2__abc_52155_new_n20533_), .B(sqrto_122_), .Y(u2__abc_52155_new_n20546_));
AND2X2 AND2X2_10346 ( .A(u2__abc_52155_new_n20547_), .B(u2__abc_52155_new_n20545_), .Y(u2__abc_52155_new_n20548_));
AND2X2 AND2X2_10347 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3689_), .Y(u2__abc_52155_new_n20550_));
AND2X2 AND2X2_10348 ( .A(u2__abc_52155_new_n20551_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20552_));
AND2X2 AND2X2_10349 ( .A(u2__abc_52155_new_n20549_), .B(u2__abc_52155_new_n20552_), .Y(u2__abc_52155_new_n20553_));
AND2X2 AND2X2_1035 ( .A(u2__abc_52155_new_n4097_), .B(u2_remHi_65_), .Y(u2__abc_52155_new_n4098_));
AND2X2 AND2X2_10350 ( .A(u2__abc_52155_new_n20554_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__124_));
AND2X2 AND2X2_10351 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_124_), .Y(u2__abc_52155_new_n20556_));
AND2X2 AND2X2_10352 ( .A(u2__abc_52155_new_n20546_), .B(sqrto_123_), .Y(u2__abc_52155_new_n20558_));
AND2X2 AND2X2_10353 ( .A(u2__abc_52155_new_n20559_), .B(u2__abc_52155_new_n20557_), .Y(u2__abc_52155_new_n20560_));
AND2X2 AND2X2_10354 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3674_), .Y(u2__abc_52155_new_n20562_));
AND2X2 AND2X2_10355 ( .A(u2__abc_52155_new_n20563_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20564_));
AND2X2 AND2X2_10356 ( .A(u2__abc_52155_new_n20561_), .B(u2__abc_52155_new_n20564_), .Y(u2__abc_52155_new_n20565_));
AND2X2 AND2X2_10357 ( .A(u2__abc_52155_new_n20566_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__125_));
AND2X2 AND2X2_10358 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_125_), .Y(u2__abc_52155_new_n20568_));
AND2X2 AND2X2_10359 ( .A(u2__abc_52155_new_n20558_), .B(sqrto_124_), .Y(u2__abc_52155_new_n20570_));
AND2X2 AND2X2_1036 ( .A(u2__abc_52155_new_n4099_), .B(sqrto_65_), .Y(u2__abc_52155_new_n4100_));
AND2X2 AND2X2_10360 ( .A(u2__abc_52155_new_n20571_), .B(u2__abc_52155_new_n20569_), .Y(u2__abc_52155_new_n20572_));
AND2X2 AND2X2_10361 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3684_), .Y(u2__abc_52155_new_n20574_));
AND2X2 AND2X2_10362 ( .A(u2__abc_52155_new_n20575_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20576_));
AND2X2 AND2X2_10363 ( .A(u2__abc_52155_new_n20573_), .B(u2__abc_52155_new_n20576_), .Y(u2__abc_52155_new_n20577_));
AND2X2 AND2X2_10364 ( .A(u2__abc_52155_new_n20578_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__126_));
AND2X2 AND2X2_10365 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_126_), .Y(u2__abc_52155_new_n20580_));
AND2X2 AND2X2_10366 ( .A(u2__abc_52155_new_n20570_), .B(sqrto_125_), .Y(u2__abc_52155_new_n20581_));
AND2X2 AND2X2_10367 ( .A(u2__abc_52155_new_n20582_), .B(u2__abc_52155_new_n20583_), .Y(u2__abc_52155_new_n20584_));
AND2X2 AND2X2_10368 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5233_), .Y(u2__abc_52155_new_n20586_));
AND2X2 AND2X2_10369 ( .A(u2__abc_52155_new_n20587_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20588_));
AND2X2 AND2X2_1037 ( .A(u2__abc_52155_new_n4103_), .B(u2__abc_52155_new_n4091_), .Y(u2__abc_52155_new_n4104_));
AND2X2 AND2X2_10370 ( .A(u2__abc_52155_new_n20585_), .B(u2__abc_52155_new_n20588_), .Y(u2__abc_52155_new_n20589_));
AND2X2 AND2X2_10371 ( .A(u2__abc_52155_new_n20590_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__127_));
AND2X2 AND2X2_10372 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_127_), .Y(u2__abc_52155_new_n20592_));
AND2X2 AND2X2_10373 ( .A(u2__abc_52155_new_n20581_), .B(sqrto_126_), .Y(u2__abc_52155_new_n20594_));
AND2X2 AND2X2_10374 ( .A(u2__abc_52155_new_n20595_), .B(u2__abc_52155_new_n20593_), .Y(u2__abc_52155_new_n20596_));
AND2X2 AND2X2_10375 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5238_), .Y(u2__abc_52155_new_n20598_));
AND2X2 AND2X2_10376 ( .A(u2__abc_52155_new_n20599_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20600_));
AND2X2 AND2X2_10377 ( .A(u2__abc_52155_new_n20597_), .B(u2__abc_52155_new_n20600_), .Y(u2__abc_52155_new_n20601_));
AND2X2 AND2X2_10378 ( .A(u2__abc_52155_new_n20602_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__128_));
AND2X2 AND2X2_10379 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_128_), .Y(u2__abc_52155_new_n20604_));
AND2X2 AND2X2_1038 ( .A(u2__abc_52155_new_n4105_), .B(u2_remHi_68_), .Y(u2__abc_52155_new_n4106_));
AND2X2 AND2X2_10380 ( .A(u2__abc_52155_new_n20594_), .B(sqrto_127_), .Y(u2__abc_52155_new_n20606_));
AND2X2 AND2X2_10381 ( .A(u2__abc_52155_new_n20607_), .B(u2__abc_52155_new_n20605_), .Y(u2__abc_52155_new_n20608_));
AND2X2 AND2X2_10382 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5246_), .Y(u2__abc_52155_new_n20610_));
AND2X2 AND2X2_10383 ( .A(u2__abc_52155_new_n20611_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20612_));
AND2X2 AND2X2_10384 ( .A(u2__abc_52155_new_n20609_), .B(u2__abc_52155_new_n20612_), .Y(u2__abc_52155_new_n20613_));
AND2X2 AND2X2_10385 ( .A(u2__abc_52155_new_n20614_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__129_));
AND2X2 AND2X2_10386 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_129_), .Y(u2__abc_52155_new_n20616_));
AND2X2 AND2X2_10387 ( .A(u2__abc_52155_new_n20606_), .B(sqrto_128_), .Y(u2__abc_52155_new_n20618_));
AND2X2 AND2X2_10388 ( .A(u2__abc_52155_new_n20619_), .B(u2__abc_52155_new_n20617_), .Y(u2__abc_52155_new_n20620_));
AND2X2 AND2X2_10389 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5251_), .Y(u2__abc_52155_new_n20622_));
AND2X2 AND2X2_1039 ( .A(u2__abc_52155_new_n4107_), .B(sqrto_68_), .Y(u2__abc_52155_new_n4108_));
AND2X2 AND2X2_10390 ( .A(u2__abc_52155_new_n20623_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20624_));
AND2X2 AND2X2_10391 ( .A(u2__abc_52155_new_n20621_), .B(u2__abc_52155_new_n20624_), .Y(u2__abc_52155_new_n20625_));
AND2X2 AND2X2_10392 ( .A(u2__abc_52155_new_n20626_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__130_));
AND2X2 AND2X2_10393 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_130_), .Y(u2__abc_52155_new_n20628_));
AND2X2 AND2X2_10394 ( .A(u2__abc_52155_new_n20618_), .B(sqrto_129_), .Y(u2__abc_52155_new_n20630_));
AND2X2 AND2X2_10395 ( .A(u2__abc_52155_new_n20631_), .B(u2__abc_52155_new_n20629_), .Y(u2__abc_52155_new_n20632_));
AND2X2 AND2X2_10396 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5275_), .Y(u2__abc_52155_new_n20634_));
AND2X2 AND2X2_10397 ( .A(u2__abc_52155_new_n20635_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20636_));
AND2X2 AND2X2_10398 ( .A(u2__abc_52155_new_n20633_), .B(u2__abc_52155_new_n20636_), .Y(u2__abc_52155_new_n20637_));
AND2X2 AND2X2_10399 ( .A(u2__abc_52155_new_n20638_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__131_));
AND2X2 AND2X2_104 ( .A(_abc_73687_new_n912_), .B(_abc_73687_new_n911_), .Y(\o[139] ));
AND2X2 AND2X2_1040 ( .A(u2__abc_52155_new_n4110_), .B(u2_remHi_69_), .Y(u2__abc_52155_new_n4111_));
AND2X2 AND2X2_10400 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_131_), .Y(u2__abc_52155_new_n20640_));
AND2X2 AND2X2_10401 ( .A(u2__abc_52155_new_n20630_), .B(sqrto_130_), .Y(u2__abc_52155_new_n20642_));
AND2X2 AND2X2_10402 ( .A(u2__abc_52155_new_n20643_), .B(u2__abc_52155_new_n20641_), .Y(u2__abc_52155_new_n20644_));
AND2X2 AND2X2_10403 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5270_), .Y(u2__abc_52155_new_n20646_));
AND2X2 AND2X2_10404 ( .A(u2__abc_52155_new_n20647_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20648_));
AND2X2 AND2X2_10405 ( .A(u2__abc_52155_new_n20645_), .B(u2__abc_52155_new_n20648_), .Y(u2__abc_52155_new_n20649_));
AND2X2 AND2X2_10406 ( .A(u2__abc_52155_new_n20650_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__132_));
AND2X2 AND2X2_10407 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_132_), .Y(u2__abc_52155_new_n20652_));
AND2X2 AND2X2_10408 ( .A(u2__abc_52155_new_n20642_), .B(sqrto_131_), .Y(u2__abc_52155_new_n20654_));
AND2X2 AND2X2_10409 ( .A(u2__abc_52155_new_n20655_), .B(u2__abc_52155_new_n20653_), .Y(u2__abc_52155_new_n20656_));
AND2X2 AND2X2_1041 ( .A(u2__abc_52155_new_n4112_), .B(sqrto_69_), .Y(u2__abc_52155_new_n4113_));
AND2X2 AND2X2_10410 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5259_), .Y(u2__abc_52155_new_n20658_));
AND2X2 AND2X2_10411 ( .A(u2__abc_52155_new_n20659_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20660_));
AND2X2 AND2X2_10412 ( .A(u2__abc_52155_new_n20657_), .B(u2__abc_52155_new_n20660_), .Y(u2__abc_52155_new_n20661_));
AND2X2 AND2X2_10413 ( .A(u2__abc_52155_new_n20662_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__133_));
AND2X2 AND2X2_10414 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_133_), .Y(u2__abc_52155_new_n20664_));
AND2X2 AND2X2_10415 ( .A(u2__abc_52155_new_n20654_), .B(sqrto_132_), .Y(u2__abc_52155_new_n20666_));
AND2X2 AND2X2_10416 ( .A(u2__abc_52155_new_n20667_), .B(u2__abc_52155_new_n20665_), .Y(u2__abc_52155_new_n20668_));
AND2X2 AND2X2_10417 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5264_), .Y(u2__abc_52155_new_n20670_));
AND2X2 AND2X2_10418 ( .A(u2__abc_52155_new_n20671_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20672_));
AND2X2 AND2X2_10419 ( .A(u2__abc_52155_new_n20669_), .B(u2__abc_52155_new_n20672_), .Y(u2__abc_52155_new_n20673_));
AND2X2 AND2X2_1042 ( .A(u2__abc_52155_new_n4116_), .B(u2_remHi_67_), .Y(u2__abc_52155_new_n4117_));
AND2X2 AND2X2_10420 ( .A(u2__abc_52155_new_n20674_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__134_));
AND2X2 AND2X2_10421 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_134_), .Y(u2__abc_52155_new_n20676_));
AND2X2 AND2X2_10422 ( .A(u2__abc_52155_new_n20666_), .B(sqrto_133_), .Y(u2__abc_52155_new_n20678_));
AND2X2 AND2X2_10423 ( .A(u2__abc_52155_new_n20679_), .B(u2__abc_52155_new_n20677_), .Y(u2__abc_52155_new_n20680_));
AND2X2 AND2X2_10424 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5185_), .Y(u2__abc_52155_new_n20682_));
AND2X2 AND2X2_10425 ( .A(u2__abc_52155_new_n20683_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20684_));
AND2X2 AND2X2_10426 ( .A(u2__abc_52155_new_n20681_), .B(u2__abc_52155_new_n20684_), .Y(u2__abc_52155_new_n20685_));
AND2X2 AND2X2_10427 ( .A(u2__abc_52155_new_n20686_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__135_));
AND2X2 AND2X2_10428 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_135_), .Y(u2__abc_52155_new_n20688_));
AND2X2 AND2X2_10429 ( .A(u2__abc_52155_new_n20678_), .B(sqrto_134_), .Y(u2__abc_52155_new_n20690_));
AND2X2 AND2X2_1043 ( .A(u2__abc_52155_new_n4118_), .B(sqrto_67_), .Y(u2__abc_52155_new_n4119_));
AND2X2 AND2X2_10430 ( .A(u2__abc_52155_new_n20691_), .B(u2__abc_52155_new_n20689_), .Y(u2__abc_52155_new_n20692_));
AND2X2 AND2X2_10431 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5192_), .Y(u2__abc_52155_new_n20694_));
AND2X2 AND2X2_10432 ( .A(u2__abc_52155_new_n20695_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20696_));
AND2X2 AND2X2_10433 ( .A(u2__abc_52155_new_n20693_), .B(u2__abc_52155_new_n20696_), .Y(u2__abc_52155_new_n20697_));
AND2X2 AND2X2_10434 ( .A(u2__abc_52155_new_n20698_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__136_));
AND2X2 AND2X2_10435 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_136_), .Y(u2__abc_52155_new_n20700_));
AND2X2 AND2X2_10436 ( .A(u2__abc_52155_new_n20690_), .B(sqrto_135_), .Y(u2__abc_52155_new_n20701_));
AND2X2 AND2X2_10437 ( .A(u2__abc_52155_new_n20702_), .B(u2__abc_52155_new_n20703_), .Y(u2__abc_52155_new_n20704_));
AND2X2 AND2X2_10438 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5173_), .Y(u2__abc_52155_new_n20706_));
AND2X2 AND2X2_10439 ( .A(u2__abc_52155_new_n20707_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20708_));
AND2X2 AND2X2_1044 ( .A(u2__abc_52155_new_n4121_), .B(u2_remHi_66_), .Y(u2__abc_52155_new_n4122_));
AND2X2 AND2X2_10440 ( .A(u2__abc_52155_new_n20705_), .B(u2__abc_52155_new_n20708_), .Y(u2__abc_52155_new_n20709_));
AND2X2 AND2X2_10441 ( .A(u2__abc_52155_new_n20710_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__137_));
AND2X2 AND2X2_10442 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_137_), .Y(u2__abc_52155_new_n20712_));
AND2X2 AND2X2_10443 ( .A(u2__abc_52155_new_n20701_), .B(sqrto_136_), .Y(u2__abc_52155_new_n20714_));
AND2X2 AND2X2_10444 ( .A(u2__abc_52155_new_n20715_), .B(u2__abc_52155_new_n20713_), .Y(u2__abc_52155_new_n20716_));
AND2X2 AND2X2_10445 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5178_), .Y(u2__abc_52155_new_n20718_));
AND2X2 AND2X2_10446 ( .A(u2__abc_52155_new_n20719_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20720_));
AND2X2 AND2X2_10447 ( .A(u2__abc_52155_new_n20717_), .B(u2__abc_52155_new_n20720_), .Y(u2__abc_52155_new_n20721_));
AND2X2 AND2X2_10448 ( .A(u2__abc_52155_new_n20722_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__138_));
AND2X2 AND2X2_10449 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_138_), .Y(u2__abc_52155_new_n20724_));
AND2X2 AND2X2_1045 ( .A(u2__abc_52155_new_n4123_), .B(sqrto_66_), .Y(u2__abc_52155_new_n4124_));
AND2X2 AND2X2_10450 ( .A(u2__abc_52155_new_n20714_), .B(sqrto_137_), .Y(u2__abc_52155_new_n20726_));
AND2X2 AND2X2_10451 ( .A(u2__abc_52155_new_n20727_), .B(u2__abc_52155_new_n20725_), .Y(u2__abc_52155_new_n20728_));
AND2X2 AND2X2_10452 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5223_), .Y(u2__abc_52155_new_n20730_));
AND2X2 AND2X2_10453 ( .A(u2__abc_52155_new_n20731_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20732_));
AND2X2 AND2X2_10454 ( .A(u2__abc_52155_new_n20729_), .B(u2__abc_52155_new_n20732_), .Y(u2__abc_52155_new_n20733_));
AND2X2 AND2X2_10455 ( .A(u2__abc_52155_new_n20734_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__139_));
AND2X2 AND2X2_10456 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_139_), .Y(u2__abc_52155_new_n20736_));
AND2X2 AND2X2_10457 ( .A(u2__abc_52155_new_n20726_), .B(sqrto_138_), .Y(u2__abc_52155_new_n20738_));
AND2X2 AND2X2_10458 ( .A(u2__abc_52155_new_n20739_), .B(u2__abc_52155_new_n20737_), .Y(u2__abc_52155_new_n20740_));
AND2X2 AND2X2_10459 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5216_), .Y(u2__abc_52155_new_n20742_));
AND2X2 AND2X2_1046 ( .A(u2__abc_52155_new_n4128_), .B(u2__abc_52155_new_n4104_), .Y(u2__abc_52155_new_n4129_));
AND2X2 AND2X2_10460 ( .A(u2__abc_52155_new_n20743_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20744_));
AND2X2 AND2X2_10461 ( .A(u2__abc_52155_new_n20741_), .B(u2__abc_52155_new_n20744_), .Y(u2__abc_52155_new_n20745_));
AND2X2 AND2X2_10462 ( .A(u2__abc_52155_new_n20746_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__140_));
AND2X2 AND2X2_10463 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_140_), .Y(u2__abc_52155_new_n20748_));
AND2X2 AND2X2_10464 ( .A(u2__abc_52155_new_n20738_), .B(sqrto_139_), .Y(u2__abc_52155_new_n20749_));
AND2X2 AND2X2_10465 ( .A(u2__abc_52155_new_n20750_), .B(u2__abc_52155_new_n20751_), .Y(u2__abc_52155_new_n20752_));
AND2X2 AND2X2_10466 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5201_), .Y(u2__abc_52155_new_n20754_));
AND2X2 AND2X2_10467 ( .A(u2__abc_52155_new_n20755_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20756_));
AND2X2 AND2X2_10468 ( .A(u2__abc_52155_new_n20753_), .B(u2__abc_52155_new_n20756_), .Y(u2__abc_52155_new_n20757_));
AND2X2 AND2X2_10469 ( .A(u2__abc_52155_new_n20758_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__141_));
AND2X2 AND2X2_1047 ( .A(u2__abc_52155_new_n4129_), .B(u2__abc_52155_new_n4078_), .Y(u2__abc_52155_new_n4130_));
AND2X2 AND2X2_10470 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_141_), .Y(u2__abc_52155_new_n20760_));
AND2X2 AND2X2_10471 ( .A(u2__abc_52155_new_n20749_), .B(sqrto_140_), .Y(u2__abc_52155_new_n20762_));
AND2X2 AND2X2_10472 ( .A(u2__abc_52155_new_n20763_), .B(u2__abc_52155_new_n20761_), .Y(u2__abc_52155_new_n20764_));
AND2X2 AND2X2_10473 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5208_), .Y(u2__abc_52155_new_n20766_));
AND2X2 AND2X2_10474 ( .A(u2__abc_52155_new_n20767_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20768_));
AND2X2 AND2X2_10475 ( .A(u2__abc_52155_new_n20765_), .B(u2__abc_52155_new_n20768_), .Y(u2__abc_52155_new_n20769_));
AND2X2 AND2X2_10476 ( .A(u2__abc_52155_new_n20770_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__142_));
AND2X2 AND2X2_10477 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_142_), .Y(u2__abc_52155_new_n20772_));
AND2X2 AND2X2_10478 ( .A(u2__abc_52155_new_n20762_), .B(sqrto_141_), .Y(u2__abc_52155_new_n20773_));
AND2X2 AND2X2_10479 ( .A(u2__abc_52155_new_n20774_), .B(u2__abc_52155_new_n20775_), .Y(u2__abc_52155_new_n20776_));
AND2X2 AND2X2_1048 ( .A(u2__abc_52155_new_n4130_), .B(u2__abc_52155_new_n4018_), .Y(u2__abc_52155_new_n4131_));
AND2X2 AND2X2_10480 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5162_), .Y(u2__abc_52155_new_n20778_));
AND2X2 AND2X2_10481 ( .A(u2__abc_52155_new_n20779_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20780_));
AND2X2 AND2X2_10482 ( .A(u2__abc_52155_new_n20777_), .B(u2__abc_52155_new_n20780_), .Y(u2__abc_52155_new_n20781_));
AND2X2 AND2X2_10483 ( .A(u2__abc_52155_new_n20782_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__143_));
AND2X2 AND2X2_10484 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_143_), .Y(u2__abc_52155_new_n20784_));
AND2X2 AND2X2_10485 ( .A(u2__abc_52155_new_n20773_), .B(sqrto_142_), .Y(u2__abc_52155_new_n20786_));
AND2X2 AND2X2_10486 ( .A(u2__abc_52155_new_n20787_), .B(u2__abc_52155_new_n20785_), .Y(u2__abc_52155_new_n20788_));
AND2X2 AND2X2_10487 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5155_), .Y(u2__abc_52155_new_n20790_));
AND2X2 AND2X2_10488 ( .A(u2__abc_52155_new_n20791_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20792_));
AND2X2 AND2X2_10489 ( .A(u2__abc_52155_new_n20789_), .B(u2__abc_52155_new_n20792_), .Y(u2__abc_52155_new_n20793_));
AND2X2 AND2X2_1049 ( .A(u2__abc_52155_new_n4131_), .B(u2__abc_52155_new_n3894_), .Y(u2__abc_52155_new_n4132_));
AND2X2 AND2X2_10490 ( .A(u2__abc_52155_new_n20794_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__144_));
AND2X2 AND2X2_10491 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_144_), .Y(u2__abc_52155_new_n20796_));
AND2X2 AND2X2_10492 ( .A(u2__abc_52155_new_n20786_), .B(sqrto_143_), .Y(u2__abc_52155_new_n20798_));
AND2X2 AND2X2_10493 ( .A(u2__abc_52155_new_n20799_), .B(u2__abc_52155_new_n20797_), .Y(u2__abc_52155_new_n20800_));
AND2X2 AND2X2_10494 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5143_), .Y(u2__abc_52155_new_n20802_));
AND2X2 AND2X2_10495 ( .A(u2__abc_52155_new_n20803_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20804_));
AND2X2 AND2X2_10496 ( .A(u2__abc_52155_new_n20801_), .B(u2__abc_52155_new_n20804_), .Y(u2__abc_52155_new_n20805_));
AND2X2 AND2X2_10497 ( .A(u2__abc_52155_new_n20806_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__145_));
AND2X2 AND2X2_10498 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_145_), .Y(u2__abc_52155_new_n20808_));
AND2X2 AND2X2_10499 ( .A(u2__abc_52155_new_n20798_), .B(sqrto_144_), .Y(u2__abc_52155_new_n20810_));
AND2X2 AND2X2_105 ( .A(_abc_73687_new_n915_), .B(_abc_73687_new_n914_), .Y(\o[140] ));
AND2X2 AND2X2_1050 ( .A(u2__abc_52155_new_n4138_), .B(u2__abc_52155_new_n4089_), .Y(u2__abc_52155_new_n4139_));
AND2X2 AND2X2_10500 ( .A(u2__abc_52155_new_n20811_), .B(u2__abc_52155_new_n20809_), .Y(u2__abc_52155_new_n20812_));
AND2X2 AND2X2_10501 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5148_), .Y(u2__abc_52155_new_n20814_));
AND2X2 AND2X2_10502 ( .A(u2__abc_52155_new_n20815_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20816_));
AND2X2 AND2X2_10503 ( .A(u2__abc_52155_new_n20813_), .B(u2__abc_52155_new_n20816_), .Y(u2__abc_52155_new_n20817_));
AND2X2 AND2X2_10504 ( .A(u2__abc_52155_new_n20818_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__146_));
AND2X2 AND2X2_10505 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_146_), .Y(u2__abc_52155_new_n20820_));
AND2X2 AND2X2_10506 ( .A(u2__abc_52155_new_n20810_), .B(sqrto_145_), .Y(u2__abc_52155_new_n20822_));
AND2X2 AND2X2_10507 ( .A(u2__abc_52155_new_n20823_), .B(u2__abc_52155_new_n20821_), .Y(u2__abc_52155_new_n20824_));
AND2X2 AND2X2_10508 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5134_), .Y(u2__abc_52155_new_n20826_));
AND2X2 AND2X2_10509 ( .A(u2__abc_52155_new_n20827_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20828_));
AND2X2 AND2X2_1051 ( .A(u2__abc_52155_new_n4143_), .B(u2__abc_52155_new_n4141_), .Y(u2__abc_52155_new_n4144_));
AND2X2 AND2X2_10510 ( .A(u2__abc_52155_new_n20825_), .B(u2__abc_52155_new_n20828_), .Y(u2__abc_52155_new_n20829_));
AND2X2 AND2X2_10511 ( .A(u2__abc_52155_new_n20830_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__147_));
AND2X2 AND2X2_10512 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_147_), .Y(u2__abc_52155_new_n20832_));
AND2X2 AND2X2_10513 ( .A(u2__abc_52155_new_n20822_), .B(sqrto_146_), .Y(u2__abc_52155_new_n20834_));
AND2X2 AND2X2_10514 ( .A(u2__abc_52155_new_n20835_), .B(u2__abc_52155_new_n20833_), .Y(u2__abc_52155_new_n20836_));
AND2X2 AND2X2_10515 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5127_), .Y(u2__abc_52155_new_n20838_));
AND2X2 AND2X2_10516 ( .A(u2__abc_52155_new_n20839_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20840_));
AND2X2 AND2X2_10517 ( .A(u2__abc_52155_new_n20837_), .B(u2__abc_52155_new_n20840_), .Y(u2__abc_52155_new_n20841_));
AND2X2 AND2X2_10518 ( .A(u2__abc_52155_new_n20842_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__148_));
AND2X2 AND2X2_10519 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_148_), .Y(u2__abc_52155_new_n20844_));
AND2X2 AND2X2_1052 ( .A(u2__abc_52155_new_n4140_), .B(u2__abc_52155_new_n4144_), .Y(u2__abc_52155_new_n4145_));
AND2X2 AND2X2_10520 ( .A(u2__abc_52155_new_n20834_), .B(sqrto_147_), .Y(u2__abc_52155_new_n20845_));
AND2X2 AND2X2_10521 ( .A(u2__abc_52155_new_n20846_), .B(u2__abc_52155_new_n20847_), .Y(u2__abc_52155_new_n20848_));
AND2X2 AND2X2_10522 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5112_), .Y(u2__abc_52155_new_n20850_));
AND2X2 AND2X2_10523 ( .A(u2__abc_52155_new_n20851_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20852_));
AND2X2 AND2X2_10524 ( .A(u2__abc_52155_new_n20849_), .B(u2__abc_52155_new_n20852_), .Y(u2__abc_52155_new_n20853_));
AND2X2 AND2X2_10525 ( .A(u2__abc_52155_new_n20854_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__149_));
AND2X2 AND2X2_10526 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_149_), .Y(u2__abc_52155_new_n20856_));
AND2X2 AND2X2_10527 ( .A(u2__abc_52155_new_n20845_), .B(sqrto_148_), .Y(u2__abc_52155_new_n20858_));
AND2X2 AND2X2_10528 ( .A(u2__abc_52155_new_n20859_), .B(u2__abc_52155_new_n20857_), .Y(u2__abc_52155_new_n20860_));
AND2X2 AND2X2_10529 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5119_), .Y(u2__abc_52155_new_n20862_));
AND2X2 AND2X2_1053 ( .A(u2__abc_52155_new_n4149_), .B(u2__abc_52155_new_n4147_), .Y(u2__abc_52155_new_n4150_));
AND2X2 AND2X2_10530 ( .A(u2__abc_52155_new_n20863_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20864_));
AND2X2 AND2X2_10531 ( .A(u2__abc_52155_new_n20861_), .B(u2__abc_52155_new_n20864_), .Y(u2__abc_52155_new_n20865_));
AND2X2 AND2X2_10532 ( .A(u2__abc_52155_new_n20866_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__150_));
AND2X2 AND2X2_10533 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_150_), .Y(u2__abc_52155_new_n20868_));
AND2X2 AND2X2_10534 ( .A(u2__abc_52155_new_n20858_), .B(sqrto_149_), .Y(u2__abc_52155_new_n20869_));
AND2X2 AND2X2_10535 ( .A(u2__abc_52155_new_n20870_), .B(u2__abc_52155_new_n20871_), .Y(u2__abc_52155_new_n20872_));
AND2X2 AND2X2_10536 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5071_), .Y(u2__abc_52155_new_n20874_));
AND2X2 AND2X2_10537 ( .A(u2__abc_52155_new_n20875_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20876_));
AND2X2 AND2X2_10538 ( .A(u2__abc_52155_new_n20873_), .B(u2__abc_52155_new_n20876_), .Y(u2__abc_52155_new_n20877_));
AND2X2 AND2X2_10539 ( .A(u2__abc_52155_new_n20878_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__151_));
AND2X2 AND2X2_1054 ( .A(u2__abc_52155_new_n4152_), .B(u2__abc_52155_new_n4108_), .Y(u2__abc_52155_new_n4153_));
AND2X2 AND2X2_10540 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_151_), .Y(u2__abc_52155_new_n20880_));
AND2X2 AND2X2_10541 ( .A(u2__abc_52155_new_n20869_), .B(sqrto_150_), .Y(u2__abc_52155_new_n20882_));
AND2X2 AND2X2_10542 ( .A(u2__abc_52155_new_n20883_), .B(u2__abc_52155_new_n20881_), .Y(u2__abc_52155_new_n20884_));
AND2X2 AND2X2_10543 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5064_), .Y(u2__abc_52155_new_n20886_));
AND2X2 AND2X2_10544 ( .A(u2__abc_52155_new_n20887_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20888_));
AND2X2 AND2X2_10545 ( .A(u2__abc_52155_new_n20885_), .B(u2__abc_52155_new_n20888_), .Y(u2__abc_52155_new_n20889_));
AND2X2 AND2X2_10546 ( .A(u2__abc_52155_new_n20890_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__152_));
AND2X2 AND2X2_10547 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_152_), .Y(u2__abc_52155_new_n20892_));
AND2X2 AND2X2_10548 ( .A(u2__abc_52155_new_n20882_), .B(sqrto_151_), .Y(u2__abc_52155_new_n20894_));
AND2X2 AND2X2_10549 ( .A(u2__abc_52155_new_n20895_), .B(u2__abc_52155_new_n20893_), .Y(u2__abc_52155_new_n20896_));
AND2X2 AND2X2_1055 ( .A(u2__abc_52155_new_n4151_), .B(u2__abc_52155_new_n4155_), .Y(u2__abc_52155_new_n4156_));
AND2X2 AND2X2_10550 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5049_), .Y(u2__abc_52155_new_n20898_));
AND2X2 AND2X2_10551 ( .A(u2__abc_52155_new_n20899_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20900_));
AND2X2 AND2X2_10552 ( .A(u2__abc_52155_new_n20897_), .B(u2__abc_52155_new_n20900_), .Y(u2__abc_52155_new_n20901_));
AND2X2 AND2X2_10553 ( .A(u2__abc_52155_new_n20902_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__153_));
AND2X2 AND2X2_10554 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_153_), .Y(u2__abc_52155_new_n20904_));
AND2X2 AND2X2_10555 ( .A(u2__abc_52155_new_n20894_), .B(sqrto_152_), .Y(u2__abc_52155_new_n20906_));
AND2X2 AND2X2_10556 ( .A(u2__abc_52155_new_n20907_), .B(u2__abc_52155_new_n20905_), .Y(u2__abc_52155_new_n20908_));
AND2X2 AND2X2_10557 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5056_), .Y(u2__abc_52155_new_n20910_));
AND2X2 AND2X2_10558 ( .A(u2__abc_52155_new_n20911_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20912_));
AND2X2 AND2X2_10559 ( .A(u2__abc_52155_new_n20909_), .B(u2__abc_52155_new_n20912_), .Y(u2__abc_52155_new_n20913_));
AND2X2 AND2X2_1056 ( .A(u2__abc_52155_new_n4146_), .B(u2__abc_52155_new_n4156_), .Y(u2__abc_52155_new_n4157_));
AND2X2 AND2X2_10560 ( .A(u2__abc_52155_new_n20914_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__154_));
AND2X2 AND2X2_10561 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_154_), .Y(u2__abc_52155_new_n20916_));
AND2X2 AND2X2_10562 ( .A(u2__abc_52155_new_n20906_), .B(sqrto_153_), .Y(u2__abc_52155_new_n20917_));
AND2X2 AND2X2_10563 ( .A(u2__abc_52155_new_n20918_), .B(u2__abc_52155_new_n20919_), .Y(u2__abc_52155_new_n20920_));
AND2X2 AND2X2_10564 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5102_), .Y(u2__abc_52155_new_n20922_));
AND2X2 AND2X2_10565 ( .A(u2__abc_52155_new_n20923_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20924_));
AND2X2 AND2X2_10566 ( .A(u2__abc_52155_new_n20921_), .B(u2__abc_52155_new_n20924_), .Y(u2__abc_52155_new_n20925_));
AND2X2 AND2X2_10567 ( .A(u2__abc_52155_new_n20926_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__155_));
AND2X2 AND2X2_10568 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_155_), .Y(u2__abc_52155_new_n20928_));
AND2X2 AND2X2_10569 ( .A(u2__abc_52155_new_n20917_), .B(sqrto_154_), .Y(u2__abc_52155_new_n20930_));
AND2X2 AND2X2_1057 ( .A(u2__abc_52155_new_n4160_), .B(u2__abc_52155_new_n4031_), .Y(u2__abc_52155_new_n4161_));
AND2X2 AND2X2_10570 ( .A(u2__abc_52155_new_n20931_), .B(u2__abc_52155_new_n20929_), .Y(u2__abc_52155_new_n20932_));
AND2X2 AND2X2_10571 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5095_), .Y(u2__abc_52155_new_n20934_));
AND2X2 AND2X2_10572 ( .A(u2__abc_52155_new_n20935_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20936_));
AND2X2 AND2X2_10573 ( .A(u2__abc_52155_new_n20933_), .B(u2__abc_52155_new_n20936_), .Y(u2__abc_52155_new_n20937_));
AND2X2 AND2X2_10574 ( .A(u2__abc_52155_new_n20938_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__156_));
AND2X2 AND2X2_10575 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_156_), .Y(u2__abc_52155_new_n20940_));
AND2X2 AND2X2_10576 ( .A(u2__abc_52155_new_n20930_), .B(sqrto_155_), .Y(u2__abc_52155_new_n20942_));
AND2X2 AND2X2_10577 ( .A(u2__abc_52155_new_n20943_), .B(u2__abc_52155_new_n20941_), .Y(u2__abc_52155_new_n20944_));
AND2X2 AND2X2_10578 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5080_), .Y(u2__abc_52155_new_n20946_));
AND2X2 AND2X2_10579 ( .A(u2__abc_52155_new_n20947_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20948_));
AND2X2 AND2X2_1058 ( .A(u2__abc_52155_new_n4163_), .B(u2__abc_52155_new_n4037_), .Y(u2__abc_52155_new_n4164_));
AND2X2 AND2X2_10580 ( .A(u2__abc_52155_new_n20945_), .B(u2__abc_52155_new_n20948_), .Y(u2__abc_52155_new_n20949_));
AND2X2 AND2X2_10581 ( .A(u2__abc_52155_new_n20950_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__157_));
AND2X2 AND2X2_10582 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_157_), .Y(u2__abc_52155_new_n20952_));
AND2X2 AND2X2_10583 ( .A(u2__abc_52155_new_n20942_), .B(sqrto_156_), .Y(u2__abc_52155_new_n20954_));
AND2X2 AND2X2_10584 ( .A(u2__abc_52155_new_n20955_), .B(u2__abc_52155_new_n20953_), .Y(u2__abc_52155_new_n20956_));
AND2X2 AND2X2_10585 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5087_), .Y(u2__abc_52155_new_n20958_));
AND2X2 AND2X2_10586 ( .A(u2__abc_52155_new_n20959_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20960_));
AND2X2 AND2X2_10587 ( .A(u2__abc_52155_new_n20957_), .B(u2__abc_52155_new_n20960_), .Y(u2__abc_52155_new_n20961_));
AND2X2 AND2X2_10588 ( .A(u2__abc_52155_new_n20962_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__158_));
AND2X2 AND2X2_10589 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_158_), .Y(u2__abc_52155_new_n20964_));
AND2X2 AND2X2_1059 ( .A(u2__abc_52155_new_n4162_), .B(u2__abc_52155_new_n4166_), .Y(u2__abc_52155_new_n4167_));
AND2X2 AND2X2_10590 ( .A(u2__abc_52155_new_n20954_), .B(sqrto_157_), .Y(u2__abc_52155_new_n20965_));
AND2X2 AND2X2_10591 ( .A(u2__abc_52155_new_n20966_), .B(u2__abc_52155_new_n20967_), .Y(u2__abc_52155_new_n20968_));
AND2X2 AND2X2_10592 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5006_), .Y(u2__abc_52155_new_n20970_));
AND2X2 AND2X2_10593 ( .A(u2__abc_52155_new_n20971_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20972_));
AND2X2 AND2X2_10594 ( .A(u2__abc_52155_new_n20969_), .B(u2__abc_52155_new_n20972_), .Y(u2__abc_52155_new_n20973_));
AND2X2 AND2X2_10595 ( .A(u2__abc_52155_new_n20974_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__159_));
AND2X2 AND2X2_10596 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_159_), .Y(u2__abc_52155_new_n20976_));
AND2X2 AND2X2_10597 ( .A(u2__abc_52155_new_n20965_), .B(sqrto_158_), .Y(u2__abc_52155_new_n20978_));
AND2X2 AND2X2_10598 ( .A(u2__abc_52155_new_n20979_), .B(u2__abc_52155_new_n20977_), .Y(u2__abc_52155_new_n20980_));
AND2X2 AND2X2_10599 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4999_), .Y(u2__abc_52155_new_n20982_));
AND2X2 AND2X2_106 ( .A(_abc_73687_new_n918_), .B(_abc_73687_new_n917_), .Y(\o[141] ));
AND2X2 AND2X2_1060 ( .A(u2__abc_52155_new_n4064_), .B(u2__abc_52155_new_n4073_), .Y(u2__abc_52155_new_n4169_));
AND2X2 AND2X2_10600 ( .A(u2__abc_52155_new_n20983_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20984_));
AND2X2 AND2X2_10601 ( .A(u2__abc_52155_new_n20981_), .B(u2__abc_52155_new_n20984_), .Y(u2__abc_52155_new_n20985_));
AND2X2 AND2X2_10602 ( .A(u2__abc_52155_new_n20986_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__160_));
AND2X2 AND2X2_10603 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_160_), .Y(u2__abc_52155_new_n20988_));
AND2X2 AND2X2_10604 ( .A(u2__abc_52155_new_n20978_), .B(sqrto_159_), .Y(u2__abc_52155_new_n20990_));
AND2X2 AND2X2_10605 ( .A(u2__abc_52155_new_n20991_), .B(u2__abc_52155_new_n20989_), .Y(u2__abc_52155_new_n20992_));
AND2X2 AND2X2_10606 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4987_), .Y(u2__abc_52155_new_n20994_));
AND2X2 AND2X2_10607 ( .A(u2__abc_52155_new_n20995_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n20996_));
AND2X2 AND2X2_10608 ( .A(u2__abc_52155_new_n20993_), .B(u2__abc_52155_new_n20996_), .Y(u2__abc_52155_new_n20997_));
AND2X2 AND2X2_10609 ( .A(u2__abc_52155_new_n20998_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__161_));
AND2X2 AND2X2_1061 ( .A(u2__abc_52155_new_n4170_), .B(u2__abc_52155_new_n4061_), .Y(u2__abc_52155_new_n4171_));
AND2X2 AND2X2_10610 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_161_), .Y(u2__abc_52155_new_n21000_));
AND2X2 AND2X2_10611 ( .A(u2__abc_52155_new_n20990_), .B(sqrto_160_), .Y(u2__abc_52155_new_n21002_));
AND2X2 AND2X2_10612 ( .A(u2__abc_52155_new_n21003_), .B(u2__abc_52155_new_n21001_), .Y(u2__abc_52155_new_n21004_));
AND2X2 AND2X2_10613 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4992_), .Y(u2__abc_52155_new_n21006_));
AND2X2 AND2X2_10614 ( .A(u2__abc_52155_new_n21007_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21008_));
AND2X2 AND2X2_10615 ( .A(u2__abc_52155_new_n21005_), .B(u2__abc_52155_new_n21008_), .Y(u2__abc_52155_new_n21009_));
AND2X2 AND2X2_10616 ( .A(u2__abc_52155_new_n21010_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__162_));
AND2X2 AND2X2_10617 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_162_), .Y(u2__abc_52155_new_n21012_));
AND2X2 AND2X2_10618 ( .A(u2__abc_52155_new_n21002_), .B(sqrto_161_), .Y(u2__abc_52155_new_n21014_));
AND2X2 AND2X2_10619 ( .A(u2__abc_52155_new_n21015_), .B(u2__abc_52155_new_n21013_), .Y(u2__abc_52155_new_n21016_));
AND2X2 AND2X2_1062 ( .A(u2__abc_52155_new_n4056_), .B(u2__abc_52155_new_n4051_), .Y(u2__abc_52155_new_n4172_));
AND2X2 AND2X2_10620 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5037_), .Y(u2__abc_52155_new_n21018_));
AND2X2 AND2X2_10621 ( .A(u2__abc_52155_new_n21019_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21020_));
AND2X2 AND2X2_10622 ( .A(u2__abc_52155_new_n21017_), .B(u2__abc_52155_new_n21020_), .Y(u2__abc_52155_new_n21021_));
AND2X2 AND2X2_10623 ( .A(u2__abc_52155_new_n21022_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__163_));
AND2X2 AND2X2_10624 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_163_), .Y(u2__abc_52155_new_n21024_));
AND2X2 AND2X2_10625 ( .A(u2__abc_52155_new_n21014_), .B(sqrto_162_), .Y(u2__abc_52155_new_n21026_));
AND2X2 AND2X2_10626 ( .A(u2__abc_52155_new_n21027_), .B(u2__abc_52155_new_n21025_), .Y(u2__abc_52155_new_n21028_));
AND2X2 AND2X2_10627 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5030_), .Y(u2__abc_52155_new_n21030_));
AND2X2 AND2X2_10628 ( .A(u2__abc_52155_new_n21031_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21032_));
AND2X2 AND2X2_10629 ( .A(u2__abc_52155_new_n21029_), .B(u2__abc_52155_new_n21032_), .Y(u2__abc_52155_new_n21033_));
AND2X2 AND2X2_1063 ( .A(u2__abc_52155_new_n4168_), .B(u2__abc_52155_new_n4175_), .Y(u2__abc_52155_new_n4176_));
AND2X2 AND2X2_10630 ( .A(u2__abc_52155_new_n21034_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__164_));
AND2X2 AND2X2_10631 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_164_), .Y(u2__abc_52155_new_n21036_));
AND2X2 AND2X2_10632 ( .A(u2__abc_52155_new_n21026_), .B(sqrto_163_), .Y(u2__abc_52155_new_n21037_));
AND2X2 AND2X2_10633 ( .A(u2__abc_52155_new_n21038_), .B(u2__abc_52155_new_n21039_), .Y(u2__abc_52155_new_n21040_));
AND2X2 AND2X2_10634 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5015_), .Y(u2__abc_52155_new_n21042_));
AND2X2 AND2X2_10635 ( .A(u2__abc_52155_new_n21043_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21044_));
AND2X2 AND2X2_10636 ( .A(u2__abc_52155_new_n21041_), .B(u2__abc_52155_new_n21044_), .Y(u2__abc_52155_new_n21045_));
AND2X2 AND2X2_10637 ( .A(u2__abc_52155_new_n21046_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__165_));
AND2X2 AND2X2_10638 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_165_), .Y(u2__abc_52155_new_n21048_));
AND2X2 AND2X2_10639 ( .A(u2__abc_52155_new_n21037_), .B(sqrto_164_), .Y(u2__abc_52155_new_n21050_));
AND2X2 AND2X2_1064 ( .A(u2__abc_52155_new_n4158_), .B(u2__abc_52155_new_n4176_), .Y(u2__abc_52155_new_n4177_));
AND2X2 AND2X2_10640 ( .A(u2__abc_52155_new_n21051_), .B(u2__abc_52155_new_n21049_), .Y(u2__abc_52155_new_n21052_));
AND2X2 AND2X2_10641 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5022_), .Y(u2__abc_52155_new_n21054_));
AND2X2 AND2X2_10642 ( .A(u2__abc_52155_new_n21055_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21056_));
AND2X2 AND2X2_10643 ( .A(u2__abc_52155_new_n21053_), .B(u2__abc_52155_new_n21056_), .Y(u2__abc_52155_new_n21057_));
AND2X2 AND2X2_10644 ( .A(u2__abc_52155_new_n21058_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__166_));
AND2X2 AND2X2_10645 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_166_), .Y(u2__abc_52155_new_n21060_));
AND2X2 AND2X2_10646 ( .A(u2__abc_52155_new_n21050_), .B(sqrto_165_), .Y(u2__abc_52155_new_n21061_));
AND2X2 AND2X2_10647 ( .A(u2__abc_52155_new_n21062_), .B(u2__abc_52155_new_n21063_), .Y(u2__abc_52155_new_n21064_));
AND2X2 AND2X2_10648 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4977_), .Y(u2__abc_52155_new_n21066_));
AND2X2 AND2X2_10649 ( .A(u2__abc_52155_new_n21067_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21068_));
AND2X2 AND2X2_1065 ( .A(u2__abc_52155_new_n4181_), .B(u2__abc_52155_new_n3970_), .Y(u2__abc_52155_new_n4182_));
AND2X2 AND2X2_10650 ( .A(u2__abc_52155_new_n21065_), .B(u2__abc_52155_new_n21068_), .Y(u2__abc_52155_new_n21069_));
AND2X2 AND2X2_10651 ( .A(u2__abc_52155_new_n21070_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__167_));
AND2X2 AND2X2_10652 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_167_), .Y(u2__abc_52155_new_n21072_));
AND2X2 AND2X2_10653 ( .A(u2__abc_52155_new_n21061_), .B(sqrto_166_), .Y(u2__abc_52155_new_n21074_));
AND2X2 AND2X2_10654 ( .A(u2__abc_52155_new_n21075_), .B(u2__abc_52155_new_n21073_), .Y(u2__abc_52155_new_n21076_));
AND2X2 AND2X2_10655 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4970_), .Y(u2__abc_52155_new_n21078_));
AND2X2 AND2X2_10656 ( .A(u2__abc_52155_new_n21079_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21080_));
AND2X2 AND2X2_10657 ( .A(u2__abc_52155_new_n21077_), .B(u2__abc_52155_new_n21080_), .Y(u2__abc_52155_new_n21081_));
AND2X2 AND2X2_10658 ( .A(u2__abc_52155_new_n21082_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__168_));
AND2X2 AND2X2_10659 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_168_), .Y(u2__abc_52155_new_n21084_));
AND2X2 AND2X2_1066 ( .A(u2__abc_52155_new_n4184_), .B(u2__abc_52155_new_n3976_), .Y(u2__abc_52155_new_n4185_));
AND2X2 AND2X2_10660 ( .A(u2__abc_52155_new_n21074_), .B(sqrto_167_), .Y(u2__abc_52155_new_n21086_));
AND2X2 AND2X2_10661 ( .A(u2__abc_52155_new_n21087_), .B(u2__abc_52155_new_n21085_), .Y(u2__abc_52155_new_n21088_));
AND2X2 AND2X2_10662 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4955_), .Y(u2__abc_52155_new_n21090_));
AND2X2 AND2X2_10663 ( .A(u2__abc_52155_new_n21091_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21092_));
AND2X2 AND2X2_10664 ( .A(u2__abc_52155_new_n21089_), .B(u2__abc_52155_new_n21092_), .Y(u2__abc_52155_new_n21093_));
AND2X2 AND2X2_10665 ( .A(u2__abc_52155_new_n21094_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__169_));
AND2X2 AND2X2_10666 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_169_), .Y(u2__abc_52155_new_n21096_));
AND2X2 AND2X2_10667 ( .A(u2__abc_52155_new_n21086_), .B(sqrto_168_), .Y(u2__abc_52155_new_n21098_));
AND2X2 AND2X2_10668 ( .A(u2__abc_52155_new_n21099_), .B(u2__abc_52155_new_n21097_), .Y(u2__abc_52155_new_n21100_));
AND2X2 AND2X2_10669 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4962_), .Y(u2__abc_52155_new_n21102_));
AND2X2 AND2X2_1067 ( .A(u2__abc_52155_new_n4183_), .B(u2__abc_52155_new_n4187_), .Y(u2__abc_52155_new_n4188_));
AND2X2 AND2X2_10670 ( .A(u2__abc_52155_new_n21103_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21104_));
AND2X2 AND2X2_10671 ( .A(u2__abc_52155_new_n21101_), .B(u2__abc_52155_new_n21104_), .Y(u2__abc_52155_new_n21105_));
AND2X2 AND2X2_10672 ( .A(u2__abc_52155_new_n21106_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__170_));
AND2X2 AND2X2_10673 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_170_), .Y(u2__abc_52155_new_n21108_));
AND2X2 AND2X2_10674 ( .A(u2__abc_52155_new_n21098_), .B(sqrto_169_), .Y(u2__abc_52155_new_n21109_));
AND2X2 AND2X2_10675 ( .A(u2__abc_52155_new_n21110_), .B(u2__abc_52155_new_n21111_), .Y(u2__abc_52155_new_n21112_));
AND2X2 AND2X2_10676 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4946_), .Y(u2__abc_52155_new_n21114_));
AND2X2 AND2X2_10677 ( .A(u2__abc_52155_new_n21115_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21116_));
AND2X2 AND2X2_10678 ( .A(u2__abc_52155_new_n21113_), .B(u2__abc_52155_new_n21116_), .Y(u2__abc_52155_new_n21117_));
AND2X2 AND2X2_10679 ( .A(u2__abc_52155_new_n21118_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__171_));
AND2X2 AND2X2_1068 ( .A(u2__abc_52155_new_n4003_), .B(u2__abc_52155_new_n4012_), .Y(u2__abc_52155_new_n4190_));
AND2X2 AND2X2_10680 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_171_), .Y(u2__abc_52155_new_n21120_));
AND2X2 AND2X2_10681 ( .A(u2__abc_52155_new_n21109_), .B(sqrto_170_), .Y(u2__abc_52155_new_n21122_));
AND2X2 AND2X2_10682 ( .A(u2__abc_52155_new_n21123_), .B(u2__abc_52155_new_n21121_), .Y(u2__abc_52155_new_n21124_));
AND2X2 AND2X2_10683 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4939_), .Y(u2__abc_52155_new_n21126_));
AND2X2 AND2X2_10684 ( .A(u2__abc_52155_new_n21127_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21128_));
AND2X2 AND2X2_10685 ( .A(u2__abc_52155_new_n21125_), .B(u2__abc_52155_new_n21128_), .Y(u2__abc_52155_new_n21129_));
AND2X2 AND2X2_10686 ( .A(u2__abc_52155_new_n21130_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__172_));
AND2X2 AND2X2_10687 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_172_), .Y(u2__abc_52155_new_n21132_));
AND2X2 AND2X2_10688 ( .A(u2__abc_52155_new_n21122_), .B(sqrto_171_), .Y(u2__abc_52155_new_n21134_));
AND2X2 AND2X2_10689 ( .A(u2__abc_52155_new_n21135_), .B(u2__abc_52155_new_n21133_), .Y(u2__abc_52155_new_n21136_));
AND2X2 AND2X2_1069 ( .A(u2__abc_52155_new_n4191_), .B(u2__abc_52155_new_n4000_), .Y(u2__abc_52155_new_n4192_));
AND2X2 AND2X2_10690 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4924_), .Y(u2__abc_52155_new_n21138_));
AND2X2 AND2X2_10691 ( .A(u2__abc_52155_new_n21139_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21140_));
AND2X2 AND2X2_10692 ( .A(u2__abc_52155_new_n21137_), .B(u2__abc_52155_new_n21140_), .Y(u2__abc_52155_new_n21141_));
AND2X2 AND2X2_10693 ( .A(u2__abc_52155_new_n21142_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__173_));
AND2X2 AND2X2_10694 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_173_), .Y(u2__abc_52155_new_n21144_));
AND2X2 AND2X2_10695 ( .A(u2__abc_52155_new_n21134_), .B(sqrto_172_), .Y(u2__abc_52155_new_n21146_));
AND2X2 AND2X2_10696 ( .A(u2__abc_52155_new_n21147_), .B(u2__abc_52155_new_n21145_), .Y(u2__abc_52155_new_n21148_));
AND2X2 AND2X2_10697 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4931_), .Y(u2__abc_52155_new_n21150_));
AND2X2 AND2X2_10698 ( .A(u2__abc_52155_new_n21151_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21152_));
AND2X2 AND2X2_10699 ( .A(u2__abc_52155_new_n21149_), .B(u2__abc_52155_new_n21152_), .Y(u2__abc_52155_new_n21153_));
AND2X2 AND2X2_107 ( .A(_abc_73687_new_n921_), .B(_abc_73687_new_n920_), .Y(\o[142] ));
AND2X2 AND2X2_1070 ( .A(u2__abc_52155_new_n3995_), .B(u2__abc_52155_new_n3990_), .Y(u2__abc_52155_new_n4193_));
AND2X2 AND2X2_10700 ( .A(u2__abc_52155_new_n21154_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__174_));
AND2X2 AND2X2_10701 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_174_), .Y(u2__abc_52155_new_n21156_));
AND2X2 AND2X2_10702 ( .A(u2__abc_52155_new_n21146_), .B(sqrto_173_), .Y(u2__abc_52155_new_n21157_));
AND2X2 AND2X2_10703 ( .A(u2__abc_52155_new_n21158_), .B(u2__abc_52155_new_n21159_), .Y(u2__abc_52155_new_n21160_));
AND2X2 AND2X2_10704 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4906_), .Y(u2__abc_52155_new_n21162_));
AND2X2 AND2X2_10705 ( .A(u2__abc_52155_new_n21163_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21164_));
AND2X2 AND2X2_10706 ( .A(u2__abc_52155_new_n21161_), .B(u2__abc_52155_new_n21164_), .Y(u2__abc_52155_new_n21165_));
AND2X2 AND2X2_10707 ( .A(u2__abc_52155_new_n21166_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__175_));
AND2X2 AND2X2_10708 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_175_), .Y(u2__abc_52155_new_n21168_));
AND2X2 AND2X2_10709 ( .A(u2__abc_52155_new_n21157_), .B(sqrto_174_), .Y(u2__abc_52155_new_n21170_));
AND2X2 AND2X2_1071 ( .A(u2__abc_52155_new_n4189_), .B(u2__abc_52155_new_n4196_), .Y(u2__abc_52155_new_n4197_));
AND2X2 AND2X2_10710 ( .A(u2__abc_52155_new_n21171_), .B(u2__abc_52155_new_n21169_), .Y(u2__abc_52155_new_n21172_));
AND2X2 AND2X2_10711 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4913_), .Y(u2__abc_52155_new_n21174_));
AND2X2 AND2X2_10712 ( .A(u2__abc_52155_new_n21175_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21176_));
AND2X2 AND2X2_10713 ( .A(u2__abc_52155_new_n21173_), .B(u2__abc_52155_new_n21176_), .Y(u2__abc_52155_new_n21177_));
AND2X2 AND2X2_10714 ( .A(u2__abc_52155_new_n21178_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__176_));
AND2X2 AND2X2_10715 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_176_), .Y(u2__abc_52155_new_n21180_));
AND2X2 AND2X2_10716 ( .A(u2__abc_52155_new_n21170_), .B(sqrto_175_), .Y(u2__abc_52155_new_n21182_));
AND2X2 AND2X2_10717 ( .A(u2__abc_52155_new_n21183_), .B(u2__abc_52155_new_n21181_), .Y(u2__abc_52155_new_n21184_));
AND2X2 AND2X2_10718 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4891_), .Y(u2__abc_52155_new_n21186_));
AND2X2 AND2X2_10719 ( .A(u2__abc_52155_new_n21187_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21188_));
AND2X2 AND2X2_1072 ( .A(u2__abc_52155_new_n3943_), .B(u2__abc_52155_new_n3952_), .Y(u2__abc_52155_new_n4199_));
AND2X2 AND2X2_10720 ( .A(u2__abc_52155_new_n21185_), .B(u2__abc_52155_new_n21188_), .Y(u2__abc_52155_new_n21189_));
AND2X2 AND2X2_10721 ( .A(u2__abc_52155_new_n21190_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__177_));
AND2X2 AND2X2_10722 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_177_), .Y(u2__abc_52155_new_n21192_));
AND2X2 AND2X2_10723 ( .A(u2__abc_52155_new_n21182_), .B(sqrto_176_), .Y(u2__abc_52155_new_n21194_));
AND2X2 AND2X2_10724 ( .A(u2__abc_52155_new_n21195_), .B(u2__abc_52155_new_n21193_), .Y(u2__abc_52155_new_n21196_));
AND2X2 AND2X2_10725 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4898_), .Y(u2__abc_52155_new_n21198_));
AND2X2 AND2X2_10726 ( .A(u2__abc_52155_new_n21199_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21200_));
AND2X2 AND2X2_10727 ( .A(u2__abc_52155_new_n21197_), .B(u2__abc_52155_new_n21200_), .Y(u2__abc_52155_new_n21201_));
AND2X2 AND2X2_10728 ( .A(u2__abc_52155_new_n21202_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__178_));
AND2X2 AND2X2_10729 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_178_), .Y(u2__abc_52155_new_n21204_));
AND2X2 AND2X2_1073 ( .A(u2__abc_52155_new_n4200_), .B(u2__abc_52155_new_n3940_), .Y(u2__abc_52155_new_n4201_));
AND2X2 AND2X2_10730 ( .A(u2__abc_52155_new_n21194_), .B(sqrto_177_), .Y(u2__abc_52155_new_n21205_));
AND2X2 AND2X2_10731 ( .A(u2__abc_52155_new_n21206_), .B(u2__abc_52155_new_n21207_), .Y(u2__abc_52155_new_n21208_));
AND2X2 AND2X2_10732 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4882_), .Y(u2__abc_52155_new_n21210_));
AND2X2 AND2X2_10733 ( .A(u2__abc_52155_new_n21211_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21212_));
AND2X2 AND2X2_10734 ( .A(u2__abc_52155_new_n21209_), .B(u2__abc_52155_new_n21212_), .Y(u2__abc_52155_new_n21213_));
AND2X2 AND2X2_10735 ( .A(u2__abc_52155_new_n21214_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__179_));
AND2X2 AND2X2_10736 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_179_), .Y(u2__abc_52155_new_n21216_));
AND2X2 AND2X2_10737 ( .A(u2__abc_52155_new_n21205_), .B(sqrto_178_), .Y(u2__abc_52155_new_n21218_));
AND2X2 AND2X2_10738 ( .A(u2__abc_52155_new_n21219_), .B(u2__abc_52155_new_n21217_), .Y(u2__abc_52155_new_n21220_));
AND2X2 AND2X2_10739 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4875_), .Y(u2__abc_52155_new_n21222_));
AND2X2 AND2X2_1074 ( .A(u2__abc_52155_new_n3935_), .B(u2__abc_52155_new_n3930_), .Y(u2__abc_52155_new_n4202_));
AND2X2 AND2X2_10740 ( .A(u2__abc_52155_new_n21223_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21224_));
AND2X2 AND2X2_10741 ( .A(u2__abc_52155_new_n21221_), .B(u2__abc_52155_new_n21224_), .Y(u2__abc_52155_new_n21225_));
AND2X2 AND2X2_10742 ( .A(u2__abc_52155_new_n21226_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__180_));
AND2X2 AND2X2_10743 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_180_), .Y(u2__abc_52155_new_n21228_));
AND2X2 AND2X2_10744 ( .A(u2__abc_52155_new_n21218_), .B(sqrto_179_), .Y(u2__abc_52155_new_n21230_));
AND2X2 AND2X2_10745 ( .A(u2__abc_52155_new_n21231_), .B(u2__abc_52155_new_n21229_), .Y(u2__abc_52155_new_n21232_));
AND2X2 AND2X2_10746 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4860_), .Y(u2__abc_52155_new_n21234_));
AND2X2 AND2X2_10747 ( .A(u2__abc_52155_new_n21235_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21236_));
AND2X2 AND2X2_10748 ( .A(u2__abc_52155_new_n21233_), .B(u2__abc_52155_new_n21236_), .Y(u2__abc_52155_new_n21237_));
AND2X2 AND2X2_10749 ( .A(u2__abc_52155_new_n21238_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__181_));
AND2X2 AND2X2_1075 ( .A(u2__abc_52155_new_n4204_), .B(u2__abc_52155_new_n3925_), .Y(u2__abc_52155_new_n4205_));
AND2X2 AND2X2_10750 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_181_), .Y(u2__abc_52155_new_n21240_));
AND2X2 AND2X2_10751 ( .A(u2__abc_52155_new_n21230_), .B(sqrto_180_), .Y(u2__abc_52155_new_n21242_));
AND2X2 AND2X2_10752 ( .A(u2__abc_52155_new_n21243_), .B(u2__abc_52155_new_n21241_), .Y(u2__abc_52155_new_n21244_));
AND2X2 AND2X2_10753 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4867_), .Y(u2__abc_52155_new_n21246_));
AND2X2 AND2X2_10754 ( .A(u2__abc_52155_new_n21247_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21248_));
AND2X2 AND2X2_10755 ( .A(u2__abc_52155_new_n21245_), .B(u2__abc_52155_new_n21248_), .Y(u2__abc_52155_new_n21249_));
AND2X2 AND2X2_10756 ( .A(u2__abc_52155_new_n21250_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__182_));
AND2X2 AND2X2_10757 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_182_), .Y(u2__abc_52155_new_n21252_));
AND2X2 AND2X2_10758 ( .A(u2__abc_52155_new_n21242_), .B(sqrto_181_), .Y(u2__abc_52155_new_n21253_));
AND2X2 AND2X2_10759 ( .A(u2__abc_52155_new_n21254_), .B(u2__abc_52155_new_n21255_), .Y(u2__abc_52155_new_n21256_));
AND2X2 AND2X2_1076 ( .A(u2__abc_52155_new_n3912_), .B(u2__abc_52155_new_n3921_), .Y(u2__abc_52155_new_n4206_));
AND2X2 AND2X2_10760 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4797_), .Y(u2__abc_52155_new_n21258_));
AND2X2 AND2X2_10761 ( .A(u2__abc_52155_new_n21259_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21260_));
AND2X2 AND2X2_10762 ( .A(u2__abc_52155_new_n21257_), .B(u2__abc_52155_new_n21260_), .Y(u2__abc_52155_new_n21261_));
AND2X2 AND2X2_10763 ( .A(u2__abc_52155_new_n21262_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__183_));
AND2X2 AND2X2_10764 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_183_), .Y(u2__abc_52155_new_n21264_));
AND2X2 AND2X2_10765 ( .A(u2__abc_52155_new_n21253_), .B(sqrto_182_), .Y(u2__abc_52155_new_n21266_));
AND2X2 AND2X2_10766 ( .A(u2__abc_52155_new_n21267_), .B(u2__abc_52155_new_n21265_), .Y(u2__abc_52155_new_n21268_));
AND2X2 AND2X2_10767 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4804_), .Y(u2__abc_52155_new_n21270_));
AND2X2 AND2X2_10768 ( .A(u2__abc_52155_new_n21271_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21272_));
AND2X2 AND2X2_10769 ( .A(u2__abc_52155_new_n21269_), .B(u2__abc_52155_new_n21272_), .Y(u2__abc_52155_new_n21273_));
AND2X2 AND2X2_1077 ( .A(u2__abc_52155_new_n4207_), .B(u2__abc_52155_new_n3909_), .Y(u2__abc_52155_new_n4208_));
AND2X2 AND2X2_10770 ( .A(u2__abc_52155_new_n21274_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__184_));
AND2X2 AND2X2_10771 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_184_), .Y(u2__abc_52155_new_n21276_));
AND2X2 AND2X2_10772 ( .A(u2__abc_52155_new_n21266_), .B(sqrto_183_), .Y(u2__abc_52155_new_n21278_));
AND2X2 AND2X2_10773 ( .A(u2__abc_52155_new_n21279_), .B(u2__abc_52155_new_n21277_), .Y(u2__abc_52155_new_n21280_));
AND2X2 AND2X2_10774 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4812_), .Y(u2__abc_52155_new_n21282_));
AND2X2 AND2X2_10775 ( .A(u2__abc_52155_new_n21283_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21284_));
AND2X2 AND2X2_10776 ( .A(u2__abc_52155_new_n21281_), .B(u2__abc_52155_new_n21284_), .Y(u2__abc_52155_new_n21285_));
AND2X2 AND2X2_10777 ( .A(u2__abc_52155_new_n21286_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__185_));
AND2X2 AND2X2_10778 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_185_), .Y(u2__abc_52155_new_n21288_));
AND2X2 AND2X2_10779 ( .A(u2__abc_52155_new_n21278_), .B(sqrto_184_), .Y(u2__abc_52155_new_n21290_));
AND2X2 AND2X2_1078 ( .A(u2__abc_52155_new_n3904_), .B(u2__abc_52155_new_n3899_), .Y(u2__abc_52155_new_n4209_));
AND2X2 AND2X2_10780 ( .A(u2__abc_52155_new_n21291_), .B(u2__abc_52155_new_n21289_), .Y(u2__abc_52155_new_n21292_));
AND2X2 AND2X2_10781 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4819_), .Y(u2__abc_52155_new_n21294_));
AND2X2 AND2X2_10782 ( .A(u2__abc_52155_new_n21295_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21296_));
AND2X2 AND2X2_10783 ( .A(u2__abc_52155_new_n21293_), .B(u2__abc_52155_new_n21296_), .Y(u2__abc_52155_new_n21297_));
AND2X2 AND2X2_10784 ( .A(u2__abc_52155_new_n21298_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__186_));
AND2X2 AND2X2_10785 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_186_), .Y(u2__abc_52155_new_n21300_));
AND2X2 AND2X2_10786 ( .A(u2__abc_52155_new_n21290_), .B(sqrto_185_), .Y(u2__abc_52155_new_n21301_));
AND2X2 AND2X2_10787 ( .A(u2__abc_52155_new_n21302_), .B(u2__abc_52155_new_n21303_), .Y(u2__abc_52155_new_n21304_));
AND2X2 AND2X2_10788 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4850_), .Y(u2__abc_52155_new_n21306_));
AND2X2 AND2X2_10789 ( .A(u2__abc_52155_new_n21307_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21308_));
AND2X2 AND2X2_1079 ( .A(u2__abc_52155_new_n4198_), .B(u2__abc_52155_new_n4213_), .Y(u2__abc_52155_new_n4214_));
AND2X2 AND2X2_10790 ( .A(u2__abc_52155_new_n21305_), .B(u2__abc_52155_new_n21308_), .Y(u2__abc_52155_new_n21309_));
AND2X2 AND2X2_10791 ( .A(u2__abc_52155_new_n21310_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__187_));
AND2X2 AND2X2_10792 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_187_), .Y(u2__abc_52155_new_n21312_));
AND2X2 AND2X2_10793 ( .A(u2__abc_52155_new_n21301_), .B(sqrto_186_), .Y(u2__abc_52155_new_n21314_));
AND2X2 AND2X2_10794 ( .A(u2__abc_52155_new_n21315_), .B(u2__abc_52155_new_n21313_), .Y(u2__abc_52155_new_n21316_));
AND2X2 AND2X2_10795 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4843_), .Y(u2__abc_52155_new_n21318_));
AND2X2 AND2X2_10796 ( .A(u2__abc_52155_new_n21319_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21320_));
AND2X2 AND2X2_10797 ( .A(u2__abc_52155_new_n21317_), .B(u2__abc_52155_new_n21320_), .Y(u2__abc_52155_new_n21321_));
AND2X2 AND2X2_10798 ( .A(u2__abc_52155_new_n21322_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__188_));
AND2X2 AND2X2_10799 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_188_), .Y(u2__abc_52155_new_n21324_));
AND2X2 AND2X2_108 ( .A(_abc_73687_new_n924_), .B(_abc_73687_new_n923_), .Y(\o[143] ));
AND2X2 AND2X2_1080 ( .A(u2__abc_52155_new_n4178_), .B(u2__abc_52155_new_n4214_), .Y(u2__abc_52155_new_n4215_));
AND2X2 AND2X2_10800 ( .A(u2__abc_52155_new_n21314_), .B(sqrto_187_), .Y(u2__abc_52155_new_n21326_));
AND2X2 AND2X2_10801 ( .A(u2__abc_52155_new_n21327_), .B(u2__abc_52155_new_n21325_), .Y(u2__abc_52155_new_n21328_));
AND2X2 AND2X2_10802 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4828_), .Y(u2__abc_52155_new_n21330_));
AND2X2 AND2X2_10803 ( .A(u2__abc_52155_new_n21331_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21332_));
AND2X2 AND2X2_10804 ( .A(u2__abc_52155_new_n21329_), .B(u2__abc_52155_new_n21332_), .Y(u2__abc_52155_new_n21333_));
AND2X2 AND2X2_10805 ( .A(u2__abc_52155_new_n21334_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__189_));
AND2X2 AND2X2_10806 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_189_), .Y(u2__abc_52155_new_n21336_));
AND2X2 AND2X2_10807 ( .A(u2__abc_52155_new_n21326_), .B(sqrto_188_), .Y(u2__abc_52155_new_n21338_));
AND2X2 AND2X2_10808 ( .A(u2__abc_52155_new_n21339_), .B(u2__abc_52155_new_n21337_), .Y(u2__abc_52155_new_n21340_));
AND2X2 AND2X2_10809 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4835_), .Y(u2__abc_52155_new_n21342_));
AND2X2 AND2X2_1081 ( .A(u2__abc_52155_new_n4220_), .B(u2__abc_52155_new_n3850_), .Y(u2__abc_52155_new_n4221_));
AND2X2 AND2X2_10810 ( .A(u2__abc_52155_new_n21343_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21344_));
AND2X2 AND2X2_10811 ( .A(u2__abc_52155_new_n21341_), .B(u2__abc_52155_new_n21344_), .Y(u2__abc_52155_new_n21345_));
AND2X2 AND2X2_10812 ( .A(u2__abc_52155_new_n21346_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__190_));
AND2X2 AND2X2_10813 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_190_), .Y(u2__abc_52155_new_n21348_));
AND2X2 AND2X2_10814 ( .A(u2__abc_52155_new_n21338_), .B(sqrto_189_), .Y(u2__abc_52155_new_n21349_));
AND2X2 AND2X2_10815 ( .A(u2__abc_52155_new_n21350_), .B(u2__abc_52155_new_n21351_), .Y(u2__abc_52155_new_n21352_));
AND2X2 AND2X2_10816 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4777_), .Y(u2__abc_52155_new_n21354_));
AND2X2 AND2X2_10817 ( .A(u2__abc_52155_new_n21355_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21356_));
AND2X2 AND2X2_10818 ( .A(u2__abc_52155_new_n21353_), .B(u2__abc_52155_new_n21356_), .Y(u2__abc_52155_new_n21357_));
AND2X2 AND2X2_10819 ( .A(u2__abc_52155_new_n21358_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__191_));
AND2X2 AND2X2_1082 ( .A(u2__abc_52155_new_n4223_), .B(u2__abc_52155_new_n3836_), .Y(u2__abc_52155_new_n4224_));
AND2X2 AND2X2_10820 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_191_), .Y(u2__abc_52155_new_n21360_));
AND2X2 AND2X2_10821 ( .A(u2__abc_52155_new_n21349_), .B(sqrto_190_), .Y(u2__abc_52155_new_n21362_));
AND2X2 AND2X2_10822 ( .A(u2__abc_52155_new_n21363_), .B(u2__abc_52155_new_n21361_), .Y(u2__abc_52155_new_n21364_));
AND2X2 AND2X2_10823 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4784_), .Y(u2__abc_52155_new_n21366_));
AND2X2 AND2X2_10824 ( .A(u2__abc_52155_new_n21367_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21368_));
AND2X2 AND2X2_10825 ( .A(u2__abc_52155_new_n21365_), .B(u2__abc_52155_new_n21368_), .Y(u2__abc_52155_new_n21369_));
AND2X2 AND2X2_10826 ( .A(u2__abc_52155_new_n21370_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__192_));
AND2X2 AND2X2_10827 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_192_), .Y(u2__abc_52155_new_n21372_));
AND2X2 AND2X2_10828 ( .A(u2__abc_52155_new_n21362_), .B(sqrto_191_), .Y(u2__abc_52155_new_n21373_));
AND2X2 AND2X2_10829 ( .A(u2__abc_52155_new_n21374_), .B(u2__abc_52155_new_n21375_), .Y(u2__abc_52155_new_n21376_));
AND2X2 AND2X2_1083 ( .A(u2__abc_52155_new_n4222_), .B(u2__abc_52155_new_n4226_), .Y(u2__abc_52155_new_n4227_));
AND2X2 AND2X2_10830 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4765_), .Y(u2__abc_52155_new_n21378_));
AND2X2 AND2X2_10831 ( .A(u2__abc_52155_new_n21379_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21380_));
AND2X2 AND2X2_10832 ( .A(u2__abc_52155_new_n21377_), .B(u2__abc_52155_new_n21380_), .Y(u2__abc_52155_new_n21381_));
AND2X2 AND2X2_10833 ( .A(u2__abc_52155_new_n21382_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__193_));
AND2X2 AND2X2_10834 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_193_), .Y(u2__abc_52155_new_n21384_));
AND2X2 AND2X2_10835 ( .A(u2__abc_52155_new_n21373_), .B(sqrto_192_), .Y(u2__abc_52155_new_n21386_));
AND2X2 AND2X2_10836 ( .A(u2__abc_52155_new_n21387_), .B(u2__abc_52155_new_n21385_), .Y(u2__abc_52155_new_n21388_));
AND2X2 AND2X2_10837 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4770_), .Y(u2__abc_52155_new_n21390_));
AND2X2 AND2X2_10838 ( .A(u2__abc_52155_new_n21391_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21392_));
AND2X2 AND2X2_10839 ( .A(u2__abc_52155_new_n21389_), .B(u2__abc_52155_new_n21392_), .Y(u2__abc_52155_new_n21393_));
AND2X2 AND2X2_1084 ( .A(u2__abc_52155_new_n3878_), .B(u2__abc_52155_new_n3887_), .Y(u2__abc_52155_new_n4229_));
AND2X2 AND2X2_10840 ( .A(u2__abc_52155_new_n21394_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__194_));
AND2X2 AND2X2_10841 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_194_), .Y(u2__abc_52155_new_n21396_));
AND2X2 AND2X2_10842 ( .A(u2__abc_52155_new_n21386_), .B(sqrto_193_), .Y(u2__abc_52155_new_n21398_));
AND2X2 AND2X2_10843 ( .A(u2__abc_52155_new_n21399_), .B(u2__abc_52155_new_n21397_), .Y(u2__abc_52155_new_n21400_));
AND2X2 AND2X2_10844 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4756_), .Y(u2__abc_52155_new_n21402_));
AND2X2 AND2X2_10845 ( .A(u2__abc_52155_new_n21403_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21404_));
AND2X2 AND2X2_10846 ( .A(u2__abc_52155_new_n21401_), .B(u2__abc_52155_new_n21404_), .Y(u2__abc_52155_new_n21405_));
AND2X2 AND2X2_10847 ( .A(u2__abc_52155_new_n21406_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__195_));
AND2X2 AND2X2_10848 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_195_), .Y(u2__abc_52155_new_n21408_));
AND2X2 AND2X2_10849 ( .A(u2__abc_52155_new_n21398_), .B(sqrto_194_), .Y(u2__abc_52155_new_n21410_));
AND2X2 AND2X2_1085 ( .A(u2__abc_52155_new_n4230_), .B(u2__abc_52155_new_n3875_), .Y(u2__abc_52155_new_n4231_));
AND2X2 AND2X2_10850 ( .A(u2__abc_52155_new_n21411_), .B(u2__abc_52155_new_n21409_), .Y(u2__abc_52155_new_n21412_));
AND2X2 AND2X2_10851 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4749_), .Y(u2__abc_52155_new_n21414_));
AND2X2 AND2X2_10852 ( .A(u2__abc_52155_new_n21415_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21416_));
AND2X2 AND2X2_10853 ( .A(u2__abc_52155_new_n21413_), .B(u2__abc_52155_new_n21416_), .Y(u2__abc_52155_new_n21417_));
AND2X2 AND2X2_10854 ( .A(u2__abc_52155_new_n21418_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__196_));
AND2X2 AND2X2_10855 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_196_), .Y(u2__abc_52155_new_n21420_));
AND2X2 AND2X2_10856 ( .A(u2__abc_52155_new_n21410_), .B(sqrto_195_), .Y(u2__abc_52155_new_n21421_));
AND2X2 AND2X2_10857 ( .A(u2__abc_52155_new_n21422_), .B(u2__abc_52155_new_n21423_), .Y(u2__abc_52155_new_n21424_));
AND2X2 AND2X2_10858 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4734_), .Y(u2__abc_52155_new_n21426_));
AND2X2 AND2X2_10859 ( .A(u2__abc_52155_new_n21427_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21428_));
AND2X2 AND2X2_1086 ( .A(u2__abc_52155_new_n3870_), .B(u2__abc_52155_new_n3865_), .Y(u2__abc_52155_new_n4232_));
AND2X2 AND2X2_10860 ( .A(u2__abc_52155_new_n21425_), .B(u2__abc_52155_new_n21428_), .Y(u2__abc_52155_new_n21429_));
AND2X2 AND2X2_10861 ( .A(u2__abc_52155_new_n21430_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__197_));
AND2X2 AND2X2_10862 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_197_), .Y(u2__abc_52155_new_n21432_));
AND2X2 AND2X2_10863 ( .A(u2__abc_52155_new_n21421_), .B(sqrto_196_), .Y(u2__abc_52155_new_n21434_));
AND2X2 AND2X2_10864 ( .A(u2__abc_52155_new_n21435_), .B(u2__abc_52155_new_n21433_), .Y(u2__abc_52155_new_n21436_));
AND2X2 AND2X2_10865 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4741_), .Y(u2__abc_52155_new_n21438_));
AND2X2 AND2X2_10866 ( .A(u2__abc_52155_new_n21439_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21440_));
AND2X2 AND2X2_10867 ( .A(u2__abc_52155_new_n21437_), .B(u2__abc_52155_new_n21440_), .Y(u2__abc_52155_new_n21441_));
AND2X2 AND2X2_10868 ( .A(u2__abc_52155_new_n21442_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__198_));
AND2X2 AND2X2_10869 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_198_), .Y(u2__abc_52155_new_n21444_));
AND2X2 AND2X2_1087 ( .A(u2__abc_52155_new_n4228_), .B(u2__abc_52155_new_n4235_), .Y(u2__abc_52155_new_n4236_));
AND2X2 AND2X2_10870 ( .A(u2__abc_52155_new_n21434_), .B(sqrto_197_), .Y(u2__abc_52155_new_n21445_));
AND2X2 AND2X2_10871 ( .A(u2__abc_52155_new_n21446_), .B(u2__abc_52155_new_n21447_), .Y(u2__abc_52155_new_n21448_));
AND2X2 AND2X2_10872 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4693_), .Y(u2__abc_52155_new_n21450_));
AND2X2 AND2X2_10873 ( .A(u2__abc_52155_new_n21451_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21452_));
AND2X2 AND2X2_10874 ( .A(u2__abc_52155_new_n21449_), .B(u2__abc_52155_new_n21452_), .Y(u2__abc_52155_new_n21453_));
AND2X2 AND2X2_10875 ( .A(u2__abc_52155_new_n21454_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__199_));
AND2X2 AND2X2_10876 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_199_), .Y(u2__abc_52155_new_n21456_));
AND2X2 AND2X2_10877 ( .A(u2__abc_52155_new_n21445_), .B(sqrto_198_), .Y(u2__abc_52155_new_n21458_));
AND2X2 AND2X2_10878 ( .A(u2__abc_52155_new_n21459_), .B(u2__abc_52155_new_n21457_), .Y(u2__abc_52155_new_n21460_));
AND2X2 AND2X2_10879 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4686_), .Y(u2__abc_52155_new_n21462_));
AND2X2 AND2X2_1088 ( .A(u2__abc_52155_new_n3787_), .B(u2__abc_52155_new_n3796_), .Y(u2__abc_52155_new_n4238_));
AND2X2 AND2X2_10880 ( .A(u2__abc_52155_new_n21463_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21464_));
AND2X2 AND2X2_10881 ( .A(u2__abc_52155_new_n21461_), .B(u2__abc_52155_new_n21464_), .Y(u2__abc_52155_new_n21465_));
AND2X2 AND2X2_10882 ( .A(u2__abc_52155_new_n21466_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__200_));
AND2X2 AND2X2_10883 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_200_), .Y(u2__abc_52155_new_n21468_));
AND2X2 AND2X2_10884 ( .A(u2__abc_52155_new_n21458_), .B(sqrto_199_), .Y(u2__abc_52155_new_n21470_));
AND2X2 AND2X2_10885 ( .A(u2__abc_52155_new_n21471_), .B(u2__abc_52155_new_n21469_), .Y(u2__abc_52155_new_n21472_));
AND2X2 AND2X2_10886 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4671_), .Y(u2__abc_52155_new_n21474_));
AND2X2 AND2X2_10887 ( .A(u2__abc_52155_new_n21475_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21476_));
AND2X2 AND2X2_10888 ( .A(u2__abc_52155_new_n21473_), .B(u2__abc_52155_new_n21476_), .Y(u2__abc_52155_new_n21477_));
AND2X2 AND2X2_10889 ( .A(u2__abc_52155_new_n21478_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__201_));
AND2X2 AND2X2_1089 ( .A(u2__abc_52155_new_n4239_), .B(u2__abc_52155_new_n3784_), .Y(u2__abc_52155_new_n4240_));
AND2X2 AND2X2_10890 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_201_), .Y(u2__abc_52155_new_n21480_));
AND2X2 AND2X2_10891 ( .A(u2__abc_52155_new_n21470_), .B(sqrto_200_), .Y(u2__abc_52155_new_n21482_));
AND2X2 AND2X2_10892 ( .A(u2__abc_52155_new_n21483_), .B(u2__abc_52155_new_n21481_), .Y(u2__abc_52155_new_n21484_));
AND2X2 AND2X2_10893 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4678_), .Y(u2__abc_52155_new_n21486_));
AND2X2 AND2X2_10894 ( .A(u2__abc_52155_new_n21487_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21488_));
AND2X2 AND2X2_10895 ( .A(u2__abc_52155_new_n21485_), .B(u2__abc_52155_new_n21488_), .Y(u2__abc_52155_new_n21489_));
AND2X2 AND2X2_10896 ( .A(u2__abc_52155_new_n21490_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__202_));
AND2X2 AND2X2_10897 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_202_), .Y(u2__abc_52155_new_n21492_));
AND2X2 AND2X2_10898 ( .A(u2__abc_52155_new_n21482_), .B(sqrto_201_), .Y(u2__abc_52155_new_n21493_));
AND2X2 AND2X2_10899 ( .A(u2__abc_52155_new_n21494_), .B(u2__abc_52155_new_n21495_), .Y(u2__abc_52155_new_n21496_));
AND2X2 AND2X2_109 ( .A(_abc_73687_new_n927_), .B(_abc_73687_new_n926_), .Y(\o[144] ));
AND2X2 AND2X2_1090 ( .A(u2__abc_52155_new_n3779_), .B(u2__abc_52155_new_n3774_), .Y(u2__abc_52155_new_n4241_));
AND2X2 AND2X2_10900 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4724_), .Y(u2__abc_52155_new_n21498_));
AND2X2 AND2X2_10901 ( .A(u2__abc_52155_new_n21499_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21500_));
AND2X2 AND2X2_10902 ( .A(u2__abc_52155_new_n21497_), .B(u2__abc_52155_new_n21500_), .Y(u2__abc_52155_new_n21501_));
AND2X2 AND2X2_10903 ( .A(u2__abc_52155_new_n21502_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__203_));
AND2X2 AND2X2_10904 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_203_), .Y(u2__abc_52155_new_n21504_));
AND2X2 AND2X2_10905 ( .A(u2__abc_52155_new_n21493_), .B(sqrto_202_), .Y(u2__abc_52155_new_n21506_));
AND2X2 AND2X2_10906 ( .A(u2__abc_52155_new_n21507_), .B(u2__abc_52155_new_n21505_), .Y(u2__abc_52155_new_n21508_));
AND2X2 AND2X2_10907 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4717_), .Y(u2__abc_52155_new_n21510_));
AND2X2 AND2X2_10908 ( .A(u2__abc_52155_new_n21511_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21512_));
AND2X2 AND2X2_10909 ( .A(u2__abc_52155_new_n21509_), .B(u2__abc_52155_new_n21512_), .Y(u2__abc_52155_new_n21513_));
AND2X2 AND2X2_1091 ( .A(u2__abc_52155_new_n4243_), .B(u2__abc_52155_new_n3831_), .Y(u2__abc_52155_new_n4244_));
AND2X2 AND2X2_10910 ( .A(u2__abc_52155_new_n21514_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__204_));
AND2X2 AND2X2_10911 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_204_), .Y(u2__abc_52155_new_n21516_));
AND2X2 AND2X2_10912 ( .A(u2__abc_52155_new_n21506_), .B(sqrto_203_), .Y(u2__abc_52155_new_n21518_));
AND2X2 AND2X2_10913 ( .A(u2__abc_52155_new_n21519_), .B(u2__abc_52155_new_n21517_), .Y(u2__abc_52155_new_n21520_));
AND2X2 AND2X2_10914 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4702_), .Y(u2__abc_52155_new_n21522_));
AND2X2 AND2X2_10915 ( .A(u2__abc_52155_new_n21523_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21524_));
AND2X2 AND2X2_10916 ( .A(u2__abc_52155_new_n21521_), .B(u2__abc_52155_new_n21524_), .Y(u2__abc_52155_new_n21525_));
AND2X2 AND2X2_10917 ( .A(u2__abc_52155_new_n21526_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__205_));
AND2X2 AND2X2_10918 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_205_), .Y(u2__abc_52155_new_n21528_));
AND2X2 AND2X2_10919 ( .A(u2__abc_52155_new_n21518_), .B(sqrto_204_), .Y(u2__abc_52155_new_n21530_));
AND2X2 AND2X2_1092 ( .A(u2__abc_52155_new_n3818_), .B(u2__abc_52155_new_n3827_), .Y(u2__abc_52155_new_n4245_));
AND2X2 AND2X2_10920 ( .A(u2__abc_52155_new_n21531_), .B(u2__abc_52155_new_n21529_), .Y(u2__abc_52155_new_n21532_));
AND2X2 AND2X2_10921 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4709_), .Y(u2__abc_52155_new_n21534_));
AND2X2 AND2X2_10922 ( .A(u2__abc_52155_new_n21535_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21536_));
AND2X2 AND2X2_10923 ( .A(u2__abc_52155_new_n21533_), .B(u2__abc_52155_new_n21536_), .Y(u2__abc_52155_new_n21537_));
AND2X2 AND2X2_10924 ( .A(u2__abc_52155_new_n21538_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__206_));
AND2X2 AND2X2_10925 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_206_), .Y(u2__abc_52155_new_n21540_));
AND2X2 AND2X2_10926 ( .A(u2__abc_52155_new_n21530_), .B(sqrto_205_), .Y(u2__abc_52155_new_n21541_));
AND2X2 AND2X2_10927 ( .A(u2__abc_52155_new_n21542_), .B(u2__abc_52155_new_n21543_), .Y(u2__abc_52155_new_n21544_));
AND2X2 AND2X2_10928 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4622_), .Y(u2__abc_52155_new_n21546_));
AND2X2 AND2X2_10929 ( .A(u2__abc_52155_new_n21547_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21548_));
AND2X2 AND2X2_1093 ( .A(u2__abc_52155_new_n4246_), .B(u2__abc_52155_new_n3815_), .Y(u2__abc_52155_new_n4247_));
AND2X2 AND2X2_10930 ( .A(u2__abc_52155_new_n21545_), .B(u2__abc_52155_new_n21548_), .Y(u2__abc_52155_new_n21549_));
AND2X2 AND2X2_10931 ( .A(u2__abc_52155_new_n21550_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__207_));
AND2X2 AND2X2_10932 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_207_), .Y(u2__abc_52155_new_n21552_));
AND2X2 AND2X2_10933 ( .A(u2__abc_52155_new_n21541_), .B(sqrto_206_), .Y(u2__abc_52155_new_n21554_));
AND2X2 AND2X2_10934 ( .A(u2__abc_52155_new_n21555_), .B(u2__abc_52155_new_n21553_), .Y(u2__abc_52155_new_n21556_));
AND2X2 AND2X2_10935 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4629_), .Y(u2__abc_52155_new_n21558_));
AND2X2 AND2X2_10936 ( .A(u2__abc_52155_new_n21559_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21560_));
AND2X2 AND2X2_10937 ( .A(u2__abc_52155_new_n21557_), .B(u2__abc_52155_new_n21560_), .Y(u2__abc_52155_new_n21561_));
AND2X2 AND2X2_10938 ( .A(u2__abc_52155_new_n21562_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__208_));
AND2X2 AND2X2_10939 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_208_), .Y(u2__abc_52155_new_n21564_));
AND2X2 AND2X2_1094 ( .A(u2__abc_52155_new_n3810_), .B(u2__abc_52155_new_n3805_), .Y(u2__abc_52155_new_n4248_));
AND2X2 AND2X2_10940 ( .A(u2__abc_52155_new_n21554_), .B(sqrto_207_), .Y(u2__abc_52155_new_n21566_));
AND2X2 AND2X2_10941 ( .A(u2__abc_52155_new_n21567_), .B(u2__abc_52155_new_n21565_), .Y(u2__abc_52155_new_n21568_));
AND2X2 AND2X2_10942 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4607_), .Y(u2__abc_52155_new_n21570_));
AND2X2 AND2X2_10943 ( .A(u2__abc_52155_new_n21571_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21572_));
AND2X2 AND2X2_10944 ( .A(u2__abc_52155_new_n21569_), .B(u2__abc_52155_new_n21572_), .Y(u2__abc_52155_new_n21573_));
AND2X2 AND2X2_10945 ( .A(u2__abc_52155_new_n21574_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__209_));
AND2X2 AND2X2_10946 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_209_), .Y(u2__abc_52155_new_n21576_));
AND2X2 AND2X2_10947 ( .A(u2__abc_52155_new_n21566_), .B(sqrto_208_), .Y(u2__abc_52155_new_n21578_));
AND2X2 AND2X2_10948 ( .A(u2__abc_52155_new_n21579_), .B(u2__abc_52155_new_n21577_), .Y(u2__abc_52155_new_n21580_));
AND2X2 AND2X2_10949 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4614_), .Y(u2__abc_52155_new_n21582_));
AND2X2 AND2X2_1095 ( .A(u2__abc_52155_new_n4237_), .B(u2__abc_52155_new_n4252_), .Y(u2__abc_52155_new_n4253_));
AND2X2 AND2X2_10950 ( .A(u2__abc_52155_new_n21583_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21584_));
AND2X2 AND2X2_10951 ( .A(u2__abc_52155_new_n21581_), .B(u2__abc_52155_new_n21584_), .Y(u2__abc_52155_new_n21585_));
AND2X2 AND2X2_10952 ( .A(u2__abc_52155_new_n21586_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__210_));
AND2X2 AND2X2_10953 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_210_), .Y(u2__abc_52155_new_n21588_));
AND2X2 AND2X2_10954 ( .A(u2__abc_52155_new_n21578_), .B(sqrto_209_), .Y(u2__abc_52155_new_n21589_));
AND2X2 AND2X2_10955 ( .A(u2__abc_52155_new_n21590_), .B(u2__abc_52155_new_n21591_), .Y(u2__abc_52155_new_n21592_));
AND2X2 AND2X2_10956 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4660_), .Y(u2__abc_52155_new_n21594_));
AND2X2 AND2X2_10957 ( .A(u2__abc_52155_new_n21595_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21596_));
AND2X2 AND2X2_10958 ( .A(u2__abc_52155_new_n21593_), .B(u2__abc_52155_new_n21596_), .Y(u2__abc_52155_new_n21597_));
AND2X2 AND2X2_10959 ( .A(u2__abc_52155_new_n21598_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__211_));
AND2X2 AND2X2_1096 ( .A(u2__abc_52155_new_n3652_), .B(u2__abc_52155_new_n3647_), .Y(u2__abc_52155_new_n4255_));
AND2X2 AND2X2_10960 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_211_), .Y(u2__abc_52155_new_n21600_));
AND2X2 AND2X2_10961 ( .A(u2__abc_52155_new_n21589_), .B(sqrto_210_), .Y(u2__abc_52155_new_n21602_));
AND2X2 AND2X2_10962 ( .A(u2__abc_52155_new_n21603_), .B(u2__abc_52155_new_n21601_), .Y(u2__abc_52155_new_n21604_));
AND2X2 AND2X2_10963 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4653_), .Y(u2__abc_52155_new_n21606_));
AND2X2 AND2X2_10964 ( .A(u2__abc_52155_new_n21607_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21608_));
AND2X2 AND2X2_10965 ( .A(u2__abc_52155_new_n21605_), .B(u2__abc_52155_new_n21608_), .Y(u2__abc_52155_new_n21609_));
AND2X2 AND2X2_10966 ( .A(u2__abc_52155_new_n21610_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__212_));
AND2X2 AND2X2_10967 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_212_), .Y(u2__abc_52155_new_n21612_));
AND2X2 AND2X2_10968 ( .A(u2__abc_52155_new_n21602_), .B(sqrto_211_), .Y(u2__abc_52155_new_n21614_));
AND2X2 AND2X2_10969 ( .A(u2__abc_52155_new_n21615_), .B(u2__abc_52155_new_n21613_), .Y(u2__abc_52155_new_n21616_));
AND2X2 AND2X2_1097 ( .A(u2__abc_52155_new_n4256_), .B(u2__abc_52155_new_n3672_), .Y(u2__abc_52155_new_n4257_));
AND2X2 AND2X2_10970 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4638_), .Y(u2__abc_52155_new_n21618_));
AND2X2 AND2X2_10971 ( .A(u2__abc_52155_new_n21619_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21620_));
AND2X2 AND2X2_10972 ( .A(u2__abc_52155_new_n21617_), .B(u2__abc_52155_new_n21620_), .Y(u2__abc_52155_new_n21621_));
AND2X2 AND2X2_10973 ( .A(u2__abc_52155_new_n21622_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__213_));
AND2X2 AND2X2_10974 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_213_), .Y(u2__abc_52155_new_n21624_));
AND2X2 AND2X2_10975 ( .A(u2__abc_52155_new_n21614_), .B(sqrto_212_), .Y(u2__abc_52155_new_n21626_));
AND2X2 AND2X2_10976 ( .A(u2__abc_52155_new_n21627_), .B(u2__abc_52155_new_n21625_), .Y(u2__abc_52155_new_n21628_));
AND2X2 AND2X2_10977 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4645_), .Y(u2__abc_52155_new_n21630_));
AND2X2 AND2X2_10978 ( .A(u2__abc_52155_new_n21631_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21632_));
AND2X2 AND2X2_10979 ( .A(u2__abc_52155_new_n21629_), .B(u2__abc_52155_new_n21632_), .Y(u2__abc_52155_new_n21633_));
AND2X2 AND2X2_1098 ( .A(u2__abc_52155_new_n3667_), .B(u2__abc_52155_new_n3662_), .Y(u2__abc_52155_new_n4258_));
AND2X2 AND2X2_10980 ( .A(u2__abc_52155_new_n21634_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__214_));
AND2X2 AND2X2_10981 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_214_), .Y(u2__abc_52155_new_n21636_));
AND2X2 AND2X2_10982 ( .A(u2__abc_52155_new_n21626_), .B(sqrto_213_), .Y(u2__abc_52155_new_n21637_));
AND2X2 AND2X2_10983 ( .A(u2__abc_52155_new_n21638_), .B(u2__abc_52155_new_n21639_), .Y(u2__abc_52155_new_n21640_));
AND2X2 AND2X2_10984 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4559_), .Y(u2__abc_52155_new_n21642_));
AND2X2 AND2X2_10985 ( .A(u2__abc_52155_new_n21643_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21644_));
AND2X2 AND2X2_10986 ( .A(u2__abc_52155_new_n21641_), .B(u2__abc_52155_new_n21644_), .Y(u2__abc_52155_new_n21645_));
AND2X2 AND2X2_10987 ( .A(u2__abc_52155_new_n21646_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__215_));
AND2X2 AND2X2_10988 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_215_), .Y(u2__abc_52155_new_n21648_));
AND2X2 AND2X2_10989 ( .A(u2__abc_52155_new_n21637_), .B(sqrto_214_), .Y(u2__abc_52155_new_n21650_));
AND2X2 AND2X2_1099 ( .A(u2__abc_52155_new_n4260_), .B(u2__abc_52155_new_n3704_), .Y(u2__abc_52155_new_n4261_));
AND2X2 AND2X2_10990 ( .A(u2__abc_52155_new_n21651_), .B(u2__abc_52155_new_n21649_), .Y(u2__abc_52155_new_n21652_));
AND2X2 AND2X2_10991 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4566_), .Y(u2__abc_52155_new_n21654_));
AND2X2 AND2X2_10992 ( .A(u2__abc_52155_new_n21655_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21656_));
AND2X2 AND2X2_10993 ( .A(u2__abc_52155_new_n21653_), .B(u2__abc_52155_new_n21656_), .Y(u2__abc_52155_new_n21657_));
AND2X2 AND2X2_10994 ( .A(u2__abc_52155_new_n21658_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__216_));
AND2X2 AND2X2_10995 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_216_), .Y(u2__abc_52155_new_n21660_));
AND2X2 AND2X2_10996 ( .A(u2__abc_52155_new_n21650_), .B(sqrto_215_), .Y(u2__abc_52155_new_n21662_));
AND2X2 AND2X2_10997 ( .A(u2__abc_52155_new_n21663_), .B(u2__abc_52155_new_n21661_), .Y(u2__abc_52155_new_n21664_));
AND2X2 AND2X2_10998 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4544_), .Y(u2__abc_52155_new_n21666_));
AND2X2 AND2X2_10999 ( .A(u2__abc_52155_new_n21667_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21668_));
AND2X2 AND2X2_11 ( .A(_abc_73687_new_n753_), .B(sqrto_10_), .Y(\o[46] ));
AND2X2 AND2X2_110 ( .A(_abc_73687_new_n930_), .B(_abc_73687_new_n929_), .Y(\o[145] ));
AND2X2 AND2X2_1100 ( .A(u2__abc_52155_new_n3686_), .B(u2__abc_52155_new_n3678_), .Y(u2__abc_52155_new_n4262_));
AND2X2 AND2X2_11000 ( .A(u2__abc_52155_new_n21665_), .B(u2__abc_52155_new_n21668_), .Y(u2__abc_52155_new_n21669_));
AND2X2 AND2X2_11001 ( .A(u2__abc_52155_new_n21670_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__217_));
AND2X2 AND2X2_11002 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_217_), .Y(u2__abc_52155_new_n21672_));
AND2X2 AND2X2_11003 ( .A(u2__abc_52155_new_n21662_), .B(sqrto_216_), .Y(u2__abc_52155_new_n21674_));
AND2X2 AND2X2_11004 ( .A(u2__abc_52155_new_n21675_), .B(u2__abc_52155_new_n21673_), .Y(u2__abc_52155_new_n21676_));
AND2X2 AND2X2_11005 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4551_), .Y(u2__abc_52155_new_n21678_));
AND2X2 AND2X2_11006 ( .A(u2__abc_52155_new_n21679_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21680_));
AND2X2 AND2X2_11007 ( .A(u2__abc_52155_new_n21677_), .B(u2__abc_52155_new_n21680_), .Y(u2__abc_52155_new_n21681_));
AND2X2 AND2X2_11008 ( .A(u2__abc_52155_new_n21682_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__218_));
AND2X2 AND2X2_11009 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_218_), .Y(u2__abc_52155_new_n21684_));
AND2X2 AND2X2_1101 ( .A(u2__abc_52155_new_n3691_), .B(u2__abc_52155_new_n3700_), .Y(u2__abc_52155_new_n4264_));
AND2X2 AND2X2_11010 ( .A(u2__abc_52155_new_n21674_), .B(sqrto_217_), .Y(u2__abc_52155_new_n21685_));
AND2X2 AND2X2_11011 ( .A(u2__abc_52155_new_n21686_), .B(u2__abc_52155_new_n21687_), .Y(u2__abc_52155_new_n21688_));
AND2X2 AND2X2_11012 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4597_), .Y(u2__abc_52155_new_n21690_));
AND2X2 AND2X2_11013 ( .A(u2__abc_52155_new_n21691_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21692_));
AND2X2 AND2X2_11014 ( .A(u2__abc_52155_new_n21689_), .B(u2__abc_52155_new_n21692_), .Y(u2__abc_52155_new_n21693_));
AND2X2 AND2X2_11015 ( .A(u2__abc_52155_new_n21694_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__219_));
AND2X2 AND2X2_11016 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_219_), .Y(u2__abc_52155_new_n21696_));
AND2X2 AND2X2_11017 ( .A(u2__abc_52155_new_n21685_), .B(sqrto_218_), .Y(u2__abc_52155_new_n21698_));
AND2X2 AND2X2_11018 ( .A(u2__abc_52155_new_n21699_), .B(u2__abc_52155_new_n21697_), .Y(u2__abc_52155_new_n21700_));
AND2X2 AND2X2_11019 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4590_), .Y(u2__abc_52155_new_n21702_));
AND2X2 AND2X2_1102 ( .A(u2__abc_52155_new_n4265_), .B(u2__abc_52155_new_n3688_), .Y(u2__abc_52155_new_n4266_));
AND2X2 AND2X2_11020 ( .A(u2__abc_52155_new_n21703_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21704_));
AND2X2 AND2X2_11021 ( .A(u2__abc_52155_new_n21701_), .B(u2__abc_52155_new_n21704_), .Y(u2__abc_52155_new_n21705_));
AND2X2 AND2X2_11022 ( .A(u2__abc_52155_new_n21706_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__220_));
AND2X2 AND2X2_11023 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_220_), .Y(u2__abc_52155_new_n21708_));
AND2X2 AND2X2_11024 ( .A(u2__abc_52155_new_n21698_), .B(sqrto_219_), .Y(u2__abc_52155_new_n21710_));
AND2X2 AND2X2_11025 ( .A(u2__abc_52155_new_n21711_), .B(u2__abc_52155_new_n21709_), .Y(u2__abc_52155_new_n21712_));
AND2X2 AND2X2_11026 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4575_), .Y(u2__abc_52155_new_n21714_));
AND2X2 AND2X2_11027 ( .A(u2__abc_52155_new_n21715_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21716_));
AND2X2 AND2X2_11028 ( .A(u2__abc_52155_new_n21713_), .B(u2__abc_52155_new_n21716_), .Y(u2__abc_52155_new_n21717_));
AND2X2 AND2X2_11029 ( .A(u2__abc_52155_new_n21718_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__221_));
AND2X2 AND2X2_1103 ( .A(u2__abc_52155_new_n3715_), .B(u2__abc_52155_new_n3710_), .Y(u2__abc_52155_new_n4269_));
AND2X2 AND2X2_11030 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_221_), .Y(u2__abc_52155_new_n21720_));
AND2X2 AND2X2_11031 ( .A(u2__abc_52155_new_n21710_), .B(sqrto_220_), .Y(u2__abc_52155_new_n21722_));
AND2X2 AND2X2_11032 ( .A(u2__abc_52155_new_n21723_), .B(u2__abc_52155_new_n21721_), .Y(u2__abc_52155_new_n21724_));
AND2X2 AND2X2_11033 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4582_), .Y(u2__abc_52155_new_n21726_));
AND2X2 AND2X2_11034 ( .A(u2__abc_52155_new_n21727_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21728_));
AND2X2 AND2X2_11035 ( .A(u2__abc_52155_new_n21725_), .B(u2__abc_52155_new_n21728_), .Y(u2__abc_52155_new_n21729_));
AND2X2 AND2X2_11036 ( .A(u2__abc_52155_new_n21730_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__222_));
AND2X2 AND2X2_11037 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_222_), .Y(u2__abc_52155_new_n21732_));
AND2X2 AND2X2_11038 ( .A(u2__abc_52155_new_n21722_), .B(sqrto_221_), .Y(u2__abc_52155_new_n21733_));
AND2X2 AND2X2_11039 ( .A(u2__abc_52155_new_n21734_), .B(u2__abc_52155_new_n21735_), .Y(u2__abc_52155_new_n21736_));
AND2X2 AND2X2_1104 ( .A(u2__abc_52155_new_n4270_), .B(u2__abc_52155_new_n3735_), .Y(u2__abc_52155_new_n4271_));
AND2X2 AND2X2_11040 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4501_), .Y(u2__abc_52155_new_n21738_));
AND2X2 AND2X2_11041 ( .A(u2__abc_52155_new_n21739_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21740_));
AND2X2 AND2X2_11042 ( .A(u2__abc_52155_new_n21737_), .B(u2__abc_52155_new_n21740_), .Y(u2__abc_52155_new_n21741_));
AND2X2 AND2X2_11043 ( .A(u2__abc_52155_new_n21742_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__223_));
AND2X2 AND2X2_11044 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_223_), .Y(u2__abc_52155_new_n21744_));
AND2X2 AND2X2_11045 ( .A(u2__abc_52155_new_n21733_), .B(sqrto_222_), .Y(u2__abc_52155_new_n21746_));
AND2X2 AND2X2_11046 ( .A(u2__abc_52155_new_n21747_), .B(u2__abc_52155_new_n21745_), .Y(u2__abc_52155_new_n21748_));
AND2X2 AND2X2_11047 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4494_), .Y(u2__abc_52155_new_n21750_));
AND2X2 AND2X2_11048 ( .A(u2__abc_52155_new_n21751_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21752_));
AND2X2 AND2X2_11049 ( .A(u2__abc_52155_new_n21749_), .B(u2__abc_52155_new_n21752_), .Y(u2__abc_52155_new_n21753_));
AND2X2 AND2X2_1105 ( .A(u2__abc_52155_new_n3730_), .B(u2__abc_52155_new_n3725_), .Y(u2__abc_52155_new_n4272_));
AND2X2 AND2X2_11050 ( .A(u2__abc_52155_new_n21754_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__224_));
AND2X2 AND2X2_11051 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_224_), .Y(u2__abc_52155_new_n21756_));
AND2X2 AND2X2_11052 ( .A(u2__abc_52155_new_n21746_), .B(sqrto_223_), .Y(u2__abc_52155_new_n21757_));
AND2X2 AND2X2_11053 ( .A(u2__abc_52155_new_n21758_), .B(u2__abc_52155_new_n21759_), .Y(u2__abc_52155_new_n21760_));
AND2X2 AND2X2_11054 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4479_), .Y(u2__abc_52155_new_n21762_));
AND2X2 AND2X2_11055 ( .A(u2__abc_52155_new_n21763_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21764_));
AND2X2 AND2X2_11056 ( .A(u2__abc_52155_new_n21761_), .B(u2__abc_52155_new_n21764_), .Y(u2__abc_52155_new_n21765_));
AND2X2 AND2X2_11057 ( .A(u2__abc_52155_new_n21766_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__225_));
AND2X2 AND2X2_11058 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_225_), .Y(u2__abc_52155_new_n21768_));
AND2X2 AND2X2_11059 ( .A(u2__abc_52155_new_n21757_), .B(sqrto_224_), .Y(u2__abc_52155_new_n21770_));
AND2X2 AND2X2_1106 ( .A(u2__abc_52155_new_n4274_), .B(u2__abc_52155_new_n3767_), .Y(u2__abc_52155_new_n4275_));
AND2X2 AND2X2_11060 ( .A(u2__abc_52155_new_n21771_), .B(u2__abc_52155_new_n21769_), .Y(u2__abc_52155_new_n21772_));
AND2X2 AND2X2_11061 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4486_), .Y(u2__abc_52155_new_n21774_));
AND2X2 AND2X2_11062 ( .A(u2__abc_52155_new_n21775_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21776_));
AND2X2 AND2X2_11063 ( .A(u2__abc_52155_new_n21773_), .B(u2__abc_52155_new_n21776_), .Y(u2__abc_52155_new_n21777_));
AND2X2 AND2X2_11064 ( .A(u2__abc_52155_new_n21778_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__226_));
AND2X2 AND2X2_11065 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_226_), .Y(u2__abc_52155_new_n21780_));
AND2X2 AND2X2_11066 ( .A(u2__abc_52155_new_n21770_), .B(sqrto_225_), .Y(u2__abc_52155_new_n21781_));
AND2X2 AND2X2_11067 ( .A(u2__abc_52155_new_n21782_), .B(u2__abc_52155_new_n21783_), .Y(u2__abc_52155_new_n21784_));
AND2X2 AND2X2_11068 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4532_), .Y(u2__abc_52155_new_n21786_));
AND2X2 AND2X2_11069 ( .A(u2__abc_52155_new_n21787_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21788_));
AND2X2 AND2X2_1107 ( .A(u2__abc_52155_new_n3746_), .B(u2__abc_52155_new_n3741_), .Y(u2__abc_52155_new_n4276_));
AND2X2 AND2X2_11070 ( .A(u2__abc_52155_new_n21785_), .B(u2__abc_52155_new_n21788_), .Y(u2__abc_52155_new_n21789_));
AND2X2 AND2X2_11071 ( .A(u2__abc_52155_new_n21790_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__227_));
AND2X2 AND2X2_11072 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_227_), .Y(u2__abc_52155_new_n21792_));
AND2X2 AND2X2_11073 ( .A(u2__abc_52155_new_n21781_), .B(u2_o_226_), .Y(u2__abc_52155_new_n21794_));
AND2X2 AND2X2_11074 ( .A(u2__abc_52155_new_n21795_), .B(u2__abc_52155_new_n21793_), .Y(u2__abc_52155_new_n21796_));
AND2X2 AND2X2_11075 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4525_), .Y(u2__abc_52155_new_n21798_));
AND2X2 AND2X2_11076 ( .A(u2__abc_52155_new_n21799_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21800_));
AND2X2 AND2X2_11077 ( .A(u2__abc_52155_new_n21797_), .B(u2__abc_52155_new_n21800_), .Y(u2__abc_52155_new_n21801_));
AND2X2 AND2X2_11078 ( .A(u2__abc_52155_new_n21802_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__228_));
AND2X2 AND2X2_11079 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_228_), .Y(u2__abc_52155_new_n21804_));
AND2X2 AND2X2_1108 ( .A(u2__abc_52155_new_n3754_), .B(u2__abc_52155_new_n3763_), .Y(u2__abc_52155_new_n4278_));
AND2X2 AND2X2_11080 ( .A(u2__abc_52155_new_n21794_), .B(u2_o_227_), .Y(u2__abc_52155_new_n21806_));
AND2X2 AND2X2_11081 ( .A(u2__abc_52155_new_n21807_), .B(u2__abc_52155_new_n21805_), .Y(u2__abc_52155_new_n21808_));
AND2X2 AND2X2_11082 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4510_), .Y(u2__abc_52155_new_n21810_));
AND2X2 AND2X2_11083 ( .A(u2__abc_52155_new_n21811_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21812_));
AND2X2 AND2X2_11084 ( .A(u2__abc_52155_new_n21809_), .B(u2__abc_52155_new_n21812_), .Y(u2__abc_52155_new_n21813_));
AND2X2 AND2X2_11085 ( .A(u2__abc_52155_new_n21814_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__229_));
AND2X2 AND2X2_11086 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_229_), .Y(u2__abc_52155_new_n21816_));
AND2X2 AND2X2_11087 ( .A(u2__abc_52155_new_n21806_), .B(u2_o_228_), .Y(u2__abc_52155_new_n21818_));
AND2X2 AND2X2_11088 ( .A(u2__abc_52155_new_n21819_), .B(u2__abc_52155_new_n21817_), .Y(u2__abc_52155_new_n21820_));
AND2X2 AND2X2_11089 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4517_), .Y(u2__abc_52155_new_n21822_));
AND2X2 AND2X2_1109 ( .A(u2__abc_52155_new_n4279_), .B(u2__abc_52155_new_n3751_), .Y(u2__abc_52155_new_n4280_));
AND2X2 AND2X2_11090 ( .A(u2__abc_52155_new_n21823_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21824_));
AND2X2 AND2X2_11091 ( .A(u2__abc_52155_new_n21821_), .B(u2__abc_52155_new_n21824_), .Y(u2__abc_52155_new_n21825_));
AND2X2 AND2X2_11092 ( .A(u2__abc_52155_new_n21826_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__230_));
AND2X2 AND2X2_11093 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_230_), .Y(u2__abc_52155_new_n21828_));
AND2X2 AND2X2_11094 ( .A(u2__abc_52155_new_n21818_), .B(u2_o_229_), .Y(u2__abc_52155_new_n21829_));
AND2X2 AND2X2_11095 ( .A(u2__abc_52155_new_n21830_), .B(u2__abc_52155_new_n21831_), .Y(u2__abc_52155_new_n21832_));
AND2X2 AND2X2_11096 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4469_), .Y(u2__abc_52155_new_n21834_));
AND2X2 AND2X2_11097 ( .A(u2__abc_52155_new_n21835_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21836_));
AND2X2 AND2X2_11098 ( .A(u2__abc_52155_new_n21833_), .B(u2__abc_52155_new_n21836_), .Y(u2__abc_52155_new_n21837_));
AND2X2 AND2X2_11099 ( .A(u2__abc_52155_new_n21838_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__231_));
AND2X2 AND2X2_111 ( .A(_abc_73687_new_n933_), .B(_abc_73687_new_n932_), .Y(\o[146] ));
AND2X2 AND2X2_1110 ( .A(u2__abc_52155_new_n4282_), .B(u2__abc_52155_new_n3705_), .Y(u2__abc_52155_new_n4283_));
AND2X2 AND2X2_11100 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_231_), .Y(u2__abc_52155_new_n21840_));
AND2X2 AND2X2_11101 ( .A(u2__abc_52155_new_n21829_), .B(u2_o_230_), .Y(u2__abc_52155_new_n21842_));
AND2X2 AND2X2_11102 ( .A(u2__abc_52155_new_n21843_), .B(u2__abc_52155_new_n21841_), .Y(u2__abc_52155_new_n21844_));
AND2X2 AND2X2_11103 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4462_), .Y(u2__abc_52155_new_n21846_));
AND2X2 AND2X2_11104 ( .A(u2__abc_52155_new_n21847_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21848_));
AND2X2 AND2X2_11105 ( .A(u2__abc_52155_new_n21845_), .B(u2__abc_52155_new_n21848_), .Y(u2__abc_52155_new_n21849_));
AND2X2 AND2X2_11106 ( .A(u2__abc_52155_new_n21850_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__232_));
AND2X2 AND2X2_11107 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_232_), .Y(u2__abc_52155_new_n21852_));
AND2X2 AND2X2_11108 ( .A(u2__abc_52155_new_n21842_), .B(u2_o_231_), .Y(u2__abc_52155_new_n21854_));
AND2X2 AND2X2_11109 ( .A(u2__abc_52155_new_n21855_), .B(u2__abc_52155_new_n21853_), .Y(u2__abc_52155_new_n21856_));
AND2X2 AND2X2_1111 ( .A(u2__abc_52155_new_n4254_), .B(u2__abc_52155_new_n4285_), .Y(u2__abc_52155_new_n4286_));
AND2X2 AND2X2_11110 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4447_), .Y(u2__abc_52155_new_n21858_));
AND2X2 AND2X2_11111 ( .A(u2__abc_52155_new_n21859_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21860_));
AND2X2 AND2X2_11112 ( .A(u2__abc_52155_new_n21857_), .B(u2__abc_52155_new_n21860_), .Y(u2__abc_52155_new_n21861_));
AND2X2 AND2X2_11113 ( .A(u2__abc_52155_new_n21862_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__233_));
AND2X2 AND2X2_11114 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_233_), .Y(u2__abc_52155_new_n21864_));
AND2X2 AND2X2_11115 ( .A(u2__abc_52155_new_n21854_), .B(u2_o_232_), .Y(u2__abc_52155_new_n21866_));
AND2X2 AND2X2_11116 ( .A(u2__abc_52155_new_n21867_), .B(u2__abc_52155_new_n21865_), .Y(u2__abc_52155_new_n21868_));
AND2X2 AND2X2_11117 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4454_), .Y(u2__abc_52155_new_n21870_));
AND2X2 AND2X2_11118 ( .A(u2__abc_52155_new_n21871_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21872_));
AND2X2 AND2X2_11119 ( .A(u2__abc_52155_new_n21869_), .B(u2__abc_52155_new_n21872_), .Y(u2__abc_52155_new_n21873_));
AND2X2 AND2X2_1112 ( .A(u2__abc_52155_new_n4216_), .B(u2__abc_52155_new_n4286_), .Y(u2__abc_52155_new_n4287_));
AND2X2 AND2X2_11120 ( .A(u2__abc_52155_new_n21874_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__234_));
AND2X2 AND2X2_11121 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_234_), .Y(u2__abc_52155_new_n21876_));
AND2X2 AND2X2_11122 ( .A(u2__abc_52155_new_n21866_), .B(u2_o_233_), .Y(u2__abc_52155_new_n21877_));
AND2X2 AND2X2_11123 ( .A(u2__abc_52155_new_n21878_), .B(u2__abc_52155_new_n21879_), .Y(u2__abc_52155_new_n21880_));
AND2X2 AND2X2_11124 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4438_), .Y(u2__abc_52155_new_n21882_));
AND2X2 AND2X2_11125 ( .A(u2__abc_52155_new_n21883_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21884_));
AND2X2 AND2X2_11126 ( .A(u2__abc_52155_new_n21881_), .B(u2__abc_52155_new_n21884_), .Y(u2__abc_52155_new_n21885_));
AND2X2 AND2X2_11127 ( .A(u2__abc_52155_new_n21886_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__235_));
AND2X2 AND2X2_11128 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_235_), .Y(u2__abc_52155_new_n21888_));
AND2X2 AND2X2_11129 ( .A(u2__abc_52155_new_n21877_), .B(u2_o_234_), .Y(u2__abc_52155_new_n21890_));
AND2X2 AND2X2_1113 ( .A(u2__abc_52155_new_n4134_), .B(u2__abc_52155_new_n4287_), .Y(u2__abc_52155_new_n4288_));
AND2X2 AND2X2_11130 ( .A(u2__abc_52155_new_n21891_), .B(u2__abc_52155_new_n21889_), .Y(u2__abc_52155_new_n21892_));
AND2X2 AND2X2_11131 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4431_), .Y(u2__abc_52155_new_n21894_));
AND2X2 AND2X2_11132 ( .A(u2__abc_52155_new_n21895_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21896_));
AND2X2 AND2X2_11133 ( .A(u2__abc_52155_new_n21893_), .B(u2__abc_52155_new_n21896_), .Y(u2__abc_52155_new_n21897_));
AND2X2 AND2X2_11134 ( .A(u2__abc_52155_new_n21898_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__236_));
AND2X2 AND2X2_11135 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_236_), .Y(u2__abc_52155_new_n21900_));
AND2X2 AND2X2_11136 ( .A(u2__abc_52155_new_n21890_), .B(u2_o_235_), .Y(u2__abc_52155_new_n21902_));
AND2X2 AND2X2_11137 ( .A(u2__abc_52155_new_n21903_), .B(u2__abc_52155_new_n21901_), .Y(u2__abc_52155_new_n21904_));
AND2X2 AND2X2_11138 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4416_), .Y(u2__abc_52155_new_n21906_));
AND2X2 AND2X2_11139 ( .A(u2__abc_52155_new_n21907_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21908_));
AND2X2 AND2X2_1114 ( .A(u2__abc_52155_new_n4289_), .B(u2_remHi_246_), .Y(u2__abc_52155_new_n4290_));
AND2X2 AND2X2_11140 ( .A(u2__abc_52155_new_n21905_), .B(u2__abc_52155_new_n21908_), .Y(u2__abc_52155_new_n21909_));
AND2X2 AND2X2_11141 ( .A(u2__abc_52155_new_n21910_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__237_));
AND2X2 AND2X2_11142 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_237_), .Y(u2__abc_52155_new_n21912_));
AND2X2 AND2X2_11143 ( .A(u2__abc_52155_new_n21902_), .B(u2_o_236_), .Y(u2__abc_52155_new_n21914_));
AND2X2 AND2X2_11144 ( .A(u2__abc_52155_new_n21915_), .B(u2__abc_52155_new_n21913_), .Y(u2__abc_52155_new_n21916_));
AND2X2 AND2X2_11145 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4423_), .Y(u2__abc_52155_new_n21918_));
AND2X2 AND2X2_11146 ( .A(u2__abc_52155_new_n21919_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21920_));
AND2X2 AND2X2_11147 ( .A(u2__abc_52155_new_n21917_), .B(u2__abc_52155_new_n21920_), .Y(u2__abc_52155_new_n21921_));
AND2X2 AND2X2_11148 ( .A(u2__abc_52155_new_n21922_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__238_));
AND2X2 AND2X2_11149 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_238_), .Y(u2__abc_52155_new_n21924_));
AND2X2 AND2X2_1115 ( .A(u2__abc_52155_new_n4292_), .B(u2_o_246_), .Y(u2__abc_52155_new_n4293_));
AND2X2 AND2X2_11150 ( .A(u2__abc_52155_new_n21914_), .B(u2_o_237_), .Y(u2__abc_52155_new_n21925_));
AND2X2 AND2X2_11151 ( .A(u2__abc_52155_new_n21926_), .B(u2__abc_52155_new_n21927_), .Y(u2__abc_52155_new_n21928_));
AND2X2 AND2X2_11152 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4352_), .Y(u2__abc_52155_new_n21930_));
AND2X2 AND2X2_11153 ( .A(u2__abc_52155_new_n21931_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21932_));
AND2X2 AND2X2_11154 ( .A(u2__abc_52155_new_n21929_), .B(u2__abc_52155_new_n21932_), .Y(u2__abc_52155_new_n21933_));
AND2X2 AND2X2_11155 ( .A(u2__abc_52155_new_n21934_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__239_));
AND2X2 AND2X2_11156 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_239_), .Y(u2__abc_52155_new_n21936_));
AND2X2 AND2X2_11157 ( .A(u2__abc_52155_new_n21925_), .B(u2_o_238_), .Y(u2__abc_52155_new_n21938_));
AND2X2 AND2X2_11158 ( .A(u2__abc_52155_new_n21939_), .B(u2__abc_52155_new_n21937_), .Y(u2__abc_52155_new_n21940_));
AND2X2 AND2X2_11159 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4359_), .Y(u2__abc_52155_new_n21942_));
AND2X2 AND2X2_1116 ( .A(u2__abc_52155_new_n4291_), .B(u2__abc_52155_new_n4294_), .Y(u2__abc_52155_new_n4295_));
AND2X2 AND2X2_11160 ( .A(u2__abc_52155_new_n21943_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21944_));
AND2X2 AND2X2_11161 ( .A(u2__abc_52155_new_n21941_), .B(u2__abc_52155_new_n21944_), .Y(u2__abc_52155_new_n21945_));
AND2X2 AND2X2_11162 ( .A(u2__abc_52155_new_n21946_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__240_));
AND2X2 AND2X2_11163 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_240_), .Y(u2__abc_52155_new_n21948_));
AND2X2 AND2X2_11164 ( .A(u2__abc_52155_new_n21938_), .B(u2_o_239_), .Y(u2__abc_52155_new_n21949_));
AND2X2 AND2X2_11165 ( .A(u2__abc_52155_new_n21950_), .B(u2__abc_52155_new_n21951_), .Y(u2__abc_52155_new_n21952_));
AND2X2 AND2X2_11166 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4367_), .Y(u2__abc_52155_new_n21954_));
AND2X2 AND2X2_11167 ( .A(u2__abc_52155_new_n21955_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21956_));
AND2X2 AND2X2_11168 ( .A(u2__abc_52155_new_n21953_), .B(u2__abc_52155_new_n21956_), .Y(u2__abc_52155_new_n21957_));
AND2X2 AND2X2_11169 ( .A(u2__abc_52155_new_n21958_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__241_));
AND2X2 AND2X2_1117 ( .A(u2__abc_52155_new_n4296_), .B(u2_remHi_247_), .Y(u2__abc_52155_new_n4297_));
AND2X2 AND2X2_11170 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_241_), .Y(u2__abc_52155_new_n21960_));
AND2X2 AND2X2_11171 ( .A(u2__abc_52155_new_n21949_), .B(u2_o_240_), .Y(u2__abc_52155_new_n21962_));
AND2X2 AND2X2_11172 ( .A(u2__abc_52155_new_n21963_), .B(u2__abc_52155_new_n21961_), .Y(u2__abc_52155_new_n21964_));
AND2X2 AND2X2_11173 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4374_), .Y(u2__abc_52155_new_n21966_));
AND2X2 AND2X2_11174 ( .A(u2__abc_52155_new_n21967_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21968_));
AND2X2 AND2X2_11175 ( .A(u2__abc_52155_new_n21965_), .B(u2__abc_52155_new_n21968_), .Y(u2__abc_52155_new_n21969_));
AND2X2 AND2X2_11176 ( .A(u2__abc_52155_new_n21970_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__242_));
AND2X2 AND2X2_11177 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_242_), .Y(u2__abc_52155_new_n21972_));
AND2X2 AND2X2_11178 ( .A(u2__abc_52155_new_n21962_), .B(u2_o_241_), .Y(u2__abc_52155_new_n21973_));
AND2X2 AND2X2_11179 ( .A(u2__abc_52155_new_n21974_), .B(u2__abc_52155_new_n21975_), .Y(u2__abc_52155_new_n21976_));
AND2X2 AND2X2_1118 ( .A(u2__abc_52155_new_n4299_), .B(u2_o_247_), .Y(u2__abc_52155_new_n4300_));
AND2X2 AND2X2_11180 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4405_), .Y(u2__abc_52155_new_n21978_));
AND2X2 AND2X2_11181 ( .A(u2__abc_52155_new_n21979_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21980_));
AND2X2 AND2X2_11182 ( .A(u2__abc_52155_new_n21977_), .B(u2__abc_52155_new_n21980_), .Y(u2__abc_52155_new_n21981_));
AND2X2 AND2X2_11183 ( .A(u2__abc_52155_new_n21982_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__243_));
AND2X2 AND2X2_11184 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_243_), .Y(u2__abc_52155_new_n21984_));
AND2X2 AND2X2_11185 ( .A(u2__abc_52155_new_n21973_), .B(u2_o_242_), .Y(u2__abc_52155_new_n21986_));
AND2X2 AND2X2_11186 ( .A(u2__abc_52155_new_n21987_), .B(u2__abc_52155_new_n21985_), .Y(u2__abc_52155_new_n21988_));
AND2X2 AND2X2_11187 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4398_), .Y(u2__abc_52155_new_n21990_));
AND2X2 AND2X2_11188 ( .A(u2__abc_52155_new_n21991_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n21992_));
AND2X2 AND2X2_11189 ( .A(u2__abc_52155_new_n21989_), .B(u2__abc_52155_new_n21992_), .Y(u2__abc_52155_new_n21993_));
AND2X2 AND2X2_1119 ( .A(u2__abc_52155_new_n4298_), .B(u2__abc_52155_new_n4301_), .Y(u2__abc_52155_new_n4302_));
AND2X2 AND2X2_11190 ( .A(u2__abc_52155_new_n21994_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__244_));
AND2X2 AND2X2_11191 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_244_), .Y(u2__abc_52155_new_n21996_));
AND2X2 AND2X2_11192 ( .A(u2__abc_52155_new_n21986_), .B(u2_o_243_), .Y(u2__abc_52155_new_n21998_));
AND2X2 AND2X2_11193 ( .A(u2__abc_52155_new_n21999_), .B(u2__abc_52155_new_n21997_), .Y(u2__abc_52155_new_n22000_));
AND2X2 AND2X2_11194 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4383_), .Y(u2__abc_52155_new_n22002_));
AND2X2 AND2X2_11195 ( .A(u2__abc_52155_new_n22003_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22004_));
AND2X2 AND2X2_11196 ( .A(u2__abc_52155_new_n22001_), .B(u2__abc_52155_new_n22004_), .Y(u2__abc_52155_new_n22005_));
AND2X2 AND2X2_11197 ( .A(u2__abc_52155_new_n22006_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__245_));
AND2X2 AND2X2_11198 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_245_), .Y(u2__abc_52155_new_n22008_));
AND2X2 AND2X2_11199 ( .A(u2__abc_52155_new_n21998_), .B(u2_o_244_), .Y(u2__abc_52155_new_n22010_));
AND2X2 AND2X2_112 ( .A(_abc_73687_new_n936_), .B(_abc_73687_new_n935_), .Y(\o[147] ));
AND2X2 AND2X2_1120 ( .A(u2__abc_52155_new_n4295_), .B(u2__abc_52155_new_n4302_), .Y(u2__abc_52155_new_n4303_));
AND2X2 AND2X2_11200 ( .A(u2__abc_52155_new_n22011_), .B(u2__abc_52155_new_n22009_), .Y(u2__abc_52155_new_n22012_));
AND2X2 AND2X2_11201 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4390_), .Y(u2__abc_52155_new_n22014_));
AND2X2 AND2X2_11202 ( .A(u2__abc_52155_new_n22015_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22016_));
AND2X2 AND2X2_11203 ( .A(u2__abc_52155_new_n22013_), .B(u2__abc_52155_new_n22016_), .Y(u2__abc_52155_new_n22017_));
AND2X2 AND2X2_11204 ( .A(u2__abc_52155_new_n22018_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__246_));
AND2X2 AND2X2_11205 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_246_), .Y(u2__abc_52155_new_n22020_));
AND2X2 AND2X2_11206 ( .A(u2__abc_52155_new_n22010_), .B(u2_o_245_), .Y(u2__abc_52155_new_n22021_));
AND2X2 AND2X2_11207 ( .A(u2__abc_52155_new_n22022_), .B(u2__abc_52155_new_n22023_), .Y(u2__abc_52155_new_n22024_));
AND2X2 AND2X2_11208 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4289_), .Y(u2__abc_52155_new_n22026_));
AND2X2 AND2X2_11209 ( .A(u2__abc_52155_new_n22027_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22028_));
AND2X2 AND2X2_1121 ( .A(u2__abc_52155_new_n4304_), .B(u2_remHi_248_), .Y(u2__abc_52155_new_n4305_));
AND2X2 AND2X2_11210 ( .A(u2__abc_52155_new_n22025_), .B(u2__abc_52155_new_n22028_), .Y(u2__abc_52155_new_n22029_));
AND2X2 AND2X2_11211 ( .A(u2__abc_52155_new_n22030_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__247_));
AND2X2 AND2X2_11212 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_247_), .Y(u2__abc_52155_new_n22032_));
AND2X2 AND2X2_11213 ( .A(u2__abc_52155_new_n22021_), .B(u2_o_246_), .Y(u2__abc_52155_new_n22034_));
AND2X2 AND2X2_11214 ( .A(u2__abc_52155_new_n22035_), .B(u2__abc_52155_new_n22033_), .Y(u2__abc_52155_new_n22036_));
AND2X2 AND2X2_11215 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4296_), .Y(u2__abc_52155_new_n22038_));
AND2X2 AND2X2_11216 ( .A(u2__abc_52155_new_n22039_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22040_));
AND2X2 AND2X2_11217 ( .A(u2__abc_52155_new_n22037_), .B(u2__abc_52155_new_n22040_), .Y(u2__abc_52155_new_n22041_));
AND2X2 AND2X2_11218 ( .A(u2__abc_52155_new_n22042_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__248_));
AND2X2 AND2X2_11219 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_248_), .Y(u2__abc_52155_new_n22044_));
AND2X2 AND2X2_1122 ( .A(u2__abc_52155_new_n4307_), .B(u2_o_248_), .Y(u2__abc_52155_new_n4308_));
AND2X2 AND2X2_11220 ( .A(u2__abc_52155_new_n22034_), .B(u2_o_247_), .Y(u2__abc_52155_new_n22045_));
AND2X2 AND2X2_11221 ( .A(u2__abc_52155_new_n22046_), .B(u2__abc_52155_new_n22047_), .Y(u2__abc_52155_new_n22048_));
AND2X2 AND2X2_11222 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4304_), .Y(u2__abc_52155_new_n22050_));
AND2X2 AND2X2_11223 ( .A(u2__abc_52155_new_n22051_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22052_));
AND2X2 AND2X2_11224 ( .A(u2__abc_52155_new_n22049_), .B(u2__abc_52155_new_n22052_), .Y(u2__abc_52155_new_n22053_));
AND2X2 AND2X2_11225 ( .A(u2__abc_52155_new_n22054_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__249_));
AND2X2 AND2X2_11226 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_249_), .Y(u2__abc_52155_new_n22056_));
AND2X2 AND2X2_11227 ( .A(u2__abc_52155_new_n22045_), .B(u2_o_248_), .Y(u2__abc_52155_new_n22058_));
AND2X2 AND2X2_11228 ( .A(u2__abc_52155_new_n22059_), .B(u2__abc_52155_new_n22057_), .Y(u2__abc_52155_new_n22060_));
AND2X2 AND2X2_11229 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4311_), .Y(u2__abc_52155_new_n22062_));
AND2X2 AND2X2_1123 ( .A(u2__abc_52155_new_n4306_), .B(u2__abc_52155_new_n4309_), .Y(u2__abc_52155_new_n4310_));
AND2X2 AND2X2_11230 ( .A(u2__abc_52155_new_n22063_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22064_));
AND2X2 AND2X2_11231 ( .A(u2__abc_52155_new_n22061_), .B(u2__abc_52155_new_n22064_), .Y(u2__abc_52155_new_n22065_));
AND2X2 AND2X2_11232 ( .A(u2__abc_52155_new_n22066_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__250_));
AND2X2 AND2X2_11233 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_250_), .Y(u2__abc_52155_new_n22068_));
AND2X2 AND2X2_11234 ( .A(u2__abc_52155_new_n22058_), .B(u2_o_249_), .Y(u2__abc_52155_new_n22069_));
AND2X2 AND2X2_11235 ( .A(u2__abc_52155_new_n22070_), .B(u2__abc_52155_new_n22071_), .Y(u2__abc_52155_new_n22072_));
AND2X2 AND2X2_11236 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4342_), .Y(u2__abc_52155_new_n22074_));
AND2X2 AND2X2_11237 ( .A(u2__abc_52155_new_n22075_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22076_));
AND2X2 AND2X2_11238 ( .A(u2__abc_52155_new_n22073_), .B(u2__abc_52155_new_n22076_), .Y(u2__abc_52155_new_n22077_));
AND2X2 AND2X2_11239 ( .A(u2__abc_52155_new_n22078_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__251_));
AND2X2 AND2X2_1124 ( .A(u2__abc_52155_new_n4311_), .B(u2_remHi_249_), .Y(u2__abc_52155_new_n4312_));
AND2X2 AND2X2_11240 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_251_), .Y(u2__abc_52155_new_n22080_));
AND2X2 AND2X2_11241 ( .A(u2__abc_52155_new_n22069_), .B(u2_o_250_), .Y(u2__abc_52155_new_n22082_));
AND2X2 AND2X2_11242 ( .A(u2__abc_52155_new_n22083_), .B(u2__abc_52155_new_n22081_), .Y(u2__abc_52155_new_n22084_));
AND2X2 AND2X2_11243 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4335_), .Y(u2__abc_52155_new_n22086_));
AND2X2 AND2X2_11244 ( .A(u2__abc_52155_new_n22087_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22088_));
AND2X2 AND2X2_11245 ( .A(u2__abc_52155_new_n22085_), .B(u2__abc_52155_new_n22088_), .Y(u2__abc_52155_new_n22089_));
AND2X2 AND2X2_11246 ( .A(u2__abc_52155_new_n22090_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__252_));
AND2X2 AND2X2_11247 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_252_), .Y(u2__abc_52155_new_n22092_));
AND2X2 AND2X2_11248 ( .A(u2__abc_52155_new_n22082_), .B(u2_o_251_), .Y(u2__abc_52155_new_n22093_));
AND2X2 AND2X2_11249 ( .A(u2__abc_52155_new_n22094_), .B(u2__abc_52155_new_n22095_), .Y(u2__abc_52155_new_n22096_));
AND2X2 AND2X2_1125 ( .A(u2__abc_52155_new_n4314_), .B(u2_o_249_), .Y(u2__abc_52155_new_n4315_));
AND2X2 AND2X2_11250 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4320_), .Y(u2__abc_52155_new_n22098_));
AND2X2 AND2X2_11251 ( .A(u2__abc_52155_new_n22099_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22100_));
AND2X2 AND2X2_11252 ( .A(u2__abc_52155_new_n22097_), .B(u2__abc_52155_new_n22100_), .Y(u2__abc_52155_new_n22101_));
AND2X2 AND2X2_11253 ( .A(u2__abc_52155_new_n22102_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__253_));
AND2X2 AND2X2_11254 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_253_), .Y(u2__abc_52155_new_n22104_));
AND2X2 AND2X2_11255 ( .A(u2__abc_52155_new_n22093_), .B(u2_o_252_), .Y(u2__abc_52155_new_n22106_));
AND2X2 AND2X2_11256 ( .A(u2__abc_52155_new_n22107_), .B(u2__abc_52155_new_n22105_), .Y(u2__abc_52155_new_n22108_));
AND2X2 AND2X2_11257 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4330_), .Y(u2__abc_52155_new_n22110_));
AND2X2 AND2X2_11258 ( .A(u2__abc_52155_new_n22111_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22112_));
AND2X2 AND2X2_11259 ( .A(u2__abc_52155_new_n22109_), .B(u2__abc_52155_new_n22112_), .Y(u2__abc_52155_new_n22113_));
AND2X2 AND2X2_1126 ( .A(u2__abc_52155_new_n4313_), .B(u2__abc_52155_new_n4316_), .Y(u2__abc_52155_new_n4317_));
AND2X2 AND2X2_11260 ( .A(u2__abc_52155_new_n22114_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__254_));
AND2X2 AND2X2_11261 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_254_), .Y(u2__abc_52155_new_n22116_));
AND2X2 AND2X2_11262 ( .A(u2__abc_52155_new_n22106_), .B(u2_o_253_), .Y(u2__abc_52155_new_n22117_));
AND2X2 AND2X2_11263 ( .A(u2__abc_52155_new_n22118_), .B(u2__abc_52155_new_n22119_), .Y(u2__abc_52155_new_n22120_));
AND2X2 AND2X2_11264 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6542_), .Y(u2__abc_52155_new_n22122_));
AND2X2 AND2X2_11265 ( .A(u2__abc_52155_new_n22123_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22124_));
AND2X2 AND2X2_11266 ( .A(u2__abc_52155_new_n22121_), .B(u2__abc_52155_new_n22124_), .Y(u2__abc_52155_new_n22125_));
AND2X2 AND2X2_11267 ( .A(u2__abc_52155_new_n22126_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__255_));
AND2X2 AND2X2_11268 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_255_), .Y(u2__abc_52155_new_n22128_));
AND2X2 AND2X2_11269 ( .A(u2__abc_52155_new_n22117_), .B(u2_o_254_), .Y(u2__abc_52155_new_n22130_));
AND2X2 AND2X2_1127 ( .A(u2__abc_52155_new_n4310_), .B(u2__abc_52155_new_n4317_), .Y(u2__abc_52155_new_n4318_));
AND2X2 AND2X2_11270 ( .A(u2__abc_52155_new_n22131_), .B(u2__abc_52155_new_n22129_), .Y(u2__abc_52155_new_n22132_));
AND2X2 AND2X2_11271 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6549_), .Y(u2__abc_52155_new_n22134_));
AND2X2 AND2X2_11272 ( .A(u2__abc_52155_new_n22135_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22136_));
AND2X2 AND2X2_11273 ( .A(u2__abc_52155_new_n22133_), .B(u2__abc_52155_new_n22136_), .Y(u2__abc_52155_new_n22137_));
AND2X2 AND2X2_11274 ( .A(u2__abc_52155_new_n22138_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__256_));
AND2X2 AND2X2_11275 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_256_), .Y(u2__abc_52155_new_n22140_));
AND2X2 AND2X2_11276 ( .A(u2__abc_52155_new_n22130_), .B(u2_o_255_), .Y(u2__abc_52155_new_n22141_));
AND2X2 AND2X2_11277 ( .A(u2__abc_52155_new_n22142_), .B(u2__abc_52155_new_n22143_), .Y(u2__abc_52155_new_n22144_));
AND2X2 AND2X2_11278 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6554_), .Y(u2__abc_52155_new_n22146_));
AND2X2 AND2X2_11279 ( .A(u2__abc_52155_new_n22147_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22148_));
AND2X2 AND2X2_1128 ( .A(u2__abc_52155_new_n4303_), .B(u2__abc_52155_new_n4318_), .Y(u2__abc_52155_new_n4319_));
AND2X2 AND2X2_11280 ( .A(u2__abc_52155_new_n22145_), .B(u2__abc_52155_new_n22148_), .Y(u2__abc_52155_new_n22149_));
AND2X2 AND2X2_11281 ( .A(u2__abc_52155_new_n22150_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__257_));
AND2X2 AND2X2_11282 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_257_), .Y(u2__abc_52155_new_n22152_));
AND2X2 AND2X2_11283 ( .A(u2__abc_52155_new_n22141_), .B(u2_o_256_), .Y(u2__abc_52155_new_n22154_));
AND2X2 AND2X2_11284 ( .A(u2__abc_52155_new_n22155_), .B(u2__abc_52155_new_n22153_), .Y(u2__abc_52155_new_n22156_));
AND2X2 AND2X2_11285 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6561_), .Y(u2__abc_52155_new_n22158_));
AND2X2 AND2X2_11286 ( .A(u2__abc_52155_new_n22159_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22160_));
AND2X2 AND2X2_11287 ( .A(u2__abc_52155_new_n22157_), .B(u2__abc_52155_new_n22160_), .Y(u2__abc_52155_new_n22161_));
AND2X2 AND2X2_11288 ( .A(u2__abc_52155_new_n22162_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__258_));
AND2X2 AND2X2_11289 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_258_), .Y(u2__abc_52155_new_n22164_));
AND2X2 AND2X2_1129 ( .A(u2__abc_52155_new_n4320_), .B(u2_remHi_252_), .Y(u2__abc_52155_new_n4321_));
AND2X2 AND2X2_11290 ( .A(u2__abc_52155_new_n22154_), .B(u2_o_257_), .Y(u2__abc_52155_new_n22166_));
AND2X2 AND2X2_11291 ( .A(u2__abc_52155_new_n22167_), .B(u2__abc_52155_new_n22165_), .Y(u2__abc_52155_new_n22168_));
AND2X2 AND2X2_11292 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6585_), .Y(u2__abc_52155_new_n22170_));
AND2X2 AND2X2_11293 ( .A(u2__abc_52155_new_n22171_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22172_));
AND2X2 AND2X2_11294 ( .A(u2__abc_52155_new_n22169_), .B(u2__abc_52155_new_n22172_), .Y(u2__abc_52155_new_n22173_));
AND2X2 AND2X2_11295 ( .A(u2__abc_52155_new_n22174_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__259_));
AND2X2 AND2X2_11296 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_259_), .Y(u2__abc_52155_new_n22176_));
AND2X2 AND2X2_11297 ( .A(u2__abc_52155_new_n22166_), .B(u2_o_258_), .Y(u2__abc_52155_new_n22178_));
AND2X2 AND2X2_11298 ( .A(u2__abc_52155_new_n22179_), .B(u2__abc_52155_new_n22177_), .Y(u2__abc_52155_new_n22180_));
AND2X2 AND2X2_11299 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6592_), .Y(u2__abc_52155_new_n22182_));
AND2X2 AND2X2_113 ( .A(_abc_73687_new_n939_), .B(_abc_73687_new_n938_), .Y(\o[148] ));
AND2X2 AND2X2_1130 ( .A(u2__abc_52155_new_n4323_), .B(u2_o_252_), .Y(u2__abc_52155_new_n4324_));
AND2X2 AND2X2_11300 ( .A(u2__abc_52155_new_n22183_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22184_));
AND2X2 AND2X2_11301 ( .A(u2__abc_52155_new_n22181_), .B(u2__abc_52155_new_n22184_), .Y(u2__abc_52155_new_n22185_));
AND2X2 AND2X2_11302 ( .A(u2__abc_52155_new_n22186_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__260_));
AND2X2 AND2X2_11303 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_260_), .Y(u2__abc_52155_new_n22188_));
AND2X2 AND2X2_11304 ( .A(u2__abc_52155_new_n22178_), .B(u2_o_259_), .Y(u2__abc_52155_new_n22189_));
AND2X2 AND2X2_11305 ( .A(u2__abc_52155_new_n22190_), .B(u2__abc_52155_new_n22191_), .Y(u2__abc_52155_new_n22192_));
AND2X2 AND2X2_11306 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6570_), .Y(u2__abc_52155_new_n22194_));
AND2X2 AND2X2_11307 ( .A(u2__abc_52155_new_n22195_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22196_));
AND2X2 AND2X2_11308 ( .A(u2__abc_52155_new_n22193_), .B(u2__abc_52155_new_n22196_), .Y(u2__abc_52155_new_n22197_));
AND2X2 AND2X2_11309 ( .A(u2__abc_52155_new_n22198_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__261_));
AND2X2 AND2X2_1131 ( .A(u2__abc_52155_new_n4322_), .B(u2__abc_52155_new_n4325_), .Y(u2__abc_52155_new_n4326_));
AND2X2 AND2X2_11310 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_261_), .Y(u2__abc_52155_new_n22200_));
AND2X2 AND2X2_11311 ( .A(u2__abc_52155_new_n22189_), .B(u2_o_260_), .Y(u2__abc_52155_new_n22202_));
AND2X2 AND2X2_11312 ( .A(u2__abc_52155_new_n22203_), .B(u2__abc_52155_new_n22201_), .Y(u2__abc_52155_new_n22204_));
AND2X2 AND2X2_11313 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6577_), .Y(u2__abc_52155_new_n22206_));
AND2X2 AND2X2_11314 ( .A(u2__abc_52155_new_n22207_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22208_));
AND2X2 AND2X2_11315 ( .A(u2__abc_52155_new_n22205_), .B(u2__abc_52155_new_n22208_), .Y(u2__abc_52155_new_n22209_));
AND2X2 AND2X2_11316 ( .A(u2__abc_52155_new_n22210_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__262_));
AND2X2 AND2X2_11317 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_262_), .Y(u2__abc_52155_new_n22212_));
AND2X2 AND2X2_11318 ( .A(u2__abc_52155_new_n22202_), .B(u2_o_261_), .Y(u2__abc_52155_new_n22213_));
AND2X2 AND2X2_11319 ( .A(u2__abc_52155_new_n22214_), .B(u2__abc_52155_new_n22215_), .Y(u2__abc_52155_new_n22216_));
AND2X2 AND2X2_1132 ( .A(u2__abc_52155_new_n4327_), .B(u2_o_253_), .Y(u2__abc_52155_new_n4328_));
AND2X2 AND2X2_11320 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6525_), .Y(u2__abc_52155_new_n22218_));
AND2X2 AND2X2_11321 ( .A(u2__abc_52155_new_n22219_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22220_));
AND2X2 AND2X2_11322 ( .A(u2__abc_52155_new_n22217_), .B(u2__abc_52155_new_n22220_), .Y(u2__abc_52155_new_n22221_));
AND2X2 AND2X2_11323 ( .A(u2__abc_52155_new_n22222_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__263_));
AND2X2 AND2X2_11324 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_263_), .Y(u2__abc_52155_new_n22224_));
AND2X2 AND2X2_11325 ( .A(u2__abc_52155_new_n22213_), .B(u2_o_262_), .Y(u2__abc_52155_new_n22226_));
AND2X2 AND2X2_11326 ( .A(u2__abc_52155_new_n22227_), .B(u2__abc_52155_new_n22225_), .Y(u2__abc_52155_new_n22228_));
AND2X2 AND2X2_11327 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6532_), .Y(u2__abc_52155_new_n22230_));
AND2X2 AND2X2_11328 ( .A(u2__abc_52155_new_n22231_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22232_));
AND2X2 AND2X2_11329 ( .A(u2__abc_52155_new_n22229_), .B(u2__abc_52155_new_n22232_), .Y(u2__abc_52155_new_n22233_));
AND2X2 AND2X2_1133 ( .A(u2__abc_52155_new_n4330_), .B(u2_remHi_253_), .Y(u2__abc_52155_new_n4331_));
AND2X2 AND2X2_11330 ( .A(u2__abc_52155_new_n22234_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__264_));
AND2X2 AND2X2_11331 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_264_), .Y(u2__abc_52155_new_n22236_));
AND2X2 AND2X2_11332 ( .A(u2__abc_52155_new_n22226_), .B(u2_o_263_), .Y(u2__abc_52155_new_n22238_));
AND2X2 AND2X2_11333 ( .A(u2__abc_52155_new_n22239_), .B(u2__abc_52155_new_n22237_), .Y(u2__abc_52155_new_n22240_));
AND2X2 AND2X2_11334 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6507_), .Y(u2__abc_52155_new_n22242_));
AND2X2 AND2X2_11335 ( .A(u2__abc_52155_new_n22243_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22244_));
AND2X2 AND2X2_11336 ( .A(u2__abc_52155_new_n22241_), .B(u2__abc_52155_new_n22244_), .Y(u2__abc_52155_new_n22245_));
AND2X2 AND2X2_11337 ( .A(u2__abc_52155_new_n22246_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__265_));
AND2X2 AND2X2_11338 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_265_), .Y(u2__abc_52155_new_n22248_));
AND2X2 AND2X2_11339 ( .A(u2__abc_52155_new_n22238_), .B(u2_o_264_), .Y(u2__abc_52155_new_n22250_));
AND2X2 AND2X2_1134 ( .A(u2__abc_52155_new_n4329_), .B(u2__abc_52155_new_n4332_), .Y(u2__abc_52155_new_n4333_));
AND2X2 AND2X2_11340 ( .A(u2__abc_52155_new_n22251_), .B(u2__abc_52155_new_n22249_), .Y(u2__abc_52155_new_n22252_));
AND2X2 AND2X2_11341 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6514_), .Y(u2__abc_52155_new_n22254_));
AND2X2 AND2X2_11342 ( .A(u2__abc_52155_new_n22255_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22256_));
AND2X2 AND2X2_11343 ( .A(u2__abc_52155_new_n22253_), .B(u2__abc_52155_new_n22256_), .Y(u2__abc_52155_new_n22257_));
AND2X2 AND2X2_11344 ( .A(u2__abc_52155_new_n22258_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__266_));
AND2X2 AND2X2_11345 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_266_), .Y(u2__abc_52155_new_n22260_));
AND2X2 AND2X2_11346 ( .A(u2__abc_52155_new_n22250_), .B(u2_o_265_), .Y(u2__abc_52155_new_n22261_));
AND2X2 AND2X2_11347 ( .A(u2__abc_52155_new_n22262_), .B(u2__abc_52155_new_n22263_), .Y(u2__abc_52155_new_n22264_));
AND2X2 AND2X2_11348 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6491_), .Y(u2__abc_52155_new_n22266_));
AND2X2 AND2X2_11349 ( .A(u2__abc_52155_new_n22267_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22268_));
AND2X2 AND2X2_1135 ( .A(u2__abc_52155_new_n4326_), .B(u2__abc_52155_new_n4333_), .Y(u2__abc_52155_new_n4334_));
AND2X2 AND2X2_11350 ( .A(u2__abc_52155_new_n22265_), .B(u2__abc_52155_new_n22268_), .Y(u2__abc_52155_new_n22269_));
AND2X2 AND2X2_11351 ( .A(u2__abc_52155_new_n22270_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__267_));
AND2X2 AND2X2_11352 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_267_), .Y(u2__abc_52155_new_n22272_));
AND2X2 AND2X2_11353 ( .A(u2__abc_52155_new_n22261_), .B(u2_o_266_), .Y(u2__abc_52155_new_n22274_));
AND2X2 AND2X2_11354 ( .A(u2__abc_52155_new_n22275_), .B(u2__abc_52155_new_n22273_), .Y(u2__abc_52155_new_n22276_));
AND2X2 AND2X2_11355 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6498_), .Y(u2__abc_52155_new_n22278_));
AND2X2 AND2X2_11356 ( .A(u2__abc_52155_new_n22279_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22280_));
AND2X2 AND2X2_11357 ( .A(u2__abc_52155_new_n22277_), .B(u2__abc_52155_new_n22280_), .Y(u2__abc_52155_new_n22281_));
AND2X2 AND2X2_11358 ( .A(u2__abc_52155_new_n22282_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__268_));
AND2X2 AND2X2_11359 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_268_), .Y(u2__abc_52155_new_n22284_));
AND2X2 AND2X2_1136 ( .A(u2__abc_52155_new_n4335_), .B(u2_remHi_251_), .Y(u2__abc_52155_new_n4336_));
AND2X2 AND2X2_11360 ( .A(u2__abc_52155_new_n22274_), .B(u2_o_267_), .Y(u2__abc_52155_new_n22286_));
AND2X2 AND2X2_11361 ( .A(u2__abc_52155_new_n22287_), .B(u2__abc_52155_new_n22285_), .Y(u2__abc_52155_new_n22288_));
AND2X2 AND2X2_11362 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6479_), .Y(u2__abc_52155_new_n22290_));
AND2X2 AND2X2_11363 ( .A(u2__abc_52155_new_n22291_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22292_));
AND2X2 AND2X2_11364 ( .A(u2__abc_52155_new_n22289_), .B(u2__abc_52155_new_n22292_), .Y(u2__abc_52155_new_n22293_));
AND2X2 AND2X2_11365 ( .A(u2__abc_52155_new_n22294_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__269_));
AND2X2 AND2X2_11366 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_269_), .Y(u2__abc_52155_new_n22296_));
AND2X2 AND2X2_11367 ( .A(u2__abc_52155_new_n22286_), .B(u2_o_268_), .Y(u2__abc_52155_new_n22298_));
AND2X2 AND2X2_11368 ( .A(u2__abc_52155_new_n22299_), .B(u2__abc_52155_new_n22297_), .Y(u2__abc_52155_new_n22300_));
AND2X2 AND2X2_11369 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6486_), .Y(u2__abc_52155_new_n22302_));
AND2X2 AND2X2_1137 ( .A(u2__abc_52155_new_n4338_), .B(u2_o_251_), .Y(u2__abc_52155_new_n4339_));
AND2X2 AND2X2_11370 ( .A(u2__abc_52155_new_n22303_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22304_));
AND2X2 AND2X2_11371 ( .A(u2__abc_52155_new_n22301_), .B(u2__abc_52155_new_n22304_), .Y(u2__abc_52155_new_n22305_));
AND2X2 AND2X2_11372 ( .A(u2__abc_52155_new_n22306_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__270_));
AND2X2 AND2X2_11373 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_270_), .Y(u2__abc_52155_new_n22308_));
AND2X2 AND2X2_11374 ( .A(u2__abc_52155_new_n22298_), .B(u2_o_269_), .Y(u2__abc_52155_new_n22309_));
AND2X2 AND2X2_11375 ( .A(u2__abc_52155_new_n22310_), .B(u2__abc_52155_new_n22311_), .Y(u2__abc_52155_new_n22312_));
AND2X2 AND2X2_11376 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6427_), .Y(u2__abc_52155_new_n22314_));
AND2X2 AND2X2_11377 ( .A(u2__abc_52155_new_n22315_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22316_));
AND2X2 AND2X2_11378 ( .A(u2__abc_52155_new_n22313_), .B(u2__abc_52155_new_n22316_), .Y(u2__abc_52155_new_n22317_));
AND2X2 AND2X2_11379 ( .A(u2__abc_52155_new_n22318_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__271_));
AND2X2 AND2X2_1138 ( .A(u2__abc_52155_new_n4337_), .B(u2__abc_52155_new_n4340_), .Y(u2__abc_52155_new_n4341_));
AND2X2 AND2X2_11380 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_271_), .Y(u2__abc_52155_new_n22320_));
AND2X2 AND2X2_11381 ( .A(u2__abc_52155_new_n22309_), .B(u2_o_270_), .Y(u2__abc_52155_new_n22322_));
AND2X2 AND2X2_11382 ( .A(u2__abc_52155_new_n22323_), .B(u2__abc_52155_new_n22321_), .Y(u2__abc_52155_new_n22324_));
AND2X2 AND2X2_11383 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6434_), .Y(u2__abc_52155_new_n22326_));
AND2X2 AND2X2_11384 ( .A(u2__abc_52155_new_n22327_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22328_));
AND2X2 AND2X2_11385 ( .A(u2__abc_52155_new_n22325_), .B(u2__abc_52155_new_n22328_), .Y(u2__abc_52155_new_n22329_));
AND2X2 AND2X2_11386 ( .A(u2__abc_52155_new_n22330_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__272_));
AND2X2 AND2X2_11387 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_272_), .Y(u2__abc_52155_new_n22332_));
AND2X2 AND2X2_11388 ( .A(u2__abc_52155_new_n22322_), .B(u2_o_271_), .Y(u2__abc_52155_new_n22334_));
AND2X2 AND2X2_11389 ( .A(u2__abc_52155_new_n22335_), .B(u2__abc_52155_new_n22333_), .Y(u2__abc_52155_new_n22336_));
AND2X2 AND2X2_1139 ( .A(u2__abc_52155_new_n4342_), .B(u2_remHi_250_), .Y(u2__abc_52155_new_n4343_));
AND2X2 AND2X2_11390 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6412_), .Y(u2__abc_52155_new_n22338_));
AND2X2 AND2X2_11391 ( .A(u2__abc_52155_new_n22339_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22340_));
AND2X2 AND2X2_11392 ( .A(u2__abc_52155_new_n22337_), .B(u2__abc_52155_new_n22340_), .Y(u2__abc_52155_new_n22341_));
AND2X2 AND2X2_11393 ( .A(u2__abc_52155_new_n22342_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__273_));
AND2X2 AND2X2_11394 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_273_), .Y(u2__abc_52155_new_n22344_));
AND2X2 AND2X2_11395 ( .A(u2__abc_52155_new_n22334_), .B(u2_o_272_), .Y(u2__abc_52155_new_n22346_));
AND2X2 AND2X2_11396 ( .A(u2__abc_52155_new_n22347_), .B(u2__abc_52155_new_n22345_), .Y(u2__abc_52155_new_n22348_));
AND2X2 AND2X2_11397 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6419_), .Y(u2__abc_52155_new_n22350_));
AND2X2 AND2X2_11398 ( .A(u2__abc_52155_new_n22351_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22352_));
AND2X2 AND2X2_11399 ( .A(u2__abc_52155_new_n22349_), .B(u2__abc_52155_new_n22352_), .Y(u2__abc_52155_new_n22353_));
AND2X2 AND2X2_114 ( .A(_abc_73687_new_n942_), .B(_abc_73687_new_n941_), .Y(\o[149] ));
AND2X2 AND2X2_1140 ( .A(u2__abc_52155_new_n4345_), .B(u2_o_250_), .Y(u2__abc_52155_new_n4346_));
AND2X2 AND2X2_11400 ( .A(u2__abc_52155_new_n22354_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__274_));
AND2X2 AND2X2_11401 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_274_), .Y(u2__abc_52155_new_n22356_));
AND2X2 AND2X2_11402 ( .A(u2__abc_52155_new_n22346_), .B(u2_o_273_), .Y(u2__abc_52155_new_n22357_));
AND2X2 AND2X2_11403 ( .A(u2__abc_52155_new_n22358_), .B(u2__abc_52155_new_n22359_), .Y(u2__abc_52155_new_n22360_));
AND2X2 AND2X2_11404 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6458_), .Y(u2__abc_52155_new_n22362_));
AND2X2 AND2X2_11405 ( .A(u2__abc_52155_new_n22363_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22364_));
AND2X2 AND2X2_11406 ( .A(u2__abc_52155_new_n22361_), .B(u2__abc_52155_new_n22364_), .Y(u2__abc_52155_new_n22365_));
AND2X2 AND2X2_11407 ( .A(u2__abc_52155_new_n22366_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__275_));
AND2X2 AND2X2_11408 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_275_), .Y(u2__abc_52155_new_n22368_));
AND2X2 AND2X2_11409 ( .A(u2__abc_52155_new_n22357_), .B(u2_o_274_), .Y(u2__abc_52155_new_n22370_));
AND2X2 AND2X2_1141 ( .A(u2__abc_52155_new_n4344_), .B(u2__abc_52155_new_n4347_), .Y(u2__abc_52155_new_n4348_));
AND2X2 AND2X2_11410 ( .A(u2__abc_52155_new_n22371_), .B(u2__abc_52155_new_n22369_), .Y(u2__abc_52155_new_n22372_));
AND2X2 AND2X2_11411 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6465_), .Y(u2__abc_52155_new_n22374_));
AND2X2 AND2X2_11412 ( .A(u2__abc_52155_new_n22375_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22376_));
AND2X2 AND2X2_11413 ( .A(u2__abc_52155_new_n22373_), .B(u2__abc_52155_new_n22376_), .Y(u2__abc_52155_new_n22377_));
AND2X2 AND2X2_11414 ( .A(u2__abc_52155_new_n22378_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__276_));
AND2X2 AND2X2_11415 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_276_), .Y(u2__abc_52155_new_n22380_));
AND2X2 AND2X2_11416 ( .A(u2__abc_52155_new_n22370_), .B(u2_o_275_), .Y(u2__abc_52155_new_n22382_));
AND2X2 AND2X2_11417 ( .A(u2__abc_52155_new_n22383_), .B(u2__abc_52155_new_n22381_), .Y(u2__abc_52155_new_n22384_));
AND2X2 AND2X2_11418 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6443_), .Y(u2__abc_52155_new_n22386_));
AND2X2 AND2X2_11419 ( .A(u2__abc_52155_new_n22387_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22388_));
AND2X2 AND2X2_1142 ( .A(u2__abc_52155_new_n4341_), .B(u2__abc_52155_new_n4348_), .Y(u2__abc_52155_new_n4349_));
AND2X2 AND2X2_11420 ( .A(u2__abc_52155_new_n22385_), .B(u2__abc_52155_new_n22388_), .Y(u2__abc_52155_new_n22389_));
AND2X2 AND2X2_11421 ( .A(u2__abc_52155_new_n22390_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__277_));
AND2X2 AND2X2_11422 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_277_), .Y(u2__abc_52155_new_n22392_));
AND2X2 AND2X2_11423 ( .A(u2__abc_52155_new_n22382_), .B(u2_o_276_), .Y(u2__abc_52155_new_n22394_));
AND2X2 AND2X2_11424 ( .A(u2__abc_52155_new_n22395_), .B(u2__abc_52155_new_n22393_), .Y(u2__abc_52155_new_n22396_));
AND2X2 AND2X2_11425 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6450_), .Y(u2__abc_52155_new_n22398_));
AND2X2 AND2X2_11426 ( .A(u2__abc_52155_new_n22399_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22400_));
AND2X2 AND2X2_11427 ( .A(u2__abc_52155_new_n22397_), .B(u2__abc_52155_new_n22400_), .Y(u2__abc_52155_new_n22401_));
AND2X2 AND2X2_11428 ( .A(u2__abc_52155_new_n22402_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__278_));
AND2X2 AND2X2_11429 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_278_), .Y(u2__abc_52155_new_n22404_));
AND2X2 AND2X2_1143 ( .A(u2__abc_52155_new_n4334_), .B(u2__abc_52155_new_n4349_), .Y(u2__abc_52155_new_n4350_));
AND2X2 AND2X2_11430 ( .A(u2__abc_52155_new_n22394_), .B(u2_o_277_), .Y(u2__abc_52155_new_n22405_));
AND2X2 AND2X2_11431 ( .A(u2__abc_52155_new_n22406_), .B(u2__abc_52155_new_n22407_), .Y(u2__abc_52155_new_n22408_));
AND2X2 AND2X2_11432 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6364_), .Y(u2__abc_52155_new_n22410_));
AND2X2 AND2X2_11433 ( .A(u2__abc_52155_new_n22411_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22412_));
AND2X2 AND2X2_11434 ( .A(u2__abc_52155_new_n22409_), .B(u2__abc_52155_new_n22412_), .Y(u2__abc_52155_new_n22413_));
AND2X2 AND2X2_11435 ( .A(u2__abc_52155_new_n22414_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__279_));
AND2X2 AND2X2_11436 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_279_), .Y(u2__abc_52155_new_n22416_));
AND2X2 AND2X2_11437 ( .A(u2__abc_52155_new_n22405_), .B(u2_o_278_), .Y(u2__abc_52155_new_n22418_));
AND2X2 AND2X2_11438 ( .A(u2__abc_52155_new_n22419_), .B(u2__abc_52155_new_n22417_), .Y(u2__abc_52155_new_n22420_));
AND2X2 AND2X2_11439 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6371_), .Y(u2__abc_52155_new_n22422_));
AND2X2 AND2X2_1144 ( .A(u2__abc_52155_new_n4319_), .B(u2__abc_52155_new_n4350_), .Y(u2__abc_52155_new_n4351_));
AND2X2 AND2X2_11440 ( .A(u2__abc_52155_new_n22423_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22424_));
AND2X2 AND2X2_11441 ( .A(u2__abc_52155_new_n22421_), .B(u2__abc_52155_new_n22424_), .Y(u2__abc_52155_new_n22425_));
AND2X2 AND2X2_11442 ( .A(u2__abc_52155_new_n22426_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__280_));
AND2X2 AND2X2_11443 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_280_), .Y(u2__abc_52155_new_n22428_));
AND2X2 AND2X2_11444 ( .A(u2__abc_52155_new_n22418_), .B(u2_o_279_), .Y(u2__abc_52155_new_n22430_));
AND2X2 AND2X2_11445 ( .A(u2__abc_52155_new_n22431_), .B(u2__abc_52155_new_n22429_), .Y(u2__abc_52155_new_n22432_));
AND2X2 AND2X2_11446 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6349_), .Y(u2__abc_52155_new_n22434_));
AND2X2 AND2X2_11447 ( .A(u2__abc_52155_new_n22435_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22436_));
AND2X2 AND2X2_11448 ( .A(u2__abc_52155_new_n22433_), .B(u2__abc_52155_new_n22436_), .Y(u2__abc_52155_new_n22437_));
AND2X2 AND2X2_11449 ( .A(u2__abc_52155_new_n22438_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__281_));
AND2X2 AND2X2_1145 ( .A(u2__abc_52155_new_n4352_), .B(u2_remHi_238_), .Y(u2__abc_52155_new_n4353_));
AND2X2 AND2X2_11450 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_281_), .Y(u2__abc_52155_new_n22440_));
AND2X2 AND2X2_11451 ( .A(u2__abc_52155_new_n22430_), .B(u2_o_280_), .Y(u2__abc_52155_new_n22442_));
AND2X2 AND2X2_11452 ( .A(u2__abc_52155_new_n22443_), .B(u2__abc_52155_new_n22441_), .Y(u2__abc_52155_new_n22444_));
AND2X2 AND2X2_11453 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6356_), .Y(u2__abc_52155_new_n22446_));
AND2X2 AND2X2_11454 ( .A(u2__abc_52155_new_n22447_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22448_));
AND2X2 AND2X2_11455 ( .A(u2__abc_52155_new_n22445_), .B(u2__abc_52155_new_n22448_), .Y(u2__abc_52155_new_n22449_));
AND2X2 AND2X2_11456 ( .A(u2__abc_52155_new_n22450_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__282_));
AND2X2 AND2X2_11457 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_282_), .Y(u2__abc_52155_new_n22452_));
AND2X2 AND2X2_11458 ( .A(u2__abc_52155_new_n22442_), .B(u2_o_281_), .Y(u2__abc_52155_new_n22453_));
AND2X2 AND2X2_11459 ( .A(u2__abc_52155_new_n22454_), .B(u2__abc_52155_new_n22455_), .Y(u2__abc_52155_new_n22456_));
AND2X2 AND2X2_1146 ( .A(u2__abc_52155_new_n4355_), .B(u2_o_238_), .Y(u2__abc_52155_new_n4356_));
AND2X2 AND2X2_11460 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6395_), .Y(u2__abc_52155_new_n22458_));
AND2X2 AND2X2_11461 ( .A(u2__abc_52155_new_n22459_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22460_));
AND2X2 AND2X2_11462 ( .A(u2__abc_52155_new_n22457_), .B(u2__abc_52155_new_n22460_), .Y(u2__abc_52155_new_n22461_));
AND2X2 AND2X2_11463 ( .A(u2__abc_52155_new_n22462_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__283_));
AND2X2 AND2X2_11464 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_283_), .Y(u2__abc_52155_new_n22464_));
AND2X2 AND2X2_11465 ( .A(u2__abc_52155_new_n22453_), .B(u2_o_282_), .Y(u2__abc_52155_new_n22466_));
AND2X2 AND2X2_11466 ( .A(u2__abc_52155_new_n22467_), .B(u2__abc_52155_new_n22465_), .Y(u2__abc_52155_new_n22468_));
AND2X2 AND2X2_11467 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6402_), .Y(u2__abc_52155_new_n22470_));
AND2X2 AND2X2_11468 ( .A(u2__abc_52155_new_n22471_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22472_));
AND2X2 AND2X2_11469 ( .A(u2__abc_52155_new_n22469_), .B(u2__abc_52155_new_n22472_), .Y(u2__abc_52155_new_n22473_));
AND2X2 AND2X2_1147 ( .A(u2__abc_52155_new_n4354_), .B(u2__abc_52155_new_n4357_), .Y(u2__abc_52155_new_n4358_));
AND2X2 AND2X2_11470 ( .A(u2__abc_52155_new_n22474_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__284_));
AND2X2 AND2X2_11471 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_284_), .Y(u2__abc_52155_new_n22476_));
AND2X2 AND2X2_11472 ( .A(u2__abc_52155_new_n22466_), .B(u2_o_283_), .Y(u2__abc_52155_new_n22478_));
AND2X2 AND2X2_11473 ( .A(u2__abc_52155_new_n22479_), .B(u2__abc_52155_new_n22477_), .Y(u2__abc_52155_new_n22480_));
AND2X2 AND2X2_11474 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6380_), .Y(u2__abc_52155_new_n22482_));
AND2X2 AND2X2_11475 ( .A(u2__abc_52155_new_n22483_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22484_));
AND2X2 AND2X2_11476 ( .A(u2__abc_52155_new_n22481_), .B(u2__abc_52155_new_n22484_), .Y(u2__abc_52155_new_n22485_));
AND2X2 AND2X2_11477 ( .A(u2__abc_52155_new_n22486_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__285_));
AND2X2 AND2X2_11478 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_285_), .Y(u2__abc_52155_new_n22488_));
AND2X2 AND2X2_11479 ( .A(u2__abc_52155_new_n22478_), .B(u2_o_284_), .Y(u2__abc_52155_new_n22490_));
AND2X2 AND2X2_1148 ( .A(u2__abc_52155_new_n4359_), .B(u2_remHi_239_), .Y(u2__abc_52155_new_n4360_));
AND2X2 AND2X2_11480 ( .A(u2__abc_52155_new_n22491_), .B(u2__abc_52155_new_n22489_), .Y(u2__abc_52155_new_n22492_));
AND2X2 AND2X2_11481 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6387_), .Y(u2__abc_52155_new_n22494_));
AND2X2 AND2X2_11482 ( .A(u2__abc_52155_new_n22495_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22496_));
AND2X2 AND2X2_11483 ( .A(u2__abc_52155_new_n22493_), .B(u2__abc_52155_new_n22496_), .Y(u2__abc_52155_new_n22497_));
AND2X2 AND2X2_11484 ( .A(u2__abc_52155_new_n22498_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__286_));
AND2X2 AND2X2_11485 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_286_), .Y(u2__abc_52155_new_n22500_));
AND2X2 AND2X2_11486 ( .A(u2__abc_52155_new_n22490_), .B(u2_o_285_), .Y(u2__abc_52155_new_n22501_));
AND2X2 AND2X2_11487 ( .A(u2__abc_52155_new_n22502_), .B(u2__abc_52155_new_n22503_), .Y(u2__abc_52155_new_n22504_));
AND2X2 AND2X2_11488 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6299_), .Y(u2__abc_52155_new_n22506_));
AND2X2 AND2X2_11489 ( .A(u2__abc_52155_new_n22507_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22508_));
AND2X2 AND2X2_1149 ( .A(u2__abc_52155_new_n4362_), .B(u2_o_239_), .Y(u2__abc_52155_new_n4363_));
AND2X2 AND2X2_11490 ( .A(u2__abc_52155_new_n22505_), .B(u2__abc_52155_new_n22508_), .Y(u2__abc_52155_new_n22509_));
AND2X2 AND2X2_11491 ( .A(u2__abc_52155_new_n22510_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__287_));
AND2X2 AND2X2_11492 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_287_), .Y(u2__abc_52155_new_n22512_));
AND2X2 AND2X2_11493 ( .A(u2__abc_52155_new_n22501_), .B(u2_o_286_), .Y(u2__abc_52155_new_n22514_));
AND2X2 AND2X2_11494 ( .A(u2__abc_52155_new_n22515_), .B(u2__abc_52155_new_n22513_), .Y(u2__abc_52155_new_n22516_));
AND2X2 AND2X2_11495 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6306_), .Y(u2__abc_52155_new_n22518_));
AND2X2 AND2X2_11496 ( .A(u2__abc_52155_new_n22519_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22520_));
AND2X2 AND2X2_11497 ( .A(u2__abc_52155_new_n22517_), .B(u2__abc_52155_new_n22520_), .Y(u2__abc_52155_new_n22521_));
AND2X2 AND2X2_11498 ( .A(u2__abc_52155_new_n22522_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__288_));
AND2X2 AND2X2_11499 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_288_), .Y(u2__abc_52155_new_n22524_));
AND2X2 AND2X2_115 ( .A(_abc_73687_new_n945_), .B(_abc_73687_new_n944_), .Y(\o[150] ));
AND2X2 AND2X2_1150 ( .A(u2__abc_52155_new_n4361_), .B(u2__abc_52155_new_n4364_), .Y(u2__abc_52155_new_n4365_));
AND2X2 AND2X2_11500 ( .A(u2__abc_52155_new_n22514_), .B(u2_o_287_), .Y(u2__abc_52155_new_n22525_));
AND2X2 AND2X2_11501 ( .A(u2__abc_52155_new_n22526_), .B(u2__abc_52155_new_n22527_), .Y(u2__abc_52155_new_n22528_));
AND2X2 AND2X2_11502 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6284_), .Y(u2__abc_52155_new_n22530_));
AND2X2 AND2X2_11503 ( .A(u2__abc_52155_new_n22531_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22532_));
AND2X2 AND2X2_11504 ( .A(u2__abc_52155_new_n22529_), .B(u2__abc_52155_new_n22532_), .Y(u2__abc_52155_new_n22533_));
AND2X2 AND2X2_11505 ( .A(u2__abc_52155_new_n22534_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__289_));
AND2X2 AND2X2_11506 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_289_), .Y(u2__abc_52155_new_n22536_));
AND2X2 AND2X2_11507 ( .A(u2__abc_52155_new_n22525_), .B(u2_o_288_), .Y(u2__abc_52155_new_n22538_));
AND2X2 AND2X2_11508 ( .A(u2__abc_52155_new_n22539_), .B(u2__abc_52155_new_n22537_), .Y(u2__abc_52155_new_n22540_));
AND2X2 AND2X2_11509 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6291_), .Y(u2__abc_52155_new_n22542_));
AND2X2 AND2X2_1151 ( .A(u2__abc_52155_new_n4358_), .B(u2__abc_52155_new_n4365_), .Y(u2__abc_52155_new_n4366_));
AND2X2 AND2X2_11510 ( .A(u2__abc_52155_new_n22543_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22544_));
AND2X2 AND2X2_11511 ( .A(u2__abc_52155_new_n22541_), .B(u2__abc_52155_new_n22544_), .Y(u2__abc_52155_new_n22545_));
AND2X2 AND2X2_11512 ( .A(u2__abc_52155_new_n22546_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__290_));
AND2X2 AND2X2_11513 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_290_), .Y(u2__abc_52155_new_n22548_));
AND2X2 AND2X2_11514 ( .A(u2__abc_52155_new_n22538_), .B(u2_o_289_), .Y(u2__abc_52155_new_n22549_));
AND2X2 AND2X2_11515 ( .A(u2__abc_52155_new_n22550_), .B(u2__abc_52155_new_n22551_), .Y(u2__abc_52155_new_n22552_));
AND2X2 AND2X2_11516 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6330_), .Y(u2__abc_52155_new_n22554_));
AND2X2 AND2X2_11517 ( .A(u2__abc_52155_new_n22555_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22556_));
AND2X2 AND2X2_11518 ( .A(u2__abc_52155_new_n22553_), .B(u2__abc_52155_new_n22556_), .Y(u2__abc_52155_new_n22557_));
AND2X2 AND2X2_11519 ( .A(u2__abc_52155_new_n22558_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__291_));
AND2X2 AND2X2_1152 ( .A(u2__abc_52155_new_n4367_), .B(u2_remHi_240_), .Y(u2__abc_52155_new_n4368_));
AND2X2 AND2X2_11520 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_291_), .Y(u2__abc_52155_new_n22560_));
AND2X2 AND2X2_11521 ( .A(u2__abc_52155_new_n22549_), .B(u2_o_290_), .Y(u2__abc_52155_new_n22562_));
AND2X2 AND2X2_11522 ( .A(u2__abc_52155_new_n22563_), .B(u2__abc_52155_new_n22561_), .Y(u2__abc_52155_new_n22564_));
AND2X2 AND2X2_11523 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6337_), .Y(u2__abc_52155_new_n22566_));
AND2X2 AND2X2_11524 ( .A(u2__abc_52155_new_n22567_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22568_));
AND2X2 AND2X2_11525 ( .A(u2__abc_52155_new_n22565_), .B(u2__abc_52155_new_n22568_), .Y(u2__abc_52155_new_n22569_));
AND2X2 AND2X2_11526 ( .A(u2__abc_52155_new_n22570_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__292_));
AND2X2 AND2X2_11527 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_292_), .Y(u2__abc_52155_new_n22572_));
AND2X2 AND2X2_11528 ( .A(u2__abc_52155_new_n22562_), .B(u2_o_291_), .Y(u2__abc_52155_new_n22574_));
AND2X2 AND2X2_11529 ( .A(u2__abc_52155_new_n22575_), .B(u2__abc_52155_new_n22573_), .Y(u2__abc_52155_new_n22576_));
AND2X2 AND2X2_1153 ( .A(u2__abc_52155_new_n4370_), .B(u2_o_240_), .Y(u2__abc_52155_new_n4371_));
AND2X2 AND2X2_11530 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6315_), .Y(u2__abc_52155_new_n22578_));
AND2X2 AND2X2_11531 ( .A(u2__abc_52155_new_n22579_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22580_));
AND2X2 AND2X2_11532 ( .A(u2__abc_52155_new_n22577_), .B(u2__abc_52155_new_n22580_), .Y(u2__abc_52155_new_n22581_));
AND2X2 AND2X2_11533 ( .A(u2__abc_52155_new_n22582_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__293_));
AND2X2 AND2X2_11534 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_293_), .Y(u2__abc_52155_new_n22584_));
AND2X2 AND2X2_11535 ( .A(u2__abc_52155_new_n22574_), .B(u2_o_292_), .Y(u2__abc_52155_new_n22586_));
AND2X2 AND2X2_11536 ( .A(u2__abc_52155_new_n22587_), .B(u2__abc_52155_new_n22585_), .Y(u2__abc_52155_new_n22588_));
AND2X2 AND2X2_11537 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6322_), .Y(u2__abc_52155_new_n22590_));
AND2X2 AND2X2_11538 ( .A(u2__abc_52155_new_n22591_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22592_));
AND2X2 AND2X2_11539 ( .A(u2__abc_52155_new_n22589_), .B(u2__abc_52155_new_n22592_), .Y(u2__abc_52155_new_n22593_));
AND2X2 AND2X2_1154 ( .A(u2__abc_52155_new_n4369_), .B(u2__abc_52155_new_n4372_), .Y(u2__abc_52155_new_n4373_));
AND2X2 AND2X2_11540 ( .A(u2__abc_52155_new_n22594_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__294_));
AND2X2 AND2X2_11541 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_294_), .Y(u2__abc_52155_new_n22596_));
AND2X2 AND2X2_11542 ( .A(u2__abc_52155_new_n22586_), .B(u2_o_293_), .Y(u2__abc_52155_new_n22597_));
AND2X2 AND2X2_11543 ( .A(u2__abc_52155_new_n22598_), .B(u2__abc_52155_new_n22599_), .Y(u2__abc_52155_new_n22600_));
AND2X2 AND2X2_11544 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6224_), .Y(u2__abc_52155_new_n22602_));
AND2X2 AND2X2_11545 ( .A(u2__abc_52155_new_n22603_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22604_));
AND2X2 AND2X2_11546 ( .A(u2__abc_52155_new_n22601_), .B(u2__abc_52155_new_n22604_), .Y(u2__abc_52155_new_n22605_));
AND2X2 AND2X2_11547 ( .A(u2__abc_52155_new_n22606_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__295_));
AND2X2 AND2X2_11548 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_295_), .Y(u2__abc_52155_new_n22608_));
AND2X2 AND2X2_11549 ( .A(u2__abc_52155_new_n22597_), .B(u2_o_294_), .Y(u2__abc_52155_new_n22610_));
AND2X2 AND2X2_1155 ( .A(u2__abc_52155_new_n4374_), .B(u2_remHi_241_), .Y(u2__abc_52155_new_n4375_));
AND2X2 AND2X2_11550 ( .A(u2__abc_52155_new_n22611_), .B(u2__abc_52155_new_n22609_), .Y(u2__abc_52155_new_n22612_));
AND2X2 AND2X2_11551 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6231_), .Y(u2__abc_52155_new_n22614_));
AND2X2 AND2X2_11552 ( .A(u2__abc_52155_new_n22615_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22616_));
AND2X2 AND2X2_11553 ( .A(u2__abc_52155_new_n22613_), .B(u2__abc_52155_new_n22616_), .Y(u2__abc_52155_new_n22617_));
AND2X2 AND2X2_11554 ( .A(u2__abc_52155_new_n22618_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__296_));
AND2X2 AND2X2_11555 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_296_), .Y(u2__abc_52155_new_n22620_));
AND2X2 AND2X2_11556 ( .A(u2__abc_52155_new_n22610_), .B(u2_o_295_), .Y(u2__abc_52155_new_n22622_));
AND2X2 AND2X2_11557 ( .A(u2__abc_52155_new_n22623_), .B(u2__abc_52155_new_n22621_), .Y(u2__abc_52155_new_n22624_));
AND2X2 AND2X2_11558 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6236_), .Y(u2__abc_52155_new_n22626_));
AND2X2 AND2X2_11559 ( .A(u2__abc_52155_new_n22627_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22628_));
AND2X2 AND2X2_1156 ( .A(u2__abc_52155_new_n4377_), .B(u2_o_241_), .Y(u2__abc_52155_new_n4378_));
AND2X2 AND2X2_11560 ( .A(u2__abc_52155_new_n22625_), .B(u2__abc_52155_new_n22628_), .Y(u2__abc_52155_new_n22629_));
AND2X2 AND2X2_11561 ( .A(u2__abc_52155_new_n22630_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__297_));
AND2X2 AND2X2_11562 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_297_), .Y(u2__abc_52155_new_n22632_));
AND2X2 AND2X2_11563 ( .A(u2__abc_52155_new_n22622_), .B(u2_o_296_), .Y(u2__abc_52155_new_n22634_));
AND2X2 AND2X2_11564 ( .A(u2__abc_52155_new_n22635_), .B(u2__abc_52155_new_n22633_), .Y(u2__abc_52155_new_n22636_));
AND2X2 AND2X2_11565 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6243_), .Y(u2__abc_52155_new_n22638_));
AND2X2 AND2X2_11566 ( .A(u2__abc_52155_new_n22639_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22640_));
AND2X2 AND2X2_11567 ( .A(u2__abc_52155_new_n22637_), .B(u2__abc_52155_new_n22640_), .Y(u2__abc_52155_new_n22641_));
AND2X2 AND2X2_11568 ( .A(u2__abc_52155_new_n22642_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__298_));
AND2X2 AND2X2_11569 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_298_), .Y(u2__abc_52155_new_n22644_));
AND2X2 AND2X2_1157 ( .A(u2__abc_52155_new_n4376_), .B(u2__abc_52155_new_n4379_), .Y(u2__abc_52155_new_n4380_));
AND2X2 AND2X2_11570 ( .A(u2__abc_52155_new_n22634_), .B(u2_o_297_), .Y(u2__abc_52155_new_n22645_));
AND2X2 AND2X2_11571 ( .A(u2__abc_52155_new_n22646_), .B(u2__abc_52155_new_n22647_), .Y(u2__abc_52155_new_n22648_));
AND2X2 AND2X2_11572 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6267_), .Y(u2__abc_52155_new_n22650_));
AND2X2 AND2X2_11573 ( .A(u2__abc_52155_new_n22651_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22652_));
AND2X2 AND2X2_11574 ( .A(u2__abc_52155_new_n22649_), .B(u2__abc_52155_new_n22652_), .Y(u2__abc_52155_new_n22653_));
AND2X2 AND2X2_11575 ( .A(u2__abc_52155_new_n22654_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__299_));
AND2X2 AND2X2_11576 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_299_), .Y(u2__abc_52155_new_n22656_));
AND2X2 AND2X2_11577 ( .A(u2__abc_52155_new_n22645_), .B(u2_o_298_), .Y(u2__abc_52155_new_n22658_));
AND2X2 AND2X2_11578 ( .A(u2__abc_52155_new_n22659_), .B(u2__abc_52155_new_n22657_), .Y(u2__abc_52155_new_n22660_));
AND2X2 AND2X2_11579 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6274_), .Y(u2__abc_52155_new_n22662_));
AND2X2 AND2X2_1158 ( .A(u2__abc_52155_new_n4373_), .B(u2__abc_52155_new_n4380_), .Y(u2__abc_52155_new_n4381_));
AND2X2 AND2X2_11580 ( .A(u2__abc_52155_new_n22663_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22664_));
AND2X2 AND2X2_11581 ( .A(u2__abc_52155_new_n22661_), .B(u2__abc_52155_new_n22664_), .Y(u2__abc_52155_new_n22665_));
AND2X2 AND2X2_11582 ( .A(u2__abc_52155_new_n22666_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__300_));
AND2X2 AND2X2_11583 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_300_), .Y(u2__abc_52155_new_n22668_));
AND2X2 AND2X2_11584 ( .A(u2__abc_52155_new_n22658_), .B(u2_o_299_), .Y(u2__abc_52155_new_n22670_));
AND2X2 AND2X2_11585 ( .A(u2__abc_52155_new_n22671_), .B(u2__abc_52155_new_n22669_), .Y(u2__abc_52155_new_n22672_));
AND2X2 AND2X2_11586 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6252_), .Y(u2__abc_52155_new_n22674_));
AND2X2 AND2X2_11587 ( .A(u2__abc_52155_new_n22675_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22676_));
AND2X2 AND2X2_11588 ( .A(u2__abc_52155_new_n22673_), .B(u2__abc_52155_new_n22676_), .Y(u2__abc_52155_new_n22677_));
AND2X2 AND2X2_11589 ( .A(u2__abc_52155_new_n22678_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__301_));
AND2X2 AND2X2_1159 ( .A(u2__abc_52155_new_n4366_), .B(u2__abc_52155_new_n4381_), .Y(u2__abc_52155_new_n4382_));
AND2X2 AND2X2_11590 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_301_), .Y(u2__abc_52155_new_n22680_));
AND2X2 AND2X2_11591 ( .A(u2__abc_52155_new_n22670_), .B(u2_o_300_), .Y(u2__abc_52155_new_n22682_));
AND2X2 AND2X2_11592 ( .A(u2__abc_52155_new_n22683_), .B(u2__abc_52155_new_n22681_), .Y(u2__abc_52155_new_n22684_));
AND2X2 AND2X2_11593 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6259_), .Y(u2__abc_52155_new_n22686_));
AND2X2 AND2X2_11594 ( .A(u2__abc_52155_new_n22687_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22688_));
AND2X2 AND2X2_11595 ( .A(u2__abc_52155_new_n22685_), .B(u2__abc_52155_new_n22688_), .Y(u2__abc_52155_new_n22689_));
AND2X2 AND2X2_11596 ( .A(u2__abc_52155_new_n22690_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__302_));
AND2X2 AND2X2_11597 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_302_), .Y(u2__abc_52155_new_n22692_));
AND2X2 AND2X2_11598 ( .A(u2__abc_52155_new_n22682_), .B(u2_o_301_), .Y(u2__abc_52155_new_n22693_));
AND2X2 AND2X2_11599 ( .A(u2__abc_52155_new_n22694_), .B(u2__abc_52155_new_n22695_), .Y(u2__abc_52155_new_n22696_));
AND2X2 AND2X2_116 ( .A(_abc_73687_new_n948_), .B(_abc_73687_new_n947_), .Y(\o[151] ));
AND2X2 AND2X2_1160 ( .A(u2__abc_52155_new_n4383_), .B(u2_remHi_244_), .Y(u2__abc_52155_new_n4384_));
AND2X2 AND2X2_11600 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6160_), .Y(u2__abc_52155_new_n22698_));
AND2X2 AND2X2_11601 ( .A(u2__abc_52155_new_n22699_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22700_));
AND2X2 AND2X2_11602 ( .A(u2__abc_52155_new_n22697_), .B(u2__abc_52155_new_n22700_), .Y(u2__abc_52155_new_n22701_));
AND2X2 AND2X2_11603 ( .A(u2__abc_52155_new_n22702_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__303_));
AND2X2 AND2X2_11604 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_303_), .Y(u2__abc_52155_new_n22704_));
AND2X2 AND2X2_11605 ( .A(u2__abc_52155_new_n22693_), .B(u2_o_302_), .Y(u2__abc_52155_new_n22706_));
AND2X2 AND2X2_11606 ( .A(u2__abc_52155_new_n22707_), .B(u2__abc_52155_new_n22705_), .Y(u2__abc_52155_new_n22708_));
AND2X2 AND2X2_11607 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6167_), .Y(u2__abc_52155_new_n22710_));
AND2X2 AND2X2_11608 ( .A(u2__abc_52155_new_n22711_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22712_));
AND2X2 AND2X2_11609 ( .A(u2__abc_52155_new_n22709_), .B(u2__abc_52155_new_n22712_), .Y(u2__abc_52155_new_n22713_));
AND2X2 AND2X2_1161 ( .A(u2__abc_52155_new_n4386_), .B(u2_o_244_), .Y(u2__abc_52155_new_n4387_));
AND2X2 AND2X2_11610 ( .A(u2__abc_52155_new_n22714_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__304_));
AND2X2 AND2X2_11611 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_304_), .Y(u2__abc_52155_new_n22716_));
AND2X2 AND2X2_11612 ( .A(u2__abc_52155_new_n22706_), .B(u2_o_303_), .Y(u2__abc_52155_new_n22717_));
AND2X2 AND2X2_11613 ( .A(u2__abc_52155_new_n22718_), .B(u2__abc_52155_new_n22719_), .Y(u2__abc_52155_new_n22720_));
AND2X2 AND2X2_11614 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6172_), .Y(u2__abc_52155_new_n22722_));
AND2X2 AND2X2_11615 ( .A(u2__abc_52155_new_n22723_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22724_));
AND2X2 AND2X2_11616 ( .A(u2__abc_52155_new_n22721_), .B(u2__abc_52155_new_n22724_), .Y(u2__abc_52155_new_n22725_));
AND2X2 AND2X2_11617 ( .A(u2__abc_52155_new_n22726_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__305_));
AND2X2 AND2X2_11618 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_305_), .Y(u2__abc_52155_new_n22728_));
AND2X2 AND2X2_11619 ( .A(u2__abc_52155_new_n22717_), .B(u2_o_304_), .Y(u2__abc_52155_new_n22730_));
AND2X2 AND2X2_1162 ( .A(u2__abc_52155_new_n4385_), .B(u2__abc_52155_new_n4388_), .Y(u2__abc_52155_new_n4389_));
AND2X2 AND2X2_11620 ( .A(u2__abc_52155_new_n22731_), .B(u2__abc_52155_new_n22729_), .Y(u2__abc_52155_new_n22732_));
AND2X2 AND2X2_11621 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6179_), .Y(u2__abc_52155_new_n22734_));
AND2X2 AND2X2_11622 ( .A(u2__abc_52155_new_n22735_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22736_));
AND2X2 AND2X2_11623 ( .A(u2__abc_52155_new_n22733_), .B(u2__abc_52155_new_n22736_), .Y(u2__abc_52155_new_n22737_));
AND2X2 AND2X2_11624 ( .A(u2__abc_52155_new_n22738_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__306_));
AND2X2 AND2X2_11625 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_306_), .Y(u2__abc_52155_new_n22740_));
AND2X2 AND2X2_11626 ( .A(u2__abc_52155_new_n22730_), .B(u2_o_305_), .Y(u2__abc_52155_new_n22741_));
AND2X2 AND2X2_11627 ( .A(u2__abc_52155_new_n22742_), .B(u2__abc_52155_new_n22743_), .Y(u2__abc_52155_new_n22744_));
AND2X2 AND2X2_11628 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6210_), .Y(u2__abc_52155_new_n22746_));
AND2X2 AND2X2_11629 ( .A(u2__abc_52155_new_n22747_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22748_));
AND2X2 AND2X2_1163 ( .A(u2__abc_52155_new_n4390_), .B(u2_remHi_245_), .Y(u2__abc_52155_new_n4391_));
AND2X2 AND2X2_11630 ( .A(u2__abc_52155_new_n22745_), .B(u2__abc_52155_new_n22748_), .Y(u2__abc_52155_new_n22749_));
AND2X2 AND2X2_11631 ( .A(u2__abc_52155_new_n22750_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__307_));
AND2X2 AND2X2_11632 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_307_), .Y(u2__abc_52155_new_n22752_));
AND2X2 AND2X2_11633 ( .A(u2__abc_52155_new_n22741_), .B(u2_o_306_), .Y(u2__abc_52155_new_n22754_));
AND2X2 AND2X2_11634 ( .A(u2__abc_52155_new_n22755_), .B(u2__abc_52155_new_n22753_), .Y(u2__abc_52155_new_n22756_));
AND2X2 AND2X2_11635 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6203_), .Y(u2__abc_52155_new_n22758_));
AND2X2 AND2X2_11636 ( .A(u2__abc_52155_new_n22759_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22760_));
AND2X2 AND2X2_11637 ( .A(u2__abc_52155_new_n22757_), .B(u2__abc_52155_new_n22760_), .Y(u2__abc_52155_new_n22761_));
AND2X2 AND2X2_11638 ( .A(u2__abc_52155_new_n22762_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__308_));
AND2X2 AND2X2_11639 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_308_), .Y(u2__abc_52155_new_n22764_));
AND2X2 AND2X2_1164 ( .A(u2__abc_52155_new_n4393_), .B(u2_o_245_), .Y(u2__abc_52155_new_n4394_));
AND2X2 AND2X2_11640 ( .A(u2__abc_52155_new_n22754_), .B(u2_o_307_), .Y(u2__abc_52155_new_n22766_));
AND2X2 AND2X2_11641 ( .A(u2__abc_52155_new_n22767_), .B(u2__abc_52155_new_n22765_), .Y(u2__abc_52155_new_n22768_));
AND2X2 AND2X2_11642 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6188_), .Y(u2__abc_52155_new_n22770_));
AND2X2 AND2X2_11643 ( .A(u2__abc_52155_new_n22771_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22772_));
AND2X2 AND2X2_11644 ( .A(u2__abc_52155_new_n22769_), .B(u2__abc_52155_new_n22772_), .Y(u2__abc_52155_new_n22773_));
AND2X2 AND2X2_11645 ( .A(u2__abc_52155_new_n22774_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__309_));
AND2X2 AND2X2_11646 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_309_), .Y(u2__abc_52155_new_n22776_));
AND2X2 AND2X2_11647 ( .A(u2__abc_52155_new_n22766_), .B(u2_o_308_), .Y(u2__abc_52155_new_n22778_));
AND2X2 AND2X2_11648 ( .A(u2__abc_52155_new_n22779_), .B(u2__abc_52155_new_n22777_), .Y(u2__abc_52155_new_n22780_));
AND2X2 AND2X2_11649 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6195_), .Y(u2__abc_52155_new_n22782_));
AND2X2 AND2X2_1165 ( .A(u2__abc_52155_new_n4392_), .B(u2__abc_52155_new_n4395_), .Y(u2__abc_52155_new_n4396_));
AND2X2 AND2X2_11650 ( .A(u2__abc_52155_new_n22783_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22784_));
AND2X2 AND2X2_11651 ( .A(u2__abc_52155_new_n22781_), .B(u2__abc_52155_new_n22784_), .Y(u2__abc_52155_new_n22785_));
AND2X2 AND2X2_11652 ( .A(u2__abc_52155_new_n22786_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__310_));
AND2X2 AND2X2_11653 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_310_), .Y(u2__abc_52155_new_n22788_));
AND2X2 AND2X2_11654 ( .A(u2__abc_52155_new_n22778_), .B(u2_o_309_), .Y(u2__abc_52155_new_n22789_));
AND2X2 AND2X2_11655 ( .A(u2__abc_52155_new_n22790_), .B(u2__abc_52155_new_n22791_), .Y(u2__abc_52155_new_n22792_));
AND2X2 AND2X2_11656 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6109_), .Y(u2__abc_52155_new_n22794_));
AND2X2 AND2X2_11657 ( .A(u2__abc_52155_new_n22795_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22796_));
AND2X2 AND2X2_11658 ( .A(u2__abc_52155_new_n22793_), .B(u2__abc_52155_new_n22796_), .Y(u2__abc_52155_new_n22797_));
AND2X2 AND2X2_11659 ( .A(u2__abc_52155_new_n22798_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__311_));
AND2X2 AND2X2_1166 ( .A(u2__abc_52155_new_n4389_), .B(u2__abc_52155_new_n4396_), .Y(u2__abc_52155_new_n4397_));
AND2X2 AND2X2_11660 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_311_), .Y(u2__abc_52155_new_n22800_));
AND2X2 AND2X2_11661 ( .A(u2__abc_52155_new_n22789_), .B(u2_o_310_), .Y(u2__abc_52155_new_n22802_));
AND2X2 AND2X2_11662 ( .A(u2__abc_52155_new_n22803_), .B(u2__abc_52155_new_n22801_), .Y(u2__abc_52155_new_n22804_));
AND2X2 AND2X2_11663 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6116_), .Y(u2__abc_52155_new_n22806_));
AND2X2 AND2X2_11664 ( .A(u2__abc_52155_new_n22807_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22808_));
AND2X2 AND2X2_11665 ( .A(u2__abc_52155_new_n22805_), .B(u2__abc_52155_new_n22808_), .Y(u2__abc_52155_new_n22809_));
AND2X2 AND2X2_11666 ( .A(u2__abc_52155_new_n22810_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__312_));
AND2X2 AND2X2_11667 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_312_), .Y(u2__abc_52155_new_n22812_));
AND2X2 AND2X2_11668 ( .A(u2__abc_52155_new_n22802_), .B(u2_o_311_), .Y(u2__abc_52155_new_n22813_));
AND2X2 AND2X2_11669 ( .A(u2__abc_52155_new_n22814_), .B(u2__abc_52155_new_n22815_), .Y(u2__abc_52155_new_n22816_));
AND2X2 AND2X2_1167 ( .A(u2__abc_52155_new_n4398_), .B(u2_remHi_243_), .Y(u2__abc_52155_new_n4399_));
AND2X2 AND2X2_11670 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6094_), .Y(u2__abc_52155_new_n22818_));
AND2X2 AND2X2_11671 ( .A(u2__abc_52155_new_n22819_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22820_));
AND2X2 AND2X2_11672 ( .A(u2__abc_52155_new_n22817_), .B(u2__abc_52155_new_n22820_), .Y(u2__abc_52155_new_n22821_));
AND2X2 AND2X2_11673 ( .A(u2__abc_52155_new_n22822_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__313_));
AND2X2 AND2X2_11674 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_313_), .Y(u2__abc_52155_new_n22824_));
AND2X2 AND2X2_11675 ( .A(u2__abc_52155_new_n22813_), .B(u2_o_312_), .Y(u2__abc_52155_new_n22826_));
AND2X2 AND2X2_11676 ( .A(u2__abc_52155_new_n22827_), .B(u2__abc_52155_new_n22825_), .Y(u2__abc_52155_new_n22828_));
AND2X2 AND2X2_11677 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6101_), .Y(u2__abc_52155_new_n22830_));
AND2X2 AND2X2_11678 ( .A(u2__abc_52155_new_n22831_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22832_));
AND2X2 AND2X2_11679 ( .A(u2__abc_52155_new_n22829_), .B(u2__abc_52155_new_n22832_), .Y(u2__abc_52155_new_n22833_));
AND2X2 AND2X2_1168 ( .A(u2__abc_52155_new_n4401_), .B(u2_o_243_), .Y(u2__abc_52155_new_n4402_));
AND2X2 AND2X2_11680 ( .A(u2__abc_52155_new_n22834_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__314_));
AND2X2 AND2X2_11681 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_314_), .Y(u2__abc_52155_new_n22836_));
AND2X2 AND2X2_11682 ( .A(u2__abc_52155_new_n22826_), .B(u2_o_313_), .Y(u2__abc_52155_new_n22837_));
AND2X2 AND2X2_11683 ( .A(u2__abc_52155_new_n22838_), .B(u2__abc_52155_new_n22839_), .Y(u2__abc_52155_new_n22840_));
AND2X2 AND2X2_11684 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6140_), .Y(u2__abc_52155_new_n22842_));
AND2X2 AND2X2_11685 ( .A(u2__abc_52155_new_n22843_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22844_));
AND2X2 AND2X2_11686 ( .A(u2__abc_52155_new_n22841_), .B(u2__abc_52155_new_n22844_), .Y(u2__abc_52155_new_n22845_));
AND2X2 AND2X2_11687 ( .A(u2__abc_52155_new_n22846_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__315_));
AND2X2 AND2X2_11688 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_315_), .Y(u2__abc_52155_new_n22848_));
AND2X2 AND2X2_11689 ( .A(u2__abc_52155_new_n22837_), .B(u2_o_314_), .Y(u2__abc_52155_new_n22850_));
AND2X2 AND2X2_1169 ( .A(u2__abc_52155_new_n4400_), .B(u2__abc_52155_new_n4403_), .Y(u2__abc_52155_new_n4404_));
AND2X2 AND2X2_11690 ( .A(u2__abc_52155_new_n22851_), .B(u2__abc_52155_new_n22849_), .Y(u2__abc_52155_new_n22852_));
AND2X2 AND2X2_11691 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6147_), .Y(u2__abc_52155_new_n22854_));
AND2X2 AND2X2_11692 ( .A(u2__abc_52155_new_n22855_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22856_));
AND2X2 AND2X2_11693 ( .A(u2__abc_52155_new_n22853_), .B(u2__abc_52155_new_n22856_), .Y(u2__abc_52155_new_n22857_));
AND2X2 AND2X2_11694 ( .A(u2__abc_52155_new_n22858_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__316_));
AND2X2 AND2X2_11695 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_316_), .Y(u2__abc_52155_new_n22860_));
AND2X2 AND2X2_11696 ( .A(u2__abc_52155_new_n22850_), .B(u2_o_315_), .Y(u2__abc_52155_new_n22861_));
AND2X2 AND2X2_11697 ( .A(u2__abc_52155_new_n22862_), .B(u2__abc_52155_new_n22863_), .Y(u2__abc_52155_new_n22864_));
AND2X2 AND2X2_11698 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6125_), .Y(u2__abc_52155_new_n22866_));
AND2X2 AND2X2_11699 ( .A(u2__abc_52155_new_n22867_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22868_));
AND2X2 AND2X2_117 ( .A(_abc_73687_new_n951_), .B(_abc_73687_new_n950_), .Y(\o[152] ));
AND2X2 AND2X2_1170 ( .A(u2__abc_52155_new_n4405_), .B(u2_remHi_242_), .Y(u2__abc_52155_new_n4406_));
AND2X2 AND2X2_11700 ( .A(u2__abc_52155_new_n22865_), .B(u2__abc_52155_new_n22868_), .Y(u2__abc_52155_new_n22869_));
AND2X2 AND2X2_11701 ( .A(u2__abc_52155_new_n22870_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__317_));
AND2X2 AND2X2_11702 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_317_), .Y(u2__abc_52155_new_n22872_));
AND2X2 AND2X2_11703 ( .A(u2__abc_52155_new_n22861_), .B(u2_o_316_), .Y(u2__abc_52155_new_n22874_));
AND2X2 AND2X2_11704 ( .A(u2__abc_52155_new_n22875_), .B(u2__abc_52155_new_n22873_), .Y(u2__abc_52155_new_n22876_));
AND2X2 AND2X2_11705 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6132_), .Y(u2__abc_52155_new_n22878_));
AND2X2 AND2X2_11706 ( .A(u2__abc_52155_new_n22879_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22880_));
AND2X2 AND2X2_11707 ( .A(u2__abc_52155_new_n22877_), .B(u2__abc_52155_new_n22880_), .Y(u2__abc_52155_new_n22881_));
AND2X2 AND2X2_11708 ( .A(u2__abc_52155_new_n22882_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__318_));
AND2X2 AND2X2_11709 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_318_), .Y(u2__abc_52155_new_n22884_));
AND2X2 AND2X2_1171 ( .A(u2__abc_52155_new_n4408_), .B(u2_o_242_), .Y(u2__abc_52155_new_n4409_));
AND2X2 AND2X2_11710 ( .A(u2__abc_52155_new_n22874_), .B(u2_o_317_), .Y(u2__abc_52155_new_n22885_));
AND2X2 AND2X2_11711 ( .A(u2__abc_52155_new_n22886_), .B(u2__abc_52155_new_n22887_), .Y(u2__abc_52155_new_n22888_));
AND2X2 AND2X2_11712 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6062_), .Y(u2__abc_52155_new_n22890_));
AND2X2 AND2X2_11713 ( .A(u2__abc_52155_new_n22891_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22892_));
AND2X2 AND2X2_11714 ( .A(u2__abc_52155_new_n22889_), .B(u2__abc_52155_new_n22892_), .Y(u2__abc_52155_new_n22893_));
AND2X2 AND2X2_11715 ( .A(u2__abc_52155_new_n22894_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__319_));
AND2X2 AND2X2_11716 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_319_), .Y(u2__abc_52155_new_n22896_));
AND2X2 AND2X2_11717 ( .A(u2__abc_52155_new_n22885_), .B(u2_o_318_), .Y(u2__abc_52155_new_n22898_));
AND2X2 AND2X2_11718 ( .A(u2__abc_52155_new_n22899_), .B(u2__abc_52155_new_n22897_), .Y(u2__abc_52155_new_n22900_));
AND2X2 AND2X2_11719 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6069_), .Y(u2__abc_52155_new_n22902_));
AND2X2 AND2X2_1172 ( .A(u2__abc_52155_new_n4407_), .B(u2__abc_52155_new_n4410_), .Y(u2__abc_52155_new_n4411_));
AND2X2 AND2X2_11720 ( .A(u2__abc_52155_new_n22903_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22904_));
AND2X2 AND2X2_11721 ( .A(u2__abc_52155_new_n22901_), .B(u2__abc_52155_new_n22904_), .Y(u2__abc_52155_new_n22905_));
AND2X2 AND2X2_11722 ( .A(u2__abc_52155_new_n22906_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__320_));
AND2X2 AND2X2_11723 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_320_), .Y(u2__abc_52155_new_n22908_));
AND2X2 AND2X2_11724 ( .A(u2__abc_52155_new_n22898_), .B(u2_o_319_), .Y(u2__abc_52155_new_n22909_));
AND2X2 AND2X2_11725 ( .A(u2__abc_52155_new_n22910_), .B(u2__abc_52155_new_n22911_), .Y(u2__abc_52155_new_n22912_));
AND2X2 AND2X2_11726 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6074_), .Y(u2__abc_52155_new_n22914_));
AND2X2 AND2X2_11727 ( .A(u2__abc_52155_new_n22915_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22916_));
AND2X2 AND2X2_11728 ( .A(u2__abc_52155_new_n22913_), .B(u2__abc_52155_new_n22916_), .Y(u2__abc_52155_new_n22917_));
AND2X2 AND2X2_11729 ( .A(u2__abc_52155_new_n22918_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__321_));
AND2X2 AND2X2_1173 ( .A(u2__abc_52155_new_n4404_), .B(u2__abc_52155_new_n4411_), .Y(u2__abc_52155_new_n4412_));
AND2X2 AND2X2_11730 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_321_), .Y(u2__abc_52155_new_n22920_));
AND2X2 AND2X2_11731 ( .A(u2__abc_52155_new_n22909_), .B(u2_o_320_), .Y(u2__abc_52155_new_n22922_));
AND2X2 AND2X2_11732 ( .A(u2__abc_52155_new_n22923_), .B(u2__abc_52155_new_n22921_), .Y(u2__abc_52155_new_n22924_));
AND2X2 AND2X2_11733 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6081_), .Y(u2__abc_52155_new_n22926_));
AND2X2 AND2X2_11734 ( .A(u2__abc_52155_new_n22927_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22928_));
AND2X2 AND2X2_11735 ( .A(u2__abc_52155_new_n22925_), .B(u2__abc_52155_new_n22928_), .Y(u2__abc_52155_new_n22929_));
AND2X2 AND2X2_11736 ( .A(u2__abc_52155_new_n22930_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__322_));
AND2X2 AND2X2_11737 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_322_), .Y(u2__abc_52155_new_n22932_));
AND2X2 AND2X2_11738 ( .A(u2__abc_52155_new_n22922_), .B(u2_o_321_), .Y(u2__abc_52155_new_n22933_));
AND2X2 AND2X2_11739 ( .A(u2__abc_52155_new_n22934_), .B(u2__abc_52155_new_n22935_), .Y(u2__abc_52155_new_n22936_));
AND2X2 AND2X2_1174 ( .A(u2__abc_52155_new_n4397_), .B(u2__abc_52155_new_n4412_), .Y(u2__abc_52155_new_n4413_));
AND2X2 AND2X2_11740 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6043_), .Y(u2__abc_52155_new_n22938_));
AND2X2 AND2X2_11741 ( .A(u2__abc_52155_new_n22939_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22940_));
AND2X2 AND2X2_11742 ( .A(u2__abc_52155_new_n22937_), .B(u2__abc_52155_new_n22940_), .Y(u2__abc_52155_new_n22941_));
AND2X2 AND2X2_11743 ( .A(u2__abc_52155_new_n22942_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__323_));
AND2X2 AND2X2_11744 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_323_), .Y(u2__abc_52155_new_n22944_));
AND2X2 AND2X2_11745 ( .A(u2__abc_52155_new_n22933_), .B(u2_o_322_), .Y(u2__abc_52155_new_n22946_));
AND2X2 AND2X2_11746 ( .A(u2__abc_52155_new_n22947_), .B(u2__abc_52155_new_n22945_), .Y(u2__abc_52155_new_n22948_));
AND2X2 AND2X2_11747 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6050_), .Y(u2__abc_52155_new_n22950_));
AND2X2 AND2X2_11748 ( .A(u2__abc_52155_new_n22951_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22952_));
AND2X2 AND2X2_11749 ( .A(u2__abc_52155_new_n22949_), .B(u2__abc_52155_new_n22952_), .Y(u2__abc_52155_new_n22953_));
AND2X2 AND2X2_1175 ( .A(u2__abc_52155_new_n4382_), .B(u2__abc_52155_new_n4413_), .Y(u2__abc_52155_new_n4414_));
AND2X2 AND2X2_11750 ( .A(u2__abc_52155_new_n22954_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__324_));
AND2X2 AND2X2_11751 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_324_), .Y(u2__abc_52155_new_n22956_));
AND2X2 AND2X2_11752 ( .A(u2__abc_52155_new_n22946_), .B(u2_o_323_), .Y(u2__abc_52155_new_n22958_));
AND2X2 AND2X2_11753 ( .A(u2__abc_52155_new_n22959_), .B(u2__abc_52155_new_n22957_), .Y(u2__abc_52155_new_n22960_));
AND2X2 AND2X2_11754 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6031_), .Y(u2__abc_52155_new_n22962_));
AND2X2 AND2X2_11755 ( .A(u2__abc_52155_new_n22963_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22964_));
AND2X2 AND2X2_11756 ( .A(u2__abc_52155_new_n22961_), .B(u2__abc_52155_new_n22964_), .Y(u2__abc_52155_new_n22965_));
AND2X2 AND2X2_11757 ( .A(u2__abc_52155_new_n22966_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__325_));
AND2X2 AND2X2_11758 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_325_), .Y(u2__abc_52155_new_n22968_));
AND2X2 AND2X2_11759 ( .A(u2__abc_52155_new_n22958_), .B(u2_o_324_), .Y(u2__abc_52155_new_n22970_));
AND2X2 AND2X2_1176 ( .A(u2__abc_52155_new_n4351_), .B(u2__abc_52155_new_n4414_), .Y(u2__abc_52155_new_n4415_));
AND2X2 AND2X2_11760 ( .A(u2__abc_52155_new_n22971_), .B(u2__abc_52155_new_n22969_), .Y(u2__abc_52155_new_n22972_));
AND2X2 AND2X2_11761 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6038_), .Y(u2__abc_52155_new_n22974_));
AND2X2 AND2X2_11762 ( .A(u2__abc_52155_new_n22975_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22976_));
AND2X2 AND2X2_11763 ( .A(u2__abc_52155_new_n22973_), .B(u2__abc_52155_new_n22976_), .Y(u2__abc_52155_new_n22977_));
AND2X2 AND2X2_11764 ( .A(u2__abc_52155_new_n22978_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__326_));
AND2X2 AND2X2_11765 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_326_), .Y(u2__abc_52155_new_n22980_));
AND2X2 AND2X2_11766 ( .A(u2__abc_52155_new_n22970_), .B(u2_o_325_), .Y(u2__abc_52155_new_n22981_));
AND2X2 AND2X2_11767 ( .A(u2__abc_52155_new_n22982_), .B(u2__abc_52155_new_n22983_), .Y(u2__abc_52155_new_n22984_));
AND2X2 AND2X2_11768 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5968_), .Y(u2__abc_52155_new_n22986_));
AND2X2 AND2X2_11769 ( .A(u2__abc_52155_new_n22987_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n22988_));
AND2X2 AND2X2_1177 ( .A(u2__abc_52155_new_n4416_), .B(u2_remHi_236_), .Y(u2__abc_52155_new_n4417_));
AND2X2 AND2X2_11770 ( .A(u2__abc_52155_new_n22985_), .B(u2__abc_52155_new_n22988_), .Y(u2__abc_52155_new_n22989_));
AND2X2 AND2X2_11771 ( .A(u2__abc_52155_new_n22990_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__327_));
AND2X2 AND2X2_11772 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_327_), .Y(u2__abc_52155_new_n22992_));
AND2X2 AND2X2_11773 ( .A(u2__abc_52155_new_n22981_), .B(u2_o_326_), .Y(u2__abc_52155_new_n22994_));
AND2X2 AND2X2_11774 ( .A(u2__abc_52155_new_n22995_), .B(u2__abc_52155_new_n22993_), .Y(u2__abc_52155_new_n22996_));
AND2X2 AND2X2_11775 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5975_), .Y(u2__abc_52155_new_n22998_));
AND2X2 AND2X2_11776 ( .A(u2__abc_52155_new_n22999_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23000_));
AND2X2 AND2X2_11777 ( .A(u2__abc_52155_new_n22997_), .B(u2__abc_52155_new_n23000_), .Y(u2__abc_52155_new_n23001_));
AND2X2 AND2X2_11778 ( .A(u2__abc_52155_new_n23002_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__328_));
AND2X2 AND2X2_11779 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_328_), .Y(u2__abc_52155_new_n23004_));
AND2X2 AND2X2_1178 ( .A(u2__abc_52155_new_n4419_), .B(u2_o_236_), .Y(u2__abc_52155_new_n4420_));
AND2X2 AND2X2_11780 ( .A(u2__abc_52155_new_n22994_), .B(u2_o_327_), .Y(u2__abc_52155_new_n23006_));
AND2X2 AND2X2_11781 ( .A(u2__abc_52155_new_n23007_), .B(u2__abc_52155_new_n23005_), .Y(u2__abc_52155_new_n23008_));
AND2X2 AND2X2_11782 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5980_), .Y(u2__abc_52155_new_n23010_));
AND2X2 AND2X2_11783 ( .A(u2__abc_52155_new_n23011_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23012_));
AND2X2 AND2X2_11784 ( .A(u2__abc_52155_new_n23009_), .B(u2__abc_52155_new_n23012_), .Y(u2__abc_52155_new_n23013_));
AND2X2 AND2X2_11785 ( .A(u2__abc_52155_new_n23014_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__329_));
AND2X2 AND2X2_11786 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_329_), .Y(u2__abc_52155_new_n23016_));
AND2X2 AND2X2_11787 ( .A(u2__abc_52155_new_n23006_), .B(u2_o_328_), .Y(u2__abc_52155_new_n23018_));
AND2X2 AND2X2_11788 ( .A(u2__abc_52155_new_n23019_), .B(u2__abc_52155_new_n23017_), .Y(u2__abc_52155_new_n23020_));
AND2X2 AND2X2_11789 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5987_), .Y(u2__abc_52155_new_n23022_));
AND2X2 AND2X2_1179 ( .A(u2__abc_52155_new_n4418_), .B(u2__abc_52155_new_n4421_), .Y(u2__abc_52155_new_n4422_));
AND2X2 AND2X2_11790 ( .A(u2__abc_52155_new_n23023_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23024_));
AND2X2 AND2X2_11791 ( .A(u2__abc_52155_new_n23021_), .B(u2__abc_52155_new_n23024_), .Y(u2__abc_52155_new_n23025_));
AND2X2 AND2X2_11792 ( .A(u2__abc_52155_new_n23026_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__330_));
AND2X2 AND2X2_11793 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_330_), .Y(u2__abc_52155_new_n23028_));
AND2X2 AND2X2_11794 ( .A(u2__abc_52155_new_n23018_), .B(u2_o_329_), .Y(u2__abc_52155_new_n23029_));
AND2X2 AND2X2_11795 ( .A(u2__abc_52155_new_n23030_), .B(u2__abc_52155_new_n23031_), .Y(u2__abc_52155_new_n23032_));
AND2X2 AND2X2_11796 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6011_), .Y(u2__abc_52155_new_n23034_));
AND2X2 AND2X2_11797 ( .A(u2__abc_52155_new_n23035_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23036_));
AND2X2 AND2X2_11798 ( .A(u2__abc_52155_new_n23033_), .B(u2__abc_52155_new_n23036_), .Y(u2__abc_52155_new_n23037_));
AND2X2 AND2X2_11799 ( .A(u2__abc_52155_new_n23038_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__331_));
AND2X2 AND2X2_118 ( .A(_abc_73687_new_n954_), .B(_abc_73687_new_n953_), .Y(\o[153] ));
AND2X2 AND2X2_1180 ( .A(u2__abc_52155_new_n4423_), .B(u2_remHi_237_), .Y(u2__abc_52155_new_n4424_));
AND2X2 AND2X2_11800 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_331_), .Y(u2__abc_52155_new_n23040_));
AND2X2 AND2X2_11801 ( .A(u2__abc_52155_new_n23029_), .B(u2_o_330_), .Y(u2__abc_52155_new_n23042_));
AND2X2 AND2X2_11802 ( .A(u2__abc_52155_new_n23043_), .B(u2__abc_52155_new_n23041_), .Y(u2__abc_52155_new_n23044_));
AND2X2 AND2X2_11803 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6018_), .Y(u2__abc_52155_new_n23046_));
AND2X2 AND2X2_11804 ( .A(u2__abc_52155_new_n23047_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23048_));
AND2X2 AND2X2_11805 ( .A(u2__abc_52155_new_n23045_), .B(u2__abc_52155_new_n23048_), .Y(u2__abc_52155_new_n23049_));
AND2X2 AND2X2_11806 ( .A(u2__abc_52155_new_n23050_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__332_));
AND2X2 AND2X2_11807 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_332_), .Y(u2__abc_52155_new_n23052_));
AND2X2 AND2X2_11808 ( .A(u2__abc_52155_new_n23042_), .B(u2_o_331_), .Y(u2__abc_52155_new_n23054_));
AND2X2 AND2X2_11809 ( .A(u2__abc_52155_new_n23055_), .B(u2__abc_52155_new_n23053_), .Y(u2__abc_52155_new_n23056_));
AND2X2 AND2X2_1181 ( .A(u2__abc_52155_new_n4426_), .B(u2_o_237_), .Y(u2__abc_52155_new_n4427_));
AND2X2 AND2X2_11810 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5996_), .Y(u2__abc_52155_new_n23058_));
AND2X2 AND2X2_11811 ( .A(u2__abc_52155_new_n23059_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23060_));
AND2X2 AND2X2_11812 ( .A(u2__abc_52155_new_n23057_), .B(u2__abc_52155_new_n23060_), .Y(u2__abc_52155_new_n23061_));
AND2X2 AND2X2_11813 ( .A(u2__abc_52155_new_n23062_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__333_));
AND2X2 AND2X2_11814 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_333_), .Y(u2__abc_52155_new_n23064_));
AND2X2 AND2X2_11815 ( .A(u2__abc_52155_new_n23054_), .B(u2_o_332_), .Y(u2__abc_52155_new_n23066_));
AND2X2 AND2X2_11816 ( .A(u2__abc_52155_new_n23067_), .B(u2__abc_52155_new_n23065_), .Y(u2__abc_52155_new_n23068_));
AND2X2 AND2X2_11817 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6003_), .Y(u2__abc_52155_new_n23070_));
AND2X2 AND2X2_11818 ( .A(u2__abc_52155_new_n23071_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23072_));
AND2X2 AND2X2_11819 ( .A(u2__abc_52155_new_n23069_), .B(u2__abc_52155_new_n23072_), .Y(u2__abc_52155_new_n23073_));
AND2X2 AND2X2_1182 ( .A(u2__abc_52155_new_n4425_), .B(u2__abc_52155_new_n4428_), .Y(u2__abc_52155_new_n4429_));
AND2X2 AND2X2_11820 ( .A(u2__abc_52155_new_n23074_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__334_));
AND2X2 AND2X2_11821 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_334_), .Y(u2__abc_52155_new_n23076_));
AND2X2 AND2X2_11822 ( .A(u2__abc_52155_new_n23066_), .B(u2_o_333_), .Y(u2__abc_52155_new_n23077_));
AND2X2 AND2X2_11823 ( .A(u2__abc_52155_new_n23078_), .B(u2__abc_52155_new_n23079_), .Y(u2__abc_52155_new_n23080_));
AND2X2 AND2X2_11824 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5916_), .Y(u2__abc_52155_new_n23082_));
AND2X2 AND2X2_11825 ( .A(u2__abc_52155_new_n23083_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23084_));
AND2X2 AND2X2_11826 ( .A(u2__abc_52155_new_n23081_), .B(u2__abc_52155_new_n23084_), .Y(u2__abc_52155_new_n23085_));
AND2X2 AND2X2_11827 ( .A(u2__abc_52155_new_n23086_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__335_));
AND2X2 AND2X2_11828 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_335_), .Y(u2__abc_52155_new_n23088_));
AND2X2 AND2X2_11829 ( .A(u2__abc_52155_new_n23077_), .B(u2_o_334_), .Y(u2__abc_52155_new_n23090_));
AND2X2 AND2X2_1183 ( .A(u2__abc_52155_new_n4422_), .B(u2__abc_52155_new_n4429_), .Y(u2__abc_52155_new_n4430_));
AND2X2 AND2X2_11830 ( .A(u2__abc_52155_new_n23091_), .B(u2__abc_52155_new_n23089_), .Y(u2__abc_52155_new_n23092_));
AND2X2 AND2X2_11831 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5923_), .Y(u2__abc_52155_new_n23094_));
AND2X2 AND2X2_11832 ( .A(u2__abc_52155_new_n23095_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23096_));
AND2X2 AND2X2_11833 ( .A(u2__abc_52155_new_n23093_), .B(u2__abc_52155_new_n23096_), .Y(u2__abc_52155_new_n23097_));
AND2X2 AND2X2_11834 ( .A(u2__abc_52155_new_n23098_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__336_));
AND2X2 AND2X2_11835 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_336_), .Y(u2__abc_52155_new_n23100_));
AND2X2 AND2X2_11836 ( .A(u2__abc_52155_new_n23090_), .B(u2_o_335_), .Y(u2__abc_52155_new_n23101_));
AND2X2 AND2X2_11837 ( .A(u2__abc_52155_new_n23102_), .B(u2__abc_52155_new_n23103_), .Y(u2__abc_52155_new_n23104_));
AND2X2 AND2X2_11838 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5901_), .Y(u2__abc_52155_new_n23106_));
AND2X2 AND2X2_11839 ( .A(u2__abc_52155_new_n23107_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23108_));
AND2X2 AND2X2_1184 ( .A(u2__abc_52155_new_n4431_), .B(u2_remHi_235_), .Y(u2__abc_52155_new_n4432_));
AND2X2 AND2X2_11840 ( .A(u2__abc_52155_new_n23105_), .B(u2__abc_52155_new_n23108_), .Y(u2__abc_52155_new_n23109_));
AND2X2 AND2X2_11841 ( .A(u2__abc_52155_new_n23110_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__337_));
AND2X2 AND2X2_11842 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_337_), .Y(u2__abc_52155_new_n23112_));
AND2X2 AND2X2_11843 ( .A(u2__abc_52155_new_n23101_), .B(u2_o_336_), .Y(u2__abc_52155_new_n23114_));
AND2X2 AND2X2_11844 ( .A(u2__abc_52155_new_n23115_), .B(u2__abc_52155_new_n23113_), .Y(u2__abc_52155_new_n23116_));
AND2X2 AND2X2_11845 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5908_), .Y(u2__abc_52155_new_n23118_));
AND2X2 AND2X2_11846 ( .A(u2__abc_52155_new_n23119_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23120_));
AND2X2 AND2X2_11847 ( .A(u2__abc_52155_new_n23117_), .B(u2__abc_52155_new_n23120_), .Y(u2__abc_52155_new_n23121_));
AND2X2 AND2X2_11848 ( .A(u2__abc_52155_new_n23122_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__338_));
AND2X2 AND2X2_11849 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_338_), .Y(u2__abc_52155_new_n23124_));
AND2X2 AND2X2_1185 ( .A(u2__abc_52155_new_n4434_), .B(u2_o_235_), .Y(u2__abc_52155_new_n4435_));
AND2X2 AND2X2_11850 ( .A(u2__abc_52155_new_n23114_), .B(u2_o_337_), .Y(u2__abc_52155_new_n23125_));
AND2X2 AND2X2_11851 ( .A(u2__abc_52155_new_n23126_), .B(u2__abc_52155_new_n23127_), .Y(u2__abc_52155_new_n23128_));
AND2X2 AND2X2_11852 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5947_), .Y(u2__abc_52155_new_n23130_));
AND2X2 AND2X2_11853 ( .A(u2__abc_52155_new_n23131_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23132_));
AND2X2 AND2X2_11854 ( .A(u2__abc_52155_new_n23129_), .B(u2__abc_52155_new_n23132_), .Y(u2__abc_52155_new_n23133_));
AND2X2 AND2X2_11855 ( .A(u2__abc_52155_new_n23134_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__339_));
AND2X2 AND2X2_11856 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_339_), .Y(u2__abc_52155_new_n23136_));
AND2X2 AND2X2_11857 ( .A(u2__abc_52155_new_n23125_), .B(u2_o_338_), .Y(u2__abc_52155_new_n23138_));
AND2X2 AND2X2_11858 ( .A(u2__abc_52155_new_n23139_), .B(u2__abc_52155_new_n23137_), .Y(u2__abc_52155_new_n23140_));
AND2X2 AND2X2_11859 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5954_), .Y(u2__abc_52155_new_n23142_));
AND2X2 AND2X2_1186 ( .A(u2__abc_52155_new_n4433_), .B(u2__abc_52155_new_n4436_), .Y(u2__abc_52155_new_n4437_));
AND2X2 AND2X2_11860 ( .A(u2__abc_52155_new_n23143_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23144_));
AND2X2 AND2X2_11861 ( .A(u2__abc_52155_new_n23141_), .B(u2__abc_52155_new_n23144_), .Y(u2__abc_52155_new_n23145_));
AND2X2 AND2X2_11862 ( .A(u2__abc_52155_new_n23146_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__340_));
AND2X2 AND2X2_11863 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_340_), .Y(u2__abc_52155_new_n23148_));
AND2X2 AND2X2_11864 ( .A(u2__abc_52155_new_n23138_), .B(u2_o_339_), .Y(u2__abc_52155_new_n23150_));
AND2X2 AND2X2_11865 ( .A(u2__abc_52155_new_n23151_), .B(u2__abc_52155_new_n23149_), .Y(u2__abc_52155_new_n23152_));
AND2X2 AND2X2_11866 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5932_), .Y(u2__abc_52155_new_n23154_));
AND2X2 AND2X2_11867 ( .A(u2__abc_52155_new_n23155_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23156_));
AND2X2 AND2X2_11868 ( .A(u2__abc_52155_new_n23153_), .B(u2__abc_52155_new_n23156_), .Y(u2__abc_52155_new_n23157_));
AND2X2 AND2X2_11869 ( .A(u2__abc_52155_new_n23158_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__341_));
AND2X2 AND2X2_1187 ( .A(u2__abc_52155_new_n4438_), .B(u2_remHi_234_), .Y(u2__abc_52155_new_n4439_));
AND2X2 AND2X2_11870 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_341_), .Y(u2__abc_52155_new_n23160_));
AND2X2 AND2X2_11871 ( .A(u2__abc_52155_new_n23150_), .B(u2_o_340_), .Y(u2__abc_52155_new_n23162_));
AND2X2 AND2X2_11872 ( .A(u2__abc_52155_new_n23163_), .B(u2__abc_52155_new_n23161_), .Y(u2__abc_52155_new_n23164_));
AND2X2 AND2X2_11873 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5939_), .Y(u2__abc_52155_new_n23166_));
AND2X2 AND2X2_11874 ( .A(u2__abc_52155_new_n23167_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23168_));
AND2X2 AND2X2_11875 ( .A(u2__abc_52155_new_n23165_), .B(u2__abc_52155_new_n23168_), .Y(u2__abc_52155_new_n23169_));
AND2X2 AND2X2_11876 ( .A(u2__abc_52155_new_n23170_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__342_));
AND2X2 AND2X2_11877 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_342_), .Y(u2__abc_52155_new_n23172_));
AND2X2 AND2X2_11878 ( .A(u2__abc_52155_new_n23162_), .B(u2_o_341_), .Y(u2__abc_52155_new_n23173_));
AND2X2 AND2X2_11879 ( .A(u2__abc_52155_new_n23174_), .B(u2__abc_52155_new_n23175_), .Y(u2__abc_52155_new_n23176_));
AND2X2 AND2X2_1188 ( .A(u2__abc_52155_new_n4441_), .B(u2_o_234_), .Y(u2__abc_52155_new_n4442_));
AND2X2 AND2X2_11880 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5853_), .Y(u2__abc_52155_new_n23178_));
AND2X2 AND2X2_11881 ( .A(u2__abc_52155_new_n23179_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23180_));
AND2X2 AND2X2_11882 ( .A(u2__abc_52155_new_n23177_), .B(u2__abc_52155_new_n23180_), .Y(u2__abc_52155_new_n23181_));
AND2X2 AND2X2_11883 ( .A(u2__abc_52155_new_n23182_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__343_));
AND2X2 AND2X2_11884 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_343_), .Y(u2__abc_52155_new_n23184_));
AND2X2 AND2X2_11885 ( .A(u2__abc_52155_new_n23173_), .B(u2_o_342_), .Y(u2__abc_52155_new_n23186_));
AND2X2 AND2X2_11886 ( .A(u2__abc_52155_new_n23187_), .B(u2__abc_52155_new_n23185_), .Y(u2__abc_52155_new_n23188_));
AND2X2 AND2X2_11887 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5860_), .Y(u2__abc_52155_new_n23190_));
AND2X2 AND2X2_11888 ( .A(u2__abc_52155_new_n23191_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23192_));
AND2X2 AND2X2_11889 ( .A(u2__abc_52155_new_n23189_), .B(u2__abc_52155_new_n23192_), .Y(u2__abc_52155_new_n23193_));
AND2X2 AND2X2_1189 ( .A(u2__abc_52155_new_n4440_), .B(u2__abc_52155_new_n4443_), .Y(u2__abc_52155_new_n4444_));
AND2X2 AND2X2_11890 ( .A(u2__abc_52155_new_n23194_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__344_));
AND2X2 AND2X2_11891 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_344_), .Y(u2__abc_52155_new_n23196_));
AND2X2 AND2X2_11892 ( .A(u2__abc_52155_new_n23186_), .B(u2_o_343_), .Y(u2__abc_52155_new_n23197_));
AND2X2 AND2X2_11893 ( .A(u2__abc_52155_new_n23198_), .B(u2__abc_52155_new_n23199_), .Y(u2__abc_52155_new_n23200_));
AND2X2 AND2X2_11894 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5838_), .Y(u2__abc_52155_new_n23202_));
AND2X2 AND2X2_11895 ( .A(u2__abc_52155_new_n23203_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23204_));
AND2X2 AND2X2_11896 ( .A(u2__abc_52155_new_n23201_), .B(u2__abc_52155_new_n23204_), .Y(u2__abc_52155_new_n23205_));
AND2X2 AND2X2_11897 ( .A(u2__abc_52155_new_n23206_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__345_));
AND2X2 AND2X2_11898 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_345_), .Y(u2__abc_52155_new_n23208_));
AND2X2 AND2X2_11899 ( .A(u2__abc_52155_new_n23197_), .B(u2_o_344_), .Y(u2__abc_52155_new_n23210_));
AND2X2 AND2X2_119 ( .A(_abc_73687_new_n957_), .B(_abc_73687_new_n956_), .Y(\o[154] ));
AND2X2 AND2X2_1190 ( .A(u2__abc_52155_new_n4437_), .B(u2__abc_52155_new_n4444_), .Y(u2__abc_52155_new_n4445_));
AND2X2 AND2X2_11900 ( .A(u2__abc_52155_new_n23211_), .B(u2__abc_52155_new_n23209_), .Y(u2__abc_52155_new_n23212_));
AND2X2 AND2X2_11901 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5845_), .Y(u2__abc_52155_new_n23214_));
AND2X2 AND2X2_11902 ( .A(u2__abc_52155_new_n23215_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23216_));
AND2X2 AND2X2_11903 ( .A(u2__abc_52155_new_n23213_), .B(u2__abc_52155_new_n23216_), .Y(u2__abc_52155_new_n23217_));
AND2X2 AND2X2_11904 ( .A(u2__abc_52155_new_n23218_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__346_));
AND2X2 AND2X2_11905 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_346_), .Y(u2__abc_52155_new_n23220_));
AND2X2 AND2X2_11906 ( .A(u2__abc_52155_new_n23210_), .B(u2_o_345_), .Y(u2__abc_52155_new_n23221_));
AND2X2 AND2X2_11907 ( .A(u2__abc_52155_new_n23222_), .B(u2__abc_52155_new_n23223_), .Y(u2__abc_52155_new_n23224_));
AND2X2 AND2X2_11908 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5884_), .Y(u2__abc_52155_new_n23226_));
AND2X2 AND2X2_11909 ( .A(u2__abc_52155_new_n23227_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23228_));
AND2X2 AND2X2_1191 ( .A(u2__abc_52155_new_n4430_), .B(u2__abc_52155_new_n4445_), .Y(u2__abc_52155_new_n4446_));
AND2X2 AND2X2_11910 ( .A(u2__abc_52155_new_n23225_), .B(u2__abc_52155_new_n23228_), .Y(u2__abc_52155_new_n23229_));
AND2X2 AND2X2_11911 ( .A(u2__abc_52155_new_n23230_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__347_));
AND2X2 AND2X2_11912 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_347_), .Y(u2__abc_52155_new_n23232_));
AND2X2 AND2X2_11913 ( .A(u2__abc_52155_new_n23221_), .B(u2_o_346_), .Y(u2__abc_52155_new_n23234_));
AND2X2 AND2X2_11914 ( .A(u2__abc_52155_new_n23235_), .B(u2__abc_52155_new_n23233_), .Y(u2__abc_52155_new_n23236_));
AND2X2 AND2X2_11915 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5891_), .Y(u2__abc_52155_new_n23238_));
AND2X2 AND2X2_11916 ( .A(u2__abc_52155_new_n23239_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23240_));
AND2X2 AND2X2_11917 ( .A(u2__abc_52155_new_n23237_), .B(u2__abc_52155_new_n23240_), .Y(u2__abc_52155_new_n23241_));
AND2X2 AND2X2_11918 ( .A(u2__abc_52155_new_n23242_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__348_));
AND2X2 AND2X2_11919 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_348_), .Y(u2__abc_52155_new_n23244_));
AND2X2 AND2X2_1192 ( .A(u2__abc_52155_new_n4447_), .B(u2_remHi_232_), .Y(u2__abc_52155_new_n4448_));
AND2X2 AND2X2_11920 ( .A(u2__abc_52155_new_n23234_), .B(u2_o_347_), .Y(u2__abc_52155_new_n23245_));
AND2X2 AND2X2_11921 ( .A(u2__abc_52155_new_n23246_), .B(u2__abc_52155_new_n23247_), .Y(u2__abc_52155_new_n23248_));
AND2X2 AND2X2_11922 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5869_), .Y(u2__abc_52155_new_n23250_));
AND2X2 AND2X2_11923 ( .A(u2__abc_52155_new_n23251_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23252_));
AND2X2 AND2X2_11924 ( .A(u2__abc_52155_new_n23249_), .B(u2__abc_52155_new_n23252_), .Y(u2__abc_52155_new_n23253_));
AND2X2 AND2X2_11925 ( .A(u2__abc_52155_new_n23254_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__349_));
AND2X2 AND2X2_11926 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_349_), .Y(u2__abc_52155_new_n23256_));
AND2X2 AND2X2_11927 ( .A(u2__abc_52155_new_n23245_), .B(u2_o_348_), .Y(u2__abc_52155_new_n23258_));
AND2X2 AND2X2_11928 ( .A(u2__abc_52155_new_n23259_), .B(u2__abc_52155_new_n23257_), .Y(u2__abc_52155_new_n23260_));
AND2X2 AND2X2_11929 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5876_), .Y(u2__abc_52155_new_n23262_));
AND2X2 AND2X2_1193 ( .A(u2__abc_52155_new_n4450_), .B(u2_o_232_), .Y(u2__abc_52155_new_n4451_));
AND2X2 AND2X2_11930 ( .A(u2__abc_52155_new_n23263_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23264_));
AND2X2 AND2X2_11931 ( .A(u2__abc_52155_new_n23261_), .B(u2__abc_52155_new_n23264_), .Y(u2__abc_52155_new_n23265_));
AND2X2 AND2X2_11932 ( .A(u2__abc_52155_new_n23266_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__350_));
AND2X2 AND2X2_11933 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_350_), .Y(u2__abc_52155_new_n23268_));
AND2X2 AND2X2_11934 ( .A(u2__abc_52155_new_n23258_), .B(u2_o_349_), .Y(u2__abc_52155_new_n23269_));
AND2X2 AND2X2_11935 ( .A(u2__abc_52155_new_n23270_), .B(u2__abc_52155_new_n23271_), .Y(u2__abc_52155_new_n23272_));
AND2X2 AND2X2_11936 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5788_), .Y(u2__abc_52155_new_n23274_));
AND2X2 AND2X2_11937 ( .A(u2__abc_52155_new_n23275_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23276_));
AND2X2 AND2X2_11938 ( .A(u2__abc_52155_new_n23273_), .B(u2__abc_52155_new_n23276_), .Y(u2__abc_52155_new_n23277_));
AND2X2 AND2X2_11939 ( .A(u2__abc_52155_new_n23278_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__351_));
AND2X2 AND2X2_1194 ( .A(u2__abc_52155_new_n4449_), .B(u2__abc_52155_new_n4452_), .Y(u2__abc_52155_new_n4453_));
AND2X2 AND2X2_11940 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_351_), .Y(u2__abc_52155_new_n23280_));
AND2X2 AND2X2_11941 ( .A(u2__abc_52155_new_n23269_), .B(u2_o_350_), .Y(u2__abc_52155_new_n23282_));
AND2X2 AND2X2_11942 ( .A(u2__abc_52155_new_n23283_), .B(u2__abc_52155_new_n23281_), .Y(u2__abc_52155_new_n23284_));
AND2X2 AND2X2_11943 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5795_), .Y(u2__abc_52155_new_n23286_));
AND2X2 AND2X2_11944 ( .A(u2__abc_52155_new_n23287_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23288_));
AND2X2 AND2X2_11945 ( .A(u2__abc_52155_new_n23285_), .B(u2__abc_52155_new_n23288_), .Y(u2__abc_52155_new_n23289_));
AND2X2 AND2X2_11946 ( .A(u2__abc_52155_new_n23290_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__352_));
AND2X2 AND2X2_11947 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_352_), .Y(u2__abc_52155_new_n23292_));
AND2X2 AND2X2_11948 ( .A(u2__abc_52155_new_n23282_), .B(u2_o_351_), .Y(u2__abc_52155_new_n23293_));
AND2X2 AND2X2_11949 ( .A(u2__abc_52155_new_n23294_), .B(u2__abc_52155_new_n23295_), .Y(u2__abc_52155_new_n23296_));
AND2X2 AND2X2_1195 ( .A(u2__abc_52155_new_n4454_), .B(u2_remHi_233_), .Y(u2__abc_52155_new_n4455_));
AND2X2 AND2X2_11950 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5773_), .Y(u2__abc_52155_new_n23298_));
AND2X2 AND2X2_11951 ( .A(u2__abc_52155_new_n23299_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23300_));
AND2X2 AND2X2_11952 ( .A(u2__abc_52155_new_n23297_), .B(u2__abc_52155_new_n23300_), .Y(u2__abc_52155_new_n23301_));
AND2X2 AND2X2_11953 ( .A(u2__abc_52155_new_n23302_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__353_));
AND2X2 AND2X2_11954 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_353_), .Y(u2__abc_52155_new_n23304_));
AND2X2 AND2X2_11955 ( .A(u2__abc_52155_new_n23293_), .B(u2_o_352_), .Y(u2__abc_52155_new_n23306_));
AND2X2 AND2X2_11956 ( .A(u2__abc_52155_new_n23307_), .B(u2__abc_52155_new_n23305_), .Y(u2__abc_52155_new_n23308_));
AND2X2 AND2X2_11957 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5780_), .Y(u2__abc_52155_new_n23310_));
AND2X2 AND2X2_11958 ( .A(u2__abc_52155_new_n23311_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23312_));
AND2X2 AND2X2_11959 ( .A(u2__abc_52155_new_n23309_), .B(u2__abc_52155_new_n23312_), .Y(u2__abc_52155_new_n23313_));
AND2X2 AND2X2_1196 ( .A(u2__abc_52155_new_n4457_), .B(u2_o_233_), .Y(u2__abc_52155_new_n4458_));
AND2X2 AND2X2_11960 ( .A(u2__abc_52155_new_n23314_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__354_));
AND2X2 AND2X2_11961 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_354_), .Y(u2__abc_52155_new_n23316_));
AND2X2 AND2X2_11962 ( .A(u2__abc_52155_new_n23306_), .B(u2_o_353_), .Y(u2__abc_52155_new_n23317_));
AND2X2 AND2X2_11963 ( .A(u2__abc_52155_new_n23318_), .B(u2__abc_52155_new_n23319_), .Y(u2__abc_52155_new_n23320_));
AND2X2 AND2X2_11964 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5819_), .Y(u2__abc_52155_new_n23322_));
AND2X2 AND2X2_11965 ( .A(u2__abc_52155_new_n23323_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23324_));
AND2X2 AND2X2_11966 ( .A(u2__abc_52155_new_n23321_), .B(u2__abc_52155_new_n23324_), .Y(u2__abc_52155_new_n23325_));
AND2X2 AND2X2_11967 ( .A(u2__abc_52155_new_n23326_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__355_));
AND2X2 AND2X2_11968 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_355_), .Y(u2__abc_52155_new_n23328_));
AND2X2 AND2X2_11969 ( .A(u2__abc_52155_new_n23317_), .B(u2_o_354_), .Y(u2__abc_52155_new_n23330_));
AND2X2 AND2X2_1197 ( .A(u2__abc_52155_new_n4456_), .B(u2__abc_52155_new_n4459_), .Y(u2__abc_52155_new_n4460_));
AND2X2 AND2X2_11970 ( .A(u2__abc_52155_new_n23331_), .B(u2__abc_52155_new_n23329_), .Y(u2__abc_52155_new_n23332_));
AND2X2 AND2X2_11971 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5826_), .Y(u2__abc_52155_new_n23334_));
AND2X2 AND2X2_11972 ( .A(u2__abc_52155_new_n23335_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23336_));
AND2X2 AND2X2_11973 ( .A(u2__abc_52155_new_n23333_), .B(u2__abc_52155_new_n23336_), .Y(u2__abc_52155_new_n23337_));
AND2X2 AND2X2_11974 ( .A(u2__abc_52155_new_n23338_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__356_));
AND2X2 AND2X2_11975 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_356_), .Y(u2__abc_52155_new_n23340_));
AND2X2 AND2X2_11976 ( .A(u2__abc_52155_new_n23330_), .B(u2_o_355_), .Y(u2__abc_52155_new_n23342_));
AND2X2 AND2X2_11977 ( .A(u2__abc_52155_new_n23343_), .B(u2__abc_52155_new_n23341_), .Y(u2__abc_52155_new_n23344_));
AND2X2 AND2X2_11978 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5804_), .Y(u2__abc_52155_new_n23346_));
AND2X2 AND2X2_11979 ( .A(u2__abc_52155_new_n23347_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23348_));
AND2X2 AND2X2_1198 ( .A(u2__abc_52155_new_n4453_), .B(u2__abc_52155_new_n4460_), .Y(u2__abc_52155_new_n4461_));
AND2X2 AND2X2_11980 ( .A(u2__abc_52155_new_n23345_), .B(u2__abc_52155_new_n23348_), .Y(u2__abc_52155_new_n23349_));
AND2X2 AND2X2_11981 ( .A(u2__abc_52155_new_n23350_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__357_));
AND2X2 AND2X2_11982 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_357_), .Y(u2__abc_52155_new_n23352_));
AND2X2 AND2X2_11983 ( .A(u2__abc_52155_new_n23342_), .B(u2_o_356_), .Y(u2__abc_52155_new_n23354_));
AND2X2 AND2X2_11984 ( .A(u2__abc_52155_new_n23355_), .B(u2__abc_52155_new_n23353_), .Y(u2__abc_52155_new_n23356_));
AND2X2 AND2X2_11985 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5811_), .Y(u2__abc_52155_new_n23358_));
AND2X2 AND2X2_11986 ( .A(u2__abc_52155_new_n23359_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23360_));
AND2X2 AND2X2_11987 ( .A(u2__abc_52155_new_n23357_), .B(u2__abc_52155_new_n23360_), .Y(u2__abc_52155_new_n23361_));
AND2X2 AND2X2_11988 ( .A(u2__abc_52155_new_n23362_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__358_));
AND2X2 AND2X2_11989 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_358_), .Y(u2__abc_52155_new_n23364_));
AND2X2 AND2X2_1199 ( .A(u2__abc_52155_new_n4462_), .B(u2_remHi_231_), .Y(u2__abc_52155_new_n4463_));
AND2X2 AND2X2_11990 ( .A(u2__abc_52155_new_n23354_), .B(u2_o_357_), .Y(u2__abc_52155_new_n23365_));
AND2X2 AND2X2_11991 ( .A(u2__abc_52155_new_n23366_), .B(u2__abc_52155_new_n23367_), .Y(u2__abc_52155_new_n23368_));
AND2X2 AND2X2_11992 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5713_), .Y(u2__abc_52155_new_n23370_));
AND2X2 AND2X2_11993 ( .A(u2__abc_52155_new_n23371_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23372_));
AND2X2 AND2X2_11994 ( .A(u2__abc_52155_new_n23369_), .B(u2__abc_52155_new_n23372_), .Y(u2__abc_52155_new_n23373_));
AND2X2 AND2X2_11995 ( .A(u2__abc_52155_new_n23374_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__359_));
AND2X2 AND2X2_11996 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_359_), .Y(u2__abc_52155_new_n23376_));
AND2X2 AND2X2_11997 ( .A(u2__abc_52155_new_n23365_), .B(u2_o_358_), .Y(u2__abc_52155_new_n23378_));
AND2X2 AND2X2_11998 ( .A(u2__abc_52155_new_n23379_), .B(u2__abc_52155_new_n23377_), .Y(u2__abc_52155_new_n23380_));
AND2X2 AND2X2_11999 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5720_), .Y(u2__abc_52155_new_n23382_));
AND2X2 AND2X2_12 ( .A(_abc_73687_new_n753_), .B(sqrto_11_), .Y(\o[47] ));
AND2X2 AND2X2_120 ( .A(_abc_73687_new_n960_), .B(_abc_73687_new_n959_), .Y(\o[155] ));
AND2X2 AND2X2_1200 ( .A(u2__abc_52155_new_n4465_), .B(u2_o_231_), .Y(u2__abc_52155_new_n4466_));
AND2X2 AND2X2_12000 ( .A(u2__abc_52155_new_n23383_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23384_));
AND2X2 AND2X2_12001 ( .A(u2__abc_52155_new_n23381_), .B(u2__abc_52155_new_n23384_), .Y(u2__abc_52155_new_n23385_));
AND2X2 AND2X2_12002 ( .A(u2__abc_52155_new_n23386_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__360_));
AND2X2 AND2X2_12003 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_360_), .Y(u2__abc_52155_new_n23388_));
AND2X2 AND2X2_12004 ( .A(u2__abc_52155_new_n23378_), .B(u2_o_359_), .Y(u2__abc_52155_new_n23389_));
AND2X2 AND2X2_12005 ( .A(u2__abc_52155_new_n23390_), .B(u2__abc_52155_new_n23391_), .Y(u2__abc_52155_new_n23392_));
AND2X2 AND2X2_12006 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5725_), .Y(u2__abc_52155_new_n23394_));
AND2X2 AND2X2_12007 ( .A(u2__abc_52155_new_n23395_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23396_));
AND2X2 AND2X2_12008 ( .A(u2__abc_52155_new_n23393_), .B(u2__abc_52155_new_n23396_), .Y(u2__abc_52155_new_n23397_));
AND2X2 AND2X2_12009 ( .A(u2__abc_52155_new_n23398_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__361_));
AND2X2 AND2X2_1201 ( .A(u2__abc_52155_new_n4464_), .B(u2__abc_52155_new_n4467_), .Y(u2__abc_52155_new_n4468_));
AND2X2 AND2X2_12010 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_361_), .Y(u2__abc_52155_new_n23400_));
AND2X2 AND2X2_12011 ( .A(u2__abc_52155_new_n23389_), .B(u2_o_360_), .Y(u2__abc_52155_new_n23402_));
AND2X2 AND2X2_12012 ( .A(u2__abc_52155_new_n23403_), .B(u2__abc_52155_new_n23401_), .Y(u2__abc_52155_new_n23404_));
AND2X2 AND2X2_12013 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5732_), .Y(u2__abc_52155_new_n23406_));
AND2X2 AND2X2_12014 ( .A(u2__abc_52155_new_n23407_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23408_));
AND2X2 AND2X2_12015 ( .A(u2__abc_52155_new_n23405_), .B(u2__abc_52155_new_n23408_), .Y(u2__abc_52155_new_n23409_));
AND2X2 AND2X2_12016 ( .A(u2__abc_52155_new_n23410_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__362_));
AND2X2 AND2X2_12017 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_362_), .Y(u2__abc_52155_new_n23412_));
AND2X2 AND2X2_12018 ( .A(u2__abc_52155_new_n23402_), .B(u2_o_361_), .Y(u2__abc_52155_new_n23413_));
AND2X2 AND2X2_12019 ( .A(u2__abc_52155_new_n23414_), .B(u2__abc_52155_new_n23415_), .Y(u2__abc_52155_new_n23416_));
AND2X2 AND2X2_1202 ( .A(u2__abc_52155_new_n4469_), .B(u2_remHi_230_), .Y(u2__abc_52155_new_n4470_));
AND2X2 AND2X2_12020 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5756_), .Y(u2__abc_52155_new_n23418_));
AND2X2 AND2X2_12021 ( .A(u2__abc_52155_new_n23419_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23420_));
AND2X2 AND2X2_12022 ( .A(u2__abc_52155_new_n23417_), .B(u2__abc_52155_new_n23420_), .Y(u2__abc_52155_new_n23421_));
AND2X2 AND2X2_12023 ( .A(u2__abc_52155_new_n23422_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__363_));
AND2X2 AND2X2_12024 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_363_), .Y(u2__abc_52155_new_n23424_));
AND2X2 AND2X2_12025 ( .A(u2__abc_52155_new_n23413_), .B(u2_o_362_), .Y(u2__abc_52155_new_n23426_));
AND2X2 AND2X2_12026 ( .A(u2__abc_52155_new_n23427_), .B(u2__abc_52155_new_n23425_), .Y(u2__abc_52155_new_n23428_));
AND2X2 AND2X2_12027 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5763_), .Y(u2__abc_52155_new_n23430_));
AND2X2 AND2X2_12028 ( .A(u2__abc_52155_new_n23431_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23432_));
AND2X2 AND2X2_12029 ( .A(u2__abc_52155_new_n23429_), .B(u2__abc_52155_new_n23432_), .Y(u2__abc_52155_new_n23433_));
AND2X2 AND2X2_1203 ( .A(u2__abc_52155_new_n4472_), .B(u2_o_230_), .Y(u2__abc_52155_new_n4473_));
AND2X2 AND2X2_12030 ( .A(u2__abc_52155_new_n23434_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__364_));
AND2X2 AND2X2_12031 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_364_), .Y(u2__abc_52155_new_n23436_));
AND2X2 AND2X2_12032 ( .A(u2__abc_52155_new_n23426_), .B(u2_o_363_), .Y(u2__abc_52155_new_n23437_));
AND2X2 AND2X2_12033 ( .A(u2__abc_52155_new_n23438_), .B(u2__abc_52155_new_n23439_), .Y(u2__abc_52155_new_n23440_));
AND2X2 AND2X2_12034 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5741_), .Y(u2__abc_52155_new_n23442_));
AND2X2 AND2X2_12035 ( .A(u2__abc_52155_new_n23443_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23444_));
AND2X2 AND2X2_12036 ( .A(u2__abc_52155_new_n23441_), .B(u2__abc_52155_new_n23444_), .Y(u2__abc_52155_new_n23445_));
AND2X2 AND2X2_12037 ( .A(u2__abc_52155_new_n23446_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__365_));
AND2X2 AND2X2_12038 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_365_), .Y(u2__abc_52155_new_n23448_));
AND2X2 AND2X2_12039 ( .A(u2__abc_52155_new_n23437_), .B(u2_o_364_), .Y(u2__abc_52155_new_n23450_));
AND2X2 AND2X2_1204 ( .A(u2__abc_52155_new_n4471_), .B(u2__abc_52155_new_n4474_), .Y(u2__abc_52155_new_n4475_));
AND2X2 AND2X2_12040 ( .A(u2__abc_52155_new_n23451_), .B(u2__abc_52155_new_n23449_), .Y(u2__abc_52155_new_n23452_));
AND2X2 AND2X2_12041 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5748_), .Y(u2__abc_52155_new_n23454_));
AND2X2 AND2X2_12042 ( .A(u2__abc_52155_new_n23455_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23456_));
AND2X2 AND2X2_12043 ( .A(u2__abc_52155_new_n23453_), .B(u2__abc_52155_new_n23456_), .Y(u2__abc_52155_new_n23457_));
AND2X2 AND2X2_12044 ( .A(u2__abc_52155_new_n23458_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__366_));
AND2X2 AND2X2_12045 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_366_), .Y(u2__abc_52155_new_n23460_));
AND2X2 AND2X2_12046 ( .A(u2__abc_52155_new_n23450_), .B(u2_o_365_), .Y(u2__abc_52155_new_n23461_));
AND2X2 AND2X2_12047 ( .A(u2__abc_52155_new_n23462_), .B(u2__abc_52155_new_n23463_), .Y(u2__abc_52155_new_n23464_));
AND2X2 AND2X2_12048 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5661_), .Y(u2__abc_52155_new_n23466_));
AND2X2 AND2X2_12049 ( .A(u2__abc_52155_new_n23467_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23468_));
AND2X2 AND2X2_1205 ( .A(u2__abc_52155_new_n4468_), .B(u2__abc_52155_new_n4475_), .Y(u2__abc_52155_new_n4476_));
AND2X2 AND2X2_12050 ( .A(u2__abc_52155_new_n23465_), .B(u2__abc_52155_new_n23468_), .Y(u2__abc_52155_new_n23469_));
AND2X2 AND2X2_12051 ( .A(u2__abc_52155_new_n23470_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__367_));
AND2X2 AND2X2_12052 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_367_), .Y(u2__abc_52155_new_n23472_));
AND2X2 AND2X2_12053 ( .A(u2__abc_52155_new_n23461_), .B(u2_o_366_), .Y(u2__abc_52155_new_n23474_));
AND2X2 AND2X2_12054 ( .A(u2__abc_52155_new_n23475_), .B(u2__abc_52155_new_n23473_), .Y(u2__abc_52155_new_n23476_));
AND2X2 AND2X2_12055 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5668_), .Y(u2__abc_52155_new_n23478_));
AND2X2 AND2X2_12056 ( .A(u2__abc_52155_new_n23479_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23480_));
AND2X2 AND2X2_12057 ( .A(u2__abc_52155_new_n23477_), .B(u2__abc_52155_new_n23480_), .Y(u2__abc_52155_new_n23481_));
AND2X2 AND2X2_12058 ( .A(u2__abc_52155_new_n23482_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__368_));
AND2X2 AND2X2_12059 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_368_), .Y(u2__abc_52155_new_n23484_));
AND2X2 AND2X2_1206 ( .A(u2__abc_52155_new_n4461_), .B(u2__abc_52155_new_n4476_), .Y(u2__abc_52155_new_n4477_));
AND2X2 AND2X2_12060 ( .A(u2__abc_52155_new_n23474_), .B(u2_o_367_), .Y(u2__abc_52155_new_n23485_));
AND2X2 AND2X2_12061 ( .A(u2__abc_52155_new_n23486_), .B(u2__abc_52155_new_n23487_), .Y(u2__abc_52155_new_n23488_));
AND2X2 AND2X2_12062 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5646_), .Y(u2__abc_52155_new_n23490_));
AND2X2 AND2X2_12063 ( .A(u2__abc_52155_new_n23491_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23492_));
AND2X2 AND2X2_12064 ( .A(u2__abc_52155_new_n23489_), .B(u2__abc_52155_new_n23492_), .Y(u2__abc_52155_new_n23493_));
AND2X2 AND2X2_12065 ( .A(u2__abc_52155_new_n23494_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__369_));
AND2X2 AND2X2_12066 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_369_), .Y(u2__abc_52155_new_n23496_));
AND2X2 AND2X2_12067 ( .A(u2__abc_52155_new_n23485_), .B(u2_o_368_), .Y(u2__abc_52155_new_n23498_));
AND2X2 AND2X2_12068 ( .A(u2__abc_52155_new_n23499_), .B(u2__abc_52155_new_n23497_), .Y(u2__abc_52155_new_n23500_));
AND2X2 AND2X2_12069 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5653_), .Y(u2__abc_52155_new_n23502_));
AND2X2 AND2X2_1207 ( .A(u2__abc_52155_new_n4446_), .B(u2__abc_52155_new_n4477_), .Y(u2__abc_52155_new_n4478_));
AND2X2 AND2X2_12070 ( .A(u2__abc_52155_new_n23503_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23504_));
AND2X2 AND2X2_12071 ( .A(u2__abc_52155_new_n23501_), .B(u2__abc_52155_new_n23504_), .Y(u2__abc_52155_new_n23505_));
AND2X2 AND2X2_12072 ( .A(u2__abc_52155_new_n23506_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__370_));
AND2X2 AND2X2_12073 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_370_), .Y(u2__abc_52155_new_n23508_));
AND2X2 AND2X2_12074 ( .A(u2__abc_52155_new_n23498_), .B(u2_o_369_), .Y(u2__abc_52155_new_n23509_));
AND2X2 AND2X2_12075 ( .A(u2__abc_52155_new_n23510_), .B(u2__abc_52155_new_n23511_), .Y(u2__abc_52155_new_n23512_));
AND2X2 AND2X2_12076 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5699_), .Y(u2__abc_52155_new_n23514_));
AND2X2 AND2X2_12077 ( .A(u2__abc_52155_new_n23515_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23516_));
AND2X2 AND2X2_12078 ( .A(u2__abc_52155_new_n23513_), .B(u2__abc_52155_new_n23516_), .Y(u2__abc_52155_new_n23517_));
AND2X2 AND2X2_12079 ( .A(u2__abc_52155_new_n23518_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__371_));
AND2X2 AND2X2_1208 ( .A(u2__abc_52155_new_n4479_), .B(u2_remHi_224_), .Y(u2__abc_52155_new_n4480_));
AND2X2 AND2X2_12080 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_371_), .Y(u2__abc_52155_new_n23520_));
AND2X2 AND2X2_12081 ( .A(u2__abc_52155_new_n23509_), .B(u2_o_370_), .Y(u2__abc_52155_new_n23522_));
AND2X2 AND2X2_12082 ( .A(u2__abc_52155_new_n23523_), .B(u2__abc_52155_new_n23521_), .Y(u2__abc_52155_new_n23524_));
AND2X2 AND2X2_12083 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5692_), .Y(u2__abc_52155_new_n23526_));
AND2X2 AND2X2_12084 ( .A(u2__abc_52155_new_n23527_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23528_));
AND2X2 AND2X2_12085 ( .A(u2__abc_52155_new_n23525_), .B(u2__abc_52155_new_n23528_), .Y(u2__abc_52155_new_n23529_));
AND2X2 AND2X2_12086 ( .A(u2__abc_52155_new_n23530_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__372_));
AND2X2 AND2X2_12087 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_372_), .Y(u2__abc_52155_new_n23532_));
AND2X2 AND2X2_12088 ( .A(u2__abc_52155_new_n23522_), .B(u2_o_371_), .Y(u2__abc_52155_new_n23533_));
AND2X2 AND2X2_12089 ( .A(u2__abc_52155_new_n23534_), .B(u2__abc_52155_new_n23535_), .Y(u2__abc_52155_new_n23536_));
AND2X2 AND2X2_1209 ( .A(u2__abc_52155_new_n4482_), .B(sqrto_224_), .Y(u2__abc_52155_new_n4483_));
AND2X2 AND2X2_12090 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5677_), .Y(u2__abc_52155_new_n23538_));
AND2X2 AND2X2_12091 ( .A(u2__abc_52155_new_n23539_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23540_));
AND2X2 AND2X2_12092 ( .A(u2__abc_52155_new_n23537_), .B(u2__abc_52155_new_n23540_), .Y(u2__abc_52155_new_n23541_));
AND2X2 AND2X2_12093 ( .A(u2__abc_52155_new_n23542_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__373_));
AND2X2 AND2X2_12094 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_373_), .Y(u2__abc_52155_new_n23544_));
AND2X2 AND2X2_12095 ( .A(u2__abc_52155_new_n23533_), .B(u2_o_372_), .Y(u2__abc_52155_new_n23546_));
AND2X2 AND2X2_12096 ( .A(u2__abc_52155_new_n23547_), .B(u2__abc_52155_new_n23545_), .Y(u2__abc_52155_new_n23548_));
AND2X2 AND2X2_12097 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5684_), .Y(u2__abc_52155_new_n23550_));
AND2X2 AND2X2_12098 ( .A(u2__abc_52155_new_n23551_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23552_));
AND2X2 AND2X2_12099 ( .A(u2__abc_52155_new_n23549_), .B(u2__abc_52155_new_n23552_), .Y(u2__abc_52155_new_n23553_));
AND2X2 AND2X2_121 ( .A(_abc_73687_new_n963_), .B(_abc_73687_new_n962_), .Y(\o[156] ));
AND2X2 AND2X2_1210 ( .A(u2__abc_52155_new_n4481_), .B(u2__abc_52155_new_n4484_), .Y(u2__abc_52155_new_n4485_));
AND2X2 AND2X2_12100 ( .A(u2__abc_52155_new_n23554_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__374_));
AND2X2 AND2X2_12101 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_374_), .Y(u2__abc_52155_new_n23556_));
AND2X2 AND2X2_12102 ( .A(u2__abc_52155_new_n23546_), .B(u2_o_373_), .Y(u2__abc_52155_new_n23557_));
AND2X2 AND2X2_12103 ( .A(u2__abc_52155_new_n23558_), .B(u2__abc_52155_new_n23559_), .Y(u2__abc_52155_new_n23560_));
AND2X2 AND2X2_12104 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5617_), .Y(u2__abc_52155_new_n23562_));
AND2X2 AND2X2_12105 ( .A(u2__abc_52155_new_n23563_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23564_));
AND2X2 AND2X2_12106 ( .A(u2__abc_52155_new_n23561_), .B(u2__abc_52155_new_n23564_), .Y(u2__abc_52155_new_n23565_));
AND2X2 AND2X2_12107 ( .A(u2__abc_52155_new_n23566_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__375_));
AND2X2 AND2X2_12108 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_375_), .Y(u2__abc_52155_new_n23568_));
AND2X2 AND2X2_12109 ( .A(u2__abc_52155_new_n23557_), .B(u2_o_374_), .Y(u2__abc_52155_new_n23570_));
AND2X2 AND2X2_1211 ( .A(u2__abc_52155_new_n4486_), .B(u2_remHi_225_), .Y(u2__abc_52155_new_n4487_));
AND2X2 AND2X2_12110 ( .A(u2__abc_52155_new_n23571_), .B(u2__abc_52155_new_n23569_), .Y(u2__abc_52155_new_n23572_));
AND2X2 AND2X2_12111 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5624_), .Y(u2__abc_52155_new_n23574_));
AND2X2 AND2X2_12112 ( .A(u2__abc_52155_new_n23575_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23576_));
AND2X2 AND2X2_12113 ( .A(u2__abc_52155_new_n23573_), .B(u2__abc_52155_new_n23576_), .Y(u2__abc_52155_new_n23577_));
AND2X2 AND2X2_12114 ( .A(u2__abc_52155_new_n23578_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__376_));
AND2X2 AND2X2_12115 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_376_), .Y(u2__abc_52155_new_n23580_));
AND2X2 AND2X2_12116 ( .A(u2__abc_52155_new_n23570_), .B(u2_o_375_), .Y(u2__abc_52155_new_n23581_));
AND2X2 AND2X2_12117 ( .A(u2__abc_52155_new_n23582_), .B(u2__abc_52155_new_n23583_), .Y(u2__abc_52155_new_n23584_));
AND2X2 AND2X2_12118 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5629_), .Y(u2__abc_52155_new_n23586_));
AND2X2 AND2X2_12119 ( .A(u2__abc_52155_new_n23587_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23588_));
AND2X2 AND2X2_1212 ( .A(u2__abc_52155_new_n4489_), .B(sqrto_225_), .Y(u2__abc_52155_new_n4490_));
AND2X2 AND2X2_12120 ( .A(u2__abc_52155_new_n23585_), .B(u2__abc_52155_new_n23588_), .Y(u2__abc_52155_new_n23589_));
AND2X2 AND2X2_12121 ( .A(u2__abc_52155_new_n23590_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__377_));
AND2X2 AND2X2_12122 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_377_), .Y(u2__abc_52155_new_n23592_));
AND2X2 AND2X2_12123 ( .A(u2__abc_52155_new_n23581_), .B(u2_o_376_), .Y(u2__abc_52155_new_n23594_));
AND2X2 AND2X2_12124 ( .A(u2__abc_52155_new_n23595_), .B(u2__abc_52155_new_n23593_), .Y(u2__abc_52155_new_n23596_));
AND2X2 AND2X2_12125 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5636_), .Y(u2__abc_52155_new_n23598_));
AND2X2 AND2X2_12126 ( .A(u2__abc_52155_new_n23599_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23600_));
AND2X2 AND2X2_12127 ( .A(u2__abc_52155_new_n23597_), .B(u2__abc_52155_new_n23600_), .Y(u2__abc_52155_new_n23601_));
AND2X2 AND2X2_12128 ( .A(u2__abc_52155_new_n23602_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__378_));
AND2X2 AND2X2_12129 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_378_), .Y(u2__abc_52155_new_n23604_));
AND2X2 AND2X2_1213 ( .A(u2__abc_52155_new_n4488_), .B(u2__abc_52155_new_n4491_), .Y(u2__abc_52155_new_n4492_));
AND2X2 AND2X2_12130 ( .A(u2__abc_52155_new_n23594_), .B(u2_o_377_), .Y(u2__abc_52155_new_n23605_));
AND2X2 AND2X2_12131 ( .A(u2__abc_52155_new_n23606_), .B(u2__abc_52155_new_n23607_), .Y(u2__abc_52155_new_n23608_));
AND2X2 AND2X2_12132 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5598_), .Y(u2__abc_52155_new_n23610_));
AND2X2 AND2X2_12133 ( .A(u2__abc_52155_new_n23611_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23612_));
AND2X2 AND2X2_12134 ( .A(u2__abc_52155_new_n23609_), .B(u2__abc_52155_new_n23612_), .Y(u2__abc_52155_new_n23613_));
AND2X2 AND2X2_12135 ( .A(u2__abc_52155_new_n23614_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__379_));
AND2X2 AND2X2_12136 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_379_), .Y(u2__abc_52155_new_n23616_));
AND2X2 AND2X2_12137 ( .A(u2__abc_52155_new_n23605_), .B(u2_o_378_), .Y(u2__abc_52155_new_n23618_));
AND2X2 AND2X2_12138 ( .A(u2__abc_52155_new_n23619_), .B(u2__abc_52155_new_n23617_), .Y(u2__abc_52155_new_n23620_));
AND2X2 AND2X2_12139 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5605_), .Y(u2__abc_52155_new_n23622_));
AND2X2 AND2X2_1214 ( .A(u2__abc_52155_new_n4485_), .B(u2__abc_52155_new_n4492_), .Y(u2__abc_52155_new_n4493_));
AND2X2 AND2X2_12140 ( .A(u2__abc_52155_new_n23623_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23624_));
AND2X2 AND2X2_12141 ( .A(u2__abc_52155_new_n23621_), .B(u2__abc_52155_new_n23624_), .Y(u2__abc_52155_new_n23625_));
AND2X2 AND2X2_12142 ( .A(u2__abc_52155_new_n23626_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__380_));
AND2X2 AND2X2_12143 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_380_), .Y(u2__abc_52155_new_n23628_));
AND2X2 AND2X2_12144 ( .A(u2__abc_52155_new_n23618_), .B(u2_o_379_), .Y(u2__abc_52155_new_n23629_));
AND2X2 AND2X2_12145 ( .A(u2__abc_52155_new_n23630_), .B(u2__abc_52155_new_n23631_), .Y(u2__abc_52155_new_n23632_));
AND2X2 AND2X2_12146 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5583_), .Y(u2__abc_52155_new_n23634_));
AND2X2 AND2X2_12147 ( .A(u2__abc_52155_new_n23635_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23636_));
AND2X2 AND2X2_12148 ( .A(u2__abc_52155_new_n23633_), .B(u2__abc_52155_new_n23636_), .Y(u2__abc_52155_new_n23637_));
AND2X2 AND2X2_12149 ( .A(u2__abc_52155_new_n23638_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__381_));
AND2X2 AND2X2_1215 ( .A(u2__abc_52155_new_n4494_), .B(u2_remHi_223_), .Y(u2__abc_52155_new_n4495_));
AND2X2 AND2X2_12150 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_381_), .Y(u2__abc_52155_new_n23640_));
AND2X2 AND2X2_12151 ( .A(u2__abc_52155_new_n23629_), .B(u2_o_380_), .Y(u2__abc_52155_new_n23642_));
AND2X2 AND2X2_12152 ( .A(u2__abc_52155_new_n23643_), .B(u2__abc_52155_new_n23641_), .Y(u2__abc_52155_new_n23644_));
AND2X2 AND2X2_12153 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5593_), .Y(u2__abc_52155_new_n23646_));
AND2X2 AND2X2_12154 ( .A(u2__abc_52155_new_n23647_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23648_));
AND2X2 AND2X2_12155 ( .A(u2__abc_52155_new_n23645_), .B(u2__abc_52155_new_n23648_), .Y(u2__abc_52155_new_n23649_));
AND2X2 AND2X2_12156 ( .A(u2__abc_52155_new_n23650_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__382_));
AND2X2 AND2X2_12157 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_382_), .Y(u2__abc_52155_new_n23652_));
AND2X2 AND2X2_12158 ( .A(u2__abc_52155_new_n23642_), .B(u2_o_381_), .Y(u2__abc_52155_new_n23653_));
AND2X2 AND2X2_12159 ( .A(u2__abc_52155_new_n23654_), .B(u2__abc_52155_new_n23655_), .Y(u2__abc_52155_new_n23656_));
AND2X2 AND2X2_1216 ( .A(u2__abc_52155_new_n4497_), .B(sqrto_223_), .Y(u2__abc_52155_new_n4498_));
AND2X2 AND2X2_12160 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7235_), .Y(u2__abc_52155_new_n23658_));
AND2X2 AND2X2_12161 ( .A(u2__abc_52155_new_n23659_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23660_));
AND2X2 AND2X2_12162 ( .A(u2__abc_52155_new_n23657_), .B(u2__abc_52155_new_n23660_), .Y(u2__abc_52155_new_n23661_));
AND2X2 AND2X2_12163 ( .A(u2__abc_52155_new_n23662_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__383_));
AND2X2 AND2X2_12164 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_383_), .Y(u2__abc_52155_new_n23664_));
AND2X2 AND2X2_12165 ( .A(u2__abc_52155_new_n23653_), .B(u2_o_382_), .Y(u2__abc_52155_new_n23666_));
AND2X2 AND2X2_12166 ( .A(u2__abc_52155_new_n23667_), .B(u2__abc_52155_new_n23665_), .Y(u2__abc_52155_new_n23668_));
AND2X2 AND2X2_12167 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7231_), .Y(u2__abc_52155_new_n23670_));
AND2X2 AND2X2_12168 ( .A(u2__abc_52155_new_n23671_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23672_));
AND2X2 AND2X2_12169 ( .A(u2__abc_52155_new_n23669_), .B(u2__abc_52155_new_n23672_), .Y(u2__abc_52155_new_n23673_));
AND2X2 AND2X2_1217 ( .A(u2__abc_52155_new_n4496_), .B(u2__abc_52155_new_n4499_), .Y(u2__abc_52155_new_n4500_));
AND2X2 AND2X2_12170 ( .A(u2__abc_52155_new_n23674_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__384_));
AND2X2 AND2X2_12171 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_384_), .Y(u2__abc_52155_new_n23676_));
AND2X2 AND2X2_12172 ( .A(u2__abc_52155_new_n23666_), .B(u2_o_383_), .Y(u2__abc_52155_new_n23677_));
AND2X2 AND2X2_12173 ( .A(u2__abc_52155_new_n23678_), .B(u2__abc_52155_new_n23679_), .Y(u2__abc_52155_new_n23680_));
AND2X2 AND2X2_12174 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7213_), .Y(u2__abc_52155_new_n23682_));
AND2X2 AND2X2_12175 ( .A(u2__abc_52155_new_n23683_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23684_));
AND2X2 AND2X2_12176 ( .A(u2__abc_52155_new_n23681_), .B(u2__abc_52155_new_n23684_), .Y(u2__abc_52155_new_n23685_));
AND2X2 AND2X2_12177 ( .A(u2__abc_52155_new_n23686_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__385_));
AND2X2 AND2X2_12178 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_385_), .Y(u2__abc_52155_new_n23688_));
AND2X2 AND2X2_12179 ( .A(u2__abc_52155_new_n23677_), .B(u2_o_384_), .Y(u2__abc_52155_new_n23690_));
AND2X2 AND2X2_1218 ( .A(u2__abc_52155_new_n4501_), .B(u2_remHi_222_), .Y(u2__abc_52155_new_n4502_));
AND2X2 AND2X2_12180 ( .A(u2__abc_52155_new_n23691_), .B(u2__abc_52155_new_n23689_), .Y(u2__abc_52155_new_n23692_));
AND2X2 AND2X2_12181 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7223_), .Y(u2__abc_52155_new_n23694_));
AND2X2 AND2X2_12182 ( .A(u2__abc_52155_new_n23695_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23696_));
AND2X2 AND2X2_12183 ( .A(u2__abc_52155_new_n23693_), .B(u2__abc_52155_new_n23696_), .Y(u2__abc_52155_new_n23697_));
AND2X2 AND2X2_12184 ( .A(u2__abc_52155_new_n23698_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__386_));
AND2X2 AND2X2_12185 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_386_), .Y(u2__abc_52155_new_n23700_));
AND2X2 AND2X2_12186 ( .A(u2__abc_52155_new_n23690_), .B(u2_o_385_), .Y(u2__abc_52155_new_n23701_));
AND2X2 AND2X2_12187 ( .A(u2__abc_52155_new_n23702_), .B(u2__abc_52155_new_n23703_), .Y(u2__abc_52155_new_n23704_));
AND2X2 AND2X2_12188 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7204_), .Y(u2__abc_52155_new_n23706_));
AND2X2 AND2X2_12189 ( .A(u2__abc_52155_new_n23707_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23708_));
AND2X2 AND2X2_1219 ( .A(u2__abc_52155_new_n4504_), .B(sqrto_222_), .Y(u2__abc_52155_new_n4505_));
AND2X2 AND2X2_12190 ( .A(u2__abc_52155_new_n23705_), .B(u2__abc_52155_new_n23708_), .Y(u2__abc_52155_new_n23709_));
AND2X2 AND2X2_12191 ( .A(u2__abc_52155_new_n23710_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__387_));
AND2X2 AND2X2_12192 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_387_), .Y(u2__abc_52155_new_n23712_));
AND2X2 AND2X2_12193 ( .A(u2__abc_52155_new_n23701_), .B(u2_o_386_), .Y(u2__abc_52155_new_n23714_));
AND2X2 AND2X2_12194 ( .A(u2__abc_52155_new_n23715_), .B(u2__abc_52155_new_n23713_), .Y(u2__abc_52155_new_n23716_));
AND2X2 AND2X2_12195 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7200_), .Y(u2__abc_52155_new_n23718_));
AND2X2 AND2X2_12196 ( .A(u2__abc_52155_new_n23719_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23720_));
AND2X2 AND2X2_12197 ( .A(u2__abc_52155_new_n23717_), .B(u2__abc_52155_new_n23720_), .Y(u2__abc_52155_new_n23721_));
AND2X2 AND2X2_12198 ( .A(u2__abc_52155_new_n23722_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__388_));
AND2X2 AND2X2_12199 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_388_), .Y(u2__abc_52155_new_n23724_));
AND2X2 AND2X2_122 ( .A(_abc_73687_new_n966_), .B(_abc_73687_new_n965_), .Y(\o[157] ));
AND2X2 AND2X2_1220 ( .A(u2__abc_52155_new_n4503_), .B(u2__abc_52155_new_n4506_), .Y(u2__abc_52155_new_n4507_));
AND2X2 AND2X2_12200 ( .A(u2__abc_52155_new_n23714_), .B(u2_o_387_), .Y(u2__abc_52155_new_n23726_));
AND2X2 AND2X2_12201 ( .A(u2__abc_52155_new_n23727_), .B(u2__abc_52155_new_n23725_), .Y(u2__abc_52155_new_n23728_));
AND2X2 AND2X2_12202 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7182_), .Y(u2__abc_52155_new_n23730_));
AND2X2 AND2X2_12203 ( .A(u2__abc_52155_new_n23731_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23732_));
AND2X2 AND2X2_12204 ( .A(u2__abc_52155_new_n23729_), .B(u2__abc_52155_new_n23732_), .Y(u2__abc_52155_new_n23733_));
AND2X2 AND2X2_12205 ( .A(u2__abc_52155_new_n23734_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__389_));
AND2X2 AND2X2_12206 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_389_), .Y(u2__abc_52155_new_n23736_));
AND2X2 AND2X2_12207 ( .A(u2__abc_52155_new_n23726_), .B(u2_o_388_), .Y(u2__abc_52155_new_n23738_));
AND2X2 AND2X2_12208 ( .A(u2__abc_52155_new_n23739_), .B(u2__abc_52155_new_n23737_), .Y(u2__abc_52155_new_n23740_));
AND2X2 AND2X2_12209 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7189_), .Y(u2__abc_52155_new_n23742_));
AND2X2 AND2X2_1221 ( .A(u2__abc_52155_new_n4500_), .B(u2__abc_52155_new_n4507_), .Y(u2__abc_52155_new_n4508_));
AND2X2 AND2X2_12210 ( .A(u2__abc_52155_new_n23743_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23744_));
AND2X2 AND2X2_12211 ( .A(u2__abc_52155_new_n23741_), .B(u2__abc_52155_new_n23744_), .Y(u2__abc_52155_new_n23745_));
AND2X2 AND2X2_12212 ( .A(u2__abc_52155_new_n23746_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__390_));
AND2X2 AND2X2_12213 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_390_), .Y(u2__abc_52155_new_n23748_));
AND2X2 AND2X2_12214 ( .A(u2__abc_52155_new_n23738_), .B(u2_o_389_), .Y(u2__abc_52155_new_n23749_));
AND2X2 AND2X2_12215 ( .A(u2__abc_52155_new_n23750_), .B(u2__abc_52155_new_n23751_), .Y(u2__abc_52155_new_n23752_));
AND2X2 AND2X2_12216 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7387_), .Y(u2__abc_52155_new_n23754_));
AND2X2 AND2X2_12217 ( .A(u2__abc_52155_new_n23755_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23756_));
AND2X2 AND2X2_12218 ( .A(u2__abc_52155_new_n23753_), .B(u2__abc_52155_new_n23756_), .Y(u2__abc_52155_new_n23757_));
AND2X2 AND2X2_12219 ( .A(u2__abc_52155_new_n23758_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__391_));
AND2X2 AND2X2_1222 ( .A(u2__abc_52155_new_n4493_), .B(u2__abc_52155_new_n4508_), .Y(u2__abc_52155_new_n4509_));
AND2X2 AND2X2_12220 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_391_), .Y(u2__abc_52155_new_n23760_));
AND2X2 AND2X2_12221 ( .A(u2__abc_52155_new_n23749_), .B(u2_o_390_), .Y(u2__abc_52155_new_n23762_));
AND2X2 AND2X2_12222 ( .A(u2__abc_52155_new_n23763_), .B(u2__abc_52155_new_n23761_), .Y(u2__abc_52155_new_n23764_));
AND2X2 AND2X2_12223 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7397_), .Y(u2__abc_52155_new_n23766_));
AND2X2 AND2X2_12224 ( .A(u2__abc_52155_new_n23767_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23768_));
AND2X2 AND2X2_12225 ( .A(u2__abc_52155_new_n23765_), .B(u2__abc_52155_new_n23768_), .Y(u2__abc_52155_new_n23769_));
AND2X2 AND2X2_12226 ( .A(u2__abc_52155_new_n23770_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__392_));
AND2X2 AND2X2_12227 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_392_), .Y(u2__abc_52155_new_n23772_));
AND2X2 AND2X2_12228 ( .A(u2__abc_52155_new_n23762_), .B(u2_o_391_), .Y(u2__abc_52155_new_n23774_));
AND2X2 AND2X2_12229 ( .A(u2__abc_52155_new_n23775_), .B(u2__abc_52155_new_n23773_), .Y(u2__abc_52155_new_n23776_));
AND2X2 AND2X2_1223 ( .A(u2__abc_52155_new_n4510_), .B(u2_remHi_228_), .Y(u2__abc_52155_new_n4511_));
AND2X2 AND2X2_12230 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7372_), .Y(u2__abc_52155_new_n23778_));
AND2X2 AND2X2_12231 ( .A(u2__abc_52155_new_n23779_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23780_));
AND2X2 AND2X2_12232 ( .A(u2__abc_52155_new_n23777_), .B(u2__abc_52155_new_n23780_), .Y(u2__abc_52155_new_n23781_));
AND2X2 AND2X2_12233 ( .A(u2__abc_52155_new_n23782_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__393_));
AND2X2 AND2X2_12234 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_393_), .Y(u2__abc_52155_new_n23784_));
AND2X2 AND2X2_12235 ( .A(u2__abc_52155_new_n23774_), .B(u2_o_392_), .Y(u2__abc_52155_new_n23786_));
AND2X2 AND2X2_12236 ( .A(u2__abc_52155_new_n23787_), .B(u2__abc_52155_new_n23785_), .Y(u2__abc_52155_new_n23788_));
AND2X2 AND2X2_12237 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7382_), .Y(u2__abc_52155_new_n23790_));
AND2X2 AND2X2_12238 ( .A(u2__abc_52155_new_n23791_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23792_));
AND2X2 AND2X2_12239 ( .A(u2__abc_52155_new_n23789_), .B(u2__abc_52155_new_n23792_), .Y(u2__abc_52155_new_n23793_));
AND2X2 AND2X2_1224 ( .A(u2__abc_52155_new_n4513_), .B(u2_o_228_), .Y(u2__abc_52155_new_n4514_));
AND2X2 AND2X2_12240 ( .A(u2__abc_52155_new_n23794_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__394_));
AND2X2 AND2X2_12241 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_394_), .Y(u2__abc_52155_new_n23796_));
AND2X2 AND2X2_12242 ( .A(u2__abc_52155_new_n23786_), .B(u2_o_393_), .Y(u2__abc_52155_new_n23797_));
AND2X2 AND2X2_12243 ( .A(u2__abc_52155_new_n23798_), .B(u2__abc_52155_new_n23799_), .Y(u2__abc_52155_new_n23800_));
AND2X2 AND2X2_12244 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7425_), .Y(u2__abc_52155_new_n23802_));
AND2X2 AND2X2_12245 ( .A(u2__abc_52155_new_n23803_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23804_));
AND2X2 AND2X2_12246 ( .A(u2__abc_52155_new_n23801_), .B(u2__abc_52155_new_n23804_), .Y(u2__abc_52155_new_n23805_));
AND2X2 AND2X2_12247 ( .A(u2__abc_52155_new_n23806_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__395_));
AND2X2 AND2X2_12248 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_395_), .Y(u2__abc_52155_new_n23808_));
AND2X2 AND2X2_12249 ( .A(u2__abc_52155_new_n23797_), .B(u2_o_394_), .Y(u2__abc_52155_new_n23810_));
AND2X2 AND2X2_1225 ( .A(u2__abc_52155_new_n4512_), .B(u2__abc_52155_new_n4515_), .Y(u2__abc_52155_new_n4516_));
AND2X2 AND2X2_12250 ( .A(u2__abc_52155_new_n23811_), .B(u2__abc_52155_new_n23809_), .Y(u2__abc_52155_new_n23812_));
AND2X2 AND2X2_12251 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7421_), .Y(u2__abc_52155_new_n23814_));
AND2X2 AND2X2_12252 ( .A(u2__abc_52155_new_n23815_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23816_));
AND2X2 AND2X2_12253 ( .A(u2__abc_52155_new_n23813_), .B(u2__abc_52155_new_n23816_), .Y(u2__abc_52155_new_n23817_));
AND2X2 AND2X2_12254 ( .A(u2__abc_52155_new_n23818_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__396_));
AND2X2 AND2X2_12255 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_396_), .Y(u2__abc_52155_new_n23820_));
AND2X2 AND2X2_12256 ( .A(u2__abc_52155_new_n23810_), .B(u2_o_395_), .Y(u2__abc_52155_new_n23822_));
AND2X2 AND2X2_12257 ( .A(u2__abc_52155_new_n23823_), .B(u2__abc_52155_new_n23821_), .Y(u2__abc_52155_new_n23824_));
AND2X2 AND2X2_12258 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7403_), .Y(u2__abc_52155_new_n23826_));
AND2X2 AND2X2_12259 ( .A(u2__abc_52155_new_n23827_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23828_));
AND2X2 AND2X2_1226 ( .A(u2__abc_52155_new_n4517_), .B(u2_remHi_229_), .Y(u2__abc_52155_new_n4518_));
AND2X2 AND2X2_12260 ( .A(u2__abc_52155_new_n23825_), .B(u2__abc_52155_new_n23828_), .Y(u2__abc_52155_new_n23829_));
AND2X2 AND2X2_12261 ( .A(u2__abc_52155_new_n23830_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__397_));
AND2X2 AND2X2_12262 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_397_), .Y(u2__abc_52155_new_n23832_));
AND2X2 AND2X2_12263 ( .A(u2__abc_52155_new_n23822_), .B(u2_o_396_), .Y(u2__abc_52155_new_n23834_));
AND2X2 AND2X2_12264 ( .A(u2__abc_52155_new_n23835_), .B(u2__abc_52155_new_n23833_), .Y(u2__abc_52155_new_n23836_));
AND2X2 AND2X2_12265 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7410_), .Y(u2__abc_52155_new_n23838_));
AND2X2 AND2X2_12266 ( .A(u2__abc_52155_new_n23839_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23840_));
AND2X2 AND2X2_12267 ( .A(u2__abc_52155_new_n23837_), .B(u2__abc_52155_new_n23840_), .Y(u2__abc_52155_new_n23841_));
AND2X2 AND2X2_12268 ( .A(u2__abc_52155_new_n23842_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__398_));
AND2X2 AND2X2_12269 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_398_), .Y(u2__abc_52155_new_n23844_));
AND2X2 AND2X2_1227 ( .A(u2__abc_52155_new_n4520_), .B(u2_o_229_), .Y(u2__abc_52155_new_n4521_));
AND2X2 AND2X2_12270 ( .A(u2__abc_52155_new_n23834_), .B(u2_o_397_), .Y(u2__abc_52155_new_n23845_));
AND2X2 AND2X2_12271 ( .A(u2__abc_52155_new_n23846_), .B(u2__abc_52155_new_n23847_), .Y(u2__abc_52155_new_n23848_));
AND2X2 AND2X2_12272 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7308_), .Y(u2__abc_52155_new_n23850_));
AND2X2 AND2X2_12273 ( .A(u2__abc_52155_new_n23851_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23852_));
AND2X2 AND2X2_12274 ( .A(u2__abc_52155_new_n23849_), .B(u2__abc_52155_new_n23852_), .Y(u2__abc_52155_new_n23853_));
AND2X2 AND2X2_12275 ( .A(u2__abc_52155_new_n23854_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__399_));
AND2X2 AND2X2_12276 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_399_), .Y(u2__abc_52155_new_n23856_));
AND2X2 AND2X2_12277 ( .A(u2__abc_52155_new_n23845_), .B(u2_o_398_), .Y(u2__abc_52155_new_n23858_));
AND2X2 AND2X2_12278 ( .A(u2__abc_52155_new_n23859_), .B(u2__abc_52155_new_n23857_), .Y(u2__abc_52155_new_n23860_));
AND2X2 AND2X2_12279 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7318_), .Y(u2__abc_52155_new_n23862_));
AND2X2 AND2X2_1228 ( .A(u2__abc_52155_new_n4519_), .B(u2__abc_52155_new_n4522_), .Y(u2__abc_52155_new_n4523_));
AND2X2 AND2X2_12280 ( .A(u2__abc_52155_new_n23863_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23864_));
AND2X2 AND2X2_12281 ( .A(u2__abc_52155_new_n23861_), .B(u2__abc_52155_new_n23864_), .Y(u2__abc_52155_new_n23865_));
AND2X2 AND2X2_12282 ( .A(u2__abc_52155_new_n23866_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__400_));
AND2X2 AND2X2_12283 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_400_), .Y(u2__abc_52155_new_n23868_));
AND2X2 AND2X2_12284 ( .A(u2__abc_52155_new_n23858_), .B(u2_o_399_), .Y(u2__abc_52155_new_n23869_));
AND2X2 AND2X2_12285 ( .A(u2__abc_52155_new_n23870_), .B(u2__abc_52155_new_n23871_), .Y(u2__abc_52155_new_n23872_));
AND2X2 AND2X2_12286 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7323_), .Y(u2__abc_52155_new_n23874_));
AND2X2 AND2X2_12287 ( .A(u2__abc_52155_new_n23875_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23876_));
AND2X2 AND2X2_12288 ( .A(u2__abc_52155_new_n23873_), .B(u2__abc_52155_new_n23876_), .Y(u2__abc_52155_new_n23877_));
AND2X2 AND2X2_12289 ( .A(u2__abc_52155_new_n23878_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__401_));
AND2X2 AND2X2_1229 ( .A(u2__abc_52155_new_n4516_), .B(u2__abc_52155_new_n4523_), .Y(u2__abc_52155_new_n4524_));
AND2X2 AND2X2_12290 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_401_), .Y(u2__abc_52155_new_n23880_));
AND2X2 AND2X2_12291 ( .A(u2__abc_52155_new_n23869_), .B(u2_o_400_), .Y(u2__abc_52155_new_n23882_));
AND2X2 AND2X2_12292 ( .A(u2__abc_52155_new_n23883_), .B(u2__abc_52155_new_n23881_), .Y(u2__abc_52155_new_n23884_));
AND2X2 AND2X2_12293 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7333_), .Y(u2__abc_52155_new_n23886_));
AND2X2 AND2X2_12294 ( .A(u2__abc_52155_new_n23887_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23888_));
AND2X2 AND2X2_12295 ( .A(u2__abc_52155_new_n23885_), .B(u2__abc_52155_new_n23888_), .Y(u2__abc_52155_new_n23889_));
AND2X2 AND2X2_12296 ( .A(u2__abc_52155_new_n23890_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__402_));
AND2X2 AND2X2_12297 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_402_), .Y(u2__abc_52155_new_n23892_));
AND2X2 AND2X2_12298 ( .A(u2__abc_52155_new_n23882_), .B(u2_o_401_), .Y(u2__abc_52155_new_n23893_));
AND2X2 AND2X2_12299 ( .A(u2__abc_52155_new_n23894_), .B(u2__abc_52155_new_n23895_), .Y(u2__abc_52155_new_n23896_));
AND2X2 AND2X2_123 ( .A(_abc_73687_new_n969_), .B(_abc_73687_new_n968_), .Y(\o[158] ));
AND2X2 AND2X2_1230 ( .A(u2__abc_52155_new_n4525_), .B(u2_remHi_227_), .Y(u2__abc_52155_new_n4526_));
AND2X2 AND2X2_12300 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7361_), .Y(u2__abc_52155_new_n23898_));
AND2X2 AND2X2_12301 ( .A(u2__abc_52155_new_n23899_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23900_));
AND2X2 AND2X2_12302 ( .A(u2__abc_52155_new_n23897_), .B(u2__abc_52155_new_n23900_), .Y(u2__abc_52155_new_n23901_));
AND2X2 AND2X2_12303 ( .A(u2__abc_52155_new_n23902_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__403_));
AND2X2 AND2X2_12304 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_403_), .Y(u2__abc_52155_new_n23904_));
AND2X2 AND2X2_12305 ( .A(u2__abc_52155_new_n23893_), .B(u2_o_402_), .Y(u2__abc_52155_new_n23906_));
AND2X2 AND2X2_12306 ( .A(u2__abc_52155_new_n23907_), .B(u2__abc_52155_new_n23905_), .Y(u2__abc_52155_new_n23908_));
AND2X2 AND2X2_12307 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7357_), .Y(u2__abc_52155_new_n23910_));
AND2X2 AND2X2_12308 ( .A(u2__abc_52155_new_n23911_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23912_));
AND2X2 AND2X2_12309 ( .A(u2__abc_52155_new_n23909_), .B(u2__abc_52155_new_n23912_), .Y(u2__abc_52155_new_n23913_));
AND2X2 AND2X2_1231 ( .A(u2__abc_52155_new_n4528_), .B(u2_o_227_), .Y(u2__abc_52155_new_n4529_));
AND2X2 AND2X2_12310 ( .A(u2__abc_52155_new_n23914_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__404_));
AND2X2 AND2X2_12311 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_404_), .Y(u2__abc_52155_new_n23916_));
AND2X2 AND2X2_12312 ( .A(u2__abc_52155_new_n23906_), .B(u2_o_403_), .Y(u2__abc_52155_new_n23918_));
AND2X2 AND2X2_12313 ( .A(u2__abc_52155_new_n23919_), .B(u2__abc_52155_new_n23917_), .Y(u2__abc_52155_new_n23920_));
AND2X2 AND2X2_12314 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7339_), .Y(u2__abc_52155_new_n23922_));
AND2X2 AND2X2_12315 ( .A(u2__abc_52155_new_n23923_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23924_));
AND2X2 AND2X2_12316 ( .A(u2__abc_52155_new_n23921_), .B(u2__abc_52155_new_n23924_), .Y(u2__abc_52155_new_n23925_));
AND2X2 AND2X2_12317 ( .A(u2__abc_52155_new_n23926_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__405_));
AND2X2 AND2X2_12318 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_405_), .Y(u2__abc_52155_new_n23928_));
AND2X2 AND2X2_12319 ( .A(u2__abc_52155_new_n23918_), .B(u2_o_404_), .Y(u2__abc_52155_new_n23930_));
AND2X2 AND2X2_1232 ( .A(u2__abc_52155_new_n4527_), .B(u2__abc_52155_new_n4530_), .Y(u2__abc_52155_new_n4531_));
AND2X2 AND2X2_12320 ( .A(u2__abc_52155_new_n23931_), .B(u2__abc_52155_new_n23929_), .Y(u2__abc_52155_new_n23932_));
AND2X2 AND2X2_12321 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7346_), .Y(u2__abc_52155_new_n23934_));
AND2X2 AND2X2_12322 ( .A(u2__abc_52155_new_n23935_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23936_));
AND2X2 AND2X2_12323 ( .A(u2__abc_52155_new_n23933_), .B(u2__abc_52155_new_n23936_), .Y(u2__abc_52155_new_n23937_));
AND2X2 AND2X2_12324 ( .A(u2__abc_52155_new_n23938_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__406_));
AND2X2 AND2X2_12325 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_406_), .Y(u2__abc_52155_new_n23940_));
AND2X2 AND2X2_12326 ( .A(u2__abc_52155_new_n23930_), .B(u2_o_405_), .Y(u2__abc_52155_new_n23941_));
AND2X2 AND2X2_12327 ( .A(u2__abc_52155_new_n23942_), .B(u2__abc_52155_new_n23943_), .Y(u2__abc_52155_new_n23944_));
AND2X2 AND2X2_12328 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7267_), .Y(u2__abc_52155_new_n23946_));
AND2X2 AND2X2_12329 ( .A(u2__abc_52155_new_n23947_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23948_));
AND2X2 AND2X2_1233 ( .A(u2__abc_52155_new_n4532_), .B(u2_remHi_226_), .Y(u2__abc_52155_new_n4533_));
AND2X2 AND2X2_12330 ( .A(u2__abc_52155_new_n23945_), .B(u2__abc_52155_new_n23948_), .Y(u2__abc_52155_new_n23949_));
AND2X2 AND2X2_12331 ( .A(u2__abc_52155_new_n23950_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__407_));
AND2X2 AND2X2_12332 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_407_), .Y(u2__abc_52155_new_n23952_));
AND2X2 AND2X2_12333 ( .A(u2__abc_52155_new_n23941_), .B(u2_o_406_), .Y(u2__abc_52155_new_n23954_));
AND2X2 AND2X2_12334 ( .A(u2__abc_52155_new_n23955_), .B(u2__abc_52155_new_n23953_), .Y(u2__abc_52155_new_n23956_));
AND2X2 AND2X2_12335 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7263_), .Y(u2__abc_52155_new_n23958_));
AND2X2 AND2X2_12336 ( .A(u2__abc_52155_new_n23959_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23960_));
AND2X2 AND2X2_12337 ( .A(u2__abc_52155_new_n23957_), .B(u2__abc_52155_new_n23960_), .Y(u2__abc_52155_new_n23961_));
AND2X2 AND2X2_12338 ( .A(u2__abc_52155_new_n23962_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__408_));
AND2X2 AND2X2_12339 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_408_), .Y(u2__abc_52155_new_n23964_));
AND2X2 AND2X2_1234 ( .A(u2__abc_52155_new_n4535_), .B(u2_o_226_), .Y(u2__abc_52155_new_n4536_));
AND2X2 AND2X2_12340 ( .A(u2__abc_52155_new_n23954_), .B(u2_o_407_), .Y(u2__abc_52155_new_n23965_));
AND2X2 AND2X2_12341 ( .A(u2__abc_52155_new_n23966_), .B(u2__abc_52155_new_n23967_), .Y(u2__abc_52155_new_n23968_));
AND2X2 AND2X2_12342 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7245_), .Y(u2__abc_52155_new_n23970_));
AND2X2 AND2X2_12343 ( .A(u2__abc_52155_new_n23971_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23972_));
AND2X2 AND2X2_12344 ( .A(u2__abc_52155_new_n23969_), .B(u2__abc_52155_new_n23972_), .Y(u2__abc_52155_new_n23973_));
AND2X2 AND2X2_12345 ( .A(u2__abc_52155_new_n23974_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__409_));
AND2X2 AND2X2_12346 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_409_), .Y(u2__abc_52155_new_n23976_));
AND2X2 AND2X2_12347 ( .A(u2__abc_52155_new_n23965_), .B(u2_o_408_), .Y(u2__abc_52155_new_n23978_));
AND2X2 AND2X2_12348 ( .A(u2__abc_52155_new_n23979_), .B(u2__abc_52155_new_n23977_), .Y(u2__abc_52155_new_n23980_));
AND2X2 AND2X2_12349 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7255_), .Y(u2__abc_52155_new_n23982_));
AND2X2 AND2X2_1235 ( .A(u2__abc_52155_new_n4534_), .B(u2__abc_52155_new_n4537_), .Y(u2__abc_52155_new_n4538_));
AND2X2 AND2X2_12350 ( .A(u2__abc_52155_new_n23983_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23984_));
AND2X2 AND2X2_12351 ( .A(u2__abc_52155_new_n23981_), .B(u2__abc_52155_new_n23984_), .Y(u2__abc_52155_new_n23985_));
AND2X2 AND2X2_12352 ( .A(u2__abc_52155_new_n23986_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__410_));
AND2X2 AND2X2_12353 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_410_), .Y(u2__abc_52155_new_n23988_));
AND2X2 AND2X2_12354 ( .A(u2__abc_52155_new_n23978_), .B(u2_o_409_), .Y(u2__abc_52155_new_n23989_));
AND2X2 AND2X2_12355 ( .A(u2__abc_52155_new_n23990_), .B(u2__abc_52155_new_n23991_), .Y(u2__abc_52155_new_n23992_));
AND2X2 AND2X2_12356 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7298_), .Y(u2__abc_52155_new_n23994_));
AND2X2 AND2X2_12357 ( .A(u2__abc_52155_new_n23995_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n23996_));
AND2X2 AND2X2_12358 ( .A(u2__abc_52155_new_n23993_), .B(u2__abc_52155_new_n23996_), .Y(u2__abc_52155_new_n23997_));
AND2X2 AND2X2_12359 ( .A(u2__abc_52155_new_n23998_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__411_));
AND2X2 AND2X2_1236 ( .A(u2__abc_52155_new_n4531_), .B(u2__abc_52155_new_n4538_), .Y(u2__abc_52155_new_n4539_));
AND2X2 AND2X2_12360 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_411_), .Y(u2__abc_52155_new_n24000_));
AND2X2 AND2X2_12361 ( .A(u2__abc_52155_new_n23989_), .B(u2_o_410_), .Y(u2__abc_52155_new_n24002_));
AND2X2 AND2X2_12362 ( .A(u2__abc_52155_new_n24003_), .B(u2__abc_52155_new_n24001_), .Y(u2__abc_52155_new_n24004_));
AND2X2 AND2X2_12363 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7294_), .Y(u2__abc_52155_new_n24006_));
AND2X2 AND2X2_12364 ( .A(u2__abc_52155_new_n24007_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24008_));
AND2X2 AND2X2_12365 ( .A(u2__abc_52155_new_n24005_), .B(u2__abc_52155_new_n24008_), .Y(u2__abc_52155_new_n24009_));
AND2X2 AND2X2_12366 ( .A(u2__abc_52155_new_n24010_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__412_));
AND2X2 AND2X2_12367 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_412_), .Y(u2__abc_52155_new_n24012_));
AND2X2 AND2X2_12368 ( .A(u2__abc_52155_new_n24002_), .B(u2_o_411_), .Y(u2__abc_52155_new_n24013_));
AND2X2 AND2X2_12369 ( .A(u2__abc_52155_new_n24014_), .B(u2__abc_52155_new_n24015_), .Y(u2__abc_52155_new_n24016_));
AND2X2 AND2X2_1237 ( .A(u2__abc_52155_new_n4524_), .B(u2__abc_52155_new_n4539_), .Y(u2__abc_52155_new_n4540_));
AND2X2 AND2X2_12370 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7276_), .Y(u2__abc_52155_new_n24018_));
AND2X2 AND2X2_12371 ( .A(u2__abc_52155_new_n24019_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24020_));
AND2X2 AND2X2_12372 ( .A(u2__abc_52155_new_n24017_), .B(u2__abc_52155_new_n24020_), .Y(u2__abc_52155_new_n24021_));
AND2X2 AND2X2_12373 ( .A(u2__abc_52155_new_n24022_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__413_));
AND2X2 AND2X2_12374 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_413_), .Y(u2__abc_52155_new_n24024_));
AND2X2 AND2X2_12375 ( .A(u2__abc_52155_new_n24013_), .B(u2_o_412_), .Y(u2__abc_52155_new_n24026_));
AND2X2 AND2X2_12376 ( .A(u2__abc_52155_new_n24027_), .B(u2__abc_52155_new_n24025_), .Y(u2__abc_52155_new_n24028_));
AND2X2 AND2X2_12377 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7283_), .Y(u2__abc_52155_new_n24030_));
AND2X2 AND2X2_12378 ( .A(u2__abc_52155_new_n24031_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24032_));
AND2X2 AND2X2_12379 ( .A(u2__abc_52155_new_n24029_), .B(u2__abc_52155_new_n24032_), .Y(u2__abc_52155_new_n24033_));
AND2X2 AND2X2_1238 ( .A(u2__abc_52155_new_n4509_), .B(u2__abc_52155_new_n4540_), .Y(u2__abc_52155_new_n4541_));
AND2X2 AND2X2_12380 ( .A(u2__abc_52155_new_n24034_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__414_));
AND2X2 AND2X2_12381 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_414_), .Y(u2__abc_52155_new_n24036_));
AND2X2 AND2X2_12382 ( .A(u2__abc_52155_new_n24026_), .B(u2_o_413_), .Y(u2__abc_52155_new_n24037_));
AND2X2 AND2X2_12383 ( .A(u2__abc_52155_new_n24038_), .B(u2__abc_52155_new_n24039_), .Y(u2__abc_52155_new_n24040_));
AND2X2 AND2X2_12384 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7170_), .Y(u2__abc_52155_new_n24042_));
AND2X2 AND2X2_12385 ( .A(u2__abc_52155_new_n24043_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24044_));
AND2X2 AND2X2_12386 ( .A(u2__abc_52155_new_n24041_), .B(u2__abc_52155_new_n24044_), .Y(u2__abc_52155_new_n24045_));
AND2X2 AND2X2_12387 ( .A(u2__abc_52155_new_n24046_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__415_));
AND2X2 AND2X2_12388 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_415_), .Y(u2__abc_52155_new_n24048_));
AND2X2 AND2X2_12389 ( .A(u2__abc_52155_new_n24037_), .B(u2_o_414_), .Y(u2__abc_52155_new_n24050_));
AND2X2 AND2X2_1239 ( .A(u2__abc_52155_new_n4478_), .B(u2__abc_52155_new_n4541_), .Y(u2__abc_52155_new_n4542_));
AND2X2 AND2X2_12390 ( .A(u2__abc_52155_new_n24051_), .B(u2__abc_52155_new_n24049_), .Y(u2__abc_52155_new_n24052_));
AND2X2 AND2X2_12391 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7166_), .Y(u2__abc_52155_new_n24054_));
AND2X2 AND2X2_12392 ( .A(u2__abc_52155_new_n24055_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24056_));
AND2X2 AND2X2_12393 ( .A(u2__abc_52155_new_n24053_), .B(u2__abc_52155_new_n24056_), .Y(u2__abc_52155_new_n24057_));
AND2X2 AND2X2_12394 ( .A(u2__abc_52155_new_n24058_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__416_));
AND2X2 AND2X2_12395 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_416_), .Y(u2__abc_52155_new_n24060_));
AND2X2 AND2X2_12396 ( .A(u2__abc_52155_new_n24050_), .B(u2_o_415_), .Y(u2__abc_52155_new_n24061_));
AND2X2 AND2X2_12397 ( .A(u2__abc_52155_new_n24062_), .B(u2__abc_52155_new_n24063_), .Y(u2__abc_52155_new_n24064_));
AND2X2 AND2X2_12398 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7148_), .Y(u2__abc_52155_new_n24066_));
AND2X2 AND2X2_12399 ( .A(u2__abc_52155_new_n24067_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24068_));
AND2X2 AND2X2_124 ( .A(_abc_73687_new_n972_), .B(_abc_73687_new_n971_), .Y(\o[159] ));
AND2X2 AND2X2_1240 ( .A(u2__abc_52155_new_n4415_), .B(u2__abc_52155_new_n4542_), .Y(u2__abc_52155_new_n4543_));
AND2X2 AND2X2_12400 ( .A(u2__abc_52155_new_n24065_), .B(u2__abc_52155_new_n24068_), .Y(u2__abc_52155_new_n24069_));
AND2X2 AND2X2_12401 ( .A(u2__abc_52155_new_n24070_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__417_));
AND2X2 AND2X2_12402 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_417_), .Y(u2__abc_52155_new_n24072_));
AND2X2 AND2X2_12403 ( .A(u2__abc_52155_new_n24061_), .B(u2_o_416_), .Y(u2__abc_52155_new_n24074_));
AND2X2 AND2X2_12404 ( .A(u2__abc_52155_new_n24075_), .B(u2__abc_52155_new_n24073_), .Y(u2__abc_52155_new_n24076_));
AND2X2 AND2X2_12405 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7158_), .Y(u2__abc_52155_new_n24078_));
AND2X2 AND2X2_12406 ( .A(u2__abc_52155_new_n24079_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24080_));
AND2X2 AND2X2_12407 ( .A(u2__abc_52155_new_n24077_), .B(u2__abc_52155_new_n24080_), .Y(u2__abc_52155_new_n24081_));
AND2X2 AND2X2_12408 ( .A(u2__abc_52155_new_n24082_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__418_));
AND2X2 AND2X2_12409 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_418_), .Y(u2__abc_52155_new_n24084_));
AND2X2 AND2X2_1241 ( .A(u2__abc_52155_new_n4544_), .B(u2_remHi_216_), .Y(u2__abc_52155_new_n4545_));
AND2X2 AND2X2_12410 ( .A(u2__abc_52155_new_n24074_), .B(u2_o_417_), .Y(u2__abc_52155_new_n24085_));
AND2X2 AND2X2_12411 ( .A(u2__abc_52155_new_n24086_), .B(u2__abc_52155_new_n24087_), .Y(u2__abc_52155_new_n24088_));
AND2X2 AND2X2_12412 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7139_), .Y(u2__abc_52155_new_n24090_));
AND2X2 AND2X2_12413 ( .A(u2__abc_52155_new_n24091_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24092_));
AND2X2 AND2X2_12414 ( .A(u2__abc_52155_new_n24089_), .B(u2__abc_52155_new_n24092_), .Y(u2__abc_52155_new_n24093_));
AND2X2 AND2X2_12415 ( .A(u2__abc_52155_new_n24094_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__419_));
AND2X2 AND2X2_12416 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_419_), .Y(u2__abc_52155_new_n24096_));
AND2X2 AND2X2_12417 ( .A(u2__abc_52155_new_n24085_), .B(u2_o_418_), .Y(u2__abc_52155_new_n24098_));
AND2X2 AND2X2_12418 ( .A(u2__abc_52155_new_n24099_), .B(u2__abc_52155_new_n24097_), .Y(u2__abc_52155_new_n24100_));
AND2X2 AND2X2_12419 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7135_), .Y(u2__abc_52155_new_n24102_));
AND2X2 AND2X2_1242 ( .A(u2__abc_52155_new_n4547_), .B(sqrto_216_), .Y(u2__abc_52155_new_n4548_));
AND2X2 AND2X2_12420 ( .A(u2__abc_52155_new_n24103_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24104_));
AND2X2 AND2X2_12421 ( .A(u2__abc_52155_new_n24101_), .B(u2__abc_52155_new_n24104_), .Y(u2__abc_52155_new_n24105_));
AND2X2 AND2X2_12422 ( .A(u2__abc_52155_new_n24106_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__420_));
AND2X2 AND2X2_12423 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_420_), .Y(u2__abc_52155_new_n24108_));
AND2X2 AND2X2_12424 ( .A(u2__abc_52155_new_n24098_), .B(u2_o_419_), .Y(u2__abc_52155_new_n24110_));
AND2X2 AND2X2_12425 ( .A(u2__abc_52155_new_n24111_), .B(u2__abc_52155_new_n24109_), .Y(u2__abc_52155_new_n24112_));
AND2X2 AND2X2_12426 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7117_), .Y(u2__abc_52155_new_n24114_));
AND2X2 AND2X2_12427 ( .A(u2__abc_52155_new_n24115_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24116_));
AND2X2 AND2X2_12428 ( .A(u2__abc_52155_new_n24113_), .B(u2__abc_52155_new_n24116_), .Y(u2__abc_52155_new_n24117_));
AND2X2 AND2X2_12429 ( .A(u2__abc_52155_new_n24118_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__421_));
AND2X2 AND2X2_1243 ( .A(u2__abc_52155_new_n4546_), .B(u2__abc_52155_new_n4549_), .Y(u2__abc_52155_new_n4550_));
AND2X2 AND2X2_12430 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_421_), .Y(u2__abc_52155_new_n24120_));
AND2X2 AND2X2_12431 ( .A(u2__abc_52155_new_n24110_), .B(u2_o_420_), .Y(u2__abc_52155_new_n24122_));
AND2X2 AND2X2_12432 ( .A(u2__abc_52155_new_n24123_), .B(u2__abc_52155_new_n24121_), .Y(u2__abc_52155_new_n24124_));
AND2X2 AND2X2_12433 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7124_), .Y(u2__abc_52155_new_n24126_));
AND2X2 AND2X2_12434 ( .A(u2__abc_52155_new_n24127_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24128_));
AND2X2 AND2X2_12435 ( .A(u2__abc_52155_new_n24125_), .B(u2__abc_52155_new_n24128_), .Y(u2__abc_52155_new_n24129_));
AND2X2 AND2X2_12436 ( .A(u2__abc_52155_new_n24130_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__422_));
AND2X2 AND2X2_12437 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_422_), .Y(u2__abc_52155_new_n24132_));
AND2X2 AND2X2_12438 ( .A(u2__abc_52155_new_n24122_), .B(u2_o_421_), .Y(u2__abc_52155_new_n24133_));
AND2X2 AND2X2_12439 ( .A(u2__abc_52155_new_n24134_), .B(u2__abc_52155_new_n24135_), .Y(u2__abc_52155_new_n24136_));
AND2X2 AND2X2_1244 ( .A(u2__abc_52155_new_n4551_), .B(u2_remHi_217_), .Y(u2__abc_52155_new_n4552_));
AND2X2 AND2X2_12440 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7069_), .Y(u2__abc_52155_new_n24138_));
AND2X2 AND2X2_12441 ( .A(u2__abc_52155_new_n24139_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24140_));
AND2X2 AND2X2_12442 ( .A(u2__abc_52155_new_n24137_), .B(u2__abc_52155_new_n24140_), .Y(u2__abc_52155_new_n24141_));
AND2X2 AND2X2_12443 ( .A(u2__abc_52155_new_n24142_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__423_));
AND2X2 AND2X2_12444 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_423_), .Y(u2__abc_52155_new_n24144_));
AND2X2 AND2X2_12445 ( .A(u2__abc_52155_new_n24133_), .B(u2_o_422_), .Y(u2__abc_52155_new_n24146_));
AND2X2 AND2X2_12446 ( .A(u2__abc_52155_new_n24147_), .B(u2__abc_52155_new_n24145_), .Y(u2__abc_52155_new_n24148_));
AND2X2 AND2X2_12447 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7079_), .Y(u2__abc_52155_new_n24150_));
AND2X2 AND2X2_12448 ( .A(u2__abc_52155_new_n24151_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24152_));
AND2X2 AND2X2_12449 ( .A(u2__abc_52155_new_n24149_), .B(u2__abc_52155_new_n24152_), .Y(u2__abc_52155_new_n24153_));
AND2X2 AND2X2_1245 ( .A(u2__abc_52155_new_n4554_), .B(sqrto_217_), .Y(u2__abc_52155_new_n4555_));
AND2X2 AND2X2_12450 ( .A(u2__abc_52155_new_n24154_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__424_));
AND2X2 AND2X2_12451 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_424_), .Y(u2__abc_52155_new_n24156_));
AND2X2 AND2X2_12452 ( .A(u2__abc_52155_new_n24146_), .B(u2_o_423_), .Y(u2__abc_52155_new_n24157_));
AND2X2 AND2X2_12453 ( .A(u2__abc_52155_new_n24158_), .B(u2__abc_52155_new_n24159_), .Y(u2__abc_52155_new_n24160_));
AND2X2 AND2X2_12454 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7054_), .Y(u2__abc_52155_new_n24162_));
AND2X2 AND2X2_12455 ( .A(u2__abc_52155_new_n24163_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24164_));
AND2X2 AND2X2_12456 ( .A(u2__abc_52155_new_n24161_), .B(u2__abc_52155_new_n24164_), .Y(u2__abc_52155_new_n24165_));
AND2X2 AND2X2_12457 ( .A(u2__abc_52155_new_n24166_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__425_));
AND2X2 AND2X2_12458 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_425_), .Y(u2__abc_52155_new_n24168_));
AND2X2 AND2X2_12459 ( .A(u2__abc_52155_new_n24157_), .B(u2_o_424_), .Y(u2__abc_52155_new_n24170_));
AND2X2 AND2X2_1246 ( .A(u2__abc_52155_new_n4553_), .B(u2__abc_52155_new_n4556_), .Y(u2__abc_52155_new_n4557_));
AND2X2 AND2X2_12460 ( .A(u2__abc_52155_new_n24171_), .B(u2__abc_52155_new_n24169_), .Y(u2__abc_52155_new_n24172_));
AND2X2 AND2X2_12461 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7064_), .Y(u2__abc_52155_new_n24174_));
AND2X2 AND2X2_12462 ( .A(u2__abc_52155_new_n24175_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24176_));
AND2X2 AND2X2_12463 ( .A(u2__abc_52155_new_n24173_), .B(u2__abc_52155_new_n24176_), .Y(u2__abc_52155_new_n24177_));
AND2X2 AND2X2_12464 ( .A(u2__abc_52155_new_n24178_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__426_));
AND2X2 AND2X2_12465 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_426_), .Y(u2__abc_52155_new_n24180_));
AND2X2 AND2X2_12466 ( .A(u2__abc_52155_new_n24170_), .B(u2_o_425_), .Y(u2__abc_52155_new_n24181_));
AND2X2 AND2X2_12467 ( .A(u2__abc_52155_new_n24182_), .B(u2__abc_52155_new_n24183_), .Y(u2__abc_52155_new_n24184_));
AND2X2 AND2X2_12468 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7107_), .Y(u2__abc_52155_new_n24186_));
AND2X2 AND2X2_12469 ( .A(u2__abc_52155_new_n24187_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24188_));
AND2X2 AND2X2_1247 ( .A(u2__abc_52155_new_n4550_), .B(u2__abc_52155_new_n4557_), .Y(u2__abc_52155_new_n4558_));
AND2X2 AND2X2_12470 ( .A(u2__abc_52155_new_n24185_), .B(u2__abc_52155_new_n24188_), .Y(u2__abc_52155_new_n24189_));
AND2X2 AND2X2_12471 ( .A(u2__abc_52155_new_n24190_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__427_));
AND2X2 AND2X2_12472 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_427_), .Y(u2__abc_52155_new_n24192_));
AND2X2 AND2X2_12473 ( .A(u2__abc_52155_new_n24181_), .B(u2_o_426_), .Y(u2__abc_52155_new_n24194_));
AND2X2 AND2X2_12474 ( .A(u2__abc_52155_new_n24195_), .B(u2__abc_52155_new_n24193_), .Y(u2__abc_52155_new_n24196_));
AND2X2 AND2X2_12475 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7103_), .Y(u2__abc_52155_new_n24198_));
AND2X2 AND2X2_12476 ( .A(u2__abc_52155_new_n24199_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24200_));
AND2X2 AND2X2_12477 ( .A(u2__abc_52155_new_n24197_), .B(u2__abc_52155_new_n24200_), .Y(u2__abc_52155_new_n24201_));
AND2X2 AND2X2_12478 ( .A(u2__abc_52155_new_n24202_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__428_));
AND2X2 AND2X2_12479 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_428_), .Y(u2__abc_52155_new_n24204_));
AND2X2 AND2X2_1248 ( .A(u2__abc_52155_new_n4559_), .B(u2_remHi_214_), .Y(u2__abc_52155_new_n4560_));
AND2X2 AND2X2_12480 ( .A(u2__abc_52155_new_n24194_), .B(u2_o_427_), .Y(u2__abc_52155_new_n24205_));
AND2X2 AND2X2_12481 ( .A(u2__abc_52155_new_n24206_), .B(u2__abc_52155_new_n24207_), .Y(u2__abc_52155_new_n24208_));
AND2X2 AND2X2_12482 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7085_), .Y(u2__abc_52155_new_n24210_));
AND2X2 AND2X2_12483 ( .A(u2__abc_52155_new_n24211_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24212_));
AND2X2 AND2X2_12484 ( .A(u2__abc_52155_new_n24209_), .B(u2__abc_52155_new_n24212_), .Y(u2__abc_52155_new_n24213_));
AND2X2 AND2X2_12485 ( .A(u2__abc_52155_new_n24214_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__429_));
AND2X2 AND2X2_12486 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_429_), .Y(u2__abc_52155_new_n24216_));
AND2X2 AND2X2_12487 ( .A(u2__abc_52155_new_n24205_), .B(u2_o_428_), .Y(u2__abc_52155_new_n24218_));
AND2X2 AND2X2_12488 ( .A(u2__abc_52155_new_n24219_), .B(u2__abc_52155_new_n24217_), .Y(u2__abc_52155_new_n24220_));
AND2X2 AND2X2_12489 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7092_), .Y(u2__abc_52155_new_n24222_));
AND2X2 AND2X2_1249 ( .A(u2__abc_52155_new_n4562_), .B(sqrto_214_), .Y(u2__abc_52155_new_n4563_));
AND2X2 AND2X2_12490 ( .A(u2__abc_52155_new_n24223_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24224_));
AND2X2 AND2X2_12491 ( .A(u2__abc_52155_new_n24221_), .B(u2__abc_52155_new_n24224_), .Y(u2__abc_52155_new_n24225_));
AND2X2 AND2X2_12492 ( .A(u2__abc_52155_new_n24226_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__430_));
AND2X2 AND2X2_12493 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_430_), .Y(u2__abc_52155_new_n24228_));
AND2X2 AND2X2_12494 ( .A(u2__abc_52155_new_n24218_), .B(u2_o_429_), .Y(u2__abc_52155_new_n24229_));
AND2X2 AND2X2_12495 ( .A(u2__abc_52155_new_n24230_), .B(u2__abc_52155_new_n24231_), .Y(u2__abc_52155_new_n24232_));
AND2X2 AND2X2_12496 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7021_), .Y(u2__abc_52155_new_n24234_));
AND2X2 AND2X2_12497 ( .A(u2__abc_52155_new_n24235_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24236_));
AND2X2 AND2X2_12498 ( .A(u2__abc_52155_new_n24233_), .B(u2__abc_52155_new_n24236_), .Y(u2__abc_52155_new_n24237_));
AND2X2 AND2X2_12499 ( .A(u2__abc_52155_new_n24238_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__431_));
AND2X2 AND2X2_125 ( .A(_abc_73687_new_n975_), .B(_abc_73687_new_n974_), .Y(\o[160] ));
AND2X2 AND2X2_1250 ( .A(u2__abc_52155_new_n4561_), .B(u2__abc_52155_new_n4564_), .Y(u2__abc_52155_new_n4565_));
AND2X2 AND2X2_12500 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_431_), .Y(u2__abc_52155_new_n24240_));
AND2X2 AND2X2_12501 ( .A(u2__abc_52155_new_n24229_), .B(u2_o_430_), .Y(u2__abc_52155_new_n24242_));
AND2X2 AND2X2_12502 ( .A(u2__abc_52155_new_n24243_), .B(u2__abc_52155_new_n24241_), .Y(u2__abc_52155_new_n24244_));
AND2X2 AND2X2_12503 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7031_), .Y(u2__abc_52155_new_n24246_));
AND2X2 AND2X2_12504 ( .A(u2__abc_52155_new_n24247_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24248_));
AND2X2 AND2X2_12505 ( .A(u2__abc_52155_new_n24245_), .B(u2__abc_52155_new_n24248_), .Y(u2__abc_52155_new_n24249_));
AND2X2 AND2X2_12506 ( .A(u2__abc_52155_new_n24250_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__432_));
AND2X2 AND2X2_12507 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_432_), .Y(u2__abc_52155_new_n24252_));
AND2X2 AND2X2_12508 ( .A(u2__abc_52155_new_n24242_), .B(u2_o_431_), .Y(u2__abc_52155_new_n24253_));
AND2X2 AND2X2_12509 ( .A(u2__abc_52155_new_n24254_), .B(u2__abc_52155_new_n24255_), .Y(u2__abc_52155_new_n24256_));
AND2X2 AND2X2_1251 ( .A(u2__abc_52155_new_n4566_), .B(u2_remHi_215_), .Y(u2__abc_52155_new_n4567_));
AND2X2 AND2X2_12510 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7036_), .Y(u2__abc_52155_new_n24258_));
AND2X2 AND2X2_12511 ( .A(u2__abc_52155_new_n24259_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24260_));
AND2X2 AND2X2_12512 ( .A(u2__abc_52155_new_n24257_), .B(u2__abc_52155_new_n24260_), .Y(u2__abc_52155_new_n24261_));
AND2X2 AND2X2_12513 ( .A(u2__abc_52155_new_n24262_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__433_));
AND2X2 AND2X2_12514 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_433_), .Y(u2__abc_52155_new_n24264_));
AND2X2 AND2X2_12515 ( .A(u2__abc_52155_new_n24253_), .B(u2_o_432_), .Y(u2__abc_52155_new_n24266_));
AND2X2 AND2X2_12516 ( .A(u2__abc_52155_new_n24267_), .B(u2__abc_52155_new_n24265_), .Y(u2__abc_52155_new_n24268_));
AND2X2 AND2X2_12517 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7046_), .Y(u2__abc_52155_new_n24270_));
AND2X2 AND2X2_12518 ( .A(u2__abc_52155_new_n24271_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24272_));
AND2X2 AND2X2_12519 ( .A(u2__abc_52155_new_n24269_), .B(u2__abc_52155_new_n24272_), .Y(u2__abc_52155_new_n24273_));
AND2X2 AND2X2_1252 ( .A(u2__abc_52155_new_n4569_), .B(sqrto_215_), .Y(u2__abc_52155_new_n4570_));
AND2X2 AND2X2_12520 ( .A(u2__abc_52155_new_n24274_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__434_));
AND2X2 AND2X2_12521 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_434_), .Y(u2__abc_52155_new_n24276_));
AND2X2 AND2X2_12522 ( .A(u2__abc_52155_new_n24266_), .B(u2_o_433_), .Y(u2__abc_52155_new_n24277_));
AND2X2 AND2X2_12523 ( .A(u2__abc_52155_new_n24278_), .B(u2__abc_52155_new_n24279_), .Y(u2__abc_52155_new_n24280_));
AND2X2 AND2X2_12524 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7012_), .Y(u2__abc_52155_new_n24282_));
AND2X2 AND2X2_12525 ( .A(u2__abc_52155_new_n24283_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24284_));
AND2X2 AND2X2_12526 ( .A(u2__abc_52155_new_n24281_), .B(u2__abc_52155_new_n24284_), .Y(u2__abc_52155_new_n24285_));
AND2X2 AND2X2_12527 ( .A(u2__abc_52155_new_n24286_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__435_));
AND2X2 AND2X2_12528 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_435_), .Y(u2__abc_52155_new_n24288_));
AND2X2 AND2X2_12529 ( .A(u2__abc_52155_new_n24277_), .B(u2_o_434_), .Y(u2__abc_52155_new_n24290_));
AND2X2 AND2X2_1253 ( .A(u2__abc_52155_new_n4568_), .B(u2__abc_52155_new_n4571_), .Y(u2__abc_52155_new_n4572_));
AND2X2 AND2X2_12530 ( .A(u2__abc_52155_new_n24291_), .B(u2__abc_52155_new_n24289_), .Y(u2__abc_52155_new_n24292_));
AND2X2 AND2X2_12531 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7008_), .Y(u2__abc_52155_new_n24294_));
AND2X2 AND2X2_12532 ( .A(u2__abc_52155_new_n24295_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24296_));
AND2X2 AND2X2_12533 ( .A(u2__abc_52155_new_n24293_), .B(u2__abc_52155_new_n24296_), .Y(u2__abc_52155_new_n24297_));
AND2X2 AND2X2_12534 ( .A(u2__abc_52155_new_n24298_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__436_));
AND2X2 AND2X2_12535 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_436_), .Y(u2__abc_52155_new_n24300_));
AND2X2 AND2X2_12536 ( .A(u2__abc_52155_new_n24290_), .B(u2_o_435_), .Y(u2__abc_52155_new_n24301_));
AND2X2 AND2X2_12537 ( .A(u2__abc_52155_new_n24302_), .B(u2__abc_52155_new_n24303_), .Y(u2__abc_52155_new_n24304_));
AND2X2 AND2X2_12538 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6990_), .Y(u2__abc_52155_new_n24306_));
AND2X2 AND2X2_12539 ( .A(u2__abc_52155_new_n24307_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24308_));
AND2X2 AND2X2_1254 ( .A(u2__abc_52155_new_n4565_), .B(u2__abc_52155_new_n4572_), .Y(u2__abc_52155_new_n4573_));
AND2X2 AND2X2_12540 ( .A(u2__abc_52155_new_n24305_), .B(u2__abc_52155_new_n24308_), .Y(u2__abc_52155_new_n24309_));
AND2X2 AND2X2_12541 ( .A(u2__abc_52155_new_n24310_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__437_));
AND2X2 AND2X2_12542 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_437_), .Y(u2__abc_52155_new_n24312_));
AND2X2 AND2X2_12543 ( .A(u2__abc_52155_new_n24301_), .B(u2_o_436_), .Y(u2__abc_52155_new_n24314_));
AND2X2 AND2X2_12544 ( .A(u2__abc_52155_new_n24315_), .B(u2__abc_52155_new_n24313_), .Y(u2__abc_52155_new_n24316_));
AND2X2 AND2X2_12545 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6997_), .Y(u2__abc_52155_new_n24318_));
AND2X2 AND2X2_12546 ( .A(u2__abc_52155_new_n24319_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24320_));
AND2X2 AND2X2_12547 ( .A(u2__abc_52155_new_n24317_), .B(u2__abc_52155_new_n24320_), .Y(u2__abc_52155_new_n24321_));
AND2X2 AND2X2_12548 ( .A(u2__abc_52155_new_n24322_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__438_));
AND2X2 AND2X2_12549 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_438_), .Y(u2__abc_52155_new_n24324_));
AND2X2 AND2X2_1255 ( .A(u2__abc_52155_new_n4558_), .B(u2__abc_52155_new_n4573_), .Y(u2__abc_52155_new_n4574_));
AND2X2 AND2X2_12550 ( .A(u2__abc_52155_new_n24314_), .B(u2_o_437_), .Y(u2__abc_52155_new_n24325_));
AND2X2 AND2X2_12551 ( .A(u2__abc_52155_new_n24326_), .B(u2__abc_52155_new_n24327_), .Y(u2__abc_52155_new_n24328_));
AND2X2 AND2X2_12552 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6958_), .Y(u2__abc_52155_new_n24330_));
AND2X2 AND2X2_12553 ( .A(u2__abc_52155_new_n24331_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24332_));
AND2X2 AND2X2_12554 ( .A(u2__abc_52155_new_n24329_), .B(u2__abc_52155_new_n24332_), .Y(u2__abc_52155_new_n24333_));
AND2X2 AND2X2_12555 ( .A(u2__abc_52155_new_n24334_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__439_));
AND2X2 AND2X2_12556 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_439_), .Y(u2__abc_52155_new_n24336_));
AND2X2 AND2X2_12557 ( .A(u2__abc_52155_new_n24325_), .B(u2_o_438_), .Y(u2__abc_52155_new_n24338_));
AND2X2 AND2X2_12558 ( .A(u2__abc_52155_new_n24339_), .B(u2__abc_52155_new_n24337_), .Y(u2__abc_52155_new_n24340_));
AND2X2 AND2X2_12559 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6968_), .Y(u2__abc_52155_new_n24342_));
AND2X2 AND2X2_1256 ( .A(u2__abc_52155_new_n4575_), .B(u2_remHi_220_), .Y(u2__abc_52155_new_n4576_));
AND2X2 AND2X2_12560 ( .A(u2__abc_52155_new_n24343_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24344_));
AND2X2 AND2X2_12561 ( .A(u2__abc_52155_new_n24341_), .B(u2__abc_52155_new_n24344_), .Y(u2__abc_52155_new_n24345_));
AND2X2 AND2X2_12562 ( .A(u2__abc_52155_new_n24346_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__440_));
AND2X2 AND2X2_12563 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_440_), .Y(u2__abc_52155_new_n24348_));
AND2X2 AND2X2_12564 ( .A(u2__abc_52155_new_n24338_), .B(u2_o_439_), .Y(u2__abc_52155_new_n24349_));
AND2X2 AND2X2_12565 ( .A(u2__abc_52155_new_n24350_), .B(u2__abc_52155_new_n24351_), .Y(u2__abc_52155_new_n24352_));
AND2X2 AND2X2_12566 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6973_), .Y(u2__abc_52155_new_n24354_));
AND2X2 AND2X2_12567 ( .A(u2__abc_52155_new_n24355_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24356_));
AND2X2 AND2X2_12568 ( .A(u2__abc_52155_new_n24353_), .B(u2__abc_52155_new_n24356_), .Y(u2__abc_52155_new_n24357_));
AND2X2 AND2X2_12569 ( .A(u2__abc_52155_new_n24358_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__441_));
AND2X2 AND2X2_1257 ( .A(u2__abc_52155_new_n4578_), .B(sqrto_220_), .Y(u2__abc_52155_new_n4579_));
AND2X2 AND2X2_12570 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_441_), .Y(u2__abc_52155_new_n24360_));
AND2X2 AND2X2_12571 ( .A(u2__abc_52155_new_n24349_), .B(u2_o_440_), .Y(u2__abc_52155_new_n24362_));
AND2X2 AND2X2_12572 ( .A(u2__abc_52155_new_n24363_), .B(u2__abc_52155_new_n24361_), .Y(u2__abc_52155_new_n24364_));
AND2X2 AND2X2_12573 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6983_), .Y(u2__abc_52155_new_n24366_));
AND2X2 AND2X2_12574 ( .A(u2__abc_52155_new_n24367_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24368_));
AND2X2 AND2X2_12575 ( .A(u2__abc_52155_new_n24365_), .B(u2__abc_52155_new_n24368_), .Y(u2__abc_52155_new_n24369_));
AND2X2 AND2X2_12576 ( .A(u2__abc_52155_new_n24370_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__442_));
AND2X2 AND2X2_12577 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_442_), .Y(u2__abc_52155_new_n24372_));
AND2X2 AND2X2_12578 ( .A(u2__abc_52155_new_n24362_), .B(u2_o_441_), .Y(u2__abc_52155_new_n24373_));
AND2X2 AND2X2_12579 ( .A(u2__abc_52155_new_n24374_), .B(u2__abc_52155_new_n24375_), .Y(u2__abc_52155_new_n24376_));
AND2X2 AND2X2_1258 ( .A(u2__abc_52155_new_n4577_), .B(u2__abc_52155_new_n4580_), .Y(u2__abc_52155_new_n4581_));
AND2X2 AND2X2_12580 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6949_), .Y(u2__abc_52155_new_n24378_));
AND2X2 AND2X2_12581 ( .A(u2__abc_52155_new_n24379_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24380_));
AND2X2 AND2X2_12582 ( .A(u2__abc_52155_new_n24377_), .B(u2__abc_52155_new_n24380_), .Y(u2__abc_52155_new_n24381_));
AND2X2 AND2X2_12583 ( .A(u2__abc_52155_new_n24382_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__443_));
AND2X2 AND2X2_12584 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_443_), .Y(u2__abc_52155_new_n24384_));
AND2X2 AND2X2_12585 ( .A(u2__abc_52155_new_n24373_), .B(u2_o_442_), .Y(u2__abc_52155_new_n24386_));
AND2X2 AND2X2_12586 ( .A(u2__abc_52155_new_n24387_), .B(u2__abc_52155_new_n24385_), .Y(u2__abc_52155_new_n24388_));
AND2X2 AND2X2_12587 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6945_), .Y(u2__abc_52155_new_n24390_));
AND2X2 AND2X2_12588 ( .A(u2__abc_52155_new_n24391_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24392_));
AND2X2 AND2X2_12589 ( .A(u2__abc_52155_new_n24389_), .B(u2__abc_52155_new_n24392_), .Y(u2__abc_52155_new_n24393_));
AND2X2 AND2X2_1259 ( .A(u2__abc_52155_new_n4582_), .B(u2_remHi_221_), .Y(u2__abc_52155_new_n4583_));
AND2X2 AND2X2_12590 ( .A(u2__abc_52155_new_n24394_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__444_));
AND2X2 AND2X2_12591 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_444_), .Y(u2__abc_52155_new_n24396_));
AND2X2 AND2X2_12592 ( .A(u2__abc_52155_new_n24386_), .B(u2_o_443_), .Y(u2__abc_52155_new_n24397_));
AND2X2 AND2X2_12593 ( .A(u2__abc_52155_new_n24398_), .B(u2__abc_52155_new_n24399_), .Y(u2__abc_52155_new_n24400_));
AND2X2 AND2X2_12594 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6927_), .Y(u2__abc_52155_new_n24402_));
AND2X2 AND2X2_12595 ( .A(u2__abc_52155_new_n24403_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24404_));
AND2X2 AND2X2_12596 ( .A(u2__abc_52155_new_n24401_), .B(u2__abc_52155_new_n24404_), .Y(u2__abc_52155_new_n24405_));
AND2X2 AND2X2_12597 ( .A(u2__abc_52155_new_n24406_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__445_));
AND2X2 AND2X2_12598 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_445_), .Y(u2__abc_52155_new_n24408_));
AND2X2 AND2X2_12599 ( .A(u2__abc_52155_new_n24397_), .B(u2_o_444_), .Y(u2__abc_52155_new_n24410_));
AND2X2 AND2X2_126 ( .A(_abc_73687_new_n978_), .B(_abc_73687_new_n977_), .Y(\o[161] ));
AND2X2 AND2X2_1260 ( .A(u2__abc_52155_new_n4585_), .B(sqrto_221_), .Y(u2__abc_52155_new_n4586_));
AND2X2 AND2X2_12600 ( .A(u2__abc_52155_new_n24411_), .B(u2__abc_52155_new_n24409_), .Y(u2__abc_52155_new_n24412_));
AND2X2 AND2X2_12601 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6937_), .Y(u2__abc_52155_new_n24414_));
AND2X2 AND2X2_12602 ( .A(u2__abc_52155_new_n24415_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24416_));
AND2X2 AND2X2_12603 ( .A(u2__abc_52155_new_n24413_), .B(u2__abc_52155_new_n24416_), .Y(u2__abc_52155_new_n24417_));
AND2X2 AND2X2_12604 ( .A(u2__abc_52155_new_n24418_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__446_));
AND2X2 AND2X2_12605 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_446_), .Y(u2__abc_52155_new_n24420_));
AND2X2 AND2X2_12606 ( .A(u2__abc_52155_new_n24410_), .B(u2_o_445_), .Y(u2__abc_52155_new_n24421_));
AND2X2 AND2X2_12607 ( .A(u2__abc_52155_new_n24422_), .B(u2__abc_52155_new_n24423_), .Y(u2__abc_52155_new_n24424_));
AND2X2 AND2X2_12608 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3025_), .Y(u2__abc_52155_new_n24426_));
AND2X2 AND2X2_12609 ( .A(u2__abc_52155_new_n24427_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24428_));
AND2X2 AND2X2_1261 ( .A(u2__abc_52155_new_n4584_), .B(u2__abc_52155_new_n4587_), .Y(u2__abc_52155_new_n4588_));
AND2X2 AND2X2_12610 ( .A(u2__abc_52155_new_n24425_), .B(u2__abc_52155_new_n24428_), .Y(u2__abc_52155_new_n24429_));
AND2X2 AND2X2_12611 ( .A(u2__abc_52155_new_n24430_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__447_));
AND2X2 AND2X2_12612 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_447_), .Y(u2__abc_52155_new_n24432_));
AND2X2 AND2X2_12613 ( .A(u2__abc_52155_new_n24421_), .B(u2_o_446_), .Y(u2__abc_52155_new_n24434_));
AND2X2 AND2X2_12614 ( .A(u2__abc_52155_new_n24435_), .B(u2__abc_52155_new_n24433_), .Y(u2__abc_52155_new_n24436_));
AND2X2 AND2X2_12615 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3018_), .Y(u2__abc_52155_new_n24438_));
AND2X2 AND2X2_12616 ( .A(u2__abc_52155_new_n24439_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24440_));
AND2X2 AND2X2_12617 ( .A(u2__abc_52155_new_n24437_), .B(u2__abc_52155_new_n24440_), .Y(u2__abc_52155_new_n24441_));
AND2X2 AND2X2_12618 ( .A(u2__abc_52155_new_n24442_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__448_));
AND2X2 AND2X2_12619 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_448_), .Y(u2__abc_52155_new_n24444_));
AND2X2 AND2X2_1262 ( .A(u2__abc_52155_new_n4581_), .B(u2__abc_52155_new_n4588_), .Y(u2__abc_52155_new_n4589_));
AND2X2 AND2X2_12620 ( .A(u2__abc_52155_new_n24434_), .B(u2_o_447_), .Y(u2__abc_52155_new_n24446_));
AND2X2 AND2X2_12621 ( .A(u2__abc_52155_new_n24447_), .B(u2__abc_52155_new_n24445_), .Y(u2__abc_52155_new_n24448_));
AND2X2 AND2X2_12622 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3013_), .Y(u2__abc_52155_new_n24450_));
AND2X2 AND2X2_12623 ( .A(u2__abc_52155_new_n24451_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24452_));
AND2X2 AND2X2_12624 ( .A(u2__abc_52155_new_n24449_), .B(u2__abc_52155_new_n24452_), .Y(u2__abc_52155_new_n24453_));
AND2X2 AND2X2_12625 ( .A(u2__abc_52155_new_n24454_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__449_));
AND2X2 AND2X2_12626 ( .A(u2__abc_52155_new_n3002_), .B(u2_o_449_), .Y(u2__abc_52155_new_n24456_));
AND2X2 AND2X2_12627 ( .A(u2__abc_52155_new_n24446_), .B(u2_o_448_), .Y(u2__abc_52155_new_n24458_));
AND2X2 AND2X2_12628 ( .A(u2__abc_52155_new_n24459_), .B(u2__abc_52155_new_n24457_), .Y(u2__abc_52155_new_n24460_));
AND2X2 AND2X2_12629 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3007_), .Y(u2__abc_52155_new_n24462_));
AND2X2 AND2X2_1263 ( .A(u2__abc_52155_new_n4590_), .B(u2_remHi_219_), .Y(u2__abc_52155_new_n4591_));
AND2X2 AND2X2_12630 ( .A(u2__abc_52155_new_n24463_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n24464_));
AND2X2 AND2X2_12631 ( .A(u2__abc_52155_new_n24461_), .B(u2__abc_52155_new_n24464_), .Y(u2__abc_52155_new_n24465_));
AND2X2 AND2X2_12632 ( .A(u2__abc_52155_new_n24466_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__450_));
AND2X2 AND2X2_1264 ( .A(u2__abc_52155_new_n4593_), .B(sqrto_219_), .Y(u2__abc_52155_new_n4594_));
AND2X2 AND2X2_1265 ( .A(u2__abc_52155_new_n4592_), .B(u2__abc_52155_new_n4595_), .Y(u2__abc_52155_new_n4596_));
AND2X2 AND2X2_1266 ( .A(u2__abc_52155_new_n4597_), .B(u2_remHi_218_), .Y(u2__abc_52155_new_n4598_));
AND2X2 AND2X2_1267 ( .A(u2__abc_52155_new_n4600_), .B(sqrto_218_), .Y(u2__abc_52155_new_n4601_));
AND2X2 AND2X2_1268 ( .A(u2__abc_52155_new_n4599_), .B(u2__abc_52155_new_n4602_), .Y(u2__abc_52155_new_n4603_));
AND2X2 AND2X2_1269 ( .A(u2__abc_52155_new_n4596_), .B(u2__abc_52155_new_n4603_), .Y(u2__abc_52155_new_n4604_));
AND2X2 AND2X2_127 ( .A(_abc_73687_new_n981_), .B(_abc_73687_new_n980_), .Y(\o[162] ));
AND2X2 AND2X2_1270 ( .A(u2__abc_52155_new_n4589_), .B(u2__abc_52155_new_n4604_), .Y(u2__abc_52155_new_n4605_));
AND2X2 AND2X2_1271 ( .A(u2__abc_52155_new_n4574_), .B(u2__abc_52155_new_n4605_), .Y(u2__abc_52155_new_n4606_));
AND2X2 AND2X2_1272 ( .A(u2__abc_52155_new_n4607_), .B(u2_remHi_208_), .Y(u2__abc_52155_new_n4608_));
AND2X2 AND2X2_1273 ( .A(u2__abc_52155_new_n4610_), .B(sqrto_208_), .Y(u2__abc_52155_new_n4611_));
AND2X2 AND2X2_1274 ( .A(u2__abc_52155_new_n4609_), .B(u2__abc_52155_new_n4612_), .Y(u2__abc_52155_new_n4613_));
AND2X2 AND2X2_1275 ( .A(u2__abc_52155_new_n4614_), .B(u2_remHi_209_), .Y(u2__abc_52155_new_n4615_));
AND2X2 AND2X2_1276 ( .A(u2__abc_52155_new_n4617_), .B(sqrto_209_), .Y(u2__abc_52155_new_n4618_));
AND2X2 AND2X2_1277 ( .A(u2__abc_52155_new_n4616_), .B(u2__abc_52155_new_n4619_), .Y(u2__abc_52155_new_n4620_));
AND2X2 AND2X2_1278 ( .A(u2__abc_52155_new_n4613_), .B(u2__abc_52155_new_n4620_), .Y(u2__abc_52155_new_n4621_));
AND2X2 AND2X2_1279 ( .A(u2__abc_52155_new_n4622_), .B(u2_remHi_206_), .Y(u2__abc_52155_new_n4623_));
AND2X2 AND2X2_128 ( .A(_abc_73687_new_n984_), .B(_abc_73687_new_n983_), .Y(\o[163] ));
AND2X2 AND2X2_1280 ( .A(u2__abc_52155_new_n4625_), .B(sqrto_206_), .Y(u2__abc_52155_new_n4626_));
AND2X2 AND2X2_1281 ( .A(u2__abc_52155_new_n4624_), .B(u2__abc_52155_new_n4627_), .Y(u2__abc_52155_new_n4628_));
AND2X2 AND2X2_1282 ( .A(u2__abc_52155_new_n4629_), .B(u2_remHi_207_), .Y(u2__abc_52155_new_n4630_));
AND2X2 AND2X2_1283 ( .A(u2__abc_52155_new_n4632_), .B(sqrto_207_), .Y(u2__abc_52155_new_n4633_));
AND2X2 AND2X2_1284 ( .A(u2__abc_52155_new_n4631_), .B(u2__abc_52155_new_n4634_), .Y(u2__abc_52155_new_n4635_));
AND2X2 AND2X2_1285 ( .A(u2__abc_52155_new_n4628_), .B(u2__abc_52155_new_n4635_), .Y(u2__abc_52155_new_n4636_));
AND2X2 AND2X2_1286 ( .A(u2__abc_52155_new_n4621_), .B(u2__abc_52155_new_n4636_), .Y(u2__abc_52155_new_n4637_));
AND2X2 AND2X2_1287 ( .A(u2__abc_52155_new_n4638_), .B(u2_remHi_212_), .Y(u2__abc_52155_new_n4639_));
AND2X2 AND2X2_1288 ( .A(u2__abc_52155_new_n4641_), .B(sqrto_212_), .Y(u2__abc_52155_new_n4642_));
AND2X2 AND2X2_1289 ( .A(u2__abc_52155_new_n4640_), .B(u2__abc_52155_new_n4643_), .Y(u2__abc_52155_new_n4644_));
AND2X2 AND2X2_129 ( .A(_abc_73687_new_n987_), .B(_abc_73687_new_n986_), .Y(\o[164] ));
AND2X2 AND2X2_1290 ( .A(u2__abc_52155_new_n4645_), .B(u2_remHi_213_), .Y(u2__abc_52155_new_n4646_));
AND2X2 AND2X2_1291 ( .A(u2__abc_52155_new_n4648_), .B(sqrto_213_), .Y(u2__abc_52155_new_n4649_));
AND2X2 AND2X2_1292 ( .A(u2__abc_52155_new_n4647_), .B(u2__abc_52155_new_n4650_), .Y(u2__abc_52155_new_n4651_));
AND2X2 AND2X2_1293 ( .A(u2__abc_52155_new_n4644_), .B(u2__abc_52155_new_n4651_), .Y(u2__abc_52155_new_n4652_));
AND2X2 AND2X2_1294 ( .A(u2__abc_52155_new_n4653_), .B(u2_remHi_211_), .Y(u2__abc_52155_new_n4654_));
AND2X2 AND2X2_1295 ( .A(u2__abc_52155_new_n4656_), .B(sqrto_211_), .Y(u2__abc_52155_new_n4657_));
AND2X2 AND2X2_1296 ( .A(u2__abc_52155_new_n4655_), .B(u2__abc_52155_new_n4658_), .Y(u2__abc_52155_new_n4659_));
AND2X2 AND2X2_1297 ( .A(u2__abc_52155_new_n4660_), .B(u2_remHi_210_), .Y(u2__abc_52155_new_n4661_));
AND2X2 AND2X2_1298 ( .A(u2__abc_52155_new_n4663_), .B(sqrto_210_), .Y(u2__abc_52155_new_n4664_));
AND2X2 AND2X2_1299 ( .A(u2__abc_52155_new_n4662_), .B(u2__abc_52155_new_n4665_), .Y(u2__abc_52155_new_n4666_));
AND2X2 AND2X2_13 ( .A(_abc_73687_new_n753_), .B(sqrto_12_), .Y(\o[48] ));
AND2X2 AND2X2_130 ( .A(_abc_73687_new_n990_), .B(_abc_73687_new_n989_), .Y(\o[165] ));
AND2X2 AND2X2_1300 ( .A(u2__abc_52155_new_n4659_), .B(u2__abc_52155_new_n4666_), .Y(u2__abc_52155_new_n4667_));
AND2X2 AND2X2_1301 ( .A(u2__abc_52155_new_n4652_), .B(u2__abc_52155_new_n4667_), .Y(u2__abc_52155_new_n4668_));
AND2X2 AND2X2_1302 ( .A(u2__abc_52155_new_n4637_), .B(u2__abc_52155_new_n4668_), .Y(u2__abc_52155_new_n4669_));
AND2X2 AND2X2_1303 ( .A(u2__abc_52155_new_n4606_), .B(u2__abc_52155_new_n4669_), .Y(u2__abc_52155_new_n4670_));
AND2X2 AND2X2_1304 ( .A(u2__abc_52155_new_n4671_), .B(u2_remHi_200_), .Y(u2__abc_52155_new_n4672_));
AND2X2 AND2X2_1305 ( .A(u2__abc_52155_new_n4674_), .B(sqrto_200_), .Y(u2__abc_52155_new_n4675_));
AND2X2 AND2X2_1306 ( .A(u2__abc_52155_new_n4673_), .B(u2__abc_52155_new_n4676_), .Y(u2__abc_52155_new_n4677_));
AND2X2 AND2X2_1307 ( .A(u2__abc_52155_new_n4678_), .B(u2_remHi_201_), .Y(u2__abc_52155_new_n4679_));
AND2X2 AND2X2_1308 ( .A(u2__abc_52155_new_n4681_), .B(sqrto_201_), .Y(u2__abc_52155_new_n4682_));
AND2X2 AND2X2_1309 ( .A(u2__abc_52155_new_n4680_), .B(u2__abc_52155_new_n4683_), .Y(u2__abc_52155_new_n4684_));
AND2X2 AND2X2_131 ( .A(_abc_73687_new_n993_), .B(_abc_73687_new_n992_), .Y(\o[166] ));
AND2X2 AND2X2_1310 ( .A(u2__abc_52155_new_n4677_), .B(u2__abc_52155_new_n4684_), .Y(u2__abc_52155_new_n4685_));
AND2X2 AND2X2_1311 ( .A(u2__abc_52155_new_n4686_), .B(u2_remHi_199_), .Y(u2__abc_52155_new_n4687_));
AND2X2 AND2X2_1312 ( .A(u2__abc_52155_new_n4689_), .B(sqrto_199_), .Y(u2__abc_52155_new_n4690_));
AND2X2 AND2X2_1313 ( .A(u2__abc_52155_new_n4688_), .B(u2__abc_52155_new_n4691_), .Y(u2__abc_52155_new_n4692_));
AND2X2 AND2X2_1314 ( .A(u2__abc_52155_new_n4693_), .B(u2_remHi_198_), .Y(u2__abc_52155_new_n4694_));
AND2X2 AND2X2_1315 ( .A(u2__abc_52155_new_n4696_), .B(sqrto_198_), .Y(u2__abc_52155_new_n4697_));
AND2X2 AND2X2_1316 ( .A(u2__abc_52155_new_n4695_), .B(u2__abc_52155_new_n4698_), .Y(u2__abc_52155_new_n4699_));
AND2X2 AND2X2_1317 ( .A(u2__abc_52155_new_n4692_), .B(u2__abc_52155_new_n4699_), .Y(u2__abc_52155_new_n4700_));
AND2X2 AND2X2_1318 ( .A(u2__abc_52155_new_n4685_), .B(u2__abc_52155_new_n4700_), .Y(u2__abc_52155_new_n4701_));
AND2X2 AND2X2_1319 ( .A(u2__abc_52155_new_n4702_), .B(u2_remHi_204_), .Y(u2__abc_52155_new_n4703_));
AND2X2 AND2X2_132 ( .A(_abc_73687_new_n996_), .B(_abc_73687_new_n995_), .Y(\o[167] ));
AND2X2 AND2X2_1320 ( .A(u2__abc_52155_new_n4705_), .B(sqrto_204_), .Y(u2__abc_52155_new_n4706_));
AND2X2 AND2X2_1321 ( .A(u2__abc_52155_new_n4704_), .B(u2__abc_52155_new_n4707_), .Y(u2__abc_52155_new_n4708_));
AND2X2 AND2X2_1322 ( .A(u2__abc_52155_new_n4709_), .B(u2_remHi_205_), .Y(u2__abc_52155_new_n4710_));
AND2X2 AND2X2_1323 ( .A(u2__abc_52155_new_n4712_), .B(sqrto_205_), .Y(u2__abc_52155_new_n4713_));
AND2X2 AND2X2_1324 ( .A(u2__abc_52155_new_n4711_), .B(u2__abc_52155_new_n4714_), .Y(u2__abc_52155_new_n4715_));
AND2X2 AND2X2_1325 ( .A(u2__abc_52155_new_n4708_), .B(u2__abc_52155_new_n4715_), .Y(u2__abc_52155_new_n4716_));
AND2X2 AND2X2_1326 ( .A(u2__abc_52155_new_n4717_), .B(u2_remHi_203_), .Y(u2__abc_52155_new_n4718_));
AND2X2 AND2X2_1327 ( .A(u2__abc_52155_new_n4720_), .B(sqrto_203_), .Y(u2__abc_52155_new_n4721_));
AND2X2 AND2X2_1328 ( .A(u2__abc_52155_new_n4719_), .B(u2__abc_52155_new_n4722_), .Y(u2__abc_52155_new_n4723_));
AND2X2 AND2X2_1329 ( .A(u2__abc_52155_new_n4724_), .B(u2_remHi_202_), .Y(u2__abc_52155_new_n4725_));
AND2X2 AND2X2_133 ( .A(_abc_73687_new_n999_), .B(_abc_73687_new_n998_), .Y(\o[168] ));
AND2X2 AND2X2_1330 ( .A(u2__abc_52155_new_n4727_), .B(sqrto_202_), .Y(u2__abc_52155_new_n4728_));
AND2X2 AND2X2_1331 ( .A(u2__abc_52155_new_n4726_), .B(u2__abc_52155_new_n4729_), .Y(u2__abc_52155_new_n4730_));
AND2X2 AND2X2_1332 ( .A(u2__abc_52155_new_n4723_), .B(u2__abc_52155_new_n4730_), .Y(u2__abc_52155_new_n4731_));
AND2X2 AND2X2_1333 ( .A(u2__abc_52155_new_n4716_), .B(u2__abc_52155_new_n4731_), .Y(u2__abc_52155_new_n4732_));
AND2X2 AND2X2_1334 ( .A(u2__abc_52155_new_n4701_), .B(u2__abc_52155_new_n4732_), .Y(u2__abc_52155_new_n4733_));
AND2X2 AND2X2_1335 ( .A(u2__abc_52155_new_n4734_), .B(u2_remHi_196_), .Y(u2__abc_52155_new_n4735_));
AND2X2 AND2X2_1336 ( .A(u2__abc_52155_new_n4737_), .B(sqrto_196_), .Y(u2__abc_52155_new_n4738_));
AND2X2 AND2X2_1337 ( .A(u2__abc_52155_new_n4736_), .B(u2__abc_52155_new_n4739_), .Y(u2__abc_52155_new_n4740_));
AND2X2 AND2X2_1338 ( .A(u2__abc_52155_new_n4741_), .B(u2_remHi_197_), .Y(u2__abc_52155_new_n4742_));
AND2X2 AND2X2_1339 ( .A(u2__abc_52155_new_n4744_), .B(sqrto_197_), .Y(u2__abc_52155_new_n4745_));
AND2X2 AND2X2_134 ( .A(_abc_73687_new_n1002_), .B(_abc_73687_new_n1001_), .Y(\o[169] ));
AND2X2 AND2X2_1340 ( .A(u2__abc_52155_new_n4743_), .B(u2__abc_52155_new_n4746_), .Y(u2__abc_52155_new_n4747_));
AND2X2 AND2X2_1341 ( .A(u2__abc_52155_new_n4740_), .B(u2__abc_52155_new_n4747_), .Y(u2__abc_52155_new_n4748_));
AND2X2 AND2X2_1342 ( .A(u2__abc_52155_new_n4749_), .B(u2_remHi_195_), .Y(u2__abc_52155_new_n4750_));
AND2X2 AND2X2_1343 ( .A(u2__abc_52155_new_n4752_), .B(sqrto_195_), .Y(u2__abc_52155_new_n4753_));
AND2X2 AND2X2_1344 ( .A(u2__abc_52155_new_n4751_), .B(u2__abc_52155_new_n4754_), .Y(u2__abc_52155_new_n4755_));
AND2X2 AND2X2_1345 ( .A(u2__abc_52155_new_n4756_), .B(u2_remHi_194_), .Y(u2__abc_52155_new_n4757_));
AND2X2 AND2X2_1346 ( .A(u2__abc_52155_new_n4759_), .B(sqrto_194_), .Y(u2__abc_52155_new_n4760_));
AND2X2 AND2X2_1347 ( .A(u2__abc_52155_new_n4758_), .B(u2__abc_52155_new_n4761_), .Y(u2__abc_52155_new_n4762_));
AND2X2 AND2X2_1348 ( .A(u2__abc_52155_new_n4755_), .B(u2__abc_52155_new_n4762_), .Y(u2__abc_52155_new_n4763_));
AND2X2 AND2X2_1349 ( .A(u2__abc_52155_new_n4748_), .B(u2__abc_52155_new_n4763_), .Y(u2__abc_52155_new_n4764_));
AND2X2 AND2X2_135 ( .A(_abc_73687_new_n1005_), .B(_abc_73687_new_n1004_), .Y(\o[170] ));
AND2X2 AND2X2_1350 ( .A(u2__abc_52155_new_n4765_), .B(u2_remHi_192_), .Y(u2__abc_52155_new_n4766_));
AND2X2 AND2X2_1351 ( .A(u2__abc_52155_new_n4767_), .B(sqrto_192_), .Y(u2__abc_52155_new_n4768_));
AND2X2 AND2X2_1352 ( .A(u2__abc_52155_new_n4770_), .B(u2_remHi_193_), .Y(u2__abc_52155_new_n4771_));
AND2X2 AND2X2_1353 ( .A(u2__abc_52155_new_n4772_), .B(sqrto_193_), .Y(u2__abc_52155_new_n4773_));
AND2X2 AND2X2_1354 ( .A(u2__abc_52155_new_n4777_), .B(u2_remHi_190_), .Y(u2__abc_52155_new_n4778_));
AND2X2 AND2X2_1355 ( .A(u2__abc_52155_new_n4780_), .B(sqrto_190_), .Y(u2__abc_52155_new_n4781_));
AND2X2 AND2X2_1356 ( .A(u2__abc_52155_new_n4779_), .B(u2__abc_52155_new_n4782_), .Y(u2__abc_52155_new_n4783_));
AND2X2 AND2X2_1357 ( .A(u2__abc_52155_new_n4784_), .B(u2_remHi_191_), .Y(u2__abc_52155_new_n4785_));
AND2X2 AND2X2_1358 ( .A(u2__abc_52155_new_n4787_), .B(sqrto_191_), .Y(u2__abc_52155_new_n4788_));
AND2X2 AND2X2_1359 ( .A(u2__abc_52155_new_n4786_), .B(u2__abc_52155_new_n4789_), .Y(u2__abc_52155_new_n4790_));
AND2X2 AND2X2_136 ( .A(_abc_73687_new_n1008_), .B(_abc_73687_new_n1007_), .Y(\o[171] ));
AND2X2 AND2X2_1360 ( .A(u2__abc_52155_new_n4783_), .B(u2__abc_52155_new_n4790_), .Y(u2__abc_52155_new_n4791_));
AND2X2 AND2X2_1361 ( .A(u2__abc_52155_new_n4776_), .B(u2__abc_52155_new_n4791_), .Y(u2__abc_52155_new_n4792_));
AND2X2 AND2X2_1362 ( .A(u2__abc_52155_new_n4792_), .B(u2__abc_52155_new_n4764_), .Y(u2__abc_52155_new_n4793_));
AND2X2 AND2X2_1363 ( .A(u2__abc_52155_new_n4793_), .B(u2__abc_52155_new_n4733_), .Y(u2__abc_52155_new_n4794_));
AND2X2 AND2X2_1364 ( .A(u2__abc_52155_new_n4794_), .B(u2__abc_52155_new_n4670_), .Y(u2__abc_52155_new_n4795_));
AND2X2 AND2X2_1365 ( .A(u2__abc_52155_new_n4795_), .B(u2__abc_52155_new_n4543_), .Y(u2__abc_52155_new_n4796_));
AND2X2 AND2X2_1366 ( .A(u2__abc_52155_new_n4797_), .B(u2_remHi_182_), .Y(u2__abc_52155_new_n4798_));
AND2X2 AND2X2_1367 ( .A(u2__abc_52155_new_n4800_), .B(sqrto_182_), .Y(u2__abc_52155_new_n4801_));
AND2X2 AND2X2_1368 ( .A(u2__abc_52155_new_n4799_), .B(u2__abc_52155_new_n4802_), .Y(u2__abc_52155_new_n4803_));
AND2X2 AND2X2_1369 ( .A(u2__abc_52155_new_n4804_), .B(u2_remHi_183_), .Y(u2__abc_52155_new_n4805_));
AND2X2 AND2X2_137 ( .A(_abc_73687_new_n1011_), .B(_abc_73687_new_n1010_), .Y(\o[172] ));
AND2X2 AND2X2_1370 ( .A(u2__abc_52155_new_n4807_), .B(sqrto_183_), .Y(u2__abc_52155_new_n4808_));
AND2X2 AND2X2_1371 ( .A(u2__abc_52155_new_n4806_), .B(u2__abc_52155_new_n4809_), .Y(u2__abc_52155_new_n4810_));
AND2X2 AND2X2_1372 ( .A(u2__abc_52155_new_n4803_), .B(u2__abc_52155_new_n4810_), .Y(u2__abc_52155_new_n4811_));
AND2X2 AND2X2_1373 ( .A(u2__abc_52155_new_n4812_), .B(u2_remHi_184_), .Y(u2__abc_52155_new_n4813_));
AND2X2 AND2X2_1374 ( .A(u2__abc_52155_new_n4815_), .B(sqrto_184_), .Y(u2__abc_52155_new_n4816_));
AND2X2 AND2X2_1375 ( .A(u2__abc_52155_new_n4814_), .B(u2__abc_52155_new_n4817_), .Y(u2__abc_52155_new_n4818_));
AND2X2 AND2X2_1376 ( .A(u2__abc_52155_new_n4819_), .B(u2_remHi_185_), .Y(u2__abc_52155_new_n4820_));
AND2X2 AND2X2_1377 ( .A(u2__abc_52155_new_n4822_), .B(sqrto_185_), .Y(u2__abc_52155_new_n4823_));
AND2X2 AND2X2_1378 ( .A(u2__abc_52155_new_n4821_), .B(u2__abc_52155_new_n4824_), .Y(u2__abc_52155_new_n4825_));
AND2X2 AND2X2_1379 ( .A(u2__abc_52155_new_n4818_), .B(u2__abc_52155_new_n4825_), .Y(u2__abc_52155_new_n4826_));
AND2X2 AND2X2_138 ( .A(_abc_73687_new_n1014_), .B(_abc_73687_new_n1013_), .Y(\o[173] ));
AND2X2 AND2X2_1380 ( .A(u2__abc_52155_new_n4811_), .B(u2__abc_52155_new_n4826_), .Y(u2__abc_52155_new_n4827_));
AND2X2 AND2X2_1381 ( .A(u2__abc_52155_new_n4828_), .B(u2_remHi_188_), .Y(u2__abc_52155_new_n4829_));
AND2X2 AND2X2_1382 ( .A(u2__abc_52155_new_n4831_), .B(sqrto_188_), .Y(u2__abc_52155_new_n4832_));
AND2X2 AND2X2_1383 ( .A(u2__abc_52155_new_n4830_), .B(u2__abc_52155_new_n4833_), .Y(u2__abc_52155_new_n4834_));
AND2X2 AND2X2_1384 ( .A(u2__abc_52155_new_n4835_), .B(u2_remHi_189_), .Y(u2__abc_52155_new_n4836_));
AND2X2 AND2X2_1385 ( .A(u2__abc_52155_new_n4838_), .B(sqrto_189_), .Y(u2__abc_52155_new_n4839_));
AND2X2 AND2X2_1386 ( .A(u2__abc_52155_new_n4837_), .B(u2__abc_52155_new_n4840_), .Y(u2__abc_52155_new_n4841_));
AND2X2 AND2X2_1387 ( .A(u2__abc_52155_new_n4834_), .B(u2__abc_52155_new_n4841_), .Y(u2__abc_52155_new_n4842_));
AND2X2 AND2X2_1388 ( .A(u2__abc_52155_new_n4843_), .B(u2_remHi_187_), .Y(u2__abc_52155_new_n4844_));
AND2X2 AND2X2_1389 ( .A(u2__abc_52155_new_n4846_), .B(sqrto_187_), .Y(u2__abc_52155_new_n4847_));
AND2X2 AND2X2_139 ( .A(_abc_73687_new_n1017_), .B(_abc_73687_new_n1016_), .Y(\o[174] ));
AND2X2 AND2X2_1390 ( .A(u2__abc_52155_new_n4845_), .B(u2__abc_52155_new_n4848_), .Y(u2__abc_52155_new_n4849_));
AND2X2 AND2X2_1391 ( .A(u2__abc_52155_new_n4850_), .B(u2_remHi_186_), .Y(u2__abc_52155_new_n4851_));
AND2X2 AND2X2_1392 ( .A(u2__abc_52155_new_n4853_), .B(sqrto_186_), .Y(u2__abc_52155_new_n4854_));
AND2X2 AND2X2_1393 ( .A(u2__abc_52155_new_n4852_), .B(u2__abc_52155_new_n4855_), .Y(u2__abc_52155_new_n4856_));
AND2X2 AND2X2_1394 ( .A(u2__abc_52155_new_n4849_), .B(u2__abc_52155_new_n4856_), .Y(u2__abc_52155_new_n4857_));
AND2X2 AND2X2_1395 ( .A(u2__abc_52155_new_n4842_), .B(u2__abc_52155_new_n4857_), .Y(u2__abc_52155_new_n4858_));
AND2X2 AND2X2_1396 ( .A(u2__abc_52155_new_n4827_), .B(u2__abc_52155_new_n4858_), .Y(u2__abc_52155_new_n4859_));
AND2X2 AND2X2_1397 ( .A(u2__abc_52155_new_n4860_), .B(u2_remHi_180_), .Y(u2__abc_52155_new_n4861_));
AND2X2 AND2X2_1398 ( .A(u2__abc_52155_new_n4863_), .B(sqrto_180_), .Y(u2__abc_52155_new_n4864_));
AND2X2 AND2X2_1399 ( .A(u2__abc_52155_new_n4862_), .B(u2__abc_52155_new_n4865_), .Y(u2__abc_52155_new_n4866_));
AND2X2 AND2X2_14 ( .A(_abc_73687_new_n753_), .B(sqrto_13_), .Y(\o[49] ));
AND2X2 AND2X2_140 ( .A(_abc_73687_new_n1020_), .B(_abc_73687_new_n1019_), .Y(\o[175] ));
AND2X2 AND2X2_1400 ( .A(u2__abc_52155_new_n4867_), .B(u2_remHi_181_), .Y(u2__abc_52155_new_n4868_));
AND2X2 AND2X2_1401 ( .A(u2__abc_52155_new_n4870_), .B(sqrto_181_), .Y(u2__abc_52155_new_n4871_));
AND2X2 AND2X2_1402 ( .A(u2__abc_52155_new_n4869_), .B(u2__abc_52155_new_n4872_), .Y(u2__abc_52155_new_n4873_));
AND2X2 AND2X2_1403 ( .A(u2__abc_52155_new_n4866_), .B(u2__abc_52155_new_n4873_), .Y(u2__abc_52155_new_n4874_));
AND2X2 AND2X2_1404 ( .A(u2__abc_52155_new_n4875_), .B(u2_remHi_179_), .Y(u2__abc_52155_new_n4876_));
AND2X2 AND2X2_1405 ( .A(u2__abc_52155_new_n4878_), .B(sqrto_179_), .Y(u2__abc_52155_new_n4879_));
AND2X2 AND2X2_1406 ( .A(u2__abc_52155_new_n4877_), .B(u2__abc_52155_new_n4880_), .Y(u2__abc_52155_new_n4881_));
AND2X2 AND2X2_1407 ( .A(u2__abc_52155_new_n4882_), .B(u2_remHi_178_), .Y(u2__abc_52155_new_n4883_));
AND2X2 AND2X2_1408 ( .A(u2__abc_52155_new_n4885_), .B(sqrto_178_), .Y(u2__abc_52155_new_n4886_));
AND2X2 AND2X2_1409 ( .A(u2__abc_52155_new_n4884_), .B(u2__abc_52155_new_n4887_), .Y(u2__abc_52155_new_n4888_));
AND2X2 AND2X2_141 ( .A(_abc_73687_new_n1023_), .B(_abc_73687_new_n1022_), .Y(\o[176] ));
AND2X2 AND2X2_1410 ( .A(u2__abc_52155_new_n4881_), .B(u2__abc_52155_new_n4888_), .Y(u2__abc_52155_new_n4889_));
AND2X2 AND2X2_1411 ( .A(u2__abc_52155_new_n4874_), .B(u2__abc_52155_new_n4889_), .Y(u2__abc_52155_new_n4890_));
AND2X2 AND2X2_1412 ( .A(u2__abc_52155_new_n4891_), .B(u2_remHi_176_), .Y(u2__abc_52155_new_n4892_));
AND2X2 AND2X2_1413 ( .A(u2__abc_52155_new_n4894_), .B(sqrto_176_), .Y(u2__abc_52155_new_n4895_));
AND2X2 AND2X2_1414 ( .A(u2__abc_52155_new_n4893_), .B(u2__abc_52155_new_n4896_), .Y(u2__abc_52155_new_n4897_));
AND2X2 AND2X2_1415 ( .A(u2__abc_52155_new_n4898_), .B(u2_remHi_177_), .Y(u2__abc_52155_new_n4899_));
AND2X2 AND2X2_1416 ( .A(u2__abc_52155_new_n4901_), .B(sqrto_177_), .Y(u2__abc_52155_new_n4902_));
AND2X2 AND2X2_1417 ( .A(u2__abc_52155_new_n4900_), .B(u2__abc_52155_new_n4903_), .Y(u2__abc_52155_new_n4904_));
AND2X2 AND2X2_1418 ( .A(u2__abc_52155_new_n4897_), .B(u2__abc_52155_new_n4904_), .Y(u2__abc_52155_new_n4905_));
AND2X2 AND2X2_1419 ( .A(u2__abc_52155_new_n4906_), .B(u2_remHi_174_), .Y(u2__abc_52155_new_n4907_));
AND2X2 AND2X2_142 ( .A(_abc_73687_new_n1026_), .B(_abc_73687_new_n1025_), .Y(\o[177] ));
AND2X2 AND2X2_1420 ( .A(u2__abc_52155_new_n4909_), .B(sqrto_174_), .Y(u2__abc_52155_new_n4910_));
AND2X2 AND2X2_1421 ( .A(u2__abc_52155_new_n4908_), .B(u2__abc_52155_new_n4911_), .Y(u2__abc_52155_new_n4912_));
AND2X2 AND2X2_1422 ( .A(u2__abc_52155_new_n4913_), .B(u2_remHi_175_), .Y(u2__abc_52155_new_n4914_));
AND2X2 AND2X2_1423 ( .A(u2__abc_52155_new_n4916_), .B(sqrto_175_), .Y(u2__abc_52155_new_n4917_));
AND2X2 AND2X2_1424 ( .A(u2__abc_52155_new_n4915_), .B(u2__abc_52155_new_n4918_), .Y(u2__abc_52155_new_n4919_));
AND2X2 AND2X2_1425 ( .A(u2__abc_52155_new_n4912_), .B(u2__abc_52155_new_n4919_), .Y(u2__abc_52155_new_n4920_));
AND2X2 AND2X2_1426 ( .A(u2__abc_52155_new_n4905_), .B(u2__abc_52155_new_n4920_), .Y(u2__abc_52155_new_n4921_));
AND2X2 AND2X2_1427 ( .A(u2__abc_52155_new_n4890_), .B(u2__abc_52155_new_n4921_), .Y(u2__abc_52155_new_n4922_));
AND2X2 AND2X2_1428 ( .A(u2__abc_52155_new_n4859_), .B(u2__abc_52155_new_n4922_), .Y(u2__abc_52155_new_n4923_));
AND2X2 AND2X2_1429 ( .A(u2__abc_52155_new_n4924_), .B(u2_remHi_172_), .Y(u2__abc_52155_new_n4925_));
AND2X2 AND2X2_143 ( .A(_abc_73687_new_n1029_), .B(_abc_73687_new_n1028_), .Y(\o[178] ));
AND2X2 AND2X2_1430 ( .A(u2__abc_52155_new_n4927_), .B(sqrto_172_), .Y(u2__abc_52155_new_n4928_));
AND2X2 AND2X2_1431 ( .A(u2__abc_52155_new_n4926_), .B(u2__abc_52155_new_n4929_), .Y(u2__abc_52155_new_n4930_));
AND2X2 AND2X2_1432 ( .A(u2__abc_52155_new_n4931_), .B(u2_remHi_173_), .Y(u2__abc_52155_new_n4932_));
AND2X2 AND2X2_1433 ( .A(u2__abc_52155_new_n4934_), .B(sqrto_173_), .Y(u2__abc_52155_new_n4935_));
AND2X2 AND2X2_1434 ( .A(u2__abc_52155_new_n4933_), .B(u2__abc_52155_new_n4936_), .Y(u2__abc_52155_new_n4937_));
AND2X2 AND2X2_1435 ( .A(u2__abc_52155_new_n4930_), .B(u2__abc_52155_new_n4937_), .Y(u2__abc_52155_new_n4938_));
AND2X2 AND2X2_1436 ( .A(u2__abc_52155_new_n4939_), .B(u2_remHi_171_), .Y(u2__abc_52155_new_n4940_));
AND2X2 AND2X2_1437 ( .A(u2__abc_52155_new_n4942_), .B(sqrto_171_), .Y(u2__abc_52155_new_n4943_));
AND2X2 AND2X2_1438 ( .A(u2__abc_52155_new_n4941_), .B(u2__abc_52155_new_n4944_), .Y(u2__abc_52155_new_n4945_));
AND2X2 AND2X2_1439 ( .A(u2__abc_52155_new_n4946_), .B(u2_remHi_170_), .Y(u2__abc_52155_new_n4947_));
AND2X2 AND2X2_144 ( .A(_abc_73687_new_n1032_), .B(_abc_73687_new_n1031_), .Y(\o[179] ));
AND2X2 AND2X2_1440 ( .A(u2__abc_52155_new_n4949_), .B(sqrto_170_), .Y(u2__abc_52155_new_n4950_));
AND2X2 AND2X2_1441 ( .A(u2__abc_52155_new_n4948_), .B(u2__abc_52155_new_n4951_), .Y(u2__abc_52155_new_n4952_));
AND2X2 AND2X2_1442 ( .A(u2__abc_52155_new_n4945_), .B(u2__abc_52155_new_n4952_), .Y(u2__abc_52155_new_n4953_));
AND2X2 AND2X2_1443 ( .A(u2__abc_52155_new_n4938_), .B(u2__abc_52155_new_n4953_), .Y(u2__abc_52155_new_n4954_));
AND2X2 AND2X2_1444 ( .A(u2__abc_52155_new_n4955_), .B(u2_remHi_168_), .Y(u2__abc_52155_new_n4956_));
AND2X2 AND2X2_1445 ( .A(u2__abc_52155_new_n4958_), .B(sqrto_168_), .Y(u2__abc_52155_new_n4959_));
AND2X2 AND2X2_1446 ( .A(u2__abc_52155_new_n4957_), .B(u2__abc_52155_new_n4960_), .Y(u2__abc_52155_new_n4961_));
AND2X2 AND2X2_1447 ( .A(u2__abc_52155_new_n4962_), .B(u2_remHi_169_), .Y(u2__abc_52155_new_n4963_));
AND2X2 AND2X2_1448 ( .A(u2__abc_52155_new_n4965_), .B(sqrto_169_), .Y(u2__abc_52155_new_n4966_));
AND2X2 AND2X2_1449 ( .A(u2__abc_52155_new_n4964_), .B(u2__abc_52155_new_n4967_), .Y(u2__abc_52155_new_n4968_));
AND2X2 AND2X2_145 ( .A(_abc_73687_new_n1035_), .B(_abc_73687_new_n1034_), .Y(\o[180] ));
AND2X2 AND2X2_1450 ( .A(u2__abc_52155_new_n4961_), .B(u2__abc_52155_new_n4968_), .Y(u2__abc_52155_new_n4969_));
AND2X2 AND2X2_1451 ( .A(u2__abc_52155_new_n4970_), .B(u2_remHi_167_), .Y(u2__abc_52155_new_n4971_));
AND2X2 AND2X2_1452 ( .A(u2__abc_52155_new_n4973_), .B(sqrto_167_), .Y(u2__abc_52155_new_n4974_));
AND2X2 AND2X2_1453 ( .A(u2__abc_52155_new_n4972_), .B(u2__abc_52155_new_n4975_), .Y(u2__abc_52155_new_n4976_));
AND2X2 AND2X2_1454 ( .A(u2__abc_52155_new_n4977_), .B(u2_remHi_166_), .Y(u2__abc_52155_new_n4978_));
AND2X2 AND2X2_1455 ( .A(u2__abc_52155_new_n4980_), .B(sqrto_166_), .Y(u2__abc_52155_new_n4981_));
AND2X2 AND2X2_1456 ( .A(u2__abc_52155_new_n4979_), .B(u2__abc_52155_new_n4982_), .Y(u2__abc_52155_new_n4983_));
AND2X2 AND2X2_1457 ( .A(u2__abc_52155_new_n4976_), .B(u2__abc_52155_new_n4983_), .Y(u2__abc_52155_new_n4984_));
AND2X2 AND2X2_1458 ( .A(u2__abc_52155_new_n4969_), .B(u2__abc_52155_new_n4984_), .Y(u2__abc_52155_new_n4985_));
AND2X2 AND2X2_1459 ( .A(u2__abc_52155_new_n4954_), .B(u2__abc_52155_new_n4985_), .Y(u2__abc_52155_new_n4986_));
AND2X2 AND2X2_146 ( .A(_abc_73687_new_n1038_), .B(_abc_73687_new_n1037_), .Y(\o[181] ));
AND2X2 AND2X2_1460 ( .A(u2__abc_52155_new_n4987_), .B(u2_remHi_160_), .Y(u2__abc_52155_new_n4988_));
AND2X2 AND2X2_1461 ( .A(u2__abc_52155_new_n4989_), .B(sqrto_160_), .Y(u2__abc_52155_new_n4990_));
AND2X2 AND2X2_1462 ( .A(u2__abc_52155_new_n4992_), .B(u2_remHi_161_), .Y(u2__abc_52155_new_n4993_));
AND2X2 AND2X2_1463 ( .A(u2__abc_52155_new_n4994_), .B(sqrto_161_), .Y(u2__abc_52155_new_n4995_));
AND2X2 AND2X2_1464 ( .A(u2__abc_52155_new_n4999_), .B(u2_remHi_159_), .Y(u2__abc_52155_new_n5000_));
AND2X2 AND2X2_1465 ( .A(u2__abc_52155_new_n5002_), .B(sqrto_159_), .Y(u2__abc_52155_new_n5003_));
AND2X2 AND2X2_1466 ( .A(u2__abc_52155_new_n5001_), .B(u2__abc_52155_new_n5004_), .Y(u2__abc_52155_new_n5005_));
AND2X2 AND2X2_1467 ( .A(u2__abc_52155_new_n5006_), .B(u2_remHi_158_), .Y(u2__abc_52155_new_n5007_));
AND2X2 AND2X2_1468 ( .A(u2__abc_52155_new_n5009_), .B(sqrto_158_), .Y(u2__abc_52155_new_n5010_));
AND2X2 AND2X2_1469 ( .A(u2__abc_52155_new_n5008_), .B(u2__abc_52155_new_n5011_), .Y(u2__abc_52155_new_n5012_));
AND2X2 AND2X2_147 ( .A(_abc_73687_new_n1041_), .B(_abc_73687_new_n1040_), .Y(\o[182] ));
AND2X2 AND2X2_1470 ( .A(u2__abc_52155_new_n5005_), .B(u2__abc_52155_new_n5012_), .Y(u2__abc_52155_new_n5013_));
AND2X2 AND2X2_1471 ( .A(u2__abc_52155_new_n4998_), .B(u2__abc_52155_new_n5013_), .Y(u2__abc_52155_new_n5014_));
AND2X2 AND2X2_1472 ( .A(u2__abc_52155_new_n5015_), .B(u2_remHi_164_), .Y(u2__abc_52155_new_n5016_));
AND2X2 AND2X2_1473 ( .A(u2__abc_52155_new_n5018_), .B(sqrto_164_), .Y(u2__abc_52155_new_n5019_));
AND2X2 AND2X2_1474 ( .A(u2__abc_52155_new_n5017_), .B(u2__abc_52155_new_n5020_), .Y(u2__abc_52155_new_n5021_));
AND2X2 AND2X2_1475 ( .A(u2__abc_52155_new_n5022_), .B(u2_remHi_165_), .Y(u2__abc_52155_new_n5023_));
AND2X2 AND2X2_1476 ( .A(u2__abc_52155_new_n5025_), .B(sqrto_165_), .Y(u2__abc_52155_new_n5026_));
AND2X2 AND2X2_1477 ( .A(u2__abc_52155_new_n5024_), .B(u2__abc_52155_new_n5027_), .Y(u2__abc_52155_new_n5028_));
AND2X2 AND2X2_1478 ( .A(u2__abc_52155_new_n5021_), .B(u2__abc_52155_new_n5028_), .Y(u2__abc_52155_new_n5029_));
AND2X2 AND2X2_1479 ( .A(u2__abc_52155_new_n5030_), .B(u2_remHi_163_), .Y(u2__abc_52155_new_n5031_));
AND2X2 AND2X2_148 ( .A(_abc_73687_new_n1044_), .B(_abc_73687_new_n1043_), .Y(\o[183] ));
AND2X2 AND2X2_1480 ( .A(u2__abc_52155_new_n5033_), .B(sqrto_163_), .Y(u2__abc_52155_new_n5034_));
AND2X2 AND2X2_1481 ( .A(u2__abc_52155_new_n5032_), .B(u2__abc_52155_new_n5035_), .Y(u2__abc_52155_new_n5036_));
AND2X2 AND2X2_1482 ( .A(u2__abc_52155_new_n5037_), .B(u2_remHi_162_), .Y(u2__abc_52155_new_n5038_));
AND2X2 AND2X2_1483 ( .A(u2__abc_52155_new_n5040_), .B(sqrto_162_), .Y(u2__abc_52155_new_n5041_));
AND2X2 AND2X2_1484 ( .A(u2__abc_52155_new_n5039_), .B(u2__abc_52155_new_n5042_), .Y(u2__abc_52155_new_n5043_));
AND2X2 AND2X2_1485 ( .A(u2__abc_52155_new_n5036_), .B(u2__abc_52155_new_n5043_), .Y(u2__abc_52155_new_n5044_));
AND2X2 AND2X2_1486 ( .A(u2__abc_52155_new_n5029_), .B(u2__abc_52155_new_n5044_), .Y(u2__abc_52155_new_n5045_));
AND2X2 AND2X2_1487 ( .A(u2__abc_52155_new_n5014_), .B(u2__abc_52155_new_n5045_), .Y(u2__abc_52155_new_n5046_));
AND2X2 AND2X2_1488 ( .A(u2__abc_52155_new_n5046_), .B(u2__abc_52155_new_n4986_), .Y(u2__abc_52155_new_n5047_));
AND2X2 AND2X2_1489 ( .A(u2__abc_52155_new_n5047_), .B(u2__abc_52155_new_n4923_), .Y(u2__abc_52155_new_n5048_));
AND2X2 AND2X2_149 ( .A(_abc_73687_new_n1047_), .B(_abc_73687_new_n1046_), .Y(\o[184] ));
AND2X2 AND2X2_1490 ( .A(u2__abc_52155_new_n5049_), .B(u2_remHi_152_), .Y(u2__abc_52155_new_n5050_));
AND2X2 AND2X2_1491 ( .A(u2__abc_52155_new_n5052_), .B(sqrto_152_), .Y(u2__abc_52155_new_n5053_));
AND2X2 AND2X2_1492 ( .A(u2__abc_52155_new_n5051_), .B(u2__abc_52155_new_n5054_), .Y(u2__abc_52155_new_n5055_));
AND2X2 AND2X2_1493 ( .A(u2__abc_52155_new_n5056_), .B(u2_remHi_153_), .Y(u2__abc_52155_new_n5057_));
AND2X2 AND2X2_1494 ( .A(u2__abc_52155_new_n5059_), .B(sqrto_153_), .Y(u2__abc_52155_new_n5060_));
AND2X2 AND2X2_1495 ( .A(u2__abc_52155_new_n5058_), .B(u2__abc_52155_new_n5061_), .Y(u2__abc_52155_new_n5062_));
AND2X2 AND2X2_1496 ( .A(u2__abc_52155_new_n5055_), .B(u2__abc_52155_new_n5062_), .Y(u2__abc_52155_new_n5063_));
AND2X2 AND2X2_1497 ( .A(u2__abc_52155_new_n5064_), .B(u2_remHi_151_), .Y(u2__abc_52155_new_n5065_));
AND2X2 AND2X2_1498 ( .A(u2__abc_52155_new_n5067_), .B(sqrto_151_), .Y(u2__abc_52155_new_n5068_));
AND2X2 AND2X2_1499 ( .A(u2__abc_52155_new_n5066_), .B(u2__abc_52155_new_n5069_), .Y(u2__abc_52155_new_n5070_));
AND2X2 AND2X2_15 ( .A(_abc_73687_new_n753_), .B(sqrto_14_), .Y(\o[50] ));
AND2X2 AND2X2_150 ( .A(_abc_73687_new_n1050_), .B(_abc_73687_new_n1049_), .Y(\o[185] ));
AND2X2 AND2X2_1500 ( .A(u2__abc_52155_new_n5071_), .B(u2_remHi_150_), .Y(u2__abc_52155_new_n5072_));
AND2X2 AND2X2_1501 ( .A(u2__abc_52155_new_n5074_), .B(sqrto_150_), .Y(u2__abc_52155_new_n5075_));
AND2X2 AND2X2_1502 ( .A(u2__abc_52155_new_n5073_), .B(u2__abc_52155_new_n5076_), .Y(u2__abc_52155_new_n5077_));
AND2X2 AND2X2_1503 ( .A(u2__abc_52155_new_n5070_), .B(u2__abc_52155_new_n5077_), .Y(u2__abc_52155_new_n5078_));
AND2X2 AND2X2_1504 ( .A(u2__abc_52155_new_n5063_), .B(u2__abc_52155_new_n5078_), .Y(u2__abc_52155_new_n5079_));
AND2X2 AND2X2_1505 ( .A(u2__abc_52155_new_n5080_), .B(u2_remHi_156_), .Y(u2__abc_52155_new_n5081_));
AND2X2 AND2X2_1506 ( .A(u2__abc_52155_new_n5083_), .B(sqrto_156_), .Y(u2__abc_52155_new_n5084_));
AND2X2 AND2X2_1507 ( .A(u2__abc_52155_new_n5082_), .B(u2__abc_52155_new_n5085_), .Y(u2__abc_52155_new_n5086_));
AND2X2 AND2X2_1508 ( .A(u2__abc_52155_new_n5087_), .B(u2_remHi_157_), .Y(u2__abc_52155_new_n5088_));
AND2X2 AND2X2_1509 ( .A(u2__abc_52155_new_n5090_), .B(sqrto_157_), .Y(u2__abc_52155_new_n5091_));
AND2X2 AND2X2_151 ( .A(_abc_73687_new_n1053_), .B(_abc_73687_new_n1052_), .Y(\o[186] ));
AND2X2 AND2X2_1510 ( .A(u2__abc_52155_new_n5089_), .B(u2__abc_52155_new_n5092_), .Y(u2__abc_52155_new_n5093_));
AND2X2 AND2X2_1511 ( .A(u2__abc_52155_new_n5086_), .B(u2__abc_52155_new_n5093_), .Y(u2__abc_52155_new_n5094_));
AND2X2 AND2X2_1512 ( .A(u2__abc_52155_new_n5095_), .B(u2_remHi_155_), .Y(u2__abc_52155_new_n5096_));
AND2X2 AND2X2_1513 ( .A(u2__abc_52155_new_n5098_), .B(sqrto_155_), .Y(u2__abc_52155_new_n5099_));
AND2X2 AND2X2_1514 ( .A(u2__abc_52155_new_n5097_), .B(u2__abc_52155_new_n5100_), .Y(u2__abc_52155_new_n5101_));
AND2X2 AND2X2_1515 ( .A(u2__abc_52155_new_n5102_), .B(u2_remHi_154_), .Y(u2__abc_52155_new_n5103_));
AND2X2 AND2X2_1516 ( .A(u2__abc_52155_new_n5105_), .B(sqrto_154_), .Y(u2__abc_52155_new_n5106_));
AND2X2 AND2X2_1517 ( .A(u2__abc_52155_new_n5104_), .B(u2__abc_52155_new_n5107_), .Y(u2__abc_52155_new_n5108_));
AND2X2 AND2X2_1518 ( .A(u2__abc_52155_new_n5101_), .B(u2__abc_52155_new_n5108_), .Y(u2__abc_52155_new_n5109_));
AND2X2 AND2X2_1519 ( .A(u2__abc_52155_new_n5094_), .B(u2__abc_52155_new_n5109_), .Y(u2__abc_52155_new_n5110_));
AND2X2 AND2X2_152 ( .A(_abc_73687_new_n1056_), .B(_abc_73687_new_n1055_), .Y(\o[187] ));
AND2X2 AND2X2_1520 ( .A(u2__abc_52155_new_n5079_), .B(u2__abc_52155_new_n5110_), .Y(u2__abc_52155_new_n5111_));
AND2X2 AND2X2_1521 ( .A(u2__abc_52155_new_n5112_), .B(u2_remHi_148_), .Y(u2__abc_52155_new_n5113_));
AND2X2 AND2X2_1522 ( .A(u2__abc_52155_new_n5115_), .B(sqrto_148_), .Y(u2__abc_52155_new_n5116_));
AND2X2 AND2X2_1523 ( .A(u2__abc_52155_new_n5114_), .B(u2__abc_52155_new_n5117_), .Y(u2__abc_52155_new_n5118_));
AND2X2 AND2X2_1524 ( .A(u2__abc_52155_new_n5119_), .B(u2_remHi_149_), .Y(u2__abc_52155_new_n5120_));
AND2X2 AND2X2_1525 ( .A(u2__abc_52155_new_n5122_), .B(sqrto_149_), .Y(u2__abc_52155_new_n5123_));
AND2X2 AND2X2_1526 ( .A(u2__abc_52155_new_n5121_), .B(u2__abc_52155_new_n5124_), .Y(u2__abc_52155_new_n5125_));
AND2X2 AND2X2_1527 ( .A(u2__abc_52155_new_n5118_), .B(u2__abc_52155_new_n5125_), .Y(u2__abc_52155_new_n5126_));
AND2X2 AND2X2_1528 ( .A(u2__abc_52155_new_n5127_), .B(u2_remHi_147_), .Y(u2__abc_52155_new_n5128_));
AND2X2 AND2X2_1529 ( .A(u2__abc_52155_new_n5130_), .B(sqrto_147_), .Y(u2__abc_52155_new_n5131_));
AND2X2 AND2X2_153 ( .A(_abc_73687_new_n1059_), .B(_abc_73687_new_n1058_), .Y(\o[188] ));
AND2X2 AND2X2_1530 ( .A(u2__abc_52155_new_n5129_), .B(u2__abc_52155_new_n5132_), .Y(u2__abc_52155_new_n5133_));
AND2X2 AND2X2_1531 ( .A(u2__abc_52155_new_n5134_), .B(u2_remHi_146_), .Y(u2__abc_52155_new_n5135_));
AND2X2 AND2X2_1532 ( .A(u2__abc_52155_new_n5137_), .B(sqrto_146_), .Y(u2__abc_52155_new_n5138_));
AND2X2 AND2X2_1533 ( .A(u2__abc_52155_new_n5136_), .B(u2__abc_52155_new_n5139_), .Y(u2__abc_52155_new_n5140_));
AND2X2 AND2X2_1534 ( .A(u2__abc_52155_new_n5133_), .B(u2__abc_52155_new_n5140_), .Y(u2__abc_52155_new_n5141_));
AND2X2 AND2X2_1535 ( .A(u2__abc_52155_new_n5126_), .B(u2__abc_52155_new_n5141_), .Y(u2__abc_52155_new_n5142_));
AND2X2 AND2X2_1536 ( .A(u2__abc_52155_new_n5143_), .B(u2_remHi_144_), .Y(u2__abc_52155_new_n5144_));
AND2X2 AND2X2_1537 ( .A(u2__abc_52155_new_n5145_), .B(sqrto_144_), .Y(u2__abc_52155_new_n5146_));
AND2X2 AND2X2_1538 ( .A(u2__abc_52155_new_n5148_), .B(u2_remHi_145_), .Y(u2__abc_52155_new_n5149_));
AND2X2 AND2X2_1539 ( .A(u2__abc_52155_new_n5150_), .B(sqrto_145_), .Y(u2__abc_52155_new_n5151_));
AND2X2 AND2X2_154 ( .A(_abc_73687_new_n1062_), .B(_abc_73687_new_n1061_), .Y(\o[189] ));
AND2X2 AND2X2_1540 ( .A(u2__abc_52155_new_n5155_), .B(u2_remHi_143_), .Y(u2__abc_52155_new_n5156_));
AND2X2 AND2X2_1541 ( .A(u2__abc_52155_new_n5158_), .B(sqrto_143_), .Y(u2__abc_52155_new_n5159_));
AND2X2 AND2X2_1542 ( .A(u2__abc_52155_new_n5157_), .B(u2__abc_52155_new_n5160_), .Y(u2__abc_52155_new_n5161_));
AND2X2 AND2X2_1543 ( .A(u2__abc_52155_new_n5162_), .B(u2_remHi_142_), .Y(u2__abc_52155_new_n5163_));
AND2X2 AND2X2_1544 ( .A(u2__abc_52155_new_n5165_), .B(sqrto_142_), .Y(u2__abc_52155_new_n5166_));
AND2X2 AND2X2_1545 ( .A(u2__abc_52155_new_n5164_), .B(u2__abc_52155_new_n5167_), .Y(u2__abc_52155_new_n5168_));
AND2X2 AND2X2_1546 ( .A(u2__abc_52155_new_n5161_), .B(u2__abc_52155_new_n5168_), .Y(u2__abc_52155_new_n5169_));
AND2X2 AND2X2_1547 ( .A(u2__abc_52155_new_n5154_), .B(u2__abc_52155_new_n5169_), .Y(u2__abc_52155_new_n5170_));
AND2X2 AND2X2_1548 ( .A(u2__abc_52155_new_n5170_), .B(u2__abc_52155_new_n5142_), .Y(u2__abc_52155_new_n5171_));
AND2X2 AND2X2_1549 ( .A(u2__abc_52155_new_n5171_), .B(u2__abc_52155_new_n5111_), .Y(u2__abc_52155_new_n5172_));
AND2X2 AND2X2_155 ( .A(_abc_73687_new_n1065_), .B(_abc_73687_new_n1064_), .Y(\o[190] ));
AND2X2 AND2X2_1550 ( .A(u2__abc_52155_new_n5173_), .B(u2_remHi_136_), .Y(u2__abc_52155_new_n5174_));
AND2X2 AND2X2_1551 ( .A(u2__abc_52155_new_n5175_), .B(sqrto_136_), .Y(u2__abc_52155_new_n5176_));
AND2X2 AND2X2_1552 ( .A(u2__abc_52155_new_n5178_), .B(u2_remHi_137_), .Y(u2__abc_52155_new_n5179_));
AND2X2 AND2X2_1553 ( .A(u2__abc_52155_new_n5180_), .B(sqrto_137_), .Y(u2__abc_52155_new_n5181_));
AND2X2 AND2X2_1554 ( .A(u2__abc_52155_new_n5185_), .B(u2_remHi_134_), .Y(u2__abc_52155_new_n5186_));
AND2X2 AND2X2_1555 ( .A(u2__abc_52155_new_n5188_), .B(sqrto_134_), .Y(u2__abc_52155_new_n5189_));
AND2X2 AND2X2_1556 ( .A(u2__abc_52155_new_n5187_), .B(u2__abc_52155_new_n5190_), .Y(u2__abc_52155_new_n5191_));
AND2X2 AND2X2_1557 ( .A(u2__abc_52155_new_n5192_), .B(u2_remHi_135_), .Y(u2__abc_52155_new_n5193_));
AND2X2 AND2X2_1558 ( .A(u2__abc_52155_new_n5195_), .B(sqrto_135_), .Y(u2__abc_52155_new_n5196_));
AND2X2 AND2X2_1559 ( .A(u2__abc_52155_new_n5194_), .B(u2__abc_52155_new_n5197_), .Y(u2__abc_52155_new_n5198_));
AND2X2 AND2X2_156 ( .A(_abc_73687_new_n1068_), .B(_abc_73687_new_n1067_), .Y(\o[191] ));
AND2X2 AND2X2_1560 ( .A(u2__abc_52155_new_n5191_), .B(u2__abc_52155_new_n5198_), .Y(u2__abc_52155_new_n5199_));
AND2X2 AND2X2_1561 ( .A(u2__abc_52155_new_n5184_), .B(u2__abc_52155_new_n5199_), .Y(u2__abc_52155_new_n5200_));
AND2X2 AND2X2_1562 ( .A(u2__abc_52155_new_n5201_), .B(u2_remHi_140_), .Y(u2__abc_52155_new_n5202_));
AND2X2 AND2X2_1563 ( .A(u2__abc_52155_new_n5204_), .B(sqrto_140_), .Y(u2__abc_52155_new_n5205_));
AND2X2 AND2X2_1564 ( .A(u2__abc_52155_new_n5203_), .B(u2__abc_52155_new_n5206_), .Y(u2__abc_52155_new_n5207_));
AND2X2 AND2X2_1565 ( .A(u2__abc_52155_new_n5208_), .B(u2_remHi_141_), .Y(u2__abc_52155_new_n5209_));
AND2X2 AND2X2_1566 ( .A(u2__abc_52155_new_n5211_), .B(sqrto_141_), .Y(u2__abc_52155_new_n5212_));
AND2X2 AND2X2_1567 ( .A(u2__abc_52155_new_n5210_), .B(u2__abc_52155_new_n5213_), .Y(u2__abc_52155_new_n5214_));
AND2X2 AND2X2_1568 ( .A(u2__abc_52155_new_n5207_), .B(u2__abc_52155_new_n5214_), .Y(u2__abc_52155_new_n5215_));
AND2X2 AND2X2_1569 ( .A(u2__abc_52155_new_n5216_), .B(u2_remHi_139_), .Y(u2__abc_52155_new_n5217_));
AND2X2 AND2X2_157 ( .A(_abc_73687_new_n1071_), .B(_abc_73687_new_n1070_), .Y(\o[192] ));
AND2X2 AND2X2_1570 ( .A(u2__abc_52155_new_n5219_), .B(sqrto_139_), .Y(u2__abc_52155_new_n5220_));
AND2X2 AND2X2_1571 ( .A(u2__abc_52155_new_n5218_), .B(u2__abc_52155_new_n5221_), .Y(u2__abc_52155_new_n5222_));
AND2X2 AND2X2_1572 ( .A(u2__abc_52155_new_n5223_), .B(u2_remHi_138_), .Y(u2__abc_52155_new_n5224_));
AND2X2 AND2X2_1573 ( .A(u2__abc_52155_new_n5226_), .B(sqrto_138_), .Y(u2__abc_52155_new_n5227_));
AND2X2 AND2X2_1574 ( .A(u2__abc_52155_new_n5225_), .B(u2__abc_52155_new_n5228_), .Y(u2__abc_52155_new_n5229_));
AND2X2 AND2X2_1575 ( .A(u2__abc_52155_new_n5222_), .B(u2__abc_52155_new_n5229_), .Y(u2__abc_52155_new_n5230_));
AND2X2 AND2X2_1576 ( .A(u2__abc_52155_new_n5215_), .B(u2__abc_52155_new_n5230_), .Y(u2__abc_52155_new_n5231_));
AND2X2 AND2X2_1577 ( .A(u2__abc_52155_new_n5200_), .B(u2__abc_52155_new_n5231_), .Y(u2__abc_52155_new_n5232_));
AND2X2 AND2X2_1578 ( .A(u2__abc_52155_new_n5233_), .B(u2_remHi_126_), .Y(u2__abc_52155_new_n5234_));
AND2X2 AND2X2_1579 ( .A(u2__abc_52155_new_n5235_), .B(u2__abc_52155_new_n5236_), .Y(u2__abc_52155_new_n5237_));
AND2X2 AND2X2_158 ( .A(_abc_73687_new_n1074_), .B(_abc_73687_new_n1073_), .Y(\o[193] ));
AND2X2 AND2X2_1580 ( .A(u2__abc_52155_new_n5238_), .B(u2_remHi_127_), .Y(u2__abc_52155_new_n5239_));
AND2X2 AND2X2_1581 ( .A(u2__abc_52155_new_n5241_), .B(sqrto_127_), .Y(u2__abc_52155_new_n5242_));
AND2X2 AND2X2_1582 ( .A(u2__abc_52155_new_n5240_), .B(u2__abc_52155_new_n5243_), .Y(u2__abc_52155_new_n5244_));
AND2X2 AND2X2_1583 ( .A(u2__abc_52155_new_n5244_), .B(u2__abc_52155_new_n5237_), .Y(u2__abc_52155_new_n5245_));
AND2X2 AND2X2_1584 ( .A(u2__abc_52155_new_n5246_), .B(u2_remHi_128_), .Y(u2__abc_52155_new_n5247_));
AND2X2 AND2X2_1585 ( .A(u2__abc_52155_new_n5248_), .B(sqrto_128_), .Y(u2__abc_52155_new_n5249_));
AND2X2 AND2X2_1586 ( .A(u2__abc_52155_new_n5251_), .B(u2_remHi_129_), .Y(u2__abc_52155_new_n5252_));
AND2X2 AND2X2_1587 ( .A(u2__abc_52155_new_n5253_), .B(sqrto_129_), .Y(u2__abc_52155_new_n5254_));
AND2X2 AND2X2_1588 ( .A(u2__abc_52155_new_n5257_), .B(u2__abc_52155_new_n5245_), .Y(u2__abc_52155_new_n5258_));
AND2X2 AND2X2_1589 ( .A(u2__abc_52155_new_n5259_), .B(u2_remHi_132_), .Y(u2__abc_52155_new_n5260_));
AND2X2 AND2X2_159 ( .A(_abc_73687_new_n1077_), .B(_abc_73687_new_n1076_), .Y(\o[194] ));
AND2X2 AND2X2_1590 ( .A(u2__abc_52155_new_n5261_), .B(sqrto_132_), .Y(u2__abc_52155_new_n5262_));
AND2X2 AND2X2_1591 ( .A(u2__abc_52155_new_n5264_), .B(u2_remHi_133_), .Y(u2__abc_52155_new_n5265_));
AND2X2 AND2X2_1592 ( .A(u2__abc_52155_new_n5266_), .B(sqrto_133_), .Y(u2__abc_52155_new_n5267_));
AND2X2 AND2X2_1593 ( .A(u2__abc_52155_new_n5270_), .B(u2_remHi_131_), .Y(u2__abc_52155_new_n5271_));
AND2X2 AND2X2_1594 ( .A(u2__abc_52155_new_n5272_), .B(sqrto_131_), .Y(u2__abc_52155_new_n5273_));
AND2X2 AND2X2_1595 ( .A(u2__abc_52155_new_n5275_), .B(u2_remHi_130_), .Y(u2__abc_52155_new_n5276_));
AND2X2 AND2X2_1596 ( .A(u2__abc_52155_new_n5277_), .B(sqrto_130_), .Y(u2__abc_52155_new_n5278_));
AND2X2 AND2X2_1597 ( .A(u2__abc_52155_new_n5282_), .B(u2__abc_52155_new_n5258_), .Y(u2__abc_52155_new_n5283_));
AND2X2 AND2X2_1598 ( .A(u2__abc_52155_new_n5283_), .B(u2__abc_52155_new_n5232_), .Y(u2__abc_52155_new_n5284_));
AND2X2 AND2X2_1599 ( .A(u2__abc_52155_new_n5284_), .B(u2__abc_52155_new_n5172_), .Y(u2__abc_52155_new_n5285_));
AND2X2 AND2X2_16 ( .A(_abc_73687_new_n753_), .B(sqrto_15_), .Y(\o[51] ));
AND2X2 AND2X2_160 ( .A(_abc_73687_new_n1080_), .B(_abc_73687_new_n1079_), .Y(\o[195] ));
AND2X2 AND2X2_1600 ( .A(u2__abc_52155_new_n5285_), .B(u2__abc_52155_new_n5048_), .Y(u2__abc_52155_new_n5286_));
AND2X2 AND2X2_1601 ( .A(u2__abc_52155_new_n5286_), .B(u2__abc_52155_new_n4796_), .Y(u2__abc_52155_new_n5287_));
AND2X2 AND2X2_1602 ( .A(u2__abc_52155_new_n5294_), .B(u2__abc_52155_new_n5243_), .Y(u2__abc_52155_new_n5295_));
AND2X2 AND2X2_1603 ( .A(u2__abc_52155_new_n5299_), .B(u2__abc_52155_new_n5297_), .Y(u2__abc_52155_new_n5300_));
AND2X2 AND2X2_1604 ( .A(u2__abc_52155_new_n5296_), .B(u2__abc_52155_new_n5300_), .Y(u2__abc_52155_new_n5301_));
AND2X2 AND2X2_1605 ( .A(u2__abc_52155_new_n5305_), .B(u2__abc_52155_new_n5303_), .Y(u2__abc_52155_new_n5306_));
AND2X2 AND2X2_1606 ( .A(u2__abc_52155_new_n5308_), .B(u2__abc_52155_new_n5262_), .Y(u2__abc_52155_new_n5309_));
AND2X2 AND2X2_1607 ( .A(u2__abc_52155_new_n5307_), .B(u2__abc_52155_new_n5311_), .Y(u2__abc_52155_new_n5312_));
AND2X2 AND2X2_1608 ( .A(u2__abc_52155_new_n5302_), .B(u2__abc_52155_new_n5312_), .Y(u2__abc_52155_new_n5313_));
AND2X2 AND2X2_1609 ( .A(u2__abc_52155_new_n5316_), .B(u2__abc_52155_new_n5197_), .Y(u2__abc_52155_new_n5317_));
AND2X2 AND2X2_161 ( .A(_abc_73687_new_n1083_), .B(_abc_73687_new_n1082_), .Y(\o[196] ));
AND2X2 AND2X2_1610 ( .A(u2__abc_52155_new_n5319_), .B(u2__abc_52155_new_n5176_), .Y(u2__abc_52155_new_n5320_));
AND2X2 AND2X2_1611 ( .A(u2__abc_52155_new_n5318_), .B(u2__abc_52155_new_n5322_), .Y(u2__abc_52155_new_n5323_));
AND2X2 AND2X2_1612 ( .A(u2__abc_52155_new_n5218_), .B(u2__abc_52155_new_n5227_), .Y(u2__abc_52155_new_n5325_));
AND2X2 AND2X2_1613 ( .A(u2__abc_52155_new_n5326_), .B(u2__abc_52155_new_n5215_), .Y(u2__abc_52155_new_n5327_));
AND2X2 AND2X2_1614 ( .A(u2__abc_52155_new_n5210_), .B(u2__abc_52155_new_n5205_), .Y(u2__abc_52155_new_n5328_));
AND2X2 AND2X2_1615 ( .A(u2__abc_52155_new_n5324_), .B(u2__abc_52155_new_n5331_), .Y(u2__abc_52155_new_n5332_));
AND2X2 AND2X2_1616 ( .A(u2__abc_52155_new_n5314_), .B(u2__abc_52155_new_n5332_), .Y(u2__abc_52155_new_n5333_));
AND2X2 AND2X2_1617 ( .A(u2__abc_52155_new_n5337_), .B(u2__abc_52155_new_n5160_), .Y(u2__abc_52155_new_n5338_));
AND2X2 AND2X2_1618 ( .A(u2__abc_52155_new_n5340_), .B(u2__abc_52155_new_n5146_), .Y(u2__abc_52155_new_n5341_));
AND2X2 AND2X2_1619 ( .A(u2__abc_52155_new_n5339_), .B(u2__abc_52155_new_n5343_), .Y(u2__abc_52155_new_n5344_));
AND2X2 AND2X2_162 ( .A(_abc_73687_new_n1086_), .B(_abc_73687_new_n1085_), .Y(\o[197] ));
AND2X2 AND2X2_1620 ( .A(u2__abc_52155_new_n5129_), .B(u2__abc_52155_new_n5138_), .Y(u2__abc_52155_new_n5346_));
AND2X2 AND2X2_1621 ( .A(u2__abc_52155_new_n5347_), .B(u2__abc_52155_new_n5126_), .Y(u2__abc_52155_new_n5348_));
AND2X2 AND2X2_1622 ( .A(u2__abc_52155_new_n5121_), .B(u2__abc_52155_new_n5116_), .Y(u2__abc_52155_new_n5349_));
AND2X2 AND2X2_1623 ( .A(u2__abc_52155_new_n5345_), .B(u2__abc_52155_new_n5352_), .Y(u2__abc_52155_new_n5353_));
AND2X2 AND2X2_1624 ( .A(u2__abc_52155_new_n5066_), .B(u2__abc_52155_new_n5075_), .Y(u2__abc_52155_new_n5355_));
AND2X2 AND2X2_1625 ( .A(u2__abc_52155_new_n5356_), .B(u2__abc_52155_new_n5063_), .Y(u2__abc_52155_new_n5357_));
AND2X2 AND2X2_1626 ( .A(u2__abc_52155_new_n5058_), .B(u2__abc_52155_new_n5053_), .Y(u2__abc_52155_new_n5358_));
AND2X2 AND2X2_1627 ( .A(u2__abc_52155_new_n5360_), .B(u2__abc_52155_new_n5110_), .Y(u2__abc_52155_new_n5361_));
AND2X2 AND2X2_1628 ( .A(u2__abc_52155_new_n5097_), .B(u2__abc_52155_new_n5106_), .Y(u2__abc_52155_new_n5362_));
AND2X2 AND2X2_1629 ( .A(u2__abc_52155_new_n5363_), .B(u2__abc_52155_new_n5094_), .Y(u2__abc_52155_new_n5364_));
AND2X2 AND2X2_163 ( .A(_abc_73687_new_n1089_), .B(_abc_73687_new_n1088_), .Y(\o[198] ));
AND2X2 AND2X2_1630 ( .A(u2__abc_52155_new_n5089_), .B(u2__abc_52155_new_n5084_), .Y(u2__abc_52155_new_n5365_));
AND2X2 AND2X2_1631 ( .A(u2__abc_52155_new_n5354_), .B(u2__abc_52155_new_n5369_), .Y(u2__abc_52155_new_n5370_));
AND2X2 AND2X2_1632 ( .A(u2__abc_52155_new_n5334_), .B(u2__abc_52155_new_n5370_), .Y(u2__abc_52155_new_n5371_));
AND2X2 AND2X2_1633 ( .A(u2__abc_52155_new_n5376_), .B(u2__abc_52155_new_n5004_), .Y(u2__abc_52155_new_n5377_));
AND2X2 AND2X2_1634 ( .A(u2__abc_52155_new_n5379_), .B(u2__abc_52155_new_n4990_), .Y(u2__abc_52155_new_n5380_));
AND2X2 AND2X2_1635 ( .A(u2__abc_52155_new_n5378_), .B(u2__abc_52155_new_n5382_), .Y(u2__abc_52155_new_n5383_));
AND2X2 AND2X2_1636 ( .A(u2__abc_52155_new_n5032_), .B(u2__abc_52155_new_n5041_), .Y(u2__abc_52155_new_n5385_));
AND2X2 AND2X2_1637 ( .A(u2__abc_52155_new_n5386_), .B(u2__abc_52155_new_n5029_), .Y(u2__abc_52155_new_n5387_));
AND2X2 AND2X2_1638 ( .A(u2__abc_52155_new_n5024_), .B(u2__abc_52155_new_n5019_), .Y(u2__abc_52155_new_n5388_));
AND2X2 AND2X2_1639 ( .A(u2__abc_52155_new_n5384_), .B(u2__abc_52155_new_n5391_), .Y(u2__abc_52155_new_n5392_));
AND2X2 AND2X2_164 ( .A(_abc_73687_new_n1092_), .B(_abc_73687_new_n1091_), .Y(\o[199] ));
AND2X2 AND2X2_1640 ( .A(u2__abc_52155_new_n4972_), .B(u2__abc_52155_new_n4981_), .Y(u2__abc_52155_new_n5394_));
AND2X2 AND2X2_1641 ( .A(u2__abc_52155_new_n5395_), .B(u2__abc_52155_new_n4969_), .Y(u2__abc_52155_new_n5396_));
AND2X2 AND2X2_1642 ( .A(u2__abc_52155_new_n4964_), .B(u2__abc_52155_new_n4959_), .Y(u2__abc_52155_new_n5397_));
AND2X2 AND2X2_1643 ( .A(u2__abc_52155_new_n5399_), .B(u2__abc_52155_new_n4954_), .Y(u2__abc_52155_new_n5400_));
AND2X2 AND2X2_1644 ( .A(u2__abc_52155_new_n4941_), .B(u2__abc_52155_new_n4950_), .Y(u2__abc_52155_new_n5401_));
AND2X2 AND2X2_1645 ( .A(u2__abc_52155_new_n5402_), .B(u2__abc_52155_new_n4938_), .Y(u2__abc_52155_new_n5403_));
AND2X2 AND2X2_1646 ( .A(u2__abc_52155_new_n4933_), .B(u2__abc_52155_new_n4928_), .Y(u2__abc_52155_new_n5404_));
AND2X2 AND2X2_1647 ( .A(u2__abc_52155_new_n5393_), .B(u2__abc_52155_new_n5408_), .Y(u2__abc_52155_new_n5409_));
AND2X2 AND2X2_1648 ( .A(u2__abc_52155_new_n4915_), .B(u2__abc_52155_new_n4910_), .Y(u2__abc_52155_new_n5411_));
AND2X2 AND2X2_1649 ( .A(u2__abc_52155_new_n5412_), .B(u2__abc_52155_new_n4905_), .Y(u2__abc_52155_new_n5413_));
AND2X2 AND2X2_165 ( .A(_abc_73687_new_n1095_), .B(_abc_73687_new_n1094_), .Y(\o[200] ));
AND2X2 AND2X2_1650 ( .A(u2__abc_52155_new_n4900_), .B(u2__abc_52155_new_n4895_), .Y(u2__abc_52155_new_n5414_));
AND2X2 AND2X2_1651 ( .A(u2__abc_52155_new_n5416_), .B(u2__abc_52155_new_n4890_), .Y(u2__abc_52155_new_n5417_));
AND2X2 AND2X2_1652 ( .A(u2__abc_52155_new_n4869_), .B(u2__abc_52155_new_n4864_), .Y(u2__abc_52155_new_n5418_));
AND2X2 AND2X2_1653 ( .A(u2__abc_52155_new_n4877_), .B(u2__abc_52155_new_n4886_), .Y(u2__abc_52155_new_n5420_));
AND2X2 AND2X2_1654 ( .A(u2__abc_52155_new_n5421_), .B(u2__abc_52155_new_n4874_), .Y(u2__abc_52155_new_n5422_));
AND2X2 AND2X2_1655 ( .A(u2__abc_52155_new_n5424_), .B(u2__abc_52155_new_n4859_), .Y(u2__abc_52155_new_n5425_));
AND2X2 AND2X2_1656 ( .A(u2__abc_52155_new_n4806_), .B(u2__abc_52155_new_n4801_), .Y(u2__abc_52155_new_n5426_));
AND2X2 AND2X2_1657 ( .A(u2__abc_52155_new_n5427_), .B(u2__abc_52155_new_n4826_), .Y(u2__abc_52155_new_n5428_));
AND2X2 AND2X2_1658 ( .A(u2__abc_52155_new_n4821_), .B(u2__abc_52155_new_n4816_), .Y(u2__abc_52155_new_n5429_));
AND2X2 AND2X2_1659 ( .A(u2__abc_52155_new_n5431_), .B(u2__abc_52155_new_n4858_), .Y(u2__abc_52155_new_n5432_));
AND2X2 AND2X2_166 ( .A(_abc_73687_new_n1098_), .B(_abc_73687_new_n1097_), .Y(\o[201] ));
AND2X2 AND2X2_1660 ( .A(u2__abc_52155_new_n4845_), .B(u2__abc_52155_new_n4854_), .Y(u2__abc_52155_new_n5433_));
AND2X2 AND2X2_1661 ( .A(u2__abc_52155_new_n5434_), .B(u2__abc_52155_new_n4842_), .Y(u2__abc_52155_new_n5435_));
AND2X2 AND2X2_1662 ( .A(u2__abc_52155_new_n4837_), .B(u2__abc_52155_new_n4832_), .Y(u2__abc_52155_new_n5436_));
AND2X2 AND2X2_1663 ( .A(u2__abc_52155_new_n5410_), .B(u2__abc_52155_new_n5441_), .Y(u2__abc_52155_new_n5442_));
AND2X2 AND2X2_1664 ( .A(u2__abc_52155_new_n5372_), .B(u2__abc_52155_new_n5442_), .Y(u2__abc_52155_new_n5443_));
AND2X2 AND2X2_1665 ( .A(u2__abc_52155_new_n5449_), .B(u2__abc_52155_new_n4789_), .Y(u2__abc_52155_new_n5450_));
AND2X2 AND2X2_1666 ( .A(u2__abc_52155_new_n5452_), .B(u2__abc_52155_new_n4768_), .Y(u2__abc_52155_new_n5453_));
AND2X2 AND2X2_1667 ( .A(u2__abc_52155_new_n5451_), .B(u2__abc_52155_new_n5455_), .Y(u2__abc_52155_new_n5456_));
AND2X2 AND2X2_1668 ( .A(u2__abc_52155_new_n4751_), .B(u2__abc_52155_new_n4760_), .Y(u2__abc_52155_new_n5458_));
AND2X2 AND2X2_1669 ( .A(u2__abc_52155_new_n5459_), .B(u2__abc_52155_new_n4748_), .Y(u2__abc_52155_new_n5460_));
AND2X2 AND2X2_167 ( .A(_abc_73687_new_n1101_), .B(_abc_73687_new_n1100_), .Y(\o[202] ));
AND2X2 AND2X2_1670 ( .A(u2__abc_52155_new_n4743_), .B(u2__abc_52155_new_n4738_), .Y(u2__abc_52155_new_n5461_));
AND2X2 AND2X2_1671 ( .A(u2__abc_52155_new_n5457_), .B(u2__abc_52155_new_n5464_), .Y(u2__abc_52155_new_n5465_));
AND2X2 AND2X2_1672 ( .A(u2__abc_52155_new_n4688_), .B(u2__abc_52155_new_n4697_), .Y(u2__abc_52155_new_n5467_));
AND2X2 AND2X2_1673 ( .A(u2__abc_52155_new_n5468_), .B(u2__abc_52155_new_n4685_), .Y(u2__abc_52155_new_n5469_));
AND2X2 AND2X2_1674 ( .A(u2__abc_52155_new_n4680_), .B(u2__abc_52155_new_n4675_), .Y(u2__abc_52155_new_n5470_));
AND2X2 AND2X2_1675 ( .A(u2__abc_52155_new_n5472_), .B(u2__abc_52155_new_n4732_), .Y(u2__abc_52155_new_n5473_));
AND2X2 AND2X2_1676 ( .A(u2__abc_52155_new_n4719_), .B(u2__abc_52155_new_n4728_), .Y(u2__abc_52155_new_n5474_));
AND2X2 AND2X2_1677 ( .A(u2__abc_52155_new_n5475_), .B(u2__abc_52155_new_n4716_), .Y(u2__abc_52155_new_n5476_));
AND2X2 AND2X2_1678 ( .A(u2__abc_52155_new_n4711_), .B(u2__abc_52155_new_n4706_), .Y(u2__abc_52155_new_n5477_));
AND2X2 AND2X2_1679 ( .A(u2__abc_52155_new_n5466_), .B(u2__abc_52155_new_n5481_), .Y(u2__abc_52155_new_n5482_));
AND2X2 AND2X2_168 ( .A(_abc_73687_new_n1104_), .B(_abc_73687_new_n1103_), .Y(\o[203] ));
AND2X2 AND2X2_1680 ( .A(u2__abc_52155_new_n4631_), .B(u2__abc_52155_new_n4626_), .Y(u2__abc_52155_new_n5484_));
AND2X2 AND2X2_1681 ( .A(u2__abc_52155_new_n5485_), .B(u2__abc_52155_new_n4621_), .Y(u2__abc_52155_new_n5486_));
AND2X2 AND2X2_1682 ( .A(u2__abc_52155_new_n4616_), .B(u2__abc_52155_new_n4611_), .Y(u2__abc_52155_new_n5487_));
AND2X2 AND2X2_1683 ( .A(u2__abc_52155_new_n5489_), .B(u2__abc_52155_new_n4668_), .Y(u2__abc_52155_new_n5490_));
AND2X2 AND2X2_1684 ( .A(u2__abc_52155_new_n4655_), .B(u2__abc_52155_new_n4664_), .Y(u2__abc_52155_new_n5491_));
AND2X2 AND2X2_1685 ( .A(u2__abc_52155_new_n5492_), .B(u2__abc_52155_new_n4652_), .Y(u2__abc_52155_new_n5493_));
AND2X2 AND2X2_1686 ( .A(u2__abc_52155_new_n4647_), .B(u2__abc_52155_new_n4642_), .Y(u2__abc_52155_new_n5494_));
AND2X2 AND2X2_1687 ( .A(u2__abc_52155_new_n5497_), .B(u2__abc_52155_new_n4606_), .Y(u2__abc_52155_new_n5498_));
AND2X2 AND2X2_1688 ( .A(u2__abc_52155_new_n4568_), .B(u2__abc_52155_new_n4563_), .Y(u2__abc_52155_new_n5499_));
AND2X2 AND2X2_1689 ( .A(u2__abc_52155_new_n5500_), .B(u2__abc_52155_new_n4558_), .Y(u2__abc_52155_new_n5501_));
AND2X2 AND2X2_169 ( .A(_abc_73687_new_n1107_), .B(_abc_73687_new_n1106_), .Y(\o[204] ));
AND2X2 AND2X2_1690 ( .A(u2__abc_52155_new_n4553_), .B(u2__abc_52155_new_n4548_), .Y(u2__abc_52155_new_n5502_));
AND2X2 AND2X2_1691 ( .A(u2__abc_52155_new_n5504_), .B(u2__abc_52155_new_n4605_), .Y(u2__abc_52155_new_n5505_));
AND2X2 AND2X2_1692 ( .A(u2__abc_52155_new_n4584_), .B(u2__abc_52155_new_n4579_), .Y(u2__abc_52155_new_n5506_));
AND2X2 AND2X2_1693 ( .A(u2__abc_52155_new_n4592_), .B(u2__abc_52155_new_n4601_), .Y(u2__abc_52155_new_n5508_));
AND2X2 AND2X2_1694 ( .A(u2__abc_52155_new_n5509_), .B(u2__abc_52155_new_n4589_), .Y(u2__abc_52155_new_n5510_));
AND2X2 AND2X2_1695 ( .A(u2__abc_52155_new_n5483_), .B(u2__abc_52155_new_n5514_), .Y(u2__abc_52155_new_n5515_));
AND2X2 AND2X2_1696 ( .A(u2__abc_52155_new_n4496_), .B(u2__abc_52155_new_n4505_), .Y(u2__abc_52155_new_n5517_));
AND2X2 AND2X2_1697 ( .A(u2__abc_52155_new_n5518_), .B(u2__abc_52155_new_n4493_), .Y(u2__abc_52155_new_n5519_));
AND2X2 AND2X2_1698 ( .A(u2__abc_52155_new_n4488_), .B(u2__abc_52155_new_n4483_), .Y(u2__abc_52155_new_n5520_));
AND2X2 AND2X2_1699 ( .A(u2__abc_52155_new_n5522_), .B(u2__abc_52155_new_n4540_), .Y(u2__abc_52155_new_n5523_));
AND2X2 AND2X2_17 ( .A(_abc_73687_new_n753_), .B(sqrto_16_), .Y(\o[52] ));
AND2X2 AND2X2_170 ( .A(_abc_73687_new_n1110_), .B(_abc_73687_new_n1109_), .Y(\o[205] ));
AND2X2 AND2X2_1700 ( .A(u2__abc_52155_new_n4527_), .B(u2__abc_52155_new_n4536_), .Y(u2__abc_52155_new_n5524_));
AND2X2 AND2X2_1701 ( .A(u2__abc_52155_new_n5525_), .B(u2__abc_52155_new_n4524_), .Y(u2__abc_52155_new_n5526_));
AND2X2 AND2X2_1702 ( .A(u2__abc_52155_new_n4519_), .B(u2__abc_52155_new_n4514_), .Y(u2__abc_52155_new_n5527_));
AND2X2 AND2X2_1703 ( .A(u2__abc_52155_new_n5530_), .B(u2__abc_52155_new_n4478_), .Y(u2__abc_52155_new_n5531_));
AND2X2 AND2X2_1704 ( .A(u2__abc_52155_new_n4464_), .B(u2__abc_52155_new_n4473_), .Y(u2__abc_52155_new_n5532_));
AND2X2 AND2X2_1705 ( .A(u2__abc_52155_new_n5533_), .B(u2__abc_52155_new_n4461_), .Y(u2__abc_52155_new_n5534_));
AND2X2 AND2X2_1706 ( .A(u2__abc_52155_new_n4456_), .B(u2__abc_52155_new_n4451_), .Y(u2__abc_52155_new_n5535_));
AND2X2 AND2X2_1707 ( .A(u2__abc_52155_new_n5537_), .B(u2__abc_52155_new_n4446_), .Y(u2__abc_52155_new_n5538_));
AND2X2 AND2X2_1708 ( .A(u2__abc_52155_new_n4433_), .B(u2__abc_52155_new_n4442_), .Y(u2__abc_52155_new_n5539_));
AND2X2 AND2X2_1709 ( .A(u2__abc_52155_new_n5540_), .B(u2__abc_52155_new_n4430_), .Y(u2__abc_52155_new_n5541_));
AND2X2 AND2X2_171 ( .A(_abc_73687_new_n1113_), .B(_abc_73687_new_n1112_), .Y(\o[206] ));
AND2X2 AND2X2_1710 ( .A(u2__abc_52155_new_n4425_), .B(u2__abc_52155_new_n4420_), .Y(u2__abc_52155_new_n5542_));
AND2X2 AND2X2_1711 ( .A(u2__abc_52155_new_n5546_), .B(u2__abc_52155_new_n4415_), .Y(u2__abc_52155_new_n5547_));
AND2X2 AND2X2_1712 ( .A(u2__abc_52155_new_n4298_), .B(u2__abc_52155_new_n4293_), .Y(u2__abc_52155_new_n5548_));
AND2X2 AND2X2_1713 ( .A(u2__abc_52155_new_n5549_), .B(u2__abc_52155_new_n4318_), .Y(u2__abc_52155_new_n5550_));
AND2X2 AND2X2_1714 ( .A(u2__abc_52155_new_n4313_), .B(u2__abc_52155_new_n4308_), .Y(u2__abc_52155_new_n5551_));
AND2X2 AND2X2_1715 ( .A(u2__abc_52155_new_n5553_), .B(u2__abc_52155_new_n4350_), .Y(u2__abc_52155_new_n5554_));
AND2X2 AND2X2_1716 ( .A(u2__abc_52155_new_n4332_), .B(u2__abc_52155_new_n4324_), .Y(u2__abc_52155_new_n5555_));
AND2X2 AND2X2_1717 ( .A(u2__abc_52155_new_n4337_), .B(u2__abc_52155_new_n4346_), .Y(u2__abc_52155_new_n5557_));
AND2X2 AND2X2_1718 ( .A(u2__abc_52155_new_n5558_), .B(u2__abc_52155_new_n4334_), .Y(u2__abc_52155_new_n5559_));
AND2X2 AND2X2_1719 ( .A(u2__abc_52155_new_n4361_), .B(u2__abc_52155_new_n4356_), .Y(u2__abc_52155_new_n5562_));
AND2X2 AND2X2_172 ( .A(_abc_73687_new_n1116_), .B(_abc_73687_new_n1115_), .Y(\o[207] ));
AND2X2 AND2X2_1720 ( .A(u2__abc_52155_new_n5563_), .B(u2__abc_52155_new_n4381_), .Y(u2__abc_52155_new_n5564_));
AND2X2 AND2X2_1721 ( .A(u2__abc_52155_new_n4376_), .B(u2__abc_52155_new_n4371_), .Y(u2__abc_52155_new_n5565_));
AND2X2 AND2X2_1722 ( .A(u2__abc_52155_new_n5567_), .B(u2__abc_52155_new_n4413_), .Y(u2__abc_52155_new_n5568_));
AND2X2 AND2X2_1723 ( .A(u2__abc_52155_new_n4392_), .B(u2__abc_52155_new_n4387_), .Y(u2__abc_52155_new_n5569_));
AND2X2 AND2X2_1724 ( .A(u2__abc_52155_new_n4400_), .B(u2__abc_52155_new_n4409_), .Y(u2__abc_52155_new_n5571_));
AND2X2 AND2X2_1725 ( .A(u2__abc_52155_new_n5572_), .B(u2__abc_52155_new_n4397_), .Y(u2__abc_52155_new_n5573_));
AND2X2 AND2X2_1726 ( .A(u2__abc_52155_new_n5575_), .B(u2__abc_52155_new_n4351_), .Y(u2__abc_52155_new_n5576_));
AND2X2 AND2X2_1727 ( .A(u2__abc_52155_new_n5516_), .B(u2__abc_52155_new_n5579_), .Y(u2__abc_52155_new_n5580_));
AND2X2 AND2X2_1728 ( .A(u2__abc_52155_new_n5444_), .B(u2__abc_52155_new_n5580_), .Y(u2__abc_52155_new_n5581_));
AND2X2 AND2X2_1729 ( .A(u2__abc_52155_new_n5289_), .B(u2__abc_52155_new_n5581_), .Y(u2__abc_52155_new_n5582_));
AND2X2 AND2X2_173 ( .A(_abc_73687_new_n1119_), .B(_abc_73687_new_n1118_), .Y(\o[208] ));
AND2X2 AND2X2_1730 ( .A(u2__abc_52155_new_n5583_), .B(u2_remHi_380_), .Y(u2__abc_52155_new_n5584_));
AND2X2 AND2X2_1731 ( .A(u2__abc_52155_new_n5586_), .B(u2_o_380_), .Y(u2__abc_52155_new_n5587_));
AND2X2 AND2X2_1732 ( .A(u2__abc_52155_new_n5585_), .B(u2__abc_52155_new_n5588_), .Y(u2__abc_52155_new_n5589_));
AND2X2 AND2X2_1733 ( .A(u2__abc_52155_new_n5590_), .B(u2_o_381_), .Y(u2__abc_52155_new_n5591_));
AND2X2 AND2X2_1734 ( .A(u2__abc_52155_new_n5593_), .B(u2_remHi_381_), .Y(u2__abc_52155_new_n5594_));
AND2X2 AND2X2_1735 ( .A(u2__abc_52155_new_n5592_), .B(u2__abc_52155_new_n5595_), .Y(u2__abc_52155_new_n5596_));
AND2X2 AND2X2_1736 ( .A(u2__abc_52155_new_n5589_), .B(u2__abc_52155_new_n5596_), .Y(u2__abc_52155_new_n5597_));
AND2X2 AND2X2_1737 ( .A(u2__abc_52155_new_n5598_), .B(u2_remHi_378_), .Y(u2__abc_52155_new_n5599_));
AND2X2 AND2X2_1738 ( .A(u2__abc_52155_new_n5601_), .B(u2_o_378_), .Y(u2__abc_52155_new_n5602_));
AND2X2 AND2X2_1739 ( .A(u2__abc_52155_new_n5600_), .B(u2__abc_52155_new_n5603_), .Y(u2__abc_52155_new_n5604_));
AND2X2 AND2X2_174 ( .A(_abc_73687_new_n1122_), .B(_abc_73687_new_n1121_), .Y(\o[209] ));
AND2X2 AND2X2_1740 ( .A(u2__abc_52155_new_n5605_), .B(u2_remHi_379_), .Y(u2__abc_52155_new_n5606_));
AND2X2 AND2X2_1741 ( .A(u2__abc_52155_new_n5608_), .B(u2_o_379_), .Y(u2__abc_52155_new_n5609_));
AND2X2 AND2X2_1742 ( .A(u2__abc_52155_new_n5607_), .B(u2__abc_52155_new_n5610_), .Y(u2__abc_52155_new_n5611_));
AND2X2 AND2X2_1743 ( .A(u2__abc_52155_new_n5604_), .B(u2__abc_52155_new_n5611_), .Y(u2__abc_52155_new_n5612_));
AND2X2 AND2X2_1744 ( .A(u2__abc_52155_new_n5597_), .B(u2__abc_52155_new_n5612_), .Y(u2__abc_52155_new_n5613_));
AND2X2 AND2X2_1745 ( .A(u2__abc_52155_new_n5614_), .B(u2_o_374_), .Y(u2__abc_52155_new_n5615_));
AND2X2 AND2X2_1746 ( .A(u2__abc_52155_new_n5617_), .B(u2_remHi_374_), .Y(u2__abc_52155_new_n5618_));
AND2X2 AND2X2_1747 ( .A(u2__abc_52155_new_n5616_), .B(u2__abc_52155_new_n5619_), .Y(u2__abc_52155_new_n5620_));
AND2X2 AND2X2_1748 ( .A(u2__abc_52155_new_n5621_), .B(u2_o_375_), .Y(u2__abc_52155_new_n5622_));
AND2X2 AND2X2_1749 ( .A(u2__abc_52155_new_n5624_), .B(u2_remHi_375_), .Y(u2__abc_52155_new_n5625_));
AND2X2 AND2X2_175 ( .A(_abc_73687_new_n1125_), .B(_abc_73687_new_n1124_), .Y(\o[210] ));
AND2X2 AND2X2_1750 ( .A(u2__abc_52155_new_n5623_), .B(u2__abc_52155_new_n5626_), .Y(u2__abc_52155_new_n5627_));
AND2X2 AND2X2_1751 ( .A(u2__abc_52155_new_n5620_), .B(u2__abc_52155_new_n5627_), .Y(u2__abc_52155_new_n5628_));
AND2X2 AND2X2_1752 ( .A(u2__abc_52155_new_n5629_), .B(u2_remHi_376_), .Y(u2__abc_52155_new_n5630_));
AND2X2 AND2X2_1753 ( .A(u2__abc_52155_new_n5632_), .B(u2_o_376_), .Y(u2__abc_52155_new_n5633_));
AND2X2 AND2X2_1754 ( .A(u2__abc_52155_new_n5631_), .B(u2__abc_52155_new_n5634_), .Y(u2__abc_52155_new_n5635_));
AND2X2 AND2X2_1755 ( .A(u2__abc_52155_new_n5636_), .B(u2_remHi_377_), .Y(u2__abc_52155_new_n5637_));
AND2X2 AND2X2_1756 ( .A(u2__abc_52155_new_n5639_), .B(u2_o_377_), .Y(u2__abc_52155_new_n5640_));
AND2X2 AND2X2_1757 ( .A(u2__abc_52155_new_n5638_), .B(u2__abc_52155_new_n5641_), .Y(u2__abc_52155_new_n5642_));
AND2X2 AND2X2_1758 ( .A(u2__abc_52155_new_n5635_), .B(u2__abc_52155_new_n5642_), .Y(u2__abc_52155_new_n5643_));
AND2X2 AND2X2_1759 ( .A(u2__abc_52155_new_n5628_), .B(u2__abc_52155_new_n5643_), .Y(u2__abc_52155_new_n5644_));
AND2X2 AND2X2_176 ( .A(_abc_73687_new_n1128_), .B(_abc_73687_new_n1127_), .Y(\o[211] ));
AND2X2 AND2X2_1760 ( .A(u2__abc_52155_new_n5613_), .B(u2__abc_52155_new_n5644_), .Y(u2__abc_52155_new_n5645_));
AND2X2 AND2X2_1761 ( .A(u2__abc_52155_new_n5646_), .B(u2_remHi_368_), .Y(u2__abc_52155_new_n5647_));
AND2X2 AND2X2_1762 ( .A(u2__abc_52155_new_n5649_), .B(u2_o_368_), .Y(u2__abc_52155_new_n5650_));
AND2X2 AND2X2_1763 ( .A(u2__abc_52155_new_n5648_), .B(u2__abc_52155_new_n5651_), .Y(u2__abc_52155_new_n5652_));
AND2X2 AND2X2_1764 ( .A(u2__abc_52155_new_n5653_), .B(u2_remHi_369_), .Y(u2__abc_52155_new_n5654_));
AND2X2 AND2X2_1765 ( .A(u2__abc_52155_new_n5656_), .B(u2_o_369_), .Y(u2__abc_52155_new_n5657_));
AND2X2 AND2X2_1766 ( .A(u2__abc_52155_new_n5655_), .B(u2__abc_52155_new_n5658_), .Y(u2__abc_52155_new_n5659_));
AND2X2 AND2X2_1767 ( .A(u2__abc_52155_new_n5652_), .B(u2__abc_52155_new_n5659_), .Y(u2__abc_52155_new_n5660_));
AND2X2 AND2X2_1768 ( .A(u2__abc_52155_new_n5661_), .B(u2_remHi_366_), .Y(u2__abc_52155_new_n5662_));
AND2X2 AND2X2_1769 ( .A(u2__abc_52155_new_n5664_), .B(u2_o_366_), .Y(u2__abc_52155_new_n5665_));
AND2X2 AND2X2_177 ( .A(_abc_73687_new_n1131_), .B(_abc_73687_new_n1130_), .Y(\o[212] ));
AND2X2 AND2X2_1770 ( .A(u2__abc_52155_new_n5663_), .B(u2__abc_52155_new_n5666_), .Y(u2__abc_52155_new_n5667_));
AND2X2 AND2X2_1771 ( .A(u2__abc_52155_new_n5668_), .B(u2_remHi_367_), .Y(u2__abc_52155_new_n5669_));
AND2X2 AND2X2_1772 ( .A(u2__abc_52155_new_n5671_), .B(u2_o_367_), .Y(u2__abc_52155_new_n5672_));
AND2X2 AND2X2_1773 ( .A(u2__abc_52155_new_n5670_), .B(u2__abc_52155_new_n5673_), .Y(u2__abc_52155_new_n5674_));
AND2X2 AND2X2_1774 ( .A(u2__abc_52155_new_n5667_), .B(u2__abc_52155_new_n5674_), .Y(u2__abc_52155_new_n5675_));
AND2X2 AND2X2_1775 ( .A(u2__abc_52155_new_n5660_), .B(u2__abc_52155_new_n5675_), .Y(u2__abc_52155_new_n5676_));
AND2X2 AND2X2_1776 ( .A(u2__abc_52155_new_n5677_), .B(u2_remHi_372_), .Y(u2__abc_52155_new_n5678_));
AND2X2 AND2X2_1777 ( .A(u2__abc_52155_new_n5680_), .B(u2_o_372_), .Y(u2__abc_52155_new_n5681_));
AND2X2 AND2X2_1778 ( .A(u2__abc_52155_new_n5679_), .B(u2__abc_52155_new_n5682_), .Y(u2__abc_52155_new_n5683_));
AND2X2 AND2X2_1779 ( .A(u2__abc_52155_new_n5684_), .B(u2_remHi_373_), .Y(u2__abc_52155_new_n5685_));
AND2X2 AND2X2_178 ( .A(_abc_73687_new_n1134_), .B(_abc_73687_new_n1133_), .Y(\o[213] ));
AND2X2 AND2X2_1780 ( .A(u2__abc_52155_new_n5687_), .B(u2_o_373_), .Y(u2__abc_52155_new_n5688_));
AND2X2 AND2X2_1781 ( .A(u2__abc_52155_new_n5686_), .B(u2__abc_52155_new_n5689_), .Y(u2__abc_52155_new_n5690_));
AND2X2 AND2X2_1782 ( .A(u2__abc_52155_new_n5683_), .B(u2__abc_52155_new_n5690_), .Y(u2__abc_52155_new_n5691_));
AND2X2 AND2X2_1783 ( .A(u2__abc_52155_new_n5692_), .B(u2_remHi_371_), .Y(u2__abc_52155_new_n5693_));
AND2X2 AND2X2_1784 ( .A(u2__abc_52155_new_n5695_), .B(u2_o_371_), .Y(u2__abc_52155_new_n5696_));
AND2X2 AND2X2_1785 ( .A(u2__abc_52155_new_n5694_), .B(u2__abc_52155_new_n5697_), .Y(u2__abc_52155_new_n5698_));
AND2X2 AND2X2_1786 ( .A(u2__abc_52155_new_n5699_), .B(u2_remHi_370_), .Y(u2__abc_52155_new_n5700_));
AND2X2 AND2X2_1787 ( .A(u2__abc_52155_new_n5702_), .B(u2_o_370_), .Y(u2__abc_52155_new_n5703_));
AND2X2 AND2X2_1788 ( .A(u2__abc_52155_new_n5701_), .B(u2__abc_52155_new_n5704_), .Y(u2__abc_52155_new_n5705_));
AND2X2 AND2X2_1789 ( .A(u2__abc_52155_new_n5698_), .B(u2__abc_52155_new_n5705_), .Y(u2__abc_52155_new_n5706_));
AND2X2 AND2X2_179 ( .A(_abc_73687_new_n1137_), .B(_abc_73687_new_n1136_), .Y(\o[214] ));
AND2X2 AND2X2_1790 ( .A(u2__abc_52155_new_n5691_), .B(u2__abc_52155_new_n5706_), .Y(u2__abc_52155_new_n5707_));
AND2X2 AND2X2_1791 ( .A(u2__abc_52155_new_n5676_), .B(u2__abc_52155_new_n5707_), .Y(u2__abc_52155_new_n5708_));
AND2X2 AND2X2_1792 ( .A(u2__abc_52155_new_n5645_), .B(u2__abc_52155_new_n5708_), .Y(u2__abc_52155_new_n5709_));
AND2X2 AND2X2_1793 ( .A(u2__abc_52155_new_n5710_), .B(u2_o_358_), .Y(u2__abc_52155_new_n5711_));
AND2X2 AND2X2_1794 ( .A(u2__abc_52155_new_n5713_), .B(u2_remHi_358_), .Y(u2__abc_52155_new_n5714_));
AND2X2 AND2X2_1795 ( .A(u2__abc_52155_new_n5712_), .B(u2__abc_52155_new_n5715_), .Y(u2__abc_52155_new_n5716_));
AND2X2 AND2X2_1796 ( .A(u2__abc_52155_new_n5717_), .B(u2_o_359_), .Y(u2__abc_52155_new_n5718_));
AND2X2 AND2X2_1797 ( .A(u2__abc_52155_new_n5720_), .B(u2_remHi_359_), .Y(u2__abc_52155_new_n5721_));
AND2X2 AND2X2_1798 ( .A(u2__abc_52155_new_n5719_), .B(u2__abc_52155_new_n5722_), .Y(u2__abc_52155_new_n5723_));
AND2X2 AND2X2_1799 ( .A(u2__abc_52155_new_n5716_), .B(u2__abc_52155_new_n5723_), .Y(u2__abc_52155_new_n5724_));
AND2X2 AND2X2_18 ( .A(_abc_73687_new_n753_), .B(sqrto_17_), .Y(\o[53] ));
AND2X2 AND2X2_180 ( .A(_abc_73687_new_n1140_), .B(_abc_73687_new_n1139_), .Y(\o[215] ));
AND2X2 AND2X2_1800 ( .A(u2__abc_52155_new_n5725_), .B(u2_remHi_360_), .Y(u2__abc_52155_new_n5726_));
AND2X2 AND2X2_1801 ( .A(u2__abc_52155_new_n5728_), .B(u2_o_360_), .Y(u2__abc_52155_new_n5729_));
AND2X2 AND2X2_1802 ( .A(u2__abc_52155_new_n5727_), .B(u2__abc_52155_new_n5730_), .Y(u2__abc_52155_new_n5731_));
AND2X2 AND2X2_1803 ( .A(u2__abc_52155_new_n5732_), .B(u2_remHi_361_), .Y(u2__abc_52155_new_n5733_));
AND2X2 AND2X2_1804 ( .A(u2__abc_52155_new_n5735_), .B(u2_o_361_), .Y(u2__abc_52155_new_n5736_));
AND2X2 AND2X2_1805 ( .A(u2__abc_52155_new_n5734_), .B(u2__abc_52155_new_n5737_), .Y(u2__abc_52155_new_n5738_));
AND2X2 AND2X2_1806 ( .A(u2__abc_52155_new_n5731_), .B(u2__abc_52155_new_n5738_), .Y(u2__abc_52155_new_n5739_));
AND2X2 AND2X2_1807 ( .A(u2__abc_52155_new_n5724_), .B(u2__abc_52155_new_n5739_), .Y(u2__abc_52155_new_n5740_));
AND2X2 AND2X2_1808 ( .A(u2__abc_52155_new_n5741_), .B(u2_remHi_364_), .Y(u2__abc_52155_new_n5742_));
AND2X2 AND2X2_1809 ( .A(u2__abc_52155_new_n5744_), .B(u2_o_364_), .Y(u2__abc_52155_new_n5745_));
AND2X2 AND2X2_181 ( .A(_abc_73687_new_n1143_), .B(_abc_73687_new_n1142_), .Y(\o[216] ));
AND2X2 AND2X2_1810 ( .A(u2__abc_52155_new_n5743_), .B(u2__abc_52155_new_n5746_), .Y(u2__abc_52155_new_n5747_));
AND2X2 AND2X2_1811 ( .A(u2__abc_52155_new_n5748_), .B(u2_remHi_365_), .Y(u2__abc_52155_new_n5749_));
AND2X2 AND2X2_1812 ( .A(u2__abc_52155_new_n5751_), .B(u2_o_365_), .Y(u2__abc_52155_new_n5752_));
AND2X2 AND2X2_1813 ( .A(u2__abc_52155_new_n5750_), .B(u2__abc_52155_new_n5753_), .Y(u2__abc_52155_new_n5754_));
AND2X2 AND2X2_1814 ( .A(u2__abc_52155_new_n5747_), .B(u2__abc_52155_new_n5754_), .Y(u2__abc_52155_new_n5755_));
AND2X2 AND2X2_1815 ( .A(u2__abc_52155_new_n5756_), .B(u2_remHi_362_), .Y(u2__abc_52155_new_n5757_));
AND2X2 AND2X2_1816 ( .A(u2__abc_52155_new_n5759_), .B(u2_o_362_), .Y(u2__abc_52155_new_n5760_));
AND2X2 AND2X2_1817 ( .A(u2__abc_52155_new_n5758_), .B(u2__abc_52155_new_n5761_), .Y(u2__abc_52155_new_n5762_));
AND2X2 AND2X2_1818 ( .A(u2__abc_52155_new_n5763_), .B(u2_remHi_363_), .Y(u2__abc_52155_new_n5764_));
AND2X2 AND2X2_1819 ( .A(u2__abc_52155_new_n5766_), .B(u2_o_363_), .Y(u2__abc_52155_new_n5767_));
AND2X2 AND2X2_182 ( .A(_abc_73687_new_n1146_), .B(_abc_73687_new_n1145_), .Y(\o[217] ));
AND2X2 AND2X2_1820 ( .A(u2__abc_52155_new_n5765_), .B(u2__abc_52155_new_n5768_), .Y(u2__abc_52155_new_n5769_));
AND2X2 AND2X2_1821 ( .A(u2__abc_52155_new_n5762_), .B(u2__abc_52155_new_n5769_), .Y(u2__abc_52155_new_n5770_));
AND2X2 AND2X2_1822 ( .A(u2__abc_52155_new_n5755_), .B(u2__abc_52155_new_n5770_), .Y(u2__abc_52155_new_n5771_));
AND2X2 AND2X2_1823 ( .A(u2__abc_52155_new_n5740_), .B(u2__abc_52155_new_n5771_), .Y(u2__abc_52155_new_n5772_));
AND2X2 AND2X2_1824 ( .A(u2__abc_52155_new_n5773_), .B(u2_remHi_352_), .Y(u2__abc_52155_new_n5774_));
AND2X2 AND2X2_1825 ( .A(u2__abc_52155_new_n5776_), .B(u2_o_352_), .Y(u2__abc_52155_new_n5777_));
AND2X2 AND2X2_1826 ( .A(u2__abc_52155_new_n5775_), .B(u2__abc_52155_new_n5778_), .Y(u2__abc_52155_new_n5779_));
AND2X2 AND2X2_1827 ( .A(u2__abc_52155_new_n5780_), .B(u2_remHi_353_), .Y(u2__abc_52155_new_n5781_));
AND2X2 AND2X2_1828 ( .A(u2__abc_52155_new_n5783_), .B(u2_o_353_), .Y(u2__abc_52155_new_n5784_));
AND2X2 AND2X2_1829 ( .A(u2__abc_52155_new_n5782_), .B(u2__abc_52155_new_n5785_), .Y(u2__abc_52155_new_n5786_));
AND2X2 AND2X2_183 ( .A(_abc_73687_new_n1149_), .B(_abc_73687_new_n1148_), .Y(\o[218] ));
AND2X2 AND2X2_1830 ( .A(u2__abc_52155_new_n5779_), .B(u2__abc_52155_new_n5786_), .Y(u2__abc_52155_new_n5787_));
AND2X2 AND2X2_1831 ( .A(u2__abc_52155_new_n5788_), .B(u2_remHi_350_), .Y(u2__abc_52155_new_n5789_));
AND2X2 AND2X2_1832 ( .A(u2__abc_52155_new_n5791_), .B(u2_o_350_), .Y(u2__abc_52155_new_n5792_));
AND2X2 AND2X2_1833 ( .A(u2__abc_52155_new_n5790_), .B(u2__abc_52155_new_n5793_), .Y(u2__abc_52155_new_n5794_));
AND2X2 AND2X2_1834 ( .A(u2__abc_52155_new_n5795_), .B(u2_remHi_351_), .Y(u2__abc_52155_new_n5796_));
AND2X2 AND2X2_1835 ( .A(u2__abc_52155_new_n5798_), .B(u2_o_351_), .Y(u2__abc_52155_new_n5799_));
AND2X2 AND2X2_1836 ( .A(u2__abc_52155_new_n5797_), .B(u2__abc_52155_new_n5800_), .Y(u2__abc_52155_new_n5801_));
AND2X2 AND2X2_1837 ( .A(u2__abc_52155_new_n5794_), .B(u2__abc_52155_new_n5801_), .Y(u2__abc_52155_new_n5802_));
AND2X2 AND2X2_1838 ( .A(u2__abc_52155_new_n5787_), .B(u2__abc_52155_new_n5802_), .Y(u2__abc_52155_new_n5803_));
AND2X2 AND2X2_1839 ( .A(u2__abc_52155_new_n5804_), .B(u2_remHi_356_), .Y(u2__abc_52155_new_n5805_));
AND2X2 AND2X2_184 ( .A(_abc_73687_new_n1152_), .B(_abc_73687_new_n1151_), .Y(\o[219] ));
AND2X2 AND2X2_1840 ( .A(u2__abc_52155_new_n5807_), .B(u2_o_356_), .Y(u2__abc_52155_new_n5808_));
AND2X2 AND2X2_1841 ( .A(u2__abc_52155_new_n5806_), .B(u2__abc_52155_new_n5809_), .Y(u2__abc_52155_new_n5810_));
AND2X2 AND2X2_1842 ( .A(u2__abc_52155_new_n5811_), .B(u2_remHi_357_), .Y(u2__abc_52155_new_n5812_));
AND2X2 AND2X2_1843 ( .A(u2__abc_52155_new_n5814_), .B(u2_o_357_), .Y(u2__abc_52155_new_n5815_));
AND2X2 AND2X2_1844 ( .A(u2__abc_52155_new_n5813_), .B(u2__abc_52155_new_n5816_), .Y(u2__abc_52155_new_n5817_));
AND2X2 AND2X2_1845 ( .A(u2__abc_52155_new_n5810_), .B(u2__abc_52155_new_n5817_), .Y(u2__abc_52155_new_n5818_));
AND2X2 AND2X2_1846 ( .A(u2__abc_52155_new_n5819_), .B(u2_remHi_354_), .Y(u2__abc_52155_new_n5820_));
AND2X2 AND2X2_1847 ( .A(u2__abc_52155_new_n5822_), .B(u2_o_354_), .Y(u2__abc_52155_new_n5823_));
AND2X2 AND2X2_1848 ( .A(u2__abc_52155_new_n5821_), .B(u2__abc_52155_new_n5824_), .Y(u2__abc_52155_new_n5825_));
AND2X2 AND2X2_1849 ( .A(u2__abc_52155_new_n5826_), .B(u2_remHi_355_), .Y(u2__abc_52155_new_n5827_));
AND2X2 AND2X2_185 ( .A(_abc_73687_new_n1155_), .B(_abc_73687_new_n1154_), .Y(\o[220] ));
AND2X2 AND2X2_1850 ( .A(u2__abc_52155_new_n5829_), .B(u2_o_355_), .Y(u2__abc_52155_new_n5830_));
AND2X2 AND2X2_1851 ( .A(u2__abc_52155_new_n5828_), .B(u2__abc_52155_new_n5831_), .Y(u2__abc_52155_new_n5832_));
AND2X2 AND2X2_1852 ( .A(u2__abc_52155_new_n5825_), .B(u2__abc_52155_new_n5832_), .Y(u2__abc_52155_new_n5833_));
AND2X2 AND2X2_1853 ( .A(u2__abc_52155_new_n5818_), .B(u2__abc_52155_new_n5833_), .Y(u2__abc_52155_new_n5834_));
AND2X2 AND2X2_1854 ( .A(u2__abc_52155_new_n5803_), .B(u2__abc_52155_new_n5834_), .Y(u2__abc_52155_new_n5835_));
AND2X2 AND2X2_1855 ( .A(u2__abc_52155_new_n5772_), .B(u2__abc_52155_new_n5835_), .Y(u2__abc_52155_new_n5836_));
AND2X2 AND2X2_1856 ( .A(u2__abc_52155_new_n5709_), .B(u2__abc_52155_new_n5836_), .Y(u2__abc_52155_new_n5837_));
AND2X2 AND2X2_1857 ( .A(u2__abc_52155_new_n5838_), .B(u2_remHi_344_), .Y(u2__abc_52155_new_n5839_));
AND2X2 AND2X2_1858 ( .A(u2__abc_52155_new_n5841_), .B(u2_o_344_), .Y(u2__abc_52155_new_n5842_));
AND2X2 AND2X2_1859 ( .A(u2__abc_52155_new_n5840_), .B(u2__abc_52155_new_n5843_), .Y(u2__abc_52155_new_n5844_));
AND2X2 AND2X2_186 ( .A(_abc_73687_new_n1158_), .B(_abc_73687_new_n1157_), .Y(\o[221] ));
AND2X2 AND2X2_1860 ( .A(u2__abc_52155_new_n5845_), .B(u2_remHi_345_), .Y(u2__abc_52155_new_n5846_));
AND2X2 AND2X2_1861 ( .A(u2__abc_52155_new_n5848_), .B(u2_o_345_), .Y(u2__abc_52155_new_n5849_));
AND2X2 AND2X2_1862 ( .A(u2__abc_52155_new_n5847_), .B(u2__abc_52155_new_n5850_), .Y(u2__abc_52155_new_n5851_));
AND2X2 AND2X2_1863 ( .A(u2__abc_52155_new_n5844_), .B(u2__abc_52155_new_n5851_), .Y(u2__abc_52155_new_n5852_));
AND2X2 AND2X2_1864 ( .A(u2__abc_52155_new_n5853_), .B(u2_remHi_342_), .Y(u2__abc_52155_new_n5854_));
AND2X2 AND2X2_1865 ( .A(u2__abc_52155_new_n5856_), .B(u2_o_342_), .Y(u2__abc_52155_new_n5857_));
AND2X2 AND2X2_1866 ( .A(u2__abc_52155_new_n5855_), .B(u2__abc_52155_new_n5858_), .Y(u2__abc_52155_new_n5859_));
AND2X2 AND2X2_1867 ( .A(u2__abc_52155_new_n5860_), .B(u2_remHi_343_), .Y(u2__abc_52155_new_n5861_));
AND2X2 AND2X2_1868 ( .A(u2__abc_52155_new_n5863_), .B(u2_o_343_), .Y(u2__abc_52155_new_n5864_));
AND2X2 AND2X2_1869 ( .A(u2__abc_52155_new_n5862_), .B(u2__abc_52155_new_n5865_), .Y(u2__abc_52155_new_n5866_));
AND2X2 AND2X2_187 ( .A(_abc_73687_new_n1161_), .B(_abc_73687_new_n1160_), .Y(\o[222] ));
AND2X2 AND2X2_1870 ( .A(u2__abc_52155_new_n5859_), .B(u2__abc_52155_new_n5866_), .Y(u2__abc_52155_new_n5867_));
AND2X2 AND2X2_1871 ( .A(u2__abc_52155_new_n5852_), .B(u2__abc_52155_new_n5867_), .Y(u2__abc_52155_new_n5868_));
AND2X2 AND2X2_1872 ( .A(u2__abc_52155_new_n5869_), .B(u2_remHi_348_), .Y(u2__abc_52155_new_n5870_));
AND2X2 AND2X2_1873 ( .A(u2__abc_52155_new_n5872_), .B(u2_o_348_), .Y(u2__abc_52155_new_n5873_));
AND2X2 AND2X2_1874 ( .A(u2__abc_52155_new_n5871_), .B(u2__abc_52155_new_n5874_), .Y(u2__abc_52155_new_n5875_));
AND2X2 AND2X2_1875 ( .A(u2__abc_52155_new_n5876_), .B(u2_remHi_349_), .Y(u2__abc_52155_new_n5877_));
AND2X2 AND2X2_1876 ( .A(u2__abc_52155_new_n5879_), .B(u2_o_349_), .Y(u2__abc_52155_new_n5880_));
AND2X2 AND2X2_1877 ( .A(u2__abc_52155_new_n5878_), .B(u2__abc_52155_new_n5881_), .Y(u2__abc_52155_new_n5882_));
AND2X2 AND2X2_1878 ( .A(u2__abc_52155_new_n5875_), .B(u2__abc_52155_new_n5882_), .Y(u2__abc_52155_new_n5883_));
AND2X2 AND2X2_1879 ( .A(u2__abc_52155_new_n5884_), .B(u2_remHi_346_), .Y(u2__abc_52155_new_n5885_));
AND2X2 AND2X2_188 ( .A(_abc_73687_new_n1164_), .B(_abc_73687_new_n1163_), .Y(\o[223] ));
AND2X2 AND2X2_1880 ( .A(u2__abc_52155_new_n5887_), .B(u2_o_346_), .Y(u2__abc_52155_new_n5888_));
AND2X2 AND2X2_1881 ( .A(u2__abc_52155_new_n5886_), .B(u2__abc_52155_new_n5889_), .Y(u2__abc_52155_new_n5890_));
AND2X2 AND2X2_1882 ( .A(u2__abc_52155_new_n5891_), .B(u2_remHi_347_), .Y(u2__abc_52155_new_n5892_));
AND2X2 AND2X2_1883 ( .A(u2__abc_52155_new_n5894_), .B(u2_o_347_), .Y(u2__abc_52155_new_n5895_));
AND2X2 AND2X2_1884 ( .A(u2__abc_52155_new_n5893_), .B(u2__abc_52155_new_n5896_), .Y(u2__abc_52155_new_n5897_));
AND2X2 AND2X2_1885 ( .A(u2__abc_52155_new_n5890_), .B(u2__abc_52155_new_n5897_), .Y(u2__abc_52155_new_n5898_));
AND2X2 AND2X2_1886 ( .A(u2__abc_52155_new_n5883_), .B(u2__abc_52155_new_n5898_), .Y(u2__abc_52155_new_n5899_));
AND2X2 AND2X2_1887 ( .A(u2__abc_52155_new_n5868_), .B(u2__abc_52155_new_n5899_), .Y(u2__abc_52155_new_n5900_));
AND2X2 AND2X2_1888 ( .A(u2__abc_52155_new_n5901_), .B(u2_remHi_336_), .Y(u2__abc_52155_new_n5902_));
AND2X2 AND2X2_1889 ( .A(u2__abc_52155_new_n5904_), .B(u2_o_336_), .Y(u2__abc_52155_new_n5905_));
AND2X2 AND2X2_189 ( .A(_abc_73687_new_n753_), .B(sqrto_189_), .Y(\o[225] ));
AND2X2 AND2X2_1890 ( .A(u2__abc_52155_new_n5903_), .B(u2__abc_52155_new_n5906_), .Y(u2__abc_52155_new_n5907_));
AND2X2 AND2X2_1891 ( .A(u2__abc_52155_new_n5908_), .B(u2_remHi_337_), .Y(u2__abc_52155_new_n5909_));
AND2X2 AND2X2_1892 ( .A(u2__abc_52155_new_n5911_), .B(u2_o_337_), .Y(u2__abc_52155_new_n5912_));
AND2X2 AND2X2_1893 ( .A(u2__abc_52155_new_n5910_), .B(u2__abc_52155_new_n5913_), .Y(u2__abc_52155_new_n5914_));
AND2X2 AND2X2_1894 ( .A(u2__abc_52155_new_n5907_), .B(u2__abc_52155_new_n5914_), .Y(u2__abc_52155_new_n5915_));
AND2X2 AND2X2_1895 ( .A(u2__abc_52155_new_n5916_), .B(u2_remHi_334_), .Y(u2__abc_52155_new_n5917_));
AND2X2 AND2X2_1896 ( .A(u2__abc_52155_new_n5919_), .B(u2_o_334_), .Y(u2__abc_52155_new_n5920_));
AND2X2 AND2X2_1897 ( .A(u2__abc_52155_new_n5918_), .B(u2__abc_52155_new_n5921_), .Y(u2__abc_52155_new_n5922_));
AND2X2 AND2X2_1898 ( .A(u2__abc_52155_new_n5923_), .B(u2_remHi_335_), .Y(u2__abc_52155_new_n5924_));
AND2X2 AND2X2_1899 ( .A(u2__abc_52155_new_n5926_), .B(u2_o_335_), .Y(u2__abc_52155_new_n5927_));
AND2X2 AND2X2_19 ( .A(_abc_73687_new_n753_), .B(sqrto_18_), .Y(\o[54] ));
AND2X2 AND2X2_190 ( .A(\a[112] ), .B(\a[0] ), .Y(fracta1_0_));
AND2X2 AND2X2_1900 ( .A(u2__abc_52155_new_n5925_), .B(u2__abc_52155_new_n5928_), .Y(u2__abc_52155_new_n5929_));
AND2X2 AND2X2_1901 ( .A(u2__abc_52155_new_n5922_), .B(u2__abc_52155_new_n5929_), .Y(u2__abc_52155_new_n5930_));
AND2X2 AND2X2_1902 ( .A(u2__abc_52155_new_n5915_), .B(u2__abc_52155_new_n5930_), .Y(u2__abc_52155_new_n5931_));
AND2X2 AND2X2_1903 ( .A(u2__abc_52155_new_n5932_), .B(u2_remHi_340_), .Y(u2__abc_52155_new_n5933_));
AND2X2 AND2X2_1904 ( .A(u2__abc_52155_new_n5935_), .B(u2_o_340_), .Y(u2__abc_52155_new_n5936_));
AND2X2 AND2X2_1905 ( .A(u2__abc_52155_new_n5934_), .B(u2__abc_52155_new_n5937_), .Y(u2__abc_52155_new_n5938_));
AND2X2 AND2X2_1906 ( .A(u2__abc_52155_new_n5939_), .B(u2_remHi_341_), .Y(u2__abc_52155_new_n5940_));
AND2X2 AND2X2_1907 ( .A(u2__abc_52155_new_n5942_), .B(u2_o_341_), .Y(u2__abc_52155_new_n5943_));
AND2X2 AND2X2_1908 ( .A(u2__abc_52155_new_n5941_), .B(u2__abc_52155_new_n5944_), .Y(u2__abc_52155_new_n5945_));
AND2X2 AND2X2_1909 ( .A(u2__abc_52155_new_n5938_), .B(u2__abc_52155_new_n5945_), .Y(u2__abc_52155_new_n5946_));
AND2X2 AND2X2_191 ( .A(_abc_73687_new_n1171_), .B(_abc_73687_new_n1169_), .Y(fracta1_1_));
AND2X2 AND2X2_1910 ( .A(u2__abc_52155_new_n5947_), .B(u2_remHi_338_), .Y(u2__abc_52155_new_n5948_));
AND2X2 AND2X2_1911 ( .A(u2__abc_52155_new_n5950_), .B(u2_o_338_), .Y(u2__abc_52155_new_n5951_));
AND2X2 AND2X2_1912 ( .A(u2__abc_52155_new_n5949_), .B(u2__abc_52155_new_n5952_), .Y(u2__abc_52155_new_n5953_));
AND2X2 AND2X2_1913 ( .A(u2__abc_52155_new_n5954_), .B(u2_remHi_339_), .Y(u2__abc_52155_new_n5955_));
AND2X2 AND2X2_1914 ( .A(u2__abc_52155_new_n5957_), .B(u2_o_339_), .Y(u2__abc_52155_new_n5958_));
AND2X2 AND2X2_1915 ( .A(u2__abc_52155_new_n5956_), .B(u2__abc_52155_new_n5959_), .Y(u2__abc_52155_new_n5960_));
AND2X2 AND2X2_1916 ( .A(u2__abc_52155_new_n5953_), .B(u2__abc_52155_new_n5960_), .Y(u2__abc_52155_new_n5961_));
AND2X2 AND2X2_1917 ( .A(u2__abc_52155_new_n5946_), .B(u2__abc_52155_new_n5961_), .Y(u2__abc_52155_new_n5962_));
AND2X2 AND2X2_1918 ( .A(u2__abc_52155_new_n5931_), .B(u2__abc_52155_new_n5962_), .Y(u2__abc_52155_new_n5963_));
AND2X2 AND2X2_1919 ( .A(u2__abc_52155_new_n5900_), .B(u2__abc_52155_new_n5963_), .Y(u2__abc_52155_new_n5964_));
AND2X2 AND2X2_192 ( .A(_abc_73687_new_n1174_), .B(_abc_73687_new_n1173_), .Y(fracta1_2_));
AND2X2 AND2X2_1920 ( .A(u2__abc_52155_new_n5965_), .B(u2_o_326_), .Y(u2__abc_52155_new_n5966_));
AND2X2 AND2X2_1921 ( .A(u2__abc_52155_new_n5968_), .B(u2_remHi_326_), .Y(u2__abc_52155_new_n5969_));
AND2X2 AND2X2_1922 ( .A(u2__abc_52155_new_n5967_), .B(u2__abc_52155_new_n5970_), .Y(u2__abc_52155_new_n5971_));
AND2X2 AND2X2_1923 ( .A(u2__abc_52155_new_n5972_), .B(u2_o_327_), .Y(u2__abc_52155_new_n5973_));
AND2X2 AND2X2_1924 ( .A(u2__abc_52155_new_n5975_), .B(u2_remHi_327_), .Y(u2__abc_52155_new_n5976_));
AND2X2 AND2X2_1925 ( .A(u2__abc_52155_new_n5974_), .B(u2__abc_52155_new_n5977_), .Y(u2__abc_52155_new_n5978_));
AND2X2 AND2X2_1926 ( .A(u2__abc_52155_new_n5971_), .B(u2__abc_52155_new_n5978_), .Y(u2__abc_52155_new_n5979_));
AND2X2 AND2X2_1927 ( .A(u2__abc_52155_new_n5980_), .B(u2_remHi_328_), .Y(u2__abc_52155_new_n5981_));
AND2X2 AND2X2_1928 ( .A(u2__abc_52155_new_n5983_), .B(u2_o_328_), .Y(u2__abc_52155_new_n5984_));
AND2X2 AND2X2_1929 ( .A(u2__abc_52155_new_n5982_), .B(u2__abc_52155_new_n5985_), .Y(u2__abc_52155_new_n5986_));
AND2X2 AND2X2_193 ( .A(_abc_73687_new_n1177_), .B(_abc_73687_new_n1176_), .Y(fracta1_3_));
AND2X2 AND2X2_1930 ( .A(u2__abc_52155_new_n5987_), .B(u2_remHi_329_), .Y(u2__abc_52155_new_n5988_));
AND2X2 AND2X2_1931 ( .A(u2__abc_52155_new_n5990_), .B(u2_o_329_), .Y(u2__abc_52155_new_n5991_));
AND2X2 AND2X2_1932 ( .A(u2__abc_52155_new_n5989_), .B(u2__abc_52155_new_n5992_), .Y(u2__abc_52155_new_n5993_));
AND2X2 AND2X2_1933 ( .A(u2__abc_52155_new_n5986_), .B(u2__abc_52155_new_n5993_), .Y(u2__abc_52155_new_n5994_));
AND2X2 AND2X2_1934 ( .A(u2__abc_52155_new_n5979_), .B(u2__abc_52155_new_n5994_), .Y(u2__abc_52155_new_n5995_));
AND2X2 AND2X2_1935 ( .A(u2__abc_52155_new_n5996_), .B(u2_remHi_332_), .Y(u2__abc_52155_new_n5997_));
AND2X2 AND2X2_1936 ( .A(u2__abc_52155_new_n5999_), .B(u2_o_332_), .Y(u2__abc_52155_new_n6000_));
AND2X2 AND2X2_1937 ( .A(u2__abc_52155_new_n5998_), .B(u2__abc_52155_new_n6001_), .Y(u2__abc_52155_new_n6002_));
AND2X2 AND2X2_1938 ( .A(u2__abc_52155_new_n6003_), .B(u2_remHi_333_), .Y(u2__abc_52155_new_n6004_));
AND2X2 AND2X2_1939 ( .A(u2__abc_52155_new_n6006_), .B(u2_o_333_), .Y(u2__abc_52155_new_n6007_));
AND2X2 AND2X2_194 ( .A(_abc_73687_new_n1180_), .B(_abc_73687_new_n1179_), .Y(fracta1_4_));
AND2X2 AND2X2_1940 ( .A(u2__abc_52155_new_n6005_), .B(u2__abc_52155_new_n6008_), .Y(u2__abc_52155_new_n6009_));
AND2X2 AND2X2_1941 ( .A(u2__abc_52155_new_n6002_), .B(u2__abc_52155_new_n6009_), .Y(u2__abc_52155_new_n6010_));
AND2X2 AND2X2_1942 ( .A(u2__abc_52155_new_n6011_), .B(u2_remHi_330_), .Y(u2__abc_52155_new_n6012_));
AND2X2 AND2X2_1943 ( .A(u2__abc_52155_new_n6014_), .B(u2_o_330_), .Y(u2__abc_52155_new_n6015_));
AND2X2 AND2X2_1944 ( .A(u2__abc_52155_new_n6013_), .B(u2__abc_52155_new_n6016_), .Y(u2__abc_52155_new_n6017_));
AND2X2 AND2X2_1945 ( .A(u2__abc_52155_new_n6018_), .B(u2_remHi_331_), .Y(u2__abc_52155_new_n6019_));
AND2X2 AND2X2_1946 ( .A(u2__abc_52155_new_n6021_), .B(u2_o_331_), .Y(u2__abc_52155_new_n6022_));
AND2X2 AND2X2_1947 ( .A(u2__abc_52155_new_n6020_), .B(u2__abc_52155_new_n6023_), .Y(u2__abc_52155_new_n6024_));
AND2X2 AND2X2_1948 ( .A(u2__abc_52155_new_n6017_), .B(u2__abc_52155_new_n6024_), .Y(u2__abc_52155_new_n6025_));
AND2X2 AND2X2_1949 ( .A(u2__abc_52155_new_n6010_), .B(u2__abc_52155_new_n6025_), .Y(u2__abc_52155_new_n6026_));
AND2X2 AND2X2_195 ( .A(_abc_73687_new_n1183_), .B(_abc_73687_new_n1182_), .Y(fracta1_5_));
AND2X2 AND2X2_1950 ( .A(u2__abc_52155_new_n5995_), .B(u2__abc_52155_new_n6026_), .Y(u2__abc_52155_new_n6027_));
AND2X2 AND2X2_1951 ( .A(u2__abc_52155_new_n6028_), .B(u2_o_324_), .Y(u2__abc_52155_new_n6029_));
AND2X2 AND2X2_1952 ( .A(u2__abc_52155_new_n6031_), .B(u2_remHi_324_), .Y(u2__abc_52155_new_n6032_));
AND2X2 AND2X2_1953 ( .A(u2__abc_52155_new_n6030_), .B(u2__abc_52155_new_n6033_), .Y(u2__abc_52155_new_n6034_));
AND2X2 AND2X2_1954 ( .A(u2__abc_52155_new_n6035_), .B(u2_o_325_), .Y(u2__abc_52155_new_n6036_));
AND2X2 AND2X2_1955 ( .A(u2__abc_52155_new_n6038_), .B(u2_remHi_325_), .Y(u2__abc_52155_new_n6039_));
AND2X2 AND2X2_1956 ( .A(u2__abc_52155_new_n6037_), .B(u2__abc_52155_new_n6040_), .Y(u2__abc_52155_new_n6041_));
AND2X2 AND2X2_1957 ( .A(u2__abc_52155_new_n6034_), .B(u2__abc_52155_new_n6041_), .Y(u2__abc_52155_new_n6042_));
AND2X2 AND2X2_1958 ( .A(u2__abc_52155_new_n6043_), .B(u2_remHi_322_), .Y(u2__abc_52155_new_n6044_));
AND2X2 AND2X2_1959 ( .A(u2__abc_52155_new_n6046_), .B(u2_o_322_), .Y(u2__abc_52155_new_n6047_));
AND2X2 AND2X2_196 ( .A(_abc_73687_new_n1186_), .B(_abc_73687_new_n1185_), .Y(fracta1_6_));
AND2X2 AND2X2_1960 ( .A(u2__abc_52155_new_n6045_), .B(u2__abc_52155_new_n6048_), .Y(u2__abc_52155_new_n6049_));
AND2X2 AND2X2_1961 ( .A(u2__abc_52155_new_n6050_), .B(u2_remHi_323_), .Y(u2__abc_52155_new_n6051_));
AND2X2 AND2X2_1962 ( .A(u2__abc_52155_new_n6053_), .B(u2_o_323_), .Y(u2__abc_52155_new_n6054_));
AND2X2 AND2X2_1963 ( .A(u2__abc_52155_new_n6052_), .B(u2__abc_52155_new_n6055_), .Y(u2__abc_52155_new_n6056_));
AND2X2 AND2X2_1964 ( .A(u2__abc_52155_new_n6049_), .B(u2__abc_52155_new_n6056_), .Y(u2__abc_52155_new_n6057_));
AND2X2 AND2X2_1965 ( .A(u2__abc_52155_new_n6042_), .B(u2__abc_52155_new_n6057_), .Y(u2__abc_52155_new_n6058_));
AND2X2 AND2X2_1966 ( .A(u2__abc_52155_new_n6059_), .B(u2_o_318_), .Y(u2__abc_52155_new_n6060_));
AND2X2 AND2X2_1967 ( .A(u2__abc_52155_new_n6062_), .B(u2_remHi_318_), .Y(u2__abc_52155_new_n6063_));
AND2X2 AND2X2_1968 ( .A(u2__abc_52155_new_n6061_), .B(u2__abc_52155_new_n6064_), .Y(u2__abc_52155_new_n6065_));
AND2X2 AND2X2_1969 ( .A(u2__abc_52155_new_n6066_), .B(u2_o_319_), .Y(u2__abc_52155_new_n6067_));
AND2X2 AND2X2_197 ( .A(_abc_73687_new_n1189_), .B(_abc_73687_new_n1188_), .Y(fracta1_7_));
AND2X2 AND2X2_1970 ( .A(u2__abc_52155_new_n6069_), .B(u2_remHi_319_), .Y(u2__abc_52155_new_n6070_));
AND2X2 AND2X2_1971 ( .A(u2__abc_52155_new_n6068_), .B(u2__abc_52155_new_n6071_), .Y(u2__abc_52155_new_n6072_));
AND2X2 AND2X2_1972 ( .A(u2__abc_52155_new_n6065_), .B(u2__abc_52155_new_n6072_), .Y(u2__abc_52155_new_n6073_));
AND2X2 AND2X2_1973 ( .A(u2__abc_52155_new_n6074_), .B(u2_remHi_320_), .Y(u2__abc_52155_new_n6075_));
AND2X2 AND2X2_1974 ( .A(u2__abc_52155_new_n6077_), .B(u2_o_320_), .Y(u2__abc_52155_new_n6078_));
AND2X2 AND2X2_1975 ( .A(u2__abc_52155_new_n6076_), .B(u2__abc_52155_new_n6079_), .Y(u2__abc_52155_new_n6080_));
AND2X2 AND2X2_1976 ( .A(u2__abc_52155_new_n6081_), .B(u2_remHi_321_), .Y(u2__abc_52155_new_n6082_));
AND2X2 AND2X2_1977 ( .A(u2__abc_52155_new_n6084_), .B(u2_o_321_), .Y(u2__abc_52155_new_n6085_));
AND2X2 AND2X2_1978 ( .A(u2__abc_52155_new_n6083_), .B(u2__abc_52155_new_n6086_), .Y(u2__abc_52155_new_n6087_));
AND2X2 AND2X2_1979 ( .A(u2__abc_52155_new_n6080_), .B(u2__abc_52155_new_n6087_), .Y(u2__abc_52155_new_n6088_));
AND2X2 AND2X2_198 ( .A(_abc_73687_new_n1192_), .B(_abc_73687_new_n1191_), .Y(fracta1_8_));
AND2X2 AND2X2_1980 ( .A(u2__abc_52155_new_n6073_), .B(u2__abc_52155_new_n6088_), .Y(u2__abc_52155_new_n6089_));
AND2X2 AND2X2_1981 ( .A(u2__abc_52155_new_n6058_), .B(u2__abc_52155_new_n6089_), .Y(u2__abc_52155_new_n6090_));
AND2X2 AND2X2_1982 ( .A(u2__abc_52155_new_n6027_), .B(u2__abc_52155_new_n6090_), .Y(u2__abc_52155_new_n6091_));
AND2X2 AND2X2_1983 ( .A(u2__abc_52155_new_n5964_), .B(u2__abc_52155_new_n6091_), .Y(u2__abc_52155_new_n6092_));
AND2X2 AND2X2_1984 ( .A(u2__abc_52155_new_n5837_), .B(u2__abc_52155_new_n6092_), .Y(u2__abc_52155_new_n6093_));
AND2X2 AND2X2_1985 ( .A(u2__abc_52155_new_n6094_), .B(u2_remHi_312_), .Y(u2__abc_52155_new_n6095_));
AND2X2 AND2X2_1986 ( .A(u2__abc_52155_new_n6097_), .B(u2_o_312_), .Y(u2__abc_52155_new_n6098_));
AND2X2 AND2X2_1987 ( .A(u2__abc_52155_new_n6096_), .B(u2__abc_52155_new_n6099_), .Y(u2__abc_52155_new_n6100_));
AND2X2 AND2X2_1988 ( .A(u2__abc_52155_new_n6101_), .B(u2_remHi_313_), .Y(u2__abc_52155_new_n6102_));
AND2X2 AND2X2_1989 ( .A(u2__abc_52155_new_n6104_), .B(u2_o_313_), .Y(u2__abc_52155_new_n6105_));
AND2X2 AND2X2_199 ( .A(_abc_73687_new_n1195_), .B(_abc_73687_new_n1194_), .Y(fracta1_9_));
AND2X2 AND2X2_1990 ( .A(u2__abc_52155_new_n6103_), .B(u2__abc_52155_new_n6106_), .Y(u2__abc_52155_new_n6107_));
AND2X2 AND2X2_1991 ( .A(u2__abc_52155_new_n6100_), .B(u2__abc_52155_new_n6107_), .Y(u2__abc_52155_new_n6108_));
AND2X2 AND2X2_1992 ( .A(u2__abc_52155_new_n6109_), .B(u2_remHi_310_), .Y(u2__abc_52155_new_n6110_));
AND2X2 AND2X2_1993 ( .A(u2__abc_52155_new_n6112_), .B(u2_o_310_), .Y(u2__abc_52155_new_n6113_));
AND2X2 AND2X2_1994 ( .A(u2__abc_52155_new_n6111_), .B(u2__abc_52155_new_n6114_), .Y(u2__abc_52155_new_n6115_));
AND2X2 AND2X2_1995 ( .A(u2__abc_52155_new_n6116_), .B(u2_remHi_311_), .Y(u2__abc_52155_new_n6117_));
AND2X2 AND2X2_1996 ( .A(u2__abc_52155_new_n6119_), .B(u2_o_311_), .Y(u2__abc_52155_new_n6120_));
AND2X2 AND2X2_1997 ( .A(u2__abc_52155_new_n6118_), .B(u2__abc_52155_new_n6121_), .Y(u2__abc_52155_new_n6122_));
AND2X2 AND2X2_1998 ( .A(u2__abc_52155_new_n6115_), .B(u2__abc_52155_new_n6122_), .Y(u2__abc_52155_new_n6123_));
AND2X2 AND2X2_1999 ( .A(u2__abc_52155_new_n6108_), .B(u2__abc_52155_new_n6123_), .Y(u2__abc_52155_new_n6124_));
AND2X2 AND2X2_2 ( .A(_abc_73687_new_n753_), .B(sqrto_1_), .Y(\o[37] ));
AND2X2 AND2X2_20 ( .A(_abc_73687_new_n753_), .B(sqrto_19_), .Y(\o[55] ));
AND2X2 AND2X2_200 ( .A(_abc_73687_new_n1198_), .B(_abc_73687_new_n1197_), .Y(fracta1_10_));
AND2X2 AND2X2_2000 ( .A(u2__abc_52155_new_n6125_), .B(u2_remHi_316_), .Y(u2__abc_52155_new_n6126_));
AND2X2 AND2X2_2001 ( .A(u2__abc_52155_new_n6128_), .B(u2_o_316_), .Y(u2__abc_52155_new_n6129_));
AND2X2 AND2X2_2002 ( .A(u2__abc_52155_new_n6127_), .B(u2__abc_52155_new_n6130_), .Y(u2__abc_52155_new_n6131_));
AND2X2 AND2X2_2003 ( .A(u2__abc_52155_new_n6132_), .B(u2_remHi_317_), .Y(u2__abc_52155_new_n6133_));
AND2X2 AND2X2_2004 ( .A(u2__abc_52155_new_n6135_), .B(u2_o_317_), .Y(u2__abc_52155_new_n6136_));
AND2X2 AND2X2_2005 ( .A(u2__abc_52155_new_n6134_), .B(u2__abc_52155_new_n6137_), .Y(u2__abc_52155_new_n6138_));
AND2X2 AND2X2_2006 ( .A(u2__abc_52155_new_n6131_), .B(u2__abc_52155_new_n6138_), .Y(u2__abc_52155_new_n6139_));
AND2X2 AND2X2_2007 ( .A(u2__abc_52155_new_n6140_), .B(u2_remHi_314_), .Y(u2__abc_52155_new_n6141_));
AND2X2 AND2X2_2008 ( .A(u2__abc_52155_new_n6143_), .B(u2_o_314_), .Y(u2__abc_52155_new_n6144_));
AND2X2 AND2X2_2009 ( .A(u2__abc_52155_new_n6142_), .B(u2__abc_52155_new_n6145_), .Y(u2__abc_52155_new_n6146_));
AND2X2 AND2X2_201 ( .A(_abc_73687_new_n1201_), .B(_abc_73687_new_n1200_), .Y(fracta1_11_));
AND2X2 AND2X2_2010 ( .A(u2__abc_52155_new_n6147_), .B(u2_remHi_315_), .Y(u2__abc_52155_new_n6148_));
AND2X2 AND2X2_2011 ( .A(u2__abc_52155_new_n6150_), .B(u2_o_315_), .Y(u2__abc_52155_new_n6151_));
AND2X2 AND2X2_2012 ( .A(u2__abc_52155_new_n6149_), .B(u2__abc_52155_new_n6152_), .Y(u2__abc_52155_new_n6153_));
AND2X2 AND2X2_2013 ( .A(u2__abc_52155_new_n6146_), .B(u2__abc_52155_new_n6153_), .Y(u2__abc_52155_new_n6154_));
AND2X2 AND2X2_2014 ( .A(u2__abc_52155_new_n6139_), .B(u2__abc_52155_new_n6154_), .Y(u2__abc_52155_new_n6155_));
AND2X2 AND2X2_2015 ( .A(u2__abc_52155_new_n6124_), .B(u2__abc_52155_new_n6155_), .Y(u2__abc_52155_new_n6156_));
AND2X2 AND2X2_2016 ( .A(u2__abc_52155_new_n6157_), .B(u2_o_302_), .Y(u2__abc_52155_new_n6158_));
AND2X2 AND2X2_2017 ( .A(u2__abc_52155_new_n6160_), .B(u2_remHi_302_), .Y(u2__abc_52155_new_n6161_));
AND2X2 AND2X2_2018 ( .A(u2__abc_52155_new_n6159_), .B(u2__abc_52155_new_n6162_), .Y(u2__abc_52155_new_n6163_));
AND2X2 AND2X2_2019 ( .A(u2__abc_52155_new_n6164_), .B(u2_o_303_), .Y(u2__abc_52155_new_n6165_));
AND2X2 AND2X2_202 ( .A(_abc_73687_new_n1204_), .B(_abc_73687_new_n1203_), .Y(fracta1_12_));
AND2X2 AND2X2_2020 ( .A(u2__abc_52155_new_n6167_), .B(u2_remHi_303_), .Y(u2__abc_52155_new_n6168_));
AND2X2 AND2X2_2021 ( .A(u2__abc_52155_new_n6166_), .B(u2__abc_52155_new_n6169_), .Y(u2__abc_52155_new_n6170_));
AND2X2 AND2X2_2022 ( .A(u2__abc_52155_new_n6163_), .B(u2__abc_52155_new_n6170_), .Y(u2__abc_52155_new_n6171_));
AND2X2 AND2X2_2023 ( .A(u2__abc_52155_new_n6172_), .B(u2_remHi_304_), .Y(u2__abc_52155_new_n6173_));
AND2X2 AND2X2_2024 ( .A(u2__abc_52155_new_n6175_), .B(u2_o_304_), .Y(u2__abc_52155_new_n6176_));
AND2X2 AND2X2_2025 ( .A(u2__abc_52155_new_n6174_), .B(u2__abc_52155_new_n6177_), .Y(u2__abc_52155_new_n6178_));
AND2X2 AND2X2_2026 ( .A(u2__abc_52155_new_n6179_), .B(u2_remHi_305_), .Y(u2__abc_52155_new_n6180_));
AND2X2 AND2X2_2027 ( .A(u2__abc_52155_new_n6182_), .B(u2_o_305_), .Y(u2__abc_52155_new_n6183_));
AND2X2 AND2X2_2028 ( .A(u2__abc_52155_new_n6181_), .B(u2__abc_52155_new_n6184_), .Y(u2__abc_52155_new_n6185_));
AND2X2 AND2X2_2029 ( .A(u2__abc_52155_new_n6178_), .B(u2__abc_52155_new_n6185_), .Y(u2__abc_52155_new_n6186_));
AND2X2 AND2X2_203 ( .A(_abc_73687_new_n1207_), .B(_abc_73687_new_n1206_), .Y(fracta1_13_));
AND2X2 AND2X2_2030 ( .A(u2__abc_52155_new_n6171_), .B(u2__abc_52155_new_n6186_), .Y(u2__abc_52155_new_n6187_));
AND2X2 AND2X2_2031 ( .A(u2__abc_52155_new_n6188_), .B(u2_remHi_308_), .Y(u2__abc_52155_new_n6189_));
AND2X2 AND2X2_2032 ( .A(u2__abc_52155_new_n6191_), .B(u2_o_308_), .Y(u2__abc_52155_new_n6192_));
AND2X2 AND2X2_2033 ( .A(u2__abc_52155_new_n6190_), .B(u2__abc_52155_new_n6193_), .Y(u2__abc_52155_new_n6194_));
AND2X2 AND2X2_2034 ( .A(u2__abc_52155_new_n6195_), .B(u2_remHi_309_), .Y(u2__abc_52155_new_n6196_));
AND2X2 AND2X2_2035 ( .A(u2__abc_52155_new_n6198_), .B(u2_o_309_), .Y(u2__abc_52155_new_n6199_));
AND2X2 AND2X2_2036 ( .A(u2__abc_52155_new_n6197_), .B(u2__abc_52155_new_n6200_), .Y(u2__abc_52155_new_n6201_));
AND2X2 AND2X2_2037 ( .A(u2__abc_52155_new_n6194_), .B(u2__abc_52155_new_n6201_), .Y(u2__abc_52155_new_n6202_));
AND2X2 AND2X2_2038 ( .A(u2__abc_52155_new_n6203_), .B(u2_remHi_307_), .Y(u2__abc_52155_new_n6204_));
AND2X2 AND2X2_2039 ( .A(u2__abc_52155_new_n6206_), .B(u2_o_307_), .Y(u2__abc_52155_new_n6207_));
AND2X2 AND2X2_204 ( .A(_abc_73687_new_n1210_), .B(_abc_73687_new_n1209_), .Y(fracta1_14_));
AND2X2 AND2X2_2040 ( .A(u2__abc_52155_new_n6205_), .B(u2__abc_52155_new_n6208_), .Y(u2__abc_52155_new_n6209_));
AND2X2 AND2X2_2041 ( .A(u2__abc_52155_new_n6210_), .B(u2_remHi_306_), .Y(u2__abc_52155_new_n6211_));
AND2X2 AND2X2_2042 ( .A(u2__abc_52155_new_n6213_), .B(u2_o_306_), .Y(u2__abc_52155_new_n6214_));
AND2X2 AND2X2_2043 ( .A(u2__abc_52155_new_n6212_), .B(u2__abc_52155_new_n6215_), .Y(u2__abc_52155_new_n6216_));
AND2X2 AND2X2_2044 ( .A(u2__abc_52155_new_n6209_), .B(u2__abc_52155_new_n6216_), .Y(u2__abc_52155_new_n6217_));
AND2X2 AND2X2_2045 ( .A(u2__abc_52155_new_n6202_), .B(u2__abc_52155_new_n6217_), .Y(u2__abc_52155_new_n6218_));
AND2X2 AND2X2_2046 ( .A(u2__abc_52155_new_n6187_), .B(u2__abc_52155_new_n6218_), .Y(u2__abc_52155_new_n6219_));
AND2X2 AND2X2_2047 ( .A(u2__abc_52155_new_n6156_), .B(u2__abc_52155_new_n6219_), .Y(u2__abc_52155_new_n6220_));
AND2X2 AND2X2_2048 ( .A(u2__abc_52155_new_n6221_), .B(u2_o_294_), .Y(u2__abc_52155_new_n6222_));
AND2X2 AND2X2_2049 ( .A(u2__abc_52155_new_n6224_), .B(u2_remHi_294_), .Y(u2__abc_52155_new_n6225_));
AND2X2 AND2X2_205 ( .A(_abc_73687_new_n1213_), .B(_abc_73687_new_n1212_), .Y(fracta1_15_));
AND2X2 AND2X2_2050 ( .A(u2__abc_52155_new_n6223_), .B(u2__abc_52155_new_n6226_), .Y(u2__abc_52155_new_n6227_));
AND2X2 AND2X2_2051 ( .A(u2__abc_52155_new_n6228_), .B(u2_o_295_), .Y(u2__abc_52155_new_n6229_));
AND2X2 AND2X2_2052 ( .A(u2__abc_52155_new_n6231_), .B(u2_remHi_295_), .Y(u2__abc_52155_new_n6232_));
AND2X2 AND2X2_2053 ( .A(u2__abc_52155_new_n6230_), .B(u2__abc_52155_new_n6233_), .Y(u2__abc_52155_new_n6234_));
AND2X2 AND2X2_2054 ( .A(u2__abc_52155_new_n6227_), .B(u2__abc_52155_new_n6234_), .Y(u2__abc_52155_new_n6235_));
AND2X2 AND2X2_2055 ( .A(u2__abc_52155_new_n6236_), .B(u2_remHi_296_), .Y(u2__abc_52155_new_n6237_));
AND2X2 AND2X2_2056 ( .A(u2__abc_52155_new_n6239_), .B(u2_o_296_), .Y(u2__abc_52155_new_n6240_));
AND2X2 AND2X2_2057 ( .A(u2__abc_52155_new_n6238_), .B(u2__abc_52155_new_n6241_), .Y(u2__abc_52155_new_n6242_));
AND2X2 AND2X2_2058 ( .A(u2__abc_52155_new_n6243_), .B(u2_remHi_297_), .Y(u2__abc_52155_new_n6244_));
AND2X2 AND2X2_2059 ( .A(u2__abc_52155_new_n6246_), .B(u2_o_297_), .Y(u2__abc_52155_new_n6247_));
AND2X2 AND2X2_206 ( .A(_abc_73687_new_n1216_), .B(_abc_73687_new_n1215_), .Y(fracta1_16_));
AND2X2 AND2X2_2060 ( .A(u2__abc_52155_new_n6245_), .B(u2__abc_52155_new_n6248_), .Y(u2__abc_52155_new_n6249_));
AND2X2 AND2X2_2061 ( .A(u2__abc_52155_new_n6242_), .B(u2__abc_52155_new_n6249_), .Y(u2__abc_52155_new_n6250_));
AND2X2 AND2X2_2062 ( .A(u2__abc_52155_new_n6235_), .B(u2__abc_52155_new_n6250_), .Y(u2__abc_52155_new_n6251_));
AND2X2 AND2X2_2063 ( .A(u2__abc_52155_new_n6252_), .B(u2_remHi_300_), .Y(u2__abc_52155_new_n6253_));
AND2X2 AND2X2_2064 ( .A(u2__abc_52155_new_n6255_), .B(u2_o_300_), .Y(u2__abc_52155_new_n6256_));
AND2X2 AND2X2_2065 ( .A(u2__abc_52155_new_n6254_), .B(u2__abc_52155_new_n6257_), .Y(u2__abc_52155_new_n6258_));
AND2X2 AND2X2_2066 ( .A(u2__abc_52155_new_n6259_), .B(u2_remHi_301_), .Y(u2__abc_52155_new_n6260_));
AND2X2 AND2X2_2067 ( .A(u2__abc_52155_new_n6262_), .B(u2_o_301_), .Y(u2__abc_52155_new_n6263_));
AND2X2 AND2X2_2068 ( .A(u2__abc_52155_new_n6261_), .B(u2__abc_52155_new_n6264_), .Y(u2__abc_52155_new_n6265_));
AND2X2 AND2X2_2069 ( .A(u2__abc_52155_new_n6258_), .B(u2__abc_52155_new_n6265_), .Y(u2__abc_52155_new_n6266_));
AND2X2 AND2X2_207 ( .A(_abc_73687_new_n1219_), .B(_abc_73687_new_n1218_), .Y(fracta1_17_));
AND2X2 AND2X2_2070 ( .A(u2__abc_52155_new_n6267_), .B(u2_remHi_298_), .Y(u2__abc_52155_new_n6268_));
AND2X2 AND2X2_2071 ( .A(u2__abc_52155_new_n6270_), .B(u2_o_298_), .Y(u2__abc_52155_new_n6271_));
AND2X2 AND2X2_2072 ( .A(u2__abc_52155_new_n6269_), .B(u2__abc_52155_new_n6272_), .Y(u2__abc_52155_new_n6273_));
AND2X2 AND2X2_2073 ( .A(u2__abc_52155_new_n6274_), .B(u2_remHi_299_), .Y(u2__abc_52155_new_n6275_));
AND2X2 AND2X2_2074 ( .A(u2__abc_52155_new_n6277_), .B(u2_o_299_), .Y(u2__abc_52155_new_n6278_));
AND2X2 AND2X2_2075 ( .A(u2__abc_52155_new_n6276_), .B(u2__abc_52155_new_n6279_), .Y(u2__abc_52155_new_n6280_));
AND2X2 AND2X2_2076 ( .A(u2__abc_52155_new_n6273_), .B(u2__abc_52155_new_n6280_), .Y(u2__abc_52155_new_n6281_));
AND2X2 AND2X2_2077 ( .A(u2__abc_52155_new_n6266_), .B(u2__abc_52155_new_n6281_), .Y(u2__abc_52155_new_n6282_));
AND2X2 AND2X2_2078 ( .A(u2__abc_52155_new_n6251_), .B(u2__abc_52155_new_n6282_), .Y(u2__abc_52155_new_n6283_));
AND2X2 AND2X2_2079 ( .A(u2__abc_52155_new_n6284_), .B(u2_remHi_288_), .Y(u2__abc_52155_new_n6285_));
AND2X2 AND2X2_208 ( .A(_abc_73687_new_n1222_), .B(_abc_73687_new_n1221_), .Y(fracta1_18_));
AND2X2 AND2X2_2080 ( .A(u2__abc_52155_new_n6287_), .B(u2_o_288_), .Y(u2__abc_52155_new_n6288_));
AND2X2 AND2X2_2081 ( .A(u2__abc_52155_new_n6286_), .B(u2__abc_52155_new_n6289_), .Y(u2__abc_52155_new_n6290_));
AND2X2 AND2X2_2082 ( .A(u2__abc_52155_new_n6291_), .B(u2_remHi_289_), .Y(u2__abc_52155_new_n6292_));
AND2X2 AND2X2_2083 ( .A(u2__abc_52155_new_n6294_), .B(u2_o_289_), .Y(u2__abc_52155_new_n6295_));
AND2X2 AND2X2_2084 ( .A(u2__abc_52155_new_n6293_), .B(u2__abc_52155_new_n6296_), .Y(u2__abc_52155_new_n6297_));
AND2X2 AND2X2_2085 ( .A(u2__abc_52155_new_n6290_), .B(u2__abc_52155_new_n6297_), .Y(u2__abc_52155_new_n6298_));
AND2X2 AND2X2_2086 ( .A(u2__abc_52155_new_n6299_), .B(u2_remHi_286_), .Y(u2__abc_52155_new_n6300_));
AND2X2 AND2X2_2087 ( .A(u2__abc_52155_new_n6302_), .B(u2_o_286_), .Y(u2__abc_52155_new_n6303_));
AND2X2 AND2X2_2088 ( .A(u2__abc_52155_new_n6301_), .B(u2__abc_52155_new_n6304_), .Y(u2__abc_52155_new_n6305_));
AND2X2 AND2X2_2089 ( .A(u2__abc_52155_new_n6306_), .B(u2_remHi_287_), .Y(u2__abc_52155_new_n6307_));
AND2X2 AND2X2_209 ( .A(_abc_73687_new_n1225_), .B(_abc_73687_new_n1224_), .Y(fracta1_19_));
AND2X2 AND2X2_2090 ( .A(u2__abc_52155_new_n6309_), .B(u2_o_287_), .Y(u2__abc_52155_new_n6310_));
AND2X2 AND2X2_2091 ( .A(u2__abc_52155_new_n6308_), .B(u2__abc_52155_new_n6311_), .Y(u2__abc_52155_new_n6312_));
AND2X2 AND2X2_2092 ( .A(u2__abc_52155_new_n6305_), .B(u2__abc_52155_new_n6312_), .Y(u2__abc_52155_new_n6313_));
AND2X2 AND2X2_2093 ( .A(u2__abc_52155_new_n6298_), .B(u2__abc_52155_new_n6313_), .Y(u2__abc_52155_new_n6314_));
AND2X2 AND2X2_2094 ( .A(u2__abc_52155_new_n6315_), .B(u2_remHi_292_), .Y(u2__abc_52155_new_n6316_));
AND2X2 AND2X2_2095 ( .A(u2__abc_52155_new_n6318_), .B(u2_o_292_), .Y(u2__abc_52155_new_n6319_));
AND2X2 AND2X2_2096 ( .A(u2__abc_52155_new_n6317_), .B(u2__abc_52155_new_n6320_), .Y(u2__abc_52155_new_n6321_));
AND2X2 AND2X2_2097 ( .A(u2__abc_52155_new_n6322_), .B(u2_remHi_293_), .Y(u2__abc_52155_new_n6323_));
AND2X2 AND2X2_2098 ( .A(u2__abc_52155_new_n6325_), .B(u2_o_293_), .Y(u2__abc_52155_new_n6326_));
AND2X2 AND2X2_2099 ( .A(u2__abc_52155_new_n6324_), .B(u2__abc_52155_new_n6327_), .Y(u2__abc_52155_new_n6328_));
AND2X2 AND2X2_21 ( .A(_abc_73687_new_n753_), .B(sqrto_20_), .Y(\o[56] ));
AND2X2 AND2X2_210 ( .A(_abc_73687_new_n1228_), .B(_abc_73687_new_n1227_), .Y(fracta1_20_));
AND2X2 AND2X2_2100 ( .A(u2__abc_52155_new_n6321_), .B(u2__abc_52155_new_n6328_), .Y(u2__abc_52155_new_n6329_));
AND2X2 AND2X2_2101 ( .A(u2__abc_52155_new_n6330_), .B(u2_remHi_290_), .Y(u2__abc_52155_new_n6331_));
AND2X2 AND2X2_2102 ( .A(u2__abc_52155_new_n6333_), .B(u2_o_290_), .Y(u2__abc_52155_new_n6334_));
AND2X2 AND2X2_2103 ( .A(u2__abc_52155_new_n6332_), .B(u2__abc_52155_new_n6335_), .Y(u2__abc_52155_new_n6336_));
AND2X2 AND2X2_2104 ( .A(u2__abc_52155_new_n6337_), .B(u2_remHi_291_), .Y(u2__abc_52155_new_n6338_));
AND2X2 AND2X2_2105 ( .A(u2__abc_52155_new_n6340_), .B(u2_o_291_), .Y(u2__abc_52155_new_n6341_));
AND2X2 AND2X2_2106 ( .A(u2__abc_52155_new_n6339_), .B(u2__abc_52155_new_n6342_), .Y(u2__abc_52155_new_n6343_));
AND2X2 AND2X2_2107 ( .A(u2__abc_52155_new_n6336_), .B(u2__abc_52155_new_n6343_), .Y(u2__abc_52155_new_n6344_));
AND2X2 AND2X2_2108 ( .A(u2__abc_52155_new_n6329_), .B(u2__abc_52155_new_n6344_), .Y(u2__abc_52155_new_n6345_));
AND2X2 AND2X2_2109 ( .A(u2__abc_52155_new_n6314_), .B(u2__abc_52155_new_n6345_), .Y(u2__abc_52155_new_n6346_));
AND2X2 AND2X2_211 ( .A(_abc_73687_new_n1231_), .B(_abc_73687_new_n1230_), .Y(fracta1_21_));
AND2X2 AND2X2_2110 ( .A(u2__abc_52155_new_n6283_), .B(u2__abc_52155_new_n6346_), .Y(u2__abc_52155_new_n6347_));
AND2X2 AND2X2_2111 ( .A(u2__abc_52155_new_n6220_), .B(u2__abc_52155_new_n6347_), .Y(u2__abc_52155_new_n6348_));
AND2X2 AND2X2_2112 ( .A(u2__abc_52155_new_n6349_), .B(u2_remHi_280_), .Y(u2__abc_52155_new_n6350_));
AND2X2 AND2X2_2113 ( .A(u2__abc_52155_new_n6352_), .B(u2_o_280_), .Y(u2__abc_52155_new_n6353_));
AND2X2 AND2X2_2114 ( .A(u2__abc_52155_new_n6351_), .B(u2__abc_52155_new_n6354_), .Y(u2__abc_52155_new_n6355_));
AND2X2 AND2X2_2115 ( .A(u2__abc_52155_new_n6356_), .B(u2_remHi_281_), .Y(u2__abc_52155_new_n6357_));
AND2X2 AND2X2_2116 ( .A(u2__abc_52155_new_n6359_), .B(u2_o_281_), .Y(u2__abc_52155_new_n6360_));
AND2X2 AND2X2_2117 ( .A(u2__abc_52155_new_n6358_), .B(u2__abc_52155_new_n6361_), .Y(u2__abc_52155_new_n6362_));
AND2X2 AND2X2_2118 ( .A(u2__abc_52155_new_n6355_), .B(u2__abc_52155_new_n6362_), .Y(u2__abc_52155_new_n6363_));
AND2X2 AND2X2_2119 ( .A(u2__abc_52155_new_n6364_), .B(u2_remHi_278_), .Y(u2__abc_52155_new_n6365_));
AND2X2 AND2X2_212 ( .A(_abc_73687_new_n1234_), .B(_abc_73687_new_n1233_), .Y(fracta1_22_));
AND2X2 AND2X2_2120 ( .A(u2__abc_52155_new_n6367_), .B(u2_o_278_), .Y(u2__abc_52155_new_n6368_));
AND2X2 AND2X2_2121 ( .A(u2__abc_52155_new_n6366_), .B(u2__abc_52155_new_n6369_), .Y(u2__abc_52155_new_n6370_));
AND2X2 AND2X2_2122 ( .A(u2__abc_52155_new_n6371_), .B(u2_remHi_279_), .Y(u2__abc_52155_new_n6372_));
AND2X2 AND2X2_2123 ( .A(u2__abc_52155_new_n6374_), .B(u2_o_279_), .Y(u2__abc_52155_new_n6375_));
AND2X2 AND2X2_2124 ( .A(u2__abc_52155_new_n6373_), .B(u2__abc_52155_new_n6376_), .Y(u2__abc_52155_new_n6377_));
AND2X2 AND2X2_2125 ( .A(u2__abc_52155_new_n6370_), .B(u2__abc_52155_new_n6377_), .Y(u2__abc_52155_new_n6378_));
AND2X2 AND2X2_2126 ( .A(u2__abc_52155_new_n6363_), .B(u2__abc_52155_new_n6378_), .Y(u2__abc_52155_new_n6379_));
AND2X2 AND2X2_2127 ( .A(u2__abc_52155_new_n6380_), .B(u2_remHi_284_), .Y(u2__abc_52155_new_n6381_));
AND2X2 AND2X2_2128 ( .A(u2__abc_52155_new_n6383_), .B(u2_o_284_), .Y(u2__abc_52155_new_n6384_));
AND2X2 AND2X2_2129 ( .A(u2__abc_52155_new_n6382_), .B(u2__abc_52155_new_n6385_), .Y(u2__abc_52155_new_n6386_));
AND2X2 AND2X2_213 ( .A(_abc_73687_new_n1237_), .B(_abc_73687_new_n1236_), .Y(fracta1_23_));
AND2X2 AND2X2_2130 ( .A(u2__abc_52155_new_n6387_), .B(u2_remHi_285_), .Y(u2__abc_52155_new_n6388_));
AND2X2 AND2X2_2131 ( .A(u2__abc_52155_new_n6390_), .B(u2_o_285_), .Y(u2__abc_52155_new_n6391_));
AND2X2 AND2X2_2132 ( .A(u2__abc_52155_new_n6389_), .B(u2__abc_52155_new_n6392_), .Y(u2__abc_52155_new_n6393_));
AND2X2 AND2X2_2133 ( .A(u2__abc_52155_new_n6386_), .B(u2__abc_52155_new_n6393_), .Y(u2__abc_52155_new_n6394_));
AND2X2 AND2X2_2134 ( .A(u2__abc_52155_new_n6395_), .B(u2_remHi_282_), .Y(u2__abc_52155_new_n6396_));
AND2X2 AND2X2_2135 ( .A(u2__abc_52155_new_n6398_), .B(u2_o_282_), .Y(u2__abc_52155_new_n6399_));
AND2X2 AND2X2_2136 ( .A(u2__abc_52155_new_n6397_), .B(u2__abc_52155_new_n6400_), .Y(u2__abc_52155_new_n6401_));
AND2X2 AND2X2_2137 ( .A(u2__abc_52155_new_n6402_), .B(u2_remHi_283_), .Y(u2__abc_52155_new_n6403_));
AND2X2 AND2X2_2138 ( .A(u2__abc_52155_new_n6405_), .B(u2_o_283_), .Y(u2__abc_52155_new_n6406_));
AND2X2 AND2X2_2139 ( .A(u2__abc_52155_new_n6404_), .B(u2__abc_52155_new_n6407_), .Y(u2__abc_52155_new_n6408_));
AND2X2 AND2X2_214 ( .A(_abc_73687_new_n1240_), .B(_abc_73687_new_n1239_), .Y(fracta1_24_));
AND2X2 AND2X2_2140 ( .A(u2__abc_52155_new_n6401_), .B(u2__abc_52155_new_n6408_), .Y(u2__abc_52155_new_n6409_));
AND2X2 AND2X2_2141 ( .A(u2__abc_52155_new_n6394_), .B(u2__abc_52155_new_n6409_), .Y(u2__abc_52155_new_n6410_));
AND2X2 AND2X2_2142 ( .A(u2__abc_52155_new_n6379_), .B(u2__abc_52155_new_n6410_), .Y(u2__abc_52155_new_n6411_));
AND2X2 AND2X2_2143 ( .A(u2__abc_52155_new_n6412_), .B(u2_remHi_272_), .Y(u2__abc_52155_new_n6413_));
AND2X2 AND2X2_2144 ( .A(u2__abc_52155_new_n6415_), .B(u2_o_272_), .Y(u2__abc_52155_new_n6416_));
AND2X2 AND2X2_2145 ( .A(u2__abc_52155_new_n6414_), .B(u2__abc_52155_new_n6417_), .Y(u2__abc_52155_new_n6418_));
AND2X2 AND2X2_2146 ( .A(u2__abc_52155_new_n6419_), .B(u2_remHi_273_), .Y(u2__abc_52155_new_n6420_));
AND2X2 AND2X2_2147 ( .A(u2__abc_52155_new_n6422_), .B(u2_o_273_), .Y(u2__abc_52155_new_n6423_));
AND2X2 AND2X2_2148 ( .A(u2__abc_52155_new_n6421_), .B(u2__abc_52155_new_n6424_), .Y(u2__abc_52155_new_n6425_));
AND2X2 AND2X2_2149 ( .A(u2__abc_52155_new_n6418_), .B(u2__abc_52155_new_n6425_), .Y(u2__abc_52155_new_n6426_));
AND2X2 AND2X2_215 ( .A(_abc_73687_new_n1243_), .B(_abc_73687_new_n1242_), .Y(fracta1_25_));
AND2X2 AND2X2_2150 ( .A(u2__abc_52155_new_n6427_), .B(u2_remHi_270_), .Y(u2__abc_52155_new_n6428_));
AND2X2 AND2X2_2151 ( .A(u2__abc_52155_new_n6430_), .B(u2_o_270_), .Y(u2__abc_52155_new_n6431_));
AND2X2 AND2X2_2152 ( .A(u2__abc_52155_new_n6429_), .B(u2__abc_52155_new_n6432_), .Y(u2__abc_52155_new_n6433_));
AND2X2 AND2X2_2153 ( .A(u2__abc_52155_new_n6434_), .B(u2_remHi_271_), .Y(u2__abc_52155_new_n6435_));
AND2X2 AND2X2_2154 ( .A(u2__abc_52155_new_n6437_), .B(u2_o_271_), .Y(u2__abc_52155_new_n6438_));
AND2X2 AND2X2_2155 ( .A(u2__abc_52155_new_n6436_), .B(u2__abc_52155_new_n6439_), .Y(u2__abc_52155_new_n6440_));
AND2X2 AND2X2_2156 ( .A(u2__abc_52155_new_n6433_), .B(u2__abc_52155_new_n6440_), .Y(u2__abc_52155_new_n6441_));
AND2X2 AND2X2_2157 ( .A(u2__abc_52155_new_n6426_), .B(u2__abc_52155_new_n6441_), .Y(u2__abc_52155_new_n6442_));
AND2X2 AND2X2_2158 ( .A(u2__abc_52155_new_n6443_), .B(u2_remHi_276_), .Y(u2__abc_52155_new_n6444_));
AND2X2 AND2X2_2159 ( .A(u2__abc_52155_new_n6446_), .B(u2_o_276_), .Y(u2__abc_52155_new_n6447_));
AND2X2 AND2X2_216 ( .A(_abc_73687_new_n1246_), .B(_abc_73687_new_n1245_), .Y(fracta1_26_));
AND2X2 AND2X2_2160 ( .A(u2__abc_52155_new_n6445_), .B(u2__abc_52155_new_n6448_), .Y(u2__abc_52155_new_n6449_));
AND2X2 AND2X2_2161 ( .A(u2__abc_52155_new_n6450_), .B(u2_remHi_277_), .Y(u2__abc_52155_new_n6451_));
AND2X2 AND2X2_2162 ( .A(u2__abc_52155_new_n6453_), .B(u2_o_277_), .Y(u2__abc_52155_new_n6454_));
AND2X2 AND2X2_2163 ( .A(u2__abc_52155_new_n6452_), .B(u2__abc_52155_new_n6455_), .Y(u2__abc_52155_new_n6456_));
AND2X2 AND2X2_2164 ( .A(u2__abc_52155_new_n6449_), .B(u2__abc_52155_new_n6456_), .Y(u2__abc_52155_new_n6457_));
AND2X2 AND2X2_2165 ( .A(u2__abc_52155_new_n6458_), .B(u2_remHi_274_), .Y(u2__abc_52155_new_n6459_));
AND2X2 AND2X2_2166 ( .A(u2__abc_52155_new_n6461_), .B(u2_o_274_), .Y(u2__abc_52155_new_n6462_));
AND2X2 AND2X2_2167 ( .A(u2__abc_52155_new_n6460_), .B(u2__abc_52155_new_n6463_), .Y(u2__abc_52155_new_n6464_));
AND2X2 AND2X2_2168 ( .A(u2__abc_52155_new_n6465_), .B(u2_remHi_275_), .Y(u2__abc_52155_new_n6466_));
AND2X2 AND2X2_2169 ( .A(u2__abc_52155_new_n6468_), .B(u2_o_275_), .Y(u2__abc_52155_new_n6469_));
AND2X2 AND2X2_217 ( .A(_abc_73687_new_n1249_), .B(_abc_73687_new_n1248_), .Y(fracta1_27_));
AND2X2 AND2X2_2170 ( .A(u2__abc_52155_new_n6467_), .B(u2__abc_52155_new_n6470_), .Y(u2__abc_52155_new_n6471_));
AND2X2 AND2X2_2171 ( .A(u2__abc_52155_new_n6464_), .B(u2__abc_52155_new_n6471_), .Y(u2__abc_52155_new_n6472_));
AND2X2 AND2X2_2172 ( .A(u2__abc_52155_new_n6457_), .B(u2__abc_52155_new_n6472_), .Y(u2__abc_52155_new_n6473_));
AND2X2 AND2X2_2173 ( .A(u2__abc_52155_new_n6442_), .B(u2__abc_52155_new_n6473_), .Y(u2__abc_52155_new_n6474_));
AND2X2 AND2X2_2174 ( .A(u2__abc_52155_new_n6411_), .B(u2__abc_52155_new_n6474_), .Y(u2__abc_52155_new_n6475_));
AND2X2 AND2X2_2175 ( .A(u2__abc_52155_new_n6476_), .B(u2_o_268_), .Y(u2__abc_52155_new_n6477_));
AND2X2 AND2X2_2176 ( .A(u2__abc_52155_new_n6479_), .B(u2_remHi_268_), .Y(u2__abc_52155_new_n6480_));
AND2X2 AND2X2_2177 ( .A(u2__abc_52155_new_n6478_), .B(u2__abc_52155_new_n6481_), .Y(u2__abc_52155_new_n6482_));
AND2X2 AND2X2_2178 ( .A(u2__abc_52155_new_n6483_), .B(u2_o_269_), .Y(u2__abc_52155_new_n6484_));
AND2X2 AND2X2_2179 ( .A(u2__abc_52155_new_n6486_), .B(u2_remHi_269_), .Y(u2__abc_52155_new_n6487_));
AND2X2 AND2X2_218 ( .A(_abc_73687_new_n1252_), .B(_abc_73687_new_n1251_), .Y(fracta1_28_));
AND2X2 AND2X2_2180 ( .A(u2__abc_52155_new_n6485_), .B(u2__abc_52155_new_n6488_), .Y(u2__abc_52155_new_n6489_));
AND2X2 AND2X2_2181 ( .A(u2__abc_52155_new_n6482_), .B(u2__abc_52155_new_n6489_), .Y(u2__abc_52155_new_n6490_));
AND2X2 AND2X2_2182 ( .A(u2__abc_52155_new_n6491_), .B(u2_remHi_266_), .Y(u2__abc_52155_new_n6492_));
AND2X2 AND2X2_2183 ( .A(u2__abc_52155_new_n6494_), .B(u2_o_266_), .Y(u2__abc_52155_new_n6495_));
AND2X2 AND2X2_2184 ( .A(u2__abc_52155_new_n6493_), .B(u2__abc_52155_new_n6496_), .Y(u2__abc_52155_new_n6497_));
AND2X2 AND2X2_2185 ( .A(u2__abc_52155_new_n6498_), .B(u2_remHi_267_), .Y(u2__abc_52155_new_n6499_));
AND2X2 AND2X2_2186 ( .A(u2__abc_52155_new_n6501_), .B(u2_o_267_), .Y(u2__abc_52155_new_n6502_));
AND2X2 AND2X2_2187 ( .A(u2__abc_52155_new_n6500_), .B(u2__abc_52155_new_n6503_), .Y(u2__abc_52155_new_n6504_));
AND2X2 AND2X2_2188 ( .A(u2__abc_52155_new_n6497_), .B(u2__abc_52155_new_n6504_), .Y(u2__abc_52155_new_n6505_));
AND2X2 AND2X2_2189 ( .A(u2__abc_52155_new_n6490_), .B(u2__abc_52155_new_n6505_), .Y(u2__abc_52155_new_n6506_));
AND2X2 AND2X2_219 ( .A(_abc_73687_new_n1255_), .B(_abc_73687_new_n1254_), .Y(fracta1_29_));
AND2X2 AND2X2_2190 ( .A(u2__abc_52155_new_n6507_), .B(u2_remHi_264_), .Y(u2__abc_52155_new_n6508_));
AND2X2 AND2X2_2191 ( .A(u2__abc_52155_new_n6510_), .B(u2_o_264_), .Y(u2__abc_52155_new_n6511_));
AND2X2 AND2X2_2192 ( .A(u2__abc_52155_new_n6509_), .B(u2__abc_52155_new_n6512_), .Y(u2__abc_52155_new_n6513_));
AND2X2 AND2X2_2193 ( .A(u2__abc_52155_new_n6514_), .B(u2_remHi_265_), .Y(u2__abc_52155_new_n6515_));
AND2X2 AND2X2_2194 ( .A(u2__abc_52155_new_n6517_), .B(u2_o_265_), .Y(u2__abc_52155_new_n6518_));
AND2X2 AND2X2_2195 ( .A(u2__abc_52155_new_n6516_), .B(u2__abc_52155_new_n6519_), .Y(u2__abc_52155_new_n6520_));
AND2X2 AND2X2_2196 ( .A(u2__abc_52155_new_n6513_), .B(u2__abc_52155_new_n6520_), .Y(u2__abc_52155_new_n6521_));
AND2X2 AND2X2_2197 ( .A(u2__abc_52155_new_n6522_), .B(u2_o_262_), .Y(u2__abc_52155_new_n6523_));
AND2X2 AND2X2_2198 ( .A(u2__abc_52155_new_n6525_), .B(u2_remHi_262_), .Y(u2__abc_52155_new_n6526_));
AND2X2 AND2X2_2199 ( .A(u2__abc_52155_new_n6524_), .B(u2__abc_52155_new_n6527_), .Y(u2__abc_52155_new_n6528_));
AND2X2 AND2X2_22 ( .A(_abc_73687_new_n753_), .B(sqrto_21_), .Y(\o[57] ));
AND2X2 AND2X2_220 ( .A(_abc_73687_new_n1258_), .B(_abc_73687_new_n1257_), .Y(fracta1_30_));
AND2X2 AND2X2_2200 ( .A(u2__abc_52155_new_n6529_), .B(u2_o_263_), .Y(u2__abc_52155_new_n6530_));
AND2X2 AND2X2_2201 ( .A(u2__abc_52155_new_n6532_), .B(u2_remHi_263_), .Y(u2__abc_52155_new_n6533_));
AND2X2 AND2X2_2202 ( .A(u2__abc_52155_new_n6531_), .B(u2__abc_52155_new_n6534_), .Y(u2__abc_52155_new_n6535_));
AND2X2 AND2X2_2203 ( .A(u2__abc_52155_new_n6528_), .B(u2__abc_52155_new_n6535_), .Y(u2__abc_52155_new_n6536_));
AND2X2 AND2X2_2204 ( .A(u2__abc_52155_new_n6521_), .B(u2__abc_52155_new_n6536_), .Y(u2__abc_52155_new_n6537_));
AND2X2 AND2X2_2205 ( .A(u2__abc_52155_new_n6506_), .B(u2__abc_52155_new_n6537_), .Y(u2__abc_52155_new_n6538_));
AND2X2 AND2X2_2206 ( .A(u2__abc_52155_new_n6539_), .B(u2_o_254_), .Y(u2__abc_52155_new_n6540_));
AND2X2 AND2X2_2207 ( .A(u2__abc_52155_new_n6542_), .B(u2_remHi_254_), .Y(u2__abc_52155_new_n6543_));
AND2X2 AND2X2_2208 ( .A(u2__abc_52155_new_n6541_), .B(u2__abc_52155_new_n6544_), .Y(u2__abc_52155_new_n6545_));
AND2X2 AND2X2_2209 ( .A(u2__abc_52155_new_n6546_), .B(u2_o_255_), .Y(u2__abc_52155_new_n6547_));
AND2X2 AND2X2_221 ( .A(_abc_73687_new_n1261_), .B(_abc_73687_new_n1260_), .Y(fracta1_31_));
AND2X2 AND2X2_2210 ( .A(u2__abc_52155_new_n6549_), .B(u2_remHi_255_), .Y(u2__abc_52155_new_n6550_));
AND2X2 AND2X2_2211 ( .A(u2__abc_52155_new_n6548_), .B(u2__abc_52155_new_n6551_), .Y(u2__abc_52155_new_n6552_));
AND2X2 AND2X2_2212 ( .A(u2__abc_52155_new_n6545_), .B(u2__abc_52155_new_n6552_), .Y(u2__abc_52155_new_n6553_));
AND2X2 AND2X2_2213 ( .A(u2__abc_52155_new_n6554_), .B(u2_remHi_256_), .Y(u2__abc_52155_new_n6555_));
AND2X2 AND2X2_2214 ( .A(u2__abc_52155_new_n6557_), .B(u2_o_256_), .Y(u2__abc_52155_new_n6558_));
AND2X2 AND2X2_2215 ( .A(u2__abc_52155_new_n6556_), .B(u2__abc_52155_new_n6559_), .Y(u2__abc_52155_new_n6560_));
AND2X2 AND2X2_2216 ( .A(u2__abc_52155_new_n6561_), .B(u2_remHi_257_), .Y(u2__abc_52155_new_n6562_));
AND2X2 AND2X2_2217 ( .A(u2__abc_52155_new_n6564_), .B(u2_o_257_), .Y(u2__abc_52155_new_n6565_));
AND2X2 AND2X2_2218 ( .A(u2__abc_52155_new_n6563_), .B(u2__abc_52155_new_n6566_), .Y(u2__abc_52155_new_n6567_));
AND2X2 AND2X2_2219 ( .A(u2__abc_52155_new_n6560_), .B(u2__abc_52155_new_n6567_), .Y(u2__abc_52155_new_n6568_));
AND2X2 AND2X2_222 ( .A(_abc_73687_new_n1264_), .B(_abc_73687_new_n1263_), .Y(fracta1_32_));
AND2X2 AND2X2_2220 ( .A(u2__abc_52155_new_n6553_), .B(u2__abc_52155_new_n6568_), .Y(u2__abc_52155_new_n6569_));
AND2X2 AND2X2_2221 ( .A(u2__abc_52155_new_n6570_), .B(u2_remHi_260_), .Y(u2__abc_52155_new_n6571_));
AND2X2 AND2X2_2222 ( .A(u2__abc_52155_new_n6573_), .B(u2_o_260_), .Y(u2__abc_52155_new_n6574_));
AND2X2 AND2X2_2223 ( .A(u2__abc_52155_new_n6572_), .B(u2__abc_52155_new_n6575_), .Y(u2__abc_52155_new_n6576_));
AND2X2 AND2X2_2224 ( .A(u2__abc_52155_new_n6577_), .B(u2_remHi_261_), .Y(u2__abc_52155_new_n6578_));
AND2X2 AND2X2_2225 ( .A(u2__abc_52155_new_n6580_), .B(u2_o_261_), .Y(u2__abc_52155_new_n6581_));
AND2X2 AND2X2_2226 ( .A(u2__abc_52155_new_n6579_), .B(u2__abc_52155_new_n6582_), .Y(u2__abc_52155_new_n6583_));
AND2X2 AND2X2_2227 ( .A(u2__abc_52155_new_n6576_), .B(u2__abc_52155_new_n6583_), .Y(u2__abc_52155_new_n6584_));
AND2X2 AND2X2_2228 ( .A(u2__abc_52155_new_n6585_), .B(u2_remHi_258_), .Y(u2__abc_52155_new_n6586_));
AND2X2 AND2X2_2229 ( .A(u2__abc_52155_new_n6588_), .B(u2_o_258_), .Y(u2__abc_52155_new_n6589_));
AND2X2 AND2X2_223 ( .A(_abc_73687_new_n1267_), .B(_abc_73687_new_n1266_), .Y(fracta1_33_));
AND2X2 AND2X2_2230 ( .A(u2__abc_52155_new_n6587_), .B(u2__abc_52155_new_n6590_), .Y(u2__abc_52155_new_n6591_));
AND2X2 AND2X2_2231 ( .A(u2__abc_52155_new_n6592_), .B(u2_remHi_259_), .Y(u2__abc_52155_new_n6593_));
AND2X2 AND2X2_2232 ( .A(u2__abc_52155_new_n6595_), .B(u2_o_259_), .Y(u2__abc_52155_new_n6596_));
AND2X2 AND2X2_2233 ( .A(u2__abc_52155_new_n6594_), .B(u2__abc_52155_new_n6597_), .Y(u2__abc_52155_new_n6598_));
AND2X2 AND2X2_2234 ( .A(u2__abc_52155_new_n6591_), .B(u2__abc_52155_new_n6598_), .Y(u2__abc_52155_new_n6599_));
AND2X2 AND2X2_2235 ( .A(u2__abc_52155_new_n6584_), .B(u2__abc_52155_new_n6599_), .Y(u2__abc_52155_new_n6600_));
AND2X2 AND2X2_2236 ( .A(u2__abc_52155_new_n6569_), .B(u2__abc_52155_new_n6600_), .Y(u2__abc_52155_new_n6601_));
AND2X2 AND2X2_2237 ( .A(u2__abc_52155_new_n6538_), .B(u2__abc_52155_new_n6601_), .Y(u2__abc_52155_new_n6602_));
AND2X2 AND2X2_2238 ( .A(u2__abc_52155_new_n6475_), .B(u2__abc_52155_new_n6602_), .Y(u2__abc_52155_new_n6603_));
AND2X2 AND2X2_2239 ( .A(u2__abc_52155_new_n6348_), .B(u2__abc_52155_new_n6603_), .Y(u2__abc_52155_new_n6604_));
AND2X2 AND2X2_224 ( .A(_abc_73687_new_n1270_), .B(_abc_73687_new_n1269_), .Y(fracta1_34_));
AND2X2 AND2X2_2240 ( .A(u2__abc_52155_new_n6093_), .B(u2__abc_52155_new_n6604_), .Y(u2__abc_52155_new_n6605_));
AND2X2 AND2X2_2241 ( .A(u2__abc_52155_new_n6448_), .B(u2__abc_52155_new_n6455_), .Y(u2__abc_52155_new_n6611_));
AND2X2 AND2X2_2242 ( .A(u2__abc_52155_new_n6463_), .B(u2__abc_52155_new_n6470_), .Y(u2__abc_52155_new_n6613_));
AND2X2 AND2X2_2243 ( .A(u2__abc_52155_new_n6432_), .B(u2__abc_52155_new_n6439_), .Y(u2__abc_52155_new_n6615_));
AND2X2 AND2X2_2244 ( .A(u2__abc_52155_new_n6421_), .B(u2__abc_52155_new_n6416_), .Y(u2__abc_52155_new_n6618_));
AND2X2 AND2X2_2245 ( .A(u2__abc_52155_new_n6617_), .B(u2__abc_52155_new_n6620_), .Y(u2__abc_52155_new_n6621_));
AND2X2 AND2X2_2246 ( .A(u2__abc_52155_new_n6622_), .B(u2__abc_52155_new_n6613_), .Y(u2__abc_52155_new_n6623_));
AND2X2 AND2X2_2247 ( .A(u2__abc_52155_new_n6626_), .B(u2__abc_52155_new_n6612_), .Y(u2__abc_52155_new_n6627_));
AND2X2 AND2X2_2248 ( .A(u2__abc_52155_new_n6541_), .B(u2__abc_52155_new_n6548_), .Y(u2__abc_52155_new_n6633_));
AND2X2 AND2X2_2249 ( .A(u2__abc_52155_new_n6563_), .B(u2__abc_52155_new_n6558_), .Y(u2__abc_52155_new_n6636_));
AND2X2 AND2X2_225 ( .A(_abc_73687_new_n1273_), .B(_abc_73687_new_n1272_), .Y(fracta1_35_));
AND2X2 AND2X2_2250 ( .A(u2__abc_52155_new_n6635_), .B(u2__abc_52155_new_n6638_), .Y(u2__abc_52155_new_n6639_));
AND2X2 AND2X2_2251 ( .A(u2__abc_52155_new_n6590_), .B(u2__abc_52155_new_n6597_), .Y(u2__abc_52155_new_n6642_));
AND2X2 AND2X2_2252 ( .A(u2__abc_52155_new_n6579_), .B(u2__abc_52155_new_n6574_), .Y(u2__abc_52155_new_n6645_));
AND2X2 AND2X2_2253 ( .A(u2__abc_52155_new_n6644_), .B(u2__abc_52155_new_n6647_), .Y(u2__abc_52155_new_n6648_));
AND2X2 AND2X2_2254 ( .A(u2__abc_52155_new_n6640_), .B(u2__abc_52155_new_n6648_), .Y(u2__abc_52155_new_n6649_));
AND2X2 AND2X2_2255 ( .A(u2__abc_52155_new_n6524_), .B(u2__abc_52155_new_n6531_), .Y(u2__abc_52155_new_n6653_));
AND2X2 AND2X2_2256 ( .A(u2__abc_52155_new_n6516_), .B(u2__abc_52155_new_n6511_), .Y(u2__abc_52155_new_n6656_));
AND2X2 AND2X2_2257 ( .A(u2__abc_52155_new_n6655_), .B(u2__abc_52155_new_n6658_), .Y(u2__abc_52155_new_n6659_));
AND2X2 AND2X2_2258 ( .A(u2__abc_52155_new_n6478_), .B(u2__abc_52155_new_n6485_), .Y(u2__abc_52155_new_n6661_));
AND2X2 AND2X2_2259 ( .A(u2__abc_52155_new_n6496_), .B(u2__abc_52155_new_n6503_), .Y(u2__abc_52155_new_n6664_));
AND2X2 AND2X2_226 ( .A(_abc_73687_new_n1276_), .B(_abc_73687_new_n1275_), .Y(fracta1_36_));
AND2X2 AND2X2_2260 ( .A(u2__abc_52155_new_n6666_), .B(u2__abc_52155_new_n6662_), .Y(u2__abc_52155_new_n6667_));
AND2X2 AND2X2_2261 ( .A(u2__abc_52155_new_n6660_), .B(u2__abc_52155_new_n6667_), .Y(u2__abc_52155_new_n6668_));
AND2X2 AND2X2_2262 ( .A(u2__abc_52155_new_n6650_), .B(u2__abc_52155_new_n6668_), .Y(u2__abc_52155_new_n6669_));
AND2X2 AND2X2_2263 ( .A(u2__abc_52155_new_n6369_), .B(u2__abc_52155_new_n6376_), .Y(u2__abc_52155_new_n6673_));
AND2X2 AND2X2_2264 ( .A(u2__abc_52155_new_n6358_), .B(u2__abc_52155_new_n6353_), .Y(u2__abc_52155_new_n6676_));
AND2X2 AND2X2_2265 ( .A(u2__abc_52155_new_n6675_), .B(u2__abc_52155_new_n6678_), .Y(u2__abc_52155_new_n6679_));
AND2X2 AND2X2_2266 ( .A(u2__abc_52155_new_n6400_), .B(u2__abc_52155_new_n6407_), .Y(u2__abc_52155_new_n6682_));
AND2X2 AND2X2_2267 ( .A(u2__abc_52155_new_n6385_), .B(u2__abc_52155_new_n6392_), .Y(u2__abc_52155_new_n6685_));
AND2X2 AND2X2_2268 ( .A(u2__abc_52155_new_n6684_), .B(u2__abc_52155_new_n6686_), .Y(u2__abc_52155_new_n6687_));
AND2X2 AND2X2_2269 ( .A(u2__abc_52155_new_n6680_), .B(u2__abc_52155_new_n6687_), .Y(u2__abc_52155_new_n6688_));
AND2X2 AND2X2_227 ( .A(_abc_73687_new_n1279_), .B(_abc_73687_new_n1278_), .Y(fracta1_37_));
AND2X2 AND2X2_2270 ( .A(u2__abc_52155_new_n6670_), .B(u2__abc_52155_new_n6688_), .Y(u2__abc_52155_new_n6689_));
AND2X2 AND2X2_2271 ( .A(u2__abc_52155_new_n6689_), .B(u2__abc_52155_new_n6628_), .Y(u2__abc_52155_new_n6690_));
AND2X2 AND2X2_2272 ( .A(u2__abc_52155_new_n6208_), .B(u2__abc_52155_new_n6215_), .Y(u2__abc_52155_new_n6693_));
AND2X2 AND2X2_2273 ( .A(u2__abc_52155_new_n6159_), .B(u2__abc_52155_new_n6166_), .Y(u2__abc_52155_new_n6695_));
AND2X2 AND2X2_2274 ( .A(u2__abc_52155_new_n6181_), .B(u2__abc_52155_new_n6176_), .Y(u2__abc_52155_new_n6698_));
AND2X2 AND2X2_2275 ( .A(u2__abc_52155_new_n6697_), .B(u2__abc_52155_new_n6700_), .Y(u2__abc_52155_new_n6701_));
AND2X2 AND2X2_2276 ( .A(u2__abc_52155_new_n6702_), .B(u2__abc_52155_new_n6693_), .Y(u2__abc_52155_new_n6703_));
AND2X2 AND2X2_2277 ( .A(u2__abc_52155_new_n6705_), .B(u2__abc_52155_new_n6193_), .Y(u2__abc_52155_new_n6706_));
AND2X2 AND2X2_2278 ( .A(u2__abc_52155_new_n6707_), .B(u2__abc_52155_new_n6200_), .Y(u2__abc_52155_new_n6708_));
AND2X2 AND2X2_2279 ( .A(u2__abc_52155_new_n6145_), .B(u2__abc_52155_new_n6152_), .Y(u2__abc_52155_new_n6710_));
AND2X2 AND2X2_228 ( .A(_abc_73687_new_n1282_), .B(_abc_73687_new_n1281_), .Y(fracta1_38_));
AND2X2 AND2X2_2280 ( .A(u2__abc_52155_new_n6114_), .B(u2__abc_52155_new_n6121_), .Y(u2__abc_52155_new_n6711_));
AND2X2 AND2X2_2281 ( .A(u2__abc_52155_new_n6713_), .B(u2__abc_52155_new_n6099_), .Y(u2__abc_52155_new_n6714_));
AND2X2 AND2X2_2282 ( .A(u2__abc_52155_new_n6715_), .B(u2__abc_52155_new_n6106_), .Y(u2__abc_52155_new_n6716_));
AND2X2 AND2X2_2283 ( .A(u2__abc_52155_new_n6717_), .B(u2__abc_52155_new_n6710_), .Y(u2__abc_52155_new_n6718_));
AND2X2 AND2X2_2284 ( .A(u2__abc_52155_new_n6720_), .B(u2__abc_52155_new_n6130_), .Y(u2__abc_52155_new_n6721_));
AND2X2 AND2X2_2285 ( .A(u2__abc_52155_new_n6722_), .B(u2__abc_52155_new_n6137_), .Y(u2__abc_52155_new_n6723_));
AND2X2 AND2X2_2286 ( .A(u2__abc_52155_new_n6289_), .B(u2__abc_52155_new_n6296_), .Y(u2__abc_52155_new_n6727_));
AND2X2 AND2X2_2287 ( .A(u2__abc_52155_new_n6304_), .B(u2__abc_52155_new_n6311_), .Y(u2__abc_52155_new_n6730_));
AND2X2 AND2X2_2288 ( .A(u2__abc_52155_new_n6732_), .B(u2__abc_52155_new_n6728_), .Y(u2__abc_52155_new_n6733_));
AND2X2 AND2X2_2289 ( .A(u2__abc_52155_new_n6335_), .B(u2__abc_52155_new_n6342_), .Y(u2__abc_52155_new_n6736_));
AND2X2 AND2X2_229 ( .A(_abc_73687_new_n1285_), .B(_abc_73687_new_n1284_), .Y(fracta1_39_));
AND2X2 AND2X2_2290 ( .A(u2__abc_52155_new_n6324_), .B(u2__abc_52155_new_n6319_), .Y(u2__abc_52155_new_n6739_));
AND2X2 AND2X2_2291 ( .A(u2__abc_52155_new_n6738_), .B(u2__abc_52155_new_n6741_), .Y(u2__abc_52155_new_n6742_));
AND2X2 AND2X2_2292 ( .A(u2__abc_52155_new_n6734_), .B(u2__abc_52155_new_n6742_), .Y(u2__abc_52155_new_n6743_));
AND2X2 AND2X2_2293 ( .A(u2__abc_52155_new_n6223_), .B(u2__abc_52155_new_n6230_), .Y(u2__abc_52155_new_n6747_));
AND2X2 AND2X2_2294 ( .A(u2__abc_52155_new_n6245_), .B(u2__abc_52155_new_n6240_), .Y(u2__abc_52155_new_n6750_));
AND2X2 AND2X2_2295 ( .A(u2__abc_52155_new_n6749_), .B(u2__abc_52155_new_n6752_), .Y(u2__abc_52155_new_n6753_));
AND2X2 AND2X2_2296 ( .A(u2__abc_52155_new_n6272_), .B(u2__abc_52155_new_n6279_), .Y(u2__abc_52155_new_n6756_));
AND2X2 AND2X2_2297 ( .A(u2__abc_52155_new_n6261_), .B(u2__abc_52155_new_n6256_), .Y(u2__abc_52155_new_n6759_));
AND2X2 AND2X2_2298 ( .A(u2__abc_52155_new_n6758_), .B(u2__abc_52155_new_n6761_), .Y(u2__abc_52155_new_n6762_));
AND2X2 AND2X2_2299 ( .A(u2__abc_52155_new_n6754_), .B(u2__abc_52155_new_n6762_), .Y(u2__abc_52155_new_n6763_));
AND2X2 AND2X2_23 ( .A(_abc_73687_new_n753_), .B(sqrto_22_), .Y(\o[58] ));
AND2X2 AND2X2_230 ( .A(_abc_73687_new_n1288_), .B(_abc_73687_new_n1287_), .Y(fracta1_40_));
AND2X2 AND2X2_2300 ( .A(u2__abc_52155_new_n6744_), .B(u2__abc_52155_new_n6763_), .Y(u2__abc_52155_new_n6764_));
AND2X2 AND2X2_2301 ( .A(u2__abc_52155_new_n6723_), .B(u2__abc_52155_new_n6765_), .Y(u2__abc_52155_new_n6766_));
AND2X2 AND2X2_2302 ( .A(u2__abc_52155_new_n6766_), .B(u2__abc_52155_new_n6709_), .Y(u2__abc_52155_new_n6767_));
AND2X2 AND2X2_2303 ( .A(u2__abc_52155_new_n6767_), .B(u2__abc_52155_new_n6691_), .Y(u2__abc_52155_new_n6768_));
AND2X2 AND2X2_2304 ( .A(u2__abc_52155_new_n6061_), .B(u2__abc_52155_new_n6068_), .Y(u2__abc_52155_new_n6775_));
AND2X2 AND2X2_2305 ( .A(u2__abc_52155_new_n6778_), .B(u2__abc_52155_new_n6086_), .Y(u2__abc_52155_new_n6779_));
AND2X2 AND2X2_2306 ( .A(u2__abc_52155_new_n6777_), .B(u2__abc_52155_new_n6779_), .Y(u2__abc_52155_new_n6780_));
AND2X2 AND2X2_2307 ( .A(u2__abc_52155_new_n6030_), .B(u2__abc_52155_new_n6037_), .Y(u2__abc_52155_new_n6782_));
AND2X2 AND2X2_2308 ( .A(u2__abc_52155_new_n6048_), .B(u2__abc_52155_new_n6055_), .Y(u2__abc_52155_new_n6785_));
AND2X2 AND2X2_2309 ( .A(u2__abc_52155_new_n6787_), .B(u2__abc_52155_new_n6783_), .Y(u2__abc_52155_new_n6788_));
AND2X2 AND2X2_231 ( .A(_abc_73687_new_n1291_), .B(_abc_73687_new_n1290_), .Y(fracta1_41_));
AND2X2 AND2X2_2310 ( .A(u2__abc_52155_new_n6781_), .B(u2__abc_52155_new_n6788_), .Y(u2__abc_52155_new_n6789_));
AND2X2 AND2X2_2311 ( .A(u2__abc_52155_new_n5967_), .B(u2__abc_52155_new_n5974_), .Y(u2__abc_52155_new_n6793_));
AND2X2 AND2X2_2312 ( .A(u2__abc_52155_new_n5989_), .B(u2__abc_52155_new_n5984_), .Y(u2__abc_52155_new_n6796_));
AND2X2 AND2X2_2313 ( .A(u2__abc_52155_new_n6795_), .B(u2__abc_52155_new_n6798_), .Y(u2__abc_52155_new_n6799_));
AND2X2 AND2X2_2314 ( .A(u2__abc_52155_new_n6016_), .B(u2__abc_52155_new_n6023_), .Y(u2__abc_52155_new_n6802_));
AND2X2 AND2X2_2315 ( .A(u2__abc_52155_new_n6001_), .B(u2__abc_52155_new_n6008_), .Y(u2__abc_52155_new_n6805_));
AND2X2 AND2X2_2316 ( .A(u2__abc_52155_new_n6804_), .B(u2__abc_52155_new_n6806_), .Y(u2__abc_52155_new_n6807_));
AND2X2 AND2X2_2317 ( .A(u2__abc_52155_new_n6800_), .B(u2__abc_52155_new_n6807_), .Y(u2__abc_52155_new_n6808_));
AND2X2 AND2X2_2318 ( .A(u2__abc_52155_new_n6790_), .B(u2__abc_52155_new_n6808_), .Y(u2__abc_52155_new_n6809_));
AND2X2 AND2X2_2319 ( .A(u2__abc_52155_new_n5858_), .B(u2__abc_52155_new_n5865_), .Y(u2__abc_52155_new_n6813_));
AND2X2 AND2X2_232 ( .A(_abc_73687_new_n1294_), .B(_abc_73687_new_n1293_), .Y(fracta1_42_));
AND2X2 AND2X2_2320 ( .A(u2__abc_52155_new_n5847_), .B(u2__abc_52155_new_n5842_), .Y(u2__abc_52155_new_n6816_));
AND2X2 AND2X2_2321 ( .A(u2__abc_52155_new_n6815_), .B(u2__abc_52155_new_n6818_), .Y(u2__abc_52155_new_n6819_));
AND2X2 AND2X2_2322 ( .A(u2__abc_52155_new_n5889_), .B(u2__abc_52155_new_n5896_), .Y(u2__abc_52155_new_n6822_));
AND2X2 AND2X2_2323 ( .A(u2__abc_52155_new_n5878_), .B(u2__abc_52155_new_n5873_), .Y(u2__abc_52155_new_n6825_));
AND2X2 AND2X2_2324 ( .A(u2__abc_52155_new_n6824_), .B(u2__abc_52155_new_n6827_), .Y(u2__abc_52155_new_n6828_));
AND2X2 AND2X2_2325 ( .A(u2__abc_52155_new_n6820_), .B(u2__abc_52155_new_n6828_), .Y(u2__abc_52155_new_n6829_));
AND2X2 AND2X2_2326 ( .A(u2__abc_52155_new_n5941_), .B(u2__abc_52155_new_n5936_), .Y(u2__abc_52155_new_n6831_));
AND2X2 AND2X2_2327 ( .A(u2__abc_52155_new_n5952_), .B(u2__abc_52155_new_n5959_), .Y(u2__abc_52155_new_n6834_));
AND2X2 AND2X2_2328 ( .A(u2__abc_52155_new_n5906_), .B(u2__abc_52155_new_n5913_), .Y(u2__abc_52155_new_n6835_));
AND2X2 AND2X2_2329 ( .A(u2__abc_52155_new_n5921_), .B(u2__abc_52155_new_n5928_), .Y(u2__abc_52155_new_n6838_));
AND2X2 AND2X2_233 ( .A(_abc_73687_new_n1297_), .B(_abc_73687_new_n1296_), .Y(fracta1_43_));
AND2X2 AND2X2_2330 ( .A(u2__abc_52155_new_n6840_), .B(u2__abc_52155_new_n6836_), .Y(u2__abc_52155_new_n6841_));
AND2X2 AND2X2_2331 ( .A(u2__abc_52155_new_n6842_), .B(u2__abc_52155_new_n6834_), .Y(u2__abc_52155_new_n6843_));
AND2X2 AND2X2_2332 ( .A(u2__abc_52155_new_n6846_), .B(u2__abc_52155_new_n6833_), .Y(u2__abc_52155_new_n6847_));
AND2X2 AND2X2_2333 ( .A(u2__abc_52155_new_n6848_), .B(u2__abc_52155_new_n6829_), .Y(u2__abc_52155_new_n6849_));
AND2X2 AND2X2_2334 ( .A(u2__abc_52155_new_n6849_), .B(u2__abc_52155_new_n6810_), .Y(u2__abc_52155_new_n6850_));
AND2X2 AND2X2_2335 ( .A(u2__abc_52155_new_n5697_), .B(u2__abc_52155_new_n5704_), .Y(u2__abc_52155_new_n6853_));
AND2X2 AND2X2_2336 ( .A(u2__abc_52155_new_n5651_), .B(u2__abc_52155_new_n5658_), .Y(u2__abc_52155_new_n6856_));
AND2X2 AND2X2_2337 ( .A(u2__abc_52155_new_n5666_), .B(u2__abc_52155_new_n5673_), .Y(u2__abc_52155_new_n6859_));
AND2X2 AND2X2_2338 ( .A(u2__abc_52155_new_n6861_), .B(u2__abc_52155_new_n6857_), .Y(u2__abc_52155_new_n6862_));
AND2X2 AND2X2_2339 ( .A(u2__abc_52155_new_n6863_), .B(u2__abc_52155_new_n6854_), .Y(u2__abc_52155_new_n6864_));
AND2X2 AND2X2_234 ( .A(_abc_73687_new_n1300_), .B(_abc_73687_new_n1299_), .Y(fracta1_44_));
AND2X2 AND2X2_2340 ( .A(u2__abc_52155_new_n6865_), .B(u2__abc_52155_new_n5682_), .Y(u2__abc_52155_new_n6866_));
AND2X2 AND2X2_2341 ( .A(u2__abc_52155_new_n6867_), .B(u2__abc_52155_new_n5689_), .Y(u2__abc_52155_new_n6868_));
AND2X2 AND2X2_2342 ( .A(u2__abc_52155_new_n5761_), .B(u2__abc_52155_new_n5768_), .Y(u2__abc_52155_new_n6871_));
AND2X2 AND2X2_2343 ( .A(u2__abc_52155_new_n5730_), .B(u2__abc_52155_new_n5737_), .Y(u2__abc_52155_new_n6872_));
AND2X2 AND2X2_2344 ( .A(u2__abc_52155_new_n5712_), .B(u2__abc_52155_new_n5719_), .Y(u2__abc_52155_new_n6873_));
AND2X2 AND2X2_2345 ( .A(u2__abc_52155_new_n6875_), .B(u2__abc_52155_new_n6872_), .Y(u2__abc_52155_new_n6876_));
AND2X2 AND2X2_2346 ( .A(u2__abc_52155_new_n6878_), .B(u2__abc_52155_new_n6871_), .Y(u2__abc_52155_new_n6879_));
AND2X2 AND2X2_2347 ( .A(u2__abc_52155_new_n6881_), .B(u2__abc_52155_new_n5746_), .Y(u2__abc_52155_new_n6882_));
AND2X2 AND2X2_2348 ( .A(u2__abc_52155_new_n6883_), .B(u2__abc_52155_new_n5753_), .Y(u2__abc_52155_new_n6884_));
AND2X2 AND2X2_2349 ( .A(u2__abc_52155_new_n5809_), .B(u2__abc_52155_new_n5816_), .Y(u2__abc_52155_new_n6885_));
AND2X2 AND2X2_235 ( .A(_abc_73687_new_n1303_), .B(_abc_73687_new_n1302_), .Y(fracta1_45_));
AND2X2 AND2X2_2350 ( .A(u2__abc_52155_new_n5824_), .B(u2__abc_52155_new_n5831_), .Y(u2__abc_52155_new_n6886_));
AND2X2 AND2X2_2351 ( .A(u2__abc_52155_new_n5778_), .B(u2__abc_52155_new_n5785_), .Y(u2__abc_52155_new_n6887_));
AND2X2 AND2X2_2352 ( .A(u2__abc_52155_new_n5793_), .B(u2__abc_52155_new_n5800_), .Y(u2__abc_52155_new_n6890_));
AND2X2 AND2X2_2353 ( .A(u2__abc_52155_new_n6892_), .B(u2__abc_52155_new_n6888_), .Y(u2__abc_52155_new_n6893_));
AND2X2 AND2X2_2354 ( .A(u2__abc_52155_new_n6894_), .B(u2__abc_52155_new_n6886_), .Y(u2__abc_52155_new_n6895_));
AND2X2 AND2X2_2355 ( .A(u2__abc_52155_new_n6897_), .B(u2__abc_52155_new_n6885_), .Y(u2__abc_52155_new_n6898_));
AND2X2 AND2X2_2356 ( .A(u2__abc_52155_new_n5772_), .B(u2__abc_52155_new_n5813_), .Y(u2__abc_52155_new_n6899_));
AND2X2 AND2X2_2357 ( .A(u2__abc_52155_new_n6901_), .B(u2__abc_52155_new_n6884_), .Y(u2__abc_52155_new_n6902_));
AND2X2 AND2X2_2358 ( .A(u2__abc_52155_new_n5634_), .B(u2__abc_52155_new_n5641_), .Y(u2__abc_52155_new_n6905_));
AND2X2 AND2X2_2359 ( .A(u2__abc_52155_new_n5616_), .B(u2__abc_52155_new_n5623_), .Y(u2__abc_52155_new_n6908_));
AND2X2 AND2X2_236 ( .A(_abc_73687_new_n1306_), .B(_abc_73687_new_n1305_), .Y(fracta1_46_));
AND2X2 AND2X2_2360 ( .A(u2__abc_52155_new_n6910_), .B(u2__abc_52155_new_n6906_), .Y(u2__abc_52155_new_n6911_));
AND2X2 AND2X2_2361 ( .A(u2__abc_52155_new_n5603_), .B(u2__abc_52155_new_n5610_), .Y(u2__abc_52155_new_n6914_));
AND2X2 AND2X2_2362 ( .A(u2__abc_52155_new_n5595_), .B(u2__abc_52155_new_n5587_), .Y(u2__abc_52155_new_n6917_));
AND2X2 AND2X2_2363 ( .A(u2__abc_52155_new_n6916_), .B(u2__abc_52155_new_n6919_), .Y(u2__abc_52155_new_n6920_));
AND2X2 AND2X2_2364 ( .A(u2__abc_52155_new_n6912_), .B(u2__abc_52155_new_n6920_), .Y(u2__abc_52155_new_n6921_));
AND2X2 AND2X2_2365 ( .A(u2__abc_52155_new_n6903_), .B(u2__abc_52155_new_n6921_), .Y(u2__abc_52155_new_n6922_));
AND2X2 AND2X2_2366 ( .A(u2__abc_52155_new_n6922_), .B(u2__abc_52155_new_n6869_), .Y(u2__abc_52155_new_n6923_));
AND2X2 AND2X2_2367 ( .A(u2__abc_52155_new_n6923_), .B(u2__abc_52155_new_n6851_), .Y(u2__abc_52155_new_n6924_));
AND2X2 AND2X2_2368 ( .A(u2__abc_52155_new_n6769_), .B(u2__abc_52155_new_n6924_), .Y(u2__abc_52155_new_n6925_));
AND2X2 AND2X2_2369 ( .A(u2__abc_52155_new_n6607_), .B(u2__abc_52155_new_n6925_), .Y(u2__abc_52155_new_n6926_));
AND2X2 AND2X2_237 ( .A(_abc_73687_new_n1309_), .B(_abc_73687_new_n1308_), .Y(fracta1_47_));
AND2X2 AND2X2_2370 ( .A(u2__abc_52155_new_n6927_), .B(u2_remHi_444_), .Y(u2__abc_52155_new_n6928_));
AND2X2 AND2X2_2371 ( .A(u2__abc_52155_new_n6930_), .B(u2_o_444_), .Y(u2__abc_52155_new_n6931_));
AND2X2 AND2X2_2372 ( .A(u2__abc_52155_new_n6929_), .B(u2__abc_52155_new_n6932_), .Y(u2__abc_52155_new_n6933_));
AND2X2 AND2X2_2373 ( .A(u2__abc_52155_new_n6934_), .B(u2_o_445_), .Y(u2__abc_52155_new_n6935_));
AND2X2 AND2X2_2374 ( .A(u2__abc_52155_new_n6937_), .B(u2_remHi_445_), .Y(u2__abc_52155_new_n6938_));
AND2X2 AND2X2_2375 ( .A(u2__abc_52155_new_n6936_), .B(u2__abc_52155_new_n6939_), .Y(u2__abc_52155_new_n6940_));
AND2X2 AND2X2_2376 ( .A(u2__abc_52155_new_n6933_), .B(u2__abc_52155_new_n6940_), .Y(u2__abc_52155_new_n6941_));
AND2X2 AND2X2_2377 ( .A(u2__abc_52155_new_n6942_), .B(u2_o_443_), .Y(u2__abc_52155_new_n6943_));
AND2X2 AND2X2_2378 ( .A(u2__abc_52155_new_n6945_), .B(u2_remHi_443_), .Y(u2__abc_52155_new_n6946_));
AND2X2 AND2X2_2379 ( .A(u2__abc_52155_new_n6944_), .B(u2__abc_52155_new_n6947_), .Y(u2__abc_52155_new_n6948_));
AND2X2 AND2X2_238 ( .A(_abc_73687_new_n1312_), .B(_abc_73687_new_n1311_), .Y(fracta1_48_));
AND2X2 AND2X2_2380 ( .A(u2__abc_52155_new_n6949_), .B(u2_remHi_442_), .Y(u2__abc_52155_new_n6950_));
AND2X2 AND2X2_2381 ( .A(u2__abc_52155_new_n6952_), .B(u2_o_442_), .Y(u2__abc_52155_new_n6953_));
AND2X2 AND2X2_2382 ( .A(u2__abc_52155_new_n6951_), .B(u2__abc_52155_new_n6954_), .Y(u2__abc_52155_new_n6955_));
AND2X2 AND2X2_2383 ( .A(u2__abc_52155_new_n6948_), .B(u2__abc_52155_new_n6955_), .Y(u2__abc_52155_new_n6956_));
AND2X2 AND2X2_2384 ( .A(u2__abc_52155_new_n6941_), .B(u2__abc_52155_new_n6956_), .Y(u2__abc_52155_new_n6957_));
AND2X2 AND2X2_2385 ( .A(u2__abc_52155_new_n6958_), .B(u2_remHi_438_), .Y(u2__abc_52155_new_n6959_));
AND2X2 AND2X2_2386 ( .A(u2__abc_52155_new_n6961_), .B(u2_o_438_), .Y(u2__abc_52155_new_n6962_));
AND2X2 AND2X2_2387 ( .A(u2__abc_52155_new_n6960_), .B(u2__abc_52155_new_n6963_), .Y(u2__abc_52155_new_n6964_));
AND2X2 AND2X2_2388 ( .A(u2__abc_52155_new_n6965_), .B(u2_o_439_), .Y(u2__abc_52155_new_n6966_));
AND2X2 AND2X2_2389 ( .A(u2__abc_52155_new_n6968_), .B(u2_remHi_439_), .Y(u2__abc_52155_new_n6969_));
AND2X2 AND2X2_239 ( .A(_abc_73687_new_n1315_), .B(_abc_73687_new_n1314_), .Y(fracta1_49_));
AND2X2 AND2X2_2390 ( .A(u2__abc_52155_new_n6967_), .B(u2__abc_52155_new_n6970_), .Y(u2__abc_52155_new_n6971_));
AND2X2 AND2X2_2391 ( .A(u2__abc_52155_new_n6964_), .B(u2__abc_52155_new_n6971_), .Y(u2__abc_52155_new_n6972_));
AND2X2 AND2X2_2392 ( .A(u2__abc_52155_new_n6973_), .B(u2_remHi_440_), .Y(u2__abc_52155_new_n6974_));
AND2X2 AND2X2_2393 ( .A(u2__abc_52155_new_n6976_), .B(u2_o_440_), .Y(u2__abc_52155_new_n6977_));
AND2X2 AND2X2_2394 ( .A(u2__abc_52155_new_n6975_), .B(u2__abc_52155_new_n6978_), .Y(u2__abc_52155_new_n6979_));
AND2X2 AND2X2_2395 ( .A(u2__abc_52155_new_n6980_), .B(u2_o_441_), .Y(u2__abc_52155_new_n6981_));
AND2X2 AND2X2_2396 ( .A(u2__abc_52155_new_n6983_), .B(u2_remHi_441_), .Y(u2__abc_52155_new_n6984_));
AND2X2 AND2X2_2397 ( .A(u2__abc_52155_new_n6982_), .B(u2__abc_52155_new_n6985_), .Y(u2__abc_52155_new_n6986_));
AND2X2 AND2X2_2398 ( .A(u2__abc_52155_new_n6979_), .B(u2__abc_52155_new_n6986_), .Y(u2__abc_52155_new_n6987_));
AND2X2 AND2X2_2399 ( .A(u2__abc_52155_new_n6972_), .B(u2__abc_52155_new_n6987_), .Y(u2__abc_52155_new_n6988_));
AND2X2 AND2X2_24 ( .A(_abc_73687_new_n753_), .B(sqrto_23_), .Y(\o[59] ));
AND2X2 AND2X2_240 ( .A(_abc_73687_new_n1318_), .B(_abc_73687_new_n1317_), .Y(fracta1_50_));
AND2X2 AND2X2_2400 ( .A(u2__abc_52155_new_n6957_), .B(u2__abc_52155_new_n6988_), .Y(u2__abc_52155_new_n6989_));
AND2X2 AND2X2_2401 ( .A(u2__abc_52155_new_n6990_), .B(u2_remHi_436_), .Y(u2__abc_52155_new_n6991_));
AND2X2 AND2X2_2402 ( .A(u2__abc_52155_new_n6993_), .B(u2_o_436_), .Y(u2__abc_52155_new_n6994_));
AND2X2 AND2X2_2403 ( .A(u2__abc_52155_new_n6992_), .B(u2__abc_52155_new_n6995_), .Y(u2__abc_52155_new_n6996_));
AND2X2 AND2X2_2404 ( .A(u2__abc_52155_new_n6997_), .B(u2_remHi_437_), .Y(u2__abc_52155_new_n6998_));
AND2X2 AND2X2_2405 ( .A(u2__abc_52155_new_n7000_), .B(u2_o_437_), .Y(u2__abc_52155_new_n7001_));
AND2X2 AND2X2_2406 ( .A(u2__abc_52155_new_n6999_), .B(u2__abc_52155_new_n7002_), .Y(u2__abc_52155_new_n7003_));
AND2X2 AND2X2_2407 ( .A(u2__abc_52155_new_n6996_), .B(u2__abc_52155_new_n7003_), .Y(u2__abc_52155_new_n7004_));
AND2X2 AND2X2_2408 ( .A(u2__abc_52155_new_n7005_), .B(u2_o_435_), .Y(u2__abc_52155_new_n7006_));
AND2X2 AND2X2_2409 ( .A(u2__abc_52155_new_n7008_), .B(u2_remHi_435_), .Y(u2__abc_52155_new_n7009_));
AND2X2 AND2X2_241 ( .A(_abc_73687_new_n1321_), .B(_abc_73687_new_n1320_), .Y(fracta1_51_));
AND2X2 AND2X2_2410 ( .A(u2__abc_52155_new_n7007_), .B(u2__abc_52155_new_n7010_), .Y(u2__abc_52155_new_n7011_));
AND2X2 AND2X2_2411 ( .A(u2__abc_52155_new_n7012_), .B(u2_remHi_434_), .Y(u2__abc_52155_new_n7013_));
AND2X2 AND2X2_2412 ( .A(u2__abc_52155_new_n7015_), .B(u2_o_434_), .Y(u2__abc_52155_new_n7016_));
AND2X2 AND2X2_2413 ( .A(u2__abc_52155_new_n7014_), .B(u2__abc_52155_new_n7017_), .Y(u2__abc_52155_new_n7018_));
AND2X2 AND2X2_2414 ( .A(u2__abc_52155_new_n7011_), .B(u2__abc_52155_new_n7018_), .Y(u2__abc_52155_new_n7019_));
AND2X2 AND2X2_2415 ( .A(u2__abc_52155_new_n7004_), .B(u2__abc_52155_new_n7019_), .Y(u2__abc_52155_new_n7020_));
AND2X2 AND2X2_2416 ( .A(u2__abc_52155_new_n7021_), .B(u2_remHi_430_), .Y(u2__abc_52155_new_n7022_));
AND2X2 AND2X2_2417 ( .A(u2__abc_52155_new_n7024_), .B(u2_o_430_), .Y(u2__abc_52155_new_n7025_));
AND2X2 AND2X2_2418 ( .A(u2__abc_52155_new_n7023_), .B(u2__abc_52155_new_n7026_), .Y(u2__abc_52155_new_n7027_));
AND2X2 AND2X2_2419 ( .A(u2__abc_52155_new_n7028_), .B(u2_o_431_), .Y(u2__abc_52155_new_n7029_));
AND2X2 AND2X2_242 ( .A(_abc_73687_new_n1324_), .B(_abc_73687_new_n1323_), .Y(fracta1_52_));
AND2X2 AND2X2_2420 ( .A(u2__abc_52155_new_n7031_), .B(u2_remHi_431_), .Y(u2__abc_52155_new_n7032_));
AND2X2 AND2X2_2421 ( .A(u2__abc_52155_new_n7030_), .B(u2__abc_52155_new_n7033_), .Y(u2__abc_52155_new_n7034_));
AND2X2 AND2X2_2422 ( .A(u2__abc_52155_new_n7027_), .B(u2__abc_52155_new_n7034_), .Y(u2__abc_52155_new_n7035_));
AND2X2 AND2X2_2423 ( .A(u2__abc_52155_new_n7036_), .B(u2_remHi_432_), .Y(u2__abc_52155_new_n7037_));
AND2X2 AND2X2_2424 ( .A(u2__abc_52155_new_n7039_), .B(u2_o_432_), .Y(u2__abc_52155_new_n7040_));
AND2X2 AND2X2_2425 ( .A(u2__abc_52155_new_n7038_), .B(u2__abc_52155_new_n7041_), .Y(u2__abc_52155_new_n7042_));
AND2X2 AND2X2_2426 ( .A(u2__abc_52155_new_n7043_), .B(u2_o_433_), .Y(u2__abc_52155_new_n7044_));
AND2X2 AND2X2_2427 ( .A(u2__abc_52155_new_n7046_), .B(u2_remHi_433_), .Y(u2__abc_52155_new_n7047_));
AND2X2 AND2X2_2428 ( .A(u2__abc_52155_new_n7045_), .B(u2__abc_52155_new_n7048_), .Y(u2__abc_52155_new_n7049_));
AND2X2 AND2X2_2429 ( .A(u2__abc_52155_new_n7042_), .B(u2__abc_52155_new_n7049_), .Y(u2__abc_52155_new_n7050_));
AND2X2 AND2X2_243 ( .A(_abc_73687_new_n1327_), .B(_abc_73687_new_n1326_), .Y(fracta1_53_));
AND2X2 AND2X2_2430 ( .A(u2__abc_52155_new_n7035_), .B(u2__abc_52155_new_n7050_), .Y(u2__abc_52155_new_n7051_));
AND2X2 AND2X2_2431 ( .A(u2__abc_52155_new_n7020_), .B(u2__abc_52155_new_n7051_), .Y(u2__abc_52155_new_n7052_));
AND2X2 AND2X2_2432 ( .A(u2__abc_52155_new_n6989_), .B(u2__abc_52155_new_n7052_), .Y(u2__abc_52155_new_n7053_));
AND2X2 AND2X2_2433 ( .A(u2__abc_52155_new_n7054_), .B(u2_remHi_424_), .Y(u2__abc_52155_new_n7055_));
AND2X2 AND2X2_2434 ( .A(u2__abc_52155_new_n7057_), .B(u2_o_424_), .Y(u2__abc_52155_new_n7058_));
AND2X2 AND2X2_2435 ( .A(u2__abc_52155_new_n7056_), .B(u2__abc_52155_new_n7059_), .Y(u2__abc_52155_new_n7060_));
AND2X2 AND2X2_2436 ( .A(u2__abc_52155_new_n7061_), .B(u2_o_425_), .Y(u2__abc_52155_new_n7062_));
AND2X2 AND2X2_2437 ( .A(u2__abc_52155_new_n7064_), .B(u2_remHi_425_), .Y(u2__abc_52155_new_n7065_));
AND2X2 AND2X2_2438 ( .A(u2__abc_52155_new_n7063_), .B(u2__abc_52155_new_n7066_), .Y(u2__abc_52155_new_n7067_));
AND2X2 AND2X2_2439 ( .A(u2__abc_52155_new_n7060_), .B(u2__abc_52155_new_n7067_), .Y(u2__abc_52155_new_n7068_));
AND2X2 AND2X2_244 ( .A(_abc_73687_new_n1330_), .B(_abc_73687_new_n1329_), .Y(fracta1_54_));
AND2X2 AND2X2_2440 ( .A(u2__abc_52155_new_n7069_), .B(u2_remHi_422_), .Y(u2__abc_52155_new_n7070_));
AND2X2 AND2X2_2441 ( .A(u2__abc_52155_new_n7072_), .B(u2_o_422_), .Y(u2__abc_52155_new_n7073_));
AND2X2 AND2X2_2442 ( .A(u2__abc_52155_new_n7071_), .B(u2__abc_52155_new_n7074_), .Y(u2__abc_52155_new_n7075_));
AND2X2 AND2X2_2443 ( .A(u2__abc_52155_new_n7076_), .B(u2_o_423_), .Y(u2__abc_52155_new_n7077_));
AND2X2 AND2X2_2444 ( .A(u2__abc_52155_new_n7079_), .B(u2_remHi_423_), .Y(u2__abc_52155_new_n7080_));
AND2X2 AND2X2_2445 ( .A(u2__abc_52155_new_n7078_), .B(u2__abc_52155_new_n7081_), .Y(u2__abc_52155_new_n7082_));
AND2X2 AND2X2_2446 ( .A(u2__abc_52155_new_n7075_), .B(u2__abc_52155_new_n7082_), .Y(u2__abc_52155_new_n7083_));
AND2X2 AND2X2_2447 ( .A(u2__abc_52155_new_n7068_), .B(u2__abc_52155_new_n7083_), .Y(u2__abc_52155_new_n7084_));
AND2X2 AND2X2_2448 ( .A(u2__abc_52155_new_n7085_), .B(u2_remHi_428_), .Y(u2__abc_52155_new_n7086_));
AND2X2 AND2X2_2449 ( .A(u2__abc_52155_new_n7088_), .B(u2_o_428_), .Y(u2__abc_52155_new_n7089_));
AND2X2 AND2X2_245 ( .A(_abc_73687_new_n1333_), .B(_abc_73687_new_n1332_), .Y(fracta1_55_));
AND2X2 AND2X2_2450 ( .A(u2__abc_52155_new_n7087_), .B(u2__abc_52155_new_n7090_), .Y(u2__abc_52155_new_n7091_));
AND2X2 AND2X2_2451 ( .A(u2__abc_52155_new_n7092_), .B(u2_remHi_429_), .Y(u2__abc_52155_new_n7093_));
AND2X2 AND2X2_2452 ( .A(u2__abc_52155_new_n7095_), .B(u2_o_429_), .Y(u2__abc_52155_new_n7096_));
AND2X2 AND2X2_2453 ( .A(u2__abc_52155_new_n7094_), .B(u2__abc_52155_new_n7097_), .Y(u2__abc_52155_new_n7098_));
AND2X2 AND2X2_2454 ( .A(u2__abc_52155_new_n7091_), .B(u2__abc_52155_new_n7098_), .Y(u2__abc_52155_new_n7099_));
AND2X2 AND2X2_2455 ( .A(u2__abc_52155_new_n7100_), .B(u2_o_427_), .Y(u2__abc_52155_new_n7101_));
AND2X2 AND2X2_2456 ( .A(u2__abc_52155_new_n7103_), .B(u2_remHi_427_), .Y(u2__abc_52155_new_n7104_));
AND2X2 AND2X2_2457 ( .A(u2__abc_52155_new_n7102_), .B(u2__abc_52155_new_n7105_), .Y(u2__abc_52155_new_n7106_));
AND2X2 AND2X2_2458 ( .A(u2__abc_52155_new_n7107_), .B(u2_remHi_426_), .Y(u2__abc_52155_new_n7108_));
AND2X2 AND2X2_2459 ( .A(u2__abc_52155_new_n7110_), .B(u2_o_426_), .Y(u2__abc_52155_new_n7111_));
AND2X2 AND2X2_246 ( .A(_abc_73687_new_n1336_), .B(_abc_73687_new_n1335_), .Y(fracta1_56_));
AND2X2 AND2X2_2460 ( .A(u2__abc_52155_new_n7109_), .B(u2__abc_52155_new_n7112_), .Y(u2__abc_52155_new_n7113_));
AND2X2 AND2X2_2461 ( .A(u2__abc_52155_new_n7106_), .B(u2__abc_52155_new_n7113_), .Y(u2__abc_52155_new_n7114_));
AND2X2 AND2X2_2462 ( .A(u2__abc_52155_new_n7099_), .B(u2__abc_52155_new_n7114_), .Y(u2__abc_52155_new_n7115_));
AND2X2 AND2X2_2463 ( .A(u2__abc_52155_new_n7084_), .B(u2__abc_52155_new_n7115_), .Y(u2__abc_52155_new_n7116_));
AND2X2 AND2X2_2464 ( .A(u2__abc_52155_new_n7117_), .B(u2_remHi_420_), .Y(u2__abc_52155_new_n7118_));
AND2X2 AND2X2_2465 ( .A(u2__abc_52155_new_n7120_), .B(u2_o_420_), .Y(u2__abc_52155_new_n7121_));
AND2X2 AND2X2_2466 ( .A(u2__abc_52155_new_n7119_), .B(u2__abc_52155_new_n7122_), .Y(u2__abc_52155_new_n7123_));
AND2X2 AND2X2_2467 ( .A(u2__abc_52155_new_n7124_), .B(u2_remHi_421_), .Y(u2__abc_52155_new_n7125_));
AND2X2 AND2X2_2468 ( .A(u2__abc_52155_new_n7127_), .B(u2_o_421_), .Y(u2__abc_52155_new_n7128_));
AND2X2 AND2X2_2469 ( .A(u2__abc_52155_new_n7126_), .B(u2__abc_52155_new_n7129_), .Y(u2__abc_52155_new_n7130_));
AND2X2 AND2X2_247 ( .A(_abc_73687_new_n1339_), .B(_abc_73687_new_n1338_), .Y(fracta1_57_));
AND2X2 AND2X2_2470 ( .A(u2__abc_52155_new_n7123_), .B(u2__abc_52155_new_n7130_), .Y(u2__abc_52155_new_n7131_));
AND2X2 AND2X2_2471 ( .A(u2__abc_52155_new_n7132_), .B(u2_o_419_), .Y(u2__abc_52155_new_n7133_));
AND2X2 AND2X2_2472 ( .A(u2__abc_52155_new_n7135_), .B(u2_remHi_419_), .Y(u2__abc_52155_new_n7136_));
AND2X2 AND2X2_2473 ( .A(u2__abc_52155_new_n7134_), .B(u2__abc_52155_new_n7137_), .Y(u2__abc_52155_new_n7138_));
AND2X2 AND2X2_2474 ( .A(u2__abc_52155_new_n7139_), .B(u2_remHi_418_), .Y(u2__abc_52155_new_n7140_));
AND2X2 AND2X2_2475 ( .A(u2__abc_52155_new_n7142_), .B(u2_o_418_), .Y(u2__abc_52155_new_n7143_));
AND2X2 AND2X2_2476 ( .A(u2__abc_52155_new_n7141_), .B(u2__abc_52155_new_n7144_), .Y(u2__abc_52155_new_n7145_));
AND2X2 AND2X2_2477 ( .A(u2__abc_52155_new_n7138_), .B(u2__abc_52155_new_n7145_), .Y(u2__abc_52155_new_n7146_));
AND2X2 AND2X2_2478 ( .A(u2__abc_52155_new_n7131_), .B(u2__abc_52155_new_n7146_), .Y(u2__abc_52155_new_n7147_));
AND2X2 AND2X2_2479 ( .A(u2__abc_52155_new_n7148_), .B(u2_remHi_416_), .Y(u2__abc_52155_new_n7149_));
AND2X2 AND2X2_248 ( .A(_abc_73687_new_n1342_), .B(_abc_73687_new_n1341_), .Y(fracta1_58_));
AND2X2 AND2X2_2480 ( .A(u2__abc_52155_new_n7151_), .B(u2_o_416_), .Y(u2__abc_52155_new_n7152_));
AND2X2 AND2X2_2481 ( .A(u2__abc_52155_new_n7150_), .B(u2__abc_52155_new_n7153_), .Y(u2__abc_52155_new_n7154_));
AND2X2 AND2X2_2482 ( .A(u2__abc_52155_new_n7155_), .B(u2_o_417_), .Y(u2__abc_52155_new_n7156_));
AND2X2 AND2X2_2483 ( .A(u2__abc_52155_new_n7158_), .B(u2_remHi_417_), .Y(u2__abc_52155_new_n7159_));
AND2X2 AND2X2_2484 ( .A(u2__abc_52155_new_n7157_), .B(u2__abc_52155_new_n7160_), .Y(u2__abc_52155_new_n7161_));
AND2X2 AND2X2_2485 ( .A(u2__abc_52155_new_n7154_), .B(u2__abc_52155_new_n7161_), .Y(u2__abc_52155_new_n7162_));
AND2X2 AND2X2_2486 ( .A(u2__abc_52155_new_n7163_), .B(u2_o_415_), .Y(u2__abc_52155_new_n7164_));
AND2X2 AND2X2_2487 ( .A(u2__abc_52155_new_n7166_), .B(u2_remHi_415_), .Y(u2__abc_52155_new_n7167_));
AND2X2 AND2X2_2488 ( .A(u2__abc_52155_new_n7165_), .B(u2__abc_52155_new_n7168_), .Y(u2__abc_52155_new_n7169_));
AND2X2 AND2X2_2489 ( .A(u2__abc_52155_new_n7170_), .B(u2_remHi_414_), .Y(u2__abc_52155_new_n7171_));
AND2X2 AND2X2_249 ( .A(_abc_73687_new_n1345_), .B(_abc_73687_new_n1344_), .Y(fracta1_59_));
AND2X2 AND2X2_2490 ( .A(u2__abc_52155_new_n7173_), .B(u2_o_414_), .Y(u2__abc_52155_new_n7174_));
AND2X2 AND2X2_2491 ( .A(u2__abc_52155_new_n7172_), .B(u2__abc_52155_new_n7175_), .Y(u2__abc_52155_new_n7176_));
AND2X2 AND2X2_2492 ( .A(u2__abc_52155_new_n7169_), .B(u2__abc_52155_new_n7176_), .Y(u2__abc_52155_new_n7177_));
AND2X2 AND2X2_2493 ( .A(u2__abc_52155_new_n7162_), .B(u2__abc_52155_new_n7177_), .Y(u2__abc_52155_new_n7178_));
AND2X2 AND2X2_2494 ( .A(u2__abc_52155_new_n7147_), .B(u2__abc_52155_new_n7178_), .Y(u2__abc_52155_new_n7179_));
AND2X2 AND2X2_2495 ( .A(u2__abc_52155_new_n7116_), .B(u2__abc_52155_new_n7179_), .Y(u2__abc_52155_new_n7180_));
AND2X2 AND2X2_2496 ( .A(u2__abc_52155_new_n7053_), .B(u2__abc_52155_new_n7180_), .Y(u2__abc_52155_new_n7181_));
AND2X2 AND2X2_2497 ( .A(u2__abc_52155_new_n7182_), .B(u2_remHi_388_), .Y(u2__abc_52155_new_n7183_));
AND2X2 AND2X2_2498 ( .A(u2__abc_52155_new_n7185_), .B(u2_o_388_), .Y(u2__abc_52155_new_n7186_));
AND2X2 AND2X2_2499 ( .A(u2__abc_52155_new_n7184_), .B(u2__abc_52155_new_n7187_), .Y(u2__abc_52155_new_n7188_));
AND2X2 AND2X2_25 ( .A(_abc_73687_new_n753_), .B(sqrto_24_), .Y(\o[60] ));
AND2X2 AND2X2_250 ( .A(_abc_73687_new_n1348_), .B(_abc_73687_new_n1347_), .Y(fracta1_60_));
AND2X2 AND2X2_2500 ( .A(u2__abc_52155_new_n7189_), .B(u2_remHi_389_), .Y(u2__abc_52155_new_n7190_));
AND2X2 AND2X2_2501 ( .A(u2__abc_52155_new_n7192_), .B(u2_o_389_), .Y(u2__abc_52155_new_n7193_));
AND2X2 AND2X2_2502 ( .A(u2__abc_52155_new_n7191_), .B(u2__abc_52155_new_n7194_), .Y(u2__abc_52155_new_n7195_));
AND2X2 AND2X2_2503 ( .A(u2__abc_52155_new_n7188_), .B(u2__abc_52155_new_n7195_), .Y(u2__abc_52155_new_n7196_));
AND2X2 AND2X2_2504 ( .A(u2__abc_52155_new_n7197_), .B(u2_o_387_), .Y(u2__abc_52155_new_n7198_));
AND2X2 AND2X2_2505 ( .A(u2__abc_52155_new_n7200_), .B(u2_remHi_387_), .Y(u2__abc_52155_new_n7201_));
AND2X2 AND2X2_2506 ( .A(u2__abc_52155_new_n7199_), .B(u2__abc_52155_new_n7202_), .Y(u2__abc_52155_new_n7203_));
AND2X2 AND2X2_2507 ( .A(u2__abc_52155_new_n7204_), .B(u2_remHi_386_), .Y(u2__abc_52155_new_n7205_));
AND2X2 AND2X2_2508 ( .A(u2__abc_52155_new_n7207_), .B(u2_o_386_), .Y(u2__abc_52155_new_n7208_));
AND2X2 AND2X2_2509 ( .A(u2__abc_52155_new_n7206_), .B(u2__abc_52155_new_n7209_), .Y(u2__abc_52155_new_n7210_));
AND2X2 AND2X2_251 ( .A(_abc_73687_new_n1351_), .B(_abc_73687_new_n1350_), .Y(fracta1_61_));
AND2X2 AND2X2_2510 ( .A(u2__abc_52155_new_n7203_), .B(u2__abc_52155_new_n7210_), .Y(u2__abc_52155_new_n7211_));
AND2X2 AND2X2_2511 ( .A(u2__abc_52155_new_n7196_), .B(u2__abc_52155_new_n7211_), .Y(u2__abc_52155_new_n7212_));
AND2X2 AND2X2_2512 ( .A(u2__abc_52155_new_n7213_), .B(u2_remHi_384_), .Y(u2__abc_52155_new_n7214_));
AND2X2 AND2X2_2513 ( .A(u2__abc_52155_new_n7216_), .B(u2_o_384_), .Y(u2__abc_52155_new_n7217_));
AND2X2 AND2X2_2514 ( .A(u2__abc_52155_new_n7215_), .B(u2__abc_52155_new_n7218_), .Y(u2__abc_52155_new_n7219_));
AND2X2 AND2X2_2515 ( .A(u2__abc_52155_new_n7220_), .B(u2_o_385_), .Y(u2__abc_52155_new_n7221_));
AND2X2 AND2X2_2516 ( .A(u2__abc_52155_new_n7223_), .B(u2_remHi_385_), .Y(u2__abc_52155_new_n7224_));
AND2X2 AND2X2_2517 ( .A(u2__abc_52155_new_n7222_), .B(u2__abc_52155_new_n7225_), .Y(u2__abc_52155_new_n7226_));
AND2X2 AND2X2_2518 ( .A(u2__abc_52155_new_n7219_), .B(u2__abc_52155_new_n7226_), .Y(u2__abc_52155_new_n7227_));
AND2X2 AND2X2_2519 ( .A(u2__abc_52155_new_n7228_), .B(u2_o_383_), .Y(u2__abc_52155_new_n7229_));
AND2X2 AND2X2_252 ( .A(_abc_73687_new_n1354_), .B(_abc_73687_new_n1353_), .Y(fracta1_62_));
AND2X2 AND2X2_2520 ( .A(u2__abc_52155_new_n7231_), .B(u2_remHi_383_), .Y(u2__abc_52155_new_n7232_));
AND2X2 AND2X2_2521 ( .A(u2__abc_52155_new_n7230_), .B(u2__abc_52155_new_n7233_), .Y(u2__abc_52155_new_n7234_));
AND2X2 AND2X2_2522 ( .A(u2__abc_52155_new_n7235_), .B(u2_remHi_382_), .Y(u2__abc_52155_new_n7236_));
AND2X2 AND2X2_2523 ( .A(u2__abc_52155_new_n7238_), .B(u2_o_382_), .Y(u2__abc_52155_new_n7239_));
AND2X2 AND2X2_2524 ( .A(u2__abc_52155_new_n7237_), .B(u2__abc_52155_new_n7240_), .Y(u2__abc_52155_new_n7241_));
AND2X2 AND2X2_2525 ( .A(u2__abc_52155_new_n7234_), .B(u2__abc_52155_new_n7241_), .Y(u2__abc_52155_new_n7242_));
AND2X2 AND2X2_2526 ( .A(u2__abc_52155_new_n7227_), .B(u2__abc_52155_new_n7242_), .Y(u2__abc_52155_new_n7243_));
AND2X2 AND2X2_2527 ( .A(u2__abc_52155_new_n7212_), .B(u2__abc_52155_new_n7243_), .Y(u2__abc_52155_new_n7244_));
AND2X2 AND2X2_2528 ( .A(u2__abc_52155_new_n7245_), .B(u2_remHi_408_), .Y(u2__abc_52155_new_n7246_));
AND2X2 AND2X2_2529 ( .A(u2__abc_52155_new_n7248_), .B(u2_o_408_), .Y(u2__abc_52155_new_n7249_));
AND2X2 AND2X2_253 ( .A(_abc_73687_new_n1357_), .B(_abc_73687_new_n1356_), .Y(fracta1_63_));
AND2X2 AND2X2_2530 ( .A(u2__abc_52155_new_n7247_), .B(u2__abc_52155_new_n7250_), .Y(u2__abc_52155_new_n7251_));
AND2X2 AND2X2_2531 ( .A(u2__abc_52155_new_n7252_), .B(u2_o_409_), .Y(u2__abc_52155_new_n7253_));
AND2X2 AND2X2_2532 ( .A(u2__abc_52155_new_n7255_), .B(u2_remHi_409_), .Y(u2__abc_52155_new_n7256_));
AND2X2 AND2X2_2533 ( .A(u2__abc_52155_new_n7254_), .B(u2__abc_52155_new_n7257_), .Y(u2__abc_52155_new_n7258_));
AND2X2 AND2X2_2534 ( .A(u2__abc_52155_new_n7251_), .B(u2__abc_52155_new_n7258_), .Y(u2__abc_52155_new_n7259_));
AND2X2 AND2X2_2535 ( .A(u2__abc_52155_new_n7260_), .B(u2_o_407_), .Y(u2__abc_52155_new_n7261_));
AND2X2 AND2X2_2536 ( .A(u2__abc_52155_new_n7263_), .B(u2_remHi_407_), .Y(u2__abc_52155_new_n7264_));
AND2X2 AND2X2_2537 ( .A(u2__abc_52155_new_n7262_), .B(u2__abc_52155_new_n7265_), .Y(u2__abc_52155_new_n7266_));
AND2X2 AND2X2_2538 ( .A(u2__abc_52155_new_n7267_), .B(u2_remHi_406_), .Y(u2__abc_52155_new_n7268_));
AND2X2 AND2X2_2539 ( .A(u2__abc_52155_new_n7270_), .B(u2_o_406_), .Y(u2__abc_52155_new_n7271_));
AND2X2 AND2X2_254 ( .A(_abc_73687_new_n1360_), .B(_abc_73687_new_n1359_), .Y(fracta1_64_));
AND2X2 AND2X2_2540 ( .A(u2__abc_52155_new_n7269_), .B(u2__abc_52155_new_n7272_), .Y(u2__abc_52155_new_n7273_));
AND2X2 AND2X2_2541 ( .A(u2__abc_52155_new_n7266_), .B(u2__abc_52155_new_n7273_), .Y(u2__abc_52155_new_n7274_));
AND2X2 AND2X2_2542 ( .A(u2__abc_52155_new_n7259_), .B(u2__abc_52155_new_n7274_), .Y(u2__abc_52155_new_n7275_));
AND2X2 AND2X2_2543 ( .A(u2__abc_52155_new_n7276_), .B(u2_remHi_412_), .Y(u2__abc_52155_new_n7277_));
AND2X2 AND2X2_2544 ( .A(u2__abc_52155_new_n7279_), .B(u2_o_412_), .Y(u2__abc_52155_new_n7280_));
AND2X2 AND2X2_2545 ( .A(u2__abc_52155_new_n7278_), .B(u2__abc_52155_new_n7281_), .Y(u2__abc_52155_new_n7282_));
AND2X2 AND2X2_2546 ( .A(u2__abc_52155_new_n7283_), .B(u2_remHi_413_), .Y(u2__abc_52155_new_n7284_));
AND2X2 AND2X2_2547 ( .A(u2__abc_52155_new_n7286_), .B(u2_o_413_), .Y(u2__abc_52155_new_n7287_));
AND2X2 AND2X2_2548 ( .A(u2__abc_52155_new_n7285_), .B(u2__abc_52155_new_n7288_), .Y(u2__abc_52155_new_n7289_));
AND2X2 AND2X2_2549 ( .A(u2__abc_52155_new_n7282_), .B(u2__abc_52155_new_n7289_), .Y(u2__abc_52155_new_n7290_));
AND2X2 AND2X2_255 ( .A(_abc_73687_new_n1363_), .B(_abc_73687_new_n1362_), .Y(fracta1_65_));
AND2X2 AND2X2_2550 ( .A(u2__abc_52155_new_n7291_), .B(u2_o_411_), .Y(u2__abc_52155_new_n7292_));
AND2X2 AND2X2_2551 ( .A(u2__abc_52155_new_n7294_), .B(u2_remHi_411_), .Y(u2__abc_52155_new_n7295_));
AND2X2 AND2X2_2552 ( .A(u2__abc_52155_new_n7293_), .B(u2__abc_52155_new_n7296_), .Y(u2__abc_52155_new_n7297_));
AND2X2 AND2X2_2553 ( .A(u2__abc_52155_new_n7298_), .B(u2_remHi_410_), .Y(u2__abc_52155_new_n7299_));
AND2X2 AND2X2_2554 ( .A(u2__abc_52155_new_n7301_), .B(u2_o_410_), .Y(u2__abc_52155_new_n7302_));
AND2X2 AND2X2_2555 ( .A(u2__abc_52155_new_n7300_), .B(u2__abc_52155_new_n7303_), .Y(u2__abc_52155_new_n7304_));
AND2X2 AND2X2_2556 ( .A(u2__abc_52155_new_n7297_), .B(u2__abc_52155_new_n7304_), .Y(u2__abc_52155_new_n7305_));
AND2X2 AND2X2_2557 ( .A(u2__abc_52155_new_n7290_), .B(u2__abc_52155_new_n7305_), .Y(u2__abc_52155_new_n7306_));
AND2X2 AND2X2_2558 ( .A(u2__abc_52155_new_n7275_), .B(u2__abc_52155_new_n7306_), .Y(u2__abc_52155_new_n7307_));
AND2X2 AND2X2_2559 ( .A(u2__abc_52155_new_n7308_), .B(u2_remHi_398_), .Y(u2__abc_52155_new_n7309_));
AND2X2 AND2X2_256 ( .A(_abc_73687_new_n1366_), .B(_abc_73687_new_n1365_), .Y(fracta1_66_));
AND2X2 AND2X2_2560 ( .A(u2__abc_52155_new_n7311_), .B(u2_o_398_), .Y(u2__abc_52155_new_n7312_));
AND2X2 AND2X2_2561 ( .A(u2__abc_52155_new_n7310_), .B(u2__abc_52155_new_n7313_), .Y(u2__abc_52155_new_n7314_));
AND2X2 AND2X2_2562 ( .A(u2__abc_52155_new_n7315_), .B(u2_o_399_), .Y(u2__abc_52155_new_n7316_));
AND2X2 AND2X2_2563 ( .A(u2__abc_52155_new_n7318_), .B(u2_remHi_399_), .Y(u2__abc_52155_new_n7319_));
AND2X2 AND2X2_2564 ( .A(u2__abc_52155_new_n7317_), .B(u2__abc_52155_new_n7320_), .Y(u2__abc_52155_new_n7321_));
AND2X2 AND2X2_2565 ( .A(u2__abc_52155_new_n7314_), .B(u2__abc_52155_new_n7321_), .Y(u2__abc_52155_new_n7322_));
AND2X2 AND2X2_2566 ( .A(u2__abc_52155_new_n7323_), .B(u2_remHi_400_), .Y(u2__abc_52155_new_n7324_));
AND2X2 AND2X2_2567 ( .A(u2__abc_52155_new_n7326_), .B(u2_o_400_), .Y(u2__abc_52155_new_n7327_));
AND2X2 AND2X2_2568 ( .A(u2__abc_52155_new_n7325_), .B(u2__abc_52155_new_n7328_), .Y(u2__abc_52155_new_n7329_));
AND2X2 AND2X2_2569 ( .A(u2__abc_52155_new_n7330_), .B(u2_o_401_), .Y(u2__abc_52155_new_n7331_));
AND2X2 AND2X2_257 ( .A(_abc_73687_new_n1369_), .B(_abc_73687_new_n1368_), .Y(fracta1_67_));
AND2X2 AND2X2_2570 ( .A(u2__abc_52155_new_n7333_), .B(u2_remHi_401_), .Y(u2__abc_52155_new_n7334_));
AND2X2 AND2X2_2571 ( .A(u2__abc_52155_new_n7332_), .B(u2__abc_52155_new_n7335_), .Y(u2__abc_52155_new_n7336_));
AND2X2 AND2X2_2572 ( .A(u2__abc_52155_new_n7329_), .B(u2__abc_52155_new_n7336_), .Y(u2__abc_52155_new_n7337_));
AND2X2 AND2X2_2573 ( .A(u2__abc_52155_new_n7322_), .B(u2__abc_52155_new_n7337_), .Y(u2__abc_52155_new_n7338_));
AND2X2 AND2X2_2574 ( .A(u2__abc_52155_new_n7339_), .B(u2_remHi_404_), .Y(u2__abc_52155_new_n7340_));
AND2X2 AND2X2_2575 ( .A(u2__abc_52155_new_n7342_), .B(u2_o_404_), .Y(u2__abc_52155_new_n7343_));
AND2X2 AND2X2_2576 ( .A(u2__abc_52155_new_n7341_), .B(u2__abc_52155_new_n7344_), .Y(u2__abc_52155_new_n7345_));
AND2X2 AND2X2_2577 ( .A(u2__abc_52155_new_n7346_), .B(u2_remHi_405_), .Y(u2__abc_52155_new_n7347_));
AND2X2 AND2X2_2578 ( .A(u2__abc_52155_new_n7349_), .B(u2_o_405_), .Y(u2__abc_52155_new_n7350_));
AND2X2 AND2X2_2579 ( .A(u2__abc_52155_new_n7348_), .B(u2__abc_52155_new_n7351_), .Y(u2__abc_52155_new_n7352_));
AND2X2 AND2X2_258 ( .A(_abc_73687_new_n1372_), .B(_abc_73687_new_n1371_), .Y(fracta1_68_));
AND2X2 AND2X2_2580 ( .A(u2__abc_52155_new_n7345_), .B(u2__abc_52155_new_n7352_), .Y(u2__abc_52155_new_n7353_));
AND2X2 AND2X2_2581 ( .A(u2__abc_52155_new_n7354_), .B(u2_o_403_), .Y(u2__abc_52155_new_n7355_));
AND2X2 AND2X2_2582 ( .A(u2__abc_52155_new_n7357_), .B(u2_remHi_403_), .Y(u2__abc_52155_new_n7358_));
AND2X2 AND2X2_2583 ( .A(u2__abc_52155_new_n7356_), .B(u2__abc_52155_new_n7359_), .Y(u2__abc_52155_new_n7360_));
AND2X2 AND2X2_2584 ( .A(u2__abc_52155_new_n7361_), .B(u2_remHi_402_), .Y(u2__abc_52155_new_n7362_));
AND2X2 AND2X2_2585 ( .A(u2__abc_52155_new_n7364_), .B(u2_o_402_), .Y(u2__abc_52155_new_n7365_));
AND2X2 AND2X2_2586 ( .A(u2__abc_52155_new_n7363_), .B(u2__abc_52155_new_n7366_), .Y(u2__abc_52155_new_n7367_));
AND2X2 AND2X2_2587 ( .A(u2__abc_52155_new_n7360_), .B(u2__abc_52155_new_n7367_), .Y(u2__abc_52155_new_n7368_));
AND2X2 AND2X2_2588 ( .A(u2__abc_52155_new_n7353_), .B(u2__abc_52155_new_n7368_), .Y(u2__abc_52155_new_n7369_));
AND2X2 AND2X2_2589 ( .A(u2__abc_52155_new_n7338_), .B(u2__abc_52155_new_n7369_), .Y(u2__abc_52155_new_n7370_));
AND2X2 AND2X2_259 ( .A(_abc_73687_new_n1375_), .B(_abc_73687_new_n1374_), .Y(fracta1_69_));
AND2X2 AND2X2_2590 ( .A(u2__abc_52155_new_n7307_), .B(u2__abc_52155_new_n7370_), .Y(u2__abc_52155_new_n7371_));
AND2X2 AND2X2_2591 ( .A(u2__abc_52155_new_n7372_), .B(u2_remHi_392_), .Y(u2__abc_52155_new_n7373_));
AND2X2 AND2X2_2592 ( .A(u2__abc_52155_new_n7375_), .B(u2_o_392_), .Y(u2__abc_52155_new_n7376_));
AND2X2 AND2X2_2593 ( .A(u2__abc_52155_new_n7374_), .B(u2__abc_52155_new_n7377_), .Y(u2__abc_52155_new_n7378_));
AND2X2 AND2X2_2594 ( .A(u2__abc_52155_new_n7379_), .B(u2_o_393_), .Y(u2__abc_52155_new_n7380_));
AND2X2 AND2X2_2595 ( .A(u2__abc_52155_new_n7382_), .B(u2_remHi_393_), .Y(u2__abc_52155_new_n7383_));
AND2X2 AND2X2_2596 ( .A(u2__abc_52155_new_n7381_), .B(u2__abc_52155_new_n7384_), .Y(u2__abc_52155_new_n7385_));
AND2X2 AND2X2_2597 ( .A(u2__abc_52155_new_n7378_), .B(u2__abc_52155_new_n7385_), .Y(u2__abc_52155_new_n7386_));
AND2X2 AND2X2_2598 ( .A(u2__abc_52155_new_n7387_), .B(u2_remHi_390_), .Y(u2__abc_52155_new_n7388_));
AND2X2 AND2X2_2599 ( .A(u2__abc_52155_new_n7390_), .B(u2_o_390_), .Y(u2__abc_52155_new_n7391_));
AND2X2 AND2X2_26 ( .A(_abc_73687_new_n753_), .B(sqrto_25_), .Y(\o[61] ));
AND2X2 AND2X2_260 ( .A(_abc_73687_new_n1378_), .B(_abc_73687_new_n1377_), .Y(fracta1_70_));
AND2X2 AND2X2_2600 ( .A(u2__abc_52155_new_n7389_), .B(u2__abc_52155_new_n7392_), .Y(u2__abc_52155_new_n7393_));
AND2X2 AND2X2_2601 ( .A(u2__abc_52155_new_n7394_), .B(u2_o_391_), .Y(u2__abc_52155_new_n7395_));
AND2X2 AND2X2_2602 ( .A(u2__abc_52155_new_n7397_), .B(u2_remHi_391_), .Y(u2__abc_52155_new_n7398_));
AND2X2 AND2X2_2603 ( .A(u2__abc_52155_new_n7396_), .B(u2__abc_52155_new_n7399_), .Y(u2__abc_52155_new_n7400_));
AND2X2 AND2X2_2604 ( .A(u2__abc_52155_new_n7393_), .B(u2__abc_52155_new_n7400_), .Y(u2__abc_52155_new_n7401_));
AND2X2 AND2X2_2605 ( .A(u2__abc_52155_new_n7386_), .B(u2__abc_52155_new_n7401_), .Y(u2__abc_52155_new_n7402_));
AND2X2 AND2X2_2606 ( .A(u2__abc_52155_new_n7403_), .B(u2_remHi_396_), .Y(u2__abc_52155_new_n7404_));
AND2X2 AND2X2_2607 ( .A(u2__abc_52155_new_n7406_), .B(u2_o_396_), .Y(u2__abc_52155_new_n7407_));
AND2X2 AND2X2_2608 ( .A(u2__abc_52155_new_n7405_), .B(u2__abc_52155_new_n7408_), .Y(u2__abc_52155_new_n7409_));
AND2X2 AND2X2_2609 ( .A(u2__abc_52155_new_n7410_), .B(u2_remHi_397_), .Y(u2__abc_52155_new_n7411_));
AND2X2 AND2X2_261 ( .A(_abc_73687_new_n1381_), .B(_abc_73687_new_n1380_), .Y(fracta1_71_));
AND2X2 AND2X2_2610 ( .A(u2__abc_52155_new_n7413_), .B(u2_o_397_), .Y(u2__abc_52155_new_n7414_));
AND2X2 AND2X2_2611 ( .A(u2__abc_52155_new_n7412_), .B(u2__abc_52155_new_n7415_), .Y(u2__abc_52155_new_n7416_));
AND2X2 AND2X2_2612 ( .A(u2__abc_52155_new_n7409_), .B(u2__abc_52155_new_n7416_), .Y(u2__abc_52155_new_n7417_));
AND2X2 AND2X2_2613 ( .A(u2__abc_52155_new_n7418_), .B(u2_o_395_), .Y(u2__abc_52155_new_n7419_));
AND2X2 AND2X2_2614 ( .A(u2__abc_52155_new_n7421_), .B(u2_remHi_395_), .Y(u2__abc_52155_new_n7422_));
AND2X2 AND2X2_2615 ( .A(u2__abc_52155_new_n7420_), .B(u2__abc_52155_new_n7423_), .Y(u2__abc_52155_new_n7424_));
AND2X2 AND2X2_2616 ( .A(u2__abc_52155_new_n7425_), .B(u2_remHi_394_), .Y(u2__abc_52155_new_n7426_));
AND2X2 AND2X2_2617 ( .A(u2__abc_52155_new_n7428_), .B(u2_o_394_), .Y(u2__abc_52155_new_n7429_));
AND2X2 AND2X2_2618 ( .A(u2__abc_52155_new_n7427_), .B(u2__abc_52155_new_n7430_), .Y(u2__abc_52155_new_n7431_));
AND2X2 AND2X2_2619 ( .A(u2__abc_52155_new_n7424_), .B(u2__abc_52155_new_n7431_), .Y(u2__abc_52155_new_n7432_));
AND2X2 AND2X2_262 ( .A(_abc_73687_new_n1384_), .B(_abc_73687_new_n1383_), .Y(fracta1_72_));
AND2X2 AND2X2_2620 ( .A(u2__abc_52155_new_n7417_), .B(u2__abc_52155_new_n7432_), .Y(u2__abc_52155_new_n7433_));
AND2X2 AND2X2_2621 ( .A(u2__abc_52155_new_n7402_), .B(u2__abc_52155_new_n7433_), .Y(u2__abc_52155_new_n7434_));
AND2X2 AND2X2_2622 ( .A(u2__abc_52155_new_n7371_), .B(u2__abc_52155_new_n7434_), .Y(u2__abc_52155_new_n7435_));
AND2X2 AND2X2_2623 ( .A(u2__abc_52155_new_n7435_), .B(u2__abc_52155_new_n7244_), .Y(u2__abc_52155_new_n7436_));
AND2X2 AND2X2_2624 ( .A(u2__abc_52155_new_n7436_), .B(u2__abc_52155_new_n7181_), .Y(u2__abc_52155_new_n7437_));
AND2X2 AND2X2_2625 ( .A(u2__abc_52155_new_n7233_), .B(u2__abc_52155_new_n7239_), .Y(u2__abc_52155_new_n7440_));
AND2X2 AND2X2_2626 ( .A(u2__abc_52155_new_n7441_), .B(u2__abc_52155_new_n7227_), .Y(u2__abc_52155_new_n7442_));
AND2X2 AND2X2_2627 ( .A(u2__abc_52155_new_n7225_), .B(u2__abc_52155_new_n7217_), .Y(u2__abc_52155_new_n7443_));
AND2X2 AND2X2_2628 ( .A(u2__abc_52155_new_n7445_), .B(u2__abc_52155_new_n7212_), .Y(u2__abc_52155_new_n7446_));
AND2X2 AND2X2_2629 ( .A(u2__abc_52155_new_n7202_), .B(u2__abc_52155_new_n7208_), .Y(u2__abc_52155_new_n7447_));
AND2X2 AND2X2_263 ( .A(_abc_73687_new_n1387_), .B(_abc_73687_new_n1386_), .Y(fracta1_73_));
AND2X2 AND2X2_2630 ( .A(u2__abc_52155_new_n7448_), .B(u2__abc_52155_new_n7196_), .Y(u2__abc_52155_new_n7449_));
AND2X2 AND2X2_2631 ( .A(u2__abc_52155_new_n7191_), .B(u2__abc_52155_new_n7186_), .Y(u2__abc_52155_new_n7450_));
AND2X2 AND2X2_2632 ( .A(u2__abc_52155_new_n7453_), .B(u2__abc_52155_new_n7434_), .Y(u2__abc_52155_new_n7454_));
AND2X2 AND2X2_2633 ( .A(u2__abc_52155_new_n7423_), .B(u2__abc_52155_new_n7429_), .Y(u2__abc_52155_new_n7455_));
AND2X2 AND2X2_2634 ( .A(u2__abc_52155_new_n7456_), .B(u2__abc_52155_new_n7417_), .Y(u2__abc_52155_new_n7457_));
AND2X2 AND2X2_2635 ( .A(u2__abc_52155_new_n7412_), .B(u2__abc_52155_new_n7407_), .Y(u2__abc_52155_new_n7458_));
AND2X2 AND2X2_2636 ( .A(u2__abc_52155_new_n7399_), .B(u2__abc_52155_new_n7391_), .Y(u2__abc_52155_new_n7461_));
AND2X2 AND2X2_2637 ( .A(u2__abc_52155_new_n7462_), .B(u2__abc_52155_new_n7386_), .Y(u2__abc_52155_new_n7463_));
AND2X2 AND2X2_2638 ( .A(u2__abc_52155_new_n7384_), .B(u2__abc_52155_new_n7376_), .Y(u2__abc_52155_new_n7464_));
AND2X2 AND2X2_2639 ( .A(u2__abc_52155_new_n7466_), .B(u2__abc_52155_new_n7433_), .Y(u2__abc_52155_new_n7467_));
AND2X2 AND2X2_264 ( .A(_abc_73687_new_n1390_), .B(_abc_73687_new_n1389_), .Y(fracta1_74_));
AND2X2 AND2X2_2640 ( .A(u2__abc_52155_new_n7469_), .B(u2__abc_52155_new_n7371_), .Y(u2__abc_52155_new_n7470_));
AND2X2 AND2X2_2641 ( .A(u2__abc_52155_new_n7265_), .B(u2__abc_52155_new_n7271_), .Y(u2__abc_52155_new_n7471_));
AND2X2 AND2X2_2642 ( .A(u2__abc_52155_new_n7472_), .B(u2__abc_52155_new_n7259_), .Y(u2__abc_52155_new_n7473_));
AND2X2 AND2X2_2643 ( .A(u2__abc_52155_new_n7257_), .B(u2__abc_52155_new_n7249_), .Y(u2__abc_52155_new_n7474_));
AND2X2 AND2X2_2644 ( .A(u2__abc_52155_new_n7476_), .B(u2__abc_52155_new_n7306_), .Y(u2__abc_52155_new_n7477_));
AND2X2 AND2X2_2645 ( .A(u2__abc_52155_new_n7296_), .B(u2__abc_52155_new_n7302_), .Y(u2__abc_52155_new_n7478_));
AND2X2 AND2X2_2646 ( .A(u2__abc_52155_new_n7479_), .B(u2__abc_52155_new_n7290_), .Y(u2__abc_52155_new_n7480_));
AND2X2 AND2X2_2647 ( .A(u2__abc_52155_new_n7285_), .B(u2__abc_52155_new_n7280_), .Y(u2__abc_52155_new_n7481_));
AND2X2 AND2X2_2648 ( .A(u2__abc_52155_new_n7320_), .B(u2__abc_52155_new_n7312_), .Y(u2__abc_52155_new_n7485_));
AND2X2 AND2X2_2649 ( .A(u2__abc_52155_new_n7486_), .B(u2__abc_52155_new_n7337_), .Y(u2__abc_52155_new_n7487_));
AND2X2 AND2X2_265 ( .A(_abc_73687_new_n1393_), .B(_abc_73687_new_n1392_), .Y(fracta1_75_));
AND2X2 AND2X2_2650 ( .A(u2__abc_52155_new_n7335_), .B(u2__abc_52155_new_n7327_), .Y(u2__abc_52155_new_n7488_));
AND2X2 AND2X2_2651 ( .A(u2__abc_52155_new_n7490_), .B(u2__abc_52155_new_n7369_), .Y(u2__abc_52155_new_n7491_));
AND2X2 AND2X2_2652 ( .A(u2__abc_52155_new_n7359_), .B(u2__abc_52155_new_n7365_), .Y(u2__abc_52155_new_n7492_));
AND2X2 AND2X2_2653 ( .A(u2__abc_52155_new_n7493_), .B(u2__abc_52155_new_n7353_), .Y(u2__abc_52155_new_n7494_));
AND2X2 AND2X2_2654 ( .A(u2__abc_52155_new_n7348_), .B(u2__abc_52155_new_n7343_), .Y(u2__abc_52155_new_n7495_));
AND2X2 AND2X2_2655 ( .A(u2__abc_52155_new_n7498_), .B(u2__abc_52155_new_n7307_), .Y(u2__abc_52155_new_n7499_));
AND2X2 AND2X2_2656 ( .A(u2__abc_52155_new_n7501_), .B(u2__abc_52155_new_n7181_), .Y(u2__abc_52155_new_n7502_));
AND2X2 AND2X2_2657 ( .A(u2__abc_52155_new_n7168_), .B(u2__abc_52155_new_n7174_), .Y(u2__abc_52155_new_n7503_));
AND2X2 AND2X2_2658 ( .A(u2__abc_52155_new_n7504_), .B(u2__abc_52155_new_n7162_), .Y(u2__abc_52155_new_n7505_));
AND2X2 AND2X2_2659 ( .A(u2__abc_52155_new_n7160_), .B(u2__abc_52155_new_n7152_), .Y(u2__abc_52155_new_n7506_));
AND2X2 AND2X2_266 ( .A(_abc_73687_new_n1396_), .B(_abc_73687_new_n1395_), .Y(fracta1_76_));
AND2X2 AND2X2_2660 ( .A(u2__abc_52155_new_n7508_), .B(u2__abc_52155_new_n7147_), .Y(u2__abc_52155_new_n7509_));
AND2X2 AND2X2_2661 ( .A(u2__abc_52155_new_n7137_), .B(u2__abc_52155_new_n7143_), .Y(u2__abc_52155_new_n7510_));
AND2X2 AND2X2_2662 ( .A(u2__abc_52155_new_n7511_), .B(u2__abc_52155_new_n7131_), .Y(u2__abc_52155_new_n7512_));
AND2X2 AND2X2_2663 ( .A(u2__abc_52155_new_n7126_), .B(u2__abc_52155_new_n7121_), .Y(u2__abc_52155_new_n7513_));
AND2X2 AND2X2_2664 ( .A(u2__abc_52155_new_n7516_), .B(u2__abc_52155_new_n7116_), .Y(u2__abc_52155_new_n7517_));
AND2X2 AND2X2_2665 ( .A(u2__abc_52155_new_n7081_), .B(u2__abc_52155_new_n7073_), .Y(u2__abc_52155_new_n7518_));
AND2X2 AND2X2_2666 ( .A(u2__abc_52155_new_n7519_), .B(u2__abc_52155_new_n7068_), .Y(u2__abc_52155_new_n7520_));
AND2X2 AND2X2_2667 ( .A(u2__abc_52155_new_n7066_), .B(u2__abc_52155_new_n7058_), .Y(u2__abc_52155_new_n7521_));
AND2X2 AND2X2_2668 ( .A(u2__abc_52155_new_n7523_), .B(u2__abc_52155_new_n7115_), .Y(u2__abc_52155_new_n7524_));
AND2X2 AND2X2_2669 ( .A(u2__abc_52155_new_n7105_), .B(u2__abc_52155_new_n7111_), .Y(u2__abc_52155_new_n7525_));
AND2X2 AND2X2_267 ( .A(_abc_73687_new_n1399_), .B(_abc_73687_new_n1398_), .Y(fracta1_77_));
AND2X2 AND2X2_2670 ( .A(u2__abc_52155_new_n7526_), .B(u2__abc_52155_new_n7099_), .Y(u2__abc_52155_new_n7527_));
AND2X2 AND2X2_2671 ( .A(u2__abc_52155_new_n7094_), .B(u2__abc_52155_new_n7089_), .Y(u2__abc_52155_new_n7528_));
AND2X2 AND2X2_2672 ( .A(u2__abc_52155_new_n7532_), .B(u2__abc_52155_new_n7053_), .Y(u2__abc_52155_new_n7533_));
AND2X2 AND2X2_2673 ( .A(u2__abc_52155_new_n6970_), .B(u2__abc_52155_new_n6962_), .Y(u2__abc_52155_new_n7534_));
AND2X2 AND2X2_2674 ( .A(u2__abc_52155_new_n7535_), .B(u2__abc_52155_new_n6987_), .Y(u2__abc_52155_new_n7536_));
AND2X2 AND2X2_2675 ( .A(u2__abc_52155_new_n6985_), .B(u2__abc_52155_new_n6977_), .Y(u2__abc_52155_new_n7537_));
AND2X2 AND2X2_2676 ( .A(u2__abc_52155_new_n7539_), .B(u2__abc_52155_new_n6957_), .Y(u2__abc_52155_new_n7540_));
AND2X2 AND2X2_2677 ( .A(u2__abc_52155_new_n6947_), .B(u2__abc_52155_new_n6953_), .Y(u2__abc_52155_new_n7541_));
AND2X2 AND2X2_2678 ( .A(u2__abc_52155_new_n7542_), .B(u2__abc_52155_new_n6941_), .Y(u2__abc_52155_new_n7543_));
AND2X2 AND2X2_2679 ( .A(u2__abc_52155_new_n6939_), .B(u2__abc_52155_new_n6931_), .Y(u2__abc_52155_new_n7544_));
AND2X2 AND2X2_268 ( .A(_abc_73687_new_n1402_), .B(_abc_73687_new_n1401_), .Y(fracta1_78_));
AND2X2 AND2X2_2680 ( .A(u2__abc_52155_new_n7033_), .B(u2__abc_52155_new_n7025_), .Y(u2__abc_52155_new_n7548_));
AND2X2 AND2X2_2681 ( .A(u2__abc_52155_new_n7549_), .B(u2__abc_52155_new_n7050_), .Y(u2__abc_52155_new_n7550_));
AND2X2 AND2X2_2682 ( .A(u2__abc_52155_new_n7048_), .B(u2__abc_52155_new_n7040_), .Y(u2__abc_52155_new_n7551_));
AND2X2 AND2X2_2683 ( .A(u2__abc_52155_new_n7553_), .B(u2__abc_52155_new_n7020_), .Y(u2__abc_52155_new_n7554_));
AND2X2 AND2X2_2684 ( .A(u2__abc_52155_new_n7010_), .B(u2__abc_52155_new_n7016_), .Y(u2__abc_52155_new_n7555_));
AND2X2 AND2X2_2685 ( .A(u2__abc_52155_new_n7556_), .B(u2__abc_52155_new_n7004_), .Y(u2__abc_52155_new_n7557_));
AND2X2 AND2X2_2686 ( .A(u2__abc_52155_new_n7003_), .B(u2__abc_52155_new_n6994_), .Y(u2__abc_52155_new_n7558_));
AND2X2 AND2X2_2687 ( .A(u2__abc_52155_new_n7561_), .B(u2__abc_52155_new_n6989_), .Y(u2__abc_52155_new_n7562_));
AND2X2 AND2X2_2688 ( .A(u2__abc_52155_new_n7439_), .B(u2__abc_52155_new_n7566_), .Y(u2__abc_52155_new_n7567_));
AND2X2 AND2X2_2689 ( .A(u2__abc_52155_new_n3023_), .B(u2__abc_52155_new_n3030_), .Y(u2__abc_52155_new_n7569_));
AND2X2 AND2X2_269 ( .A(_abc_73687_new_n1405_), .B(_abc_73687_new_n1404_), .Y(fracta1_79_));
AND2X2 AND2X2_2690 ( .A(u2__abc_52155_new_n7571_), .B(u2__abc_52155_new_n3017_), .Y(u2__abc_52155_new_n7572_));
AND2X2 AND2X2_2691 ( .A(u2__abc_52155_new_n3009_), .B(u2__abc_52155_new_n3012_), .Y(u2__abc_52155_new_n7573_));
AND2X2 AND2X2_2692 ( .A(u2__abc_52155_new_n7568_), .B(u2__abc_52155_new_n7576_), .Y(u2__abc_52155_new_n7577_));
AND2X2 AND2X2_2693 ( .A(u2__abc_52155_new_n4130_), .B(u2__abc_52155_new_n3893_), .Y(u2__abc_52155_new_n7578_));
AND2X2 AND2X2_2694 ( .A(u2__abc_52155_new_n4542_), .B(u2__abc_52155_new_n4923_), .Y(u2__abc_52155_new_n7579_));
AND2X2 AND2X2_2695 ( .A(u2__abc_52155_new_n7578_), .B(u2__abc_52155_new_n7579_), .Y(u2__abc_52155_new_n7580_));
AND2X2 AND2X2_2696 ( .A(u2__abc_52155_new_n4792_), .B(u2__abc_52155_new_n7147_), .Y(u2__abc_52155_new_n7581_));
AND2X2 AND2X2_2697 ( .A(u2__abc_52155_new_n7581_), .B(u2__abc_52155_new_n7178_), .Y(u2__abc_52155_new_n7582_));
AND2X2 AND2X2_2698 ( .A(u2__abc_52155_new_n7584_), .B(u2__abc_52155_new_n7585_), .Y(u2__abc_52155_new_n7586_));
AND2X2 AND2X2_2699 ( .A(u2__abc_52155_new_n7586_), .B(u2_remHiShift_0_), .Y(u2__abc_52155_new_n7587_));
AND2X2 AND2X2_27 ( .A(_abc_73687_new_n753_), .B(sqrto_26_), .Y(\o[62] ));
AND2X2 AND2X2_270 ( .A(_abc_73687_new_n1408_), .B(_abc_73687_new_n1407_), .Y(fracta1_80_));
AND2X2 AND2X2_2700 ( .A(u2__abc_52155_new_n7583_), .B(u2__abc_52155_new_n7587_), .Y(u2__abc_52155_new_n7588_));
AND2X2 AND2X2_2701 ( .A(u2__abc_52155_new_n7588_), .B(u2__abc_52155_new_n3033_), .Y(u2__abc_52155_new_n7589_));
AND2X2 AND2X2_2702 ( .A(u2__abc_52155_new_n7590_), .B(u2__abc_52155_new_n4764_), .Y(u2__abc_52155_new_n7591_));
AND2X2 AND2X2_2703 ( .A(u2__abc_52155_new_n7591_), .B(u2__abc_52155_new_n7589_), .Y(u2__abc_52155_new_n7592_));
AND2X2 AND2X2_2704 ( .A(u2__abc_52155_new_n7592_), .B(u2__abc_52155_new_n7582_), .Y(u2__abc_52155_new_n7593_));
AND2X2 AND2X2_2705 ( .A(u2__abc_52155_new_n3278_), .B(u2__abc_52155_new_n3446_), .Y(u2__abc_52155_new_n7594_));
AND2X2 AND2X2_2706 ( .A(u2__abc_52155_new_n7593_), .B(u2__abc_52155_new_n7594_), .Y(u2__abc_52155_new_n7595_));
AND2X2 AND2X2_2707 ( .A(u2__abc_52155_new_n7595_), .B(u2__abc_52155_new_n7580_), .Y(u2__abc_52155_new_n7596_));
AND2X2 AND2X2_2708 ( .A(u2__abc_52155_new_n6091_), .B(u2__abc_52155_new_n6475_), .Y(u2__abc_52155_new_n7597_));
AND2X2 AND2X2_2709 ( .A(u2__abc_52155_new_n7597_), .B(u2__abc_52155_new_n7053_), .Y(u2__abc_52155_new_n7598_));
AND2X2 AND2X2_271 ( .A(_abc_73687_new_n1411_), .B(_abc_73687_new_n1410_), .Y(fracta1_81_));
AND2X2 AND2X2_2710 ( .A(u2__abc_52155_new_n5047_), .B(u2__abc_52155_new_n5709_), .Y(u2__abc_52155_new_n7599_));
AND2X2 AND2X2_2711 ( .A(u2__abc_52155_new_n5836_), .B(u2__abc_52155_new_n5964_), .Y(u2__abc_52155_new_n7600_));
AND2X2 AND2X2_2712 ( .A(u2__abc_52155_new_n7599_), .B(u2__abc_52155_new_n7600_), .Y(u2__abc_52155_new_n7601_));
AND2X2 AND2X2_2713 ( .A(u2__abc_52155_new_n7601_), .B(u2__abc_52155_new_n7598_), .Y(u2__abc_52155_new_n7602_));
AND2X2 AND2X2_2714 ( .A(u2__abc_52155_new_n7596_), .B(u2__abc_52155_new_n7602_), .Y(u2__abc_52155_new_n7603_));
AND2X2 AND2X2_2715 ( .A(u2__abc_52155_new_n7116_), .B(u2__abc_52155_new_n7244_), .Y(u2__abc_52155_new_n7604_));
AND2X2 AND2X2_2716 ( .A(u2__abc_52155_new_n6602_), .B(u2__abc_52155_new_n7604_), .Y(u2__abc_52155_new_n7605_));
AND2X2 AND2X2_2717 ( .A(u2__abc_52155_new_n5285_), .B(u2__abc_52155_new_n7605_), .Y(u2__abc_52155_new_n7606_));
AND2X2 AND2X2_2718 ( .A(u2__abc_52155_new_n7606_), .B(u2__abc_52155_new_n7435_), .Y(u2__abc_52155_new_n7607_));
AND2X2 AND2X2_2719 ( .A(u2__abc_52155_new_n3768_), .B(u2__abc_52155_new_n3957_), .Y(u2__abc_52155_new_n7608_));
AND2X2 AND2X2_272 ( .A(_abc_73687_new_n1414_), .B(_abc_73687_new_n1413_), .Y(fracta1_82_));
AND2X2 AND2X2_2720 ( .A(u2__abc_52155_new_n4017_), .B(u2__abc_52155_new_n4351_), .Y(u2__abc_52155_new_n7609_));
AND2X2 AND2X2_2721 ( .A(u2__abc_52155_new_n7609_), .B(u2__abc_52155_new_n7608_), .Y(u2__abc_52155_new_n7610_));
AND2X2 AND2X2_2722 ( .A(u2__abc_52155_new_n3506_), .B(u2__abc_52155_new_n3089_), .Y(u2__abc_52155_new_n7611_));
AND2X2 AND2X2_2723 ( .A(u2__abc_52155_new_n3557_), .B(u2__abc_52155_new_n3705_), .Y(u2__abc_52155_new_n7612_));
AND2X2 AND2X2_2724 ( .A(u2__abc_52155_new_n7612_), .B(u2__abc_52155_new_n7611_), .Y(u2__abc_52155_new_n7613_));
AND2X2 AND2X2_2725 ( .A(u2__abc_52155_new_n7613_), .B(u2__abc_52155_new_n7610_), .Y(u2__abc_52155_new_n7614_));
AND2X2 AND2X2_2726 ( .A(u2__abc_52155_new_n4414_), .B(u2__abc_52155_new_n4606_), .Y(u2__abc_52155_new_n7615_));
AND2X2 AND2X2_2727 ( .A(u2__abc_52155_new_n4669_), .B(u2__abc_52155_new_n4733_), .Y(u2__abc_52155_new_n7616_));
AND2X2 AND2X2_2728 ( .A(u2__abc_52155_new_n7615_), .B(u2__abc_52155_new_n7616_), .Y(u2__abc_52155_new_n7617_));
AND2X2 AND2X2_2729 ( .A(u2__abc_52155_new_n6348_), .B(u2__abc_52155_new_n7617_), .Y(u2__abc_52155_new_n7618_));
AND2X2 AND2X2_273 ( .A(_abc_73687_new_n1417_), .B(_abc_73687_new_n1416_), .Y(fracta1_83_));
AND2X2 AND2X2_2730 ( .A(u2__abc_52155_new_n7614_), .B(u2__abc_52155_new_n7618_), .Y(u2__abc_52155_new_n7619_));
AND2X2 AND2X2_2731 ( .A(u2__abc_52155_new_n7619_), .B(u2__abc_52155_new_n7607_), .Y(u2__abc_52155_new_n7620_));
AND2X2 AND2X2_2732 ( .A(u2__abc_52155_new_n7603_), .B(u2__abc_52155_new_n7620_), .Y(u2__abc_52155_new_n7621_));
AND2X2 AND2X2_2733 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHiShift_0_), .Y(u2__abc_52155_new_n7624_));
AND2X2 AND2X2_2734 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7625_), .Y(u2__abc_52155_new_n7626_));
AND2X2 AND2X2_2735 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3116_), .Y(u2__abc_52155_new_n7629_));
AND2X2 AND2X2_2736 ( .A(u2__abc_52155_new_n7630_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7631_));
AND2X2 AND2X2_2737 ( .A(u2__abc_52155_new_n7628_), .B(u2__abc_52155_new_n7631_), .Y(u2__abc_52155_new_n7632_));
AND2X2 AND2X2_2738 ( .A(u2__abc_52155_new_n7633_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__0_));
AND2X2 AND2X2_2739 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_1_), .Y(u2__abc_52155_new_n7635_));
AND2X2 AND2X2_274 ( .A(_abc_73687_new_n1420_), .B(_abc_73687_new_n1419_), .Y(fracta1_84_));
AND2X2 AND2X2_2740 ( .A(u2__abc_52155_new_n7636_), .B(u2__abc_52155_new_n7637_), .Y(u2__abc_52155_new_n7638_));
AND2X2 AND2X2_2741 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7638_), .Y(u2__abc_52155_new_n7639_));
AND2X2 AND2X2_2742 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHiShift_1_), .Y(u2__abc_52155_new_n7640_));
AND2X2 AND2X2_2743 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3119_), .Y(u2__abc_52155_new_n7643_));
AND2X2 AND2X2_2744 ( .A(u2__abc_52155_new_n7644_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7645_));
AND2X2 AND2X2_2745 ( .A(u2__abc_52155_new_n7642_), .B(u2__abc_52155_new_n7645_), .Y(u2__abc_52155_new_n7646_));
AND2X2 AND2X2_2746 ( .A(u2__abc_52155_new_n7647_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__1_));
AND2X2 AND2X2_2747 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_2_), .Y(u2__abc_52155_new_n7649_));
AND2X2 AND2X2_2748 ( .A(u2__abc_52155_new_n7636_), .B(u2__abc_52155_new_n7584_), .Y(u2__abc_52155_new_n7651_));
AND2X2 AND2X2_2749 ( .A(u2__abc_52155_new_n7652_), .B(u2__abc_52155_new_n7650_), .Y(u2__abc_52155_new_n7653_));
AND2X2 AND2X2_275 ( .A(_abc_73687_new_n1423_), .B(_abc_73687_new_n1422_), .Y(fracta1_85_));
AND2X2 AND2X2_2750 ( .A(u2__abc_52155_new_n7654_), .B(u2__abc_52155_new_n7655_), .Y(u2__abc_52155_new_n7656_));
AND2X2 AND2X2_2751 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7656_), .Y(u2__abc_52155_new_n7657_));
AND2X2 AND2X2_2752 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_0_), .Y(u2__abc_52155_new_n7658_));
AND2X2 AND2X2_2753 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3109_), .Y(u2__abc_52155_new_n7661_));
AND2X2 AND2X2_2754 ( .A(u2__abc_52155_new_n7662_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7663_));
AND2X2 AND2X2_2755 ( .A(u2__abc_52155_new_n7660_), .B(u2__abc_52155_new_n7663_), .Y(u2__abc_52155_new_n7664_));
AND2X2 AND2X2_2756 ( .A(u2__abc_52155_new_n7665_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__2_));
AND2X2 AND2X2_2757 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_3_), .Y(u2__abc_52155_new_n7667_));
AND2X2 AND2X2_2758 ( .A(u2__abc_52155_new_n7668_), .B(u2__abc_52155_new_n3115_), .Y(u2__abc_52155_new_n7671_));
AND2X2 AND2X2_2759 ( .A(u2__abc_52155_new_n7652_), .B(u2__abc_52155_new_n7583_), .Y(u2__abc_52155_new_n7672_));
AND2X2 AND2X2_276 ( .A(_abc_73687_new_n1426_), .B(_abc_73687_new_n1425_), .Y(fracta1_86_));
AND2X2 AND2X2_2760 ( .A(u2__abc_52155_new_n7674_), .B(u2__abc_52155_new_n7670_), .Y(u2__abc_52155_new_n7675_));
AND2X2 AND2X2_2761 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7675_), .Y(u2__abc_52155_new_n7676_));
AND2X2 AND2X2_2762 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_1_), .Y(u2__abc_52155_new_n7677_));
AND2X2 AND2X2_2763 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3104_), .Y(u2__abc_52155_new_n7680_));
AND2X2 AND2X2_2764 ( .A(u2__abc_52155_new_n7681_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7682_));
AND2X2 AND2X2_2765 ( .A(u2__abc_52155_new_n7679_), .B(u2__abc_52155_new_n7682_), .Y(u2__abc_52155_new_n7683_));
AND2X2 AND2X2_2766 ( .A(u2__abc_52155_new_n7684_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__3_));
AND2X2 AND2X2_2767 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_4_), .Y(u2__abc_52155_new_n7686_));
AND2X2 AND2X2_2768 ( .A(u2__abc_52155_new_n7688_), .B(u2__abc_52155_new_n7687_), .Y(u2__abc_52155_new_n7690_));
AND2X2 AND2X2_2769 ( .A(u2__abc_52155_new_n7691_), .B(u2__abc_52155_new_n7689_), .Y(u2__abc_52155_new_n7692_));
AND2X2 AND2X2_277 ( .A(_abc_73687_new_n1429_), .B(_abc_73687_new_n1428_), .Y(fracta1_87_));
AND2X2 AND2X2_2770 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7692_), .Y(u2__abc_52155_new_n7693_));
AND2X2 AND2X2_2771 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_2_), .Y(u2__abc_52155_new_n7694_));
AND2X2 AND2X2_2772 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3093_), .Y(u2__abc_52155_new_n7697_));
AND2X2 AND2X2_2773 ( .A(u2__abc_52155_new_n7698_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7699_));
AND2X2 AND2X2_2774 ( .A(u2__abc_52155_new_n7696_), .B(u2__abc_52155_new_n7699_), .Y(u2__abc_52155_new_n7700_));
AND2X2 AND2X2_2775 ( .A(u2__abc_52155_new_n7701_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__4_));
AND2X2 AND2X2_2776 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_5_), .Y(u2__abc_52155_new_n7703_));
AND2X2 AND2X2_2777 ( .A(u2__abc_52155_new_n7691_), .B(u2__abc_52155_new_n7705_), .Y(u2__abc_52155_new_n7706_));
AND2X2 AND2X2_2778 ( .A(u2__abc_52155_new_n7708_), .B(u2__abc_52155_new_n7709_), .Y(u2__abc_52155_new_n7710_));
AND2X2 AND2X2_2779 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7710_), .Y(u2__abc_52155_new_n7711_));
AND2X2 AND2X2_278 ( .A(_abc_73687_new_n1432_), .B(_abc_73687_new_n1431_), .Y(fracta1_88_));
AND2X2 AND2X2_2780 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_3_), .Y(u2__abc_52155_new_n7712_));
AND2X2 AND2X2_2781 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3096_), .Y(u2__abc_52155_new_n7715_));
AND2X2 AND2X2_2782 ( .A(u2__abc_52155_new_n7716_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7717_));
AND2X2 AND2X2_2783 ( .A(u2__abc_52155_new_n7714_), .B(u2__abc_52155_new_n7717_), .Y(u2__abc_52155_new_n7718_));
AND2X2 AND2X2_2784 ( .A(u2__abc_52155_new_n7719_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__5_));
AND2X2 AND2X2_2785 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_6_), .Y(u2__abc_52155_new_n7721_));
AND2X2 AND2X2_2786 ( .A(u2__abc_52155_new_n7690_), .B(u2__abc_52155_new_n7704_), .Y(u2__abc_52155_new_n7723_));
AND2X2 AND2X2_2787 ( .A(u2__abc_52155_new_n7724_), .B(u2__abc_52155_new_n3134_), .Y(u2__abc_52155_new_n7725_));
AND2X2 AND2X2_2788 ( .A(u2__abc_52155_new_n7726_), .B(u2__abc_52155_new_n7722_), .Y(u2__abc_52155_new_n7728_));
AND2X2 AND2X2_2789 ( .A(u2__abc_52155_new_n7729_), .B(u2__abc_52155_new_n7727_), .Y(u2__abc_52155_new_n7730_));
AND2X2 AND2X2_279 ( .A(_abc_73687_new_n1435_), .B(_abc_73687_new_n1434_), .Y(fracta1_89_));
AND2X2 AND2X2_2790 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7730_), .Y(u2__abc_52155_new_n7731_));
AND2X2 AND2X2_2791 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_4_), .Y(u2__abc_52155_new_n7732_));
AND2X2 AND2X2_2792 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3082_), .Y(u2__abc_52155_new_n7735_));
AND2X2 AND2X2_2793 ( .A(u2__abc_52155_new_n7736_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7737_));
AND2X2 AND2X2_2794 ( .A(u2__abc_52155_new_n7734_), .B(u2__abc_52155_new_n7737_), .Y(u2__abc_52155_new_n7738_));
AND2X2 AND2X2_2795 ( .A(u2__abc_52155_new_n7739_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__6_));
AND2X2 AND2X2_2796 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_7_), .Y(u2__abc_52155_new_n7741_));
AND2X2 AND2X2_2797 ( .A(u2__abc_52155_new_n7729_), .B(u2__abc_52155_new_n7743_), .Y(u2__abc_52155_new_n7744_));
AND2X2 AND2X2_2798 ( .A(u2__abc_52155_new_n7746_), .B(u2__abc_52155_new_n7747_), .Y(u2__abc_52155_new_n7748_));
AND2X2 AND2X2_2799 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7748_), .Y(u2__abc_52155_new_n7749_));
AND2X2 AND2X2_28 ( .A(_abc_73687_new_n753_), .B(sqrto_27_), .Y(\o[63] ));
AND2X2 AND2X2_280 ( .A(_abc_73687_new_n1438_), .B(_abc_73687_new_n1437_), .Y(fracta1_90_));
AND2X2 AND2X2_2800 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_5_), .Y(u2__abc_52155_new_n7750_));
AND2X2 AND2X2_2801 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n7753_), .Y(u2__abc_52155_new_n7754_));
AND2X2 AND2X2_2802 ( .A(u2__abc_52155_new_n7755_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7756_));
AND2X2 AND2X2_2803 ( .A(u2__abc_52155_new_n7752_), .B(u2__abc_52155_new_n7756_), .Y(u2__abc_52155_new_n7757_));
AND2X2 AND2X2_2804 ( .A(u2__abc_52155_new_n7758_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__7_));
AND2X2 AND2X2_2805 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_8_), .Y(u2__abc_52155_new_n7760_));
AND2X2 AND2X2_2806 ( .A(u2__abc_52155_new_n7688_), .B(u2__abc_52155_new_n7590_), .Y(u2__abc_52155_new_n7761_));
AND2X2 AND2X2_2807 ( .A(u2__abc_52155_new_n7762_), .B(u2__abc_52155_new_n7725_), .Y(u2__abc_52155_new_n7763_));
AND2X2 AND2X2_2808 ( .A(u2__abc_52155_new_n3139_), .B(u2__abc_52155_new_n3092_), .Y(u2__abc_52155_new_n7764_));
AND2X2 AND2X2_2809 ( .A(u2__abc_52155_new_n7767_), .B(u2__abc_52155_new_n3086_), .Y(u2__abc_52155_new_n7768_));
AND2X2 AND2X2_281 ( .A(_abc_73687_new_n1441_), .B(_abc_73687_new_n1440_), .Y(fracta1_91_));
AND2X2 AND2X2_2810 ( .A(u2__abc_52155_new_n7769_), .B(u2__abc_52155_new_n7770_), .Y(u2__abc_52155_new_n7771_));
AND2X2 AND2X2_2811 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7771_), .Y(u2__abc_52155_new_n7772_));
AND2X2 AND2X2_2812 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_6_), .Y(u2__abc_52155_new_n7773_));
AND2X2 AND2X2_2813 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3065_), .Y(u2__abc_52155_new_n7776_));
AND2X2 AND2X2_2814 ( .A(u2__abc_52155_new_n7777_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7778_));
AND2X2 AND2X2_2815 ( .A(u2__abc_52155_new_n7775_), .B(u2__abc_52155_new_n7778_), .Y(u2__abc_52155_new_n7779_));
AND2X2 AND2X2_2816 ( .A(u2__abc_52155_new_n7780_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__8_));
AND2X2 AND2X2_2817 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_9_), .Y(u2__abc_52155_new_n7782_));
AND2X2 AND2X2_2818 ( .A(u2__abc_52155_new_n7769_), .B(u2__abc_52155_new_n3083_), .Y(u2__abc_52155_new_n7784_));
AND2X2 AND2X2_2819 ( .A(u2__abc_52155_new_n7785_), .B(u2__abc_52155_new_n7783_), .Y(u2__abc_52155_new_n7786_));
AND2X2 AND2X2_282 ( .A(_abc_73687_new_n1444_), .B(_abc_73687_new_n1443_), .Y(fracta1_92_));
AND2X2 AND2X2_2820 ( .A(u2__abc_52155_new_n7784_), .B(u2__abc_52155_new_n3081_), .Y(u2__abc_52155_new_n7787_));
AND2X2 AND2X2_2821 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7788_), .Y(u2__abc_52155_new_n7789_));
AND2X2 AND2X2_2822 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_7_), .Y(u2__abc_52155_new_n7790_));
AND2X2 AND2X2_2823 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3072_), .Y(u2__abc_52155_new_n7793_));
AND2X2 AND2X2_2824 ( .A(u2__abc_52155_new_n7794_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7795_));
AND2X2 AND2X2_2825 ( .A(u2__abc_52155_new_n7792_), .B(u2__abc_52155_new_n7795_), .Y(u2__abc_52155_new_n7796_));
AND2X2 AND2X2_2826 ( .A(u2__abc_52155_new_n7797_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__9_));
AND2X2 AND2X2_2827 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_10_), .Y(u2__abc_52155_new_n7799_));
AND2X2 AND2X2_2828 ( .A(u2__abc_52155_new_n3079_), .B(u2__abc_52155_new_n3083_), .Y(u2__abc_52155_new_n7800_));
AND2X2 AND2X2_2829 ( .A(u2__abc_52155_new_n7801_), .B(u2__abc_52155_new_n3080_), .Y(u2__abc_52155_new_n7802_));
AND2X2 AND2X2_283 ( .A(_abc_73687_new_n1447_), .B(_abc_73687_new_n1446_), .Y(fracta1_93_));
AND2X2 AND2X2_2830 ( .A(u2__abc_52155_new_n7767_), .B(u2__abc_52155_new_n3087_), .Y(u2__abc_52155_new_n7803_));
AND2X2 AND2X2_2831 ( .A(u2__abc_52155_new_n7804_), .B(u2__abc_52155_new_n3068_), .Y(u2__abc_52155_new_n7806_));
AND2X2 AND2X2_2832 ( .A(u2__abc_52155_new_n7807_), .B(u2__abc_52155_new_n7805_), .Y(u2__abc_52155_new_n7808_));
AND2X2 AND2X2_2833 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7808_), .Y(u2__abc_52155_new_n7809_));
AND2X2 AND2X2_2834 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_8_), .Y(u2__abc_52155_new_n7810_));
AND2X2 AND2X2_2835 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3057_), .Y(u2__abc_52155_new_n7813_));
AND2X2 AND2X2_2836 ( .A(u2__abc_52155_new_n7814_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7815_));
AND2X2 AND2X2_2837 ( .A(u2__abc_52155_new_n7812_), .B(u2__abc_52155_new_n7815_), .Y(u2__abc_52155_new_n7816_));
AND2X2 AND2X2_2838 ( .A(u2__abc_52155_new_n7817_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__10_));
AND2X2 AND2X2_2839 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_11_), .Y(u2__abc_52155_new_n7819_));
AND2X2 AND2X2_284 ( .A(_abc_73687_new_n1450_), .B(_abc_73687_new_n1449_), .Y(fracta1_94_));
AND2X2 AND2X2_2840 ( .A(u2__abc_52155_new_n7807_), .B(u2__abc_52155_new_n7821_), .Y(u2__abc_52155_new_n7822_));
AND2X2 AND2X2_2841 ( .A(u2__abc_52155_new_n7823_), .B(u2__abc_52155_new_n7820_), .Y(u2__abc_52155_new_n7824_));
AND2X2 AND2X2_2842 ( .A(u2__abc_52155_new_n7822_), .B(u2__abc_52155_new_n3075_), .Y(u2__abc_52155_new_n7825_));
AND2X2 AND2X2_2843 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7826_), .Y(u2__abc_52155_new_n7827_));
AND2X2 AND2X2_2844 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_9_), .Y(u2__abc_52155_new_n7828_));
AND2X2 AND2X2_2845 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3051_), .Y(u2__abc_52155_new_n7831_));
AND2X2 AND2X2_2846 ( .A(u2__abc_52155_new_n7832_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7833_));
AND2X2 AND2X2_2847 ( .A(u2__abc_52155_new_n7830_), .B(u2__abc_52155_new_n7833_), .Y(u2__abc_52155_new_n7834_));
AND2X2 AND2X2_2848 ( .A(u2__abc_52155_new_n7835_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__11_));
AND2X2 AND2X2_2849 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_12_), .Y(u2__abc_52155_new_n7837_));
AND2X2 AND2X2_285 ( .A(_abc_73687_new_n1453_), .B(_abc_73687_new_n1452_), .Y(fracta1_95_));
AND2X2 AND2X2_2850 ( .A(u2__abc_52155_new_n7821_), .B(u2__abc_52155_new_n3071_), .Y(u2__abc_52155_new_n7838_));
AND2X2 AND2X2_2851 ( .A(u2__abc_52155_new_n7807_), .B(u2__abc_52155_new_n7838_), .Y(u2__abc_52155_new_n7839_));
AND2X2 AND2X2_2852 ( .A(u2__abc_52155_new_n7841_), .B(u2__abc_52155_new_n3060_), .Y(u2__abc_52155_new_n7843_));
AND2X2 AND2X2_2853 ( .A(u2__abc_52155_new_n7844_), .B(u2__abc_52155_new_n7842_), .Y(u2__abc_52155_new_n7845_));
AND2X2 AND2X2_2854 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7845_), .Y(u2__abc_52155_new_n7846_));
AND2X2 AND2X2_2855 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_10_), .Y(u2__abc_52155_new_n7847_));
AND2X2 AND2X2_2856 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3037_), .Y(u2__abc_52155_new_n7850_));
AND2X2 AND2X2_2857 ( .A(u2__abc_52155_new_n7851_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7852_));
AND2X2 AND2X2_2858 ( .A(u2__abc_52155_new_n7849_), .B(u2__abc_52155_new_n7852_), .Y(u2__abc_52155_new_n7853_));
AND2X2 AND2X2_2859 ( .A(u2__abc_52155_new_n7854_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__12_));
AND2X2 AND2X2_286 ( .A(_abc_73687_new_n1456_), .B(_abc_73687_new_n1455_), .Y(fracta1_96_));
AND2X2 AND2X2_2860 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_13_), .Y(u2__abc_52155_new_n7856_));
AND2X2 AND2X2_2861 ( .A(u2__abc_52155_new_n7844_), .B(u2__abc_52155_new_n7857_), .Y(u2__abc_52155_new_n7858_));
AND2X2 AND2X2_2862 ( .A(u2__abc_52155_new_n7858_), .B(u2__abc_52155_new_n3054_), .Y(u2__abc_52155_new_n7859_));
AND2X2 AND2X2_2863 ( .A(u2__abc_52155_new_n7861_), .B(u2__abc_52155_new_n7860_), .Y(u2__abc_52155_new_n7862_));
AND2X2 AND2X2_2864 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7863_), .Y(u2__abc_52155_new_n7864_));
AND2X2 AND2X2_2865 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_11_), .Y(u2__abc_52155_new_n7865_));
AND2X2 AND2X2_2866 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3041_), .Y(u2__abc_52155_new_n7868_));
AND2X2 AND2X2_2867 ( .A(u2__abc_52155_new_n7869_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7870_));
AND2X2 AND2X2_2868 ( .A(u2__abc_52155_new_n7867_), .B(u2__abc_52155_new_n7870_), .Y(u2__abc_52155_new_n7871_));
AND2X2 AND2X2_2869 ( .A(u2__abc_52155_new_n7872_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__13_));
AND2X2 AND2X2_287 ( .A(_abc_73687_new_n1459_), .B(_abc_73687_new_n1458_), .Y(fracta1_97_));
AND2X2 AND2X2_2870 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_14_), .Y(u2__abc_52155_new_n7874_));
AND2X2 AND2X2_2871 ( .A(u2__abc_52155_new_n3054_), .B(u2__abc_52155_new_n3056_), .Y(u2__abc_52155_new_n7877_));
AND2X2 AND2X2_2872 ( .A(u2__abc_52155_new_n7876_), .B(u2__abc_52155_new_n7879_), .Y(u2__abc_52155_new_n7880_));
AND2X2 AND2X2_2873 ( .A(u2__abc_52155_new_n7881_), .B(u2__abc_52155_new_n3040_), .Y(u2__abc_52155_new_n7883_));
AND2X2 AND2X2_2874 ( .A(u2__abc_52155_new_n7884_), .B(u2__abc_52155_new_n7882_), .Y(u2__abc_52155_new_n7885_));
AND2X2 AND2X2_2875 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7885_), .Y(u2__abc_52155_new_n7886_));
AND2X2 AND2X2_2876 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_12_), .Y(u2__abc_52155_new_n7887_));
AND2X2 AND2X2_2877 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n7890_), .Y(u2__abc_52155_new_n7891_));
AND2X2 AND2X2_2878 ( .A(u2__abc_52155_new_n7892_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7893_));
AND2X2 AND2X2_2879 ( .A(u2__abc_52155_new_n7889_), .B(u2__abc_52155_new_n7893_), .Y(u2__abc_52155_new_n7894_));
AND2X2 AND2X2_288 ( .A(_abc_73687_new_n1462_), .B(_abc_73687_new_n1461_), .Y(fracta1_98_));
AND2X2 AND2X2_2880 ( .A(u2__abc_52155_new_n7895_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__14_));
AND2X2 AND2X2_2881 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_15_), .Y(u2__abc_52155_new_n7897_));
AND2X2 AND2X2_2882 ( .A(u2__abc_52155_new_n7884_), .B(u2__abc_52155_new_n7898_), .Y(u2__abc_52155_new_n7899_));
AND2X2 AND2X2_2883 ( .A(u2__abc_52155_new_n7901_), .B(u2__abc_52155_new_n7902_), .Y(u2__abc_52155_new_n7903_));
AND2X2 AND2X2_2884 ( .A(u2__abc_52155_new_n7904_), .B(u2__abc_52155_new_n7905_), .Y(u2__abc_52155_new_n7906_));
AND2X2 AND2X2_2885 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3247_), .Y(u2__abc_52155_new_n7908_));
AND2X2 AND2X2_2886 ( .A(u2__abc_52155_new_n7909_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7910_));
AND2X2 AND2X2_2887 ( .A(u2__abc_52155_new_n7907_), .B(u2__abc_52155_new_n7910_), .Y(u2__abc_52155_new_n7911_));
AND2X2 AND2X2_2888 ( .A(u2__abc_52155_new_n7912_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__15_));
AND2X2 AND2X2_2889 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_16_), .Y(u2__abc_52155_new_n7914_));
AND2X2 AND2X2_289 ( .A(_abc_73687_new_n1465_), .B(_abc_73687_new_n1464_), .Y(fracta1_99_));
AND2X2 AND2X2_2890 ( .A(u2__abc_52155_new_n7767_), .B(u2__abc_52155_new_n3089_), .Y(u2__abc_52155_new_n7915_));
AND2X2 AND2X2_2891 ( .A(u2__abc_52155_new_n7802_), .B(u2__abc_52155_new_n3076_), .Y(u2__abc_52155_new_n7918_));
AND2X2 AND2X2_2892 ( .A(u2__abc_52155_new_n7919_), .B(u2__abc_52155_new_n7917_), .Y(u2__abc_52155_new_n7920_));
AND2X2 AND2X2_2893 ( .A(u2__abc_52155_new_n7878_), .B(u2__abc_52155_new_n3047_), .Y(u2__abc_52155_new_n7922_));
AND2X2 AND2X2_2894 ( .A(u2__abc_52155_new_n3046_), .B(u2__abc_52155_new_n3036_), .Y(u2__abc_52155_new_n7923_));
AND2X2 AND2X2_2895 ( .A(u2__abc_52155_new_n7921_), .B(u2__abc_52155_new_n7926_), .Y(u2__abc_52155_new_n7927_));
AND2X2 AND2X2_2896 ( .A(u2__abc_52155_new_n7916_), .B(u2__abc_52155_new_n7927_), .Y(u2__abc_52155_new_n7928_));
AND2X2 AND2X2_2897 ( .A(u2__abc_52155_new_n7929_), .B(u2__abc_52155_new_n3243_), .Y(u2__abc_52155_new_n7931_));
AND2X2 AND2X2_2898 ( .A(u2__abc_52155_new_n7932_), .B(u2__abc_52155_new_n7930_), .Y(u2__abc_52155_new_n7933_));
AND2X2 AND2X2_2899 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7933_), .Y(u2__abc_52155_new_n7934_));
AND2X2 AND2X2_29 ( .A(_abc_73687_new_n753_), .B(sqrto_28_), .Y(\o[64] ));
AND2X2 AND2X2_290 ( .A(_abc_73687_new_n1468_), .B(_abc_73687_new_n1467_), .Y(fracta1_100_));
AND2X2 AND2X2_2900 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_14_), .Y(u2__abc_52155_new_n7935_));
AND2X2 AND2X2_2901 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3229_), .Y(u2__abc_52155_new_n7938_));
AND2X2 AND2X2_2902 ( .A(u2__abc_52155_new_n7939_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7940_));
AND2X2 AND2X2_2903 ( .A(u2__abc_52155_new_n7937_), .B(u2__abc_52155_new_n7940_), .Y(u2__abc_52155_new_n7941_));
AND2X2 AND2X2_2904 ( .A(u2__abc_52155_new_n7942_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__16_));
AND2X2 AND2X2_2905 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_17_), .Y(u2__abc_52155_new_n7944_));
AND2X2 AND2X2_2906 ( .A(u2__abc_52155_new_n7932_), .B(u2__abc_52155_new_n3241_), .Y(u2__abc_52155_new_n7946_));
AND2X2 AND2X2_2907 ( .A(u2__abc_52155_new_n7947_), .B(u2__abc_52155_new_n7945_), .Y(u2__abc_52155_new_n7948_));
AND2X2 AND2X2_2908 ( .A(u2__abc_52155_new_n7946_), .B(u2__abc_52155_new_n3250_), .Y(u2__abc_52155_new_n7949_));
AND2X2 AND2X2_2909 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7950_), .Y(u2__abc_52155_new_n7951_));
AND2X2 AND2X2_291 ( .A(_abc_73687_new_n1471_), .B(_abc_73687_new_n1470_), .Y(fracta1_101_));
AND2X2 AND2X2_2910 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_15_), .Y(u2__abc_52155_new_n7952_));
AND2X2 AND2X2_2911 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3234_), .Y(u2__abc_52155_new_n7955_));
AND2X2 AND2X2_2912 ( .A(u2__abc_52155_new_n7956_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7957_));
AND2X2 AND2X2_2913 ( .A(u2__abc_52155_new_n7954_), .B(u2__abc_52155_new_n7957_), .Y(u2__abc_52155_new_n7958_));
AND2X2 AND2X2_2914 ( .A(u2__abc_52155_new_n7959_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__17_));
AND2X2 AND2X2_2915 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_18_), .Y(u2__abc_52155_new_n7961_));
AND2X2 AND2X2_2916 ( .A(u2__abc_52155_new_n7947_), .B(u2__abc_52155_new_n3249_), .Y(u2__abc_52155_new_n7963_));
AND2X2 AND2X2_2917 ( .A(u2__abc_52155_new_n7964_), .B(u2__abc_52155_new_n7962_), .Y(u2__abc_52155_new_n7966_));
AND2X2 AND2X2_2918 ( .A(u2__abc_52155_new_n7967_), .B(u2__abc_52155_new_n7965_), .Y(u2__abc_52155_new_n7968_));
AND2X2 AND2X2_2919 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7968_), .Y(u2__abc_52155_new_n7969_));
AND2X2 AND2X2_292 ( .A(_abc_73687_new_n1474_), .B(_abc_73687_new_n1473_), .Y(fracta1_102_));
AND2X2 AND2X2_2920 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_16_), .Y(u2__abc_52155_new_n7970_));
AND2X2 AND2X2_2921 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3271_), .Y(u2__abc_52155_new_n7973_));
AND2X2 AND2X2_2922 ( .A(u2__abc_52155_new_n7974_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7975_));
AND2X2 AND2X2_2923 ( .A(u2__abc_52155_new_n7972_), .B(u2__abc_52155_new_n7975_), .Y(u2__abc_52155_new_n7976_));
AND2X2 AND2X2_2924 ( .A(u2__abc_52155_new_n7977_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__18_));
AND2X2 AND2X2_2925 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_19_), .Y(u2__abc_52155_new_n7979_));
AND2X2 AND2X2_2926 ( .A(u2__abc_52155_new_n7967_), .B(u2__abc_52155_new_n7980_), .Y(u2__abc_52155_new_n7981_));
AND2X2 AND2X2_2927 ( .A(u2__abc_52155_new_n7982_), .B(u2__abc_52155_new_n3236_), .Y(u2__abc_52155_new_n7983_));
AND2X2 AND2X2_2928 ( .A(u2__abc_52155_new_n7981_), .B(u2__abc_52155_new_n7984_), .Y(u2__abc_52155_new_n7985_));
AND2X2 AND2X2_2929 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n7986_), .Y(u2__abc_52155_new_n7987_));
AND2X2 AND2X2_293 ( .A(_abc_73687_new_n1477_), .B(_abc_73687_new_n1476_), .Y(fracta1_103_));
AND2X2 AND2X2_2930 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_17_), .Y(u2__abc_52155_new_n7988_));
AND2X2 AND2X2_2931 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3266_), .Y(u2__abc_52155_new_n7991_));
AND2X2 AND2X2_2932 ( .A(u2__abc_52155_new_n7992_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n7993_));
AND2X2 AND2X2_2933 ( .A(u2__abc_52155_new_n7990_), .B(u2__abc_52155_new_n7993_), .Y(u2__abc_52155_new_n7994_));
AND2X2 AND2X2_2934 ( .A(u2__abc_52155_new_n7995_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__19_));
AND2X2 AND2X2_2935 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_20_), .Y(u2__abc_52155_new_n7997_));
AND2X2 AND2X2_2936 ( .A(u2__abc_52155_new_n3241_), .B(u2__abc_52155_new_n3246_), .Y(u2__abc_52155_new_n7999_));
AND2X2 AND2X2_2937 ( .A(u2__abc_52155_new_n3285_), .B(u2__abc_52155_new_n3228_), .Y(u2__abc_52155_new_n8002_));
AND2X2 AND2X2_2938 ( .A(u2__abc_52155_new_n8001_), .B(u2__abc_52155_new_n8004_), .Y(u2__abc_52155_new_n8005_));
AND2X2 AND2X2_2939 ( .A(u2__abc_52155_new_n7929_), .B(u2__abc_52155_new_n3252_), .Y(u2__abc_52155_new_n8007_));
AND2X2 AND2X2_294 ( .A(_abc_73687_new_n1480_), .B(_abc_73687_new_n1479_), .Y(fracta1_104_));
AND2X2 AND2X2_2940 ( .A(u2__abc_52155_new_n8008_), .B(u2__abc_52155_new_n7998_), .Y(u2__abc_52155_new_n8010_));
AND2X2 AND2X2_2941 ( .A(u2__abc_52155_new_n8011_), .B(u2__abc_52155_new_n8009_), .Y(u2__abc_52155_new_n8012_));
AND2X2 AND2X2_2942 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n8012_), .Y(u2__abc_52155_new_n8013_));
AND2X2 AND2X2_2943 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_18_), .Y(u2__abc_52155_new_n8014_));
AND2X2 AND2X2_2944 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3255_), .Y(u2__abc_52155_new_n8017_));
AND2X2 AND2X2_2945 ( .A(u2__abc_52155_new_n8018_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8019_));
AND2X2 AND2X2_2946 ( .A(u2__abc_52155_new_n8016_), .B(u2__abc_52155_new_n8019_), .Y(u2__abc_52155_new_n8020_));
AND2X2 AND2X2_2947 ( .A(u2__abc_52155_new_n8021_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__20_));
AND2X2 AND2X2_2948 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_21_), .Y(u2__abc_52155_new_n8023_));
AND2X2 AND2X2_2949 ( .A(u2__abc_52155_new_n8011_), .B(u2__abc_52155_new_n8025_), .Y(u2__abc_52155_new_n8026_));
AND2X2 AND2X2_295 ( .A(_abc_73687_new_n1483_), .B(_abc_73687_new_n1482_), .Y(fracta1_105_));
AND2X2 AND2X2_2950 ( .A(u2__abc_52155_new_n8028_), .B(u2__abc_52155_new_n8029_), .Y(u2__abc_52155_new_n8030_));
AND2X2 AND2X2_2951 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n8030_), .Y(u2__abc_52155_new_n8031_));
AND2X2 AND2X2_2952 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_19_), .Y(u2__abc_52155_new_n8032_));
AND2X2 AND2X2_2953 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3260_), .Y(u2__abc_52155_new_n8035_));
AND2X2 AND2X2_2954 ( .A(u2__abc_52155_new_n8036_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8037_));
AND2X2 AND2X2_2955 ( .A(u2__abc_52155_new_n8034_), .B(u2__abc_52155_new_n8037_), .Y(u2__abc_52155_new_n8038_));
AND2X2 AND2X2_2956 ( .A(u2__abc_52155_new_n8039_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__21_));
AND2X2 AND2X2_2957 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_22_), .Y(u2__abc_52155_new_n8041_));
AND2X2 AND2X2_2958 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_20_), .Y(u2__abc_52155_new_n8042_));
AND2X2 AND2X2_2959 ( .A(u2__abc_52155_new_n8011_), .B(u2__abc_52155_new_n8045_), .Y(u2__abc_52155_new_n8046_));
AND2X2 AND2X2_296 ( .A(_abc_73687_new_n1486_), .B(_abc_73687_new_n1485_), .Y(fracta1_106_));
AND2X2 AND2X2_2960 ( .A(u2__abc_52155_new_n8048_), .B(u2__abc_52155_new_n8043_), .Y(u2__abc_52155_new_n8050_));
AND2X2 AND2X2_2961 ( .A(u2__abc_52155_new_n8051_), .B(u2__abc_52155_new_n8049_), .Y(u2__abc_52155_new_n8052_));
AND2X2 AND2X2_2962 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n8052_), .Y(u2__abc_52155_new_n8053_));
AND2X2 AND2X2_2963 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3189_), .Y(u2__abc_52155_new_n8056_));
AND2X2 AND2X2_2964 ( .A(u2__abc_52155_new_n8057_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8058_));
AND2X2 AND2X2_2965 ( .A(u2__abc_52155_new_n8055_), .B(u2__abc_52155_new_n8058_), .Y(u2__abc_52155_new_n8059_));
AND2X2 AND2X2_2966 ( .A(u2__abc_52155_new_n8060_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__22_));
AND2X2 AND2X2_2967 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_23_), .Y(u2__abc_52155_new_n8062_));
AND2X2 AND2X2_2968 ( .A(u2__abc_52155_new_n8051_), .B(u2__abc_52155_new_n8064_), .Y(u2__abc_52155_new_n8065_));
AND2X2 AND2X2_2969 ( .A(u2__abc_52155_new_n8066_), .B(u2__abc_52155_new_n3262_), .Y(u2__abc_52155_new_n8067_));
AND2X2 AND2X2_297 ( .A(_abc_73687_new_n1489_), .B(_abc_73687_new_n1488_), .Y(fracta1_107_));
AND2X2 AND2X2_2970 ( .A(u2__abc_52155_new_n8065_), .B(u2__abc_52155_new_n8068_), .Y(u2__abc_52155_new_n8069_));
AND2X2 AND2X2_2971 ( .A(u2__abc_52155_new_n8071_), .B(u2__abc_52155_new_n8063_), .Y(u2__abc_52155_new_n8072_));
AND2X2 AND2X2_2972 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3182_), .Y(u2__abc_52155_new_n8074_));
AND2X2 AND2X2_2973 ( .A(u2__abc_52155_new_n8075_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8076_));
AND2X2 AND2X2_2974 ( .A(u2__abc_52155_new_n8073_), .B(u2__abc_52155_new_n8076_), .Y(u2__abc_52155_new_n8077_));
AND2X2 AND2X2_2975 ( .A(u2__abc_52155_new_n8078_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__23_));
AND2X2 AND2X2_2976 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_24_), .Y(u2__abc_52155_new_n8080_));
AND2X2 AND2X2_2977 ( .A(u2__abc_52155_new_n7929_), .B(u2__abc_52155_new_n3277_), .Y(u2__abc_52155_new_n8081_));
AND2X2 AND2X2_2978 ( .A(u2__abc_52155_new_n8006_), .B(u2__abc_52155_new_n3276_), .Y(u2__abc_52155_new_n8083_));
AND2X2 AND2X2_2979 ( .A(u2__abc_52155_new_n8087_), .B(u2__abc_52155_new_n3296_), .Y(u2__abc_52155_new_n8088_));
AND2X2 AND2X2_298 ( .A(_abc_73687_new_n1492_), .B(_abc_73687_new_n1491_), .Y(fracta1_108_));
AND2X2 AND2X2_2980 ( .A(u2__abc_52155_new_n8086_), .B(u2__abc_52155_new_n8088_), .Y(u2__abc_52155_new_n8089_));
AND2X2 AND2X2_2981 ( .A(u2__abc_52155_new_n8084_), .B(u2__abc_52155_new_n8089_), .Y(u2__abc_52155_new_n8090_));
AND2X2 AND2X2_2982 ( .A(u2__abc_52155_new_n8082_), .B(u2__abc_52155_new_n8090_), .Y(u2__abc_52155_new_n8091_));
AND2X2 AND2X2_2983 ( .A(u2__abc_52155_new_n8092_), .B(u2__abc_52155_new_n3192_), .Y(u2__abc_52155_new_n8094_));
AND2X2 AND2X2_2984 ( .A(u2__abc_52155_new_n8095_), .B(u2__abc_52155_new_n8093_), .Y(u2__abc_52155_new_n8096_));
AND2X2 AND2X2_2985 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n8096_), .Y(u2__abc_52155_new_n8097_));
AND2X2 AND2X2_2986 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_22_), .Y(u2__abc_52155_new_n8098_));
AND2X2 AND2X2_2987 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3169_), .Y(u2__abc_52155_new_n8101_));
AND2X2 AND2X2_2988 ( .A(u2__abc_52155_new_n8102_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8103_));
AND2X2 AND2X2_2989 ( .A(u2__abc_52155_new_n8100_), .B(u2__abc_52155_new_n8103_), .Y(u2__abc_52155_new_n8104_));
AND2X2 AND2X2_299 ( .A(_abc_73687_new_n1495_), .B(_abc_73687_new_n1494_), .Y(fracta1_109_));
AND2X2 AND2X2_2990 ( .A(u2__abc_52155_new_n8105_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__24_));
AND2X2 AND2X2_2991 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_25_), .Y(u2__abc_52155_new_n8107_));
AND2X2 AND2X2_2992 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_23_), .Y(u2__abc_52155_new_n8108_));
AND2X2 AND2X2_2993 ( .A(u2__abc_52155_new_n8095_), .B(u2__abc_52155_new_n3188_), .Y(u2__abc_52155_new_n8109_));
AND2X2 AND2X2_2994 ( .A(u2__abc_52155_new_n8111_), .B(u2__abc_52155_new_n8113_), .Y(u2__abc_52155_new_n8114_));
AND2X2 AND2X2_2995 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n8114_), .Y(u2__abc_52155_new_n8115_));
AND2X2 AND2X2_2996 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3174_), .Y(u2__abc_52155_new_n8118_));
AND2X2 AND2X2_2997 ( .A(u2__abc_52155_new_n8119_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8120_));
AND2X2 AND2X2_2998 ( .A(u2__abc_52155_new_n8117_), .B(u2__abc_52155_new_n8120_), .Y(u2__abc_52155_new_n8121_));
AND2X2 AND2X2_2999 ( .A(u2__abc_52155_new_n8122_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__25_));
AND2X2 AND2X2_3 ( .A(_abc_73687_new_n753_), .B(sqrto_2_), .Y(\o[38] ));
AND2X2 AND2X2_30 ( .A(_abc_73687_new_n753_), .B(sqrto_29_), .Y(\o[65] ));
AND2X2 AND2X2_300 ( .A(_abc_73687_new_n1498_), .B(_abc_73687_new_n1497_), .Y(fracta1_110_));
AND2X2 AND2X2_3000 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_26_), .Y(u2__abc_52155_new_n8124_));
AND2X2 AND2X2_3001 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_24_), .Y(u2__abc_52155_new_n8125_));
AND2X2 AND2X2_3002 ( .A(u2__abc_52155_new_n3181_), .B(u2__abc_52155_new_n3188_), .Y(u2__abc_52155_new_n8127_));
AND2X2 AND2X2_3003 ( .A(u2__abc_52155_new_n8095_), .B(u2__abc_52155_new_n8127_), .Y(u2__abc_52155_new_n8128_));
AND2X2 AND2X2_3004 ( .A(u2__abc_52155_new_n8130_), .B(u2__abc_52155_new_n8126_), .Y(u2__abc_52155_new_n8132_));
AND2X2 AND2X2_3005 ( .A(u2__abc_52155_new_n8133_), .B(u2__abc_52155_new_n8131_), .Y(u2__abc_52155_new_n8134_));
AND2X2 AND2X2_3006 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n8134_), .Y(u2__abc_52155_new_n8135_));
AND2X2 AND2X2_3007 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3220_), .Y(u2__abc_52155_new_n8138_));
AND2X2 AND2X2_3008 ( .A(u2__abc_52155_new_n8139_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8140_));
AND2X2 AND2X2_3009 ( .A(u2__abc_52155_new_n8137_), .B(u2__abc_52155_new_n8140_), .Y(u2__abc_52155_new_n8141_));
AND2X2 AND2X2_301 ( .A(_abc_73687_new_n1501_), .B(_abc_73687_new_n1500_), .Y(fracta1_111_));
AND2X2 AND2X2_3010 ( .A(u2__abc_52155_new_n8142_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__26_));
AND2X2 AND2X2_3011 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_27_), .Y(u2__abc_52155_new_n8144_));
AND2X2 AND2X2_3012 ( .A(u2__abc_52155_new_n8133_), .B(u2__abc_52155_new_n8145_), .Y(u2__abc_52155_new_n8146_));
AND2X2 AND2X2_3013 ( .A(u2__abc_52155_new_n8147_), .B(u2__abc_52155_new_n3176_), .Y(u2__abc_52155_new_n8148_));
AND2X2 AND2X2_3014 ( .A(u2__abc_52155_new_n8146_), .B(u2__abc_52155_new_n8149_), .Y(u2__abc_52155_new_n8150_));
AND2X2 AND2X2_3015 ( .A(u2__abc_52155_new_n8151_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8152_));
AND2X2 AND2X2_3016 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_25_), .Y(u2__abc_52155_new_n8153_));
AND2X2 AND2X2_3017 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3213_), .Y(u2__abc_52155_new_n8156_));
AND2X2 AND2X2_3018 ( .A(u2__abc_52155_new_n8157_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8158_));
AND2X2 AND2X2_3019 ( .A(u2__abc_52155_new_n8155_), .B(u2__abc_52155_new_n8158_), .Y(u2__abc_52155_new_n8159_));
AND2X2 AND2X2_302 ( .A(_abc_73687_new_n1504_), .B(_abc_73687_new_n1503_), .Y(fracta1_112_));
AND2X2 AND2X2_3020 ( .A(u2__abc_52155_new_n8160_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__27_));
AND2X2 AND2X2_3021 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_28_), .Y(u2__abc_52155_new_n8162_));
AND2X2 AND2X2_3022 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_26_), .Y(u2__abc_52155_new_n8163_));
AND2X2 AND2X2_3023 ( .A(u2__abc_52155_new_n8092_), .B(u2__abc_52155_new_n3194_), .Y(u2__abc_52155_new_n8164_));
AND2X2 AND2X2_3024 ( .A(u2__abc_52155_new_n8168_), .B(u2__abc_52155_new_n3307_), .Y(u2__abc_52155_new_n8169_));
AND2X2 AND2X2_3025 ( .A(u2__abc_52155_new_n8167_), .B(u2__abc_52155_new_n8169_), .Y(u2__abc_52155_new_n8170_));
AND2X2 AND2X2_3026 ( .A(u2__abc_52155_new_n8165_), .B(u2__abc_52155_new_n8170_), .Y(u2__abc_52155_new_n8171_));
AND2X2 AND2X2_3027 ( .A(u2__abc_52155_new_n8172_), .B(u2__abc_52155_new_n3223_), .Y(u2__abc_52155_new_n8174_));
AND2X2 AND2X2_3028 ( .A(u2__abc_52155_new_n8175_), .B(u2__abc_52155_new_n8173_), .Y(u2__abc_52155_new_n8176_));
AND2X2 AND2X2_3029 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n8176_), .Y(u2__abc_52155_new_n8177_));
AND2X2 AND2X2_303 ( .A(_abc_73687_new_n1170_), .B(fracta_112_), .Y(fracta1_113_));
AND2X2 AND2X2_3030 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3198_), .Y(u2__abc_52155_new_n8180_));
AND2X2 AND2X2_3031 ( .A(u2__abc_52155_new_n8181_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8182_));
AND2X2 AND2X2_3032 ( .A(u2__abc_52155_new_n8179_), .B(u2__abc_52155_new_n8182_), .Y(u2__abc_52155_new_n8183_));
AND2X2 AND2X2_3033 ( .A(u2__abc_52155_new_n8184_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__28_));
AND2X2 AND2X2_3034 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_29_), .Y(u2__abc_52155_new_n8186_));
AND2X2 AND2X2_3035 ( .A(u2__abc_52155_new_n8175_), .B(u2__abc_52155_new_n3219_), .Y(u2__abc_52155_new_n8189_));
AND2X2 AND2X2_3036 ( .A(u2__abc_52155_new_n8190_), .B(u2__abc_52155_new_n8188_), .Y(u2__abc_52155_new_n8191_));
AND2X2 AND2X2_3037 ( .A(u2__abc_52155_new_n8189_), .B(u2__abc_52155_new_n3216_), .Y(u2__abc_52155_new_n8192_));
AND2X2 AND2X2_3038 ( .A(u2__abc_52155_new_n8194_), .B(u2__abc_52155_new_n8187_), .Y(u2__abc_52155_new_n8195_));
AND2X2 AND2X2_3039 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3202_), .Y(u2__abc_52155_new_n8197_));
AND2X2 AND2X2_304 ( .A(\a[112] ), .B(\a[113] ), .Y(_abc_73687_new_n1507_));
AND2X2 AND2X2_3040 ( .A(u2__abc_52155_new_n8198_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8199_));
AND2X2 AND2X2_3041 ( .A(u2__abc_52155_new_n8196_), .B(u2__abc_52155_new_n8199_), .Y(u2__abc_52155_new_n8200_));
AND2X2 AND2X2_3042 ( .A(u2__abc_52155_new_n8201_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__29_));
AND2X2 AND2X2_3043 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_30_), .Y(u2__abc_52155_new_n8203_));
AND2X2 AND2X2_3044 ( .A(u2__abc_52155_new_n3212_), .B(u2__abc_52155_new_n3219_), .Y(u2__abc_52155_new_n8204_));
AND2X2 AND2X2_3045 ( .A(u2__abc_52155_new_n8175_), .B(u2__abc_52155_new_n8204_), .Y(u2__abc_52155_new_n8205_));
AND2X2 AND2X2_3046 ( .A(u2__abc_52155_new_n8207_), .B(u2__abc_52155_new_n3201_), .Y(u2__abc_52155_new_n8209_));
AND2X2 AND2X2_3047 ( .A(u2__abc_52155_new_n8210_), .B(u2__abc_52155_new_n8208_), .Y(u2__abc_52155_new_n8211_));
AND2X2 AND2X2_3048 ( .A(u2__abc_52155_new_n8212_), .B(u2__abc_52155_new_n8213_), .Y(u2__abc_52155_new_n8214_));
AND2X2 AND2X2_3049 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n8216_), .Y(u2__abc_52155_new_n8217_));
AND2X2 AND2X2_305 ( .A(_abc_73687_new_n1170_), .B(_abc_73687_new_n1508_), .Y(_abc_73687_new_n1509_));
AND2X2 AND2X2_3050 ( .A(u2__abc_52155_new_n8218_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8219_));
AND2X2 AND2X2_3051 ( .A(u2__abc_52155_new_n8215_), .B(u2__abc_52155_new_n8219_), .Y(u2__abc_52155_new_n8220_));
AND2X2 AND2X2_3052 ( .A(u2__abc_52155_new_n8221_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__30_));
AND2X2 AND2X2_3053 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_31_), .Y(u2__abc_52155_new_n8223_));
AND2X2 AND2X2_3054 ( .A(u2__abc_52155_new_n8210_), .B(u2__abc_52155_new_n3197_), .Y(u2__abc_52155_new_n8224_));
AND2X2 AND2X2_3055 ( .A(u2__abc_52155_new_n8226_), .B(u2__abc_52155_new_n8228_), .Y(u2__abc_52155_new_n8229_));
AND2X2 AND2X2_3056 ( .A(u2__abc_52155_new_n8229_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8230_));
AND2X2 AND2X2_3057 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_29_), .Y(u2__abc_52155_new_n8231_));
AND2X2 AND2X2_3058 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3527_), .Y(u2__abc_52155_new_n8234_));
AND2X2 AND2X2_3059 ( .A(u2__abc_52155_new_n8235_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8236_));
AND2X2 AND2X2_306 ( .A(_abc_73687_new_n1510_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1511_));
AND2X2 AND2X2_3060 ( .A(u2__abc_52155_new_n8233_), .B(u2__abc_52155_new_n8236_), .Y(u2__abc_52155_new_n8237_));
AND2X2 AND2X2_3061 ( .A(u2__abc_52155_new_n8238_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__31_));
AND2X2 AND2X2_3062 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_32_), .Y(u2__abc_52155_new_n8240_));
AND2X2 AND2X2_3063 ( .A(u2__abc_52155_new_n8242_), .B(u2__abc_52155_new_n3209_), .Y(u2__abc_52155_new_n8243_));
AND2X2 AND2X2_3064 ( .A(u2__abc_52155_new_n3204_), .B(u2__abc_52155_new_n3196_), .Y(u2__abc_52155_new_n8244_));
AND2X2 AND2X2_3065 ( .A(u2__abc_52155_new_n8172_), .B(u2__abc_52155_new_n3225_), .Y(u2__abc_52155_new_n8247_));
AND2X2 AND2X2_3066 ( .A(u2__abc_52155_new_n8248_), .B(u2__abc_52155_new_n3523_), .Y(u2__abc_52155_new_n8249_));
AND2X2 AND2X2_3067 ( .A(u2__abc_52155_new_n8250_), .B(u2__abc_52155_new_n8251_), .Y(u2__abc_52155_new_n8252_));
AND2X2 AND2X2_3068 ( .A(u2__abc_52155_new_n7622_), .B(u2__abc_52155_new_n8252_), .Y(u2__abc_52155_new_n8253_));
AND2X2 AND2X2_3069 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_30_), .Y(u2__abc_52155_new_n8254_));
AND2X2 AND2X2_307 ( .A(aNan), .B(\a[112] ), .Y(_abc_73687_new_n1512_));
AND2X2 AND2X2_3070 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3509_), .Y(u2__abc_52155_new_n8257_));
AND2X2 AND2X2_3071 ( .A(u2__abc_52155_new_n8258_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8259_));
AND2X2 AND2X2_3072 ( .A(u2__abc_52155_new_n8256_), .B(u2__abc_52155_new_n8259_), .Y(u2__abc_52155_new_n8260_));
AND2X2 AND2X2_3073 ( .A(u2__abc_52155_new_n8261_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__32_));
AND2X2 AND2X2_3074 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_33_), .Y(u2__abc_52155_new_n8263_));
AND2X2 AND2X2_3075 ( .A(u2__abc_52155_new_n8250_), .B(u2__abc_52155_new_n3521_), .Y(u2__abc_52155_new_n8265_));
AND2X2 AND2X2_3076 ( .A(u2__abc_52155_new_n8268_), .B(u2__abc_52155_new_n8266_), .Y(u2__abc_52155_new_n8269_));
AND2X2 AND2X2_3077 ( .A(u2__abc_52155_new_n8269_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8270_));
AND2X2 AND2X2_3078 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_31_), .Y(u2__abc_52155_new_n8271_));
AND2X2 AND2X2_3079 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3514_), .Y(u2__abc_52155_new_n8274_));
AND2X2 AND2X2_308 ( .A(_abc_73687_new_n1517_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1518_));
AND2X2 AND2X2_3080 ( .A(u2__abc_52155_new_n8275_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8276_));
AND2X2 AND2X2_3081 ( .A(u2__abc_52155_new_n8273_), .B(u2__abc_52155_new_n8276_), .Y(u2__abc_52155_new_n8277_));
AND2X2 AND2X2_3082 ( .A(u2__abc_52155_new_n8278_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__33_));
AND2X2 AND2X2_3083 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_34_), .Y(u2__abc_52155_new_n8280_));
AND2X2 AND2X2_3084 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_32_), .Y(u2__abc_52155_new_n8281_));
AND2X2 AND2X2_3085 ( .A(u2__abc_52155_new_n8267_), .B(u2__abc_52155_new_n3529_), .Y(u2__abc_52155_new_n8283_));
AND2X2 AND2X2_3086 ( .A(u2__abc_52155_new_n8284_), .B(u2__abc_52155_new_n8282_), .Y(u2__abc_52155_new_n8286_));
AND2X2 AND2X2_3087 ( .A(u2__abc_52155_new_n8287_), .B(u2__abc_52155_new_n8285_), .Y(u2__abc_52155_new_n8288_));
AND2X2 AND2X2_3088 ( .A(u2__abc_52155_new_n8288_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8289_));
AND2X2 AND2X2_3089 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3551_), .Y(u2__abc_52155_new_n8292_));
AND2X2 AND2X2_309 ( .A(_abc_73687_new_n1519_), .B(_abc_73687_new_n1515_), .Y(\o[227] ));
AND2X2 AND2X2_3090 ( .A(u2__abc_52155_new_n8293_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8294_));
AND2X2 AND2X2_3091 ( .A(u2__abc_52155_new_n8291_), .B(u2__abc_52155_new_n8294_), .Y(u2__abc_52155_new_n8295_));
AND2X2 AND2X2_3092 ( .A(u2__abc_52155_new_n8296_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__34_));
AND2X2 AND2X2_3093 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_35_), .Y(u2__abc_52155_new_n8298_));
AND2X2 AND2X2_3094 ( .A(u2__abc_52155_new_n8287_), .B(u2__abc_52155_new_n8300_), .Y(u2__abc_52155_new_n8301_));
AND2X2 AND2X2_3095 ( .A(u2__abc_52155_new_n8301_), .B(u2__abc_52155_new_n8299_), .Y(u2__abc_52155_new_n8302_));
AND2X2 AND2X2_3096 ( .A(u2__abc_52155_new_n8303_), .B(u2__abc_52155_new_n3516_), .Y(u2__abc_52155_new_n8304_));
AND2X2 AND2X2_3097 ( .A(u2__abc_52155_new_n8305_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8306_));
AND2X2 AND2X2_3098 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_33_), .Y(u2__abc_52155_new_n8307_));
AND2X2 AND2X2_3099 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3546_), .Y(u2__abc_52155_new_n8310_));
AND2X2 AND2X2_31 ( .A(_abc_73687_new_n753_), .B(sqrto_30_), .Y(\o[66] ));
AND2X2 AND2X2_310 ( .A(_abc_73687_new_n753_), .B(_abc_73687_new_n1521_), .Y(_abc_73687_new_n1522_));
AND2X2 AND2X2_3100 ( .A(u2__abc_52155_new_n8311_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8312_));
AND2X2 AND2X2_3101 ( .A(u2__abc_52155_new_n8309_), .B(u2__abc_52155_new_n8312_), .Y(u2__abc_52155_new_n8313_));
AND2X2 AND2X2_3102 ( .A(u2__abc_52155_new_n8314_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__35_));
AND2X2 AND2X2_3103 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_36_), .Y(u2__abc_52155_new_n8316_));
AND2X2 AND2X2_3104 ( .A(u2__abc_52155_new_n3521_), .B(u2__abc_52155_new_n3526_), .Y(u2__abc_52155_new_n8318_));
AND2X2 AND2X2_3105 ( .A(u2__abc_52155_new_n3567_), .B(u2__abc_52155_new_n3508_), .Y(u2__abc_52155_new_n8321_));
AND2X2 AND2X2_3106 ( .A(u2__abc_52155_new_n8320_), .B(u2__abc_52155_new_n8323_), .Y(u2__abc_52155_new_n8324_));
AND2X2 AND2X2_3107 ( .A(u2__abc_52155_new_n8248_), .B(u2__abc_52155_new_n3532_), .Y(u2__abc_52155_new_n8326_));
AND2X2 AND2X2_3108 ( .A(u2__abc_52155_new_n8327_), .B(u2__abc_52155_new_n8317_), .Y(u2__abc_52155_new_n8329_));
AND2X2 AND2X2_3109 ( .A(u2__abc_52155_new_n8330_), .B(u2__abc_52155_new_n8328_), .Y(u2__abc_52155_new_n8331_));
AND2X2 AND2X2_311 ( .A(_abc_73687_new_n1524_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1525_));
AND2X2 AND2X2_3110 ( .A(u2__abc_52155_new_n8332_), .B(u2__abc_52155_new_n8333_), .Y(u2__abc_52155_new_n8334_));
AND2X2 AND2X2_3111 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3535_), .Y(u2__abc_52155_new_n8336_));
AND2X2 AND2X2_3112 ( .A(u2__abc_52155_new_n8337_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8338_));
AND2X2 AND2X2_3113 ( .A(u2__abc_52155_new_n8335_), .B(u2__abc_52155_new_n8338_), .Y(u2__abc_52155_new_n8339_));
AND2X2 AND2X2_3114 ( .A(u2__abc_52155_new_n8340_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__36_));
AND2X2 AND2X2_3115 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_37_), .Y(u2__abc_52155_new_n8342_));
AND2X2 AND2X2_3116 ( .A(u2__abc_52155_new_n8330_), .B(u2__abc_52155_new_n8344_), .Y(u2__abc_52155_new_n8345_));
AND2X2 AND2X2_3117 ( .A(u2__abc_52155_new_n8347_), .B(u2__abc_52155_new_n8348_), .Y(u2__abc_52155_new_n8349_));
AND2X2 AND2X2_3118 ( .A(u2__abc_52155_new_n8349_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8350_));
AND2X2 AND2X2_3119 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_35_), .Y(u2__abc_52155_new_n8351_));
AND2X2 AND2X2_312 ( .A(_abc_73687_new_n1528_), .B(_abc_73687_new_n1529_), .Y(\o[228] ));
AND2X2 AND2X2_3120 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3540_), .Y(u2__abc_52155_new_n8354_));
AND2X2 AND2X2_3121 ( .A(u2__abc_52155_new_n8355_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8356_));
AND2X2 AND2X2_3122 ( .A(u2__abc_52155_new_n8353_), .B(u2__abc_52155_new_n8356_), .Y(u2__abc_52155_new_n8357_));
AND2X2 AND2X2_3123 ( .A(u2__abc_52155_new_n8358_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__37_));
AND2X2 AND2X2_3124 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_38_), .Y(u2__abc_52155_new_n8360_));
AND2X2 AND2X2_3125 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_36_), .Y(u2__abc_52155_new_n8361_));
AND2X2 AND2X2_3126 ( .A(u2__abc_52155_new_n8330_), .B(u2__abc_52155_new_n8364_), .Y(u2__abc_52155_new_n8365_));
AND2X2 AND2X2_3127 ( .A(u2__abc_52155_new_n8367_), .B(u2__abc_52155_new_n8362_), .Y(u2__abc_52155_new_n8369_));
AND2X2 AND2X2_3128 ( .A(u2__abc_52155_new_n8370_), .B(u2__abc_52155_new_n8368_), .Y(u2__abc_52155_new_n8371_));
AND2X2 AND2X2_3129 ( .A(u2__abc_52155_new_n8371_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8372_));
AND2X2 AND2X2_313 ( .A(\a[114] ), .B(\a[115] ), .Y(_abc_73687_new_n1531_));
AND2X2 AND2X2_3130 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3462_), .Y(u2__abc_52155_new_n8375_));
AND2X2 AND2X2_3131 ( .A(u2__abc_52155_new_n8376_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8377_));
AND2X2 AND2X2_3132 ( .A(u2__abc_52155_new_n8374_), .B(u2__abc_52155_new_n8377_), .Y(u2__abc_52155_new_n8378_));
AND2X2 AND2X2_3133 ( .A(u2__abc_52155_new_n8379_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__38_));
AND2X2 AND2X2_3134 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_39_), .Y(u2__abc_52155_new_n8381_));
AND2X2 AND2X2_3135 ( .A(u2__abc_52155_new_n8370_), .B(u2__abc_52155_new_n8382_), .Y(u2__abc_52155_new_n8383_));
AND2X2 AND2X2_3136 ( .A(u2__abc_52155_new_n8387_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8388_));
AND2X2 AND2X2_3137 ( .A(u2__abc_52155_new_n8388_), .B(u2__abc_52155_new_n8384_), .Y(u2__abc_52155_new_n8389_));
AND2X2 AND2X2_3138 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_37_), .Y(u2__abc_52155_new_n8390_));
AND2X2 AND2X2_3139 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3469_), .Y(u2__abc_52155_new_n8393_));
AND2X2 AND2X2_314 ( .A(_abc_73687_new_n1507_), .B(_abc_73687_new_n1531_), .Y(_abc_73687_new_n1532_));
AND2X2 AND2X2_3140 ( .A(u2__abc_52155_new_n8394_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8395_));
AND2X2 AND2X2_3141 ( .A(u2__abc_52155_new_n8392_), .B(u2__abc_52155_new_n8395_), .Y(u2__abc_52155_new_n8396_));
AND2X2 AND2X2_3142 ( .A(u2__abc_52155_new_n8397_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__39_));
AND2X2 AND2X2_3143 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_40_), .Y(u2__abc_52155_new_n8399_));
AND2X2 AND2X2_3144 ( .A(u2__abc_52155_new_n8325_), .B(u2__abc_52155_new_n3556_), .Y(u2__abc_52155_new_n8400_));
AND2X2 AND2X2_3145 ( .A(u2__abc_52155_new_n8404_), .B(u2__abc_52155_new_n3578_), .Y(u2__abc_52155_new_n8405_));
AND2X2 AND2X2_3146 ( .A(u2__abc_52155_new_n8403_), .B(u2__abc_52155_new_n8405_), .Y(u2__abc_52155_new_n8406_));
AND2X2 AND2X2_3147 ( .A(u2__abc_52155_new_n8401_), .B(u2__abc_52155_new_n8406_), .Y(u2__abc_52155_new_n8407_));
AND2X2 AND2X2_3148 ( .A(u2__abc_52155_new_n8248_), .B(u2__abc_52155_new_n3557_), .Y(u2__abc_52155_new_n8409_));
AND2X2 AND2X2_3149 ( .A(u2__abc_52155_new_n8410_), .B(u2__abc_52155_new_n3465_), .Y(u2__abc_52155_new_n8412_));
AND2X2 AND2X2_315 ( .A(_abc_73687_new_n1516_), .B(_abc_73687_new_n1521_), .Y(_abc_73687_new_n1533_));
AND2X2 AND2X2_3150 ( .A(u2__abc_52155_new_n8413_), .B(u2__abc_52155_new_n8411_), .Y(u2__abc_52155_new_n8414_));
AND2X2 AND2X2_3151 ( .A(u2__abc_52155_new_n8415_), .B(u2__abc_52155_new_n8416_), .Y(u2__abc_52155_new_n8417_));
AND2X2 AND2X2_3152 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3449_), .Y(u2__abc_52155_new_n8419_));
AND2X2 AND2X2_3153 ( .A(u2__abc_52155_new_n8420_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8421_));
AND2X2 AND2X2_3154 ( .A(u2__abc_52155_new_n8418_), .B(u2__abc_52155_new_n8421_), .Y(u2__abc_52155_new_n8422_));
AND2X2 AND2X2_3155 ( .A(u2__abc_52155_new_n8423_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__40_));
AND2X2 AND2X2_3156 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_41_), .Y(u2__abc_52155_new_n8425_));
AND2X2 AND2X2_3157 ( .A(u2__abc_52155_new_n8413_), .B(u2__abc_52155_new_n3461_), .Y(u2__abc_52155_new_n8427_));
AND2X2 AND2X2_3158 ( .A(u2__abc_52155_new_n8428_), .B(u2__abc_52155_new_n8426_), .Y(u2__abc_52155_new_n8429_));
AND2X2 AND2X2_3159 ( .A(u2__abc_52155_new_n8427_), .B(u2__abc_52155_new_n3472_), .Y(u2__abc_52155_new_n8430_));
AND2X2 AND2X2_316 ( .A(_abc_73687_new_n1509_), .B(_abc_73687_new_n1533_), .Y(_abc_73687_new_n1534_));
AND2X2 AND2X2_3160 ( .A(u2__abc_52155_new_n8431_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8432_));
AND2X2 AND2X2_3161 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_39_), .Y(u2__abc_52155_new_n8433_));
AND2X2 AND2X2_3162 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3454_), .Y(u2__abc_52155_new_n8436_));
AND2X2 AND2X2_3163 ( .A(u2__abc_52155_new_n8437_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8438_));
AND2X2 AND2X2_3164 ( .A(u2__abc_52155_new_n8435_), .B(u2__abc_52155_new_n8438_), .Y(u2__abc_52155_new_n8439_));
AND2X2 AND2X2_3165 ( .A(u2__abc_52155_new_n8440_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__41_));
AND2X2 AND2X2_3166 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_42_), .Y(u2__abc_52155_new_n8442_));
AND2X2 AND2X2_3167 ( .A(u2__abc_52155_new_n8428_), .B(u2__abc_52155_new_n3471_), .Y(u2__abc_52155_new_n8444_));
AND2X2 AND2X2_3168 ( .A(u2__abc_52155_new_n8445_), .B(u2__abc_52155_new_n8443_), .Y(u2__abc_52155_new_n8447_));
AND2X2 AND2X2_3169 ( .A(u2__abc_52155_new_n8448_), .B(u2__abc_52155_new_n8446_), .Y(u2__abc_52155_new_n8449_));
AND2X2 AND2X2_317 ( .A(_abc_73687_new_n1532_), .B(\a[116] ), .Y(_abc_73687_new_n1536_));
AND2X2 AND2X2_3170 ( .A(u2__abc_52155_new_n8450_), .B(u2__abc_52155_new_n8451_), .Y(u2__abc_52155_new_n8452_));
AND2X2 AND2X2_3171 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3500_), .Y(u2__abc_52155_new_n8454_));
AND2X2 AND2X2_3172 ( .A(u2__abc_52155_new_n8455_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8456_));
AND2X2 AND2X2_3173 ( .A(u2__abc_52155_new_n8453_), .B(u2__abc_52155_new_n8456_), .Y(u2__abc_52155_new_n8457_));
AND2X2 AND2X2_3174 ( .A(u2__abc_52155_new_n8458_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__42_));
AND2X2 AND2X2_3175 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_43_), .Y(u2__abc_52155_new_n8460_));
AND2X2 AND2X2_3176 ( .A(u2__abc_52155_new_n8448_), .B(u2__abc_52155_new_n8461_), .Y(u2__abc_52155_new_n8462_));
AND2X2 AND2X2_3177 ( .A(u2__abc_52155_new_n8466_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8467_));
AND2X2 AND2X2_3178 ( .A(u2__abc_52155_new_n8467_), .B(u2__abc_52155_new_n8463_), .Y(u2__abc_52155_new_n8468_));
AND2X2 AND2X2_3179 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_41_), .Y(u2__abc_52155_new_n8469_));
AND2X2 AND2X2_318 ( .A(_abc_73687_new_n1538_), .B(_abc_73687_new_n1537_), .Y(_abc_73687_new_n1539_));
AND2X2 AND2X2_3180 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3493_), .Y(u2__abc_52155_new_n8472_));
AND2X2 AND2X2_3181 ( .A(u2__abc_52155_new_n8473_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8474_));
AND2X2 AND2X2_3182 ( .A(u2__abc_52155_new_n8471_), .B(u2__abc_52155_new_n8474_), .Y(u2__abc_52155_new_n8475_));
AND2X2 AND2X2_3183 ( .A(u2__abc_52155_new_n8476_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__43_));
AND2X2 AND2X2_3184 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_44_), .Y(u2__abc_52155_new_n8478_));
AND2X2 AND2X2_3185 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_42_), .Y(u2__abc_52155_new_n8479_));
AND2X2 AND2X2_3186 ( .A(u2__abc_52155_new_n3461_), .B(u2__abc_52155_new_n3468_), .Y(u2__abc_52155_new_n8480_));
AND2X2 AND2X2_3187 ( .A(u2__abc_52155_new_n8483_), .B(u2__abc_52155_new_n3589_), .Y(u2__abc_52155_new_n8484_));
AND2X2 AND2X2_3188 ( .A(u2__abc_52155_new_n8482_), .B(u2__abc_52155_new_n8484_), .Y(u2__abc_52155_new_n8485_));
AND2X2 AND2X2_3189 ( .A(u2__abc_52155_new_n8410_), .B(u2__abc_52155_new_n3474_), .Y(u2__abc_52155_new_n8487_));
AND2X2 AND2X2_319 ( .A(_abc_73687_new_n1540_), .B(_abc_73687_new_n1535_), .Y(_abc_73687_new_n1541_));
AND2X2 AND2X2_3190 ( .A(u2__abc_52155_new_n8488_), .B(u2__abc_52155_new_n3503_), .Y(u2__abc_52155_new_n8490_));
AND2X2 AND2X2_3191 ( .A(u2__abc_52155_new_n8491_), .B(u2__abc_52155_new_n8489_), .Y(u2__abc_52155_new_n8492_));
AND2X2 AND2X2_3192 ( .A(u2__abc_52155_new_n8492_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8493_));
AND2X2 AND2X2_3193 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3478_), .Y(u2__abc_52155_new_n8496_));
AND2X2 AND2X2_3194 ( .A(u2__abc_52155_new_n8497_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8498_));
AND2X2 AND2X2_3195 ( .A(u2__abc_52155_new_n8495_), .B(u2__abc_52155_new_n8498_), .Y(u2__abc_52155_new_n8499_));
AND2X2 AND2X2_3196 ( .A(u2__abc_52155_new_n8500_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__44_));
AND2X2 AND2X2_3197 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_45_), .Y(u2__abc_52155_new_n8502_));
AND2X2 AND2X2_3198 ( .A(u2__abc_52155_new_n8491_), .B(u2__abc_52155_new_n3499_), .Y(u2__abc_52155_new_n8503_));
AND2X2 AND2X2_3199 ( .A(u2__abc_52155_new_n8503_), .B(u2__abc_52155_new_n3496_), .Y(u2__abc_52155_new_n8504_));
AND2X2 AND2X2_32 ( .A(_abc_73687_new_n753_), .B(sqrto_31_), .Y(\o[67] ));
AND2X2 AND2X2_320 ( .A(_abc_73687_new_n1542_), .B(\a[116] ), .Y(_abc_73687_new_n1543_));
AND2X2 AND2X2_3200 ( .A(u2__abc_52155_new_n8506_), .B(u2__abc_52155_new_n8505_), .Y(u2__abc_52155_new_n8507_));
AND2X2 AND2X2_3201 ( .A(u2__abc_52155_new_n8508_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8509_));
AND2X2 AND2X2_3202 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_43_), .Y(u2__abc_52155_new_n8510_));
AND2X2 AND2X2_3203 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3485_), .Y(u2__abc_52155_new_n8513_));
AND2X2 AND2X2_3204 ( .A(u2__abc_52155_new_n8514_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8515_));
AND2X2 AND2X2_3205 ( .A(u2__abc_52155_new_n8512_), .B(u2__abc_52155_new_n8515_), .Y(u2__abc_52155_new_n8516_));
AND2X2 AND2X2_3206 ( .A(u2__abc_52155_new_n8517_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__45_));
AND2X2 AND2X2_3207 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_46_), .Y(u2__abc_52155_new_n8519_));
AND2X2 AND2X2_3208 ( .A(u2__abc_52155_new_n3492_), .B(u2__abc_52155_new_n3499_), .Y(u2__abc_52155_new_n8520_));
AND2X2 AND2X2_3209 ( .A(u2__abc_52155_new_n8491_), .B(u2__abc_52155_new_n8520_), .Y(u2__abc_52155_new_n8521_));
AND2X2 AND2X2_321 ( .A(_abc_73687_new_n1544_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1545_));
AND2X2 AND2X2_3210 ( .A(u2__abc_52155_new_n8523_), .B(u2__abc_52155_new_n3481_), .Y(u2__abc_52155_new_n8524_));
AND2X2 AND2X2_3211 ( .A(u2__abc_52155_new_n8525_), .B(u2__abc_52155_new_n8526_), .Y(u2__abc_52155_new_n8527_));
AND2X2 AND2X2_3212 ( .A(u2__abc_52155_new_n8527_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8528_));
AND2X2 AND2X2_3213 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_44_), .Y(u2__abc_52155_new_n8529_));
AND2X2 AND2X2_3214 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3408_), .Y(u2__abc_52155_new_n8532_));
AND2X2 AND2X2_3215 ( .A(u2__abc_52155_new_n8533_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8534_));
AND2X2 AND2X2_3216 ( .A(u2__abc_52155_new_n8531_), .B(u2__abc_52155_new_n8534_), .Y(u2__abc_52155_new_n8535_));
AND2X2 AND2X2_3217 ( .A(u2__abc_52155_new_n8536_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__46_));
AND2X2 AND2X2_3218 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_47_), .Y(u2__abc_52155_new_n8538_));
AND2X2 AND2X2_3219 ( .A(u2__abc_52155_new_n8525_), .B(u2__abc_52155_new_n3477_), .Y(u2__abc_52155_new_n8540_));
AND2X2 AND2X2_322 ( .A(aNan), .B(\a[115] ), .Y(_abc_73687_new_n1546_));
AND2X2 AND2X2_3220 ( .A(u2__abc_52155_new_n8543_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8544_));
AND2X2 AND2X2_3221 ( .A(u2__abc_52155_new_n8544_), .B(u2__abc_52155_new_n8541_), .Y(u2__abc_52155_new_n8545_));
AND2X2 AND2X2_3222 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_45_), .Y(u2__abc_52155_new_n8546_));
AND2X2 AND2X2_3223 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3401_), .Y(u2__abc_52155_new_n8549_));
AND2X2 AND2X2_3224 ( .A(u2__abc_52155_new_n8550_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8551_));
AND2X2 AND2X2_3225 ( .A(u2__abc_52155_new_n8548_), .B(u2__abc_52155_new_n8551_), .Y(u2__abc_52155_new_n8552_));
AND2X2 AND2X2_3226 ( .A(u2__abc_52155_new_n8553_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__47_));
AND2X2 AND2X2_3227 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_48_), .Y(u2__abc_52155_new_n8555_));
AND2X2 AND2X2_3228 ( .A(u2__abc_52155_new_n8248_), .B(u2__abc_52155_new_n3558_), .Y(u2__abc_52155_new_n8556_));
AND2X2 AND2X2_3229 ( .A(u2__abc_52155_new_n8408_), .B(u2__abc_52155_new_n3506_), .Y(u2__abc_52155_new_n8557_));
AND2X2 AND2X2_323 ( .A(_abc_73687_new_n1549_), .B(_abc_73687_new_n1548_), .Y(_abc_73687_new_n1550_));
AND2X2 AND2X2_3230 ( .A(u2__abc_52155_new_n8486_), .B(u2__abc_52155_new_n3505_), .Y(u2__abc_52155_new_n8558_));
AND2X2 AND2X2_3231 ( .A(u2__abc_52155_new_n8560_), .B(u2__abc_52155_new_n3489_), .Y(u2__abc_52155_new_n8561_));
AND2X2 AND2X2_3232 ( .A(u2__abc_52155_new_n3487_), .B(u2__abc_52155_new_n3476_), .Y(u2__abc_52155_new_n8562_));
AND2X2 AND2X2_3233 ( .A(u2__abc_52155_new_n8567_), .B(u2__abc_52155_new_n3411_), .Y(u2__abc_52155_new_n8569_));
AND2X2 AND2X2_3234 ( .A(u2__abc_52155_new_n8570_), .B(u2__abc_52155_new_n8568_), .Y(u2__abc_52155_new_n8571_));
AND2X2 AND2X2_3235 ( .A(u2__abc_52155_new_n8572_), .B(u2__abc_52155_new_n8573_), .Y(u2__abc_52155_new_n8574_));
AND2X2 AND2X2_3236 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3388_), .Y(u2__abc_52155_new_n8576_));
AND2X2 AND2X2_3237 ( .A(u2__abc_52155_new_n8577_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8578_));
AND2X2 AND2X2_3238 ( .A(u2__abc_52155_new_n8575_), .B(u2__abc_52155_new_n8578_), .Y(u2__abc_52155_new_n8579_));
AND2X2 AND2X2_3239 ( .A(u2__abc_52155_new_n8580_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__48_));
AND2X2 AND2X2_324 ( .A(_abc_73687_new_n1536_), .B(\a[117] ), .Y(_abc_73687_new_n1551_));
AND2X2 AND2X2_3240 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_49_), .Y(u2__abc_52155_new_n8582_));
AND2X2 AND2X2_3241 ( .A(u2__abc_52155_new_n8570_), .B(u2__abc_52155_new_n3407_), .Y(u2__abc_52155_new_n8583_));
AND2X2 AND2X2_3242 ( .A(u2__abc_52155_new_n8585_), .B(u2__abc_52155_new_n8587_), .Y(u2__abc_52155_new_n8588_));
AND2X2 AND2X2_3243 ( .A(u2__abc_52155_new_n8588_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8589_));
AND2X2 AND2X2_3244 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_47_), .Y(u2__abc_52155_new_n8590_));
AND2X2 AND2X2_3245 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3393_), .Y(u2__abc_52155_new_n8593_));
AND2X2 AND2X2_3246 ( .A(u2__abc_52155_new_n8594_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8595_));
AND2X2 AND2X2_3247 ( .A(u2__abc_52155_new_n8592_), .B(u2__abc_52155_new_n8595_), .Y(u2__abc_52155_new_n8596_));
AND2X2 AND2X2_3248 ( .A(u2__abc_52155_new_n8597_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__49_));
AND2X2 AND2X2_3249 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_50_), .Y(u2__abc_52155_new_n8599_));
AND2X2 AND2X2_325 ( .A(_abc_73687_new_n1552_), .B(_abc_73687_new_n1541_), .Y(_abc_73687_new_n1553_));
AND2X2 AND2X2_3250 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_48_), .Y(u2__abc_52155_new_n8600_));
AND2X2 AND2X2_3251 ( .A(u2__abc_52155_new_n3400_), .B(u2__abc_52155_new_n3407_), .Y(u2__abc_52155_new_n8602_));
AND2X2 AND2X2_3252 ( .A(u2__abc_52155_new_n8570_), .B(u2__abc_52155_new_n8602_), .Y(u2__abc_52155_new_n8603_));
AND2X2 AND2X2_3253 ( .A(u2__abc_52155_new_n8605_), .B(u2__abc_52155_new_n8601_), .Y(u2__abc_52155_new_n8607_));
AND2X2 AND2X2_3254 ( .A(u2__abc_52155_new_n8608_), .B(u2__abc_52155_new_n8606_), .Y(u2__abc_52155_new_n8609_));
AND2X2 AND2X2_3255 ( .A(u2__abc_52155_new_n8609_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8610_));
AND2X2 AND2X2_3256 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3439_), .Y(u2__abc_52155_new_n8613_));
AND2X2 AND2X2_3257 ( .A(u2__abc_52155_new_n8614_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8615_));
AND2X2 AND2X2_3258 ( .A(u2__abc_52155_new_n8612_), .B(u2__abc_52155_new_n8615_), .Y(u2__abc_52155_new_n8616_));
AND2X2 AND2X2_3259 ( .A(u2__abc_52155_new_n8617_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__50_));
AND2X2 AND2X2_326 ( .A(_abc_73687_new_n1554_), .B(_abc_73687_new_n1555_), .Y(_abc_73687_new_n1556_));
AND2X2 AND2X2_3260 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_51_), .Y(u2__abc_52155_new_n8619_));
AND2X2 AND2X2_3261 ( .A(u2__abc_52155_new_n8608_), .B(u2__abc_52155_new_n8620_), .Y(u2__abc_52155_new_n8621_));
AND2X2 AND2X2_3262 ( .A(u2__abc_52155_new_n8625_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8626_));
AND2X2 AND2X2_3263 ( .A(u2__abc_52155_new_n8626_), .B(u2__abc_52155_new_n8622_), .Y(u2__abc_52155_new_n8627_));
AND2X2 AND2X2_3264 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_49_), .Y(u2__abc_52155_new_n8628_));
AND2X2 AND2X2_3265 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3432_), .Y(u2__abc_52155_new_n8631_));
AND2X2 AND2X2_3266 ( .A(u2__abc_52155_new_n8632_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8633_));
AND2X2 AND2X2_3267 ( .A(u2__abc_52155_new_n8630_), .B(u2__abc_52155_new_n8633_), .Y(u2__abc_52155_new_n8634_));
AND2X2 AND2X2_3268 ( .A(u2__abc_52155_new_n8635_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__51_));
AND2X2 AND2X2_3269 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_52_), .Y(u2__abc_52155_new_n8637_));
AND2X2 AND2X2_327 ( .A(_abc_73687_new_n1558_), .B(_abc_73687_new_n1559_), .Y(\o[230] ));
AND2X2 AND2X2_3270 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_50_), .Y(u2__abc_52155_new_n8638_));
AND2X2 AND2X2_3271 ( .A(u2__abc_52155_new_n8641_), .B(u2__abc_52155_new_n3610_), .Y(u2__abc_52155_new_n8642_));
AND2X2 AND2X2_3272 ( .A(u2__abc_52155_new_n8640_), .B(u2__abc_52155_new_n8642_), .Y(u2__abc_52155_new_n8643_));
AND2X2 AND2X2_3273 ( .A(u2__abc_52155_new_n8567_), .B(u2__abc_52155_new_n3413_), .Y(u2__abc_52155_new_n8645_));
AND2X2 AND2X2_3274 ( .A(u2__abc_52155_new_n8646_), .B(u2__abc_52155_new_n3442_), .Y(u2__abc_52155_new_n8648_));
AND2X2 AND2X2_3275 ( .A(u2__abc_52155_new_n8649_), .B(u2__abc_52155_new_n8647_), .Y(u2__abc_52155_new_n8650_));
AND2X2 AND2X2_3276 ( .A(u2__abc_52155_new_n8650_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8651_));
AND2X2 AND2X2_3277 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3417_), .Y(u2__abc_52155_new_n8654_));
AND2X2 AND2X2_3278 ( .A(u2__abc_52155_new_n8655_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8656_));
AND2X2 AND2X2_3279 ( .A(u2__abc_52155_new_n8653_), .B(u2__abc_52155_new_n8656_), .Y(u2__abc_52155_new_n8657_));
AND2X2 AND2X2_328 ( .A(aNan), .B(\a[117] ), .Y(_abc_73687_new_n1561_));
AND2X2 AND2X2_3280 ( .A(u2__abc_52155_new_n8658_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__52_));
AND2X2 AND2X2_3281 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_53_), .Y(u2__abc_52155_new_n8660_));
AND2X2 AND2X2_3282 ( .A(u2__abc_52155_new_n8649_), .B(u2__abc_52155_new_n3438_), .Y(u2__abc_52155_new_n8661_));
AND2X2 AND2X2_3283 ( .A(u2__abc_52155_new_n8661_), .B(u2__abc_52155_new_n3435_), .Y(u2__abc_52155_new_n8662_));
AND2X2 AND2X2_3284 ( .A(u2__abc_52155_new_n8664_), .B(u2__abc_52155_new_n8663_), .Y(u2__abc_52155_new_n8665_));
AND2X2 AND2X2_3285 ( .A(u2__abc_52155_new_n8666_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8667_));
AND2X2 AND2X2_3286 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_51_), .Y(u2__abc_52155_new_n8668_));
AND2X2 AND2X2_3287 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3424_), .Y(u2__abc_52155_new_n8671_));
AND2X2 AND2X2_3288 ( .A(u2__abc_52155_new_n8672_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8673_));
AND2X2 AND2X2_3289 ( .A(u2__abc_52155_new_n8670_), .B(u2__abc_52155_new_n8673_), .Y(u2__abc_52155_new_n8674_));
AND2X2 AND2X2_329 ( .A(_abc_73687_new_n1551_), .B(\a[118] ), .Y(_abc_73687_new_n1562_));
AND2X2 AND2X2_3290 ( .A(u2__abc_52155_new_n8675_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__53_));
AND2X2 AND2X2_3291 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_54_), .Y(u2__abc_52155_new_n8677_));
AND2X2 AND2X2_3292 ( .A(u2__abc_52155_new_n3431_), .B(u2__abc_52155_new_n3438_), .Y(u2__abc_52155_new_n8678_));
AND2X2 AND2X2_3293 ( .A(u2__abc_52155_new_n8649_), .B(u2__abc_52155_new_n8678_), .Y(u2__abc_52155_new_n8679_));
AND2X2 AND2X2_3294 ( .A(u2__abc_52155_new_n8681_), .B(u2__abc_52155_new_n3420_), .Y(u2__abc_52155_new_n8682_));
AND2X2 AND2X2_3295 ( .A(u2__abc_52155_new_n8683_), .B(u2__abc_52155_new_n8684_), .Y(u2__abc_52155_new_n8685_));
AND2X2 AND2X2_3296 ( .A(u2__abc_52155_new_n8685_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8686_));
AND2X2 AND2X2_3297 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_52_), .Y(u2__abc_52155_new_n8687_));
AND2X2 AND2X2_3298 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3341_), .Y(u2__abc_52155_new_n8690_));
AND2X2 AND2X2_3299 ( .A(u2__abc_52155_new_n8691_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8692_));
AND2X2 AND2X2_33 ( .A(_abc_73687_new_n753_), .B(sqrto_32_), .Y(\o[68] ));
AND2X2 AND2X2_330 ( .A(_abc_73687_new_n1564_), .B(_abc_73687_new_n1563_), .Y(_abc_73687_new_n1565_));
AND2X2 AND2X2_3300 ( .A(u2__abc_52155_new_n8689_), .B(u2__abc_52155_new_n8692_), .Y(u2__abc_52155_new_n8693_));
AND2X2 AND2X2_3301 ( .A(u2__abc_52155_new_n8694_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__54_));
AND2X2 AND2X2_3302 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_55_), .Y(u2__abc_52155_new_n8696_));
AND2X2 AND2X2_3303 ( .A(u2__abc_52155_new_n8683_), .B(u2__abc_52155_new_n3416_), .Y(u2__abc_52155_new_n8698_));
AND2X2 AND2X2_3304 ( .A(u2__abc_52155_new_n8701_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8702_));
AND2X2 AND2X2_3305 ( .A(u2__abc_52155_new_n8702_), .B(u2__abc_52155_new_n8699_), .Y(u2__abc_52155_new_n8703_));
AND2X2 AND2X2_3306 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_53_), .Y(u2__abc_52155_new_n8704_));
AND2X2 AND2X2_3307 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3348_), .Y(u2__abc_52155_new_n8707_));
AND2X2 AND2X2_3308 ( .A(u2__abc_52155_new_n8708_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8709_));
AND2X2 AND2X2_3309 ( .A(u2__abc_52155_new_n8706_), .B(u2__abc_52155_new_n8709_), .Y(u2__abc_52155_new_n8710_));
AND2X2 AND2X2_331 ( .A(_abc_73687_new_n1553_), .B(_abc_73687_new_n1566_), .Y(_abc_73687_new_n1567_));
AND2X2 AND2X2_3310 ( .A(u2__abc_52155_new_n8711_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__55_));
AND2X2 AND2X2_3311 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_56_), .Y(u2__abc_52155_new_n8713_));
AND2X2 AND2X2_3312 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_54_), .Y(u2__abc_52155_new_n8714_));
AND2X2 AND2X2_3313 ( .A(u2__abc_52155_new_n8644_), .B(u2__abc_52155_new_n3444_), .Y(u2__abc_52155_new_n8715_));
AND2X2 AND2X2_3314 ( .A(u2__abc_52155_new_n8717_), .B(u2__abc_52155_new_n3428_), .Y(u2__abc_52155_new_n8718_));
AND2X2 AND2X2_3315 ( .A(u2__abc_52155_new_n3426_), .B(u2__abc_52155_new_n3415_), .Y(u2__abc_52155_new_n8719_));
AND2X2 AND2X2_3316 ( .A(u2__abc_52155_new_n8567_), .B(u2__abc_52155_new_n3445_), .Y(u2__abc_52155_new_n8723_));
AND2X2 AND2X2_3317 ( .A(u2__abc_52155_new_n8724_), .B(u2__abc_52155_new_n3344_), .Y(u2__abc_52155_new_n8726_));
AND2X2 AND2X2_3318 ( .A(u2__abc_52155_new_n8727_), .B(u2__abc_52155_new_n8725_), .Y(u2__abc_52155_new_n8728_));
AND2X2 AND2X2_3319 ( .A(u2__abc_52155_new_n8728_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8729_));
AND2X2 AND2X2_332 ( .A(_abc_73687_new_n1568_), .B(_abc_73687_new_n1569_), .Y(_abc_73687_new_n1570_));
AND2X2 AND2X2_3320 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3326_), .Y(u2__abc_52155_new_n8732_));
AND2X2 AND2X2_3321 ( .A(u2__abc_52155_new_n8733_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8734_));
AND2X2 AND2X2_3322 ( .A(u2__abc_52155_new_n8731_), .B(u2__abc_52155_new_n8734_), .Y(u2__abc_52155_new_n8735_));
AND2X2 AND2X2_3323 ( .A(u2__abc_52155_new_n8736_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__56_));
AND2X2 AND2X2_3324 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_57_), .Y(u2__abc_52155_new_n8738_));
AND2X2 AND2X2_3325 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_55_), .Y(u2__abc_52155_new_n8739_));
AND2X2 AND2X2_3326 ( .A(u2__abc_52155_new_n8727_), .B(u2__abc_52155_new_n3340_), .Y(u2__abc_52155_new_n8742_));
AND2X2 AND2X2_3327 ( .A(u2__abc_52155_new_n8745_), .B(u2__abc_52155_new_n8743_), .Y(u2__abc_52155_new_n8746_));
AND2X2 AND2X2_3328 ( .A(u2__abc_52155_new_n8746_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8747_));
AND2X2 AND2X2_3329 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3333_), .Y(u2__abc_52155_new_n8749_));
AND2X2 AND2X2_333 ( .A(_abc_73687_new_n1571_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1572_));
AND2X2 AND2X2_3330 ( .A(u2__abc_52155_new_n8750_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8751_));
AND2X2 AND2X2_3331 ( .A(u2__abc_52155_new_n8748_), .B(u2__abc_52155_new_n8751_), .Y(u2__abc_52155_new_n8752_));
AND2X2 AND2X2_3332 ( .A(u2__abc_52155_new_n8753_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__57_));
AND2X2 AND2X2_3333 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_58_), .Y(u2__abc_52155_new_n8755_));
AND2X2 AND2X2_3334 ( .A(u2__abc_52155_new_n3340_), .B(u2__abc_52155_new_n3347_), .Y(u2__abc_52155_new_n8756_));
AND2X2 AND2X2_3335 ( .A(u2__abc_52155_new_n8724_), .B(u2__abc_52155_new_n3352_), .Y(u2__abc_52155_new_n8759_));
AND2X2 AND2X2_3336 ( .A(u2__abc_52155_new_n8760_), .B(u2__abc_52155_new_n3329_), .Y(u2__abc_52155_new_n8761_));
AND2X2 AND2X2_3337 ( .A(u2__abc_52155_new_n8762_), .B(u2__abc_52155_new_n8763_), .Y(u2__abc_52155_new_n8764_));
AND2X2 AND2X2_3338 ( .A(u2__abc_52155_new_n8764_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8765_));
AND2X2 AND2X2_3339 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_56_), .Y(u2__abc_52155_new_n8766_));
AND2X2 AND2X2_334 ( .A(_abc_73687_new_n1576_), .B(_abc_73687_new_n1575_), .Y(_abc_73687_new_n1577_));
AND2X2 AND2X2_3340 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3379_), .Y(u2__abc_52155_new_n8769_));
AND2X2 AND2X2_3341 ( .A(u2__abc_52155_new_n8770_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8771_));
AND2X2 AND2X2_3342 ( .A(u2__abc_52155_new_n8768_), .B(u2__abc_52155_new_n8771_), .Y(u2__abc_52155_new_n8772_));
AND2X2 AND2X2_3343 ( .A(u2__abc_52155_new_n8773_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__58_));
AND2X2 AND2X2_3344 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_59_), .Y(u2__abc_52155_new_n8775_));
AND2X2 AND2X2_3345 ( .A(u2__abc_52155_new_n8762_), .B(u2__abc_52155_new_n3325_), .Y(u2__abc_52155_new_n8777_));
AND2X2 AND2X2_3346 ( .A(u2__abc_52155_new_n8780_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8781_));
AND2X2 AND2X2_3347 ( .A(u2__abc_52155_new_n8781_), .B(u2__abc_52155_new_n8778_), .Y(u2__abc_52155_new_n8782_));
AND2X2 AND2X2_3348 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_57_), .Y(u2__abc_52155_new_n8783_));
AND2X2 AND2X2_3349 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3372_), .Y(u2__abc_52155_new_n8786_));
AND2X2 AND2X2_335 ( .A(_abc_73687_new_n1562_), .B(\a[119] ), .Y(_abc_73687_new_n1578_));
AND2X2 AND2X2_3350 ( .A(u2__abc_52155_new_n8787_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8788_));
AND2X2 AND2X2_3351 ( .A(u2__abc_52155_new_n8785_), .B(u2__abc_52155_new_n8788_), .Y(u2__abc_52155_new_n8789_));
AND2X2 AND2X2_3352 ( .A(u2__abc_52155_new_n8790_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__59_));
AND2X2 AND2X2_3353 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_60_), .Y(u2__abc_52155_new_n8792_));
AND2X2 AND2X2_3354 ( .A(u2__abc_52155_new_n8758_), .B(u2__abc_52155_new_n3337_), .Y(u2__abc_52155_new_n8793_));
AND2X2 AND2X2_3355 ( .A(u2__abc_52155_new_n3335_), .B(u2__abc_52155_new_n3324_), .Y(u2__abc_52155_new_n8794_));
AND2X2 AND2X2_3356 ( .A(u2__abc_52155_new_n8724_), .B(u2__abc_52155_new_n3353_), .Y(u2__abc_52155_new_n8797_));
AND2X2 AND2X2_3357 ( .A(u2__abc_52155_new_n8798_), .B(u2__abc_52155_new_n3382_), .Y(u2__abc_52155_new_n8799_));
AND2X2 AND2X2_3358 ( .A(u2__abc_52155_new_n8800_), .B(u2__abc_52155_new_n8801_), .Y(u2__abc_52155_new_n8802_));
AND2X2 AND2X2_3359 ( .A(u2__abc_52155_new_n8802_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8803_));
AND2X2 AND2X2_336 ( .A(_abc_73687_new_n1574_), .B(_abc_73687_new_n1580_), .Y(_abc_73687_new_n1581_));
AND2X2 AND2X2_3360 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_58_), .Y(u2__abc_52155_new_n8804_));
AND2X2 AND2X2_3361 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3357_), .Y(u2__abc_52155_new_n8807_));
AND2X2 AND2X2_3362 ( .A(u2__abc_52155_new_n8808_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8809_));
AND2X2 AND2X2_3363 ( .A(u2__abc_52155_new_n8806_), .B(u2__abc_52155_new_n8809_), .Y(u2__abc_52155_new_n8810_));
AND2X2 AND2X2_3364 ( .A(u2__abc_52155_new_n8811_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__60_));
AND2X2 AND2X2_3365 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_61_), .Y(u2__abc_52155_new_n8813_));
AND2X2 AND2X2_3366 ( .A(u2__abc_52155_new_n8800_), .B(u2__abc_52155_new_n3378_), .Y(u2__abc_52155_new_n8814_));
AND2X2 AND2X2_3367 ( .A(u2__abc_52155_new_n8815_), .B(u2__abc_52155_new_n3375_), .Y(u2__abc_52155_new_n8817_));
AND2X2 AND2X2_3368 ( .A(u2__abc_52155_new_n8818_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8819_));
AND2X2 AND2X2_3369 ( .A(u2__abc_52155_new_n8819_), .B(u2__abc_52155_new_n8816_), .Y(u2__abc_52155_new_n8820_));
AND2X2 AND2X2_337 ( .A(_abc_73687_new_n1567_), .B(_abc_73687_new_n1579_), .Y(_abc_73687_new_n1582_));
AND2X2 AND2X2_3370 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_59_), .Y(u2__abc_52155_new_n8821_));
AND2X2 AND2X2_3371 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3361_), .Y(u2__abc_52155_new_n8824_));
AND2X2 AND2X2_3372 ( .A(u2__abc_52155_new_n8825_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8826_));
AND2X2 AND2X2_3373 ( .A(u2__abc_52155_new_n8823_), .B(u2__abc_52155_new_n8826_), .Y(u2__abc_52155_new_n8827_));
AND2X2 AND2X2_3374 ( .A(u2__abc_52155_new_n8828_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__61_));
AND2X2 AND2X2_3375 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_62_), .Y(u2__abc_52155_new_n8830_));
AND2X2 AND2X2_3376 ( .A(u2__abc_52155_new_n8818_), .B(u2__abc_52155_new_n3371_), .Y(u2__abc_52155_new_n8831_));
AND2X2 AND2X2_3377 ( .A(u2__abc_52155_new_n8832_), .B(u2__abc_52155_new_n3360_), .Y(u2__abc_52155_new_n8833_));
AND2X2 AND2X2_3378 ( .A(u2__abc_52155_new_n8835_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8836_));
AND2X2 AND2X2_3379 ( .A(u2__abc_52155_new_n8836_), .B(u2__abc_52155_new_n8834_), .Y(u2__abc_52155_new_n8837_));
AND2X2 AND2X2_338 ( .A(_abc_73687_new_n1583_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1584_));
AND2X2 AND2X2_3380 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_60_), .Y(u2__abc_52155_new_n8838_));
AND2X2 AND2X2_3381 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n8841_), .Y(u2__abc_52155_new_n8842_));
AND2X2 AND2X2_3382 ( .A(u2__abc_52155_new_n8843_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8844_));
AND2X2 AND2X2_3383 ( .A(u2__abc_52155_new_n8840_), .B(u2__abc_52155_new_n8844_), .Y(u2__abc_52155_new_n8845_));
AND2X2 AND2X2_3384 ( .A(u2__abc_52155_new_n8846_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__62_));
AND2X2 AND2X2_3385 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_63_), .Y(u2__abc_52155_new_n8848_));
AND2X2 AND2X2_3386 ( .A(u2__abc_52155_new_n8834_), .B(u2__abc_52155_new_n3356_), .Y(u2__abc_52155_new_n8850_));
AND2X2 AND2X2_3387 ( .A(u2__abc_52155_new_n8853_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8854_));
AND2X2 AND2X2_3388 ( .A(u2__abc_52155_new_n8854_), .B(u2__abc_52155_new_n8851_), .Y(u2__abc_52155_new_n8855_));
AND2X2 AND2X2_3389 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_61_), .Y(u2__abc_52155_new_n8856_));
AND2X2 AND2X2_339 ( .A(aNan), .B(\a[118] ), .Y(_abc_73687_new_n1585_));
AND2X2 AND2X2_3390 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4087_), .Y(u2__abc_52155_new_n8859_));
AND2X2 AND2X2_3391 ( .A(u2__abc_52155_new_n8860_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8861_));
AND2X2 AND2X2_3392 ( .A(u2__abc_52155_new_n8858_), .B(u2__abc_52155_new_n8861_), .Y(u2__abc_52155_new_n8862_));
AND2X2 AND2X2_3393 ( .A(u2__abc_52155_new_n8863_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__63_));
AND2X2 AND2X2_3394 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_64_), .Y(u2__abc_52155_new_n8865_));
AND2X2 AND2X2_3395 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_62_), .Y(u2__abc_52155_new_n8866_));
AND2X2 AND2X2_3396 ( .A(u2__abc_52155_new_n8722_), .B(u2__abc_52155_new_n3385_), .Y(u2__abc_52155_new_n8867_));
AND2X2 AND2X2_3397 ( .A(u2__abc_52155_new_n8796_), .B(u2__abc_52155_new_n3384_), .Y(u2__abc_52155_new_n8868_));
AND2X2 AND2X2_3398 ( .A(u2__abc_52155_new_n8869_), .B(u2__abc_52155_new_n3374_), .Y(u2__abc_52155_new_n8870_));
AND2X2 AND2X2_3399 ( .A(u2__abc_52155_new_n3368_), .B(u2__abc_52155_new_n8870_), .Y(u2__abc_52155_new_n8871_));
AND2X2 AND2X2_34 ( .A(_abc_73687_new_n753_), .B(sqrto_33_), .Y(\o[69] ));
AND2X2 AND2X2_340 ( .A(aNan), .B(\a[119] ), .Y(_abc_73687_new_n1587_));
AND2X2 AND2X2_3400 ( .A(u2__abc_52155_new_n3363_), .B(u2__abc_52155_new_n3355_), .Y(u2__abc_52155_new_n8872_));
AND2X2 AND2X2_3401 ( .A(u2__abc_52155_new_n8567_), .B(u2__abc_52155_new_n3446_), .Y(u2__abc_52155_new_n8877_));
AND2X2 AND2X2_3402 ( .A(u2__abc_52155_new_n8878_), .B(u2__abc_52155_new_n4083_), .Y(u2__abc_52155_new_n8880_));
AND2X2 AND2X2_3403 ( .A(u2__abc_52155_new_n8881_), .B(u2__abc_52155_new_n8879_), .Y(u2__abc_52155_new_n8882_));
AND2X2 AND2X2_3404 ( .A(u2__abc_52155_new_n8882_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8883_));
AND2X2 AND2X2_3405 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n4094_), .Y(u2__abc_52155_new_n8886_));
AND2X2 AND2X2_3406 ( .A(u2__abc_52155_new_n8887_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8888_));
AND2X2 AND2X2_3407 ( .A(u2__abc_52155_new_n8885_), .B(u2__abc_52155_new_n8888_), .Y(u2__abc_52155_new_n8889_));
AND2X2 AND2X2_3408 ( .A(u2__abc_52155_new_n8890_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__64_));
AND2X2 AND2X2_3409 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_65_), .Y(u2__abc_52155_new_n8892_));
AND2X2 AND2X2_341 ( .A(_abc_73687_new_n1578_), .B(\a[120] ), .Y(_abc_73687_new_n1588_));
AND2X2 AND2X2_3410 ( .A(u2__abc_52155_new_n8881_), .B(u2__abc_52155_new_n4081_), .Y(u2__abc_52155_new_n8893_));
AND2X2 AND2X2_3411 ( .A(u2__abc_52155_new_n8897_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8898_));
AND2X2 AND2X2_3412 ( .A(u2__abc_52155_new_n8898_), .B(u2__abc_52155_new_n8895_), .Y(u2__abc_52155_new_n8899_));
AND2X2 AND2X2_3413 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_63_), .Y(u2__abc_52155_new_n8900_));
AND2X2 AND2X2_3414 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n4099_), .Y(u2__abc_52155_new_n8903_));
AND2X2 AND2X2_3415 ( .A(u2__abc_52155_new_n8904_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8905_));
AND2X2 AND2X2_3416 ( .A(u2__abc_52155_new_n8902_), .B(u2__abc_52155_new_n8905_), .Y(u2__abc_52155_new_n8906_));
AND2X2 AND2X2_3417 ( .A(u2__abc_52155_new_n8907_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__65_));
AND2X2 AND2X2_3418 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_66_), .Y(u2__abc_52155_new_n8909_));
AND2X2 AND2X2_3419 ( .A(u2__abc_52155_new_n8911_), .B(u2__abc_52155_new_n4086_), .Y(u2__abc_52155_new_n8912_));
AND2X2 AND2X2_342 ( .A(_abc_73687_new_n1590_), .B(_abc_73687_new_n1589_), .Y(_abc_73687_new_n1591_));
AND2X2 AND2X2_3420 ( .A(u2__abc_52155_new_n8878_), .B(u2__abc_52155_new_n4091_), .Y(u2__abc_52155_new_n8914_));
AND2X2 AND2X2_3421 ( .A(u2__abc_52155_new_n8915_), .B(u2__abc_52155_new_n8910_), .Y(u2__abc_52155_new_n8917_));
AND2X2 AND2X2_3422 ( .A(u2__abc_52155_new_n8918_), .B(u2__abc_52155_new_n8916_), .Y(u2__abc_52155_new_n8919_));
AND2X2 AND2X2_3423 ( .A(u2__abc_52155_new_n8920_), .B(u2__abc_52155_new_n8921_), .Y(u2__abc_52155_new_n8922_));
AND2X2 AND2X2_3424 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n4123_), .Y(u2__abc_52155_new_n8924_));
AND2X2 AND2X2_3425 ( .A(u2__abc_52155_new_n8925_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8926_));
AND2X2 AND2X2_3426 ( .A(u2__abc_52155_new_n8923_), .B(u2__abc_52155_new_n8926_), .Y(u2__abc_52155_new_n8927_));
AND2X2 AND2X2_3427 ( .A(u2__abc_52155_new_n8928_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__66_));
AND2X2 AND2X2_3428 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_67_), .Y(u2__abc_52155_new_n8930_));
AND2X2 AND2X2_3429 ( .A(u2__abc_52155_new_n8918_), .B(u2__abc_52155_new_n8931_), .Y(u2__abc_52155_new_n8932_));
AND2X2 AND2X2_343 ( .A(_abc_73687_new_n1582_), .B(_abc_73687_new_n1592_), .Y(_abc_73687_new_n1593_));
AND2X2 AND2X2_3430 ( .A(u2__abc_52155_new_n8936_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8937_));
AND2X2 AND2X2_3431 ( .A(u2__abc_52155_new_n8937_), .B(u2__abc_52155_new_n8933_), .Y(u2__abc_52155_new_n8938_));
AND2X2 AND2X2_3432 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_65_), .Y(u2__abc_52155_new_n8939_));
AND2X2 AND2X2_3433 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4118_), .Y(u2__abc_52155_new_n8942_));
AND2X2 AND2X2_3434 ( .A(u2__abc_52155_new_n8943_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8944_));
AND2X2 AND2X2_3435 ( .A(u2__abc_52155_new_n8941_), .B(u2__abc_52155_new_n8944_), .Y(u2__abc_52155_new_n8945_));
AND2X2 AND2X2_3436 ( .A(u2__abc_52155_new_n8946_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__67_));
AND2X2 AND2X2_3437 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_68_), .Y(u2__abc_52155_new_n8948_));
AND2X2 AND2X2_3438 ( .A(u2__abc_52155_new_n8913_), .B(u2__abc_52155_new_n4103_), .Y(u2__abc_52155_new_n8950_));
AND2X2 AND2X2_3439 ( .A(u2__abc_52155_new_n4141_), .B(u2__abc_52155_new_n4093_), .Y(u2__abc_52155_new_n8951_));
AND2X2 AND2X2_344 ( .A(_abc_73687_new_n1594_), .B(_abc_73687_new_n1595_), .Y(_abc_73687_new_n1596_));
AND2X2 AND2X2_3440 ( .A(u2__abc_52155_new_n8878_), .B(u2__abc_52155_new_n4104_), .Y(u2__abc_52155_new_n8954_));
AND2X2 AND2X2_3441 ( .A(u2__abc_52155_new_n8955_), .B(u2__abc_52155_new_n8949_), .Y(u2__abc_52155_new_n8957_));
AND2X2 AND2X2_3442 ( .A(u2__abc_52155_new_n8958_), .B(u2__abc_52155_new_n8956_), .Y(u2__abc_52155_new_n8959_));
AND2X2 AND2X2_3443 ( .A(u2__abc_52155_new_n8960_), .B(u2__abc_52155_new_n8961_), .Y(u2__abc_52155_new_n8962_));
AND2X2 AND2X2_3444 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n4107_), .Y(u2__abc_52155_new_n8964_));
AND2X2 AND2X2_3445 ( .A(u2__abc_52155_new_n8965_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8966_));
AND2X2 AND2X2_3446 ( .A(u2__abc_52155_new_n8963_), .B(u2__abc_52155_new_n8966_), .Y(u2__abc_52155_new_n8967_));
AND2X2 AND2X2_3447 ( .A(u2__abc_52155_new_n8968_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__68_));
AND2X2 AND2X2_3448 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_69_), .Y(u2__abc_52155_new_n8970_));
AND2X2 AND2X2_3449 ( .A(u2__abc_52155_new_n8958_), .B(u2__abc_52155_new_n8972_), .Y(u2__abc_52155_new_n8973_));
AND2X2 AND2X2_345 ( .A(_abc_73687_new_n1597_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1598_));
AND2X2 AND2X2_3450 ( .A(u2__abc_52155_new_n8974_), .B(u2__abc_52155_new_n8971_), .Y(u2__abc_52155_new_n8975_));
AND2X2 AND2X2_3451 ( .A(u2__abc_52155_new_n8976_), .B(u2__abc_52155_new_n8977_), .Y(u2__abc_52155_new_n8978_));
AND2X2 AND2X2_3452 ( .A(u2__abc_52155_new_n8978_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8979_));
AND2X2 AND2X2_3453 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_67_), .Y(u2__abc_52155_new_n8980_));
AND2X2 AND2X2_3454 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4112_), .Y(u2__abc_52155_new_n8983_));
AND2X2 AND2X2_3455 ( .A(u2__abc_52155_new_n8984_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n8985_));
AND2X2 AND2X2_3456 ( .A(u2__abc_52155_new_n8982_), .B(u2__abc_52155_new_n8985_), .Y(u2__abc_52155_new_n8986_));
AND2X2 AND2X2_3457 ( .A(u2__abc_52155_new_n8987_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__69_));
AND2X2 AND2X2_3458 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_70_), .Y(u2__abc_52155_new_n8989_));
AND2X2 AND2X2_3459 ( .A(u2__abc_52155_new_n8991_), .B(u2__abc_52155_new_n8990_), .Y(u2__abc_52155_new_n8992_));
AND2X2 AND2X2_346 ( .A(_abc_73687_new_n1588_), .B(\a[121] ), .Y(_abc_73687_new_n1600_));
AND2X2 AND2X2_3460 ( .A(u2__abc_52155_new_n8994_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n8995_));
AND2X2 AND2X2_3461 ( .A(u2__abc_52155_new_n8995_), .B(u2__abc_52155_new_n8993_), .Y(u2__abc_52155_new_n8996_));
AND2X2 AND2X2_3462 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_68_), .Y(u2__abc_52155_new_n8997_));
AND2X2 AND2X2_3463 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4022_), .Y(u2__abc_52155_new_n9000_));
AND2X2 AND2X2_3464 ( .A(u2__abc_52155_new_n9001_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9002_));
AND2X2 AND2X2_3465 ( .A(u2__abc_52155_new_n8999_), .B(u2__abc_52155_new_n9002_), .Y(u2__abc_52155_new_n9003_));
AND2X2 AND2X2_3466 ( .A(u2__abc_52155_new_n9004_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__70_));
AND2X2 AND2X2_3467 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_71_), .Y(u2__abc_52155_new_n9006_));
AND2X2 AND2X2_3468 ( .A(u2__abc_52155_new_n8993_), .B(u2__abc_52155_new_n9007_), .Y(u2__abc_52155_new_n9008_));
AND2X2 AND2X2_3469 ( .A(u2__abc_52155_new_n9012_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9013_));
AND2X2 AND2X2_347 ( .A(_abc_73687_new_n1602_), .B(_abc_73687_new_n1601_), .Y(_abc_73687_new_n1603_));
AND2X2 AND2X2_3470 ( .A(u2__abc_52155_new_n9013_), .B(u2__abc_52155_new_n9009_), .Y(u2__abc_52155_new_n9014_));
AND2X2 AND2X2_3471 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_69_), .Y(u2__abc_52155_new_n9015_));
AND2X2 AND2X2_3472 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4029_), .Y(u2__abc_52155_new_n9018_));
AND2X2 AND2X2_3473 ( .A(u2__abc_52155_new_n9019_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9020_));
AND2X2 AND2X2_3474 ( .A(u2__abc_52155_new_n9017_), .B(u2__abc_52155_new_n9020_), .Y(u2__abc_52155_new_n9021_));
AND2X2 AND2X2_3475 ( .A(u2__abc_52155_new_n9022_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__71_));
AND2X2 AND2X2_3476 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_72_), .Y(u2__abc_52155_new_n9024_));
AND2X2 AND2X2_3477 ( .A(u2__abc_52155_new_n8953_), .B(u2__abc_52155_new_n4128_), .Y(u2__abc_52155_new_n9025_));
AND2X2 AND2X2_3478 ( .A(u2__abc_52155_new_n9028_), .B(u2__abc_52155_new_n4147_), .Y(u2__abc_52155_new_n9029_));
AND2X2 AND2X2_3479 ( .A(u2__abc_52155_new_n9027_), .B(u2__abc_52155_new_n9029_), .Y(u2__abc_52155_new_n9030_));
AND2X2 AND2X2_348 ( .A(_abc_73687_new_n1593_), .B(_abc_73687_new_n1604_), .Y(_abc_73687_new_n1605_));
AND2X2 AND2X2_3480 ( .A(u2__abc_52155_new_n9032_), .B(u2__abc_52155_new_n4152_), .Y(u2__abc_52155_new_n9033_));
AND2X2 AND2X2_3481 ( .A(u2__abc_52155_new_n9031_), .B(u2__abc_52155_new_n9033_), .Y(u2__abc_52155_new_n9034_));
AND2X2 AND2X2_3482 ( .A(u2__abc_52155_new_n9026_), .B(u2__abc_52155_new_n9034_), .Y(u2__abc_52155_new_n9035_));
AND2X2 AND2X2_3483 ( .A(u2__abc_52155_new_n8878_), .B(u2__abc_52155_new_n4129_), .Y(u2__abc_52155_new_n9037_));
AND2X2 AND2X2_3484 ( .A(u2__abc_52155_new_n9038_), .B(u2__abc_52155_new_n4025_), .Y(u2__abc_52155_new_n9040_));
AND2X2 AND2X2_3485 ( .A(u2__abc_52155_new_n9041_), .B(u2__abc_52155_new_n9039_), .Y(u2__abc_52155_new_n9042_));
AND2X2 AND2X2_3486 ( .A(u2__abc_52155_new_n9043_), .B(u2__abc_52155_new_n9044_), .Y(u2__abc_52155_new_n9045_));
AND2X2 AND2X2_3487 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n4036_), .Y(u2__abc_52155_new_n9047_));
AND2X2 AND2X2_3488 ( .A(u2__abc_52155_new_n9048_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9049_));
AND2X2 AND2X2_3489 ( .A(u2__abc_52155_new_n9046_), .B(u2__abc_52155_new_n9049_), .Y(u2__abc_52155_new_n9050_));
AND2X2 AND2X2_349 ( .A(_abc_73687_new_n1606_), .B(_abc_73687_new_n1607_), .Y(_abc_73687_new_n1608_));
AND2X2 AND2X2_3490 ( .A(u2__abc_52155_new_n9051_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__72_));
AND2X2 AND2X2_3491 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_73_), .Y(u2__abc_52155_new_n9053_));
AND2X2 AND2X2_3492 ( .A(u2__abc_52155_new_n9041_), .B(u2__abc_52155_new_n4021_), .Y(u2__abc_52155_new_n9055_));
AND2X2 AND2X2_3493 ( .A(u2__abc_52155_new_n9058_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9059_));
AND2X2 AND2X2_3494 ( .A(u2__abc_52155_new_n9059_), .B(u2__abc_52155_new_n9056_), .Y(u2__abc_52155_new_n9060_));
AND2X2 AND2X2_3495 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_71_), .Y(u2__abc_52155_new_n9061_));
AND2X2 AND2X2_3496 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4041_), .Y(u2__abc_52155_new_n9064_));
AND2X2 AND2X2_3497 ( .A(u2__abc_52155_new_n9065_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9066_));
AND2X2 AND2X2_3498 ( .A(u2__abc_52155_new_n9063_), .B(u2__abc_52155_new_n9066_), .Y(u2__abc_52155_new_n9067_));
AND2X2 AND2X2_3499 ( .A(u2__abc_52155_new_n9068_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__73_));
AND2X2 AND2X2_35 ( .A(_abc_73687_new_n753_), .B(sqrto_34_), .Y(\o[70] ));
AND2X2 AND2X2_350 ( .A(_abc_73687_new_n1609_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1610_));
AND2X2 AND2X2_3500 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_74_), .Y(u2__abc_52155_new_n9070_));
AND2X2 AND2X2_3501 ( .A(u2__abc_52155_new_n9072_), .B(u2__abc_52155_new_n4028_), .Y(u2__abc_52155_new_n9073_));
AND2X2 AND2X2_3502 ( .A(u2__abc_52155_new_n9038_), .B(u2__abc_52155_new_n4033_), .Y(u2__abc_52155_new_n9075_));
AND2X2 AND2X2_3503 ( .A(u2__abc_52155_new_n9076_), .B(u2__abc_52155_new_n9071_), .Y(u2__abc_52155_new_n9077_));
AND2X2 AND2X2_3504 ( .A(u2__abc_52155_new_n9078_), .B(u2__abc_52155_new_n9079_), .Y(u2__abc_52155_new_n9080_));
AND2X2 AND2X2_3505 ( .A(u2__abc_52155_new_n9080_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9081_));
AND2X2 AND2X2_3506 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_72_), .Y(u2__abc_52155_new_n9082_));
AND2X2 AND2X2_3507 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4072_), .Y(u2__abc_52155_new_n9085_));
AND2X2 AND2X2_3508 ( .A(u2__abc_52155_new_n9086_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9087_));
AND2X2 AND2X2_3509 ( .A(u2__abc_52155_new_n9084_), .B(u2__abc_52155_new_n9087_), .Y(u2__abc_52155_new_n9088_));
AND2X2 AND2X2_351 ( .A(aNan), .B(\a[120] ), .Y(_abc_73687_new_n1611_));
AND2X2 AND2X2_3510 ( .A(u2__abc_52155_new_n9089_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__74_));
AND2X2 AND2X2_3511 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_75_), .Y(u2__abc_52155_new_n9091_));
AND2X2 AND2X2_3512 ( .A(u2__abc_52155_new_n9078_), .B(u2__abc_52155_new_n9092_), .Y(u2__abc_52155_new_n9093_));
AND2X2 AND2X2_3513 ( .A(u2__abc_52155_new_n9097_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9098_));
AND2X2 AND2X2_3514 ( .A(u2__abc_52155_new_n9098_), .B(u2__abc_52155_new_n9094_), .Y(u2__abc_52155_new_n9099_));
AND2X2 AND2X2_3515 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_73_), .Y(u2__abc_52155_new_n9100_));
AND2X2 AND2X2_3516 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4065_), .Y(u2__abc_52155_new_n9103_));
AND2X2 AND2X2_3517 ( .A(u2__abc_52155_new_n9104_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9105_));
AND2X2 AND2X2_3518 ( .A(u2__abc_52155_new_n9102_), .B(u2__abc_52155_new_n9105_), .Y(u2__abc_52155_new_n9106_));
AND2X2 AND2X2_3519 ( .A(u2__abc_52155_new_n9107_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__75_));
AND2X2 AND2X2_352 ( .A(aNan), .B(\a[121] ), .Y(_abc_73687_new_n1613_));
AND2X2 AND2X2_3520 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_76_), .Y(u2__abc_52155_new_n9109_));
AND2X2 AND2X2_3521 ( .A(u2__abc_52155_new_n9074_), .B(u2__abc_52155_new_n4045_), .Y(u2__abc_52155_new_n9110_));
AND2X2 AND2X2_3522 ( .A(u2__abc_52155_new_n9112_), .B(u2__abc_52155_new_n4163_), .Y(u2__abc_52155_new_n9113_));
AND2X2 AND2X2_3523 ( .A(u2__abc_52155_new_n9111_), .B(u2__abc_52155_new_n9113_), .Y(u2__abc_52155_new_n9114_));
AND2X2 AND2X2_3524 ( .A(u2__abc_52155_new_n9038_), .B(u2__abc_52155_new_n4046_), .Y(u2__abc_52155_new_n9116_));
AND2X2 AND2X2_3525 ( .A(u2__abc_52155_new_n9117_), .B(u2__abc_52155_new_n4075_), .Y(u2__abc_52155_new_n9118_));
AND2X2 AND2X2_3526 ( .A(u2__abc_52155_new_n9119_), .B(u2__abc_52155_new_n9120_), .Y(u2__abc_52155_new_n9121_));
AND2X2 AND2X2_3527 ( .A(u2__abc_52155_new_n9121_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9122_));
AND2X2 AND2X2_3528 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_74_), .Y(u2__abc_52155_new_n9123_));
AND2X2 AND2X2_3529 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4050_), .Y(u2__abc_52155_new_n9126_));
AND2X2 AND2X2_353 ( .A(_abc_73687_new_n1600_), .B(\a[122] ), .Y(_abc_73687_new_n1614_));
AND2X2 AND2X2_3530 ( .A(u2__abc_52155_new_n9127_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9128_));
AND2X2 AND2X2_3531 ( .A(u2__abc_52155_new_n9125_), .B(u2__abc_52155_new_n9128_), .Y(u2__abc_52155_new_n9129_));
AND2X2 AND2X2_3532 ( .A(u2__abc_52155_new_n9130_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__76_));
AND2X2 AND2X2_3533 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_77_), .Y(u2__abc_52155_new_n9132_));
AND2X2 AND2X2_3534 ( .A(u2__abc_52155_new_n9119_), .B(u2__abc_52155_new_n4071_), .Y(u2__abc_52155_new_n9133_));
AND2X2 AND2X2_3535 ( .A(u2__abc_52155_new_n9134_), .B(u2__abc_52155_new_n4068_), .Y(u2__abc_52155_new_n9135_));
AND2X2 AND2X2_3536 ( .A(u2__abc_52155_new_n9137_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9138_));
AND2X2 AND2X2_3537 ( .A(u2__abc_52155_new_n9138_), .B(u2__abc_52155_new_n9136_), .Y(u2__abc_52155_new_n9139_));
AND2X2 AND2X2_3538 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_75_), .Y(u2__abc_52155_new_n9140_));
AND2X2 AND2X2_3539 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4057_), .Y(u2__abc_52155_new_n9143_));
AND2X2 AND2X2_354 ( .A(_abc_73687_new_n1616_), .B(_abc_73687_new_n1615_), .Y(_abc_73687_new_n1617_));
AND2X2 AND2X2_3540 ( .A(u2__abc_52155_new_n9144_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9145_));
AND2X2 AND2X2_3541 ( .A(u2__abc_52155_new_n9142_), .B(u2__abc_52155_new_n9145_), .Y(u2__abc_52155_new_n9146_));
AND2X2 AND2X2_3542 ( .A(u2__abc_52155_new_n9147_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__77_));
AND2X2 AND2X2_3543 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_78_), .Y(u2__abc_52155_new_n9149_));
AND2X2 AND2X2_3544 ( .A(u2__abc_52155_new_n9136_), .B(u2__abc_52155_new_n4064_), .Y(u2__abc_52155_new_n9150_));
AND2X2 AND2X2_3545 ( .A(u2__abc_52155_new_n9151_), .B(u2__abc_52155_new_n4053_), .Y(u2__abc_52155_new_n9152_));
AND2X2 AND2X2_3546 ( .A(u2__abc_52155_new_n9154_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9155_));
AND2X2 AND2X2_3547 ( .A(u2__abc_52155_new_n9155_), .B(u2__abc_52155_new_n9153_), .Y(u2__abc_52155_new_n9156_));
AND2X2 AND2X2_3548 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_76_), .Y(u2__abc_52155_new_n9157_));
AND2X2 AND2X2_3549 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3961_), .Y(u2__abc_52155_new_n9160_));
AND2X2 AND2X2_355 ( .A(_abc_73687_new_n1605_), .B(_abc_73687_new_n1618_), .Y(_abc_73687_new_n1619_));
AND2X2 AND2X2_3550 ( .A(u2__abc_52155_new_n9161_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9162_));
AND2X2 AND2X2_3551 ( .A(u2__abc_52155_new_n9159_), .B(u2__abc_52155_new_n9162_), .Y(u2__abc_52155_new_n9163_));
AND2X2 AND2X2_3552 ( .A(u2__abc_52155_new_n9164_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__78_));
AND2X2 AND2X2_3553 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_79_), .Y(u2__abc_52155_new_n9166_));
AND2X2 AND2X2_3554 ( .A(u2__abc_52155_new_n9153_), .B(u2__abc_52155_new_n4049_), .Y(u2__abc_52155_new_n9168_));
AND2X2 AND2X2_3555 ( .A(u2__abc_52155_new_n9171_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9172_));
AND2X2 AND2X2_3556 ( .A(u2__abc_52155_new_n9172_), .B(u2__abc_52155_new_n9169_), .Y(u2__abc_52155_new_n9173_));
AND2X2 AND2X2_3557 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_77_), .Y(u2__abc_52155_new_n9174_));
AND2X2 AND2X2_3558 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3968_), .Y(u2__abc_52155_new_n9177_));
AND2X2 AND2X2_3559 ( .A(u2__abc_52155_new_n9178_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9179_));
AND2X2 AND2X2_356 ( .A(_abc_73687_new_n1620_), .B(_abc_73687_new_n1621_), .Y(_abc_73687_new_n1622_));
AND2X2 AND2X2_3560 ( .A(u2__abc_52155_new_n9176_), .B(u2__abc_52155_new_n9179_), .Y(u2__abc_52155_new_n9180_));
AND2X2 AND2X2_3561 ( .A(u2__abc_52155_new_n9181_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__79_));
AND2X2 AND2X2_3562 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_80_), .Y(u2__abc_52155_new_n9183_));
AND2X2 AND2X2_3563 ( .A(u2__abc_52155_new_n9036_), .B(u2__abc_52155_new_n4078_), .Y(u2__abc_52155_new_n9184_));
AND2X2 AND2X2_3564 ( .A(u2__abc_52155_new_n9115_), .B(u2__abc_52155_new_n4077_), .Y(u2__abc_52155_new_n9185_));
AND2X2 AND2X2_3565 ( .A(u2__abc_52155_new_n4059_), .B(u2__abc_52155_new_n4048_), .Y(u2__abc_52155_new_n9186_));
AND2X2 AND2X2_3566 ( .A(u2__abc_52155_new_n9188_), .B(u2__abc_52155_new_n4067_), .Y(u2__abc_52155_new_n9189_));
AND2X2 AND2X2_3567 ( .A(u2__abc_52155_new_n4061_), .B(u2__abc_52155_new_n9189_), .Y(u2__abc_52155_new_n9190_));
AND2X2 AND2X2_3568 ( .A(u2__abc_52155_new_n8878_), .B(u2__abc_52155_new_n4130_), .Y(u2__abc_52155_new_n9194_));
AND2X2 AND2X2_3569 ( .A(u2__abc_52155_new_n9195_), .B(u2__abc_52155_new_n3964_), .Y(u2__abc_52155_new_n9197_));
AND2X2 AND2X2_357 ( .A(_abc_73687_new_n1623_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1624_));
AND2X2 AND2X2_3570 ( .A(u2__abc_52155_new_n9198_), .B(u2__abc_52155_new_n9196_), .Y(u2__abc_52155_new_n9199_));
AND2X2 AND2X2_3571 ( .A(u2__abc_52155_new_n9200_), .B(u2__abc_52155_new_n9201_), .Y(u2__abc_52155_new_n9202_));
AND2X2 AND2X2_3572 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3975_), .Y(u2__abc_52155_new_n9204_));
AND2X2 AND2X2_3573 ( .A(u2__abc_52155_new_n9205_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9206_));
AND2X2 AND2X2_3574 ( .A(u2__abc_52155_new_n9203_), .B(u2__abc_52155_new_n9206_), .Y(u2__abc_52155_new_n9207_));
AND2X2 AND2X2_3575 ( .A(u2__abc_52155_new_n9208_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__80_));
AND2X2 AND2X2_3576 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_81_), .Y(u2__abc_52155_new_n9210_));
AND2X2 AND2X2_3577 ( .A(u2__abc_52155_new_n9198_), .B(u2__abc_52155_new_n3960_), .Y(u2__abc_52155_new_n9212_));
AND2X2 AND2X2_3578 ( .A(u2__abc_52155_new_n9215_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9216_));
AND2X2 AND2X2_3579 ( .A(u2__abc_52155_new_n9216_), .B(u2__abc_52155_new_n9213_), .Y(u2__abc_52155_new_n9217_));
AND2X2 AND2X2_358 ( .A(\a[120] ), .B(\a[121] ), .Y(_abc_73687_new_n1628_));
AND2X2 AND2X2_3580 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_79_), .Y(u2__abc_52155_new_n9218_));
AND2X2 AND2X2_3581 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3980_), .Y(u2__abc_52155_new_n9221_));
AND2X2 AND2X2_3582 ( .A(u2__abc_52155_new_n9222_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9223_));
AND2X2 AND2X2_3583 ( .A(u2__abc_52155_new_n9220_), .B(u2__abc_52155_new_n9223_), .Y(u2__abc_52155_new_n9224_));
AND2X2 AND2X2_3584 ( .A(u2__abc_52155_new_n9225_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__81_));
AND2X2 AND2X2_3585 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_82_), .Y(u2__abc_52155_new_n9227_));
AND2X2 AND2X2_3586 ( .A(u2__abc_52155_new_n9229_), .B(u2__abc_52155_new_n3967_), .Y(u2__abc_52155_new_n9230_));
AND2X2 AND2X2_3587 ( .A(u2__abc_52155_new_n9195_), .B(u2__abc_52155_new_n3972_), .Y(u2__abc_52155_new_n9232_));
AND2X2 AND2X2_3588 ( .A(u2__abc_52155_new_n9233_), .B(u2__abc_52155_new_n9228_), .Y(u2__abc_52155_new_n9234_));
AND2X2 AND2X2_3589 ( .A(u2__abc_52155_new_n9235_), .B(u2__abc_52155_new_n9236_), .Y(u2__abc_52155_new_n9237_));
AND2X2 AND2X2_359 ( .A(_abc_73687_new_n1578_), .B(_abc_73687_new_n1628_), .Y(_abc_73687_new_n1629_));
AND2X2 AND2X2_3590 ( .A(u2__abc_52155_new_n9237_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9238_));
AND2X2 AND2X2_3591 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_80_), .Y(u2__abc_52155_new_n9239_));
AND2X2 AND2X2_3592 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4011_), .Y(u2__abc_52155_new_n9242_));
AND2X2 AND2X2_3593 ( .A(u2__abc_52155_new_n9243_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9244_));
AND2X2 AND2X2_3594 ( .A(u2__abc_52155_new_n9241_), .B(u2__abc_52155_new_n9244_), .Y(u2__abc_52155_new_n9245_));
AND2X2 AND2X2_3595 ( .A(u2__abc_52155_new_n9246_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__82_));
AND2X2 AND2X2_3596 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_83_), .Y(u2__abc_52155_new_n9248_));
AND2X2 AND2X2_3597 ( .A(u2__abc_52155_new_n9235_), .B(u2__abc_52155_new_n9249_), .Y(u2__abc_52155_new_n9250_));
AND2X2 AND2X2_3598 ( .A(u2__abc_52155_new_n9254_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9255_));
AND2X2 AND2X2_3599 ( .A(u2__abc_52155_new_n9255_), .B(u2__abc_52155_new_n9251_), .Y(u2__abc_52155_new_n9256_));
AND2X2 AND2X2_36 ( .A(_abc_73687_new_n753_), .B(sqrto_35_), .Y(\o[71] ));
AND2X2 AND2X2_360 ( .A(_abc_73687_new_n1629_), .B(\a[122] ), .Y(_abc_73687_new_n1630_));
AND2X2 AND2X2_3600 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_81_), .Y(u2__abc_52155_new_n9257_));
AND2X2 AND2X2_3601 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4004_), .Y(u2__abc_52155_new_n9260_));
AND2X2 AND2X2_3602 ( .A(u2__abc_52155_new_n9261_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9262_));
AND2X2 AND2X2_3603 ( .A(u2__abc_52155_new_n9259_), .B(u2__abc_52155_new_n9262_), .Y(u2__abc_52155_new_n9263_));
AND2X2 AND2X2_3604 ( .A(u2__abc_52155_new_n9264_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__83_));
AND2X2 AND2X2_3605 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_84_), .Y(u2__abc_52155_new_n9266_));
AND2X2 AND2X2_3606 ( .A(u2__abc_52155_new_n9231_), .B(u2__abc_52155_new_n3984_), .Y(u2__abc_52155_new_n9267_));
AND2X2 AND2X2_3607 ( .A(u2__abc_52155_new_n9269_), .B(u2__abc_52155_new_n4184_), .Y(u2__abc_52155_new_n9270_));
AND2X2 AND2X2_3608 ( .A(u2__abc_52155_new_n9268_), .B(u2__abc_52155_new_n9270_), .Y(u2__abc_52155_new_n9271_));
AND2X2 AND2X2_3609 ( .A(u2__abc_52155_new_n9195_), .B(u2__abc_52155_new_n3985_), .Y(u2__abc_52155_new_n9273_));
AND2X2 AND2X2_361 ( .A(_abc_73687_new_n1631_), .B(_abc_73687_new_n1627_), .Y(_abc_73687_new_n1632_));
AND2X2 AND2X2_3610 ( .A(u2__abc_52155_new_n9274_), .B(u2__abc_52155_new_n4014_), .Y(u2__abc_52155_new_n9275_));
AND2X2 AND2X2_3611 ( .A(u2__abc_52155_new_n9276_), .B(u2__abc_52155_new_n9277_), .Y(u2__abc_52155_new_n9278_));
AND2X2 AND2X2_3612 ( .A(u2__abc_52155_new_n9278_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9279_));
AND2X2 AND2X2_3613 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_82_), .Y(u2__abc_52155_new_n9280_));
AND2X2 AND2X2_3614 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3989_), .Y(u2__abc_52155_new_n9283_));
AND2X2 AND2X2_3615 ( .A(u2__abc_52155_new_n9284_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9285_));
AND2X2 AND2X2_3616 ( .A(u2__abc_52155_new_n9282_), .B(u2__abc_52155_new_n9285_), .Y(u2__abc_52155_new_n9286_));
AND2X2 AND2X2_3617 ( .A(u2__abc_52155_new_n9287_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__84_));
AND2X2 AND2X2_3618 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_85_), .Y(u2__abc_52155_new_n9289_));
AND2X2 AND2X2_3619 ( .A(u2__abc_52155_new_n9276_), .B(u2__abc_52155_new_n4010_), .Y(u2__abc_52155_new_n9290_));
AND2X2 AND2X2_362 ( .A(_abc_73687_new_n1630_), .B(\a[123] ), .Y(_abc_73687_new_n1633_));
AND2X2 AND2X2_3620 ( .A(u2__abc_52155_new_n9290_), .B(u2__abc_52155_new_n4007_), .Y(u2__abc_52155_new_n9291_));
AND2X2 AND2X2_3621 ( .A(u2__abc_52155_new_n9293_), .B(u2__abc_52155_new_n9292_), .Y(u2__abc_52155_new_n9294_));
AND2X2 AND2X2_3622 ( .A(u2__abc_52155_new_n9295_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9296_));
AND2X2 AND2X2_3623 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_83_), .Y(u2__abc_52155_new_n9297_));
AND2X2 AND2X2_3624 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3996_), .Y(u2__abc_52155_new_n9300_));
AND2X2 AND2X2_3625 ( .A(u2__abc_52155_new_n9301_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9302_));
AND2X2 AND2X2_3626 ( .A(u2__abc_52155_new_n9299_), .B(u2__abc_52155_new_n9302_), .Y(u2__abc_52155_new_n9303_));
AND2X2 AND2X2_3627 ( .A(u2__abc_52155_new_n9304_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__85_));
AND2X2 AND2X2_3628 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_86_), .Y(u2__abc_52155_new_n9306_));
AND2X2 AND2X2_3629 ( .A(u2__abc_52155_new_n4003_), .B(u2__abc_52155_new_n4010_), .Y(u2__abc_52155_new_n9307_));
AND2X2 AND2X2_363 ( .A(_abc_73687_new_n1626_), .B(_abc_73687_new_n1635_), .Y(_abc_73687_new_n1636_));
AND2X2 AND2X2_3630 ( .A(u2__abc_52155_new_n9276_), .B(u2__abc_52155_new_n9307_), .Y(u2__abc_52155_new_n9308_));
AND2X2 AND2X2_3631 ( .A(u2__abc_52155_new_n9310_), .B(u2__abc_52155_new_n3992_), .Y(u2__abc_52155_new_n9311_));
AND2X2 AND2X2_3632 ( .A(u2__abc_52155_new_n9313_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9314_));
AND2X2 AND2X2_3633 ( .A(u2__abc_52155_new_n9314_), .B(u2__abc_52155_new_n9312_), .Y(u2__abc_52155_new_n9315_));
AND2X2 AND2X2_3634 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_84_), .Y(u2__abc_52155_new_n9316_));
AND2X2 AND2X2_3635 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3951_), .Y(u2__abc_52155_new_n9319_));
AND2X2 AND2X2_3636 ( .A(u2__abc_52155_new_n9320_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9321_));
AND2X2 AND2X2_3637 ( .A(u2__abc_52155_new_n9318_), .B(u2__abc_52155_new_n9321_), .Y(u2__abc_52155_new_n9322_));
AND2X2 AND2X2_3638 ( .A(u2__abc_52155_new_n9323_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__86_));
AND2X2 AND2X2_3639 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_87_), .Y(u2__abc_52155_new_n9325_));
AND2X2 AND2X2_364 ( .A(_abc_73687_new_n1619_), .B(_abc_73687_new_n1634_), .Y(_abc_73687_new_n1637_));
AND2X2 AND2X2_3640 ( .A(u2__abc_52155_new_n9312_), .B(u2__abc_52155_new_n3988_), .Y(u2__abc_52155_new_n9327_));
AND2X2 AND2X2_3641 ( .A(u2__abc_52155_new_n9330_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9331_));
AND2X2 AND2X2_3642 ( .A(u2__abc_52155_new_n9331_), .B(u2__abc_52155_new_n9328_), .Y(u2__abc_52155_new_n9332_));
AND2X2 AND2X2_3643 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_85_), .Y(u2__abc_52155_new_n9333_));
AND2X2 AND2X2_3644 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3944_), .Y(u2__abc_52155_new_n9336_));
AND2X2 AND2X2_3645 ( .A(u2__abc_52155_new_n9337_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9338_));
AND2X2 AND2X2_3646 ( .A(u2__abc_52155_new_n9335_), .B(u2__abc_52155_new_n9338_), .Y(u2__abc_52155_new_n9339_));
AND2X2 AND2X2_3647 ( .A(u2__abc_52155_new_n9340_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__87_));
AND2X2 AND2X2_3648 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_88_), .Y(u2__abc_52155_new_n9342_));
AND2X2 AND2X2_3649 ( .A(u2__abc_52155_new_n9272_), .B(u2__abc_52155_new_n4016_), .Y(u2__abc_52155_new_n9343_));
AND2X2 AND2X2_365 ( .A(_abc_73687_new_n1638_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1639_));
AND2X2 AND2X2_3650 ( .A(u2__abc_52155_new_n3988_), .B(u2__abc_52155_new_n3995_), .Y(u2__abc_52155_new_n9345_));
AND2X2 AND2X2_3651 ( .A(u2__abc_52155_new_n9348_), .B(u2__abc_52155_new_n4000_), .Y(u2__abc_52155_new_n9349_));
AND2X2 AND2X2_3652 ( .A(u2__abc_52155_new_n9350_), .B(u2__abc_52155_new_n9346_), .Y(u2__abc_52155_new_n9351_));
AND2X2 AND2X2_3653 ( .A(u2__abc_52155_new_n9344_), .B(u2__abc_52155_new_n9351_), .Y(u2__abc_52155_new_n9352_));
AND2X2 AND2X2_3654 ( .A(u2__abc_52155_new_n9195_), .B(u2__abc_52155_new_n4017_), .Y(u2__abc_52155_new_n9354_));
AND2X2 AND2X2_3655 ( .A(u2__abc_52155_new_n9355_), .B(u2__abc_52155_new_n3954_), .Y(u2__abc_52155_new_n9356_));
AND2X2 AND2X2_3656 ( .A(u2__abc_52155_new_n9357_), .B(u2__abc_52155_new_n9358_), .Y(u2__abc_52155_new_n9359_));
AND2X2 AND2X2_3657 ( .A(u2__abc_52155_new_n9359_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9360_));
AND2X2 AND2X2_3658 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_86_), .Y(u2__abc_52155_new_n9361_));
AND2X2 AND2X2_3659 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3929_), .Y(u2__abc_52155_new_n9364_));
AND2X2 AND2X2_366 ( .A(aNan), .B(\a[122] ), .Y(_abc_73687_new_n1640_));
AND2X2 AND2X2_3660 ( .A(u2__abc_52155_new_n9365_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9366_));
AND2X2 AND2X2_3661 ( .A(u2__abc_52155_new_n9363_), .B(u2__abc_52155_new_n9366_), .Y(u2__abc_52155_new_n9367_));
AND2X2 AND2X2_3662 ( .A(u2__abc_52155_new_n9368_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__88_));
AND2X2 AND2X2_3663 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_89_), .Y(u2__abc_52155_new_n9370_));
AND2X2 AND2X2_3664 ( .A(u2__abc_52155_new_n9357_), .B(u2__abc_52155_new_n3950_), .Y(u2__abc_52155_new_n9371_));
AND2X2 AND2X2_3665 ( .A(u2__abc_52155_new_n9375_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9376_));
AND2X2 AND2X2_3666 ( .A(u2__abc_52155_new_n9376_), .B(u2__abc_52155_new_n9373_), .Y(u2__abc_52155_new_n9377_));
AND2X2 AND2X2_3667 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_87_), .Y(u2__abc_52155_new_n9378_));
AND2X2 AND2X2_3668 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3936_), .Y(u2__abc_52155_new_n9381_));
AND2X2 AND2X2_3669 ( .A(u2__abc_52155_new_n9382_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9383_));
AND2X2 AND2X2_367 ( .A(aNan), .B(\a[123] ), .Y(_abc_73687_new_n1642_));
AND2X2 AND2X2_3670 ( .A(u2__abc_52155_new_n9380_), .B(u2__abc_52155_new_n9383_), .Y(u2__abc_52155_new_n9384_));
AND2X2 AND2X2_3671 ( .A(u2__abc_52155_new_n9385_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__89_));
AND2X2 AND2X2_3672 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_90_), .Y(u2__abc_52155_new_n9387_));
AND2X2 AND2X2_3673 ( .A(u2__abc_52155_new_n3943_), .B(u2__abc_52155_new_n3950_), .Y(u2__abc_52155_new_n9388_));
AND2X2 AND2X2_3674 ( .A(u2__abc_52155_new_n9355_), .B(u2__abc_52155_new_n3955_), .Y(u2__abc_52155_new_n9391_));
AND2X2 AND2X2_3675 ( .A(u2__abc_52155_new_n9392_), .B(u2__abc_52155_new_n3932_), .Y(u2__abc_52155_new_n9393_));
AND2X2 AND2X2_3676 ( .A(u2__abc_52155_new_n9395_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9396_));
AND2X2 AND2X2_3677 ( .A(u2__abc_52155_new_n9396_), .B(u2__abc_52155_new_n9394_), .Y(u2__abc_52155_new_n9397_));
AND2X2 AND2X2_3678 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_88_), .Y(u2__abc_52155_new_n9398_));
AND2X2 AND2X2_3679 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3920_), .Y(u2__abc_52155_new_n9401_));
AND2X2 AND2X2_368 ( .A(_abc_73687_new_n1633_), .B(_abc_73687_new_n1643_), .Y(_abc_73687_new_n1644_));
AND2X2 AND2X2_3680 ( .A(u2__abc_52155_new_n9402_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9403_));
AND2X2 AND2X2_3681 ( .A(u2__abc_52155_new_n9400_), .B(u2__abc_52155_new_n9403_), .Y(u2__abc_52155_new_n9404_));
AND2X2 AND2X2_3682 ( .A(u2__abc_52155_new_n9405_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__90_));
AND2X2 AND2X2_3683 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_91_), .Y(u2__abc_52155_new_n9407_));
AND2X2 AND2X2_3684 ( .A(u2__abc_52155_new_n9394_), .B(u2__abc_52155_new_n3928_), .Y(u2__abc_52155_new_n9409_));
AND2X2 AND2X2_3685 ( .A(u2__abc_52155_new_n9412_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9413_));
AND2X2 AND2X2_3686 ( .A(u2__abc_52155_new_n9413_), .B(u2__abc_52155_new_n9410_), .Y(u2__abc_52155_new_n9414_));
AND2X2 AND2X2_3687 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_89_), .Y(u2__abc_52155_new_n9415_));
AND2X2 AND2X2_3688 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3913_), .Y(u2__abc_52155_new_n9418_));
AND2X2 AND2X2_3689 ( .A(u2__abc_52155_new_n9419_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9420_));
AND2X2 AND2X2_369 ( .A(_abc_73687_new_n1645_), .B(_abc_73687_new_n1646_), .Y(_abc_73687_new_n1647_));
AND2X2 AND2X2_3690 ( .A(u2__abc_52155_new_n9417_), .B(u2__abc_52155_new_n9420_), .Y(u2__abc_52155_new_n9421_));
AND2X2 AND2X2_3691 ( .A(u2__abc_52155_new_n9422_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__91_));
AND2X2 AND2X2_3692 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_92_), .Y(u2__abc_52155_new_n9424_));
AND2X2 AND2X2_3693 ( .A(u2__abc_52155_new_n3928_), .B(u2__abc_52155_new_n3935_), .Y(u2__abc_52155_new_n9425_));
AND2X2 AND2X2_3694 ( .A(u2__abc_52155_new_n9394_), .B(u2__abc_52155_new_n9425_), .Y(u2__abc_52155_new_n9426_));
AND2X2 AND2X2_3695 ( .A(u2__abc_52155_new_n9428_), .B(u2__abc_52155_new_n3923_), .Y(u2__abc_52155_new_n9429_));
AND2X2 AND2X2_3696 ( .A(u2__abc_52155_new_n9431_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9432_));
AND2X2 AND2X2_3697 ( .A(u2__abc_52155_new_n9432_), .B(u2__abc_52155_new_n9430_), .Y(u2__abc_52155_new_n9433_));
AND2X2 AND2X2_3698 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_90_), .Y(u2__abc_52155_new_n9434_));
AND2X2 AND2X2_3699 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3898_), .Y(u2__abc_52155_new_n9437_));
AND2X2 AND2X2_37 ( .A(_abc_73687_new_n753_), .B(sqrto_36_), .Y(\o[72] ));
AND2X2 AND2X2_370 ( .A(_abc_73687_new_n1637_), .B(_abc_73687_new_n1647_), .Y(_abc_73687_new_n1648_));
AND2X2 AND2X2_3700 ( .A(u2__abc_52155_new_n9438_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9439_));
AND2X2 AND2X2_3701 ( .A(u2__abc_52155_new_n9436_), .B(u2__abc_52155_new_n9439_), .Y(u2__abc_52155_new_n9440_));
AND2X2 AND2X2_3702 ( .A(u2__abc_52155_new_n9441_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__92_));
AND2X2 AND2X2_3703 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_93_), .Y(u2__abc_52155_new_n9443_));
AND2X2 AND2X2_3704 ( .A(u2__abc_52155_new_n9430_), .B(u2__abc_52155_new_n3919_), .Y(u2__abc_52155_new_n9444_));
AND2X2 AND2X2_3705 ( .A(u2__abc_52155_new_n9444_), .B(u2__abc_52155_new_n3916_), .Y(u2__abc_52155_new_n9445_));
AND2X2 AND2X2_3706 ( .A(u2__abc_52155_new_n9447_), .B(u2__abc_52155_new_n9446_), .Y(u2__abc_52155_new_n9448_));
AND2X2 AND2X2_3707 ( .A(u2__abc_52155_new_n9449_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9450_));
AND2X2 AND2X2_3708 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_91_), .Y(u2__abc_52155_new_n9451_));
AND2X2 AND2X2_3709 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3905_), .Y(u2__abc_52155_new_n9454_));
AND2X2 AND2X2_371 ( .A(_abc_73687_new_n1649_), .B(_abc_73687_new_n1650_), .Y(_abc_73687_new_n1651_));
AND2X2 AND2X2_3710 ( .A(u2__abc_52155_new_n9455_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9456_));
AND2X2 AND2X2_3711 ( .A(u2__abc_52155_new_n9453_), .B(u2__abc_52155_new_n9456_), .Y(u2__abc_52155_new_n9457_));
AND2X2 AND2X2_3712 ( .A(u2__abc_52155_new_n9458_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__93_));
AND2X2 AND2X2_3713 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_94_), .Y(u2__abc_52155_new_n9460_));
AND2X2 AND2X2_3714 ( .A(u2__abc_52155_new_n3912_), .B(u2__abc_52155_new_n3919_), .Y(u2__abc_52155_new_n9461_));
AND2X2 AND2X2_3715 ( .A(u2__abc_52155_new_n9430_), .B(u2__abc_52155_new_n9461_), .Y(u2__abc_52155_new_n9462_));
AND2X2 AND2X2_3716 ( .A(u2__abc_52155_new_n9464_), .B(u2__abc_52155_new_n3901_), .Y(u2__abc_52155_new_n9465_));
AND2X2 AND2X2_3717 ( .A(u2__abc_52155_new_n9467_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9468_));
AND2X2 AND2X2_3718 ( .A(u2__abc_52155_new_n9468_), .B(u2__abc_52155_new_n9466_), .Y(u2__abc_52155_new_n9469_));
AND2X2 AND2X2_3719 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_92_), .Y(u2__abc_52155_new_n9470_));
AND2X2 AND2X2_372 ( .A(_abc_73687_new_n1652_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1653_));
AND2X2 AND2X2_3720 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3855_), .Y(u2__abc_52155_new_n9473_));
AND2X2 AND2X2_3721 ( .A(u2__abc_52155_new_n9474_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9475_));
AND2X2 AND2X2_3722 ( .A(u2__abc_52155_new_n9472_), .B(u2__abc_52155_new_n9475_), .Y(u2__abc_52155_new_n9476_));
AND2X2 AND2X2_3723 ( .A(u2__abc_52155_new_n9477_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__94_));
AND2X2 AND2X2_3724 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_95_), .Y(u2__abc_52155_new_n9479_));
AND2X2 AND2X2_3725 ( .A(u2__abc_52155_new_n9466_), .B(u2__abc_52155_new_n3897_), .Y(u2__abc_52155_new_n9480_));
AND2X2 AND2X2_3726 ( .A(u2__abc_52155_new_n9480_), .B(u2__abc_52155_new_n3908_), .Y(u2__abc_52155_new_n9481_));
AND2X2 AND2X2_3727 ( .A(u2__abc_52155_new_n9483_), .B(u2__abc_52155_new_n9482_), .Y(u2__abc_52155_new_n9484_));
AND2X2 AND2X2_3728 ( .A(u2__abc_52155_new_n9485_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9486_));
AND2X2 AND2X2_3729 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_93_), .Y(u2__abc_52155_new_n9487_));
AND2X2 AND2X2_373 ( .A(_abc_73687_new_n1633_), .B(\a[124] ), .Y(_abc_73687_new_n1657_));
AND2X2 AND2X2_3730 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3848_), .Y(u2__abc_52155_new_n9490_));
AND2X2 AND2X2_3731 ( .A(u2__abc_52155_new_n9491_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9492_));
AND2X2 AND2X2_3732 ( .A(u2__abc_52155_new_n9489_), .B(u2__abc_52155_new_n9492_), .Y(u2__abc_52155_new_n9493_));
AND2X2 AND2X2_3733 ( .A(u2__abc_52155_new_n9494_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__95_));
AND2X2 AND2X2_3734 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_96_), .Y(u2__abc_52155_new_n9496_));
AND2X2 AND2X2_3735 ( .A(u2__abc_52155_new_n9193_), .B(u2__abc_52155_new_n4018_), .Y(u2__abc_52155_new_n9497_));
AND2X2 AND2X2_3736 ( .A(u2__abc_52155_new_n9353_), .B(u2__abc_52155_new_n3957_), .Y(u2__abc_52155_new_n9499_));
AND2X2 AND2X2_3737 ( .A(u2__abc_52155_new_n9390_), .B(u2__abc_52155_new_n3940_), .Y(u2__abc_52155_new_n9502_));
AND2X2 AND2X2_3738 ( .A(u2__abc_52155_new_n9503_), .B(u2__abc_52155_new_n9501_), .Y(u2__abc_52155_new_n9504_));
AND2X2 AND2X2_3739 ( .A(u2__abc_52155_new_n9505_), .B(u2__abc_52155_new_n3925_), .Y(u2__abc_52155_new_n9506_));
AND2X2 AND2X2_374 ( .A(_abc_73687_new_n1658_), .B(_abc_73687_new_n1656_), .Y(_abc_73687_new_n1659_));
AND2X2 AND2X2_3740 ( .A(u2__abc_52155_new_n9509_), .B(u2__abc_52155_new_n3909_), .Y(u2__abc_52155_new_n9510_));
AND2X2 AND2X2_3741 ( .A(u2__abc_52155_new_n3897_), .B(u2__abc_52155_new_n3904_), .Y(u2__abc_52155_new_n9512_));
AND2X2 AND2X2_3742 ( .A(u2__abc_52155_new_n9511_), .B(u2__abc_52155_new_n9513_), .Y(u2__abc_52155_new_n9514_));
AND2X2 AND2X2_3743 ( .A(u2__abc_52155_new_n9507_), .B(u2__abc_52155_new_n9514_), .Y(u2__abc_52155_new_n9515_));
AND2X2 AND2X2_3744 ( .A(u2__abc_52155_new_n9500_), .B(u2__abc_52155_new_n9515_), .Y(u2__abc_52155_new_n9516_));
AND2X2 AND2X2_3745 ( .A(u2__abc_52155_new_n9498_), .B(u2__abc_52155_new_n9516_), .Y(u2__abc_52155_new_n9517_));
AND2X2 AND2X2_3746 ( .A(u2__abc_52155_new_n8878_), .B(u2__abc_52155_new_n4131_), .Y(u2__abc_52155_new_n9519_));
AND2X2 AND2X2_3747 ( .A(u2__abc_52155_new_n9520_), .B(u2__abc_52155_new_n3858_), .Y(u2__abc_52155_new_n9522_));
AND2X2 AND2X2_3748 ( .A(u2__abc_52155_new_n9523_), .B(u2__abc_52155_new_n9521_), .Y(u2__abc_52155_new_n9524_));
AND2X2 AND2X2_3749 ( .A(u2__abc_52155_new_n9525_), .B(u2__abc_52155_new_n9526_), .Y(u2__abc_52155_new_n9527_));
AND2X2 AND2X2_375 ( .A(_abc_73687_new_n1657_), .B(\a[125] ), .Y(_abc_73687_new_n1660_));
AND2X2 AND2X2_3750 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n3835_), .Y(u2__abc_52155_new_n9529_));
AND2X2 AND2X2_3751 ( .A(u2__abc_52155_new_n9530_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9531_));
AND2X2 AND2X2_3752 ( .A(u2__abc_52155_new_n9528_), .B(u2__abc_52155_new_n9531_), .Y(u2__abc_52155_new_n9532_));
AND2X2 AND2X2_3753 ( .A(u2__abc_52155_new_n9533_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__96_));
AND2X2 AND2X2_3754 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_97_), .Y(u2__abc_52155_new_n9535_));
AND2X2 AND2X2_3755 ( .A(u2__abc_52155_new_n9523_), .B(u2__abc_52155_new_n3854_), .Y(u2__abc_52155_new_n9536_));
AND2X2 AND2X2_3756 ( .A(u2__abc_52155_new_n9536_), .B(u2__abc_52155_new_n3851_), .Y(u2__abc_52155_new_n9537_));
AND2X2 AND2X2_3757 ( .A(u2__abc_52155_new_n9539_), .B(u2__abc_52155_new_n9538_), .Y(u2__abc_52155_new_n9540_));
AND2X2 AND2X2_3758 ( .A(u2__abc_52155_new_n9541_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9542_));
AND2X2 AND2X2_3759 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_95_), .Y(u2__abc_52155_new_n9543_));
AND2X2 AND2X2_376 ( .A(_abc_73687_new_n1655_), .B(_abc_73687_new_n1662_), .Y(_abc_73687_new_n1663_));
AND2X2 AND2X2_3760 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3840_), .Y(u2__abc_52155_new_n9546_));
AND2X2 AND2X2_3761 ( .A(u2__abc_52155_new_n9547_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9548_));
AND2X2 AND2X2_3762 ( .A(u2__abc_52155_new_n9545_), .B(u2__abc_52155_new_n9548_), .Y(u2__abc_52155_new_n9549_));
AND2X2 AND2X2_3763 ( .A(u2__abc_52155_new_n9550_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__97_));
AND2X2 AND2X2_3764 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_98_), .Y(u2__abc_52155_new_n9552_));
AND2X2 AND2X2_3765 ( .A(u2__abc_52155_new_n3847_), .B(u2__abc_52155_new_n3854_), .Y(u2__abc_52155_new_n9554_));
AND2X2 AND2X2_3766 ( .A(u2__abc_52155_new_n9523_), .B(u2__abc_52155_new_n9554_), .Y(u2__abc_52155_new_n9555_));
AND2X2 AND2X2_3767 ( .A(u2__abc_52155_new_n9557_), .B(u2__abc_52155_new_n9553_), .Y(u2__abc_52155_new_n9558_));
AND2X2 AND2X2_3768 ( .A(u2__abc_52155_new_n9559_), .B(u2__abc_52155_new_n9560_), .Y(u2__abc_52155_new_n9561_));
AND2X2 AND2X2_3769 ( .A(u2__abc_52155_new_n9561_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9562_));
AND2X2 AND2X2_377 ( .A(_abc_73687_new_n1648_), .B(_abc_73687_new_n1661_), .Y(_abc_73687_new_n1664_));
AND2X2 AND2X2_3770 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_96_), .Y(u2__abc_52155_new_n9563_));
AND2X2 AND2X2_3771 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3886_), .Y(u2__abc_52155_new_n9566_));
AND2X2 AND2X2_3772 ( .A(u2__abc_52155_new_n9567_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9568_));
AND2X2 AND2X2_3773 ( .A(u2__abc_52155_new_n9565_), .B(u2__abc_52155_new_n9568_), .Y(u2__abc_52155_new_n9569_));
AND2X2 AND2X2_3774 ( .A(u2__abc_52155_new_n9570_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__98_));
AND2X2 AND2X2_3775 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_99_), .Y(u2__abc_52155_new_n9572_));
AND2X2 AND2X2_3776 ( .A(u2__abc_52155_new_n9559_), .B(u2__abc_52155_new_n9573_), .Y(u2__abc_52155_new_n9574_));
AND2X2 AND2X2_3777 ( .A(u2__abc_52155_new_n9578_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9579_));
AND2X2 AND2X2_3778 ( .A(u2__abc_52155_new_n9579_), .B(u2__abc_52155_new_n9575_), .Y(u2__abc_52155_new_n9580_));
AND2X2 AND2X2_3779 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_97_), .Y(u2__abc_52155_new_n9581_));
AND2X2 AND2X2_378 ( .A(_abc_73687_new_n1665_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1666_));
AND2X2 AND2X2_3780 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3879_), .Y(u2__abc_52155_new_n9584_));
AND2X2 AND2X2_3781 ( .A(u2__abc_52155_new_n9585_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9586_));
AND2X2 AND2X2_3782 ( .A(u2__abc_52155_new_n9583_), .B(u2__abc_52155_new_n9586_), .Y(u2__abc_52155_new_n9587_));
AND2X2 AND2X2_3783 ( .A(u2__abc_52155_new_n9588_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__99_));
AND2X2 AND2X2_3784 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_100_), .Y(u2__abc_52155_new_n9590_));
AND2X2 AND2X2_3785 ( .A(u2__abc_52155_new_n9593_), .B(u2__abc_52155_new_n4223_), .Y(u2__abc_52155_new_n9594_));
AND2X2 AND2X2_3786 ( .A(u2__abc_52155_new_n9592_), .B(u2__abc_52155_new_n9594_), .Y(u2__abc_52155_new_n9595_));
AND2X2 AND2X2_3787 ( .A(u2__abc_52155_new_n9520_), .B(u2__abc_52155_new_n3860_), .Y(u2__abc_52155_new_n9597_));
AND2X2 AND2X2_3788 ( .A(u2__abc_52155_new_n9598_), .B(u2__abc_52155_new_n3889_), .Y(u2__abc_52155_new_n9599_));
AND2X2 AND2X2_3789 ( .A(u2__abc_52155_new_n9600_), .B(u2__abc_52155_new_n9601_), .Y(u2__abc_52155_new_n9602_));
AND2X2 AND2X2_379 ( .A(aNan), .B(\a[124] ), .Y(_abc_73687_new_n1667_));
AND2X2 AND2X2_3790 ( .A(u2__abc_52155_new_n9602_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9603_));
AND2X2 AND2X2_3791 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_98_), .Y(u2__abc_52155_new_n9604_));
AND2X2 AND2X2_3792 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3864_), .Y(u2__abc_52155_new_n9607_));
AND2X2 AND2X2_3793 ( .A(u2__abc_52155_new_n9608_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9609_));
AND2X2 AND2X2_3794 ( .A(u2__abc_52155_new_n9606_), .B(u2__abc_52155_new_n9609_), .Y(u2__abc_52155_new_n9610_));
AND2X2 AND2X2_3795 ( .A(u2__abc_52155_new_n9611_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__100_));
AND2X2 AND2X2_3796 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_101_), .Y(u2__abc_52155_new_n9613_));
AND2X2 AND2X2_3797 ( .A(u2__abc_52155_new_n9600_), .B(u2__abc_52155_new_n3885_), .Y(u2__abc_52155_new_n9614_));
AND2X2 AND2X2_3798 ( .A(u2__abc_52155_new_n9614_), .B(u2__abc_52155_new_n3882_), .Y(u2__abc_52155_new_n9615_));
AND2X2 AND2X2_3799 ( .A(u2__abc_52155_new_n9617_), .B(u2__abc_52155_new_n9616_), .Y(u2__abc_52155_new_n9618_));
AND2X2 AND2X2_38 ( .A(_abc_73687_new_n753_), .B(sqrto_37_), .Y(\o[73] ));
AND2X2 AND2X2_380 ( .A(_abc_73687_new_n1660_), .B(_abc_73687_new_n1670_), .Y(_abc_73687_new_n1672_));
AND2X2 AND2X2_3800 ( .A(u2__abc_52155_new_n9619_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9620_));
AND2X2 AND2X2_3801 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_99_), .Y(u2__abc_52155_new_n9621_));
AND2X2 AND2X2_3802 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3871_), .Y(u2__abc_52155_new_n9624_));
AND2X2 AND2X2_3803 ( .A(u2__abc_52155_new_n9625_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9626_));
AND2X2 AND2X2_3804 ( .A(u2__abc_52155_new_n9623_), .B(u2__abc_52155_new_n9626_), .Y(u2__abc_52155_new_n9627_));
AND2X2 AND2X2_3805 ( .A(u2__abc_52155_new_n9628_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__101_));
AND2X2 AND2X2_3806 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_102_), .Y(u2__abc_52155_new_n9630_));
AND2X2 AND2X2_3807 ( .A(u2__abc_52155_new_n3878_), .B(u2__abc_52155_new_n3885_), .Y(u2__abc_52155_new_n9631_));
AND2X2 AND2X2_3808 ( .A(u2__abc_52155_new_n9600_), .B(u2__abc_52155_new_n9631_), .Y(u2__abc_52155_new_n9632_));
AND2X2 AND2X2_3809 ( .A(u2__abc_52155_new_n9634_), .B(u2__abc_52155_new_n3867_), .Y(u2__abc_52155_new_n9635_));
AND2X2 AND2X2_381 ( .A(_abc_73687_new_n1673_), .B(_abc_73687_new_n1671_), .Y(_abc_73687_new_n1674_));
AND2X2 AND2X2_3810 ( .A(u2__abc_52155_new_n9637_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9638_));
AND2X2 AND2X2_3811 ( .A(u2__abc_52155_new_n9638_), .B(u2__abc_52155_new_n9636_), .Y(u2__abc_52155_new_n9639_));
AND2X2 AND2X2_3812 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_100_), .Y(u2__abc_52155_new_n9640_));
AND2X2 AND2X2_3813 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3795_), .Y(u2__abc_52155_new_n9643_));
AND2X2 AND2X2_3814 ( .A(u2__abc_52155_new_n9644_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9645_));
AND2X2 AND2X2_3815 ( .A(u2__abc_52155_new_n9642_), .B(u2__abc_52155_new_n9645_), .Y(u2__abc_52155_new_n9646_));
AND2X2 AND2X2_3816 ( .A(u2__abc_52155_new_n9647_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__102_));
AND2X2 AND2X2_3817 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_103_), .Y(u2__abc_52155_new_n9649_));
AND2X2 AND2X2_3818 ( .A(u2__abc_52155_new_n9636_), .B(u2__abc_52155_new_n3863_), .Y(u2__abc_52155_new_n9651_));
AND2X2 AND2X2_3819 ( .A(u2__abc_52155_new_n9654_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9655_));
AND2X2 AND2X2_382 ( .A(_abc_73687_new_n1664_), .B(_abc_73687_new_n1674_), .Y(_abc_73687_new_n1676_));
AND2X2 AND2X2_3820 ( .A(u2__abc_52155_new_n9655_), .B(u2__abc_52155_new_n9652_), .Y(u2__abc_52155_new_n9656_));
AND2X2 AND2X2_3821 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_101_), .Y(u2__abc_52155_new_n9657_));
AND2X2 AND2X2_3822 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3788_), .Y(u2__abc_52155_new_n9660_));
AND2X2 AND2X2_3823 ( .A(u2__abc_52155_new_n9661_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9662_));
AND2X2 AND2X2_3824 ( .A(u2__abc_52155_new_n9659_), .B(u2__abc_52155_new_n9662_), .Y(u2__abc_52155_new_n9663_));
AND2X2 AND2X2_3825 ( .A(u2__abc_52155_new_n9664_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__103_));
AND2X2 AND2X2_3826 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_104_), .Y(u2__abc_52155_new_n9666_));
AND2X2 AND2X2_3827 ( .A(u2__abc_52155_new_n9596_), .B(u2__abc_52155_new_n3891_), .Y(u2__abc_52155_new_n9667_));
AND2X2 AND2X2_3828 ( .A(u2__abc_52155_new_n9669_), .B(u2__abc_52155_new_n3875_), .Y(u2__abc_52155_new_n9670_));
AND2X2 AND2X2_3829 ( .A(u2__abc_52155_new_n3873_), .B(u2__abc_52155_new_n3862_), .Y(u2__abc_52155_new_n9671_));
AND2X2 AND2X2_383 ( .A(_abc_73687_new_n1677_), .B(_abc_73687_new_n1675_), .Y(_abc_73687_new_n1678_));
AND2X2 AND2X2_3830 ( .A(u2__abc_52155_new_n9520_), .B(u2__abc_52155_new_n3892_), .Y(u2__abc_52155_new_n9675_));
AND2X2 AND2X2_3831 ( .A(u2__abc_52155_new_n9676_), .B(u2__abc_52155_new_n3798_), .Y(u2__abc_52155_new_n9677_));
AND2X2 AND2X2_3832 ( .A(u2__abc_52155_new_n9678_), .B(u2__abc_52155_new_n9679_), .Y(u2__abc_52155_new_n9680_));
AND2X2 AND2X2_3833 ( .A(u2__abc_52155_new_n9680_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9681_));
AND2X2 AND2X2_3834 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_102_), .Y(u2__abc_52155_new_n9682_));
AND2X2 AND2X2_3835 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3773_), .Y(u2__abc_52155_new_n9685_));
AND2X2 AND2X2_3836 ( .A(u2__abc_52155_new_n9686_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9687_));
AND2X2 AND2X2_3837 ( .A(u2__abc_52155_new_n9684_), .B(u2__abc_52155_new_n9687_), .Y(u2__abc_52155_new_n9688_));
AND2X2 AND2X2_3838 ( .A(u2__abc_52155_new_n9689_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__104_));
AND2X2 AND2X2_3839 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_105_), .Y(u2__abc_52155_new_n9691_));
AND2X2 AND2X2_384 ( .A(_abc_73687_new_n1679_), .B(_abc_73687_new_n1669_), .Y(\o[239] ));
AND2X2 AND2X2_3840 ( .A(u2__abc_52155_new_n9678_), .B(u2__abc_52155_new_n3794_), .Y(u2__abc_52155_new_n9692_));
AND2X2 AND2X2_3841 ( .A(u2__abc_52155_new_n9692_), .B(u2__abc_52155_new_n3791_), .Y(u2__abc_52155_new_n9693_));
AND2X2 AND2X2_3842 ( .A(u2__abc_52155_new_n9695_), .B(u2__abc_52155_new_n9694_), .Y(u2__abc_52155_new_n9696_));
AND2X2 AND2X2_3843 ( .A(u2__abc_52155_new_n9697_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9698_));
AND2X2 AND2X2_3844 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_103_), .Y(u2__abc_52155_new_n9699_));
AND2X2 AND2X2_3845 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3780_), .Y(u2__abc_52155_new_n9702_));
AND2X2 AND2X2_3846 ( .A(u2__abc_52155_new_n9703_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9704_));
AND2X2 AND2X2_3847 ( .A(u2__abc_52155_new_n9701_), .B(u2__abc_52155_new_n9704_), .Y(u2__abc_52155_new_n9705_));
AND2X2 AND2X2_3848 ( .A(u2__abc_52155_new_n9706_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__105_));
AND2X2 AND2X2_3849 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_106_), .Y(u2__abc_52155_new_n9708_));
AND2X2 AND2X2_385 ( .A(_abc_73687_new_n1614_), .B(\a[123] ), .Y(_abc_73687_new_n1681_));
AND2X2 AND2X2_3850 ( .A(u2__abc_52155_new_n3787_), .B(u2__abc_52155_new_n3794_), .Y(u2__abc_52155_new_n9709_));
AND2X2 AND2X2_3851 ( .A(u2__abc_52155_new_n9678_), .B(u2__abc_52155_new_n9709_), .Y(u2__abc_52155_new_n9710_));
AND2X2 AND2X2_3852 ( .A(u2__abc_52155_new_n9712_), .B(u2__abc_52155_new_n3776_), .Y(u2__abc_52155_new_n9713_));
AND2X2 AND2X2_3853 ( .A(u2__abc_52155_new_n9715_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9716_));
AND2X2 AND2X2_3854 ( .A(u2__abc_52155_new_n9716_), .B(u2__abc_52155_new_n9714_), .Y(u2__abc_52155_new_n9717_));
AND2X2 AND2X2_3855 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_104_), .Y(u2__abc_52155_new_n9718_));
AND2X2 AND2X2_3856 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3826_), .Y(u2__abc_52155_new_n9721_));
AND2X2 AND2X2_3857 ( .A(u2__abc_52155_new_n9722_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9723_));
AND2X2 AND2X2_3858 ( .A(u2__abc_52155_new_n9720_), .B(u2__abc_52155_new_n9723_), .Y(u2__abc_52155_new_n9724_));
AND2X2 AND2X2_3859 ( .A(u2__abc_52155_new_n9725_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__106_));
AND2X2 AND2X2_386 ( .A(_abc_73687_new_n1681_), .B(\a[124] ), .Y(_abc_73687_new_n1682_));
AND2X2 AND2X2_3860 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_107_), .Y(u2__abc_52155_new_n9727_));
AND2X2 AND2X2_3861 ( .A(u2__abc_52155_new_n9714_), .B(u2__abc_52155_new_n3772_), .Y(u2__abc_52155_new_n9729_));
AND2X2 AND2X2_3862 ( .A(u2__abc_52155_new_n9732_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9733_));
AND2X2 AND2X2_3863 ( .A(u2__abc_52155_new_n9733_), .B(u2__abc_52155_new_n9730_), .Y(u2__abc_52155_new_n9734_));
AND2X2 AND2X2_3864 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_105_), .Y(u2__abc_52155_new_n9735_));
AND2X2 AND2X2_3865 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3819_), .Y(u2__abc_52155_new_n9738_));
AND2X2 AND2X2_3866 ( .A(u2__abc_52155_new_n9739_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9740_));
AND2X2 AND2X2_3867 ( .A(u2__abc_52155_new_n9737_), .B(u2__abc_52155_new_n9740_), .Y(u2__abc_52155_new_n9741_));
AND2X2 AND2X2_3868 ( .A(u2__abc_52155_new_n9742_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__107_));
AND2X2 AND2X2_3869 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_108_), .Y(u2__abc_52155_new_n9744_));
AND2X2 AND2X2_387 ( .A(_abc_73687_new_n1682_), .B(\a[125] ), .Y(_abc_73687_new_n1683_));
AND2X2 AND2X2_3870 ( .A(u2__abc_52155_new_n9746_), .B(u2__abc_52155_new_n3784_), .Y(u2__abc_52155_new_n9747_));
AND2X2 AND2X2_3871 ( .A(u2__abc_52155_new_n3782_), .B(u2__abc_52155_new_n3771_), .Y(u2__abc_52155_new_n9748_));
AND2X2 AND2X2_3872 ( .A(u2__abc_52155_new_n9676_), .B(u2__abc_52155_new_n3800_), .Y(u2__abc_52155_new_n9751_));
AND2X2 AND2X2_3873 ( .A(u2__abc_52155_new_n9752_), .B(u2__abc_52155_new_n3829_), .Y(u2__abc_52155_new_n9753_));
AND2X2 AND2X2_3874 ( .A(u2__abc_52155_new_n9755_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9756_));
AND2X2 AND2X2_3875 ( .A(u2__abc_52155_new_n9756_), .B(u2__abc_52155_new_n9754_), .Y(u2__abc_52155_new_n9757_));
AND2X2 AND2X2_3876 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_106_), .Y(u2__abc_52155_new_n9758_));
AND2X2 AND2X2_3877 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3804_), .Y(u2__abc_52155_new_n9761_));
AND2X2 AND2X2_3878 ( .A(u2__abc_52155_new_n9762_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9763_));
AND2X2 AND2X2_3879 ( .A(u2__abc_52155_new_n9760_), .B(u2__abc_52155_new_n9763_), .Y(u2__abc_52155_new_n9764_));
AND2X2 AND2X2_388 ( .A(_abc_73687_new_n1684_), .B(\a[126] ), .Y(_abc_73687_new_n1685_));
AND2X2 AND2X2_3880 ( .A(u2__abc_52155_new_n9765_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__108_));
AND2X2 AND2X2_3881 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_109_), .Y(u2__abc_52155_new_n9767_));
AND2X2 AND2X2_3882 ( .A(u2__abc_52155_new_n9754_), .B(u2__abc_52155_new_n3825_), .Y(u2__abc_52155_new_n9768_));
AND2X2 AND2X2_3883 ( .A(u2__abc_52155_new_n9768_), .B(u2__abc_52155_new_n3822_), .Y(u2__abc_52155_new_n9769_));
AND2X2 AND2X2_3884 ( .A(u2__abc_52155_new_n9771_), .B(u2__abc_52155_new_n9770_), .Y(u2__abc_52155_new_n9772_));
AND2X2 AND2X2_3885 ( .A(u2__abc_52155_new_n9773_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9774_));
AND2X2 AND2X2_3886 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_107_), .Y(u2__abc_52155_new_n9775_));
AND2X2 AND2X2_3887 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3811_), .Y(u2__abc_52155_new_n9778_));
AND2X2 AND2X2_3888 ( .A(u2__abc_52155_new_n9779_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9780_));
AND2X2 AND2X2_3889 ( .A(u2__abc_52155_new_n9777_), .B(u2__abc_52155_new_n9780_), .Y(u2__abc_52155_new_n9781_));
AND2X2 AND2X2_389 ( .A(_abc_73687_new_n1686_), .B(_abc_73687_new_n753_), .Y(_abc_73687_new_n1687_));
AND2X2 AND2X2_3890 ( .A(u2__abc_52155_new_n9782_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__109_));
AND2X2 AND2X2_3891 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_110_), .Y(u2__abc_52155_new_n9784_));
AND2X2 AND2X2_3892 ( .A(u2__abc_52155_new_n3818_), .B(u2__abc_52155_new_n3825_), .Y(u2__abc_52155_new_n9785_));
AND2X2 AND2X2_3893 ( .A(u2__abc_52155_new_n9754_), .B(u2__abc_52155_new_n9785_), .Y(u2__abc_52155_new_n9786_));
AND2X2 AND2X2_3894 ( .A(u2__abc_52155_new_n9788_), .B(u2__abc_52155_new_n3807_), .Y(u2__abc_52155_new_n9789_));
AND2X2 AND2X2_3895 ( .A(u2__abc_52155_new_n9791_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9792_));
AND2X2 AND2X2_3896 ( .A(u2__abc_52155_new_n9792_), .B(u2__abc_52155_new_n9790_), .Y(u2__abc_52155_new_n9793_));
AND2X2 AND2X2_3897 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_108_), .Y(u2__abc_52155_new_n9794_));
AND2X2 AND2X2_3898 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3709_), .Y(u2__abc_52155_new_n9797_));
AND2X2 AND2X2_3899 ( .A(u2__abc_52155_new_n9798_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9799_));
AND2X2 AND2X2_39 ( .A(_abc_73687_new_n753_), .B(sqrto_38_), .Y(\o[74] ));
AND2X2 AND2X2_390 ( .A(aNan), .B(\a[127] ), .Y(\o[241] ));
AND2X2 AND2X2_3900 ( .A(u2__abc_52155_new_n9796_), .B(u2__abc_52155_new_n9799_), .Y(u2__abc_52155_new_n9800_));
AND2X2 AND2X2_3901 ( .A(u2__abc_52155_new_n9801_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__110_));
AND2X2 AND2X2_3902 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_111_), .Y(u2__abc_52155_new_n9803_));
AND2X2 AND2X2_3903 ( .A(u2__abc_52155_new_n9790_), .B(u2__abc_52155_new_n3803_), .Y(u2__abc_52155_new_n9804_));
AND2X2 AND2X2_3904 ( .A(u2__abc_52155_new_n9804_), .B(u2__abc_52155_new_n3814_), .Y(u2__abc_52155_new_n9805_));
AND2X2 AND2X2_3905 ( .A(u2__abc_52155_new_n9807_), .B(u2__abc_52155_new_n9806_), .Y(u2__abc_52155_new_n9808_));
AND2X2 AND2X2_3906 ( .A(u2__abc_52155_new_n9809_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9810_));
AND2X2 AND2X2_3907 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_109_), .Y(u2__abc_52155_new_n9811_));
AND2X2 AND2X2_3908 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3716_), .Y(u2__abc_52155_new_n9814_));
AND2X2 AND2X2_3909 ( .A(u2__abc_52155_new_n9815_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9816_));
AND2X2 AND2X2_391 ( .A(\a[121] ), .B(\a[122] ), .Y(u1__abc_51895_new_n152_));
AND2X2 AND2X2_3910 ( .A(u2__abc_52155_new_n9813_), .B(u2__abc_52155_new_n9816_), .Y(u2__abc_52155_new_n9817_));
AND2X2 AND2X2_3911 ( .A(u2__abc_52155_new_n9818_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__111_));
AND2X2 AND2X2_3912 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_112_), .Y(u2__abc_52155_new_n9820_));
AND2X2 AND2X2_3913 ( .A(u2__abc_52155_new_n9674_), .B(u2__abc_52155_new_n3832_), .Y(u2__abc_52155_new_n9821_));
AND2X2 AND2X2_3914 ( .A(u2__abc_52155_new_n9750_), .B(u2__abc_52155_new_n3831_), .Y(u2__abc_52155_new_n9822_));
AND2X2 AND2X2_3915 ( .A(u2__abc_52155_new_n9824_), .B(u2__abc_52155_new_n3815_), .Y(u2__abc_52155_new_n9825_));
AND2X2 AND2X2_3916 ( .A(u2__abc_52155_new_n3813_), .B(u2__abc_52155_new_n3802_), .Y(u2__abc_52155_new_n9826_));
AND2X2 AND2X2_3917 ( .A(u2__abc_52155_new_n9520_), .B(u2__abc_52155_new_n3893_), .Y(u2__abc_52155_new_n9831_));
AND2X2 AND2X2_3918 ( .A(u2__abc_52155_new_n9832_), .B(u2__abc_52155_new_n3712_), .Y(u2__abc_52155_new_n9833_));
AND2X2 AND2X2_3919 ( .A(u2__abc_52155_new_n9834_), .B(u2__abc_52155_new_n9835_), .Y(u2__abc_52155_new_n9836_));
AND2X2 AND2X2_392 ( .A(\a[119] ), .B(\a[120] ), .Y(u1__abc_51895_new_n153_));
AND2X2 AND2X2_3920 ( .A(u2__abc_52155_new_n9836_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9837_));
AND2X2 AND2X2_3921 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_110_), .Y(u2__abc_52155_new_n9838_));
AND2X2 AND2X2_3922 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3724_), .Y(u2__abc_52155_new_n9841_));
AND2X2 AND2X2_3923 ( .A(u2__abc_52155_new_n9842_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9843_));
AND2X2 AND2X2_3924 ( .A(u2__abc_52155_new_n9840_), .B(u2__abc_52155_new_n9843_), .Y(u2__abc_52155_new_n9844_));
AND2X2 AND2X2_3925 ( .A(u2__abc_52155_new_n9845_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__112_));
AND2X2 AND2X2_3926 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_113_), .Y(u2__abc_52155_new_n9847_));
AND2X2 AND2X2_3927 ( .A(u2__abc_52155_new_n9834_), .B(u2__abc_52155_new_n3708_), .Y(u2__abc_52155_new_n9849_));
AND2X2 AND2X2_3928 ( .A(u2__abc_52155_new_n9852_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9853_));
AND2X2 AND2X2_3929 ( .A(u2__abc_52155_new_n9853_), .B(u2__abc_52155_new_n9850_), .Y(u2__abc_52155_new_n9854_));
AND2X2 AND2X2_393 ( .A(u1__abc_51895_new_n152_), .B(u1__abc_51895_new_n153_), .Y(u1__abc_51895_new_n154_));
AND2X2 AND2X2_3930 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_111_), .Y(u2__abc_52155_new_n9855_));
AND2X2 AND2X2_3931 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3731_), .Y(u2__abc_52155_new_n9858_));
AND2X2 AND2X2_3932 ( .A(u2__abc_52155_new_n9859_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9860_));
AND2X2 AND2X2_3933 ( .A(u2__abc_52155_new_n9857_), .B(u2__abc_52155_new_n9860_), .Y(u2__abc_52155_new_n9861_));
AND2X2 AND2X2_3934 ( .A(u2__abc_52155_new_n9862_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__113_));
AND2X2 AND2X2_3935 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_114_), .Y(u2__abc_52155_new_n9864_));
AND2X2 AND2X2_3936 ( .A(u2__abc_52155_new_n9865_), .B(u2__abc_52155_new_n3715_), .Y(u2__abc_52155_new_n9866_));
AND2X2 AND2X2_3937 ( .A(u2__abc_52155_new_n9832_), .B(u2__abc_52155_new_n3720_), .Y(u2__abc_52155_new_n9868_));
AND2X2 AND2X2_3938 ( .A(u2__abc_52155_new_n9869_), .B(u2__abc_52155_new_n3727_), .Y(u2__abc_52155_new_n9870_));
AND2X2 AND2X2_3939 ( .A(u2__abc_52155_new_n9872_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9873_));
AND2X2 AND2X2_394 ( .A(\a[125] ), .B(\a[126] ), .Y(u1__abc_51895_new_n155_));
AND2X2 AND2X2_3940 ( .A(u2__abc_52155_new_n9873_), .B(u2__abc_52155_new_n9871_), .Y(u2__abc_52155_new_n9874_));
AND2X2 AND2X2_3941 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_112_), .Y(u2__abc_52155_new_n9875_));
AND2X2 AND2X2_3942 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3762_), .Y(u2__abc_52155_new_n9878_));
AND2X2 AND2X2_3943 ( .A(u2__abc_52155_new_n9879_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9880_));
AND2X2 AND2X2_3944 ( .A(u2__abc_52155_new_n9877_), .B(u2__abc_52155_new_n9880_), .Y(u2__abc_52155_new_n9881_));
AND2X2 AND2X2_3945 ( .A(u2__abc_52155_new_n9882_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__114_));
AND2X2 AND2X2_3946 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_115_), .Y(u2__abc_52155_new_n9884_));
AND2X2 AND2X2_3947 ( .A(u2__abc_52155_new_n9871_), .B(u2__abc_52155_new_n3723_), .Y(u2__abc_52155_new_n9886_));
AND2X2 AND2X2_3948 ( .A(u2__abc_52155_new_n9889_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9890_));
AND2X2 AND2X2_3949 ( .A(u2__abc_52155_new_n9890_), .B(u2__abc_52155_new_n9887_), .Y(u2__abc_52155_new_n9891_));
AND2X2 AND2X2_395 ( .A(\a[123] ), .B(\a[124] ), .Y(u1__abc_51895_new_n156_));
AND2X2 AND2X2_3950 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_113_), .Y(u2__abc_52155_new_n9892_));
AND2X2 AND2X2_3951 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3755_), .Y(u2__abc_52155_new_n9895_));
AND2X2 AND2X2_3952 ( .A(u2__abc_52155_new_n9896_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9897_));
AND2X2 AND2X2_3953 ( .A(u2__abc_52155_new_n9894_), .B(u2__abc_52155_new_n9897_), .Y(u2__abc_52155_new_n9898_));
AND2X2 AND2X2_3954 ( .A(u2__abc_52155_new_n9899_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__115_));
AND2X2 AND2X2_3955 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_116_), .Y(u2__abc_52155_new_n9901_));
AND2X2 AND2X2_3956 ( .A(u2__abc_52155_new_n9867_), .B(u2__abc_52155_new_n3735_), .Y(u2__abc_52155_new_n9902_));
AND2X2 AND2X2_3957 ( .A(u2__abc_52155_new_n3733_), .B(u2__abc_52155_new_n3722_), .Y(u2__abc_52155_new_n9903_));
AND2X2 AND2X2_3958 ( .A(u2__abc_52155_new_n9832_), .B(u2__abc_52155_new_n3736_), .Y(u2__abc_52155_new_n9906_));
AND2X2 AND2X2_3959 ( .A(u2__abc_52155_new_n9907_), .B(u2__abc_52155_new_n3765_), .Y(u2__abc_52155_new_n9908_));
AND2X2 AND2X2_396 ( .A(u1__abc_51895_new_n155_), .B(u1__abc_51895_new_n156_), .Y(u1__abc_51895_new_n157_));
AND2X2 AND2X2_3960 ( .A(u2__abc_52155_new_n9910_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9911_));
AND2X2 AND2X2_3961 ( .A(u2__abc_52155_new_n9911_), .B(u2__abc_52155_new_n9909_), .Y(u2__abc_52155_new_n9912_));
AND2X2 AND2X2_3962 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_114_), .Y(u2__abc_52155_new_n9913_));
AND2X2 AND2X2_3963 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3740_), .Y(u2__abc_52155_new_n9916_));
AND2X2 AND2X2_3964 ( .A(u2__abc_52155_new_n9917_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9918_));
AND2X2 AND2X2_3965 ( .A(u2__abc_52155_new_n9915_), .B(u2__abc_52155_new_n9918_), .Y(u2__abc_52155_new_n9919_));
AND2X2 AND2X2_3966 ( .A(u2__abc_52155_new_n9920_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__116_));
AND2X2 AND2X2_3967 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_117_), .Y(u2__abc_52155_new_n9922_));
AND2X2 AND2X2_3968 ( .A(u2__abc_52155_new_n9909_), .B(u2__abc_52155_new_n3761_), .Y(u2__abc_52155_new_n9923_));
AND2X2 AND2X2_3969 ( .A(u2__abc_52155_new_n9924_), .B(u2__abc_52155_new_n3758_), .Y(u2__abc_52155_new_n9925_));
AND2X2 AND2X2_397 ( .A(u1__abc_51895_new_n154_), .B(u1__abc_51895_new_n157_), .Y(u1__abc_51895_new_n158_));
AND2X2 AND2X2_3970 ( .A(u2__abc_52155_new_n9927_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9928_));
AND2X2 AND2X2_3971 ( .A(u2__abc_52155_new_n9928_), .B(u2__abc_52155_new_n9926_), .Y(u2__abc_52155_new_n9929_));
AND2X2 AND2X2_3972 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_115_), .Y(u2__abc_52155_new_n9930_));
AND2X2 AND2X2_3973 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3747_), .Y(u2__abc_52155_new_n9933_));
AND2X2 AND2X2_3974 ( .A(u2__abc_52155_new_n9934_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9935_));
AND2X2 AND2X2_3975 ( .A(u2__abc_52155_new_n9932_), .B(u2__abc_52155_new_n9935_), .Y(u2__abc_52155_new_n9936_));
AND2X2 AND2X2_3976 ( .A(u2__abc_52155_new_n9937_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__117_));
AND2X2 AND2X2_3977 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_118_), .Y(u2__abc_52155_new_n9939_));
AND2X2 AND2X2_3978 ( .A(u2__abc_52155_new_n9926_), .B(u2__abc_52155_new_n3754_), .Y(u2__abc_52155_new_n9940_));
AND2X2 AND2X2_3979 ( .A(u2__abc_52155_new_n9941_), .B(u2__abc_52155_new_n3743_), .Y(u2__abc_52155_new_n9942_));
AND2X2 AND2X2_398 ( .A(\a[113] ), .B(\a[114] ), .Y(u1__abc_51895_new_n159_));
AND2X2 AND2X2_3980 ( .A(u2__abc_52155_new_n9944_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9945_));
AND2X2 AND2X2_3981 ( .A(u2__abc_52155_new_n9945_), .B(u2__abc_52155_new_n9943_), .Y(u2__abc_52155_new_n9946_));
AND2X2 AND2X2_3982 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_116_), .Y(u2__abc_52155_new_n9947_));
AND2X2 AND2X2_3983 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3646_), .Y(u2__abc_52155_new_n9950_));
AND2X2 AND2X2_3984 ( .A(u2__abc_52155_new_n9951_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9952_));
AND2X2 AND2X2_3985 ( .A(u2__abc_52155_new_n9949_), .B(u2__abc_52155_new_n9952_), .Y(u2__abc_52155_new_n9953_));
AND2X2 AND2X2_3986 ( .A(u2__abc_52155_new_n9954_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__118_));
AND2X2 AND2X2_3987 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_119_), .Y(u2__abc_52155_new_n9956_));
AND2X2 AND2X2_3988 ( .A(u2__abc_52155_new_n9943_), .B(u2__abc_52155_new_n3739_), .Y(u2__abc_52155_new_n9957_));
AND2X2 AND2X2_3989 ( .A(u2__abc_52155_new_n9957_), .B(u2__abc_52155_new_n3750_), .Y(u2__abc_52155_new_n9958_));
AND2X2 AND2X2_399 ( .A(u1__abc_51895_new_n159_), .B(\a[112] ), .Y(u1__abc_51895_new_n160_));
AND2X2 AND2X2_3990 ( .A(u2__abc_52155_new_n9960_), .B(u2__abc_52155_new_n9959_), .Y(u2__abc_52155_new_n9961_));
AND2X2 AND2X2_3991 ( .A(u2__abc_52155_new_n9962_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9963_));
AND2X2 AND2X2_3992 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_117_), .Y(u2__abc_52155_new_n9964_));
AND2X2 AND2X2_3993 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3653_), .Y(u2__abc_52155_new_n9967_));
AND2X2 AND2X2_3994 ( .A(u2__abc_52155_new_n9968_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9969_));
AND2X2 AND2X2_3995 ( .A(u2__abc_52155_new_n9966_), .B(u2__abc_52155_new_n9969_), .Y(u2__abc_52155_new_n9970_));
AND2X2 AND2X2_3996 ( .A(u2__abc_52155_new_n9971_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__119_));
AND2X2 AND2X2_3997 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_120_), .Y(u2__abc_52155_new_n9973_));
AND2X2 AND2X2_3998 ( .A(u2__abc_52155_new_n9905_), .B(u2__abc_52155_new_n3767_), .Y(u2__abc_52155_new_n9974_));
AND2X2 AND2X2_3999 ( .A(u2__abc_52155_new_n9975_), .B(u2__abc_52155_new_n3757_), .Y(u2__abc_52155_new_n9976_));
AND2X2 AND2X2_4 ( .A(_abc_73687_new_n753_), .B(sqrto_3_), .Y(\o[39] ));
AND2X2 AND2X2_40 ( .A(_abc_73687_new_n753_), .B(sqrto_39_), .Y(\o[75] ));
AND2X2 AND2X2_400 ( .A(\a[117] ), .B(\a[118] ), .Y(u1__abc_51895_new_n161_));
AND2X2 AND2X2_4000 ( .A(u2__abc_52155_new_n3751_), .B(u2__abc_52155_new_n9976_), .Y(u2__abc_52155_new_n9977_));
AND2X2 AND2X2_4001 ( .A(u2__abc_52155_new_n3749_), .B(u2__abc_52155_new_n3738_), .Y(u2__abc_52155_new_n9978_));
AND2X2 AND2X2_4002 ( .A(u2__abc_52155_new_n9832_), .B(u2__abc_52155_new_n3768_), .Y(u2__abc_52155_new_n9982_));
AND2X2 AND2X2_4003 ( .A(u2__abc_52155_new_n9983_), .B(u2__abc_52155_new_n3649_), .Y(u2__abc_52155_new_n9984_));
AND2X2 AND2X2_4004 ( .A(u2__abc_52155_new_n9986_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n9987_));
AND2X2 AND2X2_4005 ( .A(u2__abc_52155_new_n9987_), .B(u2__abc_52155_new_n9985_), .Y(u2__abc_52155_new_n9988_));
AND2X2 AND2X2_4006 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_118_), .Y(u2__abc_52155_new_n9989_));
AND2X2 AND2X2_4007 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3661_), .Y(u2__abc_52155_new_n9992_));
AND2X2 AND2X2_4008 ( .A(u2__abc_52155_new_n9993_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n9994_));
AND2X2 AND2X2_4009 ( .A(u2__abc_52155_new_n9991_), .B(u2__abc_52155_new_n9994_), .Y(u2__abc_52155_new_n9995_));
AND2X2 AND2X2_401 ( .A(\a[115] ), .B(\a[116] ), .Y(u1__abc_51895_new_n162_));
AND2X2 AND2X2_4010 ( .A(u2__abc_52155_new_n9996_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__120_));
AND2X2 AND2X2_4011 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_121_), .Y(u2__abc_52155_new_n9998_));
AND2X2 AND2X2_4012 ( .A(u2__abc_52155_new_n9985_), .B(u2__abc_52155_new_n3645_), .Y(u2__abc_52155_new_n10000_));
AND2X2 AND2X2_4013 ( .A(u2__abc_52155_new_n10003_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10004_));
AND2X2 AND2X2_4014 ( .A(u2__abc_52155_new_n10004_), .B(u2__abc_52155_new_n10001_), .Y(u2__abc_52155_new_n10005_));
AND2X2 AND2X2_4015 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_119_), .Y(u2__abc_52155_new_n10006_));
AND2X2 AND2X2_4016 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3668_), .Y(u2__abc_52155_new_n10009_));
AND2X2 AND2X2_4017 ( .A(u2__abc_52155_new_n10010_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10011_));
AND2X2 AND2X2_4018 ( .A(u2__abc_52155_new_n10008_), .B(u2__abc_52155_new_n10011_), .Y(u2__abc_52155_new_n10012_));
AND2X2 AND2X2_4019 ( .A(u2__abc_52155_new_n10013_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__121_));
AND2X2 AND2X2_402 ( .A(u1__abc_51895_new_n161_), .B(u1__abc_51895_new_n162_), .Y(u1__abc_51895_new_n163_));
AND2X2 AND2X2_4020 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_122_), .Y(u2__abc_52155_new_n10015_));
AND2X2 AND2X2_4021 ( .A(u2__abc_52155_new_n10016_), .B(u2__abc_52155_new_n3652_), .Y(u2__abc_52155_new_n10017_));
AND2X2 AND2X2_4022 ( .A(u2__abc_52155_new_n9983_), .B(u2__abc_52155_new_n3657_), .Y(u2__abc_52155_new_n10019_));
AND2X2 AND2X2_4023 ( .A(u2__abc_52155_new_n10020_), .B(u2__abc_52155_new_n3664_), .Y(u2__abc_52155_new_n10021_));
AND2X2 AND2X2_4024 ( .A(u2__abc_52155_new_n10023_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10024_));
AND2X2 AND2X2_4025 ( .A(u2__abc_52155_new_n10024_), .B(u2__abc_52155_new_n10022_), .Y(u2__abc_52155_new_n10025_));
AND2X2 AND2X2_4026 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_120_), .Y(u2__abc_52155_new_n10026_));
AND2X2 AND2X2_4027 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3699_), .Y(u2__abc_52155_new_n10029_));
AND2X2 AND2X2_4028 ( .A(u2__abc_52155_new_n10030_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10031_));
AND2X2 AND2X2_4029 ( .A(u2__abc_52155_new_n10028_), .B(u2__abc_52155_new_n10031_), .Y(u2__abc_52155_new_n10032_));
AND2X2 AND2X2_403 ( .A(u1__abc_51895_new_n163_), .B(u1__abc_51895_new_n160_), .Y(u1__abc_51895_new_n164_));
AND2X2 AND2X2_4030 ( .A(u2__abc_52155_new_n10033_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__122_));
AND2X2 AND2X2_4031 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_123_), .Y(u2__abc_52155_new_n10035_));
AND2X2 AND2X2_4032 ( .A(u2__abc_52155_new_n10022_), .B(u2__abc_52155_new_n3660_), .Y(u2__abc_52155_new_n10036_));
AND2X2 AND2X2_4033 ( .A(u2__abc_52155_new_n10036_), .B(u2__abc_52155_new_n3671_), .Y(u2__abc_52155_new_n10037_));
AND2X2 AND2X2_4034 ( .A(u2__abc_52155_new_n10039_), .B(u2__abc_52155_new_n10038_), .Y(u2__abc_52155_new_n10040_));
AND2X2 AND2X2_4035 ( .A(u2__abc_52155_new_n10041_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10042_));
AND2X2 AND2X2_4036 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_121_), .Y(u2__abc_52155_new_n10043_));
AND2X2 AND2X2_4037 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3692_), .Y(u2__abc_52155_new_n10046_));
AND2X2 AND2X2_4038 ( .A(u2__abc_52155_new_n10047_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10048_));
AND2X2 AND2X2_4039 ( .A(u2__abc_52155_new_n10045_), .B(u2__abc_52155_new_n10048_), .Y(u2__abc_52155_new_n10049_));
AND2X2 AND2X2_404 ( .A(u1__abc_51895_new_n158_), .B(u1__abc_51895_new_n164_), .Y(u1_xinf));
AND2X2 AND2X2_4040 ( .A(u2__abc_52155_new_n10050_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__123_));
AND2X2 AND2X2_4041 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_124_), .Y(u2__abc_52155_new_n10052_));
AND2X2 AND2X2_4042 ( .A(u2__abc_52155_new_n10018_), .B(u2__abc_52155_new_n3672_), .Y(u2__abc_52155_new_n10053_));
AND2X2 AND2X2_4043 ( .A(u2__abc_52155_new_n3670_), .B(u2__abc_52155_new_n3659_), .Y(u2__abc_52155_new_n10054_));
AND2X2 AND2X2_4044 ( .A(u2__abc_52155_new_n9983_), .B(u2__abc_52155_new_n3673_), .Y(u2__abc_52155_new_n10057_));
AND2X2 AND2X2_4045 ( .A(u2__abc_52155_new_n10058_), .B(u2__abc_52155_new_n3702_), .Y(u2__abc_52155_new_n10059_));
AND2X2 AND2X2_4046 ( .A(u2__abc_52155_new_n10061_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10062_));
AND2X2 AND2X2_4047 ( .A(u2__abc_52155_new_n10062_), .B(u2__abc_52155_new_n10060_), .Y(u2__abc_52155_new_n10063_));
AND2X2 AND2X2_4048 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_122_), .Y(u2__abc_52155_new_n10064_));
AND2X2 AND2X2_4049 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3677_), .Y(u2__abc_52155_new_n10067_));
AND2X2 AND2X2_405 ( .A(u1__abc_51895_new_n166_), .B(u1__abc_51895_new_n167_), .Y(u1__abc_51895_new_n168_));
AND2X2 AND2X2_4050 ( .A(u2__abc_52155_new_n10068_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10069_));
AND2X2 AND2X2_4051 ( .A(u2__abc_52155_new_n10066_), .B(u2__abc_52155_new_n10069_), .Y(u2__abc_52155_new_n10070_));
AND2X2 AND2X2_4052 ( .A(u2__abc_52155_new_n10071_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__124_));
AND2X2 AND2X2_4053 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_125_), .Y(u2__abc_52155_new_n10073_));
AND2X2 AND2X2_4054 ( .A(u2__abc_52155_new_n10060_), .B(u2__abc_52155_new_n3698_), .Y(u2__abc_52155_new_n10074_));
AND2X2 AND2X2_4055 ( .A(u2__abc_52155_new_n10074_), .B(u2__abc_52155_new_n3695_), .Y(u2__abc_52155_new_n10075_));
AND2X2 AND2X2_4056 ( .A(u2__abc_52155_new_n10077_), .B(u2__abc_52155_new_n10076_), .Y(u2__abc_52155_new_n10078_));
AND2X2 AND2X2_4057 ( .A(u2__abc_52155_new_n10079_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10080_));
AND2X2 AND2X2_4058 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_123_), .Y(u2__abc_52155_new_n10081_));
AND2X2 AND2X2_4059 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3681_), .Y(u2__abc_52155_new_n10084_));
AND2X2 AND2X2_406 ( .A(u1__abc_51895_new_n169_), .B(u1__abc_51895_new_n170_), .Y(u1__abc_51895_new_n171_));
AND2X2 AND2X2_4060 ( .A(u2__abc_52155_new_n10085_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10086_));
AND2X2 AND2X2_4061 ( .A(u2__abc_52155_new_n10083_), .B(u2__abc_52155_new_n10086_), .Y(u2__abc_52155_new_n10087_));
AND2X2 AND2X2_4062 ( .A(u2__abc_52155_new_n10088_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__125_));
AND2X2 AND2X2_4063 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_126_), .Y(u2__abc_52155_new_n10090_));
AND2X2 AND2X2_4064 ( .A(u2__abc_52155_new_n3691_), .B(u2__abc_52155_new_n3698_), .Y(u2__abc_52155_new_n10091_));
AND2X2 AND2X2_4065 ( .A(u2__abc_52155_new_n10060_), .B(u2__abc_52155_new_n10091_), .Y(u2__abc_52155_new_n10092_));
AND2X2 AND2X2_4066 ( .A(u2__abc_52155_new_n10094_), .B(u2__abc_52155_new_n3680_), .Y(u2__abc_52155_new_n10095_));
AND2X2 AND2X2_4067 ( .A(u2__abc_52155_new_n10097_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10098_));
AND2X2 AND2X2_4068 ( .A(u2__abc_52155_new_n10098_), .B(u2__abc_52155_new_n10096_), .Y(u2__abc_52155_new_n10099_));
AND2X2 AND2X2_4069 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_124_), .Y(u2__abc_52155_new_n10100_));
AND2X2 AND2X2_407 ( .A(u1__abc_51895_new_n168_), .B(u1__abc_51895_new_n171_), .Y(u1__abc_51895_new_n172_));
AND2X2 AND2X2_4070 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n10103_), .Y(u2__abc_52155_new_n10104_));
AND2X2 AND2X2_4071 ( .A(u2__abc_52155_new_n10105_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10106_));
AND2X2 AND2X2_4072 ( .A(u2__abc_52155_new_n10102_), .B(u2__abc_52155_new_n10106_), .Y(u2__abc_52155_new_n10107_));
AND2X2 AND2X2_4073 ( .A(u2__abc_52155_new_n10108_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__126_));
AND2X2 AND2X2_4074 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_127_), .Y(u2__abc_52155_new_n10110_));
AND2X2 AND2X2_4075 ( .A(u2__abc_52155_new_n10096_), .B(u2__abc_52155_new_n3676_), .Y(u2__abc_52155_new_n10111_));
AND2X2 AND2X2_4076 ( .A(u2__abc_52155_new_n10111_), .B(u2__abc_52155_new_n3687_), .Y(u2__abc_52155_new_n10112_));
AND2X2 AND2X2_4077 ( .A(u2__abc_52155_new_n10114_), .B(u2__abc_52155_new_n10113_), .Y(u2__abc_52155_new_n10115_));
AND2X2 AND2X2_4078 ( .A(u2__abc_52155_new_n10116_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10117_));
AND2X2 AND2X2_4079 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_125_), .Y(u2__abc_52155_new_n10118_));
AND2X2 AND2X2_408 ( .A(u1__abc_51895_new_n173_), .B(u1__abc_51895_new_n174_), .Y(u1__abc_51895_new_n175_));
AND2X2 AND2X2_4080 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5241_), .Y(u2__abc_52155_new_n10121_));
AND2X2 AND2X2_4081 ( .A(u2__abc_52155_new_n10122_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10123_));
AND2X2 AND2X2_4082 ( .A(u2__abc_52155_new_n10120_), .B(u2__abc_52155_new_n10123_), .Y(u2__abc_52155_new_n10124_));
AND2X2 AND2X2_4083 ( .A(u2__abc_52155_new_n10125_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__127_));
AND2X2 AND2X2_4084 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_128_), .Y(u2__abc_52155_new_n10127_));
AND2X2 AND2X2_4085 ( .A(u2__abc_52155_new_n8878_), .B(u2__abc_52155_new_n4132_), .Y(u2__abc_52155_new_n10128_));
AND2X2 AND2X2_4086 ( .A(u2__abc_52155_new_n9518_), .B(u2__abc_52155_new_n3894_), .Y(u2__abc_52155_new_n10130_));
AND2X2 AND2X2_4087 ( .A(u2__abc_52155_new_n9830_), .B(u2__abc_52155_new_n3769_), .Y(u2__abc_52155_new_n10132_));
AND2X2 AND2X2_4088 ( .A(u2__abc_52155_new_n9981_), .B(u2__abc_52155_new_n3705_), .Y(u2__abc_52155_new_n10134_));
AND2X2 AND2X2_4089 ( .A(u2__abc_52155_new_n10056_), .B(u2__abc_52155_new_n3704_), .Y(u2__abc_52155_new_n10136_));
AND2X2 AND2X2_409 ( .A(u1__abc_51895_new_n176_), .B(u1__abc_51895_new_n177_), .Y(u1__abc_51895_new_n178_));
AND2X2 AND2X2_4090 ( .A(u2__abc_52155_new_n3676_), .B(u2__abc_52155_new_n3686_), .Y(u2__abc_52155_new_n10138_));
AND2X2 AND2X2_4091 ( .A(u2__abc_52155_new_n10141_), .B(u2__abc_52155_new_n3688_), .Y(u2__abc_52155_new_n10142_));
AND2X2 AND2X2_4092 ( .A(u2__abc_52155_new_n10143_), .B(u2__abc_52155_new_n10139_), .Y(u2__abc_52155_new_n10144_));
AND2X2 AND2X2_4093 ( .A(u2__abc_52155_new_n10137_), .B(u2__abc_52155_new_n10144_), .Y(u2__abc_52155_new_n10145_));
AND2X2 AND2X2_4094 ( .A(u2__abc_52155_new_n10135_), .B(u2__abc_52155_new_n10145_), .Y(u2__abc_52155_new_n10146_));
AND2X2 AND2X2_4095 ( .A(u2__abc_52155_new_n10133_), .B(u2__abc_52155_new_n10146_), .Y(u2__abc_52155_new_n10147_));
AND2X2 AND2X2_4096 ( .A(u2__abc_52155_new_n10131_), .B(u2__abc_52155_new_n10147_), .Y(u2__abc_52155_new_n10148_));
AND2X2 AND2X2_4097 ( .A(u2__abc_52155_new_n10129_), .B(u2__abc_52155_new_n10148_), .Y(u2__abc_52155_new_n10149_));
AND2X2 AND2X2_4098 ( .A(u2__abc_52155_new_n10150_), .B(u2__abc_52155_new_n5237_), .Y(u2__abc_52155_new_n10151_));
AND2X2 AND2X2_4099 ( .A(u2__abc_52155_new_n10152_), .B(u2__abc_52155_new_n10153_), .Y(u2__abc_52155_new_n10154_));
AND2X2 AND2X2_41 ( .A(_abc_73687_new_n753_), .B(sqrto_40_), .Y(\o[76] ));
AND2X2 AND2X2_410 ( .A(u1__abc_51895_new_n175_), .B(u1__abc_51895_new_n178_), .Y(u1__abc_51895_new_n179_));
AND2X2 AND2X2_4100 ( .A(u2__abc_52155_new_n10155_), .B(u2__abc_52155_new_n10156_), .Y(u2__abc_52155_new_n10157_));
AND2X2 AND2X2_4101 ( .A(u2__abc_52155_new_n2993_), .B(u2__abc_52155_new_n5248_), .Y(u2__abc_52155_new_n10159_));
AND2X2 AND2X2_4102 ( .A(u2__abc_52155_new_n10160_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10161_));
AND2X2 AND2X2_4103 ( .A(u2__abc_52155_new_n10158_), .B(u2__abc_52155_new_n10161_), .Y(u2__abc_52155_new_n10162_));
AND2X2 AND2X2_4104 ( .A(u2__abc_52155_new_n10163_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__128_));
AND2X2 AND2X2_4105 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_129_), .Y(u2__abc_52155_new_n10165_));
AND2X2 AND2X2_4106 ( .A(u2__abc_52155_new_n10152_), .B(u2__abc_52155_new_n5235_), .Y(u2__abc_52155_new_n10167_));
AND2X2 AND2X2_4107 ( .A(u2__abc_52155_new_n10170_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10171_));
AND2X2 AND2X2_4108 ( .A(u2__abc_52155_new_n10171_), .B(u2__abc_52155_new_n10168_), .Y(u2__abc_52155_new_n10172_));
AND2X2 AND2X2_4109 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_127_), .Y(u2__abc_52155_new_n10173_));
AND2X2 AND2X2_411 ( .A(u1__abc_51895_new_n172_), .B(u1__abc_51895_new_n179_), .Y(u1__abc_51895_new_n180_));
AND2X2 AND2X2_4110 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5253_), .Y(u2__abc_52155_new_n10176_));
AND2X2 AND2X2_4111 ( .A(u2__abc_52155_new_n10177_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10178_));
AND2X2 AND2X2_4112 ( .A(u2__abc_52155_new_n10175_), .B(u2__abc_52155_new_n10178_), .Y(u2__abc_52155_new_n10179_));
AND2X2 AND2X2_4113 ( .A(u2__abc_52155_new_n10180_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__129_));
AND2X2 AND2X2_4114 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_130_), .Y(u2__abc_52155_new_n10182_));
AND2X2 AND2X2_4115 ( .A(u2__abc_52155_new_n10184_), .B(u2__abc_52155_new_n5240_), .Y(u2__abc_52155_new_n10185_));
AND2X2 AND2X2_4116 ( .A(u2__abc_52155_new_n10150_), .B(u2__abc_52155_new_n5245_), .Y(u2__abc_52155_new_n10187_));
AND2X2 AND2X2_4117 ( .A(u2__abc_52155_new_n10188_), .B(u2__abc_52155_new_n10183_), .Y(u2__abc_52155_new_n10189_));
AND2X2 AND2X2_4118 ( .A(u2__abc_52155_new_n10190_), .B(u2__abc_52155_new_n10191_), .Y(u2__abc_52155_new_n10192_));
AND2X2 AND2X2_4119 ( .A(u2__abc_52155_new_n10192_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10193_));
AND2X2 AND2X2_412 ( .A(u1__abc_51895_new_n181_), .B(u1__abc_51895_new_n182_), .Y(u1__abc_51895_new_n183_));
AND2X2 AND2X2_4120 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_128_), .Y(u2__abc_52155_new_n10194_));
AND2X2 AND2X2_4121 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5277_), .Y(u2__abc_52155_new_n10197_));
AND2X2 AND2X2_4122 ( .A(u2__abc_52155_new_n10198_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10199_));
AND2X2 AND2X2_4123 ( .A(u2__abc_52155_new_n10196_), .B(u2__abc_52155_new_n10199_), .Y(u2__abc_52155_new_n10200_));
AND2X2 AND2X2_4124 ( .A(u2__abc_52155_new_n10201_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__130_));
AND2X2 AND2X2_4125 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_131_), .Y(u2__abc_52155_new_n10203_));
AND2X2 AND2X2_4126 ( .A(u2__abc_52155_new_n10190_), .B(u2__abc_52155_new_n10204_), .Y(u2__abc_52155_new_n10205_));
AND2X2 AND2X2_4127 ( .A(u2__abc_52155_new_n10209_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10210_));
AND2X2 AND2X2_4128 ( .A(u2__abc_52155_new_n10210_), .B(u2__abc_52155_new_n10206_), .Y(u2__abc_52155_new_n10211_));
AND2X2 AND2X2_4129 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_129_), .Y(u2__abc_52155_new_n10212_));
AND2X2 AND2X2_413 ( .A(u1__abc_51895_new_n184_), .B(u1__abc_51895_new_n185_), .Y(u1__abc_51895_new_n186_));
AND2X2 AND2X2_4130 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5272_), .Y(u2__abc_52155_new_n10215_));
AND2X2 AND2X2_4131 ( .A(u2__abc_52155_new_n10216_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10217_));
AND2X2 AND2X2_4132 ( .A(u2__abc_52155_new_n10214_), .B(u2__abc_52155_new_n10217_), .Y(u2__abc_52155_new_n10218_));
AND2X2 AND2X2_4133 ( .A(u2__abc_52155_new_n10219_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__131_));
AND2X2 AND2X2_4134 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_132_), .Y(u2__abc_52155_new_n10221_));
AND2X2 AND2X2_4135 ( .A(u2__abc_52155_new_n10186_), .B(u2__abc_52155_new_n5257_), .Y(u2__abc_52155_new_n10223_));
AND2X2 AND2X2_4136 ( .A(u2__abc_52155_new_n5297_), .B(u2__abc_52155_new_n5247_), .Y(u2__abc_52155_new_n10224_));
AND2X2 AND2X2_4137 ( .A(u2__abc_52155_new_n10150_), .B(u2__abc_52155_new_n5258_), .Y(u2__abc_52155_new_n10227_));
AND2X2 AND2X2_4138 ( .A(u2__abc_52155_new_n10228_), .B(u2__abc_52155_new_n10222_), .Y(u2__abc_52155_new_n10229_));
AND2X2 AND2X2_4139 ( .A(u2__abc_52155_new_n10230_), .B(u2__abc_52155_new_n10231_), .Y(u2__abc_52155_new_n10232_));
AND2X2 AND2X2_414 ( .A(u1__abc_51895_new_n183_), .B(u1__abc_51895_new_n186_), .Y(u1__abc_51895_new_n187_));
AND2X2 AND2X2_4140 ( .A(u2__abc_52155_new_n10232_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10233_));
AND2X2 AND2X2_4141 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_130_), .Y(u2__abc_52155_new_n10234_));
AND2X2 AND2X2_4142 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5261_), .Y(u2__abc_52155_new_n10237_));
AND2X2 AND2X2_4143 ( .A(u2__abc_52155_new_n10238_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10239_));
AND2X2 AND2X2_4144 ( .A(u2__abc_52155_new_n10236_), .B(u2__abc_52155_new_n10239_), .Y(u2__abc_52155_new_n10240_));
AND2X2 AND2X2_4145 ( .A(u2__abc_52155_new_n10241_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__132_));
AND2X2 AND2X2_4146 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_133_), .Y(u2__abc_52155_new_n10243_));
AND2X2 AND2X2_4147 ( .A(u2__abc_52155_new_n10230_), .B(u2__abc_52155_new_n10245_), .Y(u2__abc_52155_new_n10246_));
AND2X2 AND2X2_4148 ( .A(u2__abc_52155_new_n10246_), .B(u2__abc_52155_new_n10244_), .Y(u2__abc_52155_new_n10247_));
AND2X2 AND2X2_4149 ( .A(u2__abc_52155_new_n10248_), .B(u2__abc_52155_new_n5274_), .Y(u2__abc_52155_new_n10249_));
AND2X2 AND2X2_415 ( .A(u1__abc_51895_new_n188_), .B(u1__abc_51895_new_n189_), .Y(u1__abc_51895_new_n190_));
AND2X2 AND2X2_4150 ( .A(u2__abc_52155_new_n10250_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10251_));
AND2X2 AND2X2_4151 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_131_), .Y(u2__abc_52155_new_n10252_));
AND2X2 AND2X2_4152 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5266_), .Y(u2__abc_52155_new_n10255_));
AND2X2 AND2X2_4153 ( .A(u2__abc_52155_new_n10256_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10257_));
AND2X2 AND2X2_4154 ( .A(u2__abc_52155_new_n10254_), .B(u2__abc_52155_new_n10257_), .Y(u2__abc_52155_new_n10258_));
AND2X2 AND2X2_4155 ( .A(u2__abc_52155_new_n10259_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__133_));
AND2X2 AND2X2_4156 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_134_), .Y(u2__abc_52155_new_n10261_));
AND2X2 AND2X2_4157 ( .A(u2__abc_52155_new_n10230_), .B(u2__abc_52155_new_n10264_), .Y(u2__abc_52155_new_n10265_));
AND2X2 AND2X2_4158 ( .A(u2__abc_52155_new_n10267_), .B(u2__abc_52155_new_n10262_), .Y(u2__abc_52155_new_n10268_));
AND2X2 AND2X2_4159 ( .A(u2__abc_52155_new_n10270_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10271_));
AND2X2 AND2X2_416 ( .A(u1__abc_51895_new_n191_), .B(u1__abc_51895_new_n192_), .Y(u1__abc_51895_new_n193_));
AND2X2 AND2X2_4160 ( .A(u2__abc_52155_new_n10271_), .B(u2__abc_52155_new_n10269_), .Y(u2__abc_52155_new_n10272_));
AND2X2 AND2X2_4161 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_132_), .Y(u2__abc_52155_new_n10273_));
AND2X2 AND2X2_4162 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5188_), .Y(u2__abc_52155_new_n10276_));
AND2X2 AND2X2_4163 ( .A(u2__abc_52155_new_n10277_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10278_));
AND2X2 AND2X2_4164 ( .A(u2__abc_52155_new_n10275_), .B(u2__abc_52155_new_n10278_), .Y(u2__abc_52155_new_n10279_));
AND2X2 AND2X2_4165 ( .A(u2__abc_52155_new_n10280_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__134_));
AND2X2 AND2X2_4166 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_135_), .Y(u2__abc_52155_new_n10282_));
AND2X2 AND2X2_4167 ( .A(u2__abc_52155_new_n10269_), .B(u2__abc_52155_new_n10283_), .Y(u2__abc_52155_new_n10284_));
AND2X2 AND2X2_4168 ( .A(u2__abc_52155_new_n10288_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10289_));
AND2X2 AND2X2_4169 ( .A(u2__abc_52155_new_n10289_), .B(u2__abc_52155_new_n10285_), .Y(u2__abc_52155_new_n10290_));
AND2X2 AND2X2_417 ( .A(u1__abc_51895_new_n190_), .B(u1__abc_51895_new_n193_), .Y(u1__abc_51895_new_n194_));
AND2X2 AND2X2_4170 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_133_), .Y(u2__abc_52155_new_n10291_));
AND2X2 AND2X2_4171 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5195_), .Y(u2__abc_52155_new_n10294_));
AND2X2 AND2X2_4172 ( .A(u2__abc_52155_new_n10295_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10296_));
AND2X2 AND2X2_4173 ( .A(u2__abc_52155_new_n10293_), .B(u2__abc_52155_new_n10296_), .Y(u2__abc_52155_new_n10297_));
AND2X2 AND2X2_4174 ( .A(u2__abc_52155_new_n10298_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__135_));
AND2X2 AND2X2_4175 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_136_), .Y(u2__abc_52155_new_n10300_));
AND2X2 AND2X2_4176 ( .A(u2__abc_52155_new_n10226_), .B(u2__abc_52155_new_n5282_), .Y(u2__abc_52155_new_n10301_));
AND2X2 AND2X2_4177 ( .A(u2__abc_52155_new_n10305_), .B(u2__abc_52155_new_n5308_), .Y(u2__abc_52155_new_n10306_));
AND2X2 AND2X2_4178 ( .A(u2__abc_52155_new_n10304_), .B(u2__abc_52155_new_n10306_), .Y(u2__abc_52155_new_n10307_));
AND2X2 AND2X2_4179 ( .A(u2__abc_52155_new_n10302_), .B(u2__abc_52155_new_n10307_), .Y(u2__abc_52155_new_n10308_));
AND2X2 AND2X2_418 ( .A(u1__abc_51895_new_n187_), .B(u1__abc_51895_new_n194_), .Y(u1__abc_51895_new_n195_));
AND2X2 AND2X2_4180 ( .A(u2__abc_52155_new_n10150_), .B(u2__abc_52155_new_n5283_), .Y(u2__abc_52155_new_n10310_));
AND2X2 AND2X2_4181 ( .A(u2__abc_52155_new_n10311_), .B(u2__abc_52155_new_n5191_), .Y(u2__abc_52155_new_n10312_));
AND2X2 AND2X2_4182 ( .A(u2__abc_52155_new_n10313_), .B(u2__abc_52155_new_n10314_), .Y(u2__abc_52155_new_n10315_));
AND2X2 AND2X2_4183 ( .A(u2__abc_52155_new_n10315_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10316_));
AND2X2 AND2X2_4184 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_134_), .Y(u2__abc_52155_new_n10317_));
AND2X2 AND2X2_4185 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5175_), .Y(u2__abc_52155_new_n10320_));
AND2X2 AND2X2_4186 ( .A(u2__abc_52155_new_n10321_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10322_));
AND2X2 AND2X2_4187 ( .A(u2__abc_52155_new_n10319_), .B(u2__abc_52155_new_n10322_), .Y(u2__abc_52155_new_n10323_));
AND2X2 AND2X2_4188 ( .A(u2__abc_52155_new_n10324_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__136_));
AND2X2 AND2X2_4189 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_137_), .Y(u2__abc_52155_new_n10326_));
AND2X2 AND2X2_419 ( .A(u1__abc_51895_new_n180_), .B(u1__abc_51895_new_n195_), .Y(u1__abc_51895_new_n196_));
AND2X2 AND2X2_4190 ( .A(u2__abc_52155_new_n10313_), .B(u2__abc_52155_new_n5187_), .Y(u2__abc_52155_new_n10328_));
AND2X2 AND2X2_4191 ( .A(u2__abc_52155_new_n10329_), .B(u2__abc_52155_new_n10327_), .Y(u2__abc_52155_new_n10330_));
AND2X2 AND2X2_4192 ( .A(u2__abc_52155_new_n10328_), .B(u2__abc_52155_new_n5198_), .Y(u2__abc_52155_new_n10331_));
AND2X2 AND2X2_4193 ( .A(u2__abc_52155_new_n10332_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10333_));
AND2X2 AND2X2_4194 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_135_), .Y(u2__abc_52155_new_n10334_));
AND2X2 AND2X2_4195 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5180_), .Y(u2__abc_52155_new_n10337_));
AND2X2 AND2X2_4196 ( .A(u2__abc_52155_new_n10338_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10339_));
AND2X2 AND2X2_4197 ( .A(u2__abc_52155_new_n10336_), .B(u2__abc_52155_new_n10339_), .Y(u2__abc_52155_new_n10340_));
AND2X2 AND2X2_4198 ( .A(u2__abc_52155_new_n10341_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__137_));
AND2X2 AND2X2_4199 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_138_), .Y(u2__abc_52155_new_n10343_));
AND2X2 AND2X2_42 ( .A(_abc_73687_new_n753_), .B(sqrto_41_), .Y(\o[77] ));
AND2X2 AND2X2_420 ( .A(u1__abc_51895_new_n197_), .B(u1__abc_51895_new_n198_), .Y(u1__abc_51895_new_n199_));
AND2X2 AND2X2_4200 ( .A(u2__abc_52155_new_n10329_), .B(u2__abc_52155_new_n5197_), .Y(u2__abc_52155_new_n10345_));
AND2X2 AND2X2_4201 ( .A(u2__abc_52155_new_n10346_), .B(u2__abc_52155_new_n10344_), .Y(u2__abc_52155_new_n10347_));
AND2X2 AND2X2_4202 ( .A(u2__abc_52155_new_n10349_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10350_));
AND2X2 AND2X2_4203 ( .A(u2__abc_52155_new_n10350_), .B(u2__abc_52155_new_n10348_), .Y(u2__abc_52155_new_n10351_));
AND2X2 AND2X2_4204 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_136_), .Y(u2__abc_52155_new_n10352_));
AND2X2 AND2X2_4205 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5226_), .Y(u2__abc_52155_new_n10355_));
AND2X2 AND2X2_4206 ( .A(u2__abc_52155_new_n10356_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10357_));
AND2X2 AND2X2_4207 ( .A(u2__abc_52155_new_n10354_), .B(u2__abc_52155_new_n10357_), .Y(u2__abc_52155_new_n10358_));
AND2X2 AND2X2_4208 ( .A(u2__abc_52155_new_n10359_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__138_));
AND2X2 AND2X2_4209 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_139_), .Y(u2__abc_52155_new_n10361_));
AND2X2 AND2X2_421 ( .A(u1__abc_51895_new_n200_), .B(u1__abc_51895_new_n201_), .Y(u1__abc_51895_new_n202_));
AND2X2 AND2X2_4210 ( .A(u2__abc_52155_new_n10348_), .B(u2__abc_52155_new_n10362_), .Y(u2__abc_52155_new_n10363_));
AND2X2 AND2X2_4211 ( .A(u2__abc_52155_new_n10367_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10368_));
AND2X2 AND2X2_4212 ( .A(u2__abc_52155_new_n10368_), .B(u2__abc_52155_new_n10364_), .Y(u2__abc_52155_new_n10369_));
AND2X2 AND2X2_4213 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_137_), .Y(u2__abc_52155_new_n10370_));
AND2X2 AND2X2_4214 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5219_), .Y(u2__abc_52155_new_n10373_));
AND2X2 AND2X2_4215 ( .A(u2__abc_52155_new_n10374_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10375_));
AND2X2 AND2X2_4216 ( .A(u2__abc_52155_new_n10372_), .B(u2__abc_52155_new_n10375_), .Y(u2__abc_52155_new_n10376_));
AND2X2 AND2X2_4217 ( .A(u2__abc_52155_new_n10377_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__139_));
AND2X2 AND2X2_4218 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_140_), .Y(u2__abc_52155_new_n10379_));
AND2X2 AND2X2_4219 ( .A(u2__abc_52155_new_n5187_), .B(u2__abc_52155_new_n5194_), .Y(u2__abc_52155_new_n10380_));
AND2X2 AND2X2_422 ( .A(u1__abc_51895_new_n199_), .B(u1__abc_51895_new_n202_), .Y(u1__abc_51895_new_n203_));
AND2X2 AND2X2_4220 ( .A(u2__abc_52155_new_n10383_), .B(u2__abc_52155_new_n5319_), .Y(u2__abc_52155_new_n10384_));
AND2X2 AND2X2_4221 ( .A(u2__abc_52155_new_n10382_), .B(u2__abc_52155_new_n10384_), .Y(u2__abc_52155_new_n10385_));
AND2X2 AND2X2_4222 ( .A(u2__abc_52155_new_n10311_), .B(u2__abc_52155_new_n5200_), .Y(u2__abc_52155_new_n10387_));
AND2X2 AND2X2_4223 ( .A(u2__abc_52155_new_n10388_), .B(u2__abc_52155_new_n5229_), .Y(u2__abc_52155_new_n10389_));
AND2X2 AND2X2_4224 ( .A(u2__abc_52155_new_n10391_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10392_));
AND2X2 AND2X2_4225 ( .A(u2__abc_52155_new_n10392_), .B(u2__abc_52155_new_n10390_), .Y(u2__abc_52155_new_n10393_));
AND2X2 AND2X2_4226 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_138_), .Y(u2__abc_52155_new_n10394_));
AND2X2 AND2X2_4227 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5204_), .Y(u2__abc_52155_new_n10397_));
AND2X2 AND2X2_4228 ( .A(u2__abc_52155_new_n10398_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10399_));
AND2X2 AND2X2_4229 ( .A(u2__abc_52155_new_n10396_), .B(u2__abc_52155_new_n10399_), .Y(u2__abc_52155_new_n10400_));
AND2X2 AND2X2_423 ( .A(u1__abc_51895_new_n204_), .B(u1__abc_51895_new_n205_), .Y(u1__abc_51895_new_n206_));
AND2X2 AND2X2_4230 ( .A(u2__abc_52155_new_n10401_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__140_));
AND2X2 AND2X2_4231 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_141_), .Y(u2__abc_52155_new_n10403_));
AND2X2 AND2X2_4232 ( .A(u2__abc_52155_new_n10390_), .B(u2__abc_52155_new_n5225_), .Y(u2__abc_52155_new_n10404_));
AND2X2 AND2X2_4233 ( .A(u2__abc_52155_new_n10404_), .B(u2__abc_52155_new_n5222_), .Y(u2__abc_52155_new_n10405_));
AND2X2 AND2X2_4234 ( .A(u2__abc_52155_new_n10407_), .B(u2__abc_52155_new_n10406_), .Y(u2__abc_52155_new_n10408_));
AND2X2 AND2X2_4235 ( .A(u2__abc_52155_new_n10409_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10410_));
AND2X2 AND2X2_4236 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_139_), .Y(u2__abc_52155_new_n10411_));
AND2X2 AND2X2_4237 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5211_), .Y(u2__abc_52155_new_n10414_));
AND2X2 AND2X2_4238 ( .A(u2__abc_52155_new_n10415_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10416_));
AND2X2 AND2X2_4239 ( .A(u2__abc_52155_new_n10413_), .B(u2__abc_52155_new_n10416_), .Y(u2__abc_52155_new_n10417_));
AND2X2 AND2X2_424 ( .A(u1__abc_51895_new_n207_), .B(u1__abc_51895_new_n208_), .Y(u1__abc_51895_new_n209_));
AND2X2 AND2X2_4240 ( .A(u2__abc_52155_new_n10418_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__141_));
AND2X2 AND2X2_4241 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_142_), .Y(u2__abc_52155_new_n10420_));
AND2X2 AND2X2_4242 ( .A(u2__abc_52155_new_n5218_), .B(u2__abc_52155_new_n5225_), .Y(u2__abc_52155_new_n10421_));
AND2X2 AND2X2_4243 ( .A(u2__abc_52155_new_n10390_), .B(u2__abc_52155_new_n10421_), .Y(u2__abc_52155_new_n10422_));
AND2X2 AND2X2_4244 ( .A(u2__abc_52155_new_n10424_), .B(u2__abc_52155_new_n5207_), .Y(u2__abc_52155_new_n10425_));
AND2X2 AND2X2_4245 ( .A(u2__abc_52155_new_n10427_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10428_));
AND2X2 AND2X2_4246 ( .A(u2__abc_52155_new_n10428_), .B(u2__abc_52155_new_n10426_), .Y(u2__abc_52155_new_n10429_));
AND2X2 AND2X2_4247 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_140_), .Y(u2__abc_52155_new_n10430_));
AND2X2 AND2X2_4248 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5165_), .Y(u2__abc_52155_new_n10433_));
AND2X2 AND2X2_4249 ( .A(u2__abc_52155_new_n10434_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10435_));
AND2X2 AND2X2_425 ( .A(u1__abc_51895_new_n206_), .B(u1__abc_51895_new_n209_), .Y(u1__abc_51895_new_n210_));
AND2X2 AND2X2_4250 ( .A(u2__abc_52155_new_n10432_), .B(u2__abc_52155_new_n10435_), .Y(u2__abc_52155_new_n10436_));
AND2X2 AND2X2_4251 ( .A(u2__abc_52155_new_n10437_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__142_));
AND2X2 AND2X2_4252 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_143_), .Y(u2__abc_52155_new_n10439_));
AND2X2 AND2X2_4253 ( .A(u2__abc_52155_new_n10426_), .B(u2__abc_52155_new_n5203_), .Y(u2__abc_52155_new_n10440_));
AND2X2 AND2X2_4254 ( .A(u2__abc_52155_new_n10440_), .B(u2__abc_52155_new_n5214_), .Y(u2__abc_52155_new_n10441_));
AND2X2 AND2X2_4255 ( .A(u2__abc_52155_new_n10443_), .B(u2__abc_52155_new_n10442_), .Y(u2__abc_52155_new_n10444_));
AND2X2 AND2X2_4256 ( .A(u2__abc_52155_new_n10445_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10446_));
AND2X2 AND2X2_4257 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_141_), .Y(u2__abc_52155_new_n10447_));
AND2X2 AND2X2_4258 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5158_), .Y(u2__abc_52155_new_n10450_));
AND2X2 AND2X2_4259 ( .A(u2__abc_52155_new_n10451_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10452_));
AND2X2 AND2X2_426 ( .A(u1__abc_51895_new_n203_), .B(u1__abc_51895_new_n210_), .Y(u1__abc_51895_new_n211_));
AND2X2 AND2X2_4260 ( .A(u2__abc_52155_new_n10449_), .B(u2__abc_52155_new_n10452_), .Y(u2__abc_52155_new_n10453_));
AND2X2 AND2X2_4261 ( .A(u2__abc_52155_new_n10454_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__143_));
AND2X2 AND2X2_4262 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_144_), .Y(u2__abc_52155_new_n10456_));
AND2X2 AND2X2_4263 ( .A(u2__abc_52155_new_n10309_), .B(u2__abc_52155_new_n5232_), .Y(u2__abc_52155_new_n10457_));
AND2X2 AND2X2_4264 ( .A(u2__abc_52155_new_n10386_), .B(u2__abc_52155_new_n5231_), .Y(u2__abc_52155_new_n10458_));
AND2X2 AND2X2_4265 ( .A(u2__abc_52155_new_n10460_), .B(u2__abc_52155_new_n5215_), .Y(u2__abc_52155_new_n10461_));
AND2X2 AND2X2_4266 ( .A(u2__abc_52155_new_n5213_), .B(u2__abc_52155_new_n5202_), .Y(u2__abc_52155_new_n10462_));
AND2X2 AND2X2_4267 ( .A(u2__abc_52155_new_n10150_), .B(u2__abc_52155_new_n5284_), .Y(u2__abc_52155_new_n10467_));
AND2X2 AND2X2_4268 ( .A(u2__abc_52155_new_n10468_), .B(u2__abc_52155_new_n5168_), .Y(u2__abc_52155_new_n10469_));
AND2X2 AND2X2_4269 ( .A(u2__abc_52155_new_n10470_), .B(u2__abc_52155_new_n10471_), .Y(u2__abc_52155_new_n10472_));
AND2X2 AND2X2_427 ( .A(u1__abc_51895_new_n212_), .B(u1__abc_51895_new_n213_), .Y(u1__abc_51895_new_n214_));
AND2X2 AND2X2_4270 ( .A(u2__abc_52155_new_n10472_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10473_));
AND2X2 AND2X2_4271 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_142_), .Y(u2__abc_52155_new_n10474_));
AND2X2 AND2X2_4272 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5145_), .Y(u2__abc_52155_new_n10477_));
AND2X2 AND2X2_4273 ( .A(u2__abc_52155_new_n10478_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10479_));
AND2X2 AND2X2_4274 ( .A(u2__abc_52155_new_n10476_), .B(u2__abc_52155_new_n10479_), .Y(u2__abc_52155_new_n10480_));
AND2X2 AND2X2_4275 ( .A(u2__abc_52155_new_n10481_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__144_));
AND2X2 AND2X2_4276 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_145_), .Y(u2__abc_52155_new_n10483_));
AND2X2 AND2X2_4277 ( .A(u2__abc_52155_new_n10470_), .B(u2__abc_52155_new_n5164_), .Y(u2__abc_52155_new_n10485_));
AND2X2 AND2X2_4278 ( .A(u2__abc_52155_new_n10486_), .B(u2__abc_52155_new_n10484_), .Y(u2__abc_52155_new_n10487_));
AND2X2 AND2X2_4279 ( .A(u2__abc_52155_new_n10485_), .B(u2__abc_52155_new_n5161_), .Y(u2__abc_52155_new_n10488_));
AND2X2 AND2X2_428 ( .A(u1__abc_51895_new_n215_), .B(u1__abc_51895_new_n216_), .Y(u1__abc_51895_new_n217_));
AND2X2 AND2X2_4280 ( .A(u2__abc_52155_new_n10489_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10490_));
AND2X2 AND2X2_4281 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_143_), .Y(u2__abc_52155_new_n10491_));
AND2X2 AND2X2_4282 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5150_), .Y(u2__abc_52155_new_n10494_));
AND2X2 AND2X2_4283 ( .A(u2__abc_52155_new_n10495_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10496_));
AND2X2 AND2X2_4284 ( .A(u2__abc_52155_new_n10493_), .B(u2__abc_52155_new_n10496_), .Y(u2__abc_52155_new_n10497_));
AND2X2 AND2X2_4285 ( .A(u2__abc_52155_new_n10498_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__145_));
AND2X2 AND2X2_4286 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_146_), .Y(u2__abc_52155_new_n10500_));
AND2X2 AND2X2_4287 ( .A(u2__abc_52155_new_n10486_), .B(u2__abc_52155_new_n5160_), .Y(u2__abc_52155_new_n10502_));
AND2X2 AND2X2_4288 ( .A(u2__abc_52155_new_n10503_), .B(u2__abc_52155_new_n10501_), .Y(u2__abc_52155_new_n10504_));
AND2X2 AND2X2_4289 ( .A(u2__abc_52155_new_n10506_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10507_));
AND2X2 AND2X2_429 ( .A(u1__abc_51895_new_n214_), .B(u1__abc_51895_new_n217_), .Y(u1__abc_51895_new_n218_));
AND2X2 AND2X2_4290 ( .A(u2__abc_52155_new_n10507_), .B(u2__abc_52155_new_n10505_), .Y(u2__abc_52155_new_n10508_));
AND2X2 AND2X2_4291 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_144_), .Y(u2__abc_52155_new_n10509_));
AND2X2 AND2X2_4292 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5137_), .Y(u2__abc_52155_new_n10512_));
AND2X2 AND2X2_4293 ( .A(u2__abc_52155_new_n10513_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10514_));
AND2X2 AND2X2_4294 ( .A(u2__abc_52155_new_n10511_), .B(u2__abc_52155_new_n10514_), .Y(u2__abc_52155_new_n10515_));
AND2X2 AND2X2_4295 ( .A(u2__abc_52155_new_n10516_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__146_));
AND2X2 AND2X2_4296 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_147_), .Y(u2__abc_52155_new_n10518_));
AND2X2 AND2X2_4297 ( .A(u2__abc_52155_new_n10505_), .B(u2__abc_52155_new_n10519_), .Y(u2__abc_52155_new_n10520_));
AND2X2 AND2X2_4298 ( .A(u2__abc_52155_new_n10524_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10525_));
AND2X2 AND2X2_4299 ( .A(u2__abc_52155_new_n10525_), .B(u2__abc_52155_new_n10521_), .Y(u2__abc_52155_new_n10526_));
AND2X2 AND2X2_43 ( .A(_abc_73687_new_n753_), .B(sqrto_42_), .Y(\o[78] ));
AND2X2 AND2X2_430 ( .A(u1__abc_51895_new_n219_), .B(u1__abc_51895_new_n220_), .Y(u1__abc_51895_new_n221_));
AND2X2 AND2X2_4300 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_145_), .Y(u2__abc_52155_new_n10527_));
AND2X2 AND2X2_4301 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5130_), .Y(u2__abc_52155_new_n10530_));
AND2X2 AND2X2_4302 ( .A(u2__abc_52155_new_n10531_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10532_));
AND2X2 AND2X2_4303 ( .A(u2__abc_52155_new_n10529_), .B(u2__abc_52155_new_n10532_), .Y(u2__abc_52155_new_n10533_));
AND2X2 AND2X2_4304 ( .A(u2__abc_52155_new_n10534_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__147_));
AND2X2 AND2X2_4305 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_148_), .Y(u2__abc_52155_new_n10536_));
AND2X2 AND2X2_4306 ( .A(u2__abc_52155_new_n10519_), .B(u2__abc_52155_new_n5340_), .Y(u2__abc_52155_new_n10537_));
AND2X2 AND2X2_4307 ( .A(u2__abc_52155_new_n10505_), .B(u2__abc_52155_new_n10537_), .Y(u2__abc_52155_new_n10538_));
AND2X2 AND2X2_4308 ( .A(u2__abc_52155_new_n10540_), .B(u2__abc_52155_new_n5140_), .Y(u2__abc_52155_new_n10541_));
AND2X2 AND2X2_4309 ( .A(u2__abc_52155_new_n10543_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10544_));
AND2X2 AND2X2_431 ( .A(u1__abc_51895_new_n222_), .B(u1__abc_51895_new_n223_), .Y(u1__abc_51895_new_n224_));
AND2X2 AND2X2_4310 ( .A(u2__abc_52155_new_n10544_), .B(u2__abc_52155_new_n10542_), .Y(u2__abc_52155_new_n10545_));
AND2X2 AND2X2_4311 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_146_), .Y(u2__abc_52155_new_n10546_));
AND2X2 AND2X2_4312 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5115_), .Y(u2__abc_52155_new_n10549_));
AND2X2 AND2X2_4313 ( .A(u2__abc_52155_new_n10550_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10551_));
AND2X2 AND2X2_4314 ( .A(u2__abc_52155_new_n10548_), .B(u2__abc_52155_new_n10551_), .Y(u2__abc_52155_new_n10552_));
AND2X2 AND2X2_4315 ( .A(u2__abc_52155_new_n10553_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__148_));
AND2X2 AND2X2_4316 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_149_), .Y(u2__abc_52155_new_n10555_));
AND2X2 AND2X2_4317 ( .A(u2__abc_52155_new_n10542_), .B(u2__abc_52155_new_n5136_), .Y(u2__abc_52155_new_n10556_));
AND2X2 AND2X2_4318 ( .A(u2__abc_52155_new_n10557_), .B(u2__abc_52155_new_n5133_), .Y(u2__abc_52155_new_n10558_));
AND2X2 AND2X2_4319 ( .A(u2__abc_52155_new_n10560_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10561_));
AND2X2 AND2X2_432 ( .A(u1__abc_51895_new_n221_), .B(u1__abc_51895_new_n224_), .Y(u1__abc_51895_new_n225_));
AND2X2 AND2X2_4320 ( .A(u2__abc_52155_new_n10561_), .B(u2__abc_52155_new_n10559_), .Y(u2__abc_52155_new_n10562_));
AND2X2 AND2X2_4321 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_147_), .Y(u2__abc_52155_new_n10563_));
AND2X2 AND2X2_4322 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5122_), .Y(u2__abc_52155_new_n10566_));
AND2X2 AND2X2_4323 ( .A(u2__abc_52155_new_n10567_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10568_));
AND2X2 AND2X2_4324 ( .A(u2__abc_52155_new_n10565_), .B(u2__abc_52155_new_n10568_), .Y(u2__abc_52155_new_n10569_));
AND2X2 AND2X2_4325 ( .A(u2__abc_52155_new_n10570_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__149_));
AND2X2 AND2X2_4326 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_150_), .Y(u2__abc_52155_new_n10572_));
AND2X2 AND2X2_4327 ( .A(u2__abc_52155_new_n10559_), .B(u2__abc_52155_new_n5129_), .Y(u2__abc_52155_new_n10573_));
AND2X2 AND2X2_4328 ( .A(u2__abc_52155_new_n10574_), .B(u2__abc_52155_new_n5118_), .Y(u2__abc_52155_new_n10575_));
AND2X2 AND2X2_4329 ( .A(u2__abc_52155_new_n10577_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10578_));
AND2X2 AND2X2_433 ( .A(u1__abc_51895_new_n218_), .B(u1__abc_51895_new_n225_), .Y(u1__abc_51895_new_n226_));
AND2X2 AND2X2_4330 ( .A(u2__abc_52155_new_n10578_), .B(u2__abc_52155_new_n10576_), .Y(u2__abc_52155_new_n10579_));
AND2X2 AND2X2_4331 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_148_), .Y(u2__abc_52155_new_n10580_));
AND2X2 AND2X2_4332 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5074_), .Y(u2__abc_52155_new_n10583_));
AND2X2 AND2X2_4333 ( .A(u2__abc_52155_new_n10584_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10585_));
AND2X2 AND2X2_4334 ( .A(u2__abc_52155_new_n10582_), .B(u2__abc_52155_new_n10585_), .Y(u2__abc_52155_new_n10586_));
AND2X2 AND2X2_4335 ( .A(u2__abc_52155_new_n10587_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__150_));
AND2X2 AND2X2_4336 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_151_), .Y(u2__abc_52155_new_n10589_));
AND2X2 AND2X2_4337 ( .A(u2__abc_52155_new_n10576_), .B(u2__abc_52155_new_n5114_), .Y(u2__abc_52155_new_n10590_));
AND2X2 AND2X2_4338 ( .A(u2__abc_52155_new_n10590_), .B(u2__abc_52155_new_n5125_), .Y(u2__abc_52155_new_n10591_));
AND2X2 AND2X2_4339 ( .A(u2__abc_52155_new_n10593_), .B(u2__abc_52155_new_n10592_), .Y(u2__abc_52155_new_n10594_));
AND2X2 AND2X2_434 ( .A(u1__abc_51895_new_n211_), .B(u1__abc_51895_new_n226_), .Y(u1__abc_51895_new_n227_));
AND2X2 AND2X2_4340 ( .A(u2__abc_52155_new_n10595_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10596_));
AND2X2 AND2X2_4341 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_149_), .Y(u2__abc_52155_new_n10597_));
AND2X2 AND2X2_4342 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5067_), .Y(u2__abc_52155_new_n10600_));
AND2X2 AND2X2_4343 ( .A(u2__abc_52155_new_n10601_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10602_));
AND2X2 AND2X2_4344 ( .A(u2__abc_52155_new_n10599_), .B(u2__abc_52155_new_n10602_), .Y(u2__abc_52155_new_n10603_));
AND2X2 AND2X2_4345 ( .A(u2__abc_52155_new_n10604_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__151_));
AND2X2 AND2X2_4346 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_152_), .Y(u2__abc_52155_new_n10606_));
AND2X2 AND2X2_4347 ( .A(u2__abc_52155_new_n5157_), .B(u2__abc_52155_new_n5164_), .Y(u2__abc_52155_new_n10608_));
AND2X2 AND2X2_4348 ( .A(u2__abc_52155_new_n10610_), .B(u2__abc_52155_new_n10607_), .Y(u2__abc_52155_new_n10611_));
AND2X2 AND2X2_4349 ( .A(u2__abc_52155_new_n5129_), .B(u2__abc_52155_new_n5136_), .Y(u2__abc_52155_new_n10613_));
AND2X2 AND2X2_435 ( .A(u1__abc_51895_new_n228_), .B(u1__abc_51895_new_n229_), .Y(u1__abc_51895_new_n230_));
AND2X2 AND2X2_4350 ( .A(u2__abc_52155_new_n10612_), .B(u2__abc_52155_new_n10613_), .Y(u2__abc_52155_new_n10614_));
AND2X2 AND2X2_4351 ( .A(u2__abc_52155_new_n10616_), .B(u2__abc_52155_new_n5114_), .Y(u2__abc_52155_new_n10617_));
AND2X2 AND2X2_4352 ( .A(u2__abc_52155_new_n10618_), .B(u2__abc_52155_new_n5121_), .Y(u2__abc_52155_new_n10619_));
AND2X2 AND2X2_4353 ( .A(u2__abc_52155_new_n10468_), .B(u2__abc_52155_new_n5171_), .Y(u2__abc_52155_new_n10621_));
AND2X2 AND2X2_4354 ( .A(u2__abc_52155_new_n10622_), .B(u2__abc_52155_new_n5077_), .Y(u2__abc_52155_new_n10623_));
AND2X2 AND2X2_4355 ( .A(u2__abc_52155_new_n10625_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10626_));
AND2X2 AND2X2_4356 ( .A(u2__abc_52155_new_n10626_), .B(u2__abc_52155_new_n10624_), .Y(u2__abc_52155_new_n10627_));
AND2X2 AND2X2_4357 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_150_), .Y(u2__abc_52155_new_n10628_));
AND2X2 AND2X2_4358 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5052_), .Y(u2__abc_52155_new_n10631_));
AND2X2 AND2X2_4359 ( .A(u2__abc_52155_new_n10632_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10633_));
AND2X2 AND2X2_436 ( .A(u1__abc_51895_new_n231_), .B(u1__abc_51895_new_n232_), .Y(u1__abc_51895_new_n233_));
AND2X2 AND2X2_4360 ( .A(u2__abc_52155_new_n10630_), .B(u2__abc_52155_new_n10633_), .Y(u2__abc_52155_new_n10634_));
AND2X2 AND2X2_4361 ( .A(u2__abc_52155_new_n10635_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__152_));
AND2X2 AND2X2_4362 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_153_), .Y(u2__abc_52155_new_n10637_));
AND2X2 AND2X2_4363 ( .A(u2__abc_52155_new_n10624_), .B(u2__abc_52155_new_n5073_), .Y(u2__abc_52155_new_n10638_));
AND2X2 AND2X2_4364 ( .A(u2__abc_52155_new_n10638_), .B(u2__abc_52155_new_n5070_), .Y(u2__abc_52155_new_n10639_));
AND2X2 AND2X2_4365 ( .A(u2__abc_52155_new_n10641_), .B(u2__abc_52155_new_n10640_), .Y(u2__abc_52155_new_n10642_));
AND2X2 AND2X2_4366 ( .A(u2__abc_52155_new_n10643_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10644_));
AND2X2 AND2X2_4367 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_151_), .Y(u2__abc_52155_new_n10645_));
AND2X2 AND2X2_4368 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5059_), .Y(u2__abc_52155_new_n10648_));
AND2X2 AND2X2_4369 ( .A(u2__abc_52155_new_n10649_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10650_));
AND2X2 AND2X2_437 ( .A(u1__abc_51895_new_n230_), .B(u1__abc_51895_new_n233_), .Y(u1__abc_51895_new_n234_));
AND2X2 AND2X2_4370 ( .A(u2__abc_52155_new_n10647_), .B(u2__abc_52155_new_n10650_), .Y(u2__abc_52155_new_n10651_));
AND2X2 AND2X2_4371 ( .A(u2__abc_52155_new_n10652_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__153_));
AND2X2 AND2X2_4372 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_154_), .Y(u2__abc_52155_new_n10654_));
AND2X2 AND2X2_4373 ( .A(u2__abc_52155_new_n5066_), .B(u2__abc_52155_new_n5073_), .Y(u2__abc_52155_new_n10655_));
AND2X2 AND2X2_4374 ( .A(u2__abc_52155_new_n10624_), .B(u2__abc_52155_new_n10655_), .Y(u2__abc_52155_new_n10656_));
AND2X2 AND2X2_4375 ( .A(u2__abc_52155_new_n10658_), .B(u2__abc_52155_new_n5055_), .Y(u2__abc_52155_new_n10659_));
AND2X2 AND2X2_4376 ( .A(u2__abc_52155_new_n10661_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10662_));
AND2X2 AND2X2_4377 ( .A(u2__abc_52155_new_n10662_), .B(u2__abc_52155_new_n10660_), .Y(u2__abc_52155_new_n10663_));
AND2X2 AND2X2_4378 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_152_), .Y(u2__abc_52155_new_n10664_));
AND2X2 AND2X2_4379 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5105_), .Y(u2__abc_52155_new_n10667_));
AND2X2 AND2X2_438 ( .A(u1__abc_51895_new_n235_), .B(u1__abc_51895_new_n236_), .Y(u1__abc_51895_new_n237_));
AND2X2 AND2X2_4380 ( .A(u2__abc_52155_new_n10668_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10669_));
AND2X2 AND2X2_4381 ( .A(u2__abc_52155_new_n10666_), .B(u2__abc_52155_new_n10669_), .Y(u2__abc_52155_new_n10670_));
AND2X2 AND2X2_4382 ( .A(u2__abc_52155_new_n10671_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__154_));
AND2X2 AND2X2_4383 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_155_), .Y(u2__abc_52155_new_n10673_));
AND2X2 AND2X2_4384 ( .A(u2__abc_52155_new_n10660_), .B(u2__abc_52155_new_n5051_), .Y(u2__abc_52155_new_n10674_));
AND2X2 AND2X2_4385 ( .A(u2__abc_52155_new_n10674_), .B(u2__abc_52155_new_n5062_), .Y(u2__abc_52155_new_n10675_));
AND2X2 AND2X2_4386 ( .A(u2__abc_52155_new_n10677_), .B(u2__abc_52155_new_n10676_), .Y(u2__abc_52155_new_n10678_));
AND2X2 AND2X2_4387 ( .A(u2__abc_52155_new_n10679_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10680_));
AND2X2 AND2X2_4388 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_153_), .Y(u2__abc_52155_new_n10681_));
AND2X2 AND2X2_4389 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5098_), .Y(u2__abc_52155_new_n10684_));
AND2X2 AND2X2_439 ( .A(u1__abc_51895_new_n238_), .B(u1__abc_51895_new_n239_), .Y(u1__abc_51895_new_n240_));
AND2X2 AND2X2_4390 ( .A(u2__abc_52155_new_n10685_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10686_));
AND2X2 AND2X2_4391 ( .A(u2__abc_52155_new_n10683_), .B(u2__abc_52155_new_n10686_), .Y(u2__abc_52155_new_n10687_));
AND2X2 AND2X2_4392 ( .A(u2__abc_52155_new_n10688_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__155_));
AND2X2 AND2X2_4393 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_156_), .Y(u2__abc_52155_new_n10690_));
AND2X2 AND2X2_4394 ( .A(u2__abc_52155_new_n10692_), .B(u2__abc_52155_new_n5063_), .Y(u2__abc_52155_new_n10693_));
AND2X2 AND2X2_4395 ( .A(u2__abc_52155_new_n5061_), .B(u2__abc_52155_new_n5050_), .Y(u2__abc_52155_new_n10694_));
AND2X2 AND2X2_4396 ( .A(u2__abc_52155_new_n10622_), .B(u2__abc_52155_new_n5079_), .Y(u2__abc_52155_new_n10697_));
AND2X2 AND2X2_4397 ( .A(u2__abc_52155_new_n10698_), .B(u2__abc_52155_new_n5108_), .Y(u2__abc_52155_new_n10699_));
AND2X2 AND2X2_4398 ( .A(u2__abc_52155_new_n10701_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10702_));
AND2X2 AND2X2_4399 ( .A(u2__abc_52155_new_n10702_), .B(u2__abc_52155_new_n10700_), .Y(u2__abc_52155_new_n10703_));
AND2X2 AND2X2_44 ( .A(_abc_73687_new_n753_), .B(sqrto_43_), .Y(\o[79] ));
AND2X2 AND2X2_440 ( .A(u1__abc_51895_new_n237_), .B(u1__abc_51895_new_n240_), .Y(u1__abc_51895_new_n241_));
AND2X2 AND2X2_4400 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_154_), .Y(u2__abc_52155_new_n10704_));
AND2X2 AND2X2_4401 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5083_), .Y(u2__abc_52155_new_n10707_));
AND2X2 AND2X2_4402 ( .A(u2__abc_52155_new_n10708_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10709_));
AND2X2 AND2X2_4403 ( .A(u2__abc_52155_new_n10706_), .B(u2__abc_52155_new_n10709_), .Y(u2__abc_52155_new_n10710_));
AND2X2 AND2X2_4404 ( .A(u2__abc_52155_new_n10711_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__156_));
AND2X2 AND2X2_4405 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_157_), .Y(u2__abc_52155_new_n10713_));
AND2X2 AND2X2_4406 ( .A(u2__abc_52155_new_n10700_), .B(u2__abc_52155_new_n5104_), .Y(u2__abc_52155_new_n10714_));
AND2X2 AND2X2_4407 ( .A(u2__abc_52155_new_n10714_), .B(u2__abc_52155_new_n5101_), .Y(u2__abc_52155_new_n10715_));
AND2X2 AND2X2_4408 ( .A(u2__abc_52155_new_n10717_), .B(u2__abc_52155_new_n10716_), .Y(u2__abc_52155_new_n10718_));
AND2X2 AND2X2_4409 ( .A(u2__abc_52155_new_n10719_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10720_));
AND2X2 AND2X2_441 ( .A(u1__abc_51895_new_n234_), .B(u1__abc_51895_new_n241_), .Y(u1__abc_51895_new_n242_));
AND2X2 AND2X2_4410 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_155_), .Y(u2__abc_52155_new_n10721_));
AND2X2 AND2X2_4411 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5090_), .Y(u2__abc_52155_new_n10724_));
AND2X2 AND2X2_4412 ( .A(u2__abc_52155_new_n10725_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10726_));
AND2X2 AND2X2_4413 ( .A(u2__abc_52155_new_n10723_), .B(u2__abc_52155_new_n10726_), .Y(u2__abc_52155_new_n10727_));
AND2X2 AND2X2_4414 ( .A(u2__abc_52155_new_n10728_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__157_));
AND2X2 AND2X2_4415 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_158_), .Y(u2__abc_52155_new_n10730_));
AND2X2 AND2X2_4416 ( .A(u2__abc_52155_new_n5097_), .B(u2__abc_52155_new_n5104_), .Y(u2__abc_52155_new_n10731_));
AND2X2 AND2X2_4417 ( .A(u2__abc_52155_new_n10700_), .B(u2__abc_52155_new_n10731_), .Y(u2__abc_52155_new_n10732_));
AND2X2 AND2X2_4418 ( .A(u2__abc_52155_new_n10734_), .B(u2__abc_52155_new_n5086_), .Y(u2__abc_52155_new_n10735_));
AND2X2 AND2X2_4419 ( .A(u2__abc_52155_new_n10737_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10738_));
AND2X2 AND2X2_442 ( .A(u1__abc_51895_new_n243_), .B(u1__abc_51895_new_n244_), .Y(u1__abc_51895_new_n245_));
AND2X2 AND2X2_4420 ( .A(u2__abc_52155_new_n10738_), .B(u2__abc_52155_new_n10736_), .Y(u2__abc_52155_new_n10739_));
AND2X2 AND2X2_4421 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_156_), .Y(u2__abc_52155_new_n10740_));
AND2X2 AND2X2_4422 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5009_), .Y(u2__abc_52155_new_n10743_));
AND2X2 AND2X2_4423 ( .A(u2__abc_52155_new_n10744_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10745_));
AND2X2 AND2X2_4424 ( .A(u2__abc_52155_new_n10742_), .B(u2__abc_52155_new_n10745_), .Y(u2__abc_52155_new_n10746_));
AND2X2 AND2X2_4425 ( .A(u2__abc_52155_new_n10747_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__158_));
AND2X2 AND2X2_4426 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_159_), .Y(u2__abc_52155_new_n10749_));
AND2X2 AND2X2_4427 ( .A(u2__abc_52155_new_n10736_), .B(u2__abc_52155_new_n5082_), .Y(u2__abc_52155_new_n10750_));
AND2X2 AND2X2_4428 ( .A(u2__abc_52155_new_n10750_), .B(u2__abc_52155_new_n5093_), .Y(u2__abc_52155_new_n10751_));
AND2X2 AND2X2_4429 ( .A(u2__abc_52155_new_n10753_), .B(u2__abc_52155_new_n10752_), .Y(u2__abc_52155_new_n10754_));
AND2X2 AND2X2_443 ( .A(u1__abc_51895_new_n246_), .B(u1__abc_51895_new_n247_), .Y(u1__abc_51895_new_n248_));
AND2X2 AND2X2_4430 ( .A(u2__abc_52155_new_n10755_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10756_));
AND2X2 AND2X2_4431 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_157_), .Y(u2__abc_52155_new_n10757_));
AND2X2 AND2X2_4432 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5002_), .Y(u2__abc_52155_new_n10760_));
AND2X2 AND2X2_4433 ( .A(u2__abc_52155_new_n10761_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10762_));
AND2X2 AND2X2_4434 ( .A(u2__abc_52155_new_n10759_), .B(u2__abc_52155_new_n10762_), .Y(u2__abc_52155_new_n10763_));
AND2X2 AND2X2_4435 ( .A(u2__abc_52155_new_n10764_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__159_));
AND2X2 AND2X2_4436 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_160_), .Y(u2__abc_52155_new_n10766_));
AND2X2 AND2X2_4437 ( .A(u2__abc_52155_new_n10620_), .B(u2__abc_52155_new_n5111_), .Y(u2__abc_52155_new_n10767_));
AND2X2 AND2X2_4438 ( .A(u2__abc_52155_new_n10466_), .B(u2__abc_52155_new_n5172_), .Y(u2__abc_52155_new_n10768_));
AND2X2 AND2X2_4439 ( .A(u2__abc_52155_new_n10696_), .B(u2__abc_52155_new_n5110_), .Y(u2__abc_52155_new_n10769_));
AND2X2 AND2X2_444 ( .A(u1__abc_51895_new_n245_), .B(u1__abc_51895_new_n248_), .Y(u1__abc_51895_new_n249_));
AND2X2 AND2X2_4440 ( .A(u2__abc_52155_new_n10771_), .B(u2__abc_52155_new_n5094_), .Y(u2__abc_52155_new_n10772_));
AND2X2 AND2X2_4441 ( .A(u2__abc_52155_new_n5092_), .B(u2__abc_52155_new_n5081_), .Y(u2__abc_52155_new_n10773_));
AND2X2 AND2X2_4442 ( .A(u2__abc_52155_new_n10150_), .B(u2__abc_52155_new_n5285_), .Y(u2__abc_52155_new_n10779_));
AND2X2 AND2X2_4443 ( .A(u2__abc_52155_new_n10780_), .B(u2__abc_52155_new_n5012_), .Y(u2__abc_52155_new_n10781_));
AND2X2 AND2X2_4444 ( .A(u2__abc_52155_new_n10782_), .B(u2__abc_52155_new_n10783_), .Y(u2__abc_52155_new_n10784_));
AND2X2 AND2X2_4445 ( .A(u2__abc_52155_new_n10784_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10785_));
AND2X2 AND2X2_4446 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_158_), .Y(u2__abc_52155_new_n10786_));
AND2X2 AND2X2_4447 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4989_), .Y(u2__abc_52155_new_n10789_));
AND2X2 AND2X2_4448 ( .A(u2__abc_52155_new_n10790_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10791_));
AND2X2 AND2X2_4449 ( .A(u2__abc_52155_new_n10788_), .B(u2__abc_52155_new_n10791_), .Y(u2__abc_52155_new_n10792_));
AND2X2 AND2X2_445 ( .A(u1__abc_51895_new_n250_), .B(u1__abc_51895_new_n251_), .Y(u1__abc_51895_new_n252_));
AND2X2 AND2X2_4450 ( .A(u2__abc_52155_new_n10793_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__160_));
AND2X2 AND2X2_4451 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_161_), .Y(u2__abc_52155_new_n10795_));
AND2X2 AND2X2_4452 ( .A(u2__abc_52155_new_n10782_), .B(u2__abc_52155_new_n5008_), .Y(u2__abc_52155_new_n10796_));
AND2X2 AND2X2_4453 ( .A(u2__abc_52155_new_n10796_), .B(u2__abc_52155_new_n5005_), .Y(u2__abc_52155_new_n10797_));
AND2X2 AND2X2_4454 ( .A(u2__abc_52155_new_n10799_), .B(u2__abc_52155_new_n10798_), .Y(u2__abc_52155_new_n10800_));
AND2X2 AND2X2_4455 ( .A(u2__abc_52155_new_n10801_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10802_));
AND2X2 AND2X2_4456 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_159_), .Y(u2__abc_52155_new_n10803_));
AND2X2 AND2X2_4457 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4994_), .Y(u2__abc_52155_new_n10806_));
AND2X2 AND2X2_4458 ( .A(u2__abc_52155_new_n10807_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10808_));
AND2X2 AND2X2_4459 ( .A(u2__abc_52155_new_n10805_), .B(u2__abc_52155_new_n10808_), .Y(u2__abc_52155_new_n10809_));
AND2X2 AND2X2_446 ( .A(u1__abc_51895_new_n253_), .B(u1__abc_51895_new_n254_), .Y(u1__abc_51895_new_n255_));
AND2X2 AND2X2_4460 ( .A(u2__abc_52155_new_n10810_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__161_));
AND2X2 AND2X2_4461 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_162_), .Y(u2__abc_52155_new_n10812_));
AND2X2 AND2X2_4462 ( .A(u2__abc_52155_new_n5001_), .B(u2__abc_52155_new_n5008_), .Y(u2__abc_52155_new_n10814_));
AND2X2 AND2X2_4463 ( .A(u2__abc_52155_new_n10782_), .B(u2__abc_52155_new_n10814_), .Y(u2__abc_52155_new_n10815_));
AND2X2 AND2X2_4464 ( .A(u2__abc_52155_new_n10817_), .B(u2__abc_52155_new_n10813_), .Y(u2__abc_52155_new_n10818_));
AND2X2 AND2X2_4465 ( .A(u2__abc_52155_new_n10820_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10821_));
AND2X2 AND2X2_4466 ( .A(u2__abc_52155_new_n10821_), .B(u2__abc_52155_new_n10819_), .Y(u2__abc_52155_new_n10822_));
AND2X2 AND2X2_4467 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_160_), .Y(u2__abc_52155_new_n10823_));
AND2X2 AND2X2_4468 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5040_), .Y(u2__abc_52155_new_n10826_));
AND2X2 AND2X2_4469 ( .A(u2__abc_52155_new_n10827_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10828_));
AND2X2 AND2X2_447 ( .A(u1__abc_51895_new_n252_), .B(u1__abc_51895_new_n255_), .Y(u1__abc_51895_new_n256_));
AND2X2 AND2X2_4470 ( .A(u2__abc_52155_new_n10825_), .B(u2__abc_52155_new_n10828_), .Y(u2__abc_52155_new_n10829_));
AND2X2 AND2X2_4471 ( .A(u2__abc_52155_new_n10830_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__162_));
AND2X2 AND2X2_4472 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_163_), .Y(u2__abc_52155_new_n10832_));
AND2X2 AND2X2_4473 ( .A(u2__abc_52155_new_n10819_), .B(u2__abc_52155_new_n10833_), .Y(u2__abc_52155_new_n10834_));
AND2X2 AND2X2_4474 ( .A(u2__abc_52155_new_n10838_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10839_));
AND2X2 AND2X2_4475 ( .A(u2__abc_52155_new_n10839_), .B(u2__abc_52155_new_n10835_), .Y(u2__abc_52155_new_n10840_));
AND2X2 AND2X2_4476 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_161_), .Y(u2__abc_52155_new_n10841_));
AND2X2 AND2X2_4477 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5033_), .Y(u2__abc_52155_new_n10844_));
AND2X2 AND2X2_4478 ( .A(u2__abc_52155_new_n10845_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10846_));
AND2X2 AND2X2_4479 ( .A(u2__abc_52155_new_n10843_), .B(u2__abc_52155_new_n10846_), .Y(u2__abc_52155_new_n10847_));
AND2X2 AND2X2_448 ( .A(u1__abc_51895_new_n249_), .B(u1__abc_51895_new_n256_), .Y(u1__abc_51895_new_n257_));
AND2X2 AND2X2_4480 ( .A(u2__abc_52155_new_n10848_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__163_));
AND2X2 AND2X2_4481 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_164_), .Y(u2__abc_52155_new_n10850_));
AND2X2 AND2X2_4482 ( .A(u2__abc_52155_new_n10853_), .B(u2__abc_52155_new_n5379_), .Y(u2__abc_52155_new_n10854_));
AND2X2 AND2X2_4483 ( .A(u2__abc_52155_new_n10852_), .B(u2__abc_52155_new_n10854_), .Y(u2__abc_52155_new_n10855_));
AND2X2 AND2X2_4484 ( .A(u2__abc_52155_new_n10780_), .B(u2__abc_52155_new_n5014_), .Y(u2__abc_52155_new_n10857_));
AND2X2 AND2X2_4485 ( .A(u2__abc_52155_new_n10858_), .B(u2__abc_52155_new_n5043_), .Y(u2__abc_52155_new_n10859_));
AND2X2 AND2X2_4486 ( .A(u2__abc_52155_new_n10861_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10862_));
AND2X2 AND2X2_4487 ( .A(u2__abc_52155_new_n10862_), .B(u2__abc_52155_new_n10860_), .Y(u2__abc_52155_new_n10863_));
AND2X2 AND2X2_4488 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_162_), .Y(u2__abc_52155_new_n10864_));
AND2X2 AND2X2_4489 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5018_), .Y(u2__abc_52155_new_n10867_));
AND2X2 AND2X2_449 ( .A(u1__abc_51895_new_n242_), .B(u1__abc_51895_new_n257_), .Y(u1__abc_51895_new_n258_));
AND2X2 AND2X2_4490 ( .A(u2__abc_52155_new_n10868_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10869_));
AND2X2 AND2X2_4491 ( .A(u2__abc_52155_new_n10866_), .B(u2__abc_52155_new_n10869_), .Y(u2__abc_52155_new_n10870_));
AND2X2 AND2X2_4492 ( .A(u2__abc_52155_new_n10871_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__164_));
AND2X2 AND2X2_4493 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_165_), .Y(u2__abc_52155_new_n10873_));
AND2X2 AND2X2_4494 ( .A(u2__abc_52155_new_n10860_), .B(u2__abc_52155_new_n5039_), .Y(u2__abc_52155_new_n10874_));
AND2X2 AND2X2_4495 ( .A(u2__abc_52155_new_n10875_), .B(u2__abc_52155_new_n5036_), .Y(u2__abc_52155_new_n10876_));
AND2X2 AND2X2_4496 ( .A(u2__abc_52155_new_n10878_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10879_));
AND2X2 AND2X2_4497 ( .A(u2__abc_52155_new_n10879_), .B(u2__abc_52155_new_n10877_), .Y(u2__abc_52155_new_n10880_));
AND2X2 AND2X2_4498 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_163_), .Y(u2__abc_52155_new_n10881_));
AND2X2 AND2X2_4499 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5025_), .Y(u2__abc_52155_new_n10884_));
AND2X2 AND2X2_45 ( .A(_abc_73687_new_n753_), .B(sqrto_44_), .Y(\o[80] ));
AND2X2 AND2X2_450 ( .A(u1__abc_51895_new_n227_), .B(u1__abc_51895_new_n258_), .Y(u1__abc_51895_new_n259_));
AND2X2 AND2X2_4500 ( .A(u2__abc_52155_new_n10885_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10886_));
AND2X2 AND2X2_4501 ( .A(u2__abc_52155_new_n10883_), .B(u2__abc_52155_new_n10886_), .Y(u2__abc_52155_new_n10887_));
AND2X2 AND2X2_4502 ( .A(u2__abc_52155_new_n10888_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__165_));
AND2X2 AND2X2_4503 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_166_), .Y(u2__abc_52155_new_n10890_));
AND2X2 AND2X2_4504 ( .A(u2__abc_52155_new_n10877_), .B(u2__abc_52155_new_n5032_), .Y(u2__abc_52155_new_n10891_));
AND2X2 AND2X2_4505 ( .A(u2__abc_52155_new_n10892_), .B(u2__abc_52155_new_n5021_), .Y(u2__abc_52155_new_n10893_));
AND2X2 AND2X2_4506 ( .A(u2__abc_52155_new_n10895_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10896_));
AND2X2 AND2X2_4507 ( .A(u2__abc_52155_new_n10896_), .B(u2__abc_52155_new_n10894_), .Y(u2__abc_52155_new_n10897_));
AND2X2 AND2X2_4508 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_164_), .Y(u2__abc_52155_new_n10898_));
AND2X2 AND2X2_4509 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4980_), .Y(u2__abc_52155_new_n10901_));
AND2X2 AND2X2_451 ( .A(u1__abc_51895_new_n259_), .B(u1__abc_51895_new_n196_), .Y(u1__abc_51895_new_n260_));
AND2X2 AND2X2_4510 ( .A(u2__abc_52155_new_n10902_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10903_));
AND2X2 AND2X2_4511 ( .A(u2__abc_52155_new_n10900_), .B(u2__abc_52155_new_n10903_), .Y(u2__abc_52155_new_n10904_));
AND2X2 AND2X2_4512 ( .A(u2__abc_52155_new_n10905_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__166_));
AND2X2 AND2X2_4513 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_167_), .Y(u2__abc_52155_new_n10907_));
AND2X2 AND2X2_4514 ( .A(u2__abc_52155_new_n10894_), .B(u2__abc_52155_new_n5017_), .Y(u2__abc_52155_new_n10908_));
AND2X2 AND2X2_4515 ( .A(u2__abc_52155_new_n10908_), .B(u2__abc_52155_new_n5028_), .Y(u2__abc_52155_new_n10909_));
AND2X2 AND2X2_4516 ( .A(u2__abc_52155_new_n10911_), .B(u2__abc_52155_new_n10910_), .Y(u2__abc_52155_new_n10912_));
AND2X2 AND2X2_4517 ( .A(u2__abc_52155_new_n10913_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10914_));
AND2X2 AND2X2_4518 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_165_), .Y(u2__abc_52155_new_n10915_));
AND2X2 AND2X2_4519 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4973_), .Y(u2__abc_52155_new_n10918_));
AND2X2 AND2X2_452 ( .A(u1__abc_51895_new_n261_), .B(u1__abc_51895_new_n262_), .Y(u1__abc_51895_new_n263_));
AND2X2 AND2X2_4520 ( .A(u2__abc_52155_new_n10919_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10920_));
AND2X2 AND2X2_4521 ( .A(u2__abc_52155_new_n10917_), .B(u2__abc_52155_new_n10920_), .Y(u2__abc_52155_new_n10921_));
AND2X2 AND2X2_4522 ( .A(u2__abc_52155_new_n10922_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__167_));
AND2X2 AND2X2_4523 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_168_), .Y(u2__abc_52155_new_n10924_));
AND2X2 AND2X2_4524 ( .A(u2__abc_52155_new_n10856_), .B(u2__abc_52155_new_n5045_), .Y(u2__abc_52155_new_n10925_));
AND2X2 AND2X2_4525 ( .A(u2__abc_52155_new_n10926_), .B(u2__abc_52155_new_n5035_), .Y(u2__abc_52155_new_n10927_));
AND2X2 AND2X2_4526 ( .A(u2__abc_52155_new_n5029_), .B(u2__abc_52155_new_n10927_), .Y(u2__abc_52155_new_n10928_));
AND2X2 AND2X2_4527 ( .A(u2__abc_52155_new_n5027_), .B(u2__abc_52155_new_n5016_), .Y(u2__abc_52155_new_n10929_));
AND2X2 AND2X2_4528 ( .A(u2__abc_52155_new_n10780_), .B(u2__abc_52155_new_n5046_), .Y(u2__abc_52155_new_n10933_));
AND2X2 AND2X2_4529 ( .A(u2__abc_52155_new_n10934_), .B(u2__abc_52155_new_n4983_), .Y(u2__abc_52155_new_n10935_));
AND2X2 AND2X2_453 ( .A(u1__abc_51895_new_n264_), .B(u1__abc_51895_new_n265_), .Y(u1__abc_51895_new_n266_));
AND2X2 AND2X2_4530 ( .A(u2__abc_52155_new_n10937_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10938_));
AND2X2 AND2X2_4531 ( .A(u2__abc_52155_new_n10938_), .B(u2__abc_52155_new_n10936_), .Y(u2__abc_52155_new_n10939_));
AND2X2 AND2X2_4532 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_166_), .Y(u2__abc_52155_new_n10940_));
AND2X2 AND2X2_4533 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4958_), .Y(u2__abc_52155_new_n10943_));
AND2X2 AND2X2_4534 ( .A(u2__abc_52155_new_n10944_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10945_));
AND2X2 AND2X2_4535 ( .A(u2__abc_52155_new_n10942_), .B(u2__abc_52155_new_n10945_), .Y(u2__abc_52155_new_n10946_));
AND2X2 AND2X2_4536 ( .A(u2__abc_52155_new_n10947_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__168_));
AND2X2 AND2X2_4537 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_169_), .Y(u2__abc_52155_new_n10949_));
AND2X2 AND2X2_4538 ( .A(u2__abc_52155_new_n10936_), .B(u2__abc_52155_new_n4979_), .Y(u2__abc_52155_new_n10951_));
AND2X2 AND2X2_4539 ( .A(u2__abc_52155_new_n10952_), .B(u2__abc_52155_new_n10950_), .Y(u2__abc_52155_new_n10953_));
AND2X2 AND2X2_454 ( .A(u1__abc_51895_new_n263_), .B(u1__abc_51895_new_n266_), .Y(u1__abc_51895_new_n267_));
AND2X2 AND2X2_4540 ( .A(u2__abc_52155_new_n10951_), .B(u2__abc_52155_new_n4976_), .Y(u2__abc_52155_new_n10954_));
AND2X2 AND2X2_4541 ( .A(u2__abc_52155_new_n10955_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10956_));
AND2X2 AND2X2_4542 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_167_), .Y(u2__abc_52155_new_n10957_));
AND2X2 AND2X2_4543 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4965_), .Y(u2__abc_52155_new_n10960_));
AND2X2 AND2X2_4544 ( .A(u2__abc_52155_new_n10961_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10962_));
AND2X2 AND2X2_4545 ( .A(u2__abc_52155_new_n10959_), .B(u2__abc_52155_new_n10962_), .Y(u2__abc_52155_new_n10963_));
AND2X2 AND2X2_4546 ( .A(u2__abc_52155_new_n10964_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__169_));
AND2X2 AND2X2_4547 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_170_), .Y(u2__abc_52155_new_n10966_));
AND2X2 AND2X2_4548 ( .A(u2__abc_52155_new_n4972_), .B(u2__abc_52155_new_n4979_), .Y(u2__abc_52155_new_n10967_));
AND2X2 AND2X2_4549 ( .A(u2__abc_52155_new_n10934_), .B(u2__abc_52155_new_n4984_), .Y(u2__abc_52155_new_n10970_));
AND2X2 AND2X2_455 ( .A(u1__abc_51895_new_n268_), .B(u1__abc_51895_new_n269_), .Y(u1__abc_51895_new_n270_));
AND2X2 AND2X2_4550 ( .A(u2__abc_52155_new_n10971_), .B(u2__abc_52155_new_n4961_), .Y(u2__abc_52155_new_n10972_));
AND2X2 AND2X2_4551 ( .A(u2__abc_52155_new_n10974_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10975_));
AND2X2 AND2X2_4552 ( .A(u2__abc_52155_new_n10975_), .B(u2__abc_52155_new_n10973_), .Y(u2__abc_52155_new_n10976_));
AND2X2 AND2X2_4553 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_168_), .Y(u2__abc_52155_new_n10977_));
AND2X2 AND2X2_4554 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4949_), .Y(u2__abc_52155_new_n10980_));
AND2X2 AND2X2_4555 ( .A(u2__abc_52155_new_n10981_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10982_));
AND2X2 AND2X2_4556 ( .A(u2__abc_52155_new_n10979_), .B(u2__abc_52155_new_n10982_), .Y(u2__abc_52155_new_n10983_));
AND2X2 AND2X2_4557 ( .A(u2__abc_52155_new_n10984_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__170_));
AND2X2 AND2X2_4558 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_171_), .Y(u2__abc_52155_new_n10986_));
AND2X2 AND2X2_4559 ( .A(u2__abc_52155_new_n10973_), .B(u2__abc_52155_new_n4957_), .Y(u2__abc_52155_new_n10987_));
AND2X2 AND2X2_456 ( .A(u1__abc_51895_new_n271_), .B(u1__abc_51895_new_n272_), .Y(u1__abc_51895_new_n273_));
AND2X2 AND2X2_4560 ( .A(u2__abc_52155_new_n10987_), .B(u2__abc_52155_new_n4968_), .Y(u2__abc_52155_new_n10988_));
AND2X2 AND2X2_4561 ( .A(u2__abc_52155_new_n10990_), .B(u2__abc_52155_new_n10989_), .Y(u2__abc_52155_new_n10991_));
AND2X2 AND2X2_4562 ( .A(u2__abc_52155_new_n10992_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n10993_));
AND2X2 AND2X2_4563 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_169_), .Y(u2__abc_52155_new_n10994_));
AND2X2 AND2X2_4564 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4942_), .Y(u2__abc_52155_new_n10997_));
AND2X2 AND2X2_4565 ( .A(u2__abc_52155_new_n10998_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n10999_));
AND2X2 AND2X2_4566 ( .A(u2__abc_52155_new_n10996_), .B(u2__abc_52155_new_n10999_), .Y(u2__abc_52155_new_n11000_));
AND2X2 AND2X2_4567 ( .A(u2__abc_52155_new_n11001_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__171_));
AND2X2 AND2X2_4568 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_172_), .Y(u2__abc_52155_new_n11003_));
AND2X2 AND2X2_4569 ( .A(u2__abc_52155_new_n4957_), .B(u2__abc_52155_new_n4964_), .Y(u2__abc_52155_new_n11004_));
AND2X2 AND2X2_457 ( .A(u1__abc_51895_new_n270_), .B(u1__abc_51895_new_n273_), .Y(u1__abc_51895_new_n274_));
AND2X2 AND2X2_4570 ( .A(u2__abc_52155_new_n10973_), .B(u2__abc_52155_new_n11004_), .Y(u2__abc_52155_new_n11005_));
AND2X2 AND2X2_4571 ( .A(u2__abc_52155_new_n11007_), .B(u2__abc_52155_new_n4952_), .Y(u2__abc_52155_new_n11008_));
AND2X2 AND2X2_4572 ( .A(u2__abc_52155_new_n11010_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11011_));
AND2X2 AND2X2_4573 ( .A(u2__abc_52155_new_n11011_), .B(u2__abc_52155_new_n11009_), .Y(u2__abc_52155_new_n11012_));
AND2X2 AND2X2_4574 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_170_), .Y(u2__abc_52155_new_n11013_));
AND2X2 AND2X2_4575 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4927_), .Y(u2__abc_52155_new_n11016_));
AND2X2 AND2X2_4576 ( .A(u2__abc_52155_new_n11017_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11018_));
AND2X2 AND2X2_4577 ( .A(u2__abc_52155_new_n11015_), .B(u2__abc_52155_new_n11018_), .Y(u2__abc_52155_new_n11019_));
AND2X2 AND2X2_4578 ( .A(u2__abc_52155_new_n11020_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__172_));
AND2X2 AND2X2_4579 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_173_), .Y(u2__abc_52155_new_n11022_));
AND2X2 AND2X2_458 ( .A(u1__abc_51895_new_n267_), .B(u1__abc_51895_new_n274_), .Y(u1__abc_51895_new_n275_));
AND2X2 AND2X2_4580 ( .A(u2__abc_52155_new_n11009_), .B(u2__abc_52155_new_n4948_), .Y(u2__abc_52155_new_n11023_));
AND2X2 AND2X2_4581 ( .A(u2__abc_52155_new_n11023_), .B(u2__abc_52155_new_n4945_), .Y(u2__abc_52155_new_n11024_));
AND2X2 AND2X2_4582 ( .A(u2__abc_52155_new_n11026_), .B(u2__abc_52155_new_n11025_), .Y(u2__abc_52155_new_n11027_));
AND2X2 AND2X2_4583 ( .A(u2__abc_52155_new_n11028_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11029_));
AND2X2 AND2X2_4584 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_171_), .Y(u2__abc_52155_new_n11030_));
AND2X2 AND2X2_4585 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4934_), .Y(u2__abc_52155_new_n11033_));
AND2X2 AND2X2_4586 ( .A(u2__abc_52155_new_n11034_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11035_));
AND2X2 AND2X2_4587 ( .A(u2__abc_52155_new_n11032_), .B(u2__abc_52155_new_n11035_), .Y(u2__abc_52155_new_n11036_));
AND2X2 AND2X2_4588 ( .A(u2__abc_52155_new_n11037_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__173_));
AND2X2 AND2X2_4589 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_174_), .Y(u2__abc_52155_new_n11039_));
AND2X2 AND2X2_459 ( .A(u1__abc_51895_new_n276_), .B(u1__abc_51895_new_n277_), .Y(u1__abc_51895_new_n278_));
AND2X2 AND2X2_4590 ( .A(u2__abc_52155_new_n4941_), .B(u2__abc_52155_new_n4948_), .Y(u2__abc_52155_new_n11040_));
AND2X2 AND2X2_4591 ( .A(u2__abc_52155_new_n11009_), .B(u2__abc_52155_new_n11040_), .Y(u2__abc_52155_new_n11041_));
AND2X2 AND2X2_4592 ( .A(u2__abc_52155_new_n11043_), .B(u2__abc_52155_new_n4930_), .Y(u2__abc_52155_new_n11044_));
AND2X2 AND2X2_4593 ( .A(u2__abc_52155_new_n11046_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11047_));
AND2X2 AND2X2_4594 ( .A(u2__abc_52155_new_n11047_), .B(u2__abc_52155_new_n11045_), .Y(u2__abc_52155_new_n11048_));
AND2X2 AND2X2_4595 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_172_), .Y(u2__abc_52155_new_n11049_));
AND2X2 AND2X2_4596 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4909_), .Y(u2__abc_52155_new_n11052_));
AND2X2 AND2X2_4597 ( .A(u2__abc_52155_new_n11053_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11054_));
AND2X2 AND2X2_4598 ( .A(u2__abc_52155_new_n11051_), .B(u2__abc_52155_new_n11054_), .Y(u2__abc_52155_new_n11055_));
AND2X2 AND2X2_4599 ( .A(u2__abc_52155_new_n11056_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__174_));
AND2X2 AND2X2_46 ( .A(_abc_73687_new_n753_), .B(sqrto_45_), .Y(\o[81] ));
AND2X2 AND2X2_460 ( .A(u1__abc_51895_new_n279_), .B(u1__abc_51895_new_n280_), .Y(u1__abc_51895_new_n281_));
AND2X2 AND2X2_4600 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_175_), .Y(u2__abc_52155_new_n11058_));
AND2X2 AND2X2_4601 ( .A(u2__abc_52155_new_n11045_), .B(u2__abc_52155_new_n4926_), .Y(u2__abc_52155_new_n11059_));
AND2X2 AND2X2_4602 ( .A(u2__abc_52155_new_n11059_), .B(u2__abc_52155_new_n4937_), .Y(u2__abc_52155_new_n11060_));
AND2X2 AND2X2_4603 ( .A(u2__abc_52155_new_n11062_), .B(u2__abc_52155_new_n11061_), .Y(u2__abc_52155_new_n11063_));
AND2X2 AND2X2_4604 ( .A(u2__abc_52155_new_n11064_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11065_));
AND2X2 AND2X2_4605 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_173_), .Y(u2__abc_52155_new_n11066_));
AND2X2 AND2X2_4606 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4916_), .Y(u2__abc_52155_new_n11069_));
AND2X2 AND2X2_4607 ( .A(u2__abc_52155_new_n11070_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11071_));
AND2X2 AND2X2_4608 ( .A(u2__abc_52155_new_n11068_), .B(u2__abc_52155_new_n11071_), .Y(u2__abc_52155_new_n11072_));
AND2X2 AND2X2_4609 ( .A(u2__abc_52155_new_n11073_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__175_));
AND2X2 AND2X2_461 ( .A(u1__abc_51895_new_n278_), .B(u1__abc_51895_new_n281_), .Y(u1__abc_51895_new_n282_));
AND2X2 AND2X2_4610 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_176_), .Y(u2__abc_52155_new_n11075_));
AND2X2 AND2X2_4611 ( .A(u2__abc_52155_new_n10932_), .B(u2__abc_52155_new_n4986_), .Y(u2__abc_52155_new_n11076_));
AND2X2 AND2X2_4612 ( .A(u2__abc_52155_new_n10969_), .B(u2__abc_52155_new_n4969_), .Y(u2__abc_52155_new_n11079_));
AND2X2 AND2X2_4613 ( .A(u2__abc_52155_new_n11080_), .B(u2__abc_52155_new_n11078_), .Y(u2__abc_52155_new_n11081_));
AND2X2 AND2X2_4614 ( .A(u2__abc_52155_new_n11082_), .B(u2__abc_52155_new_n4954_), .Y(u2__abc_52155_new_n11083_));
AND2X2 AND2X2_4615 ( .A(u2__abc_52155_new_n11086_), .B(u2__abc_52155_new_n4938_), .Y(u2__abc_52155_new_n11087_));
AND2X2 AND2X2_4616 ( .A(u2__abc_52155_new_n4926_), .B(u2__abc_52155_new_n4933_), .Y(u2__abc_52155_new_n11089_));
AND2X2 AND2X2_4617 ( .A(u2__abc_52155_new_n11088_), .B(u2__abc_52155_new_n11090_), .Y(u2__abc_52155_new_n11091_));
AND2X2 AND2X2_4618 ( .A(u2__abc_52155_new_n11084_), .B(u2__abc_52155_new_n11091_), .Y(u2__abc_52155_new_n11092_));
AND2X2 AND2X2_4619 ( .A(u2__abc_52155_new_n11077_), .B(u2__abc_52155_new_n11092_), .Y(u2__abc_52155_new_n11093_));
AND2X2 AND2X2_462 ( .A(u1__abc_51895_new_n283_), .B(u1__abc_51895_new_n284_), .Y(u1__abc_51895_new_n285_));
AND2X2 AND2X2_4620 ( .A(u2__abc_52155_new_n10780_), .B(u2__abc_52155_new_n5047_), .Y(u2__abc_52155_new_n11095_));
AND2X2 AND2X2_4621 ( .A(u2__abc_52155_new_n11096_), .B(u2__abc_52155_new_n4912_), .Y(u2__abc_52155_new_n11097_));
AND2X2 AND2X2_4622 ( .A(u2__abc_52155_new_n11099_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11100_));
AND2X2 AND2X2_4623 ( .A(u2__abc_52155_new_n11100_), .B(u2__abc_52155_new_n11098_), .Y(u2__abc_52155_new_n11101_));
AND2X2 AND2X2_4624 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_174_), .Y(u2__abc_52155_new_n11102_));
AND2X2 AND2X2_4625 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4894_), .Y(u2__abc_52155_new_n11105_));
AND2X2 AND2X2_4626 ( .A(u2__abc_52155_new_n11106_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11107_));
AND2X2 AND2X2_4627 ( .A(u2__abc_52155_new_n11104_), .B(u2__abc_52155_new_n11107_), .Y(u2__abc_52155_new_n11108_));
AND2X2 AND2X2_4628 ( .A(u2__abc_52155_new_n11109_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__176_));
AND2X2 AND2X2_4629 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_177_), .Y(u2__abc_52155_new_n11111_));
AND2X2 AND2X2_463 ( .A(u1__abc_51895_new_n286_), .B(u1__abc_51895_new_n287_), .Y(u1__abc_51895_new_n288_));
AND2X2 AND2X2_4630 ( .A(u2__abc_52155_new_n11098_), .B(u2__abc_52155_new_n4908_), .Y(u2__abc_52155_new_n11113_));
AND2X2 AND2X2_4631 ( .A(u2__abc_52155_new_n11116_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11117_));
AND2X2 AND2X2_4632 ( .A(u2__abc_52155_new_n11117_), .B(u2__abc_52155_new_n11114_), .Y(u2__abc_52155_new_n11118_));
AND2X2 AND2X2_4633 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_175_), .Y(u2__abc_52155_new_n11119_));
AND2X2 AND2X2_4634 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4901_), .Y(u2__abc_52155_new_n11122_));
AND2X2 AND2X2_4635 ( .A(u2__abc_52155_new_n11123_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11124_));
AND2X2 AND2X2_4636 ( .A(u2__abc_52155_new_n11121_), .B(u2__abc_52155_new_n11124_), .Y(u2__abc_52155_new_n11125_));
AND2X2 AND2X2_4637 ( .A(u2__abc_52155_new_n11126_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__177_));
AND2X2 AND2X2_4638 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_178_), .Y(u2__abc_52155_new_n11128_));
AND2X2 AND2X2_4639 ( .A(u2__abc_52155_new_n11129_), .B(u2__abc_52155_new_n4915_), .Y(u2__abc_52155_new_n11130_));
AND2X2 AND2X2_464 ( .A(u1__abc_51895_new_n285_), .B(u1__abc_51895_new_n288_), .Y(u1__abc_51895_new_n289_));
AND2X2 AND2X2_4640 ( .A(u2__abc_52155_new_n11096_), .B(u2__abc_52155_new_n4920_), .Y(u2__abc_52155_new_n11132_));
AND2X2 AND2X2_4641 ( .A(u2__abc_52155_new_n11133_), .B(u2__abc_52155_new_n4897_), .Y(u2__abc_52155_new_n11134_));
AND2X2 AND2X2_4642 ( .A(u2__abc_52155_new_n11136_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11137_));
AND2X2 AND2X2_4643 ( .A(u2__abc_52155_new_n11137_), .B(u2__abc_52155_new_n11135_), .Y(u2__abc_52155_new_n11138_));
AND2X2 AND2X2_4644 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_176_), .Y(u2__abc_52155_new_n11139_));
AND2X2 AND2X2_4645 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4885_), .Y(u2__abc_52155_new_n11142_));
AND2X2 AND2X2_4646 ( .A(u2__abc_52155_new_n11143_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11144_));
AND2X2 AND2X2_4647 ( .A(u2__abc_52155_new_n11141_), .B(u2__abc_52155_new_n11144_), .Y(u2__abc_52155_new_n11145_));
AND2X2 AND2X2_4648 ( .A(u2__abc_52155_new_n11146_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__178_));
AND2X2 AND2X2_4649 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_179_), .Y(u2__abc_52155_new_n11148_));
AND2X2 AND2X2_465 ( .A(u1__abc_51895_new_n282_), .B(u1__abc_51895_new_n289_), .Y(u1__abc_51895_new_n290_));
AND2X2 AND2X2_4650 ( .A(u2__abc_52155_new_n11135_), .B(u2__abc_52155_new_n4893_), .Y(u2__abc_52155_new_n11149_));
AND2X2 AND2X2_4651 ( .A(u2__abc_52155_new_n11149_), .B(u2__abc_52155_new_n4904_), .Y(u2__abc_52155_new_n11150_));
AND2X2 AND2X2_4652 ( .A(u2__abc_52155_new_n11152_), .B(u2__abc_52155_new_n11151_), .Y(u2__abc_52155_new_n11153_));
AND2X2 AND2X2_4653 ( .A(u2__abc_52155_new_n11154_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11155_));
AND2X2 AND2X2_4654 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_177_), .Y(u2__abc_52155_new_n11156_));
AND2X2 AND2X2_4655 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4878_), .Y(u2__abc_52155_new_n11159_));
AND2X2 AND2X2_4656 ( .A(u2__abc_52155_new_n11160_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11161_));
AND2X2 AND2X2_4657 ( .A(u2__abc_52155_new_n11158_), .B(u2__abc_52155_new_n11161_), .Y(u2__abc_52155_new_n11162_));
AND2X2 AND2X2_4658 ( .A(u2__abc_52155_new_n11163_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__179_));
AND2X2 AND2X2_4659 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_180_), .Y(u2__abc_52155_new_n11165_));
AND2X2 AND2X2_466 ( .A(u1__abc_51895_new_n275_), .B(u1__abc_51895_new_n290_), .Y(u1__abc_51895_new_n291_));
AND2X2 AND2X2_4660 ( .A(u2__abc_52155_new_n4893_), .B(u2__abc_52155_new_n4900_), .Y(u2__abc_52155_new_n11166_));
AND2X2 AND2X2_4661 ( .A(u2__abc_52155_new_n11135_), .B(u2__abc_52155_new_n11166_), .Y(u2__abc_52155_new_n11167_));
AND2X2 AND2X2_4662 ( .A(u2__abc_52155_new_n11169_), .B(u2__abc_52155_new_n4888_), .Y(u2__abc_52155_new_n11170_));
AND2X2 AND2X2_4663 ( .A(u2__abc_52155_new_n11172_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11173_));
AND2X2 AND2X2_4664 ( .A(u2__abc_52155_new_n11173_), .B(u2__abc_52155_new_n11171_), .Y(u2__abc_52155_new_n11174_));
AND2X2 AND2X2_4665 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_178_), .Y(u2__abc_52155_new_n11175_));
AND2X2 AND2X2_4666 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4863_), .Y(u2__abc_52155_new_n11178_));
AND2X2 AND2X2_4667 ( .A(u2__abc_52155_new_n11179_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11180_));
AND2X2 AND2X2_4668 ( .A(u2__abc_52155_new_n11177_), .B(u2__abc_52155_new_n11180_), .Y(u2__abc_52155_new_n11181_));
AND2X2 AND2X2_4669 ( .A(u2__abc_52155_new_n11182_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__180_));
AND2X2 AND2X2_467 ( .A(u1__abc_51895_new_n292_), .B(u1__abc_51895_new_n293_), .Y(u1__abc_51895_new_n294_));
AND2X2 AND2X2_4670 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_181_), .Y(u2__abc_52155_new_n11184_));
AND2X2 AND2X2_4671 ( .A(u2__abc_52155_new_n11171_), .B(u2__abc_52155_new_n4884_), .Y(u2__abc_52155_new_n11185_));
AND2X2 AND2X2_4672 ( .A(u2__abc_52155_new_n11185_), .B(u2__abc_52155_new_n4881_), .Y(u2__abc_52155_new_n11186_));
AND2X2 AND2X2_4673 ( .A(u2__abc_52155_new_n11188_), .B(u2__abc_52155_new_n11187_), .Y(u2__abc_52155_new_n11189_));
AND2X2 AND2X2_4674 ( .A(u2__abc_52155_new_n11190_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11191_));
AND2X2 AND2X2_4675 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_179_), .Y(u2__abc_52155_new_n11192_));
AND2X2 AND2X2_4676 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4870_), .Y(u2__abc_52155_new_n11195_));
AND2X2 AND2X2_4677 ( .A(u2__abc_52155_new_n11196_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11197_));
AND2X2 AND2X2_4678 ( .A(u2__abc_52155_new_n11194_), .B(u2__abc_52155_new_n11197_), .Y(u2__abc_52155_new_n11198_));
AND2X2 AND2X2_4679 ( .A(u2__abc_52155_new_n11199_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__181_));
AND2X2 AND2X2_468 ( .A(u1__abc_51895_new_n295_), .B(u1__abc_51895_new_n296_), .Y(u1__abc_51895_new_n297_));
AND2X2 AND2X2_4680 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_182_), .Y(u2__abc_52155_new_n11201_));
AND2X2 AND2X2_4681 ( .A(u2__abc_52155_new_n4877_), .B(u2__abc_52155_new_n4884_), .Y(u2__abc_52155_new_n11202_));
AND2X2 AND2X2_4682 ( .A(u2__abc_52155_new_n11171_), .B(u2__abc_52155_new_n11202_), .Y(u2__abc_52155_new_n11203_));
AND2X2 AND2X2_4683 ( .A(u2__abc_52155_new_n11205_), .B(u2__abc_52155_new_n4866_), .Y(u2__abc_52155_new_n11206_));
AND2X2 AND2X2_4684 ( .A(u2__abc_52155_new_n11208_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11209_));
AND2X2 AND2X2_4685 ( .A(u2__abc_52155_new_n11209_), .B(u2__abc_52155_new_n11207_), .Y(u2__abc_52155_new_n11210_));
AND2X2 AND2X2_4686 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_180_), .Y(u2__abc_52155_new_n11211_));
AND2X2 AND2X2_4687 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4800_), .Y(u2__abc_52155_new_n11214_));
AND2X2 AND2X2_4688 ( .A(u2__abc_52155_new_n11215_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11216_));
AND2X2 AND2X2_4689 ( .A(u2__abc_52155_new_n11213_), .B(u2__abc_52155_new_n11216_), .Y(u2__abc_52155_new_n11217_));
AND2X2 AND2X2_469 ( .A(u1__abc_51895_new_n294_), .B(u1__abc_51895_new_n297_), .Y(u1__abc_51895_new_n298_));
AND2X2 AND2X2_4690 ( .A(u2__abc_52155_new_n11218_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__182_));
AND2X2 AND2X2_4691 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_183_), .Y(u2__abc_52155_new_n11220_));
AND2X2 AND2X2_4692 ( .A(u2__abc_52155_new_n11207_), .B(u2__abc_52155_new_n4862_), .Y(u2__abc_52155_new_n11221_));
AND2X2 AND2X2_4693 ( .A(u2__abc_52155_new_n11221_), .B(u2__abc_52155_new_n4873_), .Y(u2__abc_52155_new_n11222_));
AND2X2 AND2X2_4694 ( .A(u2__abc_52155_new_n11224_), .B(u2__abc_52155_new_n11223_), .Y(u2__abc_52155_new_n11225_));
AND2X2 AND2X2_4695 ( .A(u2__abc_52155_new_n11226_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11227_));
AND2X2 AND2X2_4696 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_181_), .Y(u2__abc_52155_new_n11228_));
AND2X2 AND2X2_4697 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4807_), .Y(u2__abc_52155_new_n11231_));
AND2X2 AND2X2_4698 ( .A(u2__abc_52155_new_n11232_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11233_));
AND2X2 AND2X2_4699 ( .A(u2__abc_52155_new_n11230_), .B(u2__abc_52155_new_n11233_), .Y(u2__abc_52155_new_n11234_));
AND2X2 AND2X2_47 ( .A(_abc_73687_new_n753_), .B(sqrto_46_), .Y(\o[82] ));
AND2X2 AND2X2_470 ( .A(u1__abc_51895_new_n299_), .B(u1__abc_51895_new_n300_), .Y(u1__abc_51895_new_n301_));
AND2X2 AND2X2_4700 ( .A(u2__abc_52155_new_n11235_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__183_));
AND2X2 AND2X2_4701 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_184_), .Y(u2__abc_52155_new_n11237_));
AND2X2 AND2X2_4702 ( .A(u2__abc_52155_new_n11131_), .B(u2__abc_52155_new_n4905_), .Y(u2__abc_52155_new_n11239_));
AND2X2 AND2X2_4703 ( .A(u2__abc_52155_new_n11240_), .B(u2__abc_52155_new_n11238_), .Y(u2__abc_52155_new_n11241_));
AND2X2 AND2X2_4704 ( .A(u2__abc_52155_new_n11242_), .B(u2__abc_52155_new_n4890_), .Y(u2__abc_52155_new_n11243_));
AND2X2 AND2X2_4705 ( .A(u2__abc_52155_new_n11245_), .B(u2__abc_52155_new_n4874_), .Y(u2__abc_52155_new_n11246_));
AND2X2 AND2X2_4706 ( .A(u2__abc_52155_new_n4872_), .B(u2__abc_52155_new_n4861_), .Y(u2__abc_52155_new_n11247_));
AND2X2 AND2X2_4707 ( .A(u2__abc_52155_new_n11096_), .B(u2__abc_52155_new_n4922_), .Y(u2__abc_52155_new_n11251_));
AND2X2 AND2X2_4708 ( .A(u2__abc_52155_new_n11252_), .B(u2__abc_52155_new_n4803_), .Y(u2__abc_52155_new_n11253_));
AND2X2 AND2X2_4709 ( .A(u2__abc_52155_new_n11255_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11256_));
AND2X2 AND2X2_471 ( .A(u1__abc_51895_new_n302_), .B(u1__abc_51895_new_n303_), .Y(u1__abc_51895_new_n304_));
AND2X2 AND2X2_4710 ( .A(u2__abc_52155_new_n11256_), .B(u2__abc_52155_new_n11254_), .Y(u2__abc_52155_new_n11257_));
AND2X2 AND2X2_4711 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_182_), .Y(u2__abc_52155_new_n11258_));
AND2X2 AND2X2_4712 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4815_), .Y(u2__abc_52155_new_n11261_));
AND2X2 AND2X2_4713 ( .A(u2__abc_52155_new_n11262_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11263_));
AND2X2 AND2X2_4714 ( .A(u2__abc_52155_new_n11260_), .B(u2__abc_52155_new_n11263_), .Y(u2__abc_52155_new_n11264_));
AND2X2 AND2X2_4715 ( .A(u2__abc_52155_new_n11265_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__184_));
AND2X2 AND2X2_4716 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_185_), .Y(u2__abc_52155_new_n11267_));
AND2X2 AND2X2_4717 ( .A(u2__abc_52155_new_n11254_), .B(u2__abc_52155_new_n4799_), .Y(u2__abc_52155_new_n11268_));
AND2X2 AND2X2_4718 ( .A(u2__abc_52155_new_n11268_), .B(u2__abc_52155_new_n4810_), .Y(u2__abc_52155_new_n11269_));
AND2X2 AND2X2_4719 ( .A(u2__abc_52155_new_n11271_), .B(u2__abc_52155_new_n11270_), .Y(u2__abc_52155_new_n11272_));
AND2X2 AND2X2_472 ( .A(u1__abc_51895_new_n301_), .B(u1__abc_51895_new_n304_), .Y(u1__abc_51895_new_n305_));
AND2X2 AND2X2_4720 ( .A(u2__abc_52155_new_n11273_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11274_));
AND2X2 AND2X2_4721 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_183_), .Y(u2__abc_52155_new_n11275_));
AND2X2 AND2X2_4722 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4822_), .Y(u2__abc_52155_new_n11278_));
AND2X2 AND2X2_4723 ( .A(u2__abc_52155_new_n11279_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11280_));
AND2X2 AND2X2_4724 ( .A(u2__abc_52155_new_n11277_), .B(u2__abc_52155_new_n11280_), .Y(u2__abc_52155_new_n11281_));
AND2X2 AND2X2_4725 ( .A(u2__abc_52155_new_n11282_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__185_));
AND2X2 AND2X2_4726 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_186_), .Y(u2__abc_52155_new_n11284_));
AND2X2 AND2X2_4727 ( .A(u2__abc_52155_new_n11285_), .B(u2__abc_52155_new_n4806_), .Y(u2__abc_52155_new_n11286_));
AND2X2 AND2X2_4728 ( .A(u2__abc_52155_new_n11252_), .B(u2__abc_52155_new_n4811_), .Y(u2__abc_52155_new_n11288_));
AND2X2 AND2X2_4729 ( .A(u2__abc_52155_new_n11289_), .B(u2__abc_52155_new_n4818_), .Y(u2__abc_52155_new_n11290_));
AND2X2 AND2X2_473 ( .A(u1__abc_51895_new_n298_), .B(u1__abc_51895_new_n305_), .Y(u1__abc_51895_new_n306_));
AND2X2 AND2X2_4730 ( .A(u2__abc_52155_new_n11292_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11293_));
AND2X2 AND2X2_4731 ( .A(u2__abc_52155_new_n11293_), .B(u2__abc_52155_new_n11291_), .Y(u2__abc_52155_new_n11294_));
AND2X2 AND2X2_4732 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_184_), .Y(u2__abc_52155_new_n11295_));
AND2X2 AND2X2_4733 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4853_), .Y(u2__abc_52155_new_n11298_));
AND2X2 AND2X2_4734 ( .A(u2__abc_52155_new_n11299_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11300_));
AND2X2 AND2X2_4735 ( .A(u2__abc_52155_new_n11297_), .B(u2__abc_52155_new_n11300_), .Y(u2__abc_52155_new_n11301_));
AND2X2 AND2X2_4736 ( .A(u2__abc_52155_new_n11302_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__186_));
AND2X2 AND2X2_4737 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_187_), .Y(u2__abc_52155_new_n11304_));
AND2X2 AND2X2_4738 ( .A(u2__abc_52155_new_n11291_), .B(u2__abc_52155_new_n4814_), .Y(u2__abc_52155_new_n11305_));
AND2X2 AND2X2_4739 ( .A(u2__abc_52155_new_n11305_), .B(u2__abc_52155_new_n4825_), .Y(u2__abc_52155_new_n11306_));
AND2X2 AND2X2_474 ( .A(u1__abc_51895_new_n307_), .B(u1__abc_51895_new_n308_), .Y(u1__abc_51895_new_n309_));
AND2X2 AND2X2_4740 ( .A(u2__abc_52155_new_n11308_), .B(u2__abc_52155_new_n11307_), .Y(u2__abc_52155_new_n11309_));
AND2X2 AND2X2_4741 ( .A(u2__abc_52155_new_n11310_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11311_));
AND2X2 AND2X2_4742 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_185_), .Y(u2__abc_52155_new_n11312_));
AND2X2 AND2X2_4743 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4846_), .Y(u2__abc_52155_new_n11315_));
AND2X2 AND2X2_4744 ( .A(u2__abc_52155_new_n11316_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11317_));
AND2X2 AND2X2_4745 ( .A(u2__abc_52155_new_n11314_), .B(u2__abc_52155_new_n11317_), .Y(u2__abc_52155_new_n11318_));
AND2X2 AND2X2_4746 ( .A(u2__abc_52155_new_n11319_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__187_));
AND2X2 AND2X2_4747 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_188_), .Y(u2__abc_52155_new_n11321_));
AND2X2 AND2X2_4748 ( .A(u2__abc_52155_new_n11287_), .B(u2__abc_52155_new_n4826_), .Y(u2__abc_52155_new_n11322_));
AND2X2 AND2X2_4749 ( .A(u2__abc_52155_new_n4824_), .B(u2__abc_52155_new_n4813_), .Y(u2__abc_52155_new_n11323_));
AND2X2 AND2X2_475 ( .A(u1__abc_51895_new_n310_), .B(u1__abc_51895_new_n311_), .Y(u1__abc_51895_new_n312_));
AND2X2 AND2X2_4750 ( .A(u2__abc_52155_new_n11252_), .B(u2__abc_52155_new_n4827_), .Y(u2__abc_52155_new_n11326_));
AND2X2 AND2X2_4751 ( .A(u2__abc_52155_new_n11327_), .B(u2__abc_52155_new_n4856_), .Y(u2__abc_52155_new_n11328_));
AND2X2 AND2X2_4752 ( .A(u2__abc_52155_new_n11330_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11331_));
AND2X2 AND2X2_4753 ( .A(u2__abc_52155_new_n11331_), .B(u2__abc_52155_new_n11329_), .Y(u2__abc_52155_new_n11332_));
AND2X2 AND2X2_4754 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_186_), .Y(u2__abc_52155_new_n11333_));
AND2X2 AND2X2_4755 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4831_), .Y(u2__abc_52155_new_n11336_));
AND2X2 AND2X2_4756 ( .A(u2__abc_52155_new_n11337_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11338_));
AND2X2 AND2X2_4757 ( .A(u2__abc_52155_new_n11335_), .B(u2__abc_52155_new_n11338_), .Y(u2__abc_52155_new_n11339_));
AND2X2 AND2X2_4758 ( .A(u2__abc_52155_new_n11340_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__188_));
AND2X2 AND2X2_4759 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_189_), .Y(u2__abc_52155_new_n11342_));
AND2X2 AND2X2_476 ( .A(u1__abc_51895_new_n309_), .B(u1__abc_51895_new_n312_), .Y(u1__abc_51895_new_n313_));
AND2X2 AND2X2_4760 ( .A(u2__abc_52155_new_n11329_), .B(u2__abc_52155_new_n4852_), .Y(u2__abc_52155_new_n11343_));
AND2X2 AND2X2_4761 ( .A(u2__abc_52155_new_n11343_), .B(u2__abc_52155_new_n4849_), .Y(u2__abc_52155_new_n11344_));
AND2X2 AND2X2_4762 ( .A(u2__abc_52155_new_n11346_), .B(u2__abc_52155_new_n11345_), .Y(u2__abc_52155_new_n11347_));
AND2X2 AND2X2_4763 ( .A(u2__abc_52155_new_n11348_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11349_));
AND2X2 AND2X2_4764 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_187_), .Y(u2__abc_52155_new_n11350_));
AND2X2 AND2X2_4765 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4838_), .Y(u2__abc_52155_new_n11353_));
AND2X2 AND2X2_4766 ( .A(u2__abc_52155_new_n11354_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11355_));
AND2X2 AND2X2_4767 ( .A(u2__abc_52155_new_n11352_), .B(u2__abc_52155_new_n11355_), .Y(u2__abc_52155_new_n11356_));
AND2X2 AND2X2_4768 ( .A(u2__abc_52155_new_n11357_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__189_));
AND2X2 AND2X2_4769 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_190_), .Y(u2__abc_52155_new_n11359_));
AND2X2 AND2X2_477 ( .A(u1__abc_51895_new_n314_), .B(u1__abc_51895_new_n315_), .Y(u1__abc_51895_new_n316_));
AND2X2 AND2X2_4770 ( .A(u2__abc_52155_new_n4845_), .B(u2__abc_52155_new_n4852_), .Y(u2__abc_52155_new_n11360_));
AND2X2 AND2X2_4771 ( .A(u2__abc_52155_new_n11329_), .B(u2__abc_52155_new_n11360_), .Y(u2__abc_52155_new_n11361_));
AND2X2 AND2X2_4772 ( .A(u2__abc_52155_new_n11363_), .B(u2__abc_52155_new_n4834_), .Y(u2__abc_52155_new_n11364_));
AND2X2 AND2X2_4773 ( .A(u2__abc_52155_new_n11366_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11367_));
AND2X2 AND2X2_4774 ( .A(u2__abc_52155_new_n11367_), .B(u2__abc_52155_new_n11365_), .Y(u2__abc_52155_new_n11368_));
AND2X2 AND2X2_4775 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_188_), .Y(u2__abc_52155_new_n11369_));
AND2X2 AND2X2_4776 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4780_), .Y(u2__abc_52155_new_n11372_));
AND2X2 AND2X2_4777 ( .A(u2__abc_52155_new_n11373_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11374_));
AND2X2 AND2X2_4778 ( .A(u2__abc_52155_new_n11371_), .B(u2__abc_52155_new_n11374_), .Y(u2__abc_52155_new_n11375_));
AND2X2 AND2X2_4779 ( .A(u2__abc_52155_new_n11376_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__190_));
AND2X2 AND2X2_478 ( .A(u1__abc_51895_new_n317_), .B(u1__abc_51895_new_n318_), .Y(u1__abc_51895_new_n319_));
AND2X2 AND2X2_4780 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_191_), .Y(u2__abc_52155_new_n11378_));
AND2X2 AND2X2_4781 ( .A(u2__abc_52155_new_n11365_), .B(u2__abc_52155_new_n4830_), .Y(u2__abc_52155_new_n11379_));
AND2X2 AND2X2_4782 ( .A(u2__abc_52155_new_n11379_), .B(u2__abc_52155_new_n4841_), .Y(u2__abc_52155_new_n11380_));
AND2X2 AND2X2_4783 ( .A(u2__abc_52155_new_n11382_), .B(u2__abc_52155_new_n11381_), .Y(u2__abc_52155_new_n11383_));
AND2X2 AND2X2_4784 ( .A(u2__abc_52155_new_n11384_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11385_));
AND2X2 AND2X2_4785 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_189_), .Y(u2__abc_52155_new_n11386_));
AND2X2 AND2X2_4786 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4787_), .Y(u2__abc_52155_new_n11389_));
AND2X2 AND2X2_4787 ( .A(u2__abc_52155_new_n11390_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11391_));
AND2X2 AND2X2_4788 ( .A(u2__abc_52155_new_n11388_), .B(u2__abc_52155_new_n11391_), .Y(u2__abc_52155_new_n11392_));
AND2X2 AND2X2_4789 ( .A(u2__abc_52155_new_n11393_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__191_));
AND2X2 AND2X2_479 ( .A(u1__abc_51895_new_n316_), .B(u1__abc_51895_new_n319_), .Y(u1__abc_51895_new_n320_));
AND2X2 AND2X2_4790 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_192_), .Y(u2__abc_52155_new_n11395_));
AND2X2 AND2X2_4791 ( .A(u2__abc_52155_new_n10778_), .B(u2__abc_52155_new_n5048_), .Y(u2__abc_52155_new_n11396_));
AND2X2 AND2X2_4792 ( .A(u2__abc_52155_new_n11094_), .B(u2__abc_52155_new_n4923_), .Y(u2__abc_52155_new_n11397_));
AND2X2 AND2X2_4793 ( .A(u2__abc_52155_new_n11250_), .B(u2__abc_52155_new_n4859_), .Y(u2__abc_52155_new_n11398_));
AND2X2 AND2X2_4794 ( .A(u2__abc_52155_new_n11325_), .B(u2__abc_52155_new_n4858_), .Y(u2__abc_52155_new_n11399_));
AND2X2 AND2X2_4795 ( .A(u2__abc_52155_new_n11401_), .B(u2__abc_52155_new_n4842_), .Y(u2__abc_52155_new_n11402_));
AND2X2 AND2X2_4796 ( .A(u2__abc_52155_new_n4840_), .B(u2__abc_52155_new_n4829_), .Y(u2__abc_52155_new_n11403_));
AND2X2 AND2X2_4797 ( .A(u2__abc_52155_new_n10150_), .B(u2__abc_52155_new_n5286_), .Y(u2__abc_52155_new_n11410_));
AND2X2 AND2X2_4798 ( .A(u2__abc_52155_new_n11411_), .B(u2__abc_52155_new_n4783_), .Y(u2__abc_52155_new_n11412_));
AND2X2 AND2X2_4799 ( .A(u2__abc_52155_new_n11413_), .B(u2__abc_52155_new_n11414_), .Y(u2__abc_52155_new_n11415_));
AND2X2 AND2X2_48 ( .A(_abc_73687_new_n753_), .B(sqrto_47_), .Y(\o[83] ));
AND2X2 AND2X2_480 ( .A(u1__abc_51895_new_n313_), .B(u1__abc_51895_new_n320_), .Y(u1__abc_51895_new_n321_));
AND2X2 AND2X2_4800 ( .A(u2__abc_52155_new_n11415_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11416_));
AND2X2 AND2X2_4801 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_190_), .Y(u2__abc_52155_new_n11417_));
AND2X2 AND2X2_4802 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4767_), .Y(u2__abc_52155_new_n11420_));
AND2X2 AND2X2_4803 ( .A(u2__abc_52155_new_n11421_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11422_));
AND2X2 AND2X2_4804 ( .A(u2__abc_52155_new_n11419_), .B(u2__abc_52155_new_n11422_), .Y(u2__abc_52155_new_n11423_));
AND2X2 AND2X2_4805 ( .A(u2__abc_52155_new_n11424_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__192_));
AND2X2 AND2X2_4806 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_193_), .Y(u2__abc_52155_new_n11426_));
AND2X2 AND2X2_4807 ( .A(u2__abc_52155_new_n11413_), .B(u2__abc_52155_new_n4779_), .Y(u2__abc_52155_new_n11428_));
AND2X2 AND2X2_4808 ( .A(u2__abc_52155_new_n11429_), .B(u2__abc_52155_new_n11427_), .Y(u2__abc_52155_new_n11430_));
AND2X2 AND2X2_4809 ( .A(u2__abc_52155_new_n11428_), .B(u2__abc_52155_new_n4790_), .Y(u2__abc_52155_new_n11431_));
AND2X2 AND2X2_481 ( .A(u1__abc_51895_new_n306_), .B(u1__abc_51895_new_n321_), .Y(u1__abc_51895_new_n322_));
AND2X2 AND2X2_4810 ( .A(u2__abc_52155_new_n11432_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11433_));
AND2X2 AND2X2_4811 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_191_), .Y(u2__abc_52155_new_n11434_));
AND2X2 AND2X2_4812 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4772_), .Y(u2__abc_52155_new_n11437_));
AND2X2 AND2X2_4813 ( .A(u2__abc_52155_new_n11438_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11439_));
AND2X2 AND2X2_4814 ( .A(u2__abc_52155_new_n11436_), .B(u2__abc_52155_new_n11439_), .Y(u2__abc_52155_new_n11440_));
AND2X2 AND2X2_4815 ( .A(u2__abc_52155_new_n11441_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__193_));
AND2X2 AND2X2_4816 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_194_), .Y(u2__abc_52155_new_n11443_));
AND2X2 AND2X2_4817 ( .A(u2__abc_52155_new_n11429_), .B(u2__abc_52155_new_n4789_), .Y(u2__abc_52155_new_n11445_));
AND2X2 AND2X2_4818 ( .A(u2__abc_52155_new_n11446_), .B(u2__abc_52155_new_n11444_), .Y(u2__abc_52155_new_n11447_));
AND2X2 AND2X2_4819 ( .A(u2__abc_52155_new_n11449_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11450_));
AND2X2 AND2X2_482 ( .A(u1__abc_51895_new_n291_), .B(u1__abc_51895_new_n322_), .Y(u1__abc_51895_new_n323_));
AND2X2 AND2X2_4820 ( .A(u2__abc_52155_new_n11450_), .B(u2__abc_52155_new_n11448_), .Y(u2__abc_52155_new_n11451_));
AND2X2 AND2X2_4821 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_192_), .Y(u2__abc_52155_new_n11452_));
AND2X2 AND2X2_4822 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4759_), .Y(u2__abc_52155_new_n11455_));
AND2X2 AND2X2_4823 ( .A(u2__abc_52155_new_n11456_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11457_));
AND2X2 AND2X2_4824 ( .A(u2__abc_52155_new_n11454_), .B(u2__abc_52155_new_n11457_), .Y(u2__abc_52155_new_n11458_));
AND2X2 AND2X2_4825 ( .A(u2__abc_52155_new_n11459_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__194_));
AND2X2 AND2X2_4826 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_195_), .Y(u2__abc_52155_new_n11461_));
AND2X2 AND2X2_4827 ( .A(u2__abc_52155_new_n11448_), .B(u2__abc_52155_new_n11462_), .Y(u2__abc_52155_new_n11463_));
AND2X2 AND2X2_4828 ( .A(u2__abc_52155_new_n11467_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11468_));
AND2X2 AND2X2_4829 ( .A(u2__abc_52155_new_n11468_), .B(u2__abc_52155_new_n11464_), .Y(u2__abc_52155_new_n11469_));
AND2X2 AND2X2_483 ( .A(u1__abc_51895_new_n324_), .B(u1__abc_51895_new_n325_), .Y(u1__abc_51895_new_n326_));
AND2X2 AND2X2_4830 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_193_), .Y(u2__abc_52155_new_n11470_));
AND2X2 AND2X2_4831 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4752_), .Y(u2__abc_52155_new_n11473_));
AND2X2 AND2X2_4832 ( .A(u2__abc_52155_new_n11474_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11475_));
AND2X2 AND2X2_4833 ( .A(u2__abc_52155_new_n11472_), .B(u2__abc_52155_new_n11475_), .Y(u2__abc_52155_new_n11476_));
AND2X2 AND2X2_4834 ( .A(u2__abc_52155_new_n11477_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__195_));
AND2X2 AND2X2_4835 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_196_), .Y(u2__abc_52155_new_n11479_));
AND2X2 AND2X2_4836 ( .A(u2__abc_52155_new_n4779_), .B(u2__abc_52155_new_n4786_), .Y(u2__abc_52155_new_n11480_));
AND2X2 AND2X2_4837 ( .A(u2__abc_52155_new_n11483_), .B(u2__abc_52155_new_n5452_), .Y(u2__abc_52155_new_n11484_));
AND2X2 AND2X2_4838 ( .A(u2__abc_52155_new_n11482_), .B(u2__abc_52155_new_n11484_), .Y(u2__abc_52155_new_n11485_));
AND2X2 AND2X2_4839 ( .A(u2__abc_52155_new_n11411_), .B(u2__abc_52155_new_n4792_), .Y(u2__abc_52155_new_n11487_));
AND2X2 AND2X2_484 ( .A(u1__abc_51895_new_n327_), .B(u1__abc_51895_new_n328_), .Y(u1__abc_51895_new_n329_));
AND2X2 AND2X2_4840 ( .A(u2__abc_52155_new_n11488_), .B(u2__abc_52155_new_n4762_), .Y(u2__abc_52155_new_n11489_));
AND2X2 AND2X2_4841 ( .A(u2__abc_52155_new_n11491_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11492_));
AND2X2 AND2X2_4842 ( .A(u2__abc_52155_new_n11492_), .B(u2__abc_52155_new_n11490_), .Y(u2__abc_52155_new_n11493_));
AND2X2 AND2X2_4843 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_194_), .Y(u2__abc_52155_new_n11494_));
AND2X2 AND2X2_4844 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4737_), .Y(u2__abc_52155_new_n11497_));
AND2X2 AND2X2_4845 ( .A(u2__abc_52155_new_n11498_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11499_));
AND2X2 AND2X2_4846 ( .A(u2__abc_52155_new_n11496_), .B(u2__abc_52155_new_n11499_), .Y(u2__abc_52155_new_n11500_));
AND2X2 AND2X2_4847 ( .A(u2__abc_52155_new_n11501_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__196_));
AND2X2 AND2X2_4848 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_197_), .Y(u2__abc_52155_new_n11503_));
AND2X2 AND2X2_4849 ( .A(u2__abc_52155_new_n11490_), .B(u2__abc_52155_new_n4758_), .Y(u2__abc_52155_new_n11504_));
AND2X2 AND2X2_485 ( .A(u1__abc_51895_new_n326_), .B(u1__abc_51895_new_n329_), .Y(u1__abc_51895_new_n330_));
AND2X2 AND2X2_4850 ( .A(u2__abc_52155_new_n11505_), .B(u2__abc_52155_new_n4755_), .Y(u2__abc_52155_new_n11506_));
AND2X2 AND2X2_4851 ( .A(u2__abc_52155_new_n11508_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11509_));
AND2X2 AND2X2_4852 ( .A(u2__abc_52155_new_n11509_), .B(u2__abc_52155_new_n11507_), .Y(u2__abc_52155_new_n11510_));
AND2X2 AND2X2_4853 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_195_), .Y(u2__abc_52155_new_n11511_));
AND2X2 AND2X2_4854 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4744_), .Y(u2__abc_52155_new_n11514_));
AND2X2 AND2X2_4855 ( .A(u2__abc_52155_new_n11515_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11516_));
AND2X2 AND2X2_4856 ( .A(u2__abc_52155_new_n11513_), .B(u2__abc_52155_new_n11516_), .Y(u2__abc_52155_new_n11517_));
AND2X2 AND2X2_4857 ( .A(u2__abc_52155_new_n11518_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__197_));
AND2X2 AND2X2_4858 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_198_), .Y(u2__abc_52155_new_n11520_));
AND2X2 AND2X2_4859 ( .A(u2__abc_52155_new_n11507_), .B(u2__abc_52155_new_n4751_), .Y(u2__abc_52155_new_n11521_));
AND2X2 AND2X2_486 ( .A(u1__abc_51895_new_n331_), .B(u1__abc_51895_new_n332_), .Y(u1__abc_51895_new_n333_));
AND2X2 AND2X2_4860 ( .A(u2__abc_52155_new_n11522_), .B(u2__abc_52155_new_n4740_), .Y(u2__abc_52155_new_n11523_));
AND2X2 AND2X2_4861 ( .A(u2__abc_52155_new_n11525_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11526_));
AND2X2 AND2X2_4862 ( .A(u2__abc_52155_new_n11526_), .B(u2__abc_52155_new_n11524_), .Y(u2__abc_52155_new_n11527_));
AND2X2 AND2X2_4863 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_196_), .Y(u2__abc_52155_new_n11528_));
AND2X2 AND2X2_4864 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4696_), .Y(u2__abc_52155_new_n11531_));
AND2X2 AND2X2_4865 ( .A(u2__abc_52155_new_n11532_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11533_));
AND2X2 AND2X2_4866 ( .A(u2__abc_52155_new_n11530_), .B(u2__abc_52155_new_n11533_), .Y(u2__abc_52155_new_n11534_));
AND2X2 AND2X2_4867 ( .A(u2__abc_52155_new_n11535_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__198_));
AND2X2 AND2X2_4868 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_199_), .Y(u2__abc_52155_new_n11537_));
AND2X2 AND2X2_4869 ( .A(u2__abc_52155_new_n11524_), .B(u2__abc_52155_new_n4736_), .Y(u2__abc_52155_new_n11538_));
AND2X2 AND2X2_487 ( .A(u1__abc_51895_new_n334_), .B(u1__abc_51895_new_n335_), .Y(u1__abc_51895_new_n336_));
AND2X2 AND2X2_4870 ( .A(u2__abc_52155_new_n11538_), .B(u2__abc_52155_new_n4747_), .Y(u2__abc_52155_new_n11539_));
AND2X2 AND2X2_4871 ( .A(u2__abc_52155_new_n11541_), .B(u2__abc_52155_new_n11540_), .Y(u2__abc_52155_new_n11542_));
AND2X2 AND2X2_4872 ( .A(u2__abc_52155_new_n11543_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11544_));
AND2X2 AND2X2_4873 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_197_), .Y(u2__abc_52155_new_n11545_));
AND2X2 AND2X2_4874 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4689_), .Y(u2__abc_52155_new_n11548_));
AND2X2 AND2X2_4875 ( .A(u2__abc_52155_new_n11549_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11550_));
AND2X2 AND2X2_4876 ( .A(u2__abc_52155_new_n11547_), .B(u2__abc_52155_new_n11550_), .Y(u2__abc_52155_new_n11551_));
AND2X2 AND2X2_4877 ( .A(u2__abc_52155_new_n11552_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__199_));
AND2X2 AND2X2_4878 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_200_), .Y(u2__abc_52155_new_n11554_));
AND2X2 AND2X2_4879 ( .A(u2__abc_52155_new_n11486_), .B(u2__abc_52155_new_n4764_), .Y(u2__abc_52155_new_n11555_));
AND2X2 AND2X2_488 ( .A(u1__abc_51895_new_n333_), .B(u1__abc_51895_new_n336_), .Y(u1__abc_51895_new_n337_));
AND2X2 AND2X2_4880 ( .A(u2__abc_52155_new_n11556_), .B(u2__abc_52155_new_n4754_), .Y(u2__abc_52155_new_n11557_));
AND2X2 AND2X2_4881 ( .A(u2__abc_52155_new_n4748_), .B(u2__abc_52155_new_n11557_), .Y(u2__abc_52155_new_n11558_));
AND2X2 AND2X2_4882 ( .A(u2__abc_52155_new_n4746_), .B(u2__abc_52155_new_n4735_), .Y(u2__abc_52155_new_n11559_));
AND2X2 AND2X2_4883 ( .A(u2__abc_52155_new_n11411_), .B(u2__abc_52155_new_n4793_), .Y(u2__abc_52155_new_n11563_));
AND2X2 AND2X2_4884 ( .A(u2__abc_52155_new_n11564_), .B(u2__abc_52155_new_n4699_), .Y(u2__abc_52155_new_n11565_));
AND2X2 AND2X2_4885 ( .A(u2__abc_52155_new_n11567_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11568_));
AND2X2 AND2X2_4886 ( .A(u2__abc_52155_new_n11568_), .B(u2__abc_52155_new_n11566_), .Y(u2__abc_52155_new_n11569_));
AND2X2 AND2X2_4887 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_198_), .Y(u2__abc_52155_new_n11570_));
AND2X2 AND2X2_4888 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4674_), .Y(u2__abc_52155_new_n11573_));
AND2X2 AND2X2_4889 ( .A(u2__abc_52155_new_n11574_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11575_));
AND2X2 AND2X2_489 ( .A(u1__abc_51895_new_n330_), .B(u1__abc_51895_new_n337_), .Y(u1__abc_51895_new_n338_));
AND2X2 AND2X2_4890 ( .A(u2__abc_52155_new_n11572_), .B(u2__abc_52155_new_n11575_), .Y(u2__abc_52155_new_n11576_));
AND2X2 AND2X2_4891 ( .A(u2__abc_52155_new_n11577_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__200_));
AND2X2 AND2X2_4892 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_201_), .Y(u2__abc_52155_new_n11579_));
AND2X2 AND2X2_4893 ( .A(u2__abc_52155_new_n11566_), .B(u2__abc_52155_new_n4695_), .Y(u2__abc_52155_new_n11580_));
AND2X2 AND2X2_4894 ( .A(u2__abc_52155_new_n11580_), .B(u2__abc_52155_new_n4692_), .Y(u2__abc_52155_new_n11581_));
AND2X2 AND2X2_4895 ( .A(u2__abc_52155_new_n11583_), .B(u2__abc_52155_new_n11582_), .Y(u2__abc_52155_new_n11584_));
AND2X2 AND2X2_4896 ( .A(u2__abc_52155_new_n11585_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11586_));
AND2X2 AND2X2_4897 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_199_), .Y(u2__abc_52155_new_n11587_));
AND2X2 AND2X2_4898 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4681_), .Y(u2__abc_52155_new_n11590_));
AND2X2 AND2X2_4899 ( .A(u2__abc_52155_new_n11591_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11592_));
AND2X2 AND2X2_49 ( .A(_abc_73687_new_n753_), .B(sqrto_48_), .Y(\o[84] ));
AND2X2 AND2X2_490 ( .A(u1__abc_51895_new_n339_), .B(u1__abc_51895_new_n340_), .Y(u1__abc_51895_new_n341_));
AND2X2 AND2X2_4900 ( .A(u2__abc_52155_new_n11589_), .B(u2__abc_52155_new_n11592_), .Y(u2__abc_52155_new_n11593_));
AND2X2 AND2X2_4901 ( .A(u2__abc_52155_new_n11594_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__201_));
AND2X2 AND2X2_4902 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_202_), .Y(u2__abc_52155_new_n11596_));
AND2X2 AND2X2_4903 ( .A(u2__abc_52155_new_n4688_), .B(u2__abc_52155_new_n4695_), .Y(u2__abc_52155_new_n11597_));
AND2X2 AND2X2_4904 ( .A(u2__abc_52155_new_n11566_), .B(u2__abc_52155_new_n11597_), .Y(u2__abc_52155_new_n11598_));
AND2X2 AND2X2_4905 ( .A(u2__abc_52155_new_n11600_), .B(u2__abc_52155_new_n4677_), .Y(u2__abc_52155_new_n11601_));
AND2X2 AND2X2_4906 ( .A(u2__abc_52155_new_n11603_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11604_));
AND2X2 AND2X2_4907 ( .A(u2__abc_52155_new_n11604_), .B(u2__abc_52155_new_n11602_), .Y(u2__abc_52155_new_n11605_));
AND2X2 AND2X2_4908 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_200_), .Y(u2__abc_52155_new_n11606_));
AND2X2 AND2X2_4909 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4727_), .Y(u2__abc_52155_new_n11609_));
AND2X2 AND2X2_491 ( .A(u1__abc_51895_new_n342_), .B(u1__abc_51895_new_n343_), .Y(u1__abc_51895_new_n344_));
AND2X2 AND2X2_4910 ( .A(u2__abc_52155_new_n11610_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11611_));
AND2X2 AND2X2_4911 ( .A(u2__abc_52155_new_n11608_), .B(u2__abc_52155_new_n11611_), .Y(u2__abc_52155_new_n11612_));
AND2X2 AND2X2_4912 ( .A(u2__abc_52155_new_n11613_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__202_));
AND2X2 AND2X2_4913 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_203_), .Y(u2__abc_52155_new_n11615_));
AND2X2 AND2X2_4914 ( .A(u2__abc_52155_new_n11602_), .B(u2__abc_52155_new_n4673_), .Y(u2__abc_52155_new_n11616_));
AND2X2 AND2X2_4915 ( .A(u2__abc_52155_new_n11616_), .B(u2__abc_52155_new_n4684_), .Y(u2__abc_52155_new_n11617_));
AND2X2 AND2X2_4916 ( .A(u2__abc_52155_new_n11619_), .B(u2__abc_52155_new_n11618_), .Y(u2__abc_52155_new_n11620_));
AND2X2 AND2X2_4917 ( .A(u2__abc_52155_new_n11621_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11622_));
AND2X2 AND2X2_4918 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_201_), .Y(u2__abc_52155_new_n11623_));
AND2X2 AND2X2_4919 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4720_), .Y(u2__abc_52155_new_n11626_));
AND2X2 AND2X2_492 ( .A(u1__abc_51895_new_n341_), .B(u1__abc_51895_new_n344_), .Y(u1__abc_51895_new_n345_));
AND2X2 AND2X2_4920 ( .A(u2__abc_52155_new_n11627_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11628_));
AND2X2 AND2X2_4921 ( .A(u2__abc_52155_new_n11625_), .B(u2__abc_52155_new_n11628_), .Y(u2__abc_52155_new_n11629_));
AND2X2 AND2X2_4922 ( .A(u2__abc_52155_new_n11630_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__203_));
AND2X2 AND2X2_4923 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_204_), .Y(u2__abc_52155_new_n11632_));
AND2X2 AND2X2_4924 ( .A(u2__abc_52155_new_n11634_), .B(u2__abc_52155_new_n4685_), .Y(u2__abc_52155_new_n11635_));
AND2X2 AND2X2_4925 ( .A(u2__abc_52155_new_n4683_), .B(u2__abc_52155_new_n4672_), .Y(u2__abc_52155_new_n11636_));
AND2X2 AND2X2_4926 ( .A(u2__abc_52155_new_n11564_), .B(u2__abc_52155_new_n4701_), .Y(u2__abc_52155_new_n11639_));
AND2X2 AND2X2_4927 ( .A(u2__abc_52155_new_n11640_), .B(u2__abc_52155_new_n4730_), .Y(u2__abc_52155_new_n11641_));
AND2X2 AND2X2_4928 ( .A(u2__abc_52155_new_n11643_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11644_));
AND2X2 AND2X2_4929 ( .A(u2__abc_52155_new_n11644_), .B(u2__abc_52155_new_n11642_), .Y(u2__abc_52155_new_n11645_));
AND2X2 AND2X2_493 ( .A(u1__abc_51895_new_n346_), .B(u1__abc_51895_new_n347_), .Y(u1__abc_51895_new_n348_));
AND2X2 AND2X2_4930 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_202_), .Y(u2__abc_52155_new_n11646_));
AND2X2 AND2X2_4931 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4705_), .Y(u2__abc_52155_new_n11649_));
AND2X2 AND2X2_4932 ( .A(u2__abc_52155_new_n11650_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11651_));
AND2X2 AND2X2_4933 ( .A(u2__abc_52155_new_n11648_), .B(u2__abc_52155_new_n11651_), .Y(u2__abc_52155_new_n11652_));
AND2X2 AND2X2_4934 ( .A(u2__abc_52155_new_n11653_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__204_));
AND2X2 AND2X2_4935 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_205_), .Y(u2__abc_52155_new_n11655_));
AND2X2 AND2X2_4936 ( .A(u2__abc_52155_new_n11642_), .B(u2__abc_52155_new_n4726_), .Y(u2__abc_52155_new_n11656_));
AND2X2 AND2X2_4937 ( .A(u2__abc_52155_new_n11656_), .B(u2__abc_52155_new_n4723_), .Y(u2__abc_52155_new_n11657_));
AND2X2 AND2X2_4938 ( .A(u2__abc_52155_new_n11659_), .B(u2__abc_52155_new_n11658_), .Y(u2__abc_52155_new_n11660_));
AND2X2 AND2X2_4939 ( .A(u2__abc_52155_new_n11661_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11662_));
AND2X2 AND2X2_494 ( .A(u1__abc_51895_new_n349_), .B(u1__abc_51895_new_n350_), .Y(u1__abc_51895_new_n351_));
AND2X2 AND2X2_4940 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_203_), .Y(u2__abc_52155_new_n11663_));
AND2X2 AND2X2_4941 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4712_), .Y(u2__abc_52155_new_n11666_));
AND2X2 AND2X2_4942 ( .A(u2__abc_52155_new_n11667_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11668_));
AND2X2 AND2X2_4943 ( .A(u2__abc_52155_new_n11665_), .B(u2__abc_52155_new_n11668_), .Y(u2__abc_52155_new_n11669_));
AND2X2 AND2X2_4944 ( .A(u2__abc_52155_new_n11670_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__205_));
AND2X2 AND2X2_4945 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_206_), .Y(u2__abc_52155_new_n11672_));
AND2X2 AND2X2_4946 ( .A(u2__abc_52155_new_n4719_), .B(u2__abc_52155_new_n4726_), .Y(u2__abc_52155_new_n11673_));
AND2X2 AND2X2_4947 ( .A(u2__abc_52155_new_n11642_), .B(u2__abc_52155_new_n11673_), .Y(u2__abc_52155_new_n11674_));
AND2X2 AND2X2_4948 ( .A(u2__abc_52155_new_n11676_), .B(u2__abc_52155_new_n4708_), .Y(u2__abc_52155_new_n11677_));
AND2X2 AND2X2_4949 ( .A(u2__abc_52155_new_n11679_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11680_));
AND2X2 AND2X2_495 ( .A(u1__abc_51895_new_n348_), .B(u1__abc_51895_new_n351_), .Y(u1__abc_51895_new_n352_));
AND2X2 AND2X2_4950 ( .A(u2__abc_52155_new_n11680_), .B(u2__abc_52155_new_n11678_), .Y(u2__abc_52155_new_n11681_));
AND2X2 AND2X2_4951 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_204_), .Y(u2__abc_52155_new_n11682_));
AND2X2 AND2X2_4952 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4625_), .Y(u2__abc_52155_new_n11685_));
AND2X2 AND2X2_4953 ( .A(u2__abc_52155_new_n11686_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11687_));
AND2X2 AND2X2_4954 ( .A(u2__abc_52155_new_n11684_), .B(u2__abc_52155_new_n11687_), .Y(u2__abc_52155_new_n11688_));
AND2X2 AND2X2_4955 ( .A(u2__abc_52155_new_n11689_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__206_));
AND2X2 AND2X2_4956 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_207_), .Y(u2__abc_52155_new_n11691_));
AND2X2 AND2X2_4957 ( .A(u2__abc_52155_new_n11678_), .B(u2__abc_52155_new_n4704_), .Y(u2__abc_52155_new_n11692_));
AND2X2 AND2X2_4958 ( .A(u2__abc_52155_new_n11692_), .B(u2__abc_52155_new_n4715_), .Y(u2__abc_52155_new_n11693_));
AND2X2 AND2X2_4959 ( .A(u2__abc_52155_new_n11695_), .B(u2__abc_52155_new_n11694_), .Y(u2__abc_52155_new_n11696_));
AND2X2 AND2X2_496 ( .A(u1__abc_51895_new_n345_), .B(u1__abc_51895_new_n352_), .Y(u1__abc_51895_new_n353_));
AND2X2 AND2X2_4960 ( .A(u2__abc_52155_new_n11697_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11698_));
AND2X2 AND2X2_4961 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_205_), .Y(u2__abc_52155_new_n11699_));
AND2X2 AND2X2_4962 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4632_), .Y(u2__abc_52155_new_n11702_));
AND2X2 AND2X2_4963 ( .A(u2__abc_52155_new_n11703_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11704_));
AND2X2 AND2X2_4964 ( .A(u2__abc_52155_new_n11701_), .B(u2__abc_52155_new_n11704_), .Y(u2__abc_52155_new_n11705_));
AND2X2 AND2X2_4965 ( .A(u2__abc_52155_new_n11706_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__207_));
AND2X2 AND2X2_4966 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_208_), .Y(u2__abc_52155_new_n11708_));
AND2X2 AND2X2_4967 ( .A(u2__abc_52155_new_n11562_), .B(u2__abc_52155_new_n4733_), .Y(u2__abc_52155_new_n11709_));
AND2X2 AND2X2_4968 ( .A(u2__abc_52155_new_n11638_), .B(u2__abc_52155_new_n4732_), .Y(u2__abc_52155_new_n11710_));
AND2X2 AND2X2_4969 ( .A(u2__abc_52155_new_n11712_), .B(u2__abc_52155_new_n4716_), .Y(u2__abc_52155_new_n11713_));
AND2X2 AND2X2_497 ( .A(u1__abc_51895_new_n338_), .B(u1__abc_51895_new_n353_), .Y(u1__abc_51895_new_n354_));
AND2X2 AND2X2_4970 ( .A(u2__abc_52155_new_n4714_), .B(u2__abc_52155_new_n4703_), .Y(u2__abc_52155_new_n11714_));
AND2X2 AND2X2_4971 ( .A(u2__abc_52155_new_n11411_), .B(u2__abc_52155_new_n4794_), .Y(u2__abc_52155_new_n11719_));
AND2X2 AND2X2_4972 ( .A(u2__abc_52155_new_n11720_), .B(u2__abc_52155_new_n4628_), .Y(u2__abc_52155_new_n11721_));
AND2X2 AND2X2_4973 ( .A(u2__abc_52155_new_n11723_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11724_));
AND2X2 AND2X2_4974 ( .A(u2__abc_52155_new_n11724_), .B(u2__abc_52155_new_n11722_), .Y(u2__abc_52155_new_n11725_));
AND2X2 AND2X2_4975 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_206_), .Y(u2__abc_52155_new_n11726_));
AND2X2 AND2X2_4976 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4610_), .Y(u2__abc_52155_new_n11729_));
AND2X2 AND2X2_4977 ( .A(u2__abc_52155_new_n11730_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11731_));
AND2X2 AND2X2_4978 ( .A(u2__abc_52155_new_n11728_), .B(u2__abc_52155_new_n11731_), .Y(u2__abc_52155_new_n11732_));
AND2X2 AND2X2_4979 ( .A(u2__abc_52155_new_n11733_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__208_));
AND2X2 AND2X2_498 ( .A(u1__abc_51895_new_n355_), .B(u1__abc_51895_new_n356_), .Y(u1__abc_51895_new_n357_));
AND2X2 AND2X2_4980 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_209_), .Y(u2__abc_52155_new_n11735_));
AND2X2 AND2X2_4981 ( .A(u2__abc_52155_new_n11722_), .B(u2__abc_52155_new_n4624_), .Y(u2__abc_52155_new_n11737_));
AND2X2 AND2X2_4982 ( .A(u2__abc_52155_new_n11738_), .B(u2__abc_52155_new_n11736_), .Y(u2__abc_52155_new_n11739_));
AND2X2 AND2X2_4983 ( .A(u2__abc_52155_new_n11737_), .B(u2__abc_52155_new_n4635_), .Y(u2__abc_52155_new_n11740_));
AND2X2 AND2X2_4984 ( .A(u2__abc_52155_new_n11741_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11742_));
AND2X2 AND2X2_4985 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_207_), .Y(u2__abc_52155_new_n11743_));
AND2X2 AND2X2_4986 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4617_), .Y(u2__abc_52155_new_n11746_));
AND2X2 AND2X2_4987 ( .A(u2__abc_52155_new_n11747_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11748_));
AND2X2 AND2X2_4988 ( .A(u2__abc_52155_new_n11745_), .B(u2__abc_52155_new_n11748_), .Y(u2__abc_52155_new_n11749_));
AND2X2 AND2X2_4989 ( .A(u2__abc_52155_new_n11750_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__209_));
AND2X2 AND2X2_499 ( .A(u1__abc_51895_new_n358_), .B(u1__abc_51895_new_n359_), .Y(u1__abc_51895_new_n360_));
AND2X2 AND2X2_4990 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_210_), .Y(u2__abc_52155_new_n11752_));
AND2X2 AND2X2_4991 ( .A(u2__abc_52155_new_n4624_), .B(u2__abc_52155_new_n4631_), .Y(u2__abc_52155_new_n11753_));
AND2X2 AND2X2_4992 ( .A(u2__abc_52155_new_n11720_), .B(u2__abc_52155_new_n4636_), .Y(u2__abc_52155_new_n11756_));
AND2X2 AND2X2_4993 ( .A(u2__abc_52155_new_n11757_), .B(u2__abc_52155_new_n4613_), .Y(u2__abc_52155_new_n11758_));
AND2X2 AND2X2_4994 ( .A(u2__abc_52155_new_n11760_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11761_));
AND2X2 AND2X2_4995 ( .A(u2__abc_52155_new_n11761_), .B(u2__abc_52155_new_n11759_), .Y(u2__abc_52155_new_n11762_));
AND2X2 AND2X2_4996 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_208_), .Y(u2__abc_52155_new_n11763_));
AND2X2 AND2X2_4997 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4663_), .Y(u2__abc_52155_new_n11766_));
AND2X2 AND2X2_4998 ( .A(u2__abc_52155_new_n11767_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11768_));
AND2X2 AND2X2_4999 ( .A(u2__abc_52155_new_n11765_), .B(u2__abc_52155_new_n11768_), .Y(u2__abc_52155_new_n11769_));
AND2X2 AND2X2_5 ( .A(_abc_73687_new_n753_), .B(sqrto_4_), .Y(\o[40] ));
AND2X2 AND2X2_50 ( .A(_abc_73687_new_n753_), .B(sqrto_49_), .Y(\o[85] ));
AND2X2 AND2X2_500 ( .A(u1__abc_51895_new_n357_), .B(u1__abc_51895_new_n360_), .Y(u1__abc_51895_new_n361_));
AND2X2 AND2X2_5000 ( .A(u2__abc_52155_new_n11770_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__210_));
AND2X2 AND2X2_5001 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_211_), .Y(u2__abc_52155_new_n11772_));
AND2X2 AND2X2_5002 ( .A(u2__abc_52155_new_n11759_), .B(u2__abc_52155_new_n4609_), .Y(u2__abc_52155_new_n11773_));
AND2X2 AND2X2_5003 ( .A(u2__abc_52155_new_n11773_), .B(u2__abc_52155_new_n4620_), .Y(u2__abc_52155_new_n11774_));
AND2X2 AND2X2_5004 ( .A(u2__abc_52155_new_n11776_), .B(u2__abc_52155_new_n11775_), .Y(u2__abc_52155_new_n11777_));
AND2X2 AND2X2_5005 ( .A(u2__abc_52155_new_n11778_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11779_));
AND2X2 AND2X2_5006 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_209_), .Y(u2__abc_52155_new_n11780_));
AND2X2 AND2X2_5007 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4656_), .Y(u2__abc_52155_new_n11783_));
AND2X2 AND2X2_5008 ( .A(u2__abc_52155_new_n11784_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11785_));
AND2X2 AND2X2_5009 ( .A(u2__abc_52155_new_n11782_), .B(u2__abc_52155_new_n11785_), .Y(u2__abc_52155_new_n11786_));
AND2X2 AND2X2_501 ( .A(u1__abc_51895_new_n362_), .B(u1__abc_51895_new_n363_), .Y(u1__abc_51895_new_n364_));
AND2X2 AND2X2_5010 ( .A(u2__abc_52155_new_n11787_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__211_));
AND2X2 AND2X2_5011 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_212_), .Y(u2__abc_52155_new_n11789_));
AND2X2 AND2X2_5012 ( .A(u2__abc_52155_new_n11755_), .B(u2__abc_52155_new_n4621_), .Y(u2__abc_52155_new_n11790_));
AND2X2 AND2X2_5013 ( .A(u2__abc_52155_new_n4619_), .B(u2__abc_52155_new_n4608_), .Y(u2__abc_52155_new_n11791_));
AND2X2 AND2X2_5014 ( .A(u2__abc_52155_new_n11720_), .B(u2__abc_52155_new_n4637_), .Y(u2__abc_52155_new_n11794_));
AND2X2 AND2X2_5015 ( .A(u2__abc_52155_new_n11795_), .B(u2__abc_52155_new_n4666_), .Y(u2__abc_52155_new_n11796_));
AND2X2 AND2X2_5016 ( .A(u2__abc_52155_new_n11798_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11799_));
AND2X2 AND2X2_5017 ( .A(u2__abc_52155_new_n11799_), .B(u2__abc_52155_new_n11797_), .Y(u2__abc_52155_new_n11800_));
AND2X2 AND2X2_5018 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_210_), .Y(u2__abc_52155_new_n11801_));
AND2X2 AND2X2_5019 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4641_), .Y(u2__abc_52155_new_n11804_));
AND2X2 AND2X2_502 ( .A(u1__abc_51895_new_n365_), .B(u1__abc_51895_new_n366_), .Y(u1__abc_51895_new_n367_));
AND2X2 AND2X2_5020 ( .A(u2__abc_52155_new_n11805_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11806_));
AND2X2 AND2X2_5021 ( .A(u2__abc_52155_new_n11803_), .B(u2__abc_52155_new_n11806_), .Y(u2__abc_52155_new_n11807_));
AND2X2 AND2X2_5022 ( .A(u2__abc_52155_new_n11808_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__212_));
AND2X2 AND2X2_5023 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_213_), .Y(u2__abc_52155_new_n11810_));
AND2X2 AND2X2_5024 ( .A(u2__abc_52155_new_n11797_), .B(u2__abc_52155_new_n4662_), .Y(u2__abc_52155_new_n11811_));
AND2X2 AND2X2_5025 ( .A(u2__abc_52155_new_n11812_), .B(u2__abc_52155_new_n4659_), .Y(u2__abc_52155_new_n11813_));
AND2X2 AND2X2_5026 ( .A(u2__abc_52155_new_n11815_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11816_));
AND2X2 AND2X2_5027 ( .A(u2__abc_52155_new_n11816_), .B(u2__abc_52155_new_n11814_), .Y(u2__abc_52155_new_n11817_));
AND2X2 AND2X2_5028 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_211_), .Y(u2__abc_52155_new_n11818_));
AND2X2 AND2X2_5029 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4648_), .Y(u2__abc_52155_new_n11821_));
AND2X2 AND2X2_503 ( .A(u1__abc_51895_new_n364_), .B(u1__abc_51895_new_n367_), .Y(u1__abc_51895_new_n368_));
AND2X2 AND2X2_5030 ( .A(u2__abc_52155_new_n11822_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11823_));
AND2X2 AND2X2_5031 ( .A(u2__abc_52155_new_n11820_), .B(u2__abc_52155_new_n11823_), .Y(u2__abc_52155_new_n11824_));
AND2X2 AND2X2_5032 ( .A(u2__abc_52155_new_n11825_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__213_));
AND2X2 AND2X2_5033 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_214_), .Y(u2__abc_52155_new_n11827_));
AND2X2 AND2X2_5034 ( .A(u2__abc_52155_new_n11814_), .B(u2__abc_52155_new_n4655_), .Y(u2__abc_52155_new_n11828_));
AND2X2 AND2X2_5035 ( .A(u2__abc_52155_new_n11829_), .B(u2__abc_52155_new_n4644_), .Y(u2__abc_52155_new_n11830_));
AND2X2 AND2X2_5036 ( .A(u2__abc_52155_new_n11832_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11833_));
AND2X2 AND2X2_5037 ( .A(u2__abc_52155_new_n11833_), .B(u2__abc_52155_new_n11831_), .Y(u2__abc_52155_new_n11834_));
AND2X2 AND2X2_5038 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_212_), .Y(u2__abc_52155_new_n11835_));
AND2X2 AND2X2_5039 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4562_), .Y(u2__abc_52155_new_n11838_));
AND2X2 AND2X2_504 ( .A(u1__abc_51895_new_n361_), .B(u1__abc_51895_new_n368_), .Y(u1__abc_51895_new_n369_));
AND2X2 AND2X2_5040 ( .A(u2__abc_52155_new_n11839_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11840_));
AND2X2 AND2X2_5041 ( .A(u2__abc_52155_new_n11837_), .B(u2__abc_52155_new_n11840_), .Y(u2__abc_52155_new_n11841_));
AND2X2 AND2X2_5042 ( .A(u2__abc_52155_new_n11842_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__214_));
AND2X2 AND2X2_5043 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_215_), .Y(u2__abc_52155_new_n11844_));
AND2X2 AND2X2_5044 ( .A(u2__abc_52155_new_n11831_), .B(u2__abc_52155_new_n4640_), .Y(u2__abc_52155_new_n11845_));
AND2X2 AND2X2_5045 ( .A(u2__abc_52155_new_n11845_), .B(u2__abc_52155_new_n4651_), .Y(u2__abc_52155_new_n11846_));
AND2X2 AND2X2_5046 ( .A(u2__abc_52155_new_n11848_), .B(u2__abc_52155_new_n11847_), .Y(u2__abc_52155_new_n11849_));
AND2X2 AND2X2_5047 ( .A(u2__abc_52155_new_n11850_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11851_));
AND2X2 AND2X2_5048 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_213_), .Y(u2__abc_52155_new_n11852_));
AND2X2 AND2X2_5049 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4569_), .Y(u2__abc_52155_new_n11855_));
AND2X2 AND2X2_505 ( .A(u1__abc_51895_new_n370_), .B(u1__abc_51895_new_n371_), .Y(u1__abc_51895_new_n372_));
AND2X2 AND2X2_5050 ( .A(u2__abc_52155_new_n11856_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11857_));
AND2X2 AND2X2_5051 ( .A(u2__abc_52155_new_n11854_), .B(u2__abc_52155_new_n11857_), .Y(u2__abc_52155_new_n11858_));
AND2X2 AND2X2_5052 ( .A(u2__abc_52155_new_n11859_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__215_));
AND2X2 AND2X2_5053 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_216_), .Y(u2__abc_52155_new_n11861_));
AND2X2 AND2X2_5054 ( .A(u2__abc_52155_new_n11793_), .B(u2__abc_52155_new_n4668_), .Y(u2__abc_52155_new_n11862_));
AND2X2 AND2X2_5055 ( .A(u2__abc_52155_new_n11863_), .B(u2__abc_52155_new_n4658_), .Y(u2__abc_52155_new_n11864_));
AND2X2 AND2X2_5056 ( .A(u2__abc_52155_new_n4652_), .B(u2__abc_52155_new_n11864_), .Y(u2__abc_52155_new_n11865_));
AND2X2 AND2X2_5057 ( .A(u2__abc_52155_new_n4650_), .B(u2__abc_52155_new_n4639_), .Y(u2__abc_52155_new_n11866_));
AND2X2 AND2X2_5058 ( .A(u2__abc_52155_new_n11720_), .B(u2__abc_52155_new_n4669_), .Y(u2__abc_52155_new_n11870_));
AND2X2 AND2X2_5059 ( .A(u2__abc_52155_new_n11871_), .B(u2__abc_52155_new_n4565_), .Y(u2__abc_52155_new_n11872_));
AND2X2 AND2X2_506 ( .A(u1__abc_51895_new_n373_), .B(u1__abc_51895_new_n374_), .Y(u1__abc_51895_new_n375_));
AND2X2 AND2X2_5060 ( .A(u2__abc_52155_new_n11874_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11875_));
AND2X2 AND2X2_5061 ( .A(u2__abc_52155_new_n11875_), .B(u2__abc_52155_new_n11873_), .Y(u2__abc_52155_new_n11876_));
AND2X2 AND2X2_5062 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_214_), .Y(u2__abc_52155_new_n11877_));
AND2X2 AND2X2_5063 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4547_), .Y(u2__abc_52155_new_n11880_));
AND2X2 AND2X2_5064 ( .A(u2__abc_52155_new_n11881_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11882_));
AND2X2 AND2X2_5065 ( .A(u2__abc_52155_new_n11879_), .B(u2__abc_52155_new_n11882_), .Y(u2__abc_52155_new_n11883_));
AND2X2 AND2X2_5066 ( .A(u2__abc_52155_new_n11884_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__216_));
AND2X2 AND2X2_5067 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_217_), .Y(u2__abc_52155_new_n11886_));
AND2X2 AND2X2_5068 ( .A(u2__abc_52155_new_n11873_), .B(u2__abc_52155_new_n4561_), .Y(u2__abc_52155_new_n11888_));
AND2X2 AND2X2_5069 ( .A(u2__abc_52155_new_n11889_), .B(u2__abc_52155_new_n11887_), .Y(u2__abc_52155_new_n11890_));
AND2X2 AND2X2_507 ( .A(u1__abc_51895_new_n372_), .B(u1__abc_51895_new_n375_), .Y(u1__abc_51895_new_n376_));
AND2X2 AND2X2_5070 ( .A(u2__abc_52155_new_n11888_), .B(u2__abc_52155_new_n4572_), .Y(u2__abc_52155_new_n11891_));
AND2X2 AND2X2_5071 ( .A(u2__abc_52155_new_n11892_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11893_));
AND2X2 AND2X2_5072 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_215_), .Y(u2__abc_52155_new_n11894_));
AND2X2 AND2X2_5073 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4554_), .Y(u2__abc_52155_new_n11897_));
AND2X2 AND2X2_5074 ( .A(u2__abc_52155_new_n11898_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11899_));
AND2X2 AND2X2_5075 ( .A(u2__abc_52155_new_n11896_), .B(u2__abc_52155_new_n11899_), .Y(u2__abc_52155_new_n11900_));
AND2X2 AND2X2_5076 ( .A(u2__abc_52155_new_n11901_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__217_));
AND2X2 AND2X2_5077 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_218_), .Y(u2__abc_52155_new_n11903_));
AND2X2 AND2X2_5078 ( .A(u2__abc_52155_new_n4561_), .B(u2__abc_52155_new_n4568_), .Y(u2__abc_52155_new_n11904_));
AND2X2 AND2X2_5079 ( .A(u2__abc_52155_new_n11871_), .B(u2__abc_52155_new_n4573_), .Y(u2__abc_52155_new_n11907_));
AND2X2 AND2X2_508 ( .A(u1__abc_51895_new_n377_), .B(u1__abc_51895_new_n378_), .Y(u1__abc_51895_new_n379_));
AND2X2 AND2X2_5080 ( .A(u2__abc_52155_new_n11908_), .B(u2__abc_52155_new_n4550_), .Y(u2__abc_52155_new_n11909_));
AND2X2 AND2X2_5081 ( .A(u2__abc_52155_new_n11911_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11912_));
AND2X2 AND2X2_5082 ( .A(u2__abc_52155_new_n11912_), .B(u2__abc_52155_new_n11910_), .Y(u2__abc_52155_new_n11913_));
AND2X2 AND2X2_5083 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_216_), .Y(u2__abc_52155_new_n11914_));
AND2X2 AND2X2_5084 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4600_), .Y(u2__abc_52155_new_n11917_));
AND2X2 AND2X2_5085 ( .A(u2__abc_52155_new_n11918_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11919_));
AND2X2 AND2X2_5086 ( .A(u2__abc_52155_new_n11916_), .B(u2__abc_52155_new_n11919_), .Y(u2__abc_52155_new_n11920_));
AND2X2 AND2X2_5087 ( .A(u2__abc_52155_new_n11921_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__218_));
AND2X2 AND2X2_5088 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_219_), .Y(u2__abc_52155_new_n11923_));
AND2X2 AND2X2_5089 ( .A(u2__abc_52155_new_n11910_), .B(u2__abc_52155_new_n4546_), .Y(u2__abc_52155_new_n11924_));
AND2X2 AND2X2_509 ( .A(u1__abc_51895_new_n380_), .B(u1__abc_51895_new_n381_), .Y(u1__abc_51895_new_n382_));
AND2X2 AND2X2_5090 ( .A(u2__abc_52155_new_n11924_), .B(u2__abc_52155_new_n4557_), .Y(u2__abc_52155_new_n11925_));
AND2X2 AND2X2_5091 ( .A(u2__abc_52155_new_n11927_), .B(u2__abc_52155_new_n11926_), .Y(u2__abc_52155_new_n11928_));
AND2X2 AND2X2_5092 ( .A(u2__abc_52155_new_n11929_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11930_));
AND2X2 AND2X2_5093 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_217_), .Y(u2__abc_52155_new_n11931_));
AND2X2 AND2X2_5094 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4593_), .Y(u2__abc_52155_new_n11934_));
AND2X2 AND2X2_5095 ( .A(u2__abc_52155_new_n11935_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11936_));
AND2X2 AND2X2_5096 ( .A(u2__abc_52155_new_n11933_), .B(u2__abc_52155_new_n11936_), .Y(u2__abc_52155_new_n11937_));
AND2X2 AND2X2_5097 ( .A(u2__abc_52155_new_n11938_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__219_));
AND2X2 AND2X2_5098 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_220_), .Y(u2__abc_52155_new_n11940_));
AND2X2 AND2X2_5099 ( .A(u2__abc_52155_new_n11906_), .B(u2__abc_52155_new_n4558_), .Y(u2__abc_52155_new_n11941_));
AND2X2 AND2X2_51 ( .A(_abc_73687_new_n753_), .B(sqrto_50_), .Y(\o[86] ));
AND2X2 AND2X2_510 ( .A(u1__abc_51895_new_n379_), .B(u1__abc_51895_new_n382_), .Y(u1__abc_51895_new_n383_));
AND2X2 AND2X2_5100 ( .A(u2__abc_52155_new_n4556_), .B(u2__abc_52155_new_n4545_), .Y(u2__abc_52155_new_n11942_));
AND2X2 AND2X2_5101 ( .A(u2__abc_52155_new_n11871_), .B(u2__abc_52155_new_n4574_), .Y(u2__abc_52155_new_n11945_));
AND2X2 AND2X2_5102 ( .A(u2__abc_52155_new_n11946_), .B(u2__abc_52155_new_n4603_), .Y(u2__abc_52155_new_n11947_));
AND2X2 AND2X2_5103 ( .A(u2__abc_52155_new_n11949_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11950_));
AND2X2 AND2X2_5104 ( .A(u2__abc_52155_new_n11950_), .B(u2__abc_52155_new_n11948_), .Y(u2__abc_52155_new_n11951_));
AND2X2 AND2X2_5105 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_218_), .Y(u2__abc_52155_new_n11952_));
AND2X2 AND2X2_5106 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4578_), .Y(u2__abc_52155_new_n11955_));
AND2X2 AND2X2_5107 ( .A(u2__abc_52155_new_n11956_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11957_));
AND2X2 AND2X2_5108 ( .A(u2__abc_52155_new_n11954_), .B(u2__abc_52155_new_n11957_), .Y(u2__abc_52155_new_n11958_));
AND2X2 AND2X2_5109 ( .A(u2__abc_52155_new_n11959_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__220_));
AND2X2 AND2X2_511 ( .A(u1__abc_51895_new_n376_), .B(u1__abc_51895_new_n383_), .Y(u1__abc_51895_new_n384_));
AND2X2 AND2X2_5110 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_221_), .Y(u2__abc_52155_new_n11961_));
AND2X2 AND2X2_5111 ( .A(u2__abc_52155_new_n11948_), .B(u2__abc_52155_new_n4599_), .Y(u2__abc_52155_new_n11962_));
AND2X2 AND2X2_5112 ( .A(u2__abc_52155_new_n11962_), .B(u2__abc_52155_new_n4596_), .Y(u2__abc_52155_new_n11963_));
AND2X2 AND2X2_5113 ( .A(u2__abc_52155_new_n11965_), .B(u2__abc_52155_new_n11964_), .Y(u2__abc_52155_new_n11966_));
AND2X2 AND2X2_5114 ( .A(u2__abc_52155_new_n11967_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11968_));
AND2X2 AND2X2_5115 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_219_), .Y(u2__abc_52155_new_n11969_));
AND2X2 AND2X2_5116 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4585_), .Y(u2__abc_52155_new_n11972_));
AND2X2 AND2X2_5117 ( .A(u2__abc_52155_new_n11973_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11974_));
AND2X2 AND2X2_5118 ( .A(u2__abc_52155_new_n11971_), .B(u2__abc_52155_new_n11974_), .Y(u2__abc_52155_new_n11975_));
AND2X2 AND2X2_5119 ( .A(u2__abc_52155_new_n11976_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__221_));
AND2X2 AND2X2_512 ( .A(u1__abc_51895_new_n369_), .B(u1__abc_51895_new_n384_), .Y(u1__abc_51895_new_n385_));
AND2X2 AND2X2_5120 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_222_), .Y(u2__abc_52155_new_n11978_));
AND2X2 AND2X2_5121 ( .A(u2__abc_52155_new_n4592_), .B(u2__abc_52155_new_n4599_), .Y(u2__abc_52155_new_n11979_));
AND2X2 AND2X2_5122 ( .A(u2__abc_52155_new_n11948_), .B(u2__abc_52155_new_n11979_), .Y(u2__abc_52155_new_n11980_));
AND2X2 AND2X2_5123 ( .A(u2__abc_52155_new_n11982_), .B(u2__abc_52155_new_n4581_), .Y(u2__abc_52155_new_n11983_));
AND2X2 AND2X2_5124 ( .A(u2__abc_52155_new_n11985_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n11986_));
AND2X2 AND2X2_5125 ( .A(u2__abc_52155_new_n11986_), .B(u2__abc_52155_new_n11984_), .Y(u2__abc_52155_new_n11987_));
AND2X2 AND2X2_5126 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_220_), .Y(u2__abc_52155_new_n11988_));
AND2X2 AND2X2_5127 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4504_), .Y(u2__abc_52155_new_n11991_));
AND2X2 AND2X2_5128 ( .A(u2__abc_52155_new_n11992_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n11993_));
AND2X2 AND2X2_5129 ( .A(u2__abc_52155_new_n11990_), .B(u2__abc_52155_new_n11993_), .Y(u2__abc_52155_new_n11994_));
AND2X2 AND2X2_513 ( .A(u1__abc_51895_new_n354_), .B(u1__abc_51895_new_n385_), .Y(u1__abc_51895_new_n386_));
AND2X2 AND2X2_5130 ( .A(u2__abc_52155_new_n11995_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__222_));
AND2X2 AND2X2_5131 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_223_), .Y(u2__abc_52155_new_n11997_));
AND2X2 AND2X2_5132 ( .A(u2__abc_52155_new_n11984_), .B(u2__abc_52155_new_n4577_), .Y(u2__abc_52155_new_n11998_));
AND2X2 AND2X2_5133 ( .A(u2__abc_52155_new_n11998_), .B(u2__abc_52155_new_n4588_), .Y(u2__abc_52155_new_n11999_));
AND2X2 AND2X2_5134 ( .A(u2__abc_52155_new_n12001_), .B(u2__abc_52155_new_n12000_), .Y(u2__abc_52155_new_n12002_));
AND2X2 AND2X2_5135 ( .A(u2__abc_52155_new_n12003_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12004_));
AND2X2 AND2X2_5136 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_221_), .Y(u2__abc_52155_new_n12005_));
AND2X2 AND2X2_5137 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4497_), .Y(u2__abc_52155_new_n12008_));
AND2X2 AND2X2_5138 ( .A(u2__abc_52155_new_n12009_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12010_));
AND2X2 AND2X2_5139 ( .A(u2__abc_52155_new_n12007_), .B(u2__abc_52155_new_n12010_), .Y(u2__abc_52155_new_n12011_));
AND2X2 AND2X2_514 ( .A(u1__abc_51895_new_n323_), .B(u1__abc_51895_new_n386_), .Y(u1__abc_51895_new_n387_));
AND2X2 AND2X2_5140 ( .A(u2__abc_52155_new_n12012_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__223_));
AND2X2 AND2X2_5141 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_224_), .Y(u2__abc_52155_new_n12014_));
AND2X2 AND2X2_5142 ( .A(u2__abc_52155_new_n11718_), .B(u2__abc_52155_new_n4670_), .Y(u2__abc_52155_new_n12015_));
AND2X2 AND2X2_5143 ( .A(u2__abc_52155_new_n11869_), .B(u2__abc_52155_new_n4606_), .Y(u2__abc_52155_new_n12017_));
AND2X2 AND2X2_5144 ( .A(u2__abc_52155_new_n11944_), .B(u2__abc_52155_new_n4605_), .Y(u2__abc_52155_new_n12019_));
AND2X2 AND2X2_5145 ( .A(u2__abc_52155_new_n4577_), .B(u2__abc_52155_new_n4584_), .Y(u2__abc_52155_new_n12021_));
AND2X2 AND2X2_5146 ( .A(u2__abc_52155_new_n12024_), .B(u2__abc_52155_new_n4589_), .Y(u2__abc_52155_new_n12025_));
AND2X2 AND2X2_5147 ( .A(u2__abc_52155_new_n12026_), .B(u2__abc_52155_new_n12022_), .Y(u2__abc_52155_new_n12027_));
AND2X2 AND2X2_5148 ( .A(u2__abc_52155_new_n12020_), .B(u2__abc_52155_new_n12027_), .Y(u2__abc_52155_new_n12028_));
AND2X2 AND2X2_5149 ( .A(u2__abc_52155_new_n12018_), .B(u2__abc_52155_new_n12028_), .Y(u2__abc_52155_new_n12029_));
AND2X2 AND2X2_515 ( .A(u1__abc_51895_new_n387_), .B(u1__abc_51895_new_n260_), .Y(u1_mz));
AND2X2 AND2X2_5150 ( .A(u2__abc_52155_new_n12016_), .B(u2__abc_52155_new_n12029_), .Y(u2__abc_52155_new_n12030_));
AND2X2 AND2X2_5151 ( .A(u2__abc_52155_new_n11411_), .B(u2__abc_52155_new_n4795_), .Y(u2__abc_52155_new_n12032_));
AND2X2 AND2X2_5152 ( .A(u2__abc_52155_new_n12033_), .B(u2__abc_52155_new_n4507_), .Y(u2__abc_52155_new_n12034_));
AND2X2 AND2X2_5153 ( .A(u2__abc_52155_new_n12036_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12037_));
AND2X2 AND2X2_5154 ( .A(u2__abc_52155_new_n12037_), .B(u2__abc_52155_new_n12035_), .Y(u2__abc_52155_new_n12038_));
AND2X2 AND2X2_5155 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_222_), .Y(u2__abc_52155_new_n12039_));
AND2X2 AND2X2_5156 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4482_), .Y(u2__abc_52155_new_n12042_));
AND2X2 AND2X2_5157 ( .A(u2__abc_52155_new_n12043_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12044_));
AND2X2 AND2X2_5158 ( .A(u2__abc_52155_new_n12041_), .B(u2__abc_52155_new_n12044_), .Y(u2__abc_52155_new_n12045_));
AND2X2 AND2X2_5159 ( .A(u2__abc_52155_new_n12046_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__224_));
AND2X2 AND2X2_516 ( .A(u1__abc_51895_new_n392_), .B(u1_xinf), .Y(aNan));
AND2X2 AND2X2_5160 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_225_), .Y(u2__abc_52155_new_n12048_));
AND2X2 AND2X2_5161 ( .A(u2__abc_52155_new_n12035_), .B(u2__abc_52155_new_n4503_), .Y(u2__abc_52155_new_n12049_));
AND2X2 AND2X2_5162 ( .A(u2__abc_52155_new_n12049_), .B(u2__abc_52155_new_n4500_), .Y(u2__abc_52155_new_n12050_));
AND2X2 AND2X2_5163 ( .A(u2__abc_52155_new_n12052_), .B(u2__abc_52155_new_n12051_), .Y(u2__abc_52155_new_n12053_));
AND2X2 AND2X2_5164 ( .A(u2__abc_52155_new_n12054_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12055_));
AND2X2 AND2X2_5165 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_223_), .Y(u2__abc_52155_new_n12056_));
AND2X2 AND2X2_5166 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4489_), .Y(u2__abc_52155_new_n12059_));
AND2X2 AND2X2_5167 ( .A(u2__abc_52155_new_n12060_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12061_));
AND2X2 AND2X2_5168 ( .A(u2__abc_52155_new_n12058_), .B(u2__abc_52155_new_n12061_), .Y(u2__abc_52155_new_n12062_));
AND2X2 AND2X2_5169 ( .A(u2__abc_52155_new_n12063_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__225_));
AND2X2 AND2X2_517 ( .A(ld), .B(u2_state_0_), .Y(u2__abc_52155_new_n2963_));
AND2X2 AND2X2_5170 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_226_), .Y(u2__abc_52155_new_n12065_));
AND2X2 AND2X2_5171 ( .A(u2__abc_52155_new_n4496_), .B(u2__abc_52155_new_n4503_), .Y(u2__abc_52155_new_n12066_));
AND2X2 AND2X2_5172 ( .A(u2__abc_52155_new_n12035_), .B(u2__abc_52155_new_n12066_), .Y(u2__abc_52155_new_n12067_));
AND2X2 AND2X2_5173 ( .A(u2__abc_52155_new_n12069_), .B(u2__abc_52155_new_n4485_), .Y(u2__abc_52155_new_n12070_));
AND2X2 AND2X2_5174 ( .A(u2__abc_52155_new_n12072_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12073_));
AND2X2 AND2X2_5175 ( .A(u2__abc_52155_new_n12073_), .B(u2__abc_52155_new_n12071_), .Y(u2__abc_52155_new_n12074_));
AND2X2 AND2X2_5176 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_224_), .Y(u2__abc_52155_new_n12075_));
AND2X2 AND2X2_5177 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4535_), .Y(u2__abc_52155_new_n12078_));
AND2X2 AND2X2_5178 ( .A(u2__abc_52155_new_n12079_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12080_));
AND2X2 AND2X2_5179 ( .A(u2__abc_52155_new_n12077_), .B(u2__abc_52155_new_n12080_), .Y(u2__abc_52155_new_n12081_));
AND2X2 AND2X2_518 ( .A(u2__abc_52155_new_n2963_), .B(ce), .Y(u2__abc_52155_new_n2964_));
AND2X2 AND2X2_5180 ( .A(u2__abc_52155_new_n12082_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__226_));
AND2X2 AND2X2_5181 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_227_), .Y(u2__abc_52155_new_n12084_));
AND2X2 AND2X2_5182 ( .A(u2__abc_52155_new_n12071_), .B(u2__abc_52155_new_n4481_), .Y(u2__abc_52155_new_n12085_));
AND2X2 AND2X2_5183 ( .A(u2__abc_52155_new_n12085_), .B(u2__abc_52155_new_n4492_), .Y(u2__abc_52155_new_n12086_));
AND2X2 AND2X2_5184 ( .A(u2__abc_52155_new_n12088_), .B(u2__abc_52155_new_n12087_), .Y(u2__abc_52155_new_n12089_));
AND2X2 AND2X2_5185 ( .A(u2__abc_52155_new_n12090_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12091_));
AND2X2 AND2X2_5186 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_225_), .Y(u2__abc_52155_new_n12092_));
AND2X2 AND2X2_5187 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4528_), .Y(u2__abc_52155_new_n12095_));
AND2X2 AND2X2_5188 ( .A(u2__abc_52155_new_n12096_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12097_));
AND2X2 AND2X2_5189 ( .A(u2__abc_52155_new_n12094_), .B(u2__abc_52155_new_n12097_), .Y(u2__abc_52155_new_n12098_));
AND2X2 AND2X2_519 ( .A(u2__abc_52155_new_n2965_), .B(u2_cnt_7_), .Y(u2__abc_52155_new_n2966_));
AND2X2 AND2X2_5190 ( .A(u2__abc_52155_new_n12099_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__227_));
AND2X2 AND2X2_5191 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_228_), .Y(u2__abc_52155_new_n12101_));
AND2X2 AND2X2_5192 ( .A(u2__abc_52155_new_n4481_), .B(u2__abc_52155_new_n4488_), .Y(u2__abc_52155_new_n12102_));
AND2X2 AND2X2_5193 ( .A(u2__abc_52155_new_n12105_), .B(u2__abc_52155_new_n4493_), .Y(u2__abc_52155_new_n12106_));
AND2X2 AND2X2_5194 ( .A(u2__abc_52155_new_n12107_), .B(u2__abc_52155_new_n12103_), .Y(u2__abc_52155_new_n12108_));
AND2X2 AND2X2_5195 ( .A(u2__abc_52155_new_n12033_), .B(u2__abc_52155_new_n4509_), .Y(u2__abc_52155_new_n12110_));
AND2X2 AND2X2_5196 ( .A(u2__abc_52155_new_n12111_), .B(u2__abc_52155_new_n4538_), .Y(u2__abc_52155_new_n12112_));
AND2X2 AND2X2_5197 ( .A(u2__abc_52155_new_n12114_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12115_));
AND2X2 AND2X2_5198 ( .A(u2__abc_52155_new_n12115_), .B(u2__abc_52155_new_n12113_), .Y(u2__abc_52155_new_n12116_));
AND2X2 AND2X2_5199 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_226_), .Y(u2__abc_52155_new_n12117_));
AND2X2 AND2X2_52 ( .A(_abc_73687_new_n753_), .B(sqrto_51_), .Y(\o[87] ));
AND2X2 AND2X2_520 ( .A(u2_cnt_5_), .B(u2_cnt_6_), .Y(u2__abc_52155_new_n2967_));
AND2X2 AND2X2_5200 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4513_), .Y(u2__abc_52155_new_n12120_));
AND2X2 AND2X2_5201 ( .A(u2__abc_52155_new_n12121_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12122_));
AND2X2 AND2X2_5202 ( .A(u2__abc_52155_new_n12119_), .B(u2__abc_52155_new_n12122_), .Y(u2__abc_52155_new_n12123_));
AND2X2 AND2X2_5203 ( .A(u2__abc_52155_new_n12124_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__228_));
AND2X2 AND2X2_5204 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_229_), .Y(u2__abc_52155_new_n12126_));
AND2X2 AND2X2_5205 ( .A(u2__abc_52155_new_n12113_), .B(u2__abc_52155_new_n4534_), .Y(u2__abc_52155_new_n12127_));
AND2X2 AND2X2_5206 ( .A(u2__abc_52155_new_n12127_), .B(u2__abc_52155_new_n4531_), .Y(u2__abc_52155_new_n12128_));
AND2X2 AND2X2_5207 ( .A(u2__abc_52155_new_n12130_), .B(u2__abc_52155_new_n12129_), .Y(u2__abc_52155_new_n12131_));
AND2X2 AND2X2_5208 ( .A(u2__abc_52155_new_n12132_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12133_));
AND2X2 AND2X2_5209 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_227_), .Y(u2__abc_52155_new_n12134_));
AND2X2 AND2X2_521 ( .A(u2__abc_52155_new_n2966_), .B(u2__abc_52155_new_n2967_), .Y(u2__abc_52155_new_n2968_));
AND2X2 AND2X2_5210 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4520_), .Y(u2__abc_52155_new_n12137_));
AND2X2 AND2X2_5211 ( .A(u2__abc_52155_new_n12138_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12139_));
AND2X2 AND2X2_5212 ( .A(u2__abc_52155_new_n12136_), .B(u2__abc_52155_new_n12139_), .Y(u2__abc_52155_new_n12140_));
AND2X2 AND2X2_5213 ( .A(u2__abc_52155_new_n12141_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__229_));
AND2X2 AND2X2_5214 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_230_), .Y(u2__abc_52155_new_n12143_));
AND2X2 AND2X2_5215 ( .A(u2__abc_52155_new_n4527_), .B(u2__abc_52155_new_n4534_), .Y(u2__abc_52155_new_n12144_));
AND2X2 AND2X2_5216 ( .A(u2__abc_52155_new_n12113_), .B(u2__abc_52155_new_n12144_), .Y(u2__abc_52155_new_n12145_));
AND2X2 AND2X2_5217 ( .A(u2__abc_52155_new_n12147_), .B(u2__abc_52155_new_n4516_), .Y(u2__abc_52155_new_n12148_));
AND2X2 AND2X2_5218 ( .A(u2__abc_52155_new_n12150_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12151_));
AND2X2 AND2X2_5219 ( .A(u2__abc_52155_new_n12151_), .B(u2__abc_52155_new_n12149_), .Y(u2__abc_52155_new_n12152_));
AND2X2 AND2X2_522 ( .A(u2__abc_52155_new_n2971_), .B(u2_cnt_1_), .Y(u2__abc_52155_new_n2972_));
AND2X2 AND2X2_5220 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_228_), .Y(u2__abc_52155_new_n12153_));
AND2X2 AND2X2_5221 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4472_), .Y(u2__abc_52155_new_n12156_));
AND2X2 AND2X2_5222 ( .A(u2__abc_52155_new_n12157_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12158_));
AND2X2 AND2X2_5223 ( .A(u2__abc_52155_new_n12155_), .B(u2__abc_52155_new_n12158_), .Y(u2__abc_52155_new_n12159_));
AND2X2 AND2X2_5224 ( .A(u2__abc_52155_new_n12160_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__230_));
AND2X2 AND2X2_5225 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_231_), .Y(u2__abc_52155_new_n12162_));
AND2X2 AND2X2_5226 ( .A(u2__abc_52155_new_n12149_), .B(u2__abc_52155_new_n4512_), .Y(u2__abc_52155_new_n12163_));
AND2X2 AND2X2_5227 ( .A(u2__abc_52155_new_n12163_), .B(u2__abc_52155_new_n4523_), .Y(u2__abc_52155_new_n12164_));
AND2X2 AND2X2_5228 ( .A(u2__abc_52155_new_n12166_), .B(u2__abc_52155_new_n12165_), .Y(u2__abc_52155_new_n12167_));
AND2X2 AND2X2_5229 ( .A(u2__abc_52155_new_n12168_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12169_));
AND2X2 AND2X2_523 ( .A(u2__abc_52155_new_n2970_), .B(u2__abc_52155_new_n2972_), .Y(u2__abc_52155_new_n2973_));
AND2X2 AND2X2_5230 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_229_), .Y(u2__abc_52155_new_n12170_));
AND2X2 AND2X2_5231 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4465_), .Y(u2__abc_52155_new_n12173_));
AND2X2 AND2X2_5232 ( .A(u2__abc_52155_new_n12174_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12175_));
AND2X2 AND2X2_5233 ( .A(u2__abc_52155_new_n12172_), .B(u2__abc_52155_new_n12175_), .Y(u2__abc_52155_new_n12176_));
AND2X2 AND2X2_5234 ( .A(u2__abc_52155_new_n12177_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__231_));
AND2X2 AND2X2_5235 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_232_), .Y(u2__abc_52155_new_n12179_));
AND2X2 AND2X2_5236 ( .A(u2__abc_52155_new_n12109_), .B(u2__abc_52155_new_n4540_), .Y(u2__abc_52155_new_n12180_));
AND2X2 AND2X2_5237 ( .A(u2__abc_52155_new_n12182_), .B(u2__abc_52155_new_n4524_), .Y(u2__abc_52155_new_n12183_));
AND2X2 AND2X2_5238 ( .A(u2__abc_52155_new_n4522_), .B(u2__abc_52155_new_n4511_), .Y(u2__abc_52155_new_n12184_));
AND2X2 AND2X2_5239 ( .A(u2__abc_52155_new_n12033_), .B(u2__abc_52155_new_n4541_), .Y(u2__abc_52155_new_n12188_));
AND2X2 AND2X2_524 ( .A(u2__abc_52155_new_n2973_), .B(u2__abc_52155_new_n2968_), .Y(u2__abc_52155_new_n2974_));
AND2X2 AND2X2_5240 ( .A(u2__abc_52155_new_n12189_), .B(u2__abc_52155_new_n4475_), .Y(u2__abc_52155_new_n12190_));
AND2X2 AND2X2_5241 ( .A(u2__abc_52155_new_n12192_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12193_));
AND2X2 AND2X2_5242 ( .A(u2__abc_52155_new_n12193_), .B(u2__abc_52155_new_n12191_), .Y(u2__abc_52155_new_n12194_));
AND2X2 AND2X2_5243 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_230_), .Y(u2__abc_52155_new_n12195_));
AND2X2 AND2X2_5244 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4450_), .Y(u2__abc_52155_new_n12198_));
AND2X2 AND2X2_5245 ( .A(u2__abc_52155_new_n12199_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12200_));
AND2X2 AND2X2_5246 ( .A(u2__abc_52155_new_n12197_), .B(u2__abc_52155_new_n12200_), .Y(u2__abc_52155_new_n12201_));
AND2X2 AND2X2_5247 ( .A(u2__abc_52155_new_n12202_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__232_));
AND2X2 AND2X2_5248 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_233_), .Y(u2__abc_52155_new_n12204_));
AND2X2 AND2X2_5249 ( .A(u2__abc_52155_new_n12191_), .B(u2__abc_52155_new_n4471_), .Y(u2__abc_52155_new_n12206_));
AND2X2 AND2X2_525 ( .A(u2__abc_52155_new_n2974_), .B(ce), .Y(u2__abc_52155_new_n2975_));
AND2X2 AND2X2_5250 ( .A(u2__abc_52155_new_n12207_), .B(u2__abc_52155_new_n12205_), .Y(u2__abc_52155_new_n12208_));
AND2X2 AND2X2_5251 ( .A(u2__abc_52155_new_n12206_), .B(u2__abc_52155_new_n4468_), .Y(u2__abc_52155_new_n12209_));
AND2X2 AND2X2_5252 ( .A(u2__abc_52155_new_n12210_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12211_));
AND2X2 AND2X2_5253 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_231_), .Y(u2__abc_52155_new_n12212_));
AND2X2 AND2X2_5254 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4457_), .Y(u2__abc_52155_new_n12215_));
AND2X2 AND2X2_5255 ( .A(u2__abc_52155_new_n12216_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12217_));
AND2X2 AND2X2_5256 ( .A(u2__abc_52155_new_n12214_), .B(u2__abc_52155_new_n12217_), .Y(u2__abc_52155_new_n12218_));
AND2X2 AND2X2_5257 ( .A(u2__abc_52155_new_n12219_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__233_));
AND2X2 AND2X2_5258 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_234_), .Y(u2__abc_52155_new_n12221_));
AND2X2 AND2X2_5259 ( .A(u2__abc_52155_new_n4464_), .B(u2__abc_52155_new_n4471_), .Y(u2__abc_52155_new_n12222_));
AND2X2 AND2X2_526 ( .A(u2__abc_52155_new_n2976_), .B(u2_state_2_), .Y(u2__abc_52155_new_n2977_));
AND2X2 AND2X2_5260 ( .A(u2__abc_52155_new_n12189_), .B(u2__abc_52155_new_n4476_), .Y(u2__abc_52155_new_n12225_));
AND2X2 AND2X2_5261 ( .A(u2__abc_52155_new_n12226_), .B(u2__abc_52155_new_n4453_), .Y(u2__abc_52155_new_n12227_));
AND2X2 AND2X2_5262 ( .A(u2__abc_52155_new_n12229_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12230_));
AND2X2 AND2X2_5263 ( .A(u2__abc_52155_new_n12230_), .B(u2__abc_52155_new_n12228_), .Y(u2__abc_52155_new_n12231_));
AND2X2 AND2X2_5264 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_232_), .Y(u2__abc_52155_new_n12232_));
AND2X2 AND2X2_5265 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4441_), .Y(u2__abc_52155_new_n12235_));
AND2X2 AND2X2_5266 ( .A(u2__abc_52155_new_n12236_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12237_));
AND2X2 AND2X2_5267 ( .A(u2__abc_52155_new_n12234_), .B(u2__abc_52155_new_n12237_), .Y(u2__abc_52155_new_n12238_));
AND2X2 AND2X2_5268 ( .A(u2__abc_52155_new_n12239_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__234_));
AND2X2 AND2X2_5269 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_235_), .Y(u2__abc_52155_new_n12241_));
AND2X2 AND2X2_527 ( .A(u2__abc_52155_new_n2978_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_2_));
AND2X2 AND2X2_5270 ( .A(u2__abc_52155_new_n12228_), .B(u2__abc_52155_new_n4449_), .Y(u2__abc_52155_new_n12242_));
AND2X2 AND2X2_5271 ( .A(u2__abc_52155_new_n12242_), .B(u2__abc_52155_new_n4460_), .Y(u2__abc_52155_new_n12243_));
AND2X2 AND2X2_5272 ( .A(u2__abc_52155_new_n12245_), .B(u2__abc_52155_new_n12244_), .Y(u2__abc_52155_new_n12246_));
AND2X2 AND2X2_5273 ( .A(u2__abc_52155_new_n12247_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12248_));
AND2X2 AND2X2_5274 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_233_), .Y(u2__abc_52155_new_n12249_));
AND2X2 AND2X2_5275 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4434_), .Y(u2__abc_52155_new_n12252_));
AND2X2 AND2X2_5276 ( .A(u2__abc_52155_new_n12253_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12254_));
AND2X2 AND2X2_5277 ( .A(u2__abc_52155_new_n12251_), .B(u2__abc_52155_new_n12254_), .Y(u2__abc_52155_new_n12255_));
AND2X2 AND2X2_5278 ( .A(u2__abc_52155_new_n12256_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__235_));
AND2X2 AND2X2_5279 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_236_), .Y(u2__abc_52155_new_n12258_));
AND2X2 AND2X2_528 ( .A(u2__abc_52155_new_n2962_), .B(ce), .Y(u2__abc_52155_new_n2982_));
AND2X2 AND2X2_5280 ( .A(u2__abc_52155_new_n4449_), .B(u2__abc_52155_new_n4456_), .Y(u2__abc_52155_new_n12259_));
AND2X2 AND2X2_5281 ( .A(u2__abc_52155_new_n12228_), .B(u2__abc_52155_new_n12259_), .Y(u2__abc_52155_new_n12260_));
AND2X2 AND2X2_5282 ( .A(u2__abc_52155_new_n12262_), .B(u2__abc_52155_new_n4444_), .Y(u2__abc_52155_new_n12263_));
AND2X2 AND2X2_5283 ( .A(u2__abc_52155_new_n12265_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12266_));
AND2X2 AND2X2_5284 ( .A(u2__abc_52155_new_n12266_), .B(u2__abc_52155_new_n12264_), .Y(u2__abc_52155_new_n12267_));
AND2X2 AND2X2_5285 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_234_), .Y(u2__abc_52155_new_n12268_));
AND2X2 AND2X2_5286 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4419_), .Y(u2__abc_52155_new_n12271_));
AND2X2 AND2X2_5287 ( .A(u2__abc_52155_new_n12272_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12273_));
AND2X2 AND2X2_5288 ( .A(u2__abc_52155_new_n12270_), .B(u2__abc_52155_new_n12273_), .Y(u2__abc_52155_new_n12274_));
AND2X2 AND2X2_5289 ( .A(u2__abc_52155_new_n12275_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__236_));
AND2X2 AND2X2_529 ( .A(u2__abc_52155_new_n2984_), .B(u2_state_0_), .Y(u2__abc_52155_new_n2985_));
AND2X2 AND2X2_5290 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_237_), .Y(u2__abc_52155_new_n12277_));
AND2X2 AND2X2_5291 ( .A(u2__abc_52155_new_n12264_), .B(u2__abc_52155_new_n4440_), .Y(u2__abc_52155_new_n12278_));
AND2X2 AND2X2_5292 ( .A(u2__abc_52155_new_n12278_), .B(u2__abc_52155_new_n4437_), .Y(u2__abc_52155_new_n12279_));
AND2X2 AND2X2_5293 ( .A(u2__abc_52155_new_n12281_), .B(u2__abc_52155_new_n12280_), .Y(u2__abc_52155_new_n12282_));
AND2X2 AND2X2_5294 ( .A(u2__abc_52155_new_n12283_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12284_));
AND2X2 AND2X2_5295 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_235_), .Y(u2__abc_52155_new_n12285_));
AND2X2 AND2X2_5296 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4426_), .Y(u2__abc_52155_new_n12288_));
AND2X2 AND2X2_5297 ( .A(u2__abc_52155_new_n12289_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12290_));
AND2X2 AND2X2_5298 ( .A(u2__abc_52155_new_n12287_), .B(u2__abc_52155_new_n12290_), .Y(u2__abc_52155_new_n12291_));
AND2X2 AND2X2_5299 ( .A(u2__abc_52155_new_n12292_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__237_));
AND2X2 AND2X2_53 ( .A(_abc_73687_new_n753_), .B(sqrto_52_), .Y(\o[88] ));
AND2X2 AND2X2_530 ( .A(u2__abc_52155_new_n2987_), .B(u2__abc_52155_new_n2981_), .Y(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_0_));
AND2X2 AND2X2_5300 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_238_), .Y(u2__abc_52155_new_n12294_));
AND2X2 AND2X2_5301 ( .A(u2__abc_52155_new_n4433_), .B(u2__abc_52155_new_n4440_), .Y(u2__abc_52155_new_n12295_));
AND2X2 AND2X2_5302 ( .A(u2__abc_52155_new_n12264_), .B(u2__abc_52155_new_n12295_), .Y(u2__abc_52155_new_n12296_));
AND2X2 AND2X2_5303 ( .A(u2__abc_52155_new_n12298_), .B(u2__abc_52155_new_n4422_), .Y(u2__abc_52155_new_n12299_));
AND2X2 AND2X2_5304 ( .A(u2__abc_52155_new_n12301_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12302_));
AND2X2 AND2X2_5305 ( .A(u2__abc_52155_new_n12302_), .B(u2__abc_52155_new_n12300_), .Y(u2__abc_52155_new_n12303_));
AND2X2 AND2X2_5306 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_236_), .Y(u2__abc_52155_new_n12304_));
AND2X2 AND2X2_5307 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4355_), .Y(u2__abc_52155_new_n12307_));
AND2X2 AND2X2_5308 ( .A(u2__abc_52155_new_n12308_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12309_));
AND2X2 AND2X2_5309 ( .A(u2__abc_52155_new_n12306_), .B(u2__abc_52155_new_n12309_), .Y(u2__abc_52155_new_n12310_));
AND2X2 AND2X2_531 ( .A(u2__abc_52155_new_n2989_), .B(done), .Y(u2__abc_52155_new_n2990_));
AND2X2 AND2X2_5310 ( .A(u2__abc_52155_new_n12311_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__238_));
AND2X2 AND2X2_5311 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_239_), .Y(u2__abc_52155_new_n12313_));
AND2X2 AND2X2_5312 ( .A(u2__abc_52155_new_n12300_), .B(u2__abc_52155_new_n4418_), .Y(u2__abc_52155_new_n12314_));
AND2X2 AND2X2_5313 ( .A(u2__abc_52155_new_n12314_), .B(u2__abc_52155_new_n4429_), .Y(u2__abc_52155_new_n12315_));
AND2X2 AND2X2_5314 ( .A(u2__abc_52155_new_n12317_), .B(u2__abc_52155_new_n12316_), .Y(u2__abc_52155_new_n12318_));
AND2X2 AND2X2_5315 ( .A(u2__abc_52155_new_n12319_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12320_));
AND2X2 AND2X2_5316 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_237_), .Y(u2__abc_52155_new_n12321_));
AND2X2 AND2X2_5317 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4362_), .Y(u2__abc_52155_new_n12324_));
AND2X2 AND2X2_5318 ( .A(u2__abc_52155_new_n12325_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12326_));
AND2X2 AND2X2_5319 ( .A(u2__abc_52155_new_n12323_), .B(u2__abc_52155_new_n12326_), .Y(u2__abc_52155_new_n12327_));
AND2X2 AND2X2_532 ( .A(u2__abc_52155_new_n2970_), .B(u2__abc_52155_new_n2966_), .Y(u2__abc_52155_new_n2991_));
AND2X2 AND2X2_5320 ( .A(u2__abc_52155_new_n12328_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__239_));
AND2X2 AND2X2_5321 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_240_), .Y(u2__abc_52155_new_n12330_));
AND2X2 AND2X2_5322 ( .A(u2__abc_52155_new_n12187_), .B(u2__abc_52155_new_n4478_), .Y(u2__abc_52155_new_n12331_));
AND2X2 AND2X2_5323 ( .A(u2__abc_52155_new_n12224_), .B(u2__abc_52155_new_n4461_), .Y(u2__abc_52155_new_n12334_));
AND2X2 AND2X2_5324 ( .A(u2__abc_52155_new_n12335_), .B(u2__abc_52155_new_n12333_), .Y(u2__abc_52155_new_n12336_));
AND2X2 AND2X2_5325 ( .A(u2__abc_52155_new_n12337_), .B(u2__abc_52155_new_n4446_), .Y(u2__abc_52155_new_n12338_));
AND2X2 AND2X2_5326 ( .A(u2__abc_52155_new_n4418_), .B(u2__abc_52155_new_n4425_), .Y(u2__abc_52155_new_n12340_));
AND2X2 AND2X2_5327 ( .A(u2__abc_52155_new_n12343_), .B(u2__abc_52155_new_n4430_), .Y(u2__abc_52155_new_n12344_));
AND2X2 AND2X2_5328 ( .A(u2__abc_52155_new_n12345_), .B(u2__abc_52155_new_n12341_), .Y(u2__abc_52155_new_n12346_));
AND2X2 AND2X2_5329 ( .A(u2__abc_52155_new_n12339_), .B(u2__abc_52155_new_n12346_), .Y(u2__abc_52155_new_n12347_));
AND2X2 AND2X2_533 ( .A(u2__abc_52155_new_n2972_), .B(u2__abc_52155_new_n2967_), .Y(u2__abc_52155_new_n2992_));
AND2X2 AND2X2_5330 ( .A(u2__abc_52155_new_n12332_), .B(u2__abc_52155_new_n12347_), .Y(u2__abc_52155_new_n12348_));
AND2X2 AND2X2_5331 ( .A(u2__abc_52155_new_n12033_), .B(u2__abc_52155_new_n4542_), .Y(u2__abc_52155_new_n12350_));
AND2X2 AND2X2_5332 ( .A(u2__abc_52155_new_n12351_), .B(u2__abc_52155_new_n4358_), .Y(u2__abc_52155_new_n12352_));
AND2X2 AND2X2_5333 ( .A(u2__abc_52155_new_n12354_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12355_));
AND2X2 AND2X2_5334 ( .A(u2__abc_52155_new_n12355_), .B(u2__abc_52155_new_n12353_), .Y(u2__abc_52155_new_n12356_));
AND2X2 AND2X2_5335 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_238_), .Y(u2__abc_52155_new_n12357_));
AND2X2 AND2X2_5336 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4370_), .Y(u2__abc_52155_new_n12360_));
AND2X2 AND2X2_5337 ( .A(u2__abc_52155_new_n12361_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12362_));
AND2X2 AND2X2_5338 ( .A(u2__abc_52155_new_n12359_), .B(u2__abc_52155_new_n12362_), .Y(u2__abc_52155_new_n12363_));
AND2X2 AND2X2_5339 ( .A(u2__abc_52155_new_n12364_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__240_));
AND2X2 AND2X2_534 ( .A(u2__abc_52155_new_n2991_), .B(u2__abc_52155_new_n2992_), .Y(u2__abc_52155_new_n2993_));
AND2X2 AND2X2_5340 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_241_), .Y(u2__abc_52155_new_n12366_));
AND2X2 AND2X2_5341 ( .A(u2__abc_52155_new_n12353_), .B(u2__abc_52155_new_n4354_), .Y(u2__abc_52155_new_n12367_));
AND2X2 AND2X2_5342 ( .A(u2__abc_52155_new_n12367_), .B(u2__abc_52155_new_n4365_), .Y(u2__abc_52155_new_n12368_));
AND2X2 AND2X2_5343 ( .A(u2__abc_52155_new_n12370_), .B(u2__abc_52155_new_n12369_), .Y(u2__abc_52155_new_n12371_));
AND2X2 AND2X2_5344 ( .A(u2__abc_52155_new_n12372_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12373_));
AND2X2 AND2X2_5345 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_239_), .Y(u2__abc_52155_new_n12374_));
AND2X2 AND2X2_5346 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4377_), .Y(u2__abc_52155_new_n12377_));
AND2X2 AND2X2_5347 ( .A(u2__abc_52155_new_n12378_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12379_));
AND2X2 AND2X2_5348 ( .A(u2__abc_52155_new_n12376_), .B(u2__abc_52155_new_n12379_), .Y(u2__abc_52155_new_n12380_));
AND2X2 AND2X2_5349 ( .A(u2__abc_52155_new_n12381_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__241_));
AND2X2 AND2X2_535 ( .A(u2__abc_52155_new_n2993_), .B(u2_state_2_), .Y(u2__abc_52155_new_n2994_));
AND2X2 AND2X2_5350 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_242_), .Y(u2__abc_52155_new_n12383_));
AND2X2 AND2X2_5351 ( .A(u2__abc_52155_new_n12384_), .B(u2__abc_52155_new_n4361_), .Y(u2__abc_52155_new_n12385_));
AND2X2 AND2X2_5352 ( .A(u2__abc_52155_new_n12351_), .B(u2__abc_52155_new_n4366_), .Y(u2__abc_52155_new_n12387_));
AND2X2 AND2X2_5353 ( .A(u2__abc_52155_new_n12388_), .B(u2__abc_52155_new_n4373_), .Y(u2__abc_52155_new_n12389_));
AND2X2 AND2X2_5354 ( .A(u2__abc_52155_new_n12391_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12392_));
AND2X2 AND2X2_5355 ( .A(u2__abc_52155_new_n12392_), .B(u2__abc_52155_new_n12390_), .Y(u2__abc_52155_new_n12393_));
AND2X2 AND2X2_5356 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_240_), .Y(u2__abc_52155_new_n12394_));
AND2X2 AND2X2_5357 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4408_), .Y(u2__abc_52155_new_n12397_));
AND2X2 AND2X2_5358 ( .A(u2__abc_52155_new_n12398_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12399_));
AND2X2 AND2X2_5359 ( .A(u2__abc_52155_new_n12396_), .B(u2__abc_52155_new_n12399_), .Y(u2__abc_52155_new_n12400_));
AND2X2 AND2X2_536 ( .A(u2__abc_52155_new_n2994_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n2995_));
AND2X2 AND2X2_5360 ( .A(u2__abc_52155_new_n12401_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__242_));
AND2X2 AND2X2_5361 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_243_), .Y(u2__abc_52155_new_n12403_));
AND2X2 AND2X2_5362 ( .A(u2__abc_52155_new_n12390_), .B(u2__abc_52155_new_n4369_), .Y(u2__abc_52155_new_n12404_));
AND2X2 AND2X2_5363 ( .A(u2__abc_52155_new_n12404_), .B(u2__abc_52155_new_n4380_), .Y(u2__abc_52155_new_n12405_));
AND2X2 AND2X2_5364 ( .A(u2__abc_52155_new_n12407_), .B(u2__abc_52155_new_n12406_), .Y(u2__abc_52155_new_n12408_));
AND2X2 AND2X2_5365 ( .A(u2__abc_52155_new_n12409_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12410_));
AND2X2 AND2X2_5366 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_241_), .Y(u2__abc_52155_new_n12411_));
AND2X2 AND2X2_5367 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4401_), .Y(u2__abc_52155_new_n12414_));
AND2X2 AND2X2_5368 ( .A(u2__abc_52155_new_n12415_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12416_));
AND2X2 AND2X2_5369 ( .A(u2__abc_52155_new_n12413_), .B(u2__abc_52155_new_n12416_), .Y(u2__abc_52155_new_n12417_));
AND2X2 AND2X2_537 ( .A(ce), .B(u2_state_0_), .Y(u2__abc_52155_new_n2997_));
AND2X2 AND2X2_5370 ( .A(u2__abc_52155_new_n12418_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__243_));
AND2X2 AND2X2_5371 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_244_), .Y(u2__abc_52155_new_n12420_));
AND2X2 AND2X2_5372 ( .A(u2__abc_52155_new_n12386_), .B(u2__abc_52155_new_n4381_), .Y(u2__abc_52155_new_n12421_));
AND2X2 AND2X2_5373 ( .A(u2__abc_52155_new_n4379_), .B(u2__abc_52155_new_n4368_), .Y(u2__abc_52155_new_n12422_));
AND2X2 AND2X2_5374 ( .A(u2__abc_52155_new_n12351_), .B(u2__abc_52155_new_n4382_), .Y(u2__abc_52155_new_n12425_));
AND2X2 AND2X2_5375 ( .A(u2__abc_52155_new_n12426_), .B(u2__abc_52155_new_n4411_), .Y(u2__abc_52155_new_n12427_));
AND2X2 AND2X2_5376 ( .A(u2__abc_52155_new_n12429_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12430_));
AND2X2 AND2X2_5377 ( .A(u2__abc_52155_new_n12430_), .B(u2__abc_52155_new_n12428_), .Y(u2__abc_52155_new_n12431_));
AND2X2 AND2X2_5378 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_242_), .Y(u2__abc_52155_new_n12432_));
AND2X2 AND2X2_5379 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4386_), .Y(u2__abc_52155_new_n12435_));
AND2X2 AND2X2_538 ( .A(u2_state_2_), .B(ce), .Y(u2__abc_52155_new_n2999_));
AND2X2 AND2X2_5380 ( .A(u2__abc_52155_new_n12436_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12437_));
AND2X2 AND2X2_5381 ( .A(u2__abc_52155_new_n12434_), .B(u2__abc_52155_new_n12437_), .Y(u2__abc_52155_new_n12438_));
AND2X2 AND2X2_5382 ( .A(u2__abc_52155_new_n12439_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__244_));
AND2X2 AND2X2_5383 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_245_), .Y(u2__abc_52155_new_n12441_));
AND2X2 AND2X2_5384 ( .A(u2__abc_52155_new_n12428_), .B(u2__abc_52155_new_n4407_), .Y(u2__abc_52155_new_n12442_));
AND2X2 AND2X2_5385 ( .A(u2__abc_52155_new_n12443_), .B(u2__abc_52155_new_n4404_), .Y(u2__abc_52155_new_n12444_));
AND2X2 AND2X2_5386 ( .A(u2__abc_52155_new_n12446_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12447_));
AND2X2 AND2X2_5387 ( .A(u2__abc_52155_new_n12447_), .B(u2__abc_52155_new_n12445_), .Y(u2__abc_52155_new_n12448_));
AND2X2 AND2X2_5388 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_243_), .Y(u2__abc_52155_new_n12449_));
AND2X2 AND2X2_5389 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4393_), .Y(u2__abc_52155_new_n12452_));
AND2X2 AND2X2_539 ( .A(u2__abc_52155_new_n2998_), .B(u2__abc_52155_new_n3000_), .Y(u2__abc_52155_new_n3001_));
AND2X2 AND2X2_5390 ( .A(u2__abc_52155_new_n12453_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12454_));
AND2X2 AND2X2_5391 ( .A(u2__abc_52155_new_n12451_), .B(u2__abc_52155_new_n12454_), .Y(u2__abc_52155_new_n12455_));
AND2X2 AND2X2_5392 ( .A(u2__abc_52155_new_n12456_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__245_));
AND2X2 AND2X2_5393 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_246_), .Y(u2__abc_52155_new_n12458_));
AND2X2 AND2X2_5394 ( .A(u2__abc_52155_new_n12445_), .B(u2__abc_52155_new_n4400_), .Y(u2__abc_52155_new_n12459_));
AND2X2 AND2X2_5395 ( .A(u2__abc_52155_new_n12460_), .B(u2__abc_52155_new_n4389_), .Y(u2__abc_52155_new_n12461_));
AND2X2 AND2X2_5396 ( .A(u2__abc_52155_new_n12463_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12464_));
AND2X2 AND2X2_5397 ( .A(u2__abc_52155_new_n12464_), .B(u2__abc_52155_new_n12462_), .Y(u2__abc_52155_new_n12465_));
AND2X2 AND2X2_5398 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_244_), .Y(u2__abc_52155_new_n12466_));
AND2X2 AND2X2_5399 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4292_), .Y(u2__abc_52155_new_n12469_));
AND2X2 AND2X2_54 ( .A(_abc_73687_new_n753_), .B(sqrto_53_), .Y(\o[89] ));
AND2X2 AND2X2_540 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_0_), .Y(u2__abc_52155_new_n3003_));
AND2X2 AND2X2_5400 ( .A(u2__abc_52155_new_n12470_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12471_));
AND2X2 AND2X2_5401 ( .A(u2__abc_52155_new_n12468_), .B(u2__abc_52155_new_n12471_), .Y(u2__abc_52155_new_n12472_));
AND2X2 AND2X2_5402 ( .A(u2__abc_52155_new_n12473_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__246_));
AND2X2 AND2X2_5403 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_247_), .Y(u2__abc_52155_new_n12475_));
AND2X2 AND2X2_5404 ( .A(u2__abc_52155_new_n12462_), .B(u2__abc_52155_new_n4385_), .Y(u2__abc_52155_new_n12476_));
AND2X2 AND2X2_5405 ( .A(u2__abc_52155_new_n12476_), .B(u2__abc_52155_new_n4396_), .Y(u2__abc_52155_new_n12477_));
AND2X2 AND2X2_5406 ( .A(u2__abc_52155_new_n12479_), .B(u2__abc_52155_new_n12478_), .Y(u2__abc_52155_new_n12480_));
AND2X2 AND2X2_5407 ( .A(u2__abc_52155_new_n12481_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12482_));
AND2X2 AND2X2_5408 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_245_), .Y(u2__abc_52155_new_n12483_));
AND2X2 AND2X2_5409 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4299_), .Y(u2__abc_52155_new_n12486_));
AND2X2 AND2X2_541 ( .A(u2__abc_52155_new_n3004_), .B(u2_o_449_), .Y(u2__abc_52155_new_n3005_));
AND2X2 AND2X2_5410 ( .A(u2__abc_52155_new_n12487_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12488_));
AND2X2 AND2X2_5411 ( .A(u2__abc_52155_new_n12485_), .B(u2__abc_52155_new_n12488_), .Y(u2__abc_52155_new_n12489_));
AND2X2 AND2X2_5412 ( .A(u2__abc_52155_new_n12490_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__247_));
AND2X2 AND2X2_5413 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_248_), .Y(u2__abc_52155_new_n12492_));
AND2X2 AND2X2_5414 ( .A(u2__abc_52155_new_n12424_), .B(u2__abc_52155_new_n4413_), .Y(u2__abc_52155_new_n12493_));
AND2X2 AND2X2_5415 ( .A(u2__abc_52155_new_n12494_), .B(u2__abc_52155_new_n4403_), .Y(u2__abc_52155_new_n12495_));
AND2X2 AND2X2_5416 ( .A(u2__abc_52155_new_n4397_), .B(u2__abc_52155_new_n12495_), .Y(u2__abc_52155_new_n12496_));
AND2X2 AND2X2_5417 ( .A(u2__abc_52155_new_n4395_), .B(u2__abc_52155_new_n4384_), .Y(u2__abc_52155_new_n12497_));
AND2X2 AND2X2_5418 ( .A(u2__abc_52155_new_n12351_), .B(u2__abc_52155_new_n4414_), .Y(u2__abc_52155_new_n12501_));
AND2X2 AND2X2_5419 ( .A(u2__abc_52155_new_n12502_), .B(u2__abc_52155_new_n4295_), .Y(u2__abc_52155_new_n12503_));
AND2X2 AND2X2_542 ( .A(u2__abc_52155_new_n3007_), .B(u2_remHi_449_), .Y(u2__abc_52155_new_n3008_));
AND2X2 AND2X2_5420 ( .A(u2__abc_52155_new_n12505_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12506_));
AND2X2 AND2X2_5421 ( .A(u2__abc_52155_new_n12506_), .B(u2__abc_52155_new_n12504_), .Y(u2__abc_52155_new_n12507_));
AND2X2 AND2X2_5422 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_246_), .Y(u2__abc_52155_new_n12508_));
AND2X2 AND2X2_5423 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4307_), .Y(u2__abc_52155_new_n12511_));
AND2X2 AND2X2_5424 ( .A(u2__abc_52155_new_n12512_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12513_));
AND2X2 AND2X2_5425 ( .A(u2__abc_52155_new_n12510_), .B(u2__abc_52155_new_n12513_), .Y(u2__abc_52155_new_n12514_));
AND2X2 AND2X2_5426 ( .A(u2__abc_52155_new_n12515_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__248_));
AND2X2 AND2X2_5427 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_249_), .Y(u2__abc_52155_new_n12517_));
AND2X2 AND2X2_5428 ( .A(u2__abc_52155_new_n12504_), .B(u2__abc_52155_new_n4291_), .Y(u2__abc_52155_new_n12518_));
AND2X2 AND2X2_5429 ( .A(u2__abc_52155_new_n12518_), .B(u2__abc_52155_new_n4302_), .Y(u2__abc_52155_new_n12519_));
AND2X2 AND2X2_543 ( .A(u2__abc_52155_new_n3006_), .B(u2__abc_52155_new_n3009_), .Y(u2__abc_52155_new_n3010_));
AND2X2 AND2X2_5430 ( .A(u2__abc_52155_new_n12521_), .B(u2__abc_52155_new_n12520_), .Y(u2__abc_52155_new_n12522_));
AND2X2 AND2X2_5431 ( .A(u2__abc_52155_new_n12523_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12524_));
AND2X2 AND2X2_5432 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_247_), .Y(u2__abc_52155_new_n12525_));
AND2X2 AND2X2_5433 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4314_), .Y(u2__abc_52155_new_n12528_));
AND2X2 AND2X2_5434 ( .A(u2__abc_52155_new_n12529_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12530_));
AND2X2 AND2X2_5435 ( .A(u2__abc_52155_new_n12527_), .B(u2__abc_52155_new_n12530_), .Y(u2__abc_52155_new_n12531_));
AND2X2 AND2X2_5436 ( .A(u2__abc_52155_new_n12532_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__249_));
AND2X2 AND2X2_5437 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_250_), .Y(u2__abc_52155_new_n12534_));
AND2X2 AND2X2_5438 ( .A(u2__abc_52155_new_n12535_), .B(u2__abc_52155_new_n4298_), .Y(u2__abc_52155_new_n12536_));
AND2X2 AND2X2_5439 ( .A(u2__abc_52155_new_n12502_), .B(u2__abc_52155_new_n4303_), .Y(u2__abc_52155_new_n12538_));
AND2X2 AND2X2_544 ( .A(u2__abc_52155_new_n3011_), .B(u2_o_448_), .Y(u2__abc_52155_new_n3012_));
AND2X2 AND2X2_5440 ( .A(u2__abc_52155_new_n12539_), .B(u2__abc_52155_new_n4310_), .Y(u2__abc_52155_new_n12540_));
AND2X2 AND2X2_5441 ( .A(u2__abc_52155_new_n12542_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12543_));
AND2X2 AND2X2_5442 ( .A(u2__abc_52155_new_n12543_), .B(u2__abc_52155_new_n12541_), .Y(u2__abc_52155_new_n12544_));
AND2X2 AND2X2_5443 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_248_), .Y(u2__abc_52155_new_n12545_));
AND2X2 AND2X2_5444 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4345_), .Y(u2__abc_52155_new_n12548_));
AND2X2 AND2X2_5445 ( .A(u2__abc_52155_new_n12549_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12550_));
AND2X2 AND2X2_5446 ( .A(u2__abc_52155_new_n12547_), .B(u2__abc_52155_new_n12550_), .Y(u2__abc_52155_new_n12551_));
AND2X2 AND2X2_5447 ( .A(u2__abc_52155_new_n12552_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__250_));
AND2X2 AND2X2_5448 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_251_), .Y(u2__abc_52155_new_n12554_));
AND2X2 AND2X2_5449 ( .A(u2__abc_52155_new_n12541_), .B(u2__abc_52155_new_n4306_), .Y(u2__abc_52155_new_n12555_));
AND2X2 AND2X2_545 ( .A(u2__abc_52155_new_n3013_), .B(u2_remHi_448_), .Y(u2__abc_52155_new_n3014_));
AND2X2 AND2X2_5450 ( .A(u2__abc_52155_new_n12555_), .B(u2__abc_52155_new_n4317_), .Y(u2__abc_52155_new_n12556_));
AND2X2 AND2X2_5451 ( .A(u2__abc_52155_new_n12558_), .B(u2__abc_52155_new_n12557_), .Y(u2__abc_52155_new_n12559_));
AND2X2 AND2X2_5452 ( .A(u2__abc_52155_new_n12560_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12561_));
AND2X2 AND2X2_5453 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_249_), .Y(u2__abc_52155_new_n12562_));
AND2X2 AND2X2_5454 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4338_), .Y(u2__abc_52155_new_n12565_));
AND2X2 AND2X2_5455 ( .A(u2__abc_52155_new_n12566_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12567_));
AND2X2 AND2X2_5456 ( .A(u2__abc_52155_new_n12564_), .B(u2__abc_52155_new_n12567_), .Y(u2__abc_52155_new_n12568_));
AND2X2 AND2X2_5457 ( .A(u2__abc_52155_new_n12569_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__251_));
AND2X2 AND2X2_5458 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_252_), .Y(u2__abc_52155_new_n12571_));
AND2X2 AND2X2_5459 ( .A(u2__abc_52155_new_n12537_), .B(u2__abc_52155_new_n4318_), .Y(u2__abc_52155_new_n12572_));
AND2X2 AND2X2_546 ( .A(u2__abc_52155_new_n3016_), .B(u2__abc_52155_new_n3010_), .Y(u2__abc_52155_new_n3017_));
AND2X2 AND2X2_5460 ( .A(u2__abc_52155_new_n4316_), .B(u2__abc_52155_new_n4305_), .Y(u2__abc_52155_new_n12573_));
AND2X2 AND2X2_5461 ( .A(u2__abc_52155_new_n12502_), .B(u2__abc_52155_new_n4319_), .Y(u2__abc_52155_new_n12576_));
AND2X2 AND2X2_5462 ( .A(u2__abc_52155_new_n12577_), .B(u2__abc_52155_new_n4348_), .Y(u2__abc_52155_new_n12578_));
AND2X2 AND2X2_5463 ( .A(u2__abc_52155_new_n12580_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12581_));
AND2X2 AND2X2_5464 ( .A(u2__abc_52155_new_n12581_), .B(u2__abc_52155_new_n12579_), .Y(u2__abc_52155_new_n12582_));
AND2X2 AND2X2_5465 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_250_), .Y(u2__abc_52155_new_n12583_));
AND2X2 AND2X2_5466 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4323_), .Y(u2__abc_52155_new_n12586_));
AND2X2 AND2X2_5467 ( .A(u2__abc_52155_new_n12587_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12588_));
AND2X2 AND2X2_5468 ( .A(u2__abc_52155_new_n12585_), .B(u2__abc_52155_new_n12588_), .Y(u2__abc_52155_new_n12589_));
AND2X2 AND2X2_5469 ( .A(u2__abc_52155_new_n12590_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__252_));
AND2X2 AND2X2_547 ( .A(u2__abc_52155_new_n3018_), .B(u2_remHi_447_), .Y(u2__abc_52155_new_n3019_));
AND2X2 AND2X2_5470 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_253_), .Y(u2__abc_52155_new_n12592_));
AND2X2 AND2X2_5471 ( .A(u2__abc_52155_new_n12579_), .B(u2__abc_52155_new_n4344_), .Y(u2__abc_52155_new_n12593_));
AND2X2 AND2X2_5472 ( .A(u2__abc_52155_new_n12593_), .B(u2__abc_52155_new_n4341_), .Y(u2__abc_52155_new_n12594_));
AND2X2 AND2X2_5473 ( .A(u2__abc_52155_new_n12596_), .B(u2__abc_52155_new_n12595_), .Y(u2__abc_52155_new_n12597_));
AND2X2 AND2X2_5474 ( .A(u2__abc_52155_new_n12598_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12599_));
AND2X2 AND2X2_5475 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_251_), .Y(u2__abc_52155_new_n12600_));
AND2X2 AND2X2_5476 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4327_), .Y(u2__abc_52155_new_n12603_));
AND2X2 AND2X2_5477 ( .A(u2__abc_52155_new_n12604_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12605_));
AND2X2 AND2X2_5478 ( .A(u2__abc_52155_new_n12602_), .B(u2__abc_52155_new_n12605_), .Y(u2__abc_52155_new_n12606_));
AND2X2 AND2X2_5479 ( .A(u2__abc_52155_new_n12607_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__253_));
AND2X2 AND2X2_548 ( .A(u2__abc_52155_new_n3021_), .B(u2_o_447_), .Y(u2__abc_52155_new_n3022_));
AND2X2 AND2X2_5480 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_254_), .Y(u2__abc_52155_new_n12609_));
AND2X2 AND2X2_5481 ( .A(u2__abc_52155_new_n4337_), .B(u2__abc_52155_new_n4344_), .Y(u2__abc_52155_new_n12610_));
AND2X2 AND2X2_5482 ( .A(u2__abc_52155_new_n12579_), .B(u2__abc_52155_new_n12610_), .Y(u2__abc_52155_new_n12611_));
AND2X2 AND2X2_5483 ( .A(u2__abc_52155_new_n12613_), .B(u2__abc_52155_new_n4326_), .Y(u2__abc_52155_new_n12614_));
AND2X2 AND2X2_5484 ( .A(u2__abc_52155_new_n12616_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12617_));
AND2X2 AND2X2_5485 ( .A(u2__abc_52155_new_n12617_), .B(u2__abc_52155_new_n12615_), .Y(u2__abc_52155_new_n12618_));
AND2X2 AND2X2_5486 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_252_), .Y(u2__abc_52155_new_n12619_));
AND2X2 AND2X2_5487 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6539_), .Y(u2__abc_52155_new_n12622_));
AND2X2 AND2X2_5488 ( .A(u2__abc_52155_new_n12623_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12624_));
AND2X2 AND2X2_5489 ( .A(u2__abc_52155_new_n12621_), .B(u2__abc_52155_new_n12624_), .Y(u2__abc_52155_new_n12625_));
AND2X2 AND2X2_549 ( .A(u2__abc_52155_new_n3020_), .B(u2__abc_52155_new_n3023_), .Y(u2__abc_52155_new_n3024_));
AND2X2 AND2X2_5490 ( .A(u2__abc_52155_new_n12626_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__254_));
AND2X2 AND2X2_5491 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_255_), .Y(u2__abc_52155_new_n12628_));
AND2X2 AND2X2_5492 ( .A(u2__abc_52155_new_n12615_), .B(u2__abc_52155_new_n4322_), .Y(u2__abc_52155_new_n12629_));
AND2X2 AND2X2_5493 ( .A(u2__abc_52155_new_n12629_), .B(u2__abc_52155_new_n4333_), .Y(u2__abc_52155_new_n12630_));
AND2X2 AND2X2_5494 ( .A(u2__abc_52155_new_n12632_), .B(u2__abc_52155_new_n12631_), .Y(u2__abc_52155_new_n12633_));
AND2X2 AND2X2_5495 ( .A(u2__abc_52155_new_n12634_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12635_));
AND2X2 AND2X2_5496 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_253_), .Y(u2__abc_52155_new_n12636_));
AND2X2 AND2X2_5497 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6546_), .Y(u2__abc_52155_new_n12639_));
AND2X2 AND2X2_5498 ( .A(u2__abc_52155_new_n12640_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12641_));
AND2X2 AND2X2_5499 ( .A(u2__abc_52155_new_n12638_), .B(u2__abc_52155_new_n12641_), .Y(u2__abc_52155_new_n12642_));
AND2X2 AND2X2_55 ( .A(_abc_73687_new_n753_), .B(sqrto_54_), .Y(\o[90] ));
AND2X2 AND2X2_550 ( .A(u2__abc_52155_new_n3025_), .B(u2_remHi_446_), .Y(u2__abc_52155_new_n3026_));
AND2X2 AND2X2_5500 ( .A(u2__abc_52155_new_n12643_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__255_));
AND2X2 AND2X2_5501 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_256_), .Y(u2__abc_52155_new_n12645_));
AND2X2 AND2X2_5502 ( .A(u2__abc_52155_new_n10150_), .B(u2__abc_52155_new_n5287_), .Y(u2__abc_52155_new_n12646_));
AND2X2 AND2X2_5503 ( .A(u2__abc_52155_new_n11409_), .B(u2__abc_52155_new_n4796_), .Y(u2__abc_52155_new_n12647_));
AND2X2 AND2X2_5504 ( .A(u2__abc_52155_new_n12031_), .B(u2__abc_52155_new_n4543_), .Y(u2__abc_52155_new_n12648_));
AND2X2 AND2X2_5505 ( .A(u2__abc_52155_new_n12349_), .B(u2__abc_52155_new_n4415_), .Y(u2__abc_52155_new_n12649_));
AND2X2 AND2X2_5506 ( .A(u2__abc_52155_new_n12500_), .B(u2__abc_52155_new_n4351_), .Y(u2__abc_52155_new_n12650_));
AND2X2 AND2X2_5507 ( .A(u2__abc_52155_new_n12575_), .B(u2__abc_52155_new_n4350_), .Y(u2__abc_52155_new_n12651_));
AND2X2 AND2X2_5508 ( .A(u2__abc_52155_new_n12653_), .B(u2__abc_52155_new_n4334_), .Y(u2__abc_52155_new_n12654_));
AND2X2 AND2X2_5509 ( .A(u2__abc_52155_new_n4329_), .B(u2__abc_52155_new_n4321_), .Y(u2__abc_52155_new_n12655_));
AND2X2 AND2X2_551 ( .A(u2__abc_52155_new_n3028_), .B(u2_o_446_), .Y(u2__abc_52155_new_n3029_));
AND2X2 AND2X2_5510 ( .A(u2__abc_52155_new_n12663_), .B(u2__abc_52155_new_n6545_), .Y(u2__abc_52155_new_n12664_));
AND2X2 AND2X2_5511 ( .A(u2__abc_52155_new_n12666_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12667_));
AND2X2 AND2X2_5512 ( .A(u2__abc_52155_new_n12667_), .B(u2__abc_52155_new_n12665_), .Y(u2__abc_52155_new_n12668_));
AND2X2 AND2X2_5513 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_254_), .Y(u2__abc_52155_new_n12669_));
AND2X2 AND2X2_5514 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6557_), .Y(u2__abc_52155_new_n12672_));
AND2X2 AND2X2_5515 ( .A(u2__abc_52155_new_n12673_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12674_));
AND2X2 AND2X2_5516 ( .A(u2__abc_52155_new_n12671_), .B(u2__abc_52155_new_n12674_), .Y(u2__abc_52155_new_n12675_));
AND2X2 AND2X2_5517 ( .A(u2__abc_52155_new_n12676_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__256_));
AND2X2 AND2X2_5518 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_257_), .Y(u2__abc_52155_new_n12678_));
AND2X2 AND2X2_5519 ( .A(u2__abc_52155_new_n12665_), .B(u2__abc_52155_new_n6544_), .Y(u2__abc_52155_new_n12680_));
AND2X2 AND2X2_552 ( .A(u2__abc_52155_new_n3027_), .B(u2__abc_52155_new_n3030_), .Y(u2__abc_52155_new_n3031_));
AND2X2 AND2X2_5520 ( .A(u2__abc_52155_new_n12683_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12684_));
AND2X2 AND2X2_5521 ( .A(u2__abc_52155_new_n12684_), .B(u2__abc_52155_new_n12681_), .Y(u2__abc_52155_new_n12685_));
AND2X2 AND2X2_5522 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_255_), .Y(u2__abc_52155_new_n12686_));
AND2X2 AND2X2_5523 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6564_), .Y(u2__abc_52155_new_n12689_));
AND2X2 AND2X2_5524 ( .A(u2__abc_52155_new_n12690_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12691_));
AND2X2 AND2X2_5525 ( .A(u2__abc_52155_new_n12688_), .B(u2__abc_52155_new_n12691_), .Y(u2__abc_52155_new_n12692_));
AND2X2 AND2X2_5526 ( .A(u2__abc_52155_new_n12693_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__257_));
AND2X2 AND2X2_5527 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_258_), .Y(u2__abc_52155_new_n12695_));
AND2X2 AND2X2_5528 ( .A(u2__abc_52155_new_n6544_), .B(u2__abc_52155_new_n6551_), .Y(u2__abc_52155_new_n12696_));
AND2X2 AND2X2_5529 ( .A(u2__abc_52155_new_n12663_), .B(u2__abc_52155_new_n6553_), .Y(u2__abc_52155_new_n12699_));
AND2X2 AND2X2_553 ( .A(u2__abc_52155_new_n3024_), .B(u2__abc_52155_new_n3031_), .Y(u2__abc_52155_new_n3032_));
AND2X2 AND2X2_5530 ( .A(u2__abc_52155_new_n12700_), .B(u2__abc_52155_new_n6560_), .Y(u2__abc_52155_new_n12701_));
AND2X2 AND2X2_5531 ( .A(u2__abc_52155_new_n12703_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12704_));
AND2X2 AND2X2_5532 ( .A(u2__abc_52155_new_n12704_), .B(u2__abc_52155_new_n12702_), .Y(u2__abc_52155_new_n12705_));
AND2X2 AND2X2_5533 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_256_), .Y(u2__abc_52155_new_n12706_));
AND2X2 AND2X2_5534 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6588_), .Y(u2__abc_52155_new_n12709_));
AND2X2 AND2X2_5535 ( .A(u2__abc_52155_new_n12710_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12711_));
AND2X2 AND2X2_5536 ( .A(u2__abc_52155_new_n12708_), .B(u2__abc_52155_new_n12711_), .Y(u2__abc_52155_new_n12712_));
AND2X2 AND2X2_5537 ( .A(u2__abc_52155_new_n12713_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__258_));
AND2X2 AND2X2_5538 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_259_), .Y(u2__abc_52155_new_n12715_));
AND2X2 AND2X2_5539 ( .A(u2__abc_52155_new_n12702_), .B(u2__abc_52155_new_n6556_), .Y(u2__abc_52155_new_n12717_));
AND2X2 AND2X2_554 ( .A(u2__abc_52155_new_n3017_), .B(u2__abc_52155_new_n3032_), .Y(u2__abc_52155_new_n3033_));
AND2X2 AND2X2_5540 ( .A(u2__abc_52155_new_n12720_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12721_));
AND2X2 AND2X2_5541 ( .A(u2__abc_52155_new_n12721_), .B(u2__abc_52155_new_n12718_), .Y(u2__abc_52155_new_n12722_));
AND2X2 AND2X2_5542 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_257_), .Y(u2__abc_52155_new_n12723_));
AND2X2 AND2X2_5543 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6595_), .Y(u2__abc_52155_new_n12726_));
AND2X2 AND2X2_5544 ( .A(u2__abc_52155_new_n12727_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12728_));
AND2X2 AND2X2_5545 ( .A(u2__abc_52155_new_n12725_), .B(u2__abc_52155_new_n12728_), .Y(u2__abc_52155_new_n12729_));
AND2X2 AND2X2_5546 ( .A(u2__abc_52155_new_n12730_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__259_));
AND2X2 AND2X2_5547 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_260_), .Y(u2__abc_52155_new_n12732_));
AND2X2 AND2X2_5548 ( .A(u2__abc_52155_new_n12698_), .B(u2__abc_52155_new_n6568_), .Y(u2__abc_52155_new_n12733_));
AND2X2 AND2X2_5549 ( .A(u2__abc_52155_new_n6566_), .B(u2__abc_52155_new_n6555_), .Y(u2__abc_52155_new_n12734_));
AND2X2 AND2X2_555 ( .A(u2__abc_52155_new_n3035_), .B(u2_remHi_12_), .Y(u2__abc_52155_new_n3036_));
AND2X2 AND2X2_5550 ( .A(u2__abc_52155_new_n12663_), .B(u2__abc_52155_new_n6569_), .Y(u2__abc_52155_new_n12737_));
AND2X2 AND2X2_5551 ( .A(u2__abc_52155_new_n12738_), .B(u2__abc_52155_new_n6591_), .Y(u2__abc_52155_new_n12739_));
AND2X2 AND2X2_5552 ( .A(u2__abc_52155_new_n12741_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12742_));
AND2X2 AND2X2_5553 ( .A(u2__abc_52155_new_n12742_), .B(u2__abc_52155_new_n12740_), .Y(u2__abc_52155_new_n12743_));
AND2X2 AND2X2_5554 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_258_), .Y(u2__abc_52155_new_n12744_));
AND2X2 AND2X2_5555 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6573_), .Y(u2__abc_52155_new_n12747_));
AND2X2 AND2X2_5556 ( .A(u2__abc_52155_new_n12748_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12749_));
AND2X2 AND2X2_5557 ( .A(u2__abc_52155_new_n12746_), .B(u2__abc_52155_new_n12749_), .Y(u2__abc_52155_new_n12750_));
AND2X2 AND2X2_5558 ( .A(u2__abc_52155_new_n12751_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__260_));
AND2X2 AND2X2_5559 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_261_), .Y(u2__abc_52155_new_n12753_));
AND2X2 AND2X2_556 ( .A(u2__abc_52155_new_n3037_), .B(sqrto_12_), .Y(u2__abc_52155_new_n3038_));
AND2X2 AND2X2_5560 ( .A(u2__abc_52155_new_n12740_), .B(u2__abc_52155_new_n6587_), .Y(u2__abc_52155_new_n12754_));
AND2X2 AND2X2_5561 ( .A(u2__abc_52155_new_n12754_), .B(u2__abc_52155_new_n6598_), .Y(u2__abc_52155_new_n12755_));
AND2X2 AND2X2_5562 ( .A(u2__abc_52155_new_n12757_), .B(u2__abc_52155_new_n12756_), .Y(u2__abc_52155_new_n12758_));
AND2X2 AND2X2_5563 ( .A(u2__abc_52155_new_n12759_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12760_));
AND2X2 AND2X2_5564 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_259_), .Y(u2__abc_52155_new_n12761_));
AND2X2 AND2X2_5565 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6580_), .Y(u2__abc_52155_new_n12764_));
AND2X2 AND2X2_5566 ( .A(u2__abc_52155_new_n12765_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12766_));
AND2X2 AND2X2_5567 ( .A(u2__abc_52155_new_n12763_), .B(u2__abc_52155_new_n12766_), .Y(u2__abc_52155_new_n12767_));
AND2X2 AND2X2_5568 ( .A(u2__abc_52155_new_n12768_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__261_));
AND2X2 AND2X2_5569 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_262_), .Y(u2__abc_52155_new_n12770_));
AND2X2 AND2X2_557 ( .A(u2__abc_52155_new_n3041_), .B(sqrto_13_), .Y(u2__abc_52155_new_n3042_));
AND2X2 AND2X2_5570 ( .A(u2__abc_52155_new_n6587_), .B(u2__abc_52155_new_n6594_), .Y(u2__abc_52155_new_n12771_));
AND2X2 AND2X2_5571 ( .A(u2__abc_52155_new_n12740_), .B(u2__abc_52155_new_n12771_), .Y(u2__abc_52155_new_n12772_));
AND2X2 AND2X2_5572 ( .A(u2__abc_52155_new_n12774_), .B(u2__abc_52155_new_n6576_), .Y(u2__abc_52155_new_n12775_));
AND2X2 AND2X2_5573 ( .A(u2__abc_52155_new_n12777_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12778_));
AND2X2 AND2X2_5574 ( .A(u2__abc_52155_new_n12778_), .B(u2__abc_52155_new_n12776_), .Y(u2__abc_52155_new_n12779_));
AND2X2 AND2X2_5575 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_260_), .Y(u2__abc_52155_new_n12780_));
AND2X2 AND2X2_5576 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6522_), .Y(u2__abc_52155_new_n12783_));
AND2X2 AND2X2_5577 ( .A(u2__abc_52155_new_n12784_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12785_));
AND2X2 AND2X2_5578 ( .A(u2__abc_52155_new_n12782_), .B(u2__abc_52155_new_n12785_), .Y(u2__abc_52155_new_n12786_));
AND2X2 AND2X2_5579 ( .A(u2__abc_52155_new_n12787_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__262_));
AND2X2 AND2X2_558 ( .A(u2__abc_52155_new_n3043_), .B(u2_remHi_13_), .Y(u2__abc_52155_new_n3044_));
AND2X2 AND2X2_5580 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_263_), .Y(u2__abc_52155_new_n12789_));
AND2X2 AND2X2_5581 ( .A(u2__abc_52155_new_n12776_), .B(u2__abc_52155_new_n6572_), .Y(u2__abc_52155_new_n12791_));
AND2X2 AND2X2_5582 ( .A(u2__abc_52155_new_n12794_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12795_));
AND2X2 AND2X2_5583 ( .A(u2__abc_52155_new_n12795_), .B(u2__abc_52155_new_n12792_), .Y(u2__abc_52155_new_n12796_));
AND2X2 AND2X2_5584 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_261_), .Y(u2__abc_52155_new_n12797_));
AND2X2 AND2X2_5585 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6529_), .Y(u2__abc_52155_new_n12800_));
AND2X2 AND2X2_5586 ( .A(u2__abc_52155_new_n12801_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12802_));
AND2X2 AND2X2_5587 ( .A(u2__abc_52155_new_n12799_), .B(u2__abc_52155_new_n12802_), .Y(u2__abc_52155_new_n12803_));
AND2X2 AND2X2_5588 ( .A(u2__abc_52155_new_n12804_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__263_));
AND2X2 AND2X2_5589 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_264_), .Y(u2__abc_52155_new_n12806_));
AND2X2 AND2X2_559 ( .A(u2__abc_52155_new_n3040_), .B(u2__abc_52155_new_n3046_), .Y(u2__abc_52155_new_n3047_));
AND2X2 AND2X2_5590 ( .A(u2__abc_52155_new_n12736_), .B(u2__abc_52155_new_n6600_), .Y(u2__abc_52155_new_n12807_));
AND2X2 AND2X2_5591 ( .A(u2__abc_52155_new_n12811_), .B(u2__abc_52155_new_n6582_), .Y(u2__abc_52155_new_n12812_));
AND2X2 AND2X2_5592 ( .A(u2__abc_52155_new_n12810_), .B(u2__abc_52155_new_n12813_), .Y(u2__abc_52155_new_n12814_));
AND2X2 AND2X2_5593 ( .A(u2__abc_52155_new_n12808_), .B(u2__abc_52155_new_n12814_), .Y(u2__abc_52155_new_n12815_));
AND2X2 AND2X2_5594 ( .A(u2__abc_52155_new_n12663_), .B(u2__abc_52155_new_n6601_), .Y(u2__abc_52155_new_n12817_));
AND2X2 AND2X2_5595 ( .A(u2__abc_52155_new_n12818_), .B(u2__abc_52155_new_n6528_), .Y(u2__abc_52155_new_n12819_));
AND2X2 AND2X2_5596 ( .A(u2__abc_52155_new_n12821_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12822_));
AND2X2 AND2X2_5597 ( .A(u2__abc_52155_new_n12822_), .B(u2__abc_52155_new_n12820_), .Y(u2__abc_52155_new_n12823_));
AND2X2 AND2X2_5598 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_262_), .Y(u2__abc_52155_new_n12824_));
AND2X2 AND2X2_5599 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6510_), .Y(u2__abc_52155_new_n12827_));
AND2X2 AND2X2_56 ( .A(_abc_73687_new_n753_), .B(sqrto_55_), .Y(\o[91] ));
AND2X2 AND2X2_560 ( .A(u2__abc_52155_new_n3048_), .B(u2_remHi_11_), .Y(u2__abc_52155_new_n3049_));
AND2X2 AND2X2_5600 ( .A(u2__abc_52155_new_n12828_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12829_));
AND2X2 AND2X2_5601 ( .A(u2__abc_52155_new_n12826_), .B(u2__abc_52155_new_n12829_), .Y(u2__abc_52155_new_n12830_));
AND2X2 AND2X2_5602 ( .A(u2__abc_52155_new_n12831_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__264_));
AND2X2 AND2X2_5603 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_265_), .Y(u2__abc_52155_new_n12833_));
AND2X2 AND2X2_5604 ( .A(u2__abc_52155_new_n12820_), .B(u2__abc_52155_new_n6527_), .Y(u2__abc_52155_new_n12835_));
AND2X2 AND2X2_5605 ( .A(u2__abc_52155_new_n12838_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12839_));
AND2X2 AND2X2_5606 ( .A(u2__abc_52155_new_n12839_), .B(u2__abc_52155_new_n12836_), .Y(u2__abc_52155_new_n12840_));
AND2X2 AND2X2_5607 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_263_), .Y(u2__abc_52155_new_n12841_));
AND2X2 AND2X2_5608 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6517_), .Y(u2__abc_52155_new_n12844_));
AND2X2 AND2X2_5609 ( .A(u2__abc_52155_new_n12845_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12846_));
AND2X2 AND2X2_561 ( .A(u2__abc_52155_new_n3051_), .B(sqrto_11_), .Y(u2__abc_52155_new_n3052_));
AND2X2 AND2X2_5610 ( .A(u2__abc_52155_new_n12843_), .B(u2__abc_52155_new_n12846_), .Y(u2__abc_52155_new_n12847_));
AND2X2 AND2X2_5611 ( .A(u2__abc_52155_new_n12848_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__265_));
AND2X2 AND2X2_5612 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_266_), .Y(u2__abc_52155_new_n12850_));
AND2X2 AND2X2_5613 ( .A(u2__abc_52155_new_n6527_), .B(u2__abc_52155_new_n6534_), .Y(u2__abc_52155_new_n12851_));
AND2X2 AND2X2_5614 ( .A(u2__abc_52155_new_n12818_), .B(u2__abc_52155_new_n6536_), .Y(u2__abc_52155_new_n12854_));
AND2X2 AND2X2_5615 ( .A(u2__abc_52155_new_n12855_), .B(u2__abc_52155_new_n6513_), .Y(u2__abc_52155_new_n12856_));
AND2X2 AND2X2_5616 ( .A(u2__abc_52155_new_n12858_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12859_));
AND2X2 AND2X2_5617 ( .A(u2__abc_52155_new_n12859_), .B(u2__abc_52155_new_n12857_), .Y(u2__abc_52155_new_n12860_));
AND2X2 AND2X2_5618 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_264_), .Y(u2__abc_52155_new_n12861_));
AND2X2 AND2X2_5619 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6494_), .Y(u2__abc_52155_new_n12864_));
AND2X2 AND2X2_562 ( .A(u2__abc_52155_new_n3050_), .B(u2__abc_52155_new_n3053_), .Y(u2__abc_52155_new_n3054_));
AND2X2 AND2X2_5620 ( .A(u2__abc_52155_new_n12865_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12866_));
AND2X2 AND2X2_5621 ( .A(u2__abc_52155_new_n12863_), .B(u2__abc_52155_new_n12866_), .Y(u2__abc_52155_new_n12867_));
AND2X2 AND2X2_5622 ( .A(u2__abc_52155_new_n12868_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__266_));
AND2X2 AND2X2_5623 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_267_), .Y(u2__abc_52155_new_n12870_));
AND2X2 AND2X2_5624 ( .A(u2__abc_52155_new_n12857_), .B(u2__abc_52155_new_n6509_), .Y(u2__abc_52155_new_n12872_));
AND2X2 AND2X2_5625 ( .A(u2__abc_52155_new_n12875_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12876_));
AND2X2 AND2X2_5626 ( .A(u2__abc_52155_new_n12876_), .B(u2__abc_52155_new_n12873_), .Y(u2__abc_52155_new_n12877_));
AND2X2 AND2X2_5627 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_265_), .Y(u2__abc_52155_new_n12878_));
AND2X2 AND2X2_5628 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6501_), .Y(u2__abc_52155_new_n12881_));
AND2X2 AND2X2_5629 ( .A(u2__abc_52155_new_n12882_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12883_));
AND2X2 AND2X2_563 ( .A(u2__abc_52155_new_n3055_), .B(u2_remHi_10_), .Y(u2__abc_52155_new_n3056_));
AND2X2 AND2X2_5630 ( .A(u2__abc_52155_new_n12880_), .B(u2__abc_52155_new_n12883_), .Y(u2__abc_52155_new_n12884_));
AND2X2 AND2X2_5631 ( .A(u2__abc_52155_new_n12885_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__267_));
AND2X2 AND2X2_5632 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_268_), .Y(u2__abc_52155_new_n12887_));
AND2X2 AND2X2_5633 ( .A(u2__abc_52155_new_n6509_), .B(u2__abc_52155_new_n6516_), .Y(u2__abc_52155_new_n12888_));
AND2X2 AND2X2_5634 ( .A(u2__abc_52155_new_n12857_), .B(u2__abc_52155_new_n12888_), .Y(u2__abc_52155_new_n12889_));
AND2X2 AND2X2_5635 ( .A(u2__abc_52155_new_n12891_), .B(u2__abc_52155_new_n6497_), .Y(u2__abc_52155_new_n12892_));
AND2X2 AND2X2_5636 ( .A(u2__abc_52155_new_n12894_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12895_));
AND2X2 AND2X2_5637 ( .A(u2__abc_52155_new_n12895_), .B(u2__abc_52155_new_n12893_), .Y(u2__abc_52155_new_n12896_));
AND2X2 AND2X2_5638 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_266_), .Y(u2__abc_52155_new_n12897_));
AND2X2 AND2X2_5639 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6476_), .Y(u2__abc_52155_new_n12900_));
AND2X2 AND2X2_564 ( .A(u2__abc_52155_new_n3057_), .B(sqrto_10_), .Y(u2__abc_52155_new_n3058_));
AND2X2 AND2X2_5640 ( .A(u2__abc_52155_new_n12901_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12902_));
AND2X2 AND2X2_5641 ( .A(u2__abc_52155_new_n12899_), .B(u2__abc_52155_new_n12902_), .Y(u2__abc_52155_new_n12903_));
AND2X2 AND2X2_5642 ( .A(u2__abc_52155_new_n12904_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__268_));
AND2X2 AND2X2_5643 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_269_), .Y(u2__abc_52155_new_n12906_));
AND2X2 AND2X2_5644 ( .A(u2__abc_52155_new_n12893_), .B(u2__abc_52155_new_n6493_), .Y(u2__abc_52155_new_n12907_));
AND2X2 AND2X2_5645 ( .A(u2__abc_52155_new_n12907_), .B(u2__abc_52155_new_n6504_), .Y(u2__abc_52155_new_n12908_));
AND2X2 AND2X2_5646 ( .A(u2__abc_52155_new_n12910_), .B(u2__abc_52155_new_n12909_), .Y(u2__abc_52155_new_n12911_));
AND2X2 AND2X2_5647 ( .A(u2__abc_52155_new_n12912_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12913_));
AND2X2 AND2X2_5648 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_267_), .Y(u2__abc_52155_new_n12914_));
AND2X2 AND2X2_5649 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6483_), .Y(u2__abc_52155_new_n12917_));
AND2X2 AND2X2_565 ( .A(u2__abc_52155_new_n3060_), .B(u2__abc_52155_new_n3054_), .Y(u2__abc_52155_new_n3061_));
AND2X2 AND2X2_5650 ( .A(u2__abc_52155_new_n12918_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12919_));
AND2X2 AND2X2_5651 ( .A(u2__abc_52155_new_n12916_), .B(u2__abc_52155_new_n12919_), .Y(u2__abc_52155_new_n12920_));
AND2X2 AND2X2_5652 ( .A(u2__abc_52155_new_n12921_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__269_));
AND2X2 AND2X2_5653 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_270_), .Y(u2__abc_52155_new_n12923_));
AND2X2 AND2X2_5654 ( .A(u2__abc_52155_new_n6493_), .B(u2__abc_52155_new_n6500_), .Y(u2__abc_52155_new_n12924_));
AND2X2 AND2X2_5655 ( .A(u2__abc_52155_new_n12893_), .B(u2__abc_52155_new_n12924_), .Y(u2__abc_52155_new_n12925_));
AND2X2 AND2X2_5656 ( .A(u2__abc_52155_new_n12927_), .B(u2__abc_52155_new_n6482_), .Y(u2__abc_52155_new_n12928_));
AND2X2 AND2X2_5657 ( .A(u2__abc_52155_new_n12930_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12931_));
AND2X2 AND2X2_5658 ( .A(u2__abc_52155_new_n12931_), .B(u2__abc_52155_new_n12929_), .Y(u2__abc_52155_new_n12932_));
AND2X2 AND2X2_5659 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_268_), .Y(u2__abc_52155_new_n12933_));
AND2X2 AND2X2_566 ( .A(u2__abc_52155_new_n3047_), .B(u2__abc_52155_new_n3061_), .Y(u2__abc_52155_new_n3062_));
AND2X2 AND2X2_5660 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6430_), .Y(u2__abc_52155_new_n12936_));
AND2X2 AND2X2_5661 ( .A(u2__abc_52155_new_n12937_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12938_));
AND2X2 AND2X2_5662 ( .A(u2__abc_52155_new_n12935_), .B(u2__abc_52155_new_n12938_), .Y(u2__abc_52155_new_n12939_));
AND2X2 AND2X2_5663 ( .A(u2__abc_52155_new_n12940_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__270_));
AND2X2 AND2X2_5664 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_271_), .Y(u2__abc_52155_new_n12942_));
AND2X2 AND2X2_5665 ( .A(u2__abc_52155_new_n12929_), .B(u2__abc_52155_new_n6481_), .Y(u2__abc_52155_new_n12944_));
AND2X2 AND2X2_5666 ( .A(u2__abc_52155_new_n12947_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12948_));
AND2X2 AND2X2_5667 ( .A(u2__abc_52155_new_n12948_), .B(u2__abc_52155_new_n12945_), .Y(u2__abc_52155_new_n12949_));
AND2X2 AND2X2_5668 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_269_), .Y(u2__abc_52155_new_n12950_));
AND2X2 AND2X2_5669 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6437_), .Y(u2__abc_52155_new_n12953_));
AND2X2 AND2X2_567 ( .A(u2__abc_52155_new_n3063_), .B(u2_remHi_8_), .Y(u2__abc_52155_new_n3064_));
AND2X2 AND2X2_5670 ( .A(u2__abc_52155_new_n12954_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12955_));
AND2X2 AND2X2_5671 ( .A(u2__abc_52155_new_n12952_), .B(u2__abc_52155_new_n12955_), .Y(u2__abc_52155_new_n12956_));
AND2X2 AND2X2_5672 ( .A(u2__abc_52155_new_n12957_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__271_));
AND2X2 AND2X2_5673 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_272_), .Y(u2__abc_52155_new_n12959_));
AND2X2 AND2X2_5674 ( .A(u2__abc_52155_new_n12816_), .B(u2__abc_52155_new_n6538_), .Y(u2__abc_52155_new_n12960_));
AND2X2 AND2X2_5675 ( .A(u2__abc_52155_new_n12853_), .B(u2__abc_52155_new_n6521_), .Y(u2__abc_52155_new_n12963_));
AND2X2 AND2X2_5676 ( .A(u2__abc_52155_new_n12964_), .B(u2__abc_52155_new_n12962_), .Y(u2__abc_52155_new_n12965_));
AND2X2 AND2X2_5677 ( .A(u2__abc_52155_new_n6481_), .B(u2__abc_52155_new_n6488_), .Y(u2__abc_52155_new_n12967_));
AND2X2 AND2X2_5678 ( .A(u2__abc_52155_new_n12970_), .B(u2__abc_52155_new_n12968_), .Y(u2__abc_52155_new_n12971_));
AND2X2 AND2X2_5679 ( .A(u2__abc_52155_new_n12966_), .B(u2__abc_52155_new_n12971_), .Y(u2__abc_52155_new_n12972_));
AND2X2 AND2X2_568 ( .A(u2__abc_52155_new_n3065_), .B(sqrto_8_), .Y(u2__abc_52155_new_n3066_));
AND2X2 AND2X2_5680 ( .A(u2__abc_52155_new_n12961_), .B(u2__abc_52155_new_n12972_), .Y(u2__abc_52155_new_n12973_));
AND2X2 AND2X2_5681 ( .A(u2__abc_52155_new_n12663_), .B(u2__abc_52155_new_n6602_), .Y(u2__abc_52155_new_n12975_));
AND2X2 AND2X2_5682 ( .A(u2__abc_52155_new_n12976_), .B(u2__abc_52155_new_n6433_), .Y(u2__abc_52155_new_n12977_));
AND2X2 AND2X2_5683 ( .A(u2__abc_52155_new_n12979_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12980_));
AND2X2 AND2X2_5684 ( .A(u2__abc_52155_new_n12980_), .B(u2__abc_52155_new_n12978_), .Y(u2__abc_52155_new_n12981_));
AND2X2 AND2X2_5685 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_270_), .Y(u2__abc_52155_new_n12982_));
AND2X2 AND2X2_5686 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6415_), .Y(u2__abc_52155_new_n12985_));
AND2X2 AND2X2_5687 ( .A(u2__abc_52155_new_n12986_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n12987_));
AND2X2 AND2X2_5688 ( .A(u2__abc_52155_new_n12984_), .B(u2__abc_52155_new_n12987_), .Y(u2__abc_52155_new_n12988_));
AND2X2 AND2X2_5689 ( .A(u2__abc_52155_new_n12989_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__272_));
AND2X2 AND2X2_569 ( .A(u2__abc_52155_new_n3069_), .B(u2_remHi_9_), .Y(u2__abc_52155_new_n3070_));
AND2X2 AND2X2_5690 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_273_), .Y(u2__abc_52155_new_n12991_));
AND2X2 AND2X2_5691 ( .A(u2__abc_52155_new_n12978_), .B(u2__abc_52155_new_n6429_), .Y(u2__abc_52155_new_n12992_));
AND2X2 AND2X2_5692 ( .A(u2__abc_52155_new_n12992_), .B(u2__abc_52155_new_n6440_), .Y(u2__abc_52155_new_n12993_));
AND2X2 AND2X2_5693 ( .A(u2__abc_52155_new_n12995_), .B(u2__abc_52155_new_n12994_), .Y(u2__abc_52155_new_n12996_));
AND2X2 AND2X2_5694 ( .A(u2__abc_52155_new_n12997_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n12998_));
AND2X2 AND2X2_5695 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_271_), .Y(u2__abc_52155_new_n12999_));
AND2X2 AND2X2_5696 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6422_), .Y(u2__abc_52155_new_n13002_));
AND2X2 AND2X2_5697 ( .A(u2__abc_52155_new_n13003_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13004_));
AND2X2 AND2X2_5698 ( .A(u2__abc_52155_new_n13001_), .B(u2__abc_52155_new_n13004_), .Y(u2__abc_52155_new_n13005_));
AND2X2 AND2X2_5699 ( .A(u2__abc_52155_new_n13006_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__273_));
AND2X2 AND2X2_57 ( .A(_abc_73687_new_n753_), .B(sqrto_56_), .Y(\o[92] ));
AND2X2 AND2X2_570 ( .A(u2__abc_52155_new_n3072_), .B(sqrto_9_), .Y(u2__abc_52155_new_n3073_));
AND2X2 AND2X2_5700 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_274_), .Y(u2__abc_52155_new_n13008_));
AND2X2 AND2X2_5701 ( .A(u2__abc_52155_new_n6429_), .B(u2__abc_52155_new_n6436_), .Y(u2__abc_52155_new_n13009_));
AND2X2 AND2X2_5702 ( .A(u2__abc_52155_new_n12978_), .B(u2__abc_52155_new_n13009_), .Y(u2__abc_52155_new_n13010_));
AND2X2 AND2X2_5703 ( .A(u2__abc_52155_new_n13012_), .B(u2__abc_52155_new_n6418_), .Y(u2__abc_52155_new_n13013_));
AND2X2 AND2X2_5704 ( .A(u2__abc_52155_new_n13015_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13016_));
AND2X2 AND2X2_5705 ( .A(u2__abc_52155_new_n13016_), .B(u2__abc_52155_new_n13014_), .Y(u2__abc_52155_new_n13017_));
AND2X2 AND2X2_5706 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_272_), .Y(u2__abc_52155_new_n13018_));
AND2X2 AND2X2_5707 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6461_), .Y(u2__abc_52155_new_n13021_));
AND2X2 AND2X2_5708 ( .A(u2__abc_52155_new_n13022_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13023_));
AND2X2 AND2X2_5709 ( .A(u2__abc_52155_new_n13020_), .B(u2__abc_52155_new_n13023_), .Y(u2__abc_52155_new_n13024_));
AND2X2 AND2X2_571 ( .A(u2__abc_52155_new_n3071_), .B(u2__abc_52155_new_n3074_), .Y(u2__abc_52155_new_n3075_));
AND2X2 AND2X2_5710 ( .A(u2__abc_52155_new_n13025_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__274_));
AND2X2 AND2X2_5711 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_275_), .Y(u2__abc_52155_new_n13027_));
AND2X2 AND2X2_5712 ( .A(u2__abc_52155_new_n13014_), .B(u2__abc_52155_new_n6414_), .Y(u2__abc_52155_new_n13029_));
AND2X2 AND2X2_5713 ( .A(u2__abc_52155_new_n13032_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13033_));
AND2X2 AND2X2_5714 ( .A(u2__abc_52155_new_n13033_), .B(u2__abc_52155_new_n13030_), .Y(u2__abc_52155_new_n13034_));
AND2X2 AND2X2_5715 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_273_), .Y(u2__abc_52155_new_n13035_));
AND2X2 AND2X2_5716 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6468_), .Y(u2__abc_52155_new_n13038_));
AND2X2 AND2X2_5717 ( .A(u2__abc_52155_new_n13039_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13040_));
AND2X2 AND2X2_5718 ( .A(u2__abc_52155_new_n13037_), .B(u2__abc_52155_new_n13040_), .Y(u2__abc_52155_new_n13041_));
AND2X2 AND2X2_5719 ( .A(u2__abc_52155_new_n13042_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__275_));
AND2X2 AND2X2_572 ( .A(u2__abc_52155_new_n3068_), .B(u2__abc_52155_new_n3075_), .Y(u2__abc_52155_new_n3076_));
AND2X2 AND2X2_5720 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_276_), .Y(u2__abc_52155_new_n13044_));
AND2X2 AND2X2_5721 ( .A(u2__abc_52155_new_n13045_), .B(u2__abc_52155_new_n6424_), .Y(u2__abc_52155_new_n13046_));
AND2X2 AND2X2_5722 ( .A(u2__abc_52155_new_n13049_), .B(u2__abc_52155_new_n13047_), .Y(u2__abc_52155_new_n13050_));
AND2X2 AND2X2_5723 ( .A(u2__abc_52155_new_n12976_), .B(u2__abc_52155_new_n6442_), .Y(u2__abc_52155_new_n13052_));
AND2X2 AND2X2_5724 ( .A(u2__abc_52155_new_n13053_), .B(u2__abc_52155_new_n6464_), .Y(u2__abc_52155_new_n13054_));
AND2X2 AND2X2_5725 ( .A(u2__abc_52155_new_n13056_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13057_));
AND2X2 AND2X2_5726 ( .A(u2__abc_52155_new_n13057_), .B(u2__abc_52155_new_n13055_), .Y(u2__abc_52155_new_n13058_));
AND2X2 AND2X2_5727 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_274_), .Y(u2__abc_52155_new_n13059_));
AND2X2 AND2X2_5728 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6446_), .Y(u2__abc_52155_new_n13062_));
AND2X2 AND2X2_5729 ( .A(u2__abc_52155_new_n13063_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13064_));
AND2X2 AND2X2_573 ( .A(u2__abc_52155_new_n3077_), .B(u2_remHi_7_), .Y(u2__abc_52155_new_n3078_));
AND2X2 AND2X2_5730 ( .A(u2__abc_52155_new_n13061_), .B(u2__abc_52155_new_n13064_), .Y(u2__abc_52155_new_n13065_));
AND2X2 AND2X2_5731 ( .A(u2__abc_52155_new_n13066_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__276_));
AND2X2 AND2X2_5732 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_277_), .Y(u2__abc_52155_new_n13068_));
AND2X2 AND2X2_5733 ( .A(u2__abc_52155_new_n13055_), .B(u2__abc_52155_new_n6460_), .Y(u2__abc_52155_new_n13069_));
AND2X2 AND2X2_5734 ( .A(u2__abc_52155_new_n13069_), .B(u2__abc_52155_new_n6471_), .Y(u2__abc_52155_new_n13070_));
AND2X2 AND2X2_5735 ( .A(u2__abc_52155_new_n13072_), .B(u2__abc_52155_new_n13071_), .Y(u2__abc_52155_new_n13073_));
AND2X2 AND2X2_5736 ( .A(u2__abc_52155_new_n13074_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13075_));
AND2X2 AND2X2_5737 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_275_), .Y(u2__abc_52155_new_n13076_));
AND2X2 AND2X2_5738 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6453_), .Y(u2__abc_52155_new_n13079_));
AND2X2 AND2X2_5739 ( .A(u2__abc_52155_new_n13080_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13081_));
AND2X2 AND2X2_574 ( .A(u2__abc_52155_new_n3079_), .B(u2__abc_52155_new_n3080_), .Y(u2__abc_52155_new_n3081_));
AND2X2 AND2X2_5740 ( .A(u2__abc_52155_new_n13078_), .B(u2__abc_52155_new_n13081_), .Y(u2__abc_52155_new_n13082_));
AND2X2 AND2X2_5741 ( .A(u2__abc_52155_new_n13083_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__277_));
AND2X2 AND2X2_5742 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_278_), .Y(u2__abc_52155_new_n13085_));
AND2X2 AND2X2_5743 ( .A(u2__abc_52155_new_n6460_), .B(u2__abc_52155_new_n6467_), .Y(u2__abc_52155_new_n13086_));
AND2X2 AND2X2_5744 ( .A(u2__abc_52155_new_n13055_), .B(u2__abc_52155_new_n13086_), .Y(u2__abc_52155_new_n13087_));
AND2X2 AND2X2_5745 ( .A(u2__abc_52155_new_n13089_), .B(u2__abc_52155_new_n6449_), .Y(u2__abc_52155_new_n13090_));
AND2X2 AND2X2_5746 ( .A(u2__abc_52155_new_n13092_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13093_));
AND2X2 AND2X2_5747 ( .A(u2__abc_52155_new_n13093_), .B(u2__abc_52155_new_n13091_), .Y(u2__abc_52155_new_n13094_));
AND2X2 AND2X2_5748 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_276_), .Y(u2__abc_52155_new_n13095_));
AND2X2 AND2X2_5749 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6367_), .Y(u2__abc_52155_new_n13098_));
AND2X2 AND2X2_575 ( .A(u2__abc_52155_new_n3083_), .B(u2__abc_52155_new_n3085_), .Y(u2__abc_52155_new_n3086_));
AND2X2 AND2X2_5750 ( .A(u2__abc_52155_new_n13099_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13100_));
AND2X2 AND2X2_5751 ( .A(u2__abc_52155_new_n13097_), .B(u2__abc_52155_new_n13100_), .Y(u2__abc_52155_new_n13101_));
AND2X2 AND2X2_5752 ( .A(u2__abc_52155_new_n13102_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__278_));
AND2X2 AND2X2_5753 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_279_), .Y(u2__abc_52155_new_n13104_));
AND2X2 AND2X2_5754 ( .A(u2__abc_52155_new_n13091_), .B(u2__abc_52155_new_n6445_), .Y(u2__abc_52155_new_n13106_));
AND2X2 AND2X2_5755 ( .A(u2__abc_52155_new_n13109_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13110_));
AND2X2 AND2X2_5756 ( .A(u2__abc_52155_new_n13110_), .B(u2__abc_52155_new_n13107_), .Y(u2__abc_52155_new_n13111_));
AND2X2 AND2X2_5757 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_277_), .Y(u2__abc_52155_new_n13112_));
AND2X2 AND2X2_5758 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6374_), .Y(u2__abc_52155_new_n13115_));
AND2X2 AND2X2_5759 ( .A(u2__abc_52155_new_n13116_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13117_));
AND2X2 AND2X2_576 ( .A(u2__abc_52155_new_n3081_), .B(u2__abc_52155_new_n3086_), .Y(u2__abc_52155_new_n3087_));
AND2X2 AND2X2_5760 ( .A(u2__abc_52155_new_n13114_), .B(u2__abc_52155_new_n13117_), .Y(u2__abc_52155_new_n13118_));
AND2X2 AND2X2_5761 ( .A(u2__abc_52155_new_n13119_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__279_));
AND2X2 AND2X2_5762 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_280_), .Y(u2__abc_52155_new_n13121_));
AND2X2 AND2X2_5763 ( .A(u2__abc_52155_new_n13051_), .B(u2__abc_52155_new_n6473_), .Y(u2__abc_52155_new_n13122_));
AND2X2 AND2X2_5764 ( .A(u2__abc_52155_new_n6445_), .B(u2__abc_52155_new_n6452_), .Y(u2__abc_52155_new_n13126_));
AND2X2 AND2X2_5765 ( .A(u2__abc_52155_new_n13125_), .B(u2__abc_52155_new_n13127_), .Y(u2__abc_52155_new_n13128_));
AND2X2 AND2X2_5766 ( .A(u2__abc_52155_new_n13123_), .B(u2__abc_52155_new_n13128_), .Y(u2__abc_52155_new_n13129_));
AND2X2 AND2X2_5767 ( .A(u2__abc_52155_new_n12976_), .B(u2__abc_52155_new_n6474_), .Y(u2__abc_52155_new_n13131_));
AND2X2 AND2X2_5768 ( .A(u2__abc_52155_new_n13132_), .B(u2__abc_52155_new_n6370_), .Y(u2__abc_52155_new_n13133_));
AND2X2 AND2X2_5769 ( .A(u2__abc_52155_new_n13135_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13136_));
AND2X2 AND2X2_577 ( .A(u2__abc_52155_new_n3076_), .B(u2__abc_52155_new_n3087_), .Y(u2__abc_52155_new_n3088_));
AND2X2 AND2X2_5770 ( .A(u2__abc_52155_new_n13136_), .B(u2__abc_52155_new_n13134_), .Y(u2__abc_52155_new_n13137_));
AND2X2 AND2X2_5771 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_278_), .Y(u2__abc_52155_new_n13138_));
AND2X2 AND2X2_5772 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6352_), .Y(u2__abc_52155_new_n13141_));
AND2X2 AND2X2_5773 ( .A(u2__abc_52155_new_n13142_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13143_));
AND2X2 AND2X2_5774 ( .A(u2__abc_52155_new_n13140_), .B(u2__abc_52155_new_n13143_), .Y(u2__abc_52155_new_n13144_));
AND2X2 AND2X2_5775 ( .A(u2__abc_52155_new_n13145_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__280_));
AND2X2 AND2X2_5776 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_281_), .Y(u2__abc_52155_new_n13147_));
AND2X2 AND2X2_5777 ( .A(u2__abc_52155_new_n13134_), .B(u2__abc_52155_new_n6366_), .Y(u2__abc_52155_new_n13148_));
AND2X2 AND2X2_5778 ( .A(u2__abc_52155_new_n13148_), .B(u2__abc_52155_new_n6377_), .Y(u2__abc_52155_new_n13149_));
AND2X2 AND2X2_5779 ( .A(u2__abc_52155_new_n13151_), .B(u2__abc_52155_new_n13150_), .Y(u2__abc_52155_new_n13152_));
AND2X2 AND2X2_578 ( .A(u2__abc_52155_new_n3062_), .B(u2__abc_52155_new_n3088_), .Y(u2__abc_52155_new_n3089_));
AND2X2 AND2X2_5780 ( .A(u2__abc_52155_new_n13153_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13154_));
AND2X2 AND2X2_5781 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_279_), .Y(u2__abc_52155_new_n13155_));
AND2X2 AND2X2_5782 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6359_), .Y(u2__abc_52155_new_n13158_));
AND2X2 AND2X2_5783 ( .A(u2__abc_52155_new_n13159_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13160_));
AND2X2 AND2X2_5784 ( .A(u2__abc_52155_new_n13157_), .B(u2__abc_52155_new_n13160_), .Y(u2__abc_52155_new_n13161_));
AND2X2 AND2X2_5785 ( .A(u2__abc_52155_new_n13162_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__281_));
AND2X2 AND2X2_5786 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_282_), .Y(u2__abc_52155_new_n13164_));
AND2X2 AND2X2_5787 ( .A(u2__abc_52155_new_n6366_), .B(u2__abc_52155_new_n6373_), .Y(u2__abc_52155_new_n13165_));
AND2X2 AND2X2_5788 ( .A(u2__abc_52155_new_n13134_), .B(u2__abc_52155_new_n13165_), .Y(u2__abc_52155_new_n13166_));
AND2X2 AND2X2_5789 ( .A(u2__abc_52155_new_n13168_), .B(u2__abc_52155_new_n6355_), .Y(u2__abc_52155_new_n13169_));
AND2X2 AND2X2_579 ( .A(u2__abc_52155_new_n3091_), .B(u2_remHi_4_), .Y(u2__abc_52155_new_n3092_));
AND2X2 AND2X2_5790 ( .A(u2__abc_52155_new_n13171_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13172_));
AND2X2 AND2X2_5791 ( .A(u2__abc_52155_new_n13172_), .B(u2__abc_52155_new_n13170_), .Y(u2__abc_52155_new_n13173_));
AND2X2 AND2X2_5792 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_280_), .Y(u2__abc_52155_new_n13174_));
AND2X2 AND2X2_5793 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6398_), .Y(u2__abc_52155_new_n13177_));
AND2X2 AND2X2_5794 ( .A(u2__abc_52155_new_n13178_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13179_));
AND2X2 AND2X2_5795 ( .A(u2__abc_52155_new_n13176_), .B(u2__abc_52155_new_n13179_), .Y(u2__abc_52155_new_n13180_));
AND2X2 AND2X2_5796 ( .A(u2__abc_52155_new_n13181_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__282_));
AND2X2 AND2X2_5797 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_283_), .Y(u2__abc_52155_new_n13183_));
AND2X2 AND2X2_5798 ( .A(u2__abc_52155_new_n13170_), .B(u2__abc_52155_new_n6351_), .Y(u2__abc_52155_new_n13185_));
AND2X2 AND2X2_5799 ( .A(u2__abc_52155_new_n13188_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13189_));
AND2X2 AND2X2_58 ( .A(_abc_73687_new_n753_), .B(sqrto_57_), .Y(\o[93] ));
AND2X2 AND2X2_580 ( .A(u2__abc_52155_new_n3093_), .B(sqrto_4_), .Y(u2__abc_52155_new_n3094_));
AND2X2 AND2X2_5800 ( .A(u2__abc_52155_new_n13189_), .B(u2__abc_52155_new_n13186_), .Y(u2__abc_52155_new_n13190_));
AND2X2 AND2X2_5801 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_281_), .Y(u2__abc_52155_new_n13191_));
AND2X2 AND2X2_5802 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6405_), .Y(u2__abc_52155_new_n13194_));
AND2X2 AND2X2_5803 ( .A(u2__abc_52155_new_n13195_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13196_));
AND2X2 AND2X2_5804 ( .A(u2__abc_52155_new_n13193_), .B(u2__abc_52155_new_n13196_), .Y(u2__abc_52155_new_n13197_));
AND2X2 AND2X2_5805 ( .A(u2__abc_52155_new_n13198_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__283_));
AND2X2 AND2X2_5806 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_284_), .Y(u2__abc_52155_new_n13200_));
AND2X2 AND2X2_5807 ( .A(u2__abc_52155_new_n6361_), .B(u2__abc_52155_new_n6350_), .Y(u2__abc_52155_new_n13203_));
AND2X2 AND2X2_5808 ( .A(u2__abc_52155_new_n13202_), .B(u2__abc_52155_new_n13205_), .Y(u2__abc_52155_new_n13206_));
AND2X2 AND2X2_5809 ( .A(u2__abc_52155_new_n13132_), .B(u2__abc_52155_new_n6379_), .Y(u2__abc_52155_new_n13208_));
AND2X2 AND2X2_581 ( .A(u2__abc_52155_new_n3096_), .B(sqrto_5_), .Y(u2__abc_52155_new_n3097_));
AND2X2 AND2X2_5810 ( .A(u2__abc_52155_new_n13209_), .B(u2__abc_52155_new_n6401_), .Y(u2__abc_52155_new_n13210_));
AND2X2 AND2X2_5811 ( .A(u2__abc_52155_new_n13212_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13213_));
AND2X2 AND2X2_5812 ( .A(u2__abc_52155_new_n13213_), .B(u2__abc_52155_new_n13211_), .Y(u2__abc_52155_new_n13214_));
AND2X2 AND2X2_5813 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_282_), .Y(u2__abc_52155_new_n13215_));
AND2X2 AND2X2_5814 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6383_), .Y(u2__abc_52155_new_n13218_));
AND2X2 AND2X2_5815 ( .A(u2__abc_52155_new_n13219_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13220_));
AND2X2 AND2X2_5816 ( .A(u2__abc_52155_new_n13217_), .B(u2__abc_52155_new_n13220_), .Y(u2__abc_52155_new_n13221_));
AND2X2 AND2X2_5817 ( .A(u2__abc_52155_new_n13222_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__284_));
AND2X2 AND2X2_5818 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_285_), .Y(u2__abc_52155_new_n13224_));
AND2X2 AND2X2_5819 ( .A(u2__abc_52155_new_n13211_), .B(u2__abc_52155_new_n6397_), .Y(u2__abc_52155_new_n13225_));
AND2X2 AND2X2_582 ( .A(u2__abc_52155_new_n3098_), .B(u2_remHi_5_), .Y(u2__abc_52155_new_n3099_));
AND2X2 AND2X2_5820 ( .A(u2__abc_52155_new_n13225_), .B(u2__abc_52155_new_n6408_), .Y(u2__abc_52155_new_n13226_));
AND2X2 AND2X2_5821 ( .A(u2__abc_52155_new_n13228_), .B(u2__abc_52155_new_n13227_), .Y(u2__abc_52155_new_n13229_));
AND2X2 AND2X2_5822 ( .A(u2__abc_52155_new_n13230_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13231_));
AND2X2 AND2X2_5823 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_283_), .Y(u2__abc_52155_new_n13232_));
AND2X2 AND2X2_5824 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6390_), .Y(u2__abc_52155_new_n13235_));
AND2X2 AND2X2_5825 ( .A(u2__abc_52155_new_n13236_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13237_));
AND2X2 AND2X2_5826 ( .A(u2__abc_52155_new_n13234_), .B(u2__abc_52155_new_n13237_), .Y(u2__abc_52155_new_n13238_));
AND2X2 AND2X2_5827 ( .A(u2__abc_52155_new_n13239_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__285_));
AND2X2 AND2X2_5828 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_286_), .Y(u2__abc_52155_new_n13241_));
AND2X2 AND2X2_5829 ( .A(u2__abc_52155_new_n6397_), .B(u2__abc_52155_new_n6404_), .Y(u2__abc_52155_new_n13242_));
AND2X2 AND2X2_583 ( .A(u2__abc_52155_new_n3102_), .B(u2_remHi_3_), .Y(u2__abc_52155_new_n3103_));
AND2X2 AND2X2_5830 ( .A(u2__abc_52155_new_n13211_), .B(u2__abc_52155_new_n13242_), .Y(u2__abc_52155_new_n13243_));
AND2X2 AND2X2_5831 ( .A(u2__abc_52155_new_n13245_), .B(u2__abc_52155_new_n6386_), .Y(u2__abc_52155_new_n13246_));
AND2X2 AND2X2_5832 ( .A(u2__abc_52155_new_n13248_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13249_));
AND2X2 AND2X2_5833 ( .A(u2__abc_52155_new_n13249_), .B(u2__abc_52155_new_n13247_), .Y(u2__abc_52155_new_n13250_));
AND2X2 AND2X2_5834 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_284_), .Y(u2__abc_52155_new_n13251_));
AND2X2 AND2X2_5835 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6302_), .Y(u2__abc_52155_new_n13254_));
AND2X2 AND2X2_5836 ( .A(u2__abc_52155_new_n13255_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13256_));
AND2X2 AND2X2_5837 ( .A(u2__abc_52155_new_n13253_), .B(u2__abc_52155_new_n13256_), .Y(u2__abc_52155_new_n13257_));
AND2X2 AND2X2_5838 ( .A(u2__abc_52155_new_n13258_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__286_));
AND2X2 AND2X2_5839 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_287_), .Y(u2__abc_52155_new_n13260_));
AND2X2 AND2X2_584 ( .A(u2__abc_52155_new_n3104_), .B(sqrto_3_), .Y(u2__abc_52155_new_n3105_));
AND2X2 AND2X2_5840 ( .A(u2__abc_52155_new_n13247_), .B(u2__abc_52155_new_n6382_), .Y(u2__abc_52155_new_n13262_));
AND2X2 AND2X2_5841 ( .A(u2__abc_52155_new_n13265_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13266_));
AND2X2 AND2X2_5842 ( .A(u2__abc_52155_new_n13266_), .B(u2__abc_52155_new_n13263_), .Y(u2__abc_52155_new_n13267_));
AND2X2 AND2X2_5843 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_285_), .Y(u2__abc_52155_new_n13268_));
AND2X2 AND2X2_5844 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6309_), .Y(u2__abc_52155_new_n13271_));
AND2X2 AND2X2_5845 ( .A(u2__abc_52155_new_n13272_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13273_));
AND2X2 AND2X2_5846 ( .A(u2__abc_52155_new_n13270_), .B(u2__abc_52155_new_n13273_), .Y(u2__abc_52155_new_n13274_));
AND2X2 AND2X2_5847 ( .A(u2__abc_52155_new_n13275_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__287_));
AND2X2 AND2X2_5848 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_288_), .Y(u2__abc_52155_new_n13277_));
AND2X2 AND2X2_5849 ( .A(u2__abc_52155_new_n12974_), .B(u2__abc_52155_new_n6475_), .Y(u2__abc_52155_new_n13278_));
AND2X2 AND2X2_585 ( .A(u2__abc_52155_new_n3107_), .B(u2_remHi_2_), .Y(u2__abc_52155_new_n3108_));
AND2X2 AND2X2_5850 ( .A(u2__abc_52155_new_n13130_), .B(u2__abc_52155_new_n6411_), .Y(u2__abc_52155_new_n13280_));
AND2X2 AND2X2_5851 ( .A(u2__abc_52155_new_n13207_), .B(u2__abc_52155_new_n6410_), .Y(u2__abc_52155_new_n13282_));
AND2X2 AND2X2_5852 ( .A(u2__abc_52155_new_n6392_), .B(u2__abc_52155_new_n6381_), .Y(u2__abc_52155_new_n13286_));
AND2X2 AND2X2_5853 ( .A(u2__abc_52155_new_n13285_), .B(u2__abc_52155_new_n13288_), .Y(u2__abc_52155_new_n13289_));
AND2X2 AND2X2_5854 ( .A(u2__abc_52155_new_n13283_), .B(u2__abc_52155_new_n13289_), .Y(u2__abc_52155_new_n13290_));
AND2X2 AND2X2_5855 ( .A(u2__abc_52155_new_n13281_), .B(u2__abc_52155_new_n13290_), .Y(u2__abc_52155_new_n13291_));
AND2X2 AND2X2_5856 ( .A(u2__abc_52155_new_n13279_), .B(u2__abc_52155_new_n13291_), .Y(u2__abc_52155_new_n13292_));
AND2X2 AND2X2_5857 ( .A(u2__abc_52155_new_n12663_), .B(u2__abc_52155_new_n6603_), .Y(u2__abc_52155_new_n13294_));
AND2X2 AND2X2_5858 ( .A(u2__abc_52155_new_n13295_), .B(u2__abc_52155_new_n6305_), .Y(u2__abc_52155_new_n13296_));
AND2X2 AND2X2_5859 ( .A(u2__abc_52155_new_n13298_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13299_));
AND2X2 AND2X2_586 ( .A(u2__abc_52155_new_n3109_), .B(sqrto_2_), .Y(u2__abc_52155_new_n3110_));
AND2X2 AND2X2_5860 ( .A(u2__abc_52155_new_n13299_), .B(u2__abc_52155_new_n13297_), .Y(u2__abc_52155_new_n13300_));
AND2X2 AND2X2_5861 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_286_), .Y(u2__abc_52155_new_n13301_));
AND2X2 AND2X2_5862 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6287_), .Y(u2__abc_52155_new_n13304_));
AND2X2 AND2X2_5863 ( .A(u2__abc_52155_new_n13305_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13306_));
AND2X2 AND2X2_5864 ( .A(u2__abc_52155_new_n13303_), .B(u2__abc_52155_new_n13306_), .Y(u2__abc_52155_new_n13307_));
AND2X2 AND2X2_5865 ( .A(u2__abc_52155_new_n13308_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__288_));
AND2X2 AND2X2_5866 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_289_), .Y(u2__abc_52155_new_n13310_));
AND2X2 AND2X2_5867 ( .A(u2__abc_52155_new_n13297_), .B(u2__abc_52155_new_n6301_), .Y(u2__abc_52155_new_n13311_));
AND2X2 AND2X2_5868 ( .A(u2__abc_52155_new_n13311_), .B(u2__abc_52155_new_n6312_), .Y(u2__abc_52155_new_n13312_));
AND2X2 AND2X2_5869 ( .A(u2__abc_52155_new_n13314_), .B(u2__abc_52155_new_n13313_), .Y(u2__abc_52155_new_n13315_));
AND2X2 AND2X2_587 ( .A(u2__abc_52155_new_n3114_), .B(u2_remHi_0_), .Y(u2__abc_52155_new_n3115_));
AND2X2 AND2X2_5870 ( .A(u2__abc_52155_new_n13316_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13317_));
AND2X2 AND2X2_5871 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_287_), .Y(u2__abc_52155_new_n13318_));
AND2X2 AND2X2_5872 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6294_), .Y(u2__abc_52155_new_n13321_));
AND2X2 AND2X2_5873 ( .A(u2__abc_52155_new_n13322_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13323_));
AND2X2 AND2X2_5874 ( .A(u2__abc_52155_new_n13320_), .B(u2__abc_52155_new_n13323_), .Y(u2__abc_52155_new_n13324_));
AND2X2 AND2X2_5875 ( .A(u2__abc_52155_new_n13325_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__289_));
AND2X2 AND2X2_5876 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_290_), .Y(u2__abc_52155_new_n13327_));
AND2X2 AND2X2_5877 ( .A(u2__abc_52155_new_n6301_), .B(u2__abc_52155_new_n6308_), .Y(u2__abc_52155_new_n13328_));
AND2X2 AND2X2_5878 ( .A(u2__abc_52155_new_n13297_), .B(u2__abc_52155_new_n13328_), .Y(u2__abc_52155_new_n13329_));
AND2X2 AND2X2_5879 ( .A(u2__abc_52155_new_n13331_), .B(u2__abc_52155_new_n6290_), .Y(u2__abc_52155_new_n13332_));
AND2X2 AND2X2_588 ( .A(u2__abc_52155_new_n3116_), .B(sqrto_0_), .Y(u2__abc_52155_new_n3117_));
AND2X2 AND2X2_5880 ( .A(u2__abc_52155_new_n13334_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13335_));
AND2X2 AND2X2_5881 ( .A(u2__abc_52155_new_n13335_), .B(u2__abc_52155_new_n13333_), .Y(u2__abc_52155_new_n13336_));
AND2X2 AND2X2_5882 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_288_), .Y(u2__abc_52155_new_n13337_));
AND2X2 AND2X2_5883 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6333_), .Y(u2__abc_52155_new_n13340_));
AND2X2 AND2X2_5884 ( .A(u2__abc_52155_new_n13341_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13342_));
AND2X2 AND2X2_5885 ( .A(u2__abc_52155_new_n13339_), .B(u2__abc_52155_new_n13342_), .Y(u2__abc_52155_new_n13343_));
AND2X2 AND2X2_5886 ( .A(u2__abc_52155_new_n13344_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__290_));
AND2X2 AND2X2_5887 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_291_), .Y(u2__abc_52155_new_n13346_));
AND2X2 AND2X2_5888 ( .A(u2__abc_52155_new_n13333_), .B(u2__abc_52155_new_n6286_), .Y(u2__abc_52155_new_n13348_));
AND2X2 AND2X2_5889 ( .A(u2__abc_52155_new_n13351_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13352_));
AND2X2 AND2X2_589 ( .A(u2__abc_52155_new_n3119_), .B(sqrto_1_), .Y(u2__abc_52155_new_n3120_));
AND2X2 AND2X2_5890 ( .A(u2__abc_52155_new_n13352_), .B(u2__abc_52155_new_n13349_), .Y(u2__abc_52155_new_n13353_));
AND2X2 AND2X2_5891 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_289_), .Y(u2__abc_52155_new_n13354_));
AND2X2 AND2X2_5892 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6340_), .Y(u2__abc_52155_new_n13357_));
AND2X2 AND2X2_5893 ( .A(u2__abc_52155_new_n13358_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13359_));
AND2X2 AND2X2_5894 ( .A(u2__abc_52155_new_n13356_), .B(u2__abc_52155_new_n13359_), .Y(u2__abc_52155_new_n13360_));
AND2X2 AND2X2_5895 ( .A(u2__abc_52155_new_n13361_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__291_));
AND2X2 AND2X2_5896 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_292_), .Y(u2__abc_52155_new_n13363_));
AND2X2 AND2X2_5897 ( .A(u2__abc_52155_new_n6296_), .B(u2__abc_52155_new_n6285_), .Y(u2__abc_52155_new_n13366_));
AND2X2 AND2X2_5898 ( .A(u2__abc_52155_new_n13365_), .B(u2__abc_52155_new_n13368_), .Y(u2__abc_52155_new_n13369_));
AND2X2 AND2X2_5899 ( .A(u2__abc_52155_new_n13295_), .B(u2__abc_52155_new_n6314_), .Y(u2__abc_52155_new_n13371_));
AND2X2 AND2X2_59 ( .A(_abc_73687_new_n753_), .B(sqrto_58_), .Y(\o[94] ));
AND2X2 AND2X2_590 ( .A(u2__abc_52155_new_n3121_), .B(u2_remHi_1_), .Y(u2__abc_52155_new_n3122_));
AND2X2 AND2X2_5900 ( .A(u2__abc_52155_new_n13372_), .B(u2__abc_52155_new_n6336_), .Y(u2__abc_52155_new_n13373_));
AND2X2 AND2X2_5901 ( .A(u2__abc_52155_new_n13375_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13376_));
AND2X2 AND2X2_5902 ( .A(u2__abc_52155_new_n13376_), .B(u2__abc_52155_new_n13374_), .Y(u2__abc_52155_new_n13377_));
AND2X2 AND2X2_5903 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_290_), .Y(u2__abc_52155_new_n13378_));
AND2X2 AND2X2_5904 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6318_), .Y(u2__abc_52155_new_n13381_));
AND2X2 AND2X2_5905 ( .A(u2__abc_52155_new_n13382_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13383_));
AND2X2 AND2X2_5906 ( .A(u2__abc_52155_new_n13380_), .B(u2__abc_52155_new_n13383_), .Y(u2__abc_52155_new_n13384_));
AND2X2 AND2X2_5907 ( .A(u2__abc_52155_new_n13385_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__292_));
AND2X2 AND2X2_5908 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_293_), .Y(u2__abc_52155_new_n13387_));
AND2X2 AND2X2_5909 ( .A(u2__abc_52155_new_n13374_), .B(u2__abc_52155_new_n6332_), .Y(u2__abc_52155_new_n13388_));
AND2X2 AND2X2_591 ( .A(u2__abc_52155_new_n3125_), .B(u2_remHiShift_1_), .Y(u2__abc_52155_new_n3126_));
AND2X2 AND2X2_5910 ( .A(u2__abc_52155_new_n13388_), .B(u2__abc_52155_new_n6343_), .Y(u2__abc_52155_new_n13389_));
AND2X2 AND2X2_5911 ( .A(u2__abc_52155_new_n13391_), .B(u2__abc_52155_new_n13390_), .Y(u2__abc_52155_new_n13392_));
AND2X2 AND2X2_5912 ( .A(u2__abc_52155_new_n13393_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13394_));
AND2X2 AND2X2_5913 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_291_), .Y(u2__abc_52155_new_n13395_));
AND2X2 AND2X2_5914 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6325_), .Y(u2__abc_52155_new_n13398_));
AND2X2 AND2X2_5915 ( .A(u2__abc_52155_new_n13399_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13400_));
AND2X2 AND2X2_5916 ( .A(u2__abc_52155_new_n13397_), .B(u2__abc_52155_new_n13400_), .Y(u2__abc_52155_new_n13401_));
AND2X2 AND2X2_5917 ( .A(u2__abc_52155_new_n13402_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__293_));
AND2X2 AND2X2_5918 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_294_), .Y(u2__abc_52155_new_n13404_));
AND2X2 AND2X2_5919 ( .A(u2__abc_52155_new_n6332_), .B(u2__abc_52155_new_n6339_), .Y(u2__abc_52155_new_n13405_));
AND2X2 AND2X2_592 ( .A(u2__abc_52155_new_n3130_), .B(u2__abc_52155_new_n3128_), .Y(u2__abc_52155_new_n3131_));
AND2X2 AND2X2_5920 ( .A(u2__abc_52155_new_n13374_), .B(u2__abc_52155_new_n13405_), .Y(u2__abc_52155_new_n13406_));
AND2X2 AND2X2_5921 ( .A(u2__abc_52155_new_n13408_), .B(u2__abc_52155_new_n6321_), .Y(u2__abc_52155_new_n13409_));
AND2X2 AND2X2_5922 ( .A(u2__abc_52155_new_n13411_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13412_));
AND2X2 AND2X2_5923 ( .A(u2__abc_52155_new_n13412_), .B(u2__abc_52155_new_n13410_), .Y(u2__abc_52155_new_n13413_));
AND2X2 AND2X2_5924 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_292_), .Y(u2__abc_52155_new_n13414_));
AND2X2 AND2X2_5925 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6221_), .Y(u2__abc_52155_new_n13417_));
AND2X2 AND2X2_5926 ( .A(u2__abc_52155_new_n13418_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13419_));
AND2X2 AND2X2_5927 ( .A(u2__abc_52155_new_n13416_), .B(u2__abc_52155_new_n13419_), .Y(u2__abc_52155_new_n13420_));
AND2X2 AND2X2_5928 ( .A(u2__abc_52155_new_n13421_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__294_));
AND2X2 AND2X2_5929 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_295_), .Y(u2__abc_52155_new_n13423_));
AND2X2 AND2X2_593 ( .A(u2__abc_52155_new_n3127_), .B(u2__abc_52155_new_n3131_), .Y(u2__abc_52155_new_n3132_));
AND2X2 AND2X2_5930 ( .A(u2__abc_52155_new_n13410_), .B(u2__abc_52155_new_n6317_), .Y(u2__abc_52155_new_n13425_));
AND2X2 AND2X2_5931 ( .A(u2__abc_52155_new_n13428_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13429_));
AND2X2 AND2X2_5932 ( .A(u2__abc_52155_new_n13429_), .B(u2__abc_52155_new_n13426_), .Y(u2__abc_52155_new_n13430_));
AND2X2 AND2X2_5933 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_293_), .Y(u2__abc_52155_new_n13431_));
AND2X2 AND2X2_5934 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6228_), .Y(u2__abc_52155_new_n13434_));
AND2X2 AND2X2_5935 ( .A(u2__abc_52155_new_n13435_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13436_));
AND2X2 AND2X2_5936 ( .A(u2__abc_52155_new_n13433_), .B(u2__abc_52155_new_n13436_), .Y(u2__abc_52155_new_n13437_));
AND2X2 AND2X2_5937 ( .A(u2__abc_52155_new_n13438_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__295_));
AND2X2 AND2X2_5938 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_296_), .Y(u2__abc_52155_new_n13440_));
AND2X2 AND2X2_5939 ( .A(u2__abc_52155_new_n13370_), .B(u2__abc_52155_new_n6345_), .Y(u2__abc_52155_new_n13441_));
AND2X2 AND2X2_594 ( .A(u2__abc_52155_new_n3136_), .B(u2__abc_52155_new_n3134_), .Y(u2__abc_52155_new_n3137_));
AND2X2 AND2X2_5940 ( .A(u2__abc_52155_new_n6317_), .B(u2__abc_52155_new_n6324_), .Y(u2__abc_52155_new_n13445_));
AND2X2 AND2X2_5941 ( .A(u2__abc_52155_new_n13444_), .B(u2__abc_52155_new_n13446_), .Y(u2__abc_52155_new_n13447_));
AND2X2 AND2X2_5942 ( .A(u2__abc_52155_new_n13442_), .B(u2__abc_52155_new_n13447_), .Y(u2__abc_52155_new_n13448_));
AND2X2 AND2X2_5943 ( .A(u2__abc_52155_new_n13295_), .B(u2__abc_52155_new_n6346_), .Y(u2__abc_52155_new_n13450_));
AND2X2 AND2X2_5944 ( .A(u2__abc_52155_new_n13451_), .B(u2__abc_52155_new_n6227_), .Y(u2__abc_52155_new_n13452_));
AND2X2 AND2X2_5945 ( .A(u2__abc_52155_new_n13454_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13455_));
AND2X2 AND2X2_5946 ( .A(u2__abc_52155_new_n13455_), .B(u2__abc_52155_new_n13453_), .Y(u2__abc_52155_new_n13456_));
AND2X2 AND2X2_5947 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_294_), .Y(u2__abc_52155_new_n13457_));
AND2X2 AND2X2_5948 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6239_), .Y(u2__abc_52155_new_n13460_));
AND2X2 AND2X2_5949 ( .A(u2__abc_52155_new_n13461_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13462_));
AND2X2 AND2X2_595 ( .A(u2__abc_52155_new_n3141_), .B(u2__abc_52155_new_n3139_), .Y(u2__abc_52155_new_n3142_));
AND2X2 AND2X2_5950 ( .A(u2__abc_52155_new_n13459_), .B(u2__abc_52155_new_n13462_), .Y(u2__abc_52155_new_n13463_));
AND2X2 AND2X2_5951 ( .A(u2__abc_52155_new_n13464_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__296_));
AND2X2 AND2X2_5952 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_297_), .Y(u2__abc_52155_new_n13466_));
AND2X2 AND2X2_5953 ( .A(u2__abc_52155_new_n13453_), .B(u2__abc_52155_new_n6226_), .Y(u2__abc_52155_new_n13468_));
AND2X2 AND2X2_5954 ( .A(u2__abc_52155_new_n13471_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13472_));
AND2X2 AND2X2_5955 ( .A(u2__abc_52155_new_n13472_), .B(u2__abc_52155_new_n13469_), .Y(u2__abc_52155_new_n13473_));
AND2X2 AND2X2_5956 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_295_), .Y(u2__abc_52155_new_n13474_));
AND2X2 AND2X2_5957 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6246_), .Y(u2__abc_52155_new_n13477_));
AND2X2 AND2X2_5958 ( .A(u2__abc_52155_new_n13478_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13479_));
AND2X2 AND2X2_5959 ( .A(u2__abc_52155_new_n13476_), .B(u2__abc_52155_new_n13479_), .Y(u2__abc_52155_new_n13480_));
AND2X2 AND2X2_596 ( .A(u2__abc_52155_new_n3138_), .B(u2__abc_52155_new_n3142_), .Y(u2__abc_52155_new_n3143_));
AND2X2 AND2X2_5960 ( .A(u2__abc_52155_new_n13481_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__297_));
AND2X2 AND2X2_5961 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_298_), .Y(u2__abc_52155_new_n13483_));
AND2X2 AND2X2_5962 ( .A(u2__abc_52155_new_n6226_), .B(u2__abc_52155_new_n6233_), .Y(u2__abc_52155_new_n13484_));
AND2X2 AND2X2_5963 ( .A(u2__abc_52155_new_n13451_), .B(u2__abc_52155_new_n6235_), .Y(u2__abc_52155_new_n13487_));
AND2X2 AND2X2_5964 ( .A(u2__abc_52155_new_n13488_), .B(u2__abc_52155_new_n6242_), .Y(u2__abc_52155_new_n13489_));
AND2X2 AND2X2_5965 ( .A(u2__abc_52155_new_n13491_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13492_));
AND2X2 AND2X2_5966 ( .A(u2__abc_52155_new_n13492_), .B(u2__abc_52155_new_n13490_), .Y(u2__abc_52155_new_n13493_));
AND2X2 AND2X2_5967 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_296_), .Y(u2__abc_52155_new_n13494_));
AND2X2 AND2X2_5968 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6270_), .Y(u2__abc_52155_new_n13497_));
AND2X2 AND2X2_5969 ( .A(u2__abc_52155_new_n13498_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13499_));
AND2X2 AND2X2_597 ( .A(u2__abc_52155_new_n3133_), .B(u2__abc_52155_new_n3143_), .Y(u2__abc_52155_new_n3144_));
AND2X2 AND2X2_5970 ( .A(u2__abc_52155_new_n13496_), .B(u2__abc_52155_new_n13499_), .Y(u2__abc_52155_new_n13500_));
AND2X2 AND2X2_5971 ( .A(u2__abc_52155_new_n13501_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__298_));
AND2X2 AND2X2_5972 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_299_), .Y(u2__abc_52155_new_n13503_));
AND2X2 AND2X2_5973 ( .A(u2__abc_52155_new_n13490_), .B(u2__abc_52155_new_n6238_), .Y(u2__abc_52155_new_n13505_));
AND2X2 AND2X2_5974 ( .A(u2__abc_52155_new_n13508_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13509_));
AND2X2 AND2X2_5975 ( .A(u2__abc_52155_new_n13509_), .B(u2__abc_52155_new_n13506_), .Y(u2__abc_52155_new_n13510_));
AND2X2 AND2X2_5976 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_297_), .Y(u2__abc_52155_new_n13511_));
AND2X2 AND2X2_5977 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6277_), .Y(u2__abc_52155_new_n13514_));
AND2X2 AND2X2_5978 ( .A(u2__abc_52155_new_n13515_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13516_));
AND2X2 AND2X2_5979 ( .A(u2__abc_52155_new_n13513_), .B(u2__abc_52155_new_n13516_), .Y(u2__abc_52155_new_n13517_));
AND2X2 AND2X2_598 ( .A(u2__abc_52155_new_n3148_), .B(u2__abc_52155_new_n3080_), .Y(u2__abc_52155_new_n3149_));
AND2X2 AND2X2_5980 ( .A(u2__abc_52155_new_n13518_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__299_));
AND2X2 AND2X2_5981 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_300_), .Y(u2__abc_52155_new_n13520_));
AND2X2 AND2X2_5982 ( .A(u2__abc_52155_new_n13486_), .B(u2__abc_52155_new_n6250_), .Y(u2__abc_52155_new_n13521_));
AND2X2 AND2X2_5983 ( .A(u2__abc_52155_new_n6248_), .B(u2__abc_52155_new_n6237_), .Y(u2__abc_52155_new_n13522_));
AND2X2 AND2X2_5984 ( .A(u2__abc_52155_new_n13451_), .B(u2__abc_52155_new_n6251_), .Y(u2__abc_52155_new_n13525_));
AND2X2 AND2X2_5985 ( .A(u2__abc_52155_new_n13526_), .B(u2__abc_52155_new_n6273_), .Y(u2__abc_52155_new_n13527_));
AND2X2 AND2X2_5986 ( .A(u2__abc_52155_new_n13529_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13530_));
AND2X2 AND2X2_5987 ( .A(u2__abc_52155_new_n13530_), .B(u2__abc_52155_new_n13528_), .Y(u2__abc_52155_new_n13531_));
AND2X2 AND2X2_5988 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_298_), .Y(u2__abc_52155_new_n13532_));
AND2X2 AND2X2_5989 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6255_), .Y(u2__abc_52155_new_n13535_));
AND2X2 AND2X2_599 ( .A(u2__abc_52155_new_n3071_), .B(u2__abc_52155_new_n3066_), .Y(u2__abc_52155_new_n3151_));
AND2X2 AND2X2_5990 ( .A(u2__abc_52155_new_n13536_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13537_));
AND2X2 AND2X2_5991 ( .A(u2__abc_52155_new_n13534_), .B(u2__abc_52155_new_n13537_), .Y(u2__abc_52155_new_n13538_));
AND2X2 AND2X2_5992 ( .A(u2__abc_52155_new_n13539_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__300_));
AND2X2 AND2X2_5993 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_301_), .Y(u2__abc_52155_new_n13541_));
AND2X2 AND2X2_5994 ( .A(u2__abc_52155_new_n13528_), .B(u2__abc_52155_new_n6269_), .Y(u2__abc_52155_new_n13542_));
AND2X2 AND2X2_5995 ( .A(u2__abc_52155_new_n13542_), .B(u2__abc_52155_new_n6280_), .Y(u2__abc_52155_new_n13543_));
AND2X2 AND2X2_5996 ( .A(u2__abc_52155_new_n13545_), .B(u2__abc_52155_new_n13544_), .Y(u2__abc_52155_new_n13546_));
AND2X2 AND2X2_5997 ( .A(u2__abc_52155_new_n13547_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13548_));
AND2X2 AND2X2_5998 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_299_), .Y(u2__abc_52155_new_n13549_));
AND2X2 AND2X2_5999 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6262_), .Y(u2__abc_52155_new_n13552_));
AND2X2 AND2X2_6 ( .A(_abc_73687_new_n753_), .B(sqrto_5_), .Y(\o[41] ));
AND2X2 AND2X2_60 ( .A(_abc_73687_new_n753_), .B(sqrto_59_), .Y(\o[95] ));
AND2X2 AND2X2_600 ( .A(u2__abc_52155_new_n3152_), .B(u2__abc_52155_new_n3074_), .Y(u2__abc_52155_new_n3153_));
AND2X2 AND2X2_6000 ( .A(u2__abc_52155_new_n13553_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13554_));
AND2X2 AND2X2_6001 ( .A(u2__abc_52155_new_n13551_), .B(u2__abc_52155_new_n13554_), .Y(u2__abc_52155_new_n13555_));
AND2X2 AND2X2_6002 ( .A(u2__abc_52155_new_n13556_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__301_));
AND2X2 AND2X2_6003 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_302_), .Y(u2__abc_52155_new_n13558_));
AND2X2 AND2X2_6004 ( .A(u2__abc_52155_new_n6269_), .B(u2__abc_52155_new_n6276_), .Y(u2__abc_52155_new_n13559_));
AND2X2 AND2X2_6005 ( .A(u2__abc_52155_new_n13528_), .B(u2__abc_52155_new_n13559_), .Y(u2__abc_52155_new_n13560_));
AND2X2 AND2X2_6006 ( .A(u2__abc_52155_new_n13562_), .B(u2__abc_52155_new_n6258_), .Y(u2__abc_52155_new_n13563_));
AND2X2 AND2X2_6007 ( .A(u2__abc_52155_new_n13565_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13566_));
AND2X2 AND2X2_6008 ( .A(u2__abc_52155_new_n13566_), .B(u2__abc_52155_new_n13564_), .Y(u2__abc_52155_new_n13567_));
AND2X2 AND2X2_6009 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_300_), .Y(u2__abc_52155_new_n13568_));
AND2X2 AND2X2_601 ( .A(u2__abc_52155_new_n3150_), .B(u2__abc_52155_new_n3153_), .Y(u2__abc_52155_new_n3154_));
AND2X2 AND2X2_6010 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6157_), .Y(u2__abc_52155_new_n13571_));
AND2X2 AND2X2_6011 ( .A(u2__abc_52155_new_n13572_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13573_));
AND2X2 AND2X2_6012 ( .A(u2__abc_52155_new_n13570_), .B(u2__abc_52155_new_n13573_), .Y(u2__abc_52155_new_n13574_));
AND2X2 AND2X2_6013 ( .A(u2__abc_52155_new_n13575_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__302_));
AND2X2 AND2X2_6014 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_303_), .Y(u2__abc_52155_new_n13577_));
AND2X2 AND2X2_6015 ( .A(u2__abc_52155_new_n13564_), .B(u2__abc_52155_new_n6254_), .Y(u2__abc_52155_new_n13579_));
AND2X2 AND2X2_6016 ( .A(u2__abc_52155_new_n13582_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13583_));
AND2X2 AND2X2_6017 ( .A(u2__abc_52155_new_n13583_), .B(u2__abc_52155_new_n13580_), .Y(u2__abc_52155_new_n13584_));
AND2X2 AND2X2_6018 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_301_), .Y(u2__abc_52155_new_n13585_));
AND2X2 AND2X2_6019 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6164_), .Y(u2__abc_52155_new_n13588_));
AND2X2 AND2X2_602 ( .A(u2__abc_52155_new_n3046_), .B(u2__abc_52155_new_n3038_), .Y(u2__abc_52155_new_n3156_));
AND2X2 AND2X2_6020 ( .A(u2__abc_52155_new_n13589_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13590_));
AND2X2 AND2X2_6021 ( .A(u2__abc_52155_new_n13587_), .B(u2__abc_52155_new_n13590_), .Y(u2__abc_52155_new_n13591_));
AND2X2 AND2X2_6022 ( .A(u2__abc_52155_new_n13592_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__303_));
AND2X2 AND2X2_6023 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_304_), .Y(u2__abc_52155_new_n13594_));
AND2X2 AND2X2_6024 ( .A(u2__abc_52155_new_n13449_), .B(u2__abc_52155_new_n6283_), .Y(u2__abc_52155_new_n13595_));
AND2X2 AND2X2_6025 ( .A(u2__abc_52155_new_n13524_), .B(u2__abc_52155_new_n6282_), .Y(u2__abc_52155_new_n13597_));
AND2X2 AND2X2_6026 ( .A(u2__abc_52155_new_n6264_), .B(u2__abc_52155_new_n6253_), .Y(u2__abc_52155_new_n13601_));
AND2X2 AND2X2_6027 ( .A(u2__abc_52155_new_n13600_), .B(u2__abc_52155_new_n13603_), .Y(u2__abc_52155_new_n13604_));
AND2X2 AND2X2_6028 ( .A(u2__abc_52155_new_n13598_), .B(u2__abc_52155_new_n13604_), .Y(u2__abc_52155_new_n13605_));
AND2X2 AND2X2_6029 ( .A(u2__abc_52155_new_n13596_), .B(u2__abc_52155_new_n13605_), .Y(u2__abc_52155_new_n13606_));
AND2X2 AND2X2_603 ( .A(u2__abc_52155_new_n3050_), .B(u2__abc_52155_new_n3058_), .Y(u2__abc_52155_new_n3160_));
AND2X2 AND2X2_6030 ( .A(u2__abc_52155_new_n13295_), .B(u2__abc_52155_new_n6347_), .Y(u2__abc_52155_new_n13608_));
AND2X2 AND2X2_6031 ( .A(u2__abc_52155_new_n13609_), .B(u2__abc_52155_new_n6163_), .Y(u2__abc_52155_new_n13610_));
AND2X2 AND2X2_6032 ( .A(u2__abc_52155_new_n13612_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13613_));
AND2X2 AND2X2_6033 ( .A(u2__abc_52155_new_n13613_), .B(u2__abc_52155_new_n13611_), .Y(u2__abc_52155_new_n13614_));
AND2X2 AND2X2_6034 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_302_), .Y(u2__abc_52155_new_n13615_));
AND2X2 AND2X2_6035 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6175_), .Y(u2__abc_52155_new_n13618_));
AND2X2 AND2X2_6036 ( .A(u2__abc_52155_new_n13619_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13620_));
AND2X2 AND2X2_6037 ( .A(u2__abc_52155_new_n13617_), .B(u2__abc_52155_new_n13620_), .Y(u2__abc_52155_new_n13621_));
AND2X2 AND2X2_6038 ( .A(u2__abc_52155_new_n13622_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__304_));
AND2X2 AND2X2_6039 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_305_), .Y(u2__abc_52155_new_n13624_));
AND2X2 AND2X2_604 ( .A(u2__abc_52155_new_n3161_), .B(u2__abc_52155_new_n3053_), .Y(u2__abc_52155_new_n3162_));
AND2X2 AND2X2_6040 ( .A(u2__abc_52155_new_n13611_), .B(u2__abc_52155_new_n6162_), .Y(u2__abc_52155_new_n13626_));
AND2X2 AND2X2_6041 ( .A(u2__abc_52155_new_n13629_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13630_));
AND2X2 AND2X2_6042 ( .A(u2__abc_52155_new_n13630_), .B(u2__abc_52155_new_n13627_), .Y(u2__abc_52155_new_n13631_));
AND2X2 AND2X2_6043 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_303_), .Y(u2__abc_52155_new_n13632_));
AND2X2 AND2X2_6044 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6182_), .Y(u2__abc_52155_new_n13635_));
AND2X2 AND2X2_6045 ( .A(u2__abc_52155_new_n13636_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13637_));
AND2X2 AND2X2_6046 ( .A(u2__abc_52155_new_n13634_), .B(u2__abc_52155_new_n13637_), .Y(u2__abc_52155_new_n13638_));
AND2X2 AND2X2_6047 ( .A(u2__abc_52155_new_n13639_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__305_));
AND2X2 AND2X2_6048 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_306_), .Y(u2__abc_52155_new_n13641_));
AND2X2 AND2X2_6049 ( .A(u2__abc_52155_new_n6162_), .B(u2__abc_52155_new_n6169_), .Y(u2__abc_52155_new_n13642_));
AND2X2 AND2X2_605 ( .A(u2__abc_52155_new_n3163_), .B(u2__abc_52155_new_n3158_), .Y(u2__abc_52155_new_n3164_));
AND2X2 AND2X2_6050 ( .A(u2__abc_52155_new_n13609_), .B(u2__abc_52155_new_n6171_), .Y(u2__abc_52155_new_n13645_));
AND2X2 AND2X2_6051 ( .A(u2__abc_52155_new_n13646_), .B(u2__abc_52155_new_n6178_), .Y(u2__abc_52155_new_n13647_));
AND2X2 AND2X2_6052 ( .A(u2__abc_52155_new_n13649_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13650_));
AND2X2 AND2X2_6053 ( .A(u2__abc_52155_new_n13650_), .B(u2__abc_52155_new_n13648_), .Y(u2__abc_52155_new_n13651_));
AND2X2 AND2X2_6054 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_304_), .Y(u2__abc_52155_new_n13652_));
AND2X2 AND2X2_6055 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6213_), .Y(u2__abc_52155_new_n13655_));
AND2X2 AND2X2_6056 ( .A(u2__abc_52155_new_n13656_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13657_));
AND2X2 AND2X2_6057 ( .A(u2__abc_52155_new_n13654_), .B(u2__abc_52155_new_n13657_), .Y(u2__abc_52155_new_n13658_));
AND2X2 AND2X2_6058 ( .A(u2__abc_52155_new_n13659_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__306_));
AND2X2 AND2X2_6059 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_307_), .Y(u2__abc_52155_new_n13661_));
AND2X2 AND2X2_606 ( .A(u2__abc_52155_new_n3155_), .B(u2__abc_52155_new_n3164_), .Y(u2__abc_52155_new_n3165_));
AND2X2 AND2X2_6060 ( .A(u2__abc_52155_new_n13648_), .B(u2__abc_52155_new_n6174_), .Y(u2__abc_52155_new_n13663_));
AND2X2 AND2X2_6061 ( .A(u2__abc_52155_new_n13666_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13667_));
AND2X2 AND2X2_6062 ( .A(u2__abc_52155_new_n13667_), .B(u2__abc_52155_new_n13664_), .Y(u2__abc_52155_new_n13668_));
AND2X2 AND2X2_6063 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_305_), .Y(u2__abc_52155_new_n13669_));
AND2X2 AND2X2_6064 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6206_), .Y(u2__abc_52155_new_n13672_));
AND2X2 AND2X2_6065 ( .A(u2__abc_52155_new_n13673_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13674_));
AND2X2 AND2X2_6066 ( .A(u2__abc_52155_new_n13671_), .B(u2__abc_52155_new_n13674_), .Y(u2__abc_52155_new_n13675_));
AND2X2 AND2X2_6067 ( .A(u2__abc_52155_new_n13676_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__307_));
AND2X2 AND2X2_6068 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_308_), .Y(u2__abc_52155_new_n13678_));
AND2X2 AND2X2_6069 ( .A(u2__abc_52155_new_n13644_), .B(u2__abc_52155_new_n6186_), .Y(u2__abc_52155_new_n13679_));
AND2X2 AND2X2_607 ( .A(u2__abc_52155_new_n3145_), .B(u2__abc_52155_new_n3165_), .Y(u2__abc_52155_new_n3166_));
AND2X2 AND2X2_6070 ( .A(u2__abc_52155_new_n6184_), .B(u2__abc_52155_new_n6173_), .Y(u2__abc_52155_new_n13680_));
AND2X2 AND2X2_6071 ( .A(u2__abc_52155_new_n13609_), .B(u2__abc_52155_new_n6187_), .Y(u2__abc_52155_new_n13683_));
AND2X2 AND2X2_6072 ( .A(u2__abc_52155_new_n13684_), .B(u2__abc_52155_new_n6216_), .Y(u2__abc_52155_new_n13685_));
AND2X2 AND2X2_6073 ( .A(u2__abc_52155_new_n13687_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13688_));
AND2X2 AND2X2_6074 ( .A(u2__abc_52155_new_n13688_), .B(u2__abc_52155_new_n13686_), .Y(u2__abc_52155_new_n13689_));
AND2X2 AND2X2_6075 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_306_), .Y(u2__abc_52155_new_n13690_));
AND2X2 AND2X2_6076 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6191_), .Y(u2__abc_52155_new_n13693_));
AND2X2 AND2X2_6077 ( .A(u2__abc_52155_new_n13694_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13695_));
AND2X2 AND2X2_6078 ( .A(u2__abc_52155_new_n13692_), .B(u2__abc_52155_new_n13695_), .Y(u2__abc_52155_new_n13696_));
AND2X2 AND2X2_6079 ( .A(u2__abc_52155_new_n13697_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__308_));
AND2X2 AND2X2_608 ( .A(u2__abc_52155_new_n3167_), .B(u2_remHi_24_), .Y(u2__abc_52155_new_n3168_));
AND2X2 AND2X2_6080 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_309_), .Y(u2__abc_52155_new_n13699_));
AND2X2 AND2X2_6081 ( .A(u2__abc_52155_new_n13686_), .B(u2__abc_52155_new_n6212_), .Y(u2__abc_52155_new_n13700_));
AND2X2 AND2X2_6082 ( .A(u2__abc_52155_new_n13701_), .B(u2__abc_52155_new_n6209_), .Y(u2__abc_52155_new_n13702_));
AND2X2 AND2X2_6083 ( .A(u2__abc_52155_new_n13704_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13705_));
AND2X2 AND2X2_6084 ( .A(u2__abc_52155_new_n13705_), .B(u2__abc_52155_new_n13703_), .Y(u2__abc_52155_new_n13706_));
AND2X2 AND2X2_6085 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_307_), .Y(u2__abc_52155_new_n13707_));
AND2X2 AND2X2_6086 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6198_), .Y(u2__abc_52155_new_n13710_));
AND2X2 AND2X2_6087 ( .A(u2__abc_52155_new_n13711_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13712_));
AND2X2 AND2X2_6088 ( .A(u2__abc_52155_new_n13709_), .B(u2__abc_52155_new_n13712_), .Y(u2__abc_52155_new_n13713_));
AND2X2 AND2X2_6089 ( .A(u2__abc_52155_new_n13714_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__309_));
AND2X2 AND2X2_609 ( .A(u2__abc_52155_new_n3169_), .B(sqrto_24_), .Y(u2__abc_52155_new_n3170_));
AND2X2 AND2X2_6090 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_310_), .Y(u2__abc_52155_new_n13716_));
AND2X2 AND2X2_6091 ( .A(u2__abc_52155_new_n13703_), .B(u2__abc_52155_new_n6205_), .Y(u2__abc_52155_new_n13717_));
AND2X2 AND2X2_6092 ( .A(u2__abc_52155_new_n13718_), .B(u2__abc_52155_new_n6194_), .Y(u2__abc_52155_new_n13719_));
AND2X2 AND2X2_6093 ( .A(u2__abc_52155_new_n13721_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13722_));
AND2X2 AND2X2_6094 ( .A(u2__abc_52155_new_n13722_), .B(u2__abc_52155_new_n13720_), .Y(u2__abc_52155_new_n13723_));
AND2X2 AND2X2_6095 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_308_), .Y(u2__abc_52155_new_n13724_));
AND2X2 AND2X2_6096 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6112_), .Y(u2__abc_52155_new_n13727_));
AND2X2 AND2X2_6097 ( .A(u2__abc_52155_new_n13728_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13729_));
AND2X2 AND2X2_6098 ( .A(u2__abc_52155_new_n13726_), .B(u2__abc_52155_new_n13729_), .Y(u2__abc_52155_new_n13730_));
AND2X2 AND2X2_6099 ( .A(u2__abc_52155_new_n13731_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__310_));
AND2X2 AND2X2_61 ( .A(_abc_73687_new_n753_), .B(sqrto_60_), .Y(\o[96] ));
AND2X2 AND2X2_610 ( .A(u2__abc_52155_new_n3172_), .B(u2_remHi_25_), .Y(u2__abc_52155_new_n3173_));
AND2X2 AND2X2_6100 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_311_), .Y(u2__abc_52155_new_n13733_));
AND2X2 AND2X2_6101 ( .A(u2__abc_52155_new_n13720_), .B(u2__abc_52155_new_n6190_), .Y(u2__abc_52155_new_n13735_));
AND2X2 AND2X2_6102 ( .A(u2__abc_52155_new_n13738_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13739_));
AND2X2 AND2X2_6103 ( .A(u2__abc_52155_new_n13739_), .B(u2__abc_52155_new_n13736_), .Y(u2__abc_52155_new_n13740_));
AND2X2 AND2X2_6104 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_309_), .Y(u2__abc_52155_new_n13741_));
AND2X2 AND2X2_6105 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6119_), .Y(u2__abc_52155_new_n13744_));
AND2X2 AND2X2_6106 ( .A(u2__abc_52155_new_n13745_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13746_));
AND2X2 AND2X2_6107 ( .A(u2__abc_52155_new_n13743_), .B(u2__abc_52155_new_n13746_), .Y(u2__abc_52155_new_n13747_));
AND2X2 AND2X2_6108 ( .A(u2__abc_52155_new_n13748_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__311_));
AND2X2 AND2X2_6109 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_312_), .Y(u2__abc_52155_new_n13750_));
AND2X2 AND2X2_611 ( .A(u2__abc_52155_new_n3174_), .B(sqrto_25_), .Y(u2__abc_52155_new_n3175_));
AND2X2 AND2X2_6110 ( .A(u2__abc_52155_new_n13682_), .B(u2__abc_52155_new_n6218_), .Y(u2__abc_52155_new_n13751_));
AND2X2 AND2X2_6111 ( .A(u2__abc_52155_new_n6208_), .B(u2__abc_52155_new_n6211_), .Y(u2__abc_52155_new_n13752_));
AND2X2 AND2X2_6112 ( .A(u2__abc_52155_new_n13753_), .B(u2__abc_52155_new_n6202_), .Y(u2__abc_52155_new_n13754_));
AND2X2 AND2X2_6113 ( .A(u2__abc_52155_new_n6200_), .B(u2__abc_52155_new_n6189_), .Y(u2__abc_52155_new_n13755_));
AND2X2 AND2X2_6114 ( .A(u2__abc_52155_new_n13609_), .B(u2__abc_52155_new_n6219_), .Y(u2__abc_52155_new_n13759_));
AND2X2 AND2X2_6115 ( .A(u2__abc_52155_new_n13760_), .B(u2__abc_52155_new_n6115_), .Y(u2__abc_52155_new_n13761_));
AND2X2 AND2X2_6116 ( .A(u2__abc_52155_new_n13763_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13764_));
AND2X2 AND2X2_6117 ( .A(u2__abc_52155_new_n13764_), .B(u2__abc_52155_new_n13762_), .Y(u2__abc_52155_new_n13765_));
AND2X2 AND2X2_6118 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_310_), .Y(u2__abc_52155_new_n13766_));
AND2X2 AND2X2_6119 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6097_), .Y(u2__abc_52155_new_n13769_));
AND2X2 AND2X2_612 ( .A(u2__abc_52155_new_n3179_), .B(u2_remHi_23_), .Y(u2__abc_52155_new_n3180_));
AND2X2 AND2X2_6120 ( .A(u2__abc_52155_new_n13770_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13771_));
AND2X2 AND2X2_6121 ( .A(u2__abc_52155_new_n13768_), .B(u2__abc_52155_new_n13771_), .Y(u2__abc_52155_new_n13772_));
AND2X2 AND2X2_6122 ( .A(u2__abc_52155_new_n13773_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__312_));
AND2X2 AND2X2_6123 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_313_), .Y(u2__abc_52155_new_n13775_));
AND2X2 AND2X2_6124 ( .A(u2__abc_52155_new_n13762_), .B(u2__abc_52155_new_n6111_), .Y(u2__abc_52155_new_n13776_));
AND2X2 AND2X2_6125 ( .A(u2__abc_52155_new_n13776_), .B(u2__abc_52155_new_n6122_), .Y(u2__abc_52155_new_n13777_));
AND2X2 AND2X2_6126 ( .A(u2__abc_52155_new_n13779_), .B(u2__abc_52155_new_n13778_), .Y(u2__abc_52155_new_n13780_));
AND2X2 AND2X2_6127 ( .A(u2__abc_52155_new_n13781_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13782_));
AND2X2 AND2X2_6128 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_311_), .Y(u2__abc_52155_new_n13783_));
AND2X2 AND2X2_6129 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6104_), .Y(u2__abc_52155_new_n13786_));
AND2X2 AND2X2_613 ( .A(u2__abc_52155_new_n3182_), .B(sqrto_23_), .Y(u2__abc_52155_new_n3183_));
AND2X2 AND2X2_6130 ( .A(u2__abc_52155_new_n13787_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13788_));
AND2X2 AND2X2_6131 ( .A(u2__abc_52155_new_n13785_), .B(u2__abc_52155_new_n13788_), .Y(u2__abc_52155_new_n13789_));
AND2X2 AND2X2_6132 ( .A(u2__abc_52155_new_n13790_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__313_));
AND2X2 AND2X2_6133 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_314_), .Y(u2__abc_52155_new_n13792_));
AND2X2 AND2X2_6134 ( .A(u2__abc_52155_new_n6111_), .B(u2__abc_52155_new_n6118_), .Y(u2__abc_52155_new_n13793_));
AND2X2 AND2X2_6135 ( .A(u2__abc_52155_new_n13762_), .B(u2__abc_52155_new_n13793_), .Y(u2__abc_52155_new_n13794_));
AND2X2 AND2X2_6136 ( .A(u2__abc_52155_new_n13796_), .B(u2__abc_52155_new_n6100_), .Y(u2__abc_52155_new_n13797_));
AND2X2 AND2X2_6137 ( .A(u2__abc_52155_new_n13799_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13800_));
AND2X2 AND2X2_6138 ( .A(u2__abc_52155_new_n13800_), .B(u2__abc_52155_new_n13798_), .Y(u2__abc_52155_new_n13801_));
AND2X2 AND2X2_6139 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_312_), .Y(u2__abc_52155_new_n13802_));
AND2X2 AND2X2_614 ( .A(u2__abc_52155_new_n3181_), .B(u2__abc_52155_new_n3184_), .Y(u2__abc_52155_new_n3185_));
AND2X2 AND2X2_6140 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6143_), .Y(u2__abc_52155_new_n13805_));
AND2X2 AND2X2_6141 ( .A(u2__abc_52155_new_n13806_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13807_));
AND2X2 AND2X2_6142 ( .A(u2__abc_52155_new_n13804_), .B(u2__abc_52155_new_n13807_), .Y(u2__abc_52155_new_n13808_));
AND2X2 AND2X2_6143 ( .A(u2__abc_52155_new_n13809_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__314_));
AND2X2 AND2X2_6144 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_315_), .Y(u2__abc_52155_new_n13811_));
AND2X2 AND2X2_6145 ( .A(u2__abc_52155_new_n13798_), .B(u2__abc_52155_new_n6096_), .Y(u2__abc_52155_new_n13813_));
AND2X2 AND2X2_6146 ( .A(u2__abc_52155_new_n13816_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13817_));
AND2X2 AND2X2_6147 ( .A(u2__abc_52155_new_n13817_), .B(u2__abc_52155_new_n13814_), .Y(u2__abc_52155_new_n13818_));
AND2X2 AND2X2_6148 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_313_), .Y(u2__abc_52155_new_n13819_));
AND2X2 AND2X2_6149 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6150_), .Y(u2__abc_52155_new_n13822_));
AND2X2 AND2X2_615 ( .A(u2__abc_52155_new_n3186_), .B(u2_remHi_22_), .Y(u2__abc_52155_new_n3187_));
AND2X2 AND2X2_6150 ( .A(u2__abc_52155_new_n13823_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13824_));
AND2X2 AND2X2_6151 ( .A(u2__abc_52155_new_n13821_), .B(u2__abc_52155_new_n13824_), .Y(u2__abc_52155_new_n13825_));
AND2X2 AND2X2_6152 ( .A(u2__abc_52155_new_n13826_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__315_));
AND2X2 AND2X2_6153 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_316_), .Y(u2__abc_52155_new_n13828_));
AND2X2 AND2X2_6154 ( .A(u2__abc_52155_new_n6106_), .B(u2__abc_52155_new_n6095_), .Y(u2__abc_52155_new_n13832_));
AND2X2 AND2X2_6155 ( .A(u2__abc_52155_new_n13831_), .B(u2__abc_52155_new_n13834_), .Y(u2__abc_52155_new_n13835_));
AND2X2 AND2X2_6156 ( .A(u2__abc_52155_new_n13760_), .B(u2__abc_52155_new_n6124_), .Y(u2__abc_52155_new_n13837_));
AND2X2 AND2X2_6157 ( .A(u2__abc_52155_new_n13838_), .B(u2__abc_52155_new_n6146_), .Y(u2__abc_52155_new_n13839_));
AND2X2 AND2X2_6158 ( .A(u2__abc_52155_new_n13841_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13842_));
AND2X2 AND2X2_6159 ( .A(u2__abc_52155_new_n13842_), .B(u2__abc_52155_new_n13840_), .Y(u2__abc_52155_new_n13843_));
AND2X2 AND2X2_616 ( .A(u2__abc_52155_new_n3189_), .B(sqrto_22_), .Y(u2__abc_52155_new_n3190_));
AND2X2 AND2X2_6160 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_314_), .Y(u2__abc_52155_new_n13844_));
AND2X2 AND2X2_6161 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6128_), .Y(u2__abc_52155_new_n13847_));
AND2X2 AND2X2_6162 ( .A(u2__abc_52155_new_n13848_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13849_));
AND2X2 AND2X2_6163 ( .A(u2__abc_52155_new_n13846_), .B(u2__abc_52155_new_n13849_), .Y(u2__abc_52155_new_n13850_));
AND2X2 AND2X2_6164 ( .A(u2__abc_52155_new_n13851_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__316_));
AND2X2 AND2X2_6165 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_317_), .Y(u2__abc_52155_new_n13853_));
AND2X2 AND2X2_6166 ( .A(u2__abc_52155_new_n13840_), .B(u2__abc_52155_new_n6142_), .Y(u2__abc_52155_new_n13854_));
AND2X2 AND2X2_6167 ( .A(u2__abc_52155_new_n13854_), .B(u2__abc_52155_new_n6153_), .Y(u2__abc_52155_new_n13855_));
AND2X2 AND2X2_6168 ( .A(u2__abc_52155_new_n13857_), .B(u2__abc_52155_new_n13856_), .Y(u2__abc_52155_new_n13858_));
AND2X2 AND2X2_6169 ( .A(u2__abc_52155_new_n13859_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13860_));
AND2X2 AND2X2_617 ( .A(u2__abc_52155_new_n3188_), .B(u2__abc_52155_new_n3191_), .Y(u2__abc_52155_new_n3192_));
AND2X2 AND2X2_6170 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_315_), .Y(u2__abc_52155_new_n13861_));
AND2X2 AND2X2_6171 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6135_), .Y(u2__abc_52155_new_n13864_));
AND2X2 AND2X2_6172 ( .A(u2__abc_52155_new_n13865_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13866_));
AND2X2 AND2X2_6173 ( .A(u2__abc_52155_new_n13863_), .B(u2__abc_52155_new_n13866_), .Y(u2__abc_52155_new_n13867_));
AND2X2 AND2X2_6174 ( .A(u2__abc_52155_new_n13868_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__317_));
AND2X2 AND2X2_6175 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_318_), .Y(u2__abc_52155_new_n13870_));
AND2X2 AND2X2_6176 ( .A(u2__abc_52155_new_n6142_), .B(u2__abc_52155_new_n6149_), .Y(u2__abc_52155_new_n13871_));
AND2X2 AND2X2_6177 ( .A(u2__abc_52155_new_n13840_), .B(u2__abc_52155_new_n13871_), .Y(u2__abc_52155_new_n13872_));
AND2X2 AND2X2_6178 ( .A(u2__abc_52155_new_n13874_), .B(u2__abc_52155_new_n6131_), .Y(u2__abc_52155_new_n13875_));
AND2X2 AND2X2_6179 ( .A(u2__abc_52155_new_n13877_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13878_));
AND2X2 AND2X2_618 ( .A(u2__abc_52155_new_n3185_), .B(u2__abc_52155_new_n3192_), .Y(u2__abc_52155_new_n3193_));
AND2X2 AND2X2_6180 ( .A(u2__abc_52155_new_n13878_), .B(u2__abc_52155_new_n13876_), .Y(u2__abc_52155_new_n13879_));
AND2X2 AND2X2_6181 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_316_), .Y(u2__abc_52155_new_n13880_));
AND2X2 AND2X2_6182 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6059_), .Y(u2__abc_52155_new_n13883_));
AND2X2 AND2X2_6183 ( .A(u2__abc_52155_new_n13884_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13885_));
AND2X2 AND2X2_6184 ( .A(u2__abc_52155_new_n13882_), .B(u2__abc_52155_new_n13885_), .Y(u2__abc_52155_new_n13886_));
AND2X2 AND2X2_6185 ( .A(u2__abc_52155_new_n13887_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__318_));
AND2X2 AND2X2_6186 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_319_), .Y(u2__abc_52155_new_n13889_));
AND2X2 AND2X2_6187 ( .A(u2__abc_52155_new_n13876_), .B(u2__abc_52155_new_n6127_), .Y(u2__abc_52155_new_n13891_));
AND2X2 AND2X2_6188 ( .A(u2__abc_52155_new_n13894_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13895_));
AND2X2 AND2X2_6189 ( .A(u2__abc_52155_new_n13895_), .B(u2__abc_52155_new_n13892_), .Y(u2__abc_52155_new_n13896_));
AND2X2 AND2X2_619 ( .A(u2__abc_52155_new_n3178_), .B(u2__abc_52155_new_n3193_), .Y(u2__abc_52155_new_n3194_));
AND2X2 AND2X2_6190 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_317_), .Y(u2__abc_52155_new_n13897_));
AND2X2 AND2X2_6191 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6066_), .Y(u2__abc_52155_new_n13900_));
AND2X2 AND2X2_6192 ( .A(u2__abc_52155_new_n13901_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13902_));
AND2X2 AND2X2_6193 ( .A(u2__abc_52155_new_n13899_), .B(u2__abc_52155_new_n13902_), .Y(u2__abc_52155_new_n13903_));
AND2X2 AND2X2_6194 ( .A(u2__abc_52155_new_n13904_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__319_));
AND2X2 AND2X2_6195 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_320_), .Y(u2__abc_52155_new_n13906_));
AND2X2 AND2X2_6196 ( .A(u2__abc_52155_new_n13293_), .B(u2__abc_52155_new_n6348_), .Y(u2__abc_52155_new_n13907_));
AND2X2 AND2X2_6197 ( .A(u2__abc_52155_new_n13607_), .B(u2__abc_52155_new_n6220_), .Y(u2__abc_52155_new_n13909_));
AND2X2 AND2X2_6198 ( .A(u2__abc_52155_new_n13758_), .B(u2__abc_52155_new_n6156_), .Y(u2__abc_52155_new_n13911_));
AND2X2 AND2X2_6199 ( .A(u2__abc_52155_new_n13836_), .B(u2__abc_52155_new_n6155_), .Y(u2__abc_52155_new_n13913_));
AND2X2 AND2X2_62 ( .A(_abc_73687_new_n753_), .B(sqrto_61_), .Y(\o[97] ));
AND2X2 AND2X2_620 ( .A(u2__abc_52155_new_n3195_), .B(u2_remHi_28_), .Y(u2__abc_52155_new_n3196_));
AND2X2 AND2X2_6200 ( .A(u2__abc_52155_new_n6137_), .B(u2__abc_52155_new_n6126_), .Y(u2__abc_52155_new_n13918_));
AND2X2 AND2X2_6201 ( .A(u2__abc_52155_new_n13917_), .B(u2__abc_52155_new_n13920_), .Y(u2__abc_52155_new_n13921_));
AND2X2 AND2X2_6202 ( .A(u2__abc_52155_new_n13914_), .B(u2__abc_52155_new_n13921_), .Y(u2__abc_52155_new_n13922_));
AND2X2 AND2X2_6203 ( .A(u2__abc_52155_new_n13912_), .B(u2__abc_52155_new_n13922_), .Y(u2__abc_52155_new_n13923_));
AND2X2 AND2X2_6204 ( .A(u2__abc_52155_new_n13910_), .B(u2__abc_52155_new_n13923_), .Y(u2__abc_52155_new_n13924_));
AND2X2 AND2X2_6205 ( .A(u2__abc_52155_new_n13908_), .B(u2__abc_52155_new_n13924_), .Y(u2__abc_52155_new_n13925_));
AND2X2 AND2X2_6206 ( .A(u2__abc_52155_new_n12663_), .B(u2__abc_52155_new_n6604_), .Y(u2__abc_52155_new_n13927_));
AND2X2 AND2X2_6207 ( .A(u2__abc_52155_new_n13928_), .B(u2__abc_52155_new_n6065_), .Y(u2__abc_52155_new_n13929_));
AND2X2 AND2X2_6208 ( .A(u2__abc_52155_new_n13931_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13932_));
AND2X2 AND2X2_6209 ( .A(u2__abc_52155_new_n13932_), .B(u2__abc_52155_new_n13930_), .Y(u2__abc_52155_new_n13933_));
AND2X2 AND2X2_621 ( .A(u2__abc_52155_new_n3198_), .B(sqrto_28_), .Y(u2__abc_52155_new_n3199_));
AND2X2 AND2X2_6210 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_318_), .Y(u2__abc_52155_new_n13934_));
AND2X2 AND2X2_6211 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6077_), .Y(u2__abc_52155_new_n13937_));
AND2X2 AND2X2_6212 ( .A(u2__abc_52155_new_n13938_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13939_));
AND2X2 AND2X2_6213 ( .A(u2__abc_52155_new_n13936_), .B(u2__abc_52155_new_n13939_), .Y(u2__abc_52155_new_n13940_));
AND2X2 AND2X2_6214 ( .A(u2__abc_52155_new_n13941_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__320_));
AND2X2 AND2X2_6215 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_321_), .Y(u2__abc_52155_new_n13943_));
AND2X2 AND2X2_6216 ( .A(u2__abc_52155_new_n13930_), .B(u2__abc_52155_new_n6064_), .Y(u2__abc_52155_new_n13945_));
AND2X2 AND2X2_6217 ( .A(u2__abc_52155_new_n13948_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13949_));
AND2X2 AND2X2_6218 ( .A(u2__abc_52155_new_n13949_), .B(u2__abc_52155_new_n13946_), .Y(u2__abc_52155_new_n13950_));
AND2X2 AND2X2_6219 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_319_), .Y(u2__abc_52155_new_n13951_));
AND2X2 AND2X2_622 ( .A(u2__abc_52155_new_n3197_), .B(u2__abc_52155_new_n3200_), .Y(u2__abc_52155_new_n3201_));
AND2X2 AND2X2_6220 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6084_), .Y(u2__abc_52155_new_n13954_));
AND2X2 AND2X2_6221 ( .A(u2__abc_52155_new_n13955_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13956_));
AND2X2 AND2X2_6222 ( .A(u2__abc_52155_new_n13953_), .B(u2__abc_52155_new_n13956_), .Y(u2__abc_52155_new_n13957_));
AND2X2 AND2X2_6223 ( .A(u2__abc_52155_new_n13958_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__321_));
AND2X2 AND2X2_6224 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_322_), .Y(u2__abc_52155_new_n13960_));
AND2X2 AND2X2_6225 ( .A(u2__abc_52155_new_n6064_), .B(u2__abc_52155_new_n6071_), .Y(u2__abc_52155_new_n13961_));
AND2X2 AND2X2_6226 ( .A(u2__abc_52155_new_n13928_), .B(u2__abc_52155_new_n6073_), .Y(u2__abc_52155_new_n13964_));
AND2X2 AND2X2_6227 ( .A(u2__abc_52155_new_n13965_), .B(u2__abc_52155_new_n6080_), .Y(u2__abc_52155_new_n13966_));
AND2X2 AND2X2_6228 ( .A(u2__abc_52155_new_n13968_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13969_));
AND2X2 AND2X2_6229 ( .A(u2__abc_52155_new_n13969_), .B(u2__abc_52155_new_n13967_), .Y(u2__abc_52155_new_n13970_));
AND2X2 AND2X2_623 ( .A(u2__abc_52155_new_n3202_), .B(sqrto_29_), .Y(u2__abc_52155_new_n3203_));
AND2X2 AND2X2_6230 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_320_), .Y(u2__abc_52155_new_n13971_));
AND2X2 AND2X2_6231 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6046_), .Y(u2__abc_52155_new_n13974_));
AND2X2 AND2X2_6232 ( .A(u2__abc_52155_new_n13975_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13976_));
AND2X2 AND2X2_6233 ( .A(u2__abc_52155_new_n13973_), .B(u2__abc_52155_new_n13976_), .Y(u2__abc_52155_new_n13977_));
AND2X2 AND2X2_6234 ( .A(u2__abc_52155_new_n13978_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__322_));
AND2X2 AND2X2_6235 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_323_), .Y(u2__abc_52155_new_n13980_));
AND2X2 AND2X2_6236 ( .A(u2__abc_52155_new_n13967_), .B(u2__abc_52155_new_n6076_), .Y(u2__abc_52155_new_n13982_));
AND2X2 AND2X2_6237 ( .A(u2__abc_52155_new_n13985_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n13986_));
AND2X2 AND2X2_6238 ( .A(u2__abc_52155_new_n13986_), .B(u2__abc_52155_new_n13983_), .Y(u2__abc_52155_new_n13987_));
AND2X2 AND2X2_6239 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_321_), .Y(u2__abc_52155_new_n13988_));
AND2X2 AND2X2_624 ( .A(u2__abc_52155_new_n3205_), .B(u2_remHi_29_), .Y(u2__abc_52155_new_n3206_));
AND2X2 AND2X2_6240 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6053_), .Y(u2__abc_52155_new_n13991_));
AND2X2 AND2X2_6241 ( .A(u2__abc_52155_new_n13992_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n13993_));
AND2X2 AND2X2_6242 ( .A(u2__abc_52155_new_n13990_), .B(u2__abc_52155_new_n13993_), .Y(u2__abc_52155_new_n13994_));
AND2X2 AND2X2_6243 ( .A(u2__abc_52155_new_n13995_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__323_));
AND2X2 AND2X2_6244 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_324_), .Y(u2__abc_52155_new_n13997_));
AND2X2 AND2X2_6245 ( .A(u2__abc_52155_new_n13963_), .B(u2__abc_52155_new_n6088_), .Y(u2__abc_52155_new_n13998_));
AND2X2 AND2X2_6246 ( .A(u2__abc_52155_new_n6086_), .B(u2__abc_52155_new_n6075_), .Y(u2__abc_52155_new_n13999_));
AND2X2 AND2X2_6247 ( .A(u2__abc_52155_new_n13928_), .B(u2__abc_52155_new_n6089_), .Y(u2__abc_52155_new_n14002_));
AND2X2 AND2X2_6248 ( .A(u2__abc_52155_new_n14003_), .B(u2__abc_52155_new_n6049_), .Y(u2__abc_52155_new_n14004_));
AND2X2 AND2X2_6249 ( .A(u2__abc_52155_new_n14006_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14007_));
AND2X2 AND2X2_625 ( .A(u2__abc_52155_new_n3204_), .B(u2__abc_52155_new_n3207_), .Y(u2__abc_52155_new_n3208_));
AND2X2 AND2X2_6250 ( .A(u2__abc_52155_new_n14007_), .B(u2__abc_52155_new_n14005_), .Y(u2__abc_52155_new_n14008_));
AND2X2 AND2X2_6251 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_322_), .Y(u2__abc_52155_new_n14009_));
AND2X2 AND2X2_6252 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6028_), .Y(u2__abc_52155_new_n14012_));
AND2X2 AND2X2_6253 ( .A(u2__abc_52155_new_n14013_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14014_));
AND2X2 AND2X2_6254 ( .A(u2__abc_52155_new_n14011_), .B(u2__abc_52155_new_n14014_), .Y(u2__abc_52155_new_n14015_));
AND2X2 AND2X2_6255 ( .A(u2__abc_52155_new_n14016_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__324_));
AND2X2 AND2X2_6256 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_325_), .Y(u2__abc_52155_new_n14018_));
AND2X2 AND2X2_6257 ( .A(u2__abc_52155_new_n14005_), .B(u2__abc_52155_new_n6045_), .Y(u2__abc_52155_new_n14019_));
AND2X2 AND2X2_6258 ( .A(u2__abc_52155_new_n14019_), .B(u2__abc_52155_new_n6056_), .Y(u2__abc_52155_new_n14020_));
AND2X2 AND2X2_6259 ( .A(u2__abc_52155_new_n14022_), .B(u2__abc_52155_new_n14021_), .Y(u2__abc_52155_new_n14023_));
AND2X2 AND2X2_626 ( .A(u2__abc_52155_new_n3201_), .B(u2__abc_52155_new_n3208_), .Y(u2__abc_52155_new_n3209_));
AND2X2 AND2X2_6260 ( .A(u2__abc_52155_new_n14024_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14025_));
AND2X2 AND2X2_6261 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_323_), .Y(u2__abc_52155_new_n14026_));
AND2X2 AND2X2_6262 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6035_), .Y(u2__abc_52155_new_n14029_));
AND2X2 AND2X2_6263 ( .A(u2__abc_52155_new_n14030_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14031_));
AND2X2 AND2X2_6264 ( .A(u2__abc_52155_new_n14028_), .B(u2__abc_52155_new_n14031_), .Y(u2__abc_52155_new_n14032_));
AND2X2 AND2X2_6265 ( .A(u2__abc_52155_new_n14033_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__325_));
AND2X2 AND2X2_6266 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_326_), .Y(u2__abc_52155_new_n14035_));
AND2X2 AND2X2_6267 ( .A(u2__abc_52155_new_n6045_), .B(u2__abc_52155_new_n6052_), .Y(u2__abc_52155_new_n14036_));
AND2X2 AND2X2_6268 ( .A(u2__abc_52155_new_n14005_), .B(u2__abc_52155_new_n14036_), .Y(u2__abc_52155_new_n14037_));
AND2X2 AND2X2_6269 ( .A(u2__abc_52155_new_n14039_), .B(u2__abc_52155_new_n6034_), .Y(u2__abc_52155_new_n14040_));
AND2X2 AND2X2_627 ( .A(u2__abc_52155_new_n3210_), .B(u2_remHi_27_), .Y(u2__abc_52155_new_n3211_));
AND2X2 AND2X2_6270 ( .A(u2__abc_52155_new_n14042_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14043_));
AND2X2 AND2X2_6271 ( .A(u2__abc_52155_new_n14043_), .B(u2__abc_52155_new_n14041_), .Y(u2__abc_52155_new_n14044_));
AND2X2 AND2X2_6272 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_324_), .Y(u2__abc_52155_new_n14045_));
AND2X2 AND2X2_6273 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5965_), .Y(u2__abc_52155_new_n14048_));
AND2X2 AND2X2_6274 ( .A(u2__abc_52155_new_n14049_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14050_));
AND2X2 AND2X2_6275 ( .A(u2__abc_52155_new_n14047_), .B(u2__abc_52155_new_n14050_), .Y(u2__abc_52155_new_n14051_));
AND2X2 AND2X2_6276 ( .A(u2__abc_52155_new_n14052_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__326_));
AND2X2 AND2X2_6277 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_327_), .Y(u2__abc_52155_new_n14054_));
AND2X2 AND2X2_6278 ( .A(u2__abc_52155_new_n14041_), .B(u2__abc_52155_new_n6033_), .Y(u2__abc_52155_new_n14056_));
AND2X2 AND2X2_6279 ( .A(u2__abc_52155_new_n14059_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14060_));
AND2X2 AND2X2_628 ( .A(u2__abc_52155_new_n3213_), .B(sqrto_27_), .Y(u2__abc_52155_new_n3214_));
AND2X2 AND2X2_6280 ( .A(u2__abc_52155_new_n14060_), .B(u2__abc_52155_new_n14057_), .Y(u2__abc_52155_new_n14061_));
AND2X2 AND2X2_6281 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_325_), .Y(u2__abc_52155_new_n14062_));
AND2X2 AND2X2_6282 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5972_), .Y(u2__abc_52155_new_n14065_));
AND2X2 AND2X2_6283 ( .A(u2__abc_52155_new_n14066_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14067_));
AND2X2 AND2X2_6284 ( .A(u2__abc_52155_new_n14064_), .B(u2__abc_52155_new_n14067_), .Y(u2__abc_52155_new_n14068_));
AND2X2 AND2X2_6285 ( .A(u2__abc_52155_new_n14069_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__327_));
AND2X2 AND2X2_6286 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_328_), .Y(u2__abc_52155_new_n14071_));
AND2X2 AND2X2_6287 ( .A(u2__abc_52155_new_n14001_), .B(u2__abc_52155_new_n6058_), .Y(u2__abc_52155_new_n14072_));
AND2X2 AND2X2_6288 ( .A(u2__abc_52155_new_n6033_), .B(u2__abc_52155_new_n6040_), .Y(u2__abc_52155_new_n14076_));
AND2X2 AND2X2_6289 ( .A(u2__abc_52155_new_n14075_), .B(u2__abc_52155_new_n14077_), .Y(u2__abc_52155_new_n14078_));
AND2X2 AND2X2_629 ( .A(u2__abc_52155_new_n3212_), .B(u2__abc_52155_new_n3215_), .Y(u2__abc_52155_new_n3216_));
AND2X2 AND2X2_6290 ( .A(u2__abc_52155_new_n14073_), .B(u2__abc_52155_new_n14078_), .Y(u2__abc_52155_new_n14079_));
AND2X2 AND2X2_6291 ( .A(u2__abc_52155_new_n13928_), .B(u2__abc_52155_new_n6090_), .Y(u2__abc_52155_new_n14081_));
AND2X2 AND2X2_6292 ( .A(u2__abc_52155_new_n14082_), .B(u2__abc_52155_new_n5971_), .Y(u2__abc_52155_new_n14083_));
AND2X2 AND2X2_6293 ( .A(u2__abc_52155_new_n14085_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14086_));
AND2X2 AND2X2_6294 ( .A(u2__abc_52155_new_n14086_), .B(u2__abc_52155_new_n14084_), .Y(u2__abc_52155_new_n14087_));
AND2X2 AND2X2_6295 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_326_), .Y(u2__abc_52155_new_n14088_));
AND2X2 AND2X2_6296 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5983_), .Y(u2__abc_52155_new_n14091_));
AND2X2 AND2X2_6297 ( .A(u2__abc_52155_new_n14092_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14093_));
AND2X2 AND2X2_6298 ( .A(u2__abc_52155_new_n14090_), .B(u2__abc_52155_new_n14093_), .Y(u2__abc_52155_new_n14094_));
AND2X2 AND2X2_6299 ( .A(u2__abc_52155_new_n14095_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__328_));
AND2X2 AND2X2_63 ( .A(_abc_73687_new_n753_), .B(sqrto_62_), .Y(\o[98] ));
AND2X2 AND2X2_630 ( .A(u2__abc_52155_new_n3217_), .B(u2_remHi_26_), .Y(u2__abc_52155_new_n3218_));
AND2X2 AND2X2_6300 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_329_), .Y(u2__abc_52155_new_n14097_));
AND2X2 AND2X2_6301 ( .A(u2__abc_52155_new_n14084_), .B(u2__abc_52155_new_n5970_), .Y(u2__abc_52155_new_n14099_));
AND2X2 AND2X2_6302 ( .A(u2__abc_52155_new_n14102_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14103_));
AND2X2 AND2X2_6303 ( .A(u2__abc_52155_new_n14103_), .B(u2__abc_52155_new_n14100_), .Y(u2__abc_52155_new_n14104_));
AND2X2 AND2X2_6304 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_327_), .Y(u2__abc_52155_new_n14105_));
AND2X2 AND2X2_6305 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5990_), .Y(u2__abc_52155_new_n14108_));
AND2X2 AND2X2_6306 ( .A(u2__abc_52155_new_n14109_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14110_));
AND2X2 AND2X2_6307 ( .A(u2__abc_52155_new_n14107_), .B(u2__abc_52155_new_n14110_), .Y(u2__abc_52155_new_n14111_));
AND2X2 AND2X2_6308 ( .A(u2__abc_52155_new_n14112_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__329_));
AND2X2 AND2X2_6309 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_330_), .Y(u2__abc_52155_new_n14114_));
AND2X2 AND2X2_631 ( .A(u2__abc_52155_new_n3220_), .B(sqrto_26_), .Y(u2__abc_52155_new_n3221_));
AND2X2 AND2X2_6310 ( .A(u2__abc_52155_new_n5970_), .B(u2__abc_52155_new_n5977_), .Y(u2__abc_52155_new_n14115_));
AND2X2 AND2X2_6311 ( .A(u2__abc_52155_new_n14082_), .B(u2__abc_52155_new_n5979_), .Y(u2__abc_52155_new_n14118_));
AND2X2 AND2X2_6312 ( .A(u2__abc_52155_new_n14119_), .B(u2__abc_52155_new_n5986_), .Y(u2__abc_52155_new_n14120_));
AND2X2 AND2X2_6313 ( .A(u2__abc_52155_new_n14122_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14123_));
AND2X2 AND2X2_6314 ( .A(u2__abc_52155_new_n14123_), .B(u2__abc_52155_new_n14121_), .Y(u2__abc_52155_new_n14124_));
AND2X2 AND2X2_6315 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_328_), .Y(u2__abc_52155_new_n14125_));
AND2X2 AND2X2_6316 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6014_), .Y(u2__abc_52155_new_n14128_));
AND2X2 AND2X2_6317 ( .A(u2__abc_52155_new_n14129_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14130_));
AND2X2 AND2X2_6318 ( .A(u2__abc_52155_new_n14127_), .B(u2__abc_52155_new_n14130_), .Y(u2__abc_52155_new_n14131_));
AND2X2 AND2X2_6319 ( .A(u2__abc_52155_new_n14132_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__330_));
AND2X2 AND2X2_632 ( .A(u2__abc_52155_new_n3219_), .B(u2__abc_52155_new_n3222_), .Y(u2__abc_52155_new_n3223_));
AND2X2 AND2X2_6320 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_331_), .Y(u2__abc_52155_new_n14134_));
AND2X2 AND2X2_6321 ( .A(u2__abc_52155_new_n14121_), .B(u2__abc_52155_new_n5982_), .Y(u2__abc_52155_new_n14136_));
AND2X2 AND2X2_6322 ( .A(u2__abc_52155_new_n14139_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14140_));
AND2X2 AND2X2_6323 ( .A(u2__abc_52155_new_n14140_), .B(u2__abc_52155_new_n14137_), .Y(u2__abc_52155_new_n14141_));
AND2X2 AND2X2_6324 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_329_), .Y(u2__abc_52155_new_n14142_));
AND2X2 AND2X2_6325 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6021_), .Y(u2__abc_52155_new_n14145_));
AND2X2 AND2X2_6326 ( .A(u2__abc_52155_new_n14146_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14147_));
AND2X2 AND2X2_6327 ( .A(u2__abc_52155_new_n14144_), .B(u2__abc_52155_new_n14147_), .Y(u2__abc_52155_new_n14148_));
AND2X2 AND2X2_6328 ( .A(u2__abc_52155_new_n14149_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__331_));
AND2X2 AND2X2_6329 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_332_), .Y(u2__abc_52155_new_n14151_));
AND2X2 AND2X2_633 ( .A(u2__abc_52155_new_n3216_), .B(u2__abc_52155_new_n3223_), .Y(u2__abc_52155_new_n3224_));
AND2X2 AND2X2_6330 ( .A(u2__abc_52155_new_n14117_), .B(u2__abc_52155_new_n5994_), .Y(u2__abc_52155_new_n14152_));
AND2X2 AND2X2_6331 ( .A(u2__abc_52155_new_n5992_), .B(u2__abc_52155_new_n5981_), .Y(u2__abc_52155_new_n14153_));
AND2X2 AND2X2_6332 ( .A(u2__abc_52155_new_n14082_), .B(u2__abc_52155_new_n5995_), .Y(u2__abc_52155_new_n14156_));
AND2X2 AND2X2_6333 ( .A(u2__abc_52155_new_n14157_), .B(u2__abc_52155_new_n6017_), .Y(u2__abc_52155_new_n14158_));
AND2X2 AND2X2_6334 ( .A(u2__abc_52155_new_n14160_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14161_));
AND2X2 AND2X2_6335 ( .A(u2__abc_52155_new_n14161_), .B(u2__abc_52155_new_n14159_), .Y(u2__abc_52155_new_n14162_));
AND2X2 AND2X2_6336 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_330_), .Y(u2__abc_52155_new_n14163_));
AND2X2 AND2X2_6337 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5999_), .Y(u2__abc_52155_new_n14166_));
AND2X2 AND2X2_6338 ( .A(u2__abc_52155_new_n14167_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14168_));
AND2X2 AND2X2_6339 ( .A(u2__abc_52155_new_n14165_), .B(u2__abc_52155_new_n14168_), .Y(u2__abc_52155_new_n14169_));
AND2X2 AND2X2_634 ( .A(u2__abc_52155_new_n3209_), .B(u2__abc_52155_new_n3224_), .Y(u2__abc_52155_new_n3225_));
AND2X2 AND2X2_6340 ( .A(u2__abc_52155_new_n14170_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__332_));
AND2X2 AND2X2_6341 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_333_), .Y(u2__abc_52155_new_n14172_));
AND2X2 AND2X2_6342 ( .A(u2__abc_52155_new_n14159_), .B(u2__abc_52155_new_n6013_), .Y(u2__abc_52155_new_n14173_));
AND2X2 AND2X2_6343 ( .A(u2__abc_52155_new_n14173_), .B(u2__abc_52155_new_n6024_), .Y(u2__abc_52155_new_n14174_));
AND2X2 AND2X2_6344 ( .A(u2__abc_52155_new_n14176_), .B(u2__abc_52155_new_n14175_), .Y(u2__abc_52155_new_n14177_));
AND2X2 AND2X2_6345 ( .A(u2__abc_52155_new_n14178_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14179_));
AND2X2 AND2X2_6346 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_331_), .Y(u2__abc_52155_new_n14180_));
AND2X2 AND2X2_6347 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6006_), .Y(u2__abc_52155_new_n14183_));
AND2X2 AND2X2_6348 ( .A(u2__abc_52155_new_n14184_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14185_));
AND2X2 AND2X2_6349 ( .A(u2__abc_52155_new_n14182_), .B(u2__abc_52155_new_n14185_), .Y(u2__abc_52155_new_n14186_));
AND2X2 AND2X2_635 ( .A(u2__abc_52155_new_n3194_), .B(u2__abc_52155_new_n3225_), .Y(u2__abc_52155_new_n3226_));
AND2X2 AND2X2_6350 ( .A(u2__abc_52155_new_n14187_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__333_));
AND2X2 AND2X2_6351 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_334_), .Y(u2__abc_52155_new_n14189_));
AND2X2 AND2X2_6352 ( .A(u2__abc_52155_new_n6013_), .B(u2__abc_52155_new_n6020_), .Y(u2__abc_52155_new_n14190_));
AND2X2 AND2X2_6353 ( .A(u2__abc_52155_new_n14159_), .B(u2__abc_52155_new_n14190_), .Y(u2__abc_52155_new_n14191_));
AND2X2 AND2X2_6354 ( .A(u2__abc_52155_new_n14193_), .B(u2__abc_52155_new_n6002_), .Y(u2__abc_52155_new_n14194_));
AND2X2 AND2X2_6355 ( .A(u2__abc_52155_new_n14196_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14197_));
AND2X2 AND2X2_6356 ( .A(u2__abc_52155_new_n14197_), .B(u2__abc_52155_new_n14195_), .Y(u2__abc_52155_new_n14198_));
AND2X2 AND2X2_6357 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_332_), .Y(u2__abc_52155_new_n14199_));
AND2X2 AND2X2_6358 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5919_), .Y(u2__abc_52155_new_n14202_));
AND2X2 AND2X2_6359 ( .A(u2__abc_52155_new_n14203_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14204_));
AND2X2 AND2X2_636 ( .A(u2__abc_52155_new_n3227_), .B(u2_remHi_16_), .Y(u2__abc_52155_new_n3228_));
AND2X2 AND2X2_6360 ( .A(u2__abc_52155_new_n14201_), .B(u2__abc_52155_new_n14204_), .Y(u2__abc_52155_new_n14205_));
AND2X2 AND2X2_6361 ( .A(u2__abc_52155_new_n14206_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__334_));
AND2X2 AND2X2_6362 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_335_), .Y(u2__abc_52155_new_n14208_));
AND2X2 AND2X2_6363 ( .A(u2__abc_52155_new_n14195_), .B(u2__abc_52155_new_n5998_), .Y(u2__abc_52155_new_n14210_));
AND2X2 AND2X2_6364 ( .A(u2__abc_52155_new_n14213_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14214_));
AND2X2 AND2X2_6365 ( .A(u2__abc_52155_new_n14214_), .B(u2__abc_52155_new_n14211_), .Y(u2__abc_52155_new_n14215_));
AND2X2 AND2X2_6366 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_333_), .Y(u2__abc_52155_new_n14216_));
AND2X2 AND2X2_6367 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5926_), .Y(u2__abc_52155_new_n14219_));
AND2X2 AND2X2_6368 ( .A(u2__abc_52155_new_n14220_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14221_));
AND2X2 AND2X2_6369 ( .A(u2__abc_52155_new_n14218_), .B(u2__abc_52155_new_n14221_), .Y(u2__abc_52155_new_n14222_));
AND2X2 AND2X2_637 ( .A(u2__abc_52155_new_n3229_), .B(sqrto_16_), .Y(u2__abc_52155_new_n3230_));
AND2X2 AND2X2_6370 ( .A(u2__abc_52155_new_n14223_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__335_));
AND2X2 AND2X2_6371 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_336_), .Y(u2__abc_52155_new_n14225_));
AND2X2 AND2X2_6372 ( .A(u2__abc_52155_new_n14080_), .B(u2__abc_52155_new_n6027_), .Y(u2__abc_52155_new_n14226_));
AND2X2 AND2X2_6373 ( .A(u2__abc_52155_new_n14155_), .B(u2__abc_52155_new_n6026_), .Y(u2__abc_52155_new_n14228_));
AND2X2 AND2X2_6374 ( .A(u2__abc_52155_new_n6008_), .B(u2__abc_52155_new_n5997_), .Y(u2__abc_52155_new_n14232_));
AND2X2 AND2X2_6375 ( .A(u2__abc_52155_new_n14231_), .B(u2__abc_52155_new_n14234_), .Y(u2__abc_52155_new_n14235_));
AND2X2 AND2X2_6376 ( .A(u2__abc_52155_new_n14229_), .B(u2__abc_52155_new_n14235_), .Y(u2__abc_52155_new_n14236_));
AND2X2 AND2X2_6377 ( .A(u2__abc_52155_new_n14227_), .B(u2__abc_52155_new_n14236_), .Y(u2__abc_52155_new_n14237_));
AND2X2 AND2X2_6378 ( .A(u2__abc_52155_new_n13928_), .B(u2__abc_52155_new_n6091_), .Y(u2__abc_52155_new_n14239_));
AND2X2 AND2X2_6379 ( .A(u2__abc_52155_new_n14240_), .B(u2__abc_52155_new_n5922_), .Y(u2__abc_52155_new_n14241_));
AND2X2 AND2X2_638 ( .A(u2__abc_52155_new_n3232_), .B(u2_remHi_17_), .Y(u2__abc_52155_new_n3233_));
AND2X2 AND2X2_6380 ( .A(u2__abc_52155_new_n14243_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14244_));
AND2X2 AND2X2_6381 ( .A(u2__abc_52155_new_n14244_), .B(u2__abc_52155_new_n14242_), .Y(u2__abc_52155_new_n14245_));
AND2X2 AND2X2_6382 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_334_), .Y(u2__abc_52155_new_n14246_));
AND2X2 AND2X2_6383 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5904_), .Y(u2__abc_52155_new_n14249_));
AND2X2 AND2X2_6384 ( .A(u2__abc_52155_new_n14250_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14251_));
AND2X2 AND2X2_6385 ( .A(u2__abc_52155_new_n14248_), .B(u2__abc_52155_new_n14251_), .Y(u2__abc_52155_new_n14252_));
AND2X2 AND2X2_6386 ( .A(u2__abc_52155_new_n14253_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__336_));
AND2X2 AND2X2_6387 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_337_), .Y(u2__abc_52155_new_n14255_));
AND2X2 AND2X2_6388 ( .A(u2__abc_52155_new_n14242_), .B(u2__abc_52155_new_n5918_), .Y(u2__abc_52155_new_n14256_));
AND2X2 AND2X2_6389 ( .A(u2__abc_52155_new_n14256_), .B(u2__abc_52155_new_n5929_), .Y(u2__abc_52155_new_n14257_));
AND2X2 AND2X2_639 ( .A(u2__abc_52155_new_n3234_), .B(sqrto_17_), .Y(u2__abc_52155_new_n3235_));
AND2X2 AND2X2_6390 ( .A(u2__abc_52155_new_n14259_), .B(u2__abc_52155_new_n14258_), .Y(u2__abc_52155_new_n14260_));
AND2X2 AND2X2_6391 ( .A(u2__abc_52155_new_n14261_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14262_));
AND2X2 AND2X2_6392 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_335_), .Y(u2__abc_52155_new_n14263_));
AND2X2 AND2X2_6393 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5911_), .Y(u2__abc_52155_new_n14266_));
AND2X2 AND2X2_6394 ( .A(u2__abc_52155_new_n14267_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14268_));
AND2X2 AND2X2_6395 ( .A(u2__abc_52155_new_n14265_), .B(u2__abc_52155_new_n14268_), .Y(u2__abc_52155_new_n14269_));
AND2X2 AND2X2_6396 ( .A(u2__abc_52155_new_n14270_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__337_));
AND2X2 AND2X2_6397 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_338_), .Y(u2__abc_52155_new_n14272_));
AND2X2 AND2X2_6398 ( .A(u2__abc_52155_new_n5918_), .B(u2__abc_52155_new_n5925_), .Y(u2__abc_52155_new_n14273_));
AND2X2 AND2X2_6399 ( .A(u2__abc_52155_new_n14242_), .B(u2__abc_52155_new_n14273_), .Y(u2__abc_52155_new_n14274_));
AND2X2 AND2X2_64 ( .A(_abc_73687_new_n753_), .B(sqrto_63_), .Y(\o[99] ));
AND2X2 AND2X2_640 ( .A(u2__abc_52155_new_n3239_), .B(u2_remHi_14_), .Y(u2__abc_52155_new_n3240_));
AND2X2 AND2X2_6400 ( .A(u2__abc_52155_new_n14276_), .B(u2__abc_52155_new_n5907_), .Y(u2__abc_52155_new_n14277_));
AND2X2 AND2X2_6401 ( .A(u2__abc_52155_new_n14279_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14280_));
AND2X2 AND2X2_6402 ( .A(u2__abc_52155_new_n14280_), .B(u2__abc_52155_new_n14278_), .Y(u2__abc_52155_new_n14281_));
AND2X2 AND2X2_6403 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_336_), .Y(u2__abc_52155_new_n14282_));
AND2X2 AND2X2_6404 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5950_), .Y(u2__abc_52155_new_n14285_));
AND2X2 AND2X2_6405 ( .A(u2__abc_52155_new_n14286_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14287_));
AND2X2 AND2X2_6406 ( .A(u2__abc_52155_new_n14284_), .B(u2__abc_52155_new_n14287_), .Y(u2__abc_52155_new_n14288_));
AND2X2 AND2X2_6407 ( .A(u2__abc_52155_new_n14289_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__338_));
AND2X2 AND2X2_6408 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_339_), .Y(u2__abc_52155_new_n14291_));
AND2X2 AND2X2_6409 ( .A(u2__abc_52155_new_n14278_), .B(u2__abc_52155_new_n5903_), .Y(u2__abc_52155_new_n14293_));
AND2X2 AND2X2_641 ( .A(u2__abc_52155_new_n3241_), .B(u2__abc_52155_new_n3242_), .Y(u2__abc_52155_new_n3243_));
AND2X2 AND2X2_6410 ( .A(u2__abc_52155_new_n14296_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14297_));
AND2X2 AND2X2_6411 ( .A(u2__abc_52155_new_n14297_), .B(u2__abc_52155_new_n14294_), .Y(u2__abc_52155_new_n14298_));
AND2X2 AND2X2_6412 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_337_), .Y(u2__abc_52155_new_n14299_));
AND2X2 AND2X2_6413 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5957_), .Y(u2__abc_52155_new_n14302_));
AND2X2 AND2X2_6414 ( .A(u2__abc_52155_new_n14303_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14304_));
AND2X2 AND2X2_6415 ( .A(u2__abc_52155_new_n14301_), .B(u2__abc_52155_new_n14304_), .Y(u2__abc_52155_new_n14305_));
AND2X2 AND2X2_6416 ( .A(u2__abc_52155_new_n14306_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__339_));
AND2X2 AND2X2_6417 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_340_), .Y(u2__abc_52155_new_n14308_));
AND2X2 AND2X2_6418 ( .A(u2__abc_52155_new_n5913_), .B(u2__abc_52155_new_n5902_), .Y(u2__abc_52155_new_n14311_));
AND2X2 AND2X2_6419 ( .A(u2__abc_52155_new_n14310_), .B(u2__abc_52155_new_n14313_), .Y(u2__abc_52155_new_n14314_));
AND2X2 AND2X2_642 ( .A(u2__abc_52155_new_n3244_), .B(u2_remHi_15_), .Y(u2__abc_52155_new_n3245_));
AND2X2 AND2X2_6420 ( .A(u2__abc_52155_new_n14240_), .B(u2__abc_52155_new_n5931_), .Y(u2__abc_52155_new_n14316_));
AND2X2 AND2X2_6421 ( .A(u2__abc_52155_new_n14317_), .B(u2__abc_52155_new_n5953_), .Y(u2__abc_52155_new_n14318_));
AND2X2 AND2X2_6422 ( .A(u2__abc_52155_new_n14320_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14321_));
AND2X2 AND2X2_6423 ( .A(u2__abc_52155_new_n14321_), .B(u2__abc_52155_new_n14319_), .Y(u2__abc_52155_new_n14322_));
AND2X2 AND2X2_6424 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_338_), .Y(u2__abc_52155_new_n14323_));
AND2X2 AND2X2_6425 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5935_), .Y(u2__abc_52155_new_n14326_));
AND2X2 AND2X2_6426 ( .A(u2__abc_52155_new_n14327_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14328_));
AND2X2 AND2X2_6427 ( .A(u2__abc_52155_new_n14325_), .B(u2__abc_52155_new_n14328_), .Y(u2__abc_52155_new_n14329_));
AND2X2 AND2X2_6428 ( .A(u2__abc_52155_new_n14330_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__340_));
AND2X2 AND2X2_6429 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_341_), .Y(u2__abc_52155_new_n14332_));
AND2X2 AND2X2_643 ( .A(u2__abc_52155_new_n3247_), .B(sqrto_15_), .Y(u2__abc_52155_new_n3248_));
AND2X2 AND2X2_6430 ( .A(u2__abc_52155_new_n14319_), .B(u2__abc_52155_new_n5949_), .Y(u2__abc_52155_new_n14333_));
AND2X2 AND2X2_6431 ( .A(u2__abc_52155_new_n14333_), .B(u2__abc_52155_new_n5960_), .Y(u2__abc_52155_new_n14334_));
AND2X2 AND2X2_6432 ( .A(u2__abc_52155_new_n14336_), .B(u2__abc_52155_new_n14335_), .Y(u2__abc_52155_new_n14337_));
AND2X2 AND2X2_6433 ( .A(u2__abc_52155_new_n14338_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14339_));
AND2X2 AND2X2_6434 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_339_), .Y(u2__abc_52155_new_n14340_));
AND2X2 AND2X2_6435 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5942_), .Y(u2__abc_52155_new_n14343_));
AND2X2 AND2X2_6436 ( .A(u2__abc_52155_new_n14344_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14345_));
AND2X2 AND2X2_6437 ( .A(u2__abc_52155_new_n14342_), .B(u2__abc_52155_new_n14345_), .Y(u2__abc_52155_new_n14346_));
AND2X2 AND2X2_6438 ( .A(u2__abc_52155_new_n14347_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__341_));
AND2X2 AND2X2_6439 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_342_), .Y(u2__abc_52155_new_n14349_));
AND2X2 AND2X2_644 ( .A(u2__abc_52155_new_n3246_), .B(u2__abc_52155_new_n3249_), .Y(u2__abc_52155_new_n3250_));
AND2X2 AND2X2_6440 ( .A(u2__abc_52155_new_n5949_), .B(u2__abc_52155_new_n5956_), .Y(u2__abc_52155_new_n14350_));
AND2X2 AND2X2_6441 ( .A(u2__abc_52155_new_n14319_), .B(u2__abc_52155_new_n14350_), .Y(u2__abc_52155_new_n14351_));
AND2X2 AND2X2_6442 ( .A(u2__abc_52155_new_n14353_), .B(u2__abc_52155_new_n5938_), .Y(u2__abc_52155_new_n14354_));
AND2X2 AND2X2_6443 ( .A(u2__abc_52155_new_n14356_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14357_));
AND2X2 AND2X2_6444 ( .A(u2__abc_52155_new_n14357_), .B(u2__abc_52155_new_n14355_), .Y(u2__abc_52155_new_n14358_));
AND2X2 AND2X2_6445 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_340_), .Y(u2__abc_52155_new_n14359_));
AND2X2 AND2X2_6446 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5856_), .Y(u2__abc_52155_new_n14362_));
AND2X2 AND2X2_6447 ( .A(u2__abc_52155_new_n14363_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14364_));
AND2X2 AND2X2_6448 ( .A(u2__abc_52155_new_n14361_), .B(u2__abc_52155_new_n14364_), .Y(u2__abc_52155_new_n14365_));
AND2X2 AND2X2_6449 ( .A(u2__abc_52155_new_n14366_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__342_));
AND2X2 AND2X2_645 ( .A(u2__abc_52155_new_n3250_), .B(u2__abc_52155_new_n3243_), .Y(u2__abc_52155_new_n3251_));
AND2X2 AND2X2_6450 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_343_), .Y(u2__abc_52155_new_n14368_));
AND2X2 AND2X2_6451 ( .A(u2__abc_52155_new_n14355_), .B(u2__abc_52155_new_n5934_), .Y(u2__abc_52155_new_n14370_));
AND2X2 AND2X2_6452 ( .A(u2__abc_52155_new_n14373_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14374_));
AND2X2 AND2X2_6453 ( .A(u2__abc_52155_new_n14374_), .B(u2__abc_52155_new_n14371_), .Y(u2__abc_52155_new_n14375_));
AND2X2 AND2X2_6454 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_341_), .Y(u2__abc_52155_new_n14376_));
AND2X2 AND2X2_6455 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5863_), .Y(u2__abc_52155_new_n14379_));
AND2X2 AND2X2_6456 ( .A(u2__abc_52155_new_n14380_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14381_));
AND2X2 AND2X2_6457 ( .A(u2__abc_52155_new_n14378_), .B(u2__abc_52155_new_n14381_), .Y(u2__abc_52155_new_n14382_));
AND2X2 AND2X2_6458 ( .A(u2__abc_52155_new_n14383_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__343_));
AND2X2 AND2X2_6459 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_344_), .Y(u2__abc_52155_new_n14385_));
AND2X2 AND2X2_646 ( .A(u2__abc_52155_new_n3238_), .B(u2__abc_52155_new_n3251_), .Y(u2__abc_52155_new_n3252_));
AND2X2 AND2X2_6460 ( .A(u2__abc_52155_new_n14315_), .B(u2__abc_52155_new_n5962_), .Y(u2__abc_52155_new_n14386_));
AND2X2 AND2X2_6461 ( .A(u2__abc_52155_new_n5944_), .B(u2__abc_52155_new_n5933_), .Y(u2__abc_52155_new_n14390_));
AND2X2 AND2X2_6462 ( .A(u2__abc_52155_new_n14389_), .B(u2__abc_52155_new_n14392_), .Y(u2__abc_52155_new_n14393_));
AND2X2 AND2X2_6463 ( .A(u2__abc_52155_new_n14387_), .B(u2__abc_52155_new_n14393_), .Y(u2__abc_52155_new_n14394_));
AND2X2 AND2X2_6464 ( .A(u2__abc_52155_new_n14240_), .B(u2__abc_52155_new_n5963_), .Y(u2__abc_52155_new_n14396_));
AND2X2 AND2X2_6465 ( .A(u2__abc_52155_new_n14397_), .B(u2__abc_52155_new_n5859_), .Y(u2__abc_52155_new_n14398_));
AND2X2 AND2X2_6466 ( .A(u2__abc_52155_new_n14400_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14401_));
AND2X2 AND2X2_6467 ( .A(u2__abc_52155_new_n14401_), .B(u2__abc_52155_new_n14399_), .Y(u2__abc_52155_new_n14402_));
AND2X2 AND2X2_6468 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_342_), .Y(u2__abc_52155_new_n14403_));
AND2X2 AND2X2_6469 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5841_), .Y(u2__abc_52155_new_n14406_));
AND2X2 AND2X2_647 ( .A(u2__abc_52155_new_n3253_), .B(u2_remHi_20_), .Y(u2__abc_52155_new_n3254_));
AND2X2 AND2X2_6470 ( .A(u2__abc_52155_new_n14407_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14408_));
AND2X2 AND2X2_6471 ( .A(u2__abc_52155_new_n14405_), .B(u2__abc_52155_new_n14408_), .Y(u2__abc_52155_new_n14409_));
AND2X2 AND2X2_6472 ( .A(u2__abc_52155_new_n14410_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__344_));
AND2X2 AND2X2_6473 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_345_), .Y(u2__abc_52155_new_n14412_));
AND2X2 AND2X2_6474 ( .A(u2__abc_52155_new_n14399_), .B(u2__abc_52155_new_n5855_), .Y(u2__abc_52155_new_n14413_));
AND2X2 AND2X2_6475 ( .A(u2__abc_52155_new_n14413_), .B(u2__abc_52155_new_n5866_), .Y(u2__abc_52155_new_n14414_));
AND2X2 AND2X2_6476 ( .A(u2__abc_52155_new_n14416_), .B(u2__abc_52155_new_n14415_), .Y(u2__abc_52155_new_n14417_));
AND2X2 AND2X2_6477 ( .A(u2__abc_52155_new_n14418_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14419_));
AND2X2 AND2X2_6478 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_343_), .Y(u2__abc_52155_new_n14420_));
AND2X2 AND2X2_6479 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5848_), .Y(u2__abc_52155_new_n14423_));
AND2X2 AND2X2_648 ( .A(u2__abc_52155_new_n3255_), .B(sqrto_20_), .Y(u2__abc_52155_new_n3256_));
AND2X2 AND2X2_6480 ( .A(u2__abc_52155_new_n14424_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14425_));
AND2X2 AND2X2_6481 ( .A(u2__abc_52155_new_n14422_), .B(u2__abc_52155_new_n14425_), .Y(u2__abc_52155_new_n14426_));
AND2X2 AND2X2_6482 ( .A(u2__abc_52155_new_n14427_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__345_));
AND2X2 AND2X2_6483 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_346_), .Y(u2__abc_52155_new_n14429_));
AND2X2 AND2X2_6484 ( .A(u2__abc_52155_new_n5855_), .B(u2__abc_52155_new_n5862_), .Y(u2__abc_52155_new_n14430_));
AND2X2 AND2X2_6485 ( .A(u2__abc_52155_new_n14399_), .B(u2__abc_52155_new_n14430_), .Y(u2__abc_52155_new_n14431_));
AND2X2 AND2X2_6486 ( .A(u2__abc_52155_new_n14433_), .B(u2__abc_52155_new_n5844_), .Y(u2__abc_52155_new_n14434_));
AND2X2 AND2X2_6487 ( .A(u2__abc_52155_new_n14436_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14437_));
AND2X2 AND2X2_6488 ( .A(u2__abc_52155_new_n14437_), .B(u2__abc_52155_new_n14435_), .Y(u2__abc_52155_new_n14438_));
AND2X2 AND2X2_6489 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_344_), .Y(u2__abc_52155_new_n14439_));
AND2X2 AND2X2_649 ( .A(u2__abc_52155_new_n3258_), .B(u2_remHi_21_), .Y(u2__abc_52155_new_n3259_));
AND2X2 AND2X2_6490 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5887_), .Y(u2__abc_52155_new_n14442_));
AND2X2 AND2X2_6491 ( .A(u2__abc_52155_new_n14443_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14444_));
AND2X2 AND2X2_6492 ( .A(u2__abc_52155_new_n14441_), .B(u2__abc_52155_new_n14444_), .Y(u2__abc_52155_new_n14445_));
AND2X2 AND2X2_6493 ( .A(u2__abc_52155_new_n14446_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__346_));
AND2X2 AND2X2_6494 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_347_), .Y(u2__abc_52155_new_n14448_));
AND2X2 AND2X2_6495 ( .A(u2__abc_52155_new_n14435_), .B(u2__abc_52155_new_n5840_), .Y(u2__abc_52155_new_n14450_));
AND2X2 AND2X2_6496 ( .A(u2__abc_52155_new_n14453_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14454_));
AND2X2 AND2X2_6497 ( .A(u2__abc_52155_new_n14454_), .B(u2__abc_52155_new_n14451_), .Y(u2__abc_52155_new_n14455_));
AND2X2 AND2X2_6498 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_345_), .Y(u2__abc_52155_new_n14456_));
AND2X2 AND2X2_6499 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5894_), .Y(u2__abc_52155_new_n14459_));
AND2X2 AND2X2_65 ( .A(_abc_73687_new_n753_), .B(sqrto_64_), .Y(\o[100] ));
AND2X2 AND2X2_650 ( .A(u2__abc_52155_new_n3260_), .B(sqrto_21_), .Y(u2__abc_52155_new_n3261_));
AND2X2 AND2X2_6500 ( .A(u2__abc_52155_new_n14460_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14461_));
AND2X2 AND2X2_6501 ( .A(u2__abc_52155_new_n14458_), .B(u2__abc_52155_new_n14461_), .Y(u2__abc_52155_new_n14462_));
AND2X2 AND2X2_6502 ( .A(u2__abc_52155_new_n14463_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__347_));
AND2X2 AND2X2_6503 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_348_), .Y(u2__abc_52155_new_n14465_));
AND2X2 AND2X2_6504 ( .A(u2__abc_52155_new_n5850_), .B(u2__abc_52155_new_n5839_), .Y(u2__abc_52155_new_n14468_));
AND2X2 AND2X2_6505 ( .A(u2__abc_52155_new_n14467_), .B(u2__abc_52155_new_n14470_), .Y(u2__abc_52155_new_n14471_));
AND2X2 AND2X2_6506 ( .A(u2__abc_52155_new_n14397_), .B(u2__abc_52155_new_n5868_), .Y(u2__abc_52155_new_n14473_));
AND2X2 AND2X2_6507 ( .A(u2__abc_52155_new_n14474_), .B(u2__abc_52155_new_n5890_), .Y(u2__abc_52155_new_n14475_));
AND2X2 AND2X2_6508 ( .A(u2__abc_52155_new_n14477_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14478_));
AND2X2 AND2X2_6509 ( .A(u2__abc_52155_new_n14478_), .B(u2__abc_52155_new_n14476_), .Y(u2__abc_52155_new_n14479_));
AND2X2 AND2X2_651 ( .A(u2__abc_52155_new_n3264_), .B(u2_remHi_19_), .Y(u2__abc_52155_new_n3265_));
AND2X2 AND2X2_6510 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_346_), .Y(u2__abc_52155_new_n14480_));
AND2X2 AND2X2_6511 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5872_), .Y(u2__abc_52155_new_n14483_));
AND2X2 AND2X2_6512 ( .A(u2__abc_52155_new_n14484_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14485_));
AND2X2 AND2X2_6513 ( .A(u2__abc_52155_new_n14482_), .B(u2__abc_52155_new_n14485_), .Y(u2__abc_52155_new_n14486_));
AND2X2 AND2X2_6514 ( .A(u2__abc_52155_new_n14487_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__348_));
AND2X2 AND2X2_6515 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_349_), .Y(u2__abc_52155_new_n14489_));
AND2X2 AND2X2_6516 ( .A(u2__abc_52155_new_n14476_), .B(u2__abc_52155_new_n5886_), .Y(u2__abc_52155_new_n14490_));
AND2X2 AND2X2_6517 ( .A(u2__abc_52155_new_n14490_), .B(u2__abc_52155_new_n5897_), .Y(u2__abc_52155_new_n14491_));
AND2X2 AND2X2_6518 ( .A(u2__abc_52155_new_n14493_), .B(u2__abc_52155_new_n14492_), .Y(u2__abc_52155_new_n14494_));
AND2X2 AND2X2_6519 ( .A(u2__abc_52155_new_n14495_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14496_));
AND2X2 AND2X2_652 ( .A(u2__abc_52155_new_n3266_), .B(sqrto_19_), .Y(u2__abc_52155_new_n3267_));
AND2X2 AND2X2_6520 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_347_), .Y(u2__abc_52155_new_n14497_));
AND2X2 AND2X2_6521 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5879_), .Y(u2__abc_52155_new_n14500_));
AND2X2 AND2X2_6522 ( .A(u2__abc_52155_new_n14501_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14502_));
AND2X2 AND2X2_6523 ( .A(u2__abc_52155_new_n14499_), .B(u2__abc_52155_new_n14502_), .Y(u2__abc_52155_new_n14503_));
AND2X2 AND2X2_6524 ( .A(u2__abc_52155_new_n14504_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__349_));
AND2X2 AND2X2_6525 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_350_), .Y(u2__abc_52155_new_n14506_));
AND2X2 AND2X2_6526 ( .A(u2__abc_52155_new_n5886_), .B(u2__abc_52155_new_n5893_), .Y(u2__abc_52155_new_n14507_));
AND2X2 AND2X2_6527 ( .A(u2__abc_52155_new_n14476_), .B(u2__abc_52155_new_n14507_), .Y(u2__abc_52155_new_n14508_));
AND2X2 AND2X2_6528 ( .A(u2__abc_52155_new_n14510_), .B(u2__abc_52155_new_n5875_), .Y(u2__abc_52155_new_n14511_));
AND2X2 AND2X2_6529 ( .A(u2__abc_52155_new_n14513_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14514_));
AND2X2 AND2X2_653 ( .A(u2__abc_52155_new_n3269_), .B(u2_remHi_18_), .Y(u2__abc_52155_new_n3270_));
AND2X2 AND2X2_6530 ( .A(u2__abc_52155_new_n14514_), .B(u2__abc_52155_new_n14512_), .Y(u2__abc_52155_new_n14515_));
AND2X2 AND2X2_6531 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_348_), .Y(u2__abc_52155_new_n14516_));
AND2X2 AND2X2_6532 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5791_), .Y(u2__abc_52155_new_n14519_));
AND2X2 AND2X2_6533 ( .A(u2__abc_52155_new_n14520_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14521_));
AND2X2 AND2X2_6534 ( .A(u2__abc_52155_new_n14518_), .B(u2__abc_52155_new_n14521_), .Y(u2__abc_52155_new_n14522_));
AND2X2 AND2X2_6535 ( .A(u2__abc_52155_new_n14523_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__350_));
AND2X2 AND2X2_6536 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_351_), .Y(u2__abc_52155_new_n14525_));
AND2X2 AND2X2_6537 ( .A(u2__abc_52155_new_n14512_), .B(u2__abc_52155_new_n5871_), .Y(u2__abc_52155_new_n14527_));
AND2X2 AND2X2_6538 ( .A(u2__abc_52155_new_n14530_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14531_));
AND2X2 AND2X2_6539 ( .A(u2__abc_52155_new_n14531_), .B(u2__abc_52155_new_n14528_), .Y(u2__abc_52155_new_n14532_));
AND2X2 AND2X2_654 ( .A(u2__abc_52155_new_n3271_), .B(sqrto_18_), .Y(u2__abc_52155_new_n3272_));
AND2X2 AND2X2_6540 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_349_), .Y(u2__abc_52155_new_n14533_));
AND2X2 AND2X2_6541 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5798_), .Y(u2__abc_52155_new_n14536_));
AND2X2 AND2X2_6542 ( .A(u2__abc_52155_new_n14537_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14538_));
AND2X2 AND2X2_6543 ( .A(u2__abc_52155_new_n14535_), .B(u2__abc_52155_new_n14538_), .Y(u2__abc_52155_new_n14539_));
AND2X2 AND2X2_6544 ( .A(u2__abc_52155_new_n14540_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__351_));
AND2X2 AND2X2_6545 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_352_), .Y(u2__abc_52155_new_n14542_));
AND2X2 AND2X2_6546 ( .A(u2__abc_52155_new_n14238_), .B(u2__abc_52155_new_n5964_), .Y(u2__abc_52155_new_n14543_));
AND2X2 AND2X2_6547 ( .A(u2__abc_52155_new_n14395_), .B(u2__abc_52155_new_n5900_), .Y(u2__abc_52155_new_n14545_));
AND2X2 AND2X2_6548 ( .A(u2__abc_52155_new_n14472_), .B(u2__abc_52155_new_n5899_), .Y(u2__abc_52155_new_n14547_));
AND2X2 AND2X2_6549 ( .A(u2__abc_52155_new_n5881_), .B(u2__abc_52155_new_n5870_), .Y(u2__abc_52155_new_n14551_));
AND2X2 AND2X2_655 ( .A(u2__abc_52155_new_n3276_), .B(u2__abc_52155_new_n3252_), .Y(u2__abc_52155_new_n3277_));
AND2X2 AND2X2_6550 ( .A(u2__abc_52155_new_n14550_), .B(u2__abc_52155_new_n14553_), .Y(u2__abc_52155_new_n14554_));
AND2X2 AND2X2_6551 ( .A(u2__abc_52155_new_n14548_), .B(u2__abc_52155_new_n14554_), .Y(u2__abc_52155_new_n14555_));
AND2X2 AND2X2_6552 ( .A(u2__abc_52155_new_n14546_), .B(u2__abc_52155_new_n14555_), .Y(u2__abc_52155_new_n14556_));
AND2X2 AND2X2_6553 ( .A(u2__abc_52155_new_n14544_), .B(u2__abc_52155_new_n14556_), .Y(u2__abc_52155_new_n14557_));
AND2X2 AND2X2_6554 ( .A(u2__abc_52155_new_n13928_), .B(u2__abc_52155_new_n6092_), .Y(u2__abc_52155_new_n14559_));
AND2X2 AND2X2_6555 ( .A(u2__abc_52155_new_n14560_), .B(u2__abc_52155_new_n5794_), .Y(u2__abc_52155_new_n14561_));
AND2X2 AND2X2_6556 ( .A(u2__abc_52155_new_n14563_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14564_));
AND2X2 AND2X2_6557 ( .A(u2__abc_52155_new_n14564_), .B(u2__abc_52155_new_n14562_), .Y(u2__abc_52155_new_n14565_));
AND2X2 AND2X2_6558 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_350_), .Y(u2__abc_52155_new_n14566_));
AND2X2 AND2X2_6559 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5776_), .Y(u2__abc_52155_new_n14569_));
AND2X2 AND2X2_656 ( .A(u2__abc_52155_new_n3277_), .B(u2__abc_52155_new_n3226_), .Y(u2__abc_52155_new_n3278_));
AND2X2 AND2X2_6560 ( .A(u2__abc_52155_new_n14570_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14571_));
AND2X2 AND2X2_6561 ( .A(u2__abc_52155_new_n14568_), .B(u2__abc_52155_new_n14571_), .Y(u2__abc_52155_new_n14572_));
AND2X2 AND2X2_6562 ( .A(u2__abc_52155_new_n14573_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__352_));
AND2X2 AND2X2_6563 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_353_), .Y(u2__abc_52155_new_n14575_));
AND2X2 AND2X2_6564 ( .A(u2__abc_52155_new_n14562_), .B(u2__abc_52155_new_n5790_), .Y(u2__abc_52155_new_n14576_));
AND2X2 AND2X2_6565 ( .A(u2__abc_52155_new_n14576_), .B(u2__abc_52155_new_n5801_), .Y(u2__abc_52155_new_n14577_));
AND2X2 AND2X2_6566 ( .A(u2__abc_52155_new_n14579_), .B(u2__abc_52155_new_n14578_), .Y(u2__abc_52155_new_n14580_));
AND2X2 AND2X2_6567 ( .A(u2__abc_52155_new_n14581_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14582_));
AND2X2 AND2X2_6568 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_351_), .Y(u2__abc_52155_new_n14583_));
AND2X2 AND2X2_6569 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5783_), .Y(u2__abc_52155_new_n14586_));
AND2X2 AND2X2_657 ( .A(u2__abc_52155_new_n3282_), .B(u2__abc_52155_new_n3249_), .Y(u2__abc_52155_new_n3283_));
AND2X2 AND2X2_6570 ( .A(u2__abc_52155_new_n14587_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14588_));
AND2X2 AND2X2_6571 ( .A(u2__abc_52155_new_n14585_), .B(u2__abc_52155_new_n14588_), .Y(u2__abc_52155_new_n14589_));
AND2X2 AND2X2_6572 ( .A(u2__abc_52155_new_n14590_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__353_));
AND2X2 AND2X2_6573 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_354_), .Y(u2__abc_52155_new_n14592_));
AND2X2 AND2X2_6574 ( .A(u2__abc_52155_new_n5790_), .B(u2__abc_52155_new_n5797_), .Y(u2__abc_52155_new_n14593_));
AND2X2 AND2X2_6575 ( .A(u2__abc_52155_new_n14562_), .B(u2__abc_52155_new_n14593_), .Y(u2__abc_52155_new_n14594_));
AND2X2 AND2X2_6576 ( .A(u2__abc_52155_new_n14596_), .B(u2__abc_52155_new_n5779_), .Y(u2__abc_52155_new_n14597_));
AND2X2 AND2X2_6577 ( .A(u2__abc_52155_new_n14599_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14600_));
AND2X2 AND2X2_6578 ( .A(u2__abc_52155_new_n14600_), .B(u2__abc_52155_new_n14598_), .Y(u2__abc_52155_new_n14601_));
AND2X2 AND2X2_6579 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_352_), .Y(u2__abc_52155_new_n14602_));
AND2X2 AND2X2_658 ( .A(u2__abc_52155_new_n3287_), .B(u2__abc_52155_new_n3285_), .Y(u2__abc_52155_new_n3288_));
AND2X2 AND2X2_6580 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5822_), .Y(u2__abc_52155_new_n14605_));
AND2X2 AND2X2_6581 ( .A(u2__abc_52155_new_n14606_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14607_));
AND2X2 AND2X2_6582 ( .A(u2__abc_52155_new_n14604_), .B(u2__abc_52155_new_n14607_), .Y(u2__abc_52155_new_n14608_));
AND2X2 AND2X2_6583 ( .A(u2__abc_52155_new_n14609_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__354_));
AND2X2 AND2X2_6584 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_355_), .Y(u2__abc_52155_new_n14611_));
AND2X2 AND2X2_6585 ( .A(u2__abc_52155_new_n14598_), .B(u2__abc_52155_new_n5775_), .Y(u2__abc_52155_new_n14613_));
AND2X2 AND2X2_6586 ( .A(u2__abc_52155_new_n14616_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14617_));
AND2X2 AND2X2_6587 ( .A(u2__abc_52155_new_n14617_), .B(u2__abc_52155_new_n14614_), .Y(u2__abc_52155_new_n14618_));
AND2X2 AND2X2_6588 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_353_), .Y(u2__abc_52155_new_n14619_));
AND2X2 AND2X2_6589 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5829_), .Y(u2__abc_52155_new_n14622_));
AND2X2 AND2X2_659 ( .A(u2__abc_52155_new_n3284_), .B(u2__abc_52155_new_n3288_), .Y(u2__abc_52155_new_n3289_));
AND2X2 AND2X2_6590 ( .A(u2__abc_52155_new_n14623_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14624_));
AND2X2 AND2X2_6591 ( .A(u2__abc_52155_new_n14621_), .B(u2__abc_52155_new_n14624_), .Y(u2__abc_52155_new_n14625_));
AND2X2 AND2X2_6592 ( .A(u2__abc_52155_new_n14626_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__355_));
AND2X2 AND2X2_6593 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_356_), .Y(u2__abc_52155_new_n14628_));
AND2X2 AND2X2_6594 ( .A(u2__abc_52155_new_n5785_), .B(u2__abc_52155_new_n5774_), .Y(u2__abc_52155_new_n14631_));
AND2X2 AND2X2_6595 ( .A(u2__abc_52155_new_n14630_), .B(u2__abc_52155_new_n14633_), .Y(u2__abc_52155_new_n14634_));
AND2X2 AND2X2_6596 ( .A(u2__abc_52155_new_n14560_), .B(u2__abc_52155_new_n5803_), .Y(u2__abc_52155_new_n14636_));
AND2X2 AND2X2_6597 ( .A(u2__abc_52155_new_n14637_), .B(u2__abc_52155_new_n5825_), .Y(u2__abc_52155_new_n14638_));
AND2X2 AND2X2_6598 ( .A(u2__abc_52155_new_n14640_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14641_));
AND2X2 AND2X2_6599 ( .A(u2__abc_52155_new_n14641_), .B(u2__abc_52155_new_n14639_), .Y(u2__abc_52155_new_n14642_));
AND2X2 AND2X2_66 ( .A(_abc_73687_new_n753_), .B(sqrto_65_), .Y(\o[101] ));
AND2X2 AND2X2_660 ( .A(u2__abc_52155_new_n3293_), .B(u2__abc_52155_new_n3291_), .Y(u2__abc_52155_new_n3294_));
AND2X2 AND2X2_6600 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_354_), .Y(u2__abc_52155_new_n14643_));
AND2X2 AND2X2_6601 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5807_), .Y(u2__abc_52155_new_n14646_));
AND2X2 AND2X2_6602 ( .A(u2__abc_52155_new_n14647_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14648_));
AND2X2 AND2X2_6603 ( .A(u2__abc_52155_new_n14645_), .B(u2__abc_52155_new_n14648_), .Y(u2__abc_52155_new_n14649_));
AND2X2 AND2X2_6604 ( .A(u2__abc_52155_new_n14650_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__356_));
AND2X2 AND2X2_6605 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_357_), .Y(u2__abc_52155_new_n14652_));
AND2X2 AND2X2_6606 ( .A(u2__abc_52155_new_n14639_), .B(u2__abc_52155_new_n5821_), .Y(u2__abc_52155_new_n14653_));
AND2X2 AND2X2_6607 ( .A(u2__abc_52155_new_n14653_), .B(u2__abc_52155_new_n5832_), .Y(u2__abc_52155_new_n14654_));
AND2X2 AND2X2_6608 ( .A(u2__abc_52155_new_n14656_), .B(u2__abc_52155_new_n14655_), .Y(u2__abc_52155_new_n14657_));
AND2X2 AND2X2_6609 ( .A(u2__abc_52155_new_n14658_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14659_));
AND2X2 AND2X2_661 ( .A(u2__abc_52155_new_n3296_), .B(u2__abc_52155_new_n3256_), .Y(u2__abc_52155_new_n3297_));
AND2X2 AND2X2_6610 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_355_), .Y(u2__abc_52155_new_n14660_));
AND2X2 AND2X2_6611 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5814_), .Y(u2__abc_52155_new_n14663_));
AND2X2 AND2X2_6612 ( .A(u2__abc_52155_new_n14664_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14665_));
AND2X2 AND2X2_6613 ( .A(u2__abc_52155_new_n14662_), .B(u2__abc_52155_new_n14665_), .Y(u2__abc_52155_new_n14666_));
AND2X2 AND2X2_6614 ( .A(u2__abc_52155_new_n14667_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__357_));
AND2X2 AND2X2_6615 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_358_), .Y(u2__abc_52155_new_n14669_));
AND2X2 AND2X2_6616 ( .A(u2__abc_52155_new_n5821_), .B(u2__abc_52155_new_n5828_), .Y(u2__abc_52155_new_n14670_));
AND2X2 AND2X2_6617 ( .A(u2__abc_52155_new_n14639_), .B(u2__abc_52155_new_n14670_), .Y(u2__abc_52155_new_n14671_));
AND2X2 AND2X2_6618 ( .A(u2__abc_52155_new_n14673_), .B(u2__abc_52155_new_n5810_), .Y(u2__abc_52155_new_n14674_));
AND2X2 AND2X2_6619 ( .A(u2__abc_52155_new_n14676_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14677_));
AND2X2 AND2X2_662 ( .A(u2__abc_52155_new_n3295_), .B(u2__abc_52155_new_n3299_), .Y(u2__abc_52155_new_n3300_));
AND2X2 AND2X2_6620 ( .A(u2__abc_52155_new_n14677_), .B(u2__abc_52155_new_n14675_), .Y(u2__abc_52155_new_n14678_));
AND2X2 AND2X2_6621 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_356_), .Y(u2__abc_52155_new_n14679_));
AND2X2 AND2X2_6622 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5710_), .Y(u2__abc_52155_new_n14682_));
AND2X2 AND2X2_6623 ( .A(u2__abc_52155_new_n14683_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14684_));
AND2X2 AND2X2_6624 ( .A(u2__abc_52155_new_n14681_), .B(u2__abc_52155_new_n14684_), .Y(u2__abc_52155_new_n14685_));
AND2X2 AND2X2_6625 ( .A(u2__abc_52155_new_n14686_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__358_));
AND2X2 AND2X2_6626 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_359_), .Y(u2__abc_52155_new_n14688_));
AND2X2 AND2X2_6627 ( .A(u2__abc_52155_new_n14675_), .B(u2__abc_52155_new_n5806_), .Y(u2__abc_52155_new_n14690_));
AND2X2 AND2X2_6628 ( .A(u2__abc_52155_new_n14693_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14694_));
AND2X2 AND2X2_6629 ( .A(u2__abc_52155_new_n14694_), .B(u2__abc_52155_new_n14691_), .Y(u2__abc_52155_new_n14695_));
AND2X2 AND2X2_663 ( .A(u2__abc_52155_new_n3290_), .B(u2__abc_52155_new_n3300_), .Y(u2__abc_52155_new_n3301_));
AND2X2 AND2X2_6630 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_357_), .Y(u2__abc_52155_new_n14696_));
AND2X2 AND2X2_6631 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5717_), .Y(u2__abc_52155_new_n14699_));
AND2X2 AND2X2_6632 ( .A(u2__abc_52155_new_n14700_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14701_));
AND2X2 AND2X2_6633 ( .A(u2__abc_52155_new_n14698_), .B(u2__abc_52155_new_n14701_), .Y(u2__abc_52155_new_n14702_));
AND2X2 AND2X2_6634 ( .A(u2__abc_52155_new_n14703_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__359_));
AND2X2 AND2X2_6635 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_360_), .Y(u2__abc_52155_new_n14705_));
AND2X2 AND2X2_6636 ( .A(u2__abc_52155_new_n14635_), .B(u2__abc_52155_new_n5834_), .Y(u2__abc_52155_new_n14706_));
AND2X2 AND2X2_6637 ( .A(u2__abc_52155_new_n5806_), .B(u2__abc_52155_new_n5813_), .Y(u2__abc_52155_new_n14711_));
AND2X2 AND2X2_6638 ( .A(u2__abc_52155_new_n14710_), .B(u2__abc_52155_new_n14712_), .Y(u2__abc_52155_new_n14713_));
AND2X2 AND2X2_6639 ( .A(u2__abc_52155_new_n14707_), .B(u2__abc_52155_new_n14713_), .Y(u2__abc_52155_new_n14714_));
AND2X2 AND2X2_664 ( .A(u2__abc_52155_new_n3304_), .B(u2__abc_52155_new_n3184_), .Y(u2__abc_52155_new_n3305_));
AND2X2 AND2X2_6640 ( .A(u2__abc_52155_new_n14560_), .B(u2__abc_52155_new_n5835_), .Y(u2__abc_52155_new_n14716_));
AND2X2 AND2X2_6641 ( .A(u2__abc_52155_new_n14717_), .B(u2__abc_52155_new_n5716_), .Y(u2__abc_52155_new_n14718_));
AND2X2 AND2X2_6642 ( .A(u2__abc_52155_new_n14720_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14721_));
AND2X2 AND2X2_6643 ( .A(u2__abc_52155_new_n14721_), .B(u2__abc_52155_new_n14719_), .Y(u2__abc_52155_new_n14722_));
AND2X2 AND2X2_6644 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_358_), .Y(u2__abc_52155_new_n14723_));
AND2X2 AND2X2_6645 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5728_), .Y(u2__abc_52155_new_n14726_));
AND2X2 AND2X2_6646 ( .A(u2__abc_52155_new_n14727_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14728_));
AND2X2 AND2X2_6647 ( .A(u2__abc_52155_new_n14725_), .B(u2__abc_52155_new_n14728_), .Y(u2__abc_52155_new_n14729_));
AND2X2 AND2X2_6648 ( .A(u2__abc_52155_new_n14730_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__360_));
AND2X2 AND2X2_6649 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_361_), .Y(u2__abc_52155_new_n14732_));
AND2X2 AND2X2_665 ( .A(u2__abc_52155_new_n3307_), .B(u2__abc_52155_new_n3170_), .Y(u2__abc_52155_new_n3308_));
AND2X2 AND2X2_6650 ( .A(u2__abc_52155_new_n14719_), .B(u2__abc_52155_new_n5715_), .Y(u2__abc_52155_new_n14734_));
AND2X2 AND2X2_6651 ( .A(u2__abc_52155_new_n14737_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14738_));
AND2X2 AND2X2_6652 ( .A(u2__abc_52155_new_n14738_), .B(u2__abc_52155_new_n14735_), .Y(u2__abc_52155_new_n14739_));
AND2X2 AND2X2_6653 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_359_), .Y(u2__abc_52155_new_n14740_));
AND2X2 AND2X2_6654 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5735_), .Y(u2__abc_52155_new_n14743_));
AND2X2 AND2X2_6655 ( .A(u2__abc_52155_new_n14744_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14745_));
AND2X2 AND2X2_6656 ( .A(u2__abc_52155_new_n14742_), .B(u2__abc_52155_new_n14745_), .Y(u2__abc_52155_new_n14746_));
AND2X2 AND2X2_6657 ( .A(u2__abc_52155_new_n14747_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__361_));
AND2X2 AND2X2_6658 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_362_), .Y(u2__abc_52155_new_n14749_));
AND2X2 AND2X2_6659 ( .A(u2__abc_52155_new_n5715_), .B(u2__abc_52155_new_n5722_), .Y(u2__abc_52155_new_n14750_));
AND2X2 AND2X2_666 ( .A(u2__abc_52155_new_n3306_), .B(u2__abc_52155_new_n3310_), .Y(u2__abc_52155_new_n3311_));
AND2X2 AND2X2_6660 ( .A(u2__abc_52155_new_n14717_), .B(u2__abc_52155_new_n5724_), .Y(u2__abc_52155_new_n14753_));
AND2X2 AND2X2_6661 ( .A(u2__abc_52155_new_n14754_), .B(u2__abc_52155_new_n5731_), .Y(u2__abc_52155_new_n14755_));
AND2X2 AND2X2_6662 ( .A(u2__abc_52155_new_n14757_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14758_));
AND2X2 AND2X2_6663 ( .A(u2__abc_52155_new_n14758_), .B(u2__abc_52155_new_n14756_), .Y(u2__abc_52155_new_n14759_));
AND2X2 AND2X2_6664 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_360_), .Y(u2__abc_52155_new_n14760_));
AND2X2 AND2X2_6665 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5759_), .Y(u2__abc_52155_new_n14763_));
AND2X2 AND2X2_6666 ( .A(u2__abc_52155_new_n14764_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14765_));
AND2X2 AND2X2_6667 ( .A(u2__abc_52155_new_n14762_), .B(u2__abc_52155_new_n14765_), .Y(u2__abc_52155_new_n14766_));
AND2X2 AND2X2_6668 ( .A(u2__abc_52155_new_n14767_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__362_));
AND2X2 AND2X2_6669 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_363_), .Y(u2__abc_52155_new_n14769_));
AND2X2 AND2X2_667 ( .A(u2__abc_52155_new_n3207_), .B(u2__abc_52155_new_n3199_), .Y(u2__abc_52155_new_n3313_));
AND2X2 AND2X2_6670 ( .A(u2__abc_52155_new_n14756_), .B(u2__abc_52155_new_n5727_), .Y(u2__abc_52155_new_n14771_));
AND2X2 AND2X2_6671 ( .A(u2__abc_52155_new_n14774_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14775_));
AND2X2 AND2X2_6672 ( .A(u2__abc_52155_new_n14775_), .B(u2__abc_52155_new_n14772_), .Y(u2__abc_52155_new_n14776_));
AND2X2 AND2X2_6673 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_361_), .Y(u2__abc_52155_new_n14777_));
AND2X2 AND2X2_6674 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5766_), .Y(u2__abc_52155_new_n14780_));
AND2X2 AND2X2_6675 ( .A(u2__abc_52155_new_n14781_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14782_));
AND2X2 AND2X2_6676 ( .A(u2__abc_52155_new_n14779_), .B(u2__abc_52155_new_n14782_), .Y(u2__abc_52155_new_n14783_));
AND2X2 AND2X2_6677 ( .A(u2__abc_52155_new_n14784_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__363_));
AND2X2 AND2X2_6678 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_364_), .Y(u2__abc_52155_new_n14786_));
AND2X2 AND2X2_6679 ( .A(u2__abc_52155_new_n14752_), .B(u2__abc_52155_new_n5739_), .Y(u2__abc_52155_new_n14787_));
AND2X2 AND2X2_668 ( .A(u2__abc_52155_new_n3212_), .B(u2__abc_52155_new_n3221_), .Y(u2__abc_52155_new_n3315_));
AND2X2 AND2X2_6680 ( .A(u2__abc_52155_new_n5737_), .B(u2__abc_52155_new_n5726_), .Y(u2__abc_52155_new_n14788_));
AND2X2 AND2X2_6681 ( .A(u2__abc_52155_new_n14717_), .B(u2__abc_52155_new_n5740_), .Y(u2__abc_52155_new_n14791_));
AND2X2 AND2X2_6682 ( .A(u2__abc_52155_new_n14792_), .B(u2__abc_52155_new_n5762_), .Y(u2__abc_52155_new_n14793_));
AND2X2 AND2X2_6683 ( .A(u2__abc_52155_new_n14795_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14796_));
AND2X2 AND2X2_6684 ( .A(u2__abc_52155_new_n14796_), .B(u2__abc_52155_new_n14794_), .Y(u2__abc_52155_new_n14797_));
AND2X2 AND2X2_6685 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_362_), .Y(u2__abc_52155_new_n14798_));
AND2X2 AND2X2_6686 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5744_), .Y(u2__abc_52155_new_n14801_));
AND2X2 AND2X2_6687 ( .A(u2__abc_52155_new_n14802_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14803_));
AND2X2 AND2X2_6688 ( .A(u2__abc_52155_new_n14800_), .B(u2__abc_52155_new_n14803_), .Y(u2__abc_52155_new_n14804_));
AND2X2 AND2X2_6689 ( .A(u2__abc_52155_new_n14805_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__364_));
AND2X2 AND2X2_669 ( .A(u2__abc_52155_new_n3316_), .B(u2__abc_52155_new_n3209_), .Y(u2__abc_52155_new_n3317_));
AND2X2 AND2X2_6690 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_365_), .Y(u2__abc_52155_new_n14807_));
AND2X2 AND2X2_6691 ( .A(u2__abc_52155_new_n14794_), .B(u2__abc_52155_new_n5758_), .Y(u2__abc_52155_new_n14808_));
AND2X2 AND2X2_6692 ( .A(u2__abc_52155_new_n14808_), .B(u2__abc_52155_new_n5769_), .Y(u2__abc_52155_new_n14809_));
AND2X2 AND2X2_6693 ( .A(u2__abc_52155_new_n14811_), .B(u2__abc_52155_new_n14810_), .Y(u2__abc_52155_new_n14812_));
AND2X2 AND2X2_6694 ( .A(u2__abc_52155_new_n14813_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14814_));
AND2X2 AND2X2_6695 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_363_), .Y(u2__abc_52155_new_n14815_));
AND2X2 AND2X2_6696 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5751_), .Y(u2__abc_52155_new_n14818_));
AND2X2 AND2X2_6697 ( .A(u2__abc_52155_new_n14819_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14820_));
AND2X2 AND2X2_6698 ( .A(u2__abc_52155_new_n14817_), .B(u2__abc_52155_new_n14820_), .Y(u2__abc_52155_new_n14821_));
AND2X2 AND2X2_6699 ( .A(u2__abc_52155_new_n14822_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__365_));
AND2X2 AND2X2_67 ( .A(_abc_73687_new_n753_), .B(sqrto_66_), .Y(\o[102] ));
AND2X2 AND2X2_670 ( .A(u2__abc_52155_new_n3312_), .B(u2__abc_52155_new_n3319_), .Y(u2__abc_52155_new_n3320_));
AND2X2 AND2X2_6700 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_366_), .Y(u2__abc_52155_new_n14824_));
AND2X2 AND2X2_6701 ( .A(u2__abc_52155_new_n5758_), .B(u2__abc_52155_new_n5765_), .Y(u2__abc_52155_new_n14825_));
AND2X2 AND2X2_6702 ( .A(u2__abc_52155_new_n14794_), .B(u2__abc_52155_new_n14825_), .Y(u2__abc_52155_new_n14826_));
AND2X2 AND2X2_6703 ( .A(u2__abc_52155_new_n14828_), .B(u2__abc_52155_new_n5747_), .Y(u2__abc_52155_new_n14829_));
AND2X2 AND2X2_6704 ( .A(u2__abc_52155_new_n14831_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14832_));
AND2X2 AND2X2_6705 ( .A(u2__abc_52155_new_n14832_), .B(u2__abc_52155_new_n14830_), .Y(u2__abc_52155_new_n14833_));
AND2X2 AND2X2_6706 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_364_), .Y(u2__abc_52155_new_n14834_));
AND2X2 AND2X2_6707 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5664_), .Y(u2__abc_52155_new_n14837_));
AND2X2 AND2X2_6708 ( .A(u2__abc_52155_new_n14838_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14839_));
AND2X2 AND2X2_6709 ( .A(u2__abc_52155_new_n14836_), .B(u2__abc_52155_new_n14839_), .Y(u2__abc_52155_new_n14840_));
AND2X2 AND2X2_671 ( .A(u2__abc_52155_new_n3302_), .B(u2__abc_52155_new_n3320_), .Y(u2__abc_52155_new_n3321_));
AND2X2 AND2X2_6710 ( .A(u2__abc_52155_new_n14841_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__366_));
AND2X2 AND2X2_6711 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_367_), .Y(u2__abc_52155_new_n14843_));
AND2X2 AND2X2_6712 ( .A(u2__abc_52155_new_n14830_), .B(u2__abc_52155_new_n5743_), .Y(u2__abc_52155_new_n14845_));
AND2X2 AND2X2_6713 ( .A(u2__abc_52155_new_n14848_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14849_));
AND2X2 AND2X2_6714 ( .A(u2__abc_52155_new_n14849_), .B(u2__abc_52155_new_n14846_), .Y(u2__abc_52155_new_n14850_));
AND2X2 AND2X2_6715 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_365_), .Y(u2__abc_52155_new_n14851_));
AND2X2 AND2X2_6716 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5671_), .Y(u2__abc_52155_new_n14854_));
AND2X2 AND2X2_6717 ( .A(u2__abc_52155_new_n14855_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14856_));
AND2X2 AND2X2_6718 ( .A(u2__abc_52155_new_n14853_), .B(u2__abc_52155_new_n14856_), .Y(u2__abc_52155_new_n14857_));
AND2X2 AND2X2_6719 ( .A(u2__abc_52155_new_n14858_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__367_));
AND2X2 AND2X2_672 ( .A(u2__abc_52155_new_n3280_), .B(u2__abc_52155_new_n3321_), .Y(u2__abc_52155_new_n3322_));
AND2X2 AND2X2_6720 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_368_), .Y(u2__abc_52155_new_n14860_));
AND2X2 AND2X2_6721 ( .A(u2__abc_52155_new_n14715_), .B(u2__abc_52155_new_n5772_), .Y(u2__abc_52155_new_n14861_));
AND2X2 AND2X2_6722 ( .A(u2__abc_52155_new_n14790_), .B(u2__abc_52155_new_n5771_), .Y(u2__abc_52155_new_n14863_));
AND2X2 AND2X2_6723 ( .A(u2__abc_52155_new_n5753_), .B(u2__abc_52155_new_n5742_), .Y(u2__abc_52155_new_n14868_));
AND2X2 AND2X2_6724 ( .A(u2__abc_52155_new_n14867_), .B(u2__abc_52155_new_n14870_), .Y(u2__abc_52155_new_n14871_));
AND2X2 AND2X2_6725 ( .A(u2__abc_52155_new_n14864_), .B(u2__abc_52155_new_n14871_), .Y(u2__abc_52155_new_n14872_));
AND2X2 AND2X2_6726 ( .A(u2__abc_52155_new_n14862_), .B(u2__abc_52155_new_n14872_), .Y(u2__abc_52155_new_n14873_));
AND2X2 AND2X2_6727 ( .A(u2__abc_52155_new_n14560_), .B(u2__abc_52155_new_n5836_), .Y(u2__abc_52155_new_n14875_));
AND2X2 AND2X2_6728 ( .A(u2__abc_52155_new_n14876_), .B(u2__abc_52155_new_n5667_), .Y(u2__abc_52155_new_n14877_));
AND2X2 AND2X2_6729 ( .A(u2__abc_52155_new_n14879_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14880_));
AND2X2 AND2X2_673 ( .A(u2__abc_52155_new_n3323_), .B(u2_remHi_56_), .Y(u2__abc_52155_new_n3324_));
AND2X2 AND2X2_6730 ( .A(u2__abc_52155_new_n14880_), .B(u2__abc_52155_new_n14878_), .Y(u2__abc_52155_new_n14881_));
AND2X2 AND2X2_6731 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_366_), .Y(u2__abc_52155_new_n14882_));
AND2X2 AND2X2_6732 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5649_), .Y(u2__abc_52155_new_n14885_));
AND2X2 AND2X2_6733 ( .A(u2__abc_52155_new_n14886_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14887_));
AND2X2 AND2X2_6734 ( .A(u2__abc_52155_new_n14884_), .B(u2__abc_52155_new_n14887_), .Y(u2__abc_52155_new_n14888_));
AND2X2 AND2X2_6735 ( .A(u2__abc_52155_new_n14889_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__368_));
AND2X2 AND2X2_6736 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_369_), .Y(u2__abc_52155_new_n14891_));
AND2X2 AND2X2_6737 ( .A(u2__abc_52155_new_n14878_), .B(u2__abc_52155_new_n5663_), .Y(u2__abc_52155_new_n14892_));
AND2X2 AND2X2_6738 ( .A(u2__abc_52155_new_n14892_), .B(u2__abc_52155_new_n5674_), .Y(u2__abc_52155_new_n14893_));
AND2X2 AND2X2_6739 ( .A(u2__abc_52155_new_n14895_), .B(u2__abc_52155_new_n14894_), .Y(u2__abc_52155_new_n14896_));
AND2X2 AND2X2_674 ( .A(u2__abc_52155_new_n3326_), .B(sqrto_56_), .Y(u2__abc_52155_new_n3327_));
AND2X2 AND2X2_6740 ( .A(u2__abc_52155_new_n14897_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14898_));
AND2X2 AND2X2_6741 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_367_), .Y(u2__abc_52155_new_n14899_));
AND2X2 AND2X2_6742 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5656_), .Y(u2__abc_52155_new_n14902_));
AND2X2 AND2X2_6743 ( .A(u2__abc_52155_new_n14903_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14904_));
AND2X2 AND2X2_6744 ( .A(u2__abc_52155_new_n14901_), .B(u2__abc_52155_new_n14904_), .Y(u2__abc_52155_new_n14905_));
AND2X2 AND2X2_6745 ( .A(u2__abc_52155_new_n14906_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__369_));
AND2X2 AND2X2_6746 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_370_), .Y(u2__abc_52155_new_n14908_));
AND2X2 AND2X2_6747 ( .A(u2__abc_52155_new_n5663_), .B(u2__abc_52155_new_n5670_), .Y(u2__abc_52155_new_n14909_));
AND2X2 AND2X2_6748 ( .A(u2__abc_52155_new_n14878_), .B(u2__abc_52155_new_n14909_), .Y(u2__abc_52155_new_n14910_));
AND2X2 AND2X2_6749 ( .A(u2__abc_52155_new_n14912_), .B(u2__abc_52155_new_n5652_), .Y(u2__abc_52155_new_n14913_));
AND2X2 AND2X2_675 ( .A(u2__abc_52155_new_n3325_), .B(u2__abc_52155_new_n3328_), .Y(u2__abc_52155_new_n3329_));
AND2X2 AND2X2_6750 ( .A(u2__abc_52155_new_n14915_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14916_));
AND2X2 AND2X2_6751 ( .A(u2__abc_52155_new_n14916_), .B(u2__abc_52155_new_n14914_), .Y(u2__abc_52155_new_n14917_));
AND2X2 AND2X2_6752 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_368_), .Y(u2__abc_52155_new_n14918_));
AND2X2 AND2X2_6753 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5702_), .Y(u2__abc_52155_new_n14921_));
AND2X2 AND2X2_6754 ( .A(u2__abc_52155_new_n14922_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14923_));
AND2X2 AND2X2_6755 ( .A(u2__abc_52155_new_n14920_), .B(u2__abc_52155_new_n14923_), .Y(u2__abc_52155_new_n14924_));
AND2X2 AND2X2_6756 ( .A(u2__abc_52155_new_n14925_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__370_));
AND2X2 AND2X2_6757 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_371_), .Y(u2__abc_52155_new_n14927_));
AND2X2 AND2X2_6758 ( .A(u2__abc_52155_new_n14914_), .B(u2__abc_52155_new_n5648_), .Y(u2__abc_52155_new_n14929_));
AND2X2 AND2X2_6759 ( .A(u2__abc_52155_new_n14932_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14933_));
AND2X2 AND2X2_676 ( .A(u2__abc_52155_new_n3330_), .B(u2_remHi_57_), .Y(u2__abc_52155_new_n3331_));
AND2X2 AND2X2_6760 ( .A(u2__abc_52155_new_n14933_), .B(u2__abc_52155_new_n14930_), .Y(u2__abc_52155_new_n14934_));
AND2X2 AND2X2_6761 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_369_), .Y(u2__abc_52155_new_n14935_));
AND2X2 AND2X2_6762 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5695_), .Y(u2__abc_52155_new_n14938_));
AND2X2 AND2X2_6763 ( .A(u2__abc_52155_new_n14939_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14940_));
AND2X2 AND2X2_6764 ( .A(u2__abc_52155_new_n14937_), .B(u2__abc_52155_new_n14940_), .Y(u2__abc_52155_new_n14941_));
AND2X2 AND2X2_6765 ( .A(u2__abc_52155_new_n14942_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__371_));
AND2X2 AND2X2_6766 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_372_), .Y(u2__abc_52155_new_n14944_));
AND2X2 AND2X2_6767 ( .A(u2__abc_52155_new_n14945_), .B(u2__abc_52155_new_n5658_), .Y(u2__abc_52155_new_n14946_));
AND2X2 AND2X2_6768 ( .A(u2__abc_52155_new_n14949_), .B(u2__abc_52155_new_n14947_), .Y(u2__abc_52155_new_n14950_));
AND2X2 AND2X2_6769 ( .A(u2__abc_52155_new_n14876_), .B(u2__abc_52155_new_n5676_), .Y(u2__abc_52155_new_n14952_));
AND2X2 AND2X2_677 ( .A(u2__abc_52155_new_n3333_), .B(sqrto_57_), .Y(u2__abc_52155_new_n3334_));
AND2X2 AND2X2_6770 ( .A(u2__abc_52155_new_n14953_), .B(u2__abc_52155_new_n5705_), .Y(u2__abc_52155_new_n14954_));
AND2X2 AND2X2_6771 ( .A(u2__abc_52155_new_n14956_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14957_));
AND2X2 AND2X2_6772 ( .A(u2__abc_52155_new_n14957_), .B(u2__abc_52155_new_n14955_), .Y(u2__abc_52155_new_n14958_));
AND2X2 AND2X2_6773 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_370_), .Y(u2__abc_52155_new_n14959_));
AND2X2 AND2X2_6774 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5680_), .Y(u2__abc_52155_new_n14962_));
AND2X2 AND2X2_6775 ( .A(u2__abc_52155_new_n14963_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14964_));
AND2X2 AND2X2_6776 ( .A(u2__abc_52155_new_n14961_), .B(u2__abc_52155_new_n14964_), .Y(u2__abc_52155_new_n14965_));
AND2X2 AND2X2_6777 ( .A(u2__abc_52155_new_n14966_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__372_));
AND2X2 AND2X2_6778 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_373_), .Y(u2__abc_52155_new_n14968_));
AND2X2 AND2X2_6779 ( .A(u2__abc_52155_new_n14955_), .B(u2__abc_52155_new_n5701_), .Y(u2__abc_52155_new_n14969_));
AND2X2 AND2X2_678 ( .A(u2__abc_52155_new_n3332_), .B(u2__abc_52155_new_n3335_), .Y(u2__abc_52155_new_n3336_));
AND2X2 AND2X2_6780 ( .A(u2__abc_52155_new_n14970_), .B(u2__abc_52155_new_n5698_), .Y(u2__abc_52155_new_n14971_));
AND2X2 AND2X2_6781 ( .A(u2__abc_52155_new_n14973_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14974_));
AND2X2 AND2X2_6782 ( .A(u2__abc_52155_new_n14974_), .B(u2__abc_52155_new_n14972_), .Y(u2__abc_52155_new_n14975_));
AND2X2 AND2X2_6783 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_371_), .Y(u2__abc_52155_new_n14976_));
AND2X2 AND2X2_6784 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5687_), .Y(u2__abc_52155_new_n14979_));
AND2X2 AND2X2_6785 ( .A(u2__abc_52155_new_n14980_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14981_));
AND2X2 AND2X2_6786 ( .A(u2__abc_52155_new_n14978_), .B(u2__abc_52155_new_n14981_), .Y(u2__abc_52155_new_n14982_));
AND2X2 AND2X2_6787 ( .A(u2__abc_52155_new_n14983_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__373_));
AND2X2 AND2X2_6788 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_374_), .Y(u2__abc_52155_new_n14985_));
AND2X2 AND2X2_6789 ( .A(u2__abc_52155_new_n14972_), .B(u2__abc_52155_new_n5694_), .Y(u2__abc_52155_new_n14986_));
AND2X2 AND2X2_679 ( .A(u2__abc_52155_new_n3329_), .B(u2__abc_52155_new_n3336_), .Y(u2__abc_52155_new_n3337_));
AND2X2 AND2X2_6790 ( .A(u2__abc_52155_new_n14987_), .B(u2__abc_52155_new_n5683_), .Y(u2__abc_52155_new_n14988_));
AND2X2 AND2X2_6791 ( .A(u2__abc_52155_new_n14990_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n14991_));
AND2X2 AND2X2_6792 ( .A(u2__abc_52155_new_n14991_), .B(u2__abc_52155_new_n14989_), .Y(u2__abc_52155_new_n14992_));
AND2X2 AND2X2_6793 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_372_), .Y(u2__abc_52155_new_n14993_));
AND2X2 AND2X2_6794 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5614_), .Y(u2__abc_52155_new_n14996_));
AND2X2 AND2X2_6795 ( .A(u2__abc_52155_new_n14997_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n14998_));
AND2X2 AND2X2_6796 ( .A(u2__abc_52155_new_n14995_), .B(u2__abc_52155_new_n14998_), .Y(u2__abc_52155_new_n14999_));
AND2X2 AND2X2_6797 ( .A(u2__abc_52155_new_n15000_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__374_));
AND2X2 AND2X2_6798 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_375_), .Y(u2__abc_52155_new_n15002_));
AND2X2 AND2X2_6799 ( .A(u2__abc_52155_new_n14989_), .B(u2__abc_52155_new_n5679_), .Y(u2__abc_52155_new_n15004_));
AND2X2 AND2X2_68 ( .A(_abc_73687_new_n753_), .B(sqrto_67_), .Y(\o[103] ));
AND2X2 AND2X2_680 ( .A(u2__abc_52155_new_n3338_), .B(u2_remHi_54_), .Y(u2__abc_52155_new_n3339_));
AND2X2 AND2X2_6800 ( .A(u2__abc_52155_new_n15007_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15008_));
AND2X2 AND2X2_6801 ( .A(u2__abc_52155_new_n15008_), .B(u2__abc_52155_new_n15005_), .Y(u2__abc_52155_new_n15009_));
AND2X2 AND2X2_6802 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_373_), .Y(u2__abc_52155_new_n15010_));
AND2X2 AND2X2_6803 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5621_), .Y(u2__abc_52155_new_n15013_));
AND2X2 AND2X2_6804 ( .A(u2__abc_52155_new_n15014_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15015_));
AND2X2 AND2X2_6805 ( .A(u2__abc_52155_new_n15012_), .B(u2__abc_52155_new_n15015_), .Y(u2__abc_52155_new_n15016_));
AND2X2 AND2X2_6806 ( .A(u2__abc_52155_new_n15017_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__375_));
AND2X2 AND2X2_6807 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_376_), .Y(u2__abc_52155_new_n15019_));
AND2X2 AND2X2_6808 ( .A(u2__abc_52155_new_n14951_), .B(u2__abc_52155_new_n5707_), .Y(u2__abc_52155_new_n15020_));
AND2X2 AND2X2_6809 ( .A(u2__abc_52155_new_n5697_), .B(u2__abc_52155_new_n5700_), .Y(u2__abc_52155_new_n15021_));
AND2X2 AND2X2_681 ( .A(u2__abc_52155_new_n3341_), .B(sqrto_54_), .Y(u2__abc_52155_new_n3342_));
AND2X2 AND2X2_6810 ( .A(u2__abc_52155_new_n15022_), .B(u2__abc_52155_new_n5691_), .Y(u2__abc_52155_new_n15023_));
AND2X2 AND2X2_6811 ( .A(u2__abc_52155_new_n5689_), .B(u2__abc_52155_new_n5678_), .Y(u2__abc_52155_new_n15024_));
AND2X2 AND2X2_6812 ( .A(u2__abc_52155_new_n14876_), .B(u2__abc_52155_new_n5708_), .Y(u2__abc_52155_new_n15028_));
AND2X2 AND2X2_6813 ( .A(u2__abc_52155_new_n15029_), .B(u2__abc_52155_new_n5620_), .Y(u2__abc_52155_new_n15030_));
AND2X2 AND2X2_6814 ( .A(u2__abc_52155_new_n15032_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15033_));
AND2X2 AND2X2_6815 ( .A(u2__abc_52155_new_n15033_), .B(u2__abc_52155_new_n15031_), .Y(u2__abc_52155_new_n15034_));
AND2X2 AND2X2_6816 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_374_), .Y(u2__abc_52155_new_n15035_));
AND2X2 AND2X2_6817 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5632_), .Y(u2__abc_52155_new_n15038_));
AND2X2 AND2X2_6818 ( .A(u2__abc_52155_new_n15039_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15040_));
AND2X2 AND2X2_6819 ( .A(u2__abc_52155_new_n15037_), .B(u2__abc_52155_new_n15040_), .Y(u2__abc_52155_new_n15041_));
AND2X2 AND2X2_682 ( .A(u2__abc_52155_new_n3340_), .B(u2__abc_52155_new_n3343_), .Y(u2__abc_52155_new_n3344_));
AND2X2 AND2X2_6820 ( .A(u2__abc_52155_new_n15042_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__376_));
AND2X2 AND2X2_6821 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_377_), .Y(u2__abc_52155_new_n15044_));
AND2X2 AND2X2_6822 ( .A(u2__abc_52155_new_n15031_), .B(u2__abc_52155_new_n5619_), .Y(u2__abc_52155_new_n15046_));
AND2X2 AND2X2_6823 ( .A(u2__abc_52155_new_n15049_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15050_));
AND2X2 AND2X2_6824 ( .A(u2__abc_52155_new_n15050_), .B(u2__abc_52155_new_n15047_), .Y(u2__abc_52155_new_n15051_));
AND2X2 AND2X2_6825 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_375_), .Y(u2__abc_52155_new_n15052_));
AND2X2 AND2X2_6826 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5639_), .Y(u2__abc_52155_new_n15055_));
AND2X2 AND2X2_6827 ( .A(u2__abc_52155_new_n15056_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15057_));
AND2X2 AND2X2_6828 ( .A(u2__abc_52155_new_n15054_), .B(u2__abc_52155_new_n15057_), .Y(u2__abc_52155_new_n15058_));
AND2X2 AND2X2_6829 ( .A(u2__abc_52155_new_n15059_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__377_));
AND2X2 AND2X2_683 ( .A(u2__abc_52155_new_n3345_), .B(u2_remHi_55_), .Y(u2__abc_52155_new_n3346_));
AND2X2 AND2X2_6830 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_378_), .Y(u2__abc_52155_new_n15061_));
AND2X2 AND2X2_6831 ( .A(u2__abc_52155_new_n5619_), .B(u2__abc_52155_new_n5626_), .Y(u2__abc_52155_new_n15062_));
AND2X2 AND2X2_6832 ( .A(u2__abc_52155_new_n15029_), .B(u2__abc_52155_new_n5628_), .Y(u2__abc_52155_new_n15065_));
AND2X2 AND2X2_6833 ( .A(u2__abc_52155_new_n15066_), .B(u2__abc_52155_new_n5635_), .Y(u2__abc_52155_new_n15067_));
AND2X2 AND2X2_6834 ( .A(u2__abc_52155_new_n15069_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15070_));
AND2X2 AND2X2_6835 ( .A(u2__abc_52155_new_n15070_), .B(u2__abc_52155_new_n15068_), .Y(u2__abc_52155_new_n15071_));
AND2X2 AND2X2_6836 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_376_), .Y(u2__abc_52155_new_n15072_));
AND2X2 AND2X2_6837 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5601_), .Y(u2__abc_52155_new_n15075_));
AND2X2 AND2X2_6838 ( .A(u2__abc_52155_new_n15076_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15077_));
AND2X2 AND2X2_6839 ( .A(u2__abc_52155_new_n15074_), .B(u2__abc_52155_new_n15077_), .Y(u2__abc_52155_new_n15078_));
AND2X2 AND2X2_684 ( .A(u2__abc_52155_new_n3348_), .B(sqrto_55_), .Y(u2__abc_52155_new_n3349_));
AND2X2 AND2X2_6840 ( .A(u2__abc_52155_new_n15079_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__378_));
AND2X2 AND2X2_6841 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_379_), .Y(u2__abc_52155_new_n15081_));
AND2X2 AND2X2_6842 ( .A(u2__abc_52155_new_n15068_), .B(u2__abc_52155_new_n5631_), .Y(u2__abc_52155_new_n15083_));
AND2X2 AND2X2_6843 ( .A(u2__abc_52155_new_n15086_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15087_));
AND2X2 AND2X2_6844 ( .A(u2__abc_52155_new_n15087_), .B(u2__abc_52155_new_n15084_), .Y(u2__abc_52155_new_n15088_));
AND2X2 AND2X2_6845 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_377_), .Y(u2__abc_52155_new_n15089_));
AND2X2 AND2X2_6846 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5608_), .Y(u2__abc_52155_new_n15092_));
AND2X2 AND2X2_6847 ( .A(u2__abc_52155_new_n15093_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15094_));
AND2X2 AND2X2_6848 ( .A(u2__abc_52155_new_n15091_), .B(u2__abc_52155_new_n15094_), .Y(u2__abc_52155_new_n15095_));
AND2X2 AND2X2_6849 ( .A(u2__abc_52155_new_n15096_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__379_));
AND2X2 AND2X2_685 ( .A(u2__abc_52155_new_n3347_), .B(u2__abc_52155_new_n3350_), .Y(u2__abc_52155_new_n3351_));
AND2X2 AND2X2_6850 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_380_), .Y(u2__abc_52155_new_n15098_));
AND2X2 AND2X2_6851 ( .A(u2__abc_52155_new_n5641_), .B(u2__abc_52155_new_n5630_), .Y(u2__abc_52155_new_n15099_));
AND2X2 AND2X2_6852 ( .A(u2__abc_52155_new_n15066_), .B(u2__abc_52155_new_n5643_), .Y(u2__abc_52155_new_n15101_));
AND2X2 AND2X2_6853 ( .A(u2__abc_52155_new_n15102_), .B(u2__abc_52155_new_n5604_), .Y(u2__abc_52155_new_n15103_));
AND2X2 AND2X2_6854 ( .A(u2__abc_52155_new_n15105_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15106_));
AND2X2 AND2X2_6855 ( .A(u2__abc_52155_new_n15106_), .B(u2__abc_52155_new_n15104_), .Y(u2__abc_52155_new_n15107_));
AND2X2 AND2X2_6856 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_378_), .Y(u2__abc_52155_new_n15108_));
AND2X2 AND2X2_6857 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5586_), .Y(u2__abc_52155_new_n15111_));
AND2X2 AND2X2_6858 ( .A(u2__abc_52155_new_n15112_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15113_));
AND2X2 AND2X2_6859 ( .A(u2__abc_52155_new_n15110_), .B(u2__abc_52155_new_n15113_), .Y(u2__abc_52155_new_n15114_));
AND2X2 AND2X2_686 ( .A(u2__abc_52155_new_n3344_), .B(u2__abc_52155_new_n3351_), .Y(u2__abc_52155_new_n3352_));
AND2X2 AND2X2_6860 ( .A(u2__abc_52155_new_n15115_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__380_));
AND2X2 AND2X2_6861 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_381_), .Y(u2__abc_52155_new_n15117_));
AND2X2 AND2X2_6862 ( .A(u2__abc_52155_new_n15104_), .B(u2__abc_52155_new_n5600_), .Y(u2__abc_52155_new_n15118_));
AND2X2 AND2X2_6863 ( .A(u2__abc_52155_new_n15118_), .B(u2__abc_52155_new_n5611_), .Y(u2__abc_52155_new_n15119_));
AND2X2 AND2X2_6864 ( .A(u2__abc_52155_new_n15121_), .B(u2__abc_52155_new_n15120_), .Y(u2__abc_52155_new_n15122_));
AND2X2 AND2X2_6865 ( .A(u2__abc_52155_new_n15123_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15124_));
AND2X2 AND2X2_6866 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_379_), .Y(u2__abc_52155_new_n15125_));
AND2X2 AND2X2_6867 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n5590_), .Y(u2__abc_52155_new_n15128_));
AND2X2 AND2X2_6868 ( .A(u2__abc_52155_new_n15129_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15130_));
AND2X2 AND2X2_6869 ( .A(u2__abc_52155_new_n15127_), .B(u2__abc_52155_new_n15130_), .Y(u2__abc_52155_new_n15131_));
AND2X2 AND2X2_687 ( .A(u2__abc_52155_new_n3337_), .B(u2__abc_52155_new_n3352_), .Y(u2__abc_52155_new_n3353_));
AND2X2 AND2X2_6870 ( .A(u2__abc_52155_new_n15132_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__381_));
AND2X2 AND2X2_6871 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_382_), .Y(u2__abc_52155_new_n15134_));
AND2X2 AND2X2_6872 ( .A(u2__abc_52155_new_n5600_), .B(u2__abc_52155_new_n5607_), .Y(u2__abc_52155_new_n15135_));
AND2X2 AND2X2_6873 ( .A(u2__abc_52155_new_n15104_), .B(u2__abc_52155_new_n15135_), .Y(u2__abc_52155_new_n15136_));
AND2X2 AND2X2_6874 ( .A(u2__abc_52155_new_n15138_), .B(u2__abc_52155_new_n5589_), .Y(u2__abc_52155_new_n15139_));
AND2X2 AND2X2_6875 ( .A(u2__abc_52155_new_n15141_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15142_));
AND2X2 AND2X2_6876 ( .A(u2__abc_52155_new_n15142_), .B(u2__abc_52155_new_n15140_), .Y(u2__abc_52155_new_n15143_));
AND2X2 AND2X2_6877 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_380_), .Y(u2__abc_52155_new_n15144_));
AND2X2 AND2X2_6878 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7238_), .Y(u2__abc_52155_new_n15147_));
AND2X2 AND2X2_6879 ( .A(u2__abc_52155_new_n15148_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15149_));
AND2X2 AND2X2_688 ( .A(u2__abc_52155_new_n3354_), .B(u2_remHi_60_), .Y(u2__abc_52155_new_n3355_));
AND2X2 AND2X2_6880 ( .A(u2__abc_52155_new_n15146_), .B(u2__abc_52155_new_n15149_), .Y(u2__abc_52155_new_n15150_));
AND2X2 AND2X2_6881 ( .A(u2__abc_52155_new_n15151_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__382_));
AND2X2 AND2X2_6882 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_383_), .Y(u2__abc_52155_new_n15153_));
AND2X2 AND2X2_6883 ( .A(u2__abc_52155_new_n15140_), .B(u2__abc_52155_new_n5585_), .Y(u2__abc_52155_new_n15155_));
AND2X2 AND2X2_6884 ( .A(u2__abc_52155_new_n15158_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15159_));
AND2X2 AND2X2_6885 ( .A(u2__abc_52155_new_n15159_), .B(u2__abc_52155_new_n15156_), .Y(u2__abc_52155_new_n15160_));
AND2X2 AND2X2_6886 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_381_), .Y(u2__abc_52155_new_n15161_));
AND2X2 AND2X2_6887 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7228_), .Y(u2__abc_52155_new_n15164_));
AND2X2 AND2X2_6888 ( .A(u2__abc_52155_new_n15165_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15166_));
AND2X2 AND2X2_6889 ( .A(u2__abc_52155_new_n15163_), .B(u2__abc_52155_new_n15166_), .Y(u2__abc_52155_new_n15167_));
AND2X2 AND2X2_689 ( .A(u2__abc_52155_new_n3357_), .B(sqrto_60_), .Y(u2__abc_52155_new_n3358_));
AND2X2 AND2X2_6890 ( .A(u2__abc_52155_new_n15168_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__383_));
AND2X2 AND2X2_6891 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_384_), .Y(u2__abc_52155_new_n15170_));
AND2X2 AND2X2_6892 ( .A(u2__abc_52155_new_n12663_), .B(u2__abc_52155_new_n6605_), .Y(u2__abc_52155_new_n15171_));
AND2X2 AND2X2_6893 ( .A(u2__abc_52155_new_n13926_), .B(u2__abc_52155_new_n6093_), .Y(u2__abc_52155_new_n15173_));
AND2X2 AND2X2_6894 ( .A(u2__abc_52155_new_n14558_), .B(u2__abc_52155_new_n5837_), .Y(u2__abc_52155_new_n15175_));
AND2X2 AND2X2_6895 ( .A(u2__abc_52155_new_n14874_), .B(u2__abc_52155_new_n5709_), .Y(u2__abc_52155_new_n15177_));
AND2X2 AND2X2_6896 ( .A(u2__abc_52155_new_n15027_), .B(u2__abc_52155_new_n5645_), .Y(u2__abc_52155_new_n15179_));
AND2X2 AND2X2_6897 ( .A(u2__abc_52155_new_n15064_), .B(u2__abc_52155_new_n5643_), .Y(u2__abc_52155_new_n15181_));
AND2X2 AND2X2_6898 ( .A(u2__abc_52155_new_n15182_), .B(u2__abc_52155_new_n5613_), .Y(u2__abc_52155_new_n15183_));
AND2X2 AND2X2_6899 ( .A(u2__abc_52155_new_n5592_), .B(u2__abc_52155_new_n5584_), .Y(u2__abc_52155_new_n15187_));
AND2X2 AND2X2_69 ( .A(_abc_73687_new_n753_), .B(sqrto_68_), .Y(\o[104] ));
AND2X2 AND2X2_690 ( .A(u2__abc_52155_new_n3356_), .B(u2__abc_52155_new_n3359_), .Y(u2__abc_52155_new_n3360_));
AND2X2 AND2X2_6900 ( .A(u2__abc_52155_new_n15186_), .B(u2__abc_52155_new_n15189_), .Y(u2__abc_52155_new_n15190_));
AND2X2 AND2X2_6901 ( .A(u2__abc_52155_new_n15184_), .B(u2__abc_52155_new_n15190_), .Y(u2__abc_52155_new_n15191_));
AND2X2 AND2X2_6902 ( .A(u2__abc_52155_new_n15180_), .B(u2__abc_52155_new_n15191_), .Y(u2__abc_52155_new_n15192_));
AND2X2 AND2X2_6903 ( .A(u2__abc_52155_new_n15178_), .B(u2__abc_52155_new_n15192_), .Y(u2__abc_52155_new_n15193_));
AND2X2 AND2X2_6904 ( .A(u2__abc_52155_new_n15176_), .B(u2__abc_52155_new_n15193_), .Y(u2__abc_52155_new_n15194_));
AND2X2 AND2X2_6905 ( .A(u2__abc_52155_new_n15174_), .B(u2__abc_52155_new_n15194_), .Y(u2__abc_52155_new_n15195_));
AND2X2 AND2X2_6906 ( .A(u2__abc_52155_new_n15172_), .B(u2__abc_52155_new_n15195_), .Y(u2__abc_52155_new_n15196_));
AND2X2 AND2X2_6907 ( .A(u2__abc_52155_new_n15197_), .B(u2__abc_52155_new_n7241_), .Y(u2__abc_52155_new_n15198_));
AND2X2 AND2X2_6908 ( .A(u2__abc_52155_new_n15200_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15201_));
AND2X2 AND2X2_6909 ( .A(u2__abc_52155_new_n15201_), .B(u2__abc_52155_new_n15199_), .Y(u2__abc_52155_new_n15202_));
AND2X2 AND2X2_691 ( .A(u2__abc_52155_new_n3361_), .B(sqrto_61_), .Y(u2__abc_52155_new_n3362_));
AND2X2 AND2X2_6910 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_382_), .Y(u2__abc_52155_new_n15203_));
AND2X2 AND2X2_6911 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7216_), .Y(u2__abc_52155_new_n15206_));
AND2X2 AND2X2_6912 ( .A(u2__abc_52155_new_n15207_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15208_));
AND2X2 AND2X2_6913 ( .A(u2__abc_52155_new_n15205_), .B(u2__abc_52155_new_n15208_), .Y(u2__abc_52155_new_n15209_));
AND2X2 AND2X2_6914 ( .A(u2__abc_52155_new_n15210_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__384_));
AND2X2 AND2X2_6915 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_385_), .Y(u2__abc_52155_new_n15212_));
AND2X2 AND2X2_6916 ( .A(u2__abc_52155_new_n15199_), .B(u2__abc_52155_new_n7237_), .Y(u2__abc_52155_new_n15214_));
AND2X2 AND2X2_6917 ( .A(u2__abc_52155_new_n15217_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15218_));
AND2X2 AND2X2_6918 ( .A(u2__abc_52155_new_n15218_), .B(u2__abc_52155_new_n15215_), .Y(u2__abc_52155_new_n15219_));
AND2X2 AND2X2_6919 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_383_), .Y(u2__abc_52155_new_n15220_));
AND2X2 AND2X2_692 ( .A(u2__abc_52155_new_n3364_), .B(u2_remHi_61_), .Y(u2__abc_52155_new_n3365_));
AND2X2 AND2X2_6920 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7220_), .Y(u2__abc_52155_new_n15223_));
AND2X2 AND2X2_6921 ( .A(u2__abc_52155_new_n15224_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15225_));
AND2X2 AND2X2_6922 ( .A(u2__abc_52155_new_n15222_), .B(u2__abc_52155_new_n15225_), .Y(u2__abc_52155_new_n15226_));
AND2X2 AND2X2_6923 ( .A(u2__abc_52155_new_n15227_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__385_));
AND2X2 AND2X2_6924 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_386_), .Y(u2__abc_52155_new_n15229_));
AND2X2 AND2X2_6925 ( .A(u2__abc_52155_new_n7233_), .B(u2__abc_52155_new_n7237_), .Y(u2__abc_52155_new_n15230_));
AND2X2 AND2X2_6926 ( .A(u2__abc_52155_new_n15199_), .B(u2__abc_52155_new_n15230_), .Y(u2__abc_52155_new_n15231_));
AND2X2 AND2X2_6927 ( .A(u2__abc_52155_new_n15233_), .B(u2__abc_52155_new_n7219_), .Y(u2__abc_52155_new_n15234_));
AND2X2 AND2X2_6928 ( .A(u2__abc_52155_new_n15236_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15237_));
AND2X2 AND2X2_6929 ( .A(u2__abc_52155_new_n15237_), .B(u2__abc_52155_new_n15235_), .Y(u2__abc_52155_new_n15238_));
AND2X2 AND2X2_693 ( .A(u2__abc_52155_new_n3363_), .B(u2__abc_52155_new_n3366_), .Y(u2__abc_52155_new_n3367_));
AND2X2 AND2X2_6930 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_384_), .Y(u2__abc_52155_new_n15239_));
AND2X2 AND2X2_6931 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7207_), .Y(u2__abc_52155_new_n15242_));
AND2X2 AND2X2_6932 ( .A(u2__abc_52155_new_n15243_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15244_));
AND2X2 AND2X2_6933 ( .A(u2__abc_52155_new_n15241_), .B(u2__abc_52155_new_n15244_), .Y(u2__abc_52155_new_n15245_));
AND2X2 AND2X2_6934 ( .A(u2__abc_52155_new_n15246_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__386_));
AND2X2 AND2X2_6935 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_387_), .Y(u2__abc_52155_new_n15248_));
AND2X2 AND2X2_6936 ( .A(u2__abc_52155_new_n15235_), .B(u2__abc_52155_new_n7215_), .Y(u2__abc_52155_new_n15250_));
AND2X2 AND2X2_6937 ( .A(u2__abc_52155_new_n15253_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15254_));
AND2X2 AND2X2_6938 ( .A(u2__abc_52155_new_n15254_), .B(u2__abc_52155_new_n15251_), .Y(u2__abc_52155_new_n15255_));
AND2X2 AND2X2_6939 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_385_), .Y(u2__abc_52155_new_n15256_));
AND2X2 AND2X2_694 ( .A(u2__abc_52155_new_n3360_), .B(u2__abc_52155_new_n3367_), .Y(u2__abc_52155_new_n3368_));
AND2X2 AND2X2_6940 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7197_), .Y(u2__abc_52155_new_n15259_));
AND2X2 AND2X2_6941 ( .A(u2__abc_52155_new_n15260_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15261_));
AND2X2 AND2X2_6942 ( .A(u2__abc_52155_new_n15258_), .B(u2__abc_52155_new_n15261_), .Y(u2__abc_52155_new_n15262_));
AND2X2 AND2X2_6943 ( .A(u2__abc_52155_new_n15263_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__387_));
AND2X2 AND2X2_6944 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_388_), .Y(u2__abc_52155_new_n15265_));
AND2X2 AND2X2_6945 ( .A(u2__abc_52155_new_n15267_), .B(u2__abc_52155_new_n7227_), .Y(u2__abc_52155_new_n15268_));
AND2X2 AND2X2_6946 ( .A(u2__abc_52155_new_n7222_), .B(u2__abc_52155_new_n7214_), .Y(u2__abc_52155_new_n15269_));
AND2X2 AND2X2_6947 ( .A(u2__abc_52155_new_n15197_), .B(u2__abc_52155_new_n7243_), .Y(u2__abc_52155_new_n15272_));
AND2X2 AND2X2_6948 ( .A(u2__abc_52155_new_n15273_), .B(u2__abc_52155_new_n7210_), .Y(u2__abc_52155_new_n15274_));
AND2X2 AND2X2_6949 ( .A(u2__abc_52155_new_n15276_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15277_));
AND2X2 AND2X2_695 ( .A(u2__abc_52155_new_n3369_), .B(u2_remHi_59_), .Y(u2__abc_52155_new_n3370_));
AND2X2 AND2X2_6950 ( .A(u2__abc_52155_new_n15277_), .B(u2__abc_52155_new_n15275_), .Y(u2__abc_52155_new_n15278_));
AND2X2 AND2X2_6951 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_386_), .Y(u2__abc_52155_new_n15279_));
AND2X2 AND2X2_6952 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7185_), .Y(u2__abc_52155_new_n15282_));
AND2X2 AND2X2_6953 ( .A(u2__abc_52155_new_n15283_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15284_));
AND2X2 AND2X2_6954 ( .A(u2__abc_52155_new_n15281_), .B(u2__abc_52155_new_n15284_), .Y(u2__abc_52155_new_n15285_));
AND2X2 AND2X2_6955 ( .A(u2__abc_52155_new_n15286_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__388_));
AND2X2 AND2X2_6956 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_389_), .Y(u2__abc_52155_new_n15288_));
AND2X2 AND2X2_6957 ( .A(u2__abc_52155_new_n15275_), .B(u2__abc_52155_new_n7206_), .Y(u2__abc_52155_new_n15289_));
AND2X2 AND2X2_6958 ( .A(u2__abc_52155_new_n15289_), .B(u2__abc_52155_new_n7203_), .Y(u2__abc_52155_new_n15290_));
AND2X2 AND2X2_6959 ( .A(u2__abc_52155_new_n15292_), .B(u2__abc_52155_new_n15291_), .Y(u2__abc_52155_new_n15293_));
AND2X2 AND2X2_696 ( .A(u2__abc_52155_new_n3372_), .B(sqrto_59_), .Y(u2__abc_52155_new_n3373_));
AND2X2 AND2X2_6960 ( .A(u2__abc_52155_new_n15294_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15295_));
AND2X2 AND2X2_6961 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_387_), .Y(u2__abc_52155_new_n15296_));
AND2X2 AND2X2_6962 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7192_), .Y(u2__abc_52155_new_n15299_));
AND2X2 AND2X2_6963 ( .A(u2__abc_52155_new_n15300_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15301_));
AND2X2 AND2X2_6964 ( .A(u2__abc_52155_new_n15298_), .B(u2__abc_52155_new_n15301_), .Y(u2__abc_52155_new_n15302_));
AND2X2 AND2X2_6965 ( .A(u2__abc_52155_new_n15303_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__389_));
AND2X2 AND2X2_6966 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_390_), .Y(u2__abc_52155_new_n15305_));
AND2X2 AND2X2_6967 ( .A(u2__abc_52155_new_n7202_), .B(u2__abc_52155_new_n7206_), .Y(u2__abc_52155_new_n15306_));
AND2X2 AND2X2_6968 ( .A(u2__abc_52155_new_n15275_), .B(u2__abc_52155_new_n15306_), .Y(u2__abc_52155_new_n15307_));
AND2X2 AND2X2_6969 ( .A(u2__abc_52155_new_n15309_), .B(u2__abc_52155_new_n7188_), .Y(u2__abc_52155_new_n15310_));
AND2X2 AND2X2_697 ( .A(u2__abc_52155_new_n3371_), .B(u2__abc_52155_new_n3374_), .Y(u2__abc_52155_new_n3375_));
AND2X2 AND2X2_6970 ( .A(u2__abc_52155_new_n15312_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15313_));
AND2X2 AND2X2_6971 ( .A(u2__abc_52155_new_n15313_), .B(u2__abc_52155_new_n15311_), .Y(u2__abc_52155_new_n15314_));
AND2X2 AND2X2_6972 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_388_), .Y(u2__abc_52155_new_n15315_));
AND2X2 AND2X2_6973 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7390_), .Y(u2__abc_52155_new_n15318_));
AND2X2 AND2X2_6974 ( .A(u2__abc_52155_new_n15319_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15320_));
AND2X2 AND2X2_6975 ( .A(u2__abc_52155_new_n15317_), .B(u2__abc_52155_new_n15320_), .Y(u2__abc_52155_new_n15321_));
AND2X2 AND2X2_6976 ( .A(u2__abc_52155_new_n15322_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__390_));
AND2X2 AND2X2_6977 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_391_), .Y(u2__abc_52155_new_n15324_));
AND2X2 AND2X2_6978 ( .A(u2__abc_52155_new_n15311_), .B(u2__abc_52155_new_n7184_), .Y(u2__abc_52155_new_n15326_));
AND2X2 AND2X2_6979 ( .A(u2__abc_52155_new_n15329_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15330_));
AND2X2 AND2X2_698 ( .A(u2__abc_52155_new_n3376_), .B(u2_remHi_58_), .Y(u2__abc_52155_new_n3377_));
AND2X2 AND2X2_6980 ( .A(u2__abc_52155_new_n15330_), .B(u2__abc_52155_new_n15327_), .Y(u2__abc_52155_new_n15331_));
AND2X2 AND2X2_6981 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_389_), .Y(u2__abc_52155_new_n15332_));
AND2X2 AND2X2_6982 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7394_), .Y(u2__abc_52155_new_n15335_));
AND2X2 AND2X2_6983 ( .A(u2__abc_52155_new_n15336_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15337_));
AND2X2 AND2X2_6984 ( .A(u2__abc_52155_new_n15334_), .B(u2__abc_52155_new_n15337_), .Y(u2__abc_52155_new_n15338_));
AND2X2 AND2X2_6985 ( .A(u2__abc_52155_new_n15339_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__391_));
AND2X2 AND2X2_6986 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_392_), .Y(u2__abc_52155_new_n15341_));
AND2X2 AND2X2_6987 ( .A(u2__abc_52155_new_n15271_), .B(u2__abc_52155_new_n7212_), .Y(u2__abc_52155_new_n15342_));
AND2X2 AND2X2_6988 ( .A(u2__abc_52155_new_n15344_), .B(u2__abc_52155_new_n7196_), .Y(u2__abc_52155_new_n15345_));
AND2X2 AND2X2_6989 ( .A(u2__abc_52155_new_n7194_), .B(u2__abc_52155_new_n7183_), .Y(u2__abc_52155_new_n15346_));
AND2X2 AND2X2_699 ( .A(u2__abc_52155_new_n3379_), .B(sqrto_58_), .Y(u2__abc_52155_new_n3380_));
AND2X2 AND2X2_6990 ( .A(u2__abc_52155_new_n15197_), .B(u2__abc_52155_new_n7244_), .Y(u2__abc_52155_new_n15350_));
AND2X2 AND2X2_6991 ( .A(u2__abc_52155_new_n15351_), .B(u2__abc_52155_new_n7393_), .Y(u2__abc_52155_new_n15352_));
AND2X2 AND2X2_6992 ( .A(u2__abc_52155_new_n15354_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15355_));
AND2X2 AND2X2_6993 ( .A(u2__abc_52155_new_n15355_), .B(u2__abc_52155_new_n15353_), .Y(u2__abc_52155_new_n15356_));
AND2X2 AND2X2_6994 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_390_), .Y(u2__abc_52155_new_n15357_));
AND2X2 AND2X2_6995 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7375_), .Y(u2__abc_52155_new_n15360_));
AND2X2 AND2X2_6996 ( .A(u2__abc_52155_new_n15361_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15362_));
AND2X2 AND2X2_6997 ( .A(u2__abc_52155_new_n15359_), .B(u2__abc_52155_new_n15362_), .Y(u2__abc_52155_new_n15363_));
AND2X2 AND2X2_6998 ( .A(u2__abc_52155_new_n15364_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__392_));
AND2X2 AND2X2_6999 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_393_), .Y(u2__abc_52155_new_n15366_));
AND2X2 AND2X2_7 ( .A(_abc_73687_new_n753_), .B(sqrto_6_), .Y(\o[42] ));
AND2X2 AND2X2_70 ( .A(_abc_73687_new_n753_), .B(sqrto_69_), .Y(\o[105] ));
AND2X2 AND2X2_700 ( .A(u2__abc_52155_new_n3378_), .B(u2__abc_52155_new_n3381_), .Y(u2__abc_52155_new_n3382_));
AND2X2 AND2X2_7000 ( .A(u2__abc_52155_new_n15353_), .B(u2__abc_52155_new_n7389_), .Y(u2__abc_52155_new_n15368_));
AND2X2 AND2X2_7001 ( .A(u2__abc_52155_new_n15369_), .B(u2__abc_52155_new_n15367_), .Y(u2__abc_52155_new_n15370_));
AND2X2 AND2X2_7002 ( .A(u2__abc_52155_new_n15368_), .B(u2__abc_52155_new_n7400_), .Y(u2__abc_52155_new_n15371_));
AND2X2 AND2X2_7003 ( .A(u2__abc_52155_new_n15372_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15373_));
AND2X2 AND2X2_7004 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_391_), .Y(u2__abc_52155_new_n15374_));
AND2X2 AND2X2_7005 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7379_), .Y(u2__abc_52155_new_n15377_));
AND2X2 AND2X2_7006 ( .A(u2__abc_52155_new_n15378_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15379_));
AND2X2 AND2X2_7007 ( .A(u2__abc_52155_new_n15376_), .B(u2__abc_52155_new_n15379_), .Y(u2__abc_52155_new_n15380_));
AND2X2 AND2X2_7008 ( .A(u2__abc_52155_new_n15381_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__393_));
AND2X2 AND2X2_7009 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_394_), .Y(u2__abc_52155_new_n15383_));
AND2X2 AND2X2_701 ( .A(u2__abc_52155_new_n3375_), .B(u2__abc_52155_new_n3382_), .Y(u2__abc_52155_new_n3383_));
AND2X2 AND2X2_7010 ( .A(u2__abc_52155_new_n15369_), .B(u2__abc_52155_new_n7396_), .Y(u2__abc_52155_new_n15384_));
AND2X2 AND2X2_7011 ( .A(u2__abc_52155_new_n15385_), .B(u2__abc_52155_new_n7378_), .Y(u2__abc_52155_new_n15386_));
AND2X2 AND2X2_7012 ( .A(u2__abc_52155_new_n15388_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15389_));
AND2X2 AND2X2_7013 ( .A(u2__abc_52155_new_n15389_), .B(u2__abc_52155_new_n15387_), .Y(u2__abc_52155_new_n15390_));
AND2X2 AND2X2_7014 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_392_), .Y(u2__abc_52155_new_n15391_));
AND2X2 AND2X2_7015 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7428_), .Y(u2__abc_52155_new_n15394_));
AND2X2 AND2X2_7016 ( .A(u2__abc_52155_new_n15395_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15396_));
AND2X2 AND2X2_7017 ( .A(u2__abc_52155_new_n15393_), .B(u2__abc_52155_new_n15396_), .Y(u2__abc_52155_new_n15397_));
AND2X2 AND2X2_7018 ( .A(u2__abc_52155_new_n15398_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__394_));
AND2X2 AND2X2_7019 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_395_), .Y(u2__abc_52155_new_n15400_));
AND2X2 AND2X2_702 ( .A(u2__abc_52155_new_n3368_), .B(u2__abc_52155_new_n3383_), .Y(u2__abc_52155_new_n3384_));
AND2X2 AND2X2_7020 ( .A(u2__abc_52155_new_n15387_), .B(u2__abc_52155_new_n7374_), .Y(u2__abc_52155_new_n15402_));
AND2X2 AND2X2_7021 ( .A(u2__abc_52155_new_n15405_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15406_));
AND2X2 AND2X2_7022 ( .A(u2__abc_52155_new_n15406_), .B(u2__abc_52155_new_n15403_), .Y(u2__abc_52155_new_n15407_));
AND2X2 AND2X2_7023 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_393_), .Y(u2__abc_52155_new_n15408_));
AND2X2 AND2X2_7024 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7418_), .Y(u2__abc_52155_new_n15411_));
AND2X2 AND2X2_7025 ( .A(u2__abc_52155_new_n15412_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15413_));
AND2X2 AND2X2_7026 ( .A(u2__abc_52155_new_n15410_), .B(u2__abc_52155_new_n15413_), .Y(u2__abc_52155_new_n15414_));
AND2X2 AND2X2_7027 ( .A(u2__abc_52155_new_n15415_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__395_));
AND2X2 AND2X2_7028 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_396_), .Y(u2__abc_52155_new_n15417_));
AND2X2 AND2X2_7029 ( .A(u2__abc_52155_new_n7389_), .B(u2__abc_52155_new_n7399_), .Y(u2__abc_52155_new_n15418_));
AND2X2 AND2X2_703 ( .A(u2__abc_52155_new_n3353_), .B(u2__abc_52155_new_n3384_), .Y(u2__abc_52155_new_n3385_));
AND2X2 AND2X2_7030 ( .A(u2__abc_52155_new_n15420_), .B(u2__abc_52155_new_n7386_), .Y(u2__abc_52155_new_n15421_));
AND2X2 AND2X2_7031 ( .A(u2__abc_52155_new_n7381_), .B(u2__abc_52155_new_n7373_), .Y(u2__abc_52155_new_n15422_));
AND2X2 AND2X2_7032 ( .A(u2__abc_52155_new_n15351_), .B(u2__abc_52155_new_n7402_), .Y(u2__abc_52155_new_n15425_));
AND2X2 AND2X2_7033 ( .A(u2__abc_52155_new_n15426_), .B(u2__abc_52155_new_n7431_), .Y(u2__abc_52155_new_n15427_));
AND2X2 AND2X2_7034 ( .A(u2__abc_52155_new_n15429_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15430_));
AND2X2 AND2X2_7035 ( .A(u2__abc_52155_new_n15430_), .B(u2__abc_52155_new_n15428_), .Y(u2__abc_52155_new_n15431_));
AND2X2 AND2X2_7036 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_394_), .Y(u2__abc_52155_new_n15432_));
AND2X2 AND2X2_7037 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7406_), .Y(u2__abc_52155_new_n15435_));
AND2X2 AND2X2_7038 ( .A(u2__abc_52155_new_n15436_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15437_));
AND2X2 AND2X2_7039 ( .A(u2__abc_52155_new_n15434_), .B(u2__abc_52155_new_n15437_), .Y(u2__abc_52155_new_n15438_));
AND2X2 AND2X2_704 ( .A(u2__abc_52155_new_n3386_), .B(u2_remHi_48_), .Y(u2__abc_52155_new_n3387_));
AND2X2 AND2X2_7040 ( .A(u2__abc_52155_new_n15439_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__396_));
AND2X2 AND2X2_7041 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_397_), .Y(u2__abc_52155_new_n15441_));
AND2X2 AND2X2_7042 ( .A(u2__abc_52155_new_n15428_), .B(u2__abc_52155_new_n7427_), .Y(u2__abc_52155_new_n15442_));
AND2X2 AND2X2_7043 ( .A(u2__abc_52155_new_n15442_), .B(u2__abc_52155_new_n7424_), .Y(u2__abc_52155_new_n15443_));
AND2X2 AND2X2_7044 ( .A(u2__abc_52155_new_n15445_), .B(u2__abc_52155_new_n15444_), .Y(u2__abc_52155_new_n15446_));
AND2X2 AND2X2_7045 ( .A(u2__abc_52155_new_n15447_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15448_));
AND2X2 AND2X2_7046 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_395_), .Y(u2__abc_52155_new_n15449_));
AND2X2 AND2X2_7047 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7413_), .Y(u2__abc_52155_new_n15452_));
AND2X2 AND2X2_7048 ( .A(u2__abc_52155_new_n15453_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15454_));
AND2X2 AND2X2_7049 ( .A(u2__abc_52155_new_n15451_), .B(u2__abc_52155_new_n15454_), .Y(u2__abc_52155_new_n15455_));
AND2X2 AND2X2_705 ( .A(u2__abc_52155_new_n3388_), .B(sqrto_48_), .Y(u2__abc_52155_new_n3389_));
AND2X2 AND2X2_7050 ( .A(u2__abc_52155_new_n15456_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__397_));
AND2X2 AND2X2_7051 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_398_), .Y(u2__abc_52155_new_n15458_));
AND2X2 AND2X2_7052 ( .A(u2__abc_52155_new_n7423_), .B(u2__abc_52155_new_n7427_), .Y(u2__abc_52155_new_n15459_));
AND2X2 AND2X2_7053 ( .A(u2__abc_52155_new_n15428_), .B(u2__abc_52155_new_n15459_), .Y(u2__abc_52155_new_n15460_));
AND2X2 AND2X2_7054 ( .A(u2__abc_52155_new_n15462_), .B(u2__abc_52155_new_n7409_), .Y(u2__abc_52155_new_n15463_));
AND2X2 AND2X2_7055 ( .A(u2__abc_52155_new_n15465_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15466_));
AND2X2 AND2X2_7056 ( .A(u2__abc_52155_new_n15466_), .B(u2__abc_52155_new_n15464_), .Y(u2__abc_52155_new_n15467_));
AND2X2 AND2X2_7057 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_396_), .Y(u2__abc_52155_new_n15468_));
AND2X2 AND2X2_7058 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7311_), .Y(u2__abc_52155_new_n15471_));
AND2X2 AND2X2_7059 ( .A(u2__abc_52155_new_n15472_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15473_));
AND2X2 AND2X2_706 ( .A(u2__abc_52155_new_n3391_), .B(u2_remHi_49_), .Y(u2__abc_52155_new_n3392_));
AND2X2 AND2X2_7060 ( .A(u2__abc_52155_new_n15470_), .B(u2__abc_52155_new_n15473_), .Y(u2__abc_52155_new_n15474_));
AND2X2 AND2X2_7061 ( .A(u2__abc_52155_new_n15475_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__398_));
AND2X2 AND2X2_7062 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_399_), .Y(u2__abc_52155_new_n15477_));
AND2X2 AND2X2_7063 ( .A(u2__abc_52155_new_n15464_), .B(u2__abc_52155_new_n7405_), .Y(u2__abc_52155_new_n15479_));
AND2X2 AND2X2_7064 ( .A(u2__abc_52155_new_n15482_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15483_));
AND2X2 AND2X2_7065 ( .A(u2__abc_52155_new_n15483_), .B(u2__abc_52155_new_n15480_), .Y(u2__abc_52155_new_n15484_));
AND2X2 AND2X2_7066 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_397_), .Y(u2__abc_52155_new_n15485_));
AND2X2 AND2X2_7067 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7315_), .Y(u2__abc_52155_new_n15488_));
AND2X2 AND2X2_7068 ( .A(u2__abc_52155_new_n15489_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15490_));
AND2X2 AND2X2_7069 ( .A(u2__abc_52155_new_n15487_), .B(u2__abc_52155_new_n15490_), .Y(u2__abc_52155_new_n15491_));
AND2X2 AND2X2_707 ( .A(u2__abc_52155_new_n3393_), .B(sqrto_49_), .Y(u2__abc_52155_new_n3394_));
AND2X2 AND2X2_7070 ( .A(u2__abc_52155_new_n15492_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__399_));
AND2X2 AND2X2_7071 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_400_), .Y(u2__abc_52155_new_n15494_));
AND2X2 AND2X2_7072 ( .A(u2__abc_52155_new_n15424_), .B(u2__abc_52155_new_n7433_), .Y(u2__abc_52155_new_n15495_));
AND2X2 AND2X2_7073 ( .A(u2__abc_52155_new_n15497_), .B(u2__abc_52155_new_n7417_), .Y(u2__abc_52155_new_n15498_));
AND2X2 AND2X2_7074 ( .A(u2__abc_52155_new_n7415_), .B(u2__abc_52155_new_n7404_), .Y(u2__abc_52155_new_n15499_));
AND2X2 AND2X2_7075 ( .A(u2__abc_52155_new_n15351_), .B(u2__abc_52155_new_n7434_), .Y(u2__abc_52155_new_n15503_));
AND2X2 AND2X2_7076 ( .A(u2__abc_52155_new_n15504_), .B(u2__abc_52155_new_n7314_), .Y(u2__abc_52155_new_n15505_));
AND2X2 AND2X2_7077 ( .A(u2__abc_52155_new_n15507_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15508_));
AND2X2 AND2X2_7078 ( .A(u2__abc_52155_new_n15508_), .B(u2__abc_52155_new_n15506_), .Y(u2__abc_52155_new_n15509_));
AND2X2 AND2X2_7079 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_398_), .Y(u2__abc_52155_new_n15510_));
AND2X2 AND2X2_708 ( .A(u2__abc_52155_new_n3398_), .B(u2_remHi_47_), .Y(u2__abc_52155_new_n3399_));
AND2X2 AND2X2_7080 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7326_), .Y(u2__abc_52155_new_n15513_));
AND2X2 AND2X2_7081 ( .A(u2__abc_52155_new_n15514_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15515_));
AND2X2 AND2X2_7082 ( .A(u2__abc_52155_new_n15512_), .B(u2__abc_52155_new_n15515_), .Y(u2__abc_52155_new_n15516_));
AND2X2 AND2X2_7083 ( .A(u2__abc_52155_new_n15517_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__400_));
AND2X2 AND2X2_7084 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_401_), .Y(u2__abc_52155_new_n15519_));
AND2X2 AND2X2_7085 ( .A(u2__abc_52155_new_n15506_), .B(u2__abc_52155_new_n7310_), .Y(u2__abc_52155_new_n15521_));
AND2X2 AND2X2_7086 ( .A(u2__abc_52155_new_n15524_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15525_));
AND2X2 AND2X2_7087 ( .A(u2__abc_52155_new_n15525_), .B(u2__abc_52155_new_n15522_), .Y(u2__abc_52155_new_n15526_));
AND2X2 AND2X2_7088 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_399_), .Y(u2__abc_52155_new_n15527_));
AND2X2 AND2X2_7089 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7330_), .Y(u2__abc_52155_new_n15530_));
AND2X2 AND2X2_709 ( .A(u2__abc_52155_new_n3401_), .B(sqrto_47_), .Y(u2__abc_52155_new_n3402_));
AND2X2 AND2X2_7090 ( .A(u2__abc_52155_new_n15531_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15532_));
AND2X2 AND2X2_7091 ( .A(u2__abc_52155_new_n15529_), .B(u2__abc_52155_new_n15532_), .Y(u2__abc_52155_new_n15533_));
AND2X2 AND2X2_7092 ( .A(u2__abc_52155_new_n15534_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__401_));
AND2X2 AND2X2_7093 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_402_), .Y(u2__abc_52155_new_n15536_));
AND2X2 AND2X2_7094 ( .A(u2__abc_52155_new_n15537_), .B(u2__abc_52155_new_n7320_), .Y(u2__abc_52155_new_n15538_));
AND2X2 AND2X2_7095 ( .A(u2__abc_52155_new_n15504_), .B(u2__abc_52155_new_n7322_), .Y(u2__abc_52155_new_n15540_));
AND2X2 AND2X2_7096 ( .A(u2__abc_52155_new_n15541_), .B(u2__abc_52155_new_n7329_), .Y(u2__abc_52155_new_n15542_));
AND2X2 AND2X2_7097 ( .A(u2__abc_52155_new_n15544_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15545_));
AND2X2 AND2X2_7098 ( .A(u2__abc_52155_new_n15545_), .B(u2__abc_52155_new_n15543_), .Y(u2__abc_52155_new_n15546_));
AND2X2 AND2X2_7099 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_400_), .Y(u2__abc_52155_new_n15547_));
AND2X2 AND2X2_71 ( .A(_abc_73687_new_n753_), .B(sqrto_70_), .Y(\o[106] ));
AND2X2 AND2X2_710 ( .A(u2__abc_52155_new_n3400_), .B(u2__abc_52155_new_n3403_), .Y(u2__abc_52155_new_n3404_));
AND2X2 AND2X2_7100 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7364_), .Y(u2__abc_52155_new_n15550_));
AND2X2 AND2X2_7101 ( .A(u2__abc_52155_new_n15551_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15552_));
AND2X2 AND2X2_7102 ( .A(u2__abc_52155_new_n15549_), .B(u2__abc_52155_new_n15552_), .Y(u2__abc_52155_new_n15553_));
AND2X2 AND2X2_7103 ( .A(u2__abc_52155_new_n15554_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__402_));
AND2X2 AND2X2_7104 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_403_), .Y(u2__abc_52155_new_n15556_));
AND2X2 AND2X2_7105 ( .A(u2__abc_52155_new_n15543_), .B(u2__abc_52155_new_n7325_), .Y(u2__abc_52155_new_n15558_));
AND2X2 AND2X2_7106 ( .A(u2__abc_52155_new_n15561_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15562_));
AND2X2 AND2X2_7107 ( .A(u2__abc_52155_new_n15562_), .B(u2__abc_52155_new_n15559_), .Y(u2__abc_52155_new_n15563_));
AND2X2 AND2X2_7108 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_401_), .Y(u2__abc_52155_new_n15564_));
AND2X2 AND2X2_7109 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7354_), .Y(u2__abc_52155_new_n15567_));
AND2X2 AND2X2_711 ( .A(u2__abc_52155_new_n3405_), .B(u2_remHi_46_), .Y(u2__abc_52155_new_n3406_));
AND2X2 AND2X2_7110 ( .A(u2__abc_52155_new_n15568_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15569_));
AND2X2 AND2X2_7111 ( .A(u2__abc_52155_new_n15566_), .B(u2__abc_52155_new_n15569_), .Y(u2__abc_52155_new_n15570_));
AND2X2 AND2X2_7112 ( .A(u2__abc_52155_new_n15571_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__403_));
AND2X2 AND2X2_7113 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_404_), .Y(u2__abc_52155_new_n15573_));
AND2X2 AND2X2_7114 ( .A(u2__abc_52155_new_n15539_), .B(u2__abc_52155_new_n7337_), .Y(u2__abc_52155_new_n15574_));
AND2X2 AND2X2_7115 ( .A(u2__abc_52155_new_n7332_), .B(u2__abc_52155_new_n7324_), .Y(u2__abc_52155_new_n15575_));
AND2X2 AND2X2_7116 ( .A(u2__abc_52155_new_n15504_), .B(u2__abc_52155_new_n7338_), .Y(u2__abc_52155_new_n15578_));
AND2X2 AND2X2_7117 ( .A(u2__abc_52155_new_n15579_), .B(u2__abc_52155_new_n7367_), .Y(u2__abc_52155_new_n15580_));
AND2X2 AND2X2_7118 ( .A(u2__abc_52155_new_n15582_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15583_));
AND2X2 AND2X2_7119 ( .A(u2__abc_52155_new_n15583_), .B(u2__abc_52155_new_n15581_), .Y(u2__abc_52155_new_n15584_));
AND2X2 AND2X2_712 ( .A(u2__abc_52155_new_n3408_), .B(sqrto_46_), .Y(u2__abc_52155_new_n3409_));
AND2X2 AND2X2_7120 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_402_), .Y(u2__abc_52155_new_n15585_));
AND2X2 AND2X2_7121 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7342_), .Y(u2__abc_52155_new_n15588_));
AND2X2 AND2X2_7122 ( .A(u2__abc_52155_new_n15589_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15590_));
AND2X2 AND2X2_7123 ( .A(u2__abc_52155_new_n15587_), .B(u2__abc_52155_new_n15590_), .Y(u2__abc_52155_new_n15591_));
AND2X2 AND2X2_7124 ( .A(u2__abc_52155_new_n15592_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__404_));
AND2X2 AND2X2_7125 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_405_), .Y(u2__abc_52155_new_n15594_));
AND2X2 AND2X2_7126 ( .A(u2__abc_52155_new_n15581_), .B(u2__abc_52155_new_n7363_), .Y(u2__abc_52155_new_n15595_));
AND2X2 AND2X2_7127 ( .A(u2__abc_52155_new_n15595_), .B(u2__abc_52155_new_n7360_), .Y(u2__abc_52155_new_n15596_));
AND2X2 AND2X2_7128 ( .A(u2__abc_52155_new_n15598_), .B(u2__abc_52155_new_n15597_), .Y(u2__abc_52155_new_n15599_));
AND2X2 AND2X2_7129 ( .A(u2__abc_52155_new_n15600_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15601_));
AND2X2 AND2X2_713 ( .A(u2__abc_52155_new_n3407_), .B(u2__abc_52155_new_n3410_), .Y(u2__abc_52155_new_n3411_));
AND2X2 AND2X2_7130 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_403_), .Y(u2__abc_52155_new_n15602_));
AND2X2 AND2X2_7131 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7349_), .Y(u2__abc_52155_new_n15605_));
AND2X2 AND2X2_7132 ( .A(u2__abc_52155_new_n15606_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15607_));
AND2X2 AND2X2_7133 ( .A(u2__abc_52155_new_n15604_), .B(u2__abc_52155_new_n15607_), .Y(u2__abc_52155_new_n15608_));
AND2X2 AND2X2_7134 ( .A(u2__abc_52155_new_n15609_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__405_));
AND2X2 AND2X2_7135 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_406_), .Y(u2__abc_52155_new_n15611_));
AND2X2 AND2X2_7136 ( .A(u2__abc_52155_new_n7359_), .B(u2__abc_52155_new_n7363_), .Y(u2__abc_52155_new_n15612_));
AND2X2 AND2X2_7137 ( .A(u2__abc_52155_new_n15581_), .B(u2__abc_52155_new_n15612_), .Y(u2__abc_52155_new_n15613_));
AND2X2 AND2X2_7138 ( .A(u2__abc_52155_new_n15615_), .B(u2__abc_52155_new_n7345_), .Y(u2__abc_52155_new_n15616_));
AND2X2 AND2X2_7139 ( .A(u2__abc_52155_new_n15618_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15619_));
AND2X2 AND2X2_714 ( .A(u2__abc_52155_new_n3404_), .B(u2__abc_52155_new_n3411_), .Y(u2__abc_52155_new_n3412_));
AND2X2 AND2X2_7140 ( .A(u2__abc_52155_new_n15619_), .B(u2__abc_52155_new_n15617_), .Y(u2__abc_52155_new_n15620_));
AND2X2 AND2X2_7141 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_404_), .Y(u2__abc_52155_new_n15621_));
AND2X2 AND2X2_7142 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7270_), .Y(u2__abc_52155_new_n15624_));
AND2X2 AND2X2_7143 ( .A(u2__abc_52155_new_n15625_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15626_));
AND2X2 AND2X2_7144 ( .A(u2__abc_52155_new_n15623_), .B(u2__abc_52155_new_n15626_), .Y(u2__abc_52155_new_n15627_));
AND2X2 AND2X2_7145 ( .A(u2__abc_52155_new_n15628_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__406_));
AND2X2 AND2X2_7146 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_407_), .Y(u2__abc_52155_new_n15630_));
AND2X2 AND2X2_7147 ( .A(u2__abc_52155_new_n15617_), .B(u2__abc_52155_new_n7341_), .Y(u2__abc_52155_new_n15632_));
AND2X2 AND2X2_7148 ( .A(u2__abc_52155_new_n15635_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15636_));
AND2X2 AND2X2_7149 ( .A(u2__abc_52155_new_n15636_), .B(u2__abc_52155_new_n15633_), .Y(u2__abc_52155_new_n15637_));
AND2X2 AND2X2_715 ( .A(u2__abc_52155_new_n3397_), .B(u2__abc_52155_new_n3412_), .Y(u2__abc_52155_new_n3413_));
AND2X2 AND2X2_7150 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_405_), .Y(u2__abc_52155_new_n15638_));
AND2X2 AND2X2_7151 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7260_), .Y(u2__abc_52155_new_n15641_));
AND2X2 AND2X2_7152 ( .A(u2__abc_52155_new_n15642_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15643_));
AND2X2 AND2X2_7153 ( .A(u2__abc_52155_new_n15640_), .B(u2__abc_52155_new_n15643_), .Y(u2__abc_52155_new_n15644_));
AND2X2 AND2X2_7154 ( .A(u2__abc_52155_new_n15645_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__407_));
AND2X2 AND2X2_7155 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_408_), .Y(u2__abc_52155_new_n15647_));
AND2X2 AND2X2_7156 ( .A(u2__abc_52155_new_n15577_), .B(u2__abc_52155_new_n7369_), .Y(u2__abc_52155_new_n15648_));
AND2X2 AND2X2_7157 ( .A(u2__abc_52155_new_n15650_), .B(u2__abc_52155_new_n7353_), .Y(u2__abc_52155_new_n15651_));
AND2X2 AND2X2_7158 ( .A(u2__abc_52155_new_n7351_), .B(u2__abc_52155_new_n7340_), .Y(u2__abc_52155_new_n15652_));
AND2X2 AND2X2_7159 ( .A(u2__abc_52155_new_n15504_), .B(u2__abc_52155_new_n7370_), .Y(u2__abc_52155_new_n15656_));
AND2X2 AND2X2_716 ( .A(u2__abc_52155_new_n3414_), .B(u2_remHi_52_), .Y(u2__abc_52155_new_n3415_));
AND2X2 AND2X2_7160 ( .A(u2__abc_52155_new_n15657_), .B(u2__abc_52155_new_n7273_), .Y(u2__abc_52155_new_n15658_));
AND2X2 AND2X2_7161 ( .A(u2__abc_52155_new_n15660_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15661_));
AND2X2 AND2X2_7162 ( .A(u2__abc_52155_new_n15661_), .B(u2__abc_52155_new_n15659_), .Y(u2__abc_52155_new_n15662_));
AND2X2 AND2X2_7163 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_406_), .Y(u2__abc_52155_new_n15663_));
AND2X2 AND2X2_7164 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7248_), .Y(u2__abc_52155_new_n15666_));
AND2X2 AND2X2_7165 ( .A(u2__abc_52155_new_n15667_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15668_));
AND2X2 AND2X2_7166 ( .A(u2__abc_52155_new_n15665_), .B(u2__abc_52155_new_n15668_), .Y(u2__abc_52155_new_n15669_));
AND2X2 AND2X2_7167 ( .A(u2__abc_52155_new_n15670_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__408_));
AND2X2 AND2X2_7168 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_409_), .Y(u2__abc_52155_new_n15672_));
AND2X2 AND2X2_7169 ( .A(u2__abc_52155_new_n15659_), .B(u2__abc_52155_new_n7269_), .Y(u2__abc_52155_new_n15673_));
AND2X2 AND2X2_717 ( .A(u2__abc_52155_new_n3417_), .B(sqrto_52_), .Y(u2__abc_52155_new_n3418_));
AND2X2 AND2X2_7170 ( .A(u2__abc_52155_new_n15673_), .B(u2__abc_52155_new_n7266_), .Y(u2__abc_52155_new_n15674_));
AND2X2 AND2X2_7171 ( .A(u2__abc_52155_new_n15676_), .B(u2__abc_52155_new_n15675_), .Y(u2__abc_52155_new_n15677_));
AND2X2 AND2X2_7172 ( .A(u2__abc_52155_new_n15678_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15679_));
AND2X2 AND2X2_7173 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_407_), .Y(u2__abc_52155_new_n15680_));
AND2X2 AND2X2_7174 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7252_), .Y(u2__abc_52155_new_n15683_));
AND2X2 AND2X2_7175 ( .A(u2__abc_52155_new_n15684_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15685_));
AND2X2 AND2X2_7176 ( .A(u2__abc_52155_new_n15682_), .B(u2__abc_52155_new_n15685_), .Y(u2__abc_52155_new_n15686_));
AND2X2 AND2X2_7177 ( .A(u2__abc_52155_new_n15687_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__409_));
AND2X2 AND2X2_7178 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_410_), .Y(u2__abc_52155_new_n15689_));
AND2X2 AND2X2_7179 ( .A(u2__abc_52155_new_n7265_), .B(u2__abc_52155_new_n7269_), .Y(u2__abc_52155_new_n15690_));
AND2X2 AND2X2_718 ( .A(u2__abc_52155_new_n3416_), .B(u2__abc_52155_new_n3419_), .Y(u2__abc_52155_new_n3420_));
AND2X2 AND2X2_7180 ( .A(u2__abc_52155_new_n15659_), .B(u2__abc_52155_new_n15690_), .Y(u2__abc_52155_new_n15691_));
AND2X2 AND2X2_7181 ( .A(u2__abc_52155_new_n15693_), .B(u2__abc_52155_new_n7251_), .Y(u2__abc_52155_new_n15694_));
AND2X2 AND2X2_7182 ( .A(u2__abc_52155_new_n15696_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15697_));
AND2X2 AND2X2_7183 ( .A(u2__abc_52155_new_n15697_), .B(u2__abc_52155_new_n15695_), .Y(u2__abc_52155_new_n15698_));
AND2X2 AND2X2_7184 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_408_), .Y(u2__abc_52155_new_n15699_));
AND2X2 AND2X2_7185 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7301_), .Y(u2__abc_52155_new_n15702_));
AND2X2 AND2X2_7186 ( .A(u2__abc_52155_new_n15703_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15704_));
AND2X2 AND2X2_7187 ( .A(u2__abc_52155_new_n15701_), .B(u2__abc_52155_new_n15704_), .Y(u2__abc_52155_new_n15705_));
AND2X2 AND2X2_7188 ( .A(u2__abc_52155_new_n15706_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__410_));
AND2X2 AND2X2_7189 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_411_), .Y(u2__abc_52155_new_n15708_));
AND2X2 AND2X2_719 ( .A(u2__abc_52155_new_n3421_), .B(u2_remHi_53_), .Y(u2__abc_52155_new_n3422_));
AND2X2 AND2X2_7190 ( .A(u2__abc_52155_new_n15695_), .B(u2__abc_52155_new_n7247_), .Y(u2__abc_52155_new_n15710_));
AND2X2 AND2X2_7191 ( .A(u2__abc_52155_new_n15713_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15714_));
AND2X2 AND2X2_7192 ( .A(u2__abc_52155_new_n15714_), .B(u2__abc_52155_new_n15711_), .Y(u2__abc_52155_new_n15715_));
AND2X2 AND2X2_7193 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_409_), .Y(u2__abc_52155_new_n15716_));
AND2X2 AND2X2_7194 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7291_), .Y(u2__abc_52155_new_n15719_));
AND2X2 AND2X2_7195 ( .A(u2__abc_52155_new_n15720_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15721_));
AND2X2 AND2X2_7196 ( .A(u2__abc_52155_new_n15718_), .B(u2__abc_52155_new_n15721_), .Y(u2__abc_52155_new_n15722_));
AND2X2 AND2X2_7197 ( .A(u2__abc_52155_new_n15723_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__411_));
AND2X2 AND2X2_7198 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_412_), .Y(u2__abc_52155_new_n15725_));
AND2X2 AND2X2_7199 ( .A(u2__abc_52155_new_n15727_), .B(u2__abc_52155_new_n7259_), .Y(u2__abc_52155_new_n15728_));
AND2X2 AND2X2_72 ( .A(_abc_73687_new_n753_), .B(sqrto_71_), .Y(\o[107] ));
AND2X2 AND2X2_720 ( .A(u2__abc_52155_new_n3424_), .B(sqrto_53_), .Y(u2__abc_52155_new_n3425_));
AND2X2 AND2X2_7200 ( .A(u2__abc_52155_new_n7254_), .B(u2__abc_52155_new_n7246_), .Y(u2__abc_52155_new_n15729_));
AND2X2 AND2X2_7201 ( .A(u2__abc_52155_new_n15657_), .B(u2__abc_52155_new_n7275_), .Y(u2__abc_52155_new_n15732_));
AND2X2 AND2X2_7202 ( .A(u2__abc_52155_new_n15733_), .B(u2__abc_52155_new_n7304_), .Y(u2__abc_52155_new_n15734_));
AND2X2 AND2X2_7203 ( .A(u2__abc_52155_new_n15736_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15737_));
AND2X2 AND2X2_7204 ( .A(u2__abc_52155_new_n15737_), .B(u2__abc_52155_new_n15735_), .Y(u2__abc_52155_new_n15738_));
AND2X2 AND2X2_7205 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_410_), .Y(u2__abc_52155_new_n15739_));
AND2X2 AND2X2_7206 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7279_), .Y(u2__abc_52155_new_n15742_));
AND2X2 AND2X2_7207 ( .A(u2__abc_52155_new_n15743_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15744_));
AND2X2 AND2X2_7208 ( .A(u2__abc_52155_new_n15741_), .B(u2__abc_52155_new_n15744_), .Y(u2__abc_52155_new_n15745_));
AND2X2 AND2X2_7209 ( .A(u2__abc_52155_new_n15746_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__412_));
AND2X2 AND2X2_721 ( .A(u2__abc_52155_new_n3423_), .B(u2__abc_52155_new_n3426_), .Y(u2__abc_52155_new_n3427_));
AND2X2 AND2X2_7210 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_413_), .Y(u2__abc_52155_new_n15748_));
AND2X2 AND2X2_7211 ( .A(u2__abc_52155_new_n15735_), .B(u2__abc_52155_new_n7300_), .Y(u2__abc_52155_new_n15749_));
AND2X2 AND2X2_7212 ( .A(u2__abc_52155_new_n15749_), .B(u2__abc_52155_new_n7297_), .Y(u2__abc_52155_new_n15750_));
AND2X2 AND2X2_7213 ( .A(u2__abc_52155_new_n15752_), .B(u2__abc_52155_new_n15751_), .Y(u2__abc_52155_new_n15753_));
AND2X2 AND2X2_7214 ( .A(u2__abc_52155_new_n15754_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15755_));
AND2X2 AND2X2_7215 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_411_), .Y(u2__abc_52155_new_n15756_));
AND2X2 AND2X2_7216 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7286_), .Y(u2__abc_52155_new_n15759_));
AND2X2 AND2X2_7217 ( .A(u2__abc_52155_new_n15760_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15761_));
AND2X2 AND2X2_7218 ( .A(u2__abc_52155_new_n15758_), .B(u2__abc_52155_new_n15761_), .Y(u2__abc_52155_new_n15762_));
AND2X2 AND2X2_7219 ( .A(u2__abc_52155_new_n15763_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__413_));
AND2X2 AND2X2_722 ( .A(u2__abc_52155_new_n3420_), .B(u2__abc_52155_new_n3427_), .Y(u2__abc_52155_new_n3428_));
AND2X2 AND2X2_7220 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_414_), .Y(u2__abc_52155_new_n15765_));
AND2X2 AND2X2_7221 ( .A(u2__abc_52155_new_n7296_), .B(u2__abc_52155_new_n7300_), .Y(u2__abc_52155_new_n15766_));
AND2X2 AND2X2_7222 ( .A(u2__abc_52155_new_n15735_), .B(u2__abc_52155_new_n15766_), .Y(u2__abc_52155_new_n15767_));
AND2X2 AND2X2_7223 ( .A(u2__abc_52155_new_n15769_), .B(u2__abc_52155_new_n7282_), .Y(u2__abc_52155_new_n15770_));
AND2X2 AND2X2_7224 ( .A(u2__abc_52155_new_n15772_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15773_));
AND2X2 AND2X2_7225 ( .A(u2__abc_52155_new_n15773_), .B(u2__abc_52155_new_n15771_), .Y(u2__abc_52155_new_n15774_));
AND2X2 AND2X2_7226 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_412_), .Y(u2__abc_52155_new_n15775_));
AND2X2 AND2X2_7227 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7173_), .Y(u2__abc_52155_new_n15778_));
AND2X2 AND2X2_7228 ( .A(u2__abc_52155_new_n15779_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15780_));
AND2X2 AND2X2_7229 ( .A(u2__abc_52155_new_n15777_), .B(u2__abc_52155_new_n15780_), .Y(u2__abc_52155_new_n15781_));
AND2X2 AND2X2_723 ( .A(u2__abc_52155_new_n3429_), .B(u2_remHi_51_), .Y(u2__abc_52155_new_n3430_));
AND2X2 AND2X2_7230 ( .A(u2__abc_52155_new_n15782_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__414_));
AND2X2 AND2X2_7231 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_415_), .Y(u2__abc_52155_new_n15784_));
AND2X2 AND2X2_7232 ( .A(u2__abc_52155_new_n15771_), .B(u2__abc_52155_new_n7278_), .Y(u2__abc_52155_new_n15786_));
AND2X2 AND2X2_7233 ( .A(u2__abc_52155_new_n15789_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15790_));
AND2X2 AND2X2_7234 ( .A(u2__abc_52155_new_n15790_), .B(u2__abc_52155_new_n15787_), .Y(u2__abc_52155_new_n15791_));
AND2X2 AND2X2_7235 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_413_), .Y(u2__abc_52155_new_n15792_));
AND2X2 AND2X2_7236 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7163_), .Y(u2__abc_52155_new_n15795_));
AND2X2 AND2X2_7237 ( .A(u2__abc_52155_new_n15796_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15797_));
AND2X2 AND2X2_7238 ( .A(u2__abc_52155_new_n15794_), .B(u2__abc_52155_new_n15797_), .Y(u2__abc_52155_new_n15798_));
AND2X2 AND2X2_7239 ( .A(u2__abc_52155_new_n15799_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__415_));
AND2X2 AND2X2_724 ( .A(u2__abc_52155_new_n3432_), .B(sqrto_51_), .Y(u2__abc_52155_new_n3433_));
AND2X2 AND2X2_7240 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_416_), .Y(u2__abc_52155_new_n15801_));
AND2X2 AND2X2_7241 ( .A(u2__abc_52155_new_n15197_), .B(u2__abc_52155_new_n7436_), .Y(u2__abc_52155_new_n15802_));
AND2X2 AND2X2_7242 ( .A(u2__abc_52155_new_n15731_), .B(u2__abc_52155_new_n7306_), .Y(u2__abc_52155_new_n15803_));
AND2X2 AND2X2_7243 ( .A(u2__abc_52155_new_n15805_), .B(u2__abc_52155_new_n7290_), .Y(u2__abc_52155_new_n15806_));
AND2X2 AND2X2_7244 ( .A(u2__abc_52155_new_n7288_), .B(u2__abc_52155_new_n7277_), .Y(u2__abc_52155_new_n15807_));
AND2X2 AND2X2_7245 ( .A(u2__abc_52155_new_n15349_), .B(u2__abc_52155_new_n7435_), .Y(u2__abc_52155_new_n15811_));
AND2X2 AND2X2_7246 ( .A(u2__abc_52155_new_n15655_), .B(u2__abc_52155_new_n7307_), .Y(u2__abc_52155_new_n15813_));
AND2X2 AND2X2_7247 ( .A(u2__abc_52155_new_n15502_), .B(u2__abc_52155_new_n7371_), .Y(u2__abc_52155_new_n15814_));
AND2X2 AND2X2_7248 ( .A(u2__abc_52155_new_n15817_), .B(u2__abc_52155_new_n7176_), .Y(u2__abc_52155_new_n15818_));
AND2X2 AND2X2_7249 ( .A(u2__abc_52155_new_n15820_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15821_));
AND2X2 AND2X2_725 ( .A(u2__abc_52155_new_n3431_), .B(u2__abc_52155_new_n3434_), .Y(u2__abc_52155_new_n3435_));
AND2X2 AND2X2_7250 ( .A(u2__abc_52155_new_n15821_), .B(u2__abc_52155_new_n15819_), .Y(u2__abc_52155_new_n15822_));
AND2X2 AND2X2_7251 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_414_), .Y(u2__abc_52155_new_n15823_));
AND2X2 AND2X2_7252 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7151_), .Y(u2__abc_52155_new_n15826_));
AND2X2 AND2X2_7253 ( .A(u2__abc_52155_new_n15827_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15828_));
AND2X2 AND2X2_7254 ( .A(u2__abc_52155_new_n15825_), .B(u2__abc_52155_new_n15828_), .Y(u2__abc_52155_new_n15829_));
AND2X2 AND2X2_7255 ( .A(u2__abc_52155_new_n15830_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__416_));
AND2X2 AND2X2_7256 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_417_), .Y(u2__abc_52155_new_n15832_));
AND2X2 AND2X2_7257 ( .A(u2__abc_52155_new_n15819_), .B(u2__abc_52155_new_n7172_), .Y(u2__abc_52155_new_n15833_));
AND2X2 AND2X2_7258 ( .A(u2__abc_52155_new_n15833_), .B(u2__abc_52155_new_n7169_), .Y(u2__abc_52155_new_n15834_));
AND2X2 AND2X2_7259 ( .A(u2__abc_52155_new_n15836_), .B(u2__abc_52155_new_n15835_), .Y(u2__abc_52155_new_n15837_));
AND2X2 AND2X2_726 ( .A(u2__abc_52155_new_n3436_), .B(u2_remHi_50_), .Y(u2__abc_52155_new_n3437_));
AND2X2 AND2X2_7260 ( .A(u2__abc_52155_new_n15838_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15839_));
AND2X2 AND2X2_7261 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_415_), .Y(u2__abc_52155_new_n15840_));
AND2X2 AND2X2_7262 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7155_), .Y(u2__abc_52155_new_n15843_));
AND2X2 AND2X2_7263 ( .A(u2__abc_52155_new_n15844_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15845_));
AND2X2 AND2X2_7264 ( .A(u2__abc_52155_new_n15842_), .B(u2__abc_52155_new_n15845_), .Y(u2__abc_52155_new_n15846_));
AND2X2 AND2X2_7265 ( .A(u2__abc_52155_new_n15847_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__417_));
AND2X2 AND2X2_7266 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_418_), .Y(u2__abc_52155_new_n15849_));
AND2X2 AND2X2_7267 ( .A(u2__abc_52155_new_n7168_), .B(u2__abc_52155_new_n7172_), .Y(u2__abc_52155_new_n15850_));
AND2X2 AND2X2_7268 ( .A(u2__abc_52155_new_n15819_), .B(u2__abc_52155_new_n15850_), .Y(u2__abc_52155_new_n15851_));
AND2X2 AND2X2_7269 ( .A(u2__abc_52155_new_n15853_), .B(u2__abc_52155_new_n7154_), .Y(u2__abc_52155_new_n15854_));
AND2X2 AND2X2_727 ( .A(u2__abc_52155_new_n3439_), .B(sqrto_50_), .Y(u2__abc_52155_new_n3440_));
AND2X2 AND2X2_7270 ( .A(u2__abc_52155_new_n15856_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15857_));
AND2X2 AND2X2_7271 ( .A(u2__abc_52155_new_n15857_), .B(u2__abc_52155_new_n15855_), .Y(u2__abc_52155_new_n15858_));
AND2X2 AND2X2_7272 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_416_), .Y(u2__abc_52155_new_n15859_));
AND2X2 AND2X2_7273 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7142_), .Y(u2__abc_52155_new_n15862_));
AND2X2 AND2X2_7274 ( .A(u2__abc_52155_new_n15863_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15864_));
AND2X2 AND2X2_7275 ( .A(u2__abc_52155_new_n15861_), .B(u2__abc_52155_new_n15864_), .Y(u2__abc_52155_new_n15865_));
AND2X2 AND2X2_7276 ( .A(u2__abc_52155_new_n15866_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__418_));
AND2X2 AND2X2_7277 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_419_), .Y(u2__abc_52155_new_n15868_));
AND2X2 AND2X2_7278 ( .A(u2__abc_52155_new_n15855_), .B(u2__abc_52155_new_n7150_), .Y(u2__abc_52155_new_n15870_));
AND2X2 AND2X2_7279 ( .A(u2__abc_52155_new_n15873_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15874_));
AND2X2 AND2X2_728 ( .A(u2__abc_52155_new_n3438_), .B(u2__abc_52155_new_n3441_), .Y(u2__abc_52155_new_n3442_));
AND2X2 AND2X2_7280 ( .A(u2__abc_52155_new_n15874_), .B(u2__abc_52155_new_n15871_), .Y(u2__abc_52155_new_n15875_));
AND2X2 AND2X2_7281 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_417_), .Y(u2__abc_52155_new_n15876_));
AND2X2 AND2X2_7282 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7132_), .Y(u2__abc_52155_new_n15879_));
AND2X2 AND2X2_7283 ( .A(u2__abc_52155_new_n15880_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15881_));
AND2X2 AND2X2_7284 ( .A(u2__abc_52155_new_n15878_), .B(u2__abc_52155_new_n15881_), .Y(u2__abc_52155_new_n15882_));
AND2X2 AND2X2_7285 ( .A(u2__abc_52155_new_n15883_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__419_));
AND2X2 AND2X2_7286 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_420_), .Y(u2__abc_52155_new_n15885_));
AND2X2 AND2X2_7287 ( .A(u2__abc_52155_new_n15887_), .B(u2__abc_52155_new_n7162_), .Y(u2__abc_52155_new_n15888_));
AND2X2 AND2X2_7288 ( .A(u2__abc_52155_new_n7157_), .B(u2__abc_52155_new_n7149_), .Y(u2__abc_52155_new_n15889_));
AND2X2 AND2X2_7289 ( .A(u2__abc_52155_new_n15817_), .B(u2__abc_52155_new_n7178_), .Y(u2__abc_52155_new_n15892_));
AND2X2 AND2X2_729 ( .A(u2__abc_52155_new_n3435_), .B(u2__abc_52155_new_n3442_), .Y(u2__abc_52155_new_n3443_));
AND2X2 AND2X2_7290 ( .A(u2__abc_52155_new_n15893_), .B(u2__abc_52155_new_n7145_), .Y(u2__abc_52155_new_n15894_));
AND2X2 AND2X2_7291 ( .A(u2__abc_52155_new_n15896_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15897_));
AND2X2 AND2X2_7292 ( .A(u2__abc_52155_new_n15897_), .B(u2__abc_52155_new_n15895_), .Y(u2__abc_52155_new_n15898_));
AND2X2 AND2X2_7293 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_418_), .Y(u2__abc_52155_new_n15899_));
AND2X2 AND2X2_7294 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7120_), .Y(u2__abc_52155_new_n15902_));
AND2X2 AND2X2_7295 ( .A(u2__abc_52155_new_n15903_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15904_));
AND2X2 AND2X2_7296 ( .A(u2__abc_52155_new_n15901_), .B(u2__abc_52155_new_n15904_), .Y(u2__abc_52155_new_n15905_));
AND2X2 AND2X2_7297 ( .A(u2__abc_52155_new_n15906_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__420_));
AND2X2 AND2X2_7298 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_421_), .Y(u2__abc_52155_new_n15908_));
AND2X2 AND2X2_7299 ( .A(u2__abc_52155_new_n15895_), .B(u2__abc_52155_new_n7141_), .Y(u2__abc_52155_new_n15909_));
AND2X2 AND2X2_73 ( .A(_abc_73687_new_n753_), .B(sqrto_72_), .Y(\o[108] ));
AND2X2 AND2X2_730 ( .A(u2__abc_52155_new_n3428_), .B(u2__abc_52155_new_n3443_), .Y(u2__abc_52155_new_n3444_));
AND2X2 AND2X2_7300 ( .A(u2__abc_52155_new_n15909_), .B(u2__abc_52155_new_n7138_), .Y(u2__abc_52155_new_n15910_));
AND2X2 AND2X2_7301 ( .A(u2__abc_52155_new_n15912_), .B(u2__abc_52155_new_n15911_), .Y(u2__abc_52155_new_n15913_));
AND2X2 AND2X2_7302 ( .A(u2__abc_52155_new_n15914_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15915_));
AND2X2 AND2X2_7303 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_419_), .Y(u2__abc_52155_new_n15916_));
AND2X2 AND2X2_7304 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7127_), .Y(u2__abc_52155_new_n15919_));
AND2X2 AND2X2_7305 ( .A(u2__abc_52155_new_n15920_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15921_));
AND2X2 AND2X2_7306 ( .A(u2__abc_52155_new_n15918_), .B(u2__abc_52155_new_n15921_), .Y(u2__abc_52155_new_n15922_));
AND2X2 AND2X2_7307 ( .A(u2__abc_52155_new_n15923_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__421_));
AND2X2 AND2X2_7308 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_422_), .Y(u2__abc_52155_new_n15925_));
AND2X2 AND2X2_7309 ( .A(u2__abc_52155_new_n7137_), .B(u2__abc_52155_new_n7141_), .Y(u2__abc_52155_new_n15926_));
AND2X2 AND2X2_731 ( .A(u2__abc_52155_new_n3413_), .B(u2__abc_52155_new_n3444_), .Y(u2__abc_52155_new_n3445_));
AND2X2 AND2X2_7310 ( .A(u2__abc_52155_new_n15895_), .B(u2__abc_52155_new_n15926_), .Y(u2__abc_52155_new_n15927_));
AND2X2 AND2X2_7311 ( .A(u2__abc_52155_new_n15929_), .B(u2__abc_52155_new_n7123_), .Y(u2__abc_52155_new_n15930_));
AND2X2 AND2X2_7312 ( .A(u2__abc_52155_new_n15932_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15933_));
AND2X2 AND2X2_7313 ( .A(u2__abc_52155_new_n15933_), .B(u2__abc_52155_new_n15931_), .Y(u2__abc_52155_new_n15934_));
AND2X2 AND2X2_7314 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_420_), .Y(u2__abc_52155_new_n15935_));
AND2X2 AND2X2_7315 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7072_), .Y(u2__abc_52155_new_n15938_));
AND2X2 AND2X2_7316 ( .A(u2__abc_52155_new_n15939_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15940_));
AND2X2 AND2X2_7317 ( .A(u2__abc_52155_new_n15937_), .B(u2__abc_52155_new_n15940_), .Y(u2__abc_52155_new_n15941_));
AND2X2 AND2X2_7318 ( .A(u2__abc_52155_new_n15942_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__422_));
AND2X2 AND2X2_7319 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_423_), .Y(u2__abc_52155_new_n15944_));
AND2X2 AND2X2_732 ( .A(u2__abc_52155_new_n3445_), .B(u2__abc_52155_new_n3385_), .Y(u2__abc_52155_new_n3446_));
AND2X2 AND2X2_7320 ( .A(u2__abc_52155_new_n15931_), .B(u2__abc_52155_new_n7119_), .Y(u2__abc_52155_new_n15946_));
AND2X2 AND2X2_7321 ( .A(u2__abc_52155_new_n15949_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15950_));
AND2X2 AND2X2_7322 ( .A(u2__abc_52155_new_n15950_), .B(u2__abc_52155_new_n15947_), .Y(u2__abc_52155_new_n15951_));
AND2X2 AND2X2_7323 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_421_), .Y(u2__abc_52155_new_n15952_));
AND2X2 AND2X2_7324 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7076_), .Y(u2__abc_52155_new_n15955_));
AND2X2 AND2X2_7325 ( .A(u2__abc_52155_new_n15956_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15957_));
AND2X2 AND2X2_7326 ( .A(u2__abc_52155_new_n15954_), .B(u2__abc_52155_new_n15957_), .Y(u2__abc_52155_new_n15958_));
AND2X2 AND2X2_7327 ( .A(u2__abc_52155_new_n15959_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__423_));
AND2X2 AND2X2_7328 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_424_), .Y(u2__abc_52155_new_n15961_));
AND2X2 AND2X2_7329 ( .A(u2__abc_52155_new_n15891_), .B(u2__abc_52155_new_n7147_), .Y(u2__abc_52155_new_n15962_));
AND2X2 AND2X2_733 ( .A(u2__abc_52155_new_n3447_), .B(u2_remHi_40_), .Y(u2__abc_52155_new_n3448_));
AND2X2 AND2X2_7330 ( .A(u2__abc_52155_new_n15964_), .B(u2__abc_52155_new_n7131_), .Y(u2__abc_52155_new_n15965_));
AND2X2 AND2X2_7331 ( .A(u2__abc_52155_new_n7129_), .B(u2__abc_52155_new_n7118_), .Y(u2__abc_52155_new_n15966_));
AND2X2 AND2X2_7332 ( .A(u2__abc_52155_new_n15817_), .B(u2__abc_52155_new_n7179_), .Y(u2__abc_52155_new_n15970_));
AND2X2 AND2X2_7333 ( .A(u2__abc_52155_new_n15971_), .B(u2__abc_52155_new_n7075_), .Y(u2__abc_52155_new_n15972_));
AND2X2 AND2X2_7334 ( .A(u2__abc_52155_new_n15974_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15975_));
AND2X2 AND2X2_7335 ( .A(u2__abc_52155_new_n15975_), .B(u2__abc_52155_new_n15973_), .Y(u2__abc_52155_new_n15976_));
AND2X2 AND2X2_7336 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_422_), .Y(u2__abc_52155_new_n15977_));
AND2X2 AND2X2_7337 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7057_), .Y(u2__abc_52155_new_n15980_));
AND2X2 AND2X2_7338 ( .A(u2__abc_52155_new_n15981_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15982_));
AND2X2 AND2X2_7339 ( .A(u2__abc_52155_new_n15979_), .B(u2__abc_52155_new_n15982_), .Y(u2__abc_52155_new_n15983_));
AND2X2 AND2X2_734 ( .A(u2__abc_52155_new_n3449_), .B(sqrto_40_), .Y(u2__abc_52155_new_n3450_));
AND2X2 AND2X2_7340 ( .A(u2__abc_52155_new_n15984_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__424_));
AND2X2 AND2X2_7341 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_425_), .Y(u2__abc_52155_new_n15986_));
AND2X2 AND2X2_7342 ( .A(u2__abc_52155_new_n15973_), .B(u2__abc_52155_new_n7071_), .Y(u2__abc_52155_new_n15988_));
AND2X2 AND2X2_7343 ( .A(u2__abc_52155_new_n15989_), .B(u2__abc_52155_new_n15987_), .Y(u2__abc_52155_new_n15990_));
AND2X2 AND2X2_7344 ( .A(u2__abc_52155_new_n15988_), .B(u2__abc_52155_new_n7082_), .Y(u2__abc_52155_new_n15991_));
AND2X2 AND2X2_7345 ( .A(u2__abc_52155_new_n15992_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n15993_));
AND2X2 AND2X2_7346 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_423_), .Y(u2__abc_52155_new_n15994_));
AND2X2 AND2X2_7347 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7061_), .Y(u2__abc_52155_new_n15997_));
AND2X2 AND2X2_7348 ( .A(u2__abc_52155_new_n15998_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n15999_));
AND2X2 AND2X2_7349 ( .A(u2__abc_52155_new_n15996_), .B(u2__abc_52155_new_n15999_), .Y(u2__abc_52155_new_n16000_));
AND2X2 AND2X2_735 ( .A(u2__abc_52155_new_n3452_), .B(u2_remHi_41_), .Y(u2__abc_52155_new_n3453_));
AND2X2 AND2X2_7350 ( .A(u2__abc_52155_new_n16001_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__425_));
AND2X2 AND2X2_7351 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_426_), .Y(u2__abc_52155_new_n16003_));
AND2X2 AND2X2_7352 ( .A(u2__abc_52155_new_n15989_), .B(u2__abc_52155_new_n7078_), .Y(u2__abc_52155_new_n16004_));
AND2X2 AND2X2_7353 ( .A(u2__abc_52155_new_n16005_), .B(u2__abc_52155_new_n7060_), .Y(u2__abc_52155_new_n16006_));
AND2X2 AND2X2_7354 ( .A(u2__abc_52155_new_n16008_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16009_));
AND2X2 AND2X2_7355 ( .A(u2__abc_52155_new_n16009_), .B(u2__abc_52155_new_n16007_), .Y(u2__abc_52155_new_n16010_));
AND2X2 AND2X2_7356 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_424_), .Y(u2__abc_52155_new_n16011_));
AND2X2 AND2X2_7357 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7110_), .Y(u2__abc_52155_new_n16014_));
AND2X2 AND2X2_7358 ( .A(u2__abc_52155_new_n16015_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16016_));
AND2X2 AND2X2_7359 ( .A(u2__abc_52155_new_n16013_), .B(u2__abc_52155_new_n16016_), .Y(u2__abc_52155_new_n16017_));
AND2X2 AND2X2_736 ( .A(u2__abc_52155_new_n3454_), .B(sqrto_41_), .Y(u2__abc_52155_new_n3455_));
AND2X2 AND2X2_7360 ( .A(u2__abc_52155_new_n16018_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__426_));
AND2X2 AND2X2_7361 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_427_), .Y(u2__abc_52155_new_n16020_));
AND2X2 AND2X2_7362 ( .A(u2__abc_52155_new_n16007_), .B(u2__abc_52155_new_n7056_), .Y(u2__abc_52155_new_n16022_));
AND2X2 AND2X2_7363 ( .A(u2__abc_52155_new_n16025_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16026_));
AND2X2 AND2X2_7364 ( .A(u2__abc_52155_new_n16026_), .B(u2__abc_52155_new_n16023_), .Y(u2__abc_52155_new_n16027_));
AND2X2 AND2X2_7365 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_425_), .Y(u2__abc_52155_new_n16028_));
AND2X2 AND2X2_7366 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7100_), .Y(u2__abc_52155_new_n16031_));
AND2X2 AND2X2_7367 ( .A(u2__abc_52155_new_n16032_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16033_));
AND2X2 AND2X2_7368 ( .A(u2__abc_52155_new_n16030_), .B(u2__abc_52155_new_n16033_), .Y(u2__abc_52155_new_n16034_));
AND2X2 AND2X2_7369 ( .A(u2__abc_52155_new_n16035_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__427_));
AND2X2 AND2X2_737 ( .A(u2__abc_52155_new_n3459_), .B(u2_remHi_38_), .Y(u2__abc_52155_new_n3460_));
AND2X2 AND2X2_7370 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_428_), .Y(u2__abc_52155_new_n16037_));
AND2X2 AND2X2_7371 ( .A(u2__abc_52155_new_n7071_), .B(u2__abc_52155_new_n7081_), .Y(u2__abc_52155_new_n16038_));
AND2X2 AND2X2_7372 ( .A(u2__abc_52155_new_n16040_), .B(u2__abc_52155_new_n7068_), .Y(u2__abc_52155_new_n16041_));
AND2X2 AND2X2_7373 ( .A(u2__abc_52155_new_n7063_), .B(u2__abc_52155_new_n7055_), .Y(u2__abc_52155_new_n16042_));
AND2X2 AND2X2_7374 ( .A(u2__abc_52155_new_n15971_), .B(u2__abc_52155_new_n7084_), .Y(u2__abc_52155_new_n16045_));
AND2X2 AND2X2_7375 ( .A(u2__abc_52155_new_n16046_), .B(u2__abc_52155_new_n7113_), .Y(u2__abc_52155_new_n16047_));
AND2X2 AND2X2_7376 ( .A(u2__abc_52155_new_n16049_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16050_));
AND2X2 AND2X2_7377 ( .A(u2__abc_52155_new_n16050_), .B(u2__abc_52155_new_n16048_), .Y(u2__abc_52155_new_n16051_));
AND2X2 AND2X2_7378 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_426_), .Y(u2__abc_52155_new_n16052_));
AND2X2 AND2X2_7379 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7088_), .Y(u2__abc_52155_new_n16055_));
AND2X2 AND2X2_738 ( .A(u2__abc_52155_new_n3462_), .B(sqrto_38_), .Y(u2__abc_52155_new_n3463_));
AND2X2 AND2X2_7380 ( .A(u2__abc_52155_new_n16056_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16057_));
AND2X2 AND2X2_7381 ( .A(u2__abc_52155_new_n16054_), .B(u2__abc_52155_new_n16057_), .Y(u2__abc_52155_new_n16058_));
AND2X2 AND2X2_7382 ( .A(u2__abc_52155_new_n16059_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__428_));
AND2X2 AND2X2_7383 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_429_), .Y(u2__abc_52155_new_n16061_));
AND2X2 AND2X2_7384 ( .A(u2__abc_52155_new_n16048_), .B(u2__abc_52155_new_n7109_), .Y(u2__abc_52155_new_n16062_));
AND2X2 AND2X2_7385 ( .A(u2__abc_52155_new_n16062_), .B(u2__abc_52155_new_n7106_), .Y(u2__abc_52155_new_n16063_));
AND2X2 AND2X2_7386 ( .A(u2__abc_52155_new_n16065_), .B(u2__abc_52155_new_n16064_), .Y(u2__abc_52155_new_n16066_));
AND2X2 AND2X2_7387 ( .A(u2__abc_52155_new_n16067_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16068_));
AND2X2 AND2X2_7388 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_427_), .Y(u2__abc_52155_new_n16069_));
AND2X2 AND2X2_7389 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7095_), .Y(u2__abc_52155_new_n16072_));
AND2X2 AND2X2_739 ( .A(u2__abc_52155_new_n3461_), .B(u2__abc_52155_new_n3464_), .Y(u2__abc_52155_new_n3465_));
AND2X2 AND2X2_7390 ( .A(u2__abc_52155_new_n16073_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16074_));
AND2X2 AND2X2_7391 ( .A(u2__abc_52155_new_n16071_), .B(u2__abc_52155_new_n16074_), .Y(u2__abc_52155_new_n16075_));
AND2X2 AND2X2_7392 ( .A(u2__abc_52155_new_n16076_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__429_));
AND2X2 AND2X2_7393 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_430_), .Y(u2__abc_52155_new_n16078_));
AND2X2 AND2X2_7394 ( .A(u2__abc_52155_new_n7105_), .B(u2__abc_52155_new_n7109_), .Y(u2__abc_52155_new_n16079_));
AND2X2 AND2X2_7395 ( .A(u2__abc_52155_new_n16048_), .B(u2__abc_52155_new_n16079_), .Y(u2__abc_52155_new_n16080_));
AND2X2 AND2X2_7396 ( .A(u2__abc_52155_new_n16082_), .B(u2__abc_52155_new_n7091_), .Y(u2__abc_52155_new_n16083_));
AND2X2 AND2X2_7397 ( .A(u2__abc_52155_new_n16085_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16086_));
AND2X2 AND2X2_7398 ( .A(u2__abc_52155_new_n16086_), .B(u2__abc_52155_new_n16084_), .Y(u2__abc_52155_new_n16087_));
AND2X2 AND2X2_7399 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_428_), .Y(u2__abc_52155_new_n16088_));
AND2X2 AND2X2_74 ( .A(_abc_73687_new_n753_), .B(sqrto_73_), .Y(\o[109] ));
AND2X2 AND2X2_740 ( .A(u2__abc_52155_new_n3466_), .B(u2_remHi_39_), .Y(u2__abc_52155_new_n3467_));
AND2X2 AND2X2_7400 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7024_), .Y(u2__abc_52155_new_n16091_));
AND2X2 AND2X2_7401 ( .A(u2__abc_52155_new_n16092_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16093_));
AND2X2 AND2X2_7402 ( .A(u2__abc_52155_new_n16090_), .B(u2__abc_52155_new_n16093_), .Y(u2__abc_52155_new_n16094_));
AND2X2 AND2X2_7403 ( .A(u2__abc_52155_new_n16095_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__430_));
AND2X2 AND2X2_7404 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_431_), .Y(u2__abc_52155_new_n16097_));
AND2X2 AND2X2_7405 ( .A(u2__abc_52155_new_n16084_), .B(u2__abc_52155_new_n7087_), .Y(u2__abc_52155_new_n16099_));
AND2X2 AND2X2_7406 ( .A(u2__abc_52155_new_n16102_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16103_));
AND2X2 AND2X2_7407 ( .A(u2__abc_52155_new_n16103_), .B(u2__abc_52155_new_n16100_), .Y(u2__abc_52155_new_n16104_));
AND2X2 AND2X2_7408 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_429_), .Y(u2__abc_52155_new_n16105_));
AND2X2 AND2X2_7409 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7028_), .Y(u2__abc_52155_new_n16108_));
AND2X2 AND2X2_741 ( .A(u2__abc_52155_new_n3469_), .B(sqrto_39_), .Y(u2__abc_52155_new_n3470_));
AND2X2 AND2X2_7410 ( .A(u2__abc_52155_new_n16109_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16110_));
AND2X2 AND2X2_7411 ( .A(u2__abc_52155_new_n16107_), .B(u2__abc_52155_new_n16110_), .Y(u2__abc_52155_new_n16111_));
AND2X2 AND2X2_7412 ( .A(u2__abc_52155_new_n16112_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__431_));
AND2X2 AND2X2_7413 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_432_), .Y(u2__abc_52155_new_n16114_));
AND2X2 AND2X2_7414 ( .A(u2__abc_52155_new_n15969_), .B(u2__abc_52155_new_n7116_), .Y(u2__abc_52155_new_n16115_));
AND2X2 AND2X2_7415 ( .A(u2__abc_52155_new_n16044_), .B(u2__abc_52155_new_n7115_), .Y(u2__abc_52155_new_n16116_));
AND2X2 AND2X2_7416 ( .A(u2__abc_52155_new_n16118_), .B(u2__abc_52155_new_n7099_), .Y(u2__abc_52155_new_n16119_));
AND2X2 AND2X2_7417 ( .A(u2__abc_52155_new_n7097_), .B(u2__abc_52155_new_n7086_), .Y(u2__abc_52155_new_n16120_));
AND2X2 AND2X2_7418 ( .A(u2__abc_52155_new_n15817_), .B(u2__abc_52155_new_n7180_), .Y(u2__abc_52155_new_n16125_));
AND2X2 AND2X2_7419 ( .A(u2__abc_52155_new_n16126_), .B(u2__abc_52155_new_n7027_), .Y(u2__abc_52155_new_n16127_));
AND2X2 AND2X2_742 ( .A(u2__abc_52155_new_n3468_), .B(u2__abc_52155_new_n3471_), .Y(u2__abc_52155_new_n3472_));
AND2X2 AND2X2_7420 ( .A(u2__abc_52155_new_n16129_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16130_));
AND2X2 AND2X2_7421 ( .A(u2__abc_52155_new_n16130_), .B(u2__abc_52155_new_n16128_), .Y(u2__abc_52155_new_n16131_));
AND2X2 AND2X2_7422 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_430_), .Y(u2__abc_52155_new_n16132_));
AND2X2 AND2X2_7423 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7039_), .Y(u2__abc_52155_new_n16135_));
AND2X2 AND2X2_7424 ( .A(u2__abc_52155_new_n16136_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16137_));
AND2X2 AND2X2_7425 ( .A(u2__abc_52155_new_n16134_), .B(u2__abc_52155_new_n16137_), .Y(u2__abc_52155_new_n16138_));
AND2X2 AND2X2_7426 ( .A(u2__abc_52155_new_n16139_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__432_));
AND2X2 AND2X2_7427 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_433_), .Y(u2__abc_52155_new_n16141_));
AND2X2 AND2X2_7428 ( .A(u2__abc_52155_new_n16128_), .B(u2__abc_52155_new_n7023_), .Y(u2__abc_52155_new_n16143_));
AND2X2 AND2X2_7429 ( .A(u2__abc_52155_new_n16146_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16147_));
AND2X2 AND2X2_743 ( .A(u2__abc_52155_new_n3465_), .B(u2__abc_52155_new_n3472_), .Y(u2__abc_52155_new_n3473_));
AND2X2 AND2X2_7430 ( .A(u2__abc_52155_new_n16147_), .B(u2__abc_52155_new_n16144_), .Y(u2__abc_52155_new_n16148_));
AND2X2 AND2X2_7431 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_431_), .Y(u2__abc_52155_new_n16149_));
AND2X2 AND2X2_7432 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7043_), .Y(u2__abc_52155_new_n16152_));
AND2X2 AND2X2_7433 ( .A(u2__abc_52155_new_n16153_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16154_));
AND2X2 AND2X2_7434 ( .A(u2__abc_52155_new_n16151_), .B(u2__abc_52155_new_n16154_), .Y(u2__abc_52155_new_n16155_));
AND2X2 AND2X2_7435 ( .A(u2__abc_52155_new_n16156_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__433_));
AND2X2 AND2X2_7436 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_434_), .Y(u2__abc_52155_new_n16158_));
AND2X2 AND2X2_7437 ( .A(u2__abc_52155_new_n16159_), .B(u2__abc_52155_new_n7033_), .Y(u2__abc_52155_new_n16160_));
AND2X2 AND2X2_7438 ( .A(u2__abc_52155_new_n16126_), .B(u2__abc_52155_new_n7035_), .Y(u2__abc_52155_new_n16162_));
AND2X2 AND2X2_7439 ( .A(u2__abc_52155_new_n16163_), .B(u2__abc_52155_new_n7042_), .Y(u2__abc_52155_new_n16164_));
AND2X2 AND2X2_744 ( .A(u2__abc_52155_new_n3458_), .B(u2__abc_52155_new_n3473_), .Y(u2__abc_52155_new_n3474_));
AND2X2 AND2X2_7440 ( .A(u2__abc_52155_new_n16166_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16167_));
AND2X2 AND2X2_7441 ( .A(u2__abc_52155_new_n16167_), .B(u2__abc_52155_new_n16165_), .Y(u2__abc_52155_new_n16168_));
AND2X2 AND2X2_7442 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_432_), .Y(u2__abc_52155_new_n16169_));
AND2X2 AND2X2_7443 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7015_), .Y(u2__abc_52155_new_n16172_));
AND2X2 AND2X2_7444 ( .A(u2__abc_52155_new_n16173_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16174_));
AND2X2 AND2X2_7445 ( .A(u2__abc_52155_new_n16171_), .B(u2__abc_52155_new_n16174_), .Y(u2__abc_52155_new_n16175_));
AND2X2 AND2X2_7446 ( .A(u2__abc_52155_new_n16176_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__434_));
AND2X2 AND2X2_7447 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_435_), .Y(u2__abc_52155_new_n16178_));
AND2X2 AND2X2_7448 ( .A(u2__abc_52155_new_n16165_), .B(u2__abc_52155_new_n7038_), .Y(u2__abc_52155_new_n16180_));
AND2X2 AND2X2_7449 ( .A(u2__abc_52155_new_n16183_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16184_));
AND2X2 AND2X2_745 ( .A(u2__abc_52155_new_n3475_), .B(u2_remHi_44_), .Y(u2__abc_52155_new_n3476_));
AND2X2 AND2X2_7450 ( .A(u2__abc_52155_new_n16184_), .B(u2__abc_52155_new_n16181_), .Y(u2__abc_52155_new_n16185_));
AND2X2 AND2X2_7451 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_433_), .Y(u2__abc_52155_new_n16186_));
AND2X2 AND2X2_7452 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7005_), .Y(u2__abc_52155_new_n16189_));
AND2X2 AND2X2_7453 ( .A(u2__abc_52155_new_n16190_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16191_));
AND2X2 AND2X2_7454 ( .A(u2__abc_52155_new_n16188_), .B(u2__abc_52155_new_n16191_), .Y(u2__abc_52155_new_n16192_));
AND2X2 AND2X2_7455 ( .A(u2__abc_52155_new_n16193_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__435_));
AND2X2 AND2X2_7456 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_436_), .Y(u2__abc_52155_new_n16195_));
AND2X2 AND2X2_7457 ( .A(u2__abc_52155_new_n7038_), .B(u2__abc_52155_new_n7048_), .Y(u2__abc_52155_new_n16196_));
AND2X2 AND2X2_7458 ( .A(u2__abc_52155_new_n16165_), .B(u2__abc_52155_new_n16196_), .Y(u2__abc_52155_new_n16197_));
AND2X2 AND2X2_7459 ( .A(u2__abc_52155_new_n16199_), .B(u2__abc_52155_new_n7018_), .Y(u2__abc_52155_new_n16200_));
AND2X2 AND2X2_746 ( .A(u2__abc_52155_new_n3478_), .B(sqrto_44_), .Y(u2__abc_52155_new_n3479_));
AND2X2 AND2X2_7460 ( .A(u2__abc_52155_new_n16202_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16203_));
AND2X2 AND2X2_7461 ( .A(u2__abc_52155_new_n16203_), .B(u2__abc_52155_new_n16201_), .Y(u2__abc_52155_new_n16204_));
AND2X2 AND2X2_7462 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_434_), .Y(u2__abc_52155_new_n16205_));
AND2X2 AND2X2_7463 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6993_), .Y(u2__abc_52155_new_n16208_));
AND2X2 AND2X2_7464 ( .A(u2__abc_52155_new_n16209_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16210_));
AND2X2 AND2X2_7465 ( .A(u2__abc_52155_new_n16207_), .B(u2__abc_52155_new_n16210_), .Y(u2__abc_52155_new_n16211_));
AND2X2 AND2X2_7466 ( .A(u2__abc_52155_new_n16212_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__436_));
AND2X2 AND2X2_7467 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_437_), .Y(u2__abc_52155_new_n16214_));
AND2X2 AND2X2_7468 ( .A(u2__abc_52155_new_n16201_), .B(u2__abc_52155_new_n7014_), .Y(u2__abc_52155_new_n16215_));
AND2X2 AND2X2_7469 ( .A(u2__abc_52155_new_n16216_), .B(u2__abc_52155_new_n7011_), .Y(u2__abc_52155_new_n16217_));
AND2X2 AND2X2_747 ( .A(u2__abc_52155_new_n3477_), .B(u2__abc_52155_new_n3480_), .Y(u2__abc_52155_new_n3481_));
AND2X2 AND2X2_7470 ( .A(u2__abc_52155_new_n16219_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16220_));
AND2X2 AND2X2_7471 ( .A(u2__abc_52155_new_n16220_), .B(u2__abc_52155_new_n16218_), .Y(u2__abc_52155_new_n16221_));
AND2X2 AND2X2_7472 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_435_), .Y(u2__abc_52155_new_n16222_));
AND2X2 AND2X2_7473 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n7000_), .Y(u2__abc_52155_new_n16225_));
AND2X2 AND2X2_7474 ( .A(u2__abc_52155_new_n16226_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16227_));
AND2X2 AND2X2_7475 ( .A(u2__abc_52155_new_n16224_), .B(u2__abc_52155_new_n16227_), .Y(u2__abc_52155_new_n16228_));
AND2X2 AND2X2_7476 ( .A(u2__abc_52155_new_n16229_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__437_));
AND2X2 AND2X2_7477 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_438_), .Y(u2__abc_52155_new_n16231_));
AND2X2 AND2X2_7478 ( .A(u2__abc_52155_new_n16218_), .B(u2__abc_52155_new_n7010_), .Y(u2__abc_52155_new_n16232_));
AND2X2 AND2X2_7479 ( .A(u2__abc_52155_new_n16233_), .B(u2__abc_52155_new_n6996_), .Y(u2__abc_52155_new_n16234_));
AND2X2 AND2X2_748 ( .A(u2__abc_52155_new_n3482_), .B(u2_remHi_45_), .Y(u2__abc_52155_new_n3483_));
AND2X2 AND2X2_7480 ( .A(u2__abc_52155_new_n16236_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16237_));
AND2X2 AND2X2_7481 ( .A(u2__abc_52155_new_n16237_), .B(u2__abc_52155_new_n16235_), .Y(u2__abc_52155_new_n16238_));
AND2X2 AND2X2_7482 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_436_), .Y(u2__abc_52155_new_n16239_));
AND2X2 AND2X2_7483 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6961_), .Y(u2__abc_52155_new_n16242_));
AND2X2 AND2X2_7484 ( .A(u2__abc_52155_new_n16243_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16244_));
AND2X2 AND2X2_7485 ( .A(u2__abc_52155_new_n16241_), .B(u2__abc_52155_new_n16244_), .Y(u2__abc_52155_new_n16245_));
AND2X2 AND2X2_7486 ( .A(u2__abc_52155_new_n16246_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__438_));
AND2X2 AND2X2_7487 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_439_), .Y(u2__abc_52155_new_n16248_));
AND2X2 AND2X2_7488 ( .A(u2__abc_52155_new_n16235_), .B(u2__abc_52155_new_n6992_), .Y(u2__abc_52155_new_n16250_));
AND2X2 AND2X2_7489 ( .A(u2__abc_52155_new_n16253_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16254_));
AND2X2 AND2X2_749 ( .A(u2__abc_52155_new_n3485_), .B(sqrto_45_), .Y(u2__abc_52155_new_n3486_));
AND2X2 AND2X2_7490 ( .A(u2__abc_52155_new_n16254_), .B(u2__abc_52155_new_n16251_), .Y(u2__abc_52155_new_n16255_));
AND2X2 AND2X2_7491 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_437_), .Y(u2__abc_52155_new_n16256_));
AND2X2 AND2X2_7492 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6965_), .Y(u2__abc_52155_new_n16259_));
AND2X2 AND2X2_7493 ( .A(u2__abc_52155_new_n16260_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16261_));
AND2X2 AND2X2_7494 ( .A(u2__abc_52155_new_n16258_), .B(u2__abc_52155_new_n16261_), .Y(u2__abc_52155_new_n16262_));
AND2X2 AND2X2_7495 ( .A(u2__abc_52155_new_n16263_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__439_));
AND2X2 AND2X2_7496 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_440_), .Y(u2__abc_52155_new_n16265_));
AND2X2 AND2X2_7497 ( .A(u2__abc_52155_new_n16161_), .B(u2__abc_52155_new_n7050_), .Y(u2__abc_52155_new_n16267_));
AND2X2 AND2X2_7498 ( .A(u2__abc_52155_new_n16268_), .B(u2__abc_52155_new_n16266_), .Y(u2__abc_52155_new_n16269_));
AND2X2 AND2X2_7499 ( .A(u2__abc_52155_new_n16270_), .B(u2__abc_52155_new_n7020_), .Y(u2__abc_52155_new_n16271_));
AND2X2 AND2X2_75 ( .A(_abc_73687_new_n753_), .B(sqrto_74_), .Y(\o[110] ));
AND2X2 AND2X2_750 ( .A(u2__abc_52155_new_n3484_), .B(u2__abc_52155_new_n3487_), .Y(u2__abc_52155_new_n3488_));
AND2X2 AND2X2_7500 ( .A(u2__abc_52155_new_n7010_), .B(u2__abc_52155_new_n7014_), .Y(u2__abc_52155_new_n16272_));
AND2X2 AND2X2_7501 ( .A(u2__abc_52155_new_n16274_), .B(u2__abc_52155_new_n7004_), .Y(u2__abc_52155_new_n16275_));
AND2X2 AND2X2_7502 ( .A(u2__abc_52155_new_n7002_), .B(u2__abc_52155_new_n6991_), .Y(u2__abc_52155_new_n16276_));
AND2X2 AND2X2_7503 ( .A(u2__abc_52155_new_n16126_), .B(u2__abc_52155_new_n7052_), .Y(u2__abc_52155_new_n16280_));
AND2X2 AND2X2_7504 ( .A(u2__abc_52155_new_n16281_), .B(u2__abc_52155_new_n6964_), .Y(u2__abc_52155_new_n16282_));
AND2X2 AND2X2_7505 ( .A(u2__abc_52155_new_n16284_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16285_));
AND2X2 AND2X2_7506 ( .A(u2__abc_52155_new_n16285_), .B(u2__abc_52155_new_n16283_), .Y(u2__abc_52155_new_n16286_));
AND2X2 AND2X2_7507 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_438_), .Y(u2__abc_52155_new_n16287_));
AND2X2 AND2X2_7508 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6976_), .Y(u2__abc_52155_new_n16290_));
AND2X2 AND2X2_7509 ( .A(u2__abc_52155_new_n16291_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16292_));
AND2X2 AND2X2_751 ( .A(u2__abc_52155_new_n3481_), .B(u2__abc_52155_new_n3488_), .Y(u2__abc_52155_new_n3489_));
AND2X2 AND2X2_7510 ( .A(u2__abc_52155_new_n16289_), .B(u2__abc_52155_new_n16292_), .Y(u2__abc_52155_new_n16293_));
AND2X2 AND2X2_7511 ( .A(u2__abc_52155_new_n16294_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__440_));
AND2X2 AND2X2_7512 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_441_), .Y(u2__abc_52155_new_n16296_));
AND2X2 AND2X2_7513 ( .A(u2__abc_52155_new_n16283_), .B(u2__abc_52155_new_n6960_), .Y(u2__abc_52155_new_n16298_));
AND2X2 AND2X2_7514 ( .A(u2__abc_52155_new_n16301_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16302_));
AND2X2 AND2X2_7515 ( .A(u2__abc_52155_new_n16302_), .B(u2__abc_52155_new_n16299_), .Y(u2__abc_52155_new_n16303_));
AND2X2 AND2X2_7516 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_439_), .Y(u2__abc_52155_new_n16304_));
AND2X2 AND2X2_7517 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6980_), .Y(u2__abc_52155_new_n16307_));
AND2X2 AND2X2_7518 ( .A(u2__abc_52155_new_n16308_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16309_));
AND2X2 AND2X2_7519 ( .A(u2__abc_52155_new_n16306_), .B(u2__abc_52155_new_n16309_), .Y(u2__abc_52155_new_n16310_));
AND2X2 AND2X2_752 ( .A(u2__abc_52155_new_n3490_), .B(u2_remHi_43_), .Y(u2__abc_52155_new_n3491_));
AND2X2 AND2X2_7520 ( .A(u2__abc_52155_new_n16311_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__441_));
AND2X2 AND2X2_7521 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_442_), .Y(u2__abc_52155_new_n16313_));
AND2X2 AND2X2_7522 ( .A(u2__abc_52155_new_n16314_), .B(u2__abc_52155_new_n6970_), .Y(u2__abc_52155_new_n16315_));
AND2X2 AND2X2_7523 ( .A(u2__abc_52155_new_n16281_), .B(u2__abc_52155_new_n6972_), .Y(u2__abc_52155_new_n16317_));
AND2X2 AND2X2_7524 ( .A(u2__abc_52155_new_n16318_), .B(u2__abc_52155_new_n6979_), .Y(u2__abc_52155_new_n16319_));
AND2X2 AND2X2_7525 ( .A(u2__abc_52155_new_n16321_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16322_));
AND2X2 AND2X2_7526 ( .A(u2__abc_52155_new_n16322_), .B(u2__abc_52155_new_n16320_), .Y(u2__abc_52155_new_n16323_));
AND2X2 AND2X2_7527 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_440_), .Y(u2__abc_52155_new_n16324_));
AND2X2 AND2X2_7528 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6952_), .Y(u2__abc_52155_new_n16327_));
AND2X2 AND2X2_7529 ( .A(u2__abc_52155_new_n16328_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16329_));
AND2X2 AND2X2_753 ( .A(u2__abc_52155_new_n3493_), .B(sqrto_43_), .Y(u2__abc_52155_new_n3494_));
AND2X2 AND2X2_7530 ( .A(u2__abc_52155_new_n16326_), .B(u2__abc_52155_new_n16329_), .Y(u2__abc_52155_new_n16330_));
AND2X2 AND2X2_7531 ( .A(u2__abc_52155_new_n16331_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__442_));
AND2X2 AND2X2_7532 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_443_), .Y(u2__abc_52155_new_n16333_));
AND2X2 AND2X2_7533 ( .A(u2__abc_52155_new_n16320_), .B(u2__abc_52155_new_n6975_), .Y(u2__abc_52155_new_n16335_));
AND2X2 AND2X2_7534 ( .A(u2__abc_52155_new_n16338_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16339_));
AND2X2 AND2X2_7535 ( .A(u2__abc_52155_new_n16339_), .B(u2__abc_52155_new_n16336_), .Y(u2__abc_52155_new_n16340_));
AND2X2 AND2X2_7536 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_441_), .Y(u2__abc_52155_new_n16341_));
AND2X2 AND2X2_7537 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6942_), .Y(u2__abc_52155_new_n16344_));
AND2X2 AND2X2_7538 ( .A(u2__abc_52155_new_n16345_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16346_));
AND2X2 AND2X2_7539 ( .A(u2__abc_52155_new_n16343_), .B(u2__abc_52155_new_n16346_), .Y(u2__abc_52155_new_n16347_));
AND2X2 AND2X2_754 ( .A(u2__abc_52155_new_n3492_), .B(u2__abc_52155_new_n3495_), .Y(u2__abc_52155_new_n3496_));
AND2X2 AND2X2_7540 ( .A(u2__abc_52155_new_n16348_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__443_));
AND2X2 AND2X2_7541 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_444_), .Y(u2__abc_52155_new_n16350_));
AND2X2 AND2X2_7542 ( .A(u2__abc_52155_new_n16316_), .B(u2__abc_52155_new_n6987_), .Y(u2__abc_52155_new_n16351_));
AND2X2 AND2X2_7543 ( .A(u2__abc_52155_new_n6982_), .B(u2__abc_52155_new_n6974_), .Y(u2__abc_52155_new_n16352_));
AND2X2 AND2X2_7544 ( .A(u2__abc_52155_new_n16281_), .B(u2__abc_52155_new_n6988_), .Y(u2__abc_52155_new_n16355_));
AND2X2 AND2X2_7545 ( .A(u2__abc_52155_new_n16356_), .B(u2__abc_52155_new_n6955_), .Y(u2__abc_52155_new_n16357_));
AND2X2 AND2X2_7546 ( .A(u2__abc_52155_new_n16359_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16360_));
AND2X2 AND2X2_7547 ( .A(u2__abc_52155_new_n16360_), .B(u2__abc_52155_new_n16358_), .Y(u2__abc_52155_new_n16361_));
AND2X2 AND2X2_7548 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_442_), .Y(u2__abc_52155_new_n16362_));
AND2X2 AND2X2_7549 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6930_), .Y(u2__abc_52155_new_n16365_));
AND2X2 AND2X2_755 ( .A(u2__abc_52155_new_n3497_), .B(u2_remHi_42_), .Y(u2__abc_52155_new_n3498_));
AND2X2 AND2X2_7550 ( .A(u2__abc_52155_new_n16366_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16367_));
AND2X2 AND2X2_7551 ( .A(u2__abc_52155_new_n16364_), .B(u2__abc_52155_new_n16367_), .Y(u2__abc_52155_new_n16368_));
AND2X2 AND2X2_7552 ( .A(u2__abc_52155_new_n16369_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__444_));
AND2X2 AND2X2_7553 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_445_), .Y(u2__abc_52155_new_n16371_));
AND2X2 AND2X2_7554 ( .A(u2__abc_52155_new_n16358_), .B(u2__abc_52155_new_n6951_), .Y(u2__abc_52155_new_n16372_));
AND2X2 AND2X2_7555 ( .A(u2__abc_52155_new_n16372_), .B(u2__abc_52155_new_n6948_), .Y(u2__abc_52155_new_n16373_));
AND2X2 AND2X2_7556 ( .A(u2__abc_52155_new_n16375_), .B(u2__abc_52155_new_n16374_), .Y(u2__abc_52155_new_n16376_));
AND2X2 AND2X2_7557 ( .A(u2__abc_52155_new_n16377_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16378_));
AND2X2 AND2X2_7558 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_443_), .Y(u2__abc_52155_new_n16379_));
AND2X2 AND2X2_7559 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n6934_), .Y(u2__abc_52155_new_n16382_));
AND2X2 AND2X2_756 ( .A(u2__abc_52155_new_n3500_), .B(sqrto_42_), .Y(u2__abc_52155_new_n3501_));
AND2X2 AND2X2_7560 ( .A(u2__abc_52155_new_n16383_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16384_));
AND2X2 AND2X2_7561 ( .A(u2__abc_52155_new_n16381_), .B(u2__abc_52155_new_n16384_), .Y(u2__abc_52155_new_n16385_));
AND2X2 AND2X2_7562 ( .A(u2__abc_52155_new_n16386_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__445_));
AND2X2 AND2X2_7563 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_446_), .Y(u2__abc_52155_new_n16388_));
AND2X2 AND2X2_7564 ( .A(u2__abc_52155_new_n6947_), .B(u2__abc_52155_new_n6951_), .Y(u2__abc_52155_new_n16389_));
AND2X2 AND2X2_7565 ( .A(u2__abc_52155_new_n16358_), .B(u2__abc_52155_new_n16389_), .Y(u2__abc_52155_new_n16390_));
AND2X2 AND2X2_7566 ( .A(u2__abc_52155_new_n16392_), .B(u2__abc_52155_new_n6933_), .Y(u2__abc_52155_new_n16393_));
AND2X2 AND2X2_7567 ( .A(u2__abc_52155_new_n16395_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16396_));
AND2X2 AND2X2_7568 ( .A(u2__abc_52155_new_n16396_), .B(u2__abc_52155_new_n16394_), .Y(u2__abc_52155_new_n16397_));
AND2X2 AND2X2_7569 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_444_), .Y(u2__abc_52155_new_n16398_));
AND2X2 AND2X2_757 ( .A(u2__abc_52155_new_n3499_), .B(u2__abc_52155_new_n3502_), .Y(u2__abc_52155_new_n3503_));
AND2X2 AND2X2_7570 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3028_), .Y(u2__abc_52155_new_n16401_));
AND2X2 AND2X2_7571 ( .A(u2__abc_52155_new_n16402_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16403_));
AND2X2 AND2X2_7572 ( .A(u2__abc_52155_new_n16400_), .B(u2__abc_52155_new_n16403_), .Y(u2__abc_52155_new_n16404_));
AND2X2 AND2X2_7573 ( .A(u2__abc_52155_new_n16405_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__446_));
AND2X2 AND2X2_7574 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_447_), .Y(u2__abc_52155_new_n16407_));
AND2X2 AND2X2_7575 ( .A(u2__abc_52155_new_n16394_), .B(u2__abc_52155_new_n6929_), .Y(u2__abc_52155_new_n16409_));
AND2X2 AND2X2_7576 ( .A(u2__abc_52155_new_n16412_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16413_));
AND2X2 AND2X2_7577 ( .A(u2__abc_52155_new_n16413_), .B(u2__abc_52155_new_n16410_), .Y(u2__abc_52155_new_n16414_));
AND2X2 AND2X2_7578 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_445_), .Y(u2__abc_52155_new_n16415_));
AND2X2 AND2X2_7579 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3021_), .Y(u2__abc_52155_new_n16418_));
AND2X2 AND2X2_758 ( .A(u2__abc_52155_new_n3496_), .B(u2__abc_52155_new_n3503_), .Y(u2__abc_52155_new_n3504_));
AND2X2 AND2X2_7580 ( .A(u2__abc_52155_new_n16419_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16420_));
AND2X2 AND2X2_7581 ( .A(u2__abc_52155_new_n16417_), .B(u2__abc_52155_new_n16420_), .Y(u2__abc_52155_new_n16421_));
AND2X2 AND2X2_7582 ( .A(u2__abc_52155_new_n16422_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__447_));
AND2X2 AND2X2_7583 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_448_), .Y(u2__abc_52155_new_n16424_));
AND2X2 AND2X2_7584 ( .A(u2__abc_52155_new_n15817_), .B(u2__abc_52155_new_n7181_), .Y(u2__abc_52155_new_n16425_));
AND2X2 AND2X2_7585 ( .A(u2__abc_52155_new_n16124_), .B(u2__abc_52155_new_n7053_), .Y(u2__abc_52155_new_n16426_));
AND2X2 AND2X2_7586 ( .A(u2__abc_52155_new_n16279_), .B(u2__abc_52155_new_n6989_), .Y(u2__abc_52155_new_n16427_));
AND2X2 AND2X2_7587 ( .A(u2__abc_52155_new_n16354_), .B(u2__abc_52155_new_n6957_), .Y(u2__abc_52155_new_n16428_));
AND2X2 AND2X2_7588 ( .A(u2__abc_52155_new_n6936_), .B(u2__abc_52155_new_n6928_), .Y(u2__abc_52155_new_n16429_));
AND2X2 AND2X2_7589 ( .A(u2__abc_52155_new_n16432_), .B(u2__abc_52155_new_n6941_), .Y(u2__abc_52155_new_n16433_));
AND2X2 AND2X2_759 ( .A(u2__abc_52155_new_n3489_), .B(u2__abc_52155_new_n3504_), .Y(u2__abc_52155_new_n3505_));
AND2X2 AND2X2_7590 ( .A(u2__abc_52155_new_n16438_), .B(u2__abc_52155_new_n3031_), .Y(u2__abc_52155_new_n16439_));
AND2X2 AND2X2_7591 ( .A(u2__abc_52155_new_n16441_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16442_));
AND2X2 AND2X2_7592 ( .A(u2__abc_52155_new_n16442_), .B(u2__abc_52155_new_n16440_), .Y(u2__abc_52155_new_n16443_));
AND2X2 AND2X2_7593 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_446_), .Y(u2__abc_52155_new_n16444_));
AND2X2 AND2X2_7594 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3011_), .Y(u2__abc_52155_new_n16447_));
AND2X2 AND2X2_7595 ( .A(u2__abc_52155_new_n16448_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16449_));
AND2X2 AND2X2_7596 ( .A(u2__abc_52155_new_n16446_), .B(u2__abc_52155_new_n16449_), .Y(u2__abc_52155_new_n16450_));
AND2X2 AND2X2_7597 ( .A(u2__abc_52155_new_n16451_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__448_));
AND2X2 AND2X2_7598 ( .A(u2__abc_52155_new_n3002_), .B(u2_remHi_449_), .Y(u2__abc_52155_new_n16453_));
AND2X2 AND2X2_7599 ( .A(u2__abc_52155_new_n16440_), .B(u2__abc_52155_new_n3027_), .Y(u2__abc_52155_new_n16455_));
AND2X2 AND2X2_76 ( .A(_abc_73687_new_n753_), .B(sqrto_75_), .Y(\o[111] ));
AND2X2 AND2X2_760 ( .A(u2__abc_52155_new_n3474_), .B(u2__abc_52155_new_n3505_), .Y(u2__abc_52155_new_n3506_));
AND2X2 AND2X2_7600 ( .A(u2__abc_52155_new_n16458_), .B(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n16459_));
AND2X2 AND2X2_7601 ( .A(u2__abc_52155_new_n16459_), .B(u2__abc_52155_new_n16456_), .Y(u2__abc_52155_new_n16460_));
AND2X2 AND2X2_7602 ( .A(u2__abc_52155_new_n7623_), .B(u2_remHi_447_), .Y(u2__abc_52155_new_n16461_));
AND2X2 AND2X2_7603 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3004_), .Y(u2__abc_52155_new_n16464_));
AND2X2 AND2X2_7604 ( .A(u2__abc_52155_new_n16465_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n16466_));
AND2X2 AND2X2_7605 ( .A(u2__abc_52155_new_n16463_), .B(u2__abc_52155_new_n16466_), .Y(u2__abc_52155_new_n16467_));
AND2X2 AND2X2_7606 ( .A(u2__abc_52155_new_n16468_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remHi_451_0__449_));
AND2X2 AND2X2_7607 ( .A(u2__abc_52155_new_n16471_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16472_));
AND2X2 AND2X2_7608 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16472_), .Y(u2__abc_52155_new_n16473_));
AND2X2 AND2X2_7609 ( .A(u2__abc_52155_new_n16474_), .B(u2__abc_52155_new_n16475_), .Y(u2__0cnt_7_0__0_));
AND2X2 AND2X2_761 ( .A(u2__abc_52155_new_n3507_), .B(u2_remHi_32_), .Y(u2__abc_52155_new_n3508_));
AND2X2 AND2X2_7610 ( .A(u2__abc_52155_new_n2989_), .B(u2_cnt_1_), .Y(u2__abc_52155_new_n16477_));
AND2X2 AND2X2_7611 ( .A(u2__abc_52155_new_n16478_), .B(u2_cnt_0_), .Y(u2__abc_52155_new_n16479_));
AND2X2 AND2X2_7612 ( .A(u2__abc_52155_new_n16480_), .B(u2__abc_52155_new_n16472_), .Y(u2__abc_52155_new_n16481_));
AND2X2 AND2X2_7613 ( .A(u2_cnt_0_), .B(u2_cnt_1_), .Y(u2__abc_52155_new_n16484_));
AND2X2 AND2X2_7614 ( .A(u2__abc_52155_new_n16484_), .B(u2_cnt_2_), .Y(u2__abc_52155_new_n16485_));
AND2X2 AND2X2_7615 ( .A(u2__abc_52155_new_n16487_), .B(u2__abc_52155_new_n16471_), .Y(u2__abc_52155_new_n16488_));
AND2X2 AND2X2_7616 ( .A(u2__abc_52155_new_n16488_), .B(u2__abc_52155_new_n16486_), .Y(u2__abc_52155_new_n16489_));
AND2X2 AND2X2_7617 ( .A(u2__abc_52155_new_n16490_), .B(u2__abc_52155_new_n16483_), .Y(u2__0cnt_7_0__2_));
AND2X2 AND2X2_7618 ( .A(u2__abc_52155_new_n16485_), .B(ce), .Y(u2__abc_52155_new_n16492_));
AND2X2 AND2X2_7619 ( .A(u2__abc_52155_new_n16492_), .B(u2_cnt_3_), .Y(u2__abc_52155_new_n16493_));
AND2X2 AND2X2_762 ( .A(u2__abc_52155_new_n3509_), .B(sqrto_32_), .Y(u2__abc_52155_new_n3510_));
AND2X2 AND2X2_7620 ( .A(u2__abc_52155_new_n16496_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n16497_));
AND2X2 AND2X2_7621 ( .A(u2__abc_52155_new_n16495_), .B(u2__abc_52155_new_n16497_), .Y(u2__abc_52155_new_n16498_));
AND2X2 AND2X2_7622 ( .A(u2__abc_52155_new_n16498_), .B(u2__abc_52155_new_n16494_), .Y(u2__0cnt_7_0__3_));
AND2X2 AND2X2_7623 ( .A(u2__abc_52155_new_n16493_), .B(u2_cnt_4_), .Y(u2__abc_52155_new_n16500_));
AND2X2 AND2X2_7624 ( .A(u2__abc_52155_new_n16502_), .B(u2__abc_52155_new_n16497_), .Y(u2__abc_52155_new_n16503_));
AND2X2 AND2X2_7625 ( .A(u2__abc_52155_new_n16503_), .B(u2__abc_52155_new_n16501_), .Y(u2__0cnt_7_0__4_));
AND2X2 AND2X2_7626 ( .A(u2__abc_52155_new_n16500_), .B(u2_cnt_5_), .Y(u2__abc_52155_new_n16505_));
AND2X2 AND2X2_7627 ( .A(u2__abc_52155_new_n16507_), .B(u2__abc_52155_new_n16497_), .Y(u2__abc_52155_new_n16508_));
AND2X2 AND2X2_7628 ( .A(u2__abc_52155_new_n16508_), .B(u2__abc_52155_new_n16506_), .Y(u2__0cnt_7_0__5_));
AND2X2 AND2X2_7629 ( .A(u2__abc_52155_new_n16500_), .B(u2__abc_52155_new_n2967_), .Y(u2__abc_52155_new_n16511_));
AND2X2 AND2X2_763 ( .A(u2__abc_52155_new_n3512_), .B(u2_remHi_33_), .Y(u2__abc_52155_new_n3513_));
AND2X2 AND2X2_7630 ( .A(u2__abc_52155_new_n16512_), .B(u2__abc_52155_new_n16496_), .Y(u2__abc_52155_new_n16513_));
AND2X2 AND2X2_7631 ( .A(u2__abc_52155_new_n16513_), .B(u2__abc_52155_new_n16510_), .Y(u2__abc_52155_new_n16514_));
AND2X2 AND2X2_7632 ( .A(u2__abc_52155_new_n16511_), .B(u2_cnt_7_), .Y(u2__abc_52155_new_n16516_));
AND2X2 AND2X2_7633 ( .A(u2__abc_52155_new_n16518_), .B(u2__abc_52155_new_n16496_), .Y(u2__abc_52155_new_n16519_));
AND2X2 AND2X2_7634 ( .A(u2__abc_52155_new_n16519_), .B(u2__abc_52155_new_n16517_), .Y(u2__abc_52155_new_n16520_));
AND2X2 AND2X2_7635 ( .A(u2__abc_52155_new_n2962_), .B(u2_remLo_0_), .Y(u2__abc_52155_new_n16523_));
AND2X2 AND2X2_7636 ( .A(u2__abc_52155_new_n16522_), .B(u2__abc_52155_new_n16523_), .Y(u2__0remLo_451_0__0_));
AND2X2 AND2X2_7637 ( .A(u2__abc_52155_new_n2962_), .B(u2_remLo_1_), .Y(u2__abc_52155_new_n16525_));
AND2X2 AND2X2_7638 ( .A(u2__abc_52155_new_n16522_), .B(u2__abc_52155_new_n16525_), .Y(u2__0remLo_451_0__1_));
AND2X2 AND2X2_7639 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_2_), .Y(u2__abc_52155_new_n16527_));
AND2X2 AND2X2_764 ( .A(u2__abc_52155_new_n3514_), .B(sqrto_33_), .Y(u2__abc_52155_new_n3515_));
AND2X2 AND2X2_7640 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_0_), .Y(u2__abc_52155_new_n16528_));
AND2X2 AND2X2_7641 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16528_), .Y(u2__abc_52155_new_n16529_));
AND2X2 AND2X2_7642 ( .A(u2__abc_52155_new_n16530_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__2_));
AND2X2 AND2X2_7643 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_3_), .Y(u2__abc_52155_new_n16532_));
AND2X2 AND2X2_7644 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_1_), .Y(u2__abc_52155_new_n16533_));
AND2X2 AND2X2_7645 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16533_), .Y(u2__abc_52155_new_n16534_));
AND2X2 AND2X2_7646 ( .A(u2__abc_52155_new_n16535_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__3_));
AND2X2 AND2X2_7647 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_4_), .Y(u2__abc_52155_new_n16537_));
AND2X2 AND2X2_7648 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_2_), .Y(u2__abc_52155_new_n16538_));
AND2X2 AND2X2_7649 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16538_), .Y(u2__abc_52155_new_n16539_));
AND2X2 AND2X2_765 ( .A(u2__abc_52155_new_n3519_), .B(u2_remHi_30_), .Y(u2__abc_52155_new_n3520_));
AND2X2 AND2X2_7650 ( .A(u2__abc_52155_new_n16540_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__4_));
AND2X2 AND2X2_7651 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_5_), .Y(u2__abc_52155_new_n16542_));
AND2X2 AND2X2_7652 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_3_), .Y(u2__abc_52155_new_n16543_));
AND2X2 AND2X2_7653 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16543_), .Y(u2__abc_52155_new_n16544_));
AND2X2 AND2X2_7654 ( .A(u2__abc_52155_new_n16545_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__5_));
AND2X2 AND2X2_7655 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_6_), .Y(u2__abc_52155_new_n16547_));
AND2X2 AND2X2_7656 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_4_), .Y(u2__abc_52155_new_n16548_));
AND2X2 AND2X2_7657 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16548_), .Y(u2__abc_52155_new_n16549_));
AND2X2 AND2X2_7658 ( .A(u2__abc_52155_new_n16550_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__6_));
AND2X2 AND2X2_7659 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_7_), .Y(u2__abc_52155_new_n16552_));
AND2X2 AND2X2_766 ( .A(u2__abc_52155_new_n3521_), .B(u2__abc_52155_new_n3522_), .Y(u2__abc_52155_new_n3523_));
AND2X2 AND2X2_7660 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_5_), .Y(u2__abc_52155_new_n16553_));
AND2X2 AND2X2_7661 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16553_), .Y(u2__abc_52155_new_n16554_));
AND2X2 AND2X2_7662 ( .A(u2__abc_52155_new_n16555_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__7_));
AND2X2 AND2X2_7663 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_8_), .Y(u2__abc_52155_new_n16557_));
AND2X2 AND2X2_7664 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_6_), .Y(u2__abc_52155_new_n16558_));
AND2X2 AND2X2_7665 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16558_), .Y(u2__abc_52155_new_n16559_));
AND2X2 AND2X2_7666 ( .A(u2__abc_52155_new_n16560_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__8_));
AND2X2 AND2X2_7667 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_9_), .Y(u2__abc_52155_new_n16562_));
AND2X2 AND2X2_7668 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_7_), .Y(u2__abc_52155_new_n16563_));
AND2X2 AND2X2_7669 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16563_), .Y(u2__abc_52155_new_n16564_));
AND2X2 AND2X2_767 ( .A(u2__abc_52155_new_n3524_), .B(u2_remHi_31_), .Y(u2__abc_52155_new_n3525_));
AND2X2 AND2X2_7670 ( .A(u2__abc_52155_new_n16565_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__9_));
AND2X2 AND2X2_7671 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_10_), .Y(u2__abc_52155_new_n16567_));
AND2X2 AND2X2_7672 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_8_), .Y(u2__abc_52155_new_n16568_));
AND2X2 AND2X2_7673 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16568_), .Y(u2__abc_52155_new_n16569_));
AND2X2 AND2X2_7674 ( .A(u2__abc_52155_new_n16570_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__10_));
AND2X2 AND2X2_7675 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_11_), .Y(u2__abc_52155_new_n16572_));
AND2X2 AND2X2_7676 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_9_), .Y(u2__abc_52155_new_n16573_));
AND2X2 AND2X2_7677 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16573_), .Y(u2__abc_52155_new_n16574_));
AND2X2 AND2X2_7678 ( .A(u2__abc_52155_new_n16575_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__11_));
AND2X2 AND2X2_7679 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_12_), .Y(u2__abc_52155_new_n16577_));
AND2X2 AND2X2_768 ( .A(u2__abc_52155_new_n3527_), .B(sqrto_31_), .Y(u2__abc_52155_new_n3528_));
AND2X2 AND2X2_7680 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_10_), .Y(u2__abc_52155_new_n16578_));
AND2X2 AND2X2_7681 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16578_), .Y(u2__abc_52155_new_n16579_));
AND2X2 AND2X2_7682 ( .A(u2__abc_52155_new_n16580_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__12_));
AND2X2 AND2X2_7683 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_13_), .Y(u2__abc_52155_new_n16582_));
AND2X2 AND2X2_7684 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_11_), .Y(u2__abc_52155_new_n16583_));
AND2X2 AND2X2_7685 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16583_), .Y(u2__abc_52155_new_n16584_));
AND2X2 AND2X2_7686 ( .A(u2__abc_52155_new_n16585_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__13_));
AND2X2 AND2X2_7687 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_14_), .Y(u2__abc_52155_new_n16587_));
AND2X2 AND2X2_7688 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_12_), .Y(u2__abc_52155_new_n16588_));
AND2X2 AND2X2_7689 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16588_), .Y(u2__abc_52155_new_n16589_));
AND2X2 AND2X2_769 ( .A(u2__abc_52155_new_n3526_), .B(u2__abc_52155_new_n3529_), .Y(u2__abc_52155_new_n3530_));
AND2X2 AND2X2_7690 ( .A(u2__abc_52155_new_n16590_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__14_));
AND2X2 AND2X2_7691 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_15_), .Y(u2__abc_52155_new_n16592_));
AND2X2 AND2X2_7692 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_13_), .Y(u2__abc_52155_new_n16593_));
AND2X2 AND2X2_7693 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16593_), .Y(u2__abc_52155_new_n16594_));
AND2X2 AND2X2_7694 ( .A(u2__abc_52155_new_n16595_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__15_));
AND2X2 AND2X2_7695 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_16_), .Y(u2__abc_52155_new_n16597_));
AND2X2 AND2X2_7696 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_14_), .Y(u2__abc_52155_new_n16598_));
AND2X2 AND2X2_7697 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16598_), .Y(u2__abc_52155_new_n16599_));
AND2X2 AND2X2_7698 ( .A(u2__abc_52155_new_n16600_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__16_));
AND2X2 AND2X2_7699 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_17_), .Y(u2__abc_52155_new_n16602_));
AND2X2 AND2X2_77 ( .A(_abc_73687_new_n831_), .B(_abc_73687_new_n830_), .Y(\o[112] ));
AND2X2 AND2X2_770 ( .A(u2__abc_52155_new_n3530_), .B(u2__abc_52155_new_n3523_), .Y(u2__abc_52155_new_n3531_));
AND2X2 AND2X2_7700 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_15_), .Y(u2__abc_52155_new_n16603_));
AND2X2 AND2X2_7701 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16603_), .Y(u2__abc_52155_new_n16604_));
AND2X2 AND2X2_7702 ( .A(u2__abc_52155_new_n16605_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__17_));
AND2X2 AND2X2_7703 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_18_), .Y(u2__abc_52155_new_n16607_));
AND2X2 AND2X2_7704 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_16_), .Y(u2__abc_52155_new_n16608_));
AND2X2 AND2X2_7705 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16608_), .Y(u2__abc_52155_new_n16609_));
AND2X2 AND2X2_7706 ( .A(u2__abc_52155_new_n16610_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__18_));
AND2X2 AND2X2_7707 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_19_), .Y(u2__abc_52155_new_n16612_));
AND2X2 AND2X2_7708 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_17_), .Y(u2__abc_52155_new_n16613_));
AND2X2 AND2X2_7709 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16613_), .Y(u2__abc_52155_new_n16614_));
AND2X2 AND2X2_771 ( .A(u2__abc_52155_new_n3518_), .B(u2__abc_52155_new_n3531_), .Y(u2__abc_52155_new_n3532_));
AND2X2 AND2X2_7710 ( .A(u2__abc_52155_new_n16615_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__19_));
AND2X2 AND2X2_7711 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_20_), .Y(u2__abc_52155_new_n16617_));
AND2X2 AND2X2_7712 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_18_), .Y(u2__abc_52155_new_n16618_));
AND2X2 AND2X2_7713 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16618_), .Y(u2__abc_52155_new_n16619_));
AND2X2 AND2X2_7714 ( .A(u2__abc_52155_new_n16620_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__20_));
AND2X2 AND2X2_7715 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_21_), .Y(u2__abc_52155_new_n16622_));
AND2X2 AND2X2_7716 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_19_), .Y(u2__abc_52155_new_n16623_));
AND2X2 AND2X2_7717 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16623_), .Y(u2__abc_52155_new_n16624_));
AND2X2 AND2X2_7718 ( .A(u2__abc_52155_new_n16625_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__21_));
AND2X2 AND2X2_7719 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_22_), .Y(u2__abc_52155_new_n16627_));
AND2X2 AND2X2_772 ( .A(u2__abc_52155_new_n3533_), .B(u2_remHi_36_), .Y(u2__abc_52155_new_n3534_));
AND2X2 AND2X2_7720 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_20_), .Y(u2__abc_52155_new_n16628_));
AND2X2 AND2X2_7721 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16628_), .Y(u2__abc_52155_new_n16629_));
AND2X2 AND2X2_7722 ( .A(u2__abc_52155_new_n16630_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__22_));
AND2X2 AND2X2_7723 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_23_), .Y(u2__abc_52155_new_n16632_));
AND2X2 AND2X2_7724 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_21_), .Y(u2__abc_52155_new_n16633_));
AND2X2 AND2X2_7725 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16633_), .Y(u2__abc_52155_new_n16634_));
AND2X2 AND2X2_7726 ( .A(u2__abc_52155_new_n16635_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__23_));
AND2X2 AND2X2_7727 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_24_), .Y(u2__abc_52155_new_n16637_));
AND2X2 AND2X2_7728 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_22_), .Y(u2__abc_52155_new_n16638_));
AND2X2 AND2X2_7729 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16638_), .Y(u2__abc_52155_new_n16639_));
AND2X2 AND2X2_773 ( .A(u2__abc_52155_new_n3535_), .B(sqrto_36_), .Y(u2__abc_52155_new_n3536_));
AND2X2 AND2X2_7730 ( .A(u2__abc_52155_new_n16640_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__24_));
AND2X2 AND2X2_7731 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_25_), .Y(u2__abc_52155_new_n16642_));
AND2X2 AND2X2_7732 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_23_), .Y(u2__abc_52155_new_n16643_));
AND2X2 AND2X2_7733 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16643_), .Y(u2__abc_52155_new_n16644_));
AND2X2 AND2X2_7734 ( .A(u2__abc_52155_new_n16645_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__25_));
AND2X2 AND2X2_7735 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_26_), .Y(u2__abc_52155_new_n16647_));
AND2X2 AND2X2_7736 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_24_), .Y(u2__abc_52155_new_n16648_));
AND2X2 AND2X2_7737 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16648_), .Y(u2__abc_52155_new_n16649_));
AND2X2 AND2X2_7738 ( .A(u2__abc_52155_new_n16650_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__26_));
AND2X2 AND2X2_7739 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_27_), .Y(u2__abc_52155_new_n16652_));
AND2X2 AND2X2_774 ( .A(u2__abc_52155_new_n3538_), .B(u2_remHi_37_), .Y(u2__abc_52155_new_n3539_));
AND2X2 AND2X2_7740 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_25_), .Y(u2__abc_52155_new_n16653_));
AND2X2 AND2X2_7741 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16653_), .Y(u2__abc_52155_new_n16654_));
AND2X2 AND2X2_7742 ( .A(u2__abc_52155_new_n16655_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__27_));
AND2X2 AND2X2_7743 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_28_), .Y(u2__abc_52155_new_n16657_));
AND2X2 AND2X2_7744 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_26_), .Y(u2__abc_52155_new_n16658_));
AND2X2 AND2X2_7745 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16658_), .Y(u2__abc_52155_new_n16659_));
AND2X2 AND2X2_7746 ( .A(u2__abc_52155_new_n16660_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__28_));
AND2X2 AND2X2_7747 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_29_), .Y(u2__abc_52155_new_n16662_));
AND2X2 AND2X2_7748 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_27_), .Y(u2__abc_52155_new_n16663_));
AND2X2 AND2X2_7749 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16663_), .Y(u2__abc_52155_new_n16664_));
AND2X2 AND2X2_775 ( .A(u2__abc_52155_new_n3540_), .B(sqrto_37_), .Y(u2__abc_52155_new_n3541_));
AND2X2 AND2X2_7750 ( .A(u2__abc_52155_new_n16665_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__29_));
AND2X2 AND2X2_7751 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_30_), .Y(u2__abc_52155_new_n16667_));
AND2X2 AND2X2_7752 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_28_), .Y(u2__abc_52155_new_n16668_));
AND2X2 AND2X2_7753 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16668_), .Y(u2__abc_52155_new_n16669_));
AND2X2 AND2X2_7754 ( .A(u2__abc_52155_new_n16670_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__30_));
AND2X2 AND2X2_7755 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_31_), .Y(u2__abc_52155_new_n16672_));
AND2X2 AND2X2_7756 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_29_), .Y(u2__abc_52155_new_n16673_));
AND2X2 AND2X2_7757 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n16673_), .Y(u2__abc_52155_new_n16674_));
AND2X2 AND2X2_7758 ( .A(u2__abc_52155_new_n16675_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__31_));
AND2X2 AND2X2_7759 ( .A(u2__abc_52155_new_n3001_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n16677_));
AND2X2 AND2X2_776 ( .A(u2__abc_52155_new_n3544_), .B(u2_remHi_35_), .Y(u2__abc_52155_new_n3545_));
AND2X2 AND2X2_7760 ( .A(u2__abc_52155_new_n16678_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16679_));
AND2X2 AND2X2_7761 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_32_), .Y(u2__abc_52155_new_n16681_));
AND2X2 AND2X2_7762 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16682_));
AND2X2 AND2X2_7763 ( .A(u2__abc_52155_new_n16470_), .B(u2_state_2_), .Y(u2__abc_52155_new_n16683_));
AND2X2 AND2X2_7764 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_30_), .Y(u2__abc_52155_new_n16684_));
AND2X2 AND2X2_7765 ( .A(u2__abc_52155_new_n16685_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16686_));
AND2X2 AND2X2_7766 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_33_), .Y(u2__abc_52155_new_n16688_));
AND2X2 AND2X2_7767 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_31_), .Y(u2__abc_52155_new_n16689_));
AND2X2 AND2X2_7768 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16690_));
AND2X2 AND2X2_7769 ( .A(u2__abc_52155_new_n16691_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16692_));
AND2X2 AND2X2_777 ( .A(u2__abc_52155_new_n3546_), .B(sqrto_35_), .Y(u2__abc_52155_new_n3547_));
AND2X2 AND2X2_7770 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_34_), .Y(u2__abc_52155_new_n16694_));
AND2X2 AND2X2_7771 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_32_), .Y(u2__abc_52155_new_n16695_));
AND2X2 AND2X2_7772 ( .A(u2__abc_52155_new_n16696_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16697_));
AND2X2 AND2X2_7773 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_34_), .Y(u2__abc_52155_new_n16698_));
AND2X2 AND2X2_7774 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n16699_));
AND2X2 AND2X2_7775 ( .A(u2__abc_52155_new_n16700_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n16701_));
AND2X2 AND2X2_7776 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_35_), .Y(u2__abc_52155_new_n16703_));
AND2X2 AND2X2_7777 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_33_), .Y(u2__abc_52155_new_n16704_));
AND2X2 AND2X2_7778 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16705_));
AND2X2 AND2X2_7779 ( .A(u2__abc_52155_new_n16706_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16707_));
AND2X2 AND2X2_778 ( .A(u2__abc_52155_new_n3549_), .B(u2_remHi_34_), .Y(u2__abc_52155_new_n3550_));
AND2X2 AND2X2_7780 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_36_), .Y(u2__abc_52155_new_n16709_));
AND2X2 AND2X2_7781 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_34_), .Y(u2__abc_52155_new_n16710_));
AND2X2 AND2X2_7782 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16711_));
AND2X2 AND2X2_7783 ( .A(u2__abc_52155_new_n16712_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16713_));
AND2X2 AND2X2_7784 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_37_), .Y(u2__abc_52155_new_n16715_));
AND2X2 AND2X2_7785 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_35_), .Y(u2__abc_52155_new_n16716_));
AND2X2 AND2X2_7786 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16717_));
AND2X2 AND2X2_7787 ( .A(u2__abc_52155_new_n16718_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16719_));
AND2X2 AND2X2_7788 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_38_), .Y(u2__abc_52155_new_n16721_));
AND2X2 AND2X2_7789 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16722_));
AND2X2 AND2X2_779 ( .A(u2__abc_52155_new_n3551_), .B(sqrto_34_), .Y(u2__abc_52155_new_n3552_));
AND2X2 AND2X2_7790 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_36_), .Y(u2__abc_52155_new_n16723_));
AND2X2 AND2X2_7791 ( .A(u2__abc_52155_new_n16724_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16725_));
AND2X2 AND2X2_7792 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_39_), .Y(u2__abc_52155_new_n16727_));
AND2X2 AND2X2_7793 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_37_), .Y(u2__abc_52155_new_n16728_));
AND2X2 AND2X2_7794 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16729_));
AND2X2 AND2X2_7795 ( .A(u2__abc_52155_new_n16730_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16731_));
AND2X2 AND2X2_7796 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_40_), .Y(u2__abc_52155_new_n16733_));
AND2X2 AND2X2_7797 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_38_), .Y(u2__abc_52155_new_n16734_));
AND2X2 AND2X2_7798 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16735_));
AND2X2 AND2X2_7799 ( .A(u2__abc_52155_new_n16736_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16737_));
AND2X2 AND2X2_78 ( .A(_abc_73687_new_n834_), .B(_abc_73687_new_n833_), .Y(\o[113] ));
AND2X2 AND2X2_780 ( .A(u2__abc_52155_new_n3556_), .B(u2__abc_52155_new_n3532_), .Y(u2__abc_52155_new_n3557_));
AND2X2 AND2X2_7800 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_41_), .Y(u2__abc_52155_new_n16739_));
AND2X2 AND2X2_7801 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_39_), .Y(u2__abc_52155_new_n16740_));
AND2X2 AND2X2_7802 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16741_));
AND2X2 AND2X2_7803 ( .A(u2__abc_52155_new_n16742_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16743_));
AND2X2 AND2X2_7804 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_42_), .Y(u2__abc_52155_new_n16745_));
AND2X2 AND2X2_7805 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16746_));
AND2X2 AND2X2_7806 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_40_), .Y(u2__abc_52155_new_n16747_));
AND2X2 AND2X2_7807 ( .A(u2__abc_52155_new_n16748_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16749_));
AND2X2 AND2X2_7808 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_43_), .Y(u2__abc_52155_new_n16751_));
AND2X2 AND2X2_7809 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_41_), .Y(u2__abc_52155_new_n16752_));
AND2X2 AND2X2_781 ( .A(u2__abc_52155_new_n3557_), .B(u2__abc_52155_new_n3506_), .Y(u2__abc_52155_new_n3558_));
AND2X2 AND2X2_7810 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16753_));
AND2X2 AND2X2_7811 ( .A(u2__abc_52155_new_n16754_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16755_));
AND2X2 AND2X2_7812 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_44_), .Y(u2__abc_52155_new_n16757_));
AND2X2 AND2X2_7813 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_42_), .Y(u2__abc_52155_new_n16758_));
AND2X2 AND2X2_7814 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16759_));
AND2X2 AND2X2_7815 ( .A(u2__abc_52155_new_n16760_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16761_));
AND2X2 AND2X2_7816 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_45_), .Y(u2__abc_52155_new_n16763_));
AND2X2 AND2X2_7817 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_43_), .Y(u2__abc_52155_new_n16764_));
AND2X2 AND2X2_7818 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16765_));
AND2X2 AND2X2_7819 ( .A(u2__abc_52155_new_n16766_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16767_));
AND2X2 AND2X2_782 ( .A(u2__abc_52155_new_n3558_), .B(u2__abc_52155_new_n3446_), .Y(u2__abc_52155_new_n3559_));
AND2X2 AND2X2_7820 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_46_), .Y(u2__abc_52155_new_n16769_));
AND2X2 AND2X2_7821 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_44_), .Y(u2__abc_52155_new_n16770_));
AND2X2 AND2X2_7822 ( .A(u2__abc_52155_new_n16771_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16772_));
AND2X2 AND2X2_7823 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_46_), .Y(u2__abc_52155_new_n16773_));
AND2X2 AND2X2_7824 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n16774_));
AND2X2 AND2X2_7825 ( .A(u2__abc_52155_new_n16775_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n16776_));
AND2X2 AND2X2_7826 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_47_), .Y(u2__abc_52155_new_n16778_));
AND2X2 AND2X2_7827 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16779_));
AND2X2 AND2X2_7828 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_45_), .Y(u2__abc_52155_new_n16780_));
AND2X2 AND2X2_7829 ( .A(u2__abc_52155_new_n16781_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16782_));
AND2X2 AND2X2_783 ( .A(u2__abc_52155_new_n3564_), .B(u2__abc_52155_new_n3529_), .Y(u2__abc_52155_new_n3565_));
AND2X2 AND2X2_7830 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_48_), .Y(u2__abc_52155_new_n16784_));
AND2X2 AND2X2_7831 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_46_), .Y(u2__abc_52155_new_n16785_));
AND2X2 AND2X2_7832 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16786_));
AND2X2 AND2X2_7833 ( .A(u2__abc_52155_new_n16787_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16788_));
AND2X2 AND2X2_7834 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_49_), .Y(u2__abc_52155_new_n16790_));
AND2X2 AND2X2_7835 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_47_), .Y(u2__abc_52155_new_n16791_));
AND2X2 AND2X2_7836 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16792_));
AND2X2 AND2X2_7837 ( .A(u2__abc_52155_new_n16793_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16794_));
AND2X2 AND2X2_7838 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_50_), .Y(u2__abc_52155_new_n16796_));
AND2X2 AND2X2_7839 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_48_), .Y(u2__abc_52155_new_n16797_));
AND2X2 AND2X2_784 ( .A(u2__abc_52155_new_n3569_), .B(u2__abc_52155_new_n3567_), .Y(u2__abc_52155_new_n3570_));
AND2X2 AND2X2_7840 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16798_));
AND2X2 AND2X2_7841 ( .A(u2__abc_52155_new_n16799_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16800_));
AND2X2 AND2X2_7842 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_51_), .Y(u2__abc_52155_new_n16802_));
AND2X2 AND2X2_7843 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16803_));
AND2X2 AND2X2_7844 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_49_), .Y(u2__abc_52155_new_n16804_));
AND2X2 AND2X2_7845 ( .A(u2__abc_52155_new_n16805_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16806_));
AND2X2 AND2X2_7846 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_52_), .Y(u2__abc_52155_new_n16808_));
AND2X2 AND2X2_7847 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_50_), .Y(u2__abc_52155_new_n16809_));
AND2X2 AND2X2_7848 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16810_));
AND2X2 AND2X2_7849 ( .A(u2__abc_52155_new_n16811_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16812_));
AND2X2 AND2X2_785 ( .A(u2__abc_52155_new_n3566_), .B(u2__abc_52155_new_n3570_), .Y(u2__abc_52155_new_n3571_));
AND2X2 AND2X2_7850 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_53_), .Y(u2__abc_52155_new_n16814_));
AND2X2 AND2X2_7851 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_51_), .Y(u2__abc_52155_new_n16815_));
AND2X2 AND2X2_7852 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16816_));
AND2X2 AND2X2_7853 ( .A(u2__abc_52155_new_n16817_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16818_));
AND2X2 AND2X2_7854 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_54_), .Y(u2__abc_52155_new_n16820_));
AND2X2 AND2X2_7855 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_52_), .Y(u2__abc_52155_new_n16821_));
AND2X2 AND2X2_7856 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16822_));
AND2X2 AND2X2_7857 ( .A(u2__abc_52155_new_n16823_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16824_));
AND2X2 AND2X2_7858 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_55_), .Y(u2__abc_52155_new_n16826_));
AND2X2 AND2X2_7859 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_53_), .Y(u2__abc_52155_new_n16827_));
AND2X2 AND2X2_786 ( .A(u2__abc_52155_new_n3575_), .B(u2__abc_52155_new_n3573_), .Y(u2__abc_52155_new_n3576_));
AND2X2 AND2X2_7860 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16828_));
AND2X2 AND2X2_7861 ( .A(u2__abc_52155_new_n16829_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16830_));
AND2X2 AND2X2_7862 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_56_), .Y(u2__abc_52155_new_n16832_));
AND2X2 AND2X2_7863 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_54_), .Y(u2__abc_52155_new_n16833_));
AND2X2 AND2X2_7864 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16834_));
AND2X2 AND2X2_7865 ( .A(u2__abc_52155_new_n16835_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16836_));
AND2X2 AND2X2_7866 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_57_), .Y(u2__abc_52155_new_n16838_));
AND2X2 AND2X2_7867 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16839_));
AND2X2 AND2X2_7868 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_55_), .Y(u2__abc_52155_new_n16840_));
AND2X2 AND2X2_7869 ( .A(u2__abc_52155_new_n16841_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16842_));
AND2X2 AND2X2_787 ( .A(u2__abc_52155_new_n3578_), .B(u2__abc_52155_new_n3536_), .Y(u2__abc_52155_new_n3579_));
AND2X2 AND2X2_7870 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_58_), .Y(u2__abc_52155_new_n16844_));
AND2X2 AND2X2_7871 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16845_));
AND2X2 AND2X2_7872 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_56_), .Y(u2__abc_52155_new_n16846_));
AND2X2 AND2X2_7873 ( .A(u2__abc_52155_new_n16847_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16848_));
AND2X2 AND2X2_7874 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_59_), .Y(u2__abc_52155_new_n16850_));
AND2X2 AND2X2_7875 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_57_), .Y(u2__abc_52155_new_n16851_));
AND2X2 AND2X2_7876 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16852_));
AND2X2 AND2X2_7877 ( .A(u2__abc_52155_new_n16853_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16854_));
AND2X2 AND2X2_7878 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_60_), .Y(u2__abc_52155_new_n16856_));
AND2X2 AND2X2_7879 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_58_), .Y(u2__abc_52155_new_n16857_));
AND2X2 AND2X2_788 ( .A(u2__abc_52155_new_n3577_), .B(u2__abc_52155_new_n3581_), .Y(u2__abc_52155_new_n3582_));
AND2X2 AND2X2_7880 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16858_));
AND2X2 AND2X2_7881 ( .A(u2__abc_52155_new_n16859_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16860_));
AND2X2 AND2X2_7882 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_61_), .Y(u2__abc_52155_new_n16862_));
AND2X2 AND2X2_7883 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_59_), .Y(u2__abc_52155_new_n16863_));
AND2X2 AND2X2_7884 ( .A(u2__abc_52155_new_n16864_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16865_));
AND2X2 AND2X2_7885 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_61_), .Y(u2__abc_52155_new_n16866_));
AND2X2 AND2X2_7886 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n16867_));
AND2X2 AND2X2_7887 ( .A(u2__abc_52155_new_n16868_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n16869_));
AND2X2 AND2X2_7888 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_62_), .Y(u2__abc_52155_new_n16871_));
AND2X2 AND2X2_7889 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_60_), .Y(u2__abc_52155_new_n16872_));
AND2X2 AND2X2_789 ( .A(u2__abc_52155_new_n3572_), .B(u2__abc_52155_new_n3582_), .Y(u2__abc_52155_new_n3583_));
AND2X2 AND2X2_7890 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16873_));
AND2X2 AND2X2_7891 ( .A(u2__abc_52155_new_n16874_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16875_));
AND2X2 AND2X2_7892 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_63_), .Y(u2__abc_52155_new_n16877_));
AND2X2 AND2X2_7893 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16878_));
AND2X2 AND2X2_7894 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_61_), .Y(u2__abc_52155_new_n16879_));
AND2X2 AND2X2_7895 ( .A(u2__abc_52155_new_n16880_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16881_));
AND2X2 AND2X2_7896 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_64_), .Y(u2__abc_52155_new_n16883_));
AND2X2 AND2X2_7897 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16884_));
AND2X2 AND2X2_7898 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_62_), .Y(u2__abc_52155_new_n16885_));
AND2X2 AND2X2_7899 ( .A(u2__abc_52155_new_n16886_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16887_));
AND2X2 AND2X2_79 ( .A(_abc_73687_new_n837_), .B(_abc_73687_new_n836_), .Y(\o[114] ));
AND2X2 AND2X2_790 ( .A(u2__abc_52155_new_n3586_), .B(u2__abc_52155_new_n3471_), .Y(u2__abc_52155_new_n3587_));
AND2X2 AND2X2_7900 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_65_), .Y(u2__abc_52155_new_n16889_));
AND2X2 AND2X2_7901 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_63_), .Y(u2__abc_52155_new_n16890_));
AND2X2 AND2X2_7902 ( .A(u2__abc_52155_new_n16891_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16892_));
AND2X2 AND2X2_7903 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_65_), .Y(u2__abc_52155_new_n16893_));
AND2X2 AND2X2_7904 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n16894_));
AND2X2 AND2X2_7905 ( .A(u2__abc_52155_new_n16895_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n16896_));
AND2X2 AND2X2_7906 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_66_), .Y(u2__abc_52155_new_n16898_));
AND2X2 AND2X2_7907 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16899_));
AND2X2 AND2X2_7908 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_64_), .Y(u2__abc_52155_new_n16900_));
AND2X2 AND2X2_7909 ( .A(u2__abc_52155_new_n16901_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16902_));
AND2X2 AND2X2_791 ( .A(u2__abc_52155_new_n3589_), .B(u2__abc_52155_new_n3450_), .Y(u2__abc_52155_new_n3590_));
AND2X2 AND2X2_7910 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_67_), .Y(u2__abc_52155_new_n16904_));
AND2X2 AND2X2_7911 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_65_), .Y(u2__abc_52155_new_n16905_));
AND2X2 AND2X2_7912 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16906_));
AND2X2 AND2X2_7913 ( .A(u2__abc_52155_new_n16907_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16908_));
AND2X2 AND2X2_7914 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_68_), .Y(u2__abc_52155_new_n16910_));
AND2X2 AND2X2_7915 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_66_), .Y(u2__abc_52155_new_n16911_));
AND2X2 AND2X2_7916 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16912_));
AND2X2 AND2X2_7917 ( .A(u2__abc_52155_new_n16913_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16914_));
AND2X2 AND2X2_7918 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_69_), .Y(u2__abc_52155_new_n16916_));
AND2X2 AND2X2_7919 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_67_), .Y(u2__abc_52155_new_n16917_));
AND2X2 AND2X2_792 ( .A(u2__abc_52155_new_n3588_), .B(u2__abc_52155_new_n3592_), .Y(u2__abc_52155_new_n3593_));
AND2X2 AND2X2_7920 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16918_));
AND2X2 AND2X2_7921 ( .A(u2__abc_52155_new_n16919_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16920_));
AND2X2 AND2X2_7922 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_70_), .Y(u2__abc_52155_new_n16922_));
AND2X2 AND2X2_7923 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16923_));
AND2X2 AND2X2_7924 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_68_), .Y(u2__abc_52155_new_n16924_));
AND2X2 AND2X2_7925 ( .A(u2__abc_52155_new_n16925_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16926_));
AND2X2 AND2X2_7926 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_71_), .Y(u2__abc_52155_new_n16928_));
AND2X2 AND2X2_7927 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_69_), .Y(u2__abc_52155_new_n16929_));
AND2X2 AND2X2_7928 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16930_));
AND2X2 AND2X2_7929 ( .A(u2__abc_52155_new_n16931_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16932_));
AND2X2 AND2X2_793 ( .A(u2__abc_52155_new_n3492_), .B(u2__abc_52155_new_n3501_), .Y(u2__abc_52155_new_n3595_));
AND2X2 AND2X2_7930 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_72_), .Y(u2__abc_52155_new_n16934_));
AND2X2 AND2X2_7931 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_70_), .Y(u2__abc_52155_new_n16935_));
AND2X2 AND2X2_7932 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16936_));
AND2X2 AND2X2_7933 ( .A(u2__abc_52155_new_n16937_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16938_));
AND2X2 AND2X2_7934 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_73_), .Y(u2__abc_52155_new_n16940_));
AND2X2 AND2X2_7935 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_71_), .Y(u2__abc_52155_new_n16941_));
AND2X2 AND2X2_7936 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16942_));
AND2X2 AND2X2_7937 ( .A(u2__abc_52155_new_n16943_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16944_));
AND2X2 AND2X2_7938 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_74_), .Y(u2__abc_52155_new_n16946_));
AND2X2 AND2X2_7939 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_72_), .Y(u2__abc_52155_new_n16947_));
AND2X2 AND2X2_794 ( .A(u2__abc_52155_new_n3596_), .B(u2__abc_52155_new_n3489_), .Y(u2__abc_52155_new_n3597_));
AND2X2 AND2X2_7940 ( .A(u2__abc_52155_new_n16948_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16949_));
AND2X2 AND2X2_7941 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_74_), .Y(u2__abc_52155_new_n16950_));
AND2X2 AND2X2_7942 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n16951_));
AND2X2 AND2X2_7943 ( .A(u2__abc_52155_new_n16952_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n16953_));
AND2X2 AND2X2_7944 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_75_), .Y(u2__abc_52155_new_n16955_));
AND2X2 AND2X2_7945 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_73_), .Y(u2__abc_52155_new_n16956_));
AND2X2 AND2X2_7946 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16957_));
AND2X2 AND2X2_7947 ( .A(u2__abc_52155_new_n16958_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16959_));
AND2X2 AND2X2_7948 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_76_), .Y(u2__abc_52155_new_n16961_));
AND2X2 AND2X2_7949 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_74_), .Y(u2__abc_52155_new_n16962_));
AND2X2 AND2X2_795 ( .A(u2__abc_52155_new_n3484_), .B(u2__abc_52155_new_n3479_), .Y(u2__abc_52155_new_n3598_));
AND2X2 AND2X2_7950 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16963_));
AND2X2 AND2X2_7951 ( .A(u2__abc_52155_new_n16964_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16965_));
AND2X2 AND2X2_7952 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_77_), .Y(u2__abc_52155_new_n16967_));
AND2X2 AND2X2_7953 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_75_), .Y(u2__abc_52155_new_n16968_));
AND2X2 AND2X2_7954 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16969_));
AND2X2 AND2X2_7955 ( .A(u2__abc_52155_new_n16970_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16971_));
AND2X2 AND2X2_7956 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_78_), .Y(u2__abc_52155_new_n16973_));
AND2X2 AND2X2_7957 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_76_), .Y(u2__abc_52155_new_n16974_));
AND2X2 AND2X2_7958 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16975_));
AND2X2 AND2X2_7959 ( .A(u2__abc_52155_new_n16976_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16977_));
AND2X2 AND2X2_796 ( .A(u2__abc_52155_new_n3594_), .B(u2__abc_52155_new_n3601_), .Y(u2__abc_52155_new_n3602_));
AND2X2 AND2X2_7960 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_79_), .Y(u2__abc_52155_new_n16979_));
AND2X2 AND2X2_7961 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16980_));
AND2X2 AND2X2_7962 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_77_), .Y(u2__abc_52155_new_n16981_));
AND2X2 AND2X2_7963 ( .A(u2__abc_52155_new_n16982_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16983_));
AND2X2 AND2X2_7964 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_80_), .Y(u2__abc_52155_new_n16985_));
AND2X2 AND2X2_7965 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_78_), .Y(u2__abc_52155_new_n16986_));
AND2X2 AND2X2_7966 ( .A(u2__abc_52155_new_n16987_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16988_));
AND2X2 AND2X2_7967 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_80_), .Y(u2__abc_52155_new_n16989_));
AND2X2 AND2X2_7968 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n16990_));
AND2X2 AND2X2_7969 ( .A(u2__abc_52155_new_n16991_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n16992_));
AND2X2 AND2X2_797 ( .A(u2__abc_52155_new_n3584_), .B(u2__abc_52155_new_n3602_), .Y(u2__abc_52155_new_n3603_));
AND2X2 AND2X2_7970 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_81_), .Y(u2__abc_52155_new_n16994_));
AND2X2 AND2X2_7971 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_79_), .Y(u2__abc_52155_new_n16995_));
AND2X2 AND2X2_7972 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n16996_));
AND2X2 AND2X2_7973 ( .A(u2__abc_52155_new_n16997_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n16998_));
AND2X2 AND2X2_7974 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_82_), .Y(u2__abc_52155_new_n17000_));
AND2X2 AND2X2_7975 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_80_), .Y(u2__abc_52155_new_n17001_));
AND2X2 AND2X2_7976 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17002_));
AND2X2 AND2X2_7977 ( .A(u2__abc_52155_new_n17003_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17004_));
AND2X2 AND2X2_7978 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_83_), .Y(u2__abc_52155_new_n17006_));
AND2X2 AND2X2_7979 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17007_));
AND2X2 AND2X2_798 ( .A(u2__abc_52155_new_n3607_), .B(u2__abc_52155_new_n3403_), .Y(u2__abc_52155_new_n3608_));
AND2X2 AND2X2_7980 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_81_), .Y(u2__abc_52155_new_n17008_));
AND2X2 AND2X2_7981 ( .A(u2__abc_52155_new_n17009_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17010_));
AND2X2 AND2X2_7982 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_84_), .Y(u2__abc_52155_new_n17012_));
AND2X2 AND2X2_7983 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_82_), .Y(u2__abc_52155_new_n17013_));
AND2X2 AND2X2_7984 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17014_));
AND2X2 AND2X2_7985 ( .A(u2__abc_52155_new_n17015_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17016_));
AND2X2 AND2X2_7986 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_85_), .Y(u2__abc_52155_new_n17018_));
AND2X2 AND2X2_7987 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_83_), .Y(u2__abc_52155_new_n17019_));
AND2X2 AND2X2_7988 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17020_));
AND2X2 AND2X2_7989 ( .A(u2__abc_52155_new_n17021_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17022_));
AND2X2 AND2X2_799 ( .A(u2__abc_52155_new_n3610_), .B(u2__abc_52155_new_n3389_), .Y(u2__abc_52155_new_n3611_));
AND2X2 AND2X2_7990 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_86_), .Y(u2__abc_52155_new_n17024_));
AND2X2 AND2X2_7991 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_84_), .Y(u2__abc_52155_new_n17025_));
AND2X2 AND2X2_7992 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17026_));
AND2X2 AND2X2_7993 ( .A(u2__abc_52155_new_n17027_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17028_));
AND2X2 AND2X2_7994 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_87_), .Y(u2__abc_52155_new_n17030_));
AND2X2 AND2X2_7995 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_85_), .Y(u2__abc_52155_new_n17031_));
AND2X2 AND2X2_7996 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17032_));
AND2X2 AND2X2_7997 ( .A(u2__abc_52155_new_n17033_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17034_));
AND2X2 AND2X2_7998 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_88_), .Y(u2__abc_52155_new_n17036_));
AND2X2 AND2X2_7999 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_86_), .Y(u2__abc_52155_new_n17037_));
AND2X2 AND2X2_8 ( .A(_abc_73687_new_n753_), .B(sqrto_7_), .Y(\o[43] ));
AND2X2 AND2X2_80 ( .A(_abc_73687_new_n840_), .B(_abc_73687_new_n839_), .Y(\o[115] ));
AND2X2 AND2X2_800 ( .A(u2__abc_52155_new_n3609_), .B(u2__abc_52155_new_n3613_), .Y(u2__abc_52155_new_n3614_));
AND2X2 AND2X2_8000 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17038_));
AND2X2 AND2X2_8001 ( .A(u2__abc_52155_new_n17039_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17040_));
AND2X2 AND2X2_8002 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_89_), .Y(u2__abc_52155_new_n17042_));
AND2X2 AND2X2_8003 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17043_));
AND2X2 AND2X2_8004 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_87_), .Y(u2__abc_52155_new_n17044_));
AND2X2 AND2X2_8005 ( .A(u2__abc_52155_new_n17045_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17046_));
AND2X2 AND2X2_8006 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_90_), .Y(u2__abc_52155_new_n17048_));
AND2X2 AND2X2_8007 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_88_), .Y(u2__abc_52155_new_n17049_));
AND2X2 AND2X2_8008 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17050_));
AND2X2 AND2X2_8009 ( .A(u2__abc_52155_new_n17051_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17052_));
AND2X2 AND2X2_801 ( .A(u2__abc_52155_new_n3431_), .B(u2__abc_52155_new_n3440_), .Y(u2__abc_52155_new_n3616_));
AND2X2 AND2X2_8010 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_91_), .Y(u2__abc_52155_new_n17054_));
AND2X2 AND2X2_8011 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_89_), .Y(u2__abc_52155_new_n17055_));
AND2X2 AND2X2_8012 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17056_));
AND2X2 AND2X2_8013 ( .A(u2__abc_52155_new_n17057_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17058_));
AND2X2 AND2X2_8014 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_92_), .Y(u2__abc_52155_new_n17060_));
AND2X2 AND2X2_8015 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_90_), .Y(u2__abc_52155_new_n17061_));
AND2X2 AND2X2_8016 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17062_));
AND2X2 AND2X2_8017 ( .A(u2__abc_52155_new_n17063_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17064_));
AND2X2 AND2X2_8018 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_93_), .Y(u2__abc_52155_new_n17066_));
AND2X2 AND2X2_8019 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17067_));
AND2X2 AND2X2_802 ( .A(u2__abc_52155_new_n3617_), .B(u2__abc_52155_new_n3428_), .Y(u2__abc_52155_new_n3618_));
AND2X2 AND2X2_8020 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_91_), .Y(u2__abc_52155_new_n17068_));
AND2X2 AND2X2_8021 ( .A(u2__abc_52155_new_n17069_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17070_));
AND2X2 AND2X2_8022 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_94_), .Y(u2__abc_52155_new_n17072_));
AND2X2 AND2X2_8023 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_92_), .Y(u2__abc_52155_new_n17073_));
AND2X2 AND2X2_8024 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17074_));
AND2X2 AND2X2_8025 ( .A(u2__abc_52155_new_n17075_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17076_));
AND2X2 AND2X2_8026 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_95_), .Y(u2__abc_52155_new_n17078_));
AND2X2 AND2X2_8027 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17079_));
AND2X2 AND2X2_8028 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_93_), .Y(u2__abc_52155_new_n17080_));
AND2X2 AND2X2_8029 ( .A(u2__abc_52155_new_n17081_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17082_));
AND2X2 AND2X2_803 ( .A(u2__abc_52155_new_n3423_), .B(u2__abc_52155_new_n3418_), .Y(u2__abc_52155_new_n3619_));
AND2X2 AND2X2_8030 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_96_), .Y(u2__abc_52155_new_n17084_));
AND2X2 AND2X2_8031 ( .A(u2__abc_52155_new_n2964_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17085_));
AND2X2 AND2X2_8032 ( .A(u2__abc_52155_new_n17085_), .B(1'h0), .Y(u2__abc_52155_new_n17086_));
AND2X2 AND2X2_8033 ( .A(u2__abc_52155_new_n2982_), .B(u2_remLo_94_), .Y(u2__abc_52155_new_n17087_));
AND2X2 AND2X2_8034 ( .A(u2__abc_52155_new_n16683_), .B(u2__abc_52155_new_n17087_), .Y(u2__abc_52155_new_n17088_));
AND2X2 AND2X2_8035 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_97_), .Y(u2__abc_52155_new_n17091_));
AND2X2 AND2X2_8036 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_95_), .Y(u2__abc_52155_new_n17092_));
AND2X2 AND2X2_8037 ( .A(u2__abc_52155_new_n17093_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17094_));
AND2X2 AND2X2_8038 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_97_), .Y(u2__abc_52155_new_n17095_));
AND2X2 AND2X2_8039 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n17096_));
AND2X2 AND2X2_804 ( .A(u2__abc_52155_new_n3615_), .B(u2__abc_52155_new_n3622_), .Y(u2__abc_52155_new_n3623_));
AND2X2 AND2X2_8040 ( .A(u2__abc_52155_new_n17097_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17098_));
AND2X2 AND2X2_8041 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_98_), .Y(u2__abc_52155_new_n17100_));
AND2X2 AND2X2_8042 ( .A(u2__abc_52155_new_n17085_), .B(1'h0), .Y(u2__abc_52155_new_n17101_));
AND2X2 AND2X2_8043 ( .A(u2__abc_52155_new_n2982_), .B(u2_remLo_96_), .Y(u2__abc_52155_new_n17102_));
AND2X2 AND2X2_8044 ( .A(u2__abc_52155_new_n16683_), .B(u2__abc_52155_new_n17102_), .Y(u2__abc_52155_new_n17103_));
AND2X2 AND2X2_8045 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_99_), .Y(u2__abc_52155_new_n17106_));
AND2X2 AND2X2_8046 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_97_), .Y(u2__abc_52155_new_n17107_));
AND2X2 AND2X2_8047 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17108_));
AND2X2 AND2X2_8048 ( .A(u2__abc_52155_new_n17109_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17110_));
AND2X2 AND2X2_8049 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_100_), .Y(u2__abc_52155_new_n17112_));
AND2X2 AND2X2_805 ( .A(u2__abc_52155_new_n3347_), .B(u2__abc_52155_new_n3342_), .Y(u2__abc_52155_new_n3625_));
AND2X2 AND2X2_8050 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_98_), .Y(u2__abc_52155_new_n17113_));
AND2X2 AND2X2_8051 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17114_));
AND2X2 AND2X2_8052 ( .A(u2__abc_52155_new_n17115_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17116_));
AND2X2 AND2X2_8053 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_101_), .Y(u2__abc_52155_new_n17118_));
AND2X2 AND2X2_8054 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_99_), .Y(u2__abc_52155_new_n17119_));
AND2X2 AND2X2_8055 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17120_));
AND2X2 AND2X2_8056 ( .A(u2__abc_52155_new_n17121_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17122_));
AND2X2 AND2X2_8057 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_102_), .Y(u2__abc_52155_new_n17124_));
AND2X2 AND2X2_8058 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17125_));
AND2X2 AND2X2_8059 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_100_), .Y(u2__abc_52155_new_n17126_));
AND2X2 AND2X2_806 ( .A(u2__abc_52155_new_n3626_), .B(u2__abc_52155_new_n3337_), .Y(u2__abc_52155_new_n3627_));
AND2X2 AND2X2_8060 ( .A(u2__abc_52155_new_n17127_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17128_));
AND2X2 AND2X2_8061 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_103_), .Y(u2__abc_52155_new_n17130_));
AND2X2 AND2X2_8062 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_101_), .Y(u2__abc_52155_new_n17131_));
AND2X2 AND2X2_8063 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17132_));
AND2X2 AND2X2_8064 ( .A(u2__abc_52155_new_n17133_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17134_));
AND2X2 AND2X2_8065 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_104_), .Y(u2__abc_52155_new_n17136_));
AND2X2 AND2X2_8066 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_102_), .Y(u2__abc_52155_new_n17137_));
AND2X2 AND2X2_8067 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17138_));
AND2X2 AND2X2_8068 ( .A(u2__abc_52155_new_n17139_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17140_));
AND2X2 AND2X2_8069 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_105_), .Y(u2__abc_52155_new_n17142_));
AND2X2 AND2X2_807 ( .A(u2__abc_52155_new_n3332_), .B(u2__abc_52155_new_n3327_), .Y(u2__abc_52155_new_n3628_));
AND2X2 AND2X2_8070 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_103_), .Y(u2__abc_52155_new_n17143_));
AND2X2 AND2X2_8071 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17144_));
AND2X2 AND2X2_8072 ( .A(u2__abc_52155_new_n17145_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17146_));
AND2X2 AND2X2_8073 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_106_), .Y(u2__abc_52155_new_n17148_));
AND2X2 AND2X2_8074 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17149_));
AND2X2 AND2X2_8075 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_104_), .Y(u2__abc_52155_new_n17150_));
AND2X2 AND2X2_8076 ( .A(u2__abc_52155_new_n17151_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17152_));
AND2X2 AND2X2_8077 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_107_), .Y(u2__abc_52155_new_n17154_));
AND2X2 AND2X2_8078 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_105_), .Y(u2__abc_52155_new_n17155_));
AND2X2 AND2X2_8079 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17156_));
AND2X2 AND2X2_808 ( .A(u2__abc_52155_new_n3630_), .B(u2__abc_52155_new_n3384_), .Y(u2__abc_52155_new_n3631_));
AND2X2 AND2X2_8080 ( .A(u2__abc_52155_new_n17157_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17158_));
AND2X2 AND2X2_8081 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_108_), .Y(u2__abc_52155_new_n17160_));
AND2X2 AND2X2_8082 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_106_), .Y(u2__abc_52155_new_n17161_));
AND2X2 AND2X2_8083 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17162_));
AND2X2 AND2X2_8084 ( .A(u2__abc_52155_new_n17163_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17164_));
AND2X2 AND2X2_8085 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_109_), .Y(u2__abc_52155_new_n17166_));
AND2X2 AND2X2_8086 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_107_), .Y(u2__abc_52155_new_n17167_));
AND2X2 AND2X2_8087 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17168_));
AND2X2 AND2X2_8088 ( .A(u2__abc_52155_new_n17169_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17170_));
AND2X2 AND2X2_8089 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_110_), .Y(u2__abc_52155_new_n17172_));
AND2X2 AND2X2_809 ( .A(u2__abc_52155_new_n3371_), .B(u2__abc_52155_new_n3380_), .Y(u2__abc_52155_new_n3632_));
AND2X2 AND2X2_8090 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_108_), .Y(u2__abc_52155_new_n17173_));
AND2X2 AND2X2_8091 ( .A(u2__abc_52155_new_n17174_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17175_));
AND2X2 AND2X2_8092 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_110_), .Y(u2__abc_52155_new_n17176_));
AND2X2 AND2X2_8093 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n17177_));
AND2X2 AND2X2_8094 ( .A(u2__abc_52155_new_n17178_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17179_));
AND2X2 AND2X2_8095 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_111_), .Y(u2__abc_52155_new_n17181_));
AND2X2 AND2X2_8096 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_109_), .Y(u2__abc_52155_new_n17182_));
AND2X2 AND2X2_8097 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17183_));
AND2X2 AND2X2_8098 ( .A(u2__abc_52155_new_n17184_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17185_));
AND2X2 AND2X2_8099 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_112_), .Y(u2__abc_52155_new_n17187_));
AND2X2 AND2X2_81 ( .A(_abc_73687_new_n843_), .B(_abc_73687_new_n842_), .Y(\o[116] ));
AND2X2 AND2X2_810 ( .A(u2__abc_52155_new_n3633_), .B(u2__abc_52155_new_n3368_), .Y(u2__abc_52155_new_n3634_));
AND2X2 AND2X2_8100 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_110_), .Y(u2__abc_52155_new_n17188_));
AND2X2 AND2X2_8101 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17189_));
AND2X2 AND2X2_8102 ( .A(u2__abc_52155_new_n17190_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17191_));
AND2X2 AND2X2_8103 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_113_), .Y(u2__abc_52155_new_n17193_));
AND2X2 AND2X2_8104 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_111_), .Y(u2__abc_52155_new_n17194_));
AND2X2 AND2X2_8105 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17195_));
AND2X2 AND2X2_8106 ( .A(u2__abc_52155_new_n17196_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17197_));
AND2X2 AND2X2_8107 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_114_), .Y(u2__abc_52155_new_n17199_));
AND2X2 AND2X2_8108 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_112_), .Y(u2__abc_52155_new_n17200_));
AND2X2 AND2X2_8109 ( .A(u2__abc_52155_new_n17201_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17202_));
AND2X2 AND2X2_811 ( .A(u2__abc_52155_new_n3366_), .B(u2__abc_52155_new_n3358_), .Y(u2__abc_52155_new_n3635_));
AND2X2 AND2X2_8110 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_114_), .Y(u2__abc_52155_new_n17203_));
AND2X2 AND2X2_8111 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n17204_));
AND2X2 AND2X2_8112 ( .A(u2__abc_52155_new_n17205_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17206_));
AND2X2 AND2X2_8113 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_115_), .Y(u2__abc_52155_new_n17208_));
AND2X2 AND2X2_8114 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17209_));
AND2X2 AND2X2_8115 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_113_), .Y(u2__abc_52155_new_n17210_));
AND2X2 AND2X2_8116 ( .A(u2__abc_52155_new_n17211_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17212_));
AND2X2 AND2X2_8117 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_116_), .Y(u2__abc_52155_new_n17214_));
AND2X2 AND2X2_8118 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_114_), .Y(u2__abc_52155_new_n17215_));
AND2X2 AND2X2_8119 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17216_));
AND2X2 AND2X2_812 ( .A(u2__abc_52155_new_n3624_), .B(u2__abc_52155_new_n3639_), .Y(u2__abc_52155_new_n3640_));
AND2X2 AND2X2_8120 ( .A(u2__abc_52155_new_n17217_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17218_));
AND2X2 AND2X2_8121 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_117_), .Y(u2__abc_52155_new_n17220_));
AND2X2 AND2X2_8122 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_115_), .Y(u2__abc_52155_new_n17221_));
AND2X2 AND2X2_8123 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17222_));
AND2X2 AND2X2_8124 ( .A(u2__abc_52155_new_n17223_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17224_));
AND2X2 AND2X2_8125 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_118_), .Y(u2__abc_52155_new_n17226_));
AND2X2 AND2X2_8126 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_116_), .Y(u2__abc_52155_new_n17227_));
AND2X2 AND2X2_8127 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17228_));
AND2X2 AND2X2_8128 ( .A(u2__abc_52155_new_n17229_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17230_));
AND2X2 AND2X2_8129 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_119_), .Y(u2__abc_52155_new_n17232_));
AND2X2 AND2X2_813 ( .A(u2__abc_52155_new_n3604_), .B(u2__abc_52155_new_n3640_), .Y(u2__abc_52155_new_n3641_));
AND2X2 AND2X2_8130 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_117_), .Y(u2__abc_52155_new_n17233_));
AND2X2 AND2X2_8131 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17234_));
AND2X2 AND2X2_8132 ( .A(u2__abc_52155_new_n17235_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17236_));
AND2X2 AND2X2_8133 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_120_), .Y(u2__abc_52155_new_n17238_));
AND2X2 AND2X2_8134 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_118_), .Y(u2__abc_52155_new_n17239_));
AND2X2 AND2X2_8135 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17240_));
AND2X2 AND2X2_8136 ( .A(u2__abc_52155_new_n17241_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17242_));
AND2X2 AND2X2_8137 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_121_), .Y(u2__abc_52155_new_n17244_));
AND2X2 AND2X2_8138 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17245_));
AND2X2 AND2X2_8139 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_119_), .Y(u2__abc_52155_new_n17246_));
AND2X2 AND2X2_814 ( .A(u2__abc_52155_new_n3561_), .B(u2__abc_52155_new_n3641_), .Y(u2__abc_52155_new_n3642_));
AND2X2 AND2X2_8140 ( .A(u2__abc_52155_new_n17247_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17248_));
AND2X2 AND2X2_8141 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_122_), .Y(u2__abc_52155_new_n17250_));
AND2X2 AND2X2_8142 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_120_), .Y(u2__abc_52155_new_n17251_));
AND2X2 AND2X2_8143 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17252_));
AND2X2 AND2X2_8144 ( .A(u2__abc_52155_new_n17253_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17254_));
AND2X2 AND2X2_8145 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_123_), .Y(u2__abc_52155_new_n17256_));
AND2X2 AND2X2_8146 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_121_), .Y(u2__abc_52155_new_n17257_));
AND2X2 AND2X2_8147 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17258_));
AND2X2 AND2X2_8148 ( .A(u2__abc_52155_new_n17259_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17260_));
AND2X2 AND2X2_8149 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_124_), .Y(u2__abc_52155_new_n17262_));
AND2X2 AND2X2_815 ( .A(u2__abc_52155_new_n3643_), .B(u2_remHi_118_), .Y(u2__abc_52155_new_n3644_));
AND2X2 AND2X2_8150 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_122_), .Y(u2__abc_52155_new_n17263_));
AND2X2 AND2X2_8151 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17264_));
AND2X2 AND2X2_8152 ( .A(u2__abc_52155_new_n17265_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17266_));
AND2X2 AND2X2_8153 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_125_), .Y(u2__abc_52155_new_n17268_));
AND2X2 AND2X2_8154 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17269_));
AND2X2 AND2X2_8155 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_123_), .Y(u2__abc_52155_new_n17270_));
AND2X2 AND2X2_8156 ( .A(u2__abc_52155_new_n17271_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17272_));
AND2X2 AND2X2_8157 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_126_), .Y(u2__abc_52155_new_n17274_));
AND2X2 AND2X2_8158 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_124_), .Y(u2__abc_52155_new_n17275_));
AND2X2 AND2X2_8159 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17276_));
AND2X2 AND2X2_816 ( .A(u2__abc_52155_new_n3646_), .B(sqrto_118_), .Y(u2__abc_52155_new_n3647_));
AND2X2 AND2X2_8160 ( .A(u2__abc_52155_new_n17277_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17278_));
AND2X2 AND2X2_8161 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_127_), .Y(u2__abc_52155_new_n17280_));
AND2X2 AND2X2_8162 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17281_));
AND2X2 AND2X2_8163 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_125_), .Y(u2__abc_52155_new_n17282_));
AND2X2 AND2X2_8164 ( .A(u2__abc_52155_new_n17283_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17284_));
AND2X2 AND2X2_8165 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_128_), .Y(u2__abc_52155_new_n17286_));
AND2X2 AND2X2_8166 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17287_));
AND2X2 AND2X2_8167 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_126_), .Y(u2__abc_52155_new_n17288_));
AND2X2 AND2X2_8168 ( .A(u2__abc_52155_new_n17289_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17290_));
AND2X2 AND2X2_8169 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_129_), .Y(u2__abc_52155_new_n17292_));
AND2X2 AND2X2_817 ( .A(u2__abc_52155_new_n3645_), .B(u2__abc_52155_new_n3648_), .Y(u2__abc_52155_new_n3649_));
AND2X2 AND2X2_8170 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_127_), .Y(u2__abc_52155_new_n17293_));
AND2X2 AND2X2_8171 ( .A(u2__abc_52155_new_n17294_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17295_));
AND2X2 AND2X2_8172 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_129_), .Y(u2__abc_52155_new_n17296_));
AND2X2 AND2X2_8173 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n17297_));
AND2X2 AND2X2_8174 ( .A(u2__abc_52155_new_n17298_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17299_));
AND2X2 AND2X2_8175 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_130_), .Y(u2__abc_52155_new_n17301_));
AND2X2 AND2X2_8176 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17302_));
AND2X2 AND2X2_8177 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_128_), .Y(u2__abc_52155_new_n17303_));
AND2X2 AND2X2_8178 ( .A(u2__abc_52155_new_n17304_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17305_));
AND2X2 AND2X2_8179 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_131_), .Y(u2__abc_52155_new_n17307_));
AND2X2 AND2X2_818 ( .A(u2__abc_52155_new_n3650_), .B(u2_remHi_119_), .Y(u2__abc_52155_new_n3651_));
AND2X2 AND2X2_8180 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_129_), .Y(u2__abc_52155_new_n17308_));
AND2X2 AND2X2_8181 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17309_));
AND2X2 AND2X2_8182 ( .A(u2__abc_52155_new_n17310_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17311_));
AND2X2 AND2X2_8183 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_132_), .Y(u2__abc_52155_new_n17313_));
AND2X2 AND2X2_8184 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_130_), .Y(u2__abc_52155_new_n17314_));
AND2X2 AND2X2_8185 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17315_));
AND2X2 AND2X2_8186 ( .A(u2__abc_52155_new_n17316_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17317_));
AND2X2 AND2X2_8187 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_133_), .Y(u2__abc_52155_new_n17319_));
AND2X2 AND2X2_8188 ( .A(u2__abc_52155_new_n17085_), .B(1'h0), .Y(u2__abc_52155_new_n17320_));
AND2X2 AND2X2_8189 ( .A(u2__abc_52155_new_n2982_), .B(u2_remLo_131_), .Y(u2__abc_52155_new_n17321_));
AND2X2 AND2X2_819 ( .A(u2__abc_52155_new_n3653_), .B(sqrto_119_), .Y(u2__abc_52155_new_n3654_));
AND2X2 AND2X2_8190 ( .A(u2__abc_52155_new_n16683_), .B(u2__abc_52155_new_n17321_), .Y(u2__abc_52155_new_n17322_));
AND2X2 AND2X2_8191 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_134_), .Y(u2__abc_52155_new_n17325_));
AND2X2 AND2X2_8192 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17326_));
AND2X2 AND2X2_8193 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_132_), .Y(u2__abc_52155_new_n17327_));
AND2X2 AND2X2_8194 ( .A(u2__abc_52155_new_n17328_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17329_));
AND2X2 AND2X2_8195 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_135_), .Y(u2__abc_52155_new_n17331_));
AND2X2 AND2X2_8196 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_133_), .Y(u2__abc_52155_new_n17332_));
AND2X2 AND2X2_8197 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17333_));
AND2X2 AND2X2_8198 ( .A(u2__abc_52155_new_n17334_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17335_));
AND2X2 AND2X2_8199 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_136_), .Y(u2__abc_52155_new_n17337_));
AND2X2 AND2X2_82 ( .A(_abc_73687_new_n846_), .B(_abc_73687_new_n845_), .Y(\o[117] ));
AND2X2 AND2X2_820 ( .A(u2__abc_52155_new_n3652_), .B(u2__abc_52155_new_n3655_), .Y(u2__abc_52155_new_n3656_));
AND2X2 AND2X2_8200 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_134_), .Y(u2__abc_52155_new_n17338_));
AND2X2 AND2X2_8201 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17339_));
AND2X2 AND2X2_8202 ( .A(u2__abc_52155_new_n17340_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17341_));
AND2X2 AND2X2_8203 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_137_), .Y(u2__abc_52155_new_n17343_));
AND2X2 AND2X2_8204 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_135_), .Y(u2__abc_52155_new_n17344_));
AND2X2 AND2X2_8205 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17345_));
AND2X2 AND2X2_8206 ( .A(u2__abc_52155_new_n17346_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17347_));
AND2X2 AND2X2_8207 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_138_), .Y(u2__abc_52155_new_n17349_));
AND2X2 AND2X2_8208 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17350_));
AND2X2 AND2X2_8209 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_136_), .Y(u2__abc_52155_new_n17351_));
AND2X2 AND2X2_821 ( .A(u2__abc_52155_new_n3649_), .B(u2__abc_52155_new_n3656_), .Y(u2__abc_52155_new_n3657_));
AND2X2 AND2X2_8210 ( .A(u2__abc_52155_new_n17352_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17353_));
AND2X2 AND2X2_8211 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_139_), .Y(u2__abc_52155_new_n17355_));
AND2X2 AND2X2_8212 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_137_), .Y(u2__abc_52155_new_n17356_));
AND2X2 AND2X2_8213 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17357_));
AND2X2 AND2X2_8214 ( .A(u2__abc_52155_new_n17358_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17359_));
AND2X2 AND2X2_8215 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_140_), .Y(u2__abc_52155_new_n17361_));
AND2X2 AND2X2_8216 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_138_), .Y(u2__abc_52155_new_n17362_));
AND2X2 AND2X2_8217 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17363_));
AND2X2 AND2X2_8218 ( .A(u2__abc_52155_new_n17364_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17365_));
AND2X2 AND2X2_8219 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_141_), .Y(u2__abc_52155_new_n17367_));
AND2X2 AND2X2_822 ( .A(u2__abc_52155_new_n3658_), .B(u2_remHi_120_), .Y(u2__abc_52155_new_n3659_));
AND2X2 AND2X2_8220 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_139_), .Y(u2__abc_52155_new_n17368_));
AND2X2 AND2X2_8221 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17369_));
AND2X2 AND2X2_8222 ( .A(u2__abc_52155_new_n17370_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17371_));
AND2X2 AND2X2_8223 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_142_), .Y(u2__abc_52155_new_n17373_));
AND2X2 AND2X2_8224 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_140_), .Y(u2__abc_52155_new_n17374_));
AND2X2 AND2X2_8225 ( .A(u2__abc_52155_new_n17375_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17376_));
AND2X2 AND2X2_8226 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_142_), .Y(u2__abc_52155_new_n17377_));
AND2X2 AND2X2_8227 ( .A(u2__abc_52155_new_n2964_), .B(1'h0), .Y(u2__abc_52155_new_n17378_));
AND2X2 AND2X2_8228 ( .A(u2__abc_52155_new_n17379_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17380_));
AND2X2 AND2X2_8229 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_143_), .Y(u2__abc_52155_new_n17382_));
AND2X2 AND2X2_823 ( .A(u2__abc_52155_new_n3661_), .B(sqrto_120_), .Y(u2__abc_52155_new_n3662_));
AND2X2 AND2X2_8230 ( .A(u2__abc_52155_new_n2963_), .B(1'h0), .Y(u2__abc_52155_new_n17383_));
AND2X2 AND2X2_8231 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_141_), .Y(u2__abc_52155_new_n17384_));
AND2X2 AND2X2_8232 ( .A(u2__abc_52155_new_n17385_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17386_));
AND2X2 AND2X2_8233 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_144_), .Y(u2__abc_52155_new_n17388_));
AND2X2 AND2X2_8234 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_142_), .Y(u2__abc_52155_new_n17389_));
AND2X2 AND2X2_8235 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_0_), .Y(u2__abc_52155_new_n17390_));
AND2X2 AND2X2_8236 ( .A(u2__abc_52155_new_n17391_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17392_));
AND2X2 AND2X2_8237 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_145_), .Y(u2__abc_52155_new_n17394_));
AND2X2 AND2X2_8238 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_143_), .Y(u2__abc_52155_new_n17395_));
AND2X2 AND2X2_8239 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_1_), .Y(u2__abc_52155_new_n17396_));
AND2X2 AND2X2_824 ( .A(u2__abc_52155_new_n3660_), .B(u2__abc_52155_new_n3663_), .Y(u2__abc_52155_new_n3664_));
AND2X2 AND2X2_8240 ( .A(u2__abc_52155_new_n17397_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17398_));
AND2X2 AND2X2_8241 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_146_), .Y(u2__abc_52155_new_n17400_));
AND2X2 AND2X2_8242 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_144_), .Y(u2__abc_52155_new_n17401_));
AND2X2 AND2X2_8243 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_2_), .Y(u2__abc_52155_new_n17402_));
AND2X2 AND2X2_8244 ( .A(u2__abc_52155_new_n17403_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17404_));
AND2X2 AND2X2_8245 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_147_), .Y(u2__abc_52155_new_n17406_));
AND2X2 AND2X2_8246 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_3_), .Y(u2__abc_52155_new_n17407_));
AND2X2 AND2X2_8247 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_145_), .Y(u2__abc_52155_new_n17408_));
AND2X2 AND2X2_8248 ( .A(u2__abc_52155_new_n17409_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17410_));
AND2X2 AND2X2_8249 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_148_), .Y(u2__abc_52155_new_n17412_));
AND2X2 AND2X2_825 ( .A(u2__abc_52155_new_n3665_), .B(u2_remHi_121_), .Y(u2__abc_52155_new_n3666_));
AND2X2 AND2X2_8250 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_146_), .Y(u2__abc_52155_new_n17413_));
AND2X2 AND2X2_8251 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_4_), .Y(u2__abc_52155_new_n17414_));
AND2X2 AND2X2_8252 ( .A(u2__abc_52155_new_n17415_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17416_));
AND2X2 AND2X2_8253 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_149_), .Y(u2__abc_52155_new_n17418_));
AND2X2 AND2X2_8254 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_147_), .Y(u2__abc_52155_new_n17419_));
AND2X2 AND2X2_8255 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_5_), .Y(u2__abc_52155_new_n17420_));
AND2X2 AND2X2_8256 ( .A(u2__abc_52155_new_n17421_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17422_));
AND2X2 AND2X2_8257 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_150_), .Y(u2__abc_52155_new_n17424_));
AND2X2 AND2X2_8258 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_148_), .Y(u2__abc_52155_new_n17425_));
AND2X2 AND2X2_8259 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_6_), .Y(u2__abc_52155_new_n17426_));
AND2X2 AND2X2_826 ( .A(u2__abc_52155_new_n3668_), .B(sqrto_121_), .Y(u2__abc_52155_new_n3669_));
AND2X2 AND2X2_8260 ( .A(u2__abc_52155_new_n17427_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17428_));
AND2X2 AND2X2_8261 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_151_), .Y(u2__abc_52155_new_n17430_));
AND2X2 AND2X2_8262 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_149_), .Y(u2__abc_52155_new_n17431_));
AND2X2 AND2X2_8263 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_7_), .Y(u2__abc_52155_new_n17432_));
AND2X2 AND2X2_8264 ( .A(u2__abc_52155_new_n17433_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17434_));
AND2X2 AND2X2_8265 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_152_), .Y(u2__abc_52155_new_n17436_));
AND2X2 AND2X2_8266 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_150_), .Y(u2__abc_52155_new_n17437_));
AND2X2 AND2X2_8267 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_8_), .Y(u2__abc_52155_new_n17438_));
AND2X2 AND2X2_8268 ( .A(u2__abc_52155_new_n17439_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17440_));
AND2X2 AND2X2_8269 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_153_), .Y(u2__abc_52155_new_n17442_));
AND2X2 AND2X2_827 ( .A(u2__abc_52155_new_n3667_), .B(u2__abc_52155_new_n3670_), .Y(u2__abc_52155_new_n3671_));
AND2X2 AND2X2_8270 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_9_), .Y(u2__abc_52155_new_n17443_));
AND2X2 AND2X2_8271 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_151_), .Y(u2__abc_52155_new_n17444_));
AND2X2 AND2X2_8272 ( .A(u2__abc_52155_new_n17445_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17446_));
AND2X2 AND2X2_8273 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_154_), .Y(u2__abc_52155_new_n17448_));
AND2X2 AND2X2_8274 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_10_), .Y(u2__abc_52155_new_n17449_));
AND2X2 AND2X2_8275 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_152_), .Y(u2__abc_52155_new_n17450_));
AND2X2 AND2X2_8276 ( .A(u2__abc_52155_new_n17451_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17452_));
AND2X2 AND2X2_8277 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_155_), .Y(u2__abc_52155_new_n17454_));
AND2X2 AND2X2_8278 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_153_), .Y(u2__abc_52155_new_n17455_));
AND2X2 AND2X2_8279 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_11_), .Y(u2__abc_52155_new_n17456_));
AND2X2 AND2X2_828 ( .A(u2__abc_52155_new_n3664_), .B(u2__abc_52155_new_n3671_), .Y(u2__abc_52155_new_n3672_));
AND2X2 AND2X2_8280 ( .A(u2__abc_52155_new_n17457_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17458_));
AND2X2 AND2X2_8281 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_156_), .Y(u2__abc_52155_new_n17460_));
AND2X2 AND2X2_8282 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_154_), .Y(u2__abc_52155_new_n17461_));
AND2X2 AND2X2_8283 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_12_), .Y(u2__abc_52155_new_n17462_));
AND2X2 AND2X2_8284 ( .A(u2__abc_52155_new_n17463_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17464_));
AND2X2 AND2X2_8285 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_157_), .Y(u2__abc_52155_new_n17466_));
AND2X2 AND2X2_8286 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_155_), .Y(u2__abc_52155_new_n17467_));
AND2X2 AND2X2_8287 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_13_), .Y(u2__abc_52155_new_n17468_));
AND2X2 AND2X2_8288 ( .A(u2__abc_52155_new_n17469_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17470_));
AND2X2 AND2X2_8289 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_158_), .Y(u2__abc_52155_new_n17472_));
AND2X2 AND2X2_829 ( .A(u2__abc_52155_new_n3657_), .B(u2__abc_52155_new_n3672_), .Y(u2__abc_52155_new_n3673_));
AND2X2 AND2X2_8290 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_156_), .Y(u2__abc_52155_new_n17473_));
AND2X2 AND2X2_8291 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_14_), .Y(u2__abc_52155_new_n17474_));
AND2X2 AND2X2_8292 ( .A(u2__abc_52155_new_n17475_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17476_));
AND2X2 AND2X2_8293 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_159_), .Y(u2__abc_52155_new_n17478_));
AND2X2 AND2X2_8294 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_157_), .Y(u2__abc_52155_new_n17479_));
AND2X2 AND2X2_8295 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_15_), .Y(u2__abc_52155_new_n17480_));
AND2X2 AND2X2_8296 ( .A(u2__abc_52155_new_n17481_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17482_));
AND2X2 AND2X2_8297 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_160_), .Y(u2__abc_52155_new_n17484_));
AND2X2 AND2X2_8298 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_158_), .Y(u2__abc_52155_new_n17485_));
AND2X2 AND2X2_8299 ( .A(u2__abc_52155_new_n17486_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17487_));
AND2X2 AND2X2_83 ( .A(_abc_73687_new_n849_), .B(_abc_73687_new_n848_), .Y(\o[118] ));
AND2X2 AND2X2_830 ( .A(u2__abc_52155_new_n3674_), .B(u2_remHi_124_), .Y(u2__abc_52155_new_n3675_));
AND2X2 AND2X2_8300 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_160_), .Y(u2__abc_52155_new_n17488_));
AND2X2 AND2X2_8301 ( .A(u2__abc_52155_new_n2964_), .B(fracta1_16_), .Y(u2__abc_52155_new_n17489_));
AND2X2 AND2X2_8302 ( .A(u2__abc_52155_new_n17490_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17491_));
AND2X2 AND2X2_8303 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_161_), .Y(u2__abc_52155_new_n17493_));
AND2X2 AND2X2_8304 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_159_), .Y(u2__abc_52155_new_n17494_));
AND2X2 AND2X2_8305 ( .A(u2__abc_52155_new_n17495_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17496_));
AND2X2 AND2X2_8306 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_161_), .Y(u2__abc_52155_new_n17497_));
AND2X2 AND2X2_8307 ( .A(u2__abc_52155_new_n2964_), .B(fracta1_17_), .Y(u2__abc_52155_new_n17498_));
AND2X2 AND2X2_8308 ( .A(u2__abc_52155_new_n17499_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17500_));
AND2X2 AND2X2_8309 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_162_), .Y(u2__abc_52155_new_n17502_));
AND2X2 AND2X2_831 ( .A(u2__abc_52155_new_n3677_), .B(sqrto_124_), .Y(u2__abc_52155_new_n3678_));
AND2X2 AND2X2_8310 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_160_), .Y(u2__abc_52155_new_n17503_));
AND2X2 AND2X2_8311 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_18_), .Y(u2__abc_52155_new_n17504_));
AND2X2 AND2X2_8312 ( .A(u2__abc_52155_new_n17505_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17506_));
AND2X2 AND2X2_8313 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_163_), .Y(u2__abc_52155_new_n17508_));
AND2X2 AND2X2_8314 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_161_), .Y(u2__abc_52155_new_n17509_));
AND2X2 AND2X2_8315 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_19_), .Y(u2__abc_52155_new_n17510_));
AND2X2 AND2X2_8316 ( .A(u2__abc_52155_new_n17511_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17512_));
AND2X2 AND2X2_8317 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_164_), .Y(u2__abc_52155_new_n17514_));
AND2X2 AND2X2_8318 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_162_), .Y(u2__abc_52155_new_n17515_));
AND2X2 AND2X2_8319 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_20_), .Y(u2__abc_52155_new_n17516_));
AND2X2 AND2X2_832 ( .A(u2__abc_52155_new_n3676_), .B(u2__abc_52155_new_n3679_), .Y(u2__abc_52155_new_n3680_));
AND2X2 AND2X2_8320 ( .A(u2__abc_52155_new_n17517_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17518_));
AND2X2 AND2X2_8321 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_165_), .Y(u2__abc_52155_new_n17520_));
AND2X2 AND2X2_8322 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_163_), .Y(u2__abc_52155_new_n17521_));
AND2X2 AND2X2_8323 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_21_), .Y(u2__abc_52155_new_n17522_));
AND2X2 AND2X2_8324 ( .A(u2__abc_52155_new_n17523_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17524_));
AND2X2 AND2X2_8325 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_166_), .Y(u2__abc_52155_new_n17526_));
AND2X2 AND2X2_8326 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_22_), .Y(u2__abc_52155_new_n17527_));
AND2X2 AND2X2_8327 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_164_), .Y(u2__abc_52155_new_n17528_));
AND2X2 AND2X2_8328 ( .A(u2__abc_52155_new_n17529_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17530_));
AND2X2 AND2X2_8329 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_167_), .Y(u2__abc_52155_new_n17532_));
AND2X2 AND2X2_833 ( .A(u2__abc_52155_new_n3681_), .B(sqrto_125_), .Y(u2__abc_52155_new_n3682_));
AND2X2 AND2X2_8330 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_165_), .Y(u2__abc_52155_new_n17533_));
AND2X2 AND2X2_8331 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_23_), .Y(u2__abc_52155_new_n17534_));
AND2X2 AND2X2_8332 ( .A(u2__abc_52155_new_n17535_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17536_));
AND2X2 AND2X2_8333 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_168_), .Y(u2__abc_52155_new_n17538_));
AND2X2 AND2X2_8334 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_166_), .Y(u2__abc_52155_new_n17539_));
AND2X2 AND2X2_8335 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_24_), .Y(u2__abc_52155_new_n17540_));
AND2X2 AND2X2_8336 ( .A(u2__abc_52155_new_n17541_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17542_));
AND2X2 AND2X2_8337 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_169_), .Y(u2__abc_52155_new_n17544_));
AND2X2 AND2X2_8338 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_167_), .Y(u2__abc_52155_new_n17545_));
AND2X2 AND2X2_8339 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_25_), .Y(u2__abc_52155_new_n17546_));
AND2X2 AND2X2_834 ( .A(u2__abc_52155_new_n3684_), .B(u2_remHi_125_), .Y(u2__abc_52155_new_n3685_));
AND2X2 AND2X2_8340 ( .A(u2__abc_52155_new_n17547_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17548_));
AND2X2 AND2X2_8341 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_170_), .Y(u2__abc_52155_new_n17550_));
AND2X2 AND2X2_8342 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_26_), .Y(u2__abc_52155_new_n17551_));
AND2X2 AND2X2_8343 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_168_), .Y(u2__abc_52155_new_n17552_));
AND2X2 AND2X2_8344 ( .A(u2__abc_52155_new_n17553_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17554_));
AND2X2 AND2X2_8345 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_171_), .Y(u2__abc_52155_new_n17556_));
AND2X2 AND2X2_8346 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_169_), .Y(u2__abc_52155_new_n17557_));
AND2X2 AND2X2_8347 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_27_), .Y(u2__abc_52155_new_n17558_));
AND2X2 AND2X2_8348 ( .A(u2__abc_52155_new_n17559_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17560_));
AND2X2 AND2X2_8349 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_172_), .Y(u2__abc_52155_new_n17562_));
AND2X2 AND2X2_835 ( .A(u2__abc_52155_new_n3683_), .B(u2__abc_52155_new_n3686_), .Y(u2__abc_52155_new_n3687_));
AND2X2 AND2X2_8350 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_170_), .Y(u2__abc_52155_new_n17563_));
AND2X2 AND2X2_8351 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_28_), .Y(u2__abc_52155_new_n17564_));
AND2X2 AND2X2_8352 ( .A(u2__abc_52155_new_n17565_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17566_));
AND2X2 AND2X2_8353 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_173_), .Y(u2__abc_52155_new_n17568_));
AND2X2 AND2X2_8354 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_171_), .Y(u2__abc_52155_new_n17569_));
AND2X2 AND2X2_8355 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_29_), .Y(u2__abc_52155_new_n17570_));
AND2X2 AND2X2_8356 ( .A(u2__abc_52155_new_n17571_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17572_));
AND2X2 AND2X2_8357 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_174_), .Y(u2__abc_52155_new_n17574_));
AND2X2 AND2X2_8358 ( .A(u2__abc_52155_new_n17085_), .B(fracta1_30_), .Y(u2__abc_52155_new_n17575_));
AND2X2 AND2X2_8359 ( .A(u2__abc_52155_new_n2982_), .B(u2_remLo_172_), .Y(u2__abc_52155_new_n17576_));
AND2X2 AND2X2_836 ( .A(u2__abc_52155_new_n3680_), .B(u2__abc_52155_new_n3687_), .Y(u2__abc_52155_new_n3688_));
AND2X2 AND2X2_8360 ( .A(u2__abc_52155_new_n16683_), .B(u2__abc_52155_new_n17576_), .Y(u2__abc_52155_new_n17577_));
AND2X2 AND2X2_8361 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_175_), .Y(u2__abc_52155_new_n17580_));
AND2X2 AND2X2_8362 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_173_), .Y(u2__abc_52155_new_n17581_));
AND2X2 AND2X2_8363 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_31_), .Y(u2__abc_52155_new_n17582_));
AND2X2 AND2X2_8364 ( .A(u2__abc_52155_new_n17583_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17584_));
AND2X2 AND2X2_8365 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_176_), .Y(u2__abc_52155_new_n17586_));
AND2X2 AND2X2_8366 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_174_), .Y(u2__abc_52155_new_n17587_));
AND2X2 AND2X2_8367 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_32_), .Y(u2__abc_52155_new_n17588_));
AND2X2 AND2X2_8368 ( .A(u2__abc_52155_new_n17589_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17590_));
AND2X2 AND2X2_8369 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_177_), .Y(u2__abc_52155_new_n17592_));
AND2X2 AND2X2_837 ( .A(u2__abc_52155_new_n3689_), .B(u2_remHi_123_), .Y(u2__abc_52155_new_n3690_));
AND2X2 AND2X2_8370 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_175_), .Y(u2__abc_52155_new_n17593_));
AND2X2 AND2X2_8371 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_33_), .Y(u2__abc_52155_new_n17594_));
AND2X2 AND2X2_8372 ( .A(u2__abc_52155_new_n17595_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17596_));
AND2X2 AND2X2_8373 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_178_), .Y(u2__abc_52155_new_n17598_));
AND2X2 AND2X2_8374 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_176_), .Y(u2__abc_52155_new_n17599_));
AND2X2 AND2X2_8375 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_34_), .Y(u2__abc_52155_new_n17600_));
AND2X2 AND2X2_8376 ( .A(u2__abc_52155_new_n17601_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17602_));
AND2X2 AND2X2_8377 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_179_), .Y(u2__abc_52155_new_n17604_));
AND2X2 AND2X2_8378 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_177_), .Y(u2__abc_52155_new_n17605_));
AND2X2 AND2X2_8379 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_35_), .Y(u2__abc_52155_new_n17606_));
AND2X2 AND2X2_838 ( .A(u2__abc_52155_new_n3692_), .B(sqrto_123_), .Y(u2__abc_52155_new_n3693_));
AND2X2 AND2X2_8380 ( .A(u2__abc_52155_new_n17607_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17608_));
AND2X2 AND2X2_8381 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_180_), .Y(u2__abc_52155_new_n17610_));
AND2X2 AND2X2_8382 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_178_), .Y(u2__abc_52155_new_n17611_));
AND2X2 AND2X2_8383 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_36_), .Y(u2__abc_52155_new_n17612_));
AND2X2 AND2X2_8384 ( .A(u2__abc_52155_new_n17613_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17614_));
AND2X2 AND2X2_8385 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_181_), .Y(u2__abc_52155_new_n17616_));
AND2X2 AND2X2_8386 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_179_), .Y(u2__abc_52155_new_n17617_));
AND2X2 AND2X2_8387 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_37_), .Y(u2__abc_52155_new_n17618_));
AND2X2 AND2X2_8388 ( .A(u2__abc_52155_new_n17619_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17620_));
AND2X2 AND2X2_8389 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_182_), .Y(u2__abc_52155_new_n17622_));
AND2X2 AND2X2_839 ( .A(u2__abc_52155_new_n3691_), .B(u2__abc_52155_new_n3694_), .Y(u2__abc_52155_new_n3695_));
AND2X2 AND2X2_8390 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_180_), .Y(u2__abc_52155_new_n17623_));
AND2X2 AND2X2_8391 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_38_), .Y(u2__abc_52155_new_n17624_));
AND2X2 AND2X2_8392 ( .A(u2__abc_52155_new_n17625_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17626_));
AND2X2 AND2X2_8393 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_183_), .Y(u2__abc_52155_new_n17628_));
AND2X2 AND2X2_8394 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_181_), .Y(u2__abc_52155_new_n17629_));
AND2X2 AND2X2_8395 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_39_), .Y(u2__abc_52155_new_n17630_));
AND2X2 AND2X2_8396 ( .A(u2__abc_52155_new_n17631_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17632_));
AND2X2 AND2X2_8397 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_184_), .Y(u2__abc_52155_new_n17634_));
AND2X2 AND2X2_8398 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_182_), .Y(u2__abc_52155_new_n17635_));
AND2X2 AND2X2_8399 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_40_), .Y(u2__abc_52155_new_n17636_));
AND2X2 AND2X2_84 ( .A(_abc_73687_new_n852_), .B(_abc_73687_new_n851_), .Y(\o[119] ));
AND2X2 AND2X2_840 ( .A(u2__abc_52155_new_n3696_), .B(u2_remHi_122_), .Y(u2__abc_52155_new_n3697_));
AND2X2 AND2X2_8400 ( .A(u2__abc_52155_new_n17637_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17638_));
AND2X2 AND2X2_8401 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_185_), .Y(u2__abc_52155_new_n17640_));
AND2X2 AND2X2_8402 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_41_), .Y(u2__abc_52155_new_n17641_));
AND2X2 AND2X2_8403 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_183_), .Y(u2__abc_52155_new_n17642_));
AND2X2 AND2X2_8404 ( .A(u2__abc_52155_new_n17643_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17644_));
AND2X2 AND2X2_8405 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_186_), .Y(u2__abc_52155_new_n17646_));
AND2X2 AND2X2_8406 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_42_), .Y(u2__abc_52155_new_n17647_));
AND2X2 AND2X2_8407 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_184_), .Y(u2__abc_52155_new_n17648_));
AND2X2 AND2X2_8408 ( .A(u2__abc_52155_new_n17649_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17650_));
AND2X2 AND2X2_8409 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_187_), .Y(u2__abc_52155_new_n17652_));
AND2X2 AND2X2_841 ( .A(u2__abc_52155_new_n3699_), .B(sqrto_122_), .Y(u2__abc_52155_new_n3700_));
AND2X2 AND2X2_8410 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_185_), .Y(u2__abc_52155_new_n17653_));
AND2X2 AND2X2_8411 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_43_), .Y(u2__abc_52155_new_n17654_));
AND2X2 AND2X2_8412 ( .A(u2__abc_52155_new_n17655_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17656_));
AND2X2 AND2X2_8413 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_188_), .Y(u2__abc_52155_new_n17658_));
AND2X2 AND2X2_8414 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_186_), .Y(u2__abc_52155_new_n17659_));
AND2X2 AND2X2_8415 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_44_), .Y(u2__abc_52155_new_n17660_));
AND2X2 AND2X2_8416 ( .A(u2__abc_52155_new_n17661_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17662_));
AND2X2 AND2X2_8417 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_189_), .Y(u2__abc_52155_new_n17664_));
AND2X2 AND2X2_8418 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_45_), .Y(u2__abc_52155_new_n17665_));
AND2X2 AND2X2_8419 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_187_), .Y(u2__abc_52155_new_n17666_));
AND2X2 AND2X2_842 ( .A(u2__abc_52155_new_n3698_), .B(u2__abc_52155_new_n3701_), .Y(u2__abc_52155_new_n3702_));
AND2X2 AND2X2_8420 ( .A(u2__abc_52155_new_n17667_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17668_));
AND2X2 AND2X2_8421 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_190_), .Y(u2__abc_52155_new_n17670_));
AND2X2 AND2X2_8422 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_188_), .Y(u2__abc_52155_new_n17671_));
AND2X2 AND2X2_8423 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_46_), .Y(u2__abc_52155_new_n17672_));
AND2X2 AND2X2_8424 ( .A(u2__abc_52155_new_n17673_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17674_));
AND2X2 AND2X2_8425 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_191_), .Y(u2__abc_52155_new_n17676_));
AND2X2 AND2X2_8426 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_47_), .Y(u2__abc_52155_new_n17677_));
AND2X2 AND2X2_8427 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_189_), .Y(u2__abc_52155_new_n17678_));
AND2X2 AND2X2_8428 ( .A(u2__abc_52155_new_n17679_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17680_));
AND2X2 AND2X2_8429 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_192_), .Y(u2__abc_52155_new_n17682_));
AND2X2 AND2X2_843 ( .A(u2__abc_52155_new_n3695_), .B(u2__abc_52155_new_n3702_), .Y(u2__abc_52155_new_n3703_));
AND2X2 AND2X2_8430 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_48_), .Y(u2__abc_52155_new_n17683_));
AND2X2 AND2X2_8431 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_190_), .Y(u2__abc_52155_new_n17684_));
AND2X2 AND2X2_8432 ( .A(u2__abc_52155_new_n17685_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17686_));
AND2X2 AND2X2_8433 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_193_), .Y(u2__abc_52155_new_n17688_));
AND2X2 AND2X2_8434 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_191_), .Y(u2__abc_52155_new_n17689_));
AND2X2 AND2X2_8435 ( .A(u2__abc_52155_new_n17690_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17691_));
AND2X2 AND2X2_8436 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_193_), .Y(u2__abc_52155_new_n17692_));
AND2X2 AND2X2_8437 ( .A(u2__abc_52155_new_n2964_), .B(fracta1_49_), .Y(u2__abc_52155_new_n17693_));
AND2X2 AND2X2_8438 ( .A(u2__abc_52155_new_n17694_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17695_));
AND2X2 AND2X2_8439 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_194_), .Y(u2__abc_52155_new_n17697_));
AND2X2 AND2X2_844 ( .A(u2__abc_52155_new_n3688_), .B(u2__abc_52155_new_n3703_), .Y(u2__abc_52155_new_n3704_));
AND2X2 AND2X2_8440 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_192_), .Y(u2__abc_52155_new_n17698_));
AND2X2 AND2X2_8441 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_50_), .Y(u2__abc_52155_new_n17699_));
AND2X2 AND2X2_8442 ( .A(u2__abc_52155_new_n17700_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17701_));
AND2X2 AND2X2_8443 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_195_), .Y(u2__abc_52155_new_n17703_));
AND2X2 AND2X2_8444 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_193_), .Y(u2__abc_52155_new_n17704_));
AND2X2 AND2X2_8445 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_51_), .Y(u2__abc_52155_new_n17705_));
AND2X2 AND2X2_8446 ( .A(u2__abc_52155_new_n17706_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17707_));
AND2X2 AND2X2_8447 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_196_), .Y(u2__abc_52155_new_n17709_));
AND2X2 AND2X2_8448 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_194_), .Y(u2__abc_52155_new_n17710_));
AND2X2 AND2X2_8449 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_52_), .Y(u2__abc_52155_new_n17711_));
AND2X2 AND2X2_845 ( .A(u2__abc_52155_new_n3673_), .B(u2__abc_52155_new_n3704_), .Y(u2__abc_52155_new_n3705_));
AND2X2 AND2X2_8450 ( .A(u2__abc_52155_new_n17712_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17713_));
AND2X2 AND2X2_8451 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_197_), .Y(u2__abc_52155_new_n17715_));
AND2X2 AND2X2_8452 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_195_), .Y(u2__abc_52155_new_n17716_));
AND2X2 AND2X2_8453 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_53_), .Y(u2__abc_52155_new_n17717_));
AND2X2 AND2X2_8454 ( .A(u2__abc_52155_new_n17718_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17719_));
AND2X2 AND2X2_8455 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_198_), .Y(u2__abc_52155_new_n17721_));
AND2X2 AND2X2_8456 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_54_), .Y(u2__abc_52155_new_n17722_));
AND2X2 AND2X2_8457 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_196_), .Y(u2__abc_52155_new_n17723_));
AND2X2 AND2X2_8458 ( .A(u2__abc_52155_new_n17724_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17725_));
AND2X2 AND2X2_8459 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_199_), .Y(u2__abc_52155_new_n17727_));
AND2X2 AND2X2_846 ( .A(u2__abc_52155_new_n3706_), .B(u2_remHi_110_), .Y(u2__abc_52155_new_n3707_));
AND2X2 AND2X2_8460 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_197_), .Y(u2__abc_52155_new_n17728_));
AND2X2 AND2X2_8461 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_55_), .Y(u2__abc_52155_new_n17729_));
AND2X2 AND2X2_8462 ( .A(u2__abc_52155_new_n17730_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17731_));
AND2X2 AND2X2_8463 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_200_), .Y(u2__abc_52155_new_n17733_));
AND2X2 AND2X2_8464 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_198_), .Y(u2__abc_52155_new_n17734_));
AND2X2 AND2X2_8465 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_56_), .Y(u2__abc_52155_new_n17735_));
AND2X2 AND2X2_8466 ( .A(u2__abc_52155_new_n17736_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17737_));
AND2X2 AND2X2_8467 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_201_), .Y(u2__abc_52155_new_n17739_));
AND2X2 AND2X2_8468 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_199_), .Y(u2__abc_52155_new_n17740_));
AND2X2 AND2X2_8469 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_57_), .Y(u2__abc_52155_new_n17741_));
AND2X2 AND2X2_847 ( .A(u2__abc_52155_new_n3709_), .B(sqrto_110_), .Y(u2__abc_52155_new_n3710_));
AND2X2 AND2X2_8470 ( .A(u2__abc_52155_new_n17742_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17743_));
AND2X2 AND2X2_8471 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_202_), .Y(u2__abc_52155_new_n17745_));
AND2X2 AND2X2_8472 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_200_), .Y(u2__abc_52155_new_n17746_));
AND2X2 AND2X2_8473 ( .A(u2__abc_52155_new_n17747_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17748_));
AND2X2 AND2X2_8474 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_202_), .Y(u2__abc_52155_new_n17749_));
AND2X2 AND2X2_8475 ( .A(u2__abc_52155_new_n2964_), .B(fracta1_58_), .Y(u2__abc_52155_new_n17750_));
AND2X2 AND2X2_8476 ( .A(u2__abc_52155_new_n17751_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17752_));
AND2X2 AND2X2_8477 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_203_), .Y(u2__abc_52155_new_n17754_));
AND2X2 AND2X2_8478 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_201_), .Y(u2__abc_52155_new_n17755_));
AND2X2 AND2X2_8479 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_59_), .Y(u2__abc_52155_new_n17756_));
AND2X2 AND2X2_848 ( .A(u2__abc_52155_new_n3708_), .B(u2__abc_52155_new_n3711_), .Y(u2__abc_52155_new_n3712_));
AND2X2 AND2X2_8480 ( .A(u2__abc_52155_new_n17757_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17758_));
AND2X2 AND2X2_8481 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_204_), .Y(u2__abc_52155_new_n17760_));
AND2X2 AND2X2_8482 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_202_), .Y(u2__abc_52155_new_n17761_));
AND2X2 AND2X2_8483 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_60_), .Y(u2__abc_52155_new_n17762_));
AND2X2 AND2X2_8484 ( .A(u2__abc_52155_new_n17763_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17764_));
AND2X2 AND2X2_8485 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_205_), .Y(u2__abc_52155_new_n17766_));
AND2X2 AND2X2_8486 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_203_), .Y(u2__abc_52155_new_n17767_));
AND2X2 AND2X2_8487 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_61_), .Y(u2__abc_52155_new_n17768_));
AND2X2 AND2X2_8488 ( .A(u2__abc_52155_new_n17769_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17770_));
AND2X2 AND2X2_8489 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_206_), .Y(u2__abc_52155_new_n17772_));
AND2X2 AND2X2_849 ( .A(u2__abc_52155_new_n3713_), .B(u2_remHi_111_), .Y(u2__abc_52155_new_n3714_));
AND2X2 AND2X2_8490 ( .A(u2__abc_52155_new_n17085_), .B(fracta1_62_), .Y(u2__abc_52155_new_n17773_));
AND2X2 AND2X2_8491 ( .A(u2__abc_52155_new_n2982_), .B(u2_remLo_204_), .Y(u2__abc_52155_new_n17774_));
AND2X2 AND2X2_8492 ( .A(u2__abc_52155_new_n16683_), .B(u2__abc_52155_new_n17774_), .Y(u2__abc_52155_new_n17775_));
AND2X2 AND2X2_8493 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_207_), .Y(u2__abc_52155_new_n17778_));
AND2X2 AND2X2_8494 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_63_), .Y(u2__abc_52155_new_n17779_));
AND2X2 AND2X2_8495 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_205_), .Y(u2__abc_52155_new_n17780_));
AND2X2 AND2X2_8496 ( .A(u2__abc_52155_new_n17781_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17782_));
AND2X2 AND2X2_8497 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_208_), .Y(u2__abc_52155_new_n17784_));
AND2X2 AND2X2_8498 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_206_), .Y(u2__abc_52155_new_n17785_));
AND2X2 AND2X2_8499 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_64_), .Y(u2__abc_52155_new_n17786_));
AND2X2 AND2X2_85 ( .A(_abc_73687_new_n855_), .B(_abc_73687_new_n854_), .Y(\o[120] ));
AND2X2 AND2X2_850 ( .A(u2__abc_52155_new_n3716_), .B(sqrto_111_), .Y(u2__abc_52155_new_n3717_));
AND2X2 AND2X2_8500 ( .A(u2__abc_52155_new_n17787_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17788_));
AND2X2 AND2X2_8501 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_209_), .Y(u2__abc_52155_new_n17790_));
AND2X2 AND2X2_8502 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_207_), .Y(u2__abc_52155_new_n17791_));
AND2X2 AND2X2_8503 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_65_), .Y(u2__abc_52155_new_n17792_));
AND2X2 AND2X2_8504 ( .A(u2__abc_52155_new_n17793_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17794_));
AND2X2 AND2X2_8505 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_210_), .Y(u2__abc_52155_new_n17796_));
AND2X2 AND2X2_8506 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_208_), .Y(u2__abc_52155_new_n17797_));
AND2X2 AND2X2_8507 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_66_), .Y(u2__abc_52155_new_n17798_));
AND2X2 AND2X2_8508 ( .A(u2__abc_52155_new_n17799_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17800_));
AND2X2 AND2X2_8509 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_211_), .Y(u2__abc_52155_new_n17802_));
AND2X2 AND2X2_851 ( .A(u2__abc_52155_new_n3715_), .B(u2__abc_52155_new_n3718_), .Y(u2__abc_52155_new_n3719_));
AND2X2 AND2X2_8510 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_67_), .Y(u2__abc_52155_new_n17803_));
AND2X2 AND2X2_8511 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_209_), .Y(u2__abc_52155_new_n17804_));
AND2X2 AND2X2_8512 ( .A(u2__abc_52155_new_n17805_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17806_));
AND2X2 AND2X2_8513 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_212_), .Y(u2__abc_52155_new_n17808_));
AND2X2 AND2X2_8514 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_210_), .Y(u2__abc_52155_new_n17809_));
AND2X2 AND2X2_8515 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_68_), .Y(u2__abc_52155_new_n17810_));
AND2X2 AND2X2_8516 ( .A(u2__abc_52155_new_n17811_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17812_));
AND2X2 AND2X2_8517 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_213_), .Y(u2__abc_52155_new_n17814_));
AND2X2 AND2X2_8518 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_211_), .Y(u2__abc_52155_new_n17815_));
AND2X2 AND2X2_8519 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_69_), .Y(u2__abc_52155_new_n17816_));
AND2X2 AND2X2_852 ( .A(u2__abc_52155_new_n3712_), .B(u2__abc_52155_new_n3719_), .Y(u2__abc_52155_new_n3720_));
AND2X2 AND2X2_8520 ( .A(u2__abc_52155_new_n17817_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17818_));
AND2X2 AND2X2_8521 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_214_), .Y(u2__abc_52155_new_n17820_));
AND2X2 AND2X2_8522 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_212_), .Y(u2__abc_52155_new_n17821_));
AND2X2 AND2X2_8523 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_70_), .Y(u2__abc_52155_new_n17822_));
AND2X2 AND2X2_8524 ( .A(u2__abc_52155_new_n17823_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17824_));
AND2X2 AND2X2_8525 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_215_), .Y(u2__abc_52155_new_n17826_));
AND2X2 AND2X2_8526 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_213_), .Y(u2__abc_52155_new_n17827_));
AND2X2 AND2X2_8527 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_71_), .Y(u2__abc_52155_new_n17828_));
AND2X2 AND2X2_8528 ( .A(u2__abc_52155_new_n17829_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17830_));
AND2X2 AND2X2_8529 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_216_), .Y(u2__abc_52155_new_n17832_));
AND2X2 AND2X2_853 ( .A(u2__abc_52155_new_n3721_), .B(u2_remHi_112_), .Y(u2__abc_52155_new_n3722_));
AND2X2 AND2X2_8530 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_214_), .Y(u2__abc_52155_new_n17833_));
AND2X2 AND2X2_8531 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_72_), .Y(u2__abc_52155_new_n17834_));
AND2X2 AND2X2_8532 ( .A(u2__abc_52155_new_n17835_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17836_));
AND2X2 AND2X2_8533 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_217_), .Y(u2__abc_52155_new_n17838_));
AND2X2 AND2X2_8534 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_73_), .Y(u2__abc_52155_new_n17839_));
AND2X2 AND2X2_8535 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_215_), .Y(u2__abc_52155_new_n17840_));
AND2X2 AND2X2_8536 ( .A(u2__abc_52155_new_n17841_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17842_));
AND2X2 AND2X2_8537 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_218_), .Y(u2__abc_52155_new_n17844_));
AND2X2 AND2X2_8538 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_74_), .Y(u2__abc_52155_new_n17845_));
AND2X2 AND2X2_8539 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_216_), .Y(u2__abc_52155_new_n17846_));
AND2X2 AND2X2_854 ( .A(u2__abc_52155_new_n3724_), .B(sqrto_112_), .Y(u2__abc_52155_new_n3725_));
AND2X2 AND2X2_8540 ( .A(u2__abc_52155_new_n17847_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17848_));
AND2X2 AND2X2_8541 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_219_), .Y(u2__abc_52155_new_n17850_));
AND2X2 AND2X2_8542 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_217_), .Y(u2__abc_52155_new_n17851_));
AND2X2 AND2X2_8543 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_75_), .Y(u2__abc_52155_new_n17852_));
AND2X2 AND2X2_8544 ( .A(u2__abc_52155_new_n17853_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17854_));
AND2X2 AND2X2_8545 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_220_), .Y(u2__abc_52155_new_n17856_));
AND2X2 AND2X2_8546 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_218_), .Y(u2__abc_52155_new_n17857_));
AND2X2 AND2X2_8547 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_76_), .Y(u2__abc_52155_new_n17858_));
AND2X2 AND2X2_8548 ( .A(u2__abc_52155_new_n17859_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17860_));
AND2X2 AND2X2_8549 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_221_), .Y(u2__abc_52155_new_n17862_));
AND2X2 AND2X2_855 ( .A(u2__abc_52155_new_n3723_), .B(u2__abc_52155_new_n3726_), .Y(u2__abc_52155_new_n3727_));
AND2X2 AND2X2_8550 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_219_), .Y(u2__abc_52155_new_n17863_));
AND2X2 AND2X2_8551 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_77_), .Y(u2__abc_52155_new_n17864_));
AND2X2 AND2X2_8552 ( .A(u2__abc_52155_new_n17865_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17866_));
AND2X2 AND2X2_8553 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_222_), .Y(u2__abc_52155_new_n17868_));
AND2X2 AND2X2_8554 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_220_), .Y(u2__abc_52155_new_n17869_));
AND2X2 AND2X2_8555 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_78_), .Y(u2__abc_52155_new_n17870_));
AND2X2 AND2X2_8556 ( .A(u2__abc_52155_new_n17871_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17872_));
AND2X2 AND2X2_8557 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_223_), .Y(u2__abc_52155_new_n17874_));
AND2X2 AND2X2_8558 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_79_), .Y(u2__abc_52155_new_n17875_));
AND2X2 AND2X2_8559 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_221_), .Y(u2__abc_52155_new_n17876_));
AND2X2 AND2X2_856 ( .A(u2__abc_52155_new_n3728_), .B(u2_remHi_113_), .Y(u2__abc_52155_new_n3729_));
AND2X2 AND2X2_8560 ( .A(u2__abc_52155_new_n17877_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17878_));
AND2X2 AND2X2_8561 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_224_), .Y(u2__abc_52155_new_n17880_));
AND2X2 AND2X2_8562 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_222_), .Y(u2__abc_52155_new_n17881_));
AND2X2 AND2X2_8563 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_80_), .Y(u2__abc_52155_new_n17882_));
AND2X2 AND2X2_8564 ( .A(u2__abc_52155_new_n17883_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17884_));
AND2X2 AND2X2_8565 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_225_), .Y(u2__abc_52155_new_n17886_));
AND2X2 AND2X2_8566 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_223_), .Y(u2__abc_52155_new_n17887_));
AND2X2 AND2X2_8567 ( .A(u2__abc_52155_new_n17888_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17889_));
AND2X2 AND2X2_8568 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_225_), .Y(u2__abc_52155_new_n17890_));
AND2X2 AND2X2_8569 ( .A(u2__abc_52155_new_n2964_), .B(fracta1_81_), .Y(u2__abc_52155_new_n17891_));
AND2X2 AND2X2_857 ( .A(u2__abc_52155_new_n3731_), .B(sqrto_113_), .Y(u2__abc_52155_new_n3732_));
AND2X2 AND2X2_8570 ( .A(u2__abc_52155_new_n17892_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17893_));
AND2X2 AND2X2_8571 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_226_), .Y(u2__abc_52155_new_n17895_));
AND2X2 AND2X2_8572 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_224_), .Y(u2__abc_52155_new_n17896_));
AND2X2 AND2X2_8573 ( .A(u2__abc_52155_new_n17897_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17898_));
AND2X2 AND2X2_8574 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_226_), .Y(u2__abc_52155_new_n17899_));
AND2X2 AND2X2_8575 ( .A(u2__abc_52155_new_n2964_), .B(fracta1_82_), .Y(u2__abc_52155_new_n17900_));
AND2X2 AND2X2_8576 ( .A(u2__abc_52155_new_n17901_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17902_));
AND2X2 AND2X2_8577 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_227_), .Y(u2__abc_52155_new_n17904_));
AND2X2 AND2X2_8578 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_225_), .Y(u2__abc_52155_new_n17905_));
AND2X2 AND2X2_8579 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_83_), .Y(u2__abc_52155_new_n17906_));
AND2X2 AND2X2_858 ( .A(u2__abc_52155_new_n3730_), .B(u2__abc_52155_new_n3733_), .Y(u2__abc_52155_new_n3734_));
AND2X2 AND2X2_8580 ( .A(u2__abc_52155_new_n17907_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17908_));
AND2X2 AND2X2_8581 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_228_), .Y(u2__abc_52155_new_n17910_));
AND2X2 AND2X2_8582 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_226_), .Y(u2__abc_52155_new_n17911_));
AND2X2 AND2X2_8583 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_84_), .Y(u2__abc_52155_new_n17912_));
AND2X2 AND2X2_8584 ( .A(u2__abc_52155_new_n17913_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17914_));
AND2X2 AND2X2_8585 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_229_), .Y(u2__abc_52155_new_n17916_));
AND2X2 AND2X2_8586 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_227_), .Y(u2__abc_52155_new_n17917_));
AND2X2 AND2X2_8587 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_85_), .Y(u2__abc_52155_new_n17918_));
AND2X2 AND2X2_8588 ( .A(u2__abc_52155_new_n17919_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17920_));
AND2X2 AND2X2_8589 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_230_), .Y(u2__abc_52155_new_n17922_));
AND2X2 AND2X2_859 ( .A(u2__abc_52155_new_n3727_), .B(u2__abc_52155_new_n3734_), .Y(u2__abc_52155_new_n3735_));
AND2X2 AND2X2_8590 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_228_), .Y(u2__abc_52155_new_n17923_));
AND2X2 AND2X2_8591 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_86_), .Y(u2__abc_52155_new_n17924_));
AND2X2 AND2X2_8592 ( .A(u2__abc_52155_new_n17925_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17926_));
AND2X2 AND2X2_8593 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_231_), .Y(u2__abc_52155_new_n17928_));
AND2X2 AND2X2_8594 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_229_), .Y(u2__abc_52155_new_n17929_));
AND2X2 AND2X2_8595 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_87_), .Y(u2__abc_52155_new_n17930_));
AND2X2 AND2X2_8596 ( .A(u2__abc_52155_new_n17931_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17932_));
AND2X2 AND2X2_8597 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_232_), .Y(u2__abc_52155_new_n17934_));
AND2X2 AND2X2_8598 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_230_), .Y(u2__abc_52155_new_n17935_));
AND2X2 AND2X2_8599 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_88_), .Y(u2__abc_52155_new_n17936_));
AND2X2 AND2X2_86 ( .A(_abc_73687_new_n858_), .B(_abc_73687_new_n857_), .Y(\o[121] ));
AND2X2 AND2X2_860 ( .A(u2__abc_52155_new_n3720_), .B(u2__abc_52155_new_n3735_), .Y(u2__abc_52155_new_n3736_));
AND2X2 AND2X2_8600 ( .A(u2__abc_52155_new_n17937_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17938_));
AND2X2 AND2X2_8601 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_233_), .Y(u2__abc_52155_new_n17940_));
AND2X2 AND2X2_8602 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_231_), .Y(u2__abc_52155_new_n17941_));
AND2X2 AND2X2_8603 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_89_), .Y(u2__abc_52155_new_n17942_));
AND2X2 AND2X2_8604 ( .A(u2__abc_52155_new_n17943_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17944_));
AND2X2 AND2X2_8605 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_234_), .Y(u2__abc_52155_new_n17946_));
AND2X2 AND2X2_8606 ( .A(u2__abc_52155_new_n17085_), .B(fracta1_90_), .Y(u2__abc_52155_new_n17947_));
AND2X2 AND2X2_8607 ( .A(u2__abc_52155_new_n2982_), .B(u2_remLo_232_), .Y(u2__abc_52155_new_n17948_));
AND2X2 AND2X2_8608 ( .A(u2__abc_52155_new_n16683_), .B(u2__abc_52155_new_n17948_), .Y(u2__abc_52155_new_n17949_));
AND2X2 AND2X2_8609 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_235_), .Y(u2__abc_52155_new_n17952_));
AND2X2 AND2X2_861 ( .A(u2__abc_52155_new_n3737_), .B(u2_remHi_116_), .Y(u2__abc_52155_new_n3738_));
AND2X2 AND2X2_8610 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_233_), .Y(u2__abc_52155_new_n17953_));
AND2X2 AND2X2_8611 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_91_), .Y(u2__abc_52155_new_n17954_));
AND2X2 AND2X2_8612 ( .A(u2__abc_52155_new_n17955_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17956_));
AND2X2 AND2X2_8613 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_236_), .Y(u2__abc_52155_new_n17958_));
AND2X2 AND2X2_8614 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_234_), .Y(u2__abc_52155_new_n17959_));
AND2X2 AND2X2_8615 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_92_), .Y(u2__abc_52155_new_n17960_));
AND2X2 AND2X2_8616 ( .A(u2__abc_52155_new_n17961_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17962_));
AND2X2 AND2X2_8617 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_237_), .Y(u2__abc_52155_new_n17964_));
AND2X2 AND2X2_8618 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_235_), .Y(u2__abc_52155_new_n17965_));
AND2X2 AND2X2_8619 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_93_), .Y(u2__abc_52155_new_n17966_));
AND2X2 AND2X2_862 ( .A(u2__abc_52155_new_n3740_), .B(sqrto_116_), .Y(u2__abc_52155_new_n3741_));
AND2X2 AND2X2_8620 ( .A(u2__abc_52155_new_n17967_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17968_));
AND2X2 AND2X2_8621 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_238_), .Y(u2__abc_52155_new_n17970_));
AND2X2 AND2X2_8622 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_236_), .Y(u2__abc_52155_new_n17971_));
AND2X2 AND2X2_8623 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_94_), .Y(u2__abc_52155_new_n17972_));
AND2X2 AND2X2_8624 ( .A(u2__abc_52155_new_n17973_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17974_));
AND2X2 AND2X2_8625 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_239_), .Y(u2__abc_52155_new_n17976_));
AND2X2 AND2X2_8626 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_95_), .Y(u2__abc_52155_new_n17977_));
AND2X2 AND2X2_8627 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_237_), .Y(u2__abc_52155_new_n17978_));
AND2X2 AND2X2_8628 ( .A(u2__abc_52155_new_n17979_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17980_));
AND2X2 AND2X2_8629 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_240_), .Y(u2__abc_52155_new_n17982_));
AND2X2 AND2X2_863 ( .A(u2__abc_52155_new_n3739_), .B(u2__abc_52155_new_n3742_), .Y(u2__abc_52155_new_n3743_));
AND2X2 AND2X2_8630 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_238_), .Y(u2__abc_52155_new_n17983_));
AND2X2 AND2X2_8631 ( .A(u2__abc_52155_new_n17984_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17985_));
AND2X2 AND2X2_8632 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_240_), .Y(u2__abc_52155_new_n17986_));
AND2X2 AND2X2_8633 ( .A(u2__abc_52155_new_n2964_), .B(fracta1_96_), .Y(u2__abc_52155_new_n17987_));
AND2X2 AND2X2_8634 ( .A(u2__abc_52155_new_n17988_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n17989_));
AND2X2 AND2X2_8635 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_241_), .Y(u2__abc_52155_new_n17991_));
AND2X2 AND2X2_8636 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_239_), .Y(u2__abc_52155_new_n17992_));
AND2X2 AND2X2_8637 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_97_), .Y(u2__abc_52155_new_n17993_));
AND2X2 AND2X2_8638 ( .A(u2__abc_52155_new_n17994_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n17995_));
AND2X2 AND2X2_8639 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_242_), .Y(u2__abc_52155_new_n17997_));
AND2X2 AND2X2_864 ( .A(u2__abc_52155_new_n3744_), .B(u2_remHi_117_), .Y(u2__abc_52155_new_n3745_));
AND2X2 AND2X2_8640 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_240_), .Y(u2__abc_52155_new_n17998_));
AND2X2 AND2X2_8641 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_98_), .Y(u2__abc_52155_new_n17999_));
AND2X2 AND2X2_8642 ( .A(u2__abc_52155_new_n18000_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18001_));
AND2X2 AND2X2_8643 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_243_), .Y(u2__abc_52155_new_n18003_));
AND2X2 AND2X2_8644 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_99_), .Y(u2__abc_52155_new_n18004_));
AND2X2 AND2X2_8645 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_241_), .Y(u2__abc_52155_new_n18005_));
AND2X2 AND2X2_8646 ( .A(u2__abc_52155_new_n18006_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18007_));
AND2X2 AND2X2_8647 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_244_), .Y(u2__abc_52155_new_n18009_));
AND2X2 AND2X2_8648 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_242_), .Y(u2__abc_52155_new_n18010_));
AND2X2 AND2X2_8649 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_100_), .Y(u2__abc_52155_new_n18011_));
AND2X2 AND2X2_865 ( .A(u2__abc_52155_new_n3747_), .B(sqrto_117_), .Y(u2__abc_52155_new_n3748_));
AND2X2 AND2X2_8650 ( .A(u2__abc_52155_new_n18012_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18013_));
AND2X2 AND2X2_8651 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_245_), .Y(u2__abc_52155_new_n18015_));
AND2X2 AND2X2_8652 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_243_), .Y(u2__abc_52155_new_n18016_));
AND2X2 AND2X2_8653 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_101_), .Y(u2__abc_52155_new_n18017_));
AND2X2 AND2X2_8654 ( .A(u2__abc_52155_new_n18018_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18019_));
AND2X2 AND2X2_8655 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_246_), .Y(u2__abc_52155_new_n18021_));
AND2X2 AND2X2_8656 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_244_), .Y(u2__abc_52155_new_n18022_));
AND2X2 AND2X2_8657 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_102_), .Y(u2__abc_52155_new_n18023_));
AND2X2 AND2X2_8658 ( .A(u2__abc_52155_new_n18024_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18025_));
AND2X2 AND2X2_8659 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_247_), .Y(u2__abc_52155_new_n18027_));
AND2X2 AND2X2_866 ( .A(u2__abc_52155_new_n3746_), .B(u2__abc_52155_new_n3749_), .Y(u2__abc_52155_new_n3750_));
AND2X2 AND2X2_8660 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_245_), .Y(u2__abc_52155_new_n18028_));
AND2X2 AND2X2_8661 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_103_), .Y(u2__abc_52155_new_n18029_));
AND2X2 AND2X2_8662 ( .A(u2__abc_52155_new_n18030_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18031_));
AND2X2 AND2X2_8663 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_248_), .Y(u2__abc_52155_new_n18033_));
AND2X2 AND2X2_8664 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_246_), .Y(u2__abc_52155_new_n18034_));
AND2X2 AND2X2_8665 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_104_), .Y(u2__abc_52155_new_n18035_));
AND2X2 AND2X2_8666 ( .A(u2__abc_52155_new_n18036_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18037_));
AND2X2 AND2X2_8667 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_249_), .Y(u2__abc_52155_new_n18039_));
AND2X2 AND2X2_8668 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_105_), .Y(u2__abc_52155_new_n18040_));
AND2X2 AND2X2_8669 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_247_), .Y(u2__abc_52155_new_n18041_));
AND2X2 AND2X2_867 ( .A(u2__abc_52155_new_n3743_), .B(u2__abc_52155_new_n3750_), .Y(u2__abc_52155_new_n3751_));
AND2X2 AND2X2_8670 ( .A(u2__abc_52155_new_n18042_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18043_));
AND2X2 AND2X2_8671 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_250_), .Y(u2__abc_52155_new_n18045_));
AND2X2 AND2X2_8672 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_106_), .Y(u2__abc_52155_new_n18046_));
AND2X2 AND2X2_8673 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_248_), .Y(u2__abc_52155_new_n18047_));
AND2X2 AND2X2_8674 ( .A(u2__abc_52155_new_n18048_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18049_));
AND2X2 AND2X2_8675 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_251_), .Y(u2__abc_52155_new_n18051_));
AND2X2 AND2X2_8676 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_249_), .Y(u2__abc_52155_new_n18052_));
AND2X2 AND2X2_8677 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_107_), .Y(u2__abc_52155_new_n18053_));
AND2X2 AND2X2_8678 ( .A(u2__abc_52155_new_n18054_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18055_));
AND2X2 AND2X2_8679 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_252_), .Y(u2__abc_52155_new_n18057_));
AND2X2 AND2X2_868 ( .A(u2__abc_52155_new_n3752_), .B(u2_remHi_115_), .Y(u2__abc_52155_new_n3753_));
AND2X2 AND2X2_8680 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_250_), .Y(u2__abc_52155_new_n18058_));
AND2X2 AND2X2_8681 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_108_), .Y(u2__abc_52155_new_n18059_));
AND2X2 AND2X2_8682 ( .A(u2__abc_52155_new_n18060_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18061_));
AND2X2 AND2X2_8683 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_253_), .Y(u2__abc_52155_new_n18063_));
AND2X2 AND2X2_8684 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_109_), .Y(u2__abc_52155_new_n18064_));
AND2X2 AND2X2_8685 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_251_), .Y(u2__abc_52155_new_n18065_));
AND2X2 AND2X2_8686 ( .A(u2__abc_52155_new_n18066_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18067_));
AND2X2 AND2X2_8687 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_254_), .Y(u2__abc_52155_new_n18069_));
AND2X2 AND2X2_8688 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_252_), .Y(u2__abc_52155_new_n18070_));
AND2X2 AND2X2_8689 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_110_), .Y(u2__abc_52155_new_n18071_));
AND2X2 AND2X2_869 ( .A(u2__abc_52155_new_n3755_), .B(sqrto_115_), .Y(u2__abc_52155_new_n3756_));
AND2X2 AND2X2_8690 ( .A(u2__abc_52155_new_n18072_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18073_));
AND2X2 AND2X2_8691 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_255_), .Y(u2__abc_52155_new_n18075_));
AND2X2 AND2X2_8692 ( .A(u2__abc_52155_new_n2963_), .B(fracta1_111_), .Y(u2__abc_52155_new_n18076_));
AND2X2 AND2X2_8693 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_253_), .Y(u2__abc_52155_new_n18077_));
AND2X2 AND2X2_8694 ( .A(u2__abc_52155_new_n18078_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18079_));
AND2X2 AND2X2_8695 ( .A(u2__abc_52155_new_n16680_), .B(u2_remLo_256_), .Y(u2__abc_52155_new_n18081_));
AND2X2 AND2X2_8696 ( .A(u2__abc_52155_new_n17085_), .B(fracta1_112_), .Y(u2__abc_52155_new_n18082_));
AND2X2 AND2X2_8697 ( .A(u2__abc_52155_new_n2982_), .B(u2_remLo_254_), .Y(u2__abc_52155_new_n18083_));
AND2X2 AND2X2_8698 ( .A(u2__abc_52155_new_n16683_), .B(u2__abc_52155_new_n18083_), .Y(u2__abc_52155_new_n18084_));
AND2X2 AND2X2_8699 ( .A(u2__abc_52155_new_n16678_), .B(u2_remLo_257_), .Y(u2__abc_52155_new_n18087_));
AND2X2 AND2X2_87 ( .A(_abc_73687_new_n861_), .B(_abc_73687_new_n860_), .Y(\o[122] ));
AND2X2 AND2X2_870 ( .A(u2__abc_52155_new_n3754_), .B(u2__abc_52155_new_n3757_), .Y(u2__abc_52155_new_n3758_));
AND2X2 AND2X2_8700 ( .A(u2__abc_52155_new_n16683_), .B(u2_remLo_255_), .Y(u2__abc_52155_new_n18088_));
AND2X2 AND2X2_8701 ( .A(u2__abc_52155_new_n18089_), .B(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n18090_));
AND2X2 AND2X2_8702 ( .A(u2__abc_52155_new_n3001_), .B(u2_remLo_257_), .Y(u2__abc_52155_new_n18091_));
AND2X2 AND2X2_8703 ( .A(u2__abc_52155_new_n2964_), .B(fracta1_113_), .Y(u2__abc_52155_new_n18092_));
AND2X2 AND2X2_8704 ( .A(u2__abc_52155_new_n18093_), .B(u2__abc_52155_new_n2962_), .Y(u2__abc_52155_new_n18094_));
AND2X2 AND2X2_8705 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_258_), .Y(u2__abc_52155_new_n18096_));
AND2X2 AND2X2_8706 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_256_), .Y(u2__abc_52155_new_n18097_));
AND2X2 AND2X2_8707 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18097_), .Y(u2__abc_52155_new_n18098_));
AND2X2 AND2X2_8708 ( .A(u2__abc_52155_new_n18099_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__258_));
AND2X2 AND2X2_8709 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_259_), .Y(u2__abc_52155_new_n18101_));
AND2X2 AND2X2_871 ( .A(u2__abc_52155_new_n3759_), .B(u2_remHi_114_), .Y(u2__abc_52155_new_n3760_));
AND2X2 AND2X2_8710 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_257_), .Y(u2__abc_52155_new_n18102_));
AND2X2 AND2X2_8711 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18102_), .Y(u2__abc_52155_new_n18103_));
AND2X2 AND2X2_8712 ( .A(u2__abc_52155_new_n18104_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__259_));
AND2X2 AND2X2_8713 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_260_), .Y(u2__abc_52155_new_n18106_));
AND2X2 AND2X2_8714 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_258_), .Y(u2__abc_52155_new_n18107_));
AND2X2 AND2X2_8715 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18107_), .Y(u2__abc_52155_new_n18108_));
AND2X2 AND2X2_8716 ( .A(u2__abc_52155_new_n18109_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__260_));
AND2X2 AND2X2_8717 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_261_), .Y(u2__abc_52155_new_n18111_));
AND2X2 AND2X2_8718 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_259_), .Y(u2__abc_52155_new_n18112_));
AND2X2 AND2X2_8719 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18112_), .Y(u2__abc_52155_new_n18113_));
AND2X2 AND2X2_872 ( .A(u2__abc_52155_new_n3762_), .B(sqrto_114_), .Y(u2__abc_52155_new_n3763_));
AND2X2 AND2X2_8720 ( .A(u2__abc_52155_new_n18114_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__261_));
AND2X2 AND2X2_8721 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_262_), .Y(u2__abc_52155_new_n18116_));
AND2X2 AND2X2_8722 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_260_), .Y(u2__abc_52155_new_n18117_));
AND2X2 AND2X2_8723 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18117_), .Y(u2__abc_52155_new_n18118_));
AND2X2 AND2X2_8724 ( .A(u2__abc_52155_new_n18119_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__262_));
AND2X2 AND2X2_8725 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_263_), .Y(u2__abc_52155_new_n18121_));
AND2X2 AND2X2_8726 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_261_), .Y(u2__abc_52155_new_n18122_));
AND2X2 AND2X2_8727 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18122_), .Y(u2__abc_52155_new_n18123_));
AND2X2 AND2X2_8728 ( .A(u2__abc_52155_new_n18124_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__263_));
AND2X2 AND2X2_8729 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_264_), .Y(u2__abc_52155_new_n18126_));
AND2X2 AND2X2_873 ( .A(u2__abc_52155_new_n3761_), .B(u2__abc_52155_new_n3764_), .Y(u2__abc_52155_new_n3765_));
AND2X2 AND2X2_8730 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_262_), .Y(u2__abc_52155_new_n18127_));
AND2X2 AND2X2_8731 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18127_), .Y(u2__abc_52155_new_n18128_));
AND2X2 AND2X2_8732 ( .A(u2__abc_52155_new_n18129_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__264_));
AND2X2 AND2X2_8733 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_265_), .Y(u2__abc_52155_new_n18131_));
AND2X2 AND2X2_8734 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_263_), .Y(u2__abc_52155_new_n18132_));
AND2X2 AND2X2_8735 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18132_), .Y(u2__abc_52155_new_n18133_));
AND2X2 AND2X2_8736 ( .A(u2__abc_52155_new_n18134_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__265_));
AND2X2 AND2X2_8737 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_266_), .Y(u2__abc_52155_new_n18136_));
AND2X2 AND2X2_8738 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_264_), .Y(u2__abc_52155_new_n18137_));
AND2X2 AND2X2_8739 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18137_), .Y(u2__abc_52155_new_n18138_));
AND2X2 AND2X2_874 ( .A(u2__abc_52155_new_n3758_), .B(u2__abc_52155_new_n3765_), .Y(u2__abc_52155_new_n3766_));
AND2X2 AND2X2_8740 ( .A(u2__abc_52155_new_n18139_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__266_));
AND2X2 AND2X2_8741 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_267_), .Y(u2__abc_52155_new_n18141_));
AND2X2 AND2X2_8742 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_265_), .Y(u2__abc_52155_new_n18142_));
AND2X2 AND2X2_8743 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18142_), .Y(u2__abc_52155_new_n18143_));
AND2X2 AND2X2_8744 ( .A(u2__abc_52155_new_n18144_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__267_));
AND2X2 AND2X2_8745 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_268_), .Y(u2__abc_52155_new_n18146_));
AND2X2 AND2X2_8746 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_266_), .Y(u2__abc_52155_new_n18147_));
AND2X2 AND2X2_8747 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18147_), .Y(u2__abc_52155_new_n18148_));
AND2X2 AND2X2_8748 ( .A(u2__abc_52155_new_n18149_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__268_));
AND2X2 AND2X2_8749 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_269_), .Y(u2__abc_52155_new_n18151_));
AND2X2 AND2X2_875 ( .A(u2__abc_52155_new_n3751_), .B(u2__abc_52155_new_n3766_), .Y(u2__abc_52155_new_n3767_));
AND2X2 AND2X2_8750 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_267_), .Y(u2__abc_52155_new_n18152_));
AND2X2 AND2X2_8751 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18152_), .Y(u2__abc_52155_new_n18153_));
AND2X2 AND2X2_8752 ( .A(u2__abc_52155_new_n18154_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__269_));
AND2X2 AND2X2_8753 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_270_), .Y(u2__abc_52155_new_n18156_));
AND2X2 AND2X2_8754 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_268_), .Y(u2__abc_52155_new_n18157_));
AND2X2 AND2X2_8755 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18157_), .Y(u2__abc_52155_new_n18158_));
AND2X2 AND2X2_8756 ( .A(u2__abc_52155_new_n18159_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__270_));
AND2X2 AND2X2_8757 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_271_), .Y(u2__abc_52155_new_n18161_));
AND2X2 AND2X2_8758 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_269_), .Y(u2__abc_52155_new_n18162_));
AND2X2 AND2X2_8759 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18162_), .Y(u2__abc_52155_new_n18163_));
AND2X2 AND2X2_876 ( .A(u2__abc_52155_new_n3736_), .B(u2__abc_52155_new_n3767_), .Y(u2__abc_52155_new_n3768_));
AND2X2 AND2X2_8760 ( .A(u2__abc_52155_new_n18164_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__271_));
AND2X2 AND2X2_8761 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_272_), .Y(u2__abc_52155_new_n18166_));
AND2X2 AND2X2_8762 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_270_), .Y(u2__abc_52155_new_n18167_));
AND2X2 AND2X2_8763 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18167_), .Y(u2__abc_52155_new_n18168_));
AND2X2 AND2X2_8764 ( .A(u2__abc_52155_new_n18169_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__272_));
AND2X2 AND2X2_8765 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_273_), .Y(u2__abc_52155_new_n18171_));
AND2X2 AND2X2_8766 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_271_), .Y(u2__abc_52155_new_n18172_));
AND2X2 AND2X2_8767 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18172_), .Y(u2__abc_52155_new_n18173_));
AND2X2 AND2X2_8768 ( .A(u2__abc_52155_new_n18174_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__273_));
AND2X2 AND2X2_8769 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_274_), .Y(u2__abc_52155_new_n18176_));
AND2X2 AND2X2_877 ( .A(u2__abc_52155_new_n3705_), .B(u2__abc_52155_new_n3768_), .Y(u2__abc_52155_new_n3769_));
AND2X2 AND2X2_8770 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_272_), .Y(u2__abc_52155_new_n18177_));
AND2X2 AND2X2_8771 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18177_), .Y(u2__abc_52155_new_n18178_));
AND2X2 AND2X2_8772 ( .A(u2__abc_52155_new_n18179_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__274_));
AND2X2 AND2X2_8773 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_275_), .Y(u2__abc_52155_new_n18181_));
AND2X2 AND2X2_8774 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_273_), .Y(u2__abc_52155_new_n18182_));
AND2X2 AND2X2_8775 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18182_), .Y(u2__abc_52155_new_n18183_));
AND2X2 AND2X2_8776 ( .A(u2__abc_52155_new_n18184_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__275_));
AND2X2 AND2X2_8777 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_276_), .Y(u2__abc_52155_new_n18186_));
AND2X2 AND2X2_8778 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_274_), .Y(u2__abc_52155_new_n18187_));
AND2X2 AND2X2_8779 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18187_), .Y(u2__abc_52155_new_n18188_));
AND2X2 AND2X2_878 ( .A(u2__abc_52155_new_n3770_), .B(u2_remHi_104_), .Y(u2__abc_52155_new_n3771_));
AND2X2 AND2X2_8780 ( .A(u2__abc_52155_new_n18189_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__276_));
AND2X2 AND2X2_8781 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_277_), .Y(u2__abc_52155_new_n18191_));
AND2X2 AND2X2_8782 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_275_), .Y(u2__abc_52155_new_n18192_));
AND2X2 AND2X2_8783 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18192_), .Y(u2__abc_52155_new_n18193_));
AND2X2 AND2X2_8784 ( .A(u2__abc_52155_new_n18194_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__277_));
AND2X2 AND2X2_8785 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_278_), .Y(u2__abc_52155_new_n18196_));
AND2X2 AND2X2_8786 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_276_), .Y(u2__abc_52155_new_n18197_));
AND2X2 AND2X2_8787 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18197_), .Y(u2__abc_52155_new_n18198_));
AND2X2 AND2X2_8788 ( .A(u2__abc_52155_new_n18199_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__278_));
AND2X2 AND2X2_8789 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_279_), .Y(u2__abc_52155_new_n18201_));
AND2X2 AND2X2_879 ( .A(u2__abc_52155_new_n3773_), .B(sqrto_104_), .Y(u2__abc_52155_new_n3774_));
AND2X2 AND2X2_8790 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_277_), .Y(u2__abc_52155_new_n18202_));
AND2X2 AND2X2_8791 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18202_), .Y(u2__abc_52155_new_n18203_));
AND2X2 AND2X2_8792 ( .A(u2__abc_52155_new_n18204_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__279_));
AND2X2 AND2X2_8793 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_280_), .Y(u2__abc_52155_new_n18206_));
AND2X2 AND2X2_8794 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_278_), .Y(u2__abc_52155_new_n18207_));
AND2X2 AND2X2_8795 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18207_), .Y(u2__abc_52155_new_n18208_));
AND2X2 AND2X2_8796 ( .A(u2__abc_52155_new_n18209_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__280_));
AND2X2 AND2X2_8797 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_281_), .Y(u2__abc_52155_new_n18211_));
AND2X2 AND2X2_8798 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_279_), .Y(u2__abc_52155_new_n18212_));
AND2X2 AND2X2_8799 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18212_), .Y(u2__abc_52155_new_n18213_));
AND2X2 AND2X2_88 ( .A(_abc_73687_new_n864_), .B(_abc_73687_new_n863_), .Y(\o[123] ));
AND2X2 AND2X2_880 ( .A(u2__abc_52155_new_n3772_), .B(u2__abc_52155_new_n3775_), .Y(u2__abc_52155_new_n3776_));
AND2X2 AND2X2_8800 ( .A(u2__abc_52155_new_n18214_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__281_));
AND2X2 AND2X2_8801 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_282_), .Y(u2__abc_52155_new_n18216_));
AND2X2 AND2X2_8802 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_280_), .Y(u2__abc_52155_new_n18217_));
AND2X2 AND2X2_8803 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18217_), .Y(u2__abc_52155_new_n18218_));
AND2X2 AND2X2_8804 ( .A(u2__abc_52155_new_n18219_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__282_));
AND2X2 AND2X2_8805 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_283_), .Y(u2__abc_52155_new_n18221_));
AND2X2 AND2X2_8806 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_281_), .Y(u2__abc_52155_new_n18222_));
AND2X2 AND2X2_8807 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18222_), .Y(u2__abc_52155_new_n18223_));
AND2X2 AND2X2_8808 ( .A(u2__abc_52155_new_n18224_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__283_));
AND2X2 AND2X2_8809 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_284_), .Y(u2__abc_52155_new_n18226_));
AND2X2 AND2X2_881 ( .A(u2__abc_52155_new_n3777_), .B(u2_remHi_105_), .Y(u2__abc_52155_new_n3778_));
AND2X2 AND2X2_8810 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_282_), .Y(u2__abc_52155_new_n18227_));
AND2X2 AND2X2_8811 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18227_), .Y(u2__abc_52155_new_n18228_));
AND2X2 AND2X2_8812 ( .A(u2__abc_52155_new_n18229_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__284_));
AND2X2 AND2X2_8813 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_285_), .Y(u2__abc_52155_new_n18231_));
AND2X2 AND2X2_8814 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_283_), .Y(u2__abc_52155_new_n18232_));
AND2X2 AND2X2_8815 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18232_), .Y(u2__abc_52155_new_n18233_));
AND2X2 AND2X2_8816 ( .A(u2__abc_52155_new_n18234_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__285_));
AND2X2 AND2X2_8817 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_286_), .Y(u2__abc_52155_new_n18236_));
AND2X2 AND2X2_8818 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_284_), .Y(u2__abc_52155_new_n18237_));
AND2X2 AND2X2_8819 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18237_), .Y(u2__abc_52155_new_n18238_));
AND2X2 AND2X2_882 ( .A(u2__abc_52155_new_n3780_), .B(sqrto_105_), .Y(u2__abc_52155_new_n3781_));
AND2X2 AND2X2_8820 ( .A(u2__abc_52155_new_n18239_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__286_));
AND2X2 AND2X2_8821 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_287_), .Y(u2__abc_52155_new_n18241_));
AND2X2 AND2X2_8822 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_285_), .Y(u2__abc_52155_new_n18242_));
AND2X2 AND2X2_8823 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18242_), .Y(u2__abc_52155_new_n18243_));
AND2X2 AND2X2_8824 ( .A(u2__abc_52155_new_n18244_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__287_));
AND2X2 AND2X2_8825 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_288_), .Y(u2__abc_52155_new_n18246_));
AND2X2 AND2X2_8826 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_286_), .Y(u2__abc_52155_new_n18247_));
AND2X2 AND2X2_8827 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18247_), .Y(u2__abc_52155_new_n18248_));
AND2X2 AND2X2_8828 ( .A(u2__abc_52155_new_n18249_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__288_));
AND2X2 AND2X2_8829 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_289_), .Y(u2__abc_52155_new_n18251_));
AND2X2 AND2X2_883 ( .A(u2__abc_52155_new_n3779_), .B(u2__abc_52155_new_n3782_), .Y(u2__abc_52155_new_n3783_));
AND2X2 AND2X2_8830 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_287_), .Y(u2__abc_52155_new_n18252_));
AND2X2 AND2X2_8831 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18252_), .Y(u2__abc_52155_new_n18253_));
AND2X2 AND2X2_8832 ( .A(u2__abc_52155_new_n18254_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__289_));
AND2X2 AND2X2_8833 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_290_), .Y(u2__abc_52155_new_n18256_));
AND2X2 AND2X2_8834 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_288_), .Y(u2__abc_52155_new_n18257_));
AND2X2 AND2X2_8835 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18257_), .Y(u2__abc_52155_new_n18258_));
AND2X2 AND2X2_8836 ( .A(u2__abc_52155_new_n18259_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__290_));
AND2X2 AND2X2_8837 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_291_), .Y(u2__abc_52155_new_n18261_));
AND2X2 AND2X2_8838 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_289_), .Y(u2__abc_52155_new_n18262_));
AND2X2 AND2X2_8839 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18262_), .Y(u2__abc_52155_new_n18263_));
AND2X2 AND2X2_884 ( .A(u2__abc_52155_new_n3776_), .B(u2__abc_52155_new_n3783_), .Y(u2__abc_52155_new_n3784_));
AND2X2 AND2X2_8840 ( .A(u2__abc_52155_new_n18264_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__291_));
AND2X2 AND2X2_8841 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_292_), .Y(u2__abc_52155_new_n18266_));
AND2X2 AND2X2_8842 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_290_), .Y(u2__abc_52155_new_n18267_));
AND2X2 AND2X2_8843 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18267_), .Y(u2__abc_52155_new_n18268_));
AND2X2 AND2X2_8844 ( .A(u2__abc_52155_new_n18269_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__292_));
AND2X2 AND2X2_8845 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_293_), .Y(u2__abc_52155_new_n18271_));
AND2X2 AND2X2_8846 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_291_), .Y(u2__abc_52155_new_n18272_));
AND2X2 AND2X2_8847 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18272_), .Y(u2__abc_52155_new_n18273_));
AND2X2 AND2X2_8848 ( .A(u2__abc_52155_new_n18274_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__293_));
AND2X2 AND2X2_8849 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_294_), .Y(u2__abc_52155_new_n18276_));
AND2X2 AND2X2_885 ( .A(u2__abc_52155_new_n3785_), .B(u2_remHi_103_), .Y(u2__abc_52155_new_n3786_));
AND2X2 AND2X2_8850 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_292_), .Y(u2__abc_52155_new_n18277_));
AND2X2 AND2X2_8851 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18277_), .Y(u2__abc_52155_new_n18278_));
AND2X2 AND2X2_8852 ( .A(u2__abc_52155_new_n18279_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__294_));
AND2X2 AND2X2_8853 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_295_), .Y(u2__abc_52155_new_n18281_));
AND2X2 AND2X2_8854 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_293_), .Y(u2__abc_52155_new_n18282_));
AND2X2 AND2X2_8855 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18282_), .Y(u2__abc_52155_new_n18283_));
AND2X2 AND2X2_8856 ( .A(u2__abc_52155_new_n18284_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__295_));
AND2X2 AND2X2_8857 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_296_), .Y(u2__abc_52155_new_n18286_));
AND2X2 AND2X2_8858 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_294_), .Y(u2__abc_52155_new_n18287_));
AND2X2 AND2X2_8859 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18287_), .Y(u2__abc_52155_new_n18288_));
AND2X2 AND2X2_886 ( .A(u2__abc_52155_new_n3788_), .B(sqrto_103_), .Y(u2__abc_52155_new_n3789_));
AND2X2 AND2X2_8860 ( .A(u2__abc_52155_new_n18289_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__296_));
AND2X2 AND2X2_8861 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_297_), .Y(u2__abc_52155_new_n18291_));
AND2X2 AND2X2_8862 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_295_), .Y(u2__abc_52155_new_n18292_));
AND2X2 AND2X2_8863 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18292_), .Y(u2__abc_52155_new_n18293_));
AND2X2 AND2X2_8864 ( .A(u2__abc_52155_new_n18294_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__297_));
AND2X2 AND2X2_8865 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_298_), .Y(u2__abc_52155_new_n18296_));
AND2X2 AND2X2_8866 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_296_), .Y(u2__abc_52155_new_n18297_));
AND2X2 AND2X2_8867 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18297_), .Y(u2__abc_52155_new_n18298_));
AND2X2 AND2X2_8868 ( .A(u2__abc_52155_new_n18299_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__298_));
AND2X2 AND2X2_8869 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_299_), .Y(u2__abc_52155_new_n18301_));
AND2X2 AND2X2_887 ( .A(u2__abc_52155_new_n3787_), .B(u2__abc_52155_new_n3790_), .Y(u2__abc_52155_new_n3791_));
AND2X2 AND2X2_8870 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_297_), .Y(u2__abc_52155_new_n18302_));
AND2X2 AND2X2_8871 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18302_), .Y(u2__abc_52155_new_n18303_));
AND2X2 AND2X2_8872 ( .A(u2__abc_52155_new_n18304_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__299_));
AND2X2 AND2X2_8873 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_300_), .Y(u2__abc_52155_new_n18306_));
AND2X2 AND2X2_8874 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_298_), .Y(u2__abc_52155_new_n18307_));
AND2X2 AND2X2_8875 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18307_), .Y(u2__abc_52155_new_n18308_));
AND2X2 AND2X2_8876 ( .A(u2__abc_52155_new_n18309_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__300_));
AND2X2 AND2X2_8877 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_301_), .Y(u2__abc_52155_new_n18311_));
AND2X2 AND2X2_8878 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_299_), .Y(u2__abc_52155_new_n18312_));
AND2X2 AND2X2_8879 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18312_), .Y(u2__abc_52155_new_n18313_));
AND2X2 AND2X2_888 ( .A(u2__abc_52155_new_n3792_), .B(u2_remHi_102_), .Y(u2__abc_52155_new_n3793_));
AND2X2 AND2X2_8880 ( .A(u2__abc_52155_new_n18314_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__301_));
AND2X2 AND2X2_8881 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_302_), .Y(u2__abc_52155_new_n18316_));
AND2X2 AND2X2_8882 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_300_), .Y(u2__abc_52155_new_n18317_));
AND2X2 AND2X2_8883 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18317_), .Y(u2__abc_52155_new_n18318_));
AND2X2 AND2X2_8884 ( .A(u2__abc_52155_new_n18319_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__302_));
AND2X2 AND2X2_8885 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_303_), .Y(u2__abc_52155_new_n18321_));
AND2X2 AND2X2_8886 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_301_), .Y(u2__abc_52155_new_n18322_));
AND2X2 AND2X2_8887 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18322_), .Y(u2__abc_52155_new_n18323_));
AND2X2 AND2X2_8888 ( .A(u2__abc_52155_new_n18324_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__303_));
AND2X2 AND2X2_8889 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_304_), .Y(u2__abc_52155_new_n18326_));
AND2X2 AND2X2_889 ( .A(u2__abc_52155_new_n3795_), .B(sqrto_102_), .Y(u2__abc_52155_new_n3796_));
AND2X2 AND2X2_8890 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_302_), .Y(u2__abc_52155_new_n18327_));
AND2X2 AND2X2_8891 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18327_), .Y(u2__abc_52155_new_n18328_));
AND2X2 AND2X2_8892 ( .A(u2__abc_52155_new_n18329_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__304_));
AND2X2 AND2X2_8893 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_305_), .Y(u2__abc_52155_new_n18331_));
AND2X2 AND2X2_8894 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_303_), .Y(u2__abc_52155_new_n18332_));
AND2X2 AND2X2_8895 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18332_), .Y(u2__abc_52155_new_n18333_));
AND2X2 AND2X2_8896 ( .A(u2__abc_52155_new_n18334_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__305_));
AND2X2 AND2X2_8897 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_306_), .Y(u2__abc_52155_new_n18336_));
AND2X2 AND2X2_8898 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_304_), .Y(u2__abc_52155_new_n18337_));
AND2X2 AND2X2_8899 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18337_), .Y(u2__abc_52155_new_n18338_));
AND2X2 AND2X2_89 ( .A(_abc_73687_new_n867_), .B(_abc_73687_new_n866_), .Y(\o[124] ));
AND2X2 AND2X2_890 ( .A(u2__abc_52155_new_n3794_), .B(u2__abc_52155_new_n3797_), .Y(u2__abc_52155_new_n3798_));
AND2X2 AND2X2_8900 ( .A(u2__abc_52155_new_n18339_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__306_));
AND2X2 AND2X2_8901 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_307_), .Y(u2__abc_52155_new_n18341_));
AND2X2 AND2X2_8902 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_305_), .Y(u2__abc_52155_new_n18342_));
AND2X2 AND2X2_8903 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18342_), .Y(u2__abc_52155_new_n18343_));
AND2X2 AND2X2_8904 ( .A(u2__abc_52155_new_n18344_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__307_));
AND2X2 AND2X2_8905 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_308_), .Y(u2__abc_52155_new_n18346_));
AND2X2 AND2X2_8906 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_306_), .Y(u2__abc_52155_new_n18347_));
AND2X2 AND2X2_8907 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18347_), .Y(u2__abc_52155_new_n18348_));
AND2X2 AND2X2_8908 ( .A(u2__abc_52155_new_n18349_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__308_));
AND2X2 AND2X2_8909 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_309_), .Y(u2__abc_52155_new_n18351_));
AND2X2 AND2X2_891 ( .A(u2__abc_52155_new_n3791_), .B(u2__abc_52155_new_n3798_), .Y(u2__abc_52155_new_n3799_));
AND2X2 AND2X2_8910 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_307_), .Y(u2__abc_52155_new_n18352_));
AND2X2 AND2X2_8911 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18352_), .Y(u2__abc_52155_new_n18353_));
AND2X2 AND2X2_8912 ( .A(u2__abc_52155_new_n18354_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__309_));
AND2X2 AND2X2_8913 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_310_), .Y(u2__abc_52155_new_n18356_));
AND2X2 AND2X2_8914 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_308_), .Y(u2__abc_52155_new_n18357_));
AND2X2 AND2X2_8915 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18357_), .Y(u2__abc_52155_new_n18358_));
AND2X2 AND2X2_8916 ( .A(u2__abc_52155_new_n18359_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__310_));
AND2X2 AND2X2_8917 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_311_), .Y(u2__abc_52155_new_n18361_));
AND2X2 AND2X2_8918 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_309_), .Y(u2__abc_52155_new_n18362_));
AND2X2 AND2X2_8919 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18362_), .Y(u2__abc_52155_new_n18363_));
AND2X2 AND2X2_892 ( .A(u2__abc_52155_new_n3784_), .B(u2__abc_52155_new_n3799_), .Y(u2__abc_52155_new_n3800_));
AND2X2 AND2X2_8920 ( .A(u2__abc_52155_new_n18364_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__311_));
AND2X2 AND2X2_8921 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_312_), .Y(u2__abc_52155_new_n18366_));
AND2X2 AND2X2_8922 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_310_), .Y(u2__abc_52155_new_n18367_));
AND2X2 AND2X2_8923 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18367_), .Y(u2__abc_52155_new_n18368_));
AND2X2 AND2X2_8924 ( .A(u2__abc_52155_new_n18369_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__312_));
AND2X2 AND2X2_8925 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_313_), .Y(u2__abc_52155_new_n18371_));
AND2X2 AND2X2_8926 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_311_), .Y(u2__abc_52155_new_n18372_));
AND2X2 AND2X2_8927 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18372_), .Y(u2__abc_52155_new_n18373_));
AND2X2 AND2X2_8928 ( .A(u2__abc_52155_new_n18374_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__313_));
AND2X2 AND2X2_8929 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_314_), .Y(u2__abc_52155_new_n18376_));
AND2X2 AND2X2_893 ( .A(u2__abc_52155_new_n3801_), .B(u2_remHi_108_), .Y(u2__abc_52155_new_n3802_));
AND2X2 AND2X2_8930 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_312_), .Y(u2__abc_52155_new_n18377_));
AND2X2 AND2X2_8931 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18377_), .Y(u2__abc_52155_new_n18378_));
AND2X2 AND2X2_8932 ( .A(u2__abc_52155_new_n18379_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__314_));
AND2X2 AND2X2_8933 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_315_), .Y(u2__abc_52155_new_n18381_));
AND2X2 AND2X2_8934 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_313_), .Y(u2__abc_52155_new_n18382_));
AND2X2 AND2X2_8935 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18382_), .Y(u2__abc_52155_new_n18383_));
AND2X2 AND2X2_8936 ( .A(u2__abc_52155_new_n18384_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__315_));
AND2X2 AND2X2_8937 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_316_), .Y(u2__abc_52155_new_n18386_));
AND2X2 AND2X2_8938 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_314_), .Y(u2__abc_52155_new_n18387_));
AND2X2 AND2X2_8939 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18387_), .Y(u2__abc_52155_new_n18388_));
AND2X2 AND2X2_894 ( .A(u2__abc_52155_new_n3804_), .B(sqrto_108_), .Y(u2__abc_52155_new_n3805_));
AND2X2 AND2X2_8940 ( .A(u2__abc_52155_new_n18389_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__316_));
AND2X2 AND2X2_8941 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_317_), .Y(u2__abc_52155_new_n18391_));
AND2X2 AND2X2_8942 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_315_), .Y(u2__abc_52155_new_n18392_));
AND2X2 AND2X2_8943 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18392_), .Y(u2__abc_52155_new_n18393_));
AND2X2 AND2X2_8944 ( .A(u2__abc_52155_new_n18394_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__317_));
AND2X2 AND2X2_8945 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_318_), .Y(u2__abc_52155_new_n18396_));
AND2X2 AND2X2_8946 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_316_), .Y(u2__abc_52155_new_n18397_));
AND2X2 AND2X2_8947 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18397_), .Y(u2__abc_52155_new_n18398_));
AND2X2 AND2X2_8948 ( .A(u2__abc_52155_new_n18399_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__318_));
AND2X2 AND2X2_8949 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_319_), .Y(u2__abc_52155_new_n18401_));
AND2X2 AND2X2_895 ( .A(u2__abc_52155_new_n3803_), .B(u2__abc_52155_new_n3806_), .Y(u2__abc_52155_new_n3807_));
AND2X2 AND2X2_8950 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_317_), .Y(u2__abc_52155_new_n18402_));
AND2X2 AND2X2_8951 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18402_), .Y(u2__abc_52155_new_n18403_));
AND2X2 AND2X2_8952 ( .A(u2__abc_52155_new_n18404_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__319_));
AND2X2 AND2X2_8953 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_320_), .Y(u2__abc_52155_new_n18406_));
AND2X2 AND2X2_8954 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_318_), .Y(u2__abc_52155_new_n18407_));
AND2X2 AND2X2_8955 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18407_), .Y(u2__abc_52155_new_n18408_));
AND2X2 AND2X2_8956 ( .A(u2__abc_52155_new_n18409_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__320_));
AND2X2 AND2X2_8957 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_321_), .Y(u2__abc_52155_new_n18411_));
AND2X2 AND2X2_8958 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_319_), .Y(u2__abc_52155_new_n18412_));
AND2X2 AND2X2_8959 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18412_), .Y(u2__abc_52155_new_n18413_));
AND2X2 AND2X2_896 ( .A(u2__abc_52155_new_n3808_), .B(u2_remHi_109_), .Y(u2__abc_52155_new_n3809_));
AND2X2 AND2X2_8960 ( .A(u2__abc_52155_new_n18414_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__321_));
AND2X2 AND2X2_8961 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_322_), .Y(u2__abc_52155_new_n18416_));
AND2X2 AND2X2_8962 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_320_), .Y(u2__abc_52155_new_n18417_));
AND2X2 AND2X2_8963 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18417_), .Y(u2__abc_52155_new_n18418_));
AND2X2 AND2X2_8964 ( .A(u2__abc_52155_new_n18419_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__322_));
AND2X2 AND2X2_8965 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_323_), .Y(u2__abc_52155_new_n18421_));
AND2X2 AND2X2_8966 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_321_), .Y(u2__abc_52155_new_n18422_));
AND2X2 AND2X2_8967 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18422_), .Y(u2__abc_52155_new_n18423_));
AND2X2 AND2X2_8968 ( .A(u2__abc_52155_new_n18424_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__323_));
AND2X2 AND2X2_8969 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_324_), .Y(u2__abc_52155_new_n18426_));
AND2X2 AND2X2_897 ( .A(u2__abc_52155_new_n3811_), .B(sqrto_109_), .Y(u2__abc_52155_new_n3812_));
AND2X2 AND2X2_8970 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_322_), .Y(u2__abc_52155_new_n18427_));
AND2X2 AND2X2_8971 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18427_), .Y(u2__abc_52155_new_n18428_));
AND2X2 AND2X2_8972 ( .A(u2__abc_52155_new_n18429_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__324_));
AND2X2 AND2X2_8973 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_325_), .Y(u2__abc_52155_new_n18431_));
AND2X2 AND2X2_8974 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_323_), .Y(u2__abc_52155_new_n18432_));
AND2X2 AND2X2_8975 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18432_), .Y(u2__abc_52155_new_n18433_));
AND2X2 AND2X2_8976 ( .A(u2__abc_52155_new_n18434_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__325_));
AND2X2 AND2X2_8977 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_326_), .Y(u2__abc_52155_new_n18436_));
AND2X2 AND2X2_8978 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_324_), .Y(u2__abc_52155_new_n18437_));
AND2X2 AND2X2_8979 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18437_), .Y(u2__abc_52155_new_n18438_));
AND2X2 AND2X2_898 ( .A(u2__abc_52155_new_n3810_), .B(u2__abc_52155_new_n3813_), .Y(u2__abc_52155_new_n3814_));
AND2X2 AND2X2_8980 ( .A(u2__abc_52155_new_n18439_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__326_));
AND2X2 AND2X2_8981 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_327_), .Y(u2__abc_52155_new_n18441_));
AND2X2 AND2X2_8982 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_325_), .Y(u2__abc_52155_new_n18442_));
AND2X2 AND2X2_8983 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18442_), .Y(u2__abc_52155_new_n18443_));
AND2X2 AND2X2_8984 ( .A(u2__abc_52155_new_n18444_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__327_));
AND2X2 AND2X2_8985 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_328_), .Y(u2__abc_52155_new_n18446_));
AND2X2 AND2X2_8986 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_326_), .Y(u2__abc_52155_new_n18447_));
AND2X2 AND2X2_8987 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18447_), .Y(u2__abc_52155_new_n18448_));
AND2X2 AND2X2_8988 ( .A(u2__abc_52155_new_n18449_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__328_));
AND2X2 AND2X2_8989 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_329_), .Y(u2__abc_52155_new_n18451_));
AND2X2 AND2X2_899 ( .A(u2__abc_52155_new_n3807_), .B(u2__abc_52155_new_n3814_), .Y(u2__abc_52155_new_n3815_));
AND2X2 AND2X2_8990 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_327_), .Y(u2__abc_52155_new_n18452_));
AND2X2 AND2X2_8991 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18452_), .Y(u2__abc_52155_new_n18453_));
AND2X2 AND2X2_8992 ( .A(u2__abc_52155_new_n18454_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__329_));
AND2X2 AND2X2_8993 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_330_), .Y(u2__abc_52155_new_n18456_));
AND2X2 AND2X2_8994 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_328_), .Y(u2__abc_52155_new_n18457_));
AND2X2 AND2X2_8995 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18457_), .Y(u2__abc_52155_new_n18458_));
AND2X2 AND2X2_8996 ( .A(u2__abc_52155_new_n18459_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__330_));
AND2X2 AND2X2_8997 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_331_), .Y(u2__abc_52155_new_n18461_));
AND2X2 AND2X2_8998 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_329_), .Y(u2__abc_52155_new_n18462_));
AND2X2 AND2X2_8999 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18462_), .Y(u2__abc_52155_new_n18463_));
AND2X2 AND2X2_9 ( .A(_abc_73687_new_n753_), .B(sqrto_8_), .Y(\o[44] ));
AND2X2 AND2X2_90 ( .A(_abc_73687_new_n870_), .B(_abc_73687_new_n869_), .Y(\o[125] ));
AND2X2 AND2X2_900 ( .A(u2__abc_52155_new_n3816_), .B(u2_remHi_107_), .Y(u2__abc_52155_new_n3817_));
AND2X2 AND2X2_9000 ( .A(u2__abc_52155_new_n18464_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__331_));
AND2X2 AND2X2_9001 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_332_), .Y(u2__abc_52155_new_n18466_));
AND2X2 AND2X2_9002 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_330_), .Y(u2__abc_52155_new_n18467_));
AND2X2 AND2X2_9003 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18467_), .Y(u2__abc_52155_new_n18468_));
AND2X2 AND2X2_9004 ( .A(u2__abc_52155_new_n18469_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__332_));
AND2X2 AND2X2_9005 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_333_), .Y(u2__abc_52155_new_n18471_));
AND2X2 AND2X2_9006 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_331_), .Y(u2__abc_52155_new_n18472_));
AND2X2 AND2X2_9007 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18472_), .Y(u2__abc_52155_new_n18473_));
AND2X2 AND2X2_9008 ( .A(u2__abc_52155_new_n18474_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__333_));
AND2X2 AND2X2_9009 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_334_), .Y(u2__abc_52155_new_n18476_));
AND2X2 AND2X2_901 ( .A(u2__abc_52155_new_n3819_), .B(sqrto_107_), .Y(u2__abc_52155_new_n3820_));
AND2X2 AND2X2_9010 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_332_), .Y(u2__abc_52155_new_n18477_));
AND2X2 AND2X2_9011 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18477_), .Y(u2__abc_52155_new_n18478_));
AND2X2 AND2X2_9012 ( .A(u2__abc_52155_new_n18479_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__334_));
AND2X2 AND2X2_9013 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_335_), .Y(u2__abc_52155_new_n18481_));
AND2X2 AND2X2_9014 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_333_), .Y(u2__abc_52155_new_n18482_));
AND2X2 AND2X2_9015 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18482_), .Y(u2__abc_52155_new_n18483_));
AND2X2 AND2X2_9016 ( .A(u2__abc_52155_new_n18484_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__335_));
AND2X2 AND2X2_9017 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_336_), .Y(u2__abc_52155_new_n18486_));
AND2X2 AND2X2_9018 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_334_), .Y(u2__abc_52155_new_n18487_));
AND2X2 AND2X2_9019 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18487_), .Y(u2__abc_52155_new_n18488_));
AND2X2 AND2X2_902 ( .A(u2__abc_52155_new_n3818_), .B(u2__abc_52155_new_n3821_), .Y(u2__abc_52155_new_n3822_));
AND2X2 AND2X2_9020 ( .A(u2__abc_52155_new_n18489_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__336_));
AND2X2 AND2X2_9021 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_337_), .Y(u2__abc_52155_new_n18491_));
AND2X2 AND2X2_9022 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_335_), .Y(u2__abc_52155_new_n18492_));
AND2X2 AND2X2_9023 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18492_), .Y(u2__abc_52155_new_n18493_));
AND2X2 AND2X2_9024 ( .A(u2__abc_52155_new_n18494_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__337_));
AND2X2 AND2X2_9025 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_338_), .Y(u2__abc_52155_new_n18496_));
AND2X2 AND2X2_9026 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_336_), .Y(u2__abc_52155_new_n18497_));
AND2X2 AND2X2_9027 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18497_), .Y(u2__abc_52155_new_n18498_));
AND2X2 AND2X2_9028 ( .A(u2__abc_52155_new_n18499_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__338_));
AND2X2 AND2X2_9029 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_339_), .Y(u2__abc_52155_new_n18501_));
AND2X2 AND2X2_903 ( .A(u2__abc_52155_new_n3823_), .B(u2_remHi_106_), .Y(u2__abc_52155_new_n3824_));
AND2X2 AND2X2_9030 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_337_), .Y(u2__abc_52155_new_n18502_));
AND2X2 AND2X2_9031 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18502_), .Y(u2__abc_52155_new_n18503_));
AND2X2 AND2X2_9032 ( .A(u2__abc_52155_new_n18504_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__339_));
AND2X2 AND2X2_9033 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_340_), .Y(u2__abc_52155_new_n18506_));
AND2X2 AND2X2_9034 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_338_), .Y(u2__abc_52155_new_n18507_));
AND2X2 AND2X2_9035 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18507_), .Y(u2__abc_52155_new_n18508_));
AND2X2 AND2X2_9036 ( .A(u2__abc_52155_new_n18509_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__340_));
AND2X2 AND2X2_9037 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_341_), .Y(u2__abc_52155_new_n18511_));
AND2X2 AND2X2_9038 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_339_), .Y(u2__abc_52155_new_n18512_));
AND2X2 AND2X2_9039 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18512_), .Y(u2__abc_52155_new_n18513_));
AND2X2 AND2X2_904 ( .A(u2__abc_52155_new_n3826_), .B(sqrto_106_), .Y(u2__abc_52155_new_n3827_));
AND2X2 AND2X2_9040 ( .A(u2__abc_52155_new_n18514_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__341_));
AND2X2 AND2X2_9041 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_342_), .Y(u2__abc_52155_new_n18516_));
AND2X2 AND2X2_9042 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_340_), .Y(u2__abc_52155_new_n18517_));
AND2X2 AND2X2_9043 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18517_), .Y(u2__abc_52155_new_n18518_));
AND2X2 AND2X2_9044 ( .A(u2__abc_52155_new_n18519_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__342_));
AND2X2 AND2X2_9045 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_343_), .Y(u2__abc_52155_new_n18521_));
AND2X2 AND2X2_9046 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_341_), .Y(u2__abc_52155_new_n18522_));
AND2X2 AND2X2_9047 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18522_), .Y(u2__abc_52155_new_n18523_));
AND2X2 AND2X2_9048 ( .A(u2__abc_52155_new_n18524_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__343_));
AND2X2 AND2X2_9049 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_344_), .Y(u2__abc_52155_new_n18526_));
AND2X2 AND2X2_905 ( .A(u2__abc_52155_new_n3825_), .B(u2__abc_52155_new_n3828_), .Y(u2__abc_52155_new_n3829_));
AND2X2 AND2X2_9050 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_342_), .Y(u2__abc_52155_new_n18527_));
AND2X2 AND2X2_9051 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18527_), .Y(u2__abc_52155_new_n18528_));
AND2X2 AND2X2_9052 ( .A(u2__abc_52155_new_n18529_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__344_));
AND2X2 AND2X2_9053 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_345_), .Y(u2__abc_52155_new_n18531_));
AND2X2 AND2X2_9054 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_343_), .Y(u2__abc_52155_new_n18532_));
AND2X2 AND2X2_9055 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18532_), .Y(u2__abc_52155_new_n18533_));
AND2X2 AND2X2_9056 ( .A(u2__abc_52155_new_n18534_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__345_));
AND2X2 AND2X2_9057 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_346_), .Y(u2__abc_52155_new_n18536_));
AND2X2 AND2X2_9058 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_344_), .Y(u2__abc_52155_new_n18537_));
AND2X2 AND2X2_9059 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18537_), .Y(u2__abc_52155_new_n18538_));
AND2X2 AND2X2_906 ( .A(u2__abc_52155_new_n3822_), .B(u2__abc_52155_new_n3829_), .Y(u2__abc_52155_new_n3830_));
AND2X2 AND2X2_9060 ( .A(u2__abc_52155_new_n18539_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__346_));
AND2X2 AND2X2_9061 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_347_), .Y(u2__abc_52155_new_n18541_));
AND2X2 AND2X2_9062 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_345_), .Y(u2__abc_52155_new_n18542_));
AND2X2 AND2X2_9063 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18542_), .Y(u2__abc_52155_new_n18543_));
AND2X2 AND2X2_9064 ( .A(u2__abc_52155_new_n18544_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__347_));
AND2X2 AND2X2_9065 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_348_), .Y(u2__abc_52155_new_n18546_));
AND2X2 AND2X2_9066 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_346_), .Y(u2__abc_52155_new_n18547_));
AND2X2 AND2X2_9067 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18547_), .Y(u2__abc_52155_new_n18548_));
AND2X2 AND2X2_9068 ( .A(u2__abc_52155_new_n18549_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__348_));
AND2X2 AND2X2_9069 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_349_), .Y(u2__abc_52155_new_n18551_));
AND2X2 AND2X2_907 ( .A(u2__abc_52155_new_n3815_), .B(u2__abc_52155_new_n3830_), .Y(u2__abc_52155_new_n3831_));
AND2X2 AND2X2_9070 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_347_), .Y(u2__abc_52155_new_n18552_));
AND2X2 AND2X2_9071 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18552_), .Y(u2__abc_52155_new_n18553_));
AND2X2 AND2X2_9072 ( .A(u2__abc_52155_new_n18554_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__349_));
AND2X2 AND2X2_9073 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_350_), .Y(u2__abc_52155_new_n18556_));
AND2X2 AND2X2_9074 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_348_), .Y(u2__abc_52155_new_n18557_));
AND2X2 AND2X2_9075 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18557_), .Y(u2__abc_52155_new_n18558_));
AND2X2 AND2X2_9076 ( .A(u2__abc_52155_new_n18559_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__350_));
AND2X2 AND2X2_9077 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_351_), .Y(u2__abc_52155_new_n18561_));
AND2X2 AND2X2_9078 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_349_), .Y(u2__abc_52155_new_n18562_));
AND2X2 AND2X2_9079 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18562_), .Y(u2__abc_52155_new_n18563_));
AND2X2 AND2X2_908 ( .A(u2__abc_52155_new_n3800_), .B(u2__abc_52155_new_n3831_), .Y(u2__abc_52155_new_n3832_));
AND2X2 AND2X2_9080 ( .A(u2__abc_52155_new_n18564_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__351_));
AND2X2 AND2X2_9081 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_352_), .Y(u2__abc_52155_new_n18566_));
AND2X2 AND2X2_9082 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_350_), .Y(u2__abc_52155_new_n18567_));
AND2X2 AND2X2_9083 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18567_), .Y(u2__abc_52155_new_n18568_));
AND2X2 AND2X2_9084 ( .A(u2__abc_52155_new_n18569_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__352_));
AND2X2 AND2X2_9085 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_353_), .Y(u2__abc_52155_new_n18571_));
AND2X2 AND2X2_9086 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_351_), .Y(u2__abc_52155_new_n18572_));
AND2X2 AND2X2_9087 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18572_), .Y(u2__abc_52155_new_n18573_));
AND2X2 AND2X2_9088 ( .A(u2__abc_52155_new_n18574_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__353_));
AND2X2 AND2X2_9089 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_354_), .Y(u2__abc_52155_new_n18576_));
AND2X2 AND2X2_909 ( .A(u2__abc_52155_new_n3833_), .B(u2_remHi_96_), .Y(u2__abc_52155_new_n3834_));
AND2X2 AND2X2_9090 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_352_), .Y(u2__abc_52155_new_n18577_));
AND2X2 AND2X2_9091 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18577_), .Y(u2__abc_52155_new_n18578_));
AND2X2 AND2X2_9092 ( .A(u2__abc_52155_new_n18579_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__354_));
AND2X2 AND2X2_9093 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_355_), .Y(u2__abc_52155_new_n18581_));
AND2X2 AND2X2_9094 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_353_), .Y(u2__abc_52155_new_n18582_));
AND2X2 AND2X2_9095 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18582_), .Y(u2__abc_52155_new_n18583_));
AND2X2 AND2X2_9096 ( .A(u2__abc_52155_new_n18584_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__355_));
AND2X2 AND2X2_9097 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_356_), .Y(u2__abc_52155_new_n18586_));
AND2X2 AND2X2_9098 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_354_), .Y(u2__abc_52155_new_n18587_));
AND2X2 AND2X2_9099 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18587_), .Y(u2__abc_52155_new_n18588_));
AND2X2 AND2X2_91 ( .A(_abc_73687_new_n873_), .B(_abc_73687_new_n872_), .Y(\o[126] ));
AND2X2 AND2X2_910 ( .A(u2__abc_52155_new_n3835_), .B(sqrto_96_), .Y(u2__abc_52155_new_n3836_));
AND2X2 AND2X2_9100 ( .A(u2__abc_52155_new_n18589_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__356_));
AND2X2 AND2X2_9101 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_357_), .Y(u2__abc_52155_new_n18591_));
AND2X2 AND2X2_9102 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_355_), .Y(u2__abc_52155_new_n18592_));
AND2X2 AND2X2_9103 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18592_), .Y(u2__abc_52155_new_n18593_));
AND2X2 AND2X2_9104 ( .A(u2__abc_52155_new_n18594_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__357_));
AND2X2 AND2X2_9105 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_358_), .Y(u2__abc_52155_new_n18596_));
AND2X2 AND2X2_9106 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_356_), .Y(u2__abc_52155_new_n18597_));
AND2X2 AND2X2_9107 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18597_), .Y(u2__abc_52155_new_n18598_));
AND2X2 AND2X2_9108 ( .A(u2__abc_52155_new_n18599_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__358_));
AND2X2 AND2X2_9109 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_359_), .Y(u2__abc_52155_new_n18601_));
AND2X2 AND2X2_911 ( .A(u2__abc_52155_new_n3838_), .B(u2_remHi_97_), .Y(u2__abc_52155_new_n3839_));
AND2X2 AND2X2_9110 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_357_), .Y(u2__abc_52155_new_n18602_));
AND2X2 AND2X2_9111 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18602_), .Y(u2__abc_52155_new_n18603_));
AND2X2 AND2X2_9112 ( .A(u2__abc_52155_new_n18604_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__359_));
AND2X2 AND2X2_9113 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_360_), .Y(u2__abc_52155_new_n18606_));
AND2X2 AND2X2_9114 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_358_), .Y(u2__abc_52155_new_n18607_));
AND2X2 AND2X2_9115 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18607_), .Y(u2__abc_52155_new_n18608_));
AND2X2 AND2X2_9116 ( .A(u2__abc_52155_new_n18609_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__360_));
AND2X2 AND2X2_9117 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_361_), .Y(u2__abc_52155_new_n18611_));
AND2X2 AND2X2_9118 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_359_), .Y(u2__abc_52155_new_n18612_));
AND2X2 AND2X2_9119 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18612_), .Y(u2__abc_52155_new_n18613_));
AND2X2 AND2X2_912 ( .A(u2__abc_52155_new_n3840_), .B(sqrto_97_), .Y(u2__abc_52155_new_n3841_));
AND2X2 AND2X2_9120 ( .A(u2__abc_52155_new_n18614_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__361_));
AND2X2 AND2X2_9121 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_362_), .Y(u2__abc_52155_new_n18616_));
AND2X2 AND2X2_9122 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_360_), .Y(u2__abc_52155_new_n18617_));
AND2X2 AND2X2_9123 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18617_), .Y(u2__abc_52155_new_n18618_));
AND2X2 AND2X2_9124 ( .A(u2__abc_52155_new_n18619_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__362_));
AND2X2 AND2X2_9125 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_363_), .Y(u2__abc_52155_new_n18621_));
AND2X2 AND2X2_9126 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_361_), .Y(u2__abc_52155_new_n18622_));
AND2X2 AND2X2_9127 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18622_), .Y(u2__abc_52155_new_n18623_));
AND2X2 AND2X2_9128 ( .A(u2__abc_52155_new_n18624_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__363_));
AND2X2 AND2X2_9129 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_364_), .Y(u2__abc_52155_new_n18626_));
AND2X2 AND2X2_913 ( .A(u2__abc_52155_new_n3845_), .B(u2_remHi_95_), .Y(u2__abc_52155_new_n3846_));
AND2X2 AND2X2_9130 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_362_), .Y(u2__abc_52155_new_n18627_));
AND2X2 AND2X2_9131 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18627_), .Y(u2__abc_52155_new_n18628_));
AND2X2 AND2X2_9132 ( .A(u2__abc_52155_new_n18629_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__364_));
AND2X2 AND2X2_9133 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_365_), .Y(u2__abc_52155_new_n18631_));
AND2X2 AND2X2_9134 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_363_), .Y(u2__abc_52155_new_n18632_));
AND2X2 AND2X2_9135 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18632_), .Y(u2__abc_52155_new_n18633_));
AND2X2 AND2X2_9136 ( .A(u2__abc_52155_new_n18634_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__365_));
AND2X2 AND2X2_9137 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_366_), .Y(u2__abc_52155_new_n18636_));
AND2X2 AND2X2_9138 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_364_), .Y(u2__abc_52155_new_n18637_));
AND2X2 AND2X2_9139 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18637_), .Y(u2__abc_52155_new_n18638_));
AND2X2 AND2X2_914 ( .A(u2__abc_52155_new_n3848_), .B(sqrto_95_), .Y(u2__abc_52155_new_n3849_));
AND2X2 AND2X2_9140 ( .A(u2__abc_52155_new_n18639_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__366_));
AND2X2 AND2X2_9141 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_367_), .Y(u2__abc_52155_new_n18641_));
AND2X2 AND2X2_9142 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_365_), .Y(u2__abc_52155_new_n18642_));
AND2X2 AND2X2_9143 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18642_), .Y(u2__abc_52155_new_n18643_));
AND2X2 AND2X2_9144 ( .A(u2__abc_52155_new_n18644_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__367_));
AND2X2 AND2X2_9145 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_368_), .Y(u2__abc_52155_new_n18646_));
AND2X2 AND2X2_9146 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_366_), .Y(u2__abc_52155_new_n18647_));
AND2X2 AND2X2_9147 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18647_), .Y(u2__abc_52155_new_n18648_));
AND2X2 AND2X2_9148 ( .A(u2__abc_52155_new_n18649_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__368_));
AND2X2 AND2X2_9149 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_369_), .Y(u2__abc_52155_new_n18651_));
AND2X2 AND2X2_915 ( .A(u2__abc_52155_new_n3847_), .B(u2__abc_52155_new_n3850_), .Y(u2__abc_52155_new_n3851_));
AND2X2 AND2X2_9150 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_367_), .Y(u2__abc_52155_new_n18652_));
AND2X2 AND2X2_9151 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18652_), .Y(u2__abc_52155_new_n18653_));
AND2X2 AND2X2_9152 ( .A(u2__abc_52155_new_n18654_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__369_));
AND2X2 AND2X2_9153 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_370_), .Y(u2__abc_52155_new_n18656_));
AND2X2 AND2X2_9154 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_368_), .Y(u2__abc_52155_new_n18657_));
AND2X2 AND2X2_9155 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18657_), .Y(u2__abc_52155_new_n18658_));
AND2X2 AND2X2_9156 ( .A(u2__abc_52155_new_n18659_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__370_));
AND2X2 AND2X2_9157 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_371_), .Y(u2__abc_52155_new_n18661_));
AND2X2 AND2X2_9158 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_369_), .Y(u2__abc_52155_new_n18662_));
AND2X2 AND2X2_9159 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18662_), .Y(u2__abc_52155_new_n18663_));
AND2X2 AND2X2_916 ( .A(u2__abc_52155_new_n3852_), .B(u2_remHi_94_), .Y(u2__abc_52155_new_n3853_));
AND2X2 AND2X2_9160 ( .A(u2__abc_52155_new_n18664_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__371_));
AND2X2 AND2X2_9161 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_372_), .Y(u2__abc_52155_new_n18666_));
AND2X2 AND2X2_9162 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_370_), .Y(u2__abc_52155_new_n18667_));
AND2X2 AND2X2_9163 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18667_), .Y(u2__abc_52155_new_n18668_));
AND2X2 AND2X2_9164 ( .A(u2__abc_52155_new_n18669_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__372_));
AND2X2 AND2X2_9165 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_373_), .Y(u2__abc_52155_new_n18671_));
AND2X2 AND2X2_9166 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_371_), .Y(u2__abc_52155_new_n18672_));
AND2X2 AND2X2_9167 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18672_), .Y(u2__abc_52155_new_n18673_));
AND2X2 AND2X2_9168 ( .A(u2__abc_52155_new_n18674_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__373_));
AND2X2 AND2X2_9169 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_374_), .Y(u2__abc_52155_new_n18676_));
AND2X2 AND2X2_917 ( .A(u2__abc_52155_new_n3855_), .B(sqrto_94_), .Y(u2__abc_52155_new_n3856_));
AND2X2 AND2X2_9170 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_372_), .Y(u2__abc_52155_new_n18677_));
AND2X2 AND2X2_9171 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18677_), .Y(u2__abc_52155_new_n18678_));
AND2X2 AND2X2_9172 ( .A(u2__abc_52155_new_n18679_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__374_));
AND2X2 AND2X2_9173 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_375_), .Y(u2__abc_52155_new_n18681_));
AND2X2 AND2X2_9174 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_373_), .Y(u2__abc_52155_new_n18682_));
AND2X2 AND2X2_9175 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18682_), .Y(u2__abc_52155_new_n18683_));
AND2X2 AND2X2_9176 ( .A(u2__abc_52155_new_n18684_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__375_));
AND2X2 AND2X2_9177 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_376_), .Y(u2__abc_52155_new_n18686_));
AND2X2 AND2X2_9178 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_374_), .Y(u2__abc_52155_new_n18687_));
AND2X2 AND2X2_9179 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18687_), .Y(u2__abc_52155_new_n18688_));
AND2X2 AND2X2_918 ( .A(u2__abc_52155_new_n3854_), .B(u2__abc_52155_new_n3857_), .Y(u2__abc_52155_new_n3858_));
AND2X2 AND2X2_9180 ( .A(u2__abc_52155_new_n18689_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__376_));
AND2X2 AND2X2_9181 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_377_), .Y(u2__abc_52155_new_n18691_));
AND2X2 AND2X2_9182 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_375_), .Y(u2__abc_52155_new_n18692_));
AND2X2 AND2X2_9183 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18692_), .Y(u2__abc_52155_new_n18693_));
AND2X2 AND2X2_9184 ( .A(u2__abc_52155_new_n18694_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__377_));
AND2X2 AND2X2_9185 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_378_), .Y(u2__abc_52155_new_n18696_));
AND2X2 AND2X2_9186 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_376_), .Y(u2__abc_52155_new_n18697_));
AND2X2 AND2X2_9187 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18697_), .Y(u2__abc_52155_new_n18698_));
AND2X2 AND2X2_9188 ( .A(u2__abc_52155_new_n18699_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__378_));
AND2X2 AND2X2_9189 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_379_), .Y(u2__abc_52155_new_n18701_));
AND2X2 AND2X2_919 ( .A(u2__abc_52155_new_n3851_), .B(u2__abc_52155_new_n3858_), .Y(u2__abc_52155_new_n3859_));
AND2X2 AND2X2_9190 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_377_), .Y(u2__abc_52155_new_n18702_));
AND2X2 AND2X2_9191 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18702_), .Y(u2__abc_52155_new_n18703_));
AND2X2 AND2X2_9192 ( .A(u2__abc_52155_new_n18704_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__379_));
AND2X2 AND2X2_9193 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_380_), .Y(u2__abc_52155_new_n18706_));
AND2X2 AND2X2_9194 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_378_), .Y(u2__abc_52155_new_n18707_));
AND2X2 AND2X2_9195 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18707_), .Y(u2__abc_52155_new_n18708_));
AND2X2 AND2X2_9196 ( .A(u2__abc_52155_new_n18709_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__380_));
AND2X2 AND2X2_9197 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_381_), .Y(u2__abc_52155_new_n18711_));
AND2X2 AND2X2_9198 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_379_), .Y(u2__abc_52155_new_n18712_));
AND2X2 AND2X2_9199 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18712_), .Y(u2__abc_52155_new_n18713_));
AND2X2 AND2X2_92 ( .A(_abc_73687_new_n876_), .B(_abc_73687_new_n875_), .Y(\o[127] ));
AND2X2 AND2X2_920 ( .A(u2__abc_52155_new_n3844_), .B(u2__abc_52155_new_n3859_), .Y(u2__abc_52155_new_n3860_));
AND2X2 AND2X2_9200 ( .A(u2__abc_52155_new_n18714_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__381_));
AND2X2 AND2X2_9201 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_382_), .Y(u2__abc_52155_new_n18716_));
AND2X2 AND2X2_9202 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_380_), .Y(u2__abc_52155_new_n18717_));
AND2X2 AND2X2_9203 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18717_), .Y(u2__abc_52155_new_n18718_));
AND2X2 AND2X2_9204 ( .A(u2__abc_52155_new_n18719_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__382_));
AND2X2 AND2X2_9205 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_383_), .Y(u2__abc_52155_new_n18721_));
AND2X2 AND2X2_9206 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_381_), .Y(u2__abc_52155_new_n18722_));
AND2X2 AND2X2_9207 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18722_), .Y(u2__abc_52155_new_n18723_));
AND2X2 AND2X2_9208 ( .A(u2__abc_52155_new_n18724_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__383_));
AND2X2 AND2X2_9209 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_384_), .Y(u2__abc_52155_new_n18726_));
AND2X2 AND2X2_921 ( .A(u2__abc_52155_new_n3861_), .B(u2_remHi_100_), .Y(u2__abc_52155_new_n3862_));
AND2X2 AND2X2_9210 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_382_), .Y(u2__abc_52155_new_n18727_));
AND2X2 AND2X2_9211 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18727_), .Y(u2__abc_52155_new_n18728_));
AND2X2 AND2X2_9212 ( .A(u2__abc_52155_new_n18729_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__384_));
AND2X2 AND2X2_9213 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_385_), .Y(u2__abc_52155_new_n18731_));
AND2X2 AND2X2_9214 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_383_), .Y(u2__abc_52155_new_n18732_));
AND2X2 AND2X2_9215 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18732_), .Y(u2__abc_52155_new_n18733_));
AND2X2 AND2X2_9216 ( .A(u2__abc_52155_new_n18734_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__385_));
AND2X2 AND2X2_9217 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_386_), .Y(u2__abc_52155_new_n18736_));
AND2X2 AND2X2_9218 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_384_), .Y(u2__abc_52155_new_n18737_));
AND2X2 AND2X2_9219 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18737_), .Y(u2__abc_52155_new_n18738_));
AND2X2 AND2X2_922 ( .A(u2__abc_52155_new_n3864_), .B(sqrto_100_), .Y(u2__abc_52155_new_n3865_));
AND2X2 AND2X2_9220 ( .A(u2__abc_52155_new_n18739_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__386_));
AND2X2 AND2X2_9221 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_387_), .Y(u2__abc_52155_new_n18741_));
AND2X2 AND2X2_9222 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_385_), .Y(u2__abc_52155_new_n18742_));
AND2X2 AND2X2_9223 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18742_), .Y(u2__abc_52155_new_n18743_));
AND2X2 AND2X2_9224 ( .A(u2__abc_52155_new_n18744_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__387_));
AND2X2 AND2X2_9225 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_388_), .Y(u2__abc_52155_new_n18746_));
AND2X2 AND2X2_9226 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_386_), .Y(u2__abc_52155_new_n18747_));
AND2X2 AND2X2_9227 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18747_), .Y(u2__abc_52155_new_n18748_));
AND2X2 AND2X2_9228 ( .A(u2__abc_52155_new_n18749_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__388_));
AND2X2 AND2X2_9229 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_389_), .Y(u2__abc_52155_new_n18751_));
AND2X2 AND2X2_923 ( .A(u2__abc_52155_new_n3863_), .B(u2__abc_52155_new_n3866_), .Y(u2__abc_52155_new_n3867_));
AND2X2 AND2X2_9230 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_387_), .Y(u2__abc_52155_new_n18752_));
AND2X2 AND2X2_9231 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18752_), .Y(u2__abc_52155_new_n18753_));
AND2X2 AND2X2_9232 ( .A(u2__abc_52155_new_n18754_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__389_));
AND2X2 AND2X2_9233 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_390_), .Y(u2__abc_52155_new_n18756_));
AND2X2 AND2X2_9234 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_388_), .Y(u2__abc_52155_new_n18757_));
AND2X2 AND2X2_9235 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18757_), .Y(u2__abc_52155_new_n18758_));
AND2X2 AND2X2_9236 ( .A(u2__abc_52155_new_n18759_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__390_));
AND2X2 AND2X2_9237 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_391_), .Y(u2__abc_52155_new_n18761_));
AND2X2 AND2X2_9238 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_389_), .Y(u2__abc_52155_new_n18762_));
AND2X2 AND2X2_9239 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18762_), .Y(u2__abc_52155_new_n18763_));
AND2X2 AND2X2_924 ( .A(u2__abc_52155_new_n3868_), .B(u2_remHi_101_), .Y(u2__abc_52155_new_n3869_));
AND2X2 AND2X2_9240 ( .A(u2__abc_52155_new_n18764_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__391_));
AND2X2 AND2X2_9241 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_392_), .Y(u2__abc_52155_new_n18766_));
AND2X2 AND2X2_9242 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_390_), .Y(u2__abc_52155_new_n18767_));
AND2X2 AND2X2_9243 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18767_), .Y(u2__abc_52155_new_n18768_));
AND2X2 AND2X2_9244 ( .A(u2__abc_52155_new_n18769_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__392_));
AND2X2 AND2X2_9245 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_393_), .Y(u2__abc_52155_new_n18771_));
AND2X2 AND2X2_9246 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_391_), .Y(u2__abc_52155_new_n18772_));
AND2X2 AND2X2_9247 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18772_), .Y(u2__abc_52155_new_n18773_));
AND2X2 AND2X2_9248 ( .A(u2__abc_52155_new_n18774_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__393_));
AND2X2 AND2X2_9249 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_394_), .Y(u2__abc_52155_new_n18776_));
AND2X2 AND2X2_925 ( .A(u2__abc_52155_new_n3871_), .B(sqrto_101_), .Y(u2__abc_52155_new_n3872_));
AND2X2 AND2X2_9250 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_392_), .Y(u2__abc_52155_new_n18777_));
AND2X2 AND2X2_9251 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18777_), .Y(u2__abc_52155_new_n18778_));
AND2X2 AND2X2_9252 ( .A(u2__abc_52155_new_n18779_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__394_));
AND2X2 AND2X2_9253 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_395_), .Y(u2__abc_52155_new_n18781_));
AND2X2 AND2X2_9254 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_393_), .Y(u2__abc_52155_new_n18782_));
AND2X2 AND2X2_9255 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18782_), .Y(u2__abc_52155_new_n18783_));
AND2X2 AND2X2_9256 ( .A(u2__abc_52155_new_n18784_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__395_));
AND2X2 AND2X2_9257 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_396_), .Y(u2__abc_52155_new_n18786_));
AND2X2 AND2X2_9258 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_394_), .Y(u2__abc_52155_new_n18787_));
AND2X2 AND2X2_9259 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18787_), .Y(u2__abc_52155_new_n18788_));
AND2X2 AND2X2_926 ( .A(u2__abc_52155_new_n3870_), .B(u2__abc_52155_new_n3873_), .Y(u2__abc_52155_new_n3874_));
AND2X2 AND2X2_9260 ( .A(u2__abc_52155_new_n18789_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__396_));
AND2X2 AND2X2_9261 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_397_), .Y(u2__abc_52155_new_n18791_));
AND2X2 AND2X2_9262 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_395_), .Y(u2__abc_52155_new_n18792_));
AND2X2 AND2X2_9263 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18792_), .Y(u2__abc_52155_new_n18793_));
AND2X2 AND2X2_9264 ( .A(u2__abc_52155_new_n18794_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__397_));
AND2X2 AND2X2_9265 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_398_), .Y(u2__abc_52155_new_n18796_));
AND2X2 AND2X2_9266 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_396_), .Y(u2__abc_52155_new_n18797_));
AND2X2 AND2X2_9267 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18797_), .Y(u2__abc_52155_new_n18798_));
AND2X2 AND2X2_9268 ( .A(u2__abc_52155_new_n18799_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__398_));
AND2X2 AND2X2_9269 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_399_), .Y(u2__abc_52155_new_n18801_));
AND2X2 AND2X2_927 ( .A(u2__abc_52155_new_n3867_), .B(u2__abc_52155_new_n3874_), .Y(u2__abc_52155_new_n3875_));
AND2X2 AND2X2_9270 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_397_), .Y(u2__abc_52155_new_n18802_));
AND2X2 AND2X2_9271 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18802_), .Y(u2__abc_52155_new_n18803_));
AND2X2 AND2X2_9272 ( .A(u2__abc_52155_new_n18804_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__399_));
AND2X2 AND2X2_9273 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_400_), .Y(u2__abc_52155_new_n18806_));
AND2X2 AND2X2_9274 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_398_), .Y(u2__abc_52155_new_n18807_));
AND2X2 AND2X2_9275 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18807_), .Y(u2__abc_52155_new_n18808_));
AND2X2 AND2X2_9276 ( .A(u2__abc_52155_new_n18809_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__400_));
AND2X2 AND2X2_9277 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_401_), .Y(u2__abc_52155_new_n18811_));
AND2X2 AND2X2_9278 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_399_), .Y(u2__abc_52155_new_n18812_));
AND2X2 AND2X2_9279 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18812_), .Y(u2__abc_52155_new_n18813_));
AND2X2 AND2X2_928 ( .A(u2__abc_52155_new_n3876_), .B(u2_remHi_99_), .Y(u2__abc_52155_new_n3877_));
AND2X2 AND2X2_9280 ( .A(u2__abc_52155_new_n18814_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__401_));
AND2X2 AND2X2_9281 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_402_), .Y(u2__abc_52155_new_n18816_));
AND2X2 AND2X2_9282 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_400_), .Y(u2__abc_52155_new_n18817_));
AND2X2 AND2X2_9283 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18817_), .Y(u2__abc_52155_new_n18818_));
AND2X2 AND2X2_9284 ( .A(u2__abc_52155_new_n18819_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__402_));
AND2X2 AND2X2_9285 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_403_), .Y(u2__abc_52155_new_n18821_));
AND2X2 AND2X2_9286 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_401_), .Y(u2__abc_52155_new_n18822_));
AND2X2 AND2X2_9287 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18822_), .Y(u2__abc_52155_new_n18823_));
AND2X2 AND2X2_9288 ( .A(u2__abc_52155_new_n18824_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__403_));
AND2X2 AND2X2_9289 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_404_), .Y(u2__abc_52155_new_n18826_));
AND2X2 AND2X2_929 ( .A(u2__abc_52155_new_n3879_), .B(sqrto_99_), .Y(u2__abc_52155_new_n3880_));
AND2X2 AND2X2_9290 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_402_), .Y(u2__abc_52155_new_n18827_));
AND2X2 AND2X2_9291 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18827_), .Y(u2__abc_52155_new_n18828_));
AND2X2 AND2X2_9292 ( .A(u2__abc_52155_new_n18829_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__404_));
AND2X2 AND2X2_9293 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_405_), .Y(u2__abc_52155_new_n18831_));
AND2X2 AND2X2_9294 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_403_), .Y(u2__abc_52155_new_n18832_));
AND2X2 AND2X2_9295 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18832_), .Y(u2__abc_52155_new_n18833_));
AND2X2 AND2X2_9296 ( .A(u2__abc_52155_new_n18834_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__405_));
AND2X2 AND2X2_9297 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_406_), .Y(u2__abc_52155_new_n18836_));
AND2X2 AND2X2_9298 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_404_), .Y(u2__abc_52155_new_n18837_));
AND2X2 AND2X2_9299 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18837_), .Y(u2__abc_52155_new_n18838_));
AND2X2 AND2X2_93 ( .A(_abc_73687_new_n879_), .B(_abc_73687_new_n878_), .Y(\o[128] ));
AND2X2 AND2X2_930 ( .A(u2__abc_52155_new_n3878_), .B(u2__abc_52155_new_n3881_), .Y(u2__abc_52155_new_n3882_));
AND2X2 AND2X2_9300 ( .A(u2__abc_52155_new_n18839_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__406_));
AND2X2 AND2X2_9301 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_407_), .Y(u2__abc_52155_new_n18841_));
AND2X2 AND2X2_9302 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_405_), .Y(u2__abc_52155_new_n18842_));
AND2X2 AND2X2_9303 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18842_), .Y(u2__abc_52155_new_n18843_));
AND2X2 AND2X2_9304 ( .A(u2__abc_52155_new_n18844_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__407_));
AND2X2 AND2X2_9305 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_408_), .Y(u2__abc_52155_new_n18846_));
AND2X2 AND2X2_9306 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_406_), .Y(u2__abc_52155_new_n18847_));
AND2X2 AND2X2_9307 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18847_), .Y(u2__abc_52155_new_n18848_));
AND2X2 AND2X2_9308 ( .A(u2__abc_52155_new_n18849_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__408_));
AND2X2 AND2X2_9309 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_409_), .Y(u2__abc_52155_new_n18851_));
AND2X2 AND2X2_931 ( .A(u2__abc_52155_new_n3883_), .B(u2_remHi_98_), .Y(u2__abc_52155_new_n3884_));
AND2X2 AND2X2_9310 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_407_), .Y(u2__abc_52155_new_n18852_));
AND2X2 AND2X2_9311 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18852_), .Y(u2__abc_52155_new_n18853_));
AND2X2 AND2X2_9312 ( .A(u2__abc_52155_new_n18854_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__409_));
AND2X2 AND2X2_9313 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_410_), .Y(u2__abc_52155_new_n18856_));
AND2X2 AND2X2_9314 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_408_), .Y(u2__abc_52155_new_n18857_));
AND2X2 AND2X2_9315 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18857_), .Y(u2__abc_52155_new_n18858_));
AND2X2 AND2X2_9316 ( .A(u2__abc_52155_new_n18859_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__410_));
AND2X2 AND2X2_9317 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_411_), .Y(u2__abc_52155_new_n18861_));
AND2X2 AND2X2_9318 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_409_), .Y(u2__abc_52155_new_n18862_));
AND2X2 AND2X2_9319 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18862_), .Y(u2__abc_52155_new_n18863_));
AND2X2 AND2X2_932 ( .A(u2__abc_52155_new_n3886_), .B(sqrto_98_), .Y(u2__abc_52155_new_n3887_));
AND2X2 AND2X2_9320 ( .A(u2__abc_52155_new_n18864_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__411_));
AND2X2 AND2X2_9321 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_412_), .Y(u2__abc_52155_new_n18866_));
AND2X2 AND2X2_9322 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_410_), .Y(u2__abc_52155_new_n18867_));
AND2X2 AND2X2_9323 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18867_), .Y(u2__abc_52155_new_n18868_));
AND2X2 AND2X2_9324 ( .A(u2__abc_52155_new_n18869_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__412_));
AND2X2 AND2X2_9325 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_413_), .Y(u2__abc_52155_new_n18871_));
AND2X2 AND2X2_9326 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_411_), .Y(u2__abc_52155_new_n18872_));
AND2X2 AND2X2_9327 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18872_), .Y(u2__abc_52155_new_n18873_));
AND2X2 AND2X2_9328 ( .A(u2__abc_52155_new_n18874_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__413_));
AND2X2 AND2X2_9329 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_414_), .Y(u2__abc_52155_new_n18876_));
AND2X2 AND2X2_933 ( .A(u2__abc_52155_new_n3885_), .B(u2__abc_52155_new_n3888_), .Y(u2__abc_52155_new_n3889_));
AND2X2 AND2X2_9330 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_412_), .Y(u2__abc_52155_new_n18877_));
AND2X2 AND2X2_9331 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18877_), .Y(u2__abc_52155_new_n18878_));
AND2X2 AND2X2_9332 ( .A(u2__abc_52155_new_n18879_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__414_));
AND2X2 AND2X2_9333 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_415_), .Y(u2__abc_52155_new_n18881_));
AND2X2 AND2X2_9334 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_413_), .Y(u2__abc_52155_new_n18882_));
AND2X2 AND2X2_9335 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18882_), .Y(u2__abc_52155_new_n18883_));
AND2X2 AND2X2_9336 ( .A(u2__abc_52155_new_n18884_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__415_));
AND2X2 AND2X2_9337 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_416_), .Y(u2__abc_52155_new_n18886_));
AND2X2 AND2X2_9338 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_414_), .Y(u2__abc_52155_new_n18887_));
AND2X2 AND2X2_9339 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18887_), .Y(u2__abc_52155_new_n18888_));
AND2X2 AND2X2_934 ( .A(u2__abc_52155_new_n3882_), .B(u2__abc_52155_new_n3889_), .Y(u2__abc_52155_new_n3890_));
AND2X2 AND2X2_9340 ( .A(u2__abc_52155_new_n18889_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__416_));
AND2X2 AND2X2_9341 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_417_), .Y(u2__abc_52155_new_n18891_));
AND2X2 AND2X2_9342 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_415_), .Y(u2__abc_52155_new_n18892_));
AND2X2 AND2X2_9343 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18892_), .Y(u2__abc_52155_new_n18893_));
AND2X2 AND2X2_9344 ( .A(u2__abc_52155_new_n18894_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__417_));
AND2X2 AND2X2_9345 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_418_), .Y(u2__abc_52155_new_n18896_));
AND2X2 AND2X2_9346 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_416_), .Y(u2__abc_52155_new_n18897_));
AND2X2 AND2X2_9347 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18897_), .Y(u2__abc_52155_new_n18898_));
AND2X2 AND2X2_9348 ( .A(u2__abc_52155_new_n18899_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__418_));
AND2X2 AND2X2_9349 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_419_), .Y(u2__abc_52155_new_n18901_));
AND2X2 AND2X2_935 ( .A(u2__abc_52155_new_n3875_), .B(u2__abc_52155_new_n3890_), .Y(u2__abc_52155_new_n3891_));
AND2X2 AND2X2_9350 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_417_), .Y(u2__abc_52155_new_n18902_));
AND2X2 AND2X2_9351 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18902_), .Y(u2__abc_52155_new_n18903_));
AND2X2 AND2X2_9352 ( .A(u2__abc_52155_new_n18904_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__419_));
AND2X2 AND2X2_9353 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_420_), .Y(u2__abc_52155_new_n18906_));
AND2X2 AND2X2_9354 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_418_), .Y(u2__abc_52155_new_n18907_));
AND2X2 AND2X2_9355 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18907_), .Y(u2__abc_52155_new_n18908_));
AND2X2 AND2X2_9356 ( .A(u2__abc_52155_new_n18909_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__420_));
AND2X2 AND2X2_9357 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_421_), .Y(u2__abc_52155_new_n18911_));
AND2X2 AND2X2_9358 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_419_), .Y(u2__abc_52155_new_n18912_));
AND2X2 AND2X2_9359 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18912_), .Y(u2__abc_52155_new_n18913_));
AND2X2 AND2X2_936 ( .A(u2__abc_52155_new_n3860_), .B(u2__abc_52155_new_n3891_), .Y(u2__abc_52155_new_n3892_));
AND2X2 AND2X2_9360 ( .A(u2__abc_52155_new_n18914_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__421_));
AND2X2 AND2X2_9361 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_422_), .Y(u2__abc_52155_new_n18916_));
AND2X2 AND2X2_9362 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_420_), .Y(u2__abc_52155_new_n18917_));
AND2X2 AND2X2_9363 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18917_), .Y(u2__abc_52155_new_n18918_));
AND2X2 AND2X2_9364 ( .A(u2__abc_52155_new_n18919_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__422_));
AND2X2 AND2X2_9365 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_423_), .Y(u2__abc_52155_new_n18921_));
AND2X2 AND2X2_9366 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_421_), .Y(u2__abc_52155_new_n18922_));
AND2X2 AND2X2_9367 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18922_), .Y(u2__abc_52155_new_n18923_));
AND2X2 AND2X2_9368 ( .A(u2__abc_52155_new_n18924_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__423_));
AND2X2 AND2X2_9369 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_424_), .Y(u2__abc_52155_new_n18926_));
AND2X2 AND2X2_937 ( .A(u2__abc_52155_new_n3892_), .B(u2__abc_52155_new_n3832_), .Y(u2__abc_52155_new_n3893_));
AND2X2 AND2X2_9370 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_422_), .Y(u2__abc_52155_new_n18927_));
AND2X2 AND2X2_9371 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18927_), .Y(u2__abc_52155_new_n18928_));
AND2X2 AND2X2_9372 ( .A(u2__abc_52155_new_n18929_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__424_));
AND2X2 AND2X2_9373 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_425_), .Y(u2__abc_52155_new_n18931_));
AND2X2 AND2X2_9374 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_423_), .Y(u2__abc_52155_new_n18932_));
AND2X2 AND2X2_9375 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18932_), .Y(u2__abc_52155_new_n18933_));
AND2X2 AND2X2_9376 ( .A(u2__abc_52155_new_n18934_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__425_));
AND2X2 AND2X2_9377 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_426_), .Y(u2__abc_52155_new_n18936_));
AND2X2 AND2X2_9378 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_424_), .Y(u2__abc_52155_new_n18937_));
AND2X2 AND2X2_9379 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18937_), .Y(u2__abc_52155_new_n18938_));
AND2X2 AND2X2_938 ( .A(u2__abc_52155_new_n3893_), .B(u2__abc_52155_new_n3769_), .Y(u2__abc_52155_new_n3894_));
AND2X2 AND2X2_9380 ( .A(u2__abc_52155_new_n18939_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__426_));
AND2X2 AND2X2_9381 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_427_), .Y(u2__abc_52155_new_n18941_));
AND2X2 AND2X2_9382 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_425_), .Y(u2__abc_52155_new_n18942_));
AND2X2 AND2X2_9383 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18942_), .Y(u2__abc_52155_new_n18943_));
AND2X2 AND2X2_9384 ( .A(u2__abc_52155_new_n18944_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__427_));
AND2X2 AND2X2_9385 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_428_), .Y(u2__abc_52155_new_n18946_));
AND2X2 AND2X2_9386 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_426_), .Y(u2__abc_52155_new_n18947_));
AND2X2 AND2X2_9387 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18947_), .Y(u2__abc_52155_new_n18948_));
AND2X2 AND2X2_9388 ( .A(u2__abc_52155_new_n18949_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__428_));
AND2X2 AND2X2_9389 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_429_), .Y(u2__abc_52155_new_n18951_));
AND2X2 AND2X2_939 ( .A(u2__abc_52155_new_n3895_), .B(u2_remHi_92_), .Y(u2__abc_52155_new_n3896_));
AND2X2 AND2X2_9390 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_427_), .Y(u2__abc_52155_new_n18952_));
AND2X2 AND2X2_9391 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18952_), .Y(u2__abc_52155_new_n18953_));
AND2X2 AND2X2_9392 ( .A(u2__abc_52155_new_n18954_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__429_));
AND2X2 AND2X2_9393 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_430_), .Y(u2__abc_52155_new_n18956_));
AND2X2 AND2X2_9394 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_428_), .Y(u2__abc_52155_new_n18957_));
AND2X2 AND2X2_9395 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18957_), .Y(u2__abc_52155_new_n18958_));
AND2X2 AND2X2_9396 ( .A(u2__abc_52155_new_n18959_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__430_));
AND2X2 AND2X2_9397 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_431_), .Y(u2__abc_52155_new_n18961_));
AND2X2 AND2X2_9398 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_429_), .Y(u2__abc_52155_new_n18962_));
AND2X2 AND2X2_9399 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18962_), .Y(u2__abc_52155_new_n18963_));
AND2X2 AND2X2_94 ( .A(_abc_73687_new_n882_), .B(_abc_73687_new_n881_), .Y(\o[129] ));
AND2X2 AND2X2_940 ( .A(u2__abc_52155_new_n3898_), .B(sqrto_92_), .Y(u2__abc_52155_new_n3899_));
AND2X2 AND2X2_9400 ( .A(u2__abc_52155_new_n18964_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__431_));
AND2X2 AND2X2_9401 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_432_), .Y(u2__abc_52155_new_n18966_));
AND2X2 AND2X2_9402 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_430_), .Y(u2__abc_52155_new_n18967_));
AND2X2 AND2X2_9403 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18967_), .Y(u2__abc_52155_new_n18968_));
AND2X2 AND2X2_9404 ( .A(u2__abc_52155_new_n18969_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__432_));
AND2X2 AND2X2_9405 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_433_), .Y(u2__abc_52155_new_n18971_));
AND2X2 AND2X2_9406 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_431_), .Y(u2__abc_52155_new_n18972_));
AND2X2 AND2X2_9407 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18972_), .Y(u2__abc_52155_new_n18973_));
AND2X2 AND2X2_9408 ( .A(u2__abc_52155_new_n18974_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__433_));
AND2X2 AND2X2_9409 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_434_), .Y(u2__abc_52155_new_n18976_));
AND2X2 AND2X2_941 ( .A(u2__abc_52155_new_n3897_), .B(u2__abc_52155_new_n3900_), .Y(u2__abc_52155_new_n3901_));
AND2X2 AND2X2_9410 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_432_), .Y(u2__abc_52155_new_n18977_));
AND2X2 AND2X2_9411 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18977_), .Y(u2__abc_52155_new_n18978_));
AND2X2 AND2X2_9412 ( .A(u2__abc_52155_new_n18979_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__434_));
AND2X2 AND2X2_9413 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_435_), .Y(u2__abc_52155_new_n18981_));
AND2X2 AND2X2_9414 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_433_), .Y(u2__abc_52155_new_n18982_));
AND2X2 AND2X2_9415 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18982_), .Y(u2__abc_52155_new_n18983_));
AND2X2 AND2X2_9416 ( .A(u2__abc_52155_new_n18984_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__435_));
AND2X2 AND2X2_9417 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_436_), .Y(u2__abc_52155_new_n18986_));
AND2X2 AND2X2_9418 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_434_), .Y(u2__abc_52155_new_n18987_));
AND2X2 AND2X2_9419 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18987_), .Y(u2__abc_52155_new_n18988_));
AND2X2 AND2X2_942 ( .A(u2__abc_52155_new_n3902_), .B(u2_remHi_93_), .Y(u2__abc_52155_new_n3903_));
AND2X2 AND2X2_9420 ( .A(u2__abc_52155_new_n18989_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__436_));
AND2X2 AND2X2_9421 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_437_), .Y(u2__abc_52155_new_n18991_));
AND2X2 AND2X2_9422 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_435_), .Y(u2__abc_52155_new_n18992_));
AND2X2 AND2X2_9423 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18992_), .Y(u2__abc_52155_new_n18993_));
AND2X2 AND2X2_9424 ( .A(u2__abc_52155_new_n18994_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__437_));
AND2X2 AND2X2_9425 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_438_), .Y(u2__abc_52155_new_n18996_));
AND2X2 AND2X2_9426 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_436_), .Y(u2__abc_52155_new_n18997_));
AND2X2 AND2X2_9427 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n18997_), .Y(u2__abc_52155_new_n18998_));
AND2X2 AND2X2_9428 ( .A(u2__abc_52155_new_n18999_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__438_));
AND2X2 AND2X2_9429 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_439_), .Y(u2__abc_52155_new_n19001_));
AND2X2 AND2X2_943 ( .A(u2__abc_52155_new_n3905_), .B(sqrto_93_), .Y(u2__abc_52155_new_n3906_));
AND2X2 AND2X2_9430 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_437_), .Y(u2__abc_52155_new_n19002_));
AND2X2 AND2X2_9431 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19002_), .Y(u2__abc_52155_new_n19003_));
AND2X2 AND2X2_9432 ( .A(u2__abc_52155_new_n19004_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__439_));
AND2X2 AND2X2_9433 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_440_), .Y(u2__abc_52155_new_n19006_));
AND2X2 AND2X2_9434 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_438_), .Y(u2__abc_52155_new_n19007_));
AND2X2 AND2X2_9435 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19007_), .Y(u2__abc_52155_new_n19008_));
AND2X2 AND2X2_9436 ( .A(u2__abc_52155_new_n19009_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__440_));
AND2X2 AND2X2_9437 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_441_), .Y(u2__abc_52155_new_n19011_));
AND2X2 AND2X2_9438 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_439_), .Y(u2__abc_52155_new_n19012_));
AND2X2 AND2X2_9439 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19012_), .Y(u2__abc_52155_new_n19013_));
AND2X2 AND2X2_944 ( .A(u2__abc_52155_new_n3904_), .B(u2__abc_52155_new_n3907_), .Y(u2__abc_52155_new_n3908_));
AND2X2 AND2X2_9440 ( .A(u2__abc_52155_new_n19014_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__441_));
AND2X2 AND2X2_9441 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_442_), .Y(u2__abc_52155_new_n19016_));
AND2X2 AND2X2_9442 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_440_), .Y(u2__abc_52155_new_n19017_));
AND2X2 AND2X2_9443 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19017_), .Y(u2__abc_52155_new_n19018_));
AND2X2 AND2X2_9444 ( .A(u2__abc_52155_new_n19019_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__442_));
AND2X2 AND2X2_9445 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_443_), .Y(u2__abc_52155_new_n19021_));
AND2X2 AND2X2_9446 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_441_), .Y(u2__abc_52155_new_n19022_));
AND2X2 AND2X2_9447 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19022_), .Y(u2__abc_52155_new_n19023_));
AND2X2 AND2X2_9448 ( .A(u2__abc_52155_new_n19024_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__443_));
AND2X2 AND2X2_9449 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_444_), .Y(u2__abc_52155_new_n19026_));
AND2X2 AND2X2_945 ( .A(u2__abc_52155_new_n3901_), .B(u2__abc_52155_new_n3908_), .Y(u2__abc_52155_new_n3909_));
AND2X2 AND2X2_9450 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_442_), .Y(u2__abc_52155_new_n19027_));
AND2X2 AND2X2_9451 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19027_), .Y(u2__abc_52155_new_n19028_));
AND2X2 AND2X2_9452 ( .A(u2__abc_52155_new_n19029_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__444_));
AND2X2 AND2X2_9453 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_445_), .Y(u2__abc_52155_new_n19031_));
AND2X2 AND2X2_9454 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_443_), .Y(u2__abc_52155_new_n19032_));
AND2X2 AND2X2_9455 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19032_), .Y(u2__abc_52155_new_n19033_));
AND2X2 AND2X2_9456 ( .A(u2__abc_52155_new_n19034_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__445_));
AND2X2 AND2X2_9457 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_446_), .Y(u2__abc_52155_new_n19036_));
AND2X2 AND2X2_9458 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_444_), .Y(u2__abc_52155_new_n19037_));
AND2X2 AND2X2_9459 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19037_), .Y(u2__abc_52155_new_n19038_));
AND2X2 AND2X2_946 ( .A(u2__abc_52155_new_n3910_), .B(u2_remHi_91_), .Y(u2__abc_52155_new_n3911_));
AND2X2 AND2X2_9460 ( .A(u2__abc_52155_new_n19039_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__446_));
AND2X2 AND2X2_9461 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_447_), .Y(u2__abc_52155_new_n19041_));
AND2X2 AND2X2_9462 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_445_), .Y(u2__abc_52155_new_n19042_));
AND2X2 AND2X2_9463 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19042_), .Y(u2__abc_52155_new_n19043_));
AND2X2 AND2X2_9464 ( .A(u2__abc_52155_new_n19044_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__447_));
AND2X2 AND2X2_9465 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_448_), .Y(u2__abc_52155_new_n19046_));
AND2X2 AND2X2_9466 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_446_), .Y(u2__abc_52155_new_n19047_));
AND2X2 AND2X2_9467 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19047_), .Y(u2__abc_52155_new_n19048_));
AND2X2 AND2X2_9468 ( .A(u2__abc_52155_new_n19049_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__448_));
AND2X2 AND2X2_9469 ( .A(u2__abc_52155_new_n16522_), .B(u2_remLo_449_), .Y(u2__abc_52155_new_n19051_));
AND2X2 AND2X2_947 ( .A(u2__abc_52155_new_n3913_), .B(sqrto_91_), .Y(u2__abc_52155_new_n3914_));
AND2X2 AND2X2_9470 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_447_), .Y(u2__abc_52155_new_n19052_));
AND2X2 AND2X2_9471 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19052_), .Y(u2__abc_52155_new_n19053_));
AND2X2 AND2X2_9472 ( .A(u2__abc_52155_new_n19054_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__449_));
AND2X2 AND2X2_9473 ( .A(u2__abc_52155_new_n16522_), .B(u2_remHiShift_0_), .Y(u2__abc_52155_new_n19056_));
AND2X2 AND2X2_9474 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_448_), .Y(u2__abc_52155_new_n19057_));
AND2X2 AND2X2_9475 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19057_), .Y(u2__abc_52155_new_n19058_));
AND2X2 AND2X2_9476 ( .A(u2__abc_52155_new_n19059_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__450_));
AND2X2 AND2X2_9477 ( .A(u2__abc_52155_new_n16522_), .B(u2_remHiShift_1_), .Y(u2__abc_52155_new_n19061_));
AND2X2 AND2X2_9478 ( .A(u2__abc_52155_new_n2999_), .B(u2_remLo_449_), .Y(u2__abc_52155_new_n19062_));
AND2X2 AND2X2_9479 ( .A(u2__abc_52155_new_n16470_), .B(u2__abc_52155_new_n19062_), .Y(u2__abc_52155_new_n19063_));
AND2X2 AND2X2_948 ( .A(u2__abc_52155_new_n3912_), .B(u2__abc_52155_new_n3915_), .Y(u2__abc_52155_new_n3916_));
AND2X2 AND2X2_9480 ( .A(u2__abc_52155_new_n19064_), .B(u2__abc_52155_new_n2962_), .Y(u2__0remLo_451_0__451_));
AND2X2 AND2X2_9481 ( .A(u2__abc_52155_new_n2962_), .B(u2_root_0_), .Y(u2__abc_52155_new_n19066_));
AND2X2 AND2X2_9482 ( .A(u2__abc_52155_new_n16522_), .B(u2__abc_52155_new_n19066_), .Y(u2__0root_452_0__0_));
AND2X2 AND2X2_9483 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_0_), .Y(u2__abc_52155_new_n19068_));
AND2X2 AND2X2_9484 ( .A(u2__abc_52155_new_n7622_), .B(u2_root_0_), .Y(u2__abc_52155_new_n19069_));
AND2X2 AND2X2_9485 ( .A(u2__abc_52155_new_n19070_), .B(u2__abc_52155_new_n19071_), .Y(u2__abc_52155_new_n19072_));
AND2X2 AND2X2_9486 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3114_), .Y(u2__abc_52155_new_n19074_));
AND2X2 AND2X2_9487 ( .A(u2__abc_52155_new_n19075_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19076_));
AND2X2 AND2X2_9488 ( .A(u2__abc_52155_new_n19073_), .B(u2__abc_52155_new_n19076_), .Y(u2__abc_52155_new_n19077_));
AND2X2 AND2X2_9489 ( .A(u2__abc_52155_new_n19078_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__1_));
AND2X2 AND2X2_949 ( .A(u2__abc_52155_new_n3917_), .B(u2_remHi_90_), .Y(u2__abc_52155_new_n3918_));
AND2X2 AND2X2_9490 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_1_), .Y(u2__abc_52155_new_n19080_));
AND2X2 AND2X2_9491 ( .A(u2__abc_52155_new_n19069_), .B(sqrto_0_), .Y(u2__abc_52155_new_n19081_));
AND2X2 AND2X2_9492 ( .A(u2__abc_52155_new_n19082_), .B(u2__abc_52155_new_n19083_), .Y(u2__abc_52155_new_n19084_));
AND2X2 AND2X2_9493 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3121_), .Y(u2__abc_52155_new_n19086_));
AND2X2 AND2X2_9494 ( .A(u2__abc_52155_new_n19087_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19088_));
AND2X2 AND2X2_9495 ( .A(u2__abc_52155_new_n19085_), .B(u2__abc_52155_new_n19088_), .Y(u2__abc_52155_new_n19089_));
AND2X2 AND2X2_9496 ( .A(u2__abc_52155_new_n19090_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__2_));
AND2X2 AND2X2_9497 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_2_), .Y(u2__abc_52155_new_n19092_));
AND2X2 AND2X2_9498 ( .A(u2__abc_52155_new_n19081_), .B(sqrto_1_), .Y(u2__abc_52155_new_n19094_));
AND2X2 AND2X2_9499 ( .A(u2__abc_52155_new_n19095_), .B(u2__abc_52155_new_n19093_), .Y(u2__abc_52155_new_n19096_));
AND2X2 AND2X2_95 ( .A(_abc_73687_new_n885_), .B(_abc_73687_new_n884_), .Y(\o[130] ));
AND2X2 AND2X2_950 ( .A(u2__abc_52155_new_n3920_), .B(sqrto_90_), .Y(u2__abc_52155_new_n3921_));
AND2X2 AND2X2_9500 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3107_), .Y(u2__abc_52155_new_n19098_));
AND2X2 AND2X2_9501 ( .A(u2__abc_52155_new_n19099_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19100_));
AND2X2 AND2X2_9502 ( .A(u2__abc_52155_new_n19097_), .B(u2__abc_52155_new_n19100_), .Y(u2__abc_52155_new_n19101_));
AND2X2 AND2X2_9503 ( .A(u2__abc_52155_new_n19102_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__3_));
AND2X2 AND2X2_9504 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_3_), .Y(u2__abc_52155_new_n19104_));
AND2X2 AND2X2_9505 ( .A(u2__abc_52155_new_n19094_), .B(sqrto_2_), .Y(u2__abc_52155_new_n19106_));
AND2X2 AND2X2_9506 ( .A(u2__abc_52155_new_n19107_), .B(u2__abc_52155_new_n19105_), .Y(u2__abc_52155_new_n19108_));
AND2X2 AND2X2_9507 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3102_), .Y(u2__abc_52155_new_n19110_));
AND2X2 AND2X2_9508 ( .A(u2__abc_52155_new_n19111_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19112_));
AND2X2 AND2X2_9509 ( .A(u2__abc_52155_new_n19109_), .B(u2__abc_52155_new_n19112_), .Y(u2__abc_52155_new_n19113_));
AND2X2 AND2X2_951 ( .A(u2__abc_52155_new_n3919_), .B(u2__abc_52155_new_n3922_), .Y(u2__abc_52155_new_n3923_));
AND2X2 AND2X2_9510 ( .A(u2__abc_52155_new_n19114_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__4_));
AND2X2 AND2X2_9511 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_4_), .Y(u2__abc_52155_new_n19116_));
AND2X2 AND2X2_9512 ( .A(u2__abc_52155_new_n19106_), .B(sqrto_3_), .Y(u2__abc_52155_new_n19118_));
AND2X2 AND2X2_9513 ( .A(u2__abc_52155_new_n19119_), .B(u2__abc_52155_new_n19117_), .Y(u2__abc_52155_new_n19120_));
AND2X2 AND2X2_9514 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3091_), .Y(u2__abc_52155_new_n19122_));
AND2X2 AND2X2_9515 ( .A(u2__abc_52155_new_n19123_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19124_));
AND2X2 AND2X2_9516 ( .A(u2__abc_52155_new_n19121_), .B(u2__abc_52155_new_n19124_), .Y(u2__abc_52155_new_n19125_));
AND2X2 AND2X2_9517 ( .A(u2__abc_52155_new_n19126_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__5_));
AND2X2 AND2X2_9518 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_5_), .Y(u2__abc_52155_new_n19128_));
AND2X2 AND2X2_9519 ( .A(u2__abc_52155_new_n19118_), .B(sqrto_4_), .Y(u2__abc_52155_new_n19130_));
AND2X2 AND2X2_952 ( .A(u2__abc_52155_new_n3916_), .B(u2__abc_52155_new_n3923_), .Y(u2__abc_52155_new_n3924_));
AND2X2 AND2X2_9520 ( .A(u2__abc_52155_new_n19131_), .B(u2__abc_52155_new_n19129_), .Y(u2__abc_52155_new_n19132_));
AND2X2 AND2X2_9521 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3098_), .Y(u2__abc_52155_new_n19134_));
AND2X2 AND2X2_9522 ( .A(u2__abc_52155_new_n19135_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19136_));
AND2X2 AND2X2_9523 ( .A(u2__abc_52155_new_n19133_), .B(u2__abc_52155_new_n19136_), .Y(u2__abc_52155_new_n19137_));
AND2X2 AND2X2_9524 ( .A(u2__abc_52155_new_n19138_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__6_));
AND2X2 AND2X2_9525 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_6_), .Y(u2__abc_52155_new_n19140_));
AND2X2 AND2X2_9526 ( .A(u2__abc_52155_new_n19130_), .B(sqrto_5_), .Y(u2__abc_52155_new_n19142_));
AND2X2 AND2X2_9527 ( .A(u2__abc_52155_new_n19143_), .B(u2__abc_52155_new_n19141_), .Y(u2__abc_52155_new_n19144_));
AND2X2 AND2X2_9528 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3084_), .Y(u2__abc_52155_new_n19146_));
AND2X2 AND2X2_9529 ( .A(u2__abc_52155_new_n19147_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19148_));
AND2X2 AND2X2_953 ( .A(u2__abc_52155_new_n3909_), .B(u2__abc_52155_new_n3924_), .Y(u2__abc_52155_new_n3925_));
AND2X2 AND2X2_9530 ( .A(u2__abc_52155_new_n19145_), .B(u2__abc_52155_new_n19148_), .Y(u2__abc_52155_new_n19149_));
AND2X2 AND2X2_9531 ( .A(u2__abc_52155_new_n19150_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__7_));
AND2X2 AND2X2_9532 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_7_), .Y(u2__abc_52155_new_n19152_));
AND2X2 AND2X2_9533 ( .A(u2__abc_52155_new_n19142_), .B(sqrto_6_), .Y(u2__abc_52155_new_n19154_));
AND2X2 AND2X2_9534 ( .A(u2__abc_52155_new_n19155_), .B(u2__abc_52155_new_n19153_), .Y(u2__abc_52155_new_n19156_));
AND2X2 AND2X2_9535 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3077_), .Y(u2__abc_52155_new_n19158_));
AND2X2 AND2X2_9536 ( .A(u2__abc_52155_new_n19159_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19160_));
AND2X2 AND2X2_9537 ( .A(u2__abc_52155_new_n19157_), .B(u2__abc_52155_new_n19160_), .Y(u2__abc_52155_new_n19161_));
AND2X2 AND2X2_9538 ( .A(u2__abc_52155_new_n19162_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__8_));
AND2X2 AND2X2_9539 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_8_), .Y(u2__abc_52155_new_n19164_));
AND2X2 AND2X2_954 ( .A(u2__abc_52155_new_n3926_), .B(u2_remHi_88_), .Y(u2__abc_52155_new_n3927_));
AND2X2 AND2X2_9540 ( .A(u2__abc_52155_new_n19154_), .B(sqrto_7_), .Y(u2__abc_52155_new_n19166_));
AND2X2 AND2X2_9541 ( .A(u2__abc_52155_new_n19167_), .B(u2__abc_52155_new_n19165_), .Y(u2__abc_52155_new_n19168_));
AND2X2 AND2X2_9542 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3063_), .Y(u2__abc_52155_new_n19170_));
AND2X2 AND2X2_9543 ( .A(u2__abc_52155_new_n19171_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19172_));
AND2X2 AND2X2_9544 ( .A(u2__abc_52155_new_n19169_), .B(u2__abc_52155_new_n19172_), .Y(u2__abc_52155_new_n19173_));
AND2X2 AND2X2_9545 ( .A(u2__abc_52155_new_n19174_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__9_));
AND2X2 AND2X2_9546 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_9_), .Y(u2__abc_52155_new_n19176_));
AND2X2 AND2X2_9547 ( .A(u2__abc_52155_new_n19166_), .B(sqrto_8_), .Y(u2__abc_52155_new_n19178_));
AND2X2 AND2X2_9548 ( .A(u2__abc_52155_new_n19179_), .B(u2__abc_52155_new_n19177_), .Y(u2__abc_52155_new_n19180_));
AND2X2 AND2X2_9549 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3069_), .Y(u2__abc_52155_new_n19182_));
AND2X2 AND2X2_955 ( .A(u2__abc_52155_new_n3929_), .B(sqrto_88_), .Y(u2__abc_52155_new_n3930_));
AND2X2 AND2X2_9550 ( .A(u2__abc_52155_new_n19183_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19184_));
AND2X2 AND2X2_9551 ( .A(u2__abc_52155_new_n19181_), .B(u2__abc_52155_new_n19184_), .Y(u2__abc_52155_new_n19185_));
AND2X2 AND2X2_9552 ( .A(u2__abc_52155_new_n19186_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__10_));
AND2X2 AND2X2_9553 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_10_), .Y(u2__abc_52155_new_n19188_));
AND2X2 AND2X2_9554 ( .A(u2__abc_52155_new_n19178_), .B(sqrto_9_), .Y(u2__abc_52155_new_n19190_));
AND2X2 AND2X2_9555 ( .A(u2__abc_52155_new_n19191_), .B(u2__abc_52155_new_n19189_), .Y(u2__abc_52155_new_n19192_));
AND2X2 AND2X2_9556 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3055_), .Y(u2__abc_52155_new_n19194_));
AND2X2 AND2X2_9557 ( .A(u2__abc_52155_new_n19195_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19196_));
AND2X2 AND2X2_9558 ( .A(u2__abc_52155_new_n19193_), .B(u2__abc_52155_new_n19196_), .Y(u2__abc_52155_new_n19197_));
AND2X2 AND2X2_9559 ( .A(u2__abc_52155_new_n19198_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__11_));
AND2X2 AND2X2_956 ( .A(u2__abc_52155_new_n3928_), .B(u2__abc_52155_new_n3931_), .Y(u2__abc_52155_new_n3932_));
AND2X2 AND2X2_9560 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_11_), .Y(u2__abc_52155_new_n19200_));
AND2X2 AND2X2_9561 ( .A(u2__abc_52155_new_n19190_), .B(sqrto_10_), .Y(u2__abc_52155_new_n19202_));
AND2X2 AND2X2_9562 ( .A(u2__abc_52155_new_n19203_), .B(u2__abc_52155_new_n19201_), .Y(u2__abc_52155_new_n19204_));
AND2X2 AND2X2_9563 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3048_), .Y(u2__abc_52155_new_n19206_));
AND2X2 AND2X2_9564 ( .A(u2__abc_52155_new_n19207_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19208_));
AND2X2 AND2X2_9565 ( .A(u2__abc_52155_new_n19205_), .B(u2__abc_52155_new_n19208_), .Y(u2__abc_52155_new_n19209_));
AND2X2 AND2X2_9566 ( .A(u2__abc_52155_new_n19210_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__12_));
AND2X2 AND2X2_9567 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_12_), .Y(u2__abc_52155_new_n19212_));
AND2X2 AND2X2_9568 ( .A(u2__abc_52155_new_n19202_), .B(sqrto_11_), .Y(u2__abc_52155_new_n19214_));
AND2X2 AND2X2_9569 ( .A(u2__abc_52155_new_n19215_), .B(u2__abc_52155_new_n19213_), .Y(u2__abc_52155_new_n19216_));
AND2X2 AND2X2_957 ( .A(u2__abc_52155_new_n3933_), .B(u2_remHi_89_), .Y(u2__abc_52155_new_n3934_));
AND2X2 AND2X2_9570 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3035_), .Y(u2__abc_52155_new_n19218_));
AND2X2 AND2X2_9571 ( .A(u2__abc_52155_new_n19219_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19220_));
AND2X2 AND2X2_9572 ( .A(u2__abc_52155_new_n19217_), .B(u2__abc_52155_new_n19220_), .Y(u2__abc_52155_new_n19221_));
AND2X2 AND2X2_9573 ( .A(u2__abc_52155_new_n19222_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__13_));
AND2X2 AND2X2_9574 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_13_), .Y(u2__abc_52155_new_n19224_));
AND2X2 AND2X2_9575 ( .A(u2__abc_52155_new_n19214_), .B(sqrto_12_), .Y(u2__abc_52155_new_n19226_));
AND2X2 AND2X2_9576 ( .A(u2__abc_52155_new_n19227_), .B(u2__abc_52155_new_n19225_), .Y(u2__abc_52155_new_n19228_));
AND2X2 AND2X2_9577 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3043_), .Y(u2__abc_52155_new_n19230_));
AND2X2 AND2X2_9578 ( .A(u2__abc_52155_new_n19231_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19232_));
AND2X2 AND2X2_9579 ( .A(u2__abc_52155_new_n19229_), .B(u2__abc_52155_new_n19232_), .Y(u2__abc_52155_new_n19233_));
AND2X2 AND2X2_958 ( .A(u2__abc_52155_new_n3936_), .B(sqrto_89_), .Y(u2__abc_52155_new_n3937_));
AND2X2 AND2X2_9580 ( .A(u2__abc_52155_new_n19234_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__14_));
AND2X2 AND2X2_9581 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_14_), .Y(u2__abc_52155_new_n19236_));
AND2X2 AND2X2_9582 ( .A(u2__abc_52155_new_n19226_), .B(sqrto_13_), .Y(u2__abc_52155_new_n19238_));
AND2X2 AND2X2_9583 ( .A(u2__abc_52155_new_n19239_), .B(u2__abc_52155_new_n19237_), .Y(u2__abc_52155_new_n19240_));
AND2X2 AND2X2_9584 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3239_), .Y(u2__abc_52155_new_n19242_));
AND2X2 AND2X2_9585 ( .A(u2__abc_52155_new_n19243_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19244_));
AND2X2 AND2X2_9586 ( .A(u2__abc_52155_new_n19241_), .B(u2__abc_52155_new_n19244_), .Y(u2__abc_52155_new_n19245_));
AND2X2 AND2X2_9587 ( .A(u2__abc_52155_new_n19246_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__15_));
AND2X2 AND2X2_9588 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_15_), .Y(u2__abc_52155_new_n19248_));
AND2X2 AND2X2_9589 ( .A(u2__abc_52155_new_n19238_), .B(sqrto_14_), .Y(u2__abc_52155_new_n19250_));
AND2X2 AND2X2_959 ( .A(u2__abc_52155_new_n3935_), .B(u2__abc_52155_new_n3938_), .Y(u2__abc_52155_new_n3939_));
AND2X2 AND2X2_9590 ( .A(u2__abc_52155_new_n19251_), .B(u2__abc_52155_new_n19249_), .Y(u2__abc_52155_new_n19252_));
AND2X2 AND2X2_9591 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3244_), .Y(u2__abc_52155_new_n19254_));
AND2X2 AND2X2_9592 ( .A(u2__abc_52155_new_n19255_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19256_));
AND2X2 AND2X2_9593 ( .A(u2__abc_52155_new_n19253_), .B(u2__abc_52155_new_n19256_), .Y(u2__abc_52155_new_n19257_));
AND2X2 AND2X2_9594 ( .A(u2__abc_52155_new_n19258_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__16_));
AND2X2 AND2X2_9595 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_16_), .Y(u2__abc_52155_new_n19260_));
AND2X2 AND2X2_9596 ( .A(u2__abc_52155_new_n19250_), .B(sqrto_15_), .Y(u2__abc_52155_new_n19262_));
AND2X2 AND2X2_9597 ( .A(u2__abc_52155_new_n19263_), .B(u2__abc_52155_new_n19261_), .Y(u2__abc_52155_new_n19264_));
AND2X2 AND2X2_9598 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3227_), .Y(u2__abc_52155_new_n19266_));
AND2X2 AND2X2_9599 ( .A(u2__abc_52155_new_n19267_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19268_));
AND2X2 AND2X2_96 ( .A(_abc_73687_new_n888_), .B(_abc_73687_new_n887_), .Y(\o[131] ));
AND2X2 AND2X2_960 ( .A(u2__abc_52155_new_n3932_), .B(u2__abc_52155_new_n3939_), .Y(u2__abc_52155_new_n3940_));
AND2X2 AND2X2_9600 ( .A(u2__abc_52155_new_n19265_), .B(u2__abc_52155_new_n19268_), .Y(u2__abc_52155_new_n19269_));
AND2X2 AND2X2_9601 ( .A(u2__abc_52155_new_n19270_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__17_));
AND2X2 AND2X2_9602 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_17_), .Y(u2__abc_52155_new_n19272_));
AND2X2 AND2X2_9603 ( .A(u2__abc_52155_new_n19262_), .B(sqrto_16_), .Y(u2__abc_52155_new_n19274_));
AND2X2 AND2X2_9604 ( .A(u2__abc_52155_new_n19275_), .B(u2__abc_52155_new_n19273_), .Y(u2__abc_52155_new_n19276_));
AND2X2 AND2X2_9605 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3232_), .Y(u2__abc_52155_new_n19278_));
AND2X2 AND2X2_9606 ( .A(u2__abc_52155_new_n19279_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19280_));
AND2X2 AND2X2_9607 ( .A(u2__abc_52155_new_n19277_), .B(u2__abc_52155_new_n19280_), .Y(u2__abc_52155_new_n19281_));
AND2X2 AND2X2_9608 ( .A(u2__abc_52155_new_n19282_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__18_));
AND2X2 AND2X2_9609 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_18_), .Y(u2__abc_52155_new_n19284_));
AND2X2 AND2X2_961 ( .A(u2__abc_52155_new_n3941_), .B(u2_remHi_87_), .Y(u2__abc_52155_new_n3942_));
AND2X2 AND2X2_9610 ( .A(u2__abc_52155_new_n19274_), .B(sqrto_17_), .Y(u2__abc_52155_new_n19286_));
AND2X2 AND2X2_9611 ( .A(u2__abc_52155_new_n19287_), .B(u2__abc_52155_new_n19285_), .Y(u2__abc_52155_new_n19288_));
AND2X2 AND2X2_9612 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3269_), .Y(u2__abc_52155_new_n19290_));
AND2X2 AND2X2_9613 ( .A(u2__abc_52155_new_n19291_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19292_));
AND2X2 AND2X2_9614 ( .A(u2__abc_52155_new_n19289_), .B(u2__abc_52155_new_n19292_), .Y(u2__abc_52155_new_n19293_));
AND2X2 AND2X2_9615 ( .A(u2__abc_52155_new_n19294_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__19_));
AND2X2 AND2X2_9616 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_19_), .Y(u2__abc_52155_new_n19296_));
AND2X2 AND2X2_9617 ( .A(u2__abc_52155_new_n19286_), .B(sqrto_18_), .Y(u2__abc_52155_new_n19298_));
AND2X2 AND2X2_9618 ( .A(u2__abc_52155_new_n19299_), .B(u2__abc_52155_new_n19297_), .Y(u2__abc_52155_new_n19300_));
AND2X2 AND2X2_9619 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3264_), .Y(u2__abc_52155_new_n19302_));
AND2X2 AND2X2_962 ( .A(u2__abc_52155_new_n3944_), .B(sqrto_87_), .Y(u2__abc_52155_new_n3945_));
AND2X2 AND2X2_9620 ( .A(u2__abc_52155_new_n19303_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19304_));
AND2X2 AND2X2_9621 ( .A(u2__abc_52155_new_n19301_), .B(u2__abc_52155_new_n19304_), .Y(u2__abc_52155_new_n19305_));
AND2X2 AND2X2_9622 ( .A(u2__abc_52155_new_n19306_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__20_));
AND2X2 AND2X2_9623 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_20_), .Y(u2__abc_52155_new_n19308_));
AND2X2 AND2X2_9624 ( .A(u2__abc_52155_new_n19298_), .B(sqrto_19_), .Y(u2__abc_52155_new_n19310_));
AND2X2 AND2X2_9625 ( .A(u2__abc_52155_new_n19311_), .B(u2__abc_52155_new_n19309_), .Y(u2__abc_52155_new_n19312_));
AND2X2 AND2X2_9626 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3253_), .Y(u2__abc_52155_new_n19314_));
AND2X2 AND2X2_9627 ( .A(u2__abc_52155_new_n19315_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19316_));
AND2X2 AND2X2_9628 ( .A(u2__abc_52155_new_n19313_), .B(u2__abc_52155_new_n19316_), .Y(u2__abc_52155_new_n19317_));
AND2X2 AND2X2_9629 ( .A(u2__abc_52155_new_n19318_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__21_));
AND2X2 AND2X2_963 ( .A(u2__abc_52155_new_n3943_), .B(u2__abc_52155_new_n3946_), .Y(u2__abc_52155_new_n3947_));
AND2X2 AND2X2_9630 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_21_), .Y(u2__abc_52155_new_n19320_));
AND2X2 AND2X2_9631 ( .A(u2__abc_52155_new_n19310_), .B(sqrto_20_), .Y(u2__abc_52155_new_n19322_));
AND2X2 AND2X2_9632 ( .A(u2__abc_52155_new_n19323_), .B(u2__abc_52155_new_n19321_), .Y(u2__abc_52155_new_n19324_));
AND2X2 AND2X2_9633 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3258_), .Y(u2__abc_52155_new_n19326_));
AND2X2 AND2X2_9634 ( .A(u2__abc_52155_new_n19327_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19328_));
AND2X2 AND2X2_9635 ( .A(u2__abc_52155_new_n19325_), .B(u2__abc_52155_new_n19328_), .Y(u2__abc_52155_new_n19329_));
AND2X2 AND2X2_9636 ( .A(u2__abc_52155_new_n19330_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__22_));
AND2X2 AND2X2_9637 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_22_), .Y(u2__abc_52155_new_n19332_));
AND2X2 AND2X2_9638 ( .A(u2__abc_52155_new_n19322_), .B(sqrto_21_), .Y(u2__abc_52155_new_n19334_));
AND2X2 AND2X2_9639 ( .A(u2__abc_52155_new_n19335_), .B(u2__abc_52155_new_n19333_), .Y(u2__abc_52155_new_n19336_));
AND2X2 AND2X2_964 ( .A(u2__abc_52155_new_n3948_), .B(u2_remHi_86_), .Y(u2__abc_52155_new_n3949_));
AND2X2 AND2X2_9640 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3186_), .Y(u2__abc_52155_new_n19338_));
AND2X2 AND2X2_9641 ( .A(u2__abc_52155_new_n19339_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19340_));
AND2X2 AND2X2_9642 ( .A(u2__abc_52155_new_n19337_), .B(u2__abc_52155_new_n19340_), .Y(u2__abc_52155_new_n19341_));
AND2X2 AND2X2_9643 ( .A(u2__abc_52155_new_n19342_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__23_));
AND2X2 AND2X2_9644 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_23_), .Y(u2__abc_52155_new_n19344_));
AND2X2 AND2X2_9645 ( .A(u2__abc_52155_new_n19334_), .B(sqrto_22_), .Y(u2__abc_52155_new_n19346_));
AND2X2 AND2X2_9646 ( .A(u2__abc_52155_new_n19347_), .B(u2__abc_52155_new_n19345_), .Y(u2__abc_52155_new_n19348_));
AND2X2 AND2X2_9647 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3179_), .Y(u2__abc_52155_new_n19350_));
AND2X2 AND2X2_9648 ( .A(u2__abc_52155_new_n19351_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19352_));
AND2X2 AND2X2_9649 ( .A(u2__abc_52155_new_n19349_), .B(u2__abc_52155_new_n19352_), .Y(u2__abc_52155_new_n19353_));
AND2X2 AND2X2_965 ( .A(u2__abc_52155_new_n3951_), .B(sqrto_86_), .Y(u2__abc_52155_new_n3952_));
AND2X2 AND2X2_9650 ( .A(u2__abc_52155_new_n19354_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__24_));
AND2X2 AND2X2_9651 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_24_), .Y(u2__abc_52155_new_n19356_));
AND2X2 AND2X2_9652 ( .A(u2__abc_52155_new_n19346_), .B(sqrto_23_), .Y(u2__abc_52155_new_n19358_));
AND2X2 AND2X2_9653 ( .A(u2__abc_52155_new_n19359_), .B(u2__abc_52155_new_n19357_), .Y(u2__abc_52155_new_n19360_));
AND2X2 AND2X2_9654 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3167_), .Y(u2__abc_52155_new_n19362_));
AND2X2 AND2X2_9655 ( .A(u2__abc_52155_new_n19363_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19364_));
AND2X2 AND2X2_9656 ( .A(u2__abc_52155_new_n19361_), .B(u2__abc_52155_new_n19364_), .Y(u2__abc_52155_new_n19365_));
AND2X2 AND2X2_9657 ( .A(u2__abc_52155_new_n19366_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__25_));
AND2X2 AND2X2_9658 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_25_), .Y(u2__abc_52155_new_n19368_));
AND2X2 AND2X2_9659 ( .A(u2__abc_52155_new_n19358_), .B(sqrto_24_), .Y(u2__abc_52155_new_n19370_));
AND2X2 AND2X2_966 ( .A(u2__abc_52155_new_n3950_), .B(u2__abc_52155_new_n3953_), .Y(u2__abc_52155_new_n3954_));
AND2X2 AND2X2_9660 ( .A(u2__abc_52155_new_n19371_), .B(u2__abc_52155_new_n19369_), .Y(u2__abc_52155_new_n19372_));
AND2X2 AND2X2_9661 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3172_), .Y(u2__abc_52155_new_n19374_));
AND2X2 AND2X2_9662 ( .A(u2__abc_52155_new_n19375_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19376_));
AND2X2 AND2X2_9663 ( .A(u2__abc_52155_new_n19373_), .B(u2__abc_52155_new_n19376_), .Y(u2__abc_52155_new_n19377_));
AND2X2 AND2X2_9664 ( .A(u2__abc_52155_new_n19378_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__26_));
AND2X2 AND2X2_9665 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_26_), .Y(u2__abc_52155_new_n19380_));
AND2X2 AND2X2_9666 ( .A(u2__abc_52155_new_n19370_), .B(sqrto_25_), .Y(u2__abc_52155_new_n19382_));
AND2X2 AND2X2_9667 ( .A(u2__abc_52155_new_n19383_), .B(u2__abc_52155_new_n19381_), .Y(u2__abc_52155_new_n19384_));
AND2X2 AND2X2_9668 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3217_), .Y(u2__abc_52155_new_n19386_));
AND2X2 AND2X2_9669 ( .A(u2__abc_52155_new_n19387_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19388_));
AND2X2 AND2X2_967 ( .A(u2__abc_52155_new_n3947_), .B(u2__abc_52155_new_n3954_), .Y(u2__abc_52155_new_n3955_));
AND2X2 AND2X2_9670 ( .A(u2__abc_52155_new_n19385_), .B(u2__abc_52155_new_n19388_), .Y(u2__abc_52155_new_n19389_));
AND2X2 AND2X2_9671 ( .A(u2__abc_52155_new_n19390_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__27_));
AND2X2 AND2X2_9672 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_27_), .Y(u2__abc_52155_new_n19392_));
AND2X2 AND2X2_9673 ( .A(u2__abc_52155_new_n19382_), .B(sqrto_26_), .Y(u2__abc_52155_new_n19394_));
AND2X2 AND2X2_9674 ( .A(u2__abc_52155_new_n19395_), .B(u2__abc_52155_new_n19393_), .Y(u2__abc_52155_new_n19396_));
AND2X2 AND2X2_9675 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3210_), .Y(u2__abc_52155_new_n19398_));
AND2X2 AND2X2_9676 ( .A(u2__abc_52155_new_n19399_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19400_));
AND2X2 AND2X2_9677 ( .A(u2__abc_52155_new_n19397_), .B(u2__abc_52155_new_n19400_), .Y(u2__abc_52155_new_n19401_));
AND2X2 AND2X2_9678 ( .A(u2__abc_52155_new_n19402_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__28_));
AND2X2 AND2X2_9679 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_28_), .Y(u2__abc_52155_new_n19404_));
AND2X2 AND2X2_968 ( .A(u2__abc_52155_new_n3940_), .B(u2__abc_52155_new_n3955_), .Y(u2__abc_52155_new_n3956_));
AND2X2 AND2X2_9680 ( .A(u2__abc_52155_new_n19394_), .B(sqrto_27_), .Y(u2__abc_52155_new_n19406_));
AND2X2 AND2X2_9681 ( .A(u2__abc_52155_new_n19407_), .B(u2__abc_52155_new_n19405_), .Y(u2__abc_52155_new_n19408_));
AND2X2 AND2X2_9682 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3195_), .Y(u2__abc_52155_new_n19410_));
AND2X2 AND2X2_9683 ( .A(u2__abc_52155_new_n19411_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19412_));
AND2X2 AND2X2_9684 ( .A(u2__abc_52155_new_n19409_), .B(u2__abc_52155_new_n19412_), .Y(u2__abc_52155_new_n19413_));
AND2X2 AND2X2_9685 ( .A(u2__abc_52155_new_n19414_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__29_));
AND2X2 AND2X2_9686 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_29_), .Y(u2__abc_52155_new_n19416_));
AND2X2 AND2X2_9687 ( .A(u2__abc_52155_new_n19406_), .B(sqrto_28_), .Y(u2__abc_52155_new_n19418_));
AND2X2 AND2X2_9688 ( .A(u2__abc_52155_new_n19419_), .B(u2__abc_52155_new_n19417_), .Y(u2__abc_52155_new_n19420_));
AND2X2 AND2X2_9689 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3205_), .Y(u2__abc_52155_new_n19422_));
AND2X2 AND2X2_969 ( .A(u2__abc_52155_new_n3925_), .B(u2__abc_52155_new_n3956_), .Y(u2__abc_52155_new_n3957_));
AND2X2 AND2X2_9690 ( .A(u2__abc_52155_new_n19423_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19424_));
AND2X2 AND2X2_9691 ( .A(u2__abc_52155_new_n19421_), .B(u2__abc_52155_new_n19424_), .Y(u2__abc_52155_new_n19425_));
AND2X2 AND2X2_9692 ( .A(u2__abc_52155_new_n19426_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__30_));
AND2X2 AND2X2_9693 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_30_), .Y(u2__abc_52155_new_n19428_));
AND2X2 AND2X2_9694 ( .A(u2__abc_52155_new_n19418_), .B(sqrto_29_), .Y(u2__abc_52155_new_n19430_));
AND2X2 AND2X2_9695 ( .A(u2__abc_52155_new_n19431_), .B(u2__abc_52155_new_n19429_), .Y(u2__abc_52155_new_n19432_));
AND2X2 AND2X2_9696 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3519_), .Y(u2__abc_52155_new_n19434_));
AND2X2 AND2X2_9697 ( .A(u2__abc_52155_new_n19435_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19436_));
AND2X2 AND2X2_9698 ( .A(u2__abc_52155_new_n19433_), .B(u2__abc_52155_new_n19436_), .Y(u2__abc_52155_new_n19437_));
AND2X2 AND2X2_9699 ( .A(u2__abc_52155_new_n19438_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__31_));
AND2X2 AND2X2_97 ( .A(_abc_73687_new_n891_), .B(_abc_73687_new_n890_), .Y(\o[132] ));
AND2X2 AND2X2_970 ( .A(u2__abc_52155_new_n3958_), .B(u2_remHi_78_), .Y(u2__abc_52155_new_n3959_));
AND2X2 AND2X2_9700 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_31_), .Y(u2__abc_52155_new_n19440_));
AND2X2 AND2X2_9701 ( .A(u2__abc_52155_new_n19430_), .B(sqrto_30_), .Y(u2__abc_52155_new_n19442_));
AND2X2 AND2X2_9702 ( .A(u2__abc_52155_new_n19443_), .B(u2__abc_52155_new_n19441_), .Y(u2__abc_52155_new_n19444_));
AND2X2 AND2X2_9703 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3524_), .Y(u2__abc_52155_new_n19446_));
AND2X2 AND2X2_9704 ( .A(u2__abc_52155_new_n19447_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19448_));
AND2X2 AND2X2_9705 ( .A(u2__abc_52155_new_n19445_), .B(u2__abc_52155_new_n19448_), .Y(u2__abc_52155_new_n19449_));
AND2X2 AND2X2_9706 ( .A(u2__abc_52155_new_n19450_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__32_));
AND2X2 AND2X2_9707 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_32_), .Y(u2__abc_52155_new_n19452_));
AND2X2 AND2X2_9708 ( .A(u2__abc_52155_new_n19442_), .B(sqrto_31_), .Y(u2__abc_52155_new_n19454_));
AND2X2 AND2X2_9709 ( .A(u2__abc_52155_new_n19455_), .B(u2__abc_52155_new_n19453_), .Y(u2__abc_52155_new_n19456_));
AND2X2 AND2X2_971 ( .A(u2__abc_52155_new_n3961_), .B(sqrto_78_), .Y(u2__abc_52155_new_n3962_));
AND2X2 AND2X2_9710 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3507_), .Y(u2__abc_52155_new_n19458_));
AND2X2 AND2X2_9711 ( .A(u2__abc_52155_new_n19459_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19460_));
AND2X2 AND2X2_9712 ( .A(u2__abc_52155_new_n19457_), .B(u2__abc_52155_new_n19460_), .Y(u2__abc_52155_new_n19461_));
AND2X2 AND2X2_9713 ( .A(u2__abc_52155_new_n19462_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__33_));
AND2X2 AND2X2_9714 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_33_), .Y(u2__abc_52155_new_n19464_));
AND2X2 AND2X2_9715 ( .A(u2__abc_52155_new_n19454_), .B(sqrto_32_), .Y(u2__abc_52155_new_n19466_));
AND2X2 AND2X2_9716 ( .A(u2__abc_52155_new_n19467_), .B(u2__abc_52155_new_n19465_), .Y(u2__abc_52155_new_n19468_));
AND2X2 AND2X2_9717 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3512_), .Y(u2__abc_52155_new_n19470_));
AND2X2 AND2X2_9718 ( .A(u2__abc_52155_new_n19471_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19472_));
AND2X2 AND2X2_9719 ( .A(u2__abc_52155_new_n19469_), .B(u2__abc_52155_new_n19472_), .Y(u2__abc_52155_new_n19473_));
AND2X2 AND2X2_972 ( .A(u2__abc_52155_new_n3960_), .B(u2__abc_52155_new_n3963_), .Y(u2__abc_52155_new_n3964_));
AND2X2 AND2X2_9720 ( .A(u2__abc_52155_new_n19474_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__34_));
AND2X2 AND2X2_9721 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_34_), .Y(u2__abc_52155_new_n19476_));
AND2X2 AND2X2_9722 ( .A(u2__abc_52155_new_n19466_), .B(sqrto_33_), .Y(u2__abc_52155_new_n19478_));
AND2X2 AND2X2_9723 ( .A(u2__abc_52155_new_n19479_), .B(u2__abc_52155_new_n19477_), .Y(u2__abc_52155_new_n19480_));
AND2X2 AND2X2_9724 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3549_), .Y(u2__abc_52155_new_n19482_));
AND2X2 AND2X2_9725 ( .A(u2__abc_52155_new_n19483_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19484_));
AND2X2 AND2X2_9726 ( .A(u2__abc_52155_new_n19481_), .B(u2__abc_52155_new_n19484_), .Y(u2__abc_52155_new_n19485_));
AND2X2 AND2X2_9727 ( .A(u2__abc_52155_new_n19486_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__35_));
AND2X2 AND2X2_9728 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_35_), .Y(u2__abc_52155_new_n19488_));
AND2X2 AND2X2_9729 ( .A(u2__abc_52155_new_n19478_), .B(sqrto_34_), .Y(u2__abc_52155_new_n19490_));
AND2X2 AND2X2_973 ( .A(u2__abc_52155_new_n3965_), .B(u2_remHi_79_), .Y(u2__abc_52155_new_n3966_));
AND2X2 AND2X2_9730 ( .A(u2__abc_52155_new_n19491_), .B(u2__abc_52155_new_n19489_), .Y(u2__abc_52155_new_n19492_));
AND2X2 AND2X2_9731 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3544_), .Y(u2__abc_52155_new_n19494_));
AND2X2 AND2X2_9732 ( .A(u2__abc_52155_new_n19495_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19496_));
AND2X2 AND2X2_9733 ( .A(u2__abc_52155_new_n19493_), .B(u2__abc_52155_new_n19496_), .Y(u2__abc_52155_new_n19497_));
AND2X2 AND2X2_9734 ( .A(u2__abc_52155_new_n19498_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__36_));
AND2X2 AND2X2_9735 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_36_), .Y(u2__abc_52155_new_n19500_));
AND2X2 AND2X2_9736 ( .A(u2__abc_52155_new_n19490_), .B(sqrto_35_), .Y(u2__abc_52155_new_n19502_));
AND2X2 AND2X2_9737 ( .A(u2__abc_52155_new_n19503_), .B(u2__abc_52155_new_n19501_), .Y(u2__abc_52155_new_n19504_));
AND2X2 AND2X2_9738 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3533_), .Y(u2__abc_52155_new_n19506_));
AND2X2 AND2X2_9739 ( .A(u2__abc_52155_new_n19507_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19508_));
AND2X2 AND2X2_974 ( .A(u2__abc_52155_new_n3968_), .B(sqrto_79_), .Y(u2__abc_52155_new_n3969_));
AND2X2 AND2X2_9740 ( .A(u2__abc_52155_new_n19505_), .B(u2__abc_52155_new_n19508_), .Y(u2__abc_52155_new_n19509_));
AND2X2 AND2X2_9741 ( .A(u2__abc_52155_new_n19510_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__37_));
AND2X2 AND2X2_9742 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_37_), .Y(u2__abc_52155_new_n19512_));
AND2X2 AND2X2_9743 ( .A(u2__abc_52155_new_n19502_), .B(sqrto_36_), .Y(u2__abc_52155_new_n19514_));
AND2X2 AND2X2_9744 ( .A(u2__abc_52155_new_n19515_), .B(u2__abc_52155_new_n19513_), .Y(u2__abc_52155_new_n19516_));
AND2X2 AND2X2_9745 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3538_), .Y(u2__abc_52155_new_n19518_));
AND2X2 AND2X2_9746 ( .A(u2__abc_52155_new_n19519_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19520_));
AND2X2 AND2X2_9747 ( .A(u2__abc_52155_new_n19517_), .B(u2__abc_52155_new_n19520_), .Y(u2__abc_52155_new_n19521_));
AND2X2 AND2X2_9748 ( .A(u2__abc_52155_new_n19522_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__38_));
AND2X2 AND2X2_9749 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_38_), .Y(u2__abc_52155_new_n19524_));
AND2X2 AND2X2_975 ( .A(u2__abc_52155_new_n3967_), .B(u2__abc_52155_new_n3970_), .Y(u2__abc_52155_new_n3971_));
AND2X2 AND2X2_9750 ( .A(u2__abc_52155_new_n19514_), .B(sqrto_37_), .Y(u2__abc_52155_new_n19526_));
AND2X2 AND2X2_9751 ( .A(u2__abc_52155_new_n19527_), .B(u2__abc_52155_new_n19525_), .Y(u2__abc_52155_new_n19528_));
AND2X2 AND2X2_9752 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3459_), .Y(u2__abc_52155_new_n19530_));
AND2X2 AND2X2_9753 ( .A(u2__abc_52155_new_n19531_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19532_));
AND2X2 AND2X2_9754 ( .A(u2__abc_52155_new_n19529_), .B(u2__abc_52155_new_n19532_), .Y(u2__abc_52155_new_n19533_));
AND2X2 AND2X2_9755 ( .A(u2__abc_52155_new_n19534_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__39_));
AND2X2 AND2X2_9756 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_39_), .Y(u2__abc_52155_new_n19536_));
AND2X2 AND2X2_9757 ( .A(u2__abc_52155_new_n19526_), .B(sqrto_38_), .Y(u2__abc_52155_new_n19538_));
AND2X2 AND2X2_9758 ( .A(u2__abc_52155_new_n19539_), .B(u2__abc_52155_new_n19537_), .Y(u2__abc_52155_new_n19540_));
AND2X2 AND2X2_9759 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3466_), .Y(u2__abc_52155_new_n19542_));
AND2X2 AND2X2_976 ( .A(u2__abc_52155_new_n3964_), .B(u2__abc_52155_new_n3971_), .Y(u2__abc_52155_new_n3972_));
AND2X2 AND2X2_9760 ( .A(u2__abc_52155_new_n19543_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19544_));
AND2X2 AND2X2_9761 ( .A(u2__abc_52155_new_n19541_), .B(u2__abc_52155_new_n19544_), .Y(u2__abc_52155_new_n19545_));
AND2X2 AND2X2_9762 ( .A(u2__abc_52155_new_n19546_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__40_));
AND2X2 AND2X2_9763 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_40_), .Y(u2__abc_52155_new_n19548_));
AND2X2 AND2X2_9764 ( .A(u2__abc_52155_new_n19538_), .B(sqrto_39_), .Y(u2__abc_52155_new_n19550_));
AND2X2 AND2X2_9765 ( .A(u2__abc_52155_new_n19551_), .B(u2__abc_52155_new_n19549_), .Y(u2__abc_52155_new_n19552_));
AND2X2 AND2X2_9766 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3447_), .Y(u2__abc_52155_new_n19554_));
AND2X2 AND2X2_9767 ( .A(u2__abc_52155_new_n19555_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19556_));
AND2X2 AND2X2_9768 ( .A(u2__abc_52155_new_n19553_), .B(u2__abc_52155_new_n19556_), .Y(u2__abc_52155_new_n19557_));
AND2X2 AND2X2_9769 ( .A(u2__abc_52155_new_n19558_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__41_));
AND2X2 AND2X2_977 ( .A(u2__abc_52155_new_n3973_), .B(u2_remHi_80_), .Y(u2__abc_52155_new_n3974_));
AND2X2 AND2X2_9770 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_41_), .Y(u2__abc_52155_new_n19560_));
AND2X2 AND2X2_9771 ( .A(u2__abc_52155_new_n19550_), .B(sqrto_40_), .Y(u2__abc_52155_new_n19562_));
AND2X2 AND2X2_9772 ( .A(u2__abc_52155_new_n19563_), .B(u2__abc_52155_new_n19561_), .Y(u2__abc_52155_new_n19564_));
AND2X2 AND2X2_9773 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3452_), .Y(u2__abc_52155_new_n19566_));
AND2X2 AND2X2_9774 ( .A(u2__abc_52155_new_n19567_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19568_));
AND2X2 AND2X2_9775 ( .A(u2__abc_52155_new_n19565_), .B(u2__abc_52155_new_n19568_), .Y(u2__abc_52155_new_n19569_));
AND2X2 AND2X2_9776 ( .A(u2__abc_52155_new_n19570_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__42_));
AND2X2 AND2X2_9777 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_42_), .Y(u2__abc_52155_new_n19572_));
AND2X2 AND2X2_9778 ( .A(u2__abc_52155_new_n19562_), .B(sqrto_41_), .Y(u2__abc_52155_new_n19574_));
AND2X2 AND2X2_9779 ( .A(u2__abc_52155_new_n19575_), .B(u2__abc_52155_new_n19573_), .Y(u2__abc_52155_new_n19576_));
AND2X2 AND2X2_978 ( .A(u2__abc_52155_new_n3975_), .B(sqrto_80_), .Y(u2__abc_52155_new_n3976_));
AND2X2 AND2X2_9780 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3497_), .Y(u2__abc_52155_new_n19578_));
AND2X2 AND2X2_9781 ( .A(u2__abc_52155_new_n19579_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19580_));
AND2X2 AND2X2_9782 ( .A(u2__abc_52155_new_n19577_), .B(u2__abc_52155_new_n19580_), .Y(u2__abc_52155_new_n19581_));
AND2X2 AND2X2_9783 ( .A(u2__abc_52155_new_n19582_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__43_));
AND2X2 AND2X2_9784 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_43_), .Y(u2__abc_52155_new_n19584_));
AND2X2 AND2X2_9785 ( .A(u2__abc_52155_new_n19574_), .B(sqrto_42_), .Y(u2__abc_52155_new_n19586_));
AND2X2 AND2X2_9786 ( .A(u2__abc_52155_new_n19587_), .B(u2__abc_52155_new_n19585_), .Y(u2__abc_52155_new_n19588_));
AND2X2 AND2X2_9787 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3490_), .Y(u2__abc_52155_new_n19590_));
AND2X2 AND2X2_9788 ( .A(u2__abc_52155_new_n19591_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19592_));
AND2X2 AND2X2_9789 ( .A(u2__abc_52155_new_n19589_), .B(u2__abc_52155_new_n19592_), .Y(u2__abc_52155_new_n19593_));
AND2X2 AND2X2_979 ( .A(u2__abc_52155_new_n3978_), .B(u2_remHi_81_), .Y(u2__abc_52155_new_n3979_));
AND2X2 AND2X2_9790 ( .A(u2__abc_52155_new_n19594_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__44_));
AND2X2 AND2X2_9791 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_44_), .Y(u2__abc_52155_new_n19596_));
AND2X2 AND2X2_9792 ( .A(u2__abc_52155_new_n19586_), .B(sqrto_43_), .Y(u2__abc_52155_new_n19598_));
AND2X2 AND2X2_9793 ( .A(u2__abc_52155_new_n19599_), .B(u2__abc_52155_new_n19597_), .Y(u2__abc_52155_new_n19600_));
AND2X2 AND2X2_9794 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3475_), .Y(u2__abc_52155_new_n19602_));
AND2X2 AND2X2_9795 ( .A(u2__abc_52155_new_n19603_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19604_));
AND2X2 AND2X2_9796 ( .A(u2__abc_52155_new_n19601_), .B(u2__abc_52155_new_n19604_), .Y(u2__abc_52155_new_n19605_));
AND2X2 AND2X2_9797 ( .A(u2__abc_52155_new_n19606_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__45_));
AND2X2 AND2X2_9798 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_45_), .Y(u2__abc_52155_new_n19608_));
AND2X2 AND2X2_9799 ( .A(u2__abc_52155_new_n19598_), .B(sqrto_44_), .Y(u2__abc_52155_new_n19610_));
AND2X2 AND2X2_98 ( .A(_abc_73687_new_n894_), .B(_abc_73687_new_n893_), .Y(\o[133] ));
AND2X2 AND2X2_980 ( .A(u2__abc_52155_new_n3980_), .B(sqrto_81_), .Y(u2__abc_52155_new_n3981_));
AND2X2 AND2X2_9800 ( .A(u2__abc_52155_new_n19611_), .B(u2__abc_52155_new_n19609_), .Y(u2__abc_52155_new_n19612_));
AND2X2 AND2X2_9801 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3482_), .Y(u2__abc_52155_new_n19614_));
AND2X2 AND2X2_9802 ( .A(u2__abc_52155_new_n19615_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19616_));
AND2X2 AND2X2_9803 ( .A(u2__abc_52155_new_n19613_), .B(u2__abc_52155_new_n19616_), .Y(u2__abc_52155_new_n19617_));
AND2X2 AND2X2_9804 ( .A(u2__abc_52155_new_n19618_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__46_));
AND2X2 AND2X2_9805 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_46_), .Y(u2__abc_52155_new_n19620_));
AND2X2 AND2X2_9806 ( .A(u2__abc_52155_new_n19610_), .B(sqrto_45_), .Y(u2__abc_52155_new_n19622_));
AND2X2 AND2X2_9807 ( .A(u2__abc_52155_new_n19623_), .B(u2__abc_52155_new_n19621_), .Y(u2__abc_52155_new_n19624_));
AND2X2 AND2X2_9808 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3405_), .Y(u2__abc_52155_new_n19626_));
AND2X2 AND2X2_9809 ( .A(u2__abc_52155_new_n19627_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19628_));
AND2X2 AND2X2_981 ( .A(u2__abc_52155_new_n3984_), .B(u2__abc_52155_new_n3972_), .Y(u2__abc_52155_new_n3985_));
AND2X2 AND2X2_9810 ( .A(u2__abc_52155_new_n19625_), .B(u2__abc_52155_new_n19628_), .Y(u2__abc_52155_new_n19629_));
AND2X2 AND2X2_9811 ( .A(u2__abc_52155_new_n19630_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__47_));
AND2X2 AND2X2_9812 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_47_), .Y(u2__abc_52155_new_n19632_));
AND2X2 AND2X2_9813 ( .A(u2__abc_52155_new_n19622_), .B(sqrto_46_), .Y(u2__abc_52155_new_n19634_));
AND2X2 AND2X2_9814 ( .A(u2__abc_52155_new_n19635_), .B(u2__abc_52155_new_n19633_), .Y(u2__abc_52155_new_n19636_));
AND2X2 AND2X2_9815 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3398_), .Y(u2__abc_52155_new_n19638_));
AND2X2 AND2X2_9816 ( .A(u2__abc_52155_new_n19639_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19640_));
AND2X2 AND2X2_9817 ( .A(u2__abc_52155_new_n19637_), .B(u2__abc_52155_new_n19640_), .Y(u2__abc_52155_new_n19641_));
AND2X2 AND2X2_9818 ( .A(u2__abc_52155_new_n19642_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__48_));
AND2X2 AND2X2_9819 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_48_), .Y(u2__abc_52155_new_n19644_));
AND2X2 AND2X2_982 ( .A(u2__abc_52155_new_n3986_), .B(u2_remHi_84_), .Y(u2__abc_52155_new_n3987_));
AND2X2 AND2X2_9820 ( .A(u2__abc_52155_new_n19634_), .B(sqrto_47_), .Y(u2__abc_52155_new_n19646_));
AND2X2 AND2X2_9821 ( .A(u2__abc_52155_new_n19647_), .B(u2__abc_52155_new_n19645_), .Y(u2__abc_52155_new_n19648_));
AND2X2 AND2X2_9822 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3386_), .Y(u2__abc_52155_new_n19650_));
AND2X2 AND2X2_9823 ( .A(u2__abc_52155_new_n19651_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19652_));
AND2X2 AND2X2_9824 ( .A(u2__abc_52155_new_n19649_), .B(u2__abc_52155_new_n19652_), .Y(u2__abc_52155_new_n19653_));
AND2X2 AND2X2_9825 ( .A(u2__abc_52155_new_n19654_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__49_));
AND2X2 AND2X2_9826 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_49_), .Y(u2__abc_52155_new_n19656_));
AND2X2 AND2X2_9827 ( .A(u2__abc_52155_new_n19646_), .B(sqrto_48_), .Y(u2__abc_52155_new_n19658_));
AND2X2 AND2X2_9828 ( .A(u2__abc_52155_new_n19659_), .B(u2__abc_52155_new_n19657_), .Y(u2__abc_52155_new_n19660_));
AND2X2 AND2X2_9829 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3391_), .Y(u2__abc_52155_new_n19662_));
AND2X2 AND2X2_983 ( .A(u2__abc_52155_new_n3989_), .B(sqrto_84_), .Y(u2__abc_52155_new_n3990_));
AND2X2 AND2X2_9830 ( .A(u2__abc_52155_new_n19663_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19664_));
AND2X2 AND2X2_9831 ( .A(u2__abc_52155_new_n19661_), .B(u2__abc_52155_new_n19664_), .Y(u2__abc_52155_new_n19665_));
AND2X2 AND2X2_9832 ( .A(u2__abc_52155_new_n19666_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__50_));
AND2X2 AND2X2_9833 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_50_), .Y(u2__abc_52155_new_n19668_));
AND2X2 AND2X2_9834 ( .A(u2__abc_52155_new_n19658_), .B(sqrto_49_), .Y(u2__abc_52155_new_n19670_));
AND2X2 AND2X2_9835 ( .A(u2__abc_52155_new_n19671_), .B(u2__abc_52155_new_n19669_), .Y(u2__abc_52155_new_n19672_));
AND2X2 AND2X2_9836 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3436_), .Y(u2__abc_52155_new_n19674_));
AND2X2 AND2X2_9837 ( .A(u2__abc_52155_new_n19675_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19676_));
AND2X2 AND2X2_9838 ( .A(u2__abc_52155_new_n19673_), .B(u2__abc_52155_new_n19676_), .Y(u2__abc_52155_new_n19677_));
AND2X2 AND2X2_9839 ( .A(u2__abc_52155_new_n19678_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__51_));
AND2X2 AND2X2_984 ( .A(u2__abc_52155_new_n3988_), .B(u2__abc_52155_new_n3991_), .Y(u2__abc_52155_new_n3992_));
AND2X2 AND2X2_9840 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_51_), .Y(u2__abc_52155_new_n19680_));
AND2X2 AND2X2_9841 ( .A(u2__abc_52155_new_n19670_), .B(sqrto_50_), .Y(u2__abc_52155_new_n19682_));
AND2X2 AND2X2_9842 ( .A(u2__abc_52155_new_n19683_), .B(u2__abc_52155_new_n19681_), .Y(u2__abc_52155_new_n19684_));
AND2X2 AND2X2_9843 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3429_), .Y(u2__abc_52155_new_n19686_));
AND2X2 AND2X2_9844 ( .A(u2__abc_52155_new_n19687_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19688_));
AND2X2 AND2X2_9845 ( .A(u2__abc_52155_new_n19685_), .B(u2__abc_52155_new_n19688_), .Y(u2__abc_52155_new_n19689_));
AND2X2 AND2X2_9846 ( .A(u2__abc_52155_new_n19690_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__52_));
AND2X2 AND2X2_9847 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_52_), .Y(u2__abc_52155_new_n19692_));
AND2X2 AND2X2_9848 ( .A(u2__abc_52155_new_n19682_), .B(sqrto_51_), .Y(u2__abc_52155_new_n19694_));
AND2X2 AND2X2_9849 ( .A(u2__abc_52155_new_n19695_), .B(u2__abc_52155_new_n19693_), .Y(u2__abc_52155_new_n19696_));
AND2X2 AND2X2_985 ( .A(u2__abc_52155_new_n3993_), .B(u2_remHi_85_), .Y(u2__abc_52155_new_n3994_));
AND2X2 AND2X2_9850 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3414_), .Y(u2__abc_52155_new_n19698_));
AND2X2 AND2X2_9851 ( .A(u2__abc_52155_new_n19699_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19700_));
AND2X2 AND2X2_9852 ( .A(u2__abc_52155_new_n19697_), .B(u2__abc_52155_new_n19700_), .Y(u2__abc_52155_new_n19701_));
AND2X2 AND2X2_9853 ( .A(u2__abc_52155_new_n19702_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__53_));
AND2X2 AND2X2_9854 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_53_), .Y(u2__abc_52155_new_n19704_));
AND2X2 AND2X2_9855 ( .A(u2__abc_52155_new_n19694_), .B(sqrto_52_), .Y(u2__abc_52155_new_n19706_));
AND2X2 AND2X2_9856 ( .A(u2__abc_52155_new_n19707_), .B(u2__abc_52155_new_n19705_), .Y(u2__abc_52155_new_n19708_));
AND2X2 AND2X2_9857 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3421_), .Y(u2__abc_52155_new_n19710_));
AND2X2 AND2X2_9858 ( .A(u2__abc_52155_new_n19711_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19712_));
AND2X2 AND2X2_9859 ( .A(u2__abc_52155_new_n19709_), .B(u2__abc_52155_new_n19712_), .Y(u2__abc_52155_new_n19713_));
AND2X2 AND2X2_986 ( .A(u2__abc_52155_new_n3996_), .B(sqrto_85_), .Y(u2__abc_52155_new_n3997_));
AND2X2 AND2X2_9860 ( .A(u2__abc_52155_new_n19714_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__54_));
AND2X2 AND2X2_9861 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_54_), .Y(u2__abc_52155_new_n19716_));
AND2X2 AND2X2_9862 ( .A(u2__abc_52155_new_n19706_), .B(sqrto_53_), .Y(u2__abc_52155_new_n19718_));
AND2X2 AND2X2_9863 ( .A(u2__abc_52155_new_n19719_), .B(u2__abc_52155_new_n19717_), .Y(u2__abc_52155_new_n19720_));
AND2X2 AND2X2_9864 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3338_), .Y(u2__abc_52155_new_n19722_));
AND2X2 AND2X2_9865 ( .A(u2__abc_52155_new_n19723_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19724_));
AND2X2 AND2X2_9866 ( .A(u2__abc_52155_new_n19721_), .B(u2__abc_52155_new_n19724_), .Y(u2__abc_52155_new_n19725_));
AND2X2 AND2X2_9867 ( .A(u2__abc_52155_new_n19726_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__55_));
AND2X2 AND2X2_9868 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_55_), .Y(u2__abc_52155_new_n19728_));
AND2X2 AND2X2_9869 ( .A(u2__abc_52155_new_n19718_), .B(sqrto_54_), .Y(u2__abc_52155_new_n19730_));
AND2X2 AND2X2_987 ( .A(u2__abc_52155_new_n3995_), .B(u2__abc_52155_new_n3998_), .Y(u2__abc_52155_new_n3999_));
AND2X2 AND2X2_9870 ( .A(u2__abc_52155_new_n19731_), .B(u2__abc_52155_new_n19729_), .Y(u2__abc_52155_new_n19732_));
AND2X2 AND2X2_9871 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3345_), .Y(u2__abc_52155_new_n19734_));
AND2X2 AND2X2_9872 ( .A(u2__abc_52155_new_n19735_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19736_));
AND2X2 AND2X2_9873 ( .A(u2__abc_52155_new_n19733_), .B(u2__abc_52155_new_n19736_), .Y(u2__abc_52155_new_n19737_));
AND2X2 AND2X2_9874 ( .A(u2__abc_52155_new_n19738_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__56_));
AND2X2 AND2X2_9875 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_56_), .Y(u2__abc_52155_new_n19740_));
AND2X2 AND2X2_9876 ( .A(u2__abc_52155_new_n19730_), .B(sqrto_55_), .Y(u2__abc_52155_new_n19742_));
AND2X2 AND2X2_9877 ( .A(u2__abc_52155_new_n19743_), .B(u2__abc_52155_new_n19741_), .Y(u2__abc_52155_new_n19744_));
AND2X2 AND2X2_9878 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3323_), .Y(u2__abc_52155_new_n19746_));
AND2X2 AND2X2_9879 ( .A(u2__abc_52155_new_n19747_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19748_));
AND2X2 AND2X2_988 ( .A(u2__abc_52155_new_n3992_), .B(u2__abc_52155_new_n3999_), .Y(u2__abc_52155_new_n4000_));
AND2X2 AND2X2_9880 ( .A(u2__abc_52155_new_n19745_), .B(u2__abc_52155_new_n19748_), .Y(u2__abc_52155_new_n19749_));
AND2X2 AND2X2_9881 ( .A(u2__abc_52155_new_n19750_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__57_));
AND2X2 AND2X2_9882 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_57_), .Y(u2__abc_52155_new_n19752_));
AND2X2 AND2X2_9883 ( .A(u2__abc_52155_new_n19742_), .B(sqrto_56_), .Y(u2__abc_52155_new_n19754_));
AND2X2 AND2X2_9884 ( .A(u2__abc_52155_new_n19755_), .B(u2__abc_52155_new_n19753_), .Y(u2__abc_52155_new_n19756_));
AND2X2 AND2X2_9885 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3330_), .Y(u2__abc_52155_new_n19758_));
AND2X2 AND2X2_9886 ( .A(u2__abc_52155_new_n19759_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19760_));
AND2X2 AND2X2_9887 ( .A(u2__abc_52155_new_n19757_), .B(u2__abc_52155_new_n19760_), .Y(u2__abc_52155_new_n19761_));
AND2X2 AND2X2_9888 ( .A(u2__abc_52155_new_n19762_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__58_));
AND2X2 AND2X2_9889 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_58_), .Y(u2__abc_52155_new_n19764_));
AND2X2 AND2X2_989 ( .A(u2__abc_52155_new_n4001_), .B(u2_remHi_83_), .Y(u2__abc_52155_new_n4002_));
AND2X2 AND2X2_9890 ( .A(u2__abc_52155_new_n19754_), .B(sqrto_57_), .Y(u2__abc_52155_new_n19766_));
AND2X2 AND2X2_9891 ( .A(u2__abc_52155_new_n19767_), .B(u2__abc_52155_new_n19765_), .Y(u2__abc_52155_new_n19768_));
AND2X2 AND2X2_9892 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3376_), .Y(u2__abc_52155_new_n19770_));
AND2X2 AND2X2_9893 ( .A(u2__abc_52155_new_n19771_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19772_));
AND2X2 AND2X2_9894 ( .A(u2__abc_52155_new_n19769_), .B(u2__abc_52155_new_n19772_), .Y(u2__abc_52155_new_n19773_));
AND2X2 AND2X2_9895 ( .A(u2__abc_52155_new_n19774_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__59_));
AND2X2 AND2X2_9896 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_59_), .Y(u2__abc_52155_new_n19776_));
AND2X2 AND2X2_9897 ( .A(u2__abc_52155_new_n19766_), .B(sqrto_58_), .Y(u2__abc_52155_new_n19778_));
AND2X2 AND2X2_9898 ( .A(u2__abc_52155_new_n19779_), .B(u2__abc_52155_new_n19777_), .Y(u2__abc_52155_new_n19780_));
AND2X2 AND2X2_9899 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3369_), .Y(u2__abc_52155_new_n19782_));
AND2X2 AND2X2_99 ( .A(_abc_73687_new_n897_), .B(_abc_73687_new_n896_), .Y(\o[134] ));
AND2X2 AND2X2_990 ( .A(u2__abc_52155_new_n4004_), .B(sqrto_83_), .Y(u2__abc_52155_new_n4005_));
AND2X2 AND2X2_9900 ( .A(u2__abc_52155_new_n19783_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19784_));
AND2X2 AND2X2_9901 ( .A(u2__abc_52155_new_n19781_), .B(u2__abc_52155_new_n19784_), .Y(u2__abc_52155_new_n19785_));
AND2X2 AND2X2_9902 ( .A(u2__abc_52155_new_n19786_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__60_));
AND2X2 AND2X2_9903 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_60_), .Y(u2__abc_52155_new_n19788_));
AND2X2 AND2X2_9904 ( .A(u2__abc_52155_new_n19778_), .B(sqrto_59_), .Y(u2__abc_52155_new_n19790_));
AND2X2 AND2X2_9905 ( .A(u2__abc_52155_new_n19791_), .B(u2__abc_52155_new_n19789_), .Y(u2__abc_52155_new_n19792_));
AND2X2 AND2X2_9906 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3354_), .Y(u2__abc_52155_new_n19794_));
AND2X2 AND2X2_9907 ( .A(u2__abc_52155_new_n19795_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19796_));
AND2X2 AND2X2_9908 ( .A(u2__abc_52155_new_n19793_), .B(u2__abc_52155_new_n19796_), .Y(u2__abc_52155_new_n19797_));
AND2X2 AND2X2_9909 ( .A(u2__abc_52155_new_n19798_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__61_));
AND2X2 AND2X2_991 ( .A(u2__abc_52155_new_n4003_), .B(u2__abc_52155_new_n4006_), .Y(u2__abc_52155_new_n4007_));
AND2X2 AND2X2_9910 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_61_), .Y(u2__abc_52155_new_n19800_));
AND2X2 AND2X2_9911 ( .A(u2__abc_52155_new_n19790_), .B(sqrto_60_), .Y(u2__abc_52155_new_n19802_));
AND2X2 AND2X2_9912 ( .A(u2__abc_52155_new_n19803_), .B(u2__abc_52155_new_n19801_), .Y(u2__abc_52155_new_n19804_));
AND2X2 AND2X2_9913 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n3364_), .Y(u2__abc_52155_new_n19806_));
AND2X2 AND2X2_9914 ( .A(u2__abc_52155_new_n19807_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19808_));
AND2X2 AND2X2_9915 ( .A(u2__abc_52155_new_n19805_), .B(u2__abc_52155_new_n19808_), .Y(u2__abc_52155_new_n19809_));
AND2X2 AND2X2_9916 ( .A(u2__abc_52155_new_n19810_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__62_));
AND2X2 AND2X2_9917 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_62_), .Y(u2__abc_52155_new_n19812_));
AND2X2 AND2X2_9918 ( .A(u2__abc_52155_new_n19802_), .B(sqrto_61_), .Y(u2__abc_52155_new_n19814_));
AND2X2 AND2X2_9919 ( .A(u2__abc_52155_new_n19815_), .B(u2__abc_52155_new_n19813_), .Y(u2__abc_52155_new_n19816_));
AND2X2 AND2X2_992 ( .A(u2__abc_52155_new_n4008_), .B(u2_remHi_82_), .Y(u2__abc_52155_new_n4009_));
AND2X2 AND2X2_9920 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4079_), .Y(u2__abc_52155_new_n19818_));
AND2X2 AND2X2_9921 ( .A(u2__abc_52155_new_n19819_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19820_));
AND2X2 AND2X2_9922 ( .A(u2__abc_52155_new_n19817_), .B(u2__abc_52155_new_n19820_), .Y(u2__abc_52155_new_n19821_));
AND2X2 AND2X2_9923 ( .A(u2__abc_52155_new_n19822_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__63_));
AND2X2 AND2X2_9924 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_63_), .Y(u2__abc_52155_new_n19824_));
AND2X2 AND2X2_9925 ( .A(u2__abc_52155_new_n19814_), .B(sqrto_62_), .Y(u2__abc_52155_new_n19826_));
AND2X2 AND2X2_9926 ( .A(u2__abc_52155_new_n19827_), .B(u2__abc_52155_new_n19825_), .Y(u2__abc_52155_new_n19828_));
AND2X2 AND2X2_9927 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4084_), .Y(u2__abc_52155_new_n19830_));
AND2X2 AND2X2_9928 ( .A(u2__abc_52155_new_n19831_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19832_));
AND2X2 AND2X2_9929 ( .A(u2__abc_52155_new_n19829_), .B(u2__abc_52155_new_n19832_), .Y(u2__abc_52155_new_n19833_));
AND2X2 AND2X2_993 ( .A(u2__abc_52155_new_n4011_), .B(sqrto_82_), .Y(u2__abc_52155_new_n4012_));
AND2X2 AND2X2_9930 ( .A(u2__abc_52155_new_n19834_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__64_));
AND2X2 AND2X2_9931 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_64_), .Y(u2__abc_52155_new_n19836_));
AND2X2 AND2X2_9932 ( .A(u2__abc_52155_new_n19826_), .B(sqrto_63_), .Y(u2__abc_52155_new_n19838_));
AND2X2 AND2X2_9933 ( .A(u2__abc_52155_new_n19839_), .B(u2__abc_52155_new_n19837_), .Y(u2__abc_52155_new_n19840_));
AND2X2 AND2X2_9934 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4092_), .Y(u2__abc_52155_new_n19842_));
AND2X2 AND2X2_9935 ( .A(u2__abc_52155_new_n19843_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19844_));
AND2X2 AND2X2_9936 ( .A(u2__abc_52155_new_n19841_), .B(u2__abc_52155_new_n19844_), .Y(u2__abc_52155_new_n19845_));
AND2X2 AND2X2_9937 ( .A(u2__abc_52155_new_n19846_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__65_));
AND2X2 AND2X2_9938 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_65_), .Y(u2__abc_52155_new_n19848_));
AND2X2 AND2X2_9939 ( .A(u2__abc_52155_new_n19838_), .B(sqrto_64_), .Y(u2__abc_52155_new_n19850_));
AND2X2 AND2X2_994 ( .A(u2__abc_52155_new_n4010_), .B(u2__abc_52155_new_n4013_), .Y(u2__abc_52155_new_n4014_));
AND2X2 AND2X2_9940 ( .A(u2__abc_52155_new_n19851_), .B(u2__abc_52155_new_n19849_), .Y(u2__abc_52155_new_n19852_));
AND2X2 AND2X2_9941 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4097_), .Y(u2__abc_52155_new_n19854_));
AND2X2 AND2X2_9942 ( .A(u2__abc_52155_new_n19855_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19856_));
AND2X2 AND2X2_9943 ( .A(u2__abc_52155_new_n19853_), .B(u2__abc_52155_new_n19856_), .Y(u2__abc_52155_new_n19857_));
AND2X2 AND2X2_9944 ( .A(u2__abc_52155_new_n19858_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__66_));
AND2X2 AND2X2_9945 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_66_), .Y(u2__abc_52155_new_n19860_));
AND2X2 AND2X2_9946 ( .A(u2__abc_52155_new_n19850_), .B(sqrto_65_), .Y(u2__abc_52155_new_n19862_));
AND2X2 AND2X2_9947 ( .A(u2__abc_52155_new_n19863_), .B(u2__abc_52155_new_n19861_), .Y(u2__abc_52155_new_n19864_));
AND2X2 AND2X2_9948 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4121_), .Y(u2__abc_52155_new_n19866_));
AND2X2 AND2X2_9949 ( .A(u2__abc_52155_new_n19867_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19868_));
AND2X2 AND2X2_995 ( .A(u2__abc_52155_new_n4007_), .B(u2__abc_52155_new_n4014_), .Y(u2__abc_52155_new_n4015_));
AND2X2 AND2X2_9950 ( .A(u2__abc_52155_new_n19865_), .B(u2__abc_52155_new_n19868_), .Y(u2__abc_52155_new_n19869_));
AND2X2 AND2X2_9951 ( .A(u2__abc_52155_new_n19870_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__67_));
AND2X2 AND2X2_9952 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_67_), .Y(u2__abc_52155_new_n19872_));
AND2X2 AND2X2_9953 ( .A(u2__abc_52155_new_n19862_), .B(sqrto_66_), .Y(u2__abc_52155_new_n19874_));
AND2X2 AND2X2_9954 ( .A(u2__abc_52155_new_n19875_), .B(u2__abc_52155_new_n19873_), .Y(u2__abc_52155_new_n19876_));
AND2X2 AND2X2_9955 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4116_), .Y(u2__abc_52155_new_n19878_));
AND2X2 AND2X2_9956 ( .A(u2__abc_52155_new_n19879_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19880_));
AND2X2 AND2X2_9957 ( .A(u2__abc_52155_new_n19877_), .B(u2__abc_52155_new_n19880_), .Y(u2__abc_52155_new_n19881_));
AND2X2 AND2X2_9958 ( .A(u2__abc_52155_new_n19882_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__68_));
AND2X2 AND2X2_9959 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_68_), .Y(u2__abc_52155_new_n19884_));
AND2X2 AND2X2_996 ( .A(u2__abc_52155_new_n4000_), .B(u2__abc_52155_new_n4015_), .Y(u2__abc_52155_new_n4016_));
AND2X2 AND2X2_9960 ( .A(u2__abc_52155_new_n19874_), .B(sqrto_67_), .Y(u2__abc_52155_new_n19886_));
AND2X2 AND2X2_9961 ( .A(u2__abc_52155_new_n19887_), .B(u2__abc_52155_new_n19885_), .Y(u2__abc_52155_new_n19888_));
AND2X2 AND2X2_9962 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4105_), .Y(u2__abc_52155_new_n19890_));
AND2X2 AND2X2_9963 ( .A(u2__abc_52155_new_n19891_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19892_));
AND2X2 AND2X2_9964 ( .A(u2__abc_52155_new_n19889_), .B(u2__abc_52155_new_n19892_), .Y(u2__abc_52155_new_n19893_));
AND2X2 AND2X2_9965 ( .A(u2__abc_52155_new_n19894_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__69_));
AND2X2 AND2X2_9966 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_69_), .Y(u2__abc_52155_new_n19896_));
AND2X2 AND2X2_9967 ( .A(u2__abc_52155_new_n19886_), .B(sqrto_68_), .Y(u2__abc_52155_new_n19898_));
AND2X2 AND2X2_9968 ( .A(u2__abc_52155_new_n19899_), .B(u2__abc_52155_new_n19897_), .Y(u2__abc_52155_new_n19900_));
AND2X2 AND2X2_9969 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4110_), .Y(u2__abc_52155_new_n19902_));
AND2X2 AND2X2_997 ( .A(u2__abc_52155_new_n3985_), .B(u2__abc_52155_new_n4016_), .Y(u2__abc_52155_new_n4017_));
AND2X2 AND2X2_9970 ( .A(u2__abc_52155_new_n19903_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19904_));
AND2X2 AND2X2_9971 ( .A(u2__abc_52155_new_n19901_), .B(u2__abc_52155_new_n19904_), .Y(u2__abc_52155_new_n19905_));
AND2X2 AND2X2_9972 ( .A(u2__abc_52155_new_n19906_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__70_));
AND2X2 AND2X2_9973 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_70_), .Y(u2__abc_52155_new_n19908_));
AND2X2 AND2X2_9974 ( .A(u2__abc_52155_new_n19898_), .B(sqrto_69_), .Y(u2__abc_52155_new_n19910_));
AND2X2 AND2X2_9975 ( .A(u2__abc_52155_new_n19911_), .B(u2__abc_52155_new_n19909_), .Y(u2__abc_52155_new_n19912_));
AND2X2 AND2X2_9976 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4019_), .Y(u2__abc_52155_new_n19914_));
AND2X2 AND2X2_9977 ( .A(u2__abc_52155_new_n19915_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19916_));
AND2X2 AND2X2_9978 ( .A(u2__abc_52155_new_n19913_), .B(u2__abc_52155_new_n19916_), .Y(u2__abc_52155_new_n19917_));
AND2X2 AND2X2_9979 ( .A(u2__abc_52155_new_n19918_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__71_));
AND2X2 AND2X2_998 ( .A(u2__abc_52155_new_n4017_), .B(u2__abc_52155_new_n3957_), .Y(u2__abc_52155_new_n4018_));
AND2X2 AND2X2_9980 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_71_), .Y(u2__abc_52155_new_n19920_));
AND2X2 AND2X2_9981 ( .A(u2__abc_52155_new_n19910_), .B(sqrto_70_), .Y(u2__abc_52155_new_n19922_));
AND2X2 AND2X2_9982 ( .A(u2__abc_52155_new_n19923_), .B(u2__abc_52155_new_n19921_), .Y(u2__abc_52155_new_n19924_));
AND2X2 AND2X2_9983 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4026_), .Y(u2__abc_52155_new_n19926_));
AND2X2 AND2X2_9984 ( .A(u2__abc_52155_new_n19927_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19928_));
AND2X2 AND2X2_9985 ( .A(u2__abc_52155_new_n19925_), .B(u2__abc_52155_new_n19928_), .Y(u2__abc_52155_new_n19929_));
AND2X2 AND2X2_9986 ( .A(u2__abc_52155_new_n19930_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__72_));
AND2X2 AND2X2_9987 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_72_), .Y(u2__abc_52155_new_n19932_));
AND2X2 AND2X2_9988 ( .A(u2__abc_52155_new_n19922_), .B(sqrto_71_), .Y(u2__abc_52155_new_n19934_));
AND2X2 AND2X2_9989 ( .A(u2__abc_52155_new_n19935_), .B(u2__abc_52155_new_n19933_), .Y(u2__abc_52155_new_n19936_));
AND2X2 AND2X2_999 ( .A(u2__abc_52155_new_n4019_), .B(u2_remHi_70_), .Y(u2__abc_52155_new_n4020_));
AND2X2 AND2X2_9990 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4034_), .Y(u2__abc_52155_new_n19938_));
AND2X2 AND2X2_9991 ( .A(u2__abc_52155_new_n19939_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19940_));
AND2X2 AND2X2_9992 ( .A(u2__abc_52155_new_n19937_), .B(u2__abc_52155_new_n19940_), .Y(u2__abc_52155_new_n19941_));
AND2X2 AND2X2_9993 ( .A(u2__abc_52155_new_n19942_), .B(u2__abc_52155_new_n2962_), .Y(u2__0root_452_0__73_));
AND2X2 AND2X2_9994 ( .A(u2__abc_52155_new_n3002_), .B(sqrto_73_), .Y(u2__abc_52155_new_n19944_));
AND2X2 AND2X2_9995 ( .A(u2__abc_52155_new_n19934_), .B(sqrto_72_), .Y(u2__abc_52155_new_n19946_));
AND2X2 AND2X2_9996 ( .A(u2__abc_52155_new_n19947_), .B(u2__abc_52155_new_n19945_), .Y(u2__abc_52155_new_n19948_));
AND2X2 AND2X2_9997 ( .A(u2__abc_52155_new_n2974_), .B(u2__abc_52155_new_n4039_), .Y(u2__abc_52155_new_n19950_));
AND2X2 AND2X2_9998 ( .A(u2__abc_52155_new_n19951_), .B(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n19952_));
AND2X2 AND2X2_9999 ( .A(u2__abc_52155_new_n19949_), .B(u2__abc_52155_new_n19952_), .Y(u2__abc_52155_new_n19953_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_0_), .Q(u2_state_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(u2__0root_452_0__6_), .Q(sqrto_5_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk), .D(u2__0root_452_0__96_), .Q(sqrto_95_));
DFFPOSX1 DFFPOSX1_1000 ( .CLK(clk), .D(u2__0remHi_451_0__93_), .Q(u2_remHi_93_));
DFFPOSX1 DFFPOSX1_1001 ( .CLK(clk), .D(u2__0remHi_451_0__94_), .Q(u2_remHi_94_));
DFFPOSX1 DFFPOSX1_1002 ( .CLK(clk), .D(u2__0remHi_451_0__95_), .Q(u2_remHi_95_));
DFFPOSX1 DFFPOSX1_1003 ( .CLK(clk), .D(u2__0remHi_451_0__96_), .Q(u2_remHi_96_));
DFFPOSX1 DFFPOSX1_1004 ( .CLK(clk), .D(u2__0remHi_451_0__97_), .Q(u2_remHi_97_));
DFFPOSX1 DFFPOSX1_1005 ( .CLK(clk), .D(u2__0remHi_451_0__98_), .Q(u2_remHi_98_));
DFFPOSX1 DFFPOSX1_1006 ( .CLK(clk), .D(u2__0remHi_451_0__99_), .Q(u2_remHi_99_));
DFFPOSX1 DFFPOSX1_1007 ( .CLK(clk), .D(u2__0remHi_451_0__100_), .Q(u2_remHi_100_));
DFFPOSX1 DFFPOSX1_1008 ( .CLK(clk), .D(u2__0remHi_451_0__101_), .Q(u2_remHi_101_));
DFFPOSX1 DFFPOSX1_1009 ( .CLK(clk), .D(u2__0remHi_451_0__102_), .Q(u2_remHi_102_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk), .D(u2__0root_452_0__97_), .Q(sqrto_96_));
DFFPOSX1 DFFPOSX1_1010 ( .CLK(clk), .D(u2__0remHi_451_0__103_), .Q(u2_remHi_103_));
DFFPOSX1 DFFPOSX1_1011 ( .CLK(clk), .D(u2__0remHi_451_0__104_), .Q(u2_remHi_104_));
DFFPOSX1 DFFPOSX1_1012 ( .CLK(clk), .D(u2__0remHi_451_0__105_), .Q(u2_remHi_105_));
DFFPOSX1 DFFPOSX1_1013 ( .CLK(clk), .D(u2__0remHi_451_0__106_), .Q(u2_remHi_106_));
DFFPOSX1 DFFPOSX1_1014 ( .CLK(clk), .D(u2__0remHi_451_0__107_), .Q(u2_remHi_107_));
DFFPOSX1 DFFPOSX1_1015 ( .CLK(clk), .D(u2__0remHi_451_0__108_), .Q(u2_remHi_108_));
DFFPOSX1 DFFPOSX1_1016 ( .CLK(clk), .D(u2__0remHi_451_0__109_), .Q(u2_remHi_109_));
DFFPOSX1 DFFPOSX1_1017 ( .CLK(clk), .D(u2__0remHi_451_0__110_), .Q(u2_remHi_110_));
DFFPOSX1 DFFPOSX1_1018 ( .CLK(clk), .D(u2__0remHi_451_0__111_), .Q(u2_remHi_111_));
DFFPOSX1 DFFPOSX1_1019 ( .CLK(clk), .D(u2__0remHi_451_0__112_), .Q(u2_remHi_112_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk), .D(u2__0root_452_0__98_), .Q(sqrto_97_));
DFFPOSX1 DFFPOSX1_1020 ( .CLK(clk), .D(u2__0remHi_451_0__113_), .Q(u2_remHi_113_));
DFFPOSX1 DFFPOSX1_1021 ( .CLK(clk), .D(u2__0remHi_451_0__114_), .Q(u2_remHi_114_));
DFFPOSX1 DFFPOSX1_1022 ( .CLK(clk), .D(u2__0remHi_451_0__115_), .Q(u2_remHi_115_));
DFFPOSX1 DFFPOSX1_1023 ( .CLK(clk), .D(u2__0remHi_451_0__116_), .Q(u2_remHi_116_));
DFFPOSX1 DFFPOSX1_1024 ( .CLK(clk), .D(u2__0remHi_451_0__117_), .Q(u2_remHi_117_));
DFFPOSX1 DFFPOSX1_1025 ( .CLK(clk), .D(u2__0remHi_451_0__118_), .Q(u2_remHi_118_));
DFFPOSX1 DFFPOSX1_1026 ( .CLK(clk), .D(u2__0remHi_451_0__119_), .Q(u2_remHi_119_));
DFFPOSX1 DFFPOSX1_1027 ( .CLK(clk), .D(u2__0remHi_451_0__120_), .Q(u2_remHi_120_));
DFFPOSX1 DFFPOSX1_1028 ( .CLK(clk), .D(u2__0remHi_451_0__121_), .Q(u2_remHi_121_));
DFFPOSX1 DFFPOSX1_1029 ( .CLK(clk), .D(u2__0remHi_451_0__122_), .Q(u2_remHi_122_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk), .D(u2__0root_452_0__99_), .Q(sqrto_98_));
DFFPOSX1 DFFPOSX1_1030 ( .CLK(clk), .D(u2__0remHi_451_0__123_), .Q(u2_remHi_123_));
DFFPOSX1 DFFPOSX1_1031 ( .CLK(clk), .D(u2__0remHi_451_0__124_), .Q(u2_remHi_124_));
DFFPOSX1 DFFPOSX1_1032 ( .CLK(clk), .D(u2__0remHi_451_0__125_), .Q(u2_remHi_125_));
DFFPOSX1 DFFPOSX1_1033 ( .CLK(clk), .D(u2__0remHi_451_0__126_), .Q(u2_remHi_126_));
DFFPOSX1 DFFPOSX1_1034 ( .CLK(clk), .D(u2__0remHi_451_0__127_), .Q(u2_remHi_127_));
DFFPOSX1 DFFPOSX1_1035 ( .CLK(clk), .D(u2__0remHi_451_0__128_), .Q(u2_remHi_128_));
DFFPOSX1 DFFPOSX1_1036 ( .CLK(clk), .D(u2__0remHi_451_0__129_), .Q(u2_remHi_129_));
DFFPOSX1 DFFPOSX1_1037 ( .CLK(clk), .D(u2__0remHi_451_0__130_), .Q(u2_remHi_130_));
DFFPOSX1 DFFPOSX1_1038 ( .CLK(clk), .D(u2__0remHi_451_0__131_), .Q(u2_remHi_131_));
DFFPOSX1 DFFPOSX1_1039 ( .CLK(clk), .D(u2__0remHi_451_0__132_), .Q(u2_remHi_132_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk), .D(u2__0root_452_0__100_), .Q(sqrto_99_));
DFFPOSX1 DFFPOSX1_1040 ( .CLK(clk), .D(u2__0remHi_451_0__133_), .Q(u2_remHi_133_));
DFFPOSX1 DFFPOSX1_1041 ( .CLK(clk), .D(u2__0remHi_451_0__134_), .Q(u2_remHi_134_));
DFFPOSX1 DFFPOSX1_1042 ( .CLK(clk), .D(u2__0remHi_451_0__135_), .Q(u2_remHi_135_));
DFFPOSX1 DFFPOSX1_1043 ( .CLK(clk), .D(u2__0remHi_451_0__136_), .Q(u2_remHi_136_));
DFFPOSX1 DFFPOSX1_1044 ( .CLK(clk), .D(u2__0remHi_451_0__137_), .Q(u2_remHi_137_));
DFFPOSX1 DFFPOSX1_1045 ( .CLK(clk), .D(u2__0remHi_451_0__138_), .Q(u2_remHi_138_));
DFFPOSX1 DFFPOSX1_1046 ( .CLK(clk), .D(u2__0remHi_451_0__139_), .Q(u2_remHi_139_));
DFFPOSX1 DFFPOSX1_1047 ( .CLK(clk), .D(u2__0remHi_451_0__140_), .Q(u2_remHi_140_));
DFFPOSX1 DFFPOSX1_1048 ( .CLK(clk), .D(u2__0remHi_451_0__141_), .Q(u2_remHi_141_));
DFFPOSX1 DFFPOSX1_1049 ( .CLK(clk), .D(u2__0remHi_451_0__142_), .Q(u2_remHi_142_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk), .D(u2__0root_452_0__101_), .Q(sqrto_100_));
DFFPOSX1 DFFPOSX1_1050 ( .CLK(clk), .D(u2__0remHi_451_0__143_), .Q(u2_remHi_143_));
DFFPOSX1 DFFPOSX1_1051 ( .CLK(clk), .D(u2__0remHi_451_0__144_), .Q(u2_remHi_144_));
DFFPOSX1 DFFPOSX1_1052 ( .CLK(clk), .D(u2__0remHi_451_0__145_), .Q(u2_remHi_145_));
DFFPOSX1 DFFPOSX1_1053 ( .CLK(clk), .D(u2__0remHi_451_0__146_), .Q(u2_remHi_146_));
DFFPOSX1 DFFPOSX1_1054 ( .CLK(clk), .D(u2__0remHi_451_0__147_), .Q(u2_remHi_147_));
DFFPOSX1 DFFPOSX1_1055 ( .CLK(clk), .D(u2__0remHi_451_0__148_), .Q(u2_remHi_148_));
DFFPOSX1 DFFPOSX1_1056 ( .CLK(clk), .D(u2__0remHi_451_0__149_), .Q(u2_remHi_149_));
DFFPOSX1 DFFPOSX1_1057 ( .CLK(clk), .D(u2__0remHi_451_0__150_), .Q(u2_remHi_150_));
DFFPOSX1 DFFPOSX1_1058 ( .CLK(clk), .D(u2__0remHi_451_0__151_), .Q(u2_remHi_151_));
DFFPOSX1 DFFPOSX1_1059 ( .CLK(clk), .D(u2__0remHi_451_0__152_), .Q(u2_remHi_152_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk), .D(u2__0root_452_0__102_), .Q(sqrto_101_));
DFFPOSX1 DFFPOSX1_1060 ( .CLK(clk), .D(u2__0remHi_451_0__153_), .Q(u2_remHi_153_));
DFFPOSX1 DFFPOSX1_1061 ( .CLK(clk), .D(u2__0remHi_451_0__154_), .Q(u2_remHi_154_));
DFFPOSX1 DFFPOSX1_1062 ( .CLK(clk), .D(u2__0remHi_451_0__155_), .Q(u2_remHi_155_));
DFFPOSX1 DFFPOSX1_1063 ( .CLK(clk), .D(u2__0remHi_451_0__156_), .Q(u2_remHi_156_));
DFFPOSX1 DFFPOSX1_1064 ( .CLK(clk), .D(u2__0remHi_451_0__157_), .Q(u2_remHi_157_));
DFFPOSX1 DFFPOSX1_1065 ( .CLK(clk), .D(u2__0remHi_451_0__158_), .Q(u2_remHi_158_));
DFFPOSX1 DFFPOSX1_1066 ( .CLK(clk), .D(u2__0remHi_451_0__159_), .Q(u2_remHi_159_));
DFFPOSX1 DFFPOSX1_1067 ( .CLK(clk), .D(u2__0remHi_451_0__160_), .Q(u2_remHi_160_));
DFFPOSX1 DFFPOSX1_1068 ( .CLK(clk), .D(u2__0remHi_451_0__161_), .Q(u2_remHi_161_));
DFFPOSX1 DFFPOSX1_1069 ( .CLK(clk), .D(u2__0remHi_451_0__162_), .Q(u2_remHi_162_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk), .D(u2__0root_452_0__103_), .Q(sqrto_102_));
DFFPOSX1 DFFPOSX1_1070 ( .CLK(clk), .D(u2__0remHi_451_0__163_), .Q(u2_remHi_163_));
DFFPOSX1 DFFPOSX1_1071 ( .CLK(clk), .D(u2__0remHi_451_0__164_), .Q(u2_remHi_164_));
DFFPOSX1 DFFPOSX1_1072 ( .CLK(clk), .D(u2__0remHi_451_0__165_), .Q(u2_remHi_165_));
DFFPOSX1 DFFPOSX1_1073 ( .CLK(clk), .D(u2__0remHi_451_0__166_), .Q(u2_remHi_166_));
DFFPOSX1 DFFPOSX1_1074 ( .CLK(clk), .D(u2__0remHi_451_0__167_), .Q(u2_remHi_167_));
DFFPOSX1 DFFPOSX1_1075 ( .CLK(clk), .D(u2__0remHi_451_0__168_), .Q(u2_remHi_168_));
DFFPOSX1 DFFPOSX1_1076 ( .CLK(clk), .D(u2__0remHi_451_0__169_), .Q(u2_remHi_169_));
DFFPOSX1 DFFPOSX1_1077 ( .CLK(clk), .D(u2__0remHi_451_0__170_), .Q(u2_remHi_170_));
DFFPOSX1 DFFPOSX1_1078 ( .CLK(clk), .D(u2__0remHi_451_0__171_), .Q(u2_remHi_171_));
DFFPOSX1 DFFPOSX1_1079 ( .CLK(clk), .D(u2__0remHi_451_0__172_), .Q(u2_remHi_172_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk), .D(u2__0root_452_0__104_), .Q(sqrto_103_));
DFFPOSX1 DFFPOSX1_1080 ( .CLK(clk), .D(u2__0remHi_451_0__173_), .Q(u2_remHi_173_));
DFFPOSX1 DFFPOSX1_1081 ( .CLK(clk), .D(u2__0remHi_451_0__174_), .Q(u2_remHi_174_));
DFFPOSX1 DFFPOSX1_1082 ( .CLK(clk), .D(u2__0remHi_451_0__175_), .Q(u2_remHi_175_));
DFFPOSX1 DFFPOSX1_1083 ( .CLK(clk), .D(u2__0remHi_451_0__176_), .Q(u2_remHi_176_));
DFFPOSX1 DFFPOSX1_1084 ( .CLK(clk), .D(u2__0remHi_451_0__177_), .Q(u2_remHi_177_));
DFFPOSX1 DFFPOSX1_1085 ( .CLK(clk), .D(u2__0remHi_451_0__178_), .Q(u2_remHi_178_));
DFFPOSX1 DFFPOSX1_1086 ( .CLK(clk), .D(u2__0remHi_451_0__179_), .Q(u2_remHi_179_));
DFFPOSX1 DFFPOSX1_1087 ( .CLK(clk), .D(u2__0remHi_451_0__180_), .Q(u2_remHi_180_));
DFFPOSX1 DFFPOSX1_1088 ( .CLK(clk), .D(u2__0remHi_451_0__181_), .Q(u2_remHi_181_));
DFFPOSX1 DFFPOSX1_1089 ( .CLK(clk), .D(u2__0remHi_451_0__182_), .Q(u2_remHi_182_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk), .D(u2__0root_452_0__105_), .Q(sqrto_104_));
DFFPOSX1 DFFPOSX1_1090 ( .CLK(clk), .D(u2__0remHi_451_0__183_), .Q(u2_remHi_183_));
DFFPOSX1 DFFPOSX1_1091 ( .CLK(clk), .D(u2__0remHi_451_0__184_), .Q(u2_remHi_184_));
DFFPOSX1 DFFPOSX1_1092 ( .CLK(clk), .D(u2__0remHi_451_0__185_), .Q(u2_remHi_185_));
DFFPOSX1 DFFPOSX1_1093 ( .CLK(clk), .D(u2__0remHi_451_0__186_), .Q(u2_remHi_186_));
DFFPOSX1 DFFPOSX1_1094 ( .CLK(clk), .D(u2__0remHi_451_0__187_), .Q(u2_remHi_187_));
DFFPOSX1 DFFPOSX1_1095 ( .CLK(clk), .D(u2__0remHi_451_0__188_), .Q(u2_remHi_188_));
DFFPOSX1 DFFPOSX1_1096 ( .CLK(clk), .D(u2__0remHi_451_0__189_), .Q(u2_remHi_189_));
DFFPOSX1 DFFPOSX1_1097 ( .CLK(clk), .D(u2__0remHi_451_0__190_), .Q(u2_remHi_190_));
DFFPOSX1 DFFPOSX1_1098 ( .CLK(clk), .D(u2__0remHi_451_0__191_), .Q(u2_remHi_191_));
DFFPOSX1 DFFPOSX1_1099 ( .CLK(clk), .D(u2__0remHi_451_0__192_), .Q(u2_remHi_192_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(u2__0root_452_0__7_), .Q(sqrto_6_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk), .D(u2__0root_452_0__106_), .Q(sqrto_105_));
DFFPOSX1 DFFPOSX1_1100 ( .CLK(clk), .D(u2__0remHi_451_0__193_), .Q(u2_remHi_193_));
DFFPOSX1 DFFPOSX1_1101 ( .CLK(clk), .D(u2__0remHi_451_0__194_), .Q(u2_remHi_194_));
DFFPOSX1 DFFPOSX1_1102 ( .CLK(clk), .D(u2__0remHi_451_0__195_), .Q(u2_remHi_195_));
DFFPOSX1 DFFPOSX1_1103 ( .CLK(clk), .D(u2__0remHi_451_0__196_), .Q(u2_remHi_196_));
DFFPOSX1 DFFPOSX1_1104 ( .CLK(clk), .D(u2__0remHi_451_0__197_), .Q(u2_remHi_197_));
DFFPOSX1 DFFPOSX1_1105 ( .CLK(clk), .D(u2__0remHi_451_0__198_), .Q(u2_remHi_198_));
DFFPOSX1 DFFPOSX1_1106 ( .CLK(clk), .D(u2__0remHi_451_0__199_), .Q(u2_remHi_199_));
DFFPOSX1 DFFPOSX1_1107 ( .CLK(clk), .D(u2__0remHi_451_0__200_), .Q(u2_remHi_200_));
DFFPOSX1 DFFPOSX1_1108 ( .CLK(clk), .D(u2__0remHi_451_0__201_), .Q(u2_remHi_201_));
DFFPOSX1 DFFPOSX1_1109 ( .CLK(clk), .D(u2__0remHi_451_0__202_), .Q(u2_remHi_202_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk), .D(u2__0root_452_0__107_), .Q(sqrto_106_));
DFFPOSX1 DFFPOSX1_1110 ( .CLK(clk), .D(u2__0remHi_451_0__203_), .Q(u2_remHi_203_));
DFFPOSX1 DFFPOSX1_1111 ( .CLK(clk), .D(u2__0remHi_451_0__204_), .Q(u2_remHi_204_));
DFFPOSX1 DFFPOSX1_1112 ( .CLK(clk), .D(u2__0remHi_451_0__205_), .Q(u2_remHi_205_));
DFFPOSX1 DFFPOSX1_1113 ( .CLK(clk), .D(u2__0remHi_451_0__206_), .Q(u2_remHi_206_));
DFFPOSX1 DFFPOSX1_1114 ( .CLK(clk), .D(u2__0remHi_451_0__207_), .Q(u2_remHi_207_));
DFFPOSX1 DFFPOSX1_1115 ( .CLK(clk), .D(u2__0remHi_451_0__208_), .Q(u2_remHi_208_));
DFFPOSX1 DFFPOSX1_1116 ( .CLK(clk), .D(u2__0remHi_451_0__209_), .Q(u2_remHi_209_));
DFFPOSX1 DFFPOSX1_1117 ( .CLK(clk), .D(u2__0remHi_451_0__210_), .Q(u2_remHi_210_));
DFFPOSX1 DFFPOSX1_1118 ( .CLK(clk), .D(u2__0remHi_451_0__211_), .Q(u2_remHi_211_));
DFFPOSX1 DFFPOSX1_1119 ( .CLK(clk), .D(u2__0remHi_451_0__212_), .Q(u2_remHi_212_));
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk), .D(u2__0root_452_0__108_), .Q(sqrto_107_));
DFFPOSX1 DFFPOSX1_1120 ( .CLK(clk), .D(u2__0remHi_451_0__213_), .Q(u2_remHi_213_));
DFFPOSX1 DFFPOSX1_1121 ( .CLK(clk), .D(u2__0remHi_451_0__214_), .Q(u2_remHi_214_));
DFFPOSX1 DFFPOSX1_1122 ( .CLK(clk), .D(u2__0remHi_451_0__215_), .Q(u2_remHi_215_));
DFFPOSX1 DFFPOSX1_1123 ( .CLK(clk), .D(u2__0remHi_451_0__216_), .Q(u2_remHi_216_));
DFFPOSX1 DFFPOSX1_1124 ( .CLK(clk), .D(u2__0remHi_451_0__217_), .Q(u2_remHi_217_));
DFFPOSX1 DFFPOSX1_1125 ( .CLK(clk), .D(u2__0remHi_451_0__218_), .Q(u2_remHi_218_));
DFFPOSX1 DFFPOSX1_1126 ( .CLK(clk), .D(u2__0remHi_451_0__219_), .Q(u2_remHi_219_));
DFFPOSX1 DFFPOSX1_1127 ( .CLK(clk), .D(u2__0remHi_451_0__220_), .Q(u2_remHi_220_));
DFFPOSX1 DFFPOSX1_1128 ( .CLK(clk), .D(u2__0remHi_451_0__221_), .Q(u2_remHi_221_));
DFFPOSX1 DFFPOSX1_1129 ( .CLK(clk), .D(u2__0remHi_451_0__222_), .Q(u2_remHi_222_));
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk), .D(u2__0root_452_0__109_), .Q(sqrto_108_));
DFFPOSX1 DFFPOSX1_1130 ( .CLK(clk), .D(u2__0remHi_451_0__223_), .Q(u2_remHi_223_));
DFFPOSX1 DFFPOSX1_1131 ( .CLK(clk), .D(u2__0remHi_451_0__224_), .Q(u2_remHi_224_));
DFFPOSX1 DFFPOSX1_1132 ( .CLK(clk), .D(u2__0remHi_451_0__225_), .Q(u2_remHi_225_));
DFFPOSX1 DFFPOSX1_1133 ( .CLK(clk), .D(u2__0remHi_451_0__226_), .Q(u2_remHi_226_));
DFFPOSX1 DFFPOSX1_1134 ( .CLK(clk), .D(u2__0remHi_451_0__227_), .Q(u2_remHi_227_));
DFFPOSX1 DFFPOSX1_1135 ( .CLK(clk), .D(u2__0remHi_451_0__228_), .Q(u2_remHi_228_));
DFFPOSX1 DFFPOSX1_1136 ( .CLK(clk), .D(u2__0remHi_451_0__229_), .Q(u2_remHi_229_));
DFFPOSX1 DFFPOSX1_1137 ( .CLK(clk), .D(u2__0remHi_451_0__230_), .Q(u2_remHi_230_));
DFFPOSX1 DFFPOSX1_1138 ( .CLK(clk), .D(u2__0remHi_451_0__231_), .Q(u2_remHi_231_));
DFFPOSX1 DFFPOSX1_1139 ( .CLK(clk), .D(u2__0remHi_451_0__232_), .Q(u2_remHi_232_));
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk), .D(u2__0root_452_0__110_), .Q(sqrto_109_));
DFFPOSX1 DFFPOSX1_1140 ( .CLK(clk), .D(u2__0remHi_451_0__233_), .Q(u2_remHi_233_));
DFFPOSX1 DFFPOSX1_1141 ( .CLK(clk), .D(u2__0remHi_451_0__234_), .Q(u2_remHi_234_));
DFFPOSX1 DFFPOSX1_1142 ( .CLK(clk), .D(u2__0remHi_451_0__235_), .Q(u2_remHi_235_));
DFFPOSX1 DFFPOSX1_1143 ( .CLK(clk), .D(u2__0remHi_451_0__236_), .Q(u2_remHi_236_));
DFFPOSX1 DFFPOSX1_1144 ( .CLK(clk), .D(u2__0remHi_451_0__237_), .Q(u2_remHi_237_));
DFFPOSX1 DFFPOSX1_1145 ( .CLK(clk), .D(u2__0remHi_451_0__238_), .Q(u2_remHi_238_));
DFFPOSX1 DFFPOSX1_1146 ( .CLK(clk), .D(u2__0remHi_451_0__239_), .Q(u2_remHi_239_));
DFFPOSX1 DFFPOSX1_1147 ( .CLK(clk), .D(u2__0remHi_451_0__240_), .Q(u2_remHi_240_));
DFFPOSX1 DFFPOSX1_1148 ( .CLK(clk), .D(u2__0remHi_451_0__241_), .Q(u2_remHi_241_));
DFFPOSX1 DFFPOSX1_1149 ( .CLK(clk), .D(u2__0remHi_451_0__242_), .Q(u2_remHi_242_));
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk), .D(u2__0root_452_0__111_), .Q(sqrto_110_));
DFFPOSX1 DFFPOSX1_1150 ( .CLK(clk), .D(u2__0remHi_451_0__243_), .Q(u2_remHi_243_));
DFFPOSX1 DFFPOSX1_1151 ( .CLK(clk), .D(u2__0remHi_451_0__244_), .Q(u2_remHi_244_));
DFFPOSX1 DFFPOSX1_1152 ( .CLK(clk), .D(u2__0remHi_451_0__245_), .Q(u2_remHi_245_));
DFFPOSX1 DFFPOSX1_1153 ( .CLK(clk), .D(u2__0remHi_451_0__246_), .Q(u2_remHi_246_));
DFFPOSX1 DFFPOSX1_1154 ( .CLK(clk), .D(u2__0remHi_451_0__247_), .Q(u2_remHi_247_));
DFFPOSX1 DFFPOSX1_1155 ( .CLK(clk), .D(u2__0remHi_451_0__248_), .Q(u2_remHi_248_));
DFFPOSX1 DFFPOSX1_1156 ( .CLK(clk), .D(u2__0remHi_451_0__249_), .Q(u2_remHi_249_));
DFFPOSX1 DFFPOSX1_1157 ( .CLK(clk), .D(u2__0remHi_451_0__250_), .Q(u2_remHi_250_));
DFFPOSX1 DFFPOSX1_1158 ( .CLK(clk), .D(u2__0remHi_451_0__251_), .Q(u2_remHi_251_));
DFFPOSX1 DFFPOSX1_1159 ( .CLK(clk), .D(u2__0remHi_451_0__252_), .Q(u2_remHi_252_));
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk), .D(u2__0root_452_0__112_), .Q(sqrto_111_));
DFFPOSX1 DFFPOSX1_1160 ( .CLK(clk), .D(u2__0remHi_451_0__253_), .Q(u2_remHi_253_));
DFFPOSX1 DFFPOSX1_1161 ( .CLK(clk), .D(u2__0remHi_451_0__254_), .Q(u2_remHi_254_));
DFFPOSX1 DFFPOSX1_1162 ( .CLK(clk), .D(u2__0remHi_451_0__255_), .Q(u2_remHi_255_));
DFFPOSX1 DFFPOSX1_1163 ( .CLK(clk), .D(u2__0remHi_451_0__256_), .Q(u2_remHi_256_));
DFFPOSX1 DFFPOSX1_1164 ( .CLK(clk), .D(u2__0remHi_451_0__257_), .Q(u2_remHi_257_));
DFFPOSX1 DFFPOSX1_1165 ( .CLK(clk), .D(u2__0remHi_451_0__258_), .Q(u2_remHi_258_));
DFFPOSX1 DFFPOSX1_1166 ( .CLK(clk), .D(u2__0remHi_451_0__259_), .Q(u2_remHi_259_));
DFFPOSX1 DFFPOSX1_1167 ( .CLK(clk), .D(u2__0remHi_451_0__260_), .Q(u2_remHi_260_));
DFFPOSX1 DFFPOSX1_1168 ( .CLK(clk), .D(u2__0remHi_451_0__261_), .Q(u2_remHi_261_));
DFFPOSX1 DFFPOSX1_1169 ( .CLK(clk), .D(u2__0remHi_451_0__262_), .Q(u2_remHi_262_));
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk), .D(u2__0root_452_0__113_), .Q(sqrto_112_));
DFFPOSX1 DFFPOSX1_1170 ( .CLK(clk), .D(u2__0remHi_451_0__263_), .Q(u2_remHi_263_));
DFFPOSX1 DFFPOSX1_1171 ( .CLK(clk), .D(u2__0remHi_451_0__264_), .Q(u2_remHi_264_));
DFFPOSX1 DFFPOSX1_1172 ( .CLK(clk), .D(u2__0remHi_451_0__265_), .Q(u2_remHi_265_));
DFFPOSX1 DFFPOSX1_1173 ( .CLK(clk), .D(u2__0remHi_451_0__266_), .Q(u2_remHi_266_));
DFFPOSX1 DFFPOSX1_1174 ( .CLK(clk), .D(u2__0remHi_451_0__267_), .Q(u2_remHi_267_));
DFFPOSX1 DFFPOSX1_1175 ( .CLK(clk), .D(u2__0remHi_451_0__268_), .Q(u2_remHi_268_));
DFFPOSX1 DFFPOSX1_1176 ( .CLK(clk), .D(u2__0remHi_451_0__269_), .Q(u2_remHi_269_));
DFFPOSX1 DFFPOSX1_1177 ( .CLK(clk), .D(u2__0remHi_451_0__270_), .Q(u2_remHi_270_));
DFFPOSX1 DFFPOSX1_1178 ( .CLK(clk), .D(u2__0remHi_451_0__271_), .Q(u2_remHi_271_));
DFFPOSX1 DFFPOSX1_1179 ( .CLK(clk), .D(u2__0remHi_451_0__272_), .Q(u2_remHi_272_));
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk), .D(u2__0root_452_0__114_), .Q(sqrto_113_));
DFFPOSX1 DFFPOSX1_1180 ( .CLK(clk), .D(u2__0remHi_451_0__273_), .Q(u2_remHi_273_));
DFFPOSX1 DFFPOSX1_1181 ( .CLK(clk), .D(u2__0remHi_451_0__274_), .Q(u2_remHi_274_));
DFFPOSX1 DFFPOSX1_1182 ( .CLK(clk), .D(u2__0remHi_451_0__275_), .Q(u2_remHi_275_));
DFFPOSX1 DFFPOSX1_1183 ( .CLK(clk), .D(u2__0remHi_451_0__276_), .Q(u2_remHi_276_));
DFFPOSX1 DFFPOSX1_1184 ( .CLK(clk), .D(u2__0remHi_451_0__277_), .Q(u2_remHi_277_));
DFFPOSX1 DFFPOSX1_1185 ( .CLK(clk), .D(u2__0remHi_451_0__278_), .Q(u2_remHi_278_));
DFFPOSX1 DFFPOSX1_1186 ( .CLK(clk), .D(u2__0remHi_451_0__279_), .Q(u2_remHi_279_));
DFFPOSX1 DFFPOSX1_1187 ( .CLK(clk), .D(u2__0remHi_451_0__280_), .Q(u2_remHi_280_));
DFFPOSX1 DFFPOSX1_1188 ( .CLK(clk), .D(u2__0remHi_451_0__281_), .Q(u2_remHi_281_));
DFFPOSX1 DFFPOSX1_1189 ( .CLK(clk), .D(u2__0remHi_451_0__282_), .Q(u2_remHi_282_));
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk), .D(u2__0root_452_0__115_), .Q(sqrto_114_));
DFFPOSX1 DFFPOSX1_1190 ( .CLK(clk), .D(u2__0remHi_451_0__283_), .Q(u2_remHi_283_));
DFFPOSX1 DFFPOSX1_1191 ( .CLK(clk), .D(u2__0remHi_451_0__284_), .Q(u2_remHi_284_));
DFFPOSX1 DFFPOSX1_1192 ( .CLK(clk), .D(u2__0remHi_451_0__285_), .Q(u2_remHi_285_));
DFFPOSX1 DFFPOSX1_1193 ( .CLK(clk), .D(u2__0remHi_451_0__286_), .Q(u2_remHi_286_));
DFFPOSX1 DFFPOSX1_1194 ( .CLK(clk), .D(u2__0remHi_451_0__287_), .Q(u2_remHi_287_));
DFFPOSX1 DFFPOSX1_1195 ( .CLK(clk), .D(u2__0remHi_451_0__288_), .Q(u2_remHi_288_));
DFFPOSX1 DFFPOSX1_1196 ( .CLK(clk), .D(u2__0remHi_451_0__289_), .Q(u2_remHi_289_));
DFFPOSX1 DFFPOSX1_1197 ( .CLK(clk), .D(u2__0remHi_451_0__290_), .Q(u2_remHi_290_));
DFFPOSX1 DFFPOSX1_1198 ( .CLK(clk), .D(u2__0remHi_451_0__291_), .Q(u2_remHi_291_));
DFFPOSX1 DFFPOSX1_1199 ( .CLK(clk), .D(u2__0remHi_451_0__292_), .Q(u2_remHi_292_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(u2__0root_452_0__8_), .Q(sqrto_7_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk), .D(u2__0root_452_0__116_), .Q(sqrto_115_));
DFFPOSX1 DFFPOSX1_1200 ( .CLK(clk), .D(u2__0remHi_451_0__293_), .Q(u2_remHi_293_));
DFFPOSX1 DFFPOSX1_1201 ( .CLK(clk), .D(u2__0remHi_451_0__294_), .Q(u2_remHi_294_));
DFFPOSX1 DFFPOSX1_1202 ( .CLK(clk), .D(u2__0remHi_451_0__295_), .Q(u2_remHi_295_));
DFFPOSX1 DFFPOSX1_1203 ( .CLK(clk), .D(u2__0remHi_451_0__296_), .Q(u2_remHi_296_));
DFFPOSX1 DFFPOSX1_1204 ( .CLK(clk), .D(u2__0remHi_451_0__297_), .Q(u2_remHi_297_));
DFFPOSX1 DFFPOSX1_1205 ( .CLK(clk), .D(u2__0remHi_451_0__298_), .Q(u2_remHi_298_));
DFFPOSX1 DFFPOSX1_1206 ( .CLK(clk), .D(u2__0remHi_451_0__299_), .Q(u2_remHi_299_));
DFFPOSX1 DFFPOSX1_1207 ( .CLK(clk), .D(u2__0remHi_451_0__300_), .Q(u2_remHi_300_));
DFFPOSX1 DFFPOSX1_1208 ( .CLK(clk), .D(u2__0remHi_451_0__301_), .Q(u2_remHi_301_));
DFFPOSX1 DFFPOSX1_1209 ( .CLK(clk), .D(u2__0remHi_451_0__302_), .Q(u2_remHi_302_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk), .D(u2__0root_452_0__117_), .Q(sqrto_116_));
DFFPOSX1 DFFPOSX1_1210 ( .CLK(clk), .D(u2__0remHi_451_0__303_), .Q(u2_remHi_303_));
DFFPOSX1 DFFPOSX1_1211 ( .CLK(clk), .D(u2__0remHi_451_0__304_), .Q(u2_remHi_304_));
DFFPOSX1 DFFPOSX1_1212 ( .CLK(clk), .D(u2__0remHi_451_0__305_), .Q(u2_remHi_305_));
DFFPOSX1 DFFPOSX1_1213 ( .CLK(clk), .D(u2__0remHi_451_0__306_), .Q(u2_remHi_306_));
DFFPOSX1 DFFPOSX1_1214 ( .CLK(clk), .D(u2__0remHi_451_0__307_), .Q(u2_remHi_307_));
DFFPOSX1 DFFPOSX1_1215 ( .CLK(clk), .D(u2__0remHi_451_0__308_), .Q(u2_remHi_308_));
DFFPOSX1 DFFPOSX1_1216 ( .CLK(clk), .D(u2__0remHi_451_0__309_), .Q(u2_remHi_309_));
DFFPOSX1 DFFPOSX1_1217 ( .CLK(clk), .D(u2__0remHi_451_0__310_), .Q(u2_remHi_310_));
DFFPOSX1 DFFPOSX1_1218 ( .CLK(clk), .D(u2__0remHi_451_0__311_), .Q(u2_remHi_311_));
DFFPOSX1 DFFPOSX1_1219 ( .CLK(clk), .D(u2__0remHi_451_0__312_), .Q(u2_remHi_312_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk), .D(u2__0root_452_0__118_), .Q(sqrto_117_));
DFFPOSX1 DFFPOSX1_1220 ( .CLK(clk), .D(u2__0remHi_451_0__313_), .Q(u2_remHi_313_));
DFFPOSX1 DFFPOSX1_1221 ( .CLK(clk), .D(u2__0remHi_451_0__314_), .Q(u2_remHi_314_));
DFFPOSX1 DFFPOSX1_1222 ( .CLK(clk), .D(u2__0remHi_451_0__315_), .Q(u2_remHi_315_));
DFFPOSX1 DFFPOSX1_1223 ( .CLK(clk), .D(u2__0remHi_451_0__316_), .Q(u2_remHi_316_));
DFFPOSX1 DFFPOSX1_1224 ( .CLK(clk), .D(u2__0remHi_451_0__317_), .Q(u2_remHi_317_));
DFFPOSX1 DFFPOSX1_1225 ( .CLK(clk), .D(u2__0remHi_451_0__318_), .Q(u2_remHi_318_));
DFFPOSX1 DFFPOSX1_1226 ( .CLK(clk), .D(u2__0remHi_451_0__319_), .Q(u2_remHi_319_));
DFFPOSX1 DFFPOSX1_1227 ( .CLK(clk), .D(u2__0remHi_451_0__320_), .Q(u2_remHi_320_));
DFFPOSX1 DFFPOSX1_1228 ( .CLK(clk), .D(u2__0remHi_451_0__321_), .Q(u2_remHi_321_));
DFFPOSX1 DFFPOSX1_1229 ( .CLK(clk), .D(u2__0remHi_451_0__322_), .Q(u2_remHi_322_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk), .D(u2__0root_452_0__119_), .Q(sqrto_118_));
DFFPOSX1 DFFPOSX1_1230 ( .CLK(clk), .D(u2__0remHi_451_0__323_), .Q(u2_remHi_323_));
DFFPOSX1 DFFPOSX1_1231 ( .CLK(clk), .D(u2__0remHi_451_0__324_), .Q(u2_remHi_324_));
DFFPOSX1 DFFPOSX1_1232 ( .CLK(clk), .D(u2__0remHi_451_0__325_), .Q(u2_remHi_325_));
DFFPOSX1 DFFPOSX1_1233 ( .CLK(clk), .D(u2__0remHi_451_0__326_), .Q(u2_remHi_326_));
DFFPOSX1 DFFPOSX1_1234 ( .CLK(clk), .D(u2__0remHi_451_0__327_), .Q(u2_remHi_327_));
DFFPOSX1 DFFPOSX1_1235 ( .CLK(clk), .D(u2__0remHi_451_0__328_), .Q(u2_remHi_328_));
DFFPOSX1 DFFPOSX1_1236 ( .CLK(clk), .D(u2__0remHi_451_0__329_), .Q(u2_remHi_329_));
DFFPOSX1 DFFPOSX1_1237 ( .CLK(clk), .D(u2__0remHi_451_0__330_), .Q(u2_remHi_330_));
DFFPOSX1 DFFPOSX1_1238 ( .CLK(clk), .D(u2__0remHi_451_0__331_), .Q(u2_remHi_331_));
DFFPOSX1 DFFPOSX1_1239 ( .CLK(clk), .D(u2__0remHi_451_0__332_), .Q(u2_remHi_332_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk), .D(u2__0root_452_0__120_), .Q(sqrto_119_));
DFFPOSX1 DFFPOSX1_1240 ( .CLK(clk), .D(u2__0remHi_451_0__333_), .Q(u2_remHi_333_));
DFFPOSX1 DFFPOSX1_1241 ( .CLK(clk), .D(u2__0remHi_451_0__334_), .Q(u2_remHi_334_));
DFFPOSX1 DFFPOSX1_1242 ( .CLK(clk), .D(u2__0remHi_451_0__335_), .Q(u2_remHi_335_));
DFFPOSX1 DFFPOSX1_1243 ( .CLK(clk), .D(u2__0remHi_451_0__336_), .Q(u2_remHi_336_));
DFFPOSX1 DFFPOSX1_1244 ( .CLK(clk), .D(u2__0remHi_451_0__337_), .Q(u2_remHi_337_));
DFFPOSX1 DFFPOSX1_1245 ( .CLK(clk), .D(u2__0remHi_451_0__338_), .Q(u2_remHi_338_));
DFFPOSX1 DFFPOSX1_1246 ( .CLK(clk), .D(u2__0remHi_451_0__339_), .Q(u2_remHi_339_));
DFFPOSX1 DFFPOSX1_1247 ( .CLK(clk), .D(u2__0remHi_451_0__340_), .Q(u2_remHi_340_));
DFFPOSX1 DFFPOSX1_1248 ( .CLK(clk), .D(u2__0remHi_451_0__341_), .Q(u2_remHi_341_));
DFFPOSX1 DFFPOSX1_1249 ( .CLK(clk), .D(u2__0remHi_451_0__342_), .Q(u2_remHi_342_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk), .D(u2__0root_452_0__121_), .Q(sqrto_120_));
DFFPOSX1 DFFPOSX1_1250 ( .CLK(clk), .D(u2__0remHi_451_0__343_), .Q(u2_remHi_343_));
DFFPOSX1 DFFPOSX1_1251 ( .CLK(clk), .D(u2__0remHi_451_0__344_), .Q(u2_remHi_344_));
DFFPOSX1 DFFPOSX1_1252 ( .CLK(clk), .D(u2__0remHi_451_0__345_), .Q(u2_remHi_345_));
DFFPOSX1 DFFPOSX1_1253 ( .CLK(clk), .D(u2__0remHi_451_0__346_), .Q(u2_remHi_346_));
DFFPOSX1 DFFPOSX1_1254 ( .CLK(clk), .D(u2__0remHi_451_0__347_), .Q(u2_remHi_347_));
DFFPOSX1 DFFPOSX1_1255 ( .CLK(clk), .D(u2__0remHi_451_0__348_), .Q(u2_remHi_348_));
DFFPOSX1 DFFPOSX1_1256 ( .CLK(clk), .D(u2__0remHi_451_0__349_), .Q(u2_remHi_349_));
DFFPOSX1 DFFPOSX1_1257 ( .CLK(clk), .D(u2__0remHi_451_0__350_), .Q(u2_remHi_350_));
DFFPOSX1 DFFPOSX1_1258 ( .CLK(clk), .D(u2__0remHi_451_0__351_), .Q(u2_remHi_351_));
DFFPOSX1 DFFPOSX1_1259 ( .CLK(clk), .D(u2__0remHi_451_0__352_), .Q(u2_remHi_352_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk), .D(u2__0root_452_0__122_), .Q(sqrto_121_));
DFFPOSX1 DFFPOSX1_1260 ( .CLK(clk), .D(u2__0remHi_451_0__353_), .Q(u2_remHi_353_));
DFFPOSX1 DFFPOSX1_1261 ( .CLK(clk), .D(u2__0remHi_451_0__354_), .Q(u2_remHi_354_));
DFFPOSX1 DFFPOSX1_1262 ( .CLK(clk), .D(u2__0remHi_451_0__355_), .Q(u2_remHi_355_));
DFFPOSX1 DFFPOSX1_1263 ( .CLK(clk), .D(u2__0remHi_451_0__356_), .Q(u2_remHi_356_));
DFFPOSX1 DFFPOSX1_1264 ( .CLK(clk), .D(u2__0remHi_451_0__357_), .Q(u2_remHi_357_));
DFFPOSX1 DFFPOSX1_1265 ( .CLK(clk), .D(u2__0remHi_451_0__358_), .Q(u2_remHi_358_));
DFFPOSX1 DFFPOSX1_1266 ( .CLK(clk), .D(u2__0remHi_451_0__359_), .Q(u2_remHi_359_));
DFFPOSX1 DFFPOSX1_1267 ( .CLK(clk), .D(u2__0remHi_451_0__360_), .Q(u2_remHi_360_));
DFFPOSX1 DFFPOSX1_1268 ( .CLK(clk), .D(u2__0remHi_451_0__361_), .Q(u2_remHi_361_));
DFFPOSX1 DFFPOSX1_1269 ( .CLK(clk), .D(u2__0remHi_451_0__362_), .Q(u2_remHi_362_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk), .D(u2__0root_452_0__123_), .Q(sqrto_122_));
DFFPOSX1 DFFPOSX1_1270 ( .CLK(clk), .D(u2__0remHi_451_0__363_), .Q(u2_remHi_363_));
DFFPOSX1 DFFPOSX1_1271 ( .CLK(clk), .D(u2__0remHi_451_0__364_), .Q(u2_remHi_364_));
DFFPOSX1 DFFPOSX1_1272 ( .CLK(clk), .D(u2__0remHi_451_0__365_), .Q(u2_remHi_365_));
DFFPOSX1 DFFPOSX1_1273 ( .CLK(clk), .D(u2__0remHi_451_0__366_), .Q(u2_remHi_366_));
DFFPOSX1 DFFPOSX1_1274 ( .CLK(clk), .D(u2__0remHi_451_0__367_), .Q(u2_remHi_367_));
DFFPOSX1 DFFPOSX1_1275 ( .CLK(clk), .D(u2__0remHi_451_0__368_), .Q(u2_remHi_368_));
DFFPOSX1 DFFPOSX1_1276 ( .CLK(clk), .D(u2__0remHi_451_0__369_), .Q(u2_remHi_369_));
DFFPOSX1 DFFPOSX1_1277 ( .CLK(clk), .D(u2__0remHi_451_0__370_), .Q(u2_remHi_370_));
DFFPOSX1 DFFPOSX1_1278 ( .CLK(clk), .D(u2__0remHi_451_0__371_), .Q(u2_remHi_371_));
DFFPOSX1 DFFPOSX1_1279 ( .CLK(clk), .D(u2__0remHi_451_0__372_), .Q(u2_remHi_372_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk), .D(u2__0root_452_0__124_), .Q(sqrto_123_));
DFFPOSX1 DFFPOSX1_1280 ( .CLK(clk), .D(u2__0remHi_451_0__373_), .Q(u2_remHi_373_));
DFFPOSX1 DFFPOSX1_1281 ( .CLK(clk), .D(u2__0remHi_451_0__374_), .Q(u2_remHi_374_));
DFFPOSX1 DFFPOSX1_1282 ( .CLK(clk), .D(u2__0remHi_451_0__375_), .Q(u2_remHi_375_));
DFFPOSX1 DFFPOSX1_1283 ( .CLK(clk), .D(u2__0remHi_451_0__376_), .Q(u2_remHi_376_));
DFFPOSX1 DFFPOSX1_1284 ( .CLK(clk), .D(u2__0remHi_451_0__377_), .Q(u2_remHi_377_));
DFFPOSX1 DFFPOSX1_1285 ( .CLK(clk), .D(u2__0remHi_451_0__378_), .Q(u2_remHi_378_));
DFFPOSX1 DFFPOSX1_1286 ( .CLK(clk), .D(u2__0remHi_451_0__379_), .Q(u2_remHi_379_));
DFFPOSX1 DFFPOSX1_1287 ( .CLK(clk), .D(u2__0remHi_451_0__380_), .Q(u2_remHi_380_));
DFFPOSX1 DFFPOSX1_1288 ( .CLK(clk), .D(u2__0remHi_451_0__381_), .Q(u2_remHi_381_));
DFFPOSX1 DFFPOSX1_1289 ( .CLK(clk), .D(u2__0remHi_451_0__382_), .Q(u2_remHi_382_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk), .D(u2__0root_452_0__125_), .Q(sqrto_124_));
DFFPOSX1 DFFPOSX1_1290 ( .CLK(clk), .D(u2__0remHi_451_0__383_), .Q(u2_remHi_383_));
DFFPOSX1 DFFPOSX1_1291 ( .CLK(clk), .D(u2__0remHi_451_0__384_), .Q(u2_remHi_384_));
DFFPOSX1 DFFPOSX1_1292 ( .CLK(clk), .D(u2__0remHi_451_0__385_), .Q(u2_remHi_385_));
DFFPOSX1 DFFPOSX1_1293 ( .CLK(clk), .D(u2__0remHi_451_0__386_), .Q(u2_remHi_386_));
DFFPOSX1 DFFPOSX1_1294 ( .CLK(clk), .D(u2__0remHi_451_0__387_), .Q(u2_remHi_387_));
DFFPOSX1 DFFPOSX1_1295 ( .CLK(clk), .D(u2__0remHi_451_0__388_), .Q(u2_remHi_388_));
DFFPOSX1 DFFPOSX1_1296 ( .CLK(clk), .D(u2__0remHi_451_0__389_), .Q(u2_remHi_389_));
DFFPOSX1 DFFPOSX1_1297 ( .CLK(clk), .D(u2__0remHi_451_0__390_), .Q(u2_remHi_390_));
DFFPOSX1 DFFPOSX1_1298 ( .CLK(clk), .D(u2__0remHi_451_0__391_), .Q(u2_remHi_391_));
DFFPOSX1 DFFPOSX1_1299 ( .CLK(clk), .D(u2__0remHi_451_0__392_), .Q(u2_remHi_392_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(u2__0root_452_0__9_), .Q(sqrto_8_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk), .D(u2__0root_452_0__126_), .Q(sqrto_125_));
DFFPOSX1 DFFPOSX1_1300 ( .CLK(clk), .D(u2__0remHi_451_0__393_), .Q(u2_remHi_393_));
DFFPOSX1 DFFPOSX1_1301 ( .CLK(clk), .D(u2__0remHi_451_0__394_), .Q(u2_remHi_394_));
DFFPOSX1 DFFPOSX1_1302 ( .CLK(clk), .D(u2__0remHi_451_0__395_), .Q(u2_remHi_395_));
DFFPOSX1 DFFPOSX1_1303 ( .CLK(clk), .D(u2__0remHi_451_0__396_), .Q(u2_remHi_396_));
DFFPOSX1 DFFPOSX1_1304 ( .CLK(clk), .D(u2__0remHi_451_0__397_), .Q(u2_remHi_397_));
DFFPOSX1 DFFPOSX1_1305 ( .CLK(clk), .D(u2__0remHi_451_0__398_), .Q(u2_remHi_398_));
DFFPOSX1 DFFPOSX1_1306 ( .CLK(clk), .D(u2__0remHi_451_0__399_), .Q(u2_remHi_399_));
DFFPOSX1 DFFPOSX1_1307 ( .CLK(clk), .D(u2__0remHi_451_0__400_), .Q(u2_remHi_400_));
DFFPOSX1 DFFPOSX1_1308 ( .CLK(clk), .D(u2__0remHi_451_0__401_), .Q(u2_remHi_401_));
DFFPOSX1 DFFPOSX1_1309 ( .CLK(clk), .D(u2__0remHi_451_0__402_), .Q(u2_remHi_402_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk), .D(u2__0root_452_0__127_), .Q(sqrto_126_));
DFFPOSX1 DFFPOSX1_1310 ( .CLK(clk), .D(u2__0remHi_451_0__403_), .Q(u2_remHi_403_));
DFFPOSX1 DFFPOSX1_1311 ( .CLK(clk), .D(u2__0remHi_451_0__404_), .Q(u2_remHi_404_));
DFFPOSX1 DFFPOSX1_1312 ( .CLK(clk), .D(u2__0remHi_451_0__405_), .Q(u2_remHi_405_));
DFFPOSX1 DFFPOSX1_1313 ( .CLK(clk), .D(u2__0remHi_451_0__406_), .Q(u2_remHi_406_));
DFFPOSX1 DFFPOSX1_1314 ( .CLK(clk), .D(u2__0remHi_451_0__407_), .Q(u2_remHi_407_));
DFFPOSX1 DFFPOSX1_1315 ( .CLK(clk), .D(u2__0remHi_451_0__408_), .Q(u2_remHi_408_));
DFFPOSX1 DFFPOSX1_1316 ( .CLK(clk), .D(u2__0remHi_451_0__409_), .Q(u2_remHi_409_));
DFFPOSX1 DFFPOSX1_1317 ( .CLK(clk), .D(u2__0remHi_451_0__410_), .Q(u2_remHi_410_));
DFFPOSX1 DFFPOSX1_1318 ( .CLK(clk), .D(u2__0remHi_451_0__411_), .Q(u2_remHi_411_));
DFFPOSX1 DFFPOSX1_1319 ( .CLK(clk), .D(u2__0remHi_451_0__412_), .Q(u2_remHi_412_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk), .D(u2__0root_452_0__128_), .Q(sqrto_127_));
DFFPOSX1 DFFPOSX1_1320 ( .CLK(clk), .D(u2__0remHi_451_0__413_), .Q(u2_remHi_413_));
DFFPOSX1 DFFPOSX1_1321 ( .CLK(clk), .D(u2__0remHi_451_0__414_), .Q(u2_remHi_414_));
DFFPOSX1 DFFPOSX1_1322 ( .CLK(clk), .D(u2__0remHi_451_0__415_), .Q(u2_remHi_415_));
DFFPOSX1 DFFPOSX1_1323 ( .CLK(clk), .D(u2__0remHi_451_0__416_), .Q(u2_remHi_416_));
DFFPOSX1 DFFPOSX1_1324 ( .CLK(clk), .D(u2__0remHi_451_0__417_), .Q(u2_remHi_417_));
DFFPOSX1 DFFPOSX1_1325 ( .CLK(clk), .D(u2__0remHi_451_0__418_), .Q(u2_remHi_418_));
DFFPOSX1 DFFPOSX1_1326 ( .CLK(clk), .D(u2__0remHi_451_0__419_), .Q(u2_remHi_419_));
DFFPOSX1 DFFPOSX1_1327 ( .CLK(clk), .D(u2__0remHi_451_0__420_), .Q(u2_remHi_420_));
DFFPOSX1 DFFPOSX1_1328 ( .CLK(clk), .D(u2__0remHi_451_0__421_), .Q(u2_remHi_421_));
DFFPOSX1 DFFPOSX1_1329 ( .CLK(clk), .D(u2__0remHi_451_0__422_), .Q(u2_remHi_422_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk), .D(u2__0root_452_0__129_), .Q(sqrto_128_));
DFFPOSX1 DFFPOSX1_1330 ( .CLK(clk), .D(u2__0remHi_451_0__423_), .Q(u2_remHi_423_));
DFFPOSX1 DFFPOSX1_1331 ( .CLK(clk), .D(u2__0remHi_451_0__424_), .Q(u2_remHi_424_));
DFFPOSX1 DFFPOSX1_1332 ( .CLK(clk), .D(u2__0remHi_451_0__425_), .Q(u2_remHi_425_));
DFFPOSX1 DFFPOSX1_1333 ( .CLK(clk), .D(u2__0remHi_451_0__426_), .Q(u2_remHi_426_));
DFFPOSX1 DFFPOSX1_1334 ( .CLK(clk), .D(u2__0remHi_451_0__427_), .Q(u2_remHi_427_));
DFFPOSX1 DFFPOSX1_1335 ( .CLK(clk), .D(u2__0remHi_451_0__428_), .Q(u2_remHi_428_));
DFFPOSX1 DFFPOSX1_1336 ( .CLK(clk), .D(u2__0remHi_451_0__429_), .Q(u2_remHi_429_));
DFFPOSX1 DFFPOSX1_1337 ( .CLK(clk), .D(u2__0remHi_451_0__430_), .Q(u2_remHi_430_));
DFFPOSX1 DFFPOSX1_1338 ( .CLK(clk), .D(u2__0remHi_451_0__431_), .Q(u2_remHi_431_));
DFFPOSX1 DFFPOSX1_1339 ( .CLK(clk), .D(u2__0remHi_451_0__432_), .Q(u2_remHi_432_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk), .D(u2__0root_452_0__130_), .Q(sqrto_129_));
DFFPOSX1 DFFPOSX1_1340 ( .CLK(clk), .D(u2__0remHi_451_0__433_), .Q(u2_remHi_433_));
DFFPOSX1 DFFPOSX1_1341 ( .CLK(clk), .D(u2__0remHi_451_0__434_), .Q(u2_remHi_434_));
DFFPOSX1 DFFPOSX1_1342 ( .CLK(clk), .D(u2__0remHi_451_0__435_), .Q(u2_remHi_435_));
DFFPOSX1 DFFPOSX1_1343 ( .CLK(clk), .D(u2__0remHi_451_0__436_), .Q(u2_remHi_436_));
DFFPOSX1 DFFPOSX1_1344 ( .CLK(clk), .D(u2__0remHi_451_0__437_), .Q(u2_remHi_437_));
DFFPOSX1 DFFPOSX1_1345 ( .CLK(clk), .D(u2__0remHi_451_0__438_), .Q(u2_remHi_438_));
DFFPOSX1 DFFPOSX1_1346 ( .CLK(clk), .D(u2__0remHi_451_0__439_), .Q(u2_remHi_439_));
DFFPOSX1 DFFPOSX1_1347 ( .CLK(clk), .D(u2__0remHi_451_0__440_), .Q(u2_remHi_440_));
DFFPOSX1 DFFPOSX1_1348 ( .CLK(clk), .D(u2__0remHi_451_0__441_), .Q(u2_remHi_441_));
DFFPOSX1 DFFPOSX1_1349 ( .CLK(clk), .D(u2__0remHi_451_0__442_), .Q(u2_remHi_442_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk), .D(u2__0root_452_0__131_), .Q(sqrto_130_));
DFFPOSX1 DFFPOSX1_1350 ( .CLK(clk), .D(u2__0remHi_451_0__443_), .Q(u2_remHi_443_));
DFFPOSX1 DFFPOSX1_1351 ( .CLK(clk), .D(u2__0remHi_451_0__444_), .Q(u2_remHi_444_));
DFFPOSX1 DFFPOSX1_1352 ( .CLK(clk), .D(u2__0remHi_451_0__445_), .Q(u2_remHi_445_));
DFFPOSX1 DFFPOSX1_1353 ( .CLK(clk), .D(u2__0remHi_451_0__446_), .Q(u2_remHi_446_));
DFFPOSX1 DFFPOSX1_1354 ( .CLK(clk), .D(u2__0remHi_451_0__447_), .Q(u2_remHi_447_));
DFFPOSX1 DFFPOSX1_1355 ( .CLK(clk), .D(u2__0remHi_451_0__448_), .Q(u2_remHi_448_));
DFFPOSX1 DFFPOSX1_1356 ( .CLK(clk), .D(u2__0remHi_451_0__449_), .Q(u2_remHi_449_));
DFFPOSX1 DFFPOSX1_1357 ( .CLK(clk), .D(u2__0cnt_7_0__0_), .Q(u2_cnt_0_));
DFFPOSX1 DFFPOSX1_1358 ( .CLK(clk), .D(u2__0cnt_7_0__1_), .Q(u2_cnt_1_));
DFFPOSX1 DFFPOSX1_1359 ( .CLK(clk), .D(u2__0cnt_7_0__2_), .Q(u2_cnt_2_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk), .D(u2__0root_452_0__132_), .Q(sqrto_131_));
DFFPOSX1 DFFPOSX1_1360 ( .CLK(clk), .D(u2__0cnt_7_0__3_), .Q(u2_cnt_3_));
DFFPOSX1 DFFPOSX1_1361 ( .CLK(clk), .D(u2__0cnt_7_0__4_), .Q(u2_cnt_4_));
DFFPOSX1 DFFPOSX1_1362 ( .CLK(clk), .D(u2__0cnt_7_0__5_), .Q(u2_cnt_5_));
DFFPOSX1 DFFPOSX1_1363 ( .CLK(clk), .D(u2__0cnt_7_0__6_), .Q(u2_cnt_6_));
DFFPOSX1 DFFPOSX1_1364 ( .CLK(clk), .D(u2__0cnt_7_0__7_), .Q(u2_cnt_7_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk), .D(u2__0root_452_0__133_), .Q(sqrto_132_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk), .D(u2__0root_452_0__134_), .Q(sqrto_133_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk), .D(u2__0root_452_0__135_), .Q(sqrto_134_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(u2__0root_452_0__10_), .Q(sqrto_9_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk), .D(u2__0root_452_0__136_), .Q(sqrto_135_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk), .D(u2__0root_452_0__137_), .Q(sqrto_136_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk), .D(u2__0root_452_0__138_), .Q(sqrto_137_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk), .D(u2__0root_452_0__139_), .Q(sqrto_138_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk), .D(u2__0root_452_0__140_), .Q(sqrto_139_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk), .D(u2__0root_452_0__141_), .Q(sqrto_140_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk), .D(u2__0root_452_0__142_), .Q(sqrto_141_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk), .D(u2__0root_452_0__143_), .Q(sqrto_142_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk), .D(u2__0root_452_0__144_), .Q(sqrto_143_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk), .D(u2__0root_452_0__145_), .Q(sqrto_144_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(u2__0root_452_0__11_), .Q(sqrto_10_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk), .D(u2__0root_452_0__146_), .Q(sqrto_145_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk), .D(u2__0root_452_0__147_), .Q(sqrto_146_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk), .D(u2__0root_452_0__148_), .Q(sqrto_147_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk), .D(u2__0root_452_0__149_), .Q(sqrto_148_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk), .D(u2__0root_452_0__150_), .Q(sqrto_149_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk), .D(u2__0root_452_0__151_), .Q(sqrto_150_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk), .D(u2__0root_452_0__152_), .Q(sqrto_151_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk), .D(u2__0root_452_0__153_), .Q(sqrto_152_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk), .D(u2__0root_452_0__154_), .Q(sqrto_153_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk), .D(u2__0root_452_0__155_), .Q(sqrto_154_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk), .D(u2__0root_452_0__12_), .Q(sqrto_11_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk), .D(u2__0root_452_0__156_), .Q(sqrto_155_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk), .D(u2__0root_452_0__157_), .Q(sqrto_156_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk), .D(u2__0root_452_0__158_), .Q(sqrto_157_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk), .D(u2__0root_452_0__159_), .Q(sqrto_158_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk), .D(u2__0root_452_0__160_), .Q(sqrto_159_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk), .D(u2__0root_452_0__161_), .Q(sqrto_160_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk), .D(u2__0root_452_0__162_), .Q(sqrto_161_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk), .D(u2__0root_452_0__163_), .Q(sqrto_162_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk), .D(u2__0root_452_0__164_), .Q(sqrto_163_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk), .D(u2__0root_452_0__165_), .Q(sqrto_164_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk), .D(u2__0root_452_0__13_), .Q(sqrto_12_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk), .D(u2__0root_452_0__166_), .Q(sqrto_165_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk), .D(u2__0root_452_0__167_), .Q(sqrto_166_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk), .D(u2__0root_452_0__168_), .Q(sqrto_167_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk), .D(u2__0root_452_0__169_), .Q(sqrto_168_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk), .D(u2__0root_452_0__170_), .Q(sqrto_169_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk), .D(u2__0root_452_0__171_), .Q(sqrto_170_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk), .D(u2__0root_452_0__172_), .Q(sqrto_171_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk), .D(u2__0root_452_0__173_), .Q(sqrto_172_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk), .D(u2__0root_452_0__174_), .Q(sqrto_173_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk), .D(u2__0root_452_0__175_), .Q(sqrto_174_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk), .D(u2__0root_452_0__14_), .Q(sqrto_13_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk), .D(u2__0root_452_0__176_), .Q(sqrto_175_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk), .D(u2__0root_452_0__177_), .Q(sqrto_176_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk), .D(u2__0root_452_0__178_), .Q(sqrto_177_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk), .D(u2__0root_452_0__179_), .Q(sqrto_178_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk), .D(u2__0root_452_0__180_), .Q(sqrto_179_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk), .D(u2__0root_452_0__181_), .Q(sqrto_180_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(clk), .D(u2__0root_452_0__182_), .Q(sqrto_181_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(clk), .D(u2__0root_452_0__183_), .Q(sqrto_182_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(clk), .D(u2__0root_452_0__184_), .Q(sqrto_183_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(clk), .D(u2__0root_452_0__185_), .Q(sqrto_184_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk), .D(u2__0root_452_0__15_), .Q(sqrto_14_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(clk), .D(u2__0root_452_0__186_), .Q(sqrto_185_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(clk), .D(u2__0root_452_0__187_), .Q(sqrto_186_));
DFFPOSX1 DFFPOSX1_192 ( .CLK(clk), .D(u2__0root_452_0__188_), .Q(sqrto_187_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(clk), .D(u2__0root_452_0__189_), .Q(sqrto_188_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(clk), .D(u2__0root_452_0__190_), .Q(sqrto_189_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(clk), .D(u2__0root_452_0__191_), .Q(sqrto_190_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(clk), .D(u2__0root_452_0__192_), .Q(sqrto_191_));
DFFPOSX1 DFFPOSX1_197 ( .CLK(clk), .D(u2__0root_452_0__193_), .Q(sqrto_192_));
DFFPOSX1 DFFPOSX1_198 ( .CLK(clk), .D(u2__0root_452_0__194_), .Q(sqrto_193_));
DFFPOSX1 DFFPOSX1_199 ( .CLK(clk), .D(u2__0root_452_0__195_), .Q(sqrto_194_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_1_), .Q(done));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk), .D(u2__0root_452_0__16_), .Q(sqrto_15_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(clk), .D(u2__0root_452_0__196_), .Q(sqrto_195_));
DFFPOSX1 DFFPOSX1_201 ( .CLK(clk), .D(u2__0root_452_0__197_), .Q(sqrto_196_));
DFFPOSX1 DFFPOSX1_202 ( .CLK(clk), .D(u2__0root_452_0__198_), .Q(sqrto_197_));
DFFPOSX1 DFFPOSX1_203 ( .CLK(clk), .D(u2__0root_452_0__199_), .Q(sqrto_198_));
DFFPOSX1 DFFPOSX1_204 ( .CLK(clk), .D(u2__0root_452_0__200_), .Q(sqrto_199_));
DFFPOSX1 DFFPOSX1_205 ( .CLK(clk), .D(u2__0root_452_0__201_), .Q(sqrto_200_));
DFFPOSX1 DFFPOSX1_206 ( .CLK(clk), .D(u2__0root_452_0__202_), .Q(sqrto_201_));
DFFPOSX1 DFFPOSX1_207 ( .CLK(clk), .D(u2__0root_452_0__203_), .Q(sqrto_202_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(clk), .D(u2__0root_452_0__204_), .Q(sqrto_203_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(clk), .D(u2__0root_452_0__205_), .Q(sqrto_204_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk), .D(u2__0root_452_0__17_), .Q(sqrto_16_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(clk), .D(u2__0root_452_0__206_), .Q(sqrto_205_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(clk), .D(u2__0root_452_0__207_), .Q(sqrto_206_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(clk), .D(u2__0root_452_0__208_), .Q(sqrto_207_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(clk), .D(u2__0root_452_0__209_), .Q(sqrto_208_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(clk), .D(u2__0root_452_0__210_), .Q(sqrto_209_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(clk), .D(u2__0root_452_0__211_), .Q(sqrto_210_));
DFFPOSX1 DFFPOSX1_216 ( .CLK(clk), .D(u2__0root_452_0__212_), .Q(sqrto_211_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(clk), .D(u2__0root_452_0__213_), .Q(sqrto_212_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(clk), .D(u2__0root_452_0__214_), .Q(sqrto_213_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(clk), .D(u2__0root_452_0__215_), .Q(sqrto_214_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk), .D(u2__0root_452_0__18_), .Q(sqrto_17_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(clk), .D(u2__0root_452_0__216_), .Q(sqrto_215_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(clk), .D(u2__0root_452_0__217_), .Q(sqrto_216_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(clk), .D(u2__0root_452_0__218_), .Q(sqrto_217_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(clk), .D(u2__0root_452_0__219_), .Q(sqrto_218_));
DFFPOSX1 DFFPOSX1_224 ( .CLK(clk), .D(u2__0root_452_0__220_), .Q(sqrto_219_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(clk), .D(u2__0root_452_0__221_), .Q(sqrto_220_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(clk), .D(u2__0root_452_0__222_), .Q(sqrto_221_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(clk), .D(u2__0root_452_0__223_), .Q(sqrto_222_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(clk), .D(u2__0root_452_0__224_), .Q(sqrto_223_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(clk), .D(u2__0root_452_0__225_), .Q(sqrto_224_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk), .D(u2__0root_452_0__19_), .Q(sqrto_18_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(clk), .D(u2__0root_452_0__226_), .Q(sqrto_225_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(clk), .D(u2__0root_452_0__227_), .Q(u2_o_226_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(clk), .D(u2__0root_452_0__228_), .Q(u2_o_227_));
DFFPOSX1 DFFPOSX1_233 ( .CLK(clk), .D(u2__0root_452_0__229_), .Q(u2_o_228_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(clk), .D(u2__0root_452_0__230_), .Q(u2_o_229_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(clk), .D(u2__0root_452_0__231_), .Q(u2_o_230_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(clk), .D(u2__0root_452_0__232_), .Q(u2_o_231_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(clk), .D(u2__0root_452_0__233_), .Q(u2_o_232_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(clk), .D(u2__0root_452_0__234_), .Q(u2_o_233_));
DFFPOSX1 DFFPOSX1_239 ( .CLK(clk), .D(u2__0root_452_0__235_), .Q(u2_o_234_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk), .D(u2__0root_452_0__20_), .Q(sqrto_19_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(clk), .D(u2__0root_452_0__236_), .Q(u2_o_235_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(clk), .D(u2__0root_452_0__237_), .Q(u2_o_236_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(clk), .D(u2__0root_452_0__238_), .Q(u2_o_237_));
DFFPOSX1 DFFPOSX1_243 ( .CLK(clk), .D(u2__0root_452_0__239_), .Q(u2_o_238_));
DFFPOSX1 DFFPOSX1_244 ( .CLK(clk), .D(u2__0root_452_0__240_), .Q(u2_o_239_));
DFFPOSX1 DFFPOSX1_245 ( .CLK(clk), .D(u2__0root_452_0__241_), .Q(u2_o_240_));
DFFPOSX1 DFFPOSX1_246 ( .CLK(clk), .D(u2__0root_452_0__242_), .Q(u2_o_241_));
DFFPOSX1 DFFPOSX1_247 ( .CLK(clk), .D(u2__0root_452_0__243_), .Q(u2_o_242_));
DFFPOSX1 DFFPOSX1_248 ( .CLK(clk), .D(u2__0root_452_0__244_), .Q(u2_o_243_));
DFFPOSX1 DFFPOSX1_249 ( .CLK(clk), .D(u2__0root_452_0__245_), .Q(u2_o_244_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk), .D(u2__0root_452_0__21_), .Q(sqrto_20_));
DFFPOSX1 DFFPOSX1_250 ( .CLK(clk), .D(u2__0root_452_0__246_), .Q(u2_o_245_));
DFFPOSX1 DFFPOSX1_251 ( .CLK(clk), .D(u2__0root_452_0__247_), .Q(u2_o_246_));
DFFPOSX1 DFFPOSX1_252 ( .CLK(clk), .D(u2__0root_452_0__248_), .Q(u2_o_247_));
DFFPOSX1 DFFPOSX1_253 ( .CLK(clk), .D(u2__0root_452_0__249_), .Q(u2_o_248_));
DFFPOSX1 DFFPOSX1_254 ( .CLK(clk), .D(u2__0root_452_0__250_), .Q(u2_o_249_));
DFFPOSX1 DFFPOSX1_255 ( .CLK(clk), .D(u2__0root_452_0__251_), .Q(u2_o_250_));
DFFPOSX1 DFFPOSX1_256 ( .CLK(clk), .D(u2__0root_452_0__252_), .Q(u2_o_251_));
DFFPOSX1 DFFPOSX1_257 ( .CLK(clk), .D(u2__0root_452_0__253_), .Q(u2_o_252_));
DFFPOSX1 DFFPOSX1_258 ( .CLK(clk), .D(u2__0root_452_0__254_), .Q(u2_o_253_));
DFFPOSX1 DFFPOSX1_259 ( .CLK(clk), .D(u2__0root_452_0__255_), .Q(u2_o_254_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk), .D(u2__0root_452_0__22_), .Q(sqrto_21_));
DFFPOSX1 DFFPOSX1_260 ( .CLK(clk), .D(u2__0root_452_0__256_), .Q(u2_o_255_));
DFFPOSX1 DFFPOSX1_261 ( .CLK(clk), .D(u2__0root_452_0__257_), .Q(u2_o_256_));
DFFPOSX1 DFFPOSX1_262 ( .CLK(clk), .D(u2__0root_452_0__258_), .Q(u2_o_257_));
DFFPOSX1 DFFPOSX1_263 ( .CLK(clk), .D(u2__0root_452_0__259_), .Q(u2_o_258_));
DFFPOSX1 DFFPOSX1_264 ( .CLK(clk), .D(u2__0root_452_0__260_), .Q(u2_o_259_));
DFFPOSX1 DFFPOSX1_265 ( .CLK(clk), .D(u2__0root_452_0__261_), .Q(u2_o_260_));
DFFPOSX1 DFFPOSX1_266 ( .CLK(clk), .D(u2__0root_452_0__262_), .Q(u2_o_261_));
DFFPOSX1 DFFPOSX1_267 ( .CLK(clk), .D(u2__0root_452_0__263_), .Q(u2_o_262_));
DFFPOSX1 DFFPOSX1_268 ( .CLK(clk), .D(u2__0root_452_0__264_), .Q(u2_o_263_));
DFFPOSX1 DFFPOSX1_269 ( .CLK(clk), .D(u2__0root_452_0__265_), .Q(u2_o_264_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk), .D(u2__0root_452_0__23_), .Q(sqrto_22_));
DFFPOSX1 DFFPOSX1_270 ( .CLK(clk), .D(u2__0root_452_0__266_), .Q(u2_o_265_));
DFFPOSX1 DFFPOSX1_271 ( .CLK(clk), .D(u2__0root_452_0__267_), .Q(u2_o_266_));
DFFPOSX1 DFFPOSX1_272 ( .CLK(clk), .D(u2__0root_452_0__268_), .Q(u2_o_267_));
DFFPOSX1 DFFPOSX1_273 ( .CLK(clk), .D(u2__0root_452_0__269_), .Q(u2_o_268_));
DFFPOSX1 DFFPOSX1_274 ( .CLK(clk), .D(u2__0root_452_0__270_), .Q(u2_o_269_));
DFFPOSX1 DFFPOSX1_275 ( .CLK(clk), .D(u2__0root_452_0__271_), .Q(u2_o_270_));
DFFPOSX1 DFFPOSX1_276 ( .CLK(clk), .D(u2__0root_452_0__272_), .Q(u2_o_271_));
DFFPOSX1 DFFPOSX1_277 ( .CLK(clk), .D(u2__0root_452_0__273_), .Q(u2_o_272_));
DFFPOSX1 DFFPOSX1_278 ( .CLK(clk), .D(u2__0root_452_0__274_), .Q(u2_o_273_));
DFFPOSX1 DFFPOSX1_279 ( .CLK(clk), .D(u2__0root_452_0__275_), .Q(u2_o_274_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk), .D(u2__0root_452_0__24_), .Q(sqrto_23_));
DFFPOSX1 DFFPOSX1_280 ( .CLK(clk), .D(u2__0root_452_0__276_), .Q(u2_o_275_));
DFFPOSX1 DFFPOSX1_281 ( .CLK(clk), .D(u2__0root_452_0__277_), .Q(u2_o_276_));
DFFPOSX1 DFFPOSX1_282 ( .CLK(clk), .D(u2__0root_452_0__278_), .Q(u2_o_277_));
DFFPOSX1 DFFPOSX1_283 ( .CLK(clk), .D(u2__0root_452_0__279_), .Q(u2_o_278_));
DFFPOSX1 DFFPOSX1_284 ( .CLK(clk), .D(u2__0root_452_0__280_), .Q(u2_o_279_));
DFFPOSX1 DFFPOSX1_285 ( .CLK(clk), .D(u2__0root_452_0__281_), .Q(u2_o_280_));
DFFPOSX1 DFFPOSX1_286 ( .CLK(clk), .D(u2__0root_452_0__282_), .Q(u2_o_281_));
DFFPOSX1 DFFPOSX1_287 ( .CLK(clk), .D(u2__0root_452_0__283_), .Q(u2_o_282_));
DFFPOSX1 DFFPOSX1_288 ( .CLK(clk), .D(u2__0root_452_0__284_), .Q(u2_o_283_));
DFFPOSX1 DFFPOSX1_289 ( .CLK(clk), .D(u2__0root_452_0__285_), .Q(u2_o_284_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk), .D(u2__0root_452_0__25_), .Q(sqrto_24_));
DFFPOSX1 DFFPOSX1_290 ( .CLK(clk), .D(u2__0root_452_0__286_), .Q(u2_o_285_));
DFFPOSX1 DFFPOSX1_291 ( .CLK(clk), .D(u2__0root_452_0__287_), .Q(u2_o_286_));
DFFPOSX1 DFFPOSX1_292 ( .CLK(clk), .D(u2__0root_452_0__288_), .Q(u2_o_287_));
DFFPOSX1 DFFPOSX1_293 ( .CLK(clk), .D(u2__0root_452_0__289_), .Q(u2_o_288_));
DFFPOSX1 DFFPOSX1_294 ( .CLK(clk), .D(u2__0root_452_0__290_), .Q(u2_o_289_));
DFFPOSX1 DFFPOSX1_295 ( .CLK(clk), .D(u2__0root_452_0__291_), .Q(u2_o_290_));
DFFPOSX1 DFFPOSX1_296 ( .CLK(clk), .D(u2__0root_452_0__292_), .Q(u2_o_291_));
DFFPOSX1 DFFPOSX1_297 ( .CLK(clk), .D(u2__0root_452_0__293_), .Q(u2_o_292_));
DFFPOSX1 DFFPOSX1_298 ( .CLK(clk), .D(u2__0root_452_0__294_), .Q(u2_o_293_));
DFFPOSX1 DFFPOSX1_299 ( .CLK(clk), .D(u2__0root_452_0__295_), .Q(u2_o_294_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_2_), .Q(u2_state_2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk), .D(u2__0root_452_0__26_), .Q(sqrto_25_));
DFFPOSX1 DFFPOSX1_300 ( .CLK(clk), .D(u2__0root_452_0__296_), .Q(u2_o_295_));
DFFPOSX1 DFFPOSX1_301 ( .CLK(clk), .D(u2__0root_452_0__297_), .Q(u2_o_296_));
DFFPOSX1 DFFPOSX1_302 ( .CLK(clk), .D(u2__0root_452_0__298_), .Q(u2_o_297_));
DFFPOSX1 DFFPOSX1_303 ( .CLK(clk), .D(u2__0root_452_0__299_), .Q(u2_o_298_));
DFFPOSX1 DFFPOSX1_304 ( .CLK(clk), .D(u2__0root_452_0__300_), .Q(u2_o_299_));
DFFPOSX1 DFFPOSX1_305 ( .CLK(clk), .D(u2__0root_452_0__301_), .Q(u2_o_300_));
DFFPOSX1 DFFPOSX1_306 ( .CLK(clk), .D(u2__0root_452_0__302_), .Q(u2_o_301_));
DFFPOSX1 DFFPOSX1_307 ( .CLK(clk), .D(u2__0root_452_0__303_), .Q(u2_o_302_));
DFFPOSX1 DFFPOSX1_308 ( .CLK(clk), .D(u2__0root_452_0__304_), .Q(u2_o_303_));
DFFPOSX1 DFFPOSX1_309 ( .CLK(clk), .D(u2__0root_452_0__305_), .Q(u2_o_304_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk), .D(u2__0root_452_0__27_), .Q(sqrto_26_));
DFFPOSX1 DFFPOSX1_310 ( .CLK(clk), .D(u2__0root_452_0__306_), .Q(u2_o_305_));
DFFPOSX1 DFFPOSX1_311 ( .CLK(clk), .D(u2__0root_452_0__307_), .Q(u2_o_306_));
DFFPOSX1 DFFPOSX1_312 ( .CLK(clk), .D(u2__0root_452_0__308_), .Q(u2_o_307_));
DFFPOSX1 DFFPOSX1_313 ( .CLK(clk), .D(u2__0root_452_0__309_), .Q(u2_o_308_));
DFFPOSX1 DFFPOSX1_314 ( .CLK(clk), .D(u2__0root_452_0__310_), .Q(u2_o_309_));
DFFPOSX1 DFFPOSX1_315 ( .CLK(clk), .D(u2__0root_452_0__311_), .Q(u2_o_310_));
DFFPOSX1 DFFPOSX1_316 ( .CLK(clk), .D(u2__0root_452_0__312_), .Q(u2_o_311_));
DFFPOSX1 DFFPOSX1_317 ( .CLK(clk), .D(u2__0root_452_0__313_), .Q(u2_o_312_));
DFFPOSX1 DFFPOSX1_318 ( .CLK(clk), .D(u2__0root_452_0__314_), .Q(u2_o_313_));
DFFPOSX1 DFFPOSX1_319 ( .CLK(clk), .D(u2__0root_452_0__315_), .Q(u2_o_314_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk), .D(u2__0root_452_0__28_), .Q(sqrto_27_));
DFFPOSX1 DFFPOSX1_320 ( .CLK(clk), .D(u2__0root_452_0__316_), .Q(u2_o_315_));
DFFPOSX1 DFFPOSX1_321 ( .CLK(clk), .D(u2__0root_452_0__317_), .Q(u2_o_316_));
DFFPOSX1 DFFPOSX1_322 ( .CLK(clk), .D(u2__0root_452_0__318_), .Q(u2_o_317_));
DFFPOSX1 DFFPOSX1_323 ( .CLK(clk), .D(u2__0root_452_0__319_), .Q(u2_o_318_));
DFFPOSX1 DFFPOSX1_324 ( .CLK(clk), .D(u2__0root_452_0__320_), .Q(u2_o_319_));
DFFPOSX1 DFFPOSX1_325 ( .CLK(clk), .D(u2__0root_452_0__321_), .Q(u2_o_320_));
DFFPOSX1 DFFPOSX1_326 ( .CLK(clk), .D(u2__0root_452_0__322_), .Q(u2_o_321_));
DFFPOSX1 DFFPOSX1_327 ( .CLK(clk), .D(u2__0root_452_0__323_), .Q(u2_o_322_));
DFFPOSX1 DFFPOSX1_328 ( .CLK(clk), .D(u2__0root_452_0__324_), .Q(u2_o_323_));
DFFPOSX1 DFFPOSX1_329 ( .CLK(clk), .D(u2__0root_452_0__325_), .Q(u2_o_324_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk), .D(u2__0root_452_0__29_), .Q(sqrto_28_));
DFFPOSX1 DFFPOSX1_330 ( .CLK(clk), .D(u2__0root_452_0__326_), .Q(u2_o_325_));
DFFPOSX1 DFFPOSX1_331 ( .CLK(clk), .D(u2__0root_452_0__327_), .Q(u2_o_326_));
DFFPOSX1 DFFPOSX1_332 ( .CLK(clk), .D(u2__0root_452_0__328_), .Q(u2_o_327_));
DFFPOSX1 DFFPOSX1_333 ( .CLK(clk), .D(u2__0root_452_0__329_), .Q(u2_o_328_));
DFFPOSX1 DFFPOSX1_334 ( .CLK(clk), .D(u2__0root_452_0__330_), .Q(u2_o_329_));
DFFPOSX1 DFFPOSX1_335 ( .CLK(clk), .D(u2__0root_452_0__331_), .Q(u2_o_330_));
DFFPOSX1 DFFPOSX1_336 ( .CLK(clk), .D(u2__0root_452_0__332_), .Q(u2_o_331_));
DFFPOSX1 DFFPOSX1_337 ( .CLK(clk), .D(u2__0root_452_0__333_), .Q(u2_o_332_));
DFFPOSX1 DFFPOSX1_338 ( .CLK(clk), .D(u2__0root_452_0__334_), .Q(u2_o_333_));
DFFPOSX1 DFFPOSX1_339 ( .CLK(clk), .D(u2__0root_452_0__335_), .Q(u2_o_334_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk), .D(u2__0root_452_0__30_), .Q(sqrto_29_));
DFFPOSX1 DFFPOSX1_340 ( .CLK(clk), .D(u2__0root_452_0__336_), .Q(u2_o_335_));
DFFPOSX1 DFFPOSX1_341 ( .CLK(clk), .D(u2__0root_452_0__337_), .Q(u2_o_336_));
DFFPOSX1 DFFPOSX1_342 ( .CLK(clk), .D(u2__0root_452_0__338_), .Q(u2_o_337_));
DFFPOSX1 DFFPOSX1_343 ( .CLK(clk), .D(u2__0root_452_0__339_), .Q(u2_o_338_));
DFFPOSX1 DFFPOSX1_344 ( .CLK(clk), .D(u2__0root_452_0__340_), .Q(u2_o_339_));
DFFPOSX1 DFFPOSX1_345 ( .CLK(clk), .D(u2__0root_452_0__341_), .Q(u2_o_340_));
DFFPOSX1 DFFPOSX1_346 ( .CLK(clk), .D(u2__0root_452_0__342_), .Q(u2_o_341_));
DFFPOSX1 DFFPOSX1_347 ( .CLK(clk), .D(u2__0root_452_0__343_), .Q(u2_o_342_));
DFFPOSX1 DFFPOSX1_348 ( .CLK(clk), .D(u2__0root_452_0__344_), .Q(u2_o_343_));
DFFPOSX1 DFFPOSX1_349 ( .CLK(clk), .D(u2__0root_452_0__345_), .Q(u2_o_344_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk), .D(u2__0root_452_0__31_), .Q(sqrto_30_));
DFFPOSX1 DFFPOSX1_350 ( .CLK(clk), .D(u2__0root_452_0__346_), .Q(u2_o_345_));
DFFPOSX1 DFFPOSX1_351 ( .CLK(clk), .D(u2__0root_452_0__347_), .Q(u2_o_346_));
DFFPOSX1 DFFPOSX1_352 ( .CLK(clk), .D(u2__0root_452_0__348_), .Q(u2_o_347_));
DFFPOSX1 DFFPOSX1_353 ( .CLK(clk), .D(u2__0root_452_0__349_), .Q(u2_o_348_));
DFFPOSX1 DFFPOSX1_354 ( .CLK(clk), .D(u2__0root_452_0__350_), .Q(u2_o_349_));
DFFPOSX1 DFFPOSX1_355 ( .CLK(clk), .D(u2__0root_452_0__351_), .Q(u2_o_350_));
DFFPOSX1 DFFPOSX1_356 ( .CLK(clk), .D(u2__0root_452_0__352_), .Q(u2_o_351_));
DFFPOSX1 DFFPOSX1_357 ( .CLK(clk), .D(u2__0root_452_0__353_), .Q(u2_o_352_));
DFFPOSX1 DFFPOSX1_358 ( .CLK(clk), .D(u2__0root_452_0__354_), .Q(u2_o_353_));
DFFPOSX1 DFFPOSX1_359 ( .CLK(clk), .D(u2__0root_452_0__355_), .Q(u2_o_354_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk), .D(u2__0root_452_0__32_), .Q(sqrto_31_));
DFFPOSX1 DFFPOSX1_360 ( .CLK(clk), .D(u2__0root_452_0__356_), .Q(u2_o_355_));
DFFPOSX1 DFFPOSX1_361 ( .CLK(clk), .D(u2__0root_452_0__357_), .Q(u2_o_356_));
DFFPOSX1 DFFPOSX1_362 ( .CLK(clk), .D(u2__0root_452_0__358_), .Q(u2_o_357_));
DFFPOSX1 DFFPOSX1_363 ( .CLK(clk), .D(u2__0root_452_0__359_), .Q(u2_o_358_));
DFFPOSX1 DFFPOSX1_364 ( .CLK(clk), .D(u2__0root_452_0__360_), .Q(u2_o_359_));
DFFPOSX1 DFFPOSX1_365 ( .CLK(clk), .D(u2__0root_452_0__361_), .Q(u2_o_360_));
DFFPOSX1 DFFPOSX1_366 ( .CLK(clk), .D(u2__0root_452_0__362_), .Q(u2_o_361_));
DFFPOSX1 DFFPOSX1_367 ( .CLK(clk), .D(u2__0root_452_0__363_), .Q(u2_o_362_));
DFFPOSX1 DFFPOSX1_368 ( .CLK(clk), .D(u2__0root_452_0__364_), .Q(u2_o_363_));
DFFPOSX1 DFFPOSX1_369 ( .CLK(clk), .D(u2__0root_452_0__365_), .Q(u2_o_364_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk), .D(u2__0root_452_0__33_), .Q(sqrto_32_));
DFFPOSX1 DFFPOSX1_370 ( .CLK(clk), .D(u2__0root_452_0__366_), .Q(u2_o_365_));
DFFPOSX1 DFFPOSX1_371 ( .CLK(clk), .D(u2__0root_452_0__367_), .Q(u2_o_366_));
DFFPOSX1 DFFPOSX1_372 ( .CLK(clk), .D(u2__0root_452_0__368_), .Q(u2_o_367_));
DFFPOSX1 DFFPOSX1_373 ( .CLK(clk), .D(u2__0root_452_0__369_), .Q(u2_o_368_));
DFFPOSX1 DFFPOSX1_374 ( .CLK(clk), .D(u2__0root_452_0__370_), .Q(u2_o_369_));
DFFPOSX1 DFFPOSX1_375 ( .CLK(clk), .D(u2__0root_452_0__371_), .Q(u2_o_370_));
DFFPOSX1 DFFPOSX1_376 ( .CLK(clk), .D(u2__0root_452_0__372_), .Q(u2_o_371_));
DFFPOSX1 DFFPOSX1_377 ( .CLK(clk), .D(u2__0root_452_0__373_), .Q(u2_o_372_));
DFFPOSX1 DFFPOSX1_378 ( .CLK(clk), .D(u2__0root_452_0__374_), .Q(u2_o_373_));
DFFPOSX1 DFFPOSX1_379 ( .CLK(clk), .D(u2__0root_452_0__375_), .Q(u2_o_374_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk), .D(u2__0root_452_0__34_), .Q(sqrto_33_));
DFFPOSX1 DFFPOSX1_380 ( .CLK(clk), .D(u2__0root_452_0__376_), .Q(u2_o_375_));
DFFPOSX1 DFFPOSX1_381 ( .CLK(clk), .D(u2__0root_452_0__377_), .Q(u2_o_376_));
DFFPOSX1 DFFPOSX1_382 ( .CLK(clk), .D(u2__0root_452_0__378_), .Q(u2_o_377_));
DFFPOSX1 DFFPOSX1_383 ( .CLK(clk), .D(u2__0root_452_0__379_), .Q(u2_o_378_));
DFFPOSX1 DFFPOSX1_384 ( .CLK(clk), .D(u2__0root_452_0__380_), .Q(u2_o_379_));
DFFPOSX1 DFFPOSX1_385 ( .CLK(clk), .D(u2__0root_452_0__381_), .Q(u2_o_380_));
DFFPOSX1 DFFPOSX1_386 ( .CLK(clk), .D(u2__0root_452_0__382_), .Q(u2_o_381_));
DFFPOSX1 DFFPOSX1_387 ( .CLK(clk), .D(u2__0root_452_0__383_), .Q(u2_o_382_));
DFFPOSX1 DFFPOSX1_388 ( .CLK(clk), .D(u2__0root_452_0__384_), .Q(u2_o_383_));
DFFPOSX1 DFFPOSX1_389 ( .CLK(clk), .D(u2__0root_452_0__385_), .Q(u2_o_384_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk), .D(u2__0root_452_0__35_), .Q(sqrto_34_));
DFFPOSX1 DFFPOSX1_390 ( .CLK(clk), .D(u2__0root_452_0__386_), .Q(u2_o_385_));
DFFPOSX1 DFFPOSX1_391 ( .CLK(clk), .D(u2__0root_452_0__387_), .Q(u2_o_386_));
DFFPOSX1 DFFPOSX1_392 ( .CLK(clk), .D(u2__0root_452_0__388_), .Q(u2_o_387_));
DFFPOSX1 DFFPOSX1_393 ( .CLK(clk), .D(u2__0root_452_0__389_), .Q(u2_o_388_));
DFFPOSX1 DFFPOSX1_394 ( .CLK(clk), .D(u2__0root_452_0__390_), .Q(u2_o_389_));
DFFPOSX1 DFFPOSX1_395 ( .CLK(clk), .D(u2__0root_452_0__391_), .Q(u2_o_390_));
DFFPOSX1 DFFPOSX1_396 ( .CLK(clk), .D(u2__0root_452_0__392_), .Q(u2_o_391_));
DFFPOSX1 DFFPOSX1_397 ( .CLK(clk), .D(u2__0root_452_0__393_), .Q(u2_o_392_));
DFFPOSX1 DFFPOSX1_398 ( .CLK(clk), .D(u2__0root_452_0__394_), .Q(u2_o_393_));
DFFPOSX1 DFFPOSX1_399 ( .CLK(clk), .D(u2__0root_452_0__395_), .Q(u2_o_394_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(u2__0root_452_0__0_), .Q(u2_root_0_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk), .D(u2__0root_452_0__36_), .Q(sqrto_35_));
DFFPOSX1 DFFPOSX1_400 ( .CLK(clk), .D(u2__0root_452_0__396_), .Q(u2_o_395_));
DFFPOSX1 DFFPOSX1_401 ( .CLK(clk), .D(u2__0root_452_0__397_), .Q(u2_o_396_));
DFFPOSX1 DFFPOSX1_402 ( .CLK(clk), .D(u2__0root_452_0__398_), .Q(u2_o_397_));
DFFPOSX1 DFFPOSX1_403 ( .CLK(clk), .D(u2__0root_452_0__399_), .Q(u2_o_398_));
DFFPOSX1 DFFPOSX1_404 ( .CLK(clk), .D(u2__0root_452_0__400_), .Q(u2_o_399_));
DFFPOSX1 DFFPOSX1_405 ( .CLK(clk), .D(u2__0root_452_0__401_), .Q(u2_o_400_));
DFFPOSX1 DFFPOSX1_406 ( .CLK(clk), .D(u2__0root_452_0__402_), .Q(u2_o_401_));
DFFPOSX1 DFFPOSX1_407 ( .CLK(clk), .D(u2__0root_452_0__403_), .Q(u2_o_402_));
DFFPOSX1 DFFPOSX1_408 ( .CLK(clk), .D(u2__0root_452_0__404_), .Q(u2_o_403_));
DFFPOSX1 DFFPOSX1_409 ( .CLK(clk), .D(u2__0root_452_0__405_), .Q(u2_o_404_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk), .D(u2__0root_452_0__37_), .Q(sqrto_36_));
DFFPOSX1 DFFPOSX1_410 ( .CLK(clk), .D(u2__0root_452_0__406_), .Q(u2_o_405_));
DFFPOSX1 DFFPOSX1_411 ( .CLK(clk), .D(u2__0root_452_0__407_), .Q(u2_o_406_));
DFFPOSX1 DFFPOSX1_412 ( .CLK(clk), .D(u2__0root_452_0__408_), .Q(u2_o_407_));
DFFPOSX1 DFFPOSX1_413 ( .CLK(clk), .D(u2__0root_452_0__409_), .Q(u2_o_408_));
DFFPOSX1 DFFPOSX1_414 ( .CLK(clk), .D(u2__0root_452_0__410_), .Q(u2_o_409_));
DFFPOSX1 DFFPOSX1_415 ( .CLK(clk), .D(u2__0root_452_0__411_), .Q(u2_o_410_));
DFFPOSX1 DFFPOSX1_416 ( .CLK(clk), .D(u2__0root_452_0__412_), .Q(u2_o_411_));
DFFPOSX1 DFFPOSX1_417 ( .CLK(clk), .D(u2__0root_452_0__413_), .Q(u2_o_412_));
DFFPOSX1 DFFPOSX1_418 ( .CLK(clk), .D(u2__0root_452_0__414_), .Q(u2_o_413_));
DFFPOSX1 DFFPOSX1_419 ( .CLK(clk), .D(u2__0root_452_0__415_), .Q(u2_o_414_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk), .D(u2__0root_452_0__38_), .Q(sqrto_37_));
DFFPOSX1 DFFPOSX1_420 ( .CLK(clk), .D(u2__0root_452_0__416_), .Q(u2_o_415_));
DFFPOSX1 DFFPOSX1_421 ( .CLK(clk), .D(u2__0root_452_0__417_), .Q(u2_o_416_));
DFFPOSX1 DFFPOSX1_422 ( .CLK(clk), .D(u2__0root_452_0__418_), .Q(u2_o_417_));
DFFPOSX1 DFFPOSX1_423 ( .CLK(clk), .D(u2__0root_452_0__419_), .Q(u2_o_418_));
DFFPOSX1 DFFPOSX1_424 ( .CLK(clk), .D(u2__0root_452_0__420_), .Q(u2_o_419_));
DFFPOSX1 DFFPOSX1_425 ( .CLK(clk), .D(u2__0root_452_0__421_), .Q(u2_o_420_));
DFFPOSX1 DFFPOSX1_426 ( .CLK(clk), .D(u2__0root_452_0__422_), .Q(u2_o_421_));
DFFPOSX1 DFFPOSX1_427 ( .CLK(clk), .D(u2__0root_452_0__423_), .Q(u2_o_422_));
DFFPOSX1 DFFPOSX1_428 ( .CLK(clk), .D(u2__0root_452_0__424_), .Q(u2_o_423_));
DFFPOSX1 DFFPOSX1_429 ( .CLK(clk), .D(u2__0root_452_0__425_), .Q(u2_o_424_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk), .D(u2__0root_452_0__39_), .Q(sqrto_38_));
DFFPOSX1 DFFPOSX1_430 ( .CLK(clk), .D(u2__0root_452_0__426_), .Q(u2_o_425_));
DFFPOSX1 DFFPOSX1_431 ( .CLK(clk), .D(u2__0root_452_0__427_), .Q(u2_o_426_));
DFFPOSX1 DFFPOSX1_432 ( .CLK(clk), .D(u2__0root_452_0__428_), .Q(u2_o_427_));
DFFPOSX1 DFFPOSX1_433 ( .CLK(clk), .D(u2__0root_452_0__429_), .Q(u2_o_428_));
DFFPOSX1 DFFPOSX1_434 ( .CLK(clk), .D(u2__0root_452_0__430_), .Q(u2_o_429_));
DFFPOSX1 DFFPOSX1_435 ( .CLK(clk), .D(u2__0root_452_0__431_), .Q(u2_o_430_));
DFFPOSX1 DFFPOSX1_436 ( .CLK(clk), .D(u2__0root_452_0__432_), .Q(u2_o_431_));
DFFPOSX1 DFFPOSX1_437 ( .CLK(clk), .D(u2__0root_452_0__433_), .Q(u2_o_432_));
DFFPOSX1 DFFPOSX1_438 ( .CLK(clk), .D(u2__0root_452_0__434_), .Q(u2_o_433_));
DFFPOSX1 DFFPOSX1_439 ( .CLK(clk), .D(u2__0root_452_0__435_), .Q(u2_o_434_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk), .D(u2__0root_452_0__40_), .Q(sqrto_39_));
DFFPOSX1 DFFPOSX1_440 ( .CLK(clk), .D(u2__0root_452_0__436_), .Q(u2_o_435_));
DFFPOSX1 DFFPOSX1_441 ( .CLK(clk), .D(u2__0root_452_0__437_), .Q(u2_o_436_));
DFFPOSX1 DFFPOSX1_442 ( .CLK(clk), .D(u2__0root_452_0__438_), .Q(u2_o_437_));
DFFPOSX1 DFFPOSX1_443 ( .CLK(clk), .D(u2__0root_452_0__439_), .Q(u2_o_438_));
DFFPOSX1 DFFPOSX1_444 ( .CLK(clk), .D(u2__0root_452_0__440_), .Q(u2_o_439_));
DFFPOSX1 DFFPOSX1_445 ( .CLK(clk), .D(u2__0root_452_0__441_), .Q(u2_o_440_));
DFFPOSX1 DFFPOSX1_446 ( .CLK(clk), .D(u2__0root_452_0__442_), .Q(u2_o_441_));
DFFPOSX1 DFFPOSX1_447 ( .CLK(clk), .D(u2__0root_452_0__443_), .Q(u2_o_442_));
DFFPOSX1 DFFPOSX1_448 ( .CLK(clk), .D(u2__0root_452_0__444_), .Q(u2_o_443_));
DFFPOSX1 DFFPOSX1_449 ( .CLK(clk), .D(u2__0root_452_0__445_), .Q(u2_o_444_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk), .D(u2__0root_452_0__41_), .Q(sqrto_40_));
DFFPOSX1 DFFPOSX1_450 ( .CLK(clk), .D(u2__0root_452_0__446_), .Q(u2_o_445_));
DFFPOSX1 DFFPOSX1_451 ( .CLK(clk), .D(u2__0root_452_0__447_), .Q(u2_o_446_));
DFFPOSX1 DFFPOSX1_452 ( .CLK(clk), .D(u2__0root_452_0__448_), .Q(u2_o_447_));
DFFPOSX1 DFFPOSX1_453 ( .CLK(clk), .D(u2__0root_452_0__449_), .Q(u2_o_448_));
DFFPOSX1 DFFPOSX1_454 ( .CLK(clk), .D(u2__0root_452_0__450_), .Q(u2_o_449_));
DFFPOSX1 DFFPOSX1_455 ( .CLK(clk), .D(u2__0remLo_451_0__0_), .Q(u2_remLo_0_));
DFFPOSX1 DFFPOSX1_456 ( .CLK(clk), .D(u2__0remLo_451_0__1_), .Q(u2_remLo_1_));
DFFPOSX1 DFFPOSX1_457 ( .CLK(clk), .D(u2__0remLo_451_0__2_), .Q(u2_remLo_2_));
DFFPOSX1 DFFPOSX1_458 ( .CLK(clk), .D(u2__0remLo_451_0__3_), .Q(u2_remLo_3_));
DFFPOSX1 DFFPOSX1_459 ( .CLK(clk), .D(u2__0remLo_451_0__4_), .Q(u2_remLo_4_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk), .D(u2__0root_452_0__42_), .Q(sqrto_41_));
DFFPOSX1 DFFPOSX1_460 ( .CLK(clk), .D(u2__0remLo_451_0__5_), .Q(u2_remLo_5_));
DFFPOSX1 DFFPOSX1_461 ( .CLK(clk), .D(u2__0remLo_451_0__6_), .Q(u2_remLo_6_));
DFFPOSX1 DFFPOSX1_462 ( .CLK(clk), .D(u2__0remLo_451_0__7_), .Q(u2_remLo_7_));
DFFPOSX1 DFFPOSX1_463 ( .CLK(clk), .D(u2__0remLo_451_0__8_), .Q(u2_remLo_8_));
DFFPOSX1 DFFPOSX1_464 ( .CLK(clk), .D(u2__0remLo_451_0__9_), .Q(u2_remLo_9_));
DFFPOSX1 DFFPOSX1_465 ( .CLK(clk), .D(u2__0remLo_451_0__10_), .Q(u2_remLo_10_));
DFFPOSX1 DFFPOSX1_466 ( .CLK(clk), .D(u2__0remLo_451_0__11_), .Q(u2_remLo_11_));
DFFPOSX1 DFFPOSX1_467 ( .CLK(clk), .D(u2__0remLo_451_0__12_), .Q(u2_remLo_12_));
DFFPOSX1 DFFPOSX1_468 ( .CLK(clk), .D(u2__0remLo_451_0__13_), .Q(u2_remLo_13_));
DFFPOSX1 DFFPOSX1_469 ( .CLK(clk), .D(u2__0remLo_451_0__14_), .Q(u2_remLo_14_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk), .D(u2__0root_452_0__43_), .Q(sqrto_42_));
DFFPOSX1 DFFPOSX1_470 ( .CLK(clk), .D(u2__0remLo_451_0__15_), .Q(u2_remLo_15_));
DFFPOSX1 DFFPOSX1_471 ( .CLK(clk), .D(u2__0remLo_451_0__16_), .Q(u2_remLo_16_));
DFFPOSX1 DFFPOSX1_472 ( .CLK(clk), .D(u2__0remLo_451_0__17_), .Q(u2_remLo_17_));
DFFPOSX1 DFFPOSX1_473 ( .CLK(clk), .D(u2__0remLo_451_0__18_), .Q(u2_remLo_18_));
DFFPOSX1 DFFPOSX1_474 ( .CLK(clk), .D(u2__0remLo_451_0__19_), .Q(u2_remLo_19_));
DFFPOSX1 DFFPOSX1_475 ( .CLK(clk), .D(u2__0remLo_451_0__20_), .Q(u2_remLo_20_));
DFFPOSX1 DFFPOSX1_476 ( .CLK(clk), .D(u2__0remLo_451_0__21_), .Q(u2_remLo_21_));
DFFPOSX1 DFFPOSX1_477 ( .CLK(clk), .D(u2__0remLo_451_0__22_), .Q(u2_remLo_22_));
DFFPOSX1 DFFPOSX1_478 ( .CLK(clk), .D(u2__0remLo_451_0__23_), .Q(u2_remLo_23_));
DFFPOSX1 DFFPOSX1_479 ( .CLK(clk), .D(u2__0remLo_451_0__24_), .Q(u2_remLo_24_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk), .D(u2__0root_452_0__44_), .Q(sqrto_43_));
DFFPOSX1 DFFPOSX1_480 ( .CLK(clk), .D(u2__0remLo_451_0__25_), .Q(u2_remLo_25_));
DFFPOSX1 DFFPOSX1_481 ( .CLK(clk), .D(u2__0remLo_451_0__26_), .Q(u2_remLo_26_));
DFFPOSX1 DFFPOSX1_482 ( .CLK(clk), .D(u2__0remLo_451_0__27_), .Q(u2_remLo_27_));
DFFPOSX1 DFFPOSX1_483 ( .CLK(clk), .D(u2__0remLo_451_0__28_), .Q(u2_remLo_28_));
DFFPOSX1 DFFPOSX1_484 ( .CLK(clk), .D(u2__0remLo_451_0__29_), .Q(u2_remLo_29_));
DFFPOSX1 DFFPOSX1_485 ( .CLK(clk), .D(u2__0remLo_451_0__30_), .Q(u2_remLo_30_));
DFFPOSX1 DFFPOSX1_486 ( .CLK(clk), .D(u2__0remLo_451_0__31_), .Q(u2_remLo_31_));
DFFPOSX1 DFFPOSX1_487 ( .CLK(clk), .D(u2__0remLo_451_0__32_), .Q(u2_remLo_32_));
DFFPOSX1 DFFPOSX1_488 ( .CLK(clk), .D(u2__0remLo_451_0__33_), .Q(u2_remLo_33_));
DFFPOSX1 DFFPOSX1_489 ( .CLK(clk), .D(u2__0remLo_451_0__34_), .Q(u2_remLo_34_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk), .D(u2__0root_452_0__45_), .Q(sqrto_44_));
DFFPOSX1 DFFPOSX1_490 ( .CLK(clk), .D(u2__0remLo_451_0__35_), .Q(u2_remLo_35_));
DFFPOSX1 DFFPOSX1_491 ( .CLK(clk), .D(u2__0remLo_451_0__36_), .Q(u2_remLo_36_));
DFFPOSX1 DFFPOSX1_492 ( .CLK(clk), .D(u2__0remLo_451_0__37_), .Q(u2_remLo_37_));
DFFPOSX1 DFFPOSX1_493 ( .CLK(clk), .D(u2__0remLo_451_0__38_), .Q(u2_remLo_38_));
DFFPOSX1 DFFPOSX1_494 ( .CLK(clk), .D(u2__0remLo_451_0__39_), .Q(u2_remLo_39_));
DFFPOSX1 DFFPOSX1_495 ( .CLK(clk), .D(u2__0remLo_451_0__40_), .Q(u2_remLo_40_));
DFFPOSX1 DFFPOSX1_496 ( .CLK(clk), .D(u2__0remLo_451_0__41_), .Q(u2_remLo_41_));
DFFPOSX1 DFFPOSX1_497 ( .CLK(clk), .D(u2__0remLo_451_0__42_), .Q(u2_remLo_42_));
DFFPOSX1 DFFPOSX1_498 ( .CLK(clk), .D(u2__0remLo_451_0__43_), .Q(u2_remLo_43_));
DFFPOSX1 DFFPOSX1_499 ( .CLK(clk), .D(u2__0remLo_451_0__44_), .Q(u2_remLo_44_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(u2__0root_452_0__1_), .Q(sqrto_0_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk), .D(u2__0root_452_0__46_), .Q(sqrto_45_));
DFFPOSX1 DFFPOSX1_500 ( .CLK(clk), .D(u2__0remLo_451_0__45_), .Q(u2_remLo_45_));
DFFPOSX1 DFFPOSX1_501 ( .CLK(clk), .D(u2__0remLo_451_0__46_), .Q(u2_remLo_46_));
DFFPOSX1 DFFPOSX1_502 ( .CLK(clk), .D(u2__0remLo_451_0__47_), .Q(u2_remLo_47_));
DFFPOSX1 DFFPOSX1_503 ( .CLK(clk), .D(u2__0remLo_451_0__48_), .Q(u2_remLo_48_));
DFFPOSX1 DFFPOSX1_504 ( .CLK(clk), .D(u2__0remLo_451_0__49_), .Q(u2_remLo_49_));
DFFPOSX1 DFFPOSX1_505 ( .CLK(clk), .D(u2__0remLo_451_0__50_), .Q(u2_remLo_50_));
DFFPOSX1 DFFPOSX1_506 ( .CLK(clk), .D(u2__0remLo_451_0__51_), .Q(u2_remLo_51_));
DFFPOSX1 DFFPOSX1_507 ( .CLK(clk), .D(u2__0remLo_451_0__52_), .Q(u2_remLo_52_));
DFFPOSX1 DFFPOSX1_508 ( .CLK(clk), .D(u2__0remLo_451_0__53_), .Q(u2_remLo_53_));
DFFPOSX1 DFFPOSX1_509 ( .CLK(clk), .D(u2__0remLo_451_0__54_), .Q(u2_remLo_54_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk), .D(u2__0root_452_0__47_), .Q(sqrto_46_));
DFFPOSX1 DFFPOSX1_510 ( .CLK(clk), .D(u2__0remLo_451_0__55_), .Q(u2_remLo_55_));
DFFPOSX1 DFFPOSX1_511 ( .CLK(clk), .D(u2__0remLo_451_0__56_), .Q(u2_remLo_56_));
DFFPOSX1 DFFPOSX1_512 ( .CLK(clk), .D(u2__0remLo_451_0__57_), .Q(u2_remLo_57_));
DFFPOSX1 DFFPOSX1_513 ( .CLK(clk), .D(u2__0remLo_451_0__58_), .Q(u2_remLo_58_));
DFFPOSX1 DFFPOSX1_514 ( .CLK(clk), .D(u2__0remLo_451_0__59_), .Q(u2_remLo_59_));
DFFPOSX1 DFFPOSX1_515 ( .CLK(clk), .D(u2__0remLo_451_0__60_), .Q(u2_remLo_60_));
DFFPOSX1 DFFPOSX1_516 ( .CLK(clk), .D(u2__0remLo_451_0__61_), .Q(u2_remLo_61_));
DFFPOSX1 DFFPOSX1_517 ( .CLK(clk), .D(u2__0remLo_451_0__62_), .Q(u2_remLo_62_));
DFFPOSX1 DFFPOSX1_518 ( .CLK(clk), .D(u2__0remLo_451_0__63_), .Q(u2_remLo_63_));
DFFPOSX1 DFFPOSX1_519 ( .CLK(clk), .D(u2__0remLo_451_0__64_), .Q(u2_remLo_64_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk), .D(u2__0root_452_0__48_), .Q(sqrto_47_));
DFFPOSX1 DFFPOSX1_520 ( .CLK(clk), .D(u2__0remLo_451_0__65_), .Q(u2_remLo_65_));
DFFPOSX1 DFFPOSX1_521 ( .CLK(clk), .D(u2__0remLo_451_0__66_), .Q(u2_remLo_66_));
DFFPOSX1 DFFPOSX1_522 ( .CLK(clk), .D(u2__0remLo_451_0__67_), .Q(u2_remLo_67_));
DFFPOSX1 DFFPOSX1_523 ( .CLK(clk), .D(u2__0remLo_451_0__68_), .Q(u2_remLo_68_));
DFFPOSX1 DFFPOSX1_524 ( .CLK(clk), .D(u2__0remLo_451_0__69_), .Q(u2_remLo_69_));
DFFPOSX1 DFFPOSX1_525 ( .CLK(clk), .D(u2__0remLo_451_0__70_), .Q(u2_remLo_70_));
DFFPOSX1 DFFPOSX1_526 ( .CLK(clk), .D(u2__0remLo_451_0__71_), .Q(u2_remLo_71_));
DFFPOSX1 DFFPOSX1_527 ( .CLK(clk), .D(u2__0remLo_451_0__72_), .Q(u2_remLo_72_));
DFFPOSX1 DFFPOSX1_528 ( .CLK(clk), .D(u2__0remLo_451_0__73_), .Q(u2_remLo_73_));
DFFPOSX1 DFFPOSX1_529 ( .CLK(clk), .D(u2__0remLo_451_0__74_), .Q(u2_remLo_74_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk), .D(u2__0root_452_0__49_), .Q(sqrto_48_));
DFFPOSX1 DFFPOSX1_530 ( .CLK(clk), .D(u2__0remLo_451_0__75_), .Q(u2_remLo_75_));
DFFPOSX1 DFFPOSX1_531 ( .CLK(clk), .D(u2__0remLo_451_0__76_), .Q(u2_remLo_76_));
DFFPOSX1 DFFPOSX1_532 ( .CLK(clk), .D(u2__0remLo_451_0__77_), .Q(u2_remLo_77_));
DFFPOSX1 DFFPOSX1_533 ( .CLK(clk), .D(u2__0remLo_451_0__78_), .Q(u2_remLo_78_));
DFFPOSX1 DFFPOSX1_534 ( .CLK(clk), .D(u2__0remLo_451_0__79_), .Q(u2_remLo_79_));
DFFPOSX1 DFFPOSX1_535 ( .CLK(clk), .D(u2__0remLo_451_0__80_), .Q(u2_remLo_80_));
DFFPOSX1 DFFPOSX1_536 ( .CLK(clk), .D(u2__0remLo_451_0__81_), .Q(u2_remLo_81_));
DFFPOSX1 DFFPOSX1_537 ( .CLK(clk), .D(u2__0remLo_451_0__82_), .Q(u2_remLo_82_));
DFFPOSX1 DFFPOSX1_538 ( .CLK(clk), .D(u2__0remLo_451_0__83_), .Q(u2_remLo_83_));
DFFPOSX1 DFFPOSX1_539 ( .CLK(clk), .D(u2__0remLo_451_0__84_), .Q(u2_remLo_84_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk), .D(u2__0root_452_0__50_), .Q(sqrto_49_));
DFFPOSX1 DFFPOSX1_540 ( .CLK(clk), .D(u2__0remLo_451_0__85_), .Q(u2_remLo_85_));
DFFPOSX1 DFFPOSX1_541 ( .CLK(clk), .D(u2__0remLo_451_0__86_), .Q(u2_remLo_86_));
DFFPOSX1 DFFPOSX1_542 ( .CLK(clk), .D(u2__0remLo_451_0__87_), .Q(u2_remLo_87_));
DFFPOSX1 DFFPOSX1_543 ( .CLK(clk), .D(u2__0remLo_451_0__88_), .Q(u2_remLo_88_));
DFFPOSX1 DFFPOSX1_544 ( .CLK(clk), .D(u2__0remLo_451_0__89_), .Q(u2_remLo_89_));
DFFPOSX1 DFFPOSX1_545 ( .CLK(clk), .D(u2__0remLo_451_0__90_), .Q(u2_remLo_90_));
DFFPOSX1 DFFPOSX1_546 ( .CLK(clk), .D(u2__0remLo_451_0__91_), .Q(u2_remLo_91_));
DFFPOSX1 DFFPOSX1_547 ( .CLK(clk), .D(u2__0remLo_451_0__92_), .Q(u2_remLo_92_));
DFFPOSX1 DFFPOSX1_548 ( .CLK(clk), .D(u2__0remLo_451_0__93_), .Q(u2_remLo_93_));
DFFPOSX1 DFFPOSX1_549 ( .CLK(clk), .D(u2__0remLo_451_0__94_), .Q(u2_remLo_94_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk), .D(u2__0root_452_0__51_), .Q(sqrto_50_));
DFFPOSX1 DFFPOSX1_550 ( .CLK(clk), .D(u2__0remLo_451_0__95_), .Q(u2_remLo_95_));
DFFPOSX1 DFFPOSX1_551 ( .CLK(clk), .D(u2__0remLo_451_0__96_), .Q(u2_remLo_96_));
DFFPOSX1 DFFPOSX1_552 ( .CLK(clk), .D(u2__0remLo_451_0__97_), .Q(u2_remLo_97_));
DFFPOSX1 DFFPOSX1_553 ( .CLK(clk), .D(u2__0remLo_451_0__98_), .Q(u2_remLo_98_));
DFFPOSX1 DFFPOSX1_554 ( .CLK(clk), .D(u2__0remLo_451_0__99_), .Q(u2_remLo_99_));
DFFPOSX1 DFFPOSX1_555 ( .CLK(clk), .D(u2__0remLo_451_0__100_), .Q(u2_remLo_100_));
DFFPOSX1 DFFPOSX1_556 ( .CLK(clk), .D(u2__0remLo_451_0__101_), .Q(u2_remLo_101_));
DFFPOSX1 DFFPOSX1_557 ( .CLK(clk), .D(u2__0remLo_451_0__102_), .Q(u2_remLo_102_));
DFFPOSX1 DFFPOSX1_558 ( .CLK(clk), .D(u2__0remLo_451_0__103_), .Q(u2_remLo_103_));
DFFPOSX1 DFFPOSX1_559 ( .CLK(clk), .D(u2__0remLo_451_0__104_), .Q(u2_remLo_104_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk), .D(u2__0root_452_0__52_), .Q(sqrto_51_));
DFFPOSX1 DFFPOSX1_560 ( .CLK(clk), .D(u2__0remLo_451_0__105_), .Q(u2_remLo_105_));
DFFPOSX1 DFFPOSX1_561 ( .CLK(clk), .D(u2__0remLo_451_0__106_), .Q(u2_remLo_106_));
DFFPOSX1 DFFPOSX1_562 ( .CLK(clk), .D(u2__0remLo_451_0__107_), .Q(u2_remLo_107_));
DFFPOSX1 DFFPOSX1_563 ( .CLK(clk), .D(u2__0remLo_451_0__108_), .Q(u2_remLo_108_));
DFFPOSX1 DFFPOSX1_564 ( .CLK(clk), .D(u2__0remLo_451_0__109_), .Q(u2_remLo_109_));
DFFPOSX1 DFFPOSX1_565 ( .CLK(clk), .D(u2__0remLo_451_0__110_), .Q(u2_remLo_110_));
DFFPOSX1 DFFPOSX1_566 ( .CLK(clk), .D(u2__0remLo_451_0__111_), .Q(u2_remLo_111_));
DFFPOSX1 DFFPOSX1_567 ( .CLK(clk), .D(u2__0remLo_451_0__112_), .Q(u2_remLo_112_));
DFFPOSX1 DFFPOSX1_568 ( .CLK(clk), .D(u2__0remLo_451_0__113_), .Q(u2_remLo_113_));
DFFPOSX1 DFFPOSX1_569 ( .CLK(clk), .D(u2__0remLo_451_0__114_), .Q(u2_remLo_114_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk), .D(u2__0root_452_0__53_), .Q(sqrto_52_));
DFFPOSX1 DFFPOSX1_570 ( .CLK(clk), .D(u2__0remLo_451_0__115_), .Q(u2_remLo_115_));
DFFPOSX1 DFFPOSX1_571 ( .CLK(clk), .D(u2__0remLo_451_0__116_), .Q(u2_remLo_116_));
DFFPOSX1 DFFPOSX1_572 ( .CLK(clk), .D(u2__0remLo_451_0__117_), .Q(u2_remLo_117_));
DFFPOSX1 DFFPOSX1_573 ( .CLK(clk), .D(u2__0remLo_451_0__118_), .Q(u2_remLo_118_));
DFFPOSX1 DFFPOSX1_574 ( .CLK(clk), .D(u2__0remLo_451_0__119_), .Q(u2_remLo_119_));
DFFPOSX1 DFFPOSX1_575 ( .CLK(clk), .D(u2__0remLo_451_0__120_), .Q(u2_remLo_120_));
DFFPOSX1 DFFPOSX1_576 ( .CLK(clk), .D(u2__0remLo_451_0__121_), .Q(u2_remLo_121_));
DFFPOSX1 DFFPOSX1_577 ( .CLK(clk), .D(u2__0remLo_451_0__122_), .Q(u2_remLo_122_));
DFFPOSX1 DFFPOSX1_578 ( .CLK(clk), .D(u2__0remLo_451_0__123_), .Q(u2_remLo_123_));
DFFPOSX1 DFFPOSX1_579 ( .CLK(clk), .D(u2__0remLo_451_0__124_), .Q(u2_remLo_124_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk), .D(u2__0root_452_0__54_), .Q(sqrto_53_));
DFFPOSX1 DFFPOSX1_580 ( .CLK(clk), .D(u2__0remLo_451_0__125_), .Q(u2_remLo_125_));
DFFPOSX1 DFFPOSX1_581 ( .CLK(clk), .D(u2__0remLo_451_0__126_), .Q(u2_remLo_126_));
DFFPOSX1 DFFPOSX1_582 ( .CLK(clk), .D(u2__0remLo_451_0__127_), .Q(u2_remLo_127_));
DFFPOSX1 DFFPOSX1_583 ( .CLK(clk), .D(u2__0remLo_451_0__128_), .Q(u2_remLo_128_));
DFFPOSX1 DFFPOSX1_584 ( .CLK(clk), .D(u2__0remLo_451_0__129_), .Q(u2_remLo_129_));
DFFPOSX1 DFFPOSX1_585 ( .CLK(clk), .D(u2__0remLo_451_0__130_), .Q(u2_remLo_130_));
DFFPOSX1 DFFPOSX1_586 ( .CLK(clk), .D(u2__0remLo_451_0__131_), .Q(u2_remLo_131_));
DFFPOSX1 DFFPOSX1_587 ( .CLK(clk), .D(u2__0remLo_451_0__132_), .Q(u2_remLo_132_));
DFFPOSX1 DFFPOSX1_588 ( .CLK(clk), .D(u2__0remLo_451_0__133_), .Q(u2_remLo_133_));
DFFPOSX1 DFFPOSX1_589 ( .CLK(clk), .D(u2__0remLo_451_0__134_), .Q(u2_remLo_134_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk), .D(u2__0root_452_0__55_), .Q(sqrto_54_));
DFFPOSX1 DFFPOSX1_590 ( .CLK(clk), .D(u2__0remLo_451_0__135_), .Q(u2_remLo_135_));
DFFPOSX1 DFFPOSX1_591 ( .CLK(clk), .D(u2__0remLo_451_0__136_), .Q(u2_remLo_136_));
DFFPOSX1 DFFPOSX1_592 ( .CLK(clk), .D(u2__0remLo_451_0__137_), .Q(u2_remLo_137_));
DFFPOSX1 DFFPOSX1_593 ( .CLK(clk), .D(u2__0remLo_451_0__138_), .Q(u2_remLo_138_));
DFFPOSX1 DFFPOSX1_594 ( .CLK(clk), .D(u2__0remLo_451_0__139_), .Q(u2_remLo_139_));
DFFPOSX1 DFFPOSX1_595 ( .CLK(clk), .D(u2__0remLo_451_0__140_), .Q(u2_remLo_140_));
DFFPOSX1 DFFPOSX1_596 ( .CLK(clk), .D(u2__0remLo_451_0__141_), .Q(u2_remLo_141_));
DFFPOSX1 DFFPOSX1_597 ( .CLK(clk), .D(u2__0remLo_451_0__142_), .Q(u2_remLo_142_));
DFFPOSX1 DFFPOSX1_598 ( .CLK(clk), .D(u2__0remLo_451_0__143_), .Q(u2_remLo_143_));
DFFPOSX1 DFFPOSX1_599 ( .CLK(clk), .D(u2__0remLo_451_0__144_), .Q(u2_remLo_144_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(u2__0root_452_0__2_), .Q(sqrto_1_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk), .D(u2__0root_452_0__56_), .Q(sqrto_55_));
DFFPOSX1 DFFPOSX1_600 ( .CLK(clk), .D(u2__0remLo_451_0__145_), .Q(u2_remLo_145_));
DFFPOSX1 DFFPOSX1_601 ( .CLK(clk), .D(u2__0remLo_451_0__146_), .Q(u2_remLo_146_));
DFFPOSX1 DFFPOSX1_602 ( .CLK(clk), .D(u2__0remLo_451_0__147_), .Q(u2_remLo_147_));
DFFPOSX1 DFFPOSX1_603 ( .CLK(clk), .D(u2__0remLo_451_0__148_), .Q(u2_remLo_148_));
DFFPOSX1 DFFPOSX1_604 ( .CLK(clk), .D(u2__0remLo_451_0__149_), .Q(u2_remLo_149_));
DFFPOSX1 DFFPOSX1_605 ( .CLK(clk), .D(u2__0remLo_451_0__150_), .Q(u2_remLo_150_));
DFFPOSX1 DFFPOSX1_606 ( .CLK(clk), .D(u2__0remLo_451_0__151_), .Q(u2_remLo_151_));
DFFPOSX1 DFFPOSX1_607 ( .CLK(clk), .D(u2__0remLo_451_0__152_), .Q(u2_remLo_152_));
DFFPOSX1 DFFPOSX1_608 ( .CLK(clk), .D(u2__0remLo_451_0__153_), .Q(u2_remLo_153_));
DFFPOSX1 DFFPOSX1_609 ( .CLK(clk), .D(u2__0remLo_451_0__154_), .Q(u2_remLo_154_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk), .D(u2__0root_452_0__57_), .Q(sqrto_56_));
DFFPOSX1 DFFPOSX1_610 ( .CLK(clk), .D(u2__0remLo_451_0__155_), .Q(u2_remLo_155_));
DFFPOSX1 DFFPOSX1_611 ( .CLK(clk), .D(u2__0remLo_451_0__156_), .Q(u2_remLo_156_));
DFFPOSX1 DFFPOSX1_612 ( .CLK(clk), .D(u2__0remLo_451_0__157_), .Q(u2_remLo_157_));
DFFPOSX1 DFFPOSX1_613 ( .CLK(clk), .D(u2__0remLo_451_0__158_), .Q(u2_remLo_158_));
DFFPOSX1 DFFPOSX1_614 ( .CLK(clk), .D(u2__0remLo_451_0__159_), .Q(u2_remLo_159_));
DFFPOSX1 DFFPOSX1_615 ( .CLK(clk), .D(u2__0remLo_451_0__160_), .Q(u2_remLo_160_));
DFFPOSX1 DFFPOSX1_616 ( .CLK(clk), .D(u2__0remLo_451_0__161_), .Q(u2_remLo_161_));
DFFPOSX1 DFFPOSX1_617 ( .CLK(clk), .D(u2__0remLo_451_0__162_), .Q(u2_remLo_162_));
DFFPOSX1 DFFPOSX1_618 ( .CLK(clk), .D(u2__0remLo_451_0__163_), .Q(u2_remLo_163_));
DFFPOSX1 DFFPOSX1_619 ( .CLK(clk), .D(u2__0remLo_451_0__164_), .Q(u2_remLo_164_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk), .D(u2__0root_452_0__58_), .Q(sqrto_57_));
DFFPOSX1 DFFPOSX1_620 ( .CLK(clk), .D(u2__0remLo_451_0__165_), .Q(u2_remLo_165_));
DFFPOSX1 DFFPOSX1_621 ( .CLK(clk), .D(u2__0remLo_451_0__166_), .Q(u2_remLo_166_));
DFFPOSX1 DFFPOSX1_622 ( .CLK(clk), .D(u2__0remLo_451_0__167_), .Q(u2_remLo_167_));
DFFPOSX1 DFFPOSX1_623 ( .CLK(clk), .D(u2__0remLo_451_0__168_), .Q(u2_remLo_168_));
DFFPOSX1 DFFPOSX1_624 ( .CLK(clk), .D(u2__0remLo_451_0__169_), .Q(u2_remLo_169_));
DFFPOSX1 DFFPOSX1_625 ( .CLK(clk), .D(u2__0remLo_451_0__170_), .Q(u2_remLo_170_));
DFFPOSX1 DFFPOSX1_626 ( .CLK(clk), .D(u2__0remLo_451_0__171_), .Q(u2_remLo_171_));
DFFPOSX1 DFFPOSX1_627 ( .CLK(clk), .D(u2__0remLo_451_0__172_), .Q(u2_remLo_172_));
DFFPOSX1 DFFPOSX1_628 ( .CLK(clk), .D(u2__0remLo_451_0__173_), .Q(u2_remLo_173_));
DFFPOSX1 DFFPOSX1_629 ( .CLK(clk), .D(u2__0remLo_451_0__174_), .Q(u2_remLo_174_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk), .D(u2__0root_452_0__59_), .Q(sqrto_58_));
DFFPOSX1 DFFPOSX1_630 ( .CLK(clk), .D(u2__0remLo_451_0__175_), .Q(u2_remLo_175_));
DFFPOSX1 DFFPOSX1_631 ( .CLK(clk), .D(u2__0remLo_451_0__176_), .Q(u2_remLo_176_));
DFFPOSX1 DFFPOSX1_632 ( .CLK(clk), .D(u2__0remLo_451_0__177_), .Q(u2_remLo_177_));
DFFPOSX1 DFFPOSX1_633 ( .CLK(clk), .D(u2__0remLo_451_0__178_), .Q(u2_remLo_178_));
DFFPOSX1 DFFPOSX1_634 ( .CLK(clk), .D(u2__0remLo_451_0__179_), .Q(u2_remLo_179_));
DFFPOSX1 DFFPOSX1_635 ( .CLK(clk), .D(u2__0remLo_451_0__180_), .Q(u2_remLo_180_));
DFFPOSX1 DFFPOSX1_636 ( .CLK(clk), .D(u2__0remLo_451_0__181_), .Q(u2_remLo_181_));
DFFPOSX1 DFFPOSX1_637 ( .CLK(clk), .D(u2__0remLo_451_0__182_), .Q(u2_remLo_182_));
DFFPOSX1 DFFPOSX1_638 ( .CLK(clk), .D(u2__0remLo_451_0__183_), .Q(u2_remLo_183_));
DFFPOSX1 DFFPOSX1_639 ( .CLK(clk), .D(u2__0remLo_451_0__184_), .Q(u2_remLo_184_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk), .D(u2__0root_452_0__60_), .Q(sqrto_59_));
DFFPOSX1 DFFPOSX1_640 ( .CLK(clk), .D(u2__0remLo_451_0__185_), .Q(u2_remLo_185_));
DFFPOSX1 DFFPOSX1_641 ( .CLK(clk), .D(u2__0remLo_451_0__186_), .Q(u2_remLo_186_));
DFFPOSX1 DFFPOSX1_642 ( .CLK(clk), .D(u2__0remLo_451_0__187_), .Q(u2_remLo_187_));
DFFPOSX1 DFFPOSX1_643 ( .CLK(clk), .D(u2__0remLo_451_0__188_), .Q(u2_remLo_188_));
DFFPOSX1 DFFPOSX1_644 ( .CLK(clk), .D(u2__0remLo_451_0__189_), .Q(u2_remLo_189_));
DFFPOSX1 DFFPOSX1_645 ( .CLK(clk), .D(u2__0remLo_451_0__190_), .Q(u2_remLo_190_));
DFFPOSX1 DFFPOSX1_646 ( .CLK(clk), .D(u2__0remLo_451_0__191_), .Q(u2_remLo_191_));
DFFPOSX1 DFFPOSX1_647 ( .CLK(clk), .D(u2__0remLo_451_0__192_), .Q(u2_remLo_192_));
DFFPOSX1 DFFPOSX1_648 ( .CLK(clk), .D(u2__0remLo_451_0__193_), .Q(u2_remLo_193_));
DFFPOSX1 DFFPOSX1_649 ( .CLK(clk), .D(u2__0remLo_451_0__194_), .Q(u2_remLo_194_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk), .D(u2__0root_452_0__61_), .Q(sqrto_60_));
DFFPOSX1 DFFPOSX1_650 ( .CLK(clk), .D(u2__0remLo_451_0__195_), .Q(u2_remLo_195_));
DFFPOSX1 DFFPOSX1_651 ( .CLK(clk), .D(u2__0remLo_451_0__196_), .Q(u2_remLo_196_));
DFFPOSX1 DFFPOSX1_652 ( .CLK(clk), .D(u2__0remLo_451_0__197_), .Q(u2_remLo_197_));
DFFPOSX1 DFFPOSX1_653 ( .CLK(clk), .D(u2__0remLo_451_0__198_), .Q(u2_remLo_198_));
DFFPOSX1 DFFPOSX1_654 ( .CLK(clk), .D(u2__0remLo_451_0__199_), .Q(u2_remLo_199_));
DFFPOSX1 DFFPOSX1_655 ( .CLK(clk), .D(u2__0remLo_451_0__200_), .Q(u2_remLo_200_));
DFFPOSX1 DFFPOSX1_656 ( .CLK(clk), .D(u2__0remLo_451_0__201_), .Q(u2_remLo_201_));
DFFPOSX1 DFFPOSX1_657 ( .CLK(clk), .D(u2__0remLo_451_0__202_), .Q(u2_remLo_202_));
DFFPOSX1 DFFPOSX1_658 ( .CLK(clk), .D(u2__0remLo_451_0__203_), .Q(u2_remLo_203_));
DFFPOSX1 DFFPOSX1_659 ( .CLK(clk), .D(u2__0remLo_451_0__204_), .Q(u2_remLo_204_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk), .D(u2__0root_452_0__62_), .Q(sqrto_61_));
DFFPOSX1 DFFPOSX1_660 ( .CLK(clk), .D(u2__0remLo_451_0__205_), .Q(u2_remLo_205_));
DFFPOSX1 DFFPOSX1_661 ( .CLK(clk), .D(u2__0remLo_451_0__206_), .Q(u2_remLo_206_));
DFFPOSX1 DFFPOSX1_662 ( .CLK(clk), .D(u2__0remLo_451_0__207_), .Q(u2_remLo_207_));
DFFPOSX1 DFFPOSX1_663 ( .CLK(clk), .D(u2__0remLo_451_0__208_), .Q(u2_remLo_208_));
DFFPOSX1 DFFPOSX1_664 ( .CLK(clk), .D(u2__0remLo_451_0__209_), .Q(u2_remLo_209_));
DFFPOSX1 DFFPOSX1_665 ( .CLK(clk), .D(u2__0remLo_451_0__210_), .Q(u2_remLo_210_));
DFFPOSX1 DFFPOSX1_666 ( .CLK(clk), .D(u2__0remLo_451_0__211_), .Q(u2_remLo_211_));
DFFPOSX1 DFFPOSX1_667 ( .CLK(clk), .D(u2__0remLo_451_0__212_), .Q(u2_remLo_212_));
DFFPOSX1 DFFPOSX1_668 ( .CLK(clk), .D(u2__0remLo_451_0__213_), .Q(u2_remLo_213_));
DFFPOSX1 DFFPOSX1_669 ( .CLK(clk), .D(u2__0remLo_451_0__214_), .Q(u2_remLo_214_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk), .D(u2__0root_452_0__63_), .Q(sqrto_62_));
DFFPOSX1 DFFPOSX1_670 ( .CLK(clk), .D(u2__0remLo_451_0__215_), .Q(u2_remLo_215_));
DFFPOSX1 DFFPOSX1_671 ( .CLK(clk), .D(u2__0remLo_451_0__216_), .Q(u2_remLo_216_));
DFFPOSX1 DFFPOSX1_672 ( .CLK(clk), .D(u2__0remLo_451_0__217_), .Q(u2_remLo_217_));
DFFPOSX1 DFFPOSX1_673 ( .CLK(clk), .D(u2__0remLo_451_0__218_), .Q(u2_remLo_218_));
DFFPOSX1 DFFPOSX1_674 ( .CLK(clk), .D(u2__0remLo_451_0__219_), .Q(u2_remLo_219_));
DFFPOSX1 DFFPOSX1_675 ( .CLK(clk), .D(u2__0remLo_451_0__220_), .Q(u2_remLo_220_));
DFFPOSX1 DFFPOSX1_676 ( .CLK(clk), .D(u2__0remLo_451_0__221_), .Q(u2_remLo_221_));
DFFPOSX1 DFFPOSX1_677 ( .CLK(clk), .D(u2__0remLo_451_0__222_), .Q(u2_remLo_222_));
DFFPOSX1 DFFPOSX1_678 ( .CLK(clk), .D(u2__0remLo_451_0__223_), .Q(u2_remLo_223_));
DFFPOSX1 DFFPOSX1_679 ( .CLK(clk), .D(u2__0remLo_451_0__224_), .Q(u2_remLo_224_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk), .D(u2__0root_452_0__64_), .Q(sqrto_63_));
DFFPOSX1 DFFPOSX1_680 ( .CLK(clk), .D(u2__0remLo_451_0__225_), .Q(u2_remLo_225_));
DFFPOSX1 DFFPOSX1_681 ( .CLK(clk), .D(u2__0remLo_451_0__226_), .Q(u2_remLo_226_));
DFFPOSX1 DFFPOSX1_682 ( .CLK(clk), .D(u2__0remLo_451_0__227_), .Q(u2_remLo_227_));
DFFPOSX1 DFFPOSX1_683 ( .CLK(clk), .D(u2__0remLo_451_0__228_), .Q(u2_remLo_228_));
DFFPOSX1 DFFPOSX1_684 ( .CLK(clk), .D(u2__0remLo_451_0__229_), .Q(u2_remLo_229_));
DFFPOSX1 DFFPOSX1_685 ( .CLK(clk), .D(u2__0remLo_451_0__230_), .Q(u2_remLo_230_));
DFFPOSX1 DFFPOSX1_686 ( .CLK(clk), .D(u2__0remLo_451_0__231_), .Q(u2_remLo_231_));
DFFPOSX1 DFFPOSX1_687 ( .CLK(clk), .D(u2__0remLo_451_0__232_), .Q(u2_remLo_232_));
DFFPOSX1 DFFPOSX1_688 ( .CLK(clk), .D(u2__0remLo_451_0__233_), .Q(u2_remLo_233_));
DFFPOSX1 DFFPOSX1_689 ( .CLK(clk), .D(u2__0remLo_451_0__234_), .Q(u2_remLo_234_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk), .D(u2__0root_452_0__65_), .Q(sqrto_64_));
DFFPOSX1 DFFPOSX1_690 ( .CLK(clk), .D(u2__0remLo_451_0__235_), .Q(u2_remLo_235_));
DFFPOSX1 DFFPOSX1_691 ( .CLK(clk), .D(u2__0remLo_451_0__236_), .Q(u2_remLo_236_));
DFFPOSX1 DFFPOSX1_692 ( .CLK(clk), .D(u2__0remLo_451_0__237_), .Q(u2_remLo_237_));
DFFPOSX1 DFFPOSX1_693 ( .CLK(clk), .D(u2__0remLo_451_0__238_), .Q(u2_remLo_238_));
DFFPOSX1 DFFPOSX1_694 ( .CLK(clk), .D(u2__0remLo_451_0__239_), .Q(u2_remLo_239_));
DFFPOSX1 DFFPOSX1_695 ( .CLK(clk), .D(u2__0remLo_451_0__240_), .Q(u2_remLo_240_));
DFFPOSX1 DFFPOSX1_696 ( .CLK(clk), .D(u2__0remLo_451_0__241_), .Q(u2_remLo_241_));
DFFPOSX1 DFFPOSX1_697 ( .CLK(clk), .D(u2__0remLo_451_0__242_), .Q(u2_remLo_242_));
DFFPOSX1 DFFPOSX1_698 ( .CLK(clk), .D(u2__0remLo_451_0__243_), .Q(u2_remLo_243_));
DFFPOSX1 DFFPOSX1_699 ( .CLK(clk), .D(u2__0remLo_451_0__244_), .Q(u2_remLo_244_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(u2__0root_452_0__3_), .Q(sqrto_2_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk), .D(u2__0root_452_0__66_), .Q(sqrto_65_));
DFFPOSX1 DFFPOSX1_700 ( .CLK(clk), .D(u2__0remLo_451_0__245_), .Q(u2_remLo_245_));
DFFPOSX1 DFFPOSX1_701 ( .CLK(clk), .D(u2__0remLo_451_0__246_), .Q(u2_remLo_246_));
DFFPOSX1 DFFPOSX1_702 ( .CLK(clk), .D(u2__0remLo_451_0__247_), .Q(u2_remLo_247_));
DFFPOSX1 DFFPOSX1_703 ( .CLK(clk), .D(u2__0remLo_451_0__248_), .Q(u2_remLo_248_));
DFFPOSX1 DFFPOSX1_704 ( .CLK(clk), .D(u2__0remLo_451_0__249_), .Q(u2_remLo_249_));
DFFPOSX1 DFFPOSX1_705 ( .CLK(clk), .D(u2__0remLo_451_0__250_), .Q(u2_remLo_250_));
DFFPOSX1 DFFPOSX1_706 ( .CLK(clk), .D(u2__0remLo_451_0__251_), .Q(u2_remLo_251_));
DFFPOSX1 DFFPOSX1_707 ( .CLK(clk), .D(u2__0remLo_451_0__252_), .Q(u2_remLo_252_));
DFFPOSX1 DFFPOSX1_708 ( .CLK(clk), .D(u2__0remLo_451_0__253_), .Q(u2_remLo_253_));
DFFPOSX1 DFFPOSX1_709 ( .CLK(clk), .D(u2__0remLo_451_0__254_), .Q(u2_remLo_254_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk), .D(u2__0root_452_0__67_), .Q(sqrto_66_));
DFFPOSX1 DFFPOSX1_710 ( .CLK(clk), .D(u2__0remLo_451_0__255_), .Q(u2_remLo_255_));
DFFPOSX1 DFFPOSX1_711 ( .CLK(clk), .D(u2__0remLo_451_0__256_), .Q(u2_remLo_256_));
DFFPOSX1 DFFPOSX1_712 ( .CLK(clk), .D(u2__0remLo_451_0__257_), .Q(u2_remLo_257_));
DFFPOSX1 DFFPOSX1_713 ( .CLK(clk), .D(u2__0remLo_451_0__258_), .Q(u2_remLo_258_));
DFFPOSX1 DFFPOSX1_714 ( .CLK(clk), .D(u2__0remLo_451_0__259_), .Q(u2_remLo_259_));
DFFPOSX1 DFFPOSX1_715 ( .CLK(clk), .D(u2__0remLo_451_0__260_), .Q(u2_remLo_260_));
DFFPOSX1 DFFPOSX1_716 ( .CLK(clk), .D(u2__0remLo_451_0__261_), .Q(u2_remLo_261_));
DFFPOSX1 DFFPOSX1_717 ( .CLK(clk), .D(u2__0remLo_451_0__262_), .Q(u2_remLo_262_));
DFFPOSX1 DFFPOSX1_718 ( .CLK(clk), .D(u2__0remLo_451_0__263_), .Q(u2_remLo_263_));
DFFPOSX1 DFFPOSX1_719 ( .CLK(clk), .D(u2__0remLo_451_0__264_), .Q(u2_remLo_264_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk), .D(u2__0root_452_0__68_), .Q(sqrto_67_));
DFFPOSX1 DFFPOSX1_720 ( .CLK(clk), .D(u2__0remLo_451_0__265_), .Q(u2_remLo_265_));
DFFPOSX1 DFFPOSX1_721 ( .CLK(clk), .D(u2__0remLo_451_0__266_), .Q(u2_remLo_266_));
DFFPOSX1 DFFPOSX1_722 ( .CLK(clk), .D(u2__0remLo_451_0__267_), .Q(u2_remLo_267_));
DFFPOSX1 DFFPOSX1_723 ( .CLK(clk), .D(u2__0remLo_451_0__268_), .Q(u2_remLo_268_));
DFFPOSX1 DFFPOSX1_724 ( .CLK(clk), .D(u2__0remLo_451_0__269_), .Q(u2_remLo_269_));
DFFPOSX1 DFFPOSX1_725 ( .CLK(clk), .D(u2__0remLo_451_0__270_), .Q(u2_remLo_270_));
DFFPOSX1 DFFPOSX1_726 ( .CLK(clk), .D(u2__0remLo_451_0__271_), .Q(u2_remLo_271_));
DFFPOSX1 DFFPOSX1_727 ( .CLK(clk), .D(u2__0remLo_451_0__272_), .Q(u2_remLo_272_));
DFFPOSX1 DFFPOSX1_728 ( .CLK(clk), .D(u2__0remLo_451_0__273_), .Q(u2_remLo_273_));
DFFPOSX1 DFFPOSX1_729 ( .CLK(clk), .D(u2__0remLo_451_0__274_), .Q(u2_remLo_274_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk), .D(u2__0root_452_0__69_), .Q(sqrto_68_));
DFFPOSX1 DFFPOSX1_730 ( .CLK(clk), .D(u2__0remLo_451_0__275_), .Q(u2_remLo_275_));
DFFPOSX1 DFFPOSX1_731 ( .CLK(clk), .D(u2__0remLo_451_0__276_), .Q(u2_remLo_276_));
DFFPOSX1 DFFPOSX1_732 ( .CLK(clk), .D(u2__0remLo_451_0__277_), .Q(u2_remLo_277_));
DFFPOSX1 DFFPOSX1_733 ( .CLK(clk), .D(u2__0remLo_451_0__278_), .Q(u2_remLo_278_));
DFFPOSX1 DFFPOSX1_734 ( .CLK(clk), .D(u2__0remLo_451_0__279_), .Q(u2_remLo_279_));
DFFPOSX1 DFFPOSX1_735 ( .CLK(clk), .D(u2__0remLo_451_0__280_), .Q(u2_remLo_280_));
DFFPOSX1 DFFPOSX1_736 ( .CLK(clk), .D(u2__0remLo_451_0__281_), .Q(u2_remLo_281_));
DFFPOSX1 DFFPOSX1_737 ( .CLK(clk), .D(u2__0remLo_451_0__282_), .Q(u2_remLo_282_));
DFFPOSX1 DFFPOSX1_738 ( .CLK(clk), .D(u2__0remLo_451_0__283_), .Q(u2_remLo_283_));
DFFPOSX1 DFFPOSX1_739 ( .CLK(clk), .D(u2__0remLo_451_0__284_), .Q(u2_remLo_284_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk), .D(u2__0root_452_0__70_), .Q(sqrto_69_));
DFFPOSX1 DFFPOSX1_740 ( .CLK(clk), .D(u2__0remLo_451_0__285_), .Q(u2_remLo_285_));
DFFPOSX1 DFFPOSX1_741 ( .CLK(clk), .D(u2__0remLo_451_0__286_), .Q(u2_remLo_286_));
DFFPOSX1 DFFPOSX1_742 ( .CLK(clk), .D(u2__0remLo_451_0__287_), .Q(u2_remLo_287_));
DFFPOSX1 DFFPOSX1_743 ( .CLK(clk), .D(u2__0remLo_451_0__288_), .Q(u2_remLo_288_));
DFFPOSX1 DFFPOSX1_744 ( .CLK(clk), .D(u2__0remLo_451_0__289_), .Q(u2_remLo_289_));
DFFPOSX1 DFFPOSX1_745 ( .CLK(clk), .D(u2__0remLo_451_0__290_), .Q(u2_remLo_290_));
DFFPOSX1 DFFPOSX1_746 ( .CLK(clk), .D(u2__0remLo_451_0__291_), .Q(u2_remLo_291_));
DFFPOSX1 DFFPOSX1_747 ( .CLK(clk), .D(u2__0remLo_451_0__292_), .Q(u2_remLo_292_));
DFFPOSX1 DFFPOSX1_748 ( .CLK(clk), .D(u2__0remLo_451_0__293_), .Q(u2_remLo_293_));
DFFPOSX1 DFFPOSX1_749 ( .CLK(clk), .D(u2__0remLo_451_0__294_), .Q(u2_remLo_294_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk), .D(u2__0root_452_0__71_), .Q(sqrto_70_));
DFFPOSX1 DFFPOSX1_750 ( .CLK(clk), .D(u2__0remLo_451_0__295_), .Q(u2_remLo_295_));
DFFPOSX1 DFFPOSX1_751 ( .CLK(clk), .D(u2__0remLo_451_0__296_), .Q(u2_remLo_296_));
DFFPOSX1 DFFPOSX1_752 ( .CLK(clk), .D(u2__0remLo_451_0__297_), .Q(u2_remLo_297_));
DFFPOSX1 DFFPOSX1_753 ( .CLK(clk), .D(u2__0remLo_451_0__298_), .Q(u2_remLo_298_));
DFFPOSX1 DFFPOSX1_754 ( .CLK(clk), .D(u2__0remLo_451_0__299_), .Q(u2_remLo_299_));
DFFPOSX1 DFFPOSX1_755 ( .CLK(clk), .D(u2__0remLo_451_0__300_), .Q(u2_remLo_300_));
DFFPOSX1 DFFPOSX1_756 ( .CLK(clk), .D(u2__0remLo_451_0__301_), .Q(u2_remLo_301_));
DFFPOSX1 DFFPOSX1_757 ( .CLK(clk), .D(u2__0remLo_451_0__302_), .Q(u2_remLo_302_));
DFFPOSX1 DFFPOSX1_758 ( .CLK(clk), .D(u2__0remLo_451_0__303_), .Q(u2_remLo_303_));
DFFPOSX1 DFFPOSX1_759 ( .CLK(clk), .D(u2__0remLo_451_0__304_), .Q(u2_remLo_304_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk), .D(u2__0root_452_0__72_), .Q(sqrto_71_));
DFFPOSX1 DFFPOSX1_760 ( .CLK(clk), .D(u2__0remLo_451_0__305_), .Q(u2_remLo_305_));
DFFPOSX1 DFFPOSX1_761 ( .CLK(clk), .D(u2__0remLo_451_0__306_), .Q(u2_remLo_306_));
DFFPOSX1 DFFPOSX1_762 ( .CLK(clk), .D(u2__0remLo_451_0__307_), .Q(u2_remLo_307_));
DFFPOSX1 DFFPOSX1_763 ( .CLK(clk), .D(u2__0remLo_451_0__308_), .Q(u2_remLo_308_));
DFFPOSX1 DFFPOSX1_764 ( .CLK(clk), .D(u2__0remLo_451_0__309_), .Q(u2_remLo_309_));
DFFPOSX1 DFFPOSX1_765 ( .CLK(clk), .D(u2__0remLo_451_0__310_), .Q(u2_remLo_310_));
DFFPOSX1 DFFPOSX1_766 ( .CLK(clk), .D(u2__0remLo_451_0__311_), .Q(u2_remLo_311_));
DFFPOSX1 DFFPOSX1_767 ( .CLK(clk), .D(u2__0remLo_451_0__312_), .Q(u2_remLo_312_));
DFFPOSX1 DFFPOSX1_768 ( .CLK(clk), .D(u2__0remLo_451_0__313_), .Q(u2_remLo_313_));
DFFPOSX1 DFFPOSX1_769 ( .CLK(clk), .D(u2__0remLo_451_0__314_), .Q(u2_remLo_314_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk), .D(u2__0root_452_0__73_), .Q(sqrto_72_));
DFFPOSX1 DFFPOSX1_770 ( .CLK(clk), .D(u2__0remLo_451_0__315_), .Q(u2_remLo_315_));
DFFPOSX1 DFFPOSX1_771 ( .CLK(clk), .D(u2__0remLo_451_0__316_), .Q(u2_remLo_316_));
DFFPOSX1 DFFPOSX1_772 ( .CLK(clk), .D(u2__0remLo_451_0__317_), .Q(u2_remLo_317_));
DFFPOSX1 DFFPOSX1_773 ( .CLK(clk), .D(u2__0remLo_451_0__318_), .Q(u2_remLo_318_));
DFFPOSX1 DFFPOSX1_774 ( .CLK(clk), .D(u2__0remLo_451_0__319_), .Q(u2_remLo_319_));
DFFPOSX1 DFFPOSX1_775 ( .CLK(clk), .D(u2__0remLo_451_0__320_), .Q(u2_remLo_320_));
DFFPOSX1 DFFPOSX1_776 ( .CLK(clk), .D(u2__0remLo_451_0__321_), .Q(u2_remLo_321_));
DFFPOSX1 DFFPOSX1_777 ( .CLK(clk), .D(u2__0remLo_451_0__322_), .Q(u2_remLo_322_));
DFFPOSX1 DFFPOSX1_778 ( .CLK(clk), .D(u2__0remLo_451_0__323_), .Q(u2_remLo_323_));
DFFPOSX1 DFFPOSX1_779 ( .CLK(clk), .D(u2__0remLo_451_0__324_), .Q(u2_remLo_324_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk), .D(u2__0root_452_0__74_), .Q(sqrto_73_));
DFFPOSX1 DFFPOSX1_780 ( .CLK(clk), .D(u2__0remLo_451_0__325_), .Q(u2_remLo_325_));
DFFPOSX1 DFFPOSX1_781 ( .CLK(clk), .D(u2__0remLo_451_0__326_), .Q(u2_remLo_326_));
DFFPOSX1 DFFPOSX1_782 ( .CLK(clk), .D(u2__0remLo_451_0__327_), .Q(u2_remLo_327_));
DFFPOSX1 DFFPOSX1_783 ( .CLK(clk), .D(u2__0remLo_451_0__328_), .Q(u2_remLo_328_));
DFFPOSX1 DFFPOSX1_784 ( .CLK(clk), .D(u2__0remLo_451_0__329_), .Q(u2_remLo_329_));
DFFPOSX1 DFFPOSX1_785 ( .CLK(clk), .D(u2__0remLo_451_0__330_), .Q(u2_remLo_330_));
DFFPOSX1 DFFPOSX1_786 ( .CLK(clk), .D(u2__0remLo_451_0__331_), .Q(u2_remLo_331_));
DFFPOSX1 DFFPOSX1_787 ( .CLK(clk), .D(u2__0remLo_451_0__332_), .Q(u2_remLo_332_));
DFFPOSX1 DFFPOSX1_788 ( .CLK(clk), .D(u2__0remLo_451_0__333_), .Q(u2_remLo_333_));
DFFPOSX1 DFFPOSX1_789 ( .CLK(clk), .D(u2__0remLo_451_0__334_), .Q(u2_remLo_334_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk), .D(u2__0root_452_0__75_), .Q(sqrto_74_));
DFFPOSX1 DFFPOSX1_790 ( .CLK(clk), .D(u2__0remLo_451_0__335_), .Q(u2_remLo_335_));
DFFPOSX1 DFFPOSX1_791 ( .CLK(clk), .D(u2__0remLo_451_0__336_), .Q(u2_remLo_336_));
DFFPOSX1 DFFPOSX1_792 ( .CLK(clk), .D(u2__0remLo_451_0__337_), .Q(u2_remLo_337_));
DFFPOSX1 DFFPOSX1_793 ( .CLK(clk), .D(u2__0remLo_451_0__338_), .Q(u2_remLo_338_));
DFFPOSX1 DFFPOSX1_794 ( .CLK(clk), .D(u2__0remLo_451_0__339_), .Q(u2_remLo_339_));
DFFPOSX1 DFFPOSX1_795 ( .CLK(clk), .D(u2__0remLo_451_0__340_), .Q(u2_remLo_340_));
DFFPOSX1 DFFPOSX1_796 ( .CLK(clk), .D(u2__0remLo_451_0__341_), .Q(u2_remLo_341_));
DFFPOSX1 DFFPOSX1_797 ( .CLK(clk), .D(u2__0remLo_451_0__342_), .Q(u2_remLo_342_));
DFFPOSX1 DFFPOSX1_798 ( .CLK(clk), .D(u2__0remLo_451_0__343_), .Q(u2_remLo_343_));
DFFPOSX1 DFFPOSX1_799 ( .CLK(clk), .D(u2__0remLo_451_0__344_), .Q(u2_remLo_344_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(u2__0root_452_0__4_), .Q(sqrto_3_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk), .D(u2__0root_452_0__76_), .Q(sqrto_75_));
DFFPOSX1 DFFPOSX1_800 ( .CLK(clk), .D(u2__0remLo_451_0__345_), .Q(u2_remLo_345_));
DFFPOSX1 DFFPOSX1_801 ( .CLK(clk), .D(u2__0remLo_451_0__346_), .Q(u2_remLo_346_));
DFFPOSX1 DFFPOSX1_802 ( .CLK(clk), .D(u2__0remLo_451_0__347_), .Q(u2_remLo_347_));
DFFPOSX1 DFFPOSX1_803 ( .CLK(clk), .D(u2__0remLo_451_0__348_), .Q(u2_remLo_348_));
DFFPOSX1 DFFPOSX1_804 ( .CLK(clk), .D(u2__0remLo_451_0__349_), .Q(u2_remLo_349_));
DFFPOSX1 DFFPOSX1_805 ( .CLK(clk), .D(u2__0remLo_451_0__350_), .Q(u2_remLo_350_));
DFFPOSX1 DFFPOSX1_806 ( .CLK(clk), .D(u2__0remLo_451_0__351_), .Q(u2_remLo_351_));
DFFPOSX1 DFFPOSX1_807 ( .CLK(clk), .D(u2__0remLo_451_0__352_), .Q(u2_remLo_352_));
DFFPOSX1 DFFPOSX1_808 ( .CLK(clk), .D(u2__0remLo_451_0__353_), .Q(u2_remLo_353_));
DFFPOSX1 DFFPOSX1_809 ( .CLK(clk), .D(u2__0remLo_451_0__354_), .Q(u2_remLo_354_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk), .D(u2__0root_452_0__77_), .Q(sqrto_76_));
DFFPOSX1 DFFPOSX1_810 ( .CLK(clk), .D(u2__0remLo_451_0__355_), .Q(u2_remLo_355_));
DFFPOSX1 DFFPOSX1_811 ( .CLK(clk), .D(u2__0remLo_451_0__356_), .Q(u2_remLo_356_));
DFFPOSX1 DFFPOSX1_812 ( .CLK(clk), .D(u2__0remLo_451_0__357_), .Q(u2_remLo_357_));
DFFPOSX1 DFFPOSX1_813 ( .CLK(clk), .D(u2__0remLo_451_0__358_), .Q(u2_remLo_358_));
DFFPOSX1 DFFPOSX1_814 ( .CLK(clk), .D(u2__0remLo_451_0__359_), .Q(u2_remLo_359_));
DFFPOSX1 DFFPOSX1_815 ( .CLK(clk), .D(u2__0remLo_451_0__360_), .Q(u2_remLo_360_));
DFFPOSX1 DFFPOSX1_816 ( .CLK(clk), .D(u2__0remLo_451_0__361_), .Q(u2_remLo_361_));
DFFPOSX1 DFFPOSX1_817 ( .CLK(clk), .D(u2__0remLo_451_0__362_), .Q(u2_remLo_362_));
DFFPOSX1 DFFPOSX1_818 ( .CLK(clk), .D(u2__0remLo_451_0__363_), .Q(u2_remLo_363_));
DFFPOSX1 DFFPOSX1_819 ( .CLK(clk), .D(u2__0remLo_451_0__364_), .Q(u2_remLo_364_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk), .D(u2__0root_452_0__78_), .Q(sqrto_77_));
DFFPOSX1 DFFPOSX1_820 ( .CLK(clk), .D(u2__0remLo_451_0__365_), .Q(u2_remLo_365_));
DFFPOSX1 DFFPOSX1_821 ( .CLK(clk), .D(u2__0remLo_451_0__366_), .Q(u2_remLo_366_));
DFFPOSX1 DFFPOSX1_822 ( .CLK(clk), .D(u2__0remLo_451_0__367_), .Q(u2_remLo_367_));
DFFPOSX1 DFFPOSX1_823 ( .CLK(clk), .D(u2__0remLo_451_0__368_), .Q(u2_remLo_368_));
DFFPOSX1 DFFPOSX1_824 ( .CLK(clk), .D(u2__0remLo_451_0__369_), .Q(u2_remLo_369_));
DFFPOSX1 DFFPOSX1_825 ( .CLK(clk), .D(u2__0remLo_451_0__370_), .Q(u2_remLo_370_));
DFFPOSX1 DFFPOSX1_826 ( .CLK(clk), .D(u2__0remLo_451_0__371_), .Q(u2_remLo_371_));
DFFPOSX1 DFFPOSX1_827 ( .CLK(clk), .D(u2__0remLo_451_0__372_), .Q(u2_remLo_372_));
DFFPOSX1 DFFPOSX1_828 ( .CLK(clk), .D(u2__0remLo_451_0__373_), .Q(u2_remLo_373_));
DFFPOSX1 DFFPOSX1_829 ( .CLK(clk), .D(u2__0remLo_451_0__374_), .Q(u2_remLo_374_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk), .D(u2__0root_452_0__79_), .Q(sqrto_78_));
DFFPOSX1 DFFPOSX1_830 ( .CLK(clk), .D(u2__0remLo_451_0__375_), .Q(u2_remLo_375_));
DFFPOSX1 DFFPOSX1_831 ( .CLK(clk), .D(u2__0remLo_451_0__376_), .Q(u2_remLo_376_));
DFFPOSX1 DFFPOSX1_832 ( .CLK(clk), .D(u2__0remLo_451_0__377_), .Q(u2_remLo_377_));
DFFPOSX1 DFFPOSX1_833 ( .CLK(clk), .D(u2__0remLo_451_0__378_), .Q(u2_remLo_378_));
DFFPOSX1 DFFPOSX1_834 ( .CLK(clk), .D(u2__0remLo_451_0__379_), .Q(u2_remLo_379_));
DFFPOSX1 DFFPOSX1_835 ( .CLK(clk), .D(u2__0remLo_451_0__380_), .Q(u2_remLo_380_));
DFFPOSX1 DFFPOSX1_836 ( .CLK(clk), .D(u2__0remLo_451_0__381_), .Q(u2_remLo_381_));
DFFPOSX1 DFFPOSX1_837 ( .CLK(clk), .D(u2__0remLo_451_0__382_), .Q(u2_remLo_382_));
DFFPOSX1 DFFPOSX1_838 ( .CLK(clk), .D(u2__0remLo_451_0__383_), .Q(u2_remLo_383_));
DFFPOSX1 DFFPOSX1_839 ( .CLK(clk), .D(u2__0remLo_451_0__384_), .Q(u2_remLo_384_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk), .D(u2__0root_452_0__80_), .Q(sqrto_79_));
DFFPOSX1 DFFPOSX1_840 ( .CLK(clk), .D(u2__0remLo_451_0__385_), .Q(u2_remLo_385_));
DFFPOSX1 DFFPOSX1_841 ( .CLK(clk), .D(u2__0remLo_451_0__386_), .Q(u2_remLo_386_));
DFFPOSX1 DFFPOSX1_842 ( .CLK(clk), .D(u2__0remLo_451_0__387_), .Q(u2_remLo_387_));
DFFPOSX1 DFFPOSX1_843 ( .CLK(clk), .D(u2__0remLo_451_0__388_), .Q(u2_remLo_388_));
DFFPOSX1 DFFPOSX1_844 ( .CLK(clk), .D(u2__0remLo_451_0__389_), .Q(u2_remLo_389_));
DFFPOSX1 DFFPOSX1_845 ( .CLK(clk), .D(u2__0remLo_451_0__390_), .Q(u2_remLo_390_));
DFFPOSX1 DFFPOSX1_846 ( .CLK(clk), .D(u2__0remLo_451_0__391_), .Q(u2_remLo_391_));
DFFPOSX1 DFFPOSX1_847 ( .CLK(clk), .D(u2__0remLo_451_0__392_), .Q(u2_remLo_392_));
DFFPOSX1 DFFPOSX1_848 ( .CLK(clk), .D(u2__0remLo_451_0__393_), .Q(u2_remLo_393_));
DFFPOSX1 DFFPOSX1_849 ( .CLK(clk), .D(u2__0remLo_451_0__394_), .Q(u2_remLo_394_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk), .D(u2__0root_452_0__81_), .Q(sqrto_80_));
DFFPOSX1 DFFPOSX1_850 ( .CLK(clk), .D(u2__0remLo_451_0__395_), .Q(u2_remLo_395_));
DFFPOSX1 DFFPOSX1_851 ( .CLK(clk), .D(u2__0remLo_451_0__396_), .Q(u2_remLo_396_));
DFFPOSX1 DFFPOSX1_852 ( .CLK(clk), .D(u2__0remLo_451_0__397_), .Q(u2_remLo_397_));
DFFPOSX1 DFFPOSX1_853 ( .CLK(clk), .D(u2__0remLo_451_0__398_), .Q(u2_remLo_398_));
DFFPOSX1 DFFPOSX1_854 ( .CLK(clk), .D(u2__0remLo_451_0__399_), .Q(u2_remLo_399_));
DFFPOSX1 DFFPOSX1_855 ( .CLK(clk), .D(u2__0remLo_451_0__400_), .Q(u2_remLo_400_));
DFFPOSX1 DFFPOSX1_856 ( .CLK(clk), .D(u2__0remLo_451_0__401_), .Q(u2_remLo_401_));
DFFPOSX1 DFFPOSX1_857 ( .CLK(clk), .D(u2__0remLo_451_0__402_), .Q(u2_remLo_402_));
DFFPOSX1 DFFPOSX1_858 ( .CLK(clk), .D(u2__0remLo_451_0__403_), .Q(u2_remLo_403_));
DFFPOSX1 DFFPOSX1_859 ( .CLK(clk), .D(u2__0remLo_451_0__404_), .Q(u2_remLo_404_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk), .D(u2__0root_452_0__82_), .Q(sqrto_81_));
DFFPOSX1 DFFPOSX1_860 ( .CLK(clk), .D(u2__0remLo_451_0__405_), .Q(u2_remLo_405_));
DFFPOSX1 DFFPOSX1_861 ( .CLK(clk), .D(u2__0remLo_451_0__406_), .Q(u2_remLo_406_));
DFFPOSX1 DFFPOSX1_862 ( .CLK(clk), .D(u2__0remLo_451_0__407_), .Q(u2_remLo_407_));
DFFPOSX1 DFFPOSX1_863 ( .CLK(clk), .D(u2__0remLo_451_0__408_), .Q(u2_remLo_408_));
DFFPOSX1 DFFPOSX1_864 ( .CLK(clk), .D(u2__0remLo_451_0__409_), .Q(u2_remLo_409_));
DFFPOSX1 DFFPOSX1_865 ( .CLK(clk), .D(u2__0remLo_451_0__410_), .Q(u2_remLo_410_));
DFFPOSX1 DFFPOSX1_866 ( .CLK(clk), .D(u2__0remLo_451_0__411_), .Q(u2_remLo_411_));
DFFPOSX1 DFFPOSX1_867 ( .CLK(clk), .D(u2__0remLo_451_0__412_), .Q(u2_remLo_412_));
DFFPOSX1 DFFPOSX1_868 ( .CLK(clk), .D(u2__0remLo_451_0__413_), .Q(u2_remLo_413_));
DFFPOSX1 DFFPOSX1_869 ( .CLK(clk), .D(u2__0remLo_451_0__414_), .Q(u2_remLo_414_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk), .D(u2__0root_452_0__83_), .Q(sqrto_82_));
DFFPOSX1 DFFPOSX1_870 ( .CLK(clk), .D(u2__0remLo_451_0__415_), .Q(u2_remLo_415_));
DFFPOSX1 DFFPOSX1_871 ( .CLK(clk), .D(u2__0remLo_451_0__416_), .Q(u2_remLo_416_));
DFFPOSX1 DFFPOSX1_872 ( .CLK(clk), .D(u2__0remLo_451_0__417_), .Q(u2_remLo_417_));
DFFPOSX1 DFFPOSX1_873 ( .CLK(clk), .D(u2__0remLo_451_0__418_), .Q(u2_remLo_418_));
DFFPOSX1 DFFPOSX1_874 ( .CLK(clk), .D(u2__0remLo_451_0__419_), .Q(u2_remLo_419_));
DFFPOSX1 DFFPOSX1_875 ( .CLK(clk), .D(u2__0remLo_451_0__420_), .Q(u2_remLo_420_));
DFFPOSX1 DFFPOSX1_876 ( .CLK(clk), .D(u2__0remLo_451_0__421_), .Q(u2_remLo_421_));
DFFPOSX1 DFFPOSX1_877 ( .CLK(clk), .D(u2__0remLo_451_0__422_), .Q(u2_remLo_422_));
DFFPOSX1 DFFPOSX1_878 ( .CLK(clk), .D(u2__0remLo_451_0__423_), .Q(u2_remLo_423_));
DFFPOSX1 DFFPOSX1_879 ( .CLK(clk), .D(u2__0remLo_451_0__424_), .Q(u2_remLo_424_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk), .D(u2__0root_452_0__84_), .Q(sqrto_83_));
DFFPOSX1 DFFPOSX1_880 ( .CLK(clk), .D(u2__0remLo_451_0__425_), .Q(u2_remLo_425_));
DFFPOSX1 DFFPOSX1_881 ( .CLK(clk), .D(u2__0remLo_451_0__426_), .Q(u2_remLo_426_));
DFFPOSX1 DFFPOSX1_882 ( .CLK(clk), .D(u2__0remLo_451_0__427_), .Q(u2_remLo_427_));
DFFPOSX1 DFFPOSX1_883 ( .CLK(clk), .D(u2__0remLo_451_0__428_), .Q(u2_remLo_428_));
DFFPOSX1 DFFPOSX1_884 ( .CLK(clk), .D(u2__0remLo_451_0__429_), .Q(u2_remLo_429_));
DFFPOSX1 DFFPOSX1_885 ( .CLK(clk), .D(u2__0remLo_451_0__430_), .Q(u2_remLo_430_));
DFFPOSX1 DFFPOSX1_886 ( .CLK(clk), .D(u2__0remLo_451_0__431_), .Q(u2_remLo_431_));
DFFPOSX1 DFFPOSX1_887 ( .CLK(clk), .D(u2__0remLo_451_0__432_), .Q(u2_remLo_432_));
DFFPOSX1 DFFPOSX1_888 ( .CLK(clk), .D(u2__0remLo_451_0__433_), .Q(u2_remLo_433_));
DFFPOSX1 DFFPOSX1_889 ( .CLK(clk), .D(u2__0remLo_451_0__434_), .Q(u2_remLo_434_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk), .D(u2__0root_452_0__85_), .Q(sqrto_84_));
DFFPOSX1 DFFPOSX1_890 ( .CLK(clk), .D(u2__0remLo_451_0__435_), .Q(u2_remLo_435_));
DFFPOSX1 DFFPOSX1_891 ( .CLK(clk), .D(u2__0remLo_451_0__436_), .Q(u2_remLo_436_));
DFFPOSX1 DFFPOSX1_892 ( .CLK(clk), .D(u2__0remLo_451_0__437_), .Q(u2_remLo_437_));
DFFPOSX1 DFFPOSX1_893 ( .CLK(clk), .D(u2__0remLo_451_0__438_), .Q(u2_remLo_438_));
DFFPOSX1 DFFPOSX1_894 ( .CLK(clk), .D(u2__0remLo_451_0__439_), .Q(u2_remLo_439_));
DFFPOSX1 DFFPOSX1_895 ( .CLK(clk), .D(u2__0remLo_451_0__440_), .Q(u2_remLo_440_));
DFFPOSX1 DFFPOSX1_896 ( .CLK(clk), .D(u2__0remLo_451_0__441_), .Q(u2_remLo_441_));
DFFPOSX1 DFFPOSX1_897 ( .CLK(clk), .D(u2__0remLo_451_0__442_), .Q(u2_remLo_442_));
DFFPOSX1 DFFPOSX1_898 ( .CLK(clk), .D(u2__0remLo_451_0__443_), .Q(u2_remLo_443_));
DFFPOSX1 DFFPOSX1_899 ( .CLK(clk), .D(u2__0remLo_451_0__444_), .Q(u2_remLo_444_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(u2__0root_452_0__5_), .Q(sqrto_4_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk), .D(u2__0root_452_0__86_), .Q(sqrto_85_));
DFFPOSX1 DFFPOSX1_900 ( .CLK(clk), .D(u2__0remLo_451_0__445_), .Q(u2_remLo_445_));
DFFPOSX1 DFFPOSX1_901 ( .CLK(clk), .D(u2__0remLo_451_0__446_), .Q(u2_remLo_446_));
DFFPOSX1 DFFPOSX1_902 ( .CLK(clk), .D(u2__0remLo_451_0__447_), .Q(u2_remLo_447_));
DFFPOSX1 DFFPOSX1_903 ( .CLK(clk), .D(u2__0remLo_451_0__448_), .Q(u2_remLo_448_));
DFFPOSX1 DFFPOSX1_904 ( .CLK(clk), .D(u2__0remLo_451_0__449_), .Q(u2_remLo_449_));
DFFPOSX1 DFFPOSX1_905 ( .CLK(clk), .D(u2__0remLo_451_0__450_), .Q(u2_remHiShift_0_));
DFFPOSX1 DFFPOSX1_906 ( .CLK(clk), .D(u2__0remLo_451_0__451_), .Q(u2_remHiShift_1_));
DFFPOSX1 DFFPOSX1_907 ( .CLK(clk), .D(u2__0remHi_451_0__0_), .Q(u2_remHi_0_));
DFFPOSX1 DFFPOSX1_908 ( .CLK(clk), .D(u2__0remHi_451_0__1_), .Q(u2_remHi_1_));
DFFPOSX1 DFFPOSX1_909 ( .CLK(clk), .D(u2__0remHi_451_0__2_), .Q(u2_remHi_2_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk), .D(u2__0root_452_0__87_), .Q(sqrto_86_));
DFFPOSX1 DFFPOSX1_910 ( .CLK(clk), .D(u2__0remHi_451_0__3_), .Q(u2_remHi_3_));
DFFPOSX1 DFFPOSX1_911 ( .CLK(clk), .D(u2__0remHi_451_0__4_), .Q(u2_remHi_4_));
DFFPOSX1 DFFPOSX1_912 ( .CLK(clk), .D(u2__0remHi_451_0__5_), .Q(u2_remHi_5_));
DFFPOSX1 DFFPOSX1_913 ( .CLK(clk), .D(u2__0remHi_451_0__6_), .Q(u2_remHi_6_));
DFFPOSX1 DFFPOSX1_914 ( .CLK(clk), .D(u2__0remHi_451_0__7_), .Q(u2_remHi_7_));
DFFPOSX1 DFFPOSX1_915 ( .CLK(clk), .D(u2__0remHi_451_0__8_), .Q(u2_remHi_8_));
DFFPOSX1 DFFPOSX1_916 ( .CLK(clk), .D(u2__0remHi_451_0__9_), .Q(u2_remHi_9_));
DFFPOSX1 DFFPOSX1_917 ( .CLK(clk), .D(u2__0remHi_451_0__10_), .Q(u2_remHi_10_));
DFFPOSX1 DFFPOSX1_918 ( .CLK(clk), .D(u2__0remHi_451_0__11_), .Q(u2_remHi_11_));
DFFPOSX1 DFFPOSX1_919 ( .CLK(clk), .D(u2__0remHi_451_0__12_), .Q(u2_remHi_12_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk), .D(u2__0root_452_0__88_), .Q(sqrto_87_));
DFFPOSX1 DFFPOSX1_920 ( .CLK(clk), .D(u2__0remHi_451_0__13_), .Q(u2_remHi_13_));
DFFPOSX1 DFFPOSX1_921 ( .CLK(clk), .D(u2__0remHi_451_0__14_), .Q(u2_remHi_14_));
DFFPOSX1 DFFPOSX1_922 ( .CLK(clk), .D(u2__0remHi_451_0__15_), .Q(u2_remHi_15_));
DFFPOSX1 DFFPOSX1_923 ( .CLK(clk), .D(u2__0remHi_451_0__16_), .Q(u2_remHi_16_));
DFFPOSX1 DFFPOSX1_924 ( .CLK(clk), .D(u2__0remHi_451_0__17_), .Q(u2_remHi_17_));
DFFPOSX1 DFFPOSX1_925 ( .CLK(clk), .D(u2__0remHi_451_0__18_), .Q(u2_remHi_18_));
DFFPOSX1 DFFPOSX1_926 ( .CLK(clk), .D(u2__0remHi_451_0__19_), .Q(u2_remHi_19_));
DFFPOSX1 DFFPOSX1_927 ( .CLK(clk), .D(u2__0remHi_451_0__20_), .Q(u2_remHi_20_));
DFFPOSX1 DFFPOSX1_928 ( .CLK(clk), .D(u2__0remHi_451_0__21_), .Q(u2_remHi_21_));
DFFPOSX1 DFFPOSX1_929 ( .CLK(clk), .D(u2__0remHi_451_0__22_), .Q(u2_remHi_22_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk), .D(u2__0root_452_0__89_), .Q(sqrto_88_));
DFFPOSX1 DFFPOSX1_930 ( .CLK(clk), .D(u2__0remHi_451_0__23_), .Q(u2_remHi_23_));
DFFPOSX1 DFFPOSX1_931 ( .CLK(clk), .D(u2__0remHi_451_0__24_), .Q(u2_remHi_24_));
DFFPOSX1 DFFPOSX1_932 ( .CLK(clk), .D(u2__0remHi_451_0__25_), .Q(u2_remHi_25_));
DFFPOSX1 DFFPOSX1_933 ( .CLK(clk), .D(u2__0remHi_451_0__26_), .Q(u2_remHi_26_));
DFFPOSX1 DFFPOSX1_934 ( .CLK(clk), .D(u2__0remHi_451_0__27_), .Q(u2_remHi_27_));
DFFPOSX1 DFFPOSX1_935 ( .CLK(clk), .D(u2__0remHi_451_0__28_), .Q(u2_remHi_28_));
DFFPOSX1 DFFPOSX1_936 ( .CLK(clk), .D(u2__0remHi_451_0__29_), .Q(u2_remHi_29_));
DFFPOSX1 DFFPOSX1_937 ( .CLK(clk), .D(u2__0remHi_451_0__30_), .Q(u2_remHi_30_));
DFFPOSX1 DFFPOSX1_938 ( .CLK(clk), .D(u2__0remHi_451_0__31_), .Q(u2_remHi_31_));
DFFPOSX1 DFFPOSX1_939 ( .CLK(clk), .D(u2__0remHi_451_0__32_), .Q(u2_remHi_32_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk), .D(u2__0root_452_0__90_), .Q(sqrto_89_));
DFFPOSX1 DFFPOSX1_940 ( .CLK(clk), .D(u2__0remHi_451_0__33_), .Q(u2_remHi_33_));
DFFPOSX1 DFFPOSX1_941 ( .CLK(clk), .D(u2__0remHi_451_0__34_), .Q(u2_remHi_34_));
DFFPOSX1 DFFPOSX1_942 ( .CLK(clk), .D(u2__0remHi_451_0__35_), .Q(u2_remHi_35_));
DFFPOSX1 DFFPOSX1_943 ( .CLK(clk), .D(u2__0remHi_451_0__36_), .Q(u2_remHi_36_));
DFFPOSX1 DFFPOSX1_944 ( .CLK(clk), .D(u2__0remHi_451_0__37_), .Q(u2_remHi_37_));
DFFPOSX1 DFFPOSX1_945 ( .CLK(clk), .D(u2__0remHi_451_0__38_), .Q(u2_remHi_38_));
DFFPOSX1 DFFPOSX1_946 ( .CLK(clk), .D(u2__0remHi_451_0__39_), .Q(u2_remHi_39_));
DFFPOSX1 DFFPOSX1_947 ( .CLK(clk), .D(u2__0remHi_451_0__40_), .Q(u2_remHi_40_));
DFFPOSX1 DFFPOSX1_948 ( .CLK(clk), .D(u2__0remHi_451_0__41_), .Q(u2_remHi_41_));
DFFPOSX1 DFFPOSX1_949 ( .CLK(clk), .D(u2__0remHi_451_0__42_), .Q(u2_remHi_42_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk), .D(u2__0root_452_0__91_), .Q(sqrto_90_));
DFFPOSX1 DFFPOSX1_950 ( .CLK(clk), .D(u2__0remHi_451_0__43_), .Q(u2_remHi_43_));
DFFPOSX1 DFFPOSX1_951 ( .CLK(clk), .D(u2__0remHi_451_0__44_), .Q(u2_remHi_44_));
DFFPOSX1 DFFPOSX1_952 ( .CLK(clk), .D(u2__0remHi_451_0__45_), .Q(u2_remHi_45_));
DFFPOSX1 DFFPOSX1_953 ( .CLK(clk), .D(u2__0remHi_451_0__46_), .Q(u2_remHi_46_));
DFFPOSX1 DFFPOSX1_954 ( .CLK(clk), .D(u2__0remHi_451_0__47_), .Q(u2_remHi_47_));
DFFPOSX1 DFFPOSX1_955 ( .CLK(clk), .D(u2__0remHi_451_0__48_), .Q(u2_remHi_48_));
DFFPOSX1 DFFPOSX1_956 ( .CLK(clk), .D(u2__0remHi_451_0__49_), .Q(u2_remHi_49_));
DFFPOSX1 DFFPOSX1_957 ( .CLK(clk), .D(u2__0remHi_451_0__50_), .Q(u2_remHi_50_));
DFFPOSX1 DFFPOSX1_958 ( .CLK(clk), .D(u2__0remHi_451_0__51_), .Q(u2_remHi_51_));
DFFPOSX1 DFFPOSX1_959 ( .CLK(clk), .D(u2__0remHi_451_0__52_), .Q(u2_remHi_52_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk), .D(u2__0root_452_0__92_), .Q(sqrto_91_));
DFFPOSX1 DFFPOSX1_960 ( .CLK(clk), .D(u2__0remHi_451_0__53_), .Q(u2_remHi_53_));
DFFPOSX1 DFFPOSX1_961 ( .CLK(clk), .D(u2__0remHi_451_0__54_), .Q(u2_remHi_54_));
DFFPOSX1 DFFPOSX1_962 ( .CLK(clk), .D(u2__0remHi_451_0__55_), .Q(u2_remHi_55_));
DFFPOSX1 DFFPOSX1_963 ( .CLK(clk), .D(u2__0remHi_451_0__56_), .Q(u2_remHi_56_));
DFFPOSX1 DFFPOSX1_964 ( .CLK(clk), .D(u2__0remHi_451_0__57_), .Q(u2_remHi_57_));
DFFPOSX1 DFFPOSX1_965 ( .CLK(clk), .D(u2__0remHi_451_0__58_), .Q(u2_remHi_58_));
DFFPOSX1 DFFPOSX1_966 ( .CLK(clk), .D(u2__0remHi_451_0__59_), .Q(u2_remHi_59_));
DFFPOSX1 DFFPOSX1_967 ( .CLK(clk), .D(u2__0remHi_451_0__60_), .Q(u2_remHi_60_));
DFFPOSX1 DFFPOSX1_968 ( .CLK(clk), .D(u2__0remHi_451_0__61_), .Q(u2_remHi_61_));
DFFPOSX1 DFFPOSX1_969 ( .CLK(clk), .D(u2__0remHi_451_0__62_), .Q(u2_remHi_62_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk), .D(u2__0root_452_0__93_), .Q(sqrto_92_));
DFFPOSX1 DFFPOSX1_970 ( .CLK(clk), .D(u2__0remHi_451_0__63_), .Q(u2_remHi_63_));
DFFPOSX1 DFFPOSX1_971 ( .CLK(clk), .D(u2__0remHi_451_0__64_), .Q(u2_remHi_64_));
DFFPOSX1 DFFPOSX1_972 ( .CLK(clk), .D(u2__0remHi_451_0__65_), .Q(u2_remHi_65_));
DFFPOSX1 DFFPOSX1_973 ( .CLK(clk), .D(u2__0remHi_451_0__66_), .Q(u2_remHi_66_));
DFFPOSX1 DFFPOSX1_974 ( .CLK(clk), .D(u2__0remHi_451_0__67_), .Q(u2_remHi_67_));
DFFPOSX1 DFFPOSX1_975 ( .CLK(clk), .D(u2__0remHi_451_0__68_), .Q(u2_remHi_68_));
DFFPOSX1 DFFPOSX1_976 ( .CLK(clk), .D(u2__0remHi_451_0__69_), .Q(u2_remHi_69_));
DFFPOSX1 DFFPOSX1_977 ( .CLK(clk), .D(u2__0remHi_451_0__70_), .Q(u2_remHi_70_));
DFFPOSX1 DFFPOSX1_978 ( .CLK(clk), .D(u2__0remHi_451_0__71_), .Q(u2_remHi_71_));
DFFPOSX1 DFFPOSX1_979 ( .CLK(clk), .D(u2__0remHi_451_0__72_), .Q(u2_remHi_72_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk), .D(u2__0root_452_0__94_), .Q(sqrto_93_));
DFFPOSX1 DFFPOSX1_980 ( .CLK(clk), .D(u2__0remHi_451_0__73_), .Q(u2_remHi_73_));
DFFPOSX1 DFFPOSX1_981 ( .CLK(clk), .D(u2__0remHi_451_0__74_), .Q(u2_remHi_74_));
DFFPOSX1 DFFPOSX1_982 ( .CLK(clk), .D(u2__0remHi_451_0__75_), .Q(u2_remHi_75_));
DFFPOSX1 DFFPOSX1_983 ( .CLK(clk), .D(u2__0remHi_451_0__76_), .Q(u2_remHi_76_));
DFFPOSX1 DFFPOSX1_984 ( .CLK(clk), .D(u2__0remHi_451_0__77_), .Q(u2_remHi_77_));
DFFPOSX1 DFFPOSX1_985 ( .CLK(clk), .D(u2__0remHi_451_0__78_), .Q(u2_remHi_78_));
DFFPOSX1 DFFPOSX1_986 ( .CLK(clk), .D(u2__0remHi_451_0__79_), .Q(u2_remHi_79_));
DFFPOSX1 DFFPOSX1_987 ( .CLK(clk), .D(u2__0remHi_451_0__80_), .Q(u2_remHi_80_));
DFFPOSX1 DFFPOSX1_988 ( .CLK(clk), .D(u2__0remHi_451_0__81_), .Q(u2_remHi_81_));
DFFPOSX1 DFFPOSX1_989 ( .CLK(clk), .D(u2__0remHi_451_0__82_), .Q(u2_remHi_82_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk), .D(u2__0root_452_0__95_), .Q(sqrto_94_));
DFFPOSX1 DFFPOSX1_990 ( .CLK(clk), .D(u2__0remHi_451_0__83_), .Q(u2_remHi_83_));
DFFPOSX1 DFFPOSX1_991 ( .CLK(clk), .D(u2__0remHi_451_0__84_), .Q(u2_remHi_84_));
DFFPOSX1 DFFPOSX1_992 ( .CLK(clk), .D(u2__0remHi_451_0__85_), .Q(u2_remHi_85_));
DFFPOSX1 DFFPOSX1_993 ( .CLK(clk), .D(u2__0remHi_451_0__86_), .Q(u2_remHi_86_));
DFFPOSX1 DFFPOSX1_994 ( .CLK(clk), .D(u2__0remHi_451_0__87_), .Q(u2_remHi_87_));
DFFPOSX1 DFFPOSX1_995 ( .CLK(clk), .D(u2__0remHi_451_0__88_), .Q(u2_remHi_88_));
DFFPOSX1 DFFPOSX1_996 ( .CLK(clk), .D(u2__0remHi_451_0__89_), .Q(u2_remHi_89_));
DFFPOSX1 DFFPOSX1_997 ( .CLK(clk), .D(u2__0remHi_451_0__90_), .Q(u2_remHi_90_));
DFFPOSX1 DFFPOSX1_998 ( .CLK(clk), .D(u2__0remHi_451_0__91_), .Q(u2_remHi_91_));
DFFPOSX1 DFFPOSX1_999 ( .CLK(clk), .D(u2__0remHi_451_0__92_), .Q(u2_remHi_92_));
INVX1 INVX1_1 ( .A(aNan), .Y(_abc_73687_new_n753_));
INVX1 INVX1_10 ( .A(_abc_73687_new_n1532_), .Y(_abc_73687_new_n1538_));
INVX1 INVX1_100 ( .A(\a[90] ), .Y(u1__abc_51895_new_n261_));
INVX1 INVX1_1000 ( .A(u2__abc_52155_new_n4899_), .Y(u2__abc_52155_new_n4900_));
INVX1 INVX1_1001 ( .A(u2_remHi_177_), .Y(u2__abc_52155_new_n4901_));
INVX1 INVX1_1002 ( .A(u2__abc_52155_new_n4902_), .Y(u2__abc_52155_new_n4903_));
INVX1 INVX1_1003 ( .A(sqrto_174_), .Y(u2__abc_52155_new_n4906_));
INVX1 INVX1_1004 ( .A(u2__abc_52155_new_n4907_), .Y(u2__abc_52155_new_n4908_));
INVX1 INVX1_1005 ( .A(u2_remHi_174_), .Y(u2__abc_52155_new_n4909_));
INVX1 INVX1_1006 ( .A(u2__abc_52155_new_n4910_), .Y(u2__abc_52155_new_n4911_));
INVX1 INVX1_1007 ( .A(sqrto_175_), .Y(u2__abc_52155_new_n4913_));
INVX1 INVX1_1008 ( .A(u2__abc_52155_new_n4914_), .Y(u2__abc_52155_new_n4915_));
INVX1 INVX1_1009 ( .A(u2_remHi_175_), .Y(u2__abc_52155_new_n4916_));
INVX1 INVX1_101 ( .A(\a[91] ), .Y(u1__abc_51895_new_n262_));
INVX1 INVX1_1010 ( .A(u2__abc_52155_new_n4917_), .Y(u2__abc_52155_new_n4918_));
INVX1 INVX1_1011 ( .A(sqrto_172_), .Y(u2__abc_52155_new_n4924_));
INVX1 INVX1_1012 ( .A(u2__abc_52155_new_n4925_), .Y(u2__abc_52155_new_n4926_));
INVX1 INVX1_1013 ( .A(u2_remHi_172_), .Y(u2__abc_52155_new_n4927_));
INVX1 INVX1_1014 ( .A(u2__abc_52155_new_n4928_), .Y(u2__abc_52155_new_n4929_));
INVX1 INVX1_1015 ( .A(sqrto_173_), .Y(u2__abc_52155_new_n4931_));
INVX1 INVX1_1016 ( .A(u2__abc_52155_new_n4932_), .Y(u2__abc_52155_new_n4933_));
INVX1 INVX1_1017 ( .A(u2_remHi_173_), .Y(u2__abc_52155_new_n4934_));
INVX1 INVX1_1018 ( .A(u2__abc_52155_new_n4935_), .Y(u2__abc_52155_new_n4936_));
INVX1 INVX1_1019 ( .A(sqrto_171_), .Y(u2__abc_52155_new_n4939_));
INVX1 INVX1_102 ( .A(\a[88] ), .Y(u1__abc_51895_new_n264_));
INVX1 INVX1_1020 ( .A(u2__abc_52155_new_n4940_), .Y(u2__abc_52155_new_n4941_));
INVX1 INVX1_1021 ( .A(u2_remHi_171_), .Y(u2__abc_52155_new_n4942_));
INVX1 INVX1_1022 ( .A(u2__abc_52155_new_n4943_), .Y(u2__abc_52155_new_n4944_));
INVX1 INVX1_1023 ( .A(sqrto_170_), .Y(u2__abc_52155_new_n4946_));
INVX1 INVX1_1024 ( .A(u2__abc_52155_new_n4947_), .Y(u2__abc_52155_new_n4948_));
INVX1 INVX1_1025 ( .A(u2_remHi_170_), .Y(u2__abc_52155_new_n4949_));
INVX1 INVX1_1026 ( .A(u2__abc_52155_new_n4950_), .Y(u2__abc_52155_new_n4951_));
INVX1 INVX1_1027 ( .A(sqrto_168_), .Y(u2__abc_52155_new_n4955_));
INVX1 INVX1_1028 ( .A(u2__abc_52155_new_n4956_), .Y(u2__abc_52155_new_n4957_));
INVX1 INVX1_1029 ( .A(u2_remHi_168_), .Y(u2__abc_52155_new_n4958_));
INVX1 INVX1_103 ( .A(\a[89] ), .Y(u1__abc_51895_new_n265_));
INVX1 INVX1_1030 ( .A(u2__abc_52155_new_n4959_), .Y(u2__abc_52155_new_n4960_));
INVX1 INVX1_1031 ( .A(sqrto_169_), .Y(u2__abc_52155_new_n4962_));
INVX1 INVX1_1032 ( .A(u2__abc_52155_new_n4963_), .Y(u2__abc_52155_new_n4964_));
INVX1 INVX1_1033 ( .A(u2_remHi_169_), .Y(u2__abc_52155_new_n4965_));
INVX1 INVX1_1034 ( .A(u2__abc_52155_new_n4966_), .Y(u2__abc_52155_new_n4967_));
INVX1 INVX1_1035 ( .A(sqrto_167_), .Y(u2__abc_52155_new_n4970_));
INVX1 INVX1_1036 ( .A(u2__abc_52155_new_n4971_), .Y(u2__abc_52155_new_n4972_));
INVX1 INVX1_1037 ( .A(u2_remHi_167_), .Y(u2__abc_52155_new_n4973_));
INVX1 INVX1_1038 ( .A(u2__abc_52155_new_n4974_), .Y(u2__abc_52155_new_n4975_));
INVX1 INVX1_1039 ( .A(sqrto_166_), .Y(u2__abc_52155_new_n4977_));
INVX1 INVX1_104 ( .A(\a[94] ), .Y(u1__abc_51895_new_n268_));
INVX1 INVX1_1040 ( .A(u2__abc_52155_new_n4978_), .Y(u2__abc_52155_new_n4979_));
INVX1 INVX1_1041 ( .A(u2_remHi_166_), .Y(u2__abc_52155_new_n4980_));
INVX1 INVX1_1042 ( .A(u2__abc_52155_new_n4981_), .Y(u2__abc_52155_new_n4982_));
INVX1 INVX1_1043 ( .A(sqrto_160_), .Y(u2__abc_52155_new_n4987_));
INVX1 INVX1_1044 ( .A(u2_remHi_160_), .Y(u2__abc_52155_new_n4989_));
INVX1 INVX1_1045 ( .A(sqrto_161_), .Y(u2__abc_52155_new_n4992_));
INVX1 INVX1_1046 ( .A(u2_remHi_161_), .Y(u2__abc_52155_new_n4994_));
INVX1 INVX1_1047 ( .A(u2__abc_52155_new_n4997_), .Y(u2__abc_52155_new_n4998_));
INVX1 INVX1_1048 ( .A(sqrto_159_), .Y(u2__abc_52155_new_n4999_));
INVX1 INVX1_1049 ( .A(u2__abc_52155_new_n5000_), .Y(u2__abc_52155_new_n5001_));
INVX1 INVX1_105 ( .A(\a[95] ), .Y(u1__abc_51895_new_n269_));
INVX1 INVX1_1050 ( .A(u2_remHi_159_), .Y(u2__abc_52155_new_n5002_));
INVX1 INVX1_1051 ( .A(u2__abc_52155_new_n5003_), .Y(u2__abc_52155_new_n5004_));
INVX1 INVX1_1052 ( .A(sqrto_158_), .Y(u2__abc_52155_new_n5006_));
INVX1 INVX1_1053 ( .A(u2__abc_52155_new_n5007_), .Y(u2__abc_52155_new_n5008_));
INVX1 INVX1_1054 ( .A(u2_remHi_158_), .Y(u2__abc_52155_new_n5009_));
INVX1 INVX1_1055 ( .A(u2__abc_52155_new_n5010_), .Y(u2__abc_52155_new_n5011_));
INVX1 INVX1_1056 ( .A(sqrto_164_), .Y(u2__abc_52155_new_n5015_));
INVX1 INVX1_1057 ( .A(u2__abc_52155_new_n5016_), .Y(u2__abc_52155_new_n5017_));
INVX1 INVX1_1058 ( .A(u2_remHi_164_), .Y(u2__abc_52155_new_n5018_));
INVX1 INVX1_1059 ( .A(u2__abc_52155_new_n5019_), .Y(u2__abc_52155_new_n5020_));
INVX1 INVX1_106 ( .A(\a[92] ), .Y(u1__abc_51895_new_n271_));
INVX1 INVX1_1060 ( .A(sqrto_165_), .Y(u2__abc_52155_new_n5022_));
INVX1 INVX1_1061 ( .A(u2__abc_52155_new_n5023_), .Y(u2__abc_52155_new_n5024_));
INVX1 INVX1_1062 ( .A(u2_remHi_165_), .Y(u2__abc_52155_new_n5025_));
INVX1 INVX1_1063 ( .A(u2__abc_52155_new_n5026_), .Y(u2__abc_52155_new_n5027_));
INVX1 INVX1_1064 ( .A(sqrto_163_), .Y(u2__abc_52155_new_n5030_));
INVX1 INVX1_1065 ( .A(u2__abc_52155_new_n5031_), .Y(u2__abc_52155_new_n5032_));
INVX1 INVX1_1066 ( .A(u2_remHi_163_), .Y(u2__abc_52155_new_n5033_));
INVX1 INVX1_1067 ( .A(u2__abc_52155_new_n5034_), .Y(u2__abc_52155_new_n5035_));
INVX1 INVX1_1068 ( .A(sqrto_162_), .Y(u2__abc_52155_new_n5037_));
INVX1 INVX1_1069 ( .A(u2__abc_52155_new_n5038_), .Y(u2__abc_52155_new_n5039_));
INVX1 INVX1_107 ( .A(\a[93] ), .Y(u1__abc_51895_new_n272_));
INVX1 INVX1_1070 ( .A(u2_remHi_162_), .Y(u2__abc_52155_new_n5040_));
INVX1 INVX1_1071 ( .A(u2__abc_52155_new_n5041_), .Y(u2__abc_52155_new_n5042_));
INVX1 INVX1_1072 ( .A(sqrto_152_), .Y(u2__abc_52155_new_n5049_));
INVX1 INVX1_1073 ( .A(u2__abc_52155_new_n5050_), .Y(u2__abc_52155_new_n5051_));
INVX1 INVX1_1074 ( .A(u2_remHi_152_), .Y(u2__abc_52155_new_n5052_));
INVX1 INVX1_1075 ( .A(u2__abc_52155_new_n5053_), .Y(u2__abc_52155_new_n5054_));
INVX1 INVX1_1076 ( .A(sqrto_153_), .Y(u2__abc_52155_new_n5056_));
INVX1 INVX1_1077 ( .A(u2__abc_52155_new_n5057_), .Y(u2__abc_52155_new_n5058_));
INVX1 INVX1_1078 ( .A(u2_remHi_153_), .Y(u2__abc_52155_new_n5059_));
INVX1 INVX1_1079 ( .A(u2__abc_52155_new_n5060_), .Y(u2__abc_52155_new_n5061_));
INVX1 INVX1_108 ( .A(\a[82] ), .Y(u1__abc_51895_new_n276_));
INVX1 INVX1_1080 ( .A(sqrto_151_), .Y(u2__abc_52155_new_n5064_));
INVX1 INVX1_1081 ( .A(u2__abc_52155_new_n5065_), .Y(u2__abc_52155_new_n5066_));
INVX1 INVX1_1082 ( .A(u2_remHi_151_), .Y(u2__abc_52155_new_n5067_));
INVX1 INVX1_1083 ( .A(u2__abc_52155_new_n5068_), .Y(u2__abc_52155_new_n5069_));
INVX1 INVX1_1084 ( .A(sqrto_150_), .Y(u2__abc_52155_new_n5071_));
INVX1 INVX1_1085 ( .A(u2__abc_52155_new_n5072_), .Y(u2__abc_52155_new_n5073_));
INVX1 INVX1_1086 ( .A(u2_remHi_150_), .Y(u2__abc_52155_new_n5074_));
INVX1 INVX1_1087 ( .A(u2__abc_52155_new_n5075_), .Y(u2__abc_52155_new_n5076_));
INVX1 INVX1_1088 ( .A(sqrto_156_), .Y(u2__abc_52155_new_n5080_));
INVX1 INVX1_1089 ( .A(u2__abc_52155_new_n5081_), .Y(u2__abc_52155_new_n5082_));
INVX1 INVX1_109 ( .A(\a[83] ), .Y(u1__abc_51895_new_n277_));
INVX1 INVX1_1090 ( .A(u2_remHi_156_), .Y(u2__abc_52155_new_n5083_));
INVX1 INVX1_1091 ( .A(u2__abc_52155_new_n5084_), .Y(u2__abc_52155_new_n5085_));
INVX1 INVX1_1092 ( .A(sqrto_157_), .Y(u2__abc_52155_new_n5087_));
INVX1 INVX1_1093 ( .A(u2__abc_52155_new_n5088_), .Y(u2__abc_52155_new_n5089_));
INVX1 INVX1_1094 ( .A(u2_remHi_157_), .Y(u2__abc_52155_new_n5090_));
INVX1 INVX1_1095 ( .A(u2__abc_52155_new_n5091_), .Y(u2__abc_52155_new_n5092_));
INVX1 INVX1_1096 ( .A(sqrto_155_), .Y(u2__abc_52155_new_n5095_));
INVX1 INVX1_1097 ( .A(u2__abc_52155_new_n5096_), .Y(u2__abc_52155_new_n5097_));
INVX1 INVX1_1098 ( .A(u2_remHi_155_), .Y(u2__abc_52155_new_n5098_));
INVX1 INVX1_1099 ( .A(u2__abc_52155_new_n5099_), .Y(u2__abc_52155_new_n5100_));
INVX1 INVX1_11 ( .A(_abc_73687_new_n1535_), .Y(_abc_73687_new_n1542_));
INVX1 INVX1_110 ( .A(\a[80] ), .Y(u1__abc_51895_new_n279_));
INVX1 INVX1_1100 ( .A(sqrto_154_), .Y(u2__abc_52155_new_n5102_));
INVX1 INVX1_1101 ( .A(u2__abc_52155_new_n5103_), .Y(u2__abc_52155_new_n5104_));
INVX1 INVX1_1102 ( .A(u2_remHi_154_), .Y(u2__abc_52155_new_n5105_));
INVX1 INVX1_1103 ( .A(u2__abc_52155_new_n5106_), .Y(u2__abc_52155_new_n5107_));
INVX1 INVX1_1104 ( .A(sqrto_148_), .Y(u2__abc_52155_new_n5112_));
INVX1 INVX1_1105 ( .A(u2__abc_52155_new_n5113_), .Y(u2__abc_52155_new_n5114_));
INVX1 INVX1_1106 ( .A(u2_remHi_148_), .Y(u2__abc_52155_new_n5115_));
INVX1 INVX1_1107 ( .A(u2__abc_52155_new_n5116_), .Y(u2__abc_52155_new_n5117_));
INVX1 INVX1_1108 ( .A(sqrto_149_), .Y(u2__abc_52155_new_n5119_));
INVX1 INVX1_1109 ( .A(u2__abc_52155_new_n5120_), .Y(u2__abc_52155_new_n5121_));
INVX1 INVX1_111 ( .A(\a[81] ), .Y(u1__abc_51895_new_n280_));
INVX1 INVX1_1110 ( .A(u2_remHi_149_), .Y(u2__abc_52155_new_n5122_));
INVX1 INVX1_1111 ( .A(u2__abc_52155_new_n5123_), .Y(u2__abc_52155_new_n5124_));
INVX1 INVX1_1112 ( .A(sqrto_147_), .Y(u2__abc_52155_new_n5127_));
INVX1 INVX1_1113 ( .A(u2__abc_52155_new_n5128_), .Y(u2__abc_52155_new_n5129_));
INVX1 INVX1_1114 ( .A(u2_remHi_147_), .Y(u2__abc_52155_new_n5130_));
INVX1 INVX1_1115 ( .A(u2__abc_52155_new_n5131_), .Y(u2__abc_52155_new_n5132_));
INVX1 INVX1_1116 ( .A(sqrto_146_), .Y(u2__abc_52155_new_n5134_));
INVX1 INVX1_1117 ( .A(u2__abc_52155_new_n5135_), .Y(u2__abc_52155_new_n5136_));
INVX1 INVX1_1118 ( .A(u2_remHi_146_), .Y(u2__abc_52155_new_n5137_));
INVX1 INVX1_1119 ( .A(u2__abc_52155_new_n5138_), .Y(u2__abc_52155_new_n5139_));
INVX1 INVX1_112 ( .A(\a[86] ), .Y(u1__abc_51895_new_n283_));
INVX1 INVX1_1120 ( .A(sqrto_144_), .Y(u2__abc_52155_new_n5143_));
INVX1 INVX1_1121 ( .A(u2_remHi_144_), .Y(u2__abc_52155_new_n5145_));
INVX1 INVX1_1122 ( .A(sqrto_145_), .Y(u2__abc_52155_new_n5148_));
INVX1 INVX1_1123 ( .A(u2_remHi_145_), .Y(u2__abc_52155_new_n5150_));
INVX1 INVX1_1124 ( .A(u2__abc_52155_new_n5153_), .Y(u2__abc_52155_new_n5154_));
INVX1 INVX1_1125 ( .A(sqrto_143_), .Y(u2__abc_52155_new_n5155_));
INVX1 INVX1_1126 ( .A(u2__abc_52155_new_n5156_), .Y(u2__abc_52155_new_n5157_));
INVX1 INVX1_1127 ( .A(u2_remHi_143_), .Y(u2__abc_52155_new_n5158_));
INVX1 INVX1_1128 ( .A(u2__abc_52155_new_n5159_), .Y(u2__abc_52155_new_n5160_));
INVX1 INVX1_1129 ( .A(sqrto_142_), .Y(u2__abc_52155_new_n5162_));
INVX1 INVX1_113 ( .A(\a[87] ), .Y(u1__abc_51895_new_n284_));
INVX1 INVX1_1130 ( .A(u2__abc_52155_new_n5163_), .Y(u2__abc_52155_new_n5164_));
INVX1 INVX1_1131 ( .A(u2_remHi_142_), .Y(u2__abc_52155_new_n5165_));
INVX1 INVX1_1132 ( .A(u2__abc_52155_new_n5166_), .Y(u2__abc_52155_new_n5167_));
INVX1 INVX1_1133 ( .A(sqrto_136_), .Y(u2__abc_52155_new_n5173_));
INVX1 INVX1_1134 ( .A(u2_remHi_136_), .Y(u2__abc_52155_new_n5175_));
INVX1 INVX1_1135 ( .A(sqrto_137_), .Y(u2__abc_52155_new_n5178_));
INVX1 INVX1_1136 ( .A(u2_remHi_137_), .Y(u2__abc_52155_new_n5180_));
INVX1 INVX1_1137 ( .A(u2__abc_52155_new_n5183_), .Y(u2__abc_52155_new_n5184_));
INVX1 INVX1_1138 ( .A(sqrto_134_), .Y(u2__abc_52155_new_n5185_));
INVX1 INVX1_1139 ( .A(u2__abc_52155_new_n5186_), .Y(u2__abc_52155_new_n5187_));
INVX1 INVX1_114 ( .A(\a[84] ), .Y(u1__abc_51895_new_n286_));
INVX1 INVX1_1140 ( .A(u2_remHi_134_), .Y(u2__abc_52155_new_n5188_));
INVX1 INVX1_1141 ( .A(u2__abc_52155_new_n5189_), .Y(u2__abc_52155_new_n5190_));
INVX1 INVX1_1142 ( .A(sqrto_135_), .Y(u2__abc_52155_new_n5192_));
INVX1 INVX1_1143 ( .A(u2__abc_52155_new_n5193_), .Y(u2__abc_52155_new_n5194_));
INVX1 INVX1_1144 ( .A(u2_remHi_135_), .Y(u2__abc_52155_new_n5195_));
INVX1 INVX1_1145 ( .A(u2__abc_52155_new_n5196_), .Y(u2__abc_52155_new_n5197_));
INVX1 INVX1_1146 ( .A(sqrto_140_), .Y(u2__abc_52155_new_n5201_));
INVX1 INVX1_1147 ( .A(u2__abc_52155_new_n5202_), .Y(u2__abc_52155_new_n5203_));
INVX1 INVX1_1148 ( .A(u2_remHi_140_), .Y(u2__abc_52155_new_n5204_));
INVX1 INVX1_1149 ( .A(u2__abc_52155_new_n5205_), .Y(u2__abc_52155_new_n5206_));
INVX1 INVX1_115 ( .A(\a[85] ), .Y(u1__abc_51895_new_n287_));
INVX1 INVX1_1150 ( .A(sqrto_141_), .Y(u2__abc_52155_new_n5208_));
INVX1 INVX1_1151 ( .A(u2__abc_52155_new_n5209_), .Y(u2__abc_52155_new_n5210_));
INVX1 INVX1_1152 ( .A(u2_remHi_141_), .Y(u2__abc_52155_new_n5211_));
INVX1 INVX1_1153 ( .A(u2__abc_52155_new_n5212_), .Y(u2__abc_52155_new_n5213_));
INVX1 INVX1_1154 ( .A(sqrto_139_), .Y(u2__abc_52155_new_n5216_));
INVX1 INVX1_1155 ( .A(u2__abc_52155_new_n5217_), .Y(u2__abc_52155_new_n5218_));
INVX1 INVX1_1156 ( .A(u2_remHi_139_), .Y(u2__abc_52155_new_n5219_));
INVX1 INVX1_1157 ( .A(u2__abc_52155_new_n5220_), .Y(u2__abc_52155_new_n5221_));
INVX1 INVX1_1158 ( .A(sqrto_138_), .Y(u2__abc_52155_new_n5223_));
INVX1 INVX1_1159 ( .A(u2__abc_52155_new_n5224_), .Y(u2__abc_52155_new_n5225_));
INVX1 INVX1_116 ( .A(\a[106] ), .Y(u1__abc_51895_new_n292_));
INVX1 INVX1_1160 ( .A(u2_remHi_138_), .Y(u2__abc_52155_new_n5226_));
INVX1 INVX1_1161 ( .A(u2__abc_52155_new_n5227_), .Y(u2__abc_52155_new_n5228_));
INVX1 INVX1_1162 ( .A(sqrto_126_), .Y(u2__abc_52155_new_n5233_));
INVX1 INVX1_1163 ( .A(u2__abc_52155_new_n5234_), .Y(u2__abc_52155_new_n5235_));
INVX1 INVX1_1164 ( .A(sqrto_127_), .Y(u2__abc_52155_new_n5238_));
INVX1 INVX1_1165 ( .A(u2__abc_52155_new_n5239_), .Y(u2__abc_52155_new_n5240_));
INVX1 INVX1_1166 ( .A(u2_remHi_127_), .Y(u2__abc_52155_new_n5241_));
INVX1 INVX1_1167 ( .A(u2__abc_52155_new_n5242_), .Y(u2__abc_52155_new_n5243_));
INVX1 INVX1_1168 ( .A(sqrto_128_), .Y(u2__abc_52155_new_n5246_));
INVX1 INVX1_1169 ( .A(u2_remHi_128_), .Y(u2__abc_52155_new_n5248_));
INVX1 INVX1_117 ( .A(\a[107] ), .Y(u1__abc_51895_new_n293_));
INVX1 INVX1_1170 ( .A(sqrto_129_), .Y(u2__abc_52155_new_n5251_));
INVX1 INVX1_1171 ( .A(u2_remHi_129_), .Y(u2__abc_52155_new_n5253_));
INVX1 INVX1_1172 ( .A(u2__abc_52155_new_n5256_), .Y(u2__abc_52155_new_n5257_));
INVX1 INVX1_1173 ( .A(sqrto_132_), .Y(u2__abc_52155_new_n5259_));
INVX1 INVX1_1174 ( .A(u2_remHi_132_), .Y(u2__abc_52155_new_n5261_));
INVX1 INVX1_1175 ( .A(sqrto_133_), .Y(u2__abc_52155_new_n5264_));
INVX1 INVX1_1176 ( .A(u2_remHi_133_), .Y(u2__abc_52155_new_n5266_));
INVX1 INVX1_1177 ( .A(sqrto_131_), .Y(u2__abc_52155_new_n5270_));
INVX1 INVX1_1178 ( .A(u2_remHi_131_), .Y(u2__abc_52155_new_n5272_));
INVX1 INVX1_1179 ( .A(sqrto_130_), .Y(u2__abc_52155_new_n5275_));
INVX1 INVX1_118 ( .A(\a[104] ), .Y(u1__abc_51895_new_n295_));
INVX1 INVX1_1180 ( .A(u2_remHi_130_), .Y(u2__abc_52155_new_n5277_));
INVX1 INVX1_1181 ( .A(u2__abc_52155_new_n5281_), .Y(u2__abc_52155_new_n5282_));
INVX1 INVX1_1182 ( .A(u2__abc_52155_new_n5287_), .Y(u2__abc_52155_new_n5288_));
INVX1 INVX1_1183 ( .A(u2__abc_52155_new_n4796_), .Y(u2__abc_52155_new_n5290_));
INVX1 INVX1_1184 ( .A(u2__abc_52155_new_n5048_), .Y(u2__abc_52155_new_n5291_));
INVX1 INVX1_1185 ( .A(u2__abc_52155_new_n5172_), .Y(u2__abc_52155_new_n5292_));
INVX1 INVX1_1186 ( .A(u2__abc_52155_new_n5232_), .Y(u2__abc_52155_new_n5293_));
INVX1 INVX1_1187 ( .A(u2__abc_52155_new_n5254_), .Y(u2__abc_52155_new_n5297_));
INVX1 INVX1_1188 ( .A(u2__abc_52155_new_n5249_), .Y(u2__abc_52155_new_n5298_));
INVX1 INVX1_1189 ( .A(u2__abc_52155_new_n5273_), .Y(u2__abc_52155_new_n5303_));
INVX1 INVX1_119 ( .A(\a[105] ), .Y(u1__abc_51895_new_n296_));
INVX1 INVX1_1190 ( .A(u2__abc_52155_new_n5278_), .Y(u2__abc_52155_new_n5304_));
INVX1 INVX1_1191 ( .A(u2__abc_52155_new_n5265_), .Y(u2__abc_52155_new_n5308_));
INVX1 INVX1_1192 ( .A(u2__abc_52155_new_n5310_), .Y(u2__abc_52155_new_n5311_));
INVX1 INVX1_1193 ( .A(u2__abc_52155_new_n5231_), .Y(u2__abc_52155_new_n5315_));
INVX1 INVX1_1194 ( .A(u2__abc_52155_new_n5179_), .Y(u2__abc_52155_new_n5319_));
INVX1 INVX1_1195 ( .A(u2__abc_52155_new_n5321_), .Y(u2__abc_52155_new_n5322_));
INVX1 INVX1_1196 ( .A(u2__abc_52155_new_n5330_), .Y(u2__abc_52155_new_n5331_));
INVX1 INVX1_1197 ( .A(u2__abc_52155_new_n5111_), .Y(u2__abc_52155_new_n5335_));
INVX1 INVX1_1198 ( .A(u2__abc_52155_new_n5142_), .Y(u2__abc_52155_new_n5336_));
INVX1 INVX1_1199 ( .A(u2__abc_52155_new_n5149_), .Y(u2__abc_52155_new_n5340_));
INVX1 INVX1_12 ( .A(\a[117] ), .Y(_abc_73687_new_n1548_));
INVX1 INVX1_120 ( .A(\a[110] ), .Y(u1__abc_51895_new_n299_));
INVX1 INVX1_1200 ( .A(u2__abc_52155_new_n5342_), .Y(u2__abc_52155_new_n5343_));
INVX1 INVX1_1201 ( .A(u2__abc_52155_new_n5351_), .Y(u2__abc_52155_new_n5352_));
INVX1 INVX1_1202 ( .A(u2__abc_52155_new_n5368_), .Y(u2__abc_52155_new_n5369_));
INVX1 INVX1_1203 ( .A(u2__abc_52155_new_n4923_), .Y(u2__abc_52155_new_n5373_));
INVX1 INVX1_1204 ( .A(u2__abc_52155_new_n4986_), .Y(u2__abc_52155_new_n5374_));
INVX1 INVX1_1205 ( .A(u2__abc_52155_new_n5045_), .Y(u2__abc_52155_new_n5375_));
INVX1 INVX1_1206 ( .A(u2__abc_52155_new_n4993_), .Y(u2__abc_52155_new_n5379_));
INVX1 INVX1_1207 ( .A(u2__abc_52155_new_n5381_), .Y(u2__abc_52155_new_n5382_));
INVX1 INVX1_1208 ( .A(u2__abc_52155_new_n5390_), .Y(u2__abc_52155_new_n5391_));
INVX1 INVX1_1209 ( .A(u2__abc_52155_new_n5407_), .Y(u2__abc_52155_new_n5408_));
INVX1 INVX1_121 ( .A(\a[111] ), .Y(u1__abc_51895_new_n300_));
INVX1 INVX1_1210 ( .A(u2__abc_52155_new_n5440_), .Y(u2__abc_52155_new_n5441_));
INVX1 INVX1_1211 ( .A(u2__abc_52155_new_n4543_), .Y(u2__abc_52155_new_n5445_));
INVX1 INVX1_1212 ( .A(u2__abc_52155_new_n4670_), .Y(u2__abc_52155_new_n5446_));
INVX1 INVX1_1213 ( .A(u2__abc_52155_new_n4733_), .Y(u2__abc_52155_new_n5447_));
INVX1 INVX1_1214 ( .A(u2__abc_52155_new_n4764_), .Y(u2__abc_52155_new_n5448_));
INVX1 INVX1_1215 ( .A(u2__abc_52155_new_n4771_), .Y(u2__abc_52155_new_n5452_));
INVX1 INVX1_1216 ( .A(u2__abc_52155_new_n5454_), .Y(u2__abc_52155_new_n5455_));
INVX1 INVX1_1217 ( .A(u2__abc_52155_new_n5463_), .Y(u2__abc_52155_new_n5464_));
INVX1 INVX1_1218 ( .A(u2__abc_52155_new_n5480_), .Y(u2__abc_52155_new_n5481_));
INVX1 INVX1_1219 ( .A(u2__abc_52155_new_n5513_), .Y(u2__abc_52155_new_n5514_));
INVX1 INVX1_122 ( .A(\a[108] ), .Y(u1__abc_51895_new_n302_));
INVX1 INVX1_1220 ( .A(u2__abc_52155_new_n5578_), .Y(u2__abc_52155_new_n5579_));
INVX1 INVX1_1221 ( .A(u2_o_380_), .Y(u2__abc_52155_new_n5583_));
INVX1 INVX1_1222 ( .A(u2__abc_52155_new_n5584_), .Y(u2__abc_52155_new_n5585_));
INVX1 INVX1_1223 ( .A(u2_remHi_380_), .Y(u2__abc_52155_new_n5586_));
INVX1 INVX1_1224 ( .A(u2__abc_52155_new_n5587_), .Y(u2__abc_52155_new_n5588_));
INVX1 INVX1_1225 ( .A(u2_remHi_381_), .Y(u2__abc_52155_new_n5590_));
INVX1 INVX1_1226 ( .A(u2__abc_52155_new_n5591_), .Y(u2__abc_52155_new_n5592_));
INVX1 INVX1_1227 ( .A(u2_o_381_), .Y(u2__abc_52155_new_n5593_));
INVX1 INVX1_1228 ( .A(u2__abc_52155_new_n5594_), .Y(u2__abc_52155_new_n5595_));
INVX1 INVX1_1229 ( .A(u2_o_378_), .Y(u2__abc_52155_new_n5598_));
INVX1 INVX1_123 ( .A(\a[109] ), .Y(u1__abc_51895_new_n303_));
INVX1 INVX1_1230 ( .A(u2__abc_52155_new_n5599_), .Y(u2__abc_52155_new_n5600_));
INVX1 INVX1_1231 ( .A(u2_remHi_378_), .Y(u2__abc_52155_new_n5601_));
INVX1 INVX1_1232 ( .A(u2__abc_52155_new_n5602_), .Y(u2__abc_52155_new_n5603_));
INVX1 INVX1_1233 ( .A(u2_o_379_), .Y(u2__abc_52155_new_n5605_));
INVX1 INVX1_1234 ( .A(u2__abc_52155_new_n5606_), .Y(u2__abc_52155_new_n5607_));
INVX1 INVX1_1235 ( .A(u2_remHi_379_), .Y(u2__abc_52155_new_n5608_));
INVX1 INVX1_1236 ( .A(u2__abc_52155_new_n5609_), .Y(u2__abc_52155_new_n5610_));
INVX1 INVX1_1237 ( .A(u2_remHi_374_), .Y(u2__abc_52155_new_n5614_));
INVX1 INVX1_1238 ( .A(u2__abc_52155_new_n5615_), .Y(u2__abc_52155_new_n5616_));
INVX1 INVX1_1239 ( .A(u2_o_374_), .Y(u2__abc_52155_new_n5617_));
INVX1 INVX1_124 ( .A(\a[98] ), .Y(u1__abc_51895_new_n307_));
INVX1 INVX1_1240 ( .A(u2__abc_52155_new_n5618_), .Y(u2__abc_52155_new_n5619_));
INVX1 INVX1_1241 ( .A(u2_remHi_375_), .Y(u2__abc_52155_new_n5621_));
INVX1 INVX1_1242 ( .A(u2__abc_52155_new_n5622_), .Y(u2__abc_52155_new_n5623_));
INVX1 INVX1_1243 ( .A(u2_o_375_), .Y(u2__abc_52155_new_n5624_));
INVX1 INVX1_1244 ( .A(u2__abc_52155_new_n5625_), .Y(u2__abc_52155_new_n5626_));
INVX1 INVX1_1245 ( .A(u2_o_376_), .Y(u2__abc_52155_new_n5629_));
INVX1 INVX1_1246 ( .A(u2__abc_52155_new_n5630_), .Y(u2__abc_52155_new_n5631_));
INVX1 INVX1_1247 ( .A(u2_remHi_376_), .Y(u2__abc_52155_new_n5632_));
INVX1 INVX1_1248 ( .A(u2__abc_52155_new_n5633_), .Y(u2__abc_52155_new_n5634_));
INVX1 INVX1_1249 ( .A(u2_o_377_), .Y(u2__abc_52155_new_n5636_));
INVX1 INVX1_125 ( .A(\a[99] ), .Y(u1__abc_51895_new_n308_));
INVX1 INVX1_1250 ( .A(u2__abc_52155_new_n5637_), .Y(u2__abc_52155_new_n5638_));
INVX1 INVX1_1251 ( .A(u2_remHi_377_), .Y(u2__abc_52155_new_n5639_));
INVX1 INVX1_1252 ( .A(u2__abc_52155_new_n5640_), .Y(u2__abc_52155_new_n5641_));
INVX1 INVX1_1253 ( .A(u2_o_368_), .Y(u2__abc_52155_new_n5646_));
INVX1 INVX1_1254 ( .A(u2__abc_52155_new_n5647_), .Y(u2__abc_52155_new_n5648_));
INVX1 INVX1_1255 ( .A(u2_remHi_368_), .Y(u2__abc_52155_new_n5649_));
INVX1 INVX1_1256 ( .A(u2__abc_52155_new_n5650_), .Y(u2__abc_52155_new_n5651_));
INVX1 INVX1_1257 ( .A(u2_o_369_), .Y(u2__abc_52155_new_n5653_));
INVX1 INVX1_1258 ( .A(u2__abc_52155_new_n5654_), .Y(u2__abc_52155_new_n5655_));
INVX1 INVX1_1259 ( .A(u2_remHi_369_), .Y(u2__abc_52155_new_n5656_));
INVX1 INVX1_126 ( .A(\a[96] ), .Y(u1__abc_51895_new_n310_));
INVX1 INVX1_1260 ( .A(u2__abc_52155_new_n5657_), .Y(u2__abc_52155_new_n5658_));
INVX1 INVX1_1261 ( .A(u2_o_366_), .Y(u2__abc_52155_new_n5661_));
INVX1 INVX1_1262 ( .A(u2__abc_52155_new_n5662_), .Y(u2__abc_52155_new_n5663_));
INVX1 INVX1_1263 ( .A(u2_remHi_366_), .Y(u2__abc_52155_new_n5664_));
INVX1 INVX1_1264 ( .A(u2__abc_52155_new_n5665_), .Y(u2__abc_52155_new_n5666_));
INVX1 INVX1_1265 ( .A(u2_o_367_), .Y(u2__abc_52155_new_n5668_));
INVX1 INVX1_1266 ( .A(u2__abc_52155_new_n5669_), .Y(u2__abc_52155_new_n5670_));
INVX1 INVX1_1267 ( .A(u2_remHi_367_), .Y(u2__abc_52155_new_n5671_));
INVX1 INVX1_1268 ( .A(u2__abc_52155_new_n5672_), .Y(u2__abc_52155_new_n5673_));
INVX1 INVX1_1269 ( .A(u2_o_372_), .Y(u2__abc_52155_new_n5677_));
INVX1 INVX1_127 ( .A(\a[97] ), .Y(u1__abc_51895_new_n311_));
INVX1 INVX1_1270 ( .A(u2__abc_52155_new_n5678_), .Y(u2__abc_52155_new_n5679_));
INVX1 INVX1_1271 ( .A(u2_remHi_372_), .Y(u2__abc_52155_new_n5680_));
INVX1 INVX1_1272 ( .A(u2__abc_52155_new_n5681_), .Y(u2__abc_52155_new_n5682_));
INVX1 INVX1_1273 ( .A(u2_o_373_), .Y(u2__abc_52155_new_n5684_));
INVX1 INVX1_1274 ( .A(u2__abc_52155_new_n5685_), .Y(u2__abc_52155_new_n5686_));
INVX1 INVX1_1275 ( .A(u2_remHi_373_), .Y(u2__abc_52155_new_n5687_));
INVX1 INVX1_1276 ( .A(u2__abc_52155_new_n5688_), .Y(u2__abc_52155_new_n5689_));
INVX1 INVX1_1277 ( .A(u2_o_371_), .Y(u2__abc_52155_new_n5692_));
INVX1 INVX1_1278 ( .A(u2__abc_52155_new_n5693_), .Y(u2__abc_52155_new_n5694_));
INVX1 INVX1_1279 ( .A(u2_remHi_371_), .Y(u2__abc_52155_new_n5695_));
INVX1 INVX1_128 ( .A(\a[102] ), .Y(u1__abc_51895_new_n314_));
INVX1 INVX1_1280 ( .A(u2__abc_52155_new_n5696_), .Y(u2__abc_52155_new_n5697_));
INVX1 INVX1_1281 ( .A(u2_o_370_), .Y(u2__abc_52155_new_n5699_));
INVX1 INVX1_1282 ( .A(u2__abc_52155_new_n5700_), .Y(u2__abc_52155_new_n5701_));
INVX1 INVX1_1283 ( .A(u2_remHi_370_), .Y(u2__abc_52155_new_n5702_));
INVX1 INVX1_1284 ( .A(u2__abc_52155_new_n5703_), .Y(u2__abc_52155_new_n5704_));
INVX1 INVX1_1285 ( .A(u2_remHi_358_), .Y(u2__abc_52155_new_n5710_));
INVX1 INVX1_1286 ( .A(u2__abc_52155_new_n5711_), .Y(u2__abc_52155_new_n5712_));
INVX1 INVX1_1287 ( .A(u2_o_358_), .Y(u2__abc_52155_new_n5713_));
INVX1 INVX1_1288 ( .A(u2__abc_52155_new_n5714_), .Y(u2__abc_52155_new_n5715_));
INVX1 INVX1_1289 ( .A(u2_remHi_359_), .Y(u2__abc_52155_new_n5717_));
INVX1 INVX1_129 ( .A(\a[103] ), .Y(u1__abc_51895_new_n315_));
INVX1 INVX1_1290 ( .A(u2__abc_52155_new_n5718_), .Y(u2__abc_52155_new_n5719_));
INVX1 INVX1_1291 ( .A(u2_o_359_), .Y(u2__abc_52155_new_n5720_));
INVX1 INVX1_1292 ( .A(u2__abc_52155_new_n5721_), .Y(u2__abc_52155_new_n5722_));
INVX1 INVX1_1293 ( .A(u2_o_360_), .Y(u2__abc_52155_new_n5725_));
INVX1 INVX1_1294 ( .A(u2__abc_52155_new_n5726_), .Y(u2__abc_52155_new_n5727_));
INVX1 INVX1_1295 ( .A(u2_remHi_360_), .Y(u2__abc_52155_new_n5728_));
INVX1 INVX1_1296 ( .A(u2__abc_52155_new_n5729_), .Y(u2__abc_52155_new_n5730_));
INVX1 INVX1_1297 ( .A(u2_o_361_), .Y(u2__abc_52155_new_n5732_));
INVX1 INVX1_1298 ( .A(u2__abc_52155_new_n5733_), .Y(u2__abc_52155_new_n5734_));
INVX1 INVX1_1299 ( .A(u2_remHi_361_), .Y(u2__abc_52155_new_n5735_));
INVX1 INVX1_13 ( .A(_abc_73687_new_n1536_), .Y(_abc_73687_new_n1549_));
INVX1 INVX1_130 ( .A(\a[100] ), .Y(u1__abc_51895_new_n317_));
INVX1 INVX1_1300 ( .A(u2__abc_52155_new_n5736_), .Y(u2__abc_52155_new_n5737_));
INVX1 INVX1_1301 ( .A(u2_o_364_), .Y(u2__abc_52155_new_n5741_));
INVX1 INVX1_1302 ( .A(u2__abc_52155_new_n5742_), .Y(u2__abc_52155_new_n5743_));
INVX1 INVX1_1303 ( .A(u2_remHi_364_), .Y(u2__abc_52155_new_n5744_));
INVX1 INVX1_1304 ( .A(u2__abc_52155_new_n5745_), .Y(u2__abc_52155_new_n5746_));
INVX1 INVX1_1305 ( .A(u2_o_365_), .Y(u2__abc_52155_new_n5748_));
INVX1 INVX1_1306 ( .A(u2__abc_52155_new_n5749_), .Y(u2__abc_52155_new_n5750_));
INVX1 INVX1_1307 ( .A(u2_remHi_365_), .Y(u2__abc_52155_new_n5751_));
INVX1 INVX1_1308 ( .A(u2__abc_52155_new_n5752_), .Y(u2__abc_52155_new_n5753_));
INVX1 INVX1_1309 ( .A(u2_o_362_), .Y(u2__abc_52155_new_n5756_));
INVX1 INVX1_131 ( .A(\a[101] ), .Y(u1__abc_51895_new_n318_));
INVX1 INVX1_1310 ( .A(u2__abc_52155_new_n5757_), .Y(u2__abc_52155_new_n5758_));
INVX1 INVX1_1311 ( .A(u2_remHi_362_), .Y(u2__abc_52155_new_n5759_));
INVX1 INVX1_1312 ( .A(u2__abc_52155_new_n5760_), .Y(u2__abc_52155_new_n5761_));
INVX1 INVX1_1313 ( .A(u2_o_363_), .Y(u2__abc_52155_new_n5763_));
INVX1 INVX1_1314 ( .A(u2__abc_52155_new_n5764_), .Y(u2__abc_52155_new_n5765_));
INVX1 INVX1_1315 ( .A(u2_remHi_363_), .Y(u2__abc_52155_new_n5766_));
INVX1 INVX1_1316 ( .A(u2__abc_52155_new_n5767_), .Y(u2__abc_52155_new_n5768_));
INVX1 INVX1_1317 ( .A(u2_o_352_), .Y(u2__abc_52155_new_n5773_));
INVX1 INVX1_1318 ( .A(u2__abc_52155_new_n5774_), .Y(u2__abc_52155_new_n5775_));
INVX1 INVX1_1319 ( .A(u2_remHi_352_), .Y(u2__abc_52155_new_n5776_));
INVX1 INVX1_132 ( .A(\a[58] ), .Y(u1__abc_51895_new_n324_));
INVX1 INVX1_1320 ( .A(u2__abc_52155_new_n5777_), .Y(u2__abc_52155_new_n5778_));
INVX1 INVX1_1321 ( .A(u2_o_353_), .Y(u2__abc_52155_new_n5780_));
INVX1 INVX1_1322 ( .A(u2__abc_52155_new_n5781_), .Y(u2__abc_52155_new_n5782_));
INVX1 INVX1_1323 ( .A(u2_remHi_353_), .Y(u2__abc_52155_new_n5783_));
INVX1 INVX1_1324 ( .A(u2__abc_52155_new_n5784_), .Y(u2__abc_52155_new_n5785_));
INVX1 INVX1_1325 ( .A(u2_o_350_), .Y(u2__abc_52155_new_n5788_));
INVX1 INVX1_1326 ( .A(u2__abc_52155_new_n5789_), .Y(u2__abc_52155_new_n5790_));
INVX1 INVX1_1327 ( .A(u2_remHi_350_), .Y(u2__abc_52155_new_n5791_));
INVX1 INVX1_1328 ( .A(u2__abc_52155_new_n5792_), .Y(u2__abc_52155_new_n5793_));
INVX1 INVX1_1329 ( .A(u2_o_351_), .Y(u2__abc_52155_new_n5795_));
INVX1 INVX1_133 ( .A(\a[59] ), .Y(u1__abc_51895_new_n325_));
INVX1 INVX1_1330 ( .A(u2__abc_52155_new_n5796_), .Y(u2__abc_52155_new_n5797_));
INVX1 INVX1_1331 ( .A(u2_remHi_351_), .Y(u2__abc_52155_new_n5798_));
INVX1 INVX1_1332 ( .A(u2__abc_52155_new_n5799_), .Y(u2__abc_52155_new_n5800_));
INVX1 INVX1_1333 ( .A(u2_o_356_), .Y(u2__abc_52155_new_n5804_));
INVX1 INVX1_1334 ( .A(u2__abc_52155_new_n5805_), .Y(u2__abc_52155_new_n5806_));
INVX1 INVX1_1335 ( .A(u2_remHi_356_), .Y(u2__abc_52155_new_n5807_));
INVX1 INVX1_1336 ( .A(u2__abc_52155_new_n5808_), .Y(u2__abc_52155_new_n5809_));
INVX1 INVX1_1337 ( .A(u2_o_357_), .Y(u2__abc_52155_new_n5811_));
INVX1 INVX1_1338 ( .A(u2__abc_52155_new_n5812_), .Y(u2__abc_52155_new_n5813_));
INVX1 INVX1_1339 ( .A(u2_remHi_357_), .Y(u2__abc_52155_new_n5814_));
INVX1 INVX1_134 ( .A(\a[56] ), .Y(u1__abc_51895_new_n327_));
INVX1 INVX1_1340 ( .A(u2__abc_52155_new_n5815_), .Y(u2__abc_52155_new_n5816_));
INVX1 INVX1_1341 ( .A(u2_o_354_), .Y(u2__abc_52155_new_n5819_));
INVX1 INVX1_1342 ( .A(u2__abc_52155_new_n5820_), .Y(u2__abc_52155_new_n5821_));
INVX1 INVX1_1343 ( .A(u2_remHi_354_), .Y(u2__abc_52155_new_n5822_));
INVX1 INVX1_1344 ( .A(u2__abc_52155_new_n5823_), .Y(u2__abc_52155_new_n5824_));
INVX1 INVX1_1345 ( .A(u2_o_355_), .Y(u2__abc_52155_new_n5826_));
INVX1 INVX1_1346 ( .A(u2__abc_52155_new_n5827_), .Y(u2__abc_52155_new_n5828_));
INVX1 INVX1_1347 ( .A(u2_remHi_355_), .Y(u2__abc_52155_new_n5829_));
INVX1 INVX1_1348 ( .A(u2__abc_52155_new_n5830_), .Y(u2__abc_52155_new_n5831_));
INVX1 INVX1_1349 ( .A(u2_o_344_), .Y(u2__abc_52155_new_n5838_));
INVX1 INVX1_135 ( .A(\a[57] ), .Y(u1__abc_51895_new_n328_));
INVX1 INVX1_1350 ( .A(u2__abc_52155_new_n5839_), .Y(u2__abc_52155_new_n5840_));
INVX1 INVX1_1351 ( .A(u2_remHi_344_), .Y(u2__abc_52155_new_n5841_));
INVX1 INVX1_1352 ( .A(u2__abc_52155_new_n5842_), .Y(u2__abc_52155_new_n5843_));
INVX1 INVX1_1353 ( .A(u2_o_345_), .Y(u2__abc_52155_new_n5845_));
INVX1 INVX1_1354 ( .A(u2__abc_52155_new_n5846_), .Y(u2__abc_52155_new_n5847_));
INVX1 INVX1_1355 ( .A(u2_remHi_345_), .Y(u2__abc_52155_new_n5848_));
INVX1 INVX1_1356 ( .A(u2__abc_52155_new_n5849_), .Y(u2__abc_52155_new_n5850_));
INVX1 INVX1_1357 ( .A(u2_o_342_), .Y(u2__abc_52155_new_n5853_));
INVX1 INVX1_1358 ( .A(u2__abc_52155_new_n5854_), .Y(u2__abc_52155_new_n5855_));
INVX1 INVX1_1359 ( .A(u2_remHi_342_), .Y(u2__abc_52155_new_n5856_));
INVX1 INVX1_136 ( .A(\a[62] ), .Y(u1__abc_51895_new_n331_));
INVX1 INVX1_1360 ( .A(u2__abc_52155_new_n5857_), .Y(u2__abc_52155_new_n5858_));
INVX1 INVX1_1361 ( .A(u2_o_343_), .Y(u2__abc_52155_new_n5860_));
INVX1 INVX1_1362 ( .A(u2__abc_52155_new_n5861_), .Y(u2__abc_52155_new_n5862_));
INVX1 INVX1_1363 ( .A(u2_remHi_343_), .Y(u2__abc_52155_new_n5863_));
INVX1 INVX1_1364 ( .A(u2__abc_52155_new_n5864_), .Y(u2__abc_52155_new_n5865_));
INVX1 INVX1_1365 ( .A(u2_o_348_), .Y(u2__abc_52155_new_n5869_));
INVX1 INVX1_1366 ( .A(u2__abc_52155_new_n5870_), .Y(u2__abc_52155_new_n5871_));
INVX1 INVX1_1367 ( .A(u2_remHi_348_), .Y(u2__abc_52155_new_n5872_));
INVX1 INVX1_1368 ( .A(u2__abc_52155_new_n5873_), .Y(u2__abc_52155_new_n5874_));
INVX1 INVX1_1369 ( .A(u2_o_349_), .Y(u2__abc_52155_new_n5876_));
INVX1 INVX1_137 ( .A(\a[63] ), .Y(u1__abc_51895_new_n332_));
INVX1 INVX1_1370 ( .A(u2__abc_52155_new_n5877_), .Y(u2__abc_52155_new_n5878_));
INVX1 INVX1_1371 ( .A(u2_remHi_349_), .Y(u2__abc_52155_new_n5879_));
INVX1 INVX1_1372 ( .A(u2__abc_52155_new_n5880_), .Y(u2__abc_52155_new_n5881_));
INVX1 INVX1_1373 ( .A(u2_o_346_), .Y(u2__abc_52155_new_n5884_));
INVX1 INVX1_1374 ( .A(u2__abc_52155_new_n5885_), .Y(u2__abc_52155_new_n5886_));
INVX1 INVX1_1375 ( .A(u2_remHi_346_), .Y(u2__abc_52155_new_n5887_));
INVX1 INVX1_1376 ( .A(u2__abc_52155_new_n5888_), .Y(u2__abc_52155_new_n5889_));
INVX1 INVX1_1377 ( .A(u2_o_347_), .Y(u2__abc_52155_new_n5891_));
INVX1 INVX1_1378 ( .A(u2__abc_52155_new_n5892_), .Y(u2__abc_52155_new_n5893_));
INVX1 INVX1_1379 ( .A(u2_remHi_347_), .Y(u2__abc_52155_new_n5894_));
INVX1 INVX1_138 ( .A(\a[60] ), .Y(u1__abc_51895_new_n334_));
INVX1 INVX1_1380 ( .A(u2__abc_52155_new_n5895_), .Y(u2__abc_52155_new_n5896_));
INVX1 INVX1_1381 ( .A(u2_o_336_), .Y(u2__abc_52155_new_n5901_));
INVX1 INVX1_1382 ( .A(u2__abc_52155_new_n5902_), .Y(u2__abc_52155_new_n5903_));
INVX1 INVX1_1383 ( .A(u2_remHi_336_), .Y(u2__abc_52155_new_n5904_));
INVX1 INVX1_1384 ( .A(u2__abc_52155_new_n5905_), .Y(u2__abc_52155_new_n5906_));
INVX1 INVX1_1385 ( .A(u2_o_337_), .Y(u2__abc_52155_new_n5908_));
INVX1 INVX1_1386 ( .A(u2__abc_52155_new_n5909_), .Y(u2__abc_52155_new_n5910_));
INVX1 INVX1_1387 ( .A(u2_remHi_337_), .Y(u2__abc_52155_new_n5911_));
INVX1 INVX1_1388 ( .A(u2__abc_52155_new_n5912_), .Y(u2__abc_52155_new_n5913_));
INVX1 INVX1_1389 ( .A(u2_o_334_), .Y(u2__abc_52155_new_n5916_));
INVX1 INVX1_139 ( .A(\a[61] ), .Y(u1__abc_51895_new_n335_));
INVX1 INVX1_1390 ( .A(u2__abc_52155_new_n5917_), .Y(u2__abc_52155_new_n5918_));
INVX1 INVX1_1391 ( .A(u2_remHi_334_), .Y(u2__abc_52155_new_n5919_));
INVX1 INVX1_1392 ( .A(u2__abc_52155_new_n5920_), .Y(u2__abc_52155_new_n5921_));
INVX1 INVX1_1393 ( .A(u2_o_335_), .Y(u2__abc_52155_new_n5923_));
INVX1 INVX1_1394 ( .A(u2__abc_52155_new_n5924_), .Y(u2__abc_52155_new_n5925_));
INVX1 INVX1_1395 ( .A(u2_remHi_335_), .Y(u2__abc_52155_new_n5926_));
INVX1 INVX1_1396 ( .A(u2__abc_52155_new_n5927_), .Y(u2__abc_52155_new_n5928_));
INVX1 INVX1_1397 ( .A(u2_o_340_), .Y(u2__abc_52155_new_n5932_));
INVX1 INVX1_1398 ( .A(u2__abc_52155_new_n5933_), .Y(u2__abc_52155_new_n5934_));
INVX1 INVX1_1399 ( .A(u2_remHi_340_), .Y(u2__abc_52155_new_n5935_));
INVX1 INVX1_14 ( .A(_abc_73687_new_n1541_), .Y(_abc_73687_new_n1554_));
INVX1 INVX1_140 ( .A(\a[50] ), .Y(u1__abc_51895_new_n339_));
INVX1 INVX1_1400 ( .A(u2__abc_52155_new_n5936_), .Y(u2__abc_52155_new_n5937_));
INVX1 INVX1_1401 ( .A(u2_o_341_), .Y(u2__abc_52155_new_n5939_));
INVX1 INVX1_1402 ( .A(u2__abc_52155_new_n5940_), .Y(u2__abc_52155_new_n5941_));
INVX1 INVX1_1403 ( .A(u2_remHi_341_), .Y(u2__abc_52155_new_n5942_));
INVX1 INVX1_1404 ( .A(u2__abc_52155_new_n5943_), .Y(u2__abc_52155_new_n5944_));
INVX1 INVX1_1405 ( .A(u2_o_338_), .Y(u2__abc_52155_new_n5947_));
INVX1 INVX1_1406 ( .A(u2__abc_52155_new_n5948_), .Y(u2__abc_52155_new_n5949_));
INVX1 INVX1_1407 ( .A(u2_remHi_338_), .Y(u2__abc_52155_new_n5950_));
INVX1 INVX1_1408 ( .A(u2__abc_52155_new_n5951_), .Y(u2__abc_52155_new_n5952_));
INVX1 INVX1_1409 ( .A(u2_o_339_), .Y(u2__abc_52155_new_n5954_));
INVX1 INVX1_141 ( .A(\a[51] ), .Y(u1__abc_51895_new_n340_));
INVX1 INVX1_1410 ( .A(u2__abc_52155_new_n5955_), .Y(u2__abc_52155_new_n5956_));
INVX1 INVX1_1411 ( .A(u2_remHi_339_), .Y(u2__abc_52155_new_n5957_));
INVX1 INVX1_1412 ( .A(u2__abc_52155_new_n5958_), .Y(u2__abc_52155_new_n5959_));
INVX1 INVX1_1413 ( .A(u2_remHi_326_), .Y(u2__abc_52155_new_n5965_));
INVX1 INVX1_1414 ( .A(u2__abc_52155_new_n5966_), .Y(u2__abc_52155_new_n5967_));
INVX1 INVX1_1415 ( .A(u2_o_326_), .Y(u2__abc_52155_new_n5968_));
INVX1 INVX1_1416 ( .A(u2__abc_52155_new_n5969_), .Y(u2__abc_52155_new_n5970_));
INVX1 INVX1_1417 ( .A(u2_remHi_327_), .Y(u2__abc_52155_new_n5972_));
INVX1 INVX1_1418 ( .A(u2__abc_52155_new_n5973_), .Y(u2__abc_52155_new_n5974_));
INVX1 INVX1_1419 ( .A(u2_o_327_), .Y(u2__abc_52155_new_n5975_));
INVX1 INVX1_142 ( .A(\a[48] ), .Y(u1__abc_51895_new_n342_));
INVX1 INVX1_1420 ( .A(u2__abc_52155_new_n5976_), .Y(u2__abc_52155_new_n5977_));
INVX1 INVX1_1421 ( .A(u2_o_328_), .Y(u2__abc_52155_new_n5980_));
INVX1 INVX1_1422 ( .A(u2__abc_52155_new_n5981_), .Y(u2__abc_52155_new_n5982_));
INVX1 INVX1_1423 ( .A(u2_remHi_328_), .Y(u2__abc_52155_new_n5983_));
INVX1 INVX1_1424 ( .A(u2__abc_52155_new_n5984_), .Y(u2__abc_52155_new_n5985_));
INVX1 INVX1_1425 ( .A(u2_o_329_), .Y(u2__abc_52155_new_n5987_));
INVX1 INVX1_1426 ( .A(u2__abc_52155_new_n5988_), .Y(u2__abc_52155_new_n5989_));
INVX1 INVX1_1427 ( .A(u2_remHi_329_), .Y(u2__abc_52155_new_n5990_));
INVX1 INVX1_1428 ( .A(u2__abc_52155_new_n5991_), .Y(u2__abc_52155_new_n5992_));
INVX1 INVX1_1429 ( .A(u2_o_332_), .Y(u2__abc_52155_new_n5996_));
INVX1 INVX1_143 ( .A(\a[49] ), .Y(u1__abc_51895_new_n343_));
INVX1 INVX1_1430 ( .A(u2__abc_52155_new_n5997_), .Y(u2__abc_52155_new_n5998_));
INVX1 INVX1_1431 ( .A(u2_remHi_332_), .Y(u2__abc_52155_new_n5999_));
INVX1 INVX1_1432 ( .A(u2__abc_52155_new_n6000_), .Y(u2__abc_52155_new_n6001_));
INVX1 INVX1_1433 ( .A(u2_o_333_), .Y(u2__abc_52155_new_n6003_));
INVX1 INVX1_1434 ( .A(u2__abc_52155_new_n6004_), .Y(u2__abc_52155_new_n6005_));
INVX1 INVX1_1435 ( .A(u2_remHi_333_), .Y(u2__abc_52155_new_n6006_));
INVX1 INVX1_1436 ( .A(u2__abc_52155_new_n6007_), .Y(u2__abc_52155_new_n6008_));
INVX1 INVX1_1437 ( .A(u2_o_330_), .Y(u2__abc_52155_new_n6011_));
INVX1 INVX1_1438 ( .A(u2__abc_52155_new_n6012_), .Y(u2__abc_52155_new_n6013_));
INVX1 INVX1_1439 ( .A(u2_remHi_330_), .Y(u2__abc_52155_new_n6014_));
INVX1 INVX1_144 ( .A(\a[54] ), .Y(u1__abc_51895_new_n346_));
INVX1 INVX1_1440 ( .A(u2__abc_52155_new_n6015_), .Y(u2__abc_52155_new_n6016_));
INVX1 INVX1_1441 ( .A(u2_o_331_), .Y(u2__abc_52155_new_n6018_));
INVX1 INVX1_1442 ( .A(u2__abc_52155_new_n6019_), .Y(u2__abc_52155_new_n6020_));
INVX1 INVX1_1443 ( .A(u2_remHi_331_), .Y(u2__abc_52155_new_n6021_));
INVX1 INVX1_1444 ( .A(u2__abc_52155_new_n6022_), .Y(u2__abc_52155_new_n6023_));
INVX1 INVX1_1445 ( .A(u2_remHi_324_), .Y(u2__abc_52155_new_n6028_));
INVX1 INVX1_1446 ( .A(u2__abc_52155_new_n6029_), .Y(u2__abc_52155_new_n6030_));
INVX1 INVX1_1447 ( .A(u2_o_324_), .Y(u2__abc_52155_new_n6031_));
INVX1 INVX1_1448 ( .A(u2__abc_52155_new_n6032_), .Y(u2__abc_52155_new_n6033_));
INVX1 INVX1_1449 ( .A(u2_remHi_325_), .Y(u2__abc_52155_new_n6035_));
INVX1 INVX1_145 ( .A(\a[55] ), .Y(u1__abc_51895_new_n347_));
INVX1 INVX1_1450 ( .A(u2__abc_52155_new_n6036_), .Y(u2__abc_52155_new_n6037_));
INVX1 INVX1_1451 ( .A(u2_o_325_), .Y(u2__abc_52155_new_n6038_));
INVX1 INVX1_1452 ( .A(u2__abc_52155_new_n6039_), .Y(u2__abc_52155_new_n6040_));
INVX1 INVX1_1453 ( .A(u2_o_322_), .Y(u2__abc_52155_new_n6043_));
INVX1 INVX1_1454 ( .A(u2__abc_52155_new_n6044_), .Y(u2__abc_52155_new_n6045_));
INVX1 INVX1_1455 ( .A(u2_remHi_322_), .Y(u2__abc_52155_new_n6046_));
INVX1 INVX1_1456 ( .A(u2__abc_52155_new_n6047_), .Y(u2__abc_52155_new_n6048_));
INVX1 INVX1_1457 ( .A(u2_o_323_), .Y(u2__abc_52155_new_n6050_));
INVX1 INVX1_1458 ( .A(u2__abc_52155_new_n6051_), .Y(u2__abc_52155_new_n6052_));
INVX1 INVX1_1459 ( .A(u2_remHi_323_), .Y(u2__abc_52155_new_n6053_));
INVX1 INVX1_146 ( .A(\a[52] ), .Y(u1__abc_51895_new_n349_));
INVX1 INVX1_1460 ( .A(u2__abc_52155_new_n6054_), .Y(u2__abc_52155_new_n6055_));
INVX1 INVX1_1461 ( .A(u2_remHi_318_), .Y(u2__abc_52155_new_n6059_));
INVX1 INVX1_1462 ( .A(u2__abc_52155_new_n6060_), .Y(u2__abc_52155_new_n6061_));
INVX1 INVX1_1463 ( .A(u2_o_318_), .Y(u2__abc_52155_new_n6062_));
INVX1 INVX1_1464 ( .A(u2__abc_52155_new_n6063_), .Y(u2__abc_52155_new_n6064_));
INVX1 INVX1_1465 ( .A(u2_remHi_319_), .Y(u2__abc_52155_new_n6066_));
INVX1 INVX1_1466 ( .A(u2__abc_52155_new_n6067_), .Y(u2__abc_52155_new_n6068_));
INVX1 INVX1_1467 ( .A(u2_o_319_), .Y(u2__abc_52155_new_n6069_));
INVX1 INVX1_1468 ( .A(u2__abc_52155_new_n6070_), .Y(u2__abc_52155_new_n6071_));
INVX1 INVX1_1469 ( .A(u2_o_320_), .Y(u2__abc_52155_new_n6074_));
INVX1 INVX1_147 ( .A(\a[53] ), .Y(u1__abc_51895_new_n350_));
INVX1 INVX1_1470 ( .A(u2__abc_52155_new_n6075_), .Y(u2__abc_52155_new_n6076_));
INVX1 INVX1_1471 ( .A(u2_remHi_320_), .Y(u2__abc_52155_new_n6077_));
INVX1 INVX1_1472 ( .A(u2__abc_52155_new_n6078_), .Y(u2__abc_52155_new_n6079_));
INVX1 INVX1_1473 ( .A(u2_o_321_), .Y(u2__abc_52155_new_n6081_));
INVX1 INVX1_1474 ( .A(u2__abc_52155_new_n6082_), .Y(u2__abc_52155_new_n6083_));
INVX1 INVX1_1475 ( .A(u2_remHi_321_), .Y(u2__abc_52155_new_n6084_));
INVX1 INVX1_1476 ( .A(u2__abc_52155_new_n6085_), .Y(u2__abc_52155_new_n6086_));
INVX1 INVX1_1477 ( .A(u2_o_312_), .Y(u2__abc_52155_new_n6094_));
INVX1 INVX1_1478 ( .A(u2__abc_52155_new_n6095_), .Y(u2__abc_52155_new_n6096_));
INVX1 INVX1_1479 ( .A(u2_remHi_312_), .Y(u2__abc_52155_new_n6097_));
INVX1 INVX1_148 ( .A(\a[74] ), .Y(u1__abc_51895_new_n355_));
INVX1 INVX1_1480 ( .A(u2__abc_52155_new_n6098_), .Y(u2__abc_52155_new_n6099_));
INVX1 INVX1_1481 ( .A(u2_o_313_), .Y(u2__abc_52155_new_n6101_));
INVX1 INVX1_1482 ( .A(u2__abc_52155_new_n6102_), .Y(u2__abc_52155_new_n6103_));
INVX1 INVX1_1483 ( .A(u2_remHi_313_), .Y(u2__abc_52155_new_n6104_));
INVX1 INVX1_1484 ( .A(u2__abc_52155_new_n6105_), .Y(u2__abc_52155_new_n6106_));
INVX1 INVX1_1485 ( .A(u2_o_310_), .Y(u2__abc_52155_new_n6109_));
INVX1 INVX1_1486 ( .A(u2__abc_52155_new_n6110_), .Y(u2__abc_52155_new_n6111_));
INVX1 INVX1_1487 ( .A(u2_remHi_310_), .Y(u2__abc_52155_new_n6112_));
INVX1 INVX1_1488 ( .A(u2__abc_52155_new_n6113_), .Y(u2__abc_52155_new_n6114_));
INVX1 INVX1_1489 ( .A(u2_o_311_), .Y(u2__abc_52155_new_n6116_));
INVX1 INVX1_149 ( .A(\a[75] ), .Y(u1__abc_51895_new_n356_));
INVX1 INVX1_1490 ( .A(u2__abc_52155_new_n6117_), .Y(u2__abc_52155_new_n6118_));
INVX1 INVX1_1491 ( .A(u2_remHi_311_), .Y(u2__abc_52155_new_n6119_));
INVX1 INVX1_1492 ( .A(u2__abc_52155_new_n6120_), .Y(u2__abc_52155_new_n6121_));
INVX1 INVX1_1493 ( .A(u2_o_316_), .Y(u2__abc_52155_new_n6125_));
INVX1 INVX1_1494 ( .A(u2__abc_52155_new_n6126_), .Y(u2__abc_52155_new_n6127_));
INVX1 INVX1_1495 ( .A(u2_remHi_316_), .Y(u2__abc_52155_new_n6128_));
INVX1 INVX1_1496 ( .A(u2__abc_52155_new_n6129_), .Y(u2__abc_52155_new_n6130_));
INVX1 INVX1_1497 ( .A(u2_o_317_), .Y(u2__abc_52155_new_n6132_));
INVX1 INVX1_1498 ( .A(u2__abc_52155_new_n6133_), .Y(u2__abc_52155_new_n6134_));
INVX1 INVX1_1499 ( .A(u2_remHi_317_), .Y(u2__abc_52155_new_n6135_));
INVX1 INVX1_15 ( .A(_abc_73687_new_n1552_), .Y(_abc_73687_new_n1555_));
INVX1 INVX1_150 ( .A(\a[72] ), .Y(u1__abc_51895_new_n358_));
INVX1 INVX1_1500 ( .A(u2__abc_52155_new_n6136_), .Y(u2__abc_52155_new_n6137_));
INVX1 INVX1_1501 ( .A(u2_o_314_), .Y(u2__abc_52155_new_n6140_));
INVX1 INVX1_1502 ( .A(u2__abc_52155_new_n6141_), .Y(u2__abc_52155_new_n6142_));
INVX1 INVX1_1503 ( .A(u2_remHi_314_), .Y(u2__abc_52155_new_n6143_));
INVX1 INVX1_1504 ( .A(u2__abc_52155_new_n6144_), .Y(u2__abc_52155_new_n6145_));
INVX1 INVX1_1505 ( .A(u2_o_315_), .Y(u2__abc_52155_new_n6147_));
INVX1 INVX1_1506 ( .A(u2__abc_52155_new_n6148_), .Y(u2__abc_52155_new_n6149_));
INVX1 INVX1_1507 ( .A(u2_remHi_315_), .Y(u2__abc_52155_new_n6150_));
INVX1 INVX1_1508 ( .A(u2__abc_52155_new_n6151_), .Y(u2__abc_52155_new_n6152_));
INVX1 INVX1_1509 ( .A(u2_remHi_302_), .Y(u2__abc_52155_new_n6157_));
INVX1 INVX1_151 ( .A(\a[73] ), .Y(u1__abc_51895_new_n359_));
INVX1 INVX1_1510 ( .A(u2__abc_52155_new_n6158_), .Y(u2__abc_52155_new_n6159_));
INVX1 INVX1_1511 ( .A(u2_o_302_), .Y(u2__abc_52155_new_n6160_));
INVX1 INVX1_1512 ( .A(u2__abc_52155_new_n6161_), .Y(u2__abc_52155_new_n6162_));
INVX1 INVX1_1513 ( .A(u2_remHi_303_), .Y(u2__abc_52155_new_n6164_));
INVX1 INVX1_1514 ( .A(u2__abc_52155_new_n6165_), .Y(u2__abc_52155_new_n6166_));
INVX1 INVX1_1515 ( .A(u2_o_303_), .Y(u2__abc_52155_new_n6167_));
INVX1 INVX1_1516 ( .A(u2__abc_52155_new_n6168_), .Y(u2__abc_52155_new_n6169_));
INVX1 INVX1_1517 ( .A(u2_o_304_), .Y(u2__abc_52155_new_n6172_));
INVX1 INVX1_1518 ( .A(u2__abc_52155_new_n6173_), .Y(u2__abc_52155_new_n6174_));
INVX1 INVX1_1519 ( .A(u2_remHi_304_), .Y(u2__abc_52155_new_n6175_));
INVX1 INVX1_152 ( .A(\a[78] ), .Y(u1__abc_51895_new_n362_));
INVX1 INVX1_1520 ( .A(u2__abc_52155_new_n6176_), .Y(u2__abc_52155_new_n6177_));
INVX1 INVX1_1521 ( .A(u2_o_305_), .Y(u2__abc_52155_new_n6179_));
INVX1 INVX1_1522 ( .A(u2__abc_52155_new_n6180_), .Y(u2__abc_52155_new_n6181_));
INVX1 INVX1_1523 ( .A(u2_remHi_305_), .Y(u2__abc_52155_new_n6182_));
INVX1 INVX1_1524 ( .A(u2__abc_52155_new_n6183_), .Y(u2__abc_52155_new_n6184_));
INVX1 INVX1_1525 ( .A(u2_o_308_), .Y(u2__abc_52155_new_n6188_));
INVX1 INVX1_1526 ( .A(u2__abc_52155_new_n6189_), .Y(u2__abc_52155_new_n6190_));
INVX1 INVX1_1527 ( .A(u2_remHi_308_), .Y(u2__abc_52155_new_n6191_));
INVX1 INVX1_1528 ( .A(u2__abc_52155_new_n6192_), .Y(u2__abc_52155_new_n6193_));
INVX1 INVX1_1529 ( .A(u2_o_309_), .Y(u2__abc_52155_new_n6195_));
INVX1 INVX1_153 ( .A(\a[79] ), .Y(u1__abc_51895_new_n363_));
INVX1 INVX1_1530 ( .A(u2__abc_52155_new_n6196_), .Y(u2__abc_52155_new_n6197_));
INVX1 INVX1_1531 ( .A(u2_remHi_309_), .Y(u2__abc_52155_new_n6198_));
INVX1 INVX1_1532 ( .A(u2__abc_52155_new_n6199_), .Y(u2__abc_52155_new_n6200_));
INVX1 INVX1_1533 ( .A(u2_o_307_), .Y(u2__abc_52155_new_n6203_));
INVX1 INVX1_1534 ( .A(u2__abc_52155_new_n6204_), .Y(u2__abc_52155_new_n6205_));
INVX1 INVX1_1535 ( .A(u2_remHi_307_), .Y(u2__abc_52155_new_n6206_));
INVX1 INVX1_1536 ( .A(u2__abc_52155_new_n6207_), .Y(u2__abc_52155_new_n6208_));
INVX1 INVX1_1537 ( .A(u2_o_306_), .Y(u2__abc_52155_new_n6210_));
INVX1 INVX1_1538 ( .A(u2__abc_52155_new_n6211_), .Y(u2__abc_52155_new_n6212_));
INVX1 INVX1_1539 ( .A(u2_remHi_306_), .Y(u2__abc_52155_new_n6213_));
INVX1 INVX1_154 ( .A(\a[76] ), .Y(u1__abc_51895_new_n365_));
INVX1 INVX1_1540 ( .A(u2__abc_52155_new_n6214_), .Y(u2__abc_52155_new_n6215_));
INVX1 INVX1_1541 ( .A(u2_remHi_294_), .Y(u2__abc_52155_new_n6221_));
INVX1 INVX1_1542 ( .A(u2__abc_52155_new_n6222_), .Y(u2__abc_52155_new_n6223_));
INVX1 INVX1_1543 ( .A(u2_o_294_), .Y(u2__abc_52155_new_n6224_));
INVX1 INVX1_1544 ( .A(u2__abc_52155_new_n6225_), .Y(u2__abc_52155_new_n6226_));
INVX1 INVX1_1545 ( .A(u2_remHi_295_), .Y(u2__abc_52155_new_n6228_));
INVX1 INVX1_1546 ( .A(u2__abc_52155_new_n6229_), .Y(u2__abc_52155_new_n6230_));
INVX1 INVX1_1547 ( .A(u2_o_295_), .Y(u2__abc_52155_new_n6231_));
INVX1 INVX1_1548 ( .A(u2__abc_52155_new_n6232_), .Y(u2__abc_52155_new_n6233_));
INVX1 INVX1_1549 ( .A(u2_o_296_), .Y(u2__abc_52155_new_n6236_));
INVX1 INVX1_155 ( .A(\a[77] ), .Y(u1__abc_51895_new_n366_));
INVX1 INVX1_1550 ( .A(u2__abc_52155_new_n6237_), .Y(u2__abc_52155_new_n6238_));
INVX1 INVX1_1551 ( .A(u2_remHi_296_), .Y(u2__abc_52155_new_n6239_));
INVX1 INVX1_1552 ( .A(u2__abc_52155_new_n6240_), .Y(u2__abc_52155_new_n6241_));
INVX1 INVX1_1553 ( .A(u2_o_297_), .Y(u2__abc_52155_new_n6243_));
INVX1 INVX1_1554 ( .A(u2__abc_52155_new_n6244_), .Y(u2__abc_52155_new_n6245_));
INVX1 INVX1_1555 ( .A(u2_remHi_297_), .Y(u2__abc_52155_new_n6246_));
INVX1 INVX1_1556 ( .A(u2__abc_52155_new_n6247_), .Y(u2__abc_52155_new_n6248_));
INVX1 INVX1_1557 ( .A(u2_o_300_), .Y(u2__abc_52155_new_n6252_));
INVX1 INVX1_1558 ( .A(u2__abc_52155_new_n6253_), .Y(u2__abc_52155_new_n6254_));
INVX1 INVX1_1559 ( .A(u2_remHi_300_), .Y(u2__abc_52155_new_n6255_));
INVX1 INVX1_156 ( .A(\a[66] ), .Y(u1__abc_51895_new_n370_));
INVX1 INVX1_1560 ( .A(u2__abc_52155_new_n6256_), .Y(u2__abc_52155_new_n6257_));
INVX1 INVX1_1561 ( .A(u2_o_301_), .Y(u2__abc_52155_new_n6259_));
INVX1 INVX1_1562 ( .A(u2__abc_52155_new_n6260_), .Y(u2__abc_52155_new_n6261_));
INVX1 INVX1_1563 ( .A(u2_remHi_301_), .Y(u2__abc_52155_new_n6262_));
INVX1 INVX1_1564 ( .A(u2__abc_52155_new_n6263_), .Y(u2__abc_52155_new_n6264_));
INVX1 INVX1_1565 ( .A(u2_o_298_), .Y(u2__abc_52155_new_n6267_));
INVX1 INVX1_1566 ( .A(u2__abc_52155_new_n6268_), .Y(u2__abc_52155_new_n6269_));
INVX1 INVX1_1567 ( .A(u2_remHi_298_), .Y(u2__abc_52155_new_n6270_));
INVX1 INVX1_1568 ( .A(u2__abc_52155_new_n6271_), .Y(u2__abc_52155_new_n6272_));
INVX1 INVX1_1569 ( .A(u2_o_299_), .Y(u2__abc_52155_new_n6274_));
INVX1 INVX1_157 ( .A(\a[67] ), .Y(u1__abc_51895_new_n371_));
INVX1 INVX1_1570 ( .A(u2__abc_52155_new_n6275_), .Y(u2__abc_52155_new_n6276_));
INVX1 INVX1_1571 ( .A(u2_remHi_299_), .Y(u2__abc_52155_new_n6277_));
INVX1 INVX1_1572 ( .A(u2__abc_52155_new_n6278_), .Y(u2__abc_52155_new_n6279_));
INVX1 INVX1_1573 ( .A(u2_o_288_), .Y(u2__abc_52155_new_n6284_));
INVX1 INVX1_1574 ( .A(u2__abc_52155_new_n6285_), .Y(u2__abc_52155_new_n6286_));
INVX1 INVX1_1575 ( .A(u2_remHi_288_), .Y(u2__abc_52155_new_n6287_));
INVX1 INVX1_1576 ( .A(u2__abc_52155_new_n6288_), .Y(u2__abc_52155_new_n6289_));
INVX1 INVX1_1577 ( .A(u2_o_289_), .Y(u2__abc_52155_new_n6291_));
INVX1 INVX1_1578 ( .A(u2__abc_52155_new_n6292_), .Y(u2__abc_52155_new_n6293_));
INVX1 INVX1_1579 ( .A(u2_remHi_289_), .Y(u2__abc_52155_new_n6294_));
INVX1 INVX1_158 ( .A(\a[64] ), .Y(u1__abc_51895_new_n373_));
INVX1 INVX1_1580 ( .A(u2__abc_52155_new_n6295_), .Y(u2__abc_52155_new_n6296_));
INVX1 INVX1_1581 ( .A(u2_o_286_), .Y(u2__abc_52155_new_n6299_));
INVX1 INVX1_1582 ( .A(u2__abc_52155_new_n6300_), .Y(u2__abc_52155_new_n6301_));
INVX1 INVX1_1583 ( .A(u2_remHi_286_), .Y(u2__abc_52155_new_n6302_));
INVX1 INVX1_1584 ( .A(u2__abc_52155_new_n6303_), .Y(u2__abc_52155_new_n6304_));
INVX1 INVX1_1585 ( .A(u2_o_287_), .Y(u2__abc_52155_new_n6306_));
INVX1 INVX1_1586 ( .A(u2__abc_52155_new_n6307_), .Y(u2__abc_52155_new_n6308_));
INVX1 INVX1_1587 ( .A(u2_remHi_287_), .Y(u2__abc_52155_new_n6309_));
INVX1 INVX1_1588 ( .A(u2__abc_52155_new_n6310_), .Y(u2__abc_52155_new_n6311_));
INVX1 INVX1_1589 ( .A(u2_o_292_), .Y(u2__abc_52155_new_n6315_));
INVX1 INVX1_159 ( .A(\a[65] ), .Y(u1__abc_51895_new_n374_));
INVX1 INVX1_1590 ( .A(u2__abc_52155_new_n6316_), .Y(u2__abc_52155_new_n6317_));
INVX1 INVX1_1591 ( .A(u2_remHi_292_), .Y(u2__abc_52155_new_n6318_));
INVX1 INVX1_1592 ( .A(u2__abc_52155_new_n6319_), .Y(u2__abc_52155_new_n6320_));
INVX1 INVX1_1593 ( .A(u2_o_293_), .Y(u2__abc_52155_new_n6322_));
INVX1 INVX1_1594 ( .A(u2__abc_52155_new_n6323_), .Y(u2__abc_52155_new_n6324_));
INVX1 INVX1_1595 ( .A(u2_remHi_293_), .Y(u2__abc_52155_new_n6325_));
INVX1 INVX1_1596 ( .A(u2__abc_52155_new_n6326_), .Y(u2__abc_52155_new_n6327_));
INVX1 INVX1_1597 ( .A(u2_o_290_), .Y(u2__abc_52155_new_n6330_));
INVX1 INVX1_1598 ( .A(u2__abc_52155_new_n6331_), .Y(u2__abc_52155_new_n6332_));
INVX1 INVX1_1599 ( .A(u2_remHi_290_), .Y(u2__abc_52155_new_n6333_));
INVX1 INVX1_16 ( .A(\a[118] ), .Y(_abc_73687_new_n1563_));
INVX1 INVX1_160 ( .A(\a[70] ), .Y(u1__abc_51895_new_n377_));
INVX1 INVX1_1600 ( .A(u2__abc_52155_new_n6334_), .Y(u2__abc_52155_new_n6335_));
INVX1 INVX1_1601 ( .A(u2_o_291_), .Y(u2__abc_52155_new_n6337_));
INVX1 INVX1_1602 ( .A(u2__abc_52155_new_n6338_), .Y(u2__abc_52155_new_n6339_));
INVX1 INVX1_1603 ( .A(u2_remHi_291_), .Y(u2__abc_52155_new_n6340_));
INVX1 INVX1_1604 ( .A(u2__abc_52155_new_n6341_), .Y(u2__abc_52155_new_n6342_));
INVX1 INVX1_1605 ( .A(u2_o_280_), .Y(u2__abc_52155_new_n6349_));
INVX1 INVX1_1606 ( .A(u2__abc_52155_new_n6350_), .Y(u2__abc_52155_new_n6351_));
INVX1 INVX1_1607 ( .A(u2_remHi_280_), .Y(u2__abc_52155_new_n6352_));
INVX1 INVX1_1608 ( .A(u2__abc_52155_new_n6353_), .Y(u2__abc_52155_new_n6354_));
INVX1 INVX1_1609 ( .A(u2_o_281_), .Y(u2__abc_52155_new_n6356_));
INVX1 INVX1_161 ( .A(\a[71] ), .Y(u1__abc_51895_new_n378_));
INVX1 INVX1_1610 ( .A(u2__abc_52155_new_n6357_), .Y(u2__abc_52155_new_n6358_));
INVX1 INVX1_1611 ( .A(u2_remHi_281_), .Y(u2__abc_52155_new_n6359_));
INVX1 INVX1_1612 ( .A(u2__abc_52155_new_n6360_), .Y(u2__abc_52155_new_n6361_));
INVX1 INVX1_1613 ( .A(u2_o_278_), .Y(u2__abc_52155_new_n6364_));
INVX1 INVX1_1614 ( .A(u2__abc_52155_new_n6365_), .Y(u2__abc_52155_new_n6366_));
INVX1 INVX1_1615 ( .A(u2_remHi_278_), .Y(u2__abc_52155_new_n6367_));
INVX1 INVX1_1616 ( .A(u2__abc_52155_new_n6368_), .Y(u2__abc_52155_new_n6369_));
INVX1 INVX1_1617 ( .A(u2_o_279_), .Y(u2__abc_52155_new_n6371_));
INVX1 INVX1_1618 ( .A(u2__abc_52155_new_n6372_), .Y(u2__abc_52155_new_n6373_));
INVX1 INVX1_1619 ( .A(u2_remHi_279_), .Y(u2__abc_52155_new_n6374_));
INVX1 INVX1_162 ( .A(\a[68] ), .Y(u1__abc_51895_new_n380_));
INVX1 INVX1_1620 ( .A(u2__abc_52155_new_n6375_), .Y(u2__abc_52155_new_n6376_));
INVX1 INVX1_1621 ( .A(u2_o_284_), .Y(u2__abc_52155_new_n6380_));
INVX1 INVX1_1622 ( .A(u2__abc_52155_new_n6381_), .Y(u2__abc_52155_new_n6382_));
INVX1 INVX1_1623 ( .A(u2_remHi_284_), .Y(u2__abc_52155_new_n6383_));
INVX1 INVX1_1624 ( .A(u2__abc_52155_new_n6384_), .Y(u2__abc_52155_new_n6385_));
INVX1 INVX1_1625 ( .A(u2_o_285_), .Y(u2__abc_52155_new_n6387_));
INVX1 INVX1_1626 ( .A(u2__abc_52155_new_n6388_), .Y(u2__abc_52155_new_n6389_));
INVX1 INVX1_1627 ( .A(u2_remHi_285_), .Y(u2__abc_52155_new_n6390_));
INVX1 INVX1_1628 ( .A(u2__abc_52155_new_n6391_), .Y(u2__abc_52155_new_n6392_));
INVX1 INVX1_1629 ( .A(u2_o_282_), .Y(u2__abc_52155_new_n6395_));
INVX1 INVX1_163 ( .A(\a[69] ), .Y(u1__abc_51895_new_n381_));
INVX1 INVX1_1630 ( .A(u2__abc_52155_new_n6396_), .Y(u2__abc_52155_new_n6397_));
INVX1 INVX1_1631 ( .A(u2_remHi_282_), .Y(u2__abc_52155_new_n6398_));
INVX1 INVX1_1632 ( .A(u2__abc_52155_new_n6399_), .Y(u2__abc_52155_new_n6400_));
INVX1 INVX1_1633 ( .A(u2_o_283_), .Y(u2__abc_52155_new_n6402_));
INVX1 INVX1_1634 ( .A(u2__abc_52155_new_n6403_), .Y(u2__abc_52155_new_n6404_));
INVX1 INVX1_1635 ( .A(u2_remHi_283_), .Y(u2__abc_52155_new_n6405_));
INVX1 INVX1_1636 ( .A(u2__abc_52155_new_n6406_), .Y(u2__abc_52155_new_n6407_));
INVX1 INVX1_1637 ( .A(u2_o_272_), .Y(u2__abc_52155_new_n6412_));
INVX1 INVX1_1638 ( .A(u2__abc_52155_new_n6413_), .Y(u2__abc_52155_new_n6414_));
INVX1 INVX1_1639 ( .A(u2_remHi_272_), .Y(u2__abc_52155_new_n6415_));
INVX1 INVX1_164 ( .A(u1_mz), .Y(u1__abc_51895_new_n392_));
INVX1 INVX1_1640 ( .A(u2__abc_52155_new_n6416_), .Y(u2__abc_52155_new_n6417_));
INVX1 INVX1_1641 ( .A(u2_o_273_), .Y(u2__abc_52155_new_n6419_));
INVX1 INVX1_1642 ( .A(u2__abc_52155_new_n6420_), .Y(u2__abc_52155_new_n6421_));
INVX1 INVX1_1643 ( .A(u2_remHi_273_), .Y(u2__abc_52155_new_n6422_));
INVX1 INVX1_1644 ( .A(u2__abc_52155_new_n6423_), .Y(u2__abc_52155_new_n6424_));
INVX1 INVX1_1645 ( .A(u2_o_270_), .Y(u2__abc_52155_new_n6427_));
INVX1 INVX1_1646 ( .A(u2__abc_52155_new_n6428_), .Y(u2__abc_52155_new_n6429_));
INVX1 INVX1_1647 ( .A(u2_remHi_270_), .Y(u2__abc_52155_new_n6430_));
INVX1 INVX1_1648 ( .A(u2__abc_52155_new_n6431_), .Y(u2__abc_52155_new_n6432_));
INVX1 INVX1_1649 ( .A(u2_o_271_), .Y(u2__abc_52155_new_n6434_));
INVX1 INVX1_165 ( .A(rst), .Y(u2__abc_52155_new_n2962_));
INVX1 INVX1_1650 ( .A(u2__abc_52155_new_n6435_), .Y(u2__abc_52155_new_n6436_));
INVX1 INVX1_1651 ( .A(u2_remHi_271_), .Y(u2__abc_52155_new_n6437_));
INVX1 INVX1_1652 ( .A(u2__abc_52155_new_n6438_), .Y(u2__abc_52155_new_n6439_));
INVX1 INVX1_1653 ( .A(u2_o_276_), .Y(u2__abc_52155_new_n6443_));
INVX1 INVX1_1654 ( .A(u2__abc_52155_new_n6444_), .Y(u2__abc_52155_new_n6445_));
INVX1 INVX1_1655 ( .A(u2_remHi_276_), .Y(u2__abc_52155_new_n6446_));
INVX1 INVX1_1656 ( .A(u2__abc_52155_new_n6447_), .Y(u2__abc_52155_new_n6448_));
INVX1 INVX1_1657 ( .A(u2_o_277_), .Y(u2__abc_52155_new_n6450_));
INVX1 INVX1_1658 ( .A(u2__abc_52155_new_n6451_), .Y(u2__abc_52155_new_n6452_));
INVX1 INVX1_1659 ( .A(u2_remHi_277_), .Y(u2__abc_52155_new_n6453_));
INVX1 INVX1_166 ( .A(u2_cnt_4_), .Y(u2__abc_52155_new_n2965_));
INVX1 INVX1_1660 ( .A(u2__abc_52155_new_n6454_), .Y(u2__abc_52155_new_n6455_));
INVX1 INVX1_1661 ( .A(u2_o_274_), .Y(u2__abc_52155_new_n6458_));
INVX1 INVX1_1662 ( .A(u2__abc_52155_new_n6459_), .Y(u2__abc_52155_new_n6460_));
INVX1 INVX1_1663 ( .A(u2_remHi_274_), .Y(u2__abc_52155_new_n6461_));
INVX1 INVX1_1664 ( .A(u2__abc_52155_new_n6462_), .Y(u2__abc_52155_new_n6463_));
INVX1 INVX1_1665 ( .A(u2_o_275_), .Y(u2__abc_52155_new_n6465_));
INVX1 INVX1_1666 ( .A(u2__abc_52155_new_n6466_), .Y(u2__abc_52155_new_n6467_));
INVX1 INVX1_1667 ( .A(u2_remHi_275_), .Y(u2__abc_52155_new_n6468_));
INVX1 INVX1_1668 ( .A(u2__abc_52155_new_n6469_), .Y(u2__abc_52155_new_n6470_));
INVX1 INVX1_1669 ( .A(u2_remHi_268_), .Y(u2__abc_52155_new_n6476_));
INVX1 INVX1_167 ( .A(u2__abc_52155_new_n2969_), .Y(u2__abc_52155_new_n2970_));
INVX1 INVX1_1670 ( .A(u2__abc_52155_new_n6477_), .Y(u2__abc_52155_new_n6478_));
INVX1 INVX1_1671 ( .A(u2_o_268_), .Y(u2__abc_52155_new_n6479_));
INVX1 INVX1_1672 ( .A(u2__abc_52155_new_n6480_), .Y(u2__abc_52155_new_n6481_));
INVX1 INVX1_1673 ( .A(u2_remHi_269_), .Y(u2__abc_52155_new_n6483_));
INVX1 INVX1_1674 ( .A(u2__abc_52155_new_n6484_), .Y(u2__abc_52155_new_n6485_));
INVX1 INVX1_1675 ( .A(u2_o_269_), .Y(u2__abc_52155_new_n6486_));
INVX1 INVX1_1676 ( .A(u2__abc_52155_new_n6487_), .Y(u2__abc_52155_new_n6488_));
INVX1 INVX1_1677 ( .A(u2_o_266_), .Y(u2__abc_52155_new_n6491_));
INVX1 INVX1_1678 ( .A(u2__abc_52155_new_n6492_), .Y(u2__abc_52155_new_n6493_));
INVX1 INVX1_1679 ( .A(u2_remHi_266_), .Y(u2__abc_52155_new_n6494_));
INVX1 INVX1_168 ( .A(u2_cnt_0_), .Y(u2__abc_52155_new_n2971_));
INVX1 INVX1_1680 ( .A(u2__abc_52155_new_n6495_), .Y(u2__abc_52155_new_n6496_));
INVX1 INVX1_1681 ( .A(u2_o_267_), .Y(u2__abc_52155_new_n6498_));
INVX1 INVX1_1682 ( .A(u2__abc_52155_new_n6499_), .Y(u2__abc_52155_new_n6500_));
INVX1 INVX1_1683 ( .A(u2_remHi_267_), .Y(u2__abc_52155_new_n6501_));
INVX1 INVX1_1684 ( .A(u2__abc_52155_new_n6502_), .Y(u2__abc_52155_new_n6503_));
INVX1 INVX1_1685 ( .A(u2_o_264_), .Y(u2__abc_52155_new_n6507_));
INVX1 INVX1_1686 ( .A(u2__abc_52155_new_n6508_), .Y(u2__abc_52155_new_n6509_));
INVX1 INVX1_1687 ( .A(u2_remHi_264_), .Y(u2__abc_52155_new_n6510_));
INVX1 INVX1_1688 ( .A(u2__abc_52155_new_n6511_), .Y(u2__abc_52155_new_n6512_));
INVX1 INVX1_1689 ( .A(u2_o_265_), .Y(u2__abc_52155_new_n6514_));
INVX1 INVX1_169 ( .A(u2__abc_52155_new_n2975_), .Y(u2__abc_52155_new_n2976_));
INVX1 INVX1_1690 ( .A(u2__abc_52155_new_n6515_), .Y(u2__abc_52155_new_n6516_));
INVX1 INVX1_1691 ( .A(u2_remHi_265_), .Y(u2__abc_52155_new_n6517_));
INVX1 INVX1_1692 ( .A(u2__abc_52155_new_n6518_), .Y(u2__abc_52155_new_n6519_));
INVX1 INVX1_1693 ( .A(u2_remHi_262_), .Y(u2__abc_52155_new_n6522_));
INVX1 INVX1_1694 ( .A(u2__abc_52155_new_n6523_), .Y(u2__abc_52155_new_n6524_));
INVX1 INVX1_1695 ( .A(u2_o_262_), .Y(u2__abc_52155_new_n6525_));
INVX1 INVX1_1696 ( .A(u2__abc_52155_new_n6526_), .Y(u2__abc_52155_new_n6527_));
INVX1 INVX1_1697 ( .A(u2_remHi_263_), .Y(u2__abc_52155_new_n6529_));
INVX1 INVX1_1698 ( .A(u2__abc_52155_new_n6530_), .Y(u2__abc_52155_new_n6531_));
INVX1 INVX1_1699 ( .A(u2_o_263_), .Y(u2__abc_52155_new_n6532_));
INVX1 INVX1_17 ( .A(_abc_73687_new_n1551_), .Y(_abc_73687_new_n1564_));
INVX1 INVX1_170 ( .A(u2__abc_52155_new_n2982_), .Y(u2__abc_52155_new_n2983_));
INVX1 INVX1_1700 ( .A(u2__abc_52155_new_n6533_), .Y(u2__abc_52155_new_n6534_));
INVX1 INVX1_1701 ( .A(u2_remHi_254_), .Y(u2__abc_52155_new_n6539_));
INVX1 INVX1_1702 ( .A(u2__abc_52155_new_n6540_), .Y(u2__abc_52155_new_n6541_));
INVX1 INVX1_1703 ( .A(u2_o_254_), .Y(u2__abc_52155_new_n6542_));
INVX1 INVX1_1704 ( .A(u2__abc_52155_new_n6543_), .Y(u2__abc_52155_new_n6544_));
INVX1 INVX1_1705 ( .A(u2_remHi_255_), .Y(u2__abc_52155_new_n6546_));
INVX1 INVX1_1706 ( .A(u2__abc_52155_new_n6547_), .Y(u2__abc_52155_new_n6548_));
INVX1 INVX1_1707 ( .A(u2_o_255_), .Y(u2__abc_52155_new_n6549_));
INVX1 INVX1_1708 ( .A(u2__abc_52155_new_n6550_), .Y(u2__abc_52155_new_n6551_));
INVX1 INVX1_1709 ( .A(u2_o_256_), .Y(u2__abc_52155_new_n6554_));
INVX1 INVX1_171 ( .A(ld), .Y(u2__abc_52155_new_n2984_));
INVX1 INVX1_1710 ( .A(u2__abc_52155_new_n6555_), .Y(u2__abc_52155_new_n6556_));
INVX1 INVX1_1711 ( .A(u2_remHi_256_), .Y(u2__abc_52155_new_n6557_));
INVX1 INVX1_1712 ( .A(u2__abc_52155_new_n6558_), .Y(u2__abc_52155_new_n6559_));
INVX1 INVX1_1713 ( .A(u2_o_257_), .Y(u2__abc_52155_new_n6561_));
INVX1 INVX1_1714 ( .A(u2__abc_52155_new_n6562_), .Y(u2__abc_52155_new_n6563_));
INVX1 INVX1_1715 ( .A(u2_remHi_257_), .Y(u2__abc_52155_new_n6564_));
INVX1 INVX1_1716 ( .A(u2__abc_52155_new_n6565_), .Y(u2__abc_52155_new_n6566_));
INVX1 INVX1_1717 ( .A(u2_o_260_), .Y(u2__abc_52155_new_n6570_));
INVX1 INVX1_1718 ( .A(u2__abc_52155_new_n6571_), .Y(u2__abc_52155_new_n6572_));
INVX1 INVX1_1719 ( .A(u2_remHi_260_), .Y(u2__abc_52155_new_n6573_));
INVX1 INVX1_172 ( .A(u2__abc_52155_new_n2980_), .Y(u2__abc_52155_new_n2989_));
INVX1 INVX1_1720 ( .A(u2__abc_52155_new_n6574_), .Y(u2__abc_52155_new_n6575_));
INVX1 INVX1_1721 ( .A(u2_o_261_), .Y(u2__abc_52155_new_n6577_));
INVX1 INVX1_1722 ( .A(u2__abc_52155_new_n6578_), .Y(u2__abc_52155_new_n6579_));
INVX1 INVX1_1723 ( .A(u2_remHi_261_), .Y(u2__abc_52155_new_n6580_));
INVX1 INVX1_1724 ( .A(u2__abc_52155_new_n6581_), .Y(u2__abc_52155_new_n6582_));
INVX1 INVX1_1725 ( .A(u2_o_258_), .Y(u2__abc_52155_new_n6585_));
INVX1 INVX1_1726 ( .A(u2__abc_52155_new_n6586_), .Y(u2__abc_52155_new_n6587_));
INVX1 INVX1_1727 ( .A(u2_remHi_258_), .Y(u2__abc_52155_new_n6588_));
INVX1 INVX1_1728 ( .A(u2__abc_52155_new_n6589_), .Y(u2__abc_52155_new_n6590_));
INVX1 INVX1_1729 ( .A(u2_o_259_), .Y(u2__abc_52155_new_n6592_));
INVX1 INVX1_173 ( .A(u2__abc_52155_new_n2997_), .Y(u2__abc_52155_new_n2998_));
INVX1 INVX1_1730 ( .A(u2__abc_52155_new_n6593_), .Y(u2__abc_52155_new_n6594_));
INVX1 INVX1_1731 ( .A(u2_remHi_259_), .Y(u2__abc_52155_new_n6595_));
INVX1 INVX1_1732 ( .A(u2__abc_52155_new_n6596_), .Y(u2__abc_52155_new_n6597_));
INVX1 INVX1_1733 ( .A(u2__abc_52155_new_n6605_), .Y(u2__abc_52155_new_n6606_));
INVX1 INVX1_1734 ( .A(u2__abc_52155_new_n6093_), .Y(u2__abc_52155_new_n6608_));
INVX1 INVX1_1735 ( .A(u2__abc_52155_new_n6348_), .Y(u2__abc_52155_new_n6609_));
INVX1 INVX1_1736 ( .A(u2__abc_52155_new_n6411_), .Y(u2__abc_52155_new_n6610_));
INVX1 INVX1_1737 ( .A(u2__abc_52155_new_n6426_), .Y(u2__abc_52155_new_n6614_));
INVX1 INVX1_1738 ( .A(u2__abc_52155_new_n6619_), .Y(u2__abc_52155_new_n6620_));
INVX1 INVX1_1739 ( .A(u2__abc_52155_new_n6457_), .Y(u2__abc_52155_new_n6624_));
INVX1 INVX1_174 ( .A(u2__abc_52155_new_n2999_), .Y(u2__abc_52155_new_n3000_));
INVX1 INVX1_1740 ( .A(u2__abc_52155_new_n6475_), .Y(u2__abc_52155_new_n6629_));
INVX1 INVX1_1741 ( .A(u2__abc_52155_new_n6538_), .Y(u2__abc_52155_new_n6630_));
INVX1 INVX1_1742 ( .A(u2__abc_52155_new_n6600_), .Y(u2__abc_52155_new_n6631_));
INVX1 INVX1_1743 ( .A(u2__abc_52155_new_n6568_), .Y(u2__abc_52155_new_n6632_));
INVX1 INVX1_1744 ( .A(u2__abc_52155_new_n6637_), .Y(u2__abc_52155_new_n6638_));
INVX1 INVX1_1745 ( .A(u2__abc_52155_new_n6584_), .Y(u2__abc_52155_new_n6641_));
INVX1 INVX1_1746 ( .A(u2__abc_52155_new_n6646_), .Y(u2__abc_52155_new_n6647_));
INVX1 INVX1_1747 ( .A(u2__abc_52155_new_n6506_), .Y(u2__abc_52155_new_n6651_));
INVX1 INVX1_1748 ( .A(u2__abc_52155_new_n6521_), .Y(u2__abc_52155_new_n6652_));
INVX1 INVX1_1749 ( .A(u2__abc_52155_new_n6657_), .Y(u2__abc_52155_new_n6658_));
INVX1 INVX1_175 ( .A(u2_remHi_449_), .Y(u2__abc_52155_new_n3004_));
INVX1 INVX1_1750 ( .A(u2__abc_52155_new_n6490_), .Y(u2__abc_52155_new_n6663_));
INVX1 INVX1_1751 ( .A(u2__abc_52155_new_n6410_), .Y(u2__abc_52155_new_n6671_));
INVX1 INVX1_1752 ( .A(u2__abc_52155_new_n6363_), .Y(u2__abc_52155_new_n6672_));
INVX1 INVX1_1753 ( .A(u2__abc_52155_new_n6677_), .Y(u2__abc_52155_new_n6678_));
INVX1 INVX1_1754 ( .A(u2__abc_52155_new_n6394_), .Y(u2__abc_52155_new_n6681_));
INVX1 INVX1_1755 ( .A(u2__abc_52155_new_n6156_), .Y(u2__abc_52155_new_n6692_));
INVX1 INVX1_1756 ( .A(u2__abc_52155_new_n6186_), .Y(u2__abc_52155_new_n6694_));
INVX1 INVX1_1757 ( .A(u2__abc_52155_new_n6699_), .Y(u2__abc_52155_new_n6700_));
INVX1 INVX1_1758 ( .A(u2__abc_52155_new_n6220_), .Y(u2__abc_52155_new_n6724_));
INVX1 INVX1_1759 ( .A(u2__abc_52155_new_n6283_), .Y(u2__abc_52155_new_n6725_));
INVX1 INVX1_176 ( .A(u2__abc_52155_new_n3005_), .Y(u2__abc_52155_new_n3006_));
INVX1 INVX1_1760 ( .A(u2__abc_52155_new_n6345_), .Y(u2__abc_52155_new_n6726_));
INVX1 INVX1_1761 ( .A(u2__abc_52155_new_n6298_), .Y(u2__abc_52155_new_n6729_));
INVX1 INVX1_1762 ( .A(u2__abc_52155_new_n6329_), .Y(u2__abc_52155_new_n6735_));
INVX1 INVX1_1763 ( .A(u2__abc_52155_new_n6740_), .Y(u2__abc_52155_new_n6741_));
INVX1 INVX1_1764 ( .A(u2__abc_52155_new_n6282_), .Y(u2__abc_52155_new_n6745_));
INVX1 INVX1_1765 ( .A(u2__abc_52155_new_n6250_), .Y(u2__abc_52155_new_n6746_));
INVX1 INVX1_1766 ( .A(u2__abc_52155_new_n6751_), .Y(u2__abc_52155_new_n6752_));
INVX1 INVX1_1767 ( .A(u2__abc_52155_new_n6266_), .Y(u2__abc_52155_new_n6755_));
INVX1 INVX1_1768 ( .A(u2__abc_52155_new_n6760_), .Y(u2__abc_52155_new_n6761_));
INVX1 INVX1_1769 ( .A(u2__abc_52155_new_n5837_), .Y(u2__abc_52155_new_n6770_));
INVX1 INVX1_177 ( .A(u2_o_449_), .Y(u2__abc_52155_new_n3007_));
INVX1 INVX1_1770 ( .A(u2__abc_52155_new_n5964_), .Y(u2__abc_52155_new_n6771_));
INVX1 INVX1_1771 ( .A(u2__abc_52155_new_n6027_), .Y(u2__abc_52155_new_n6772_));
INVX1 INVX1_1772 ( .A(u2__abc_52155_new_n6058_), .Y(u2__abc_52155_new_n6773_));
INVX1 INVX1_1773 ( .A(u2__abc_52155_new_n6088_), .Y(u2__abc_52155_new_n6774_));
INVX1 INVX1_1774 ( .A(u2__abc_52155_new_n6042_), .Y(u2__abc_52155_new_n6784_));
INVX1 INVX1_1775 ( .A(u2__abc_52155_new_n6026_), .Y(u2__abc_52155_new_n6791_));
INVX1 INVX1_1776 ( .A(u2__abc_52155_new_n5994_), .Y(u2__abc_52155_new_n6792_));
INVX1 INVX1_1777 ( .A(u2__abc_52155_new_n6797_), .Y(u2__abc_52155_new_n6798_));
INVX1 INVX1_1778 ( .A(u2__abc_52155_new_n6010_), .Y(u2__abc_52155_new_n6801_));
INVX1 INVX1_1779 ( .A(u2__abc_52155_new_n5899_), .Y(u2__abc_52155_new_n6811_));
INVX1 INVX1_178 ( .A(u2__abc_52155_new_n3008_), .Y(u2__abc_52155_new_n3009_));
INVX1 INVX1_1780 ( .A(u2__abc_52155_new_n5852_), .Y(u2__abc_52155_new_n6812_));
INVX1 INVX1_1781 ( .A(u2__abc_52155_new_n6817_), .Y(u2__abc_52155_new_n6818_));
INVX1 INVX1_1782 ( .A(u2__abc_52155_new_n5883_), .Y(u2__abc_52155_new_n6821_));
INVX1 INVX1_1783 ( .A(u2__abc_52155_new_n6826_), .Y(u2__abc_52155_new_n6827_));
INVX1 INVX1_1784 ( .A(u2__abc_52155_new_n5900_), .Y(u2__abc_52155_new_n6830_));
INVX1 INVX1_1785 ( .A(u2__abc_52155_new_n6832_), .Y(u2__abc_52155_new_n6833_));
INVX1 INVX1_1786 ( .A(u2__abc_52155_new_n5915_), .Y(u2__abc_52155_new_n6837_));
INVX1 INVX1_1787 ( .A(u2__abc_52155_new_n5946_), .Y(u2__abc_52155_new_n6844_));
INVX1 INVX1_1788 ( .A(u2__abc_52155_new_n5645_), .Y(u2__abc_52155_new_n6852_));
INVX1 INVX1_1789 ( .A(u2__abc_52155_new_n5706_), .Y(u2__abc_52155_new_n6855_));
INVX1 INVX1_179 ( .A(u2_remHi_448_), .Y(u2__abc_52155_new_n3011_));
INVX1 INVX1_1790 ( .A(u2__abc_52155_new_n5660_), .Y(u2__abc_52155_new_n6858_));
INVX1 INVX1_1791 ( .A(u2__abc_52155_new_n5709_), .Y(u2__abc_52155_new_n6870_));
INVX1 INVX1_1792 ( .A(u2__abc_52155_new_n5787_), .Y(u2__abc_52155_new_n6889_));
INVX1 INVX1_1793 ( .A(u2__abc_52155_new_n6899_), .Y(u2__abc_52155_new_n6900_));
INVX1 INVX1_1794 ( .A(u2__abc_52155_new_n5613_), .Y(u2__abc_52155_new_n6904_));
INVX1 INVX1_1795 ( .A(u2__abc_52155_new_n5643_), .Y(u2__abc_52155_new_n6907_));
INVX1 INVX1_1796 ( .A(u2__abc_52155_new_n5597_), .Y(u2__abc_52155_new_n6913_));
INVX1 INVX1_1797 ( .A(u2__abc_52155_new_n6918_), .Y(u2__abc_52155_new_n6919_));
INVX1 INVX1_1798 ( .A(u2_o_444_), .Y(u2__abc_52155_new_n6927_));
INVX1 INVX1_1799 ( .A(u2__abc_52155_new_n6928_), .Y(u2__abc_52155_new_n6929_));
INVX1 INVX1_18 ( .A(_abc_73687_new_n1553_), .Y(_abc_73687_new_n1568_));
INVX1 INVX1_180 ( .A(u2_o_448_), .Y(u2__abc_52155_new_n3013_));
INVX1 INVX1_1800 ( .A(u2_remHi_444_), .Y(u2__abc_52155_new_n6930_));
INVX1 INVX1_1801 ( .A(u2__abc_52155_new_n6931_), .Y(u2__abc_52155_new_n6932_));
INVX1 INVX1_1802 ( .A(u2_remHi_445_), .Y(u2__abc_52155_new_n6934_));
INVX1 INVX1_1803 ( .A(u2__abc_52155_new_n6935_), .Y(u2__abc_52155_new_n6936_));
INVX1 INVX1_1804 ( .A(u2_o_445_), .Y(u2__abc_52155_new_n6937_));
INVX1 INVX1_1805 ( .A(u2__abc_52155_new_n6938_), .Y(u2__abc_52155_new_n6939_));
INVX1 INVX1_1806 ( .A(u2_remHi_443_), .Y(u2__abc_52155_new_n6942_));
INVX1 INVX1_1807 ( .A(u2__abc_52155_new_n6943_), .Y(u2__abc_52155_new_n6944_));
INVX1 INVX1_1808 ( .A(u2_o_443_), .Y(u2__abc_52155_new_n6945_));
INVX1 INVX1_1809 ( .A(u2__abc_52155_new_n6946_), .Y(u2__abc_52155_new_n6947_));
INVX1 INVX1_181 ( .A(u2__abc_52155_new_n3015_), .Y(u2__abc_52155_new_n3016_));
INVX1 INVX1_1810 ( .A(u2_o_442_), .Y(u2__abc_52155_new_n6949_));
INVX1 INVX1_1811 ( .A(u2__abc_52155_new_n6950_), .Y(u2__abc_52155_new_n6951_));
INVX1 INVX1_1812 ( .A(u2_remHi_442_), .Y(u2__abc_52155_new_n6952_));
INVX1 INVX1_1813 ( .A(u2__abc_52155_new_n6953_), .Y(u2__abc_52155_new_n6954_));
INVX1 INVX1_1814 ( .A(u2_o_438_), .Y(u2__abc_52155_new_n6958_));
INVX1 INVX1_1815 ( .A(u2__abc_52155_new_n6959_), .Y(u2__abc_52155_new_n6960_));
INVX1 INVX1_1816 ( .A(u2_remHi_438_), .Y(u2__abc_52155_new_n6961_));
INVX1 INVX1_1817 ( .A(u2__abc_52155_new_n6962_), .Y(u2__abc_52155_new_n6963_));
INVX1 INVX1_1818 ( .A(u2_remHi_439_), .Y(u2__abc_52155_new_n6965_));
INVX1 INVX1_1819 ( .A(u2__abc_52155_new_n6966_), .Y(u2__abc_52155_new_n6967_));
INVX1 INVX1_182 ( .A(u2_o_447_), .Y(u2__abc_52155_new_n3018_));
INVX1 INVX1_1820 ( .A(u2_o_439_), .Y(u2__abc_52155_new_n6968_));
INVX1 INVX1_1821 ( .A(u2__abc_52155_new_n6969_), .Y(u2__abc_52155_new_n6970_));
INVX1 INVX1_1822 ( .A(u2_o_440_), .Y(u2__abc_52155_new_n6973_));
INVX1 INVX1_1823 ( .A(u2__abc_52155_new_n6974_), .Y(u2__abc_52155_new_n6975_));
INVX1 INVX1_1824 ( .A(u2_remHi_440_), .Y(u2__abc_52155_new_n6976_));
INVX1 INVX1_1825 ( .A(u2__abc_52155_new_n6977_), .Y(u2__abc_52155_new_n6978_));
INVX1 INVX1_1826 ( .A(u2_remHi_441_), .Y(u2__abc_52155_new_n6980_));
INVX1 INVX1_1827 ( .A(u2__abc_52155_new_n6981_), .Y(u2__abc_52155_new_n6982_));
INVX1 INVX1_1828 ( .A(u2_o_441_), .Y(u2__abc_52155_new_n6983_));
INVX1 INVX1_1829 ( .A(u2__abc_52155_new_n6984_), .Y(u2__abc_52155_new_n6985_));
INVX1 INVX1_183 ( .A(u2__abc_52155_new_n3019_), .Y(u2__abc_52155_new_n3020_));
INVX1 INVX1_1830 ( .A(u2_o_436_), .Y(u2__abc_52155_new_n6990_));
INVX1 INVX1_1831 ( .A(u2__abc_52155_new_n6991_), .Y(u2__abc_52155_new_n6992_));
INVX1 INVX1_1832 ( .A(u2_remHi_436_), .Y(u2__abc_52155_new_n6993_));
INVX1 INVX1_1833 ( .A(u2__abc_52155_new_n6994_), .Y(u2__abc_52155_new_n6995_));
INVX1 INVX1_1834 ( .A(u2_o_437_), .Y(u2__abc_52155_new_n6997_));
INVX1 INVX1_1835 ( .A(u2__abc_52155_new_n6998_), .Y(u2__abc_52155_new_n6999_));
INVX1 INVX1_1836 ( .A(u2_remHi_437_), .Y(u2__abc_52155_new_n7000_));
INVX1 INVX1_1837 ( .A(u2__abc_52155_new_n7001_), .Y(u2__abc_52155_new_n7002_));
INVX1 INVX1_1838 ( .A(u2_remHi_435_), .Y(u2__abc_52155_new_n7005_));
INVX1 INVX1_1839 ( .A(u2__abc_52155_new_n7006_), .Y(u2__abc_52155_new_n7007_));
INVX1 INVX1_184 ( .A(u2_remHi_447_), .Y(u2__abc_52155_new_n3021_));
INVX1 INVX1_1840 ( .A(u2_o_435_), .Y(u2__abc_52155_new_n7008_));
INVX1 INVX1_1841 ( .A(u2__abc_52155_new_n7009_), .Y(u2__abc_52155_new_n7010_));
INVX1 INVX1_1842 ( .A(u2_o_434_), .Y(u2__abc_52155_new_n7012_));
INVX1 INVX1_1843 ( .A(u2__abc_52155_new_n7013_), .Y(u2__abc_52155_new_n7014_));
INVX1 INVX1_1844 ( .A(u2_remHi_434_), .Y(u2__abc_52155_new_n7015_));
INVX1 INVX1_1845 ( .A(u2__abc_52155_new_n7016_), .Y(u2__abc_52155_new_n7017_));
INVX1 INVX1_1846 ( .A(u2_o_430_), .Y(u2__abc_52155_new_n7021_));
INVX1 INVX1_1847 ( .A(u2__abc_52155_new_n7022_), .Y(u2__abc_52155_new_n7023_));
INVX1 INVX1_1848 ( .A(u2_remHi_430_), .Y(u2__abc_52155_new_n7024_));
INVX1 INVX1_1849 ( .A(u2__abc_52155_new_n7025_), .Y(u2__abc_52155_new_n7026_));
INVX1 INVX1_185 ( .A(u2__abc_52155_new_n3022_), .Y(u2__abc_52155_new_n3023_));
INVX1 INVX1_1850 ( .A(u2_remHi_431_), .Y(u2__abc_52155_new_n7028_));
INVX1 INVX1_1851 ( .A(u2__abc_52155_new_n7029_), .Y(u2__abc_52155_new_n7030_));
INVX1 INVX1_1852 ( .A(u2_o_431_), .Y(u2__abc_52155_new_n7031_));
INVX1 INVX1_1853 ( .A(u2__abc_52155_new_n7032_), .Y(u2__abc_52155_new_n7033_));
INVX1 INVX1_1854 ( .A(u2_o_432_), .Y(u2__abc_52155_new_n7036_));
INVX1 INVX1_1855 ( .A(u2__abc_52155_new_n7037_), .Y(u2__abc_52155_new_n7038_));
INVX1 INVX1_1856 ( .A(u2_remHi_432_), .Y(u2__abc_52155_new_n7039_));
INVX1 INVX1_1857 ( .A(u2__abc_52155_new_n7040_), .Y(u2__abc_52155_new_n7041_));
INVX1 INVX1_1858 ( .A(u2_remHi_433_), .Y(u2__abc_52155_new_n7043_));
INVX1 INVX1_1859 ( .A(u2__abc_52155_new_n7044_), .Y(u2__abc_52155_new_n7045_));
INVX1 INVX1_186 ( .A(u2_o_446_), .Y(u2__abc_52155_new_n3025_));
INVX1 INVX1_1860 ( .A(u2_o_433_), .Y(u2__abc_52155_new_n7046_));
INVX1 INVX1_1861 ( .A(u2__abc_52155_new_n7047_), .Y(u2__abc_52155_new_n7048_));
INVX1 INVX1_1862 ( .A(u2_o_424_), .Y(u2__abc_52155_new_n7054_));
INVX1 INVX1_1863 ( .A(u2__abc_52155_new_n7055_), .Y(u2__abc_52155_new_n7056_));
INVX1 INVX1_1864 ( .A(u2_remHi_424_), .Y(u2__abc_52155_new_n7057_));
INVX1 INVX1_1865 ( .A(u2__abc_52155_new_n7058_), .Y(u2__abc_52155_new_n7059_));
INVX1 INVX1_1866 ( .A(u2_remHi_425_), .Y(u2__abc_52155_new_n7061_));
INVX1 INVX1_1867 ( .A(u2__abc_52155_new_n7062_), .Y(u2__abc_52155_new_n7063_));
INVX1 INVX1_1868 ( .A(u2_o_425_), .Y(u2__abc_52155_new_n7064_));
INVX1 INVX1_1869 ( .A(u2__abc_52155_new_n7065_), .Y(u2__abc_52155_new_n7066_));
INVX1 INVX1_187 ( .A(u2__abc_52155_new_n3026_), .Y(u2__abc_52155_new_n3027_));
INVX1 INVX1_1870 ( .A(u2_o_422_), .Y(u2__abc_52155_new_n7069_));
INVX1 INVX1_1871 ( .A(u2__abc_52155_new_n7070_), .Y(u2__abc_52155_new_n7071_));
INVX1 INVX1_1872 ( .A(u2_remHi_422_), .Y(u2__abc_52155_new_n7072_));
INVX1 INVX1_1873 ( .A(u2__abc_52155_new_n7073_), .Y(u2__abc_52155_new_n7074_));
INVX1 INVX1_1874 ( .A(u2_remHi_423_), .Y(u2__abc_52155_new_n7076_));
INVX1 INVX1_1875 ( .A(u2__abc_52155_new_n7077_), .Y(u2__abc_52155_new_n7078_));
INVX1 INVX1_1876 ( .A(u2_o_423_), .Y(u2__abc_52155_new_n7079_));
INVX1 INVX1_1877 ( .A(u2__abc_52155_new_n7080_), .Y(u2__abc_52155_new_n7081_));
INVX1 INVX1_1878 ( .A(u2_o_428_), .Y(u2__abc_52155_new_n7085_));
INVX1 INVX1_1879 ( .A(u2__abc_52155_new_n7086_), .Y(u2__abc_52155_new_n7087_));
INVX1 INVX1_188 ( .A(u2_remHi_446_), .Y(u2__abc_52155_new_n3028_));
INVX1 INVX1_1880 ( .A(u2_remHi_428_), .Y(u2__abc_52155_new_n7088_));
INVX1 INVX1_1881 ( .A(u2__abc_52155_new_n7089_), .Y(u2__abc_52155_new_n7090_));
INVX1 INVX1_1882 ( .A(u2_o_429_), .Y(u2__abc_52155_new_n7092_));
INVX1 INVX1_1883 ( .A(u2__abc_52155_new_n7093_), .Y(u2__abc_52155_new_n7094_));
INVX1 INVX1_1884 ( .A(u2_remHi_429_), .Y(u2__abc_52155_new_n7095_));
INVX1 INVX1_1885 ( .A(u2__abc_52155_new_n7096_), .Y(u2__abc_52155_new_n7097_));
INVX1 INVX1_1886 ( .A(u2_remHi_427_), .Y(u2__abc_52155_new_n7100_));
INVX1 INVX1_1887 ( .A(u2__abc_52155_new_n7101_), .Y(u2__abc_52155_new_n7102_));
INVX1 INVX1_1888 ( .A(u2_o_427_), .Y(u2__abc_52155_new_n7103_));
INVX1 INVX1_1889 ( .A(u2__abc_52155_new_n7104_), .Y(u2__abc_52155_new_n7105_));
INVX1 INVX1_189 ( .A(u2__abc_52155_new_n3029_), .Y(u2__abc_52155_new_n3030_));
INVX1 INVX1_1890 ( .A(u2_o_426_), .Y(u2__abc_52155_new_n7107_));
INVX1 INVX1_1891 ( .A(u2__abc_52155_new_n7108_), .Y(u2__abc_52155_new_n7109_));
INVX1 INVX1_1892 ( .A(u2_remHi_426_), .Y(u2__abc_52155_new_n7110_));
INVX1 INVX1_1893 ( .A(u2__abc_52155_new_n7111_), .Y(u2__abc_52155_new_n7112_));
INVX1 INVX1_1894 ( .A(u2_o_420_), .Y(u2__abc_52155_new_n7117_));
INVX1 INVX1_1895 ( .A(u2__abc_52155_new_n7118_), .Y(u2__abc_52155_new_n7119_));
INVX1 INVX1_1896 ( .A(u2_remHi_420_), .Y(u2__abc_52155_new_n7120_));
INVX1 INVX1_1897 ( .A(u2__abc_52155_new_n7121_), .Y(u2__abc_52155_new_n7122_));
INVX1 INVX1_1898 ( .A(u2_o_421_), .Y(u2__abc_52155_new_n7124_));
INVX1 INVX1_1899 ( .A(u2__abc_52155_new_n7125_), .Y(u2__abc_52155_new_n7126_));
INVX1 INVX1_19 ( .A(_abc_73687_new_n1566_), .Y(_abc_73687_new_n1569_));
INVX1 INVX1_190 ( .A(u2__abc_52155_new_n3033_), .Y(u2__abc_52155_new_n3034_));
INVX1 INVX1_1900 ( .A(u2_remHi_421_), .Y(u2__abc_52155_new_n7127_));
INVX1 INVX1_1901 ( .A(u2__abc_52155_new_n7128_), .Y(u2__abc_52155_new_n7129_));
INVX1 INVX1_1902 ( .A(u2_remHi_419_), .Y(u2__abc_52155_new_n7132_));
INVX1 INVX1_1903 ( .A(u2__abc_52155_new_n7133_), .Y(u2__abc_52155_new_n7134_));
INVX1 INVX1_1904 ( .A(u2_o_419_), .Y(u2__abc_52155_new_n7135_));
INVX1 INVX1_1905 ( .A(u2__abc_52155_new_n7136_), .Y(u2__abc_52155_new_n7137_));
INVX1 INVX1_1906 ( .A(u2_o_418_), .Y(u2__abc_52155_new_n7139_));
INVX1 INVX1_1907 ( .A(u2__abc_52155_new_n7140_), .Y(u2__abc_52155_new_n7141_));
INVX1 INVX1_1908 ( .A(u2_remHi_418_), .Y(u2__abc_52155_new_n7142_));
INVX1 INVX1_1909 ( .A(u2__abc_52155_new_n7143_), .Y(u2__abc_52155_new_n7144_));
INVX1 INVX1_191 ( .A(sqrto_12_), .Y(u2__abc_52155_new_n3035_));
INVX1 INVX1_1910 ( .A(u2_o_416_), .Y(u2__abc_52155_new_n7148_));
INVX1 INVX1_1911 ( .A(u2__abc_52155_new_n7149_), .Y(u2__abc_52155_new_n7150_));
INVX1 INVX1_1912 ( .A(u2_remHi_416_), .Y(u2__abc_52155_new_n7151_));
INVX1 INVX1_1913 ( .A(u2__abc_52155_new_n7152_), .Y(u2__abc_52155_new_n7153_));
INVX1 INVX1_1914 ( .A(u2_remHi_417_), .Y(u2__abc_52155_new_n7155_));
INVX1 INVX1_1915 ( .A(u2__abc_52155_new_n7156_), .Y(u2__abc_52155_new_n7157_));
INVX1 INVX1_1916 ( .A(u2_o_417_), .Y(u2__abc_52155_new_n7158_));
INVX1 INVX1_1917 ( .A(u2__abc_52155_new_n7159_), .Y(u2__abc_52155_new_n7160_));
INVX1 INVX1_1918 ( .A(u2_remHi_415_), .Y(u2__abc_52155_new_n7163_));
INVX1 INVX1_1919 ( .A(u2__abc_52155_new_n7164_), .Y(u2__abc_52155_new_n7165_));
INVX1 INVX1_192 ( .A(u2_remHi_12_), .Y(u2__abc_52155_new_n3037_));
INVX1 INVX1_1920 ( .A(u2_o_415_), .Y(u2__abc_52155_new_n7166_));
INVX1 INVX1_1921 ( .A(u2__abc_52155_new_n7167_), .Y(u2__abc_52155_new_n7168_));
INVX1 INVX1_1922 ( .A(u2_o_414_), .Y(u2__abc_52155_new_n7170_));
INVX1 INVX1_1923 ( .A(u2__abc_52155_new_n7171_), .Y(u2__abc_52155_new_n7172_));
INVX1 INVX1_1924 ( .A(u2_remHi_414_), .Y(u2__abc_52155_new_n7173_));
INVX1 INVX1_1925 ( .A(u2__abc_52155_new_n7174_), .Y(u2__abc_52155_new_n7175_));
INVX1 INVX1_1926 ( .A(u2_o_388_), .Y(u2__abc_52155_new_n7182_));
INVX1 INVX1_1927 ( .A(u2__abc_52155_new_n7183_), .Y(u2__abc_52155_new_n7184_));
INVX1 INVX1_1928 ( .A(u2_remHi_388_), .Y(u2__abc_52155_new_n7185_));
INVX1 INVX1_1929 ( .A(u2__abc_52155_new_n7186_), .Y(u2__abc_52155_new_n7187_));
INVX1 INVX1_193 ( .A(u2__abc_52155_new_n3039_), .Y(u2__abc_52155_new_n3040_));
INVX1 INVX1_1930 ( .A(u2_o_389_), .Y(u2__abc_52155_new_n7189_));
INVX1 INVX1_1931 ( .A(u2__abc_52155_new_n7190_), .Y(u2__abc_52155_new_n7191_));
INVX1 INVX1_1932 ( .A(u2_remHi_389_), .Y(u2__abc_52155_new_n7192_));
INVX1 INVX1_1933 ( .A(u2__abc_52155_new_n7193_), .Y(u2__abc_52155_new_n7194_));
INVX1 INVX1_1934 ( .A(u2_remHi_387_), .Y(u2__abc_52155_new_n7197_));
INVX1 INVX1_1935 ( .A(u2__abc_52155_new_n7198_), .Y(u2__abc_52155_new_n7199_));
INVX1 INVX1_1936 ( .A(u2_o_387_), .Y(u2__abc_52155_new_n7200_));
INVX1 INVX1_1937 ( .A(u2__abc_52155_new_n7201_), .Y(u2__abc_52155_new_n7202_));
INVX1 INVX1_1938 ( .A(u2_o_386_), .Y(u2__abc_52155_new_n7204_));
INVX1 INVX1_1939 ( .A(u2__abc_52155_new_n7205_), .Y(u2__abc_52155_new_n7206_));
INVX1 INVX1_194 ( .A(u2_remHi_13_), .Y(u2__abc_52155_new_n3041_));
INVX1 INVX1_1940 ( .A(u2_remHi_386_), .Y(u2__abc_52155_new_n7207_));
INVX1 INVX1_1941 ( .A(u2__abc_52155_new_n7208_), .Y(u2__abc_52155_new_n7209_));
INVX1 INVX1_1942 ( .A(u2_o_384_), .Y(u2__abc_52155_new_n7213_));
INVX1 INVX1_1943 ( .A(u2__abc_52155_new_n7214_), .Y(u2__abc_52155_new_n7215_));
INVX1 INVX1_1944 ( .A(u2_remHi_384_), .Y(u2__abc_52155_new_n7216_));
INVX1 INVX1_1945 ( .A(u2__abc_52155_new_n7217_), .Y(u2__abc_52155_new_n7218_));
INVX1 INVX1_1946 ( .A(u2_remHi_385_), .Y(u2__abc_52155_new_n7220_));
INVX1 INVX1_1947 ( .A(u2__abc_52155_new_n7221_), .Y(u2__abc_52155_new_n7222_));
INVX1 INVX1_1948 ( .A(u2_o_385_), .Y(u2__abc_52155_new_n7223_));
INVX1 INVX1_1949 ( .A(u2__abc_52155_new_n7224_), .Y(u2__abc_52155_new_n7225_));
INVX1 INVX1_195 ( .A(sqrto_13_), .Y(u2__abc_52155_new_n3043_));
INVX1 INVX1_1950 ( .A(u2_remHi_383_), .Y(u2__abc_52155_new_n7228_));
INVX1 INVX1_1951 ( .A(u2__abc_52155_new_n7229_), .Y(u2__abc_52155_new_n7230_));
INVX1 INVX1_1952 ( .A(u2_o_383_), .Y(u2__abc_52155_new_n7231_));
INVX1 INVX1_1953 ( .A(u2__abc_52155_new_n7232_), .Y(u2__abc_52155_new_n7233_));
INVX1 INVX1_1954 ( .A(u2_o_382_), .Y(u2__abc_52155_new_n7235_));
INVX1 INVX1_1955 ( .A(u2__abc_52155_new_n7236_), .Y(u2__abc_52155_new_n7237_));
INVX1 INVX1_1956 ( .A(u2_remHi_382_), .Y(u2__abc_52155_new_n7238_));
INVX1 INVX1_1957 ( .A(u2__abc_52155_new_n7239_), .Y(u2__abc_52155_new_n7240_));
INVX1 INVX1_1958 ( .A(u2_o_408_), .Y(u2__abc_52155_new_n7245_));
INVX1 INVX1_1959 ( .A(u2__abc_52155_new_n7246_), .Y(u2__abc_52155_new_n7247_));
INVX1 INVX1_196 ( .A(u2__abc_52155_new_n3045_), .Y(u2__abc_52155_new_n3046_));
INVX1 INVX1_1960 ( .A(u2_remHi_408_), .Y(u2__abc_52155_new_n7248_));
INVX1 INVX1_1961 ( .A(u2__abc_52155_new_n7249_), .Y(u2__abc_52155_new_n7250_));
INVX1 INVX1_1962 ( .A(u2_remHi_409_), .Y(u2__abc_52155_new_n7252_));
INVX1 INVX1_1963 ( .A(u2__abc_52155_new_n7253_), .Y(u2__abc_52155_new_n7254_));
INVX1 INVX1_1964 ( .A(u2_o_409_), .Y(u2__abc_52155_new_n7255_));
INVX1 INVX1_1965 ( .A(u2__abc_52155_new_n7256_), .Y(u2__abc_52155_new_n7257_));
INVX1 INVX1_1966 ( .A(u2_remHi_407_), .Y(u2__abc_52155_new_n7260_));
INVX1 INVX1_1967 ( .A(u2__abc_52155_new_n7261_), .Y(u2__abc_52155_new_n7262_));
INVX1 INVX1_1968 ( .A(u2_o_407_), .Y(u2__abc_52155_new_n7263_));
INVX1 INVX1_1969 ( .A(u2__abc_52155_new_n7264_), .Y(u2__abc_52155_new_n7265_));
INVX1 INVX1_197 ( .A(sqrto_11_), .Y(u2__abc_52155_new_n3048_));
INVX1 INVX1_1970 ( .A(u2_o_406_), .Y(u2__abc_52155_new_n7267_));
INVX1 INVX1_1971 ( .A(u2__abc_52155_new_n7268_), .Y(u2__abc_52155_new_n7269_));
INVX1 INVX1_1972 ( .A(u2_remHi_406_), .Y(u2__abc_52155_new_n7270_));
INVX1 INVX1_1973 ( .A(u2__abc_52155_new_n7271_), .Y(u2__abc_52155_new_n7272_));
INVX1 INVX1_1974 ( .A(u2_o_412_), .Y(u2__abc_52155_new_n7276_));
INVX1 INVX1_1975 ( .A(u2__abc_52155_new_n7277_), .Y(u2__abc_52155_new_n7278_));
INVX1 INVX1_1976 ( .A(u2_remHi_412_), .Y(u2__abc_52155_new_n7279_));
INVX1 INVX1_1977 ( .A(u2__abc_52155_new_n7280_), .Y(u2__abc_52155_new_n7281_));
INVX1 INVX1_1978 ( .A(u2_o_413_), .Y(u2__abc_52155_new_n7283_));
INVX1 INVX1_1979 ( .A(u2__abc_52155_new_n7284_), .Y(u2__abc_52155_new_n7285_));
INVX1 INVX1_198 ( .A(u2__abc_52155_new_n3049_), .Y(u2__abc_52155_new_n3050_));
INVX1 INVX1_1980 ( .A(u2_remHi_413_), .Y(u2__abc_52155_new_n7286_));
INVX1 INVX1_1981 ( .A(u2__abc_52155_new_n7287_), .Y(u2__abc_52155_new_n7288_));
INVX1 INVX1_1982 ( .A(u2_remHi_411_), .Y(u2__abc_52155_new_n7291_));
INVX1 INVX1_1983 ( .A(u2__abc_52155_new_n7292_), .Y(u2__abc_52155_new_n7293_));
INVX1 INVX1_1984 ( .A(u2_o_411_), .Y(u2__abc_52155_new_n7294_));
INVX1 INVX1_1985 ( .A(u2__abc_52155_new_n7295_), .Y(u2__abc_52155_new_n7296_));
INVX1 INVX1_1986 ( .A(u2_o_410_), .Y(u2__abc_52155_new_n7298_));
INVX1 INVX1_1987 ( .A(u2__abc_52155_new_n7299_), .Y(u2__abc_52155_new_n7300_));
INVX1 INVX1_1988 ( .A(u2_remHi_410_), .Y(u2__abc_52155_new_n7301_));
INVX1 INVX1_1989 ( .A(u2__abc_52155_new_n7302_), .Y(u2__abc_52155_new_n7303_));
INVX1 INVX1_199 ( .A(u2_remHi_11_), .Y(u2__abc_52155_new_n3051_));
INVX1 INVX1_1990 ( .A(u2_o_398_), .Y(u2__abc_52155_new_n7308_));
INVX1 INVX1_1991 ( .A(u2__abc_52155_new_n7309_), .Y(u2__abc_52155_new_n7310_));
INVX1 INVX1_1992 ( .A(u2_remHi_398_), .Y(u2__abc_52155_new_n7311_));
INVX1 INVX1_1993 ( .A(u2__abc_52155_new_n7312_), .Y(u2__abc_52155_new_n7313_));
INVX1 INVX1_1994 ( .A(u2_remHi_399_), .Y(u2__abc_52155_new_n7315_));
INVX1 INVX1_1995 ( .A(u2__abc_52155_new_n7316_), .Y(u2__abc_52155_new_n7317_));
INVX1 INVX1_1996 ( .A(u2_o_399_), .Y(u2__abc_52155_new_n7318_));
INVX1 INVX1_1997 ( .A(u2__abc_52155_new_n7319_), .Y(u2__abc_52155_new_n7320_));
INVX1 INVX1_1998 ( .A(u2_o_400_), .Y(u2__abc_52155_new_n7323_));
INVX1 INVX1_1999 ( .A(u2__abc_52155_new_n7324_), .Y(u2__abc_52155_new_n7325_));
INVX1 INVX1_2 ( .A(\a[112] ), .Y(_abc_73687_new_n1170_));
INVX1 INVX1_20 ( .A(_abc_73687_new_n1567_), .Y(_abc_73687_new_n1574_));
INVX1 INVX1_200 ( .A(u2__abc_52155_new_n3052_), .Y(u2__abc_52155_new_n3053_));
INVX1 INVX1_2000 ( .A(u2_remHi_400_), .Y(u2__abc_52155_new_n7326_));
INVX1 INVX1_2001 ( .A(u2__abc_52155_new_n7327_), .Y(u2__abc_52155_new_n7328_));
INVX1 INVX1_2002 ( .A(u2_remHi_401_), .Y(u2__abc_52155_new_n7330_));
INVX1 INVX1_2003 ( .A(u2__abc_52155_new_n7331_), .Y(u2__abc_52155_new_n7332_));
INVX1 INVX1_2004 ( .A(u2_o_401_), .Y(u2__abc_52155_new_n7333_));
INVX1 INVX1_2005 ( .A(u2__abc_52155_new_n7334_), .Y(u2__abc_52155_new_n7335_));
INVX1 INVX1_2006 ( .A(u2_o_404_), .Y(u2__abc_52155_new_n7339_));
INVX1 INVX1_2007 ( .A(u2__abc_52155_new_n7340_), .Y(u2__abc_52155_new_n7341_));
INVX1 INVX1_2008 ( .A(u2_remHi_404_), .Y(u2__abc_52155_new_n7342_));
INVX1 INVX1_2009 ( .A(u2__abc_52155_new_n7343_), .Y(u2__abc_52155_new_n7344_));
INVX1 INVX1_201 ( .A(sqrto_10_), .Y(u2__abc_52155_new_n3055_));
INVX1 INVX1_2010 ( .A(u2_o_405_), .Y(u2__abc_52155_new_n7346_));
INVX1 INVX1_2011 ( .A(u2__abc_52155_new_n7347_), .Y(u2__abc_52155_new_n7348_));
INVX1 INVX1_2012 ( .A(u2_remHi_405_), .Y(u2__abc_52155_new_n7349_));
INVX1 INVX1_2013 ( .A(u2__abc_52155_new_n7350_), .Y(u2__abc_52155_new_n7351_));
INVX1 INVX1_2014 ( .A(u2_remHi_403_), .Y(u2__abc_52155_new_n7354_));
INVX1 INVX1_2015 ( .A(u2__abc_52155_new_n7355_), .Y(u2__abc_52155_new_n7356_));
INVX1 INVX1_2016 ( .A(u2_o_403_), .Y(u2__abc_52155_new_n7357_));
INVX1 INVX1_2017 ( .A(u2__abc_52155_new_n7358_), .Y(u2__abc_52155_new_n7359_));
INVX1 INVX1_2018 ( .A(u2_o_402_), .Y(u2__abc_52155_new_n7361_));
INVX1 INVX1_2019 ( .A(u2__abc_52155_new_n7362_), .Y(u2__abc_52155_new_n7363_));
INVX1 INVX1_202 ( .A(u2_remHi_10_), .Y(u2__abc_52155_new_n3057_));
INVX1 INVX1_2020 ( .A(u2_remHi_402_), .Y(u2__abc_52155_new_n7364_));
INVX1 INVX1_2021 ( .A(u2__abc_52155_new_n7365_), .Y(u2__abc_52155_new_n7366_));
INVX1 INVX1_2022 ( .A(u2_o_392_), .Y(u2__abc_52155_new_n7372_));
INVX1 INVX1_2023 ( .A(u2__abc_52155_new_n7373_), .Y(u2__abc_52155_new_n7374_));
INVX1 INVX1_2024 ( .A(u2_remHi_392_), .Y(u2__abc_52155_new_n7375_));
INVX1 INVX1_2025 ( .A(u2__abc_52155_new_n7376_), .Y(u2__abc_52155_new_n7377_));
INVX1 INVX1_2026 ( .A(u2_remHi_393_), .Y(u2__abc_52155_new_n7379_));
INVX1 INVX1_2027 ( .A(u2__abc_52155_new_n7380_), .Y(u2__abc_52155_new_n7381_));
INVX1 INVX1_2028 ( .A(u2_o_393_), .Y(u2__abc_52155_new_n7382_));
INVX1 INVX1_2029 ( .A(u2__abc_52155_new_n7383_), .Y(u2__abc_52155_new_n7384_));
INVX1 INVX1_203 ( .A(u2__abc_52155_new_n3059_), .Y(u2__abc_52155_new_n3060_));
INVX1 INVX1_2030 ( .A(u2_o_390_), .Y(u2__abc_52155_new_n7387_));
INVX1 INVX1_2031 ( .A(u2__abc_52155_new_n7388_), .Y(u2__abc_52155_new_n7389_));
INVX1 INVX1_2032 ( .A(u2_remHi_390_), .Y(u2__abc_52155_new_n7390_));
INVX1 INVX1_2033 ( .A(u2__abc_52155_new_n7391_), .Y(u2__abc_52155_new_n7392_));
INVX1 INVX1_2034 ( .A(u2_remHi_391_), .Y(u2__abc_52155_new_n7394_));
INVX1 INVX1_2035 ( .A(u2__abc_52155_new_n7395_), .Y(u2__abc_52155_new_n7396_));
INVX1 INVX1_2036 ( .A(u2_o_391_), .Y(u2__abc_52155_new_n7397_));
INVX1 INVX1_2037 ( .A(u2__abc_52155_new_n7398_), .Y(u2__abc_52155_new_n7399_));
INVX1 INVX1_2038 ( .A(u2_o_396_), .Y(u2__abc_52155_new_n7403_));
INVX1 INVX1_2039 ( .A(u2__abc_52155_new_n7404_), .Y(u2__abc_52155_new_n7405_));
INVX1 INVX1_204 ( .A(sqrto_8_), .Y(u2__abc_52155_new_n3063_));
INVX1 INVX1_2040 ( .A(u2_remHi_396_), .Y(u2__abc_52155_new_n7406_));
INVX1 INVX1_2041 ( .A(u2__abc_52155_new_n7407_), .Y(u2__abc_52155_new_n7408_));
INVX1 INVX1_2042 ( .A(u2_o_397_), .Y(u2__abc_52155_new_n7410_));
INVX1 INVX1_2043 ( .A(u2__abc_52155_new_n7411_), .Y(u2__abc_52155_new_n7412_));
INVX1 INVX1_2044 ( .A(u2_remHi_397_), .Y(u2__abc_52155_new_n7413_));
INVX1 INVX1_2045 ( .A(u2__abc_52155_new_n7414_), .Y(u2__abc_52155_new_n7415_));
INVX1 INVX1_2046 ( .A(u2_remHi_395_), .Y(u2__abc_52155_new_n7418_));
INVX1 INVX1_2047 ( .A(u2__abc_52155_new_n7419_), .Y(u2__abc_52155_new_n7420_));
INVX1 INVX1_2048 ( .A(u2_o_395_), .Y(u2__abc_52155_new_n7421_));
INVX1 INVX1_2049 ( .A(u2__abc_52155_new_n7422_), .Y(u2__abc_52155_new_n7423_));
INVX1 INVX1_205 ( .A(u2_remHi_8_), .Y(u2__abc_52155_new_n3065_));
INVX1 INVX1_2050 ( .A(u2_o_394_), .Y(u2__abc_52155_new_n7425_));
INVX1 INVX1_2051 ( .A(u2__abc_52155_new_n7426_), .Y(u2__abc_52155_new_n7427_));
INVX1 INVX1_2052 ( .A(u2_remHi_394_), .Y(u2__abc_52155_new_n7428_));
INVX1 INVX1_2053 ( .A(u2__abc_52155_new_n7429_), .Y(u2__abc_52155_new_n7430_));
INVX1 INVX1_2054 ( .A(u2__abc_52155_new_n7437_), .Y(u2__abc_52155_new_n7438_));
INVX1 INVX1_2055 ( .A(u2__abc_52155_new_n7565_), .Y(u2__abc_52155_new_n7566_));
INVX1 INVX1_2056 ( .A(u2__abc_52155_new_n7570_), .Y(u2__abc_52155_new_n7571_));
INVX1 INVX1_2057 ( .A(u2__abc_52155_new_n7575_), .Y(u2__abc_52155_new_n7576_));
INVX1 INVX1_2058 ( .A(u2__abc_52155_new_n3124_), .Y(u2__abc_52155_new_n7583_));
INVX1 INVX1_2059 ( .A(u2__abc_52155_new_n3126_), .Y(u2__abc_52155_new_n7584_));
INVX1 INVX1_206 ( .A(u2__abc_52155_new_n3067_), .Y(u2__abc_52155_new_n3068_));
INVX1 INVX1_2060 ( .A(u2__abc_52155_new_n3113_), .Y(u2__abc_52155_new_n7590_));
INVX1 INVX1_2061 ( .A(u2__abc_52155_new_n7622_), .Y(u2__abc_52155_new_n7623_));
INVX1 INVX1_2062 ( .A(u2_remHiShift_0_), .Y(u2__abc_52155_new_n7625_));
INVX1 INVX1_2063 ( .A(u2__abc_52155_new_n7629_), .Y(u2__abc_52155_new_n7630_));
INVX1 INVX1_2064 ( .A(u2__abc_52155_new_n7587_), .Y(u2__abc_52155_new_n7636_));
INVX1 INVX1_2065 ( .A(u2__abc_52155_new_n7643_), .Y(u2__abc_52155_new_n7644_));
INVX1 INVX1_2066 ( .A(u2__abc_52155_new_n3118_), .Y(u2__abc_52155_new_n7650_));
INVX1 INVX1_2067 ( .A(u2__abc_52155_new_n7651_), .Y(u2__abc_52155_new_n7652_));
INVX1 INVX1_2068 ( .A(u2__abc_52155_new_n7653_), .Y(u2__abc_52155_new_n7654_));
INVX1 INVX1_2069 ( .A(u2__abc_52155_new_n7661_), .Y(u2__abc_52155_new_n7662_));
INVX1 INVX1_207 ( .A(sqrto_9_), .Y(u2__abc_52155_new_n3069_));
INVX1 INVX1_2070 ( .A(u2__abc_52155_new_n3123_), .Y(u2__abc_52155_new_n7668_));
INVX1 INVX1_2071 ( .A(u2__abc_52155_new_n7673_), .Y(u2__abc_52155_new_n7674_));
INVX1 INVX1_2072 ( .A(u2__abc_52155_new_n7680_), .Y(u2__abc_52155_new_n7681_));
INVX1 INVX1_2073 ( .A(u2__abc_52155_new_n3111_), .Y(u2__abc_52155_new_n7687_));
INVX1 INVX1_2074 ( .A(u2__abc_52155_new_n7690_), .Y(u2__abc_52155_new_n7691_));
INVX1 INVX1_2075 ( .A(u2__abc_52155_new_n7697_), .Y(u2__abc_52155_new_n7698_));
INVX1 INVX1_2076 ( .A(u2__abc_52155_new_n3106_), .Y(u2__abc_52155_new_n7704_));
INVX1 INVX1_2077 ( .A(u2__abc_52155_new_n3108_), .Y(u2__abc_52155_new_n7705_));
INVX1 INVX1_2078 ( .A(u2__abc_52155_new_n7706_), .Y(u2__abc_52155_new_n7707_));
INVX1 INVX1_2079 ( .A(u2__abc_52155_new_n7715_), .Y(u2__abc_52155_new_n7716_));
INVX1 INVX1_208 ( .A(u2__abc_52155_new_n3070_), .Y(u2__abc_52155_new_n3071_));
INVX1 INVX1_2080 ( .A(u2__abc_52155_new_n3095_), .Y(u2__abc_52155_new_n7722_));
INVX1 INVX1_2081 ( .A(u2__abc_52155_new_n7728_), .Y(u2__abc_52155_new_n7729_));
INVX1 INVX1_2082 ( .A(u2__abc_52155_new_n7735_), .Y(u2__abc_52155_new_n7736_));
INVX1 INVX1_2083 ( .A(u2__abc_52155_new_n3100_), .Y(u2__abc_52155_new_n7742_));
INVX1 INVX1_2084 ( .A(u2__abc_52155_new_n3092_), .Y(u2__abc_52155_new_n7743_));
INVX1 INVX1_2085 ( .A(u2__abc_52155_new_n7744_), .Y(u2__abc_52155_new_n7745_));
INVX1 INVX1_2086 ( .A(u2_remHi_7_), .Y(u2__abc_52155_new_n7753_));
INVX1 INVX1_2087 ( .A(u2__abc_52155_new_n7754_), .Y(u2__abc_52155_new_n7755_));
INVX1 INVX1_2088 ( .A(u2__abc_52155_new_n3101_), .Y(u2__abc_52155_new_n7762_));
INVX1 INVX1_2089 ( .A(u2__abc_52155_new_n7768_), .Y(u2__abc_52155_new_n7769_));
INVX1 INVX1_209 ( .A(u2_remHi_9_), .Y(u2__abc_52155_new_n3072_));
INVX1 INVX1_2090 ( .A(u2__abc_52155_new_n7776_), .Y(u2__abc_52155_new_n7777_));
INVX1 INVX1_2091 ( .A(u2__abc_52155_new_n3081_), .Y(u2__abc_52155_new_n7783_));
INVX1 INVX1_2092 ( .A(u2__abc_52155_new_n7784_), .Y(u2__abc_52155_new_n7785_));
INVX1 INVX1_2093 ( .A(u2__abc_52155_new_n7793_), .Y(u2__abc_52155_new_n7794_));
INVX1 INVX1_2094 ( .A(u2__abc_52155_new_n7800_), .Y(u2__abc_52155_new_n7801_));
INVX1 INVX1_2095 ( .A(u2__abc_52155_new_n7806_), .Y(u2__abc_52155_new_n7807_));
INVX1 INVX1_2096 ( .A(u2__abc_52155_new_n7813_), .Y(u2__abc_52155_new_n7814_));
INVX1 INVX1_2097 ( .A(u2__abc_52155_new_n3075_), .Y(u2__abc_52155_new_n7820_));
INVX1 INVX1_2098 ( .A(u2__abc_52155_new_n3064_), .Y(u2__abc_52155_new_n7821_));
INVX1 INVX1_2099 ( .A(u2__abc_52155_new_n7822_), .Y(u2__abc_52155_new_n7823_));
INVX1 INVX1_21 ( .A(\a[119] ), .Y(_abc_73687_new_n1575_));
INVX1 INVX1_210 ( .A(u2__abc_52155_new_n3073_), .Y(u2__abc_52155_new_n3074_));
INVX1 INVX1_2100 ( .A(u2__abc_52155_new_n7831_), .Y(u2__abc_52155_new_n7832_));
INVX1 INVX1_2101 ( .A(u2__abc_52155_new_n7840_), .Y(u2__abc_52155_new_n7841_));
INVX1 INVX1_2102 ( .A(u2__abc_52155_new_n7843_), .Y(u2__abc_52155_new_n7844_));
INVX1 INVX1_2103 ( .A(u2__abc_52155_new_n7850_), .Y(u2__abc_52155_new_n7851_));
INVX1 INVX1_2104 ( .A(u2__abc_52155_new_n3056_), .Y(u2__abc_52155_new_n7857_));
INVX1 INVX1_2105 ( .A(u2__abc_52155_new_n3054_), .Y(u2__abc_52155_new_n7860_));
INVX1 INVX1_2106 ( .A(u2__abc_52155_new_n7858_), .Y(u2__abc_52155_new_n7861_));
INVX1 INVX1_2107 ( .A(u2__abc_52155_new_n7868_), .Y(u2__abc_52155_new_n7869_));
INVX1 INVX1_2108 ( .A(u2__abc_52155_new_n3061_), .Y(u2__abc_52155_new_n7875_));
INVX1 INVX1_2109 ( .A(u2__abc_52155_new_n7878_), .Y(u2__abc_52155_new_n7879_));
INVX1 INVX1_211 ( .A(sqrto_7_), .Y(u2__abc_52155_new_n3077_));
INVX1 INVX1_2110 ( .A(u2__abc_52155_new_n7880_), .Y(u2__abc_52155_new_n7881_));
INVX1 INVX1_2111 ( .A(u2__abc_52155_new_n7883_), .Y(u2__abc_52155_new_n7884_));
INVX1 INVX1_2112 ( .A(u2_remHi_14_), .Y(u2__abc_52155_new_n7890_));
INVX1 INVX1_2113 ( .A(u2__abc_52155_new_n7891_), .Y(u2__abc_52155_new_n7892_));
INVX1 INVX1_2114 ( .A(u2__abc_52155_new_n3036_), .Y(u2__abc_52155_new_n7898_));
INVX1 INVX1_2115 ( .A(u2__abc_52155_new_n7899_), .Y(u2__abc_52155_new_n7900_));
INVX1 INVX1_2116 ( .A(u2__abc_52155_new_n7908_), .Y(u2__abc_52155_new_n7909_));
INVX1 INVX1_2117 ( .A(u2__abc_52155_new_n7915_), .Y(u2__abc_52155_new_n7916_));
INVX1 INVX1_2118 ( .A(u2__abc_52155_new_n7918_), .Y(u2__abc_52155_new_n7919_));
INVX1 INVX1_2119 ( .A(u2__abc_52155_new_n7925_), .Y(u2__abc_52155_new_n7926_));
INVX1 INVX1_212 ( .A(u2__abc_52155_new_n3078_), .Y(u2__abc_52155_new_n3079_));
INVX1 INVX1_2120 ( .A(u2__abc_52155_new_n7928_), .Y(u2__abc_52155_new_n7929_));
INVX1 INVX1_2121 ( .A(u2__abc_52155_new_n7931_), .Y(u2__abc_52155_new_n7932_));
INVX1 INVX1_2122 ( .A(u2__abc_52155_new_n7938_), .Y(u2__abc_52155_new_n7939_));
INVX1 INVX1_2123 ( .A(u2__abc_52155_new_n3250_), .Y(u2__abc_52155_new_n7945_));
INVX1 INVX1_2124 ( .A(u2__abc_52155_new_n7946_), .Y(u2__abc_52155_new_n7947_));
INVX1 INVX1_2125 ( .A(u2__abc_52155_new_n7955_), .Y(u2__abc_52155_new_n7956_));
INVX1 INVX1_2126 ( .A(u2__abc_52155_new_n3231_), .Y(u2__abc_52155_new_n7962_));
INVX1 INVX1_2127 ( .A(u2__abc_52155_new_n7966_), .Y(u2__abc_52155_new_n7967_));
INVX1 INVX1_2128 ( .A(u2__abc_52155_new_n7973_), .Y(u2__abc_52155_new_n7974_));
INVX1 INVX1_2129 ( .A(u2__abc_52155_new_n3228_), .Y(u2__abc_52155_new_n7980_));
INVX1 INVX1_213 ( .A(u2_remHi_6_), .Y(u2__abc_52155_new_n3082_));
INVX1 INVX1_2130 ( .A(u2__abc_52155_new_n7981_), .Y(u2__abc_52155_new_n7982_));
INVX1 INVX1_2131 ( .A(u2__abc_52155_new_n3236_), .Y(u2__abc_52155_new_n7984_));
INVX1 INVX1_2132 ( .A(u2__abc_52155_new_n7991_), .Y(u2__abc_52155_new_n7992_));
INVX1 INVX1_2133 ( .A(u2__abc_52155_new_n3273_), .Y(u2__abc_52155_new_n7998_));
INVX1 INVX1_2134 ( .A(u2__abc_52155_new_n8003_), .Y(u2__abc_52155_new_n8004_));
INVX1 INVX1_2135 ( .A(u2__abc_52155_new_n8005_), .Y(u2__abc_52155_new_n8006_));
INVX1 INVX1_2136 ( .A(u2__abc_52155_new_n8010_), .Y(u2__abc_52155_new_n8011_));
INVX1 INVX1_2137 ( .A(u2__abc_52155_new_n8017_), .Y(u2__abc_52155_new_n8018_));
INVX1 INVX1_2138 ( .A(u2__abc_52155_new_n3268_), .Y(u2__abc_52155_new_n8024_));
INVX1 INVX1_2139 ( .A(u2__abc_52155_new_n3270_), .Y(u2__abc_52155_new_n8025_));
INVX1 INVX1_214 ( .A(sqrto_6_), .Y(u2__abc_52155_new_n3084_));
INVX1 INVX1_2140 ( .A(u2__abc_52155_new_n8026_), .Y(u2__abc_52155_new_n8027_));
INVX1 INVX1_2141 ( .A(u2__abc_52155_new_n8035_), .Y(u2__abc_52155_new_n8036_));
INVX1 INVX1_2142 ( .A(u2__abc_52155_new_n3257_), .Y(u2__abc_52155_new_n8043_));
INVX1 INVX1_2143 ( .A(u2__abc_52155_new_n8044_), .Y(u2__abc_52155_new_n8045_));
INVX1 INVX1_2144 ( .A(u2__abc_52155_new_n8047_), .Y(u2__abc_52155_new_n8048_));
INVX1 INVX1_2145 ( .A(u2__abc_52155_new_n8050_), .Y(u2__abc_52155_new_n8051_));
INVX1 INVX1_2146 ( .A(u2__abc_52155_new_n8056_), .Y(u2__abc_52155_new_n8057_));
INVX1 INVX1_2147 ( .A(u2__abc_52155_new_n3254_), .Y(u2__abc_52155_new_n8064_));
INVX1 INVX1_2148 ( .A(u2__abc_52155_new_n8065_), .Y(u2__abc_52155_new_n8066_));
INVX1 INVX1_2149 ( .A(u2__abc_52155_new_n3262_), .Y(u2__abc_52155_new_n8068_));
INVX1 INVX1_215 ( .A(u2__abc_52155_new_n3089_), .Y(u2__abc_52155_new_n3090_));
INVX1 INVX1_2150 ( .A(u2__abc_52155_new_n8074_), .Y(u2__abc_52155_new_n8075_));
INVX1 INVX1_2151 ( .A(u2__abc_52155_new_n8081_), .Y(u2__abc_52155_new_n8082_));
INVX1 INVX1_2152 ( .A(u2__abc_52155_new_n8083_), .Y(u2__abc_52155_new_n8084_));
INVX1 INVX1_2153 ( .A(u2__abc_52155_new_n8091_), .Y(u2__abc_52155_new_n8092_));
INVX1 INVX1_2154 ( .A(u2__abc_52155_new_n8094_), .Y(u2__abc_52155_new_n8095_));
INVX1 INVX1_2155 ( .A(u2__abc_52155_new_n8101_), .Y(u2__abc_52155_new_n8102_));
INVX1 INVX1_2156 ( .A(u2__abc_52155_new_n8109_), .Y(u2__abc_52155_new_n8110_));
INVX1 INVX1_2157 ( .A(u2__abc_52155_new_n3185_), .Y(u2__abc_52155_new_n8112_));
INVX1 INVX1_2158 ( .A(u2__abc_52155_new_n8118_), .Y(u2__abc_52155_new_n8119_));
INVX1 INVX1_2159 ( .A(u2__abc_52155_new_n3171_), .Y(u2__abc_52155_new_n8126_));
INVX1 INVX1_216 ( .A(sqrto_4_), .Y(u2__abc_52155_new_n3091_));
INVX1 INVX1_2160 ( .A(u2__abc_52155_new_n8129_), .Y(u2__abc_52155_new_n8130_));
INVX1 INVX1_2161 ( .A(u2__abc_52155_new_n8132_), .Y(u2__abc_52155_new_n8133_));
INVX1 INVX1_2162 ( .A(u2__abc_52155_new_n8138_), .Y(u2__abc_52155_new_n8139_));
INVX1 INVX1_2163 ( .A(u2__abc_52155_new_n3168_), .Y(u2__abc_52155_new_n8145_));
INVX1 INVX1_2164 ( .A(u2__abc_52155_new_n8146_), .Y(u2__abc_52155_new_n8147_));
INVX1 INVX1_2165 ( .A(u2__abc_52155_new_n3176_), .Y(u2__abc_52155_new_n8149_));
INVX1 INVX1_2166 ( .A(u2__abc_52155_new_n8156_), .Y(u2__abc_52155_new_n8157_));
INVX1 INVX1_2167 ( .A(u2__abc_52155_new_n8164_), .Y(u2__abc_52155_new_n8165_));
INVX1 INVX1_2168 ( .A(u2__abc_52155_new_n8171_), .Y(u2__abc_52155_new_n8172_));
INVX1 INVX1_2169 ( .A(u2__abc_52155_new_n8174_), .Y(u2__abc_52155_new_n8175_));
INVX1 INVX1_217 ( .A(u2_remHi_4_), .Y(u2__abc_52155_new_n3093_));
INVX1 INVX1_2170 ( .A(u2__abc_52155_new_n8180_), .Y(u2__abc_52155_new_n8181_));
INVX1 INVX1_2171 ( .A(u2__abc_52155_new_n3216_), .Y(u2__abc_52155_new_n8188_));
INVX1 INVX1_2172 ( .A(u2__abc_52155_new_n8189_), .Y(u2__abc_52155_new_n8190_));
INVX1 INVX1_2173 ( .A(u2__abc_52155_new_n8197_), .Y(u2__abc_52155_new_n8198_));
INVX1 INVX1_2174 ( .A(u2__abc_52155_new_n8206_), .Y(u2__abc_52155_new_n8207_));
INVX1 INVX1_2175 ( .A(u2__abc_52155_new_n8209_), .Y(u2__abc_52155_new_n8210_));
INVX1 INVX1_2176 ( .A(u2_remHi_30_), .Y(u2__abc_52155_new_n8216_));
INVX1 INVX1_2177 ( .A(u2__abc_52155_new_n8217_), .Y(u2__abc_52155_new_n8218_));
INVX1 INVX1_2178 ( .A(u2__abc_52155_new_n8224_), .Y(u2__abc_52155_new_n8225_));
INVX1 INVX1_2179 ( .A(u2__abc_52155_new_n3208_), .Y(u2__abc_52155_new_n8227_));
INVX1 INVX1_218 ( .A(u2_remHi_5_), .Y(u2__abc_52155_new_n3096_));
INVX1 INVX1_2180 ( .A(u2__abc_52155_new_n8234_), .Y(u2__abc_52155_new_n8235_));
INVX1 INVX1_2181 ( .A(u2__abc_52155_new_n8241_), .Y(u2__abc_52155_new_n8242_));
INVX1 INVX1_2182 ( .A(u2__abc_52155_new_n8249_), .Y(u2__abc_52155_new_n8250_));
INVX1 INVX1_2183 ( .A(u2__abc_52155_new_n8257_), .Y(u2__abc_52155_new_n8258_));
INVX1 INVX1_2184 ( .A(u2__abc_52155_new_n3530_), .Y(u2__abc_52155_new_n8264_));
INVX1 INVX1_2185 ( .A(u2__abc_52155_new_n8265_), .Y(u2__abc_52155_new_n8267_));
INVX1 INVX1_2186 ( .A(u2__abc_52155_new_n8274_), .Y(u2__abc_52155_new_n8275_));
INVX1 INVX1_2187 ( .A(u2__abc_52155_new_n3511_), .Y(u2__abc_52155_new_n8282_));
INVX1 INVX1_2188 ( .A(u2__abc_52155_new_n8286_), .Y(u2__abc_52155_new_n8287_));
INVX1 INVX1_2189 ( .A(u2__abc_52155_new_n8292_), .Y(u2__abc_52155_new_n8293_));
INVX1 INVX1_219 ( .A(sqrto_5_), .Y(u2__abc_52155_new_n3098_));
INVX1 INVX1_2190 ( .A(u2__abc_52155_new_n3516_), .Y(u2__abc_52155_new_n8299_));
INVX1 INVX1_2191 ( .A(u2__abc_52155_new_n3508_), .Y(u2__abc_52155_new_n8300_));
INVX1 INVX1_2192 ( .A(u2__abc_52155_new_n8301_), .Y(u2__abc_52155_new_n8303_));
INVX1 INVX1_2193 ( .A(u2__abc_52155_new_n8310_), .Y(u2__abc_52155_new_n8311_));
INVX1 INVX1_2194 ( .A(u2__abc_52155_new_n3553_), .Y(u2__abc_52155_new_n8317_));
INVX1 INVX1_2195 ( .A(u2__abc_52155_new_n8322_), .Y(u2__abc_52155_new_n8323_));
INVX1 INVX1_2196 ( .A(u2__abc_52155_new_n8324_), .Y(u2__abc_52155_new_n8325_));
INVX1 INVX1_2197 ( .A(u2__abc_52155_new_n8329_), .Y(u2__abc_52155_new_n8330_));
INVX1 INVX1_2198 ( .A(u2__abc_52155_new_n8336_), .Y(u2__abc_52155_new_n8337_));
INVX1 INVX1_2199 ( .A(u2__abc_52155_new_n3548_), .Y(u2__abc_52155_new_n8343_));
INVX1 INVX1_22 ( .A(_abc_73687_new_n1562_), .Y(_abc_73687_new_n1576_));
INVX1 INVX1_220 ( .A(sqrto_3_), .Y(u2__abc_52155_new_n3102_));
INVX1 INVX1_2200 ( .A(u2__abc_52155_new_n3550_), .Y(u2__abc_52155_new_n8344_));
INVX1 INVX1_2201 ( .A(u2__abc_52155_new_n8345_), .Y(u2__abc_52155_new_n8346_));
INVX1 INVX1_2202 ( .A(u2__abc_52155_new_n8354_), .Y(u2__abc_52155_new_n8355_));
INVX1 INVX1_2203 ( .A(u2__abc_52155_new_n3537_), .Y(u2__abc_52155_new_n8362_));
INVX1 INVX1_2204 ( .A(u2__abc_52155_new_n8363_), .Y(u2__abc_52155_new_n8364_));
INVX1 INVX1_2205 ( .A(u2__abc_52155_new_n8366_), .Y(u2__abc_52155_new_n8367_));
INVX1 INVX1_2206 ( .A(u2__abc_52155_new_n8369_), .Y(u2__abc_52155_new_n8370_));
INVX1 INVX1_2207 ( .A(u2__abc_52155_new_n8375_), .Y(u2__abc_52155_new_n8376_));
INVX1 INVX1_2208 ( .A(u2__abc_52155_new_n3534_), .Y(u2__abc_52155_new_n8382_));
INVX1 INVX1_2209 ( .A(u2__abc_52155_new_n3542_), .Y(u2__abc_52155_new_n8385_));
INVX1 INVX1_221 ( .A(u2_remHi_3_), .Y(u2__abc_52155_new_n3104_));
INVX1 INVX1_2210 ( .A(u2__abc_52155_new_n8383_), .Y(u2__abc_52155_new_n8386_));
INVX1 INVX1_2211 ( .A(u2__abc_52155_new_n8393_), .Y(u2__abc_52155_new_n8394_));
INVX1 INVX1_2212 ( .A(u2__abc_52155_new_n8400_), .Y(u2__abc_52155_new_n8401_));
INVX1 INVX1_2213 ( .A(u2__abc_52155_new_n8407_), .Y(u2__abc_52155_new_n8408_));
INVX1 INVX1_2214 ( .A(u2__abc_52155_new_n8412_), .Y(u2__abc_52155_new_n8413_));
INVX1 INVX1_2215 ( .A(u2__abc_52155_new_n8419_), .Y(u2__abc_52155_new_n8420_));
INVX1 INVX1_2216 ( .A(u2__abc_52155_new_n3472_), .Y(u2__abc_52155_new_n8426_));
INVX1 INVX1_2217 ( .A(u2__abc_52155_new_n8427_), .Y(u2__abc_52155_new_n8428_));
INVX1 INVX1_2218 ( .A(u2__abc_52155_new_n8436_), .Y(u2__abc_52155_new_n8437_));
INVX1 INVX1_2219 ( .A(u2__abc_52155_new_n3451_), .Y(u2__abc_52155_new_n8443_));
INVX1 INVX1_222 ( .A(sqrto_2_), .Y(u2__abc_52155_new_n3107_));
INVX1 INVX1_2220 ( .A(u2__abc_52155_new_n8447_), .Y(u2__abc_52155_new_n8448_));
INVX1 INVX1_2221 ( .A(u2__abc_52155_new_n8454_), .Y(u2__abc_52155_new_n8455_));
INVX1 INVX1_2222 ( .A(u2__abc_52155_new_n3448_), .Y(u2__abc_52155_new_n8461_));
INVX1 INVX1_2223 ( .A(u2__abc_52155_new_n3456_), .Y(u2__abc_52155_new_n8464_));
INVX1 INVX1_2224 ( .A(u2__abc_52155_new_n8462_), .Y(u2__abc_52155_new_n8465_));
INVX1 INVX1_2225 ( .A(u2__abc_52155_new_n8472_), .Y(u2__abc_52155_new_n8473_));
INVX1 INVX1_2226 ( .A(u2__abc_52155_new_n8485_), .Y(u2__abc_52155_new_n8486_));
INVX1 INVX1_2227 ( .A(u2__abc_52155_new_n8490_), .Y(u2__abc_52155_new_n8491_));
INVX1 INVX1_2228 ( .A(u2__abc_52155_new_n8496_), .Y(u2__abc_52155_new_n8497_));
INVX1 INVX1_2229 ( .A(u2__abc_52155_new_n3496_), .Y(u2__abc_52155_new_n8505_));
INVX1 INVX1_223 ( .A(u2_remHi_2_), .Y(u2__abc_52155_new_n3109_));
INVX1 INVX1_2230 ( .A(u2__abc_52155_new_n8503_), .Y(u2__abc_52155_new_n8506_));
INVX1 INVX1_2231 ( .A(u2__abc_52155_new_n8513_), .Y(u2__abc_52155_new_n8514_));
INVX1 INVX1_2232 ( .A(u2__abc_52155_new_n8522_), .Y(u2__abc_52155_new_n8523_));
INVX1 INVX1_2233 ( .A(u2__abc_52155_new_n8524_), .Y(u2__abc_52155_new_n8525_));
INVX1 INVX1_2234 ( .A(u2__abc_52155_new_n8532_), .Y(u2__abc_52155_new_n8533_));
INVX1 INVX1_2235 ( .A(u2__abc_52155_new_n3488_), .Y(u2__abc_52155_new_n8539_));
INVX1 INVX1_2236 ( .A(u2__abc_52155_new_n8540_), .Y(u2__abc_52155_new_n8542_));
INVX1 INVX1_2237 ( .A(u2__abc_52155_new_n8549_), .Y(u2__abc_52155_new_n8550_));
INVX1 INVX1_2238 ( .A(u2__abc_52155_new_n8559_), .Y(u2__abc_52155_new_n8560_));
INVX1 INVX1_2239 ( .A(u2__abc_52155_new_n8569_), .Y(u2__abc_52155_new_n8570_));
INVX1 INVX1_224 ( .A(sqrto_0_), .Y(u2__abc_52155_new_n3114_));
INVX1 INVX1_2240 ( .A(u2__abc_52155_new_n8576_), .Y(u2__abc_52155_new_n8577_));
INVX1 INVX1_2241 ( .A(u2__abc_52155_new_n8583_), .Y(u2__abc_52155_new_n8584_));
INVX1 INVX1_2242 ( .A(u2__abc_52155_new_n3404_), .Y(u2__abc_52155_new_n8586_));
INVX1 INVX1_2243 ( .A(u2__abc_52155_new_n8593_), .Y(u2__abc_52155_new_n8594_));
INVX1 INVX1_2244 ( .A(u2__abc_52155_new_n3390_), .Y(u2__abc_52155_new_n8601_));
INVX1 INVX1_2245 ( .A(u2__abc_52155_new_n8604_), .Y(u2__abc_52155_new_n8605_));
INVX1 INVX1_2246 ( .A(u2__abc_52155_new_n8607_), .Y(u2__abc_52155_new_n8608_));
INVX1 INVX1_2247 ( .A(u2__abc_52155_new_n8613_), .Y(u2__abc_52155_new_n8614_));
INVX1 INVX1_2248 ( .A(u2__abc_52155_new_n3387_), .Y(u2__abc_52155_new_n8620_));
INVX1 INVX1_2249 ( .A(u2__abc_52155_new_n3395_), .Y(u2__abc_52155_new_n8623_));
INVX1 INVX1_225 ( .A(u2_remHi_0_), .Y(u2__abc_52155_new_n3116_));
INVX1 INVX1_2250 ( .A(u2__abc_52155_new_n8621_), .Y(u2__abc_52155_new_n8624_));
INVX1 INVX1_2251 ( .A(u2__abc_52155_new_n8631_), .Y(u2__abc_52155_new_n8632_));
INVX1 INVX1_2252 ( .A(u2__abc_52155_new_n8643_), .Y(u2__abc_52155_new_n8644_));
INVX1 INVX1_2253 ( .A(u2__abc_52155_new_n8648_), .Y(u2__abc_52155_new_n8649_));
INVX1 INVX1_2254 ( .A(u2__abc_52155_new_n8654_), .Y(u2__abc_52155_new_n8655_));
INVX1 INVX1_2255 ( .A(u2__abc_52155_new_n3435_), .Y(u2__abc_52155_new_n8663_));
INVX1 INVX1_2256 ( .A(u2__abc_52155_new_n8661_), .Y(u2__abc_52155_new_n8664_));
INVX1 INVX1_2257 ( .A(u2__abc_52155_new_n8671_), .Y(u2__abc_52155_new_n8672_));
INVX1 INVX1_2258 ( .A(u2__abc_52155_new_n8680_), .Y(u2__abc_52155_new_n8681_));
INVX1 INVX1_2259 ( .A(u2__abc_52155_new_n8682_), .Y(u2__abc_52155_new_n8683_));
INVX1 INVX1_226 ( .A(u2_remHi_1_), .Y(u2__abc_52155_new_n3119_));
INVX1 INVX1_2260 ( .A(u2__abc_52155_new_n8690_), .Y(u2__abc_52155_new_n8691_));
INVX1 INVX1_2261 ( .A(u2__abc_52155_new_n3427_), .Y(u2__abc_52155_new_n8697_));
INVX1 INVX1_2262 ( .A(u2__abc_52155_new_n8698_), .Y(u2__abc_52155_new_n8700_));
INVX1 INVX1_2263 ( .A(u2__abc_52155_new_n8707_), .Y(u2__abc_52155_new_n8708_));
INVX1 INVX1_2264 ( .A(u2__abc_52155_new_n8716_), .Y(u2__abc_52155_new_n8717_));
INVX1 INVX1_2265 ( .A(u2__abc_52155_new_n8726_), .Y(u2__abc_52155_new_n8727_));
INVX1 INVX1_2266 ( .A(u2__abc_52155_new_n8732_), .Y(u2__abc_52155_new_n8733_));
INVX1 INVX1_2267 ( .A(u2__abc_52155_new_n3351_), .Y(u2__abc_52155_new_n8741_));
INVX1 INVX1_2268 ( .A(u2__abc_52155_new_n8742_), .Y(u2__abc_52155_new_n8744_));
INVX1 INVX1_2269 ( .A(u2__abc_52155_new_n8749_), .Y(u2__abc_52155_new_n8750_));
INVX1 INVX1_227 ( .A(sqrto_1_), .Y(u2__abc_52155_new_n3121_));
INVX1 INVX1_2270 ( .A(u2__abc_52155_new_n8757_), .Y(u2__abc_52155_new_n8758_));
INVX1 INVX1_2271 ( .A(u2__abc_52155_new_n8761_), .Y(u2__abc_52155_new_n8762_));
INVX1 INVX1_2272 ( .A(u2__abc_52155_new_n8769_), .Y(u2__abc_52155_new_n8770_));
INVX1 INVX1_2273 ( .A(u2__abc_52155_new_n3336_), .Y(u2__abc_52155_new_n8776_));
INVX1 INVX1_2274 ( .A(u2__abc_52155_new_n8777_), .Y(u2__abc_52155_new_n8779_));
INVX1 INVX1_2275 ( .A(u2__abc_52155_new_n8786_), .Y(u2__abc_52155_new_n8787_));
INVX1 INVX1_2276 ( .A(u2__abc_52155_new_n8799_), .Y(u2__abc_52155_new_n8800_));
INVX1 INVX1_2277 ( .A(u2__abc_52155_new_n8807_), .Y(u2__abc_52155_new_n8808_));
INVX1 INVX1_2278 ( .A(u2__abc_52155_new_n8814_), .Y(u2__abc_52155_new_n8815_));
INVX1 INVX1_2279 ( .A(u2__abc_52155_new_n8817_), .Y(u2__abc_52155_new_n8818_));
INVX1 INVX1_228 ( .A(u2_root_0_), .Y(u2__abc_52155_new_n3125_));
INVX1 INVX1_2280 ( .A(u2__abc_52155_new_n8824_), .Y(u2__abc_52155_new_n8825_));
INVX1 INVX1_2281 ( .A(u2__abc_52155_new_n8831_), .Y(u2__abc_52155_new_n8832_));
INVX1 INVX1_2282 ( .A(u2__abc_52155_new_n8833_), .Y(u2__abc_52155_new_n8834_));
INVX1 INVX1_2283 ( .A(u2_remHi_62_), .Y(u2__abc_52155_new_n8841_));
INVX1 INVX1_2284 ( .A(u2__abc_52155_new_n8842_), .Y(u2__abc_52155_new_n8843_));
INVX1 INVX1_2285 ( .A(u2__abc_52155_new_n3367_), .Y(u2__abc_52155_new_n8849_));
INVX1 INVX1_2286 ( .A(u2__abc_52155_new_n8850_), .Y(u2__abc_52155_new_n8852_));
INVX1 INVX1_2287 ( .A(u2__abc_52155_new_n8859_), .Y(u2__abc_52155_new_n8860_));
INVX1 INVX1_2288 ( .A(u2__abc_52155_new_n8880_), .Y(u2__abc_52155_new_n8881_));
INVX1 INVX1_2289 ( .A(u2__abc_52155_new_n8886_), .Y(u2__abc_52155_new_n8887_));
INVX1 INVX1_229 ( .A(u2__abc_52155_new_n3120_), .Y(u2__abc_52155_new_n3128_));
INVX1 INVX1_2290 ( .A(u2__abc_52155_new_n8893_), .Y(u2__abc_52155_new_n8894_));
INVX1 INVX1_2291 ( .A(u2__abc_52155_new_n4090_), .Y(u2__abc_52155_new_n8896_));
INVX1 INVX1_2292 ( .A(u2__abc_52155_new_n8903_), .Y(u2__abc_52155_new_n8904_));
INVX1 INVX1_2293 ( .A(u2__abc_52155_new_n4096_), .Y(u2__abc_52155_new_n8910_));
INVX1 INVX1_2294 ( .A(u2__abc_52155_new_n8912_), .Y(u2__abc_52155_new_n8913_));
INVX1 INVX1_2295 ( .A(u2__abc_52155_new_n8917_), .Y(u2__abc_52155_new_n8918_));
INVX1 INVX1_2296 ( .A(u2__abc_52155_new_n8924_), .Y(u2__abc_52155_new_n8925_));
INVX1 INVX1_2297 ( .A(u2__abc_52155_new_n4093_), .Y(u2__abc_52155_new_n8931_));
INVX1 INVX1_2298 ( .A(u2__abc_52155_new_n4101_), .Y(u2__abc_52155_new_n8934_));
INVX1 INVX1_2299 ( .A(u2__abc_52155_new_n8932_), .Y(u2__abc_52155_new_n8935_));
INVX1 INVX1_23 ( .A(_abc_73687_new_n1579_), .Y(_abc_73687_new_n1580_));
INVX1 INVX1_230 ( .A(u2__abc_52155_new_n3117_), .Y(u2__abc_52155_new_n3129_));
INVX1 INVX1_2300 ( .A(u2__abc_52155_new_n8942_), .Y(u2__abc_52155_new_n8943_));
INVX1 INVX1_2301 ( .A(u2__abc_52155_new_n4125_), .Y(u2__abc_52155_new_n8949_));
INVX1 INVX1_2302 ( .A(u2__abc_52155_new_n8957_), .Y(u2__abc_52155_new_n8958_));
INVX1 INVX1_2303 ( .A(u2__abc_52155_new_n8964_), .Y(u2__abc_52155_new_n8965_));
INVX1 INVX1_2304 ( .A(u2__abc_52155_new_n4120_), .Y(u2__abc_52155_new_n8971_));
INVX1 INVX1_2305 ( .A(u2__abc_52155_new_n4122_), .Y(u2__abc_52155_new_n8972_));
INVX1 INVX1_2306 ( .A(u2__abc_52155_new_n8973_), .Y(u2__abc_52155_new_n8974_));
INVX1 INVX1_2307 ( .A(u2__abc_52155_new_n8975_), .Y(u2__abc_52155_new_n8976_));
INVX1 INVX1_2308 ( .A(u2__abc_52155_new_n8983_), .Y(u2__abc_52155_new_n8984_));
INVX1 INVX1_2309 ( .A(u2__abc_52155_new_n4109_), .Y(u2__abc_52155_new_n8990_));
INVX1 INVX1_231 ( .A(u2__abc_52155_new_n3105_), .Y(u2__abc_52155_new_n3134_));
INVX1 INVX1_2310 ( .A(u2__abc_52155_new_n8992_), .Y(u2__abc_52155_new_n8993_));
INVX1 INVX1_2311 ( .A(u2__abc_52155_new_n9000_), .Y(u2__abc_52155_new_n9001_));
INVX1 INVX1_2312 ( .A(u2__abc_52155_new_n4106_), .Y(u2__abc_52155_new_n9007_));
INVX1 INVX1_2313 ( .A(u2__abc_52155_new_n4114_), .Y(u2__abc_52155_new_n9010_));
INVX1 INVX1_2314 ( .A(u2__abc_52155_new_n9008_), .Y(u2__abc_52155_new_n9011_));
INVX1 INVX1_2315 ( .A(u2__abc_52155_new_n9018_), .Y(u2__abc_52155_new_n9019_));
INVX1 INVX1_2316 ( .A(u2__abc_52155_new_n9025_), .Y(u2__abc_52155_new_n9026_));
INVX1 INVX1_2317 ( .A(u2__abc_52155_new_n4115_), .Y(u2__abc_52155_new_n9027_));
INVX1 INVX1_2318 ( .A(u2__abc_52155_new_n9030_), .Y(u2__abc_52155_new_n9031_));
INVX1 INVX1_2319 ( .A(u2__abc_52155_new_n9035_), .Y(u2__abc_52155_new_n9036_));
INVX1 INVX1_232 ( .A(u2__abc_52155_new_n3110_), .Y(u2__abc_52155_new_n3135_));
INVX1 INVX1_2320 ( .A(u2__abc_52155_new_n9040_), .Y(u2__abc_52155_new_n9041_));
INVX1 INVX1_2321 ( .A(u2__abc_52155_new_n9047_), .Y(u2__abc_52155_new_n9048_));
INVX1 INVX1_2322 ( .A(u2__abc_52155_new_n4032_), .Y(u2__abc_52155_new_n9054_));
INVX1 INVX1_2323 ( .A(u2__abc_52155_new_n9055_), .Y(u2__abc_52155_new_n9057_));
INVX1 INVX1_2324 ( .A(u2__abc_52155_new_n9064_), .Y(u2__abc_52155_new_n9065_));
INVX1 INVX1_2325 ( .A(u2__abc_52155_new_n4038_), .Y(u2__abc_52155_new_n9071_));
INVX1 INVX1_2326 ( .A(u2__abc_52155_new_n9073_), .Y(u2__abc_52155_new_n9074_));
INVX1 INVX1_2327 ( .A(u2__abc_52155_new_n9077_), .Y(u2__abc_52155_new_n9078_));
INVX1 INVX1_2328 ( .A(u2__abc_52155_new_n9085_), .Y(u2__abc_52155_new_n9086_));
INVX1 INVX1_2329 ( .A(u2__abc_52155_new_n4035_), .Y(u2__abc_52155_new_n9092_));
INVX1 INVX1_233 ( .A(u2__abc_52155_new_n3097_), .Y(u2__abc_52155_new_n3139_));
INVX1 INVX1_2330 ( .A(u2__abc_52155_new_n4043_), .Y(u2__abc_52155_new_n9095_));
INVX1 INVX1_2331 ( .A(u2__abc_52155_new_n9093_), .Y(u2__abc_52155_new_n9096_));
INVX1 INVX1_2332 ( .A(u2__abc_52155_new_n9103_), .Y(u2__abc_52155_new_n9104_));
INVX1 INVX1_2333 ( .A(u2__abc_52155_new_n9110_), .Y(u2__abc_52155_new_n9111_));
INVX1 INVX1_2334 ( .A(u2__abc_52155_new_n9114_), .Y(u2__abc_52155_new_n9115_));
INVX1 INVX1_2335 ( .A(u2__abc_52155_new_n9118_), .Y(u2__abc_52155_new_n9119_));
INVX1 INVX1_2336 ( .A(u2__abc_52155_new_n9126_), .Y(u2__abc_52155_new_n9127_));
INVX1 INVX1_2337 ( .A(u2__abc_52155_new_n9133_), .Y(u2__abc_52155_new_n9134_));
INVX1 INVX1_2338 ( .A(u2__abc_52155_new_n9135_), .Y(u2__abc_52155_new_n9136_));
INVX1 INVX1_2339 ( .A(u2__abc_52155_new_n9143_), .Y(u2__abc_52155_new_n9144_));
INVX1 INVX1_234 ( .A(u2__abc_52155_new_n3094_), .Y(u2__abc_52155_new_n3140_));
INVX1 INVX1_2340 ( .A(u2__abc_52155_new_n9150_), .Y(u2__abc_52155_new_n9151_));
INVX1 INVX1_2341 ( .A(u2__abc_52155_new_n9152_), .Y(u2__abc_52155_new_n9153_));
INVX1 INVX1_2342 ( .A(u2__abc_52155_new_n9160_), .Y(u2__abc_52155_new_n9161_));
INVX1 INVX1_2343 ( .A(u2__abc_52155_new_n4060_), .Y(u2__abc_52155_new_n9167_));
INVX1 INVX1_2344 ( .A(u2__abc_52155_new_n9168_), .Y(u2__abc_52155_new_n9170_));
INVX1 INVX1_2345 ( .A(u2__abc_52155_new_n9177_), .Y(u2__abc_52155_new_n9178_));
INVX1 INVX1_2346 ( .A(u2__abc_52155_new_n9197_), .Y(u2__abc_52155_new_n9198_));
INVX1 INVX1_2347 ( .A(u2__abc_52155_new_n9204_), .Y(u2__abc_52155_new_n9205_));
INVX1 INVX1_2348 ( .A(u2__abc_52155_new_n3971_), .Y(u2__abc_52155_new_n9211_));
INVX1 INVX1_2349 ( .A(u2__abc_52155_new_n9212_), .Y(u2__abc_52155_new_n9214_));
INVX1 INVX1_235 ( .A(u2__abc_52155_new_n3062_), .Y(u2__abc_52155_new_n3146_));
INVX1 INVX1_2350 ( .A(u2__abc_52155_new_n9221_), .Y(u2__abc_52155_new_n9222_));
INVX1 INVX1_2351 ( .A(u2__abc_52155_new_n3977_), .Y(u2__abc_52155_new_n9228_));
INVX1 INVX1_2352 ( .A(u2__abc_52155_new_n9230_), .Y(u2__abc_52155_new_n9231_));
INVX1 INVX1_2353 ( .A(u2__abc_52155_new_n9234_), .Y(u2__abc_52155_new_n9235_));
INVX1 INVX1_2354 ( .A(u2__abc_52155_new_n9242_), .Y(u2__abc_52155_new_n9243_));
INVX1 INVX1_2355 ( .A(u2__abc_52155_new_n3974_), .Y(u2__abc_52155_new_n9249_));
INVX1 INVX1_2356 ( .A(u2__abc_52155_new_n3982_), .Y(u2__abc_52155_new_n9252_));
INVX1 INVX1_2357 ( .A(u2__abc_52155_new_n9250_), .Y(u2__abc_52155_new_n9253_));
INVX1 INVX1_2358 ( .A(u2__abc_52155_new_n9260_), .Y(u2__abc_52155_new_n9261_));
INVX1 INVX1_2359 ( .A(u2__abc_52155_new_n9267_), .Y(u2__abc_52155_new_n9268_));
INVX1 INVX1_236 ( .A(u2__abc_52155_new_n3076_), .Y(u2__abc_52155_new_n3147_));
INVX1 INVX1_2360 ( .A(u2__abc_52155_new_n9271_), .Y(u2__abc_52155_new_n9272_));
INVX1 INVX1_2361 ( .A(u2__abc_52155_new_n9275_), .Y(u2__abc_52155_new_n9276_));
INVX1 INVX1_2362 ( .A(u2__abc_52155_new_n9283_), .Y(u2__abc_52155_new_n9284_));
INVX1 INVX1_2363 ( .A(u2__abc_52155_new_n4007_), .Y(u2__abc_52155_new_n9292_));
INVX1 INVX1_2364 ( .A(u2__abc_52155_new_n9290_), .Y(u2__abc_52155_new_n9293_));
INVX1 INVX1_2365 ( .A(u2__abc_52155_new_n9300_), .Y(u2__abc_52155_new_n9301_));
INVX1 INVX1_2366 ( .A(u2__abc_52155_new_n9309_), .Y(u2__abc_52155_new_n9310_));
INVX1 INVX1_2367 ( .A(u2__abc_52155_new_n9311_), .Y(u2__abc_52155_new_n9312_));
INVX1 INVX1_2368 ( .A(u2__abc_52155_new_n9319_), .Y(u2__abc_52155_new_n9320_));
INVX1 INVX1_2369 ( .A(u2__abc_52155_new_n3999_), .Y(u2__abc_52155_new_n9326_));
INVX1 INVX1_237 ( .A(u2__abc_52155_new_n3151_), .Y(u2__abc_52155_new_n3152_));
INVX1 INVX1_2370 ( .A(u2__abc_52155_new_n9327_), .Y(u2__abc_52155_new_n9329_));
INVX1 INVX1_2371 ( .A(u2__abc_52155_new_n9336_), .Y(u2__abc_52155_new_n9337_));
INVX1 INVX1_2372 ( .A(u2__abc_52155_new_n9343_), .Y(u2__abc_52155_new_n9344_));
INVX1 INVX1_2373 ( .A(u2__abc_52155_new_n9347_), .Y(u2__abc_52155_new_n9348_));
INVX1 INVX1_2374 ( .A(u2__abc_52155_new_n9349_), .Y(u2__abc_52155_new_n9350_));
INVX1 INVX1_2375 ( .A(u2__abc_52155_new_n9352_), .Y(u2__abc_52155_new_n9353_));
INVX1 INVX1_2376 ( .A(u2__abc_52155_new_n9356_), .Y(u2__abc_52155_new_n9357_));
INVX1 INVX1_2377 ( .A(u2__abc_52155_new_n9364_), .Y(u2__abc_52155_new_n9365_));
INVX1 INVX1_2378 ( .A(u2__abc_52155_new_n9371_), .Y(u2__abc_52155_new_n9372_));
INVX1 INVX1_2379 ( .A(u2__abc_52155_new_n3947_), .Y(u2__abc_52155_new_n9374_));
INVX1 INVX1_238 ( .A(u2__abc_52155_new_n3157_), .Y(u2__abc_52155_new_n3158_));
INVX1 INVX1_2380 ( .A(u2__abc_52155_new_n9381_), .Y(u2__abc_52155_new_n9382_));
INVX1 INVX1_2381 ( .A(u2__abc_52155_new_n9389_), .Y(u2__abc_52155_new_n9390_));
INVX1 INVX1_2382 ( .A(u2__abc_52155_new_n9393_), .Y(u2__abc_52155_new_n9394_));
INVX1 INVX1_2383 ( .A(u2__abc_52155_new_n9401_), .Y(u2__abc_52155_new_n9402_));
INVX1 INVX1_2384 ( .A(u2__abc_52155_new_n3939_), .Y(u2__abc_52155_new_n9408_));
INVX1 INVX1_2385 ( .A(u2__abc_52155_new_n9409_), .Y(u2__abc_52155_new_n9411_));
INVX1 INVX1_2386 ( .A(u2__abc_52155_new_n9418_), .Y(u2__abc_52155_new_n9419_));
INVX1 INVX1_2387 ( .A(u2__abc_52155_new_n9427_), .Y(u2__abc_52155_new_n9428_));
INVX1 INVX1_2388 ( .A(u2__abc_52155_new_n9429_), .Y(u2__abc_52155_new_n9430_));
INVX1 INVX1_2389 ( .A(u2__abc_52155_new_n9437_), .Y(u2__abc_52155_new_n9438_));
INVX1 INVX1_239 ( .A(u2__abc_52155_new_n3047_), .Y(u2__abc_52155_new_n3159_));
INVX1 INVX1_2390 ( .A(u2__abc_52155_new_n3916_), .Y(u2__abc_52155_new_n9446_));
INVX1 INVX1_2391 ( .A(u2__abc_52155_new_n9444_), .Y(u2__abc_52155_new_n9447_));
INVX1 INVX1_2392 ( .A(u2__abc_52155_new_n9454_), .Y(u2__abc_52155_new_n9455_));
INVX1 INVX1_2393 ( .A(u2__abc_52155_new_n9463_), .Y(u2__abc_52155_new_n9464_));
INVX1 INVX1_2394 ( .A(u2__abc_52155_new_n9465_), .Y(u2__abc_52155_new_n9466_));
INVX1 INVX1_2395 ( .A(u2__abc_52155_new_n9473_), .Y(u2__abc_52155_new_n9474_));
INVX1 INVX1_2396 ( .A(u2__abc_52155_new_n3908_), .Y(u2__abc_52155_new_n9482_));
INVX1 INVX1_2397 ( .A(u2__abc_52155_new_n9480_), .Y(u2__abc_52155_new_n9483_));
INVX1 INVX1_2398 ( .A(u2__abc_52155_new_n9490_), .Y(u2__abc_52155_new_n9491_));
INVX1 INVX1_2399 ( .A(u2__abc_52155_new_n9497_), .Y(u2__abc_52155_new_n9498_));
INVX1 INVX1_24 ( .A(\a[120] ), .Y(_abc_73687_new_n1589_));
INVX1 INVX1_240 ( .A(u2__abc_52155_new_n3160_), .Y(u2__abc_52155_new_n3161_));
INVX1 INVX1_2400 ( .A(u2__abc_52155_new_n9499_), .Y(u2__abc_52155_new_n9500_));
INVX1 INVX1_2401 ( .A(u2__abc_52155_new_n9502_), .Y(u2__abc_52155_new_n9503_));
INVX1 INVX1_2402 ( .A(u2__abc_52155_new_n9504_), .Y(u2__abc_52155_new_n9505_));
INVX1 INVX1_2403 ( .A(u2__abc_52155_new_n9506_), .Y(u2__abc_52155_new_n9507_));
INVX1 INVX1_2404 ( .A(u2__abc_52155_new_n9508_), .Y(u2__abc_52155_new_n9509_));
INVX1 INVX1_2405 ( .A(u2__abc_52155_new_n9510_), .Y(u2__abc_52155_new_n9511_));
INVX1 INVX1_2406 ( .A(u2__abc_52155_new_n9517_), .Y(u2__abc_52155_new_n9518_));
INVX1 INVX1_2407 ( .A(u2__abc_52155_new_n9522_), .Y(u2__abc_52155_new_n9523_));
INVX1 INVX1_2408 ( .A(u2__abc_52155_new_n9529_), .Y(u2__abc_52155_new_n9530_));
INVX1 INVX1_2409 ( .A(u2__abc_52155_new_n3851_), .Y(u2__abc_52155_new_n9538_));
INVX1 INVX1_241 ( .A(sqrto_24_), .Y(u2__abc_52155_new_n3167_));
INVX1 INVX1_2410 ( .A(u2__abc_52155_new_n9536_), .Y(u2__abc_52155_new_n9539_));
INVX1 INVX1_2411 ( .A(u2__abc_52155_new_n9546_), .Y(u2__abc_52155_new_n9547_));
INVX1 INVX1_2412 ( .A(u2__abc_52155_new_n3837_), .Y(u2__abc_52155_new_n9553_));
INVX1 INVX1_2413 ( .A(u2__abc_52155_new_n9556_), .Y(u2__abc_52155_new_n9557_));
INVX1 INVX1_2414 ( .A(u2__abc_52155_new_n9558_), .Y(u2__abc_52155_new_n9559_));
INVX1 INVX1_2415 ( .A(u2__abc_52155_new_n9566_), .Y(u2__abc_52155_new_n9567_));
INVX1 INVX1_2416 ( .A(u2__abc_52155_new_n3834_), .Y(u2__abc_52155_new_n9573_));
INVX1 INVX1_2417 ( .A(u2__abc_52155_new_n3842_), .Y(u2__abc_52155_new_n9576_));
INVX1 INVX1_2418 ( .A(u2__abc_52155_new_n9574_), .Y(u2__abc_52155_new_n9577_));
INVX1 INVX1_2419 ( .A(u2__abc_52155_new_n9584_), .Y(u2__abc_52155_new_n9585_));
INVX1 INVX1_242 ( .A(u2_remHi_24_), .Y(u2__abc_52155_new_n3169_));
INVX1 INVX1_2420 ( .A(u2__abc_52155_new_n9595_), .Y(u2__abc_52155_new_n9596_));
INVX1 INVX1_2421 ( .A(u2__abc_52155_new_n9599_), .Y(u2__abc_52155_new_n9600_));
INVX1 INVX1_2422 ( .A(u2__abc_52155_new_n9607_), .Y(u2__abc_52155_new_n9608_));
INVX1 INVX1_2423 ( .A(u2__abc_52155_new_n3882_), .Y(u2__abc_52155_new_n9616_));
INVX1 INVX1_2424 ( .A(u2__abc_52155_new_n9614_), .Y(u2__abc_52155_new_n9617_));
INVX1 INVX1_2425 ( .A(u2__abc_52155_new_n9624_), .Y(u2__abc_52155_new_n9625_));
INVX1 INVX1_2426 ( .A(u2__abc_52155_new_n9633_), .Y(u2__abc_52155_new_n9634_));
INVX1 INVX1_2427 ( .A(u2__abc_52155_new_n9635_), .Y(u2__abc_52155_new_n9636_));
INVX1 INVX1_2428 ( .A(u2__abc_52155_new_n9643_), .Y(u2__abc_52155_new_n9644_));
INVX1 INVX1_2429 ( .A(u2__abc_52155_new_n3874_), .Y(u2__abc_52155_new_n9650_));
INVX1 INVX1_243 ( .A(sqrto_25_), .Y(u2__abc_52155_new_n3172_));
INVX1 INVX1_2430 ( .A(u2__abc_52155_new_n9651_), .Y(u2__abc_52155_new_n9653_));
INVX1 INVX1_2431 ( .A(u2__abc_52155_new_n9660_), .Y(u2__abc_52155_new_n9661_));
INVX1 INVX1_2432 ( .A(u2__abc_52155_new_n9668_), .Y(u2__abc_52155_new_n9669_));
INVX1 INVX1_2433 ( .A(u2__abc_52155_new_n9677_), .Y(u2__abc_52155_new_n9678_));
INVX1 INVX1_2434 ( .A(u2__abc_52155_new_n9685_), .Y(u2__abc_52155_new_n9686_));
INVX1 INVX1_2435 ( .A(u2__abc_52155_new_n3791_), .Y(u2__abc_52155_new_n9694_));
INVX1 INVX1_2436 ( .A(u2__abc_52155_new_n9692_), .Y(u2__abc_52155_new_n9695_));
INVX1 INVX1_2437 ( .A(u2__abc_52155_new_n9702_), .Y(u2__abc_52155_new_n9703_));
INVX1 INVX1_2438 ( .A(u2__abc_52155_new_n9711_), .Y(u2__abc_52155_new_n9712_));
INVX1 INVX1_2439 ( .A(u2__abc_52155_new_n9713_), .Y(u2__abc_52155_new_n9714_));
INVX1 INVX1_244 ( .A(u2_remHi_25_), .Y(u2__abc_52155_new_n3174_));
INVX1 INVX1_2440 ( .A(u2__abc_52155_new_n9721_), .Y(u2__abc_52155_new_n9722_));
INVX1 INVX1_2441 ( .A(u2__abc_52155_new_n3783_), .Y(u2__abc_52155_new_n9728_));
INVX1 INVX1_2442 ( .A(u2__abc_52155_new_n9729_), .Y(u2__abc_52155_new_n9731_));
INVX1 INVX1_2443 ( .A(u2__abc_52155_new_n9738_), .Y(u2__abc_52155_new_n9739_));
INVX1 INVX1_2444 ( .A(u2__abc_52155_new_n9745_), .Y(u2__abc_52155_new_n9746_));
INVX1 INVX1_2445 ( .A(u2__abc_52155_new_n9753_), .Y(u2__abc_52155_new_n9754_));
INVX1 INVX1_2446 ( .A(u2__abc_52155_new_n9761_), .Y(u2__abc_52155_new_n9762_));
INVX1 INVX1_2447 ( .A(u2__abc_52155_new_n3822_), .Y(u2__abc_52155_new_n9770_));
INVX1 INVX1_2448 ( .A(u2__abc_52155_new_n9768_), .Y(u2__abc_52155_new_n9771_));
INVX1 INVX1_2449 ( .A(u2__abc_52155_new_n9778_), .Y(u2__abc_52155_new_n9779_));
INVX1 INVX1_245 ( .A(u2__abc_52155_new_n3177_), .Y(u2__abc_52155_new_n3178_));
INVX1 INVX1_2450 ( .A(u2__abc_52155_new_n9787_), .Y(u2__abc_52155_new_n9788_));
INVX1 INVX1_2451 ( .A(u2__abc_52155_new_n9789_), .Y(u2__abc_52155_new_n9790_));
INVX1 INVX1_2452 ( .A(u2__abc_52155_new_n9797_), .Y(u2__abc_52155_new_n9798_));
INVX1 INVX1_2453 ( .A(u2__abc_52155_new_n3814_), .Y(u2__abc_52155_new_n9806_));
INVX1 INVX1_2454 ( .A(u2__abc_52155_new_n9804_), .Y(u2__abc_52155_new_n9807_));
INVX1 INVX1_2455 ( .A(u2__abc_52155_new_n9814_), .Y(u2__abc_52155_new_n9815_));
INVX1 INVX1_2456 ( .A(u2__abc_52155_new_n9823_), .Y(u2__abc_52155_new_n9824_));
INVX1 INVX1_2457 ( .A(u2__abc_52155_new_n9833_), .Y(u2__abc_52155_new_n9834_));
INVX1 INVX1_2458 ( .A(u2__abc_52155_new_n9841_), .Y(u2__abc_52155_new_n9842_));
INVX1 INVX1_2459 ( .A(u2__abc_52155_new_n3719_), .Y(u2__abc_52155_new_n9848_));
INVX1 INVX1_246 ( .A(sqrto_23_), .Y(u2__abc_52155_new_n3179_));
INVX1 INVX1_2460 ( .A(u2__abc_52155_new_n9849_), .Y(u2__abc_52155_new_n9851_));
INVX1 INVX1_2461 ( .A(u2__abc_52155_new_n9858_), .Y(u2__abc_52155_new_n9859_));
INVX1 INVX1_2462 ( .A(u2__abc_52155_new_n9866_), .Y(u2__abc_52155_new_n9867_));
INVX1 INVX1_2463 ( .A(u2__abc_52155_new_n9870_), .Y(u2__abc_52155_new_n9871_));
INVX1 INVX1_2464 ( .A(u2__abc_52155_new_n9878_), .Y(u2__abc_52155_new_n9879_));
INVX1 INVX1_2465 ( .A(u2__abc_52155_new_n3734_), .Y(u2__abc_52155_new_n9885_));
INVX1 INVX1_2466 ( .A(u2__abc_52155_new_n9886_), .Y(u2__abc_52155_new_n9888_));
INVX1 INVX1_2467 ( .A(u2__abc_52155_new_n9895_), .Y(u2__abc_52155_new_n9896_));
INVX1 INVX1_2468 ( .A(u2__abc_52155_new_n9908_), .Y(u2__abc_52155_new_n9909_));
INVX1 INVX1_2469 ( .A(u2__abc_52155_new_n9916_), .Y(u2__abc_52155_new_n9917_));
INVX1 INVX1_247 ( .A(u2__abc_52155_new_n3180_), .Y(u2__abc_52155_new_n3181_));
INVX1 INVX1_2470 ( .A(u2__abc_52155_new_n9923_), .Y(u2__abc_52155_new_n9924_));
INVX1 INVX1_2471 ( .A(u2__abc_52155_new_n9925_), .Y(u2__abc_52155_new_n9926_));
INVX1 INVX1_2472 ( .A(u2__abc_52155_new_n9933_), .Y(u2__abc_52155_new_n9934_));
INVX1 INVX1_2473 ( .A(u2__abc_52155_new_n9940_), .Y(u2__abc_52155_new_n9941_));
INVX1 INVX1_2474 ( .A(u2__abc_52155_new_n9942_), .Y(u2__abc_52155_new_n9943_));
INVX1 INVX1_2475 ( .A(u2__abc_52155_new_n9950_), .Y(u2__abc_52155_new_n9951_));
INVX1 INVX1_2476 ( .A(u2__abc_52155_new_n3750_), .Y(u2__abc_52155_new_n9959_));
INVX1 INVX1_2477 ( .A(u2__abc_52155_new_n9957_), .Y(u2__abc_52155_new_n9960_));
INVX1 INVX1_2478 ( .A(u2__abc_52155_new_n9967_), .Y(u2__abc_52155_new_n9968_));
INVX1 INVX1_2479 ( .A(u2__abc_52155_new_n9984_), .Y(u2__abc_52155_new_n9985_));
INVX1 INVX1_248 ( .A(u2_remHi_23_), .Y(u2__abc_52155_new_n3182_));
INVX1 INVX1_2480 ( .A(u2__abc_52155_new_n9992_), .Y(u2__abc_52155_new_n9993_));
INVX1 INVX1_2481 ( .A(u2__abc_52155_new_n3656_), .Y(u2__abc_52155_new_n9999_));
INVX1 INVX1_2482 ( .A(u2__abc_52155_new_n10000_), .Y(u2__abc_52155_new_n10002_));
INVX1 INVX1_2483 ( .A(u2__abc_52155_new_n10009_), .Y(u2__abc_52155_new_n10010_));
INVX1 INVX1_2484 ( .A(u2__abc_52155_new_n10017_), .Y(u2__abc_52155_new_n10018_));
INVX1 INVX1_2485 ( .A(u2__abc_52155_new_n10021_), .Y(u2__abc_52155_new_n10022_));
INVX1 INVX1_2486 ( .A(u2__abc_52155_new_n10029_), .Y(u2__abc_52155_new_n10030_));
INVX1 INVX1_2487 ( .A(u2__abc_52155_new_n3671_), .Y(u2__abc_52155_new_n10038_));
INVX1 INVX1_2488 ( .A(u2__abc_52155_new_n10036_), .Y(u2__abc_52155_new_n10039_));
INVX1 INVX1_2489 ( .A(u2__abc_52155_new_n10046_), .Y(u2__abc_52155_new_n10047_));
INVX1 INVX1_249 ( .A(u2__abc_52155_new_n3183_), .Y(u2__abc_52155_new_n3184_));
INVX1 INVX1_2490 ( .A(u2__abc_52155_new_n10059_), .Y(u2__abc_52155_new_n10060_));
INVX1 INVX1_2491 ( .A(u2__abc_52155_new_n10067_), .Y(u2__abc_52155_new_n10068_));
INVX1 INVX1_2492 ( .A(u2__abc_52155_new_n3695_), .Y(u2__abc_52155_new_n10076_));
INVX1 INVX1_2493 ( .A(u2__abc_52155_new_n10074_), .Y(u2__abc_52155_new_n10077_));
INVX1 INVX1_2494 ( .A(u2__abc_52155_new_n10084_), .Y(u2__abc_52155_new_n10085_));
INVX1 INVX1_2495 ( .A(u2__abc_52155_new_n10093_), .Y(u2__abc_52155_new_n10094_));
INVX1 INVX1_2496 ( .A(u2__abc_52155_new_n10095_), .Y(u2__abc_52155_new_n10096_));
INVX1 INVX1_2497 ( .A(u2_remHi_126_), .Y(u2__abc_52155_new_n10103_));
INVX1 INVX1_2498 ( .A(u2__abc_52155_new_n10104_), .Y(u2__abc_52155_new_n10105_));
INVX1 INVX1_2499 ( .A(u2__abc_52155_new_n3687_), .Y(u2__abc_52155_new_n10113_));
INVX1 INVX1_25 ( .A(_abc_73687_new_n1578_), .Y(_abc_73687_new_n1590_));
INVX1 INVX1_250 ( .A(sqrto_22_), .Y(u2__abc_52155_new_n3186_));
INVX1 INVX1_2500 ( .A(u2__abc_52155_new_n10111_), .Y(u2__abc_52155_new_n10114_));
INVX1 INVX1_2501 ( .A(u2__abc_52155_new_n10121_), .Y(u2__abc_52155_new_n10122_));
INVX1 INVX1_2502 ( .A(u2__abc_52155_new_n10128_), .Y(u2__abc_52155_new_n10129_));
INVX1 INVX1_2503 ( .A(u2__abc_52155_new_n10130_), .Y(u2__abc_52155_new_n10131_));
INVX1 INVX1_2504 ( .A(u2__abc_52155_new_n10132_), .Y(u2__abc_52155_new_n10133_));
INVX1 INVX1_2505 ( .A(u2__abc_52155_new_n10134_), .Y(u2__abc_52155_new_n10135_));
INVX1 INVX1_2506 ( .A(u2__abc_52155_new_n10136_), .Y(u2__abc_52155_new_n10137_));
INVX1 INVX1_2507 ( .A(u2__abc_52155_new_n10140_), .Y(u2__abc_52155_new_n10141_));
INVX1 INVX1_2508 ( .A(u2__abc_52155_new_n10142_), .Y(u2__abc_52155_new_n10143_));
INVX1 INVX1_2509 ( .A(u2__abc_52155_new_n10149_), .Y(u2__abc_52155_new_n10150_));
INVX1 INVX1_251 ( .A(u2__abc_52155_new_n3187_), .Y(u2__abc_52155_new_n3188_));
INVX1 INVX1_2510 ( .A(u2__abc_52155_new_n10151_), .Y(u2__abc_52155_new_n10152_));
INVX1 INVX1_2511 ( .A(u2__abc_52155_new_n10159_), .Y(u2__abc_52155_new_n10160_));
INVX1 INVX1_2512 ( .A(u2__abc_52155_new_n5244_), .Y(u2__abc_52155_new_n10166_));
INVX1 INVX1_2513 ( .A(u2__abc_52155_new_n10167_), .Y(u2__abc_52155_new_n10169_));
INVX1 INVX1_2514 ( .A(u2__abc_52155_new_n10176_), .Y(u2__abc_52155_new_n10177_));
INVX1 INVX1_2515 ( .A(u2__abc_52155_new_n5250_), .Y(u2__abc_52155_new_n10183_));
INVX1 INVX1_2516 ( .A(u2__abc_52155_new_n10185_), .Y(u2__abc_52155_new_n10186_));
INVX1 INVX1_2517 ( .A(u2__abc_52155_new_n10189_), .Y(u2__abc_52155_new_n10190_));
INVX1 INVX1_2518 ( .A(u2__abc_52155_new_n10197_), .Y(u2__abc_52155_new_n10198_));
INVX1 INVX1_2519 ( .A(u2__abc_52155_new_n5247_), .Y(u2__abc_52155_new_n10204_));
INVX1 INVX1_252 ( .A(u2_remHi_22_), .Y(u2__abc_52155_new_n3189_));
INVX1 INVX1_2520 ( .A(u2__abc_52155_new_n5255_), .Y(u2__abc_52155_new_n10207_));
INVX1 INVX1_2521 ( .A(u2__abc_52155_new_n10205_), .Y(u2__abc_52155_new_n10208_));
INVX1 INVX1_2522 ( .A(u2__abc_52155_new_n10215_), .Y(u2__abc_52155_new_n10216_));
INVX1 INVX1_2523 ( .A(u2__abc_52155_new_n5279_), .Y(u2__abc_52155_new_n10222_));
INVX1 INVX1_2524 ( .A(u2__abc_52155_new_n10229_), .Y(u2__abc_52155_new_n10230_));
INVX1 INVX1_2525 ( .A(u2__abc_52155_new_n10237_), .Y(u2__abc_52155_new_n10238_));
INVX1 INVX1_2526 ( .A(u2__abc_52155_new_n5274_), .Y(u2__abc_52155_new_n10244_));
INVX1 INVX1_2527 ( .A(u2__abc_52155_new_n5276_), .Y(u2__abc_52155_new_n10245_));
INVX1 INVX1_2528 ( .A(u2__abc_52155_new_n10246_), .Y(u2__abc_52155_new_n10248_));
INVX1 INVX1_2529 ( .A(u2__abc_52155_new_n10255_), .Y(u2__abc_52155_new_n10256_));
INVX1 INVX1_253 ( .A(u2__abc_52155_new_n3190_), .Y(u2__abc_52155_new_n3191_));
INVX1 INVX1_2530 ( .A(u2__abc_52155_new_n5263_), .Y(u2__abc_52155_new_n10262_));
INVX1 INVX1_2531 ( .A(u2__abc_52155_new_n10263_), .Y(u2__abc_52155_new_n10264_));
INVX1 INVX1_2532 ( .A(u2__abc_52155_new_n10266_), .Y(u2__abc_52155_new_n10267_));
INVX1 INVX1_2533 ( .A(u2__abc_52155_new_n10268_), .Y(u2__abc_52155_new_n10269_));
INVX1 INVX1_2534 ( .A(u2__abc_52155_new_n10276_), .Y(u2__abc_52155_new_n10277_));
INVX1 INVX1_2535 ( .A(u2__abc_52155_new_n5260_), .Y(u2__abc_52155_new_n10283_));
INVX1 INVX1_2536 ( .A(u2__abc_52155_new_n5268_), .Y(u2__abc_52155_new_n10286_));
INVX1 INVX1_2537 ( .A(u2__abc_52155_new_n10284_), .Y(u2__abc_52155_new_n10287_));
INVX1 INVX1_2538 ( .A(u2__abc_52155_new_n10294_), .Y(u2__abc_52155_new_n10295_));
INVX1 INVX1_2539 ( .A(u2__abc_52155_new_n10301_), .Y(u2__abc_52155_new_n10302_));
INVX1 INVX1_254 ( .A(sqrto_28_), .Y(u2__abc_52155_new_n3195_));
INVX1 INVX1_2540 ( .A(u2__abc_52155_new_n10308_), .Y(u2__abc_52155_new_n10309_));
INVX1 INVX1_2541 ( .A(u2__abc_52155_new_n10312_), .Y(u2__abc_52155_new_n10313_));
INVX1 INVX1_2542 ( .A(u2__abc_52155_new_n10320_), .Y(u2__abc_52155_new_n10321_));
INVX1 INVX1_2543 ( .A(u2__abc_52155_new_n5198_), .Y(u2__abc_52155_new_n10327_));
INVX1 INVX1_2544 ( .A(u2__abc_52155_new_n10328_), .Y(u2__abc_52155_new_n10329_));
INVX1 INVX1_2545 ( .A(u2__abc_52155_new_n10337_), .Y(u2__abc_52155_new_n10338_));
INVX1 INVX1_2546 ( .A(u2__abc_52155_new_n5177_), .Y(u2__abc_52155_new_n10344_));
INVX1 INVX1_2547 ( .A(u2__abc_52155_new_n10347_), .Y(u2__abc_52155_new_n10348_));
INVX1 INVX1_2548 ( .A(u2__abc_52155_new_n10355_), .Y(u2__abc_52155_new_n10356_));
INVX1 INVX1_2549 ( .A(u2__abc_52155_new_n5174_), .Y(u2__abc_52155_new_n10362_));
INVX1 INVX1_255 ( .A(u2__abc_52155_new_n3196_), .Y(u2__abc_52155_new_n3197_));
INVX1 INVX1_2550 ( .A(u2__abc_52155_new_n5182_), .Y(u2__abc_52155_new_n10365_));
INVX1 INVX1_2551 ( .A(u2__abc_52155_new_n10363_), .Y(u2__abc_52155_new_n10366_));
INVX1 INVX1_2552 ( .A(u2__abc_52155_new_n10373_), .Y(u2__abc_52155_new_n10374_));
INVX1 INVX1_2553 ( .A(u2__abc_52155_new_n10385_), .Y(u2__abc_52155_new_n10386_));
INVX1 INVX1_2554 ( .A(u2__abc_52155_new_n10389_), .Y(u2__abc_52155_new_n10390_));
INVX1 INVX1_2555 ( .A(u2__abc_52155_new_n10397_), .Y(u2__abc_52155_new_n10398_));
INVX1 INVX1_2556 ( .A(u2__abc_52155_new_n5222_), .Y(u2__abc_52155_new_n10406_));
INVX1 INVX1_2557 ( .A(u2__abc_52155_new_n10404_), .Y(u2__abc_52155_new_n10407_));
INVX1 INVX1_2558 ( .A(u2__abc_52155_new_n10414_), .Y(u2__abc_52155_new_n10415_));
INVX1 INVX1_2559 ( .A(u2__abc_52155_new_n10423_), .Y(u2__abc_52155_new_n10424_));
INVX1 INVX1_256 ( .A(u2_remHi_28_), .Y(u2__abc_52155_new_n3198_));
INVX1 INVX1_2560 ( .A(u2__abc_52155_new_n10425_), .Y(u2__abc_52155_new_n10426_));
INVX1 INVX1_2561 ( .A(u2__abc_52155_new_n10433_), .Y(u2__abc_52155_new_n10434_));
INVX1 INVX1_2562 ( .A(u2__abc_52155_new_n5214_), .Y(u2__abc_52155_new_n10442_));
INVX1 INVX1_2563 ( .A(u2__abc_52155_new_n10440_), .Y(u2__abc_52155_new_n10443_));
INVX1 INVX1_2564 ( .A(u2__abc_52155_new_n10450_), .Y(u2__abc_52155_new_n10451_));
INVX1 INVX1_2565 ( .A(u2__abc_52155_new_n10459_), .Y(u2__abc_52155_new_n10460_));
INVX1 INVX1_2566 ( .A(u2__abc_52155_new_n10469_), .Y(u2__abc_52155_new_n10470_));
INVX1 INVX1_2567 ( .A(u2__abc_52155_new_n10477_), .Y(u2__abc_52155_new_n10478_));
INVX1 INVX1_2568 ( .A(u2__abc_52155_new_n5161_), .Y(u2__abc_52155_new_n10484_));
INVX1 INVX1_2569 ( .A(u2__abc_52155_new_n10485_), .Y(u2__abc_52155_new_n10486_));
INVX1 INVX1_257 ( .A(u2__abc_52155_new_n3199_), .Y(u2__abc_52155_new_n3200_));
INVX1 INVX1_2570 ( .A(u2__abc_52155_new_n10494_), .Y(u2__abc_52155_new_n10495_));
INVX1 INVX1_2571 ( .A(u2__abc_52155_new_n5147_), .Y(u2__abc_52155_new_n10501_));
INVX1 INVX1_2572 ( .A(u2__abc_52155_new_n10504_), .Y(u2__abc_52155_new_n10505_));
INVX1 INVX1_2573 ( .A(u2__abc_52155_new_n10512_), .Y(u2__abc_52155_new_n10513_));
INVX1 INVX1_2574 ( .A(u2__abc_52155_new_n5144_), .Y(u2__abc_52155_new_n10519_));
INVX1 INVX1_2575 ( .A(u2__abc_52155_new_n5152_), .Y(u2__abc_52155_new_n10522_));
INVX1 INVX1_2576 ( .A(u2__abc_52155_new_n10520_), .Y(u2__abc_52155_new_n10523_));
INVX1 INVX1_2577 ( .A(u2__abc_52155_new_n10530_), .Y(u2__abc_52155_new_n10531_));
INVX1 INVX1_2578 ( .A(u2__abc_52155_new_n10539_), .Y(u2__abc_52155_new_n10540_));
INVX1 INVX1_2579 ( .A(u2__abc_52155_new_n10541_), .Y(u2__abc_52155_new_n10542_));
INVX1 INVX1_258 ( .A(u2_remHi_29_), .Y(u2__abc_52155_new_n3202_));
INVX1 INVX1_2580 ( .A(u2__abc_52155_new_n10549_), .Y(u2__abc_52155_new_n10550_));
INVX1 INVX1_2581 ( .A(u2__abc_52155_new_n10556_), .Y(u2__abc_52155_new_n10557_));
INVX1 INVX1_2582 ( .A(u2__abc_52155_new_n10558_), .Y(u2__abc_52155_new_n10559_));
INVX1 INVX1_2583 ( .A(u2__abc_52155_new_n10566_), .Y(u2__abc_52155_new_n10567_));
INVX1 INVX1_2584 ( .A(u2__abc_52155_new_n10573_), .Y(u2__abc_52155_new_n10574_));
INVX1 INVX1_2585 ( .A(u2__abc_52155_new_n10575_), .Y(u2__abc_52155_new_n10576_));
INVX1 INVX1_2586 ( .A(u2__abc_52155_new_n10583_), .Y(u2__abc_52155_new_n10584_));
INVX1 INVX1_2587 ( .A(u2__abc_52155_new_n5125_), .Y(u2__abc_52155_new_n10592_));
INVX1 INVX1_2588 ( .A(u2__abc_52155_new_n10590_), .Y(u2__abc_52155_new_n10593_));
INVX1 INVX1_2589 ( .A(u2__abc_52155_new_n10600_), .Y(u2__abc_52155_new_n10601_));
INVX1 INVX1_259 ( .A(u2__abc_52155_new_n3203_), .Y(u2__abc_52155_new_n3204_));
INVX1 INVX1_2590 ( .A(u2__abc_52155_new_n10619_), .Y(u2__abc_52155_new_n10620_));
INVX1 INVX1_2591 ( .A(u2__abc_52155_new_n10623_), .Y(u2__abc_52155_new_n10624_));
INVX1 INVX1_2592 ( .A(u2__abc_52155_new_n10631_), .Y(u2__abc_52155_new_n10632_));
INVX1 INVX1_2593 ( .A(u2__abc_52155_new_n5070_), .Y(u2__abc_52155_new_n10640_));
INVX1 INVX1_2594 ( .A(u2__abc_52155_new_n10638_), .Y(u2__abc_52155_new_n10641_));
INVX1 INVX1_2595 ( .A(u2__abc_52155_new_n10648_), .Y(u2__abc_52155_new_n10649_));
INVX1 INVX1_2596 ( .A(u2__abc_52155_new_n10657_), .Y(u2__abc_52155_new_n10658_));
INVX1 INVX1_2597 ( .A(u2__abc_52155_new_n10659_), .Y(u2__abc_52155_new_n10660_));
INVX1 INVX1_2598 ( .A(u2__abc_52155_new_n10667_), .Y(u2__abc_52155_new_n10668_));
INVX1 INVX1_2599 ( .A(u2__abc_52155_new_n5062_), .Y(u2__abc_52155_new_n10676_));
INVX1 INVX1_26 ( .A(_abc_73687_new_n1582_), .Y(_abc_73687_new_n1594_));
INVX1 INVX1_260 ( .A(sqrto_29_), .Y(u2__abc_52155_new_n3205_));
INVX1 INVX1_2600 ( .A(u2__abc_52155_new_n10674_), .Y(u2__abc_52155_new_n10677_));
INVX1 INVX1_2601 ( .A(u2__abc_52155_new_n10684_), .Y(u2__abc_52155_new_n10685_));
INVX1 INVX1_2602 ( .A(u2__abc_52155_new_n10691_), .Y(u2__abc_52155_new_n10692_));
INVX1 INVX1_2603 ( .A(u2__abc_52155_new_n10699_), .Y(u2__abc_52155_new_n10700_));
INVX1 INVX1_2604 ( .A(u2__abc_52155_new_n10707_), .Y(u2__abc_52155_new_n10708_));
INVX1 INVX1_2605 ( .A(u2__abc_52155_new_n5101_), .Y(u2__abc_52155_new_n10716_));
INVX1 INVX1_2606 ( .A(u2__abc_52155_new_n10714_), .Y(u2__abc_52155_new_n10717_));
INVX1 INVX1_2607 ( .A(u2__abc_52155_new_n10724_), .Y(u2__abc_52155_new_n10725_));
INVX1 INVX1_2608 ( .A(u2__abc_52155_new_n10733_), .Y(u2__abc_52155_new_n10734_));
INVX1 INVX1_2609 ( .A(u2__abc_52155_new_n10735_), .Y(u2__abc_52155_new_n10736_));
INVX1 INVX1_261 ( .A(u2__abc_52155_new_n3206_), .Y(u2__abc_52155_new_n3207_));
INVX1 INVX1_2610 ( .A(u2__abc_52155_new_n10743_), .Y(u2__abc_52155_new_n10744_));
INVX1 INVX1_2611 ( .A(u2__abc_52155_new_n5093_), .Y(u2__abc_52155_new_n10752_));
INVX1 INVX1_2612 ( .A(u2__abc_52155_new_n10750_), .Y(u2__abc_52155_new_n10753_));
INVX1 INVX1_2613 ( .A(u2__abc_52155_new_n10760_), .Y(u2__abc_52155_new_n10761_));
INVX1 INVX1_2614 ( .A(u2__abc_52155_new_n10770_), .Y(u2__abc_52155_new_n10771_));
INVX1 INVX1_2615 ( .A(u2__abc_52155_new_n10781_), .Y(u2__abc_52155_new_n10782_));
INVX1 INVX1_2616 ( .A(u2__abc_52155_new_n10789_), .Y(u2__abc_52155_new_n10790_));
INVX1 INVX1_2617 ( .A(u2__abc_52155_new_n5005_), .Y(u2__abc_52155_new_n10798_));
INVX1 INVX1_2618 ( .A(u2__abc_52155_new_n10796_), .Y(u2__abc_52155_new_n10799_));
INVX1 INVX1_2619 ( .A(u2__abc_52155_new_n10806_), .Y(u2__abc_52155_new_n10807_));
INVX1 INVX1_262 ( .A(sqrto_27_), .Y(u2__abc_52155_new_n3210_));
INVX1 INVX1_2620 ( .A(u2__abc_52155_new_n4991_), .Y(u2__abc_52155_new_n10813_));
INVX1 INVX1_2621 ( .A(u2__abc_52155_new_n10816_), .Y(u2__abc_52155_new_n10817_));
INVX1 INVX1_2622 ( .A(u2__abc_52155_new_n10818_), .Y(u2__abc_52155_new_n10819_));
INVX1 INVX1_2623 ( .A(u2__abc_52155_new_n10826_), .Y(u2__abc_52155_new_n10827_));
INVX1 INVX1_2624 ( .A(u2__abc_52155_new_n4988_), .Y(u2__abc_52155_new_n10833_));
INVX1 INVX1_2625 ( .A(u2__abc_52155_new_n4996_), .Y(u2__abc_52155_new_n10836_));
INVX1 INVX1_2626 ( .A(u2__abc_52155_new_n10834_), .Y(u2__abc_52155_new_n10837_));
INVX1 INVX1_2627 ( .A(u2__abc_52155_new_n10844_), .Y(u2__abc_52155_new_n10845_));
INVX1 INVX1_2628 ( .A(u2__abc_52155_new_n10855_), .Y(u2__abc_52155_new_n10856_));
INVX1 INVX1_2629 ( .A(u2__abc_52155_new_n10859_), .Y(u2__abc_52155_new_n10860_));
INVX1 INVX1_263 ( .A(u2__abc_52155_new_n3211_), .Y(u2__abc_52155_new_n3212_));
INVX1 INVX1_2630 ( .A(u2__abc_52155_new_n10867_), .Y(u2__abc_52155_new_n10868_));
INVX1 INVX1_2631 ( .A(u2__abc_52155_new_n10874_), .Y(u2__abc_52155_new_n10875_));
INVX1 INVX1_2632 ( .A(u2__abc_52155_new_n10876_), .Y(u2__abc_52155_new_n10877_));
INVX1 INVX1_2633 ( .A(u2__abc_52155_new_n10884_), .Y(u2__abc_52155_new_n10885_));
INVX1 INVX1_2634 ( .A(u2__abc_52155_new_n10891_), .Y(u2__abc_52155_new_n10892_));
INVX1 INVX1_2635 ( .A(u2__abc_52155_new_n10893_), .Y(u2__abc_52155_new_n10894_));
INVX1 INVX1_2636 ( .A(u2__abc_52155_new_n10901_), .Y(u2__abc_52155_new_n10902_));
INVX1 INVX1_2637 ( .A(u2__abc_52155_new_n5028_), .Y(u2__abc_52155_new_n10910_));
INVX1 INVX1_2638 ( .A(u2__abc_52155_new_n10908_), .Y(u2__abc_52155_new_n10911_));
INVX1 INVX1_2639 ( .A(u2__abc_52155_new_n10918_), .Y(u2__abc_52155_new_n10919_));
INVX1 INVX1_264 ( .A(u2_remHi_27_), .Y(u2__abc_52155_new_n3213_));
INVX1 INVX1_2640 ( .A(u2__abc_52155_new_n10935_), .Y(u2__abc_52155_new_n10936_));
INVX1 INVX1_2641 ( .A(u2__abc_52155_new_n10943_), .Y(u2__abc_52155_new_n10944_));
INVX1 INVX1_2642 ( .A(u2__abc_52155_new_n4976_), .Y(u2__abc_52155_new_n10950_));
INVX1 INVX1_2643 ( .A(u2__abc_52155_new_n10951_), .Y(u2__abc_52155_new_n10952_));
INVX1 INVX1_2644 ( .A(u2__abc_52155_new_n10960_), .Y(u2__abc_52155_new_n10961_));
INVX1 INVX1_2645 ( .A(u2__abc_52155_new_n10968_), .Y(u2__abc_52155_new_n10969_));
INVX1 INVX1_2646 ( .A(u2__abc_52155_new_n10972_), .Y(u2__abc_52155_new_n10973_));
INVX1 INVX1_2647 ( .A(u2__abc_52155_new_n10980_), .Y(u2__abc_52155_new_n10981_));
INVX1 INVX1_2648 ( .A(u2__abc_52155_new_n4968_), .Y(u2__abc_52155_new_n10989_));
INVX1 INVX1_2649 ( .A(u2__abc_52155_new_n10987_), .Y(u2__abc_52155_new_n10990_));
INVX1 INVX1_265 ( .A(u2__abc_52155_new_n3214_), .Y(u2__abc_52155_new_n3215_));
INVX1 INVX1_2650 ( .A(u2__abc_52155_new_n10997_), .Y(u2__abc_52155_new_n10998_));
INVX1 INVX1_2651 ( .A(u2__abc_52155_new_n11006_), .Y(u2__abc_52155_new_n11007_));
INVX1 INVX1_2652 ( .A(u2__abc_52155_new_n11008_), .Y(u2__abc_52155_new_n11009_));
INVX1 INVX1_2653 ( .A(u2__abc_52155_new_n11016_), .Y(u2__abc_52155_new_n11017_));
INVX1 INVX1_2654 ( .A(u2__abc_52155_new_n4945_), .Y(u2__abc_52155_new_n11025_));
INVX1 INVX1_2655 ( .A(u2__abc_52155_new_n11023_), .Y(u2__abc_52155_new_n11026_));
INVX1 INVX1_2656 ( .A(u2__abc_52155_new_n11033_), .Y(u2__abc_52155_new_n11034_));
INVX1 INVX1_2657 ( .A(u2__abc_52155_new_n11042_), .Y(u2__abc_52155_new_n11043_));
INVX1 INVX1_2658 ( .A(u2__abc_52155_new_n11044_), .Y(u2__abc_52155_new_n11045_));
INVX1 INVX1_2659 ( .A(u2__abc_52155_new_n11052_), .Y(u2__abc_52155_new_n11053_));
INVX1 INVX1_266 ( .A(sqrto_26_), .Y(u2__abc_52155_new_n3217_));
INVX1 INVX1_2660 ( .A(u2__abc_52155_new_n4937_), .Y(u2__abc_52155_new_n11061_));
INVX1 INVX1_2661 ( .A(u2__abc_52155_new_n11059_), .Y(u2__abc_52155_new_n11062_));
INVX1 INVX1_2662 ( .A(u2__abc_52155_new_n11069_), .Y(u2__abc_52155_new_n11070_));
INVX1 INVX1_2663 ( .A(u2__abc_52155_new_n11076_), .Y(u2__abc_52155_new_n11077_));
INVX1 INVX1_2664 ( .A(u2__abc_52155_new_n11079_), .Y(u2__abc_52155_new_n11080_));
INVX1 INVX1_2665 ( .A(u2__abc_52155_new_n11081_), .Y(u2__abc_52155_new_n11082_));
INVX1 INVX1_2666 ( .A(u2__abc_52155_new_n11083_), .Y(u2__abc_52155_new_n11084_));
INVX1 INVX1_2667 ( .A(u2__abc_52155_new_n11085_), .Y(u2__abc_52155_new_n11086_));
INVX1 INVX1_2668 ( .A(u2__abc_52155_new_n11087_), .Y(u2__abc_52155_new_n11088_));
INVX1 INVX1_2669 ( .A(u2__abc_52155_new_n11093_), .Y(u2__abc_52155_new_n11094_));
INVX1 INVX1_267 ( .A(u2__abc_52155_new_n3218_), .Y(u2__abc_52155_new_n3219_));
INVX1 INVX1_2670 ( .A(u2__abc_52155_new_n11097_), .Y(u2__abc_52155_new_n11098_));
INVX1 INVX1_2671 ( .A(u2__abc_52155_new_n11105_), .Y(u2__abc_52155_new_n11106_));
INVX1 INVX1_2672 ( .A(u2__abc_52155_new_n4919_), .Y(u2__abc_52155_new_n11112_));
INVX1 INVX1_2673 ( .A(u2__abc_52155_new_n11113_), .Y(u2__abc_52155_new_n11115_));
INVX1 INVX1_2674 ( .A(u2__abc_52155_new_n11122_), .Y(u2__abc_52155_new_n11123_));
INVX1 INVX1_2675 ( .A(u2__abc_52155_new_n11130_), .Y(u2__abc_52155_new_n11131_));
INVX1 INVX1_2676 ( .A(u2__abc_52155_new_n11134_), .Y(u2__abc_52155_new_n11135_));
INVX1 INVX1_2677 ( .A(u2__abc_52155_new_n11142_), .Y(u2__abc_52155_new_n11143_));
INVX1 INVX1_2678 ( .A(u2__abc_52155_new_n4904_), .Y(u2__abc_52155_new_n11151_));
INVX1 INVX1_2679 ( .A(u2__abc_52155_new_n11149_), .Y(u2__abc_52155_new_n11152_));
INVX1 INVX1_268 ( .A(u2_remHi_26_), .Y(u2__abc_52155_new_n3220_));
INVX1 INVX1_2680 ( .A(u2__abc_52155_new_n11159_), .Y(u2__abc_52155_new_n11160_));
INVX1 INVX1_2681 ( .A(u2__abc_52155_new_n11168_), .Y(u2__abc_52155_new_n11169_));
INVX1 INVX1_2682 ( .A(u2__abc_52155_new_n11170_), .Y(u2__abc_52155_new_n11171_));
INVX1 INVX1_2683 ( .A(u2__abc_52155_new_n11178_), .Y(u2__abc_52155_new_n11179_));
INVX1 INVX1_2684 ( .A(u2__abc_52155_new_n4881_), .Y(u2__abc_52155_new_n11187_));
INVX1 INVX1_2685 ( .A(u2__abc_52155_new_n11185_), .Y(u2__abc_52155_new_n11188_));
INVX1 INVX1_2686 ( .A(u2__abc_52155_new_n11195_), .Y(u2__abc_52155_new_n11196_));
INVX1 INVX1_2687 ( .A(u2__abc_52155_new_n11204_), .Y(u2__abc_52155_new_n11205_));
INVX1 INVX1_2688 ( .A(u2__abc_52155_new_n11206_), .Y(u2__abc_52155_new_n11207_));
INVX1 INVX1_2689 ( .A(u2__abc_52155_new_n11214_), .Y(u2__abc_52155_new_n11215_));
INVX1 INVX1_269 ( .A(u2__abc_52155_new_n3221_), .Y(u2__abc_52155_new_n3222_));
INVX1 INVX1_2690 ( .A(u2__abc_52155_new_n4873_), .Y(u2__abc_52155_new_n11223_));
INVX1 INVX1_2691 ( .A(u2__abc_52155_new_n11221_), .Y(u2__abc_52155_new_n11224_));
INVX1 INVX1_2692 ( .A(u2__abc_52155_new_n11231_), .Y(u2__abc_52155_new_n11232_));
INVX1 INVX1_2693 ( .A(u2__abc_52155_new_n11239_), .Y(u2__abc_52155_new_n11240_));
INVX1 INVX1_2694 ( .A(u2__abc_52155_new_n11241_), .Y(u2__abc_52155_new_n11242_));
INVX1 INVX1_2695 ( .A(u2__abc_52155_new_n11244_), .Y(u2__abc_52155_new_n11245_));
INVX1 INVX1_2696 ( .A(u2__abc_52155_new_n11253_), .Y(u2__abc_52155_new_n11254_));
INVX1 INVX1_2697 ( .A(u2__abc_52155_new_n11261_), .Y(u2__abc_52155_new_n11262_));
INVX1 INVX1_2698 ( .A(u2__abc_52155_new_n4810_), .Y(u2__abc_52155_new_n11270_));
INVX1 INVX1_2699 ( .A(u2__abc_52155_new_n11268_), .Y(u2__abc_52155_new_n11271_));
INVX1 INVX1_27 ( .A(_abc_73687_new_n1592_), .Y(_abc_73687_new_n1595_));
INVX1 INVX1_270 ( .A(sqrto_16_), .Y(u2__abc_52155_new_n3227_));
INVX1 INVX1_2700 ( .A(u2__abc_52155_new_n11278_), .Y(u2__abc_52155_new_n11279_));
INVX1 INVX1_2701 ( .A(u2__abc_52155_new_n11286_), .Y(u2__abc_52155_new_n11287_));
INVX1 INVX1_2702 ( .A(u2__abc_52155_new_n11290_), .Y(u2__abc_52155_new_n11291_));
INVX1 INVX1_2703 ( .A(u2__abc_52155_new_n11298_), .Y(u2__abc_52155_new_n11299_));
INVX1 INVX1_2704 ( .A(u2__abc_52155_new_n4825_), .Y(u2__abc_52155_new_n11307_));
INVX1 INVX1_2705 ( .A(u2__abc_52155_new_n11305_), .Y(u2__abc_52155_new_n11308_));
INVX1 INVX1_2706 ( .A(u2__abc_52155_new_n11315_), .Y(u2__abc_52155_new_n11316_));
INVX1 INVX1_2707 ( .A(u2__abc_52155_new_n11328_), .Y(u2__abc_52155_new_n11329_));
INVX1 INVX1_2708 ( .A(u2__abc_52155_new_n11336_), .Y(u2__abc_52155_new_n11337_));
INVX1 INVX1_2709 ( .A(u2__abc_52155_new_n4849_), .Y(u2__abc_52155_new_n11345_));
INVX1 INVX1_271 ( .A(u2_remHi_16_), .Y(u2__abc_52155_new_n3229_));
INVX1 INVX1_2710 ( .A(u2__abc_52155_new_n11343_), .Y(u2__abc_52155_new_n11346_));
INVX1 INVX1_2711 ( .A(u2__abc_52155_new_n11353_), .Y(u2__abc_52155_new_n11354_));
INVX1 INVX1_2712 ( .A(u2__abc_52155_new_n11362_), .Y(u2__abc_52155_new_n11363_));
INVX1 INVX1_2713 ( .A(u2__abc_52155_new_n11364_), .Y(u2__abc_52155_new_n11365_));
INVX1 INVX1_2714 ( .A(u2__abc_52155_new_n11372_), .Y(u2__abc_52155_new_n11373_));
INVX1 INVX1_2715 ( .A(u2__abc_52155_new_n4841_), .Y(u2__abc_52155_new_n11381_));
INVX1 INVX1_2716 ( .A(u2__abc_52155_new_n11379_), .Y(u2__abc_52155_new_n11382_));
INVX1 INVX1_2717 ( .A(u2__abc_52155_new_n11389_), .Y(u2__abc_52155_new_n11390_));
INVX1 INVX1_2718 ( .A(u2__abc_52155_new_n11400_), .Y(u2__abc_52155_new_n11401_));
INVX1 INVX1_2719 ( .A(u2__abc_52155_new_n11412_), .Y(u2__abc_52155_new_n11413_));
INVX1 INVX1_272 ( .A(sqrto_17_), .Y(u2__abc_52155_new_n3232_));
INVX1 INVX1_2720 ( .A(u2__abc_52155_new_n11420_), .Y(u2__abc_52155_new_n11421_));
INVX1 INVX1_2721 ( .A(u2__abc_52155_new_n4790_), .Y(u2__abc_52155_new_n11427_));
INVX1 INVX1_2722 ( .A(u2__abc_52155_new_n11428_), .Y(u2__abc_52155_new_n11429_));
INVX1 INVX1_2723 ( .A(u2__abc_52155_new_n11437_), .Y(u2__abc_52155_new_n11438_));
INVX1 INVX1_2724 ( .A(u2__abc_52155_new_n4769_), .Y(u2__abc_52155_new_n11444_));
INVX1 INVX1_2725 ( .A(u2__abc_52155_new_n11447_), .Y(u2__abc_52155_new_n11448_));
INVX1 INVX1_2726 ( .A(u2__abc_52155_new_n11455_), .Y(u2__abc_52155_new_n11456_));
INVX1 INVX1_2727 ( .A(u2__abc_52155_new_n4766_), .Y(u2__abc_52155_new_n11462_));
INVX1 INVX1_2728 ( .A(u2__abc_52155_new_n4774_), .Y(u2__abc_52155_new_n11465_));
INVX1 INVX1_2729 ( .A(u2__abc_52155_new_n11463_), .Y(u2__abc_52155_new_n11466_));
INVX1 INVX1_273 ( .A(u2_remHi_17_), .Y(u2__abc_52155_new_n3234_));
INVX1 INVX1_2730 ( .A(u2__abc_52155_new_n11473_), .Y(u2__abc_52155_new_n11474_));
INVX1 INVX1_2731 ( .A(u2__abc_52155_new_n11485_), .Y(u2__abc_52155_new_n11486_));
INVX1 INVX1_2732 ( .A(u2__abc_52155_new_n11489_), .Y(u2__abc_52155_new_n11490_));
INVX1 INVX1_2733 ( .A(u2__abc_52155_new_n11497_), .Y(u2__abc_52155_new_n11498_));
INVX1 INVX1_2734 ( .A(u2__abc_52155_new_n11504_), .Y(u2__abc_52155_new_n11505_));
INVX1 INVX1_2735 ( .A(u2__abc_52155_new_n11506_), .Y(u2__abc_52155_new_n11507_));
INVX1 INVX1_2736 ( .A(u2__abc_52155_new_n11514_), .Y(u2__abc_52155_new_n11515_));
INVX1 INVX1_2737 ( .A(u2__abc_52155_new_n11521_), .Y(u2__abc_52155_new_n11522_));
INVX1 INVX1_2738 ( .A(u2__abc_52155_new_n11523_), .Y(u2__abc_52155_new_n11524_));
INVX1 INVX1_2739 ( .A(u2__abc_52155_new_n11531_), .Y(u2__abc_52155_new_n11532_));
INVX1 INVX1_274 ( .A(u2__abc_52155_new_n3237_), .Y(u2__abc_52155_new_n3238_));
INVX1 INVX1_2740 ( .A(u2__abc_52155_new_n4747_), .Y(u2__abc_52155_new_n11540_));
INVX1 INVX1_2741 ( .A(u2__abc_52155_new_n11538_), .Y(u2__abc_52155_new_n11541_));
INVX1 INVX1_2742 ( .A(u2__abc_52155_new_n11548_), .Y(u2__abc_52155_new_n11549_));
INVX1 INVX1_2743 ( .A(u2__abc_52155_new_n11565_), .Y(u2__abc_52155_new_n11566_));
INVX1 INVX1_2744 ( .A(u2__abc_52155_new_n11573_), .Y(u2__abc_52155_new_n11574_));
INVX1 INVX1_2745 ( .A(u2__abc_52155_new_n4692_), .Y(u2__abc_52155_new_n11582_));
INVX1 INVX1_2746 ( .A(u2__abc_52155_new_n11580_), .Y(u2__abc_52155_new_n11583_));
INVX1 INVX1_2747 ( .A(u2__abc_52155_new_n11590_), .Y(u2__abc_52155_new_n11591_));
INVX1 INVX1_2748 ( .A(u2__abc_52155_new_n11599_), .Y(u2__abc_52155_new_n11600_));
INVX1 INVX1_2749 ( .A(u2__abc_52155_new_n11601_), .Y(u2__abc_52155_new_n11602_));
INVX1 INVX1_275 ( .A(sqrto_14_), .Y(u2__abc_52155_new_n3239_));
INVX1 INVX1_2750 ( .A(u2__abc_52155_new_n11609_), .Y(u2__abc_52155_new_n11610_));
INVX1 INVX1_2751 ( .A(u2__abc_52155_new_n4684_), .Y(u2__abc_52155_new_n11618_));
INVX1 INVX1_2752 ( .A(u2__abc_52155_new_n11616_), .Y(u2__abc_52155_new_n11619_));
INVX1 INVX1_2753 ( .A(u2__abc_52155_new_n11626_), .Y(u2__abc_52155_new_n11627_));
INVX1 INVX1_2754 ( .A(u2__abc_52155_new_n11633_), .Y(u2__abc_52155_new_n11634_));
INVX1 INVX1_2755 ( .A(u2__abc_52155_new_n11641_), .Y(u2__abc_52155_new_n11642_));
INVX1 INVX1_2756 ( .A(u2__abc_52155_new_n11649_), .Y(u2__abc_52155_new_n11650_));
INVX1 INVX1_2757 ( .A(u2__abc_52155_new_n4723_), .Y(u2__abc_52155_new_n11658_));
INVX1 INVX1_2758 ( .A(u2__abc_52155_new_n11656_), .Y(u2__abc_52155_new_n11659_));
INVX1 INVX1_2759 ( .A(u2__abc_52155_new_n11666_), .Y(u2__abc_52155_new_n11667_));
INVX1 INVX1_276 ( .A(u2__abc_52155_new_n3240_), .Y(u2__abc_52155_new_n3241_));
INVX1 INVX1_2760 ( .A(u2__abc_52155_new_n11675_), .Y(u2__abc_52155_new_n11676_));
INVX1 INVX1_2761 ( .A(u2__abc_52155_new_n11677_), .Y(u2__abc_52155_new_n11678_));
INVX1 INVX1_2762 ( .A(u2__abc_52155_new_n11685_), .Y(u2__abc_52155_new_n11686_));
INVX1 INVX1_2763 ( .A(u2__abc_52155_new_n4715_), .Y(u2__abc_52155_new_n11694_));
INVX1 INVX1_2764 ( .A(u2__abc_52155_new_n11692_), .Y(u2__abc_52155_new_n11695_));
INVX1 INVX1_2765 ( .A(u2__abc_52155_new_n11702_), .Y(u2__abc_52155_new_n11703_));
INVX1 INVX1_2766 ( .A(u2__abc_52155_new_n11711_), .Y(u2__abc_52155_new_n11712_));
INVX1 INVX1_2767 ( .A(u2__abc_52155_new_n11721_), .Y(u2__abc_52155_new_n11722_));
INVX1 INVX1_2768 ( .A(u2__abc_52155_new_n11729_), .Y(u2__abc_52155_new_n11730_));
INVX1 INVX1_2769 ( .A(u2__abc_52155_new_n4635_), .Y(u2__abc_52155_new_n11736_));
INVX1 INVX1_277 ( .A(sqrto_15_), .Y(u2__abc_52155_new_n3244_));
INVX1 INVX1_2770 ( .A(u2__abc_52155_new_n11737_), .Y(u2__abc_52155_new_n11738_));
INVX1 INVX1_2771 ( .A(u2__abc_52155_new_n11746_), .Y(u2__abc_52155_new_n11747_));
INVX1 INVX1_2772 ( .A(u2__abc_52155_new_n11754_), .Y(u2__abc_52155_new_n11755_));
INVX1 INVX1_2773 ( .A(u2__abc_52155_new_n11758_), .Y(u2__abc_52155_new_n11759_));
INVX1 INVX1_2774 ( .A(u2__abc_52155_new_n11766_), .Y(u2__abc_52155_new_n11767_));
INVX1 INVX1_2775 ( .A(u2__abc_52155_new_n4620_), .Y(u2__abc_52155_new_n11775_));
INVX1 INVX1_2776 ( .A(u2__abc_52155_new_n11773_), .Y(u2__abc_52155_new_n11776_));
INVX1 INVX1_2777 ( .A(u2__abc_52155_new_n11783_), .Y(u2__abc_52155_new_n11784_));
INVX1 INVX1_2778 ( .A(u2__abc_52155_new_n11796_), .Y(u2__abc_52155_new_n11797_));
INVX1 INVX1_2779 ( .A(u2__abc_52155_new_n11804_), .Y(u2__abc_52155_new_n11805_));
INVX1 INVX1_278 ( .A(u2__abc_52155_new_n3245_), .Y(u2__abc_52155_new_n3246_));
INVX1 INVX1_2780 ( .A(u2__abc_52155_new_n11811_), .Y(u2__abc_52155_new_n11812_));
INVX1 INVX1_2781 ( .A(u2__abc_52155_new_n11813_), .Y(u2__abc_52155_new_n11814_));
INVX1 INVX1_2782 ( .A(u2__abc_52155_new_n11821_), .Y(u2__abc_52155_new_n11822_));
INVX1 INVX1_2783 ( .A(u2__abc_52155_new_n11828_), .Y(u2__abc_52155_new_n11829_));
INVX1 INVX1_2784 ( .A(u2__abc_52155_new_n11830_), .Y(u2__abc_52155_new_n11831_));
INVX1 INVX1_2785 ( .A(u2__abc_52155_new_n11838_), .Y(u2__abc_52155_new_n11839_));
INVX1 INVX1_2786 ( .A(u2__abc_52155_new_n4651_), .Y(u2__abc_52155_new_n11847_));
INVX1 INVX1_2787 ( .A(u2__abc_52155_new_n11845_), .Y(u2__abc_52155_new_n11848_));
INVX1 INVX1_2788 ( .A(u2__abc_52155_new_n11855_), .Y(u2__abc_52155_new_n11856_));
INVX1 INVX1_2789 ( .A(u2__abc_52155_new_n11872_), .Y(u2__abc_52155_new_n11873_));
INVX1 INVX1_279 ( .A(u2_remHi_15_), .Y(u2__abc_52155_new_n3247_));
INVX1 INVX1_2790 ( .A(u2__abc_52155_new_n11880_), .Y(u2__abc_52155_new_n11881_));
INVX1 INVX1_2791 ( .A(u2__abc_52155_new_n4572_), .Y(u2__abc_52155_new_n11887_));
INVX1 INVX1_2792 ( .A(u2__abc_52155_new_n11888_), .Y(u2__abc_52155_new_n11889_));
INVX1 INVX1_2793 ( .A(u2__abc_52155_new_n11897_), .Y(u2__abc_52155_new_n11898_));
INVX1 INVX1_2794 ( .A(u2__abc_52155_new_n11905_), .Y(u2__abc_52155_new_n11906_));
INVX1 INVX1_2795 ( .A(u2__abc_52155_new_n11909_), .Y(u2__abc_52155_new_n11910_));
INVX1 INVX1_2796 ( .A(u2__abc_52155_new_n11917_), .Y(u2__abc_52155_new_n11918_));
INVX1 INVX1_2797 ( .A(u2__abc_52155_new_n4557_), .Y(u2__abc_52155_new_n11926_));
INVX1 INVX1_2798 ( .A(u2__abc_52155_new_n11924_), .Y(u2__abc_52155_new_n11927_));
INVX1 INVX1_2799 ( .A(u2__abc_52155_new_n11934_), .Y(u2__abc_52155_new_n11935_));
INVX1 INVX1_28 ( .A(\a[121] ), .Y(_abc_73687_new_n1601_));
INVX1 INVX1_280 ( .A(u2__abc_52155_new_n3248_), .Y(u2__abc_52155_new_n3249_));
INVX1 INVX1_2800 ( .A(u2__abc_52155_new_n11947_), .Y(u2__abc_52155_new_n11948_));
INVX1 INVX1_2801 ( .A(u2__abc_52155_new_n11955_), .Y(u2__abc_52155_new_n11956_));
INVX1 INVX1_2802 ( .A(u2__abc_52155_new_n4596_), .Y(u2__abc_52155_new_n11964_));
INVX1 INVX1_2803 ( .A(u2__abc_52155_new_n11962_), .Y(u2__abc_52155_new_n11965_));
INVX1 INVX1_2804 ( .A(u2__abc_52155_new_n11972_), .Y(u2__abc_52155_new_n11973_));
INVX1 INVX1_2805 ( .A(u2__abc_52155_new_n11981_), .Y(u2__abc_52155_new_n11982_));
INVX1 INVX1_2806 ( .A(u2__abc_52155_new_n11983_), .Y(u2__abc_52155_new_n11984_));
INVX1 INVX1_2807 ( .A(u2__abc_52155_new_n11991_), .Y(u2__abc_52155_new_n11992_));
INVX1 INVX1_2808 ( .A(u2__abc_52155_new_n4588_), .Y(u2__abc_52155_new_n12000_));
INVX1 INVX1_2809 ( .A(u2__abc_52155_new_n11998_), .Y(u2__abc_52155_new_n12001_));
INVX1 INVX1_281 ( .A(sqrto_20_), .Y(u2__abc_52155_new_n3253_));
INVX1 INVX1_2810 ( .A(u2__abc_52155_new_n12008_), .Y(u2__abc_52155_new_n12009_));
INVX1 INVX1_2811 ( .A(u2__abc_52155_new_n12015_), .Y(u2__abc_52155_new_n12016_));
INVX1 INVX1_2812 ( .A(u2__abc_52155_new_n12017_), .Y(u2__abc_52155_new_n12018_));
INVX1 INVX1_2813 ( .A(u2__abc_52155_new_n12019_), .Y(u2__abc_52155_new_n12020_));
INVX1 INVX1_2814 ( .A(u2__abc_52155_new_n12023_), .Y(u2__abc_52155_new_n12024_));
INVX1 INVX1_2815 ( .A(u2__abc_52155_new_n12025_), .Y(u2__abc_52155_new_n12026_));
INVX1 INVX1_2816 ( .A(u2__abc_52155_new_n12030_), .Y(u2__abc_52155_new_n12031_));
INVX1 INVX1_2817 ( .A(u2__abc_52155_new_n12034_), .Y(u2__abc_52155_new_n12035_));
INVX1 INVX1_2818 ( .A(u2__abc_52155_new_n12042_), .Y(u2__abc_52155_new_n12043_));
INVX1 INVX1_2819 ( .A(u2__abc_52155_new_n4500_), .Y(u2__abc_52155_new_n12051_));
INVX1 INVX1_282 ( .A(u2_remHi_20_), .Y(u2__abc_52155_new_n3255_));
INVX1 INVX1_2820 ( .A(u2__abc_52155_new_n12049_), .Y(u2__abc_52155_new_n12052_));
INVX1 INVX1_2821 ( .A(u2__abc_52155_new_n12059_), .Y(u2__abc_52155_new_n12060_));
INVX1 INVX1_2822 ( .A(u2__abc_52155_new_n12068_), .Y(u2__abc_52155_new_n12069_));
INVX1 INVX1_2823 ( .A(u2__abc_52155_new_n12070_), .Y(u2__abc_52155_new_n12071_));
INVX1 INVX1_2824 ( .A(u2__abc_52155_new_n12078_), .Y(u2__abc_52155_new_n12079_));
INVX1 INVX1_2825 ( .A(u2__abc_52155_new_n4492_), .Y(u2__abc_52155_new_n12087_));
INVX1 INVX1_2826 ( .A(u2__abc_52155_new_n12085_), .Y(u2__abc_52155_new_n12088_));
INVX1 INVX1_2827 ( .A(u2__abc_52155_new_n12095_), .Y(u2__abc_52155_new_n12096_));
INVX1 INVX1_2828 ( .A(u2__abc_52155_new_n12104_), .Y(u2__abc_52155_new_n12105_));
INVX1 INVX1_2829 ( .A(u2__abc_52155_new_n12106_), .Y(u2__abc_52155_new_n12107_));
INVX1 INVX1_283 ( .A(sqrto_21_), .Y(u2__abc_52155_new_n3258_));
INVX1 INVX1_2830 ( .A(u2__abc_52155_new_n12108_), .Y(u2__abc_52155_new_n12109_));
INVX1 INVX1_2831 ( .A(u2__abc_52155_new_n12112_), .Y(u2__abc_52155_new_n12113_));
INVX1 INVX1_2832 ( .A(u2__abc_52155_new_n12120_), .Y(u2__abc_52155_new_n12121_));
INVX1 INVX1_2833 ( .A(u2__abc_52155_new_n4531_), .Y(u2__abc_52155_new_n12129_));
INVX1 INVX1_2834 ( .A(u2__abc_52155_new_n12127_), .Y(u2__abc_52155_new_n12130_));
INVX1 INVX1_2835 ( .A(u2__abc_52155_new_n12137_), .Y(u2__abc_52155_new_n12138_));
INVX1 INVX1_2836 ( .A(u2__abc_52155_new_n12146_), .Y(u2__abc_52155_new_n12147_));
INVX1 INVX1_2837 ( .A(u2__abc_52155_new_n12148_), .Y(u2__abc_52155_new_n12149_));
INVX1 INVX1_2838 ( .A(u2__abc_52155_new_n12156_), .Y(u2__abc_52155_new_n12157_));
INVX1 INVX1_2839 ( .A(u2__abc_52155_new_n4523_), .Y(u2__abc_52155_new_n12165_));
INVX1 INVX1_284 ( .A(u2_remHi_21_), .Y(u2__abc_52155_new_n3260_));
INVX1 INVX1_2840 ( .A(u2__abc_52155_new_n12163_), .Y(u2__abc_52155_new_n12166_));
INVX1 INVX1_2841 ( .A(u2__abc_52155_new_n12173_), .Y(u2__abc_52155_new_n12174_));
INVX1 INVX1_2842 ( .A(u2__abc_52155_new_n12181_), .Y(u2__abc_52155_new_n12182_));
INVX1 INVX1_2843 ( .A(u2__abc_52155_new_n12190_), .Y(u2__abc_52155_new_n12191_));
INVX1 INVX1_2844 ( .A(u2__abc_52155_new_n12198_), .Y(u2__abc_52155_new_n12199_));
INVX1 INVX1_2845 ( .A(u2__abc_52155_new_n4468_), .Y(u2__abc_52155_new_n12205_));
INVX1 INVX1_2846 ( .A(u2__abc_52155_new_n12206_), .Y(u2__abc_52155_new_n12207_));
INVX1 INVX1_2847 ( .A(u2__abc_52155_new_n12215_), .Y(u2__abc_52155_new_n12216_));
INVX1 INVX1_2848 ( .A(u2__abc_52155_new_n12223_), .Y(u2__abc_52155_new_n12224_));
INVX1 INVX1_2849 ( .A(u2__abc_52155_new_n12227_), .Y(u2__abc_52155_new_n12228_));
INVX1 INVX1_285 ( .A(sqrto_19_), .Y(u2__abc_52155_new_n3264_));
INVX1 INVX1_2850 ( .A(u2__abc_52155_new_n12235_), .Y(u2__abc_52155_new_n12236_));
INVX1 INVX1_2851 ( .A(u2__abc_52155_new_n4460_), .Y(u2__abc_52155_new_n12244_));
INVX1 INVX1_2852 ( .A(u2__abc_52155_new_n12242_), .Y(u2__abc_52155_new_n12245_));
INVX1 INVX1_2853 ( .A(u2__abc_52155_new_n12252_), .Y(u2__abc_52155_new_n12253_));
INVX1 INVX1_2854 ( .A(u2__abc_52155_new_n12261_), .Y(u2__abc_52155_new_n12262_));
INVX1 INVX1_2855 ( .A(u2__abc_52155_new_n12263_), .Y(u2__abc_52155_new_n12264_));
INVX1 INVX1_2856 ( .A(u2__abc_52155_new_n12271_), .Y(u2__abc_52155_new_n12272_));
INVX1 INVX1_2857 ( .A(u2__abc_52155_new_n4437_), .Y(u2__abc_52155_new_n12280_));
INVX1 INVX1_2858 ( .A(u2__abc_52155_new_n12278_), .Y(u2__abc_52155_new_n12281_));
INVX1 INVX1_2859 ( .A(u2__abc_52155_new_n12288_), .Y(u2__abc_52155_new_n12289_));
INVX1 INVX1_286 ( .A(u2_remHi_19_), .Y(u2__abc_52155_new_n3266_));
INVX1 INVX1_2860 ( .A(u2__abc_52155_new_n12297_), .Y(u2__abc_52155_new_n12298_));
INVX1 INVX1_2861 ( .A(u2__abc_52155_new_n12299_), .Y(u2__abc_52155_new_n12300_));
INVX1 INVX1_2862 ( .A(u2__abc_52155_new_n12307_), .Y(u2__abc_52155_new_n12308_));
INVX1 INVX1_2863 ( .A(u2__abc_52155_new_n4429_), .Y(u2__abc_52155_new_n12316_));
INVX1 INVX1_2864 ( .A(u2__abc_52155_new_n12314_), .Y(u2__abc_52155_new_n12317_));
INVX1 INVX1_2865 ( .A(u2__abc_52155_new_n12324_), .Y(u2__abc_52155_new_n12325_));
INVX1 INVX1_2866 ( .A(u2__abc_52155_new_n12331_), .Y(u2__abc_52155_new_n12332_));
INVX1 INVX1_2867 ( .A(u2__abc_52155_new_n12334_), .Y(u2__abc_52155_new_n12335_));
INVX1 INVX1_2868 ( .A(u2__abc_52155_new_n12336_), .Y(u2__abc_52155_new_n12337_));
INVX1 INVX1_2869 ( .A(u2__abc_52155_new_n12338_), .Y(u2__abc_52155_new_n12339_));
INVX1 INVX1_287 ( .A(sqrto_18_), .Y(u2__abc_52155_new_n3269_));
INVX1 INVX1_2870 ( .A(u2__abc_52155_new_n12342_), .Y(u2__abc_52155_new_n12343_));
INVX1 INVX1_2871 ( .A(u2__abc_52155_new_n12344_), .Y(u2__abc_52155_new_n12345_));
INVX1 INVX1_2872 ( .A(u2__abc_52155_new_n12348_), .Y(u2__abc_52155_new_n12349_));
INVX1 INVX1_2873 ( .A(u2__abc_52155_new_n12352_), .Y(u2__abc_52155_new_n12353_));
INVX1 INVX1_2874 ( .A(u2__abc_52155_new_n12360_), .Y(u2__abc_52155_new_n12361_));
INVX1 INVX1_2875 ( .A(u2__abc_52155_new_n4365_), .Y(u2__abc_52155_new_n12369_));
INVX1 INVX1_2876 ( .A(u2__abc_52155_new_n12367_), .Y(u2__abc_52155_new_n12370_));
INVX1 INVX1_2877 ( .A(u2__abc_52155_new_n12377_), .Y(u2__abc_52155_new_n12378_));
INVX1 INVX1_2878 ( .A(u2__abc_52155_new_n12385_), .Y(u2__abc_52155_new_n12386_));
INVX1 INVX1_2879 ( .A(u2__abc_52155_new_n12389_), .Y(u2__abc_52155_new_n12390_));
INVX1 INVX1_288 ( .A(u2_remHi_18_), .Y(u2__abc_52155_new_n3271_));
INVX1 INVX1_2880 ( .A(u2__abc_52155_new_n12397_), .Y(u2__abc_52155_new_n12398_));
INVX1 INVX1_2881 ( .A(u2__abc_52155_new_n4380_), .Y(u2__abc_52155_new_n12406_));
INVX1 INVX1_2882 ( .A(u2__abc_52155_new_n12404_), .Y(u2__abc_52155_new_n12407_));
INVX1 INVX1_2883 ( .A(u2__abc_52155_new_n12414_), .Y(u2__abc_52155_new_n12415_));
INVX1 INVX1_2884 ( .A(u2__abc_52155_new_n12427_), .Y(u2__abc_52155_new_n12428_));
INVX1 INVX1_2885 ( .A(u2__abc_52155_new_n12435_), .Y(u2__abc_52155_new_n12436_));
INVX1 INVX1_2886 ( .A(u2__abc_52155_new_n12442_), .Y(u2__abc_52155_new_n12443_));
INVX1 INVX1_2887 ( .A(u2__abc_52155_new_n12444_), .Y(u2__abc_52155_new_n12445_));
INVX1 INVX1_2888 ( .A(u2__abc_52155_new_n12452_), .Y(u2__abc_52155_new_n12453_));
INVX1 INVX1_2889 ( .A(u2__abc_52155_new_n12459_), .Y(u2__abc_52155_new_n12460_));
INVX1 INVX1_289 ( .A(u2__abc_52155_new_n3275_), .Y(u2__abc_52155_new_n3276_));
INVX1 INVX1_2890 ( .A(u2__abc_52155_new_n12461_), .Y(u2__abc_52155_new_n12462_));
INVX1 INVX1_2891 ( .A(u2__abc_52155_new_n12469_), .Y(u2__abc_52155_new_n12470_));
INVX1 INVX1_2892 ( .A(u2__abc_52155_new_n4396_), .Y(u2__abc_52155_new_n12478_));
INVX1 INVX1_2893 ( .A(u2__abc_52155_new_n12476_), .Y(u2__abc_52155_new_n12479_));
INVX1 INVX1_2894 ( .A(u2__abc_52155_new_n12486_), .Y(u2__abc_52155_new_n12487_));
INVX1 INVX1_2895 ( .A(u2__abc_52155_new_n12503_), .Y(u2__abc_52155_new_n12504_));
INVX1 INVX1_2896 ( .A(u2__abc_52155_new_n12511_), .Y(u2__abc_52155_new_n12512_));
INVX1 INVX1_2897 ( .A(u2__abc_52155_new_n4302_), .Y(u2__abc_52155_new_n12520_));
INVX1 INVX1_2898 ( .A(u2__abc_52155_new_n12518_), .Y(u2__abc_52155_new_n12521_));
INVX1 INVX1_2899 ( .A(u2__abc_52155_new_n12528_), .Y(u2__abc_52155_new_n12529_));
INVX1 INVX1_29 ( .A(_abc_73687_new_n1588_), .Y(_abc_73687_new_n1602_));
INVX1 INVX1_290 ( .A(u2__abc_52155_new_n3278_), .Y(u2__abc_52155_new_n3279_));
INVX1 INVX1_2900 ( .A(u2__abc_52155_new_n12536_), .Y(u2__abc_52155_new_n12537_));
INVX1 INVX1_2901 ( .A(u2__abc_52155_new_n12540_), .Y(u2__abc_52155_new_n12541_));
INVX1 INVX1_2902 ( .A(u2__abc_52155_new_n12548_), .Y(u2__abc_52155_new_n12549_));
INVX1 INVX1_2903 ( .A(u2__abc_52155_new_n4317_), .Y(u2__abc_52155_new_n12557_));
INVX1 INVX1_2904 ( .A(u2__abc_52155_new_n12555_), .Y(u2__abc_52155_new_n12558_));
INVX1 INVX1_2905 ( .A(u2__abc_52155_new_n12565_), .Y(u2__abc_52155_new_n12566_));
INVX1 INVX1_2906 ( .A(u2__abc_52155_new_n12578_), .Y(u2__abc_52155_new_n12579_));
INVX1 INVX1_2907 ( .A(u2__abc_52155_new_n12586_), .Y(u2__abc_52155_new_n12587_));
INVX1 INVX1_2908 ( .A(u2__abc_52155_new_n4341_), .Y(u2__abc_52155_new_n12595_));
INVX1 INVX1_2909 ( .A(u2__abc_52155_new_n12593_), .Y(u2__abc_52155_new_n12596_));
INVX1 INVX1_291 ( .A(u2__abc_52155_new_n3226_), .Y(u2__abc_52155_new_n3281_));
INVX1 INVX1_2910 ( .A(u2__abc_52155_new_n12603_), .Y(u2__abc_52155_new_n12604_));
INVX1 INVX1_2911 ( .A(u2__abc_52155_new_n12612_), .Y(u2__abc_52155_new_n12613_));
INVX1 INVX1_2912 ( .A(u2__abc_52155_new_n12614_), .Y(u2__abc_52155_new_n12615_));
INVX1 INVX1_2913 ( .A(u2__abc_52155_new_n12622_), .Y(u2__abc_52155_new_n12623_));
INVX1 INVX1_2914 ( .A(u2__abc_52155_new_n4333_), .Y(u2__abc_52155_new_n12631_));
INVX1 INVX1_2915 ( .A(u2__abc_52155_new_n12629_), .Y(u2__abc_52155_new_n12632_));
INVX1 INVX1_2916 ( .A(u2__abc_52155_new_n12639_), .Y(u2__abc_52155_new_n12640_));
INVX1 INVX1_2917 ( .A(u2__abc_52155_new_n12652_), .Y(u2__abc_52155_new_n12653_));
INVX1 INVX1_2918 ( .A(u2__abc_52155_new_n12664_), .Y(u2__abc_52155_new_n12665_));
INVX1 INVX1_2919 ( .A(u2__abc_52155_new_n12672_), .Y(u2__abc_52155_new_n12673_));
INVX1 INVX1_292 ( .A(u2__abc_52155_new_n3235_), .Y(u2__abc_52155_new_n3285_));
INVX1 INVX1_2920 ( .A(u2__abc_52155_new_n6552_), .Y(u2__abc_52155_new_n12679_));
INVX1 INVX1_2921 ( .A(u2__abc_52155_new_n12680_), .Y(u2__abc_52155_new_n12682_));
INVX1 INVX1_2922 ( .A(u2__abc_52155_new_n12689_), .Y(u2__abc_52155_new_n12690_));
INVX1 INVX1_2923 ( .A(u2__abc_52155_new_n12697_), .Y(u2__abc_52155_new_n12698_));
INVX1 INVX1_2924 ( .A(u2__abc_52155_new_n12701_), .Y(u2__abc_52155_new_n12702_));
INVX1 INVX1_2925 ( .A(u2__abc_52155_new_n12709_), .Y(u2__abc_52155_new_n12710_));
INVX1 INVX1_2926 ( .A(u2__abc_52155_new_n6567_), .Y(u2__abc_52155_new_n12716_));
INVX1 INVX1_2927 ( .A(u2__abc_52155_new_n12717_), .Y(u2__abc_52155_new_n12719_));
INVX1 INVX1_2928 ( .A(u2__abc_52155_new_n12726_), .Y(u2__abc_52155_new_n12727_));
INVX1 INVX1_2929 ( .A(u2__abc_52155_new_n12739_), .Y(u2__abc_52155_new_n12740_));
INVX1 INVX1_293 ( .A(u2__abc_52155_new_n3230_), .Y(u2__abc_52155_new_n3286_));
INVX1 INVX1_2930 ( .A(u2__abc_52155_new_n12747_), .Y(u2__abc_52155_new_n12748_));
INVX1 INVX1_2931 ( .A(u2__abc_52155_new_n6598_), .Y(u2__abc_52155_new_n12756_));
INVX1 INVX1_2932 ( .A(u2__abc_52155_new_n12754_), .Y(u2__abc_52155_new_n12757_));
INVX1 INVX1_2933 ( .A(u2__abc_52155_new_n12764_), .Y(u2__abc_52155_new_n12765_));
INVX1 INVX1_2934 ( .A(u2__abc_52155_new_n12773_), .Y(u2__abc_52155_new_n12774_));
INVX1 INVX1_2935 ( .A(u2__abc_52155_new_n12775_), .Y(u2__abc_52155_new_n12776_));
INVX1 INVX1_2936 ( .A(u2__abc_52155_new_n12783_), .Y(u2__abc_52155_new_n12784_));
INVX1 INVX1_2937 ( .A(u2__abc_52155_new_n6583_), .Y(u2__abc_52155_new_n12790_));
INVX1 INVX1_2938 ( .A(u2__abc_52155_new_n12791_), .Y(u2__abc_52155_new_n12793_));
INVX1 INVX1_2939 ( .A(u2__abc_52155_new_n12800_), .Y(u2__abc_52155_new_n12801_));
INVX1 INVX1_294 ( .A(u2__abc_52155_new_n3267_), .Y(u2__abc_52155_new_n3291_));
INVX1 INVX1_2940 ( .A(u2__abc_52155_new_n12807_), .Y(u2__abc_52155_new_n12808_));
INVX1 INVX1_2941 ( .A(u2__abc_52155_new_n12812_), .Y(u2__abc_52155_new_n12813_));
INVX1 INVX1_2942 ( .A(u2__abc_52155_new_n12815_), .Y(u2__abc_52155_new_n12816_));
INVX1 INVX1_2943 ( .A(u2__abc_52155_new_n12819_), .Y(u2__abc_52155_new_n12820_));
INVX1 INVX1_2944 ( .A(u2__abc_52155_new_n12827_), .Y(u2__abc_52155_new_n12828_));
INVX1 INVX1_2945 ( .A(u2__abc_52155_new_n6535_), .Y(u2__abc_52155_new_n12834_));
INVX1 INVX1_2946 ( .A(u2__abc_52155_new_n12835_), .Y(u2__abc_52155_new_n12837_));
INVX1 INVX1_2947 ( .A(u2__abc_52155_new_n12844_), .Y(u2__abc_52155_new_n12845_));
INVX1 INVX1_2948 ( .A(u2__abc_52155_new_n12852_), .Y(u2__abc_52155_new_n12853_));
INVX1 INVX1_2949 ( .A(u2__abc_52155_new_n12856_), .Y(u2__abc_52155_new_n12857_));
INVX1 INVX1_295 ( .A(u2__abc_52155_new_n3272_), .Y(u2__abc_52155_new_n3292_));
INVX1 INVX1_2950 ( .A(u2__abc_52155_new_n12864_), .Y(u2__abc_52155_new_n12865_));
INVX1 INVX1_2951 ( .A(u2__abc_52155_new_n6520_), .Y(u2__abc_52155_new_n12871_));
INVX1 INVX1_2952 ( .A(u2__abc_52155_new_n12872_), .Y(u2__abc_52155_new_n12874_));
INVX1 INVX1_2953 ( .A(u2__abc_52155_new_n12881_), .Y(u2__abc_52155_new_n12882_));
INVX1 INVX1_2954 ( .A(u2__abc_52155_new_n12890_), .Y(u2__abc_52155_new_n12891_));
INVX1 INVX1_2955 ( .A(u2__abc_52155_new_n12892_), .Y(u2__abc_52155_new_n12893_));
INVX1 INVX1_2956 ( .A(u2__abc_52155_new_n12900_), .Y(u2__abc_52155_new_n12901_));
INVX1 INVX1_2957 ( .A(u2__abc_52155_new_n6504_), .Y(u2__abc_52155_new_n12909_));
INVX1 INVX1_2958 ( .A(u2__abc_52155_new_n12907_), .Y(u2__abc_52155_new_n12910_));
INVX1 INVX1_2959 ( .A(u2__abc_52155_new_n12917_), .Y(u2__abc_52155_new_n12918_));
INVX1 INVX1_296 ( .A(u2__abc_52155_new_n3259_), .Y(u2__abc_52155_new_n3296_));
INVX1 INVX1_2960 ( .A(u2__abc_52155_new_n12926_), .Y(u2__abc_52155_new_n12927_));
INVX1 INVX1_2961 ( .A(u2__abc_52155_new_n12928_), .Y(u2__abc_52155_new_n12929_));
INVX1 INVX1_2962 ( .A(u2__abc_52155_new_n12936_), .Y(u2__abc_52155_new_n12937_));
INVX1 INVX1_2963 ( .A(u2__abc_52155_new_n6489_), .Y(u2__abc_52155_new_n12943_));
INVX1 INVX1_2964 ( .A(u2__abc_52155_new_n12944_), .Y(u2__abc_52155_new_n12946_));
INVX1 INVX1_2965 ( .A(u2__abc_52155_new_n12953_), .Y(u2__abc_52155_new_n12954_));
INVX1 INVX1_2966 ( .A(u2__abc_52155_new_n12960_), .Y(u2__abc_52155_new_n12961_));
INVX1 INVX1_2967 ( .A(u2__abc_52155_new_n12963_), .Y(u2__abc_52155_new_n12964_));
INVX1 INVX1_2968 ( .A(u2__abc_52155_new_n12973_), .Y(u2__abc_52155_new_n12974_));
INVX1 INVX1_2969 ( .A(u2__abc_52155_new_n12977_), .Y(u2__abc_52155_new_n12978_));
INVX1 INVX1_297 ( .A(u2__abc_52155_new_n3298_), .Y(u2__abc_52155_new_n3299_));
INVX1 INVX1_2970 ( .A(u2__abc_52155_new_n12985_), .Y(u2__abc_52155_new_n12986_));
INVX1 INVX1_2971 ( .A(u2__abc_52155_new_n6440_), .Y(u2__abc_52155_new_n12994_));
INVX1 INVX1_2972 ( .A(u2__abc_52155_new_n12992_), .Y(u2__abc_52155_new_n12995_));
INVX1 INVX1_2973 ( .A(u2__abc_52155_new_n13002_), .Y(u2__abc_52155_new_n13003_));
INVX1 INVX1_2974 ( .A(u2__abc_52155_new_n13011_), .Y(u2__abc_52155_new_n13012_));
INVX1 INVX1_2975 ( .A(u2__abc_52155_new_n13013_), .Y(u2__abc_52155_new_n13014_));
INVX1 INVX1_2976 ( .A(u2__abc_52155_new_n13021_), .Y(u2__abc_52155_new_n13022_));
INVX1 INVX1_2977 ( .A(u2__abc_52155_new_n6425_), .Y(u2__abc_52155_new_n13028_));
INVX1 INVX1_2978 ( .A(u2__abc_52155_new_n13029_), .Y(u2__abc_52155_new_n13031_));
INVX1 INVX1_2979 ( .A(u2__abc_52155_new_n13038_), .Y(u2__abc_52155_new_n13039_));
INVX1 INVX1_298 ( .A(u2__abc_52155_new_n3225_), .Y(u2__abc_52155_new_n3303_));
INVX1 INVX1_2980 ( .A(u2__abc_52155_new_n13046_), .Y(u2__abc_52155_new_n13047_));
INVX1 INVX1_2981 ( .A(u2__abc_52155_new_n13050_), .Y(u2__abc_52155_new_n13051_));
INVX1 INVX1_2982 ( .A(u2__abc_52155_new_n13054_), .Y(u2__abc_52155_new_n13055_));
INVX1 INVX1_2983 ( .A(u2__abc_52155_new_n13062_), .Y(u2__abc_52155_new_n13063_));
INVX1 INVX1_2984 ( .A(u2__abc_52155_new_n6471_), .Y(u2__abc_52155_new_n13071_));
INVX1 INVX1_2985 ( .A(u2__abc_52155_new_n13069_), .Y(u2__abc_52155_new_n13072_));
INVX1 INVX1_2986 ( .A(u2__abc_52155_new_n13079_), .Y(u2__abc_52155_new_n13080_));
INVX1 INVX1_2987 ( .A(u2__abc_52155_new_n13088_), .Y(u2__abc_52155_new_n13089_));
INVX1 INVX1_2988 ( .A(u2__abc_52155_new_n13090_), .Y(u2__abc_52155_new_n13091_));
INVX1 INVX1_2989 ( .A(u2__abc_52155_new_n13098_), .Y(u2__abc_52155_new_n13099_));
INVX1 INVX1_299 ( .A(u2__abc_52155_new_n3173_), .Y(u2__abc_52155_new_n3307_));
INVX1 INVX1_2990 ( .A(u2__abc_52155_new_n6456_), .Y(u2__abc_52155_new_n13105_));
INVX1 INVX1_2991 ( .A(u2__abc_52155_new_n13106_), .Y(u2__abc_52155_new_n13108_));
INVX1 INVX1_2992 ( .A(u2__abc_52155_new_n13115_), .Y(u2__abc_52155_new_n13116_));
INVX1 INVX1_2993 ( .A(u2__abc_52155_new_n13122_), .Y(u2__abc_52155_new_n13123_));
INVX1 INVX1_2994 ( .A(u2__abc_52155_new_n13129_), .Y(u2__abc_52155_new_n13130_));
INVX1 INVX1_2995 ( .A(u2__abc_52155_new_n13133_), .Y(u2__abc_52155_new_n13134_));
INVX1 INVX1_2996 ( .A(u2__abc_52155_new_n13141_), .Y(u2__abc_52155_new_n13142_));
INVX1 INVX1_2997 ( .A(u2__abc_52155_new_n6377_), .Y(u2__abc_52155_new_n13150_));
INVX1 INVX1_2998 ( .A(u2__abc_52155_new_n13148_), .Y(u2__abc_52155_new_n13151_));
INVX1 INVX1_2999 ( .A(u2__abc_52155_new_n13158_), .Y(u2__abc_52155_new_n13159_));
INVX1 INVX1_3 ( .A(\a[113] ), .Y(_abc_73687_new_n1508_));
INVX1 INVX1_30 ( .A(_abc_73687_new_n1593_), .Y(_abc_73687_new_n1606_));
INVX1 INVX1_300 ( .A(u2__abc_52155_new_n3309_), .Y(u2__abc_52155_new_n3310_));
INVX1 INVX1_3000 ( .A(u2__abc_52155_new_n13167_), .Y(u2__abc_52155_new_n13168_));
INVX1 INVX1_3001 ( .A(u2__abc_52155_new_n13169_), .Y(u2__abc_52155_new_n13170_));
INVX1 INVX1_3002 ( .A(u2__abc_52155_new_n13177_), .Y(u2__abc_52155_new_n13178_));
INVX1 INVX1_3003 ( .A(u2__abc_52155_new_n6362_), .Y(u2__abc_52155_new_n13184_));
INVX1 INVX1_3004 ( .A(u2__abc_52155_new_n13185_), .Y(u2__abc_52155_new_n13187_));
INVX1 INVX1_3005 ( .A(u2__abc_52155_new_n13194_), .Y(u2__abc_52155_new_n13195_));
INVX1 INVX1_3006 ( .A(u2__abc_52155_new_n13204_), .Y(u2__abc_52155_new_n13205_));
INVX1 INVX1_3007 ( .A(u2__abc_52155_new_n13206_), .Y(u2__abc_52155_new_n13207_));
INVX1 INVX1_3008 ( .A(u2__abc_52155_new_n13210_), .Y(u2__abc_52155_new_n13211_));
INVX1 INVX1_3009 ( .A(u2__abc_52155_new_n13218_), .Y(u2__abc_52155_new_n13219_));
INVX1 INVX1_301 ( .A(u2__abc_52155_new_n3318_), .Y(u2__abc_52155_new_n3319_));
INVX1 INVX1_3010 ( .A(u2__abc_52155_new_n6408_), .Y(u2__abc_52155_new_n13227_));
INVX1 INVX1_3011 ( .A(u2__abc_52155_new_n13225_), .Y(u2__abc_52155_new_n13228_));
INVX1 INVX1_3012 ( .A(u2__abc_52155_new_n13235_), .Y(u2__abc_52155_new_n13236_));
INVX1 INVX1_3013 ( .A(u2__abc_52155_new_n13244_), .Y(u2__abc_52155_new_n13245_));
INVX1 INVX1_3014 ( .A(u2__abc_52155_new_n13246_), .Y(u2__abc_52155_new_n13247_));
INVX1 INVX1_3015 ( .A(u2__abc_52155_new_n13254_), .Y(u2__abc_52155_new_n13255_));
INVX1 INVX1_3016 ( .A(u2__abc_52155_new_n6393_), .Y(u2__abc_52155_new_n13261_));
INVX1 INVX1_3017 ( .A(u2__abc_52155_new_n13262_), .Y(u2__abc_52155_new_n13264_));
INVX1 INVX1_3018 ( .A(u2__abc_52155_new_n13271_), .Y(u2__abc_52155_new_n13272_));
INVX1 INVX1_3019 ( .A(u2__abc_52155_new_n13278_), .Y(u2__abc_52155_new_n13279_));
INVX1 INVX1_302 ( .A(sqrto_56_), .Y(u2__abc_52155_new_n3323_));
INVX1 INVX1_3020 ( .A(u2__abc_52155_new_n13280_), .Y(u2__abc_52155_new_n13281_));
INVX1 INVX1_3021 ( .A(u2__abc_52155_new_n13282_), .Y(u2__abc_52155_new_n13283_));
INVX1 INVX1_3022 ( .A(u2__abc_52155_new_n13287_), .Y(u2__abc_52155_new_n13288_));
INVX1 INVX1_3023 ( .A(u2__abc_52155_new_n13292_), .Y(u2__abc_52155_new_n13293_));
INVX1 INVX1_3024 ( .A(u2__abc_52155_new_n13296_), .Y(u2__abc_52155_new_n13297_));
INVX1 INVX1_3025 ( .A(u2__abc_52155_new_n13304_), .Y(u2__abc_52155_new_n13305_));
INVX1 INVX1_3026 ( .A(u2__abc_52155_new_n6312_), .Y(u2__abc_52155_new_n13313_));
INVX1 INVX1_3027 ( .A(u2__abc_52155_new_n13311_), .Y(u2__abc_52155_new_n13314_));
INVX1 INVX1_3028 ( .A(u2__abc_52155_new_n13321_), .Y(u2__abc_52155_new_n13322_));
INVX1 INVX1_3029 ( .A(u2__abc_52155_new_n13330_), .Y(u2__abc_52155_new_n13331_));
INVX1 INVX1_303 ( .A(u2__abc_52155_new_n3324_), .Y(u2__abc_52155_new_n3325_));
INVX1 INVX1_3030 ( .A(u2__abc_52155_new_n13332_), .Y(u2__abc_52155_new_n13333_));
INVX1 INVX1_3031 ( .A(u2__abc_52155_new_n13340_), .Y(u2__abc_52155_new_n13341_));
INVX1 INVX1_3032 ( .A(u2__abc_52155_new_n6297_), .Y(u2__abc_52155_new_n13347_));
INVX1 INVX1_3033 ( .A(u2__abc_52155_new_n13348_), .Y(u2__abc_52155_new_n13350_));
INVX1 INVX1_3034 ( .A(u2__abc_52155_new_n13357_), .Y(u2__abc_52155_new_n13358_));
INVX1 INVX1_3035 ( .A(u2__abc_52155_new_n13367_), .Y(u2__abc_52155_new_n13368_));
INVX1 INVX1_3036 ( .A(u2__abc_52155_new_n13369_), .Y(u2__abc_52155_new_n13370_));
INVX1 INVX1_3037 ( .A(u2__abc_52155_new_n13373_), .Y(u2__abc_52155_new_n13374_));
INVX1 INVX1_3038 ( .A(u2__abc_52155_new_n13381_), .Y(u2__abc_52155_new_n13382_));
INVX1 INVX1_3039 ( .A(u2__abc_52155_new_n6343_), .Y(u2__abc_52155_new_n13390_));
INVX1 INVX1_304 ( .A(u2_remHi_56_), .Y(u2__abc_52155_new_n3326_));
INVX1 INVX1_3040 ( .A(u2__abc_52155_new_n13388_), .Y(u2__abc_52155_new_n13391_));
INVX1 INVX1_3041 ( .A(u2__abc_52155_new_n13398_), .Y(u2__abc_52155_new_n13399_));
INVX1 INVX1_3042 ( .A(u2__abc_52155_new_n13407_), .Y(u2__abc_52155_new_n13408_));
INVX1 INVX1_3043 ( .A(u2__abc_52155_new_n13409_), .Y(u2__abc_52155_new_n13410_));
INVX1 INVX1_3044 ( .A(u2__abc_52155_new_n13417_), .Y(u2__abc_52155_new_n13418_));
INVX1 INVX1_3045 ( .A(u2__abc_52155_new_n6328_), .Y(u2__abc_52155_new_n13424_));
INVX1 INVX1_3046 ( .A(u2__abc_52155_new_n13425_), .Y(u2__abc_52155_new_n13427_));
INVX1 INVX1_3047 ( .A(u2__abc_52155_new_n13434_), .Y(u2__abc_52155_new_n13435_));
INVX1 INVX1_3048 ( .A(u2__abc_52155_new_n13441_), .Y(u2__abc_52155_new_n13442_));
INVX1 INVX1_3049 ( .A(u2__abc_52155_new_n13448_), .Y(u2__abc_52155_new_n13449_));
INVX1 INVX1_305 ( .A(u2__abc_52155_new_n3327_), .Y(u2__abc_52155_new_n3328_));
INVX1 INVX1_3050 ( .A(u2__abc_52155_new_n13452_), .Y(u2__abc_52155_new_n13453_));
INVX1 INVX1_3051 ( .A(u2__abc_52155_new_n13460_), .Y(u2__abc_52155_new_n13461_));
INVX1 INVX1_3052 ( .A(u2__abc_52155_new_n6234_), .Y(u2__abc_52155_new_n13467_));
INVX1 INVX1_3053 ( .A(u2__abc_52155_new_n13468_), .Y(u2__abc_52155_new_n13470_));
INVX1 INVX1_3054 ( .A(u2__abc_52155_new_n13477_), .Y(u2__abc_52155_new_n13478_));
INVX1 INVX1_3055 ( .A(u2__abc_52155_new_n13485_), .Y(u2__abc_52155_new_n13486_));
INVX1 INVX1_3056 ( .A(u2__abc_52155_new_n13489_), .Y(u2__abc_52155_new_n13490_));
INVX1 INVX1_3057 ( .A(u2__abc_52155_new_n13497_), .Y(u2__abc_52155_new_n13498_));
INVX1 INVX1_3058 ( .A(u2__abc_52155_new_n6249_), .Y(u2__abc_52155_new_n13504_));
INVX1 INVX1_3059 ( .A(u2__abc_52155_new_n13505_), .Y(u2__abc_52155_new_n13507_));
INVX1 INVX1_306 ( .A(sqrto_57_), .Y(u2__abc_52155_new_n3330_));
INVX1 INVX1_3060 ( .A(u2__abc_52155_new_n13514_), .Y(u2__abc_52155_new_n13515_));
INVX1 INVX1_3061 ( .A(u2__abc_52155_new_n13527_), .Y(u2__abc_52155_new_n13528_));
INVX1 INVX1_3062 ( .A(u2__abc_52155_new_n13535_), .Y(u2__abc_52155_new_n13536_));
INVX1 INVX1_3063 ( .A(u2__abc_52155_new_n6280_), .Y(u2__abc_52155_new_n13544_));
INVX1 INVX1_3064 ( .A(u2__abc_52155_new_n13542_), .Y(u2__abc_52155_new_n13545_));
INVX1 INVX1_3065 ( .A(u2__abc_52155_new_n13552_), .Y(u2__abc_52155_new_n13553_));
INVX1 INVX1_3066 ( .A(u2__abc_52155_new_n13561_), .Y(u2__abc_52155_new_n13562_));
INVX1 INVX1_3067 ( .A(u2__abc_52155_new_n13563_), .Y(u2__abc_52155_new_n13564_));
INVX1 INVX1_3068 ( .A(u2__abc_52155_new_n13571_), .Y(u2__abc_52155_new_n13572_));
INVX1 INVX1_3069 ( .A(u2__abc_52155_new_n6265_), .Y(u2__abc_52155_new_n13578_));
INVX1 INVX1_307 ( .A(u2__abc_52155_new_n3331_), .Y(u2__abc_52155_new_n3332_));
INVX1 INVX1_3070 ( .A(u2__abc_52155_new_n13579_), .Y(u2__abc_52155_new_n13581_));
INVX1 INVX1_3071 ( .A(u2__abc_52155_new_n13588_), .Y(u2__abc_52155_new_n13589_));
INVX1 INVX1_3072 ( .A(u2__abc_52155_new_n13595_), .Y(u2__abc_52155_new_n13596_));
INVX1 INVX1_3073 ( .A(u2__abc_52155_new_n13597_), .Y(u2__abc_52155_new_n13598_));
INVX1 INVX1_3074 ( .A(u2__abc_52155_new_n13602_), .Y(u2__abc_52155_new_n13603_));
INVX1 INVX1_3075 ( .A(u2__abc_52155_new_n13606_), .Y(u2__abc_52155_new_n13607_));
INVX1 INVX1_3076 ( .A(u2__abc_52155_new_n13610_), .Y(u2__abc_52155_new_n13611_));
INVX1 INVX1_3077 ( .A(u2__abc_52155_new_n13618_), .Y(u2__abc_52155_new_n13619_));
INVX1 INVX1_3078 ( .A(u2__abc_52155_new_n6170_), .Y(u2__abc_52155_new_n13625_));
INVX1 INVX1_3079 ( .A(u2__abc_52155_new_n13626_), .Y(u2__abc_52155_new_n13628_));
INVX1 INVX1_308 ( .A(u2_remHi_57_), .Y(u2__abc_52155_new_n3333_));
INVX1 INVX1_3080 ( .A(u2__abc_52155_new_n13635_), .Y(u2__abc_52155_new_n13636_));
INVX1 INVX1_3081 ( .A(u2__abc_52155_new_n13643_), .Y(u2__abc_52155_new_n13644_));
INVX1 INVX1_3082 ( .A(u2__abc_52155_new_n13647_), .Y(u2__abc_52155_new_n13648_));
INVX1 INVX1_3083 ( .A(u2__abc_52155_new_n13655_), .Y(u2__abc_52155_new_n13656_));
INVX1 INVX1_3084 ( .A(u2__abc_52155_new_n6185_), .Y(u2__abc_52155_new_n13662_));
INVX1 INVX1_3085 ( .A(u2__abc_52155_new_n13663_), .Y(u2__abc_52155_new_n13665_));
INVX1 INVX1_3086 ( .A(u2__abc_52155_new_n13672_), .Y(u2__abc_52155_new_n13673_));
INVX1 INVX1_3087 ( .A(u2__abc_52155_new_n13685_), .Y(u2__abc_52155_new_n13686_));
INVX1 INVX1_3088 ( .A(u2__abc_52155_new_n13693_), .Y(u2__abc_52155_new_n13694_));
INVX1 INVX1_3089 ( .A(u2__abc_52155_new_n13700_), .Y(u2__abc_52155_new_n13701_));
INVX1 INVX1_309 ( .A(u2__abc_52155_new_n3334_), .Y(u2__abc_52155_new_n3335_));
INVX1 INVX1_3090 ( .A(u2__abc_52155_new_n13702_), .Y(u2__abc_52155_new_n13703_));
INVX1 INVX1_3091 ( .A(u2__abc_52155_new_n13710_), .Y(u2__abc_52155_new_n13711_));
INVX1 INVX1_3092 ( .A(u2__abc_52155_new_n13717_), .Y(u2__abc_52155_new_n13718_));
INVX1 INVX1_3093 ( .A(u2__abc_52155_new_n13719_), .Y(u2__abc_52155_new_n13720_));
INVX1 INVX1_3094 ( .A(u2__abc_52155_new_n13727_), .Y(u2__abc_52155_new_n13728_));
INVX1 INVX1_3095 ( .A(u2__abc_52155_new_n6201_), .Y(u2__abc_52155_new_n13734_));
INVX1 INVX1_3096 ( .A(u2__abc_52155_new_n13735_), .Y(u2__abc_52155_new_n13737_));
INVX1 INVX1_3097 ( .A(u2__abc_52155_new_n13744_), .Y(u2__abc_52155_new_n13745_));
INVX1 INVX1_3098 ( .A(u2__abc_52155_new_n13761_), .Y(u2__abc_52155_new_n13762_));
INVX1 INVX1_3099 ( .A(u2__abc_52155_new_n13769_), .Y(u2__abc_52155_new_n13770_));
INVX1 INVX1_31 ( .A(_abc_73687_new_n1604_), .Y(_abc_73687_new_n1607_));
INVX1 INVX1_310 ( .A(sqrto_54_), .Y(u2__abc_52155_new_n3338_));
INVX1 INVX1_3100 ( .A(u2__abc_52155_new_n6122_), .Y(u2__abc_52155_new_n13778_));
INVX1 INVX1_3101 ( .A(u2__abc_52155_new_n13776_), .Y(u2__abc_52155_new_n13779_));
INVX1 INVX1_3102 ( .A(u2__abc_52155_new_n13786_), .Y(u2__abc_52155_new_n13787_));
INVX1 INVX1_3103 ( .A(u2__abc_52155_new_n13795_), .Y(u2__abc_52155_new_n13796_));
INVX1 INVX1_3104 ( .A(u2__abc_52155_new_n13797_), .Y(u2__abc_52155_new_n13798_));
INVX1 INVX1_3105 ( .A(u2__abc_52155_new_n13805_), .Y(u2__abc_52155_new_n13806_));
INVX1 INVX1_3106 ( .A(u2__abc_52155_new_n6107_), .Y(u2__abc_52155_new_n13812_));
INVX1 INVX1_3107 ( .A(u2__abc_52155_new_n13813_), .Y(u2__abc_52155_new_n13815_));
INVX1 INVX1_3108 ( .A(u2__abc_52155_new_n13822_), .Y(u2__abc_52155_new_n13823_));
INVX1 INVX1_3109 ( .A(u2__abc_52155_new_n6108_), .Y(u2__abc_52155_new_n13829_));
INVX1 INVX1_311 ( .A(u2__abc_52155_new_n3339_), .Y(u2__abc_52155_new_n3340_));
INVX1 INVX1_3110 ( .A(u2__abc_52155_new_n13833_), .Y(u2__abc_52155_new_n13834_));
INVX1 INVX1_3111 ( .A(u2__abc_52155_new_n13835_), .Y(u2__abc_52155_new_n13836_));
INVX1 INVX1_3112 ( .A(u2__abc_52155_new_n13839_), .Y(u2__abc_52155_new_n13840_));
INVX1 INVX1_3113 ( .A(u2__abc_52155_new_n13847_), .Y(u2__abc_52155_new_n13848_));
INVX1 INVX1_3114 ( .A(u2__abc_52155_new_n6153_), .Y(u2__abc_52155_new_n13856_));
INVX1 INVX1_3115 ( .A(u2__abc_52155_new_n13854_), .Y(u2__abc_52155_new_n13857_));
INVX1 INVX1_3116 ( .A(u2__abc_52155_new_n13864_), .Y(u2__abc_52155_new_n13865_));
INVX1 INVX1_3117 ( .A(u2__abc_52155_new_n13873_), .Y(u2__abc_52155_new_n13874_));
INVX1 INVX1_3118 ( .A(u2__abc_52155_new_n13875_), .Y(u2__abc_52155_new_n13876_));
INVX1 INVX1_3119 ( .A(u2__abc_52155_new_n13883_), .Y(u2__abc_52155_new_n13884_));
INVX1 INVX1_312 ( .A(u2_remHi_54_), .Y(u2__abc_52155_new_n3341_));
INVX1 INVX1_3120 ( .A(u2__abc_52155_new_n6138_), .Y(u2__abc_52155_new_n13890_));
INVX1 INVX1_3121 ( .A(u2__abc_52155_new_n13891_), .Y(u2__abc_52155_new_n13893_));
INVX1 INVX1_3122 ( .A(u2__abc_52155_new_n13900_), .Y(u2__abc_52155_new_n13901_));
INVX1 INVX1_3123 ( .A(u2__abc_52155_new_n13907_), .Y(u2__abc_52155_new_n13908_));
INVX1 INVX1_3124 ( .A(u2__abc_52155_new_n13909_), .Y(u2__abc_52155_new_n13910_));
INVX1 INVX1_3125 ( .A(u2__abc_52155_new_n13911_), .Y(u2__abc_52155_new_n13912_));
INVX1 INVX1_3126 ( .A(u2__abc_52155_new_n13913_), .Y(u2__abc_52155_new_n13914_));
INVX1 INVX1_3127 ( .A(u2__abc_52155_new_n6139_), .Y(u2__abc_52155_new_n13915_));
INVX1 INVX1_3128 ( .A(u2__abc_52155_new_n13919_), .Y(u2__abc_52155_new_n13920_));
INVX1 INVX1_3129 ( .A(u2__abc_52155_new_n13925_), .Y(u2__abc_52155_new_n13926_));
INVX1 INVX1_313 ( .A(u2__abc_52155_new_n3342_), .Y(u2__abc_52155_new_n3343_));
INVX1 INVX1_3130 ( .A(u2__abc_52155_new_n13929_), .Y(u2__abc_52155_new_n13930_));
INVX1 INVX1_3131 ( .A(u2__abc_52155_new_n13937_), .Y(u2__abc_52155_new_n13938_));
INVX1 INVX1_3132 ( .A(u2__abc_52155_new_n6072_), .Y(u2__abc_52155_new_n13944_));
INVX1 INVX1_3133 ( .A(u2__abc_52155_new_n13945_), .Y(u2__abc_52155_new_n13947_));
INVX1 INVX1_3134 ( .A(u2__abc_52155_new_n13954_), .Y(u2__abc_52155_new_n13955_));
INVX1 INVX1_3135 ( .A(u2__abc_52155_new_n13962_), .Y(u2__abc_52155_new_n13963_));
INVX1 INVX1_3136 ( .A(u2__abc_52155_new_n13966_), .Y(u2__abc_52155_new_n13967_));
INVX1 INVX1_3137 ( .A(u2__abc_52155_new_n13974_), .Y(u2__abc_52155_new_n13975_));
INVX1 INVX1_3138 ( .A(u2__abc_52155_new_n6087_), .Y(u2__abc_52155_new_n13981_));
INVX1 INVX1_3139 ( .A(u2__abc_52155_new_n13982_), .Y(u2__abc_52155_new_n13984_));
INVX1 INVX1_314 ( .A(sqrto_55_), .Y(u2__abc_52155_new_n3345_));
INVX1 INVX1_3140 ( .A(u2__abc_52155_new_n13991_), .Y(u2__abc_52155_new_n13992_));
INVX1 INVX1_3141 ( .A(u2__abc_52155_new_n14004_), .Y(u2__abc_52155_new_n14005_));
INVX1 INVX1_3142 ( .A(u2__abc_52155_new_n14012_), .Y(u2__abc_52155_new_n14013_));
INVX1 INVX1_3143 ( .A(u2__abc_52155_new_n6056_), .Y(u2__abc_52155_new_n14021_));
INVX1 INVX1_3144 ( .A(u2__abc_52155_new_n14019_), .Y(u2__abc_52155_new_n14022_));
INVX1 INVX1_3145 ( .A(u2__abc_52155_new_n14029_), .Y(u2__abc_52155_new_n14030_));
INVX1 INVX1_3146 ( .A(u2__abc_52155_new_n14038_), .Y(u2__abc_52155_new_n14039_));
INVX1 INVX1_3147 ( .A(u2__abc_52155_new_n14040_), .Y(u2__abc_52155_new_n14041_));
INVX1 INVX1_3148 ( .A(u2__abc_52155_new_n14048_), .Y(u2__abc_52155_new_n14049_));
INVX1 INVX1_3149 ( .A(u2__abc_52155_new_n6041_), .Y(u2__abc_52155_new_n14055_));
INVX1 INVX1_315 ( .A(u2__abc_52155_new_n3346_), .Y(u2__abc_52155_new_n3347_));
INVX1 INVX1_3150 ( .A(u2__abc_52155_new_n14056_), .Y(u2__abc_52155_new_n14058_));
INVX1 INVX1_3151 ( .A(u2__abc_52155_new_n14065_), .Y(u2__abc_52155_new_n14066_));
INVX1 INVX1_3152 ( .A(u2__abc_52155_new_n14072_), .Y(u2__abc_52155_new_n14073_));
INVX1 INVX1_3153 ( .A(u2__abc_52155_new_n14079_), .Y(u2__abc_52155_new_n14080_));
INVX1 INVX1_3154 ( .A(u2__abc_52155_new_n14083_), .Y(u2__abc_52155_new_n14084_));
INVX1 INVX1_3155 ( .A(u2__abc_52155_new_n14091_), .Y(u2__abc_52155_new_n14092_));
INVX1 INVX1_3156 ( .A(u2__abc_52155_new_n5978_), .Y(u2__abc_52155_new_n14098_));
INVX1 INVX1_3157 ( .A(u2__abc_52155_new_n14099_), .Y(u2__abc_52155_new_n14101_));
INVX1 INVX1_3158 ( .A(u2__abc_52155_new_n14108_), .Y(u2__abc_52155_new_n14109_));
INVX1 INVX1_3159 ( .A(u2__abc_52155_new_n14116_), .Y(u2__abc_52155_new_n14117_));
INVX1 INVX1_316 ( .A(u2_remHi_55_), .Y(u2__abc_52155_new_n3348_));
INVX1 INVX1_3160 ( .A(u2__abc_52155_new_n14120_), .Y(u2__abc_52155_new_n14121_));
INVX1 INVX1_3161 ( .A(u2__abc_52155_new_n14128_), .Y(u2__abc_52155_new_n14129_));
INVX1 INVX1_3162 ( .A(u2__abc_52155_new_n5993_), .Y(u2__abc_52155_new_n14135_));
INVX1 INVX1_3163 ( .A(u2__abc_52155_new_n14136_), .Y(u2__abc_52155_new_n14138_));
INVX1 INVX1_3164 ( .A(u2__abc_52155_new_n14145_), .Y(u2__abc_52155_new_n14146_));
INVX1 INVX1_3165 ( .A(u2__abc_52155_new_n14158_), .Y(u2__abc_52155_new_n14159_));
INVX1 INVX1_3166 ( .A(u2__abc_52155_new_n14166_), .Y(u2__abc_52155_new_n14167_));
INVX1 INVX1_3167 ( .A(u2__abc_52155_new_n6024_), .Y(u2__abc_52155_new_n14175_));
INVX1 INVX1_3168 ( .A(u2__abc_52155_new_n14173_), .Y(u2__abc_52155_new_n14176_));
INVX1 INVX1_3169 ( .A(u2__abc_52155_new_n14183_), .Y(u2__abc_52155_new_n14184_));
INVX1 INVX1_317 ( .A(u2__abc_52155_new_n3349_), .Y(u2__abc_52155_new_n3350_));
INVX1 INVX1_3170 ( .A(u2__abc_52155_new_n14192_), .Y(u2__abc_52155_new_n14193_));
INVX1 INVX1_3171 ( .A(u2__abc_52155_new_n14194_), .Y(u2__abc_52155_new_n14195_));
INVX1 INVX1_3172 ( .A(u2__abc_52155_new_n14202_), .Y(u2__abc_52155_new_n14203_));
INVX1 INVX1_3173 ( .A(u2__abc_52155_new_n6009_), .Y(u2__abc_52155_new_n14209_));
INVX1 INVX1_3174 ( .A(u2__abc_52155_new_n14210_), .Y(u2__abc_52155_new_n14212_));
INVX1 INVX1_3175 ( .A(u2__abc_52155_new_n14219_), .Y(u2__abc_52155_new_n14220_));
INVX1 INVX1_3176 ( .A(u2__abc_52155_new_n14226_), .Y(u2__abc_52155_new_n14227_));
INVX1 INVX1_3177 ( .A(u2__abc_52155_new_n14228_), .Y(u2__abc_52155_new_n14229_));
INVX1 INVX1_3178 ( .A(u2__abc_52155_new_n14233_), .Y(u2__abc_52155_new_n14234_));
INVX1 INVX1_3179 ( .A(u2__abc_52155_new_n14237_), .Y(u2__abc_52155_new_n14238_));
INVX1 INVX1_318 ( .A(sqrto_60_), .Y(u2__abc_52155_new_n3354_));
INVX1 INVX1_3180 ( .A(u2__abc_52155_new_n14241_), .Y(u2__abc_52155_new_n14242_));
INVX1 INVX1_3181 ( .A(u2__abc_52155_new_n14249_), .Y(u2__abc_52155_new_n14250_));
INVX1 INVX1_3182 ( .A(u2__abc_52155_new_n5929_), .Y(u2__abc_52155_new_n14258_));
INVX1 INVX1_3183 ( .A(u2__abc_52155_new_n14256_), .Y(u2__abc_52155_new_n14259_));
INVX1 INVX1_3184 ( .A(u2__abc_52155_new_n14266_), .Y(u2__abc_52155_new_n14267_));
INVX1 INVX1_3185 ( .A(u2__abc_52155_new_n14275_), .Y(u2__abc_52155_new_n14276_));
INVX1 INVX1_3186 ( .A(u2__abc_52155_new_n14277_), .Y(u2__abc_52155_new_n14278_));
INVX1 INVX1_3187 ( .A(u2__abc_52155_new_n14285_), .Y(u2__abc_52155_new_n14286_));
INVX1 INVX1_3188 ( .A(u2__abc_52155_new_n5914_), .Y(u2__abc_52155_new_n14292_));
INVX1 INVX1_3189 ( .A(u2__abc_52155_new_n14293_), .Y(u2__abc_52155_new_n14295_));
INVX1 INVX1_319 ( .A(u2__abc_52155_new_n3355_), .Y(u2__abc_52155_new_n3356_));
INVX1 INVX1_3190 ( .A(u2__abc_52155_new_n14302_), .Y(u2__abc_52155_new_n14303_));
INVX1 INVX1_3191 ( .A(u2__abc_52155_new_n14312_), .Y(u2__abc_52155_new_n14313_));
INVX1 INVX1_3192 ( .A(u2__abc_52155_new_n14314_), .Y(u2__abc_52155_new_n14315_));
INVX1 INVX1_3193 ( .A(u2__abc_52155_new_n14318_), .Y(u2__abc_52155_new_n14319_));
INVX1 INVX1_3194 ( .A(u2__abc_52155_new_n14326_), .Y(u2__abc_52155_new_n14327_));
INVX1 INVX1_3195 ( .A(u2__abc_52155_new_n5960_), .Y(u2__abc_52155_new_n14335_));
INVX1 INVX1_3196 ( .A(u2__abc_52155_new_n14333_), .Y(u2__abc_52155_new_n14336_));
INVX1 INVX1_3197 ( .A(u2__abc_52155_new_n14343_), .Y(u2__abc_52155_new_n14344_));
INVX1 INVX1_3198 ( .A(u2__abc_52155_new_n14352_), .Y(u2__abc_52155_new_n14353_));
INVX1 INVX1_3199 ( .A(u2__abc_52155_new_n14354_), .Y(u2__abc_52155_new_n14355_));
INVX1 INVX1_32 ( .A(\a[122] ), .Y(_abc_73687_new_n1615_));
INVX1 INVX1_320 ( .A(u2_remHi_60_), .Y(u2__abc_52155_new_n3357_));
INVX1 INVX1_3200 ( .A(u2__abc_52155_new_n14362_), .Y(u2__abc_52155_new_n14363_));
INVX1 INVX1_3201 ( .A(u2__abc_52155_new_n5945_), .Y(u2__abc_52155_new_n14369_));
INVX1 INVX1_3202 ( .A(u2__abc_52155_new_n14370_), .Y(u2__abc_52155_new_n14372_));
INVX1 INVX1_3203 ( .A(u2__abc_52155_new_n14379_), .Y(u2__abc_52155_new_n14380_));
INVX1 INVX1_3204 ( .A(u2__abc_52155_new_n14386_), .Y(u2__abc_52155_new_n14387_));
INVX1 INVX1_3205 ( .A(u2__abc_52155_new_n14391_), .Y(u2__abc_52155_new_n14392_));
INVX1 INVX1_3206 ( .A(u2__abc_52155_new_n14394_), .Y(u2__abc_52155_new_n14395_));
INVX1 INVX1_3207 ( .A(u2__abc_52155_new_n14398_), .Y(u2__abc_52155_new_n14399_));
INVX1 INVX1_3208 ( .A(u2__abc_52155_new_n14406_), .Y(u2__abc_52155_new_n14407_));
INVX1 INVX1_3209 ( .A(u2__abc_52155_new_n5866_), .Y(u2__abc_52155_new_n14415_));
INVX1 INVX1_321 ( .A(u2__abc_52155_new_n3358_), .Y(u2__abc_52155_new_n3359_));
INVX1 INVX1_3210 ( .A(u2__abc_52155_new_n14413_), .Y(u2__abc_52155_new_n14416_));
INVX1 INVX1_3211 ( .A(u2__abc_52155_new_n14423_), .Y(u2__abc_52155_new_n14424_));
INVX1 INVX1_3212 ( .A(u2__abc_52155_new_n14432_), .Y(u2__abc_52155_new_n14433_));
INVX1 INVX1_3213 ( .A(u2__abc_52155_new_n14434_), .Y(u2__abc_52155_new_n14435_));
INVX1 INVX1_3214 ( .A(u2__abc_52155_new_n14442_), .Y(u2__abc_52155_new_n14443_));
INVX1 INVX1_3215 ( .A(u2__abc_52155_new_n5851_), .Y(u2__abc_52155_new_n14449_));
INVX1 INVX1_3216 ( .A(u2__abc_52155_new_n14450_), .Y(u2__abc_52155_new_n14452_));
INVX1 INVX1_3217 ( .A(u2__abc_52155_new_n14459_), .Y(u2__abc_52155_new_n14460_));
INVX1 INVX1_3218 ( .A(u2__abc_52155_new_n14469_), .Y(u2__abc_52155_new_n14470_));
INVX1 INVX1_3219 ( .A(u2__abc_52155_new_n14471_), .Y(u2__abc_52155_new_n14472_));
INVX1 INVX1_322 ( .A(u2_remHi_61_), .Y(u2__abc_52155_new_n3361_));
INVX1 INVX1_3220 ( .A(u2__abc_52155_new_n14475_), .Y(u2__abc_52155_new_n14476_));
INVX1 INVX1_3221 ( .A(u2__abc_52155_new_n14483_), .Y(u2__abc_52155_new_n14484_));
INVX1 INVX1_3222 ( .A(u2__abc_52155_new_n5897_), .Y(u2__abc_52155_new_n14492_));
INVX1 INVX1_3223 ( .A(u2__abc_52155_new_n14490_), .Y(u2__abc_52155_new_n14493_));
INVX1 INVX1_3224 ( .A(u2__abc_52155_new_n14500_), .Y(u2__abc_52155_new_n14501_));
INVX1 INVX1_3225 ( .A(u2__abc_52155_new_n14509_), .Y(u2__abc_52155_new_n14510_));
INVX1 INVX1_3226 ( .A(u2__abc_52155_new_n14511_), .Y(u2__abc_52155_new_n14512_));
INVX1 INVX1_3227 ( .A(u2__abc_52155_new_n14519_), .Y(u2__abc_52155_new_n14520_));
INVX1 INVX1_3228 ( .A(u2__abc_52155_new_n5882_), .Y(u2__abc_52155_new_n14526_));
INVX1 INVX1_3229 ( .A(u2__abc_52155_new_n14527_), .Y(u2__abc_52155_new_n14529_));
INVX1 INVX1_323 ( .A(u2__abc_52155_new_n3362_), .Y(u2__abc_52155_new_n3363_));
INVX1 INVX1_3230 ( .A(u2__abc_52155_new_n14536_), .Y(u2__abc_52155_new_n14537_));
INVX1 INVX1_3231 ( .A(u2__abc_52155_new_n14543_), .Y(u2__abc_52155_new_n14544_));
INVX1 INVX1_3232 ( .A(u2__abc_52155_new_n14545_), .Y(u2__abc_52155_new_n14546_));
INVX1 INVX1_3233 ( .A(u2__abc_52155_new_n14547_), .Y(u2__abc_52155_new_n14548_));
INVX1 INVX1_3234 ( .A(u2__abc_52155_new_n14552_), .Y(u2__abc_52155_new_n14553_));
INVX1 INVX1_3235 ( .A(u2__abc_52155_new_n14557_), .Y(u2__abc_52155_new_n14558_));
INVX1 INVX1_3236 ( .A(u2__abc_52155_new_n14561_), .Y(u2__abc_52155_new_n14562_));
INVX1 INVX1_3237 ( .A(u2__abc_52155_new_n14569_), .Y(u2__abc_52155_new_n14570_));
INVX1 INVX1_3238 ( .A(u2__abc_52155_new_n5801_), .Y(u2__abc_52155_new_n14578_));
INVX1 INVX1_3239 ( .A(u2__abc_52155_new_n14576_), .Y(u2__abc_52155_new_n14579_));
INVX1 INVX1_324 ( .A(sqrto_61_), .Y(u2__abc_52155_new_n3364_));
INVX1 INVX1_3240 ( .A(u2__abc_52155_new_n14586_), .Y(u2__abc_52155_new_n14587_));
INVX1 INVX1_3241 ( .A(u2__abc_52155_new_n14595_), .Y(u2__abc_52155_new_n14596_));
INVX1 INVX1_3242 ( .A(u2__abc_52155_new_n14597_), .Y(u2__abc_52155_new_n14598_));
INVX1 INVX1_3243 ( .A(u2__abc_52155_new_n14605_), .Y(u2__abc_52155_new_n14606_));
INVX1 INVX1_3244 ( .A(u2__abc_52155_new_n5786_), .Y(u2__abc_52155_new_n14612_));
INVX1 INVX1_3245 ( .A(u2__abc_52155_new_n14613_), .Y(u2__abc_52155_new_n14615_));
INVX1 INVX1_3246 ( .A(u2__abc_52155_new_n14622_), .Y(u2__abc_52155_new_n14623_));
INVX1 INVX1_3247 ( .A(u2__abc_52155_new_n14632_), .Y(u2__abc_52155_new_n14633_));
INVX1 INVX1_3248 ( .A(u2__abc_52155_new_n14634_), .Y(u2__abc_52155_new_n14635_));
INVX1 INVX1_3249 ( .A(u2__abc_52155_new_n14638_), .Y(u2__abc_52155_new_n14639_));
INVX1 INVX1_325 ( .A(u2__abc_52155_new_n3365_), .Y(u2__abc_52155_new_n3366_));
INVX1 INVX1_3250 ( .A(u2__abc_52155_new_n14646_), .Y(u2__abc_52155_new_n14647_));
INVX1 INVX1_3251 ( .A(u2__abc_52155_new_n5832_), .Y(u2__abc_52155_new_n14655_));
INVX1 INVX1_3252 ( .A(u2__abc_52155_new_n14653_), .Y(u2__abc_52155_new_n14656_));
INVX1 INVX1_3253 ( .A(u2__abc_52155_new_n14663_), .Y(u2__abc_52155_new_n14664_));
INVX1 INVX1_3254 ( .A(u2__abc_52155_new_n14672_), .Y(u2__abc_52155_new_n14673_));
INVX1 INVX1_3255 ( .A(u2__abc_52155_new_n14674_), .Y(u2__abc_52155_new_n14675_));
INVX1 INVX1_3256 ( .A(u2__abc_52155_new_n14682_), .Y(u2__abc_52155_new_n14683_));
INVX1 INVX1_3257 ( .A(u2__abc_52155_new_n5817_), .Y(u2__abc_52155_new_n14689_));
INVX1 INVX1_3258 ( .A(u2__abc_52155_new_n14690_), .Y(u2__abc_52155_new_n14692_));
INVX1 INVX1_3259 ( .A(u2__abc_52155_new_n14699_), .Y(u2__abc_52155_new_n14700_));
INVX1 INVX1_326 ( .A(sqrto_59_), .Y(u2__abc_52155_new_n3369_));
INVX1 INVX1_3260 ( .A(u2__abc_52155_new_n14706_), .Y(u2__abc_52155_new_n14707_));
INVX1 INVX1_3261 ( .A(u2__abc_52155_new_n5818_), .Y(u2__abc_52155_new_n14708_));
INVX1 INVX1_3262 ( .A(u2__abc_52155_new_n14714_), .Y(u2__abc_52155_new_n14715_));
INVX1 INVX1_3263 ( .A(u2__abc_52155_new_n14718_), .Y(u2__abc_52155_new_n14719_));
INVX1 INVX1_3264 ( .A(u2__abc_52155_new_n14726_), .Y(u2__abc_52155_new_n14727_));
INVX1 INVX1_3265 ( .A(u2__abc_52155_new_n5723_), .Y(u2__abc_52155_new_n14733_));
INVX1 INVX1_3266 ( .A(u2__abc_52155_new_n14734_), .Y(u2__abc_52155_new_n14736_));
INVX1 INVX1_3267 ( .A(u2__abc_52155_new_n14743_), .Y(u2__abc_52155_new_n14744_));
INVX1 INVX1_3268 ( .A(u2__abc_52155_new_n14751_), .Y(u2__abc_52155_new_n14752_));
INVX1 INVX1_3269 ( .A(u2__abc_52155_new_n14755_), .Y(u2__abc_52155_new_n14756_));
INVX1 INVX1_327 ( .A(u2__abc_52155_new_n3370_), .Y(u2__abc_52155_new_n3371_));
INVX1 INVX1_3270 ( .A(u2__abc_52155_new_n14763_), .Y(u2__abc_52155_new_n14764_));
INVX1 INVX1_3271 ( .A(u2__abc_52155_new_n5738_), .Y(u2__abc_52155_new_n14770_));
INVX1 INVX1_3272 ( .A(u2__abc_52155_new_n14771_), .Y(u2__abc_52155_new_n14773_));
INVX1 INVX1_3273 ( .A(u2__abc_52155_new_n14780_), .Y(u2__abc_52155_new_n14781_));
INVX1 INVX1_3274 ( .A(u2__abc_52155_new_n14793_), .Y(u2__abc_52155_new_n14794_));
INVX1 INVX1_3275 ( .A(u2__abc_52155_new_n14801_), .Y(u2__abc_52155_new_n14802_));
INVX1 INVX1_3276 ( .A(u2__abc_52155_new_n5769_), .Y(u2__abc_52155_new_n14810_));
INVX1 INVX1_3277 ( .A(u2__abc_52155_new_n14808_), .Y(u2__abc_52155_new_n14811_));
INVX1 INVX1_3278 ( .A(u2__abc_52155_new_n14818_), .Y(u2__abc_52155_new_n14819_));
INVX1 INVX1_3279 ( .A(u2__abc_52155_new_n14827_), .Y(u2__abc_52155_new_n14828_));
INVX1 INVX1_328 ( .A(u2_remHi_59_), .Y(u2__abc_52155_new_n3372_));
INVX1 INVX1_3280 ( .A(u2__abc_52155_new_n14829_), .Y(u2__abc_52155_new_n14830_));
INVX1 INVX1_3281 ( .A(u2__abc_52155_new_n14837_), .Y(u2__abc_52155_new_n14838_));
INVX1 INVX1_3282 ( .A(u2__abc_52155_new_n5754_), .Y(u2__abc_52155_new_n14844_));
INVX1 INVX1_3283 ( .A(u2__abc_52155_new_n14845_), .Y(u2__abc_52155_new_n14847_));
INVX1 INVX1_3284 ( .A(u2__abc_52155_new_n14854_), .Y(u2__abc_52155_new_n14855_));
INVX1 INVX1_3285 ( .A(u2__abc_52155_new_n14861_), .Y(u2__abc_52155_new_n14862_));
INVX1 INVX1_3286 ( .A(u2__abc_52155_new_n14863_), .Y(u2__abc_52155_new_n14864_));
INVX1 INVX1_3287 ( .A(u2__abc_52155_new_n5755_), .Y(u2__abc_52155_new_n14865_));
INVX1 INVX1_3288 ( .A(u2__abc_52155_new_n14869_), .Y(u2__abc_52155_new_n14870_));
INVX1 INVX1_3289 ( .A(u2__abc_52155_new_n14873_), .Y(u2__abc_52155_new_n14874_));
INVX1 INVX1_329 ( .A(u2__abc_52155_new_n3373_), .Y(u2__abc_52155_new_n3374_));
INVX1 INVX1_3290 ( .A(u2__abc_52155_new_n14877_), .Y(u2__abc_52155_new_n14878_));
INVX1 INVX1_3291 ( .A(u2__abc_52155_new_n14885_), .Y(u2__abc_52155_new_n14886_));
INVX1 INVX1_3292 ( .A(u2__abc_52155_new_n5674_), .Y(u2__abc_52155_new_n14894_));
INVX1 INVX1_3293 ( .A(u2__abc_52155_new_n14892_), .Y(u2__abc_52155_new_n14895_));
INVX1 INVX1_3294 ( .A(u2__abc_52155_new_n14902_), .Y(u2__abc_52155_new_n14903_));
INVX1 INVX1_3295 ( .A(u2__abc_52155_new_n14911_), .Y(u2__abc_52155_new_n14912_));
INVX1 INVX1_3296 ( .A(u2__abc_52155_new_n14913_), .Y(u2__abc_52155_new_n14914_));
INVX1 INVX1_3297 ( .A(u2__abc_52155_new_n14921_), .Y(u2__abc_52155_new_n14922_));
INVX1 INVX1_3298 ( .A(u2__abc_52155_new_n5659_), .Y(u2__abc_52155_new_n14928_));
INVX1 INVX1_3299 ( .A(u2__abc_52155_new_n14929_), .Y(u2__abc_52155_new_n14931_));
INVX1 INVX1_33 ( .A(_abc_73687_new_n1600_), .Y(_abc_73687_new_n1616_));
INVX1 INVX1_330 ( .A(sqrto_58_), .Y(u2__abc_52155_new_n3376_));
INVX1 INVX1_3300 ( .A(u2__abc_52155_new_n14938_), .Y(u2__abc_52155_new_n14939_));
INVX1 INVX1_3301 ( .A(u2__abc_52155_new_n14946_), .Y(u2__abc_52155_new_n14947_));
INVX1 INVX1_3302 ( .A(u2__abc_52155_new_n14950_), .Y(u2__abc_52155_new_n14951_));
INVX1 INVX1_3303 ( .A(u2__abc_52155_new_n14954_), .Y(u2__abc_52155_new_n14955_));
INVX1 INVX1_3304 ( .A(u2__abc_52155_new_n14962_), .Y(u2__abc_52155_new_n14963_));
INVX1 INVX1_3305 ( .A(u2__abc_52155_new_n14969_), .Y(u2__abc_52155_new_n14970_));
INVX1 INVX1_3306 ( .A(u2__abc_52155_new_n14971_), .Y(u2__abc_52155_new_n14972_));
INVX1 INVX1_3307 ( .A(u2__abc_52155_new_n14979_), .Y(u2__abc_52155_new_n14980_));
INVX1 INVX1_3308 ( .A(u2__abc_52155_new_n14986_), .Y(u2__abc_52155_new_n14987_));
INVX1 INVX1_3309 ( .A(u2__abc_52155_new_n14988_), .Y(u2__abc_52155_new_n14989_));
INVX1 INVX1_331 ( .A(u2__abc_52155_new_n3377_), .Y(u2__abc_52155_new_n3378_));
INVX1 INVX1_3310 ( .A(u2__abc_52155_new_n14996_), .Y(u2__abc_52155_new_n14997_));
INVX1 INVX1_3311 ( .A(u2__abc_52155_new_n5690_), .Y(u2__abc_52155_new_n15003_));
INVX1 INVX1_3312 ( .A(u2__abc_52155_new_n15004_), .Y(u2__abc_52155_new_n15006_));
INVX1 INVX1_3313 ( .A(u2__abc_52155_new_n15013_), .Y(u2__abc_52155_new_n15014_));
INVX1 INVX1_3314 ( .A(u2__abc_52155_new_n15030_), .Y(u2__abc_52155_new_n15031_));
INVX1 INVX1_3315 ( .A(u2__abc_52155_new_n15038_), .Y(u2__abc_52155_new_n15039_));
INVX1 INVX1_3316 ( .A(u2__abc_52155_new_n5627_), .Y(u2__abc_52155_new_n15045_));
INVX1 INVX1_3317 ( .A(u2__abc_52155_new_n15046_), .Y(u2__abc_52155_new_n15048_));
INVX1 INVX1_3318 ( .A(u2__abc_52155_new_n15055_), .Y(u2__abc_52155_new_n15056_));
INVX1 INVX1_3319 ( .A(u2__abc_52155_new_n15063_), .Y(u2__abc_52155_new_n15064_));
INVX1 INVX1_332 ( .A(u2_remHi_58_), .Y(u2__abc_52155_new_n3379_));
INVX1 INVX1_3320 ( .A(u2__abc_52155_new_n15067_), .Y(u2__abc_52155_new_n15068_));
INVX1 INVX1_3321 ( .A(u2__abc_52155_new_n15075_), .Y(u2__abc_52155_new_n15076_));
INVX1 INVX1_3322 ( .A(u2__abc_52155_new_n5642_), .Y(u2__abc_52155_new_n15082_));
INVX1 INVX1_3323 ( .A(u2__abc_52155_new_n15083_), .Y(u2__abc_52155_new_n15085_));
INVX1 INVX1_3324 ( .A(u2__abc_52155_new_n15092_), .Y(u2__abc_52155_new_n15093_));
INVX1 INVX1_3325 ( .A(u2__abc_52155_new_n15103_), .Y(u2__abc_52155_new_n15104_));
INVX1 INVX1_3326 ( .A(u2__abc_52155_new_n15111_), .Y(u2__abc_52155_new_n15112_));
INVX1 INVX1_3327 ( .A(u2__abc_52155_new_n5611_), .Y(u2__abc_52155_new_n15120_));
INVX1 INVX1_3328 ( .A(u2__abc_52155_new_n15118_), .Y(u2__abc_52155_new_n15121_));
INVX1 INVX1_3329 ( .A(u2__abc_52155_new_n15128_), .Y(u2__abc_52155_new_n15129_));
INVX1 INVX1_333 ( .A(u2__abc_52155_new_n3380_), .Y(u2__abc_52155_new_n3381_));
INVX1 INVX1_3330 ( .A(u2__abc_52155_new_n15137_), .Y(u2__abc_52155_new_n15138_));
INVX1 INVX1_3331 ( .A(u2__abc_52155_new_n15139_), .Y(u2__abc_52155_new_n15140_));
INVX1 INVX1_3332 ( .A(u2__abc_52155_new_n15147_), .Y(u2__abc_52155_new_n15148_));
INVX1 INVX1_3333 ( .A(u2__abc_52155_new_n5596_), .Y(u2__abc_52155_new_n15154_));
INVX1 INVX1_3334 ( .A(u2__abc_52155_new_n15155_), .Y(u2__abc_52155_new_n15157_));
INVX1 INVX1_3335 ( .A(u2__abc_52155_new_n15164_), .Y(u2__abc_52155_new_n15165_));
INVX1 INVX1_3336 ( .A(u2__abc_52155_new_n15171_), .Y(u2__abc_52155_new_n15172_));
INVX1 INVX1_3337 ( .A(u2__abc_52155_new_n15173_), .Y(u2__abc_52155_new_n15174_));
INVX1 INVX1_3338 ( .A(u2__abc_52155_new_n15175_), .Y(u2__abc_52155_new_n15176_));
INVX1 INVX1_3339 ( .A(u2__abc_52155_new_n15177_), .Y(u2__abc_52155_new_n15178_));
INVX1 INVX1_334 ( .A(sqrto_48_), .Y(u2__abc_52155_new_n3386_));
INVX1 INVX1_3340 ( .A(u2__abc_52155_new_n15179_), .Y(u2__abc_52155_new_n15180_));
INVX1 INVX1_3341 ( .A(u2__abc_52155_new_n15183_), .Y(u2__abc_52155_new_n15184_));
INVX1 INVX1_3342 ( .A(u2__abc_52155_new_n15188_), .Y(u2__abc_52155_new_n15189_));
INVX1 INVX1_3343 ( .A(u2__abc_52155_new_n15196_), .Y(u2__abc_52155_new_n15197_));
INVX1 INVX1_3344 ( .A(u2__abc_52155_new_n15198_), .Y(u2__abc_52155_new_n15199_));
INVX1 INVX1_3345 ( .A(u2__abc_52155_new_n15206_), .Y(u2__abc_52155_new_n15207_));
INVX1 INVX1_3346 ( .A(u2__abc_52155_new_n7234_), .Y(u2__abc_52155_new_n15213_));
INVX1 INVX1_3347 ( .A(u2__abc_52155_new_n15214_), .Y(u2__abc_52155_new_n15216_));
INVX1 INVX1_3348 ( .A(u2__abc_52155_new_n15223_), .Y(u2__abc_52155_new_n15224_));
INVX1 INVX1_3349 ( .A(u2__abc_52155_new_n15232_), .Y(u2__abc_52155_new_n15233_));
INVX1 INVX1_335 ( .A(u2_remHi_48_), .Y(u2__abc_52155_new_n3388_));
INVX1 INVX1_3350 ( .A(u2__abc_52155_new_n15234_), .Y(u2__abc_52155_new_n15235_));
INVX1 INVX1_3351 ( .A(u2__abc_52155_new_n15242_), .Y(u2__abc_52155_new_n15243_));
INVX1 INVX1_3352 ( .A(u2__abc_52155_new_n7226_), .Y(u2__abc_52155_new_n15249_));
INVX1 INVX1_3353 ( .A(u2__abc_52155_new_n15250_), .Y(u2__abc_52155_new_n15252_));
INVX1 INVX1_3354 ( .A(u2__abc_52155_new_n15259_), .Y(u2__abc_52155_new_n15260_));
INVX1 INVX1_3355 ( .A(u2__abc_52155_new_n15266_), .Y(u2__abc_52155_new_n15267_));
INVX1 INVX1_3356 ( .A(u2__abc_52155_new_n15274_), .Y(u2__abc_52155_new_n15275_));
INVX1 INVX1_3357 ( .A(u2__abc_52155_new_n15282_), .Y(u2__abc_52155_new_n15283_));
INVX1 INVX1_3358 ( .A(u2__abc_52155_new_n7203_), .Y(u2__abc_52155_new_n15291_));
INVX1 INVX1_3359 ( .A(u2__abc_52155_new_n15289_), .Y(u2__abc_52155_new_n15292_));
INVX1 INVX1_336 ( .A(sqrto_49_), .Y(u2__abc_52155_new_n3391_));
INVX1 INVX1_3360 ( .A(u2__abc_52155_new_n15299_), .Y(u2__abc_52155_new_n15300_));
INVX1 INVX1_3361 ( .A(u2__abc_52155_new_n15308_), .Y(u2__abc_52155_new_n15309_));
INVX1 INVX1_3362 ( .A(u2__abc_52155_new_n15310_), .Y(u2__abc_52155_new_n15311_));
INVX1 INVX1_3363 ( .A(u2__abc_52155_new_n15318_), .Y(u2__abc_52155_new_n15319_));
INVX1 INVX1_3364 ( .A(u2__abc_52155_new_n7195_), .Y(u2__abc_52155_new_n15325_));
INVX1 INVX1_3365 ( .A(u2__abc_52155_new_n15326_), .Y(u2__abc_52155_new_n15328_));
INVX1 INVX1_3366 ( .A(u2__abc_52155_new_n15335_), .Y(u2__abc_52155_new_n15336_));
INVX1 INVX1_3367 ( .A(u2__abc_52155_new_n15343_), .Y(u2__abc_52155_new_n15344_));
INVX1 INVX1_3368 ( .A(u2__abc_52155_new_n15352_), .Y(u2__abc_52155_new_n15353_));
INVX1 INVX1_3369 ( .A(u2__abc_52155_new_n15360_), .Y(u2__abc_52155_new_n15361_));
INVX1 INVX1_337 ( .A(u2_remHi_49_), .Y(u2__abc_52155_new_n3393_));
INVX1 INVX1_3370 ( .A(u2__abc_52155_new_n7400_), .Y(u2__abc_52155_new_n15367_));
INVX1 INVX1_3371 ( .A(u2__abc_52155_new_n15368_), .Y(u2__abc_52155_new_n15369_));
INVX1 INVX1_3372 ( .A(u2__abc_52155_new_n15377_), .Y(u2__abc_52155_new_n15378_));
INVX1 INVX1_3373 ( .A(u2__abc_52155_new_n15386_), .Y(u2__abc_52155_new_n15387_));
INVX1 INVX1_3374 ( .A(u2__abc_52155_new_n15394_), .Y(u2__abc_52155_new_n15395_));
INVX1 INVX1_3375 ( .A(u2__abc_52155_new_n7385_), .Y(u2__abc_52155_new_n15401_));
INVX1 INVX1_3376 ( .A(u2__abc_52155_new_n15402_), .Y(u2__abc_52155_new_n15404_));
INVX1 INVX1_3377 ( .A(u2__abc_52155_new_n15411_), .Y(u2__abc_52155_new_n15412_));
INVX1 INVX1_3378 ( .A(u2__abc_52155_new_n15419_), .Y(u2__abc_52155_new_n15420_));
INVX1 INVX1_3379 ( .A(u2__abc_52155_new_n15427_), .Y(u2__abc_52155_new_n15428_));
INVX1 INVX1_338 ( .A(u2__abc_52155_new_n3396_), .Y(u2__abc_52155_new_n3397_));
INVX1 INVX1_3380 ( .A(u2__abc_52155_new_n15435_), .Y(u2__abc_52155_new_n15436_));
INVX1 INVX1_3381 ( .A(u2__abc_52155_new_n7424_), .Y(u2__abc_52155_new_n15444_));
INVX1 INVX1_3382 ( .A(u2__abc_52155_new_n15442_), .Y(u2__abc_52155_new_n15445_));
INVX1 INVX1_3383 ( .A(u2__abc_52155_new_n15452_), .Y(u2__abc_52155_new_n15453_));
INVX1 INVX1_3384 ( .A(u2__abc_52155_new_n15461_), .Y(u2__abc_52155_new_n15462_));
INVX1 INVX1_3385 ( .A(u2__abc_52155_new_n15463_), .Y(u2__abc_52155_new_n15464_));
INVX1 INVX1_3386 ( .A(u2__abc_52155_new_n15471_), .Y(u2__abc_52155_new_n15472_));
INVX1 INVX1_3387 ( .A(u2__abc_52155_new_n7416_), .Y(u2__abc_52155_new_n15478_));
INVX1 INVX1_3388 ( .A(u2__abc_52155_new_n15479_), .Y(u2__abc_52155_new_n15481_));
INVX1 INVX1_3389 ( .A(u2__abc_52155_new_n15488_), .Y(u2__abc_52155_new_n15489_));
INVX1 INVX1_339 ( .A(sqrto_47_), .Y(u2__abc_52155_new_n3398_));
INVX1 INVX1_3390 ( .A(u2__abc_52155_new_n15496_), .Y(u2__abc_52155_new_n15497_));
INVX1 INVX1_3391 ( .A(u2__abc_52155_new_n15505_), .Y(u2__abc_52155_new_n15506_));
INVX1 INVX1_3392 ( .A(u2__abc_52155_new_n15513_), .Y(u2__abc_52155_new_n15514_));
INVX1 INVX1_3393 ( .A(u2__abc_52155_new_n7321_), .Y(u2__abc_52155_new_n15520_));
INVX1 INVX1_3394 ( .A(u2__abc_52155_new_n15521_), .Y(u2__abc_52155_new_n15523_));
INVX1 INVX1_3395 ( .A(u2__abc_52155_new_n15530_), .Y(u2__abc_52155_new_n15531_));
INVX1 INVX1_3396 ( .A(u2__abc_52155_new_n15538_), .Y(u2__abc_52155_new_n15539_));
INVX1 INVX1_3397 ( .A(u2__abc_52155_new_n15542_), .Y(u2__abc_52155_new_n15543_));
INVX1 INVX1_3398 ( .A(u2__abc_52155_new_n15550_), .Y(u2__abc_52155_new_n15551_));
INVX1 INVX1_3399 ( .A(u2__abc_52155_new_n7336_), .Y(u2__abc_52155_new_n15557_));
INVX1 INVX1_34 ( .A(_abc_73687_new_n1605_), .Y(_abc_73687_new_n1620_));
INVX1 INVX1_340 ( .A(u2__abc_52155_new_n3399_), .Y(u2__abc_52155_new_n3400_));
INVX1 INVX1_3400 ( .A(u2__abc_52155_new_n15558_), .Y(u2__abc_52155_new_n15560_));
INVX1 INVX1_3401 ( .A(u2__abc_52155_new_n15567_), .Y(u2__abc_52155_new_n15568_));
INVX1 INVX1_3402 ( .A(u2__abc_52155_new_n15580_), .Y(u2__abc_52155_new_n15581_));
INVX1 INVX1_3403 ( .A(u2__abc_52155_new_n15588_), .Y(u2__abc_52155_new_n15589_));
INVX1 INVX1_3404 ( .A(u2__abc_52155_new_n7360_), .Y(u2__abc_52155_new_n15597_));
INVX1 INVX1_3405 ( .A(u2__abc_52155_new_n15595_), .Y(u2__abc_52155_new_n15598_));
INVX1 INVX1_3406 ( .A(u2__abc_52155_new_n15605_), .Y(u2__abc_52155_new_n15606_));
INVX1 INVX1_3407 ( .A(u2__abc_52155_new_n15614_), .Y(u2__abc_52155_new_n15615_));
INVX1 INVX1_3408 ( .A(u2__abc_52155_new_n15616_), .Y(u2__abc_52155_new_n15617_));
INVX1 INVX1_3409 ( .A(u2__abc_52155_new_n15624_), .Y(u2__abc_52155_new_n15625_));
INVX1 INVX1_341 ( .A(u2_remHi_47_), .Y(u2__abc_52155_new_n3401_));
INVX1 INVX1_3410 ( .A(u2__abc_52155_new_n7352_), .Y(u2__abc_52155_new_n15631_));
INVX1 INVX1_3411 ( .A(u2__abc_52155_new_n15632_), .Y(u2__abc_52155_new_n15634_));
INVX1 INVX1_3412 ( .A(u2__abc_52155_new_n15641_), .Y(u2__abc_52155_new_n15642_));
INVX1 INVX1_3413 ( .A(u2__abc_52155_new_n15649_), .Y(u2__abc_52155_new_n15650_));
INVX1 INVX1_3414 ( .A(u2__abc_52155_new_n15658_), .Y(u2__abc_52155_new_n15659_));
INVX1 INVX1_3415 ( .A(u2__abc_52155_new_n15666_), .Y(u2__abc_52155_new_n15667_));
INVX1 INVX1_3416 ( .A(u2__abc_52155_new_n7266_), .Y(u2__abc_52155_new_n15675_));
INVX1 INVX1_3417 ( .A(u2__abc_52155_new_n15673_), .Y(u2__abc_52155_new_n15676_));
INVX1 INVX1_3418 ( .A(u2__abc_52155_new_n15683_), .Y(u2__abc_52155_new_n15684_));
INVX1 INVX1_3419 ( .A(u2__abc_52155_new_n15692_), .Y(u2__abc_52155_new_n15693_));
INVX1 INVX1_342 ( .A(u2__abc_52155_new_n3402_), .Y(u2__abc_52155_new_n3403_));
INVX1 INVX1_3420 ( .A(u2__abc_52155_new_n15694_), .Y(u2__abc_52155_new_n15695_));
INVX1 INVX1_3421 ( .A(u2__abc_52155_new_n15702_), .Y(u2__abc_52155_new_n15703_));
INVX1 INVX1_3422 ( .A(u2__abc_52155_new_n7258_), .Y(u2__abc_52155_new_n15709_));
INVX1 INVX1_3423 ( .A(u2__abc_52155_new_n15710_), .Y(u2__abc_52155_new_n15712_));
INVX1 INVX1_3424 ( .A(u2__abc_52155_new_n15719_), .Y(u2__abc_52155_new_n15720_));
INVX1 INVX1_3425 ( .A(u2__abc_52155_new_n15726_), .Y(u2__abc_52155_new_n15727_));
INVX1 INVX1_3426 ( .A(u2__abc_52155_new_n15734_), .Y(u2__abc_52155_new_n15735_));
INVX1 INVX1_3427 ( .A(u2__abc_52155_new_n15742_), .Y(u2__abc_52155_new_n15743_));
INVX1 INVX1_3428 ( .A(u2__abc_52155_new_n7297_), .Y(u2__abc_52155_new_n15751_));
INVX1 INVX1_3429 ( .A(u2__abc_52155_new_n15749_), .Y(u2__abc_52155_new_n15752_));
INVX1 INVX1_343 ( .A(sqrto_46_), .Y(u2__abc_52155_new_n3405_));
INVX1 INVX1_3430 ( .A(u2__abc_52155_new_n15759_), .Y(u2__abc_52155_new_n15760_));
INVX1 INVX1_3431 ( .A(u2__abc_52155_new_n15768_), .Y(u2__abc_52155_new_n15769_));
INVX1 INVX1_3432 ( .A(u2__abc_52155_new_n15770_), .Y(u2__abc_52155_new_n15771_));
INVX1 INVX1_3433 ( .A(u2__abc_52155_new_n15778_), .Y(u2__abc_52155_new_n15779_));
INVX1 INVX1_3434 ( .A(u2__abc_52155_new_n7289_), .Y(u2__abc_52155_new_n15785_));
INVX1 INVX1_3435 ( .A(u2__abc_52155_new_n15786_), .Y(u2__abc_52155_new_n15788_));
INVX1 INVX1_3436 ( .A(u2__abc_52155_new_n15795_), .Y(u2__abc_52155_new_n15796_));
INVX1 INVX1_3437 ( .A(u2__abc_52155_new_n15804_), .Y(u2__abc_52155_new_n15805_));
INVX1 INVX1_3438 ( .A(u2__abc_52155_new_n15818_), .Y(u2__abc_52155_new_n15819_));
INVX1 INVX1_3439 ( .A(u2__abc_52155_new_n15826_), .Y(u2__abc_52155_new_n15827_));
INVX1 INVX1_344 ( .A(u2__abc_52155_new_n3406_), .Y(u2__abc_52155_new_n3407_));
INVX1 INVX1_3440 ( .A(u2__abc_52155_new_n7169_), .Y(u2__abc_52155_new_n15835_));
INVX1 INVX1_3441 ( .A(u2__abc_52155_new_n15833_), .Y(u2__abc_52155_new_n15836_));
INVX1 INVX1_3442 ( .A(u2__abc_52155_new_n15843_), .Y(u2__abc_52155_new_n15844_));
INVX1 INVX1_3443 ( .A(u2__abc_52155_new_n15852_), .Y(u2__abc_52155_new_n15853_));
INVX1 INVX1_3444 ( .A(u2__abc_52155_new_n15854_), .Y(u2__abc_52155_new_n15855_));
INVX1 INVX1_3445 ( .A(u2__abc_52155_new_n15862_), .Y(u2__abc_52155_new_n15863_));
INVX1 INVX1_3446 ( .A(u2__abc_52155_new_n7161_), .Y(u2__abc_52155_new_n15869_));
INVX1 INVX1_3447 ( .A(u2__abc_52155_new_n15870_), .Y(u2__abc_52155_new_n15872_));
INVX1 INVX1_3448 ( .A(u2__abc_52155_new_n15879_), .Y(u2__abc_52155_new_n15880_));
INVX1 INVX1_3449 ( .A(u2__abc_52155_new_n15886_), .Y(u2__abc_52155_new_n15887_));
INVX1 INVX1_345 ( .A(u2_remHi_46_), .Y(u2__abc_52155_new_n3408_));
INVX1 INVX1_3450 ( .A(u2__abc_52155_new_n15894_), .Y(u2__abc_52155_new_n15895_));
INVX1 INVX1_3451 ( .A(u2__abc_52155_new_n15902_), .Y(u2__abc_52155_new_n15903_));
INVX1 INVX1_3452 ( .A(u2__abc_52155_new_n7138_), .Y(u2__abc_52155_new_n15911_));
INVX1 INVX1_3453 ( .A(u2__abc_52155_new_n15909_), .Y(u2__abc_52155_new_n15912_));
INVX1 INVX1_3454 ( .A(u2__abc_52155_new_n15919_), .Y(u2__abc_52155_new_n15920_));
INVX1 INVX1_3455 ( .A(u2__abc_52155_new_n15928_), .Y(u2__abc_52155_new_n15929_));
INVX1 INVX1_3456 ( .A(u2__abc_52155_new_n15930_), .Y(u2__abc_52155_new_n15931_));
INVX1 INVX1_3457 ( .A(u2__abc_52155_new_n15938_), .Y(u2__abc_52155_new_n15939_));
INVX1 INVX1_3458 ( .A(u2__abc_52155_new_n7130_), .Y(u2__abc_52155_new_n15945_));
INVX1 INVX1_3459 ( .A(u2__abc_52155_new_n15946_), .Y(u2__abc_52155_new_n15948_));
INVX1 INVX1_346 ( .A(u2__abc_52155_new_n3409_), .Y(u2__abc_52155_new_n3410_));
INVX1 INVX1_3460 ( .A(u2__abc_52155_new_n15955_), .Y(u2__abc_52155_new_n15956_));
INVX1 INVX1_3461 ( .A(u2__abc_52155_new_n15963_), .Y(u2__abc_52155_new_n15964_));
INVX1 INVX1_3462 ( .A(u2__abc_52155_new_n15972_), .Y(u2__abc_52155_new_n15973_));
INVX1 INVX1_3463 ( .A(u2__abc_52155_new_n15980_), .Y(u2__abc_52155_new_n15981_));
INVX1 INVX1_3464 ( .A(u2__abc_52155_new_n7082_), .Y(u2__abc_52155_new_n15987_));
INVX1 INVX1_3465 ( .A(u2__abc_52155_new_n15988_), .Y(u2__abc_52155_new_n15989_));
INVX1 INVX1_3466 ( .A(u2__abc_52155_new_n15997_), .Y(u2__abc_52155_new_n15998_));
INVX1 INVX1_3467 ( .A(u2__abc_52155_new_n16006_), .Y(u2__abc_52155_new_n16007_));
INVX1 INVX1_3468 ( .A(u2__abc_52155_new_n16014_), .Y(u2__abc_52155_new_n16015_));
INVX1 INVX1_3469 ( .A(u2__abc_52155_new_n7067_), .Y(u2__abc_52155_new_n16021_));
INVX1 INVX1_347 ( .A(sqrto_52_), .Y(u2__abc_52155_new_n3414_));
INVX1 INVX1_3470 ( .A(u2__abc_52155_new_n16022_), .Y(u2__abc_52155_new_n16024_));
INVX1 INVX1_3471 ( .A(u2__abc_52155_new_n16031_), .Y(u2__abc_52155_new_n16032_));
INVX1 INVX1_3472 ( .A(u2__abc_52155_new_n16039_), .Y(u2__abc_52155_new_n16040_));
INVX1 INVX1_3473 ( .A(u2__abc_52155_new_n16047_), .Y(u2__abc_52155_new_n16048_));
INVX1 INVX1_3474 ( .A(u2__abc_52155_new_n16055_), .Y(u2__abc_52155_new_n16056_));
INVX1 INVX1_3475 ( .A(u2__abc_52155_new_n7106_), .Y(u2__abc_52155_new_n16064_));
INVX1 INVX1_3476 ( .A(u2__abc_52155_new_n16062_), .Y(u2__abc_52155_new_n16065_));
INVX1 INVX1_3477 ( .A(u2__abc_52155_new_n16072_), .Y(u2__abc_52155_new_n16073_));
INVX1 INVX1_3478 ( .A(u2__abc_52155_new_n16081_), .Y(u2__abc_52155_new_n16082_));
INVX1 INVX1_3479 ( .A(u2__abc_52155_new_n16083_), .Y(u2__abc_52155_new_n16084_));
INVX1 INVX1_348 ( .A(u2__abc_52155_new_n3415_), .Y(u2__abc_52155_new_n3416_));
INVX1 INVX1_3480 ( .A(u2__abc_52155_new_n16091_), .Y(u2__abc_52155_new_n16092_));
INVX1 INVX1_3481 ( .A(u2__abc_52155_new_n7098_), .Y(u2__abc_52155_new_n16098_));
INVX1 INVX1_3482 ( .A(u2__abc_52155_new_n16099_), .Y(u2__abc_52155_new_n16101_));
INVX1 INVX1_3483 ( .A(u2__abc_52155_new_n16108_), .Y(u2__abc_52155_new_n16109_));
INVX1 INVX1_3484 ( .A(u2__abc_52155_new_n16117_), .Y(u2__abc_52155_new_n16118_));
INVX1 INVX1_3485 ( .A(u2__abc_52155_new_n16127_), .Y(u2__abc_52155_new_n16128_));
INVX1 INVX1_3486 ( .A(u2__abc_52155_new_n16135_), .Y(u2__abc_52155_new_n16136_));
INVX1 INVX1_3487 ( .A(u2__abc_52155_new_n7034_), .Y(u2__abc_52155_new_n16142_));
INVX1 INVX1_3488 ( .A(u2__abc_52155_new_n16143_), .Y(u2__abc_52155_new_n16145_));
INVX1 INVX1_3489 ( .A(u2__abc_52155_new_n16152_), .Y(u2__abc_52155_new_n16153_));
INVX1 INVX1_349 ( .A(u2_remHi_52_), .Y(u2__abc_52155_new_n3417_));
INVX1 INVX1_3490 ( .A(u2__abc_52155_new_n16160_), .Y(u2__abc_52155_new_n16161_));
INVX1 INVX1_3491 ( .A(u2__abc_52155_new_n16164_), .Y(u2__abc_52155_new_n16165_));
INVX1 INVX1_3492 ( .A(u2__abc_52155_new_n16172_), .Y(u2__abc_52155_new_n16173_));
INVX1 INVX1_3493 ( .A(u2__abc_52155_new_n7049_), .Y(u2__abc_52155_new_n16179_));
INVX1 INVX1_3494 ( .A(u2__abc_52155_new_n16180_), .Y(u2__abc_52155_new_n16182_));
INVX1 INVX1_3495 ( .A(u2__abc_52155_new_n16189_), .Y(u2__abc_52155_new_n16190_));
INVX1 INVX1_3496 ( .A(u2__abc_52155_new_n16198_), .Y(u2__abc_52155_new_n16199_));
INVX1 INVX1_3497 ( .A(u2__abc_52155_new_n16200_), .Y(u2__abc_52155_new_n16201_));
INVX1 INVX1_3498 ( .A(u2__abc_52155_new_n16208_), .Y(u2__abc_52155_new_n16209_));
INVX1 INVX1_3499 ( .A(u2__abc_52155_new_n16215_), .Y(u2__abc_52155_new_n16216_));
INVX1 INVX1_35 ( .A(_abc_73687_new_n1618_), .Y(_abc_73687_new_n1621_));
INVX1 INVX1_350 ( .A(u2__abc_52155_new_n3418_), .Y(u2__abc_52155_new_n3419_));
INVX1 INVX1_3500 ( .A(u2__abc_52155_new_n16217_), .Y(u2__abc_52155_new_n16218_));
INVX1 INVX1_3501 ( .A(u2__abc_52155_new_n16225_), .Y(u2__abc_52155_new_n16226_));
INVX1 INVX1_3502 ( .A(u2__abc_52155_new_n16232_), .Y(u2__abc_52155_new_n16233_));
INVX1 INVX1_3503 ( .A(u2__abc_52155_new_n16234_), .Y(u2__abc_52155_new_n16235_));
INVX1 INVX1_3504 ( .A(u2__abc_52155_new_n16242_), .Y(u2__abc_52155_new_n16243_));
INVX1 INVX1_3505 ( .A(u2__abc_52155_new_n7003_), .Y(u2__abc_52155_new_n16249_));
INVX1 INVX1_3506 ( .A(u2__abc_52155_new_n16250_), .Y(u2__abc_52155_new_n16252_));
INVX1 INVX1_3507 ( .A(u2__abc_52155_new_n16259_), .Y(u2__abc_52155_new_n16260_));
INVX1 INVX1_3508 ( .A(u2__abc_52155_new_n16267_), .Y(u2__abc_52155_new_n16268_));
INVX1 INVX1_3509 ( .A(u2__abc_52155_new_n16269_), .Y(u2__abc_52155_new_n16270_));
INVX1 INVX1_351 ( .A(sqrto_53_), .Y(u2__abc_52155_new_n3421_));
INVX1 INVX1_3510 ( .A(u2__abc_52155_new_n16273_), .Y(u2__abc_52155_new_n16274_));
INVX1 INVX1_3511 ( .A(u2__abc_52155_new_n16282_), .Y(u2__abc_52155_new_n16283_));
INVX1 INVX1_3512 ( .A(u2__abc_52155_new_n16290_), .Y(u2__abc_52155_new_n16291_));
INVX1 INVX1_3513 ( .A(u2__abc_52155_new_n6971_), .Y(u2__abc_52155_new_n16297_));
INVX1 INVX1_3514 ( .A(u2__abc_52155_new_n16298_), .Y(u2__abc_52155_new_n16300_));
INVX1 INVX1_3515 ( .A(u2__abc_52155_new_n16307_), .Y(u2__abc_52155_new_n16308_));
INVX1 INVX1_3516 ( .A(u2__abc_52155_new_n16315_), .Y(u2__abc_52155_new_n16316_));
INVX1 INVX1_3517 ( .A(u2__abc_52155_new_n16319_), .Y(u2__abc_52155_new_n16320_));
INVX1 INVX1_3518 ( .A(u2__abc_52155_new_n16327_), .Y(u2__abc_52155_new_n16328_));
INVX1 INVX1_3519 ( .A(u2__abc_52155_new_n6986_), .Y(u2__abc_52155_new_n16334_));
INVX1 INVX1_352 ( .A(u2__abc_52155_new_n3422_), .Y(u2__abc_52155_new_n3423_));
INVX1 INVX1_3520 ( .A(u2__abc_52155_new_n16335_), .Y(u2__abc_52155_new_n16337_));
INVX1 INVX1_3521 ( .A(u2__abc_52155_new_n16344_), .Y(u2__abc_52155_new_n16345_));
INVX1 INVX1_3522 ( .A(u2__abc_52155_new_n16357_), .Y(u2__abc_52155_new_n16358_));
INVX1 INVX1_3523 ( .A(u2__abc_52155_new_n16365_), .Y(u2__abc_52155_new_n16366_));
INVX1 INVX1_3524 ( .A(u2__abc_52155_new_n6948_), .Y(u2__abc_52155_new_n16374_));
INVX1 INVX1_3525 ( .A(u2__abc_52155_new_n16372_), .Y(u2__abc_52155_new_n16375_));
INVX1 INVX1_3526 ( .A(u2__abc_52155_new_n16382_), .Y(u2__abc_52155_new_n16383_));
INVX1 INVX1_3527 ( .A(u2__abc_52155_new_n16391_), .Y(u2__abc_52155_new_n16392_));
INVX1 INVX1_3528 ( .A(u2__abc_52155_new_n16393_), .Y(u2__abc_52155_new_n16394_));
INVX1 INVX1_3529 ( .A(u2__abc_52155_new_n16401_), .Y(u2__abc_52155_new_n16402_));
INVX1 INVX1_353 ( .A(u2_remHi_53_), .Y(u2__abc_52155_new_n3424_));
INVX1 INVX1_3530 ( .A(u2__abc_52155_new_n6940_), .Y(u2__abc_52155_new_n16408_));
INVX1 INVX1_3531 ( .A(u2__abc_52155_new_n16409_), .Y(u2__abc_52155_new_n16411_));
INVX1 INVX1_3532 ( .A(u2__abc_52155_new_n16418_), .Y(u2__abc_52155_new_n16419_));
INVX1 INVX1_3533 ( .A(u2__abc_52155_new_n16431_), .Y(u2__abc_52155_new_n16432_));
INVX1 INVX1_3534 ( .A(u2__abc_52155_new_n16439_), .Y(u2__abc_52155_new_n16440_));
INVX1 INVX1_3535 ( .A(u2__abc_52155_new_n16447_), .Y(u2__abc_52155_new_n16448_));
INVX1 INVX1_3536 ( .A(u2__abc_52155_new_n3024_), .Y(u2__abc_52155_new_n16454_));
INVX1 INVX1_3537 ( .A(u2__abc_52155_new_n16455_), .Y(u2__abc_52155_new_n16457_));
INVX1 INVX1_3538 ( .A(u2__abc_52155_new_n16464_), .Y(u2__abc_52155_new_n16465_));
INVX1 INVX1_3539 ( .A(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n16470_));
INVX1 INVX1_354 ( .A(u2__abc_52155_new_n3425_), .Y(u2__abc_52155_new_n3426_));
INVX1 INVX1_3540 ( .A(u2__abc_52155_new_n2963_), .Y(u2__abc_52155_new_n16471_));
INVX1 INVX1_3541 ( .A(u2_cnt_1_), .Y(u2__abc_52155_new_n16478_));
INVX1 INVX1_3542 ( .A(u2__abc_52155_new_n16485_), .Y(u2__abc_52155_new_n16486_));
INVX1 INVX1_3543 ( .A(u2__abc_52155_new_n16493_), .Y(u2__abc_52155_new_n16494_));
INVX1 INVX1_3544 ( .A(u2__abc_52155_new_n2964_), .Y(u2__abc_52155_new_n16496_));
INVX1 INVX1_3545 ( .A(u2__abc_52155_new_n16500_), .Y(u2__abc_52155_new_n16501_));
INVX1 INVX1_3546 ( .A(u2__abc_52155_new_n16505_), .Y(u2__abc_52155_new_n16506_));
INVX1 INVX1_3547 ( .A(u2__abc_52155_new_n16511_), .Y(u2__abc_52155_new_n16512_));
INVX1 INVX1_3548 ( .A(u2__abc_52155_new_n16516_), .Y(u2__abc_52155_new_n16517_));
INVX1 INVX1_3549 ( .A(u2__abc_52155_new_n19069_), .Y(u2__abc_52155_new_n19070_));
INVX1 INVX1_355 ( .A(sqrto_51_), .Y(u2__abc_52155_new_n3429_));
INVX1 INVX1_3550 ( .A(u2__abc_52155_new_n19074_), .Y(u2__abc_52155_new_n19075_));
INVX1 INVX1_3551 ( .A(u2__abc_52155_new_n19081_), .Y(u2__abc_52155_new_n19082_));
INVX1 INVX1_3552 ( .A(u2__abc_52155_new_n19086_), .Y(u2__abc_52155_new_n19087_));
INVX1 INVX1_3553 ( .A(u2__abc_52155_new_n19094_), .Y(u2__abc_52155_new_n19095_));
INVX1 INVX1_3554 ( .A(u2__abc_52155_new_n19098_), .Y(u2__abc_52155_new_n19099_));
INVX1 INVX1_3555 ( .A(u2__abc_52155_new_n19106_), .Y(u2__abc_52155_new_n19107_));
INVX1 INVX1_3556 ( .A(u2__abc_52155_new_n19110_), .Y(u2__abc_52155_new_n19111_));
INVX1 INVX1_3557 ( .A(u2__abc_52155_new_n19118_), .Y(u2__abc_52155_new_n19119_));
INVX1 INVX1_3558 ( .A(u2__abc_52155_new_n19122_), .Y(u2__abc_52155_new_n19123_));
INVX1 INVX1_3559 ( .A(u2__abc_52155_new_n19130_), .Y(u2__abc_52155_new_n19131_));
INVX1 INVX1_356 ( .A(u2__abc_52155_new_n3430_), .Y(u2__abc_52155_new_n3431_));
INVX1 INVX1_3560 ( .A(u2__abc_52155_new_n19134_), .Y(u2__abc_52155_new_n19135_));
INVX1 INVX1_3561 ( .A(u2__abc_52155_new_n19142_), .Y(u2__abc_52155_new_n19143_));
INVX1 INVX1_3562 ( .A(u2__abc_52155_new_n19146_), .Y(u2__abc_52155_new_n19147_));
INVX1 INVX1_3563 ( .A(u2__abc_52155_new_n19154_), .Y(u2__abc_52155_new_n19155_));
INVX1 INVX1_3564 ( .A(u2__abc_52155_new_n19158_), .Y(u2__abc_52155_new_n19159_));
INVX1 INVX1_3565 ( .A(u2__abc_52155_new_n19166_), .Y(u2__abc_52155_new_n19167_));
INVX1 INVX1_3566 ( .A(u2__abc_52155_new_n19170_), .Y(u2__abc_52155_new_n19171_));
INVX1 INVX1_3567 ( .A(u2__abc_52155_new_n19178_), .Y(u2__abc_52155_new_n19179_));
INVX1 INVX1_3568 ( .A(u2__abc_52155_new_n19182_), .Y(u2__abc_52155_new_n19183_));
INVX1 INVX1_3569 ( .A(u2__abc_52155_new_n19190_), .Y(u2__abc_52155_new_n19191_));
INVX1 INVX1_357 ( .A(u2_remHi_51_), .Y(u2__abc_52155_new_n3432_));
INVX1 INVX1_3570 ( .A(u2__abc_52155_new_n19194_), .Y(u2__abc_52155_new_n19195_));
INVX1 INVX1_3571 ( .A(u2__abc_52155_new_n19202_), .Y(u2__abc_52155_new_n19203_));
INVX1 INVX1_3572 ( .A(u2__abc_52155_new_n19206_), .Y(u2__abc_52155_new_n19207_));
INVX1 INVX1_3573 ( .A(u2__abc_52155_new_n19214_), .Y(u2__abc_52155_new_n19215_));
INVX1 INVX1_3574 ( .A(u2__abc_52155_new_n19218_), .Y(u2__abc_52155_new_n19219_));
INVX1 INVX1_3575 ( .A(u2__abc_52155_new_n19226_), .Y(u2__abc_52155_new_n19227_));
INVX1 INVX1_3576 ( .A(u2__abc_52155_new_n19230_), .Y(u2__abc_52155_new_n19231_));
INVX1 INVX1_3577 ( .A(u2__abc_52155_new_n19238_), .Y(u2__abc_52155_new_n19239_));
INVX1 INVX1_3578 ( .A(u2__abc_52155_new_n19242_), .Y(u2__abc_52155_new_n19243_));
INVX1 INVX1_3579 ( .A(u2__abc_52155_new_n19250_), .Y(u2__abc_52155_new_n19251_));
INVX1 INVX1_358 ( .A(u2__abc_52155_new_n3433_), .Y(u2__abc_52155_new_n3434_));
INVX1 INVX1_3580 ( .A(u2__abc_52155_new_n19254_), .Y(u2__abc_52155_new_n19255_));
INVX1 INVX1_3581 ( .A(u2__abc_52155_new_n19262_), .Y(u2__abc_52155_new_n19263_));
INVX1 INVX1_3582 ( .A(u2__abc_52155_new_n19266_), .Y(u2__abc_52155_new_n19267_));
INVX1 INVX1_3583 ( .A(u2__abc_52155_new_n19274_), .Y(u2__abc_52155_new_n19275_));
INVX1 INVX1_3584 ( .A(u2__abc_52155_new_n19278_), .Y(u2__abc_52155_new_n19279_));
INVX1 INVX1_3585 ( .A(u2__abc_52155_new_n19286_), .Y(u2__abc_52155_new_n19287_));
INVX1 INVX1_3586 ( .A(u2__abc_52155_new_n19290_), .Y(u2__abc_52155_new_n19291_));
INVX1 INVX1_3587 ( .A(u2__abc_52155_new_n19298_), .Y(u2__abc_52155_new_n19299_));
INVX1 INVX1_3588 ( .A(u2__abc_52155_new_n19302_), .Y(u2__abc_52155_new_n19303_));
INVX1 INVX1_3589 ( .A(u2__abc_52155_new_n19310_), .Y(u2__abc_52155_new_n19311_));
INVX1 INVX1_359 ( .A(sqrto_50_), .Y(u2__abc_52155_new_n3436_));
INVX1 INVX1_3590 ( .A(u2__abc_52155_new_n19314_), .Y(u2__abc_52155_new_n19315_));
INVX1 INVX1_3591 ( .A(u2__abc_52155_new_n19322_), .Y(u2__abc_52155_new_n19323_));
INVX1 INVX1_3592 ( .A(u2__abc_52155_new_n19326_), .Y(u2__abc_52155_new_n19327_));
INVX1 INVX1_3593 ( .A(u2__abc_52155_new_n19334_), .Y(u2__abc_52155_new_n19335_));
INVX1 INVX1_3594 ( .A(u2__abc_52155_new_n19338_), .Y(u2__abc_52155_new_n19339_));
INVX1 INVX1_3595 ( .A(u2__abc_52155_new_n19346_), .Y(u2__abc_52155_new_n19347_));
INVX1 INVX1_3596 ( .A(u2__abc_52155_new_n19350_), .Y(u2__abc_52155_new_n19351_));
INVX1 INVX1_3597 ( .A(u2__abc_52155_new_n19358_), .Y(u2__abc_52155_new_n19359_));
INVX1 INVX1_3598 ( .A(u2__abc_52155_new_n19362_), .Y(u2__abc_52155_new_n19363_));
INVX1 INVX1_3599 ( .A(u2__abc_52155_new_n19370_), .Y(u2__abc_52155_new_n19371_));
INVX1 INVX1_36 ( .A(_abc_73687_new_n1619_), .Y(_abc_73687_new_n1626_));
INVX1 INVX1_360 ( .A(u2__abc_52155_new_n3437_), .Y(u2__abc_52155_new_n3438_));
INVX1 INVX1_3600 ( .A(u2__abc_52155_new_n19374_), .Y(u2__abc_52155_new_n19375_));
INVX1 INVX1_3601 ( .A(u2__abc_52155_new_n19382_), .Y(u2__abc_52155_new_n19383_));
INVX1 INVX1_3602 ( .A(u2__abc_52155_new_n19386_), .Y(u2__abc_52155_new_n19387_));
INVX1 INVX1_3603 ( .A(u2__abc_52155_new_n19394_), .Y(u2__abc_52155_new_n19395_));
INVX1 INVX1_3604 ( .A(u2__abc_52155_new_n19398_), .Y(u2__abc_52155_new_n19399_));
INVX1 INVX1_3605 ( .A(u2__abc_52155_new_n19406_), .Y(u2__abc_52155_new_n19407_));
INVX1 INVX1_3606 ( .A(u2__abc_52155_new_n19410_), .Y(u2__abc_52155_new_n19411_));
INVX1 INVX1_3607 ( .A(u2__abc_52155_new_n19418_), .Y(u2__abc_52155_new_n19419_));
INVX1 INVX1_3608 ( .A(u2__abc_52155_new_n19422_), .Y(u2__abc_52155_new_n19423_));
INVX1 INVX1_3609 ( .A(u2__abc_52155_new_n19430_), .Y(u2__abc_52155_new_n19431_));
INVX1 INVX1_361 ( .A(u2_remHi_50_), .Y(u2__abc_52155_new_n3439_));
INVX1 INVX1_3610 ( .A(u2__abc_52155_new_n19434_), .Y(u2__abc_52155_new_n19435_));
INVX1 INVX1_3611 ( .A(u2__abc_52155_new_n19442_), .Y(u2__abc_52155_new_n19443_));
INVX1 INVX1_3612 ( .A(u2__abc_52155_new_n19446_), .Y(u2__abc_52155_new_n19447_));
INVX1 INVX1_3613 ( .A(u2__abc_52155_new_n19454_), .Y(u2__abc_52155_new_n19455_));
INVX1 INVX1_3614 ( .A(u2__abc_52155_new_n19458_), .Y(u2__abc_52155_new_n19459_));
INVX1 INVX1_3615 ( .A(u2__abc_52155_new_n19466_), .Y(u2__abc_52155_new_n19467_));
INVX1 INVX1_3616 ( .A(u2__abc_52155_new_n19470_), .Y(u2__abc_52155_new_n19471_));
INVX1 INVX1_3617 ( .A(u2__abc_52155_new_n19478_), .Y(u2__abc_52155_new_n19479_));
INVX1 INVX1_3618 ( .A(u2__abc_52155_new_n19482_), .Y(u2__abc_52155_new_n19483_));
INVX1 INVX1_3619 ( .A(u2__abc_52155_new_n19490_), .Y(u2__abc_52155_new_n19491_));
INVX1 INVX1_362 ( .A(u2__abc_52155_new_n3440_), .Y(u2__abc_52155_new_n3441_));
INVX1 INVX1_3620 ( .A(u2__abc_52155_new_n19494_), .Y(u2__abc_52155_new_n19495_));
INVX1 INVX1_3621 ( .A(u2__abc_52155_new_n19502_), .Y(u2__abc_52155_new_n19503_));
INVX1 INVX1_3622 ( .A(u2__abc_52155_new_n19506_), .Y(u2__abc_52155_new_n19507_));
INVX1 INVX1_3623 ( .A(u2__abc_52155_new_n19514_), .Y(u2__abc_52155_new_n19515_));
INVX1 INVX1_3624 ( .A(u2__abc_52155_new_n19518_), .Y(u2__abc_52155_new_n19519_));
INVX1 INVX1_3625 ( .A(u2__abc_52155_new_n19526_), .Y(u2__abc_52155_new_n19527_));
INVX1 INVX1_3626 ( .A(u2__abc_52155_new_n19530_), .Y(u2__abc_52155_new_n19531_));
INVX1 INVX1_3627 ( .A(u2__abc_52155_new_n19538_), .Y(u2__abc_52155_new_n19539_));
INVX1 INVX1_3628 ( .A(u2__abc_52155_new_n19542_), .Y(u2__abc_52155_new_n19543_));
INVX1 INVX1_3629 ( .A(u2__abc_52155_new_n19550_), .Y(u2__abc_52155_new_n19551_));
INVX1 INVX1_363 ( .A(sqrto_40_), .Y(u2__abc_52155_new_n3447_));
INVX1 INVX1_3630 ( .A(u2__abc_52155_new_n19554_), .Y(u2__abc_52155_new_n19555_));
INVX1 INVX1_3631 ( .A(u2__abc_52155_new_n19562_), .Y(u2__abc_52155_new_n19563_));
INVX1 INVX1_3632 ( .A(u2__abc_52155_new_n19566_), .Y(u2__abc_52155_new_n19567_));
INVX1 INVX1_3633 ( .A(u2__abc_52155_new_n19574_), .Y(u2__abc_52155_new_n19575_));
INVX1 INVX1_3634 ( .A(u2__abc_52155_new_n19578_), .Y(u2__abc_52155_new_n19579_));
INVX1 INVX1_3635 ( .A(u2__abc_52155_new_n19586_), .Y(u2__abc_52155_new_n19587_));
INVX1 INVX1_3636 ( .A(u2__abc_52155_new_n19590_), .Y(u2__abc_52155_new_n19591_));
INVX1 INVX1_3637 ( .A(u2__abc_52155_new_n19598_), .Y(u2__abc_52155_new_n19599_));
INVX1 INVX1_3638 ( .A(u2__abc_52155_new_n19602_), .Y(u2__abc_52155_new_n19603_));
INVX1 INVX1_3639 ( .A(u2__abc_52155_new_n19610_), .Y(u2__abc_52155_new_n19611_));
INVX1 INVX1_364 ( .A(u2_remHi_40_), .Y(u2__abc_52155_new_n3449_));
INVX1 INVX1_3640 ( .A(u2__abc_52155_new_n19614_), .Y(u2__abc_52155_new_n19615_));
INVX1 INVX1_3641 ( .A(u2__abc_52155_new_n19622_), .Y(u2__abc_52155_new_n19623_));
INVX1 INVX1_3642 ( .A(u2__abc_52155_new_n19626_), .Y(u2__abc_52155_new_n19627_));
INVX1 INVX1_3643 ( .A(u2__abc_52155_new_n19634_), .Y(u2__abc_52155_new_n19635_));
INVX1 INVX1_3644 ( .A(u2__abc_52155_new_n19638_), .Y(u2__abc_52155_new_n19639_));
INVX1 INVX1_3645 ( .A(u2__abc_52155_new_n19646_), .Y(u2__abc_52155_new_n19647_));
INVX1 INVX1_3646 ( .A(u2__abc_52155_new_n19650_), .Y(u2__abc_52155_new_n19651_));
INVX1 INVX1_3647 ( .A(u2__abc_52155_new_n19658_), .Y(u2__abc_52155_new_n19659_));
INVX1 INVX1_3648 ( .A(u2__abc_52155_new_n19662_), .Y(u2__abc_52155_new_n19663_));
INVX1 INVX1_3649 ( .A(u2__abc_52155_new_n19670_), .Y(u2__abc_52155_new_n19671_));
INVX1 INVX1_365 ( .A(sqrto_41_), .Y(u2__abc_52155_new_n3452_));
INVX1 INVX1_3650 ( .A(u2__abc_52155_new_n19674_), .Y(u2__abc_52155_new_n19675_));
INVX1 INVX1_3651 ( .A(u2__abc_52155_new_n19682_), .Y(u2__abc_52155_new_n19683_));
INVX1 INVX1_3652 ( .A(u2__abc_52155_new_n19686_), .Y(u2__abc_52155_new_n19687_));
INVX1 INVX1_3653 ( .A(u2__abc_52155_new_n19694_), .Y(u2__abc_52155_new_n19695_));
INVX1 INVX1_3654 ( .A(u2__abc_52155_new_n19698_), .Y(u2__abc_52155_new_n19699_));
INVX1 INVX1_3655 ( .A(u2__abc_52155_new_n19706_), .Y(u2__abc_52155_new_n19707_));
INVX1 INVX1_3656 ( .A(u2__abc_52155_new_n19710_), .Y(u2__abc_52155_new_n19711_));
INVX1 INVX1_3657 ( .A(u2__abc_52155_new_n19718_), .Y(u2__abc_52155_new_n19719_));
INVX1 INVX1_3658 ( .A(u2__abc_52155_new_n19722_), .Y(u2__abc_52155_new_n19723_));
INVX1 INVX1_3659 ( .A(u2__abc_52155_new_n19730_), .Y(u2__abc_52155_new_n19731_));
INVX1 INVX1_366 ( .A(u2_remHi_41_), .Y(u2__abc_52155_new_n3454_));
INVX1 INVX1_3660 ( .A(u2__abc_52155_new_n19734_), .Y(u2__abc_52155_new_n19735_));
INVX1 INVX1_3661 ( .A(u2__abc_52155_new_n19742_), .Y(u2__abc_52155_new_n19743_));
INVX1 INVX1_3662 ( .A(u2__abc_52155_new_n19746_), .Y(u2__abc_52155_new_n19747_));
INVX1 INVX1_3663 ( .A(u2__abc_52155_new_n19754_), .Y(u2__abc_52155_new_n19755_));
INVX1 INVX1_3664 ( .A(u2__abc_52155_new_n19758_), .Y(u2__abc_52155_new_n19759_));
INVX1 INVX1_3665 ( .A(u2__abc_52155_new_n19766_), .Y(u2__abc_52155_new_n19767_));
INVX1 INVX1_3666 ( .A(u2__abc_52155_new_n19770_), .Y(u2__abc_52155_new_n19771_));
INVX1 INVX1_3667 ( .A(u2__abc_52155_new_n19778_), .Y(u2__abc_52155_new_n19779_));
INVX1 INVX1_3668 ( .A(u2__abc_52155_new_n19782_), .Y(u2__abc_52155_new_n19783_));
INVX1 INVX1_3669 ( .A(u2__abc_52155_new_n19790_), .Y(u2__abc_52155_new_n19791_));
INVX1 INVX1_367 ( .A(u2__abc_52155_new_n3457_), .Y(u2__abc_52155_new_n3458_));
INVX1 INVX1_3670 ( .A(u2__abc_52155_new_n19794_), .Y(u2__abc_52155_new_n19795_));
INVX1 INVX1_3671 ( .A(u2__abc_52155_new_n19802_), .Y(u2__abc_52155_new_n19803_));
INVX1 INVX1_3672 ( .A(u2__abc_52155_new_n19806_), .Y(u2__abc_52155_new_n19807_));
INVX1 INVX1_3673 ( .A(u2__abc_52155_new_n19814_), .Y(u2__abc_52155_new_n19815_));
INVX1 INVX1_3674 ( .A(u2__abc_52155_new_n19818_), .Y(u2__abc_52155_new_n19819_));
INVX1 INVX1_3675 ( .A(u2__abc_52155_new_n19826_), .Y(u2__abc_52155_new_n19827_));
INVX1 INVX1_3676 ( .A(u2__abc_52155_new_n19830_), .Y(u2__abc_52155_new_n19831_));
INVX1 INVX1_3677 ( .A(u2__abc_52155_new_n19838_), .Y(u2__abc_52155_new_n19839_));
INVX1 INVX1_3678 ( .A(u2__abc_52155_new_n19842_), .Y(u2__abc_52155_new_n19843_));
INVX1 INVX1_3679 ( .A(u2__abc_52155_new_n19850_), .Y(u2__abc_52155_new_n19851_));
INVX1 INVX1_368 ( .A(sqrto_38_), .Y(u2__abc_52155_new_n3459_));
INVX1 INVX1_3680 ( .A(u2__abc_52155_new_n19854_), .Y(u2__abc_52155_new_n19855_));
INVX1 INVX1_3681 ( .A(u2__abc_52155_new_n19862_), .Y(u2__abc_52155_new_n19863_));
INVX1 INVX1_3682 ( .A(u2__abc_52155_new_n19866_), .Y(u2__abc_52155_new_n19867_));
INVX1 INVX1_3683 ( .A(u2__abc_52155_new_n19874_), .Y(u2__abc_52155_new_n19875_));
INVX1 INVX1_3684 ( .A(u2__abc_52155_new_n19878_), .Y(u2__abc_52155_new_n19879_));
INVX1 INVX1_3685 ( .A(u2__abc_52155_new_n19886_), .Y(u2__abc_52155_new_n19887_));
INVX1 INVX1_3686 ( .A(u2__abc_52155_new_n19890_), .Y(u2__abc_52155_new_n19891_));
INVX1 INVX1_3687 ( .A(u2__abc_52155_new_n19898_), .Y(u2__abc_52155_new_n19899_));
INVX1 INVX1_3688 ( .A(u2__abc_52155_new_n19902_), .Y(u2__abc_52155_new_n19903_));
INVX1 INVX1_3689 ( .A(u2__abc_52155_new_n19910_), .Y(u2__abc_52155_new_n19911_));
INVX1 INVX1_369 ( .A(u2__abc_52155_new_n3460_), .Y(u2__abc_52155_new_n3461_));
INVX1 INVX1_3690 ( .A(u2__abc_52155_new_n19914_), .Y(u2__abc_52155_new_n19915_));
INVX1 INVX1_3691 ( .A(u2__abc_52155_new_n19922_), .Y(u2__abc_52155_new_n19923_));
INVX1 INVX1_3692 ( .A(u2__abc_52155_new_n19926_), .Y(u2__abc_52155_new_n19927_));
INVX1 INVX1_3693 ( .A(u2__abc_52155_new_n19934_), .Y(u2__abc_52155_new_n19935_));
INVX1 INVX1_3694 ( .A(u2__abc_52155_new_n19938_), .Y(u2__abc_52155_new_n19939_));
INVX1 INVX1_3695 ( .A(u2__abc_52155_new_n19946_), .Y(u2__abc_52155_new_n19947_));
INVX1 INVX1_3696 ( .A(u2__abc_52155_new_n19950_), .Y(u2__abc_52155_new_n19951_));
INVX1 INVX1_3697 ( .A(u2__abc_52155_new_n19958_), .Y(u2__abc_52155_new_n19959_));
INVX1 INVX1_3698 ( .A(u2__abc_52155_new_n19962_), .Y(u2__abc_52155_new_n19963_));
INVX1 INVX1_3699 ( .A(u2__abc_52155_new_n19970_), .Y(u2__abc_52155_new_n19971_));
INVX1 INVX1_37 ( .A(\a[123] ), .Y(_abc_73687_new_n1627_));
INVX1 INVX1_370 ( .A(u2_remHi_38_), .Y(u2__abc_52155_new_n3462_));
INVX1 INVX1_3700 ( .A(u2__abc_52155_new_n19974_), .Y(u2__abc_52155_new_n19975_));
INVX1 INVX1_3701 ( .A(u2__abc_52155_new_n19982_), .Y(u2__abc_52155_new_n19983_));
INVX1 INVX1_3702 ( .A(u2__abc_52155_new_n19986_), .Y(u2__abc_52155_new_n19987_));
INVX1 INVX1_3703 ( .A(u2__abc_52155_new_n19994_), .Y(u2__abc_52155_new_n19995_));
INVX1 INVX1_3704 ( .A(u2__abc_52155_new_n19998_), .Y(u2__abc_52155_new_n19999_));
INVX1 INVX1_3705 ( .A(u2__abc_52155_new_n20006_), .Y(u2__abc_52155_new_n20007_));
INVX1 INVX1_3706 ( .A(u2__abc_52155_new_n20010_), .Y(u2__abc_52155_new_n20011_));
INVX1 INVX1_3707 ( .A(u2__abc_52155_new_n20018_), .Y(u2__abc_52155_new_n20019_));
INVX1 INVX1_3708 ( .A(u2__abc_52155_new_n20022_), .Y(u2__abc_52155_new_n20023_));
INVX1 INVX1_3709 ( .A(u2__abc_52155_new_n20029_), .Y(u2__abc_52155_new_n20030_));
INVX1 INVX1_371 ( .A(u2__abc_52155_new_n3463_), .Y(u2__abc_52155_new_n3464_));
INVX1 INVX1_3710 ( .A(u2__abc_52155_new_n20034_), .Y(u2__abc_52155_new_n20035_));
INVX1 INVX1_3711 ( .A(u2__abc_52155_new_n20042_), .Y(u2__abc_52155_new_n20043_));
INVX1 INVX1_3712 ( .A(u2__abc_52155_new_n20046_), .Y(u2__abc_52155_new_n20047_));
INVX1 INVX1_3713 ( .A(u2__abc_52155_new_n20054_), .Y(u2__abc_52155_new_n20055_));
INVX1 INVX1_3714 ( .A(u2__abc_52155_new_n20058_), .Y(u2__abc_52155_new_n20059_));
INVX1 INVX1_3715 ( .A(u2__abc_52155_new_n20066_), .Y(u2__abc_52155_new_n20067_));
INVX1 INVX1_3716 ( .A(u2__abc_52155_new_n20070_), .Y(u2__abc_52155_new_n20071_));
INVX1 INVX1_3717 ( .A(u2__abc_52155_new_n20078_), .Y(u2__abc_52155_new_n20079_));
INVX1 INVX1_3718 ( .A(u2__abc_52155_new_n20082_), .Y(u2__abc_52155_new_n20083_));
INVX1 INVX1_3719 ( .A(u2__abc_52155_new_n20090_), .Y(u2__abc_52155_new_n20091_));
INVX1 INVX1_372 ( .A(sqrto_39_), .Y(u2__abc_52155_new_n3466_));
INVX1 INVX1_3720 ( .A(u2__abc_52155_new_n20094_), .Y(u2__abc_52155_new_n20095_));
INVX1 INVX1_3721 ( .A(u2__abc_52155_new_n20102_), .Y(u2__abc_52155_new_n20103_));
INVX1 INVX1_3722 ( .A(u2__abc_52155_new_n20106_), .Y(u2__abc_52155_new_n20107_));
INVX1 INVX1_3723 ( .A(u2__abc_52155_new_n20114_), .Y(u2__abc_52155_new_n20115_));
INVX1 INVX1_3724 ( .A(u2__abc_52155_new_n20118_), .Y(u2__abc_52155_new_n20119_));
INVX1 INVX1_3725 ( .A(u2__abc_52155_new_n20125_), .Y(u2__abc_52155_new_n20126_));
INVX1 INVX1_3726 ( .A(u2__abc_52155_new_n20130_), .Y(u2__abc_52155_new_n20131_));
INVX1 INVX1_3727 ( .A(u2__abc_52155_new_n20138_), .Y(u2__abc_52155_new_n20139_));
INVX1 INVX1_3728 ( .A(u2__abc_52155_new_n20142_), .Y(u2__abc_52155_new_n20143_));
INVX1 INVX1_3729 ( .A(u2__abc_52155_new_n20150_), .Y(u2__abc_52155_new_n20151_));
INVX1 INVX1_373 ( .A(u2__abc_52155_new_n3467_), .Y(u2__abc_52155_new_n3468_));
INVX1 INVX1_3730 ( .A(u2__abc_52155_new_n20154_), .Y(u2__abc_52155_new_n20155_));
INVX1 INVX1_3731 ( .A(u2__abc_52155_new_n20162_), .Y(u2__abc_52155_new_n20163_));
INVX1 INVX1_3732 ( .A(u2__abc_52155_new_n20166_), .Y(u2__abc_52155_new_n20167_));
INVX1 INVX1_3733 ( .A(u2__abc_52155_new_n20173_), .Y(u2__abc_52155_new_n20174_));
INVX1 INVX1_3734 ( .A(u2__abc_52155_new_n20178_), .Y(u2__abc_52155_new_n20179_));
INVX1 INVX1_3735 ( .A(u2__abc_52155_new_n20186_), .Y(u2__abc_52155_new_n20187_));
INVX1 INVX1_3736 ( .A(u2__abc_52155_new_n20190_), .Y(u2__abc_52155_new_n20191_));
INVX1 INVX1_3737 ( .A(u2__abc_52155_new_n20197_), .Y(u2__abc_52155_new_n20198_));
INVX1 INVX1_3738 ( .A(u2__abc_52155_new_n20202_), .Y(u2__abc_52155_new_n20203_));
INVX1 INVX1_3739 ( .A(u2__abc_52155_new_n20210_), .Y(u2__abc_52155_new_n20211_));
INVX1 INVX1_374 ( .A(u2_remHi_39_), .Y(u2__abc_52155_new_n3469_));
INVX1 INVX1_3740 ( .A(u2__abc_52155_new_n20214_), .Y(u2__abc_52155_new_n20215_));
INVX1 INVX1_3741 ( .A(u2__abc_52155_new_n20222_), .Y(u2__abc_52155_new_n20223_));
INVX1 INVX1_3742 ( .A(u2__abc_52155_new_n20226_), .Y(u2__abc_52155_new_n20227_));
INVX1 INVX1_3743 ( .A(u2__abc_52155_new_n20234_), .Y(u2__abc_52155_new_n20235_));
INVX1 INVX1_3744 ( .A(u2__abc_52155_new_n20238_), .Y(u2__abc_52155_new_n20239_));
INVX1 INVX1_3745 ( .A(u2__abc_52155_new_n20246_), .Y(u2__abc_52155_new_n20247_));
INVX1 INVX1_3746 ( .A(u2__abc_52155_new_n20250_), .Y(u2__abc_52155_new_n20251_));
INVX1 INVX1_3747 ( .A(u2__abc_52155_new_n20258_), .Y(u2__abc_52155_new_n20259_));
INVX1 INVX1_3748 ( .A(u2__abc_52155_new_n20262_), .Y(u2__abc_52155_new_n20263_));
INVX1 INVX1_3749 ( .A(u2__abc_52155_new_n20270_), .Y(u2__abc_52155_new_n20271_));
INVX1 INVX1_375 ( .A(u2__abc_52155_new_n3470_), .Y(u2__abc_52155_new_n3471_));
INVX1 INVX1_3750 ( .A(u2__abc_52155_new_n20274_), .Y(u2__abc_52155_new_n20275_));
INVX1 INVX1_3751 ( .A(u2__abc_52155_new_n20282_), .Y(u2__abc_52155_new_n20283_));
INVX1 INVX1_3752 ( .A(u2__abc_52155_new_n20286_), .Y(u2__abc_52155_new_n20287_));
INVX1 INVX1_3753 ( .A(u2__abc_52155_new_n20294_), .Y(u2__abc_52155_new_n20295_));
INVX1 INVX1_3754 ( .A(u2__abc_52155_new_n20298_), .Y(u2__abc_52155_new_n20299_));
INVX1 INVX1_3755 ( .A(u2__abc_52155_new_n20306_), .Y(u2__abc_52155_new_n20307_));
INVX1 INVX1_3756 ( .A(u2__abc_52155_new_n20310_), .Y(u2__abc_52155_new_n20311_));
INVX1 INVX1_3757 ( .A(u2__abc_52155_new_n20317_), .Y(u2__abc_52155_new_n20318_));
INVX1 INVX1_3758 ( .A(u2__abc_52155_new_n20322_), .Y(u2__abc_52155_new_n20323_));
INVX1 INVX1_3759 ( .A(u2__abc_52155_new_n20330_), .Y(u2__abc_52155_new_n20331_));
INVX1 INVX1_376 ( .A(sqrto_44_), .Y(u2__abc_52155_new_n3475_));
INVX1 INVX1_3760 ( .A(u2__abc_52155_new_n20334_), .Y(u2__abc_52155_new_n20335_));
INVX1 INVX1_3761 ( .A(u2__abc_52155_new_n20342_), .Y(u2__abc_52155_new_n20343_));
INVX1 INVX1_3762 ( .A(u2__abc_52155_new_n20346_), .Y(u2__abc_52155_new_n20347_));
INVX1 INVX1_3763 ( .A(u2__abc_52155_new_n20354_), .Y(u2__abc_52155_new_n20355_));
INVX1 INVX1_3764 ( .A(u2__abc_52155_new_n20358_), .Y(u2__abc_52155_new_n20359_));
INVX1 INVX1_3765 ( .A(u2__abc_52155_new_n20365_), .Y(u2__abc_52155_new_n20366_));
INVX1 INVX1_3766 ( .A(u2__abc_52155_new_n20370_), .Y(u2__abc_52155_new_n20371_));
INVX1 INVX1_3767 ( .A(u2__abc_52155_new_n20378_), .Y(u2__abc_52155_new_n20379_));
INVX1 INVX1_3768 ( .A(u2__abc_52155_new_n20382_), .Y(u2__abc_52155_new_n20383_));
INVX1 INVX1_3769 ( .A(u2__abc_52155_new_n20389_), .Y(u2__abc_52155_new_n20390_));
INVX1 INVX1_377 ( .A(u2__abc_52155_new_n3476_), .Y(u2__abc_52155_new_n3477_));
INVX1 INVX1_3770 ( .A(u2__abc_52155_new_n20394_), .Y(u2__abc_52155_new_n20395_));
INVX1 INVX1_3771 ( .A(u2__abc_52155_new_n20402_), .Y(u2__abc_52155_new_n20403_));
INVX1 INVX1_3772 ( .A(u2__abc_52155_new_n20406_), .Y(u2__abc_52155_new_n20407_));
INVX1 INVX1_3773 ( .A(u2__abc_52155_new_n20414_), .Y(u2__abc_52155_new_n20415_));
INVX1 INVX1_3774 ( .A(u2__abc_52155_new_n20418_), .Y(u2__abc_52155_new_n20419_));
INVX1 INVX1_3775 ( .A(u2__abc_52155_new_n20426_), .Y(u2__abc_52155_new_n20427_));
INVX1 INVX1_3776 ( .A(u2__abc_52155_new_n20430_), .Y(u2__abc_52155_new_n20431_));
INVX1 INVX1_3777 ( .A(u2__abc_52155_new_n20438_), .Y(u2__abc_52155_new_n20439_));
INVX1 INVX1_3778 ( .A(u2__abc_52155_new_n20442_), .Y(u2__abc_52155_new_n20443_));
INVX1 INVX1_3779 ( .A(u2__abc_52155_new_n20450_), .Y(u2__abc_52155_new_n20451_));
INVX1 INVX1_378 ( .A(u2_remHi_44_), .Y(u2__abc_52155_new_n3478_));
INVX1 INVX1_3780 ( .A(u2__abc_52155_new_n20454_), .Y(u2__abc_52155_new_n20455_));
INVX1 INVX1_3781 ( .A(u2__abc_52155_new_n20461_), .Y(u2__abc_52155_new_n20462_));
INVX1 INVX1_3782 ( .A(u2__abc_52155_new_n20466_), .Y(u2__abc_52155_new_n20467_));
INVX1 INVX1_3783 ( .A(u2__abc_52155_new_n20474_), .Y(u2__abc_52155_new_n20475_));
INVX1 INVX1_3784 ( .A(u2__abc_52155_new_n20478_), .Y(u2__abc_52155_new_n20479_));
INVX1 INVX1_3785 ( .A(u2__abc_52155_new_n20485_), .Y(u2__abc_52155_new_n20486_));
INVX1 INVX1_3786 ( .A(u2__abc_52155_new_n20490_), .Y(u2__abc_52155_new_n20491_));
INVX1 INVX1_3787 ( .A(u2__abc_52155_new_n20498_), .Y(u2__abc_52155_new_n20499_));
INVX1 INVX1_3788 ( .A(u2__abc_52155_new_n20502_), .Y(u2__abc_52155_new_n20503_));
INVX1 INVX1_3789 ( .A(u2__abc_52155_new_n20510_), .Y(u2__abc_52155_new_n20511_));
INVX1 INVX1_379 ( .A(u2__abc_52155_new_n3479_), .Y(u2__abc_52155_new_n3480_));
INVX1 INVX1_3790 ( .A(u2__abc_52155_new_n20514_), .Y(u2__abc_52155_new_n20515_));
INVX1 INVX1_3791 ( .A(u2__abc_52155_new_n20522_), .Y(u2__abc_52155_new_n20523_));
INVX1 INVX1_3792 ( .A(u2__abc_52155_new_n20526_), .Y(u2__abc_52155_new_n20527_));
INVX1 INVX1_3793 ( .A(u2__abc_52155_new_n20533_), .Y(u2__abc_52155_new_n20534_));
INVX1 INVX1_3794 ( .A(u2__abc_52155_new_n20538_), .Y(u2__abc_52155_new_n20539_));
INVX1 INVX1_3795 ( .A(u2__abc_52155_new_n20546_), .Y(u2__abc_52155_new_n20547_));
INVX1 INVX1_3796 ( .A(u2__abc_52155_new_n20550_), .Y(u2__abc_52155_new_n20551_));
INVX1 INVX1_3797 ( .A(u2__abc_52155_new_n20558_), .Y(u2__abc_52155_new_n20559_));
INVX1 INVX1_3798 ( .A(u2__abc_52155_new_n20562_), .Y(u2__abc_52155_new_n20563_));
INVX1 INVX1_3799 ( .A(u2__abc_52155_new_n20570_), .Y(u2__abc_52155_new_n20571_));
INVX1 INVX1_38 ( .A(_abc_73687_new_n1630_), .Y(_abc_73687_new_n1631_));
INVX1 INVX1_380 ( .A(sqrto_45_), .Y(u2__abc_52155_new_n3482_));
INVX1 INVX1_3800 ( .A(u2__abc_52155_new_n20574_), .Y(u2__abc_52155_new_n20575_));
INVX1 INVX1_3801 ( .A(u2__abc_52155_new_n20581_), .Y(u2__abc_52155_new_n20582_));
INVX1 INVX1_3802 ( .A(u2__abc_52155_new_n20586_), .Y(u2__abc_52155_new_n20587_));
INVX1 INVX1_3803 ( .A(u2__abc_52155_new_n20594_), .Y(u2__abc_52155_new_n20595_));
INVX1 INVX1_3804 ( .A(u2__abc_52155_new_n20598_), .Y(u2__abc_52155_new_n20599_));
INVX1 INVX1_3805 ( .A(u2__abc_52155_new_n20606_), .Y(u2__abc_52155_new_n20607_));
INVX1 INVX1_3806 ( .A(u2__abc_52155_new_n20610_), .Y(u2__abc_52155_new_n20611_));
INVX1 INVX1_3807 ( .A(u2__abc_52155_new_n20618_), .Y(u2__abc_52155_new_n20619_));
INVX1 INVX1_3808 ( .A(u2__abc_52155_new_n20622_), .Y(u2__abc_52155_new_n20623_));
INVX1 INVX1_3809 ( .A(u2__abc_52155_new_n20630_), .Y(u2__abc_52155_new_n20631_));
INVX1 INVX1_381 ( .A(u2__abc_52155_new_n3483_), .Y(u2__abc_52155_new_n3484_));
INVX1 INVX1_3810 ( .A(u2__abc_52155_new_n20634_), .Y(u2__abc_52155_new_n20635_));
INVX1 INVX1_3811 ( .A(u2__abc_52155_new_n20642_), .Y(u2__abc_52155_new_n20643_));
INVX1 INVX1_3812 ( .A(u2__abc_52155_new_n20646_), .Y(u2__abc_52155_new_n20647_));
INVX1 INVX1_3813 ( .A(u2__abc_52155_new_n20654_), .Y(u2__abc_52155_new_n20655_));
INVX1 INVX1_3814 ( .A(u2__abc_52155_new_n20658_), .Y(u2__abc_52155_new_n20659_));
INVX1 INVX1_3815 ( .A(u2__abc_52155_new_n20666_), .Y(u2__abc_52155_new_n20667_));
INVX1 INVX1_3816 ( .A(u2__abc_52155_new_n20670_), .Y(u2__abc_52155_new_n20671_));
INVX1 INVX1_3817 ( .A(u2__abc_52155_new_n20678_), .Y(u2__abc_52155_new_n20679_));
INVX1 INVX1_3818 ( .A(u2__abc_52155_new_n20682_), .Y(u2__abc_52155_new_n20683_));
INVX1 INVX1_3819 ( .A(u2__abc_52155_new_n20690_), .Y(u2__abc_52155_new_n20691_));
INVX1 INVX1_382 ( .A(u2_remHi_45_), .Y(u2__abc_52155_new_n3485_));
INVX1 INVX1_3820 ( .A(u2__abc_52155_new_n20694_), .Y(u2__abc_52155_new_n20695_));
INVX1 INVX1_3821 ( .A(u2__abc_52155_new_n20701_), .Y(u2__abc_52155_new_n20702_));
INVX1 INVX1_3822 ( .A(u2__abc_52155_new_n20706_), .Y(u2__abc_52155_new_n20707_));
INVX1 INVX1_3823 ( .A(u2__abc_52155_new_n20714_), .Y(u2__abc_52155_new_n20715_));
INVX1 INVX1_3824 ( .A(u2__abc_52155_new_n20718_), .Y(u2__abc_52155_new_n20719_));
INVX1 INVX1_3825 ( .A(u2__abc_52155_new_n20726_), .Y(u2__abc_52155_new_n20727_));
INVX1 INVX1_3826 ( .A(u2__abc_52155_new_n20730_), .Y(u2__abc_52155_new_n20731_));
INVX1 INVX1_3827 ( .A(u2__abc_52155_new_n20738_), .Y(u2__abc_52155_new_n20739_));
INVX1 INVX1_3828 ( .A(u2__abc_52155_new_n20742_), .Y(u2__abc_52155_new_n20743_));
INVX1 INVX1_3829 ( .A(u2__abc_52155_new_n20749_), .Y(u2__abc_52155_new_n20750_));
INVX1 INVX1_383 ( .A(u2__abc_52155_new_n3486_), .Y(u2__abc_52155_new_n3487_));
INVX1 INVX1_3830 ( .A(u2__abc_52155_new_n20754_), .Y(u2__abc_52155_new_n20755_));
INVX1 INVX1_3831 ( .A(u2__abc_52155_new_n20762_), .Y(u2__abc_52155_new_n20763_));
INVX1 INVX1_3832 ( .A(u2__abc_52155_new_n20766_), .Y(u2__abc_52155_new_n20767_));
INVX1 INVX1_3833 ( .A(u2__abc_52155_new_n20773_), .Y(u2__abc_52155_new_n20774_));
INVX1 INVX1_3834 ( .A(u2__abc_52155_new_n20778_), .Y(u2__abc_52155_new_n20779_));
INVX1 INVX1_3835 ( .A(u2__abc_52155_new_n20786_), .Y(u2__abc_52155_new_n20787_));
INVX1 INVX1_3836 ( .A(u2__abc_52155_new_n20790_), .Y(u2__abc_52155_new_n20791_));
INVX1 INVX1_3837 ( .A(u2__abc_52155_new_n20798_), .Y(u2__abc_52155_new_n20799_));
INVX1 INVX1_3838 ( .A(u2__abc_52155_new_n20802_), .Y(u2__abc_52155_new_n20803_));
INVX1 INVX1_3839 ( .A(u2__abc_52155_new_n20810_), .Y(u2__abc_52155_new_n20811_));
INVX1 INVX1_384 ( .A(sqrto_43_), .Y(u2__abc_52155_new_n3490_));
INVX1 INVX1_3840 ( .A(u2__abc_52155_new_n20814_), .Y(u2__abc_52155_new_n20815_));
INVX1 INVX1_3841 ( .A(u2__abc_52155_new_n20822_), .Y(u2__abc_52155_new_n20823_));
INVX1 INVX1_3842 ( .A(u2__abc_52155_new_n20826_), .Y(u2__abc_52155_new_n20827_));
INVX1 INVX1_3843 ( .A(u2__abc_52155_new_n20834_), .Y(u2__abc_52155_new_n20835_));
INVX1 INVX1_3844 ( .A(u2__abc_52155_new_n20838_), .Y(u2__abc_52155_new_n20839_));
INVX1 INVX1_3845 ( .A(u2__abc_52155_new_n20845_), .Y(u2__abc_52155_new_n20846_));
INVX1 INVX1_3846 ( .A(u2__abc_52155_new_n20850_), .Y(u2__abc_52155_new_n20851_));
INVX1 INVX1_3847 ( .A(u2__abc_52155_new_n20858_), .Y(u2__abc_52155_new_n20859_));
INVX1 INVX1_3848 ( .A(u2__abc_52155_new_n20862_), .Y(u2__abc_52155_new_n20863_));
INVX1 INVX1_3849 ( .A(u2__abc_52155_new_n20869_), .Y(u2__abc_52155_new_n20870_));
INVX1 INVX1_385 ( .A(u2__abc_52155_new_n3491_), .Y(u2__abc_52155_new_n3492_));
INVX1 INVX1_3850 ( .A(u2__abc_52155_new_n20874_), .Y(u2__abc_52155_new_n20875_));
INVX1 INVX1_3851 ( .A(u2__abc_52155_new_n20882_), .Y(u2__abc_52155_new_n20883_));
INVX1 INVX1_3852 ( .A(u2__abc_52155_new_n20886_), .Y(u2__abc_52155_new_n20887_));
INVX1 INVX1_3853 ( .A(u2__abc_52155_new_n20894_), .Y(u2__abc_52155_new_n20895_));
INVX1 INVX1_3854 ( .A(u2__abc_52155_new_n20898_), .Y(u2__abc_52155_new_n20899_));
INVX1 INVX1_3855 ( .A(u2__abc_52155_new_n20906_), .Y(u2__abc_52155_new_n20907_));
INVX1 INVX1_3856 ( .A(u2__abc_52155_new_n20910_), .Y(u2__abc_52155_new_n20911_));
INVX1 INVX1_3857 ( .A(u2__abc_52155_new_n20917_), .Y(u2__abc_52155_new_n20918_));
INVX1 INVX1_3858 ( .A(u2__abc_52155_new_n20922_), .Y(u2__abc_52155_new_n20923_));
INVX1 INVX1_3859 ( .A(u2__abc_52155_new_n20930_), .Y(u2__abc_52155_new_n20931_));
INVX1 INVX1_386 ( .A(u2_remHi_43_), .Y(u2__abc_52155_new_n3493_));
INVX1 INVX1_3860 ( .A(u2__abc_52155_new_n20934_), .Y(u2__abc_52155_new_n20935_));
INVX1 INVX1_3861 ( .A(u2__abc_52155_new_n20942_), .Y(u2__abc_52155_new_n20943_));
INVX1 INVX1_3862 ( .A(u2__abc_52155_new_n20946_), .Y(u2__abc_52155_new_n20947_));
INVX1 INVX1_3863 ( .A(u2__abc_52155_new_n20954_), .Y(u2__abc_52155_new_n20955_));
INVX1 INVX1_3864 ( .A(u2__abc_52155_new_n20958_), .Y(u2__abc_52155_new_n20959_));
INVX1 INVX1_3865 ( .A(u2__abc_52155_new_n20965_), .Y(u2__abc_52155_new_n20966_));
INVX1 INVX1_3866 ( .A(u2__abc_52155_new_n20970_), .Y(u2__abc_52155_new_n20971_));
INVX1 INVX1_3867 ( .A(u2__abc_52155_new_n20978_), .Y(u2__abc_52155_new_n20979_));
INVX1 INVX1_3868 ( .A(u2__abc_52155_new_n20982_), .Y(u2__abc_52155_new_n20983_));
INVX1 INVX1_3869 ( .A(u2__abc_52155_new_n20990_), .Y(u2__abc_52155_new_n20991_));
INVX1 INVX1_387 ( .A(u2__abc_52155_new_n3494_), .Y(u2__abc_52155_new_n3495_));
INVX1 INVX1_3870 ( .A(u2__abc_52155_new_n20994_), .Y(u2__abc_52155_new_n20995_));
INVX1 INVX1_3871 ( .A(u2__abc_52155_new_n21002_), .Y(u2__abc_52155_new_n21003_));
INVX1 INVX1_3872 ( .A(u2__abc_52155_new_n21006_), .Y(u2__abc_52155_new_n21007_));
INVX1 INVX1_3873 ( .A(u2__abc_52155_new_n21014_), .Y(u2__abc_52155_new_n21015_));
INVX1 INVX1_3874 ( .A(u2__abc_52155_new_n21018_), .Y(u2__abc_52155_new_n21019_));
INVX1 INVX1_3875 ( .A(u2__abc_52155_new_n21026_), .Y(u2__abc_52155_new_n21027_));
INVX1 INVX1_3876 ( .A(u2__abc_52155_new_n21030_), .Y(u2__abc_52155_new_n21031_));
INVX1 INVX1_3877 ( .A(u2__abc_52155_new_n21037_), .Y(u2__abc_52155_new_n21038_));
INVX1 INVX1_3878 ( .A(u2__abc_52155_new_n21042_), .Y(u2__abc_52155_new_n21043_));
INVX1 INVX1_3879 ( .A(u2__abc_52155_new_n21050_), .Y(u2__abc_52155_new_n21051_));
INVX1 INVX1_388 ( .A(sqrto_42_), .Y(u2__abc_52155_new_n3497_));
INVX1 INVX1_3880 ( .A(u2__abc_52155_new_n21054_), .Y(u2__abc_52155_new_n21055_));
INVX1 INVX1_3881 ( .A(u2__abc_52155_new_n21061_), .Y(u2__abc_52155_new_n21062_));
INVX1 INVX1_3882 ( .A(u2__abc_52155_new_n21066_), .Y(u2__abc_52155_new_n21067_));
INVX1 INVX1_3883 ( .A(u2__abc_52155_new_n21074_), .Y(u2__abc_52155_new_n21075_));
INVX1 INVX1_3884 ( .A(u2__abc_52155_new_n21078_), .Y(u2__abc_52155_new_n21079_));
INVX1 INVX1_3885 ( .A(u2__abc_52155_new_n21086_), .Y(u2__abc_52155_new_n21087_));
INVX1 INVX1_3886 ( .A(u2__abc_52155_new_n21090_), .Y(u2__abc_52155_new_n21091_));
INVX1 INVX1_3887 ( .A(u2__abc_52155_new_n21098_), .Y(u2__abc_52155_new_n21099_));
INVX1 INVX1_3888 ( .A(u2__abc_52155_new_n21102_), .Y(u2__abc_52155_new_n21103_));
INVX1 INVX1_3889 ( .A(u2__abc_52155_new_n21109_), .Y(u2__abc_52155_new_n21110_));
INVX1 INVX1_389 ( .A(u2__abc_52155_new_n3498_), .Y(u2__abc_52155_new_n3499_));
INVX1 INVX1_3890 ( .A(u2__abc_52155_new_n21114_), .Y(u2__abc_52155_new_n21115_));
INVX1 INVX1_3891 ( .A(u2__abc_52155_new_n21122_), .Y(u2__abc_52155_new_n21123_));
INVX1 INVX1_3892 ( .A(u2__abc_52155_new_n21126_), .Y(u2__abc_52155_new_n21127_));
INVX1 INVX1_3893 ( .A(u2__abc_52155_new_n21134_), .Y(u2__abc_52155_new_n21135_));
INVX1 INVX1_3894 ( .A(u2__abc_52155_new_n21138_), .Y(u2__abc_52155_new_n21139_));
INVX1 INVX1_3895 ( .A(u2__abc_52155_new_n21146_), .Y(u2__abc_52155_new_n21147_));
INVX1 INVX1_3896 ( .A(u2__abc_52155_new_n21150_), .Y(u2__abc_52155_new_n21151_));
INVX1 INVX1_3897 ( .A(u2__abc_52155_new_n21157_), .Y(u2__abc_52155_new_n21158_));
INVX1 INVX1_3898 ( .A(u2__abc_52155_new_n21162_), .Y(u2__abc_52155_new_n21163_));
INVX1 INVX1_3899 ( .A(u2__abc_52155_new_n21170_), .Y(u2__abc_52155_new_n21171_));
INVX1 INVX1_39 ( .A(_abc_73687_new_n1634_), .Y(_abc_73687_new_n1635_));
INVX1 INVX1_390 ( .A(u2_remHi_42_), .Y(u2__abc_52155_new_n3500_));
INVX1 INVX1_3900 ( .A(u2__abc_52155_new_n21174_), .Y(u2__abc_52155_new_n21175_));
INVX1 INVX1_3901 ( .A(u2__abc_52155_new_n21182_), .Y(u2__abc_52155_new_n21183_));
INVX1 INVX1_3902 ( .A(u2__abc_52155_new_n21186_), .Y(u2__abc_52155_new_n21187_));
INVX1 INVX1_3903 ( .A(u2__abc_52155_new_n21194_), .Y(u2__abc_52155_new_n21195_));
INVX1 INVX1_3904 ( .A(u2__abc_52155_new_n21198_), .Y(u2__abc_52155_new_n21199_));
INVX1 INVX1_3905 ( .A(u2__abc_52155_new_n21205_), .Y(u2__abc_52155_new_n21206_));
INVX1 INVX1_3906 ( .A(u2__abc_52155_new_n21210_), .Y(u2__abc_52155_new_n21211_));
INVX1 INVX1_3907 ( .A(u2__abc_52155_new_n21218_), .Y(u2__abc_52155_new_n21219_));
INVX1 INVX1_3908 ( .A(u2__abc_52155_new_n21222_), .Y(u2__abc_52155_new_n21223_));
INVX1 INVX1_3909 ( .A(u2__abc_52155_new_n21230_), .Y(u2__abc_52155_new_n21231_));
INVX1 INVX1_391 ( .A(u2__abc_52155_new_n3501_), .Y(u2__abc_52155_new_n3502_));
INVX1 INVX1_3910 ( .A(u2__abc_52155_new_n21234_), .Y(u2__abc_52155_new_n21235_));
INVX1 INVX1_3911 ( .A(u2__abc_52155_new_n21242_), .Y(u2__abc_52155_new_n21243_));
INVX1 INVX1_3912 ( .A(u2__abc_52155_new_n21246_), .Y(u2__abc_52155_new_n21247_));
INVX1 INVX1_3913 ( .A(u2__abc_52155_new_n21253_), .Y(u2__abc_52155_new_n21254_));
INVX1 INVX1_3914 ( .A(u2__abc_52155_new_n21258_), .Y(u2__abc_52155_new_n21259_));
INVX1 INVX1_3915 ( .A(u2__abc_52155_new_n21266_), .Y(u2__abc_52155_new_n21267_));
INVX1 INVX1_3916 ( .A(u2__abc_52155_new_n21270_), .Y(u2__abc_52155_new_n21271_));
INVX1 INVX1_3917 ( .A(u2__abc_52155_new_n21278_), .Y(u2__abc_52155_new_n21279_));
INVX1 INVX1_3918 ( .A(u2__abc_52155_new_n21282_), .Y(u2__abc_52155_new_n21283_));
INVX1 INVX1_3919 ( .A(u2__abc_52155_new_n21290_), .Y(u2__abc_52155_new_n21291_));
INVX1 INVX1_392 ( .A(sqrto_32_), .Y(u2__abc_52155_new_n3507_));
INVX1 INVX1_3920 ( .A(u2__abc_52155_new_n21294_), .Y(u2__abc_52155_new_n21295_));
INVX1 INVX1_3921 ( .A(u2__abc_52155_new_n21301_), .Y(u2__abc_52155_new_n21302_));
INVX1 INVX1_3922 ( .A(u2__abc_52155_new_n21306_), .Y(u2__abc_52155_new_n21307_));
INVX1 INVX1_3923 ( .A(u2__abc_52155_new_n21314_), .Y(u2__abc_52155_new_n21315_));
INVX1 INVX1_3924 ( .A(u2__abc_52155_new_n21318_), .Y(u2__abc_52155_new_n21319_));
INVX1 INVX1_3925 ( .A(u2__abc_52155_new_n21326_), .Y(u2__abc_52155_new_n21327_));
INVX1 INVX1_3926 ( .A(u2__abc_52155_new_n21330_), .Y(u2__abc_52155_new_n21331_));
INVX1 INVX1_3927 ( .A(u2__abc_52155_new_n21338_), .Y(u2__abc_52155_new_n21339_));
INVX1 INVX1_3928 ( .A(u2__abc_52155_new_n21342_), .Y(u2__abc_52155_new_n21343_));
INVX1 INVX1_3929 ( .A(u2__abc_52155_new_n21349_), .Y(u2__abc_52155_new_n21350_));
INVX1 INVX1_393 ( .A(u2_remHi_32_), .Y(u2__abc_52155_new_n3509_));
INVX1 INVX1_3930 ( .A(u2__abc_52155_new_n21354_), .Y(u2__abc_52155_new_n21355_));
INVX1 INVX1_3931 ( .A(u2__abc_52155_new_n21362_), .Y(u2__abc_52155_new_n21363_));
INVX1 INVX1_3932 ( .A(u2__abc_52155_new_n21366_), .Y(u2__abc_52155_new_n21367_));
INVX1 INVX1_3933 ( .A(u2__abc_52155_new_n21373_), .Y(u2__abc_52155_new_n21374_));
INVX1 INVX1_3934 ( .A(u2__abc_52155_new_n21378_), .Y(u2__abc_52155_new_n21379_));
INVX1 INVX1_3935 ( .A(u2__abc_52155_new_n21386_), .Y(u2__abc_52155_new_n21387_));
INVX1 INVX1_3936 ( .A(u2__abc_52155_new_n21390_), .Y(u2__abc_52155_new_n21391_));
INVX1 INVX1_3937 ( .A(u2__abc_52155_new_n21398_), .Y(u2__abc_52155_new_n21399_));
INVX1 INVX1_3938 ( .A(u2__abc_52155_new_n21402_), .Y(u2__abc_52155_new_n21403_));
INVX1 INVX1_3939 ( .A(u2__abc_52155_new_n21410_), .Y(u2__abc_52155_new_n21411_));
INVX1 INVX1_394 ( .A(sqrto_33_), .Y(u2__abc_52155_new_n3512_));
INVX1 INVX1_3940 ( .A(u2__abc_52155_new_n21414_), .Y(u2__abc_52155_new_n21415_));
INVX1 INVX1_3941 ( .A(u2__abc_52155_new_n21421_), .Y(u2__abc_52155_new_n21422_));
INVX1 INVX1_3942 ( .A(u2__abc_52155_new_n21426_), .Y(u2__abc_52155_new_n21427_));
INVX1 INVX1_3943 ( .A(u2__abc_52155_new_n21434_), .Y(u2__abc_52155_new_n21435_));
INVX1 INVX1_3944 ( .A(u2__abc_52155_new_n21438_), .Y(u2__abc_52155_new_n21439_));
INVX1 INVX1_3945 ( .A(u2__abc_52155_new_n21445_), .Y(u2__abc_52155_new_n21446_));
INVX1 INVX1_3946 ( .A(u2__abc_52155_new_n21450_), .Y(u2__abc_52155_new_n21451_));
INVX1 INVX1_3947 ( .A(u2__abc_52155_new_n21458_), .Y(u2__abc_52155_new_n21459_));
INVX1 INVX1_3948 ( .A(u2__abc_52155_new_n21462_), .Y(u2__abc_52155_new_n21463_));
INVX1 INVX1_3949 ( .A(u2__abc_52155_new_n21470_), .Y(u2__abc_52155_new_n21471_));
INVX1 INVX1_395 ( .A(u2_remHi_33_), .Y(u2__abc_52155_new_n3514_));
INVX1 INVX1_3950 ( .A(u2__abc_52155_new_n21474_), .Y(u2__abc_52155_new_n21475_));
INVX1 INVX1_3951 ( .A(u2__abc_52155_new_n21482_), .Y(u2__abc_52155_new_n21483_));
INVX1 INVX1_3952 ( .A(u2__abc_52155_new_n21486_), .Y(u2__abc_52155_new_n21487_));
INVX1 INVX1_3953 ( .A(u2__abc_52155_new_n21493_), .Y(u2__abc_52155_new_n21494_));
INVX1 INVX1_3954 ( .A(u2__abc_52155_new_n21498_), .Y(u2__abc_52155_new_n21499_));
INVX1 INVX1_3955 ( .A(u2__abc_52155_new_n21506_), .Y(u2__abc_52155_new_n21507_));
INVX1 INVX1_3956 ( .A(u2__abc_52155_new_n21510_), .Y(u2__abc_52155_new_n21511_));
INVX1 INVX1_3957 ( .A(u2__abc_52155_new_n21518_), .Y(u2__abc_52155_new_n21519_));
INVX1 INVX1_3958 ( .A(u2__abc_52155_new_n21522_), .Y(u2__abc_52155_new_n21523_));
INVX1 INVX1_3959 ( .A(u2__abc_52155_new_n21530_), .Y(u2__abc_52155_new_n21531_));
INVX1 INVX1_396 ( .A(u2__abc_52155_new_n3517_), .Y(u2__abc_52155_new_n3518_));
INVX1 INVX1_3960 ( .A(u2__abc_52155_new_n21534_), .Y(u2__abc_52155_new_n21535_));
INVX1 INVX1_3961 ( .A(u2__abc_52155_new_n21541_), .Y(u2__abc_52155_new_n21542_));
INVX1 INVX1_3962 ( .A(u2__abc_52155_new_n21546_), .Y(u2__abc_52155_new_n21547_));
INVX1 INVX1_3963 ( .A(u2__abc_52155_new_n21554_), .Y(u2__abc_52155_new_n21555_));
INVX1 INVX1_3964 ( .A(u2__abc_52155_new_n21558_), .Y(u2__abc_52155_new_n21559_));
INVX1 INVX1_3965 ( .A(u2__abc_52155_new_n21566_), .Y(u2__abc_52155_new_n21567_));
INVX1 INVX1_3966 ( .A(u2__abc_52155_new_n21570_), .Y(u2__abc_52155_new_n21571_));
INVX1 INVX1_3967 ( .A(u2__abc_52155_new_n21578_), .Y(u2__abc_52155_new_n21579_));
INVX1 INVX1_3968 ( .A(u2__abc_52155_new_n21582_), .Y(u2__abc_52155_new_n21583_));
INVX1 INVX1_3969 ( .A(u2__abc_52155_new_n21589_), .Y(u2__abc_52155_new_n21590_));
INVX1 INVX1_397 ( .A(sqrto_30_), .Y(u2__abc_52155_new_n3519_));
INVX1 INVX1_3970 ( .A(u2__abc_52155_new_n21594_), .Y(u2__abc_52155_new_n21595_));
INVX1 INVX1_3971 ( .A(u2__abc_52155_new_n21602_), .Y(u2__abc_52155_new_n21603_));
INVX1 INVX1_3972 ( .A(u2__abc_52155_new_n21606_), .Y(u2__abc_52155_new_n21607_));
INVX1 INVX1_3973 ( .A(u2__abc_52155_new_n21614_), .Y(u2__abc_52155_new_n21615_));
INVX1 INVX1_3974 ( .A(u2__abc_52155_new_n21618_), .Y(u2__abc_52155_new_n21619_));
INVX1 INVX1_3975 ( .A(u2__abc_52155_new_n21626_), .Y(u2__abc_52155_new_n21627_));
INVX1 INVX1_3976 ( .A(u2__abc_52155_new_n21630_), .Y(u2__abc_52155_new_n21631_));
INVX1 INVX1_3977 ( .A(u2__abc_52155_new_n21637_), .Y(u2__abc_52155_new_n21638_));
INVX1 INVX1_3978 ( .A(u2__abc_52155_new_n21642_), .Y(u2__abc_52155_new_n21643_));
INVX1 INVX1_3979 ( .A(u2__abc_52155_new_n21650_), .Y(u2__abc_52155_new_n21651_));
INVX1 INVX1_398 ( .A(u2__abc_52155_new_n3520_), .Y(u2__abc_52155_new_n3521_));
INVX1 INVX1_3980 ( .A(u2__abc_52155_new_n21654_), .Y(u2__abc_52155_new_n21655_));
INVX1 INVX1_3981 ( .A(u2__abc_52155_new_n21662_), .Y(u2__abc_52155_new_n21663_));
INVX1 INVX1_3982 ( .A(u2__abc_52155_new_n21666_), .Y(u2__abc_52155_new_n21667_));
INVX1 INVX1_3983 ( .A(u2__abc_52155_new_n21674_), .Y(u2__abc_52155_new_n21675_));
INVX1 INVX1_3984 ( .A(u2__abc_52155_new_n21678_), .Y(u2__abc_52155_new_n21679_));
INVX1 INVX1_3985 ( .A(u2__abc_52155_new_n21685_), .Y(u2__abc_52155_new_n21686_));
INVX1 INVX1_3986 ( .A(u2__abc_52155_new_n21690_), .Y(u2__abc_52155_new_n21691_));
INVX1 INVX1_3987 ( .A(u2__abc_52155_new_n21698_), .Y(u2__abc_52155_new_n21699_));
INVX1 INVX1_3988 ( .A(u2__abc_52155_new_n21702_), .Y(u2__abc_52155_new_n21703_));
INVX1 INVX1_3989 ( .A(u2__abc_52155_new_n21710_), .Y(u2__abc_52155_new_n21711_));
INVX1 INVX1_399 ( .A(sqrto_31_), .Y(u2__abc_52155_new_n3524_));
INVX1 INVX1_3990 ( .A(u2__abc_52155_new_n21714_), .Y(u2__abc_52155_new_n21715_));
INVX1 INVX1_3991 ( .A(u2__abc_52155_new_n21722_), .Y(u2__abc_52155_new_n21723_));
INVX1 INVX1_3992 ( .A(u2__abc_52155_new_n21726_), .Y(u2__abc_52155_new_n21727_));
INVX1 INVX1_3993 ( .A(u2__abc_52155_new_n21733_), .Y(u2__abc_52155_new_n21734_));
INVX1 INVX1_3994 ( .A(u2__abc_52155_new_n21738_), .Y(u2__abc_52155_new_n21739_));
INVX1 INVX1_3995 ( .A(u2__abc_52155_new_n21746_), .Y(u2__abc_52155_new_n21747_));
INVX1 INVX1_3996 ( .A(u2__abc_52155_new_n21750_), .Y(u2__abc_52155_new_n21751_));
INVX1 INVX1_3997 ( .A(u2__abc_52155_new_n21757_), .Y(u2__abc_52155_new_n21758_));
INVX1 INVX1_3998 ( .A(u2__abc_52155_new_n21762_), .Y(u2__abc_52155_new_n21763_));
INVX1 INVX1_3999 ( .A(u2__abc_52155_new_n21770_), .Y(u2__abc_52155_new_n21771_));
INVX1 INVX1_4 ( .A(\a[114] ), .Y(_abc_73687_new_n1516_));
INVX1 INVX1_40 ( .A(\a[124] ), .Y(_abc_73687_new_n1643_));
INVX1 INVX1_400 ( .A(u2__abc_52155_new_n3525_), .Y(u2__abc_52155_new_n3526_));
INVX1 INVX1_4000 ( .A(u2__abc_52155_new_n21774_), .Y(u2__abc_52155_new_n21775_));
INVX1 INVX1_4001 ( .A(u2__abc_52155_new_n21781_), .Y(u2__abc_52155_new_n21782_));
INVX1 INVX1_4002 ( .A(u2__abc_52155_new_n21786_), .Y(u2__abc_52155_new_n21787_));
INVX1 INVX1_4003 ( .A(u2__abc_52155_new_n21794_), .Y(u2__abc_52155_new_n21795_));
INVX1 INVX1_4004 ( .A(u2__abc_52155_new_n21798_), .Y(u2__abc_52155_new_n21799_));
INVX1 INVX1_4005 ( .A(u2__abc_52155_new_n21806_), .Y(u2__abc_52155_new_n21807_));
INVX1 INVX1_4006 ( .A(u2__abc_52155_new_n21810_), .Y(u2__abc_52155_new_n21811_));
INVX1 INVX1_4007 ( .A(u2__abc_52155_new_n21818_), .Y(u2__abc_52155_new_n21819_));
INVX1 INVX1_4008 ( .A(u2__abc_52155_new_n21822_), .Y(u2__abc_52155_new_n21823_));
INVX1 INVX1_4009 ( .A(u2__abc_52155_new_n21829_), .Y(u2__abc_52155_new_n21830_));
INVX1 INVX1_401 ( .A(u2_remHi_31_), .Y(u2__abc_52155_new_n3527_));
INVX1 INVX1_4010 ( .A(u2__abc_52155_new_n21834_), .Y(u2__abc_52155_new_n21835_));
INVX1 INVX1_4011 ( .A(u2__abc_52155_new_n21842_), .Y(u2__abc_52155_new_n21843_));
INVX1 INVX1_4012 ( .A(u2__abc_52155_new_n21846_), .Y(u2__abc_52155_new_n21847_));
INVX1 INVX1_4013 ( .A(u2__abc_52155_new_n21854_), .Y(u2__abc_52155_new_n21855_));
INVX1 INVX1_4014 ( .A(u2__abc_52155_new_n21858_), .Y(u2__abc_52155_new_n21859_));
INVX1 INVX1_4015 ( .A(u2__abc_52155_new_n21866_), .Y(u2__abc_52155_new_n21867_));
INVX1 INVX1_4016 ( .A(u2__abc_52155_new_n21870_), .Y(u2__abc_52155_new_n21871_));
INVX1 INVX1_4017 ( .A(u2__abc_52155_new_n21877_), .Y(u2__abc_52155_new_n21878_));
INVX1 INVX1_4018 ( .A(u2__abc_52155_new_n21882_), .Y(u2__abc_52155_new_n21883_));
INVX1 INVX1_4019 ( .A(u2__abc_52155_new_n21890_), .Y(u2__abc_52155_new_n21891_));
INVX1 INVX1_402 ( .A(u2__abc_52155_new_n3528_), .Y(u2__abc_52155_new_n3529_));
INVX1 INVX1_4020 ( .A(u2__abc_52155_new_n21894_), .Y(u2__abc_52155_new_n21895_));
INVX1 INVX1_4021 ( .A(u2__abc_52155_new_n21902_), .Y(u2__abc_52155_new_n21903_));
INVX1 INVX1_4022 ( .A(u2__abc_52155_new_n21906_), .Y(u2__abc_52155_new_n21907_));
INVX1 INVX1_4023 ( .A(u2__abc_52155_new_n21914_), .Y(u2__abc_52155_new_n21915_));
INVX1 INVX1_4024 ( .A(u2__abc_52155_new_n21918_), .Y(u2__abc_52155_new_n21919_));
INVX1 INVX1_4025 ( .A(u2__abc_52155_new_n21925_), .Y(u2__abc_52155_new_n21926_));
INVX1 INVX1_4026 ( .A(u2__abc_52155_new_n21930_), .Y(u2__abc_52155_new_n21931_));
INVX1 INVX1_4027 ( .A(u2__abc_52155_new_n21938_), .Y(u2__abc_52155_new_n21939_));
INVX1 INVX1_4028 ( .A(u2__abc_52155_new_n21942_), .Y(u2__abc_52155_new_n21943_));
INVX1 INVX1_4029 ( .A(u2__abc_52155_new_n21949_), .Y(u2__abc_52155_new_n21950_));
INVX1 INVX1_403 ( .A(sqrto_36_), .Y(u2__abc_52155_new_n3533_));
INVX1 INVX1_4030 ( .A(u2__abc_52155_new_n21954_), .Y(u2__abc_52155_new_n21955_));
INVX1 INVX1_4031 ( .A(u2__abc_52155_new_n21962_), .Y(u2__abc_52155_new_n21963_));
INVX1 INVX1_4032 ( .A(u2__abc_52155_new_n21966_), .Y(u2__abc_52155_new_n21967_));
INVX1 INVX1_4033 ( .A(u2__abc_52155_new_n21973_), .Y(u2__abc_52155_new_n21974_));
INVX1 INVX1_4034 ( .A(u2__abc_52155_new_n21978_), .Y(u2__abc_52155_new_n21979_));
INVX1 INVX1_4035 ( .A(u2__abc_52155_new_n21986_), .Y(u2__abc_52155_new_n21987_));
INVX1 INVX1_4036 ( .A(u2__abc_52155_new_n21990_), .Y(u2__abc_52155_new_n21991_));
INVX1 INVX1_4037 ( .A(u2__abc_52155_new_n21998_), .Y(u2__abc_52155_new_n21999_));
INVX1 INVX1_4038 ( .A(u2__abc_52155_new_n22002_), .Y(u2__abc_52155_new_n22003_));
INVX1 INVX1_4039 ( .A(u2__abc_52155_new_n22010_), .Y(u2__abc_52155_new_n22011_));
INVX1 INVX1_404 ( .A(u2_remHi_36_), .Y(u2__abc_52155_new_n3535_));
INVX1 INVX1_4040 ( .A(u2__abc_52155_new_n22014_), .Y(u2__abc_52155_new_n22015_));
INVX1 INVX1_4041 ( .A(u2__abc_52155_new_n22021_), .Y(u2__abc_52155_new_n22022_));
INVX1 INVX1_4042 ( .A(u2__abc_52155_new_n22026_), .Y(u2__abc_52155_new_n22027_));
INVX1 INVX1_4043 ( .A(u2__abc_52155_new_n22034_), .Y(u2__abc_52155_new_n22035_));
INVX1 INVX1_4044 ( .A(u2__abc_52155_new_n22038_), .Y(u2__abc_52155_new_n22039_));
INVX1 INVX1_4045 ( .A(u2__abc_52155_new_n22045_), .Y(u2__abc_52155_new_n22046_));
INVX1 INVX1_4046 ( .A(u2__abc_52155_new_n22050_), .Y(u2__abc_52155_new_n22051_));
INVX1 INVX1_4047 ( .A(u2__abc_52155_new_n22058_), .Y(u2__abc_52155_new_n22059_));
INVX1 INVX1_4048 ( .A(u2__abc_52155_new_n22062_), .Y(u2__abc_52155_new_n22063_));
INVX1 INVX1_4049 ( .A(u2__abc_52155_new_n22069_), .Y(u2__abc_52155_new_n22070_));
INVX1 INVX1_405 ( .A(sqrto_37_), .Y(u2__abc_52155_new_n3538_));
INVX1 INVX1_4050 ( .A(u2__abc_52155_new_n22074_), .Y(u2__abc_52155_new_n22075_));
INVX1 INVX1_4051 ( .A(u2__abc_52155_new_n22082_), .Y(u2__abc_52155_new_n22083_));
INVX1 INVX1_4052 ( .A(u2__abc_52155_new_n22086_), .Y(u2__abc_52155_new_n22087_));
INVX1 INVX1_4053 ( .A(u2__abc_52155_new_n22093_), .Y(u2__abc_52155_new_n22094_));
INVX1 INVX1_4054 ( .A(u2__abc_52155_new_n22098_), .Y(u2__abc_52155_new_n22099_));
INVX1 INVX1_4055 ( .A(u2__abc_52155_new_n22106_), .Y(u2__abc_52155_new_n22107_));
INVX1 INVX1_4056 ( .A(u2__abc_52155_new_n22110_), .Y(u2__abc_52155_new_n22111_));
INVX1 INVX1_4057 ( .A(u2__abc_52155_new_n22117_), .Y(u2__abc_52155_new_n22118_));
INVX1 INVX1_4058 ( .A(u2__abc_52155_new_n22122_), .Y(u2__abc_52155_new_n22123_));
INVX1 INVX1_4059 ( .A(u2__abc_52155_new_n22130_), .Y(u2__abc_52155_new_n22131_));
INVX1 INVX1_406 ( .A(u2_remHi_37_), .Y(u2__abc_52155_new_n3540_));
INVX1 INVX1_4060 ( .A(u2__abc_52155_new_n22134_), .Y(u2__abc_52155_new_n22135_));
INVX1 INVX1_4061 ( .A(u2__abc_52155_new_n22141_), .Y(u2__abc_52155_new_n22142_));
INVX1 INVX1_4062 ( .A(u2__abc_52155_new_n22146_), .Y(u2__abc_52155_new_n22147_));
INVX1 INVX1_4063 ( .A(u2__abc_52155_new_n22154_), .Y(u2__abc_52155_new_n22155_));
INVX1 INVX1_4064 ( .A(u2__abc_52155_new_n22158_), .Y(u2__abc_52155_new_n22159_));
INVX1 INVX1_4065 ( .A(u2__abc_52155_new_n22166_), .Y(u2__abc_52155_new_n22167_));
INVX1 INVX1_4066 ( .A(u2__abc_52155_new_n22170_), .Y(u2__abc_52155_new_n22171_));
INVX1 INVX1_4067 ( .A(u2__abc_52155_new_n22178_), .Y(u2__abc_52155_new_n22179_));
INVX1 INVX1_4068 ( .A(u2__abc_52155_new_n22182_), .Y(u2__abc_52155_new_n22183_));
INVX1 INVX1_4069 ( .A(u2__abc_52155_new_n22189_), .Y(u2__abc_52155_new_n22190_));
INVX1 INVX1_407 ( .A(sqrto_35_), .Y(u2__abc_52155_new_n3544_));
INVX1 INVX1_4070 ( .A(u2__abc_52155_new_n22194_), .Y(u2__abc_52155_new_n22195_));
INVX1 INVX1_4071 ( .A(u2__abc_52155_new_n22202_), .Y(u2__abc_52155_new_n22203_));
INVX1 INVX1_4072 ( .A(u2__abc_52155_new_n22206_), .Y(u2__abc_52155_new_n22207_));
INVX1 INVX1_4073 ( .A(u2__abc_52155_new_n22213_), .Y(u2__abc_52155_new_n22214_));
INVX1 INVX1_4074 ( .A(u2__abc_52155_new_n22218_), .Y(u2__abc_52155_new_n22219_));
INVX1 INVX1_4075 ( .A(u2__abc_52155_new_n22226_), .Y(u2__abc_52155_new_n22227_));
INVX1 INVX1_4076 ( .A(u2__abc_52155_new_n22230_), .Y(u2__abc_52155_new_n22231_));
INVX1 INVX1_4077 ( .A(u2__abc_52155_new_n22238_), .Y(u2__abc_52155_new_n22239_));
INVX1 INVX1_4078 ( .A(u2__abc_52155_new_n22242_), .Y(u2__abc_52155_new_n22243_));
INVX1 INVX1_4079 ( .A(u2__abc_52155_new_n22250_), .Y(u2__abc_52155_new_n22251_));
INVX1 INVX1_408 ( .A(u2_remHi_35_), .Y(u2__abc_52155_new_n3546_));
INVX1 INVX1_4080 ( .A(u2__abc_52155_new_n22254_), .Y(u2__abc_52155_new_n22255_));
INVX1 INVX1_4081 ( .A(u2__abc_52155_new_n22261_), .Y(u2__abc_52155_new_n22262_));
INVX1 INVX1_4082 ( .A(u2__abc_52155_new_n22266_), .Y(u2__abc_52155_new_n22267_));
INVX1 INVX1_4083 ( .A(u2__abc_52155_new_n22274_), .Y(u2__abc_52155_new_n22275_));
INVX1 INVX1_4084 ( .A(u2__abc_52155_new_n22278_), .Y(u2__abc_52155_new_n22279_));
INVX1 INVX1_4085 ( .A(u2__abc_52155_new_n22286_), .Y(u2__abc_52155_new_n22287_));
INVX1 INVX1_4086 ( .A(u2__abc_52155_new_n22290_), .Y(u2__abc_52155_new_n22291_));
INVX1 INVX1_4087 ( .A(u2__abc_52155_new_n22298_), .Y(u2__abc_52155_new_n22299_));
INVX1 INVX1_4088 ( .A(u2__abc_52155_new_n22302_), .Y(u2__abc_52155_new_n22303_));
INVX1 INVX1_4089 ( .A(u2__abc_52155_new_n22309_), .Y(u2__abc_52155_new_n22310_));
INVX1 INVX1_409 ( .A(sqrto_34_), .Y(u2__abc_52155_new_n3549_));
INVX1 INVX1_4090 ( .A(u2__abc_52155_new_n22314_), .Y(u2__abc_52155_new_n22315_));
INVX1 INVX1_4091 ( .A(u2__abc_52155_new_n22322_), .Y(u2__abc_52155_new_n22323_));
INVX1 INVX1_4092 ( .A(u2__abc_52155_new_n22326_), .Y(u2__abc_52155_new_n22327_));
INVX1 INVX1_4093 ( .A(u2__abc_52155_new_n22334_), .Y(u2__abc_52155_new_n22335_));
INVX1 INVX1_4094 ( .A(u2__abc_52155_new_n22338_), .Y(u2__abc_52155_new_n22339_));
INVX1 INVX1_4095 ( .A(u2__abc_52155_new_n22346_), .Y(u2__abc_52155_new_n22347_));
INVX1 INVX1_4096 ( .A(u2__abc_52155_new_n22350_), .Y(u2__abc_52155_new_n22351_));
INVX1 INVX1_4097 ( .A(u2__abc_52155_new_n22357_), .Y(u2__abc_52155_new_n22358_));
INVX1 INVX1_4098 ( .A(u2__abc_52155_new_n22362_), .Y(u2__abc_52155_new_n22363_));
INVX1 INVX1_4099 ( .A(u2__abc_52155_new_n22370_), .Y(u2__abc_52155_new_n22371_));
INVX1 INVX1_41 ( .A(_abc_73687_new_n1644_), .Y(_abc_73687_new_n1645_));
INVX1 INVX1_410 ( .A(u2_remHi_34_), .Y(u2__abc_52155_new_n3551_));
INVX1 INVX1_4100 ( .A(u2__abc_52155_new_n22374_), .Y(u2__abc_52155_new_n22375_));
INVX1 INVX1_4101 ( .A(u2__abc_52155_new_n22382_), .Y(u2__abc_52155_new_n22383_));
INVX1 INVX1_4102 ( .A(u2__abc_52155_new_n22386_), .Y(u2__abc_52155_new_n22387_));
INVX1 INVX1_4103 ( .A(u2__abc_52155_new_n22394_), .Y(u2__abc_52155_new_n22395_));
INVX1 INVX1_4104 ( .A(u2__abc_52155_new_n22398_), .Y(u2__abc_52155_new_n22399_));
INVX1 INVX1_4105 ( .A(u2__abc_52155_new_n22405_), .Y(u2__abc_52155_new_n22406_));
INVX1 INVX1_4106 ( .A(u2__abc_52155_new_n22410_), .Y(u2__abc_52155_new_n22411_));
INVX1 INVX1_4107 ( .A(u2__abc_52155_new_n22418_), .Y(u2__abc_52155_new_n22419_));
INVX1 INVX1_4108 ( .A(u2__abc_52155_new_n22422_), .Y(u2__abc_52155_new_n22423_));
INVX1 INVX1_4109 ( .A(u2__abc_52155_new_n22430_), .Y(u2__abc_52155_new_n22431_));
INVX1 INVX1_411 ( .A(u2__abc_52155_new_n3555_), .Y(u2__abc_52155_new_n3556_));
INVX1 INVX1_4110 ( .A(u2__abc_52155_new_n22434_), .Y(u2__abc_52155_new_n22435_));
INVX1 INVX1_4111 ( .A(u2__abc_52155_new_n22442_), .Y(u2__abc_52155_new_n22443_));
INVX1 INVX1_4112 ( .A(u2__abc_52155_new_n22446_), .Y(u2__abc_52155_new_n22447_));
INVX1 INVX1_4113 ( .A(u2__abc_52155_new_n22453_), .Y(u2__abc_52155_new_n22454_));
INVX1 INVX1_4114 ( .A(u2__abc_52155_new_n22458_), .Y(u2__abc_52155_new_n22459_));
INVX1 INVX1_4115 ( .A(u2__abc_52155_new_n22466_), .Y(u2__abc_52155_new_n22467_));
INVX1 INVX1_4116 ( .A(u2__abc_52155_new_n22470_), .Y(u2__abc_52155_new_n22471_));
INVX1 INVX1_4117 ( .A(u2__abc_52155_new_n22478_), .Y(u2__abc_52155_new_n22479_));
INVX1 INVX1_4118 ( .A(u2__abc_52155_new_n22482_), .Y(u2__abc_52155_new_n22483_));
INVX1 INVX1_4119 ( .A(u2__abc_52155_new_n22490_), .Y(u2__abc_52155_new_n22491_));
INVX1 INVX1_412 ( .A(u2__abc_52155_new_n3559_), .Y(u2__abc_52155_new_n3560_));
INVX1 INVX1_4120 ( .A(u2__abc_52155_new_n22494_), .Y(u2__abc_52155_new_n22495_));
INVX1 INVX1_4121 ( .A(u2__abc_52155_new_n22501_), .Y(u2__abc_52155_new_n22502_));
INVX1 INVX1_4122 ( .A(u2__abc_52155_new_n22506_), .Y(u2__abc_52155_new_n22507_));
INVX1 INVX1_4123 ( .A(u2__abc_52155_new_n22514_), .Y(u2__abc_52155_new_n22515_));
INVX1 INVX1_4124 ( .A(u2__abc_52155_new_n22518_), .Y(u2__abc_52155_new_n22519_));
INVX1 INVX1_4125 ( .A(u2__abc_52155_new_n22525_), .Y(u2__abc_52155_new_n22526_));
INVX1 INVX1_4126 ( .A(u2__abc_52155_new_n22530_), .Y(u2__abc_52155_new_n22531_));
INVX1 INVX1_4127 ( .A(u2__abc_52155_new_n22538_), .Y(u2__abc_52155_new_n22539_));
INVX1 INVX1_4128 ( .A(u2__abc_52155_new_n22542_), .Y(u2__abc_52155_new_n22543_));
INVX1 INVX1_4129 ( .A(u2__abc_52155_new_n22549_), .Y(u2__abc_52155_new_n22550_));
INVX1 INVX1_413 ( .A(u2__abc_52155_new_n3446_), .Y(u2__abc_52155_new_n3562_));
INVX1 INVX1_4130 ( .A(u2__abc_52155_new_n22554_), .Y(u2__abc_52155_new_n22555_));
INVX1 INVX1_4131 ( .A(u2__abc_52155_new_n22562_), .Y(u2__abc_52155_new_n22563_));
INVX1 INVX1_4132 ( .A(u2__abc_52155_new_n22566_), .Y(u2__abc_52155_new_n22567_));
INVX1 INVX1_4133 ( .A(u2__abc_52155_new_n22574_), .Y(u2__abc_52155_new_n22575_));
INVX1 INVX1_4134 ( .A(u2__abc_52155_new_n22578_), .Y(u2__abc_52155_new_n22579_));
INVX1 INVX1_4135 ( .A(u2__abc_52155_new_n22586_), .Y(u2__abc_52155_new_n22587_));
INVX1 INVX1_4136 ( .A(u2__abc_52155_new_n22590_), .Y(u2__abc_52155_new_n22591_));
INVX1 INVX1_4137 ( .A(u2__abc_52155_new_n22597_), .Y(u2__abc_52155_new_n22598_));
INVX1 INVX1_4138 ( .A(u2__abc_52155_new_n22602_), .Y(u2__abc_52155_new_n22603_));
INVX1 INVX1_4139 ( .A(u2__abc_52155_new_n22610_), .Y(u2__abc_52155_new_n22611_));
INVX1 INVX1_414 ( .A(u2__abc_52155_new_n3506_), .Y(u2__abc_52155_new_n3563_));
INVX1 INVX1_4140 ( .A(u2__abc_52155_new_n22614_), .Y(u2__abc_52155_new_n22615_));
INVX1 INVX1_4141 ( .A(u2__abc_52155_new_n22622_), .Y(u2__abc_52155_new_n22623_));
INVX1 INVX1_4142 ( .A(u2__abc_52155_new_n22626_), .Y(u2__abc_52155_new_n22627_));
INVX1 INVX1_4143 ( .A(u2__abc_52155_new_n22634_), .Y(u2__abc_52155_new_n22635_));
INVX1 INVX1_4144 ( .A(u2__abc_52155_new_n22638_), .Y(u2__abc_52155_new_n22639_));
INVX1 INVX1_4145 ( .A(u2__abc_52155_new_n22645_), .Y(u2__abc_52155_new_n22646_));
INVX1 INVX1_4146 ( .A(u2__abc_52155_new_n22650_), .Y(u2__abc_52155_new_n22651_));
INVX1 INVX1_4147 ( .A(u2__abc_52155_new_n22658_), .Y(u2__abc_52155_new_n22659_));
INVX1 INVX1_4148 ( .A(u2__abc_52155_new_n22662_), .Y(u2__abc_52155_new_n22663_));
INVX1 INVX1_4149 ( .A(u2__abc_52155_new_n22670_), .Y(u2__abc_52155_new_n22671_));
INVX1 INVX1_415 ( .A(u2__abc_52155_new_n3515_), .Y(u2__abc_52155_new_n3567_));
INVX1 INVX1_4150 ( .A(u2__abc_52155_new_n22674_), .Y(u2__abc_52155_new_n22675_));
INVX1 INVX1_4151 ( .A(u2__abc_52155_new_n22682_), .Y(u2__abc_52155_new_n22683_));
INVX1 INVX1_4152 ( .A(u2__abc_52155_new_n22686_), .Y(u2__abc_52155_new_n22687_));
INVX1 INVX1_4153 ( .A(u2__abc_52155_new_n22693_), .Y(u2__abc_52155_new_n22694_));
INVX1 INVX1_4154 ( .A(u2__abc_52155_new_n22698_), .Y(u2__abc_52155_new_n22699_));
INVX1 INVX1_4155 ( .A(u2__abc_52155_new_n22706_), .Y(u2__abc_52155_new_n22707_));
INVX1 INVX1_4156 ( .A(u2__abc_52155_new_n22710_), .Y(u2__abc_52155_new_n22711_));
INVX1 INVX1_4157 ( .A(u2__abc_52155_new_n22717_), .Y(u2__abc_52155_new_n22718_));
INVX1 INVX1_4158 ( .A(u2__abc_52155_new_n22722_), .Y(u2__abc_52155_new_n22723_));
INVX1 INVX1_4159 ( .A(u2__abc_52155_new_n22730_), .Y(u2__abc_52155_new_n22731_));
INVX1 INVX1_416 ( .A(u2__abc_52155_new_n3510_), .Y(u2__abc_52155_new_n3568_));
INVX1 INVX1_4160 ( .A(u2__abc_52155_new_n22734_), .Y(u2__abc_52155_new_n22735_));
INVX1 INVX1_4161 ( .A(u2__abc_52155_new_n22741_), .Y(u2__abc_52155_new_n22742_));
INVX1 INVX1_4162 ( .A(u2__abc_52155_new_n22746_), .Y(u2__abc_52155_new_n22747_));
INVX1 INVX1_4163 ( .A(u2__abc_52155_new_n22754_), .Y(u2__abc_52155_new_n22755_));
INVX1 INVX1_4164 ( .A(u2__abc_52155_new_n22758_), .Y(u2__abc_52155_new_n22759_));
INVX1 INVX1_4165 ( .A(u2__abc_52155_new_n22766_), .Y(u2__abc_52155_new_n22767_));
INVX1 INVX1_4166 ( .A(u2__abc_52155_new_n22770_), .Y(u2__abc_52155_new_n22771_));
INVX1 INVX1_4167 ( .A(u2__abc_52155_new_n22778_), .Y(u2__abc_52155_new_n22779_));
INVX1 INVX1_4168 ( .A(u2__abc_52155_new_n22782_), .Y(u2__abc_52155_new_n22783_));
INVX1 INVX1_4169 ( .A(u2__abc_52155_new_n22789_), .Y(u2__abc_52155_new_n22790_));
INVX1 INVX1_417 ( .A(u2__abc_52155_new_n3547_), .Y(u2__abc_52155_new_n3573_));
INVX1 INVX1_4170 ( .A(u2__abc_52155_new_n22794_), .Y(u2__abc_52155_new_n22795_));
INVX1 INVX1_4171 ( .A(u2__abc_52155_new_n22802_), .Y(u2__abc_52155_new_n22803_));
INVX1 INVX1_4172 ( .A(u2__abc_52155_new_n22806_), .Y(u2__abc_52155_new_n22807_));
INVX1 INVX1_4173 ( .A(u2__abc_52155_new_n22813_), .Y(u2__abc_52155_new_n22814_));
INVX1 INVX1_4174 ( .A(u2__abc_52155_new_n22818_), .Y(u2__abc_52155_new_n22819_));
INVX1 INVX1_4175 ( .A(u2__abc_52155_new_n22826_), .Y(u2__abc_52155_new_n22827_));
INVX1 INVX1_4176 ( .A(u2__abc_52155_new_n22830_), .Y(u2__abc_52155_new_n22831_));
INVX1 INVX1_4177 ( .A(u2__abc_52155_new_n22837_), .Y(u2__abc_52155_new_n22838_));
INVX1 INVX1_4178 ( .A(u2__abc_52155_new_n22842_), .Y(u2__abc_52155_new_n22843_));
INVX1 INVX1_4179 ( .A(u2__abc_52155_new_n22850_), .Y(u2__abc_52155_new_n22851_));
INVX1 INVX1_418 ( .A(u2__abc_52155_new_n3552_), .Y(u2__abc_52155_new_n3574_));
INVX1 INVX1_4180 ( .A(u2__abc_52155_new_n22854_), .Y(u2__abc_52155_new_n22855_));
INVX1 INVX1_4181 ( .A(u2__abc_52155_new_n22861_), .Y(u2__abc_52155_new_n22862_));
INVX1 INVX1_4182 ( .A(u2__abc_52155_new_n22866_), .Y(u2__abc_52155_new_n22867_));
INVX1 INVX1_4183 ( .A(u2__abc_52155_new_n22874_), .Y(u2__abc_52155_new_n22875_));
INVX1 INVX1_4184 ( .A(u2__abc_52155_new_n22878_), .Y(u2__abc_52155_new_n22879_));
INVX1 INVX1_4185 ( .A(u2__abc_52155_new_n22885_), .Y(u2__abc_52155_new_n22886_));
INVX1 INVX1_4186 ( .A(u2__abc_52155_new_n22890_), .Y(u2__abc_52155_new_n22891_));
INVX1 INVX1_4187 ( .A(u2__abc_52155_new_n22898_), .Y(u2__abc_52155_new_n22899_));
INVX1 INVX1_4188 ( .A(u2__abc_52155_new_n22902_), .Y(u2__abc_52155_new_n22903_));
INVX1 INVX1_4189 ( .A(u2__abc_52155_new_n22909_), .Y(u2__abc_52155_new_n22910_));
INVX1 INVX1_419 ( .A(u2__abc_52155_new_n3539_), .Y(u2__abc_52155_new_n3578_));
INVX1 INVX1_4190 ( .A(u2__abc_52155_new_n22914_), .Y(u2__abc_52155_new_n22915_));
INVX1 INVX1_4191 ( .A(u2__abc_52155_new_n22922_), .Y(u2__abc_52155_new_n22923_));
INVX1 INVX1_4192 ( .A(u2__abc_52155_new_n22926_), .Y(u2__abc_52155_new_n22927_));
INVX1 INVX1_4193 ( .A(u2__abc_52155_new_n22933_), .Y(u2__abc_52155_new_n22934_));
INVX1 INVX1_4194 ( .A(u2__abc_52155_new_n22938_), .Y(u2__abc_52155_new_n22939_));
INVX1 INVX1_4195 ( .A(u2__abc_52155_new_n22946_), .Y(u2__abc_52155_new_n22947_));
INVX1 INVX1_4196 ( .A(u2__abc_52155_new_n22950_), .Y(u2__abc_52155_new_n22951_));
INVX1 INVX1_4197 ( .A(u2__abc_52155_new_n22958_), .Y(u2__abc_52155_new_n22959_));
INVX1 INVX1_4198 ( .A(u2__abc_52155_new_n22962_), .Y(u2__abc_52155_new_n22963_));
INVX1 INVX1_4199 ( .A(u2__abc_52155_new_n22970_), .Y(u2__abc_52155_new_n22971_));
INVX1 INVX1_42 ( .A(_abc_73687_new_n1637_), .Y(_abc_73687_new_n1649_));
INVX1 INVX1_420 ( .A(u2__abc_52155_new_n3580_), .Y(u2__abc_52155_new_n3581_));
INVX1 INVX1_4200 ( .A(u2__abc_52155_new_n22974_), .Y(u2__abc_52155_new_n22975_));
INVX1 INVX1_4201 ( .A(u2__abc_52155_new_n22981_), .Y(u2__abc_52155_new_n22982_));
INVX1 INVX1_4202 ( .A(u2__abc_52155_new_n22986_), .Y(u2__abc_52155_new_n22987_));
INVX1 INVX1_4203 ( .A(u2__abc_52155_new_n22994_), .Y(u2__abc_52155_new_n22995_));
INVX1 INVX1_4204 ( .A(u2__abc_52155_new_n22998_), .Y(u2__abc_52155_new_n22999_));
INVX1 INVX1_4205 ( .A(u2__abc_52155_new_n23006_), .Y(u2__abc_52155_new_n23007_));
INVX1 INVX1_4206 ( .A(u2__abc_52155_new_n23010_), .Y(u2__abc_52155_new_n23011_));
INVX1 INVX1_4207 ( .A(u2__abc_52155_new_n23018_), .Y(u2__abc_52155_new_n23019_));
INVX1 INVX1_4208 ( .A(u2__abc_52155_new_n23022_), .Y(u2__abc_52155_new_n23023_));
INVX1 INVX1_4209 ( .A(u2__abc_52155_new_n23029_), .Y(u2__abc_52155_new_n23030_));
INVX1 INVX1_421 ( .A(u2__abc_52155_new_n3505_), .Y(u2__abc_52155_new_n3585_));
INVX1 INVX1_4210 ( .A(u2__abc_52155_new_n23034_), .Y(u2__abc_52155_new_n23035_));
INVX1 INVX1_4211 ( .A(u2__abc_52155_new_n23042_), .Y(u2__abc_52155_new_n23043_));
INVX1 INVX1_4212 ( .A(u2__abc_52155_new_n23046_), .Y(u2__abc_52155_new_n23047_));
INVX1 INVX1_4213 ( .A(u2__abc_52155_new_n23054_), .Y(u2__abc_52155_new_n23055_));
INVX1 INVX1_4214 ( .A(u2__abc_52155_new_n23058_), .Y(u2__abc_52155_new_n23059_));
INVX1 INVX1_4215 ( .A(u2__abc_52155_new_n23066_), .Y(u2__abc_52155_new_n23067_));
INVX1 INVX1_4216 ( .A(u2__abc_52155_new_n23070_), .Y(u2__abc_52155_new_n23071_));
INVX1 INVX1_4217 ( .A(u2__abc_52155_new_n23077_), .Y(u2__abc_52155_new_n23078_));
INVX1 INVX1_4218 ( .A(u2__abc_52155_new_n23082_), .Y(u2__abc_52155_new_n23083_));
INVX1 INVX1_4219 ( .A(u2__abc_52155_new_n23090_), .Y(u2__abc_52155_new_n23091_));
INVX1 INVX1_422 ( .A(u2__abc_52155_new_n3453_), .Y(u2__abc_52155_new_n3589_));
INVX1 INVX1_4220 ( .A(u2__abc_52155_new_n23094_), .Y(u2__abc_52155_new_n23095_));
INVX1 INVX1_4221 ( .A(u2__abc_52155_new_n23101_), .Y(u2__abc_52155_new_n23102_));
INVX1 INVX1_4222 ( .A(u2__abc_52155_new_n23106_), .Y(u2__abc_52155_new_n23107_));
INVX1 INVX1_4223 ( .A(u2__abc_52155_new_n23114_), .Y(u2__abc_52155_new_n23115_));
INVX1 INVX1_4224 ( .A(u2__abc_52155_new_n23118_), .Y(u2__abc_52155_new_n23119_));
INVX1 INVX1_4225 ( .A(u2__abc_52155_new_n23125_), .Y(u2__abc_52155_new_n23126_));
INVX1 INVX1_4226 ( .A(u2__abc_52155_new_n23130_), .Y(u2__abc_52155_new_n23131_));
INVX1 INVX1_4227 ( .A(u2__abc_52155_new_n23138_), .Y(u2__abc_52155_new_n23139_));
INVX1 INVX1_4228 ( .A(u2__abc_52155_new_n23142_), .Y(u2__abc_52155_new_n23143_));
INVX1 INVX1_4229 ( .A(u2__abc_52155_new_n23150_), .Y(u2__abc_52155_new_n23151_));
INVX1 INVX1_423 ( .A(u2__abc_52155_new_n3591_), .Y(u2__abc_52155_new_n3592_));
INVX1 INVX1_4230 ( .A(u2__abc_52155_new_n23154_), .Y(u2__abc_52155_new_n23155_));
INVX1 INVX1_4231 ( .A(u2__abc_52155_new_n23162_), .Y(u2__abc_52155_new_n23163_));
INVX1 INVX1_4232 ( .A(u2__abc_52155_new_n23166_), .Y(u2__abc_52155_new_n23167_));
INVX1 INVX1_4233 ( .A(u2__abc_52155_new_n23173_), .Y(u2__abc_52155_new_n23174_));
INVX1 INVX1_4234 ( .A(u2__abc_52155_new_n23178_), .Y(u2__abc_52155_new_n23179_));
INVX1 INVX1_4235 ( .A(u2__abc_52155_new_n23186_), .Y(u2__abc_52155_new_n23187_));
INVX1 INVX1_4236 ( .A(u2__abc_52155_new_n23190_), .Y(u2__abc_52155_new_n23191_));
INVX1 INVX1_4237 ( .A(u2__abc_52155_new_n23197_), .Y(u2__abc_52155_new_n23198_));
INVX1 INVX1_4238 ( .A(u2__abc_52155_new_n23202_), .Y(u2__abc_52155_new_n23203_));
INVX1 INVX1_4239 ( .A(u2__abc_52155_new_n23210_), .Y(u2__abc_52155_new_n23211_));
INVX1 INVX1_424 ( .A(u2__abc_52155_new_n3600_), .Y(u2__abc_52155_new_n3601_));
INVX1 INVX1_4240 ( .A(u2__abc_52155_new_n23214_), .Y(u2__abc_52155_new_n23215_));
INVX1 INVX1_4241 ( .A(u2__abc_52155_new_n23221_), .Y(u2__abc_52155_new_n23222_));
INVX1 INVX1_4242 ( .A(u2__abc_52155_new_n23226_), .Y(u2__abc_52155_new_n23227_));
INVX1 INVX1_4243 ( .A(u2__abc_52155_new_n23234_), .Y(u2__abc_52155_new_n23235_));
INVX1 INVX1_4244 ( .A(u2__abc_52155_new_n23238_), .Y(u2__abc_52155_new_n23239_));
INVX1 INVX1_4245 ( .A(u2__abc_52155_new_n23245_), .Y(u2__abc_52155_new_n23246_));
INVX1 INVX1_4246 ( .A(u2__abc_52155_new_n23250_), .Y(u2__abc_52155_new_n23251_));
INVX1 INVX1_4247 ( .A(u2__abc_52155_new_n23258_), .Y(u2__abc_52155_new_n23259_));
INVX1 INVX1_4248 ( .A(u2__abc_52155_new_n23262_), .Y(u2__abc_52155_new_n23263_));
INVX1 INVX1_4249 ( .A(u2__abc_52155_new_n23269_), .Y(u2__abc_52155_new_n23270_));
INVX1 INVX1_425 ( .A(u2__abc_52155_new_n3385_), .Y(u2__abc_52155_new_n3605_));
INVX1 INVX1_4250 ( .A(u2__abc_52155_new_n23274_), .Y(u2__abc_52155_new_n23275_));
INVX1 INVX1_4251 ( .A(u2__abc_52155_new_n23282_), .Y(u2__abc_52155_new_n23283_));
INVX1 INVX1_4252 ( .A(u2__abc_52155_new_n23286_), .Y(u2__abc_52155_new_n23287_));
INVX1 INVX1_4253 ( .A(u2__abc_52155_new_n23293_), .Y(u2__abc_52155_new_n23294_));
INVX1 INVX1_4254 ( .A(u2__abc_52155_new_n23298_), .Y(u2__abc_52155_new_n23299_));
INVX1 INVX1_4255 ( .A(u2__abc_52155_new_n23306_), .Y(u2__abc_52155_new_n23307_));
INVX1 INVX1_4256 ( .A(u2__abc_52155_new_n23310_), .Y(u2__abc_52155_new_n23311_));
INVX1 INVX1_4257 ( .A(u2__abc_52155_new_n23317_), .Y(u2__abc_52155_new_n23318_));
INVX1 INVX1_4258 ( .A(u2__abc_52155_new_n23322_), .Y(u2__abc_52155_new_n23323_));
INVX1 INVX1_4259 ( .A(u2__abc_52155_new_n23330_), .Y(u2__abc_52155_new_n23331_));
INVX1 INVX1_426 ( .A(u2__abc_52155_new_n3444_), .Y(u2__abc_52155_new_n3606_));
INVX1 INVX1_4260 ( .A(u2__abc_52155_new_n23334_), .Y(u2__abc_52155_new_n23335_));
INVX1 INVX1_4261 ( .A(u2__abc_52155_new_n23342_), .Y(u2__abc_52155_new_n23343_));
INVX1 INVX1_4262 ( .A(u2__abc_52155_new_n23346_), .Y(u2__abc_52155_new_n23347_));
INVX1 INVX1_4263 ( .A(u2__abc_52155_new_n23354_), .Y(u2__abc_52155_new_n23355_));
INVX1 INVX1_4264 ( .A(u2__abc_52155_new_n23358_), .Y(u2__abc_52155_new_n23359_));
INVX1 INVX1_4265 ( .A(u2__abc_52155_new_n23365_), .Y(u2__abc_52155_new_n23366_));
INVX1 INVX1_4266 ( .A(u2__abc_52155_new_n23370_), .Y(u2__abc_52155_new_n23371_));
INVX1 INVX1_4267 ( .A(u2__abc_52155_new_n23378_), .Y(u2__abc_52155_new_n23379_));
INVX1 INVX1_4268 ( .A(u2__abc_52155_new_n23382_), .Y(u2__abc_52155_new_n23383_));
INVX1 INVX1_4269 ( .A(u2__abc_52155_new_n23389_), .Y(u2__abc_52155_new_n23390_));
INVX1 INVX1_427 ( .A(u2__abc_52155_new_n3392_), .Y(u2__abc_52155_new_n3610_));
INVX1 INVX1_4270 ( .A(u2__abc_52155_new_n23394_), .Y(u2__abc_52155_new_n23395_));
INVX1 INVX1_4271 ( .A(u2__abc_52155_new_n23402_), .Y(u2__abc_52155_new_n23403_));
INVX1 INVX1_4272 ( .A(u2__abc_52155_new_n23406_), .Y(u2__abc_52155_new_n23407_));
INVX1 INVX1_4273 ( .A(u2__abc_52155_new_n23413_), .Y(u2__abc_52155_new_n23414_));
INVX1 INVX1_4274 ( .A(u2__abc_52155_new_n23418_), .Y(u2__abc_52155_new_n23419_));
INVX1 INVX1_4275 ( .A(u2__abc_52155_new_n23426_), .Y(u2__abc_52155_new_n23427_));
INVX1 INVX1_4276 ( .A(u2__abc_52155_new_n23430_), .Y(u2__abc_52155_new_n23431_));
INVX1 INVX1_4277 ( .A(u2__abc_52155_new_n23437_), .Y(u2__abc_52155_new_n23438_));
INVX1 INVX1_4278 ( .A(u2__abc_52155_new_n23442_), .Y(u2__abc_52155_new_n23443_));
INVX1 INVX1_4279 ( .A(u2__abc_52155_new_n23450_), .Y(u2__abc_52155_new_n23451_));
INVX1 INVX1_428 ( .A(u2__abc_52155_new_n3612_), .Y(u2__abc_52155_new_n3613_));
INVX1 INVX1_4280 ( .A(u2__abc_52155_new_n23454_), .Y(u2__abc_52155_new_n23455_));
INVX1 INVX1_4281 ( .A(u2__abc_52155_new_n23461_), .Y(u2__abc_52155_new_n23462_));
INVX1 INVX1_4282 ( .A(u2__abc_52155_new_n23466_), .Y(u2__abc_52155_new_n23467_));
INVX1 INVX1_4283 ( .A(u2__abc_52155_new_n23474_), .Y(u2__abc_52155_new_n23475_));
INVX1 INVX1_4284 ( .A(u2__abc_52155_new_n23478_), .Y(u2__abc_52155_new_n23479_));
INVX1 INVX1_4285 ( .A(u2__abc_52155_new_n23485_), .Y(u2__abc_52155_new_n23486_));
INVX1 INVX1_4286 ( .A(u2__abc_52155_new_n23490_), .Y(u2__abc_52155_new_n23491_));
INVX1 INVX1_4287 ( .A(u2__abc_52155_new_n23498_), .Y(u2__abc_52155_new_n23499_));
INVX1 INVX1_4288 ( .A(u2__abc_52155_new_n23502_), .Y(u2__abc_52155_new_n23503_));
INVX1 INVX1_4289 ( .A(u2__abc_52155_new_n23509_), .Y(u2__abc_52155_new_n23510_));
INVX1 INVX1_429 ( .A(u2__abc_52155_new_n3621_), .Y(u2__abc_52155_new_n3622_));
INVX1 INVX1_4290 ( .A(u2__abc_52155_new_n23514_), .Y(u2__abc_52155_new_n23515_));
INVX1 INVX1_4291 ( .A(u2__abc_52155_new_n23522_), .Y(u2__abc_52155_new_n23523_));
INVX1 INVX1_4292 ( .A(u2__abc_52155_new_n23526_), .Y(u2__abc_52155_new_n23527_));
INVX1 INVX1_4293 ( .A(u2__abc_52155_new_n23533_), .Y(u2__abc_52155_new_n23534_));
INVX1 INVX1_4294 ( .A(u2__abc_52155_new_n23538_), .Y(u2__abc_52155_new_n23539_));
INVX1 INVX1_4295 ( .A(u2__abc_52155_new_n23546_), .Y(u2__abc_52155_new_n23547_));
INVX1 INVX1_4296 ( .A(u2__abc_52155_new_n23550_), .Y(u2__abc_52155_new_n23551_));
INVX1 INVX1_4297 ( .A(u2__abc_52155_new_n23557_), .Y(u2__abc_52155_new_n23558_));
INVX1 INVX1_4298 ( .A(u2__abc_52155_new_n23562_), .Y(u2__abc_52155_new_n23563_));
INVX1 INVX1_4299 ( .A(u2__abc_52155_new_n23570_), .Y(u2__abc_52155_new_n23571_));
INVX1 INVX1_43 ( .A(_abc_73687_new_n1647_), .Y(_abc_73687_new_n1650_));
INVX1 INVX1_430 ( .A(u2__abc_52155_new_n3638_), .Y(u2__abc_52155_new_n3639_));
INVX1 INVX1_4300 ( .A(u2__abc_52155_new_n23574_), .Y(u2__abc_52155_new_n23575_));
INVX1 INVX1_4301 ( .A(u2__abc_52155_new_n23581_), .Y(u2__abc_52155_new_n23582_));
INVX1 INVX1_4302 ( .A(u2__abc_52155_new_n23586_), .Y(u2__abc_52155_new_n23587_));
INVX1 INVX1_4303 ( .A(u2__abc_52155_new_n23594_), .Y(u2__abc_52155_new_n23595_));
INVX1 INVX1_4304 ( .A(u2__abc_52155_new_n23598_), .Y(u2__abc_52155_new_n23599_));
INVX1 INVX1_4305 ( .A(u2__abc_52155_new_n23605_), .Y(u2__abc_52155_new_n23606_));
INVX1 INVX1_4306 ( .A(u2__abc_52155_new_n23610_), .Y(u2__abc_52155_new_n23611_));
INVX1 INVX1_4307 ( .A(u2__abc_52155_new_n23618_), .Y(u2__abc_52155_new_n23619_));
INVX1 INVX1_4308 ( .A(u2__abc_52155_new_n23622_), .Y(u2__abc_52155_new_n23623_));
INVX1 INVX1_4309 ( .A(u2__abc_52155_new_n23629_), .Y(u2__abc_52155_new_n23630_));
INVX1 INVX1_431 ( .A(sqrto_118_), .Y(u2__abc_52155_new_n3643_));
INVX1 INVX1_4310 ( .A(u2__abc_52155_new_n23634_), .Y(u2__abc_52155_new_n23635_));
INVX1 INVX1_4311 ( .A(u2__abc_52155_new_n23642_), .Y(u2__abc_52155_new_n23643_));
INVX1 INVX1_4312 ( .A(u2__abc_52155_new_n23646_), .Y(u2__abc_52155_new_n23647_));
INVX1 INVX1_4313 ( .A(u2__abc_52155_new_n23653_), .Y(u2__abc_52155_new_n23654_));
INVX1 INVX1_4314 ( .A(u2__abc_52155_new_n23658_), .Y(u2__abc_52155_new_n23659_));
INVX1 INVX1_4315 ( .A(u2__abc_52155_new_n23666_), .Y(u2__abc_52155_new_n23667_));
INVX1 INVX1_4316 ( .A(u2__abc_52155_new_n23670_), .Y(u2__abc_52155_new_n23671_));
INVX1 INVX1_4317 ( .A(u2__abc_52155_new_n23677_), .Y(u2__abc_52155_new_n23678_));
INVX1 INVX1_4318 ( .A(u2__abc_52155_new_n23682_), .Y(u2__abc_52155_new_n23683_));
INVX1 INVX1_4319 ( .A(u2__abc_52155_new_n23690_), .Y(u2__abc_52155_new_n23691_));
INVX1 INVX1_432 ( .A(u2__abc_52155_new_n3644_), .Y(u2__abc_52155_new_n3645_));
INVX1 INVX1_4320 ( .A(u2__abc_52155_new_n23694_), .Y(u2__abc_52155_new_n23695_));
INVX1 INVX1_4321 ( .A(u2__abc_52155_new_n23701_), .Y(u2__abc_52155_new_n23702_));
INVX1 INVX1_4322 ( .A(u2__abc_52155_new_n23706_), .Y(u2__abc_52155_new_n23707_));
INVX1 INVX1_4323 ( .A(u2__abc_52155_new_n23714_), .Y(u2__abc_52155_new_n23715_));
INVX1 INVX1_4324 ( .A(u2__abc_52155_new_n23718_), .Y(u2__abc_52155_new_n23719_));
INVX1 INVX1_4325 ( .A(u2__abc_52155_new_n23726_), .Y(u2__abc_52155_new_n23727_));
INVX1 INVX1_4326 ( .A(u2__abc_52155_new_n23730_), .Y(u2__abc_52155_new_n23731_));
INVX1 INVX1_4327 ( .A(u2__abc_52155_new_n23738_), .Y(u2__abc_52155_new_n23739_));
INVX1 INVX1_4328 ( .A(u2__abc_52155_new_n23742_), .Y(u2__abc_52155_new_n23743_));
INVX1 INVX1_4329 ( .A(u2__abc_52155_new_n23749_), .Y(u2__abc_52155_new_n23750_));
INVX1 INVX1_433 ( .A(u2_remHi_118_), .Y(u2__abc_52155_new_n3646_));
INVX1 INVX1_4330 ( .A(u2__abc_52155_new_n23754_), .Y(u2__abc_52155_new_n23755_));
INVX1 INVX1_4331 ( .A(u2__abc_52155_new_n23762_), .Y(u2__abc_52155_new_n23763_));
INVX1 INVX1_4332 ( .A(u2__abc_52155_new_n23766_), .Y(u2__abc_52155_new_n23767_));
INVX1 INVX1_4333 ( .A(u2__abc_52155_new_n23774_), .Y(u2__abc_52155_new_n23775_));
INVX1 INVX1_4334 ( .A(u2__abc_52155_new_n23778_), .Y(u2__abc_52155_new_n23779_));
INVX1 INVX1_4335 ( .A(u2__abc_52155_new_n23786_), .Y(u2__abc_52155_new_n23787_));
INVX1 INVX1_4336 ( .A(u2__abc_52155_new_n23790_), .Y(u2__abc_52155_new_n23791_));
INVX1 INVX1_4337 ( .A(u2__abc_52155_new_n23797_), .Y(u2__abc_52155_new_n23798_));
INVX1 INVX1_4338 ( .A(u2__abc_52155_new_n23802_), .Y(u2__abc_52155_new_n23803_));
INVX1 INVX1_4339 ( .A(u2__abc_52155_new_n23810_), .Y(u2__abc_52155_new_n23811_));
INVX1 INVX1_434 ( .A(u2__abc_52155_new_n3647_), .Y(u2__abc_52155_new_n3648_));
INVX1 INVX1_4340 ( .A(u2__abc_52155_new_n23814_), .Y(u2__abc_52155_new_n23815_));
INVX1 INVX1_4341 ( .A(u2__abc_52155_new_n23822_), .Y(u2__abc_52155_new_n23823_));
INVX1 INVX1_4342 ( .A(u2__abc_52155_new_n23826_), .Y(u2__abc_52155_new_n23827_));
INVX1 INVX1_4343 ( .A(u2__abc_52155_new_n23834_), .Y(u2__abc_52155_new_n23835_));
INVX1 INVX1_4344 ( .A(u2__abc_52155_new_n23838_), .Y(u2__abc_52155_new_n23839_));
INVX1 INVX1_4345 ( .A(u2__abc_52155_new_n23845_), .Y(u2__abc_52155_new_n23846_));
INVX1 INVX1_4346 ( .A(u2__abc_52155_new_n23850_), .Y(u2__abc_52155_new_n23851_));
INVX1 INVX1_4347 ( .A(u2__abc_52155_new_n23858_), .Y(u2__abc_52155_new_n23859_));
INVX1 INVX1_4348 ( .A(u2__abc_52155_new_n23862_), .Y(u2__abc_52155_new_n23863_));
INVX1 INVX1_4349 ( .A(u2__abc_52155_new_n23869_), .Y(u2__abc_52155_new_n23870_));
INVX1 INVX1_435 ( .A(sqrto_119_), .Y(u2__abc_52155_new_n3650_));
INVX1 INVX1_4350 ( .A(u2__abc_52155_new_n23874_), .Y(u2__abc_52155_new_n23875_));
INVX1 INVX1_4351 ( .A(u2__abc_52155_new_n23882_), .Y(u2__abc_52155_new_n23883_));
INVX1 INVX1_4352 ( .A(u2__abc_52155_new_n23886_), .Y(u2__abc_52155_new_n23887_));
INVX1 INVX1_4353 ( .A(u2__abc_52155_new_n23893_), .Y(u2__abc_52155_new_n23894_));
INVX1 INVX1_4354 ( .A(u2__abc_52155_new_n23898_), .Y(u2__abc_52155_new_n23899_));
INVX1 INVX1_4355 ( .A(u2__abc_52155_new_n23906_), .Y(u2__abc_52155_new_n23907_));
INVX1 INVX1_4356 ( .A(u2__abc_52155_new_n23910_), .Y(u2__abc_52155_new_n23911_));
INVX1 INVX1_4357 ( .A(u2__abc_52155_new_n23918_), .Y(u2__abc_52155_new_n23919_));
INVX1 INVX1_4358 ( .A(u2__abc_52155_new_n23922_), .Y(u2__abc_52155_new_n23923_));
INVX1 INVX1_4359 ( .A(u2__abc_52155_new_n23930_), .Y(u2__abc_52155_new_n23931_));
INVX1 INVX1_436 ( .A(u2__abc_52155_new_n3651_), .Y(u2__abc_52155_new_n3652_));
INVX1 INVX1_4360 ( .A(u2__abc_52155_new_n23934_), .Y(u2__abc_52155_new_n23935_));
INVX1 INVX1_4361 ( .A(u2__abc_52155_new_n23941_), .Y(u2__abc_52155_new_n23942_));
INVX1 INVX1_4362 ( .A(u2__abc_52155_new_n23946_), .Y(u2__abc_52155_new_n23947_));
INVX1 INVX1_4363 ( .A(u2__abc_52155_new_n23954_), .Y(u2__abc_52155_new_n23955_));
INVX1 INVX1_4364 ( .A(u2__abc_52155_new_n23958_), .Y(u2__abc_52155_new_n23959_));
INVX1 INVX1_4365 ( .A(u2__abc_52155_new_n23965_), .Y(u2__abc_52155_new_n23966_));
INVX1 INVX1_4366 ( .A(u2__abc_52155_new_n23970_), .Y(u2__abc_52155_new_n23971_));
INVX1 INVX1_4367 ( .A(u2__abc_52155_new_n23978_), .Y(u2__abc_52155_new_n23979_));
INVX1 INVX1_4368 ( .A(u2__abc_52155_new_n23982_), .Y(u2__abc_52155_new_n23983_));
INVX1 INVX1_4369 ( .A(u2__abc_52155_new_n23989_), .Y(u2__abc_52155_new_n23990_));
INVX1 INVX1_437 ( .A(u2_remHi_119_), .Y(u2__abc_52155_new_n3653_));
INVX1 INVX1_4370 ( .A(u2__abc_52155_new_n23994_), .Y(u2__abc_52155_new_n23995_));
INVX1 INVX1_4371 ( .A(u2__abc_52155_new_n24002_), .Y(u2__abc_52155_new_n24003_));
INVX1 INVX1_4372 ( .A(u2__abc_52155_new_n24006_), .Y(u2__abc_52155_new_n24007_));
INVX1 INVX1_4373 ( .A(u2__abc_52155_new_n24013_), .Y(u2__abc_52155_new_n24014_));
INVX1 INVX1_4374 ( .A(u2__abc_52155_new_n24018_), .Y(u2__abc_52155_new_n24019_));
INVX1 INVX1_4375 ( .A(u2__abc_52155_new_n24026_), .Y(u2__abc_52155_new_n24027_));
INVX1 INVX1_4376 ( .A(u2__abc_52155_new_n24030_), .Y(u2__abc_52155_new_n24031_));
INVX1 INVX1_4377 ( .A(u2__abc_52155_new_n24037_), .Y(u2__abc_52155_new_n24038_));
INVX1 INVX1_4378 ( .A(u2__abc_52155_new_n24042_), .Y(u2__abc_52155_new_n24043_));
INVX1 INVX1_4379 ( .A(u2__abc_52155_new_n24050_), .Y(u2__abc_52155_new_n24051_));
INVX1 INVX1_438 ( .A(u2__abc_52155_new_n3654_), .Y(u2__abc_52155_new_n3655_));
INVX1 INVX1_4380 ( .A(u2__abc_52155_new_n24054_), .Y(u2__abc_52155_new_n24055_));
INVX1 INVX1_4381 ( .A(u2__abc_52155_new_n24061_), .Y(u2__abc_52155_new_n24062_));
INVX1 INVX1_4382 ( .A(u2__abc_52155_new_n24066_), .Y(u2__abc_52155_new_n24067_));
INVX1 INVX1_4383 ( .A(u2__abc_52155_new_n24074_), .Y(u2__abc_52155_new_n24075_));
INVX1 INVX1_4384 ( .A(u2__abc_52155_new_n24078_), .Y(u2__abc_52155_new_n24079_));
INVX1 INVX1_4385 ( .A(u2__abc_52155_new_n24085_), .Y(u2__abc_52155_new_n24086_));
INVX1 INVX1_4386 ( .A(u2__abc_52155_new_n24090_), .Y(u2__abc_52155_new_n24091_));
INVX1 INVX1_4387 ( .A(u2__abc_52155_new_n24098_), .Y(u2__abc_52155_new_n24099_));
INVX1 INVX1_4388 ( .A(u2__abc_52155_new_n24102_), .Y(u2__abc_52155_new_n24103_));
INVX1 INVX1_4389 ( .A(u2__abc_52155_new_n24110_), .Y(u2__abc_52155_new_n24111_));
INVX1 INVX1_439 ( .A(sqrto_120_), .Y(u2__abc_52155_new_n3658_));
INVX1 INVX1_4390 ( .A(u2__abc_52155_new_n24114_), .Y(u2__abc_52155_new_n24115_));
INVX1 INVX1_4391 ( .A(u2__abc_52155_new_n24122_), .Y(u2__abc_52155_new_n24123_));
INVX1 INVX1_4392 ( .A(u2__abc_52155_new_n24126_), .Y(u2__abc_52155_new_n24127_));
INVX1 INVX1_4393 ( .A(u2__abc_52155_new_n24133_), .Y(u2__abc_52155_new_n24134_));
INVX1 INVX1_4394 ( .A(u2__abc_52155_new_n24138_), .Y(u2__abc_52155_new_n24139_));
INVX1 INVX1_4395 ( .A(u2__abc_52155_new_n24146_), .Y(u2__abc_52155_new_n24147_));
INVX1 INVX1_4396 ( .A(u2__abc_52155_new_n24150_), .Y(u2__abc_52155_new_n24151_));
INVX1 INVX1_4397 ( .A(u2__abc_52155_new_n24157_), .Y(u2__abc_52155_new_n24158_));
INVX1 INVX1_4398 ( .A(u2__abc_52155_new_n24162_), .Y(u2__abc_52155_new_n24163_));
INVX1 INVX1_4399 ( .A(u2__abc_52155_new_n24170_), .Y(u2__abc_52155_new_n24171_));
INVX1 INVX1_44 ( .A(_abc_73687_new_n1648_), .Y(_abc_73687_new_n1655_));
INVX1 INVX1_440 ( .A(u2__abc_52155_new_n3659_), .Y(u2__abc_52155_new_n3660_));
INVX1 INVX1_4400 ( .A(u2__abc_52155_new_n24174_), .Y(u2__abc_52155_new_n24175_));
INVX1 INVX1_4401 ( .A(u2__abc_52155_new_n24181_), .Y(u2__abc_52155_new_n24182_));
INVX1 INVX1_4402 ( .A(u2__abc_52155_new_n24186_), .Y(u2__abc_52155_new_n24187_));
INVX1 INVX1_4403 ( .A(u2__abc_52155_new_n24194_), .Y(u2__abc_52155_new_n24195_));
INVX1 INVX1_4404 ( .A(u2__abc_52155_new_n24198_), .Y(u2__abc_52155_new_n24199_));
INVX1 INVX1_4405 ( .A(u2__abc_52155_new_n24205_), .Y(u2__abc_52155_new_n24206_));
INVX1 INVX1_4406 ( .A(u2__abc_52155_new_n24210_), .Y(u2__abc_52155_new_n24211_));
INVX1 INVX1_4407 ( .A(u2__abc_52155_new_n24218_), .Y(u2__abc_52155_new_n24219_));
INVX1 INVX1_4408 ( .A(u2__abc_52155_new_n24222_), .Y(u2__abc_52155_new_n24223_));
INVX1 INVX1_4409 ( .A(u2__abc_52155_new_n24229_), .Y(u2__abc_52155_new_n24230_));
INVX1 INVX1_441 ( .A(u2_remHi_120_), .Y(u2__abc_52155_new_n3661_));
INVX1 INVX1_4410 ( .A(u2__abc_52155_new_n24234_), .Y(u2__abc_52155_new_n24235_));
INVX1 INVX1_4411 ( .A(u2__abc_52155_new_n24242_), .Y(u2__abc_52155_new_n24243_));
INVX1 INVX1_4412 ( .A(u2__abc_52155_new_n24246_), .Y(u2__abc_52155_new_n24247_));
INVX1 INVX1_4413 ( .A(u2__abc_52155_new_n24253_), .Y(u2__abc_52155_new_n24254_));
INVX1 INVX1_4414 ( .A(u2__abc_52155_new_n24258_), .Y(u2__abc_52155_new_n24259_));
INVX1 INVX1_4415 ( .A(u2__abc_52155_new_n24266_), .Y(u2__abc_52155_new_n24267_));
INVX1 INVX1_4416 ( .A(u2__abc_52155_new_n24270_), .Y(u2__abc_52155_new_n24271_));
INVX1 INVX1_4417 ( .A(u2__abc_52155_new_n24277_), .Y(u2__abc_52155_new_n24278_));
INVX1 INVX1_4418 ( .A(u2__abc_52155_new_n24282_), .Y(u2__abc_52155_new_n24283_));
INVX1 INVX1_4419 ( .A(u2__abc_52155_new_n24290_), .Y(u2__abc_52155_new_n24291_));
INVX1 INVX1_442 ( .A(u2__abc_52155_new_n3662_), .Y(u2__abc_52155_new_n3663_));
INVX1 INVX1_4420 ( .A(u2__abc_52155_new_n24294_), .Y(u2__abc_52155_new_n24295_));
INVX1 INVX1_4421 ( .A(u2__abc_52155_new_n24301_), .Y(u2__abc_52155_new_n24302_));
INVX1 INVX1_4422 ( .A(u2__abc_52155_new_n24306_), .Y(u2__abc_52155_new_n24307_));
INVX1 INVX1_4423 ( .A(u2__abc_52155_new_n24314_), .Y(u2__abc_52155_new_n24315_));
INVX1 INVX1_4424 ( .A(u2__abc_52155_new_n24318_), .Y(u2__abc_52155_new_n24319_));
INVX1 INVX1_4425 ( .A(u2__abc_52155_new_n24325_), .Y(u2__abc_52155_new_n24326_));
INVX1 INVX1_4426 ( .A(u2__abc_52155_new_n24330_), .Y(u2__abc_52155_new_n24331_));
INVX1 INVX1_4427 ( .A(u2__abc_52155_new_n24338_), .Y(u2__abc_52155_new_n24339_));
INVX1 INVX1_4428 ( .A(u2__abc_52155_new_n24342_), .Y(u2__abc_52155_new_n24343_));
INVX1 INVX1_4429 ( .A(u2__abc_52155_new_n24349_), .Y(u2__abc_52155_new_n24350_));
INVX1 INVX1_443 ( .A(sqrto_121_), .Y(u2__abc_52155_new_n3665_));
INVX1 INVX1_4430 ( .A(u2__abc_52155_new_n24354_), .Y(u2__abc_52155_new_n24355_));
INVX1 INVX1_4431 ( .A(u2__abc_52155_new_n24362_), .Y(u2__abc_52155_new_n24363_));
INVX1 INVX1_4432 ( .A(u2__abc_52155_new_n24366_), .Y(u2__abc_52155_new_n24367_));
INVX1 INVX1_4433 ( .A(u2__abc_52155_new_n24373_), .Y(u2__abc_52155_new_n24374_));
INVX1 INVX1_4434 ( .A(u2__abc_52155_new_n24378_), .Y(u2__abc_52155_new_n24379_));
INVX1 INVX1_4435 ( .A(u2__abc_52155_new_n24386_), .Y(u2__abc_52155_new_n24387_));
INVX1 INVX1_4436 ( .A(u2__abc_52155_new_n24390_), .Y(u2__abc_52155_new_n24391_));
INVX1 INVX1_4437 ( .A(u2__abc_52155_new_n24397_), .Y(u2__abc_52155_new_n24398_));
INVX1 INVX1_4438 ( .A(u2__abc_52155_new_n24402_), .Y(u2__abc_52155_new_n24403_));
INVX1 INVX1_4439 ( .A(u2__abc_52155_new_n24410_), .Y(u2__abc_52155_new_n24411_));
INVX1 INVX1_444 ( .A(u2__abc_52155_new_n3666_), .Y(u2__abc_52155_new_n3667_));
INVX1 INVX1_4440 ( .A(u2__abc_52155_new_n24414_), .Y(u2__abc_52155_new_n24415_));
INVX1 INVX1_4441 ( .A(u2__abc_52155_new_n24421_), .Y(u2__abc_52155_new_n24422_));
INVX1 INVX1_4442 ( .A(u2__abc_52155_new_n24426_), .Y(u2__abc_52155_new_n24427_));
INVX1 INVX1_4443 ( .A(u2__abc_52155_new_n24434_), .Y(u2__abc_52155_new_n24435_));
INVX1 INVX1_4444 ( .A(u2__abc_52155_new_n24438_), .Y(u2__abc_52155_new_n24439_));
INVX1 INVX1_4445 ( .A(u2__abc_52155_new_n24446_), .Y(u2__abc_52155_new_n24447_));
INVX1 INVX1_4446 ( .A(u2__abc_52155_new_n24450_), .Y(u2__abc_52155_new_n24451_));
INVX1 INVX1_4447 ( .A(u2__abc_52155_new_n24458_), .Y(u2__abc_52155_new_n24459_));
INVX1 INVX1_4448 ( .A(u2__abc_52155_new_n24462_), .Y(u2__abc_52155_new_n24463_));
INVX1 INVX1_445 ( .A(u2_remHi_121_), .Y(u2__abc_52155_new_n3668_));
INVX1 INVX1_446 ( .A(u2__abc_52155_new_n3669_), .Y(u2__abc_52155_new_n3670_));
INVX1 INVX1_447 ( .A(sqrto_124_), .Y(u2__abc_52155_new_n3674_));
INVX1 INVX1_448 ( .A(u2__abc_52155_new_n3675_), .Y(u2__abc_52155_new_n3676_));
INVX1 INVX1_449 ( .A(u2_remHi_124_), .Y(u2__abc_52155_new_n3677_));
INVX1 INVX1_45 ( .A(\a[125] ), .Y(_abc_73687_new_n1656_));
INVX1 INVX1_450 ( .A(u2__abc_52155_new_n3678_), .Y(u2__abc_52155_new_n3679_));
INVX1 INVX1_451 ( .A(u2_remHi_125_), .Y(u2__abc_52155_new_n3681_));
INVX1 INVX1_452 ( .A(u2__abc_52155_new_n3682_), .Y(u2__abc_52155_new_n3683_));
INVX1 INVX1_453 ( .A(sqrto_125_), .Y(u2__abc_52155_new_n3684_));
INVX1 INVX1_454 ( .A(u2__abc_52155_new_n3685_), .Y(u2__abc_52155_new_n3686_));
INVX1 INVX1_455 ( .A(sqrto_123_), .Y(u2__abc_52155_new_n3689_));
INVX1 INVX1_456 ( .A(u2__abc_52155_new_n3690_), .Y(u2__abc_52155_new_n3691_));
INVX1 INVX1_457 ( .A(u2_remHi_123_), .Y(u2__abc_52155_new_n3692_));
INVX1 INVX1_458 ( .A(u2__abc_52155_new_n3693_), .Y(u2__abc_52155_new_n3694_));
INVX1 INVX1_459 ( .A(sqrto_122_), .Y(u2__abc_52155_new_n3696_));
INVX1 INVX1_46 ( .A(_abc_73687_new_n1657_), .Y(_abc_73687_new_n1658_));
INVX1 INVX1_460 ( .A(u2__abc_52155_new_n3697_), .Y(u2__abc_52155_new_n3698_));
INVX1 INVX1_461 ( .A(u2_remHi_122_), .Y(u2__abc_52155_new_n3699_));
INVX1 INVX1_462 ( .A(u2__abc_52155_new_n3700_), .Y(u2__abc_52155_new_n3701_));
INVX1 INVX1_463 ( .A(sqrto_110_), .Y(u2__abc_52155_new_n3706_));
INVX1 INVX1_464 ( .A(u2__abc_52155_new_n3707_), .Y(u2__abc_52155_new_n3708_));
INVX1 INVX1_465 ( .A(u2_remHi_110_), .Y(u2__abc_52155_new_n3709_));
INVX1 INVX1_466 ( .A(u2__abc_52155_new_n3710_), .Y(u2__abc_52155_new_n3711_));
INVX1 INVX1_467 ( .A(sqrto_111_), .Y(u2__abc_52155_new_n3713_));
INVX1 INVX1_468 ( .A(u2__abc_52155_new_n3714_), .Y(u2__abc_52155_new_n3715_));
INVX1 INVX1_469 ( .A(u2_remHi_111_), .Y(u2__abc_52155_new_n3716_));
INVX1 INVX1_47 ( .A(_abc_73687_new_n1661_), .Y(_abc_73687_new_n1662_));
INVX1 INVX1_470 ( .A(u2__abc_52155_new_n3717_), .Y(u2__abc_52155_new_n3718_));
INVX1 INVX1_471 ( .A(sqrto_112_), .Y(u2__abc_52155_new_n3721_));
INVX1 INVX1_472 ( .A(u2__abc_52155_new_n3722_), .Y(u2__abc_52155_new_n3723_));
INVX1 INVX1_473 ( .A(u2_remHi_112_), .Y(u2__abc_52155_new_n3724_));
INVX1 INVX1_474 ( .A(u2__abc_52155_new_n3725_), .Y(u2__abc_52155_new_n3726_));
INVX1 INVX1_475 ( .A(sqrto_113_), .Y(u2__abc_52155_new_n3728_));
INVX1 INVX1_476 ( .A(u2__abc_52155_new_n3729_), .Y(u2__abc_52155_new_n3730_));
INVX1 INVX1_477 ( .A(u2_remHi_113_), .Y(u2__abc_52155_new_n3731_));
INVX1 INVX1_478 ( .A(u2__abc_52155_new_n3732_), .Y(u2__abc_52155_new_n3733_));
INVX1 INVX1_479 ( .A(sqrto_116_), .Y(u2__abc_52155_new_n3737_));
INVX1 INVX1_48 ( .A(\a[126] ), .Y(_abc_73687_new_n1670_));
INVX1 INVX1_480 ( .A(u2__abc_52155_new_n3738_), .Y(u2__abc_52155_new_n3739_));
INVX1 INVX1_481 ( .A(u2_remHi_116_), .Y(u2__abc_52155_new_n3740_));
INVX1 INVX1_482 ( .A(u2__abc_52155_new_n3741_), .Y(u2__abc_52155_new_n3742_));
INVX1 INVX1_483 ( .A(sqrto_117_), .Y(u2__abc_52155_new_n3744_));
INVX1 INVX1_484 ( .A(u2__abc_52155_new_n3745_), .Y(u2__abc_52155_new_n3746_));
INVX1 INVX1_485 ( .A(u2_remHi_117_), .Y(u2__abc_52155_new_n3747_));
INVX1 INVX1_486 ( .A(u2__abc_52155_new_n3748_), .Y(u2__abc_52155_new_n3749_));
INVX1 INVX1_487 ( .A(sqrto_115_), .Y(u2__abc_52155_new_n3752_));
INVX1 INVX1_488 ( .A(u2__abc_52155_new_n3753_), .Y(u2__abc_52155_new_n3754_));
INVX1 INVX1_489 ( .A(u2_remHi_115_), .Y(u2__abc_52155_new_n3755_));
INVX1 INVX1_49 ( .A(_abc_73687_new_n1672_), .Y(_abc_73687_new_n1673_));
INVX1 INVX1_490 ( .A(u2__abc_52155_new_n3756_), .Y(u2__abc_52155_new_n3757_));
INVX1 INVX1_491 ( .A(sqrto_114_), .Y(u2__abc_52155_new_n3759_));
INVX1 INVX1_492 ( .A(u2__abc_52155_new_n3760_), .Y(u2__abc_52155_new_n3761_));
INVX1 INVX1_493 ( .A(u2_remHi_114_), .Y(u2__abc_52155_new_n3762_));
INVX1 INVX1_494 ( .A(u2__abc_52155_new_n3763_), .Y(u2__abc_52155_new_n3764_));
INVX1 INVX1_495 ( .A(sqrto_104_), .Y(u2__abc_52155_new_n3770_));
INVX1 INVX1_496 ( .A(u2__abc_52155_new_n3771_), .Y(u2__abc_52155_new_n3772_));
INVX1 INVX1_497 ( .A(u2_remHi_104_), .Y(u2__abc_52155_new_n3773_));
INVX1 INVX1_498 ( .A(u2__abc_52155_new_n3774_), .Y(u2__abc_52155_new_n3775_));
INVX1 INVX1_499 ( .A(sqrto_105_), .Y(u2__abc_52155_new_n3777_));
INVX1 INVX1_5 ( .A(\a[115] ), .Y(_abc_73687_new_n1521_));
INVX1 INVX1_50 ( .A(_abc_73687_new_n1676_), .Y(_abc_73687_new_n1677_));
INVX1 INVX1_500 ( .A(u2__abc_52155_new_n3778_), .Y(u2__abc_52155_new_n3779_));
INVX1 INVX1_501 ( .A(u2_remHi_105_), .Y(u2__abc_52155_new_n3780_));
INVX1 INVX1_502 ( .A(u2__abc_52155_new_n3781_), .Y(u2__abc_52155_new_n3782_));
INVX1 INVX1_503 ( .A(sqrto_103_), .Y(u2__abc_52155_new_n3785_));
INVX1 INVX1_504 ( .A(u2__abc_52155_new_n3786_), .Y(u2__abc_52155_new_n3787_));
INVX1 INVX1_505 ( .A(u2_remHi_103_), .Y(u2__abc_52155_new_n3788_));
INVX1 INVX1_506 ( .A(u2__abc_52155_new_n3789_), .Y(u2__abc_52155_new_n3790_));
INVX1 INVX1_507 ( .A(sqrto_102_), .Y(u2__abc_52155_new_n3792_));
INVX1 INVX1_508 ( .A(u2__abc_52155_new_n3793_), .Y(u2__abc_52155_new_n3794_));
INVX1 INVX1_509 ( .A(u2_remHi_102_), .Y(u2__abc_52155_new_n3795_));
INVX1 INVX1_51 ( .A(_abc_73687_new_n1675_), .Y(_abc_73687_new_n1686_));
INVX1 INVX1_510 ( .A(u2__abc_52155_new_n3796_), .Y(u2__abc_52155_new_n3797_));
INVX1 INVX1_511 ( .A(sqrto_108_), .Y(u2__abc_52155_new_n3801_));
INVX1 INVX1_512 ( .A(u2__abc_52155_new_n3802_), .Y(u2__abc_52155_new_n3803_));
INVX1 INVX1_513 ( .A(u2_remHi_108_), .Y(u2__abc_52155_new_n3804_));
INVX1 INVX1_514 ( .A(u2__abc_52155_new_n3805_), .Y(u2__abc_52155_new_n3806_));
INVX1 INVX1_515 ( .A(sqrto_109_), .Y(u2__abc_52155_new_n3808_));
INVX1 INVX1_516 ( .A(u2__abc_52155_new_n3809_), .Y(u2__abc_52155_new_n3810_));
INVX1 INVX1_517 ( .A(u2_remHi_109_), .Y(u2__abc_52155_new_n3811_));
INVX1 INVX1_518 ( .A(u2__abc_52155_new_n3812_), .Y(u2__abc_52155_new_n3813_));
INVX1 INVX1_519 ( .A(sqrto_107_), .Y(u2__abc_52155_new_n3816_));
INVX1 INVX1_52 ( .A(\a[10] ), .Y(u1__abc_51895_new_n166_));
INVX1 INVX1_520 ( .A(u2__abc_52155_new_n3817_), .Y(u2__abc_52155_new_n3818_));
INVX1 INVX1_521 ( .A(u2_remHi_107_), .Y(u2__abc_52155_new_n3819_));
INVX1 INVX1_522 ( .A(u2__abc_52155_new_n3820_), .Y(u2__abc_52155_new_n3821_));
INVX1 INVX1_523 ( .A(sqrto_106_), .Y(u2__abc_52155_new_n3823_));
INVX1 INVX1_524 ( .A(u2__abc_52155_new_n3824_), .Y(u2__abc_52155_new_n3825_));
INVX1 INVX1_525 ( .A(u2_remHi_106_), .Y(u2__abc_52155_new_n3826_));
INVX1 INVX1_526 ( .A(u2__abc_52155_new_n3827_), .Y(u2__abc_52155_new_n3828_));
INVX1 INVX1_527 ( .A(sqrto_96_), .Y(u2__abc_52155_new_n3833_));
INVX1 INVX1_528 ( .A(u2_remHi_96_), .Y(u2__abc_52155_new_n3835_));
INVX1 INVX1_529 ( .A(sqrto_97_), .Y(u2__abc_52155_new_n3838_));
INVX1 INVX1_53 ( .A(\a[11] ), .Y(u1__abc_51895_new_n167_));
INVX1 INVX1_530 ( .A(u2_remHi_97_), .Y(u2__abc_52155_new_n3840_));
INVX1 INVX1_531 ( .A(u2__abc_52155_new_n3843_), .Y(u2__abc_52155_new_n3844_));
INVX1 INVX1_532 ( .A(sqrto_95_), .Y(u2__abc_52155_new_n3845_));
INVX1 INVX1_533 ( .A(u2__abc_52155_new_n3846_), .Y(u2__abc_52155_new_n3847_));
INVX1 INVX1_534 ( .A(u2_remHi_95_), .Y(u2__abc_52155_new_n3848_));
INVX1 INVX1_535 ( .A(u2__abc_52155_new_n3849_), .Y(u2__abc_52155_new_n3850_));
INVX1 INVX1_536 ( .A(sqrto_94_), .Y(u2__abc_52155_new_n3852_));
INVX1 INVX1_537 ( .A(u2__abc_52155_new_n3853_), .Y(u2__abc_52155_new_n3854_));
INVX1 INVX1_538 ( .A(u2_remHi_94_), .Y(u2__abc_52155_new_n3855_));
INVX1 INVX1_539 ( .A(u2__abc_52155_new_n3856_), .Y(u2__abc_52155_new_n3857_));
INVX1 INVX1_54 ( .A(\a[8] ), .Y(u1__abc_51895_new_n169_));
INVX1 INVX1_540 ( .A(sqrto_100_), .Y(u2__abc_52155_new_n3861_));
INVX1 INVX1_541 ( .A(u2__abc_52155_new_n3862_), .Y(u2__abc_52155_new_n3863_));
INVX1 INVX1_542 ( .A(u2_remHi_100_), .Y(u2__abc_52155_new_n3864_));
INVX1 INVX1_543 ( .A(u2__abc_52155_new_n3865_), .Y(u2__abc_52155_new_n3866_));
INVX1 INVX1_544 ( .A(sqrto_101_), .Y(u2__abc_52155_new_n3868_));
INVX1 INVX1_545 ( .A(u2__abc_52155_new_n3869_), .Y(u2__abc_52155_new_n3870_));
INVX1 INVX1_546 ( .A(u2_remHi_101_), .Y(u2__abc_52155_new_n3871_));
INVX1 INVX1_547 ( .A(u2__abc_52155_new_n3872_), .Y(u2__abc_52155_new_n3873_));
INVX1 INVX1_548 ( .A(sqrto_99_), .Y(u2__abc_52155_new_n3876_));
INVX1 INVX1_549 ( .A(u2__abc_52155_new_n3877_), .Y(u2__abc_52155_new_n3878_));
INVX1 INVX1_55 ( .A(\a[9] ), .Y(u1__abc_51895_new_n170_));
INVX1 INVX1_550 ( .A(u2_remHi_99_), .Y(u2__abc_52155_new_n3879_));
INVX1 INVX1_551 ( .A(u2__abc_52155_new_n3880_), .Y(u2__abc_52155_new_n3881_));
INVX1 INVX1_552 ( .A(sqrto_98_), .Y(u2__abc_52155_new_n3883_));
INVX1 INVX1_553 ( .A(u2__abc_52155_new_n3884_), .Y(u2__abc_52155_new_n3885_));
INVX1 INVX1_554 ( .A(u2_remHi_98_), .Y(u2__abc_52155_new_n3886_));
INVX1 INVX1_555 ( .A(u2__abc_52155_new_n3887_), .Y(u2__abc_52155_new_n3888_));
INVX1 INVX1_556 ( .A(sqrto_92_), .Y(u2__abc_52155_new_n3895_));
INVX1 INVX1_557 ( .A(u2__abc_52155_new_n3896_), .Y(u2__abc_52155_new_n3897_));
INVX1 INVX1_558 ( .A(u2_remHi_92_), .Y(u2__abc_52155_new_n3898_));
INVX1 INVX1_559 ( .A(u2__abc_52155_new_n3899_), .Y(u2__abc_52155_new_n3900_));
INVX1 INVX1_56 ( .A(\a[14] ), .Y(u1__abc_51895_new_n173_));
INVX1 INVX1_560 ( .A(sqrto_93_), .Y(u2__abc_52155_new_n3902_));
INVX1 INVX1_561 ( .A(u2__abc_52155_new_n3903_), .Y(u2__abc_52155_new_n3904_));
INVX1 INVX1_562 ( .A(u2_remHi_93_), .Y(u2__abc_52155_new_n3905_));
INVX1 INVX1_563 ( .A(u2__abc_52155_new_n3906_), .Y(u2__abc_52155_new_n3907_));
INVX1 INVX1_564 ( .A(sqrto_91_), .Y(u2__abc_52155_new_n3910_));
INVX1 INVX1_565 ( .A(u2__abc_52155_new_n3911_), .Y(u2__abc_52155_new_n3912_));
INVX1 INVX1_566 ( .A(u2_remHi_91_), .Y(u2__abc_52155_new_n3913_));
INVX1 INVX1_567 ( .A(u2__abc_52155_new_n3914_), .Y(u2__abc_52155_new_n3915_));
INVX1 INVX1_568 ( .A(sqrto_90_), .Y(u2__abc_52155_new_n3917_));
INVX1 INVX1_569 ( .A(u2__abc_52155_new_n3918_), .Y(u2__abc_52155_new_n3919_));
INVX1 INVX1_57 ( .A(\a[15] ), .Y(u1__abc_51895_new_n174_));
INVX1 INVX1_570 ( .A(u2_remHi_90_), .Y(u2__abc_52155_new_n3920_));
INVX1 INVX1_571 ( .A(u2__abc_52155_new_n3921_), .Y(u2__abc_52155_new_n3922_));
INVX1 INVX1_572 ( .A(sqrto_88_), .Y(u2__abc_52155_new_n3926_));
INVX1 INVX1_573 ( .A(u2__abc_52155_new_n3927_), .Y(u2__abc_52155_new_n3928_));
INVX1 INVX1_574 ( .A(u2_remHi_88_), .Y(u2__abc_52155_new_n3929_));
INVX1 INVX1_575 ( .A(u2__abc_52155_new_n3930_), .Y(u2__abc_52155_new_n3931_));
INVX1 INVX1_576 ( .A(sqrto_89_), .Y(u2__abc_52155_new_n3933_));
INVX1 INVX1_577 ( .A(u2__abc_52155_new_n3934_), .Y(u2__abc_52155_new_n3935_));
INVX1 INVX1_578 ( .A(u2_remHi_89_), .Y(u2__abc_52155_new_n3936_));
INVX1 INVX1_579 ( .A(u2__abc_52155_new_n3937_), .Y(u2__abc_52155_new_n3938_));
INVX1 INVX1_58 ( .A(\a[12] ), .Y(u1__abc_51895_new_n176_));
INVX1 INVX1_580 ( .A(sqrto_87_), .Y(u2__abc_52155_new_n3941_));
INVX1 INVX1_581 ( .A(u2__abc_52155_new_n3942_), .Y(u2__abc_52155_new_n3943_));
INVX1 INVX1_582 ( .A(u2_remHi_87_), .Y(u2__abc_52155_new_n3944_));
INVX1 INVX1_583 ( .A(u2__abc_52155_new_n3945_), .Y(u2__abc_52155_new_n3946_));
INVX1 INVX1_584 ( .A(sqrto_86_), .Y(u2__abc_52155_new_n3948_));
INVX1 INVX1_585 ( .A(u2__abc_52155_new_n3949_), .Y(u2__abc_52155_new_n3950_));
INVX1 INVX1_586 ( .A(u2_remHi_86_), .Y(u2__abc_52155_new_n3951_));
INVX1 INVX1_587 ( .A(u2__abc_52155_new_n3952_), .Y(u2__abc_52155_new_n3953_));
INVX1 INVX1_588 ( .A(sqrto_78_), .Y(u2__abc_52155_new_n3958_));
INVX1 INVX1_589 ( .A(u2__abc_52155_new_n3959_), .Y(u2__abc_52155_new_n3960_));
INVX1 INVX1_59 ( .A(\a[13] ), .Y(u1__abc_51895_new_n177_));
INVX1 INVX1_590 ( .A(u2_remHi_78_), .Y(u2__abc_52155_new_n3961_));
INVX1 INVX1_591 ( .A(u2__abc_52155_new_n3962_), .Y(u2__abc_52155_new_n3963_));
INVX1 INVX1_592 ( .A(sqrto_79_), .Y(u2__abc_52155_new_n3965_));
INVX1 INVX1_593 ( .A(u2__abc_52155_new_n3966_), .Y(u2__abc_52155_new_n3967_));
INVX1 INVX1_594 ( .A(u2_remHi_79_), .Y(u2__abc_52155_new_n3968_));
INVX1 INVX1_595 ( .A(u2__abc_52155_new_n3969_), .Y(u2__abc_52155_new_n3970_));
INVX1 INVX1_596 ( .A(sqrto_80_), .Y(u2__abc_52155_new_n3973_));
INVX1 INVX1_597 ( .A(u2_remHi_80_), .Y(u2__abc_52155_new_n3975_));
INVX1 INVX1_598 ( .A(sqrto_81_), .Y(u2__abc_52155_new_n3978_));
INVX1 INVX1_599 ( .A(u2_remHi_81_), .Y(u2__abc_52155_new_n3980_));
INVX1 INVX1_6 ( .A(_abc_73687_new_n1522_), .Y(_abc_73687_new_n1523_));
INVX1 INVX1_60 ( .A(\a[2] ), .Y(u1__abc_51895_new_n181_));
INVX1 INVX1_600 ( .A(u2__abc_52155_new_n3983_), .Y(u2__abc_52155_new_n3984_));
INVX1 INVX1_601 ( .A(sqrto_84_), .Y(u2__abc_52155_new_n3986_));
INVX1 INVX1_602 ( .A(u2__abc_52155_new_n3987_), .Y(u2__abc_52155_new_n3988_));
INVX1 INVX1_603 ( .A(u2_remHi_84_), .Y(u2__abc_52155_new_n3989_));
INVX1 INVX1_604 ( .A(u2__abc_52155_new_n3990_), .Y(u2__abc_52155_new_n3991_));
INVX1 INVX1_605 ( .A(sqrto_85_), .Y(u2__abc_52155_new_n3993_));
INVX1 INVX1_606 ( .A(u2__abc_52155_new_n3994_), .Y(u2__abc_52155_new_n3995_));
INVX1 INVX1_607 ( .A(u2_remHi_85_), .Y(u2__abc_52155_new_n3996_));
INVX1 INVX1_608 ( .A(u2__abc_52155_new_n3997_), .Y(u2__abc_52155_new_n3998_));
INVX1 INVX1_609 ( .A(sqrto_83_), .Y(u2__abc_52155_new_n4001_));
INVX1 INVX1_61 ( .A(\a[3] ), .Y(u1__abc_51895_new_n182_));
INVX1 INVX1_610 ( .A(u2__abc_52155_new_n4002_), .Y(u2__abc_52155_new_n4003_));
INVX1 INVX1_611 ( .A(u2_remHi_83_), .Y(u2__abc_52155_new_n4004_));
INVX1 INVX1_612 ( .A(u2__abc_52155_new_n4005_), .Y(u2__abc_52155_new_n4006_));
INVX1 INVX1_613 ( .A(sqrto_82_), .Y(u2__abc_52155_new_n4008_));
INVX1 INVX1_614 ( .A(u2__abc_52155_new_n4009_), .Y(u2__abc_52155_new_n4010_));
INVX1 INVX1_615 ( .A(u2_remHi_82_), .Y(u2__abc_52155_new_n4011_));
INVX1 INVX1_616 ( .A(u2__abc_52155_new_n4012_), .Y(u2__abc_52155_new_n4013_));
INVX1 INVX1_617 ( .A(sqrto_70_), .Y(u2__abc_52155_new_n4019_));
INVX1 INVX1_618 ( .A(u2__abc_52155_new_n4020_), .Y(u2__abc_52155_new_n4021_));
INVX1 INVX1_619 ( .A(u2_remHi_70_), .Y(u2__abc_52155_new_n4022_));
INVX1 INVX1_62 ( .A(\a[0] ), .Y(u1__abc_51895_new_n184_));
INVX1 INVX1_620 ( .A(u2__abc_52155_new_n4023_), .Y(u2__abc_52155_new_n4024_));
INVX1 INVX1_621 ( .A(sqrto_71_), .Y(u2__abc_52155_new_n4026_));
INVX1 INVX1_622 ( .A(u2__abc_52155_new_n4027_), .Y(u2__abc_52155_new_n4028_));
INVX1 INVX1_623 ( .A(u2_remHi_71_), .Y(u2__abc_52155_new_n4029_));
INVX1 INVX1_624 ( .A(u2__abc_52155_new_n4030_), .Y(u2__abc_52155_new_n4031_));
INVX1 INVX1_625 ( .A(sqrto_72_), .Y(u2__abc_52155_new_n4034_));
INVX1 INVX1_626 ( .A(u2_remHi_72_), .Y(u2__abc_52155_new_n4036_));
INVX1 INVX1_627 ( .A(sqrto_73_), .Y(u2__abc_52155_new_n4039_));
INVX1 INVX1_628 ( .A(u2_remHi_73_), .Y(u2__abc_52155_new_n4041_));
INVX1 INVX1_629 ( .A(u2__abc_52155_new_n4044_), .Y(u2__abc_52155_new_n4045_));
INVX1 INVX1_63 ( .A(\a[1] ), .Y(u1__abc_51895_new_n185_));
INVX1 INVX1_630 ( .A(sqrto_76_), .Y(u2__abc_52155_new_n4047_));
INVX1 INVX1_631 ( .A(u2__abc_52155_new_n4048_), .Y(u2__abc_52155_new_n4049_));
INVX1 INVX1_632 ( .A(u2_remHi_76_), .Y(u2__abc_52155_new_n4050_));
INVX1 INVX1_633 ( .A(u2__abc_52155_new_n4051_), .Y(u2__abc_52155_new_n4052_));
INVX1 INVX1_634 ( .A(sqrto_77_), .Y(u2__abc_52155_new_n4054_));
INVX1 INVX1_635 ( .A(u2__abc_52155_new_n4055_), .Y(u2__abc_52155_new_n4056_));
INVX1 INVX1_636 ( .A(u2_remHi_77_), .Y(u2__abc_52155_new_n4057_));
INVX1 INVX1_637 ( .A(u2__abc_52155_new_n4058_), .Y(u2__abc_52155_new_n4059_));
INVX1 INVX1_638 ( .A(sqrto_75_), .Y(u2__abc_52155_new_n4062_));
INVX1 INVX1_639 ( .A(u2__abc_52155_new_n4063_), .Y(u2__abc_52155_new_n4064_));
INVX1 INVX1_64 ( .A(\a[6] ), .Y(u1__abc_51895_new_n188_));
INVX1 INVX1_640 ( .A(u2_remHi_75_), .Y(u2__abc_52155_new_n4065_));
INVX1 INVX1_641 ( .A(u2__abc_52155_new_n4066_), .Y(u2__abc_52155_new_n4067_));
INVX1 INVX1_642 ( .A(sqrto_74_), .Y(u2__abc_52155_new_n4069_));
INVX1 INVX1_643 ( .A(u2__abc_52155_new_n4070_), .Y(u2__abc_52155_new_n4071_));
INVX1 INVX1_644 ( .A(u2_remHi_74_), .Y(u2__abc_52155_new_n4072_));
INVX1 INVX1_645 ( .A(u2__abc_52155_new_n4073_), .Y(u2__abc_52155_new_n4074_));
INVX1 INVX1_646 ( .A(sqrto_62_), .Y(u2__abc_52155_new_n4079_));
INVX1 INVX1_647 ( .A(u2__abc_52155_new_n4080_), .Y(u2__abc_52155_new_n4081_));
INVX1 INVX1_648 ( .A(sqrto_63_), .Y(u2__abc_52155_new_n4084_));
INVX1 INVX1_649 ( .A(u2__abc_52155_new_n4085_), .Y(u2__abc_52155_new_n4086_));
INVX1 INVX1_65 ( .A(\a[7] ), .Y(u1__abc_51895_new_n189_));
INVX1 INVX1_650 ( .A(u2_remHi_63_), .Y(u2__abc_52155_new_n4087_));
INVX1 INVX1_651 ( .A(u2__abc_52155_new_n4088_), .Y(u2__abc_52155_new_n4089_));
INVX1 INVX1_652 ( .A(sqrto_64_), .Y(u2__abc_52155_new_n4092_));
INVX1 INVX1_653 ( .A(u2_remHi_64_), .Y(u2__abc_52155_new_n4094_));
INVX1 INVX1_654 ( .A(sqrto_65_), .Y(u2__abc_52155_new_n4097_));
INVX1 INVX1_655 ( .A(u2_remHi_65_), .Y(u2__abc_52155_new_n4099_));
INVX1 INVX1_656 ( .A(u2__abc_52155_new_n4102_), .Y(u2__abc_52155_new_n4103_));
INVX1 INVX1_657 ( .A(sqrto_68_), .Y(u2__abc_52155_new_n4105_));
INVX1 INVX1_658 ( .A(u2_remHi_68_), .Y(u2__abc_52155_new_n4107_));
INVX1 INVX1_659 ( .A(sqrto_69_), .Y(u2__abc_52155_new_n4110_));
INVX1 INVX1_66 ( .A(\a[4] ), .Y(u1__abc_51895_new_n191_));
INVX1 INVX1_660 ( .A(u2_remHi_69_), .Y(u2__abc_52155_new_n4112_));
INVX1 INVX1_661 ( .A(sqrto_67_), .Y(u2__abc_52155_new_n4116_));
INVX1 INVX1_662 ( .A(u2_remHi_67_), .Y(u2__abc_52155_new_n4118_));
INVX1 INVX1_663 ( .A(sqrto_66_), .Y(u2__abc_52155_new_n4121_));
INVX1 INVX1_664 ( .A(u2_remHi_66_), .Y(u2__abc_52155_new_n4123_));
INVX1 INVX1_665 ( .A(u2__abc_52155_new_n4127_), .Y(u2__abc_52155_new_n4128_));
INVX1 INVX1_666 ( .A(u2__abc_52155_new_n4132_), .Y(u2__abc_52155_new_n4133_));
INVX1 INVX1_667 ( .A(u2__abc_52155_new_n3894_), .Y(u2__abc_52155_new_n4135_));
INVX1 INVX1_668 ( .A(u2__abc_52155_new_n4018_), .Y(u2__abc_52155_new_n4136_));
INVX1 INVX1_669 ( .A(u2__abc_52155_new_n4078_), .Y(u2__abc_52155_new_n4137_));
INVX1 INVX1_67 ( .A(\a[5] ), .Y(u1__abc_51895_new_n192_));
INVX1 INVX1_670 ( .A(u2__abc_52155_new_n4100_), .Y(u2__abc_52155_new_n4141_));
INVX1 INVX1_671 ( .A(u2__abc_52155_new_n4095_), .Y(u2__abc_52155_new_n4142_));
INVX1 INVX1_672 ( .A(u2__abc_52155_new_n4119_), .Y(u2__abc_52155_new_n4147_));
INVX1 INVX1_673 ( .A(u2__abc_52155_new_n4124_), .Y(u2__abc_52155_new_n4148_));
INVX1 INVX1_674 ( .A(u2__abc_52155_new_n4111_), .Y(u2__abc_52155_new_n4152_));
INVX1 INVX1_675 ( .A(u2__abc_52155_new_n4154_), .Y(u2__abc_52155_new_n4155_));
INVX1 INVX1_676 ( .A(u2__abc_52155_new_n4077_), .Y(u2__abc_52155_new_n4159_));
INVX1 INVX1_677 ( .A(u2__abc_52155_new_n4040_), .Y(u2__abc_52155_new_n4163_));
INVX1 INVX1_678 ( .A(u2__abc_52155_new_n4165_), .Y(u2__abc_52155_new_n4166_));
INVX1 INVX1_679 ( .A(u2__abc_52155_new_n4174_), .Y(u2__abc_52155_new_n4175_));
INVX1 INVX1_68 ( .A(\a[26] ), .Y(u1__abc_51895_new_n197_));
INVX1 INVX1_680 ( .A(u2__abc_52155_new_n3957_), .Y(u2__abc_52155_new_n4179_));
INVX1 INVX1_681 ( .A(u2__abc_52155_new_n4016_), .Y(u2__abc_52155_new_n4180_));
INVX1 INVX1_682 ( .A(u2__abc_52155_new_n3979_), .Y(u2__abc_52155_new_n4184_));
INVX1 INVX1_683 ( .A(u2__abc_52155_new_n4186_), .Y(u2__abc_52155_new_n4187_));
INVX1 INVX1_684 ( .A(u2__abc_52155_new_n4195_), .Y(u2__abc_52155_new_n4196_));
INVX1 INVX1_685 ( .A(u2__abc_52155_new_n4212_), .Y(u2__abc_52155_new_n4213_));
INVX1 INVX1_686 ( .A(u2__abc_52155_new_n3769_), .Y(u2__abc_52155_new_n4217_));
INVX1 INVX1_687 ( .A(u2__abc_52155_new_n3832_), .Y(u2__abc_52155_new_n4218_));
INVX1 INVX1_688 ( .A(u2__abc_52155_new_n3891_), .Y(u2__abc_52155_new_n4219_));
INVX1 INVX1_689 ( .A(u2__abc_52155_new_n3839_), .Y(u2__abc_52155_new_n4223_));
INVX1 INVX1_69 ( .A(\a[27] ), .Y(u1__abc_51895_new_n198_));
INVX1 INVX1_690 ( .A(u2__abc_52155_new_n4225_), .Y(u2__abc_52155_new_n4226_));
INVX1 INVX1_691 ( .A(u2__abc_52155_new_n4234_), .Y(u2__abc_52155_new_n4235_));
INVX1 INVX1_692 ( .A(u2__abc_52155_new_n4251_), .Y(u2__abc_52155_new_n4252_));
INVX1 INVX1_693 ( .A(u2__abc_52155_new_n4284_), .Y(u2__abc_52155_new_n4285_));
INVX1 INVX1_694 ( .A(u2_o_246_), .Y(u2__abc_52155_new_n4289_));
INVX1 INVX1_695 ( .A(u2__abc_52155_new_n4290_), .Y(u2__abc_52155_new_n4291_));
INVX1 INVX1_696 ( .A(u2_remHi_246_), .Y(u2__abc_52155_new_n4292_));
INVX1 INVX1_697 ( .A(u2__abc_52155_new_n4293_), .Y(u2__abc_52155_new_n4294_));
INVX1 INVX1_698 ( .A(u2_o_247_), .Y(u2__abc_52155_new_n4296_));
INVX1 INVX1_699 ( .A(u2__abc_52155_new_n4297_), .Y(u2__abc_52155_new_n4298_));
INVX1 INVX1_7 ( .A(_abc_73687_new_n1509_), .Y(_abc_73687_new_n1524_));
INVX1 INVX1_70 ( .A(\a[24] ), .Y(u1__abc_51895_new_n200_));
INVX1 INVX1_700 ( .A(u2_remHi_247_), .Y(u2__abc_52155_new_n4299_));
INVX1 INVX1_701 ( .A(u2__abc_52155_new_n4300_), .Y(u2__abc_52155_new_n4301_));
INVX1 INVX1_702 ( .A(u2_o_248_), .Y(u2__abc_52155_new_n4304_));
INVX1 INVX1_703 ( .A(u2__abc_52155_new_n4305_), .Y(u2__abc_52155_new_n4306_));
INVX1 INVX1_704 ( .A(u2_remHi_248_), .Y(u2__abc_52155_new_n4307_));
INVX1 INVX1_705 ( .A(u2__abc_52155_new_n4308_), .Y(u2__abc_52155_new_n4309_));
INVX1 INVX1_706 ( .A(u2_o_249_), .Y(u2__abc_52155_new_n4311_));
INVX1 INVX1_707 ( .A(u2__abc_52155_new_n4312_), .Y(u2__abc_52155_new_n4313_));
INVX1 INVX1_708 ( .A(u2_remHi_249_), .Y(u2__abc_52155_new_n4314_));
INVX1 INVX1_709 ( .A(u2__abc_52155_new_n4315_), .Y(u2__abc_52155_new_n4316_));
INVX1 INVX1_71 ( .A(\a[25] ), .Y(u1__abc_51895_new_n201_));
INVX1 INVX1_710 ( .A(u2_o_252_), .Y(u2__abc_52155_new_n4320_));
INVX1 INVX1_711 ( .A(u2__abc_52155_new_n4321_), .Y(u2__abc_52155_new_n4322_));
INVX1 INVX1_712 ( .A(u2_remHi_252_), .Y(u2__abc_52155_new_n4323_));
INVX1 INVX1_713 ( .A(u2__abc_52155_new_n4324_), .Y(u2__abc_52155_new_n4325_));
INVX1 INVX1_714 ( .A(u2_remHi_253_), .Y(u2__abc_52155_new_n4327_));
INVX1 INVX1_715 ( .A(u2__abc_52155_new_n4328_), .Y(u2__abc_52155_new_n4329_));
INVX1 INVX1_716 ( .A(u2_o_253_), .Y(u2__abc_52155_new_n4330_));
INVX1 INVX1_717 ( .A(u2__abc_52155_new_n4331_), .Y(u2__abc_52155_new_n4332_));
INVX1 INVX1_718 ( .A(u2_o_251_), .Y(u2__abc_52155_new_n4335_));
INVX1 INVX1_719 ( .A(u2__abc_52155_new_n4336_), .Y(u2__abc_52155_new_n4337_));
INVX1 INVX1_72 ( .A(\a[30] ), .Y(u1__abc_51895_new_n204_));
INVX1 INVX1_720 ( .A(u2_remHi_251_), .Y(u2__abc_52155_new_n4338_));
INVX1 INVX1_721 ( .A(u2__abc_52155_new_n4339_), .Y(u2__abc_52155_new_n4340_));
INVX1 INVX1_722 ( .A(u2_o_250_), .Y(u2__abc_52155_new_n4342_));
INVX1 INVX1_723 ( .A(u2__abc_52155_new_n4343_), .Y(u2__abc_52155_new_n4344_));
INVX1 INVX1_724 ( .A(u2_remHi_250_), .Y(u2__abc_52155_new_n4345_));
INVX1 INVX1_725 ( .A(u2__abc_52155_new_n4346_), .Y(u2__abc_52155_new_n4347_));
INVX1 INVX1_726 ( .A(u2_o_238_), .Y(u2__abc_52155_new_n4352_));
INVX1 INVX1_727 ( .A(u2__abc_52155_new_n4353_), .Y(u2__abc_52155_new_n4354_));
INVX1 INVX1_728 ( .A(u2_remHi_238_), .Y(u2__abc_52155_new_n4355_));
INVX1 INVX1_729 ( .A(u2__abc_52155_new_n4356_), .Y(u2__abc_52155_new_n4357_));
INVX1 INVX1_73 ( .A(\a[31] ), .Y(u1__abc_51895_new_n205_));
INVX1 INVX1_730 ( .A(u2_o_239_), .Y(u2__abc_52155_new_n4359_));
INVX1 INVX1_731 ( .A(u2__abc_52155_new_n4360_), .Y(u2__abc_52155_new_n4361_));
INVX1 INVX1_732 ( .A(u2_remHi_239_), .Y(u2__abc_52155_new_n4362_));
INVX1 INVX1_733 ( .A(u2__abc_52155_new_n4363_), .Y(u2__abc_52155_new_n4364_));
INVX1 INVX1_734 ( .A(u2_o_240_), .Y(u2__abc_52155_new_n4367_));
INVX1 INVX1_735 ( .A(u2__abc_52155_new_n4368_), .Y(u2__abc_52155_new_n4369_));
INVX1 INVX1_736 ( .A(u2_remHi_240_), .Y(u2__abc_52155_new_n4370_));
INVX1 INVX1_737 ( .A(u2__abc_52155_new_n4371_), .Y(u2__abc_52155_new_n4372_));
INVX1 INVX1_738 ( .A(u2_o_241_), .Y(u2__abc_52155_new_n4374_));
INVX1 INVX1_739 ( .A(u2__abc_52155_new_n4375_), .Y(u2__abc_52155_new_n4376_));
INVX1 INVX1_74 ( .A(\a[28] ), .Y(u1__abc_51895_new_n207_));
INVX1 INVX1_740 ( .A(u2_remHi_241_), .Y(u2__abc_52155_new_n4377_));
INVX1 INVX1_741 ( .A(u2__abc_52155_new_n4378_), .Y(u2__abc_52155_new_n4379_));
INVX1 INVX1_742 ( .A(u2_o_244_), .Y(u2__abc_52155_new_n4383_));
INVX1 INVX1_743 ( .A(u2__abc_52155_new_n4384_), .Y(u2__abc_52155_new_n4385_));
INVX1 INVX1_744 ( .A(u2_remHi_244_), .Y(u2__abc_52155_new_n4386_));
INVX1 INVX1_745 ( .A(u2__abc_52155_new_n4387_), .Y(u2__abc_52155_new_n4388_));
INVX1 INVX1_746 ( .A(u2_o_245_), .Y(u2__abc_52155_new_n4390_));
INVX1 INVX1_747 ( .A(u2__abc_52155_new_n4391_), .Y(u2__abc_52155_new_n4392_));
INVX1 INVX1_748 ( .A(u2_remHi_245_), .Y(u2__abc_52155_new_n4393_));
INVX1 INVX1_749 ( .A(u2__abc_52155_new_n4394_), .Y(u2__abc_52155_new_n4395_));
INVX1 INVX1_75 ( .A(\a[29] ), .Y(u1__abc_51895_new_n208_));
INVX1 INVX1_750 ( .A(u2_o_243_), .Y(u2__abc_52155_new_n4398_));
INVX1 INVX1_751 ( .A(u2__abc_52155_new_n4399_), .Y(u2__abc_52155_new_n4400_));
INVX1 INVX1_752 ( .A(u2_remHi_243_), .Y(u2__abc_52155_new_n4401_));
INVX1 INVX1_753 ( .A(u2__abc_52155_new_n4402_), .Y(u2__abc_52155_new_n4403_));
INVX1 INVX1_754 ( .A(u2_o_242_), .Y(u2__abc_52155_new_n4405_));
INVX1 INVX1_755 ( .A(u2__abc_52155_new_n4406_), .Y(u2__abc_52155_new_n4407_));
INVX1 INVX1_756 ( .A(u2_remHi_242_), .Y(u2__abc_52155_new_n4408_));
INVX1 INVX1_757 ( .A(u2__abc_52155_new_n4409_), .Y(u2__abc_52155_new_n4410_));
INVX1 INVX1_758 ( .A(u2_o_236_), .Y(u2__abc_52155_new_n4416_));
INVX1 INVX1_759 ( .A(u2__abc_52155_new_n4417_), .Y(u2__abc_52155_new_n4418_));
INVX1 INVX1_76 ( .A(\a[18] ), .Y(u1__abc_51895_new_n212_));
INVX1 INVX1_760 ( .A(u2_remHi_236_), .Y(u2__abc_52155_new_n4419_));
INVX1 INVX1_761 ( .A(u2__abc_52155_new_n4420_), .Y(u2__abc_52155_new_n4421_));
INVX1 INVX1_762 ( .A(u2_o_237_), .Y(u2__abc_52155_new_n4423_));
INVX1 INVX1_763 ( .A(u2__abc_52155_new_n4424_), .Y(u2__abc_52155_new_n4425_));
INVX1 INVX1_764 ( .A(u2_remHi_237_), .Y(u2__abc_52155_new_n4426_));
INVX1 INVX1_765 ( .A(u2__abc_52155_new_n4427_), .Y(u2__abc_52155_new_n4428_));
INVX1 INVX1_766 ( .A(u2_o_235_), .Y(u2__abc_52155_new_n4431_));
INVX1 INVX1_767 ( .A(u2__abc_52155_new_n4432_), .Y(u2__abc_52155_new_n4433_));
INVX1 INVX1_768 ( .A(u2_remHi_235_), .Y(u2__abc_52155_new_n4434_));
INVX1 INVX1_769 ( .A(u2__abc_52155_new_n4435_), .Y(u2__abc_52155_new_n4436_));
INVX1 INVX1_77 ( .A(\a[19] ), .Y(u1__abc_51895_new_n213_));
INVX1 INVX1_770 ( .A(u2_o_234_), .Y(u2__abc_52155_new_n4438_));
INVX1 INVX1_771 ( .A(u2__abc_52155_new_n4439_), .Y(u2__abc_52155_new_n4440_));
INVX1 INVX1_772 ( .A(u2_remHi_234_), .Y(u2__abc_52155_new_n4441_));
INVX1 INVX1_773 ( .A(u2__abc_52155_new_n4442_), .Y(u2__abc_52155_new_n4443_));
INVX1 INVX1_774 ( .A(u2_o_232_), .Y(u2__abc_52155_new_n4447_));
INVX1 INVX1_775 ( .A(u2__abc_52155_new_n4448_), .Y(u2__abc_52155_new_n4449_));
INVX1 INVX1_776 ( .A(u2_remHi_232_), .Y(u2__abc_52155_new_n4450_));
INVX1 INVX1_777 ( .A(u2__abc_52155_new_n4451_), .Y(u2__abc_52155_new_n4452_));
INVX1 INVX1_778 ( .A(u2_o_233_), .Y(u2__abc_52155_new_n4454_));
INVX1 INVX1_779 ( .A(u2__abc_52155_new_n4455_), .Y(u2__abc_52155_new_n4456_));
INVX1 INVX1_78 ( .A(\a[16] ), .Y(u1__abc_51895_new_n215_));
INVX1 INVX1_780 ( .A(u2_remHi_233_), .Y(u2__abc_52155_new_n4457_));
INVX1 INVX1_781 ( .A(u2__abc_52155_new_n4458_), .Y(u2__abc_52155_new_n4459_));
INVX1 INVX1_782 ( .A(u2_o_231_), .Y(u2__abc_52155_new_n4462_));
INVX1 INVX1_783 ( .A(u2__abc_52155_new_n4463_), .Y(u2__abc_52155_new_n4464_));
INVX1 INVX1_784 ( .A(u2_remHi_231_), .Y(u2__abc_52155_new_n4465_));
INVX1 INVX1_785 ( .A(u2__abc_52155_new_n4466_), .Y(u2__abc_52155_new_n4467_));
INVX1 INVX1_786 ( .A(u2_o_230_), .Y(u2__abc_52155_new_n4469_));
INVX1 INVX1_787 ( .A(u2__abc_52155_new_n4470_), .Y(u2__abc_52155_new_n4471_));
INVX1 INVX1_788 ( .A(u2_remHi_230_), .Y(u2__abc_52155_new_n4472_));
INVX1 INVX1_789 ( .A(u2__abc_52155_new_n4473_), .Y(u2__abc_52155_new_n4474_));
INVX1 INVX1_79 ( .A(\a[17] ), .Y(u1__abc_51895_new_n216_));
INVX1 INVX1_790 ( .A(sqrto_224_), .Y(u2__abc_52155_new_n4479_));
INVX1 INVX1_791 ( .A(u2__abc_52155_new_n4480_), .Y(u2__abc_52155_new_n4481_));
INVX1 INVX1_792 ( .A(u2_remHi_224_), .Y(u2__abc_52155_new_n4482_));
INVX1 INVX1_793 ( .A(u2__abc_52155_new_n4483_), .Y(u2__abc_52155_new_n4484_));
INVX1 INVX1_794 ( .A(sqrto_225_), .Y(u2__abc_52155_new_n4486_));
INVX1 INVX1_795 ( .A(u2__abc_52155_new_n4487_), .Y(u2__abc_52155_new_n4488_));
INVX1 INVX1_796 ( .A(u2_remHi_225_), .Y(u2__abc_52155_new_n4489_));
INVX1 INVX1_797 ( .A(u2__abc_52155_new_n4490_), .Y(u2__abc_52155_new_n4491_));
INVX1 INVX1_798 ( .A(sqrto_223_), .Y(u2__abc_52155_new_n4494_));
INVX1 INVX1_799 ( .A(u2__abc_52155_new_n4495_), .Y(u2__abc_52155_new_n4496_));
INVX1 INVX1_8 ( .A(_abc_73687_new_n1526_), .Y(_abc_73687_new_n1527_));
INVX1 INVX1_80 ( .A(\a[22] ), .Y(u1__abc_51895_new_n219_));
INVX1 INVX1_800 ( .A(u2_remHi_223_), .Y(u2__abc_52155_new_n4497_));
INVX1 INVX1_801 ( .A(u2__abc_52155_new_n4498_), .Y(u2__abc_52155_new_n4499_));
INVX1 INVX1_802 ( .A(sqrto_222_), .Y(u2__abc_52155_new_n4501_));
INVX1 INVX1_803 ( .A(u2__abc_52155_new_n4502_), .Y(u2__abc_52155_new_n4503_));
INVX1 INVX1_804 ( .A(u2_remHi_222_), .Y(u2__abc_52155_new_n4504_));
INVX1 INVX1_805 ( .A(u2__abc_52155_new_n4505_), .Y(u2__abc_52155_new_n4506_));
INVX1 INVX1_806 ( .A(u2_o_228_), .Y(u2__abc_52155_new_n4510_));
INVX1 INVX1_807 ( .A(u2__abc_52155_new_n4511_), .Y(u2__abc_52155_new_n4512_));
INVX1 INVX1_808 ( .A(u2_remHi_228_), .Y(u2__abc_52155_new_n4513_));
INVX1 INVX1_809 ( .A(u2__abc_52155_new_n4514_), .Y(u2__abc_52155_new_n4515_));
INVX1 INVX1_81 ( .A(\a[23] ), .Y(u1__abc_51895_new_n220_));
INVX1 INVX1_810 ( .A(u2_o_229_), .Y(u2__abc_52155_new_n4517_));
INVX1 INVX1_811 ( .A(u2__abc_52155_new_n4518_), .Y(u2__abc_52155_new_n4519_));
INVX1 INVX1_812 ( .A(u2_remHi_229_), .Y(u2__abc_52155_new_n4520_));
INVX1 INVX1_813 ( .A(u2__abc_52155_new_n4521_), .Y(u2__abc_52155_new_n4522_));
INVX1 INVX1_814 ( .A(u2_o_227_), .Y(u2__abc_52155_new_n4525_));
INVX1 INVX1_815 ( .A(u2__abc_52155_new_n4526_), .Y(u2__abc_52155_new_n4527_));
INVX1 INVX1_816 ( .A(u2_remHi_227_), .Y(u2__abc_52155_new_n4528_));
INVX1 INVX1_817 ( .A(u2__abc_52155_new_n4529_), .Y(u2__abc_52155_new_n4530_));
INVX1 INVX1_818 ( .A(u2_o_226_), .Y(u2__abc_52155_new_n4532_));
INVX1 INVX1_819 ( .A(u2__abc_52155_new_n4533_), .Y(u2__abc_52155_new_n4534_));
INVX1 INVX1_82 ( .A(\a[20] ), .Y(u1__abc_51895_new_n222_));
INVX1 INVX1_820 ( .A(u2_remHi_226_), .Y(u2__abc_52155_new_n4535_));
INVX1 INVX1_821 ( .A(u2__abc_52155_new_n4536_), .Y(u2__abc_52155_new_n4537_));
INVX1 INVX1_822 ( .A(sqrto_216_), .Y(u2__abc_52155_new_n4544_));
INVX1 INVX1_823 ( .A(u2__abc_52155_new_n4545_), .Y(u2__abc_52155_new_n4546_));
INVX1 INVX1_824 ( .A(u2_remHi_216_), .Y(u2__abc_52155_new_n4547_));
INVX1 INVX1_825 ( .A(u2__abc_52155_new_n4548_), .Y(u2__abc_52155_new_n4549_));
INVX1 INVX1_826 ( .A(sqrto_217_), .Y(u2__abc_52155_new_n4551_));
INVX1 INVX1_827 ( .A(u2__abc_52155_new_n4552_), .Y(u2__abc_52155_new_n4553_));
INVX1 INVX1_828 ( .A(u2_remHi_217_), .Y(u2__abc_52155_new_n4554_));
INVX1 INVX1_829 ( .A(u2__abc_52155_new_n4555_), .Y(u2__abc_52155_new_n4556_));
INVX1 INVX1_83 ( .A(\a[21] ), .Y(u1__abc_51895_new_n223_));
INVX1 INVX1_830 ( .A(sqrto_214_), .Y(u2__abc_52155_new_n4559_));
INVX1 INVX1_831 ( .A(u2__abc_52155_new_n4560_), .Y(u2__abc_52155_new_n4561_));
INVX1 INVX1_832 ( .A(u2_remHi_214_), .Y(u2__abc_52155_new_n4562_));
INVX1 INVX1_833 ( .A(u2__abc_52155_new_n4563_), .Y(u2__abc_52155_new_n4564_));
INVX1 INVX1_834 ( .A(sqrto_215_), .Y(u2__abc_52155_new_n4566_));
INVX1 INVX1_835 ( .A(u2__abc_52155_new_n4567_), .Y(u2__abc_52155_new_n4568_));
INVX1 INVX1_836 ( .A(u2_remHi_215_), .Y(u2__abc_52155_new_n4569_));
INVX1 INVX1_837 ( .A(u2__abc_52155_new_n4570_), .Y(u2__abc_52155_new_n4571_));
INVX1 INVX1_838 ( .A(sqrto_220_), .Y(u2__abc_52155_new_n4575_));
INVX1 INVX1_839 ( .A(u2__abc_52155_new_n4576_), .Y(u2__abc_52155_new_n4577_));
INVX1 INVX1_84 ( .A(\a[42] ), .Y(u1__abc_51895_new_n228_));
INVX1 INVX1_840 ( .A(u2_remHi_220_), .Y(u2__abc_52155_new_n4578_));
INVX1 INVX1_841 ( .A(u2__abc_52155_new_n4579_), .Y(u2__abc_52155_new_n4580_));
INVX1 INVX1_842 ( .A(sqrto_221_), .Y(u2__abc_52155_new_n4582_));
INVX1 INVX1_843 ( .A(u2__abc_52155_new_n4583_), .Y(u2__abc_52155_new_n4584_));
INVX1 INVX1_844 ( .A(u2_remHi_221_), .Y(u2__abc_52155_new_n4585_));
INVX1 INVX1_845 ( .A(u2__abc_52155_new_n4586_), .Y(u2__abc_52155_new_n4587_));
INVX1 INVX1_846 ( .A(sqrto_219_), .Y(u2__abc_52155_new_n4590_));
INVX1 INVX1_847 ( .A(u2__abc_52155_new_n4591_), .Y(u2__abc_52155_new_n4592_));
INVX1 INVX1_848 ( .A(u2_remHi_219_), .Y(u2__abc_52155_new_n4593_));
INVX1 INVX1_849 ( .A(u2__abc_52155_new_n4594_), .Y(u2__abc_52155_new_n4595_));
INVX1 INVX1_85 ( .A(\a[43] ), .Y(u1__abc_51895_new_n229_));
INVX1 INVX1_850 ( .A(sqrto_218_), .Y(u2__abc_52155_new_n4597_));
INVX1 INVX1_851 ( .A(u2__abc_52155_new_n4598_), .Y(u2__abc_52155_new_n4599_));
INVX1 INVX1_852 ( .A(u2_remHi_218_), .Y(u2__abc_52155_new_n4600_));
INVX1 INVX1_853 ( .A(u2__abc_52155_new_n4601_), .Y(u2__abc_52155_new_n4602_));
INVX1 INVX1_854 ( .A(sqrto_208_), .Y(u2__abc_52155_new_n4607_));
INVX1 INVX1_855 ( .A(u2__abc_52155_new_n4608_), .Y(u2__abc_52155_new_n4609_));
INVX1 INVX1_856 ( .A(u2_remHi_208_), .Y(u2__abc_52155_new_n4610_));
INVX1 INVX1_857 ( .A(u2__abc_52155_new_n4611_), .Y(u2__abc_52155_new_n4612_));
INVX1 INVX1_858 ( .A(sqrto_209_), .Y(u2__abc_52155_new_n4614_));
INVX1 INVX1_859 ( .A(u2__abc_52155_new_n4615_), .Y(u2__abc_52155_new_n4616_));
INVX1 INVX1_86 ( .A(\a[40] ), .Y(u1__abc_51895_new_n231_));
INVX1 INVX1_860 ( .A(u2_remHi_209_), .Y(u2__abc_52155_new_n4617_));
INVX1 INVX1_861 ( .A(u2__abc_52155_new_n4618_), .Y(u2__abc_52155_new_n4619_));
INVX1 INVX1_862 ( .A(sqrto_206_), .Y(u2__abc_52155_new_n4622_));
INVX1 INVX1_863 ( .A(u2__abc_52155_new_n4623_), .Y(u2__abc_52155_new_n4624_));
INVX1 INVX1_864 ( .A(u2_remHi_206_), .Y(u2__abc_52155_new_n4625_));
INVX1 INVX1_865 ( .A(u2__abc_52155_new_n4626_), .Y(u2__abc_52155_new_n4627_));
INVX1 INVX1_866 ( .A(sqrto_207_), .Y(u2__abc_52155_new_n4629_));
INVX1 INVX1_867 ( .A(u2__abc_52155_new_n4630_), .Y(u2__abc_52155_new_n4631_));
INVX1 INVX1_868 ( .A(u2_remHi_207_), .Y(u2__abc_52155_new_n4632_));
INVX1 INVX1_869 ( .A(u2__abc_52155_new_n4633_), .Y(u2__abc_52155_new_n4634_));
INVX1 INVX1_87 ( .A(\a[41] ), .Y(u1__abc_51895_new_n232_));
INVX1 INVX1_870 ( .A(sqrto_212_), .Y(u2__abc_52155_new_n4638_));
INVX1 INVX1_871 ( .A(u2__abc_52155_new_n4639_), .Y(u2__abc_52155_new_n4640_));
INVX1 INVX1_872 ( .A(u2_remHi_212_), .Y(u2__abc_52155_new_n4641_));
INVX1 INVX1_873 ( .A(u2__abc_52155_new_n4642_), .Y(u2__abc_52155_new_n4643_));
INVX1 INVX1_874 ( .A(sqrto_213_), .Y(u2__abc_52155_new_n4645_));
INVX1 INVX1_875 ( .A(u2__abc_52155_new_n4646_), .Y(u2__abc_52155_new_n4647_));
INVX1 INVX1_876 ( .A(u2_remHi_213_), .Y(u2__abc_52155_new_n4648_));
INVX1 INVX1_877 ( .A(u2__abc_52155_new_n4649_), .Y(u2__abc_52155_new_n4650_));
INVX1 INVX1_878 ( .A(sqrto_211_), .Y(u2__abc_52155_new_n4653_));
INVX1 INVX1_879 ( .A(u2__abc_52155_new_n4654_), .Y(u2__abc_52155_new_n4655_));
INVX1 INVX1_88 ( .A(\a[46] ), .Y(u1__abc_51895_new_n235_));
INVX1 INVX1_880 ( .A(u2_remHi_211_), .Y(u2__abc_52155_new_n4656_));
INVX1 INVX1_881 ( .A(u2__abc_52155_new_n4657_), .Y(u2__abc_52155_new_n4658_));
INVX1 INVX1_882 ( .A(sqrto_210_), .Y(u2__abc_52155_new_n4660_));
INVX1 INVX1_883 ( .A(u2__abc_52155_new_n4661_), .Y(u2__abc_52155_new_n4662_));
INVX1 INVX1_884 ( .A(u2_remHi_210_), .Y(u2__abc_52155_new_n4663_));
INVX1 INVX1_885 ( .A(u2__abc_52155_new_n4664_), .Y(u2__abc_52155_new_n4665_));
INVX1 INVX1_886 ( .A(sqrto_200_), .Y(u2__abc_52155_new_n4671_));
INVX1 INVX1_887 ( .A(u2__abc_52155_new_n4672_), .Y(u2__abc_52155_new_n4673_));
INVX1 INVX1_888 ( .A(u2_remHi_200_), .Y(u2__abc_52155_new_n4674_));
INVX1 INVX1_889 ( .A(u2__abc_52155_new_n4675_), .Y(u2__abc_52155_new_n4676_));
INVX1 INVX1_89 ( .A(\a[47] ), .Y(u1__abc_51895_new_n236_));
INVX1 INVX1_890 ( .A(sqrto_201_), .Y(u2__abc_52155_new_n4678_));
INVX1 INVX1_891 ( .A(u2__abc_52155_new_n4679_), .Y(u2__abc_52155_new_n4680_));
INVX1 INVX1_892 ( .A(u2_remHi_201_), .Y(u2__abc_52155_new_n4681_));
INVX1 INVX1_893 ( .A(u2__abc_52155_new_n4682_), .Y(u2__abc_52155_new_n4683_));
INVX1 INVX1_894 ( .A(sqrto_199_), .Y(u2__abc_52155_new_n4686_));
INVX1 INVX1_895 ( .A(u2__abc_52155_new_n4687_), .Y(u2__abc_52155_new_n4688_));
INVX1 INVX1_896 ( .A(u2_remHi_199_), .Y(u2__abc_52155_new_n4689_));
INVX1 INVX1_897 ( .A(u2__abc_52155_new_n4690_), .Y(u2__abc_52155_new_n4691_));
INVX1 INVX1_898 ( .A(sqrto_198_), .Y(u2__abc_52155_new_n4693_));
INVX1 INVX1_899 ( .A(u2__abc_52155_new_n4694_), .Y(u2__abc_52155_new_n4695_));
INVX1 INVX1_9 ( .A(\a[116] ), .Y(_abc_73687_new_n1537_));
INVX1 INVX1_90 ( .A(\a[44] ), .Y(u1__abc_51895_new_n238_));
INVX1 INVX1_900 ( .A(u2_remHi_198_), .Y(u2__abc_52155_new_n4696_));
INVX1 INVX1_901 ( .A(u2__abc_52155_new_n4697_), .Y(u2__abc_52155_new_n4698_));
INVX1 INVX1_902 ( .A(sqrto_204_), .Y(u2__abc_52155_new_n4702_));
INVX1 INVX1_903 ( .A(u2__abc_52155_new_n4703_), .Y(u2__abc_52155_new_n4704_));
INVX1 INVX1_904 ( .A(u2_remHi_204_), .Y(u2__abc_52155_new_n4705_));
INVX1 INVX1_905 ( .A(u2__abc_52155_new_n4706_), .Y(u2__abc_52155_new_n4707_));
INVX1 INVX1_906 ( .A(sqrto_205_), .Y(u2__abc_52155_new_n4709_));
INVX1 INVX1_907 ( .A(u2__abc_52155_new_n4710_), .Y(u2__abc_52155_new_n4711_));
INVX1 INVX1_908 ( .A(u2_remHi_205_), .Y(u2__abc_52155_new_n4712_));
INVX1 INVX1_909 ( .A(u2__abc_52155_new_n4713_), .Y(u2__abc_52155_new_n4714_));
INVX1 INVX1_91 ( .A(\a[45] ), .Y(u1__abc_51895_new_n239_));
INVX1 INVX1_910 ( .A(sqrto_203_), .Y(u2__abc_52155_new_n4717_));
INVX1 INVX1_911 ( .A(u2__abc_52155_new_n4718_), .Y(u2__abc_52155_new_n4719_));
INVX1 INVX1_912 ( .A(u2_remHi_203_), .Y(u2__abc_52155_new_n4720_));
INVX1 INVX1_913 ( .A(u2__abc_52155_new_n4721_), .Y(u2__abc_52155_new_n4722_));
INVX1 INVX1_914 ( .A(sqrto_202_), .Y(u2__abc_52155_new_n4724_));
INVX1 INVX1_915 ( .A(u2__abc_52155_new_n4725_), .Y(u2__abc_52155_new_n4726_));
INVX1 INVX1_916 ( .A(u2_remHi_202_), .Y(u2__abc_52155_new_n4727_));
INVX1 INVX1_917 ( .A(u2__abc_52155_new_n4728_), .Y(u2__abc_52155_new_n4729_));
INVX1 INVX1_918 ( .A(sqrto_196_), .Y(u2__abc_52155_new_n4734_));
INVX1 INVX1_919 ( .A(u2__abc_52155_new_n4735_), .Y(u2__abc_52155_new_n4736_));
INVX1 INVX1_92 ( .A(\a[34] ), .Y(u1__abc_51895_new_n243_));
INVX1 INVX1_920 ( .A(u2_remHi_196_), .Y(u2__abc_52155_new_n4737_));
INVX1 INVX1_921 ( .A(u2__abc_52155_new_n4738_), .Y(u2__abc_52155_new_n4739_));
INVX1 INVX1_922 ( .A(sqrto_197_), .Y(u2__abc_52155_new_n4741_));
INVX1 INVX1_923 ( .A(u2__abc_52155_new_n4742_), .Y(u2__abc_52155_new_n4743_));
INVX1 INVX1_924 ( .A(u2_remHi_197_), .Y(u2__abc_52155_new_n4744_));
INVX1 INVX1_925 ( .A(u2__abc_52155_new_n4745_), .Y(u2__abc_52155_new_n4746_));
INVX1 INVX1_926 ( .A(sqrto_195_), .Y(u2__abc_52155_new_n4749_));
INVX1 INVX1_927 ( .A(u2__abc_52155_new_n4750_), .Y(u2__abc_52155_new_n4751_));
INVX1 INVX1_928 ( .A(u2_remHi_195_), .Y(u2__abc_52155_new_n4752_));
INVX1 INVX1_929 ( .A(u2__abc_52155_new_n4753_), .Y(u2__abc_52155_new_n4754_));
INVX1 INVX1_93 ( .A(\a[35] ), .Y(u1__abc_51895_new_n244_));
INVX1 INVX1_930 ( .A(sqrto_194_), .Y(u2__abc_52155_new_n4756_));
INVX1 INVX1_931 ( .A(u2__abc_52155_new_n4757_), .Y(u2__abc_52155_new_n4758_));
INVX1 INVX1_932 ( .A(u2_remHi_194_), .Y(u2__abc_52155_new_n4759_));
INVX1 INVX1_933 ( .A(u2__abc_52155_new_n4760_), .Y(u2__abc_52155_new_n4761_));
INVX1 INVX1_934 ( .A(sqrto_192_), .Y(u2__abc_52155_new_n4765_));
INVX1 INVX1_935 ( .A(u2_remHi_192_), .Y(u2__abc_52155_new_n4767_));
INVX1 INVX1_936 ( .A(sqrto_193_), .Y(u2__abc_52155_new_n4770_));
INVX1 INVX1_937 ( .A(u2_remHi_193_), .Y(u2__abc_52155_new_n4772_));
INVX1 INVX1_938 ( .A(u2__abc_52155_new_n4775_), .Y(u2__abc_52155_new_n4776_));
INVX1 INVX1_939 ( .A(sqrto_190_), .Y(u2__abc_52155_new_n4777_));
INVX1 INVX1_94 ( .A(\a[32] ), .Y(u1__abc_51895_new_n246_));
INVX1 INVX1_940 ( .A(u2__abc_52155_new_n4778_), .Y(u2__abc_52155_new_n4779_));
INVX1 INVX1_941 ( .A(u2_remHi_190_), .Y(u2__abc_52155_new_n4780_));
INVX1 INVX1_942 ( .A(u2__abc_52155_new_n4781_), .Y(u2__abc_52155_new_n4782_));
INVX1 INVX1_943 ( .A(sqrto_191_), .Y(u2__abc_52155_new_n4784_));
INVX1 INVX1_944 ( .A(u2__abc_52155_new_n4785_), .Y(u2__abc_52155_new_n4786_));
INVX1 INVX1_945 ( .A(u2_remHi_191_), .Y(u2__abc_52155_new_n4787_));
INVX1 INVX1_946 ( .A(u2__abc_52155_new_n4788_), .Y(u2__abc_52155_new_n4789_));
INVX1 INVX1_947 ( .A(sqrto_182_), .Y(u2__abc_52155_new_n4797_));
INVX1 INVX1_948 ( .A(u2__abc_52155_new_n4798_), .Y(u2__abc_52155_new_n4799_));
INVX1 INVX1_949 ( .A(u2_remHi_182_), .Y(u2__abc_52155_new_n4800_));
INVX1 INVX1_95 ( .A(\a[33] ), .Y(u1__abc_51895_new_n247_));
INVX1 INVX1_950 ( .A(u2__abc_52155_new_n4801_), .Y(u2__abc_52155_new_n4802_));
INVX1 INVX1_951 ( .A(sqrto_183_), .Y(u2__abc_52155_new_n4804_));
INVX1 INVX1_952 ( .A(u2__abc_52155_new_n4805_), .Y(u2__abc_52155_new_n4806_));
INVX1 INVX1_953 ( .A(u2_remHi_183_), .Y(u2__abc_52155_new_n4807_));
INVX1 INVX1_954 ( .A(u2__abc_52155_new_n4808_), .Y(u2__abc_52155_new_n4809_));
INVX1 INVX1_955 ( .A(sqrto_184_), .Y(u2__abc_52155_new_n4812_));
INVX1 INVX1_956 ( .A(u2__abc_52155_new_n4813_), .Y(u2__abc_52155_new_n4814_));
INVX1 INVX1_957 ( .A(u2_remHi_184_), .Y(u2__abc_52155_new_n4815_));
INVX1 INVX1_958 ( .A(u2__abc_52155_new_n4816_), .Y(u2__abc_52155_new_n4817_));
INVX1 INVX1_959 ( .A(sqrto_185_), .Y(u2__abc_52155_new_n4819_));
INVX1 INVX1_96 ( .A(\a[38] ), .Y(u1__abc_51895_new_n250_));
INVX1 INVX1_960 ( .A(u2__abc_52155_new_n4820_), .Y(u2__abc_52155_new_n4821_));
INVX1 INVX1_961 ( .A(u2_remHi_185_), .Y(u2__abc_52155_new_n4822_));
INVX1 INVX1_962 ( .A(u2__abc_52155_new_n4823_), .Y(u2__abc_52155_new_n4824_));
INVX1 INVX1_963 ( .A(sqrto_188_), .Y(u2__abc_52155_new_n4828_));
INVX1 INVX1_964 ( .A(u2__abc_52155_new_n4829_), .Y(u2__abc_52155_new_n4830_));
INVX1 INVX1_965 ( .A(u2_remHi_188_), .Y(u2__abc_52155_new_n4831_));
INVX1 INVX1_966 ( .A(u2__abc_52155_new_n4832_), .Y(u2__abc_52155_new_n4833_));
INVX1 INVX1_967 ( .A(sqrto_189_), .Y(u2__abc_52155_new_n4835_));
INVX1 INVX1_968 ( .A(u2__abc_52155_new_n4836_), .Y(u2__abc_52155_new_n4837_));
INVX1 INVX1_969 ( .A(u2_remHi_189_), .Y(u2__abc_52155_new_n4838_));
INVX1 INVX1_97 ( .A(\a[39] ), .Y(u1__abc_51895_new_n251_));
INVX1 INVX1_970 ( .A(u2__abc_52155_new_n4839_), .Y(u2__abc_52155_new_n4840_));
INVX1 INVX1_971 ( .A(sqrto_187_), .Y(u2__abc_52155_new_n4843_));
INVX1 INVX1_972 ( .A(u2__abc_52155_new_n4844_), .Y(u2__abc_52155_new_n4845_));
INVX1 INVX1_973 ( .A(u2_remHi_187_), .Y(u2__abc_52155_new_n4846_));
INVX1 INVX1_974 ( .A(u2__abc_52155_new_n4847_), .Y(u2__abc_52155_new_n4848_));
INVX1 INVX1_975 ( .A(sqrto_186_), .Y(u2__abc_52155_new_n4850_));
INVX1 INVX1_976 ( .A(u2__abc_52155_new_n4851_), .Y(u2__abc_52155_new_n4852_));
INVX1 INVX1_977 ( .A(u2_remHi_186_), .Y(u2__abc_52155_new_n4853_));
INVX1 INVX1_978 ( .A(u2__abc_52155_new_n4854_), .Y(u2__abc_52155_new_n4855_));
INVX1 INVX1_979 ( .A(sqrto_180_), .Y(u2__abc_52155_new_n4860_));
INVX1 INVX1_98 ( .A(\a[36] ), .Y(u1__abc_51895_new_n253_));
INVX1 INVX1_980 ( .A(u2__abc_52155_new_n4861_), .Y(u2__abc_52155_new_n4862_));
INVX1 INVX1_981 ( .A(u2_remHi_180_), .Y(u2__abc_52155_new_n4863_));
INVX1 INVX1_982 ( .A(u2__abc_52155_new_n4864_), .Y(u2__abc_52155_new_n4865_));
INVX1 INVX1_983 ( .A(sqrto_181_), .Y(u2__abc_52155_new_n4867_));
INVX1 INVX1_984 ( .A(u2__abc_52155_new_n4868_), .Y(u2__abc_52155_new_n4869_));
INVX1 INVX1_985 ( .A(u2_remHi_181_), .Y(u2__abc_52155_new_n4870_));
INVX1 INVX1_986 ( .A(u2__abc_52155_new_n4871_), .Y(u2__abc_52155_new_n4872_));
INVX1 INVX1_987 ( .A(sqrto_179_), .Y(u2__abc_52155_new_n4875_));
INVX1 INVX1_988 ( .A(u2__abc_52155_new_n4876_), .Y(u2__abc_52155_new_n4877_));
INVX1 INVX1_989 ( .A(u2_remHi_179_), .Y(u2__abc_52155_new_n4878_));
INVX1 INVX1_99 ( .A(\a[37] ), .Y(u1__abc_51895_new_n254_));
INVX1 INVX1_990 ( .A(u2__abc_52155_new_n4879_), .Y(u2__abc_52155_new_n4880_));
INVX1 INVX1_991 ( .A(sqrto_178_), .Y(u2__abc_52155_new_n4882_));
INVX1 INVX1_992 ( .A(u2__abc_52155_new_n4883_), .Y(u2__abc_52155_new_n4884_));
INVX1 INVX1_993 ( .A(u2_remHi_178_), .Y(u2__abc_52155_new_n4885_));
INVX1 INVX1_994 ( .A(u2__abc_52155_new_n4886_), .Y(u2__abc_52155_new_n4887_));
INVX1 INVX1_995 ( .A(sqrto_176_), .Y(u2__abc_52155_new_n4891_));
INVX1 INVX1_996 ( .A(u2__abc_52155_new_n4892_), .Y(u2__abc_52155_new_n4893_));
INVX1 INVX1_997 ( .A(u2_remHi_176_), .Y(u2__abc_52155_new_n4894_));
INVX1 INVX1_998 ( .A(u2__abc_52155_new_n4895_), .Y(u2__abc_52155_new_n4896_));
INVX1 INVX1_999 ( .A(sqrto_177_), .Y(u2__abc_52155_new_n4898_));
OR2X2 OR2X2_1 ( .A(aNan), .B(sqrto_76_), .Y(_abc_73687_new_n830_));
OR2X2 OR2X2_10 ( .A(_abc_73687_new_n753_), .B(\a[4] ), .Y(_abc_73687_new_n843_));
OR2X2 OR2X2_100 ( .A(_abc_73687_new_n753_), .B(\a[49] ), .Y(_abc_73687_new_n978_));
OR2X2 OR2X2_1000 ( .A(u2__abc_52155_new_n7457_), .B(u2__abc_52155_new_n7459_), .Y(u2__abc_52155_new_n7460_));
OR2X2 OR2X2_1001 ( .A(u2__abc_52155_new_n7461_), .B(u2__abc_52155_new_n7395_), .Y(u2__abc_52155_new_n7462_));
OR2X2 OR2X2_1002 ( .A(u2__abc_52155_new_n7464_), .B(u2__abc_52155_new_n7380_), .Y(u2__abc_52155_new_n7465_));
OR2X2 OR2X2_1003 ( .A(u2__abc_52155_new_n7463_), .B(u2__abc_52155_new_n7465_), .Y(u2__abc_52155_new_n7466_));
OR2X2 OR2X2_1004 ( .A(u2__abc_52155_new_n7467_), .B(u2__abc_52155_new_n7460_), .Y(u2__abc_52155_new_n7468_));
OR2X2 OR2X2_1005 ( .A(u2__abc_52155_new_n7454_), .B(u2__abc_52155_new_n7468_), .Y(u2__abc_52155_new_n7469_));
OR2X2 OR2X2_1006 ( .A(u2__abc_52155_new_n7471_), .B(u2__abc_52155_new_n7261_), .Y(u2__abc_52155_new_n7472_));
OR2X2 OR2X2_1007 ( .A(u2__abc_52155_new_n7474_), .B(u2__abc_52155_new_n7253_), .Y(u2__abc_52155_new_n7475_));
OR2X2 OR2X2_1008 ( .A(u2__abc_52155_new_n7473_), .B(u2__abc_52155_new_n7475_), .Y(u2__abc_52155_new_n7476_));
OR2X2 OR2X2_1009 ( .A(u2__abc_52155_new_n7478_), .B(u2__abc_52155_new_n7292_), .Y(u2__abc_52155_new_n7479_));
OR2X2 OR2X2_101 ( .A(aNan), .B(sqrto_126_), .Y(_abc_73687_new_n980_));
OR2X2 OR2X2_1010 ( .A(u2__abc_52155_new_n7481_), .B(u2__abc_52155_new_n7287_), .Y(u2__abc_52155_new_n7482_));
OR2X2 OR2X2_1011 ( .A(u2__abc_52155_new_n7480_), .B(u2__abc_52155_new_n7482_), .Y(u2__abc_52155_new_n7483_));
OR2X2 OR2X2_1012 ( .A(u2__abc_52155_new_n7477_), .B(u2__abc_52155_new_n7483_), .Y(u2__abc_52155_new_n7484_));
OR2X2 OR2X2_1013 ( .A(u2__abc_52155_new_n7485_), .B(u2__abc_52155_new_n7316_), .Y(u2__abc_52155_new_n7486_));
OR2X2 OR2X2_1014 ( .A(u2__abc_52155_new_n7488_), .B(u2__abc_52155_new_n7331_), .Y(u2__abc_52155_new_n7489_));
OR2X2 OR2X2_1015 ( .A(u2__abc_52155_new_n7487_), .B(u2__abc_52155_new_n7489_), .Y(u2__abc_52155_new_n7490_));
OR2X2 OR2X2_1016 ( .A(u2__abc_52155_new_n7492_), .B(u2__abc_52155_new_n7355_), .Y(u2__abc_52155_new_n7493_));
OR2X2 OR2X2_1017 ( .A(u2__abc_52155_new_n7495_), .B(u2__abc_52155_new_n7350_), .Y(u2__abc_52155_new_n7496_));
OR2X2 OR2X2_1018 ( .A(u2__abc_52155_new_n7494_), .B(u2__abc_52155_new_n7496_), .Y(u2__abc_52155_new_n7497_));
OR2X2 OR2X2_1019 ( .A(u2__abc_52155_new_n7491_), .B(u2__abc_52155_new_n7497_), .Y(u2__abc_52155_new_n7498_));
OR2X2 OR2X2_102 ( .A(_abc_73687_new_n753_), .B(\a[50] ), .Y(_abc_73687_new_n981_));
OR2X2 OR2X2_1020 ( .A(u2__abc_52155_new_n7499_), .B(u2__abc_52155_new_n7484_), .Y(u2__abc_52155_new_n7500_));
OR2X2 OR2X2_1021 ( .A(u2__abc_52155_new_n7470_), .B(u2__abc_52155_new_n7500_), .Y(u2__abc_52155_new_n7501_));
OR2X2 OR2X2_1022 ( .A(u2__abc_52155_new_n7503_), .B(u2__abc_52155_new_n7164_), .Y(u2__abc_52155_new_n7504_));
OR2X2 OR2X2_1023 ( .A(u2__abc_52155_new_n7506_), .B(u2__abc_52155_new_n7156_), .Y(u2__abc_52155_new_n7507_));
OR2X2 OR2X2_1024 ( .A(u2__abc_52155_new_n7505_), .B(u2__abc_52155_new_n7507_), .Y(u2__abc_52155_new_n7508_));
OR2X2 OR2X2_1025 ( .A(u2__abc_52155_new_n7510_), .B(u2__abc_52155_new_n7133_), .Y(u2__abc_52155_new_n7511_));
OR2X2 OR2X2_1026 ( .A(u2__abc_52155_new_n7513_), .B(u2__abc_52155_new_n7128_), .Y(u2__abc_52155_new_n7514_));
OR2X2 OR2X2_1027 ( .A(u2__abc_52155_new_n7512_), .B(u2__abc_52155_new_n7514_), .Y(u2__abc_52155_new_n7515_));
OR2X2 OR2X2_1028 ( .A(u2__abc_52155_new_n7509_), .B(u2__abc_52155_new_n7515_), .Y(u2__abc_52155_new_n7516_));
OR2X2 OR2X2_1029 ( .A(u2__abc_52155_new_n7518_), .B(u2__abc_52155_new_n7077_), .Y(u2__abc_52155_new_n7519_));
OR2X2 OR2X2_103 ( .A(aNan), .B(sqrto_127_), .Y(_abc_73687_new_n983_));
OR2X2 OR2X2_1030 ( .A(u2__abc_52155_new_n7521_), .B(u2__abc_52155_new_n7062_), .Y(u2__abc_52155_new_n7522_));
OR2X2 OR2X2_1031 ( .A(u2__abc_52155_new_n7520_), .B(u2__abc_52155_new_n7522_), .Y(u2__abc_52155_new_n7523_));
OR2X2 OR2X2_1032 ( .A(u2__abc_52155_new_n7525_), .B(u2__abc_52155_new_n7101_), .Y(u2__abc_52155_new_n7526_));
OR2X2 OR2X2_1033 ( .A(u2__abc_52155_new_n7528_), .B(u2__abc_52155_new_n7096_), .Y(u2__abc_52155_new_n7529_));
OR2X2 OR2X2_1034 ( .A(u2__abc_52155_new_n7527_), .B(u2__abc_52155_new_n7529_), .Y(u2__abc_52155_new_n7530_));
OR2X2 OR2X2_1035 ( .A(u2__abc_52155_new_n7524_), .B(u2__abc_52155_new_n7530_), .Y(u2__abc_52155_new_n7531_));
OR2X2 OR2X2_1036 ( .A(u2__abc_52155_new_n7517_), .B(u2__abc_52155_new_n7531_), .Y(u2__abc_52155_new_n7532_));
OR2X2 OR2X2_1037 ( .A(u2__abc_52155_new_n7534_), .B(u2__abc_52155_new_n6966_), .Y(u2__abc_52155_new_n7535_));
OR2X2 OR2X2_1038 ( .A(u2__abc_52155_new_n7537_), .B(u2__abc_52155_new_n6981_), .Y(u2__abc_52155_new_n7538_));
OR2X2 OR2X2_1039 ( .A(u2__abc_52155_new_n7536_), .B(u2__abc_52155_new_n7538_), .Y(u2__abc_52155_new_n7539_));
OR2X2 OR2X2_104 ( .A(_abc_73687_new_n753_), .B(\a[51] ), .Y(_abc_73687_new_n984_));
OR2X2 OR2X2_1040 ( .A(u2__abc_52155_new_n7541_), .B(u2__abc_52155_new_n6943_), .Y(u2__abc_52155_new_n7542_));
OR2X2 OR2X2_1041 ( .A(u2__abc_52155_new_n7544_), .B(u2__abc_52155_new_n6935_), .Y(u2__abc_52155_new_n7545_));
OR2X2 OR2X2_1042 ( .A(u2__abc_52155_new_n7543_), .B(u2__abc_52155_new_n7545_), .Y(u2__abc_52155_new_n7546_));
OR2X2 OR2X2_1043 ( .A(u2__abc_52155_new_n7540_), .B(u2__abc_52155_new_n7546_), .Y(u2__abc_52155_new_n7547_));
OR2X2 OR2X2_1044 ( .A(u2__abc_52155_new_n7548_), .B(u2__abc_52155_new_n7029_), .Y(u2__abc_52155_new_n7549_));
OR2X2 OR2X2_1045 ( .A(u2__abc_52155_new_n7551_), .B(u2__abc_52155_new_n7044_), .Y(u2__abc_52155_new_n7552_));
OR2X2 OR2X2_1046 ( .A(u2__abc_52155_new_n7550_), .B(u2__abc_52155_new_n7552_), .Y(u2__abc_52155_new_n7553_));
OR2X2 OR2X2_1047 ( .A(u2__abc_52155_new_n7555_), .B(u2__abc_52155_new_n7006_), .Y(u2__abc_52155_new_n7556_));
OR2X2 OR2X2_1048 ( .A(u2__abc_52155_new_n7558_), .B(u2__abc_52155_new_n7001_), .Y(u2__abc_52155_new_n7559_));
OR2X2 OR2X2_1049 ( .A(u2__abc_52155_new_n7559_), .B(u2__abc_52155_new_n7557_), .Y(u2__abc_52155_new_n7560_));
OR2X2 OR2X2_105 ( .A(aNan), .B(sqrto_128_), .Y(_abc_73687_new_n986_));
OR2X2 OR2X2_1050 ( .A(u2__abc_52155_new_n7554_), .B(u2__abc_52155_new_n7560_), .Y(u2__abc_52155_new_n7561_));
OR2X2 OR2X2_1051 ( .A(u2__abc_52155_new_n7562_), .B(u2__abc_52155_new_n7547_), .Y(u2__abc_52155_new_n7563_));
OR2X2 OR2X2_1052 ( .A(u2__abc_52155_new_n7533_), .B(u2__abc_52155_new_n7563_), .Y(u2__abc_52155_new_n7564_));
OR2X2 OR2X2_1053 ( .A(u2__abc_52155_new_n7502_), .B(u2__abc_52155_new_n7564_), .Y(u2__abc_52155_new_n7565_));
OR2X2 OR2X2_1054 ( .A(u2__abc_52155_new_n7567_), .B(u2__abc_52155_new_n3034_), .Y(u2__abc_52155_new_n7568_));
OR2X2 OR2X2_1055 ( .A(u2__abc_52155_new_n7569_), .B(u2__abc_52155_new_n3019_), .Y(u2__abc_52155_new_n7570_));
OR2X2 OR2X2_1056 ( .A(u2__abc_52155_new_n7573_), .B(u2__abc_52155_new_n3005_), .Y(u2__abc_52155_new_n7574_));
OR2X2 OR2X2_1057 ( .A(u2__abc_52155_new_n7572_), .B(u2__abc_52155_new_n7574_), .Y(u2__abc_52155_new_n7575_));
OR2X2 OR2X2_1058 ( .A(u2__abc_52155_new_n3125_), .B(u2_remHiShift_1_), .Y(u2__abc_52155_new_n7585_));
OR2X2 OR2X2_1059 ( .A(u2__abc_52155_new_n7577_), .B(u2__abc_52155_new_n7621_), .Y(u2__abc_52155_new_n7622_));
OR2X2 OR2X2_106 ( .A(_abc_73687_new_n753_), .B(\a[52] ), .Y(_abc_73687_new_n987_));
OR2X2 OR2X2_1060 ( .A(u2__abc_52155_new_n7626_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7627_));
OR2X2 OR2X2_1061 ( .A(u2__abc_52155_new_n7627_), .B(u2__abc_52155_new_n7624_), .Y(u2__abc_52155_new_n7628_));
OR2X2 OR2X2_1062 ( .A(u2__abc_52155_new_n7632_), .B(u2__abc_52155_new_n3003_), .Y(u2__abc_52155_new_n7633_));
OR2X2 OR2X2_1063 ( .A(u2__abc_52155_new_n7586_), .B(u2_remHiShift_0_), .Y(u2__abc_52155_new_n7637_));
OR2X2 OR2X2_1064 ( .A(u2__abc_52155_new_n7640_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7641_));
OR2X2 OR2X2_1065 ( .A(u2__abc_52155_new_n7641_), .B(u2__abc_52155_new_n7639_), .Y(u2__abc_52155_new_n7642_));
OR2X2 OR2X2_1066 ( .A(u2__abc_52155_new_n7646_), .B(u2__abc_52155_new_n7635_), .Y(u2__abc_52155_new_n7647_));
OR2X2 OR2X2_1067 ( .A(u2__abc_52155_new_n7652_), .B(u2__abc_52155_new_n7650_), .Y(u2__abc_52155_new_n7655_));
OR2X2 OR2X2_1068 ( .A(u2__abc_52155_new_n7658_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7659_));
OR2X2 OR2X2_1069 ( .A(u2__abc_52155_new_n7659_), .B(u2__abc_52155_new_n7657_), .Y(u2__abc_52155_new_n7660_));
OR2X2 OR2X2_107 ( .A(aNan), .B(sqrto_129_), .Y(_abc_73687_new_n989_));
OR2X2 OR2X2_1070 ( .A(u2__abc_52155_new_n7664_), .B(u2__abc_52155_new_n7649_), .Y(u2__abc_52155_new_n7665_));
OR2X2 OR2X2_1071 ( .A(u2__abc_52155_new_n7668_), .B(u2__abc_52155_new_n3115_), .Y(u2__abc_52155_new_n7669_));
OR2X2 OR2X2_1072 ( .A(u2__abc_52155_new_n7653_), .B(u2__abc_52155_new_n7669_), .Y(u2__abc_52155_new_n7670_));
OR2X2 OR2X2_1073 ( .A(u2__abc_52155_new_n7672_), .B(u2__abc_52155_new_n7671_), .Y(u2__abc_52155_new_n7673_));
OR2X2 OR2X2_1074 ( .A(u2__abc_52155_new_n7677_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7678_));
OR2X2 OR2X2_1075 ( .A(u2__abc_52155_new_n7678_), .B(u2__abc_52155_new_n7676_), .Y(u2__abc_52155_new_n7679_));
OR2X2 OR2X2_1076 ( .A(u2__abc_52155_new_n7683_), .B(u2__abc_52155_new_n7667_), .Y(u2__abc_52155_new_n7684_));
OR2X2 OR2X2_1077 ( .A(u2__abc_52155_new_n7673_), .B(u2__abc_52155_new_n3122_), .Y(u2__abc_52155_new_n7688_));
OR2X2 OR2X2_1078 ( .A(u2__abc_52155_new_n7688_), .B(u2__abc_52155_new_n7687_), .Y(u2__abc_52155_new_n7689_));
OR2X2 OR2X2_1079 ( .A(u2__abc_52155_new_n7694_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7695_));
OR2X2 OR2X2_108 ( .A(_abc_73687_new_n753_), .B(\a[53] ), .Y(_abc_73687_new_n990_));
OR2X2 OR2X2_1080 ( .A(u2__abc_52155_new_n7695_), .B(u2__abc_52155_new_n7693_), .Y(u2__abc_52155_new_n7696_));
OR2X2 OR2X2_1081 ( .A(u2__abc_52155_new_n7700_), .B(u2__abc_52155_new_n7686_), .Y(u2__abc_52155_new_n7701_));
OR2X2 OR2X2_1082 ( .A(u2__abc_52155_new_n7707_), .B(u2__abc_52155_new_n7704_), .Y(u2__abc_52155_new_n7708_));
OR2X2 OR2X2_1083 ( .A(u2__abc_52155_new_n7706_), .B(u2__abc_52155_new_n3106_), .Y(u2__abc_52155_new_n7709_));
OR2X2 OR2X2_1084 ( .A(u2__abc_52155_new_n7712_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7713_));
OR2X2 OR2X2_1085 ( .A(u2__abc_52155_new_n7713_), .B(u2__abc_52155_new_n7711_), .Y(u2__abc_52155_new_n7714_));
OR2X2 OR2X2_1086 ( .A(u2__abc_52155_new_n7718_), .B(u2__abc_52155_new_n7703_), .Y(u2__abc_52155_new_n7719_));
OR2X2 OR2X2_1087 ( .A(u2__abc_52155_new_n3103_), .B(u2__abc_52155_new_n3108_), .Y(u2__abc_52155_new_n7724_));
OR2X2 OR2X2_1088 ( .A(u2__abc_52155_new_n7723_), .B(u2__abc_52155_new_n7725_), .Y(u2__abc_52155_new_n7726_));
OR2X2 OR2X2_1089 ( .A(u2__abc_52155_new_n7726_), .B(u2__abc_52155_new_n7722_), .Y(u2__abc_52155_new_n7727_));
OR2X2 OR2X2_109 ( .A(aNan), .B(sqrto_130_), .Y(_abc_73687_new_n992_));
OR2X2 OR2X2_1090 ( .A(u2__abc_52155_new_n7732_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7733_));
OR2X2 OR2X2_1091 ( .A(u2__abc_52155_new_n7733_), .B(u2__abc_52155_new_n7731_), .Y(u2__abc_52155_new_n7734_));
OR2X2 OR2X2_1092 ( .A(u2__abc_52155_new_n7738_), .B(u2__abc_52155_new_n7721_), .Y(u2__abc_52155_new_n7739_));
OR2X2 OR2X2_1093 ( .A(u2__abc_52155_new_n7745_), .B(u2__abc_52155_new_n7742_), .Y(u2__abc_52155_new_n7746_));
OR2X2 OR2X2_1094 ( .A(u2__abc_52155_new_n7744_), .B(u2__abc_52155_new_n3100_), .Y(u2__abc_52155_new_n7747_));
OR2X2 OR2X2_1095 ( .A(u2__abc_52155_new_n7750_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7751_));
OR2X2 OR2X2_1096 ( .A(u2__abc_52155_new_n7751_), .B(u2__abc_52155_new_n7749_), .Y(u2__abc_52155_new_n7752_));
OR2X2 OR2X2_1097 ( .A(u2__abc_52155_new_n7757_), .B(u2__abc_52155_new_n7741_), .Y(u2__abc_52155_new_n7758_));
OR2X2 OR2X2_1098 ( .A(u2__abc_52155_new_n7764_), .B(u2__abc_52155_new_n3099_), .Y(u2__abc_52155_new_n7765_));
OR2X2 OR2X2_1099 ( .A(u2__abc_52155_new_n7763_), .B(u2__abc_52155_new_n7765_), .Y(u2__abc_52155_new_n7766_));
OR2X2 OR2X2_11 ( .A(aNan), .B(sqrto_81_), .Y(_abc_73687_new_n845_));
OR2X2 OR2X2_110 ( .A(_abc_73687_new_n753_), .B(\a[54] ), .Y(_abc_73687_new_n993_));
OR2X2 OR2X2_1100 ( .A(u2__abc_52155_new_n7761_), .B(u2__abc_52155_new_n7766_), .Y(u2__abc_52155_new_n7767_));
OR2X2 OR2X2_1101 ( .A(u2__abc_52155_new_n7767_), .B(u2__abc_52155_new_n3086_), .Y(u2__abc_52155_new_n7770_));
OR2X2 OR2X2_1102 ( .A(u2__abc_52155_new_n7773_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7774_));
OR2X2 OR2X2_1103 ( .A(u2__abc_52155_new_n7774_), .B(u2__abc_52155_new_n7772_), .Y(u2__abc_52155_new_n7775_));
OR2X2 OR2X2_1104 ( .A(u2__abc_52155_new_n7779_), .B(u2__abc_52155_new_n7760_), .Y(u2__abc_52155_new_n7780_));
OR2X2 OR2X2_1105 ( .A(u2__abc_52155_new_n7786_), .B(u2__abc_52155_new_n7787_), .Y(u2__abc_52155_new_n7788_));
OR2X2 OR2X2_1106 ( .A(u2__abc_52155_new_n7790_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n7791_));
OR2X2 OR2X2_1107 ( .A(u2__abc_52155_new_n7791_), .B(u2__abc_52155_new_n7789_), .Y(u2__abc_52155_new_n7792_));
OR2X2 OR2X2_1108 ( .A(u2__abc_52155_new_n7796_), .B(u2__abc_52155_new_n7782_), .Y(u2__abc_52155_new_n7797_));
OR2X2 OR2X2_1109 ( .A(u2__abc_52155_new_n7803_), .B(u2__abc_52155_new_n7802_), .Y(u2__abc_52155_new_n7804_));
OR2X2 OR2X2_111 ( .A(aNan), .B(sqrto_131_), .Y(_abc_73687_new_n995_));
OR2X2 OR2X2_1110 ( .A(u2__abc_52155_new_n7804_), .B(u2__abc_52155_new_n3068_), .Y(u2__abc_52155_new_n7805_));
OR2X2 OR2X2_1111 ( .A(u2__abc_52155_new_n7810_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7811_));
OR2X2 OR2X2_1112 ( .A(u2__abc_52155_new_n7811_), .B(u2__abc_52155_new_n7809_), .Y(u2__abc_52155_new_n7812_));
OR2X2 OR2X2_1113 ( .A(u2__abc_52155_new_n7816_), .B(u2__abc_52155_new_n7799_), .Y(u2__abc_52155_new_n7817_));
OR2X2 OR2X2_1114 ( .A(u2__abc_52155_new_n7824_), .B(u2__abc_52155_new_n7825_), .Y(u2__abc_52155_new_n7826_));
OR2X2 OR2X2_1115 ( .A(u2__abc_52155_new_n7828_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7829_));
OR2X2 OR2X2_1116 ( .A(u2__abc_52155_new_n7829_), .B(u2__abc_52155_new_n7827_), .Y(u2__abc_52155_new_n7830_));
OR2X2 OR2X2_1117 ( .A(u2__abc_52155_new_n7834_), .B(u2__abc_52155_new_n7819_), .Y(u2__abc_52155_new_n7835_));
OR2X2 OR2X2_1118 ( .A(u2__abc_52155_new_n7839_), .B(u2__abc_52155_new_n3073_), .Y(u2__abc_52155_new_n7840_));
OR2X2 OR2X2_1119 ( .A(u2__abc_52155_new_n7841_), .B(u2__abc_52155_new_n3060_), .Y(u2__abc_52155_new_n7842_));
OR2X2 OR2X2_112 ( .A(_abc_73687_new_n753_), .B(\a[55] ), .Y(_abc_73687_new_n996_));
OR2X2 OR2X2_1120 ( .A(u2__abc_52155_new_n7847_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7848_));
OR2X2 OR2X2_1121 ( .A(u2__abc_52155_new_n7848_), .B(u2__abc_52155_new_n7846_), .Y(u2__abc_52155_new_n7849_));
OR2X2 OR2X2_1122 ( .A(u2__abc_52155_new_n7853_), .B(u2__abc_52155_new_n7837_), .Y(u2__abc_52155_new_n7854_));
OR2X2 OR2X2_1123 ( .A(u2__abc_52155_new_n7862_), .B(u2__abc_52155_new_n7859_), .Y(u2__abc_52155_new_n7863_));
OR2X2 OR2X2_1124 ( .A(u2__abc_52155_new_n7865_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n7866_));
OR2X2 OR2X2_1125 ( .A(u2__abc_52155_new_n7866_), .B(u2__abc_52155_new_n7864_), .Y(u2__abc_52155_new_n7867_));
OR2X2 OR2X2_1126 ( .A(u2__abc_52155_new_n7871_), .B(u2__abc_52155_new_n7856_), .Y(u2__abc_52155_new_n7872_));
OR2X2 OR2X2_1127 ( .A(u2__abc_52155_new_n7840_), .B(u2__abc_52155_new_n7875_), .Y(u2__abc_52155_new_n7876_));
OR2X2 OR2X2_1128 ( .A(u2__abc_52155_new_n7877_), .B(u2__abc_52155_new_n3049_), .Y(u2__abc_52155_new_n7878_));
OR2X2 OR2X2_1129 ( .A(u2__abc_52155_new_n7881_), .B(u2__abc_52155_new_n3040_), .Y(u2__abc_52155_new_n7882_));
OR2X2 OR2X2_113 ( .A(aNan), .B(sqrto_132_), .Y(_abc_73687_new_n998_));
OR2X2 OR2X2_1130 ( .A(u2__abc_52155_new_n7887_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7888_));
OR2X2 OR2X2_1131 ( .A(u2__abc_52155_new_n7888_), .B(u2__abc_52155_new_n7886_), .Y(u2__abc_52155_new_n7889_));
OR2X2 OR2X2_1132 ( .A(u2__abc_52155_new_n7894_), .B(u2__abc_52155_new_n7874_), .Y(u2__abc_52155_new_n7895_));
OR2X2 OR2X2_1133 ( .A(u2__abc_52155_new_n7900_), .B(u2__abc_52155_new_n3046_), .Y(u2__abc_52155_new_n7901_));
OR2X2 OR2X2_1134 ( .A(u2__abc_52155_new_n7899_), .B(u2__abc_52155_new_n3045_), .Y(u2__abc_52155_new_n7902_));
OR2X2 OR2X2_1135 ( .A(u2__abc_52155_new_n7623_), .B(u2__abc_52155_new_n7903_), .Y(u2__abc_52155_new_n7904_));
OR2X2 OR2X2_1136 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_13_), .Y(u2__abc_52155_new_n7905_));
OR2X2 OR2X2_1137 ( .A(u2__abc_52155_new_n7906_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n7907_));
OR2X2 OR2X2_1138 ( .A(u2__abc_52155_new_n7911_), .B(u2__abc_52155_new_n7897_), .Y(u2__abc_52155_new_n7912_));
OR2X2 OR2X2_1139 ( .A(u2__abc_52155_new_n7838_), .B(u2__abc_52155_new_n3073_), .Y(u2__abc_52155_new_n7917_));
OR2X2 OR2X2_114 ( .A(_abc_73687_new_n753_), .B(\a[56] ), .Y(_abc_73687_new_n999_));
OR2X2 OR2X2_1140 ( .A(u2__abc_52155_new_n7920_), .B(u2__abc_52155_new_n3146_), .Y(u2__abc_52155_new_n7921_));
OR2X2 OR2X2_1141 ( .A(u2__abc_52155_new_n7923_), .B(u2__abc_52155_new_n3044_), .Y(u2__abc_52155_new_n7924_));
OR2X2 OR2X2_1142 ( .A(u2__abc_52155_new_n7922_), .B(u2__abc_52155_new_n7924_), .Y(u2__abc_52155_new_n7925_));
OR2X2 OR2X2_1143 ( .A(u2__abc_52155_new_n7929_), .B(u2__abc_52155_new_n3243_), .Y(u2__abc_52155_new_n7930_));
OR2X2 OR2X2_1144 ( .A(u2__abc_52155_new_n7935_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7936_));
OR2X2 OR2X2_1145 ( .A(u2__abc_52155_new_n7936_), .B(u2__abc_52155_new_n7934_), .Y(u2__abc_52155_new_n7937_));
OR2X2 OR2X2_1146 ( .A(u2__abc_52155_new_n7941_), .B(u2__abc_52155_new_n7914_), .Y(u2__abc_52155_new_n7942_));
OR2X2 OR2X2_1147 ( .A(u2__abc_52155_new_n7948_), .B(u2__abc_52155_new_n7949_), .Y(u2__abc_52155_new_n7950_));
OR2X2 OR2X2_1148 ( .A(u2__abc_52155_new_n7952_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n7953_));
OR2X2 OR2X2_1149 ( .A(u2__abc_52155_new_n7953_), .B(u2__abc_52155_new_n7951_), .Y(u2__abc_52155_new_n7954_));
OR2X2 OR2X2_115 ( .A(aNan), .B(sqrto_133_), .Y(_abc_73687_new_n1001_));
OR2X2 OR2X2_1150 ( .A(u2__abc_52155_new_n7958_), .B(u2__abc_52155_new_n7944_), .Y(u2__abc_52155_new_n7959_));
OR2X2 OR2X2_1151 ( .A(u2__abc_52155_new_n7963_), .B(u2__abc_52155_new_n3245_), .Y(u2__abc_52155_new_n7964_));
OR2X2 OR2X2_1152 ( .A(u2__abc_52155_new_n7964_), .B(u2__abc_52155_new_n7962_), .Y(u2__abc_52155_new_n7965_));
OR2X2 OR2X2_1153 ( .A(u2__abc_52155_new_n7970_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7971_));
OR2X2 OR2X2_1154 ( .A(u2__abc_52155_new_n7971_), .B(u2__abc_52155_new_n7969_), .Y(u2__abc_52155_new_n7972_));
OR2X2 OR2X2_1155 ( .A(u2__abc_52155_new_n7976_), .B(u2__abc_52155_new_n7961_), .Y(u2__abc_52155_new_n7977_));
OR2X2 OR2X2_1156 ( .A(u2__abc_52155_new_n7983_), .B(u2__abc_52155_new_n7985_), .Y(u2__abc_52155_new_n7986_));
OR2X2 OR2X2_1157 ( .A(u2__abc_52155_new_n7988_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n7989_));
OR2X2 OR2X2_1158 ( .A(u2__abc_52155_new_n7989_), .B(u2__abc_52155_new_n7987_), .Y(u2__abc_52155_new_n7990_));
OR2X2 OR2X2_1159 ( .A(u2__abc_52155_new_n7994_), .B(u2__abc_52155_new_n7979_), .Y(u2__abc_52155_new_n7995_));
OR2X2 OR2X2_116 ( .A(_abc_73687_new_n753_), .B(\a[57] ), .Y(_abc_73687_new_n1002_));
OR2X2 OR2X2_1160 ( .A(u2__abc_52155_new_n7999_), .B(u2__abc_52155_new_n3248_), .Y(u2__abc_52155_new_n8000_));
OR2X2 OR2X2_1161 ( .A(u2__abc_52155_new_n8000_), .B(u2__abc_52155_new_n3237_), .Y(u2__abc_52155_new_n8001_));
OR2X2 OR2X2_1162 ( .A(u2__abc_52155_new_n8002_), .B(u2__abc_52155_new_n3233_), .Y(u2__abc_52155_new_n8003_));
OR2X2 OR2X2_1163 ( .A(u2__abc_52155_new_n8007_), .B(u2__abc_52155_new_n8006_), .Y(u2__abc_52155_new_n8008_));
OR2X2 OR2X2_1164 ( .A(u2__abc_52155_new_n8008_), .B(u2__abc_52155_new_n7998_), .Y(u2__abc_52155_new_n8009_));
OR2X2 OR2X2_1165 ( .A(u2__abc_52155_new_n8014_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8015_));
OR2X2 OR2X2_1166 ( .A(u2__abc_52155_new_n8015_), .B(u2__abc_52155_new_n8013_), .Y(u2__abc_52155_new_n8016_));
OR2X2 OR2X2_1167 ( .A(u2__abc_52155_new_n8020_), .B(u2__abc_52155_new_n7997_), .Y(u2__abc_52155_new_n8021_));
OR2X2 OR2X2_1168 ( .A(u2__abc_52155_new_n8027_), .B(u2__abc_52155_new_n8024_), .Y(u2__abc_52155_new_n8028_));
OR2X2 OR2X2_1169 ( .A(u2__abc_52155_new_n8026_), .B(u2__abc_52155_new_n3268_), .Y(u2__abc_52155_new_n8029_));
OR2X2 OR2X2_117 ( .A(aNan), .B(sqrto_134_), .Y(_abc_73687_new_n1004_));
OR2X2 OR2X2_1170 ( .A(u2__abc_52155_new_n8032_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8033_));
OR2X2 OR2X2_1171 ( .A(u2__abc_52155_new_n8033_), .B(u2__abc_52155_new_n8031_), .Y(u2__abc_52155_new_n8034_));
OR2X2 OR2X2_1172 ( .A(u2__abc_52155_new_n8038_), .B(u2__abc_52155_new_n8023_), .Y(u2__abc_52155_new_n8039_));
OR2X2 OR2X2_1173 ( .A(u2__abc_52155_new_n3265_), .B(u2__abc_52155_new_n3270_), .Y(u2__abc_52155_new_n8044_));
OR2X2 OR2X2_1174 ( .A(u2__abc_52155_new_n8046_), .B(u2__abc_52155_new_n3267_), .Y(u2__abc_52155_new_n8047_));
OR2X2 OR2X2_1175 ( .A(u2__abc_52155_new_n8048_), .B(u2__abc_52155_new_n8043_), .Y(u2__abc_52155_new_n8049_));
OR2X2 OR2X2_1176 ( .A(u2__abc_52155_new_n8053_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8054_));
OR2X2 OR2X2_1177 ( .A(u2__abc_52155_new_n8054_), .B(u2__abc_52155_new_n8042_), .Y(u2__abc_52155_new_n8055_));
OR2X2 OR2X2_1178 ( .A(u2__abc_52155_new_n8059_), .B(u2__abc_52155_new_n8041_), .Y(u2__abc_52155_new_n8060_));
OR2X2 OR2X2_1179 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_21_), .Y(u2__abc_52155_new_n8063_));
OR2X2 OR2X2_118 ( .A(_abc_73687_new_n753_), .B(\a[58] ), .Y(_abc_73687_new_n1005_));
OR2X2 OR2X2_1180 ( .A(u2__abc_52155_new_n8067_), .B(u2__abc_52155_new_n8069_), .Y(u2__abc_52155_new_n8070_));
OR2X2 OR2X2_1181 ( .A(u2__abc_52155_new_n7623_), .B(u2__abc_52155_new_n8070_), .Y(u2__abc_52155_new_n8071_));
OR2X2 OR2X2_1182 ( .A(u2__abc_52155_new_n8072_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8073_));
OR2X2 OR2X2_1183 ( .A(u2__abc_52155_new_n8077_), .B(u2__abc_52155_new_n8062_), .Y(u2__abc_52155_new_n8078_));
OR2X2 OR2X2_1184 ( .A(u2__abc_52155_new_n8045_), .B(u2__abc_52155_new_n3267_), .Y(u2__abc_52155_new_n8085_));
OR2X2 OR2X2_1185 ( .A(u2__abc_52155_new_n8085_), .B(u2__abc_52155_new_n3263_), .Y(u2__abc_52155_new_n8086_));
OR2X2 OR2X2_1186 ( .A(u2__abc_52155_new_n8064_), .B(u2__abc_52155_new_n3261_), .Y(u2__abc_52155_new_n8087_));
OR2X2 OR2X2_1187 ( .A(u2__abc_52155_new_n8092_), .B(u2__abc_52155_new_n3192_), .Y(u2__abc_52155_new_n8093_));
OR2X2 OR2X2_1188 ( .A(u2__abc_52155_new_n8098_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8099_));
OR2X2 OR2X2_1189 ( .A(u2__abc_52155_new_n8099_), .B(u2__abc_52155_new_n8097_), .Y(u2__abc_52155_new_n8100_));
OR2X2 OR2X2_119 ( .A(aNan), .B(sqrto_135_), .Y(_abc_73687_new_n1007_));
OR2X2 OR2X2_1190 ( .A(u2__abc_52155_new_n8104_), .B(u2__abc_52155_new_n8080_), .Y(u2__abc_52155_new_n8105_));
OR2X2 OR2X2_1191 ( .A(u2__abc_52155_new_n8110_), .B(u2__abc_52155_new_n3185_), .Y(u2__abc_52155_new_n8111_));
OR2X2 OR2X2_1192 ( .A(u2__abc_52155_new_n8109_), .B(u2__abc_52155_new_n8112_), .Y(u2__abc_52155_new_n8113_));
OR2X2 OR2X2_1193 ( .A(u2__abc_52155_new_n8115_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8116_));
OR2X2 OR2X2_1194 ( .A(u2__abc_52155_new_n8116_), .B(u2__abc_52155_new_n8108_), .Y(u2__abc_52155_new_n8117_));
OR2X2 OR2X2_1195 ( .A(u2__abc_52155_new_n8121_), .B(u2__abc_52155_new_n8107_), .Y(u2__abc_52155_new_n8122_));
OR2X2 OR2X2_1196 ( .A(u2__abc_52155_new_n8128_), .B(u2__abc_52155_new_n3183_), .Y(u2__abc_52155_new_n8129_));
OR2X2 OR2X2_1197 ( .A(u2__abc_52155_new_n8130_), .B(u2__abc_52155_new_n8126_), .Y(u2__abc_52155_new_n8131_));
OR2X2 OR2X2_1198 ( .A(u2__abc_52155_new_n8135_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8136_));
OR2X2 OR2X2_1199 ( .A(u2__abc_52155_new_n8136_), .B(u2__abc_52155_new_n8125_), .Y(u2__abc_52155_new_n8137_));
OR2X2 OR2X2_12 ( .A(_abc_73687_new_n753_), .B(\a[5] ), .Y(_abc_73687_new_n846_));
OR2X2 OR2X2_120 ( .A(_abc_73687_new_n753_), .B(\a[59] ), .Y(_abc_73687_new_n1008_));
OR2X2 OR2X2_1200 ( .A(u2__abc_52155_new_n8141_), .B(u2__abc_52155_new_n8124_), .Y(u2__abc_52155_new_n8142_));
OR2X2 OR2X2_1201 ( .A(u2__abc_52155_new_n8148_), .B(u2__abc_52155_new_n8150_), .Y(u2__abc_52155_new_n8151_));
OR2X2 OR2X2_1202 ( .A(u2__abc_52155_new_n8153_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8154_));
OR2X2 OR2X2_1203 ( .A(u2__abc_52155_new_n8154_), .B(u2__abc_52155_new_n8152_), .Y(u2__abc_52155_new_n8155_));
OR2X2 OR2X2_1204 ( .A(u2__abc_52155_new_n8159_), .B(u2__abc_52155_new_n8144_), .Y(u2__abc_52155_new_n8160_));
OR2X2 OR2X2_1205 ( .A(u2__abc_52155_new_n8127_), .B(u2__abc_52155_new_n3183_), .Y(u2__abc_52155_new_n8166_));
OR2X2 OR2X2_1206 ( .A(u2__abc_52155_new_n8166_), .B(u2__abc_52155_new_n3177_), .Y(u2__abc_52155_new_n8167_));
OR2X2 OR2X2_1207 ( .A(u2__abc_52155_new_n8145_), .B(u2__abc_52155_new_n3175_), .Y(u2__abc_52155_new_n8168_));
OR2X2 OR2X2_1208 ( .A(u2__abc_52155_new_n8172_), .B(u2__abc_52155_new_n3223_), .Y(u2__abc_52155_new_n8173_));
OR2X2 OR2X2_1209 ( .A(u2__abc_52155_new_n8177_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8178_));
OR2X2 OR2X2_121 ( .A(aNan), .B(sqrto_136_), .Y(_abc_73687_new_n1010_));
OR2X2 OR2X2_1210 ( .A(u2__abc_52155_new_n8178_), .B(u2__abc_52155_new_n8163_), .Y(u2__abc_52155_new_n8179_));
OR2X2 OR2X2_1211 ( .A(u2__abc_52155_new_n8183_), .B(u2__abc_52155_new_n8162_), .Y(u2__abc_52155_new_n8184_));
OR2X2 OR2X2_1212 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_27_), .Y(u2__abc_52155_new_n8187_));
OR2X2 OR2X2_1213 ( .A(u2__abc_52155_new_n8191_), .B(u2__abc_52155_new_n8192_), .Y(u2__abc_52155_new_n8193_));
OR2X2 OR2X2_1214 ( .A(u2__abc_52155_new_n7623_), .B(u2__abc_52155_new_n8193_), .Y(u2__abc_52155_new_n8194_));
OR2X2 OR2X2_1215 ( .A(u2__abc_52155_new_n8195_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8196_));
OR2X2 OR2X2_1216 ( .A(u2__abc_52155_new_n8200_), .B(u2__abc_52155_new_n8186_), .Y(u2__abc_52155_new_n8201_));
OR2X2 OR2X2_1217 ( .A(u2__abc_52155_new_n8205_), .B(u2__abc_52155_new_n3214_), .Y(u2__abc_52155_new_n8206_));
OR2X2 OR2X2_1218 ( .A(u2__abc_52155_new_n8207_), .B(u2__abc_52155_new_n3201_), .Y(u2__abc_52155_new_n8208_));
OR2X2 OR2X2_1219 ( .A(u2__abc_52155_new_n8211_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n8212_));
OR2X2 OR2X2_122 ( .A(_abc_73687_new_n753_), .B(\a[60] ), .Y(_abc_73687_new_n1011_));
OR2X2 OR2X2_1220 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_28_), .Y(u2__abc_52155_new_n8213_));
OR2X2 OR2X2_1221 ( .A(u2__abc_52155_new_n8214_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8215_));
OR2X2 OR2X2_1222 ( .A(u2__abc_52155_new_n8220_), .B(u2__abc_52155_new_n8203_), .Y(u2__abc_52155_new_n8221_));
OR2X2 OR2X2_1223 ( .A(u2__abc_52155_new_n8225_), .B(u2__abc_52155_new_n3208_), .Y(u2__abc_52155_new_n8226_));
OR2X2 OR2X2_1224 ( .A(u2__abc_52155_new_n8224_), .B(u2__abc_52155_new_n8227_), .Y(u2__abc_52155_new_n8228_));
OR2X2 OR2X2_1225 ( .A(u2__abc_52155_new_n8231_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8232_));
OR2X2 OR2X2_1226 ( .A(u2__abc_52155_new_n8230_), .B(u2__abc_52155_new_n8232_), .Y(u2__abc_52155_new_n8233_));
OR2X2 OR2X2_1227 ( .A(u2__abc_52155_new_n8237_), .B(u2__abc_52155_new_n8223_), .Y(u2__abc_52155_new_n8238_));
OR2X2 OR2X2_1228 ( .A(u2__abc_52155_new_n8204_), .B(u2__abc_52155_new_n3214_), .Y(u2__abc_52155_new_n8241_));
OR2X2 OR2X2_1229 ( .A(u2__abc_52155_new_n8244_), .B(u2__abc_52155_new_n3206_), .Y(u2__abc_52155_new_n8245_));
OR2X2 OR2X2_123 ( .A(aNan), .B(sqrto_137_), .Y(_abc_73687_new_n1013_));
OR2X2 OR2X2_1230 ( .A(u2__abc_52155_new_n8243_), .B(u2__abc_52155_new_n8245_), .Y(u2__abc_52155_new_n8246_));
OR2X2 OR2X2_1231 ( .A(u2__abc_52155_new_n8247_), .B(u2__abc_52155_new_n8246_), .Y(u2__abc_52155_new_n8248_));
OR2X2 OR2X2_1232 ( .A(u2__abc_52155_new_n8248_), .B(u2__abc_52155_new_n3523_), .Y(u2__abc_52155_new_n8251_));
OR2X2 OR2X2_1233 ( .A(u2__abc_52155_new_n8254_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8255_));
OR2X2 OR2X2_1234 ( .A(u2__abc_52155_new_n8255_), .B(u2__abc_52155_new_n8253_), .Y(u2__abc_52155_new_n8256_));
OR2X2 OR2X2_1235 ( .A(u2__abc_52155_new_n8260_), .B(u2__abc_52155_new_n8240_), .Y(u2__abc_52155_new_n8261_));
OR2X2 OR2X2_1236 ( .A(u2__abc_52155_new_n8265_), .B(u2__abc_52155_new_n8264_), .Y(u2__abc_52155_new_n8266_));
OR2X2 OR2X2_1237 ( .A(u2__abc_52155_new_n8267_), .B(u2__abc_52155_new_n3530_), .Y(u2__abc_52155_new_n8268_));
OR2X2 OR2X2_1238 ( .A(u2__abc_52155_new_n8271_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8272_));
OR2X2 OR2X2_1239 ( .A(u2__abc_52155_new_n8270_), .B(u2__abc_52155_new_n8272_), .Y(u2__abc_52155_new_n8273_));
OR2X2 OR2X2_124 ( .A(_abc_73687_new_n753_), .B(\a[61] ), .Y(_abc_73687_new_n1014_));
OR2X2 OR2X2_1240 ( .A(u2__abc_52155_new_n8277_), .B(u2__abc_52155_new_n8263_), .Y(u2__abc_52155_new_n8278_));
OR2X2 OR2X2_1241 ( .A(u2__abc_52155_new_n8283_), .B(u2__abc_52155_new_n3525_), .Y(u2__abc_52155_new_n8284_));
OR2X2 OR2X2_1242 ( .A(u2__abc_52155_new_n8284_), .B(u2__abc_52155_new_n8282_), .Y(u2__abc_52155_new_n8285_));
OR2X2 OR2X2_1243 ( .A(u2__abc_52155_new_n8289_), .B(u2__abc_52155_new_n8281_), .Y(u2__abc_52155_new_n8290_));
OR2X2 OR2X2_1244 ( .A(u2__abc_52155_new_n8290_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8291_));
OR2X2 OR2X2_1245 ( .A(u2__abc_52155_new_n8295_), .B(u2__abc_52155_new_n8280_), .Y(u2__abc_52155_new_n8296_));
OR2X2 OR2X2_1246 ( .A(u2__abc_52155_new_n8304_), .B(u2__abc_52155_new_n8302_), .Y(u2__abc_52155_new_n8305_));
OR2X2 OR2X2_1247 ( .A(u2__abc_52155_new_n8307_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8308_));
OR2X2 OR2X2_1248 ( .A(u2__abc_52155_new_n8306_), .B(u2__abc_52155_new_n8308_), .Y(u2__abc_52155_new_n8309_));
OR2X2 OR2X2_1249 ( .A(u2__abc_52155_new_n8313_), .B(u2__abc_52155_new_n8298_), .Y(u2__abc_52155_new_n8314_));
OR2X2 OR2X2_125 ( .A(aNan), .B(sqrto_138_), .Y(_abc_73687_new_n1016_));
OR2X2 OR2X2_1250 ( .A(u2__abc_52155_new_n8318_), .B(u2__abc_52155_new_n3528_), .Y(u2__abc_52155_new_n8319_));
OR2X2 OR2X2_1251 ( .A(u2__abc_52155_new_n8319_), .B(u2__abc_52155_new_n3517_), .Y(u2__abc_52155_new_n8320_));
OR2X2 OR2X2_1252 ( .A(u2__abc_52155_new_n8321_), .B(u2__abc_52155_new_n3513_), .Y(u2__abc_52155_new_n8322_));
OR2X2 OR2X2_1253 ( .A(u2__abc_52155_new_n8326_), .B(u2__abc_52155_new_n8325_), .Y(u2__abc_52155_new_n8327_));
OR2X2 OR2X2_1254 ( .A(u2__abc_52155_new_n8327_), .B(u2__abc_52155_new_n8317_), .Y(u2__abc_52155_new_n8328_));
OR2X2 OR2X2_1255 ( .A(u2__abc_52155_new_n8331_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n8332_));
OR2X2 OR2X2_1256 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_34_), .Y(u2__abc_52155_new_n8333_));
OR2X2 OR2X2_1257 ( .A(u2__abc_52155_new_n8334_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8335_));
OR2X2 OR2X2_1258 ( .A(u2__abc_52155_new_n8339_), .B(u2__abc_52155_new_n8316_), .Y(u2__abc_52155_new_n8340_));
OR2X2 OR2X2_1259 ( .A(u2__abc_52155_new_n8346_), .B(u2__abc_52155_new_n8343_), .Y(u2__abc_52155_new_n8347_));
OR2X2 OR2X2_126 ( .A(_abc_73687_new_n753_), .B(\a[62] ), .Y(_abc_73687_new_n1017_));
OR2X2 OR2X2_1260 ( .A(u2__abc_52155_new_n8345_), .B(u2__abc_52155_new_n3548_), .Y(u2__abc_52155_new_n8348_));
OR2X2 OR2X2_1261 ( .A(u2__abc_52155_new_n8351_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8352_));
OR2X2 OR2X2_1262 ( .A(u2__abc_52155_new_n8350_), .B(u2__abc_52155_new_n8352_), .Y(u2__abc_52155_new_n8353_));
OR2X2 OR2X2_1263 ( .A(u2__abc_52155_new_n8357_), .B(u2__abc_52155_new_n8342_), .Y(u2__abc_52155_new_n8358_));
OR2X2 OR2X2_1264 ( .A(u2__abc_52155_new_n3545_), .B(u2__abc_52155_new_n3550_), .Y(u2__abc_52155_new_n8363_));
OR2X2 OR2X2_1265 ( .A(u2__abc_52155_new_n8365_), .B(u2__abc_52155_new_n3547_), .Y(u2__abc_52155_new_n8366_));
OR2X2 OR2X2_1266 ( .A(u2__abc_52155_new_n8367_), .B(u2__abc_52155_new_n8362_), .Y(u2__abc_52155_new_n8368_));
OR2X2 OR2X2_1267 ( .A(u2__abc_52155_new_n8372_), .B(u2__abc_52155_new_n8361_), .Y(u2__abc_52155_new_n8373_));
OR2X2 OR2X2_1268 ( .A(u2__abc_52155_new_n8373_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8374_));
OR2X2 OR2X2_1269 ( .A(u2__abc_52155_new_n8378_), .B(u2__abc_52155_new_n8360_), .Y(u2__abc_52155_new_n8379_));
OR2X2 OR2X2_127 ( .A(aNan), .B(sqrto_139_), .Y(_abc_73687_new_n1019_));
OR2X2 OR2X2_1270 ( .A(u2__abc_52155_new_n8383_), .B(u2__abc_52155_new_n3542_), .Y(u2__abc_52155_new_n8384_));
OR2X2 OR2X2_1271 ( .A(u2__abc_52155_new_n8386_), .B(u2__abc_52155_new_n8385_), .Y(u2__abc_52155_new_n8387_));
OR2X2 OR2X2_1272 ( .A(u2__abc_52155_new_n8390_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8391_));
OR2X2 OR2X2_1273 ( .A(u2__abc_52155_new_n8389_), .B(u2__abc_52155_new_n8391_), .Y(u2__abc_52155_new_n8392_));
OR2X2 OR2X2_1274 ( .A(u2__abc_52155_new_n8396_), .B(u2__abc_52155_new_n8381_), .Y(u2__abc_52155_new_n8397_));
OR2X2 OR2X2_1275 ( .A(u2__abc_52155_new_n8364_), .B(u2__abc_52155_new_n3547_), .Y(u2__abc_52155_new_n8402_));
OR2X2 OR2X2_1276 ( .A(u2__abc_52155_new_n8402_), .B(u2__abc_52155_new_n3543_), .Y(u2__abc_52155_new_n8403_));
OR2X2 OR2X2_1277 ( .A(u2__abc_52155_new_n8382_), .B(u2__abc_52155_new_n3541_), .Y(u2__abc_52155_new_n8404_));
OR2X2 OR2X2_1278 ( .A(u2__abc_52155_new_n8409_), .B(u2__abc_52155_new_n8408_), .Y(u2__abc_52155_new_n8410_));
OR2X2 OR2X2_1279 ( .A(u2__abc_52155_new_n8410_), .B(u2__abc_52155_new_n3465_), .Y(u2__abc_52155_new_n8411_));
OR2X2 OR2X2_128 ( .A(_abc_73687_new_n753_), .B(\a[63] ), .Y(_abc_73687_new_n1020_));
OR2X2 OR2X2_1280 ( .A(u2__abc_52155_new_n8414_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n8415_));
OR2X2 OR2X2_1281 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_38_), .Y(u2__abc_52155_new_n8416_));
OR2X2 OR2X2_1282 ( .A(u2__abc_52155_new_n8417_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8418_));
OR2X2 OR2X2_1283 ( .A(u2__abc_52155_new_n8422_), .B(u2__abc_52155_new_n8399_), .Y(u2__abc_52155_new_n8423_));
OR2X2 OR2X2_1284 ( .A(u2__abc_52155_new_n8429_), .B(u2__abc_52155_new_n8430_), .Y(u2__abc_52155_new_n8431_));
OR2X2 OR2X2_1285 ( .A(u2__abc_52155_new_n8433_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8434_));
OR2X2 OR2X2_1286 ( .A(u2__abc_52155_new_n8432_), .B(u2__abc_52155_new_n8434_), .Y(u2__abc_52155_new_n8435_));
OR2X2 OR2X2_1287 ( .A(u2__abc_52155_new_n8439_), .B(u2__abc_52155_new_n8425_), .Y(u2__abc_52155_new_n8440_));
OR2X2 OR2X2_1288 ( .A(u2__abc_52155_new_n8444_), .B(u2__abc_52155_new_n3467_), .Y(u2__abc_52155_new_n8445_));
OR2X2 OR2X2_1289 ( .A(u2__abc_52155_new_n8445_), .B(u2__abc_52155_new_n8443_), .Y(u2__abc_52155_new_n8446_));
OR2X2 OR2X2_129 ( .A(aNan), .B(sqrto_140_), .Y(_abc_73687_new_n1022_));
OR2X2 OR2X2_1290 ( .A(u2__abc_52155_new_n8449_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n8450_));
OR2X2 OR2X2_1291 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_40_), .Y(u2__abc_52155_new_n8451_));
OR2X2 OR2X2_1292 ( .A(u2__abc_52155_new_n8452_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8453_));
OR2X2 OR2X2_1293 ( .A(u2__abc_52155_new_n8457_), .B(u2__abc_52155_new_n8442_), .Y(u2__abc_52155_new_n8458_));
OR2X2 OR2X2_1294 ( .A(u2__abc_52155_new_n8462_), .B(u2__abc_52155_new_n3456_), .Y(u2__abc_52155_new_n8463_));
OR2X2 OR2X2_1295 ( .A(u2__abc_52155_new_n8465_), .B(u2__abc_52155_new_n8464_), .Y(u2__abc_52155_new_n8466_));
OR2X2 OR2X2_1296 ( .A(u2__abc_52155_new_n8469_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8470_));
OR2X2 OR2X2_1297 ( .A(u2__abc_52155_new_n8468_), .B(u2__abc_52155_new_n8470_), .Y(u2__abc_52155_new_n8471_));
OR2X2 OR2X2_1298 ( .A(u2__abc_52155_new_n8475_), .B(u2__abc_52155_new_n8460_), .Y(u2__abc_52155_new_n8476_));
OR2X2 OR2X2_1299 ( .A(u2__abc_52155_new_n8480_), .B(u2__abc_52155_new_n3470_), .Y(u2__abc_52155_new_n8481_));
OR2X2 OR2X2_13 ( .A(aNan), .B(sqrto_82_), .Y(_abc_73687_new_n848_));
OR2X2 OR2X2_130 ( .A(_abc_73687_new_n753_), .B(\a[64] ), .Y(_abc_73687_new_n1023_));
OR2X2 OR2X2_1300 ( .A(u2__abc_52155_new_n8481_), .B(u2__abc_52155_new_n3457_), .Y(u2__abc_52155_new_n8482_));
OR2X2 OR2X2_1301 ( .A(u2__abc_52155_new_n8461_), .B(u2__abc_52155_new_n3455_), .Y(u2__abc_52155_new_n8483_));
OR2X2 OR2X2_1302 ( .A(u2__abc_52155_new_n8487_), .B(u2__abc_52155_new_n8486_), .Y(u2__abc_52155_new_n8488_));
OR2X2 OR2X2_1303 ( .A(u2__abc_52155_new_n8488_), .B(u2__abc_52155_new_n3503_), .Y(u2__abc_52155_new_n8489_));
OR2X2 OR2X2_1304 ( .A(u2__abc_52155_new_n8493_), .B(u2__abc_52155_new_n8479_), .Y(u2__abc_52155_new_n8494_));
OR2X2 OR2X2_1305 ( .A(u2__abc_52155_new_n8494_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8495_));
OR2X2 OR2X2_1306 ( .A(u2__abc_52155_new_n8499_), .B(u2__abc_52155_new_n8478_), .Y(u2__abc_52155_new_n8500_));
OR2X2 OR2X2_1307 ( .A(u2__abc_52155_new_n8507_), .B(u2__abc_52155_new_n8504_), .Y(u2__abc_52155_new_n8508_));
OR2X2 OR2X2_1308 ( .A(u2__abc_52155_new_n8510_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8511_));
OR2X2 OR2X2_1309 ( .A(u2__abc_52155_new_n8509_), .B(u2__abc_52155_new_n8511_), .Y(u2__abc_52155_new_n8512_));
OR2X2 OR2X2_131 ( .A(aNan), .B(sqrto_141_), .Y(_abc_73687_new_n1025_));
OR2X2 OR2X2_1310 ( .A(u2__abc_52155_new_n8516_), .B(u2__abc_52155_new_n8502_), .Y(u2__abc_52155_new_n8517_));
OR2X2 OR2X2_1311 ( .A(u2__abc_52155_new_n8521_), .B(u2__abc_52155_new_n3494_), .Y(u2__abc_52155_new_n8522_));
OR2X2 OR2X2_1312 ( .A(u2__abc_52155_new_n8523_), .B(u2__abc_52155_new_n3481_), .Y(u2__abc_52155_new_n8526_));
OR2X2 OR2X2_1313 ( .A(u2__abc_52155_new_n8529_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8530_));
OR2X2 OR2X2_1314 ( .A(u2__abc_52155_new_n8528_), .B(u2__abc_52155_new_n8530_), .Y(u2__abc_52155_new_n8531_));
OR2X2 OR2X2_1315 ( .A(u2__abc_52155_new_n8535_), .B(u2__abc_52155_new_n8519_), .Y(u2__abc_52155_new_n8536_));
OR2X2 OR2X2_1316 ( .A(u2__abc_52155_new_n8540_), .B(u2__abc_52155_new_n8539_), .Y(u2__abc_52155_new_n8541_));
OR2X2 OR2X2_1317 ( .A(u2__abc_52155_new_n8542_), .B(u2__abc_52155_new_n3488_), .Y(u2__abc_52155_new_n8543_));
OR2X2 OR2X2_1318 ( .A(u2__abc_52155_new_n8546_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8547_));
OR2X2 OR2X2_1319 ( .A(u2__abc_52155_new_n8545_), .B(u2__abc_52155_new_n8547_), .Y(u2__abc_52155_new_n8548_));
OR2X2 OR2X2_132 ( .A(_abc_73687_new_n753_), .B(\a[65] ), .Y(_abc_73687_new_n1026_));
OR2X2 OR2X2_1320 ( .A(u2__abc_52155_new_n8552_), .B(u2__abc_52155_new_n8538_), .Y(u2__abc_52155_new_n8553_));
OR2X2 OR2X2_1321 ( .A(u2__abc_52155_new_n8520_), .B(u2__abc_52155_new_n3494_), .Y(u2__abc_52155_new_n8559_));
OR2X2 OR2X2_1322 ( .A(u2__abc_52155_new_n8562_), .B(u2__abc_52155_new_n3483_), .Y(u2__abc_52155_new_n8563_));
OR2X2 OR2X2_1323 ( .A(u2__abc_52155_new_n8561_), .B(u2__abc_52155_new_n8563_), .Y(u2__abc_52155_new_n8564_));
OR2X2 OR2X2_1324 ( .A(u2__abc_52155_new_n8558_), .B(u2__abc_52155_new_n8564_), .Y(u2__abc_52155_new_n8565_));
OR2X2 OR2X2_1325 ( .A(u2__abc_52155_new_n8557_), .B(u2__abc_52155_new_n8565_), .Y(u2__abc_52155_new_n8566_));
OR2X2 OR2X2_1326 ( .A(u2__abc_52155_new_n8556_), .B(u2__abc_52155_new_n8566_), .Y(u2__abc_52155_new_n8567_));
OR2X2 OR2X2_1327 ( .A(u2__abc_52155_new_n8567_), .B(u2__abc_52155_new_n3411_), .Y(u2__abc_52155_new_n8568_));
OR2X2 OR2X2_1328 ( .A(u2__abc_52155_new_n8571_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n8572_));
OR2X2 OR2X2_1329 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_46_), .Y(u2__abc_52155_new_n8573_));
OR2X2 OR2X2_133 ( .A(aNan), .B(sqrto_142_), .Y(_abc_73687_new_n1028_));
OR2X2 OR2X2_1330 ( .A(u2__abc_52155_new_n8574_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8575_));
OR2X2 OR2X2_1331 ( .A(u2__abc_52155_new_n8579_), .B(u2__abc_52155_new_n8555_), .Y(u2__abc_52155_new_n8580_));
OR2X2 OR2X2_1332 ( .A(u2__abc_52155_new_n8584_), .B(u2__abc_52155_new_n3404_), .Y(u2__abc_52155_new_n8585_));
OR2X2 OR2X2_1333 ( .A(u2__abc_52155_new_n8583_), .B(u2__abc_52155_new_n8586_), .Y(u2__abc_52155_new_n8587_));
OR2X2 OR2X2_1334 ( .A(u2__abc_52155_new_n8590_), .B(u2__abc_52155_new_n2993_), .Y(u2__abc_52155_new_n8591_));
OR2X2 OR2X2_1335 ( .A(u2__abc_52155_new_n8589_), .B(u2__abc_52155_new_n8591_), .Y(u2__abc_52155_new_n8592_));
OR2X2 OR2X2_1336 ( .A(u2__abc_52155_new_n8596_), .B(u2__abc_52155_new_n8582_), .Y(u2__abc_52155_new_n8597_));
OR2X2 OR2X2_1337 ( .A(u2__abc_52155_new_n8603_), .B(u2__abc_52155_new_n3402_), .Y(u2__abc_52155_new_n8604_));
OR2X2 OR2X2_1338 ( .A(u2__abc_52155_new_n8605_), .B(u2__abc_52155_new_n8601_), .Y(u2__abc_52155_new_n8606_));
OR2X2 OR2X2_1339 ( .A(u2__abc_52155_new_n8610_), .B(u2__abc_52155_new_n8600_), .Y(u2__abc_52155_new_n8611_));
OR2X2 OR2X2_134 ( .A(_abc_73687_new_n753_), .B(\a[66] ), .Y(_abc_73687_new_n1029_));
OR2X2 OR2X2_1340 ( .A(u2__abc_52155_new_n8611_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8612_));
OR2X2 OR2X2_1341 ( .A(u2__abc_52155_new_n8616_), .B(u2__abc_52155_new_n8599_), .Y(u2__abc_52155_new_n8617_));
OR2X2 OR2X2_1342 ( .A(u2__abc_52155_new_n8621_), .B(u2__abc_52155_new_n3395_), .Y(u2__abc_52155_new_n8622_));
OR2X2 OR2X2_1343 ( .A(u2__abc_52155_new_n8624_), .B(u2__abc_52155_new_n8623_), .Y(u2__abc_52155_new_n8625_));
OR2X2 OR2X2_1344 ( .A(u2__abc_52155_new_n8628_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8629_));
OR2X2 OR2X2_1345 ( .A(u2__abc_52155_new_n8627_), .B(u2__abc_52155_new_n8629_), .Y(u2__abc_52155_new_n8630_));
OR2X2 OR2X2_1346 ( .A(u2__abc_52155_new_n8634_), .B(u2__abc_52155_new_n8619_), .Y(u2__abc_52155_new_n8635_));
OR2X2 OR2X2_1347 ( .A(u2__abc_52155_new_n8602_), .B(u2__abc_52155_new_n3402_), .Y(u2__abc_52155_new_n8639_));
OR2X2 OR2X2_1348 ( .A(u2__abc_52155_new_n8639_), .B(u2__abc_52155_new_n3396_), .Y(u2__abc_52155_new_n8640_));
OR2X2 OR2X2_1349 ( .A(u2__abc_52155_new_n8620_), .B(u2__abc_52155_new_n3394_), .Y(u2__abc_52155_new_n8641_));
OR2X2 OR2X2_135 ( .A(aNan), .B(sqrto_143_), .Y(_abc_73687_new_n1031_));
OR2X2 OR2X2_1350 ( .A(u2__abc_52155_new_n8645_), .B(u2__abc_52155_new_n8644_), .Y(u2__abc_52155_new_n8646_));
OR2X2 OR2X2_1351 ( .A(u2__abc_52155_new_n8646_), .B(u2__abc_52155_new_n3442_), .Y(u2__abc_52155_new_n8647_));
OR2X2 OR2X2_1352 ( .A(u2__abc_52155_new_n8651_), .B(u2__abc_52155_new_n8638_), .Y(u2__abc_52155_new_n8652_));
OR2X2 OR2X2_1353 ( .A(u2__abc_52155_new_n8652_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8653_));
OR2X2 OR2X2_1354 ( .A(u2__abc_52155_new_n8657_), .B(u2__abc_52155_new_n8637_), .Y(u2__abc_52155_new_n8658_));
OR2X2 OR2X2_1355 ( .A(u2__abc_52155_new_n8665_), .B(u2__abc_52155_new_n8662_), .Y(u2__abc_52155_new_n8666_));
OR2X2 OR2X2_1356 ( .A(u2__abc_52155_new_n8668_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8669_));
OR2X2 OR2X2_1357 ( .A(u2__abc_52155_new_n8667_), .B(u2__abc_52155_new_n8669_), .Y(u2__abc_52155_new_n8670_));
OR2X2 OR2X2_1358 ( .A(u2__abc_52155_new_n8674_), .B(u2__abc_52155_new_n8660_), .Y(u2__abc_52155_new_n8675_));
OR2X2 OR2X2_1359 ( .A(u2__abc_52155_new_n8679_), .B(u2__abc_52155_new_n3433_), .Y(u2__abc_52155_new_n8680_));
OR2X2 OR2X2_136 ( .A(_abc_73687_new_n753_), .B(\a[67] ), .Y(_abc_73687_new_n1032_));
OR2X2 OR2X2_1360 ( .A(u2__abc_52155_new_n8681_), .B(u2__abc_52155_new_n3420_), .Y(u2__abc_52155_new_n8684_));
OR2X2 OR2X2_1361 ( .A(u2__abc_52155_new_n8687_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8688_));
OR2X2 OR2X2_1362 ( .A(u2__abc_52155_new_n8686_), .B(u2__abc_52155_new_n8688_), .Y(u2__abc_52155_new_n8689_));
OR2X2 OR2X2_1363 ( .A(u2__abc_52155_new_n8693_), .B(u2__abc_52155_new_n8677_), .Y(u2__abc_52155_new_n8694_));
OR2X2 OR2X2_1364 ( .A(u2__abc_52155_new_n8698_), .B(u2__abc_52155_new_n8697_), .Y(u2__abc_52155_new_n8699_));
OR2X2 OR2X2_1365 ( .A(u2__abc_52155_new_n8700_), .B(u2__abc_52155_new_n3427_), .Y(u2__abc_52155_new_n8701_));
OR2X2 OR2X2_1366 ( .A(u2__abc_52155_new_n8704_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8705_));
OR2X2 OR2X2_1367 ( .A(u2__abc_52155_new_n8703_), .B(u2__abc_52155_new_n8705_), .Y(u2__abc_52155_new_n8706_));
OR2X2 OR2X2_1368 ( .A(u2__abc_52155_new_n8710_), .B(u2__abc_52155_new_n8696_), .Y(u2__abc_52155_new_n8711_));
OR2X2 OR2X2_1369 ( .A(u2__abc_52155_new_n8678_), .B(u2__abc_52155_new_n3433_), .Y(u2__abc_52155_new_n8716_));
OR2X2 OR2X2_137 ( .A(aNan), .B(sqrto_144_), .Y(_abc_73687_new_n1034_));
OR2X2 OR2X2_1370 ( .A(u2__abc_52155_new_n8719_), .B(u2__abc_52155_new_n3422_), .Y(u2__abc_52155_new_n8720_));
OR2X2 OR2X2_1371 ( .A(u2__abc_52155_new_n8718_), .B(u2__abc_52155_new_n8720_), .Y(u2__abc_52155_new_n8721_));
OR2X2 OR2X2_1372 ( .A(u2__abc_52155_new_n8715_), .B(u2__abc_52155_new_n8721_), .Y(u2__abc_52155_new_n8722_));
OR2X2 OR2X2_1373 ( .A(u2__abc_52155_new_n8723_), .B(u2__abc_52155_new_n8722_), .Y(u2__abc_52155_new_n8724_));
OR2X2 OR2X2_1374 ( .A(u2__abc_52155_new_n8724_), .B(u2__abc_52155_new_n3344_), .Y(u2__abc_52155_new_n8725_));
OR2X2 OR2X2_1375 ( .A(u2__abc_52155_new_n8729_), .B(u2__abc_52155_new_n8714_), .Y(u2__abc_52155_new_n8730_));
OR2X2 OR2X2_1376 ( .A(u2__abc_52155_new_n8730_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8731_));
OR2X2 OR2X2_1377 ( .A(u2__abc_52155_new_n8735_), .B(u2__abc_52155_new_n8713_), .Y(u2__abc_52155_new_n8736_));
OR2X2 OR2X2_1378 ( .A(u2__abc_52155_new_n8739_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8740_));
OR2X2 OR2X2_1379 ( .A(u2__abc_52155_new_n8742_), .B(u2__abc_52155_new_n8741_), .Y(u2__abc_52155_new_n8743_));
OR2X2 OR2X2_138 ( .A(_abc_73687_new_n753_), .B(\a[68] ), .Y(_abc_73687_new_n1035_));
OR2X2 OR2X2_1380 ( .A(u2__abc_52155_new_n8744_), .B(u2__abc_52155_new_n3351_), .Y(u2__abc_52155_new_n8745_));
OR2X2 OR2X2_1381 ( .A(u2__abc_52155_new_n8747_), .B(u2__abc_52155_new_n8740_), .Y(u2__abc_52155_new_n8748_));
OR2X2 OR2X2_1382 ( .A(u2__abc_52155_new_n8752_), .B(u2__abc_52155_new_n8738_), .Y(u2__abc_52155_new_n8753_));
OR2X2 OR2X2_1383 ( .A(u2__abc_52155_new_n8756_), .B(u2__abc_52155_new_n3349_), .Y(u2__abc_52155_new_n8757_));
OR2X2 OR2X2_1384 ( .A(u2__abc_52155_new_n8759_), .B(u2__abc_52155_new_n8758_), .Y(u2__abc_52155_new_n8760_));
OR2X2 OR2X2_1385 ( .A(u2__abc_52155_new_n8760_), .B(u2__abc_52155_new_n3329_), .Y(u2__abc_52155_new_n8763_));
OR2X2 OR2X2_1386 ( .A(u2__abc_52155_new_n8766_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8767_));
OR2X2 OR2X2_1387 ( .A(u2__abc_52155_new_n8765_), .B(u2__abc_52155_new_n8767_), .Y(u2__abc_52155_new_n8768_));
OR2X2 OR2X2_1388 ( .A(u2__abc_52155_new_n8772_), .B(u2__abc_52155_new_n8755_), .Y(u2__abc_52155_new_n8773_));
OR2X2 OR2X2_1389 ( .A(u2__abc_52155_new_n8777_), .B(u2__abc_52155_new_n8776_), .Y(u2__abc_52155_new_n8778_));
OR2X2 OR2X2_139 ( .A(aNan), .B(sqrto_145_), .Y(_abc_73687_new_n1037_));
OR2X2 OR2X2_1390 ( .A(u2__abc_52155_new_n8779_), .B(u2__abc_52155_new_n3336_), .Y(u2__abc_52155_new_n8780_));
OR2X2 OR2X2_1391 ( .A(u2__abc_52155_new_n8783_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8784_));
OR2X2 OR2X2_1392 ( .A(u2__abc_52155_new_n8782_), .B(u2__abc_52155_new_n8784_), .Y(u2__abc_52155_new_n8785_));
OR2X2 OR2X2_1393 ( .A(u2__abc_52155_new_n8789_), .B(u2__abc_52155_new_n8775_), .Y(u2__abc_52155_new_n8790_));
OR2X2 OR2X2_1394 ( .A(u2__abc_52155_new_n8794_), .B(u2__abc_52155_new_n3331_), .Y(u2__abc_52155_new_n8795_));
OR2X2 OR2X2_1395 ( .A(u2__abc_52155_new_n8793_), .B(u2__abc_52155_new_n8795_), .Y(u2__abc_52155_new_n8796_));
OR2X2 OR2X2_1396 ( .A(u2__abc_52155_new_n8797_), .B(u2__abc_52155_new_n8796_), .Y(u2__abc_52155_new_n8798_));
OR2X2 OR2X2_1397 ( .A(u2__abc_52155_new_n8798_), .B(u2__abc_52155_new_n3382_), .Y(u2__abc_52155_new_n8801_));
OR2X2 OR2X2_1398 ( .A(u2__abc_52155_new_n8804_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8805_));
OR2X2 OR2X2_1399 ( .A(u2__abc_52155_new_n8803_), .B(u2__abc_52155_new_n8805_), .Y(u2__abc_52155_new_n8806_));
OR2X2 OR2X2_14 ( .A(_abc_73687_new_n753_), .B(\a[6] ), .Y(_abc_73687_new_n849_));
OR2X2 OR2X2_140 ( .A(_abc_73687_new_n753_), .B(\a[69] ), .Y(_abc_73687_new_n1038_));
OR2X2 OR2X2_1400 ( .A(u2__abc_52155_new_n8810_), .B(u2__abc_52155_new_n8792_), .Y(u2__abc_52155_new_n8811_));
OR2X2 OR2X2_1401 ( .A(u2__abc_52155_new_n8815_), .B(u2__abc_52155_new_n3375_), .Y(u2__abc_52155_new_n8816_));
OR2X2 OR2X2_1402 ( .A(u2__abc_52155_new_n8821_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8822_));
OR2X2 OR2X2_1403 ( .A(u2__abc_52155_new_n8820_), .B(u2__abc_52155_new_n8822_), .Y(u2__abc_52155_new_n8823_));
OR2X2 OR2X2_1404 ( .A(u2__abc_52155_new_n8827_), .B(u2__abc_52155_new_n8813_), .Y(u2__abc_52155_new_n8828_));
OR2X2 OR2X2_1405 ( .A(u2__abc_52155_new_n8832_), .B(u2__abc_52155_new_n3360_), .Y(u2__abc_52155_new_n8835_));
OR2X2 OR2X2_1406 ( .A(u2__abc_52155_new_n8838_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8839_));
OR2X2 OR2X2_1407 ( .A(u2__abc_52155_new_n8837_), .B(u2__abc_52155_new_n8839_), .Y(u2__abc_52155_new_n8840_));
OR2X2 OR2X2_1408 ( .A(u2__abc_52155_new_n8845_), .B(u2__abc_52155_new_n8830_), .Y(u2__abc_52155_new_n8846_));
OR2X2 OR2X2_1409 ( .A(u2__abc_52155_new_n8850_), .B(u2__abc_52155_new_n8849_), .Y(u2__abc_52155_new_n8851_));
OR2X2 OR2X2_141 ( .A(aNan), .B(sqrto_146_), .Y(_abc_73687_new_n1040_));
OR2X2 OR2X2_1410 ( .A(u2__abc_52155_new_n8852_), .B(u2__abc_52155_new_n3367_), .Y(u2__abc_52155_new_n8853_));
OR2X2 OR2X2_1411 ( .A(u2__abc_52155_new_n8856_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8857_));
OR2X2 OR2X2_1412 ( .A(u2__abc_52155_new_n8855_), .B(u2__abc_52155_new_n8857_), .Y(u2__abc_52155_new_n8858_));
OR2X2 OR2X2_1413 ( .A(u2__abc_52155_new_n8862_), .B(u2__abc_52155_new_n8848_), .Y(u2__abc_52155_new_n8863_));
OR2X2 OR2X2_1414 ( .A(u2__abc_52155_new_n3370_), .B(u2__abc_52155_new_n3377_), .Y(u2__abc_52155_new_n8869_));
OR2X2 OR2X2_1415 ( .A(u2__abc_52155_new_n8872_), .B(u2__abc_52155_new_n3365_), .Y(u2__abc_52155_new_n8873_));
OR2X2 OR2X2_1416 ( .A(u2__abc_52155_new_n8871_), .B(u2__abc_52155_new_n8873_), .Y(u2__abc_52155_new_n8874_));
OR2X2 OR2X2_1417 ( .A(u2__abc_52155_new_n8868_), .B(u2__abc_52155_new_n8874_), .Y(u2__abc_52155_new_n8875_));
OR2X2 OR2X2_1418 ( .A(u2__abc_52155_new_n8867_), .B(u2__abc_52155_new_n8875_), .Y(u2__abc_52155_new_n8876_));
OR2X2 OR2X2_1419 ( .A(u2__abc_52155_new_n8877_), .B(u2__abc_52155_new_n8876_), .Y(u2__abc_52155_new_n8878_));
OR2X2 OR2X2_142 ( .A(_abc_73687_new_n753_), .B(\a[70] ), .Y(_abc_73687_new_n1041_));
OR2X2 OR2X2_1420 ( .A(u2__abc_52155_new_n8878_), .B(u2__abc_52155_new_n4083_), .Y(u2__abc_52155_new_n8879_));
OR2X2 OR2X2_1421 ( .A(u2__abc_52155_new_n8883_), .B(u2__abc_52155_new_n8866_), .Y(u2__abc_52155_new_n8884_));
OR2X2 OR2X2_1422 ( .A(u2__abc_52155_new_n8884_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8885_));
OR2X2 OR2X2_1423 ( .A(u2__abc_52155_new_n8889_), .B(u2__abc_52155_new_n8865_), .Y(u2__abc_52155_new_n8890_));
OR2X2 OR2X2_1424 ( .A(u2__abc_52155_new_n8894_), .B(u2__abc_52155_new_n4090_), .Y(u2__abc_52155_new_n8895_));
OR2X2 OR2X2_1425 ( .A(u2__abc_52155_new_n8893_), .B(u2__abc_52155_new_n8896_), .Y(u2__abc_52155_new_n8897_));
OR2X2 OR2X2_1426 ( .A(u2__abc_52155_new_n8900_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8901_));
OR2X2 OR2X2_1427 ( .A(u2__abc_52155_new_n8899_), .B(u2__abc_52155_new_n8901_), .Y(u2__abc_52155_new_n8902_));
OR2X2 OR2X2_1428 ( .A(u2__abc_52155_new_n8906_), .B(u2__abc_52155_new_n8892_), .Y(u2__abc_52155_new_n8907_));
OR2X2 OR2X2_1429 ( .A(u2__abc_52155_new_n4081_), .B(u2__abc_52155_new_n4088_), .Y(u2__abc_52155_new_n8911_));
OR2X2 OR2X2_143 ( .A(aNan), .B(sqrto_147_), .Y(_abc_73687_new_n1043_));
OR2X2 OR2X2_1430 ( .A(u2__abc_52155_new_n8914_), .B(u2__abc_52155_new_n8913_), .Y(u2__abc_52155_new_n8915_));
OR2X2 OR2X2_1431 ( .A(u2__abc_52155_new_n8915_), .B(u2__abc_52155_new_n8910_), .Y(u2__abc_52155_new_n8916_));
OR2X2 OR2X2_1432 ( .A(u2__abc_52155_new_n8919_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n8920_));
OR2X2 OR2X2_1433 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_64_), .Y(u2__abc_52155_new_n8921_));
OR2X2 OR2X2_1434 ( .A(u2__abc_52155_new_n8922_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8923_));
OR2X2 OR2X2_1435 ( .A(u2__abc_52155_new_n8927_), .B(u2__abc_52155_new_n8909_), .Y(u2__abc_52155_new_n8928_));
OR2X2 OR2X2_1436 ( .A(u2__abc_52155_new_n8932_), .B(u2__abc_52155_new_n4101_), .Y(u2__abc_52155_new_n8933_));
OR2X2 OR2X2_1437 ( .A(u2__abc_52155_new_n8935_), .B(u2__abc_52155_new_n8934_), .Y(u2__abc_52155_new_n8936_));
OR2X2 OR2X2_1438 ( .A(u2__abc_52155_new_n8939_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8940_));
OR2X2 OR2X2_1439 ( .A(u2__abc_52155_new_n8938_), .B(u2__abc_52155_new_n8940_), .Y(u2__abc_52155_new_n8941_));
OR2X2 OR2X2_144 ( .A(_abc_73687_new_n753_), .B(\a[71] ), .Y(_abc_73687_new_n1044_));
OR2X2 OR2X2_1440 ( .A(u2__abc_52155_new_n8945_), .B(u2__abc_52155_new_n8930_), .Y(u2__abc_52155_new_n8946_));
OR2X2 OR2X2_1441 ( .A(u2__abc_52155_new_n8951_), .B(u2__abc_52155_new_n4098_), .Y(u2__abc_52155_new_n8952_));
OR2X2 OR2X2_1442 ( .A(u2__abc_52155_new_n8950_), .B(u2__abc_52155_new_n8952_), .Y(u2__abc_52155_new_n8953_));
OR2X2 OR2X2_1443 ( .A(u2__abc_52155_new_n8954_), .B(u2__abc_52155_new_n8953_), .Y(u2__abc_52155_new_n8955_));
OR2X2 OR2X2_1444 ( .A(u2__abc_52155_new_n8955_), .B(u2__abc_52155_new_n8949_), .Y(u2__abc_52155_new_n8956_));
OR2X2 OR2X2_1445 ( .A(u2__abc_52155_new_n8959_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n8960_));
OR2X2 OR2X2_1446 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_66_), .Y(u2__abc_52155_new_n8961_));
OR2X2 OR2X2_1447 ( .A(u2__abc_52155_new_n8962_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8963_));
OR2X2 OR2X2_1448 ( .A(u2__abc_52155_new_n8967_), .B(u2__abc_52155_new_n8948_), .Y(u2__abc_52155_new_n8968_));
OR2X2 OR2X2_1449 ( .A(u2__abc_52155_new_n8974_), .B(u2__abc_52155_new_n8971_), .Y(u2__abc_52155_new_n8977_));
OR2X2 OR2X2_145 ( .A(aNan), .B(sqrto_148_), .Y(_abc_73687_new_n1046_));
OR2X2 OR2X2_1450 ( .A(u2__abc_52155_new_n8980_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8981_));
OR2X2 OR2X2_1451 ( .A(u2__abc_52155_new_n8979_), .B(u2__abc_52155_new_n8981_), .Y(u2__abc_52155_new_n8982_));
OR2X2 OR2X2_1452 ( .A(u2__abc_52155_new_n8986_), .B(u2__abc_52155_new_n8970_), .Y(u2__abc_52155_new_n8987_));
OR2X2 OR2X2_1453 ( .A(u2__abc_52155_new_n8975_), .B(u2__abc_52155_new_n4117_), .Y(u2__abc_52155_new_n8991_));
OR2X2 OR2X2_1454 ( .A(u2__abc_52155_new_n8991_), .B(u2__abc_52155_new_n8990_), .Y(u2__abc_52155_new_n8994_));
OR2X2 OR2X2_1455 ( .A(u2__abc_52155_new_n8997_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n8998_));
OR2X2 OR2X2_1456 ( .A(u2__abc_52155_new_n8996_), .B(u2__abc_52155_new_n8998_), .Y(u2__abc_52155_new_n8999_));
OR2X2 OR2X2_1457 ( .A(u2__abc_52155_new_n9003_), .B(u2__abc_52155_new_n8989_), .Y(u2__abc_52155_new_n9004_));
OR2X2 OR2X2_1458 ( .A(u2__abc_52155_new_n9008_), .B(u2__abc_52155_new_n4114_), .Y(u2__abc_52155_new_n9009_));
OR2X2 OR2X2_1459 ( .A(u2__abc_52155_new_n9011_), .B(u2__abc_52155_new_n9010_), .Y(u2__abc_52155_new_n9012_));
OR2X2 OR2X2_146 ( .A(_abc_73687_new_n753_), .B(\a[72] ), .Y(_abc_73687_new_n1047_));
OR2X2 OR2X2_1460 ( .A(u2__abc_52155_new_n9015_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9016_));
OR2X2 OR2X2_1461 ( .A(u2__abc_52155_new_n9014_), .B(u2__abc_52155_new_n9016_), .Y(u2__abc_52155_new_n9017_));
OR2X2 OR2X2_1462 ( .A(u2__abc_52155_new_n9021_), .B(u2__abc_52155_new_n9006_), .Y(u2__abc_52155_new_n9022_));
OR2X2 OR2X2_1463 ( .A(u2__abc_52155_new_n4117_), .B(u2__abc_52155_new_n4122_), .Y(u2__abc_52155_new_n9028_));
OR2X2 OR2X2_1464 ( .A(u2__abc_52155_new_n9007_), .B(u2__abc_52155_new_n4113_), .Y(u2__abc_52155_new_n9032_));
OR2X2 OR2X2_1465 ( .A(u2__abc_52155_new_n9037_), .B(u2__abc_52155_new_n9036_), .Y(u2__abc_52155_new_n9038_));
OR2X2 OR2X2_1466 ( .A(u2__abc_52155_new_n9038_), .B(u2__abc_52155_new_n4025_), .Y(u2__abc_52155_new_n9039_));
OR2X2 OR2X2_1467 ( .A(u2__abc_52155_new_n9042_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n9043_));
OR2X2 OR2X2_1468 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_70_), .Y(u2__abc_52155_new_n9044_));
OR2X2 OR2X2_1469 ( .A(u2__abc_52155_new_n9045_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9046_));
OR2X2 OR2X2_147 ( .A(aNan), .B(sqrto_149_), .Y(_abc_73687_new_n1049_));
OR2X2 OR2X2_1470 ( .A(u2__abc_52155_new_n9050_), .B(u2__abc_52155_new_n9024_), .Y(u2__abc_52155_new_n9051_));
OR2X2 OR2X2_1471 ( .A(u2__abc_52155_new_n9055_), .B(u2__abc_52155_new_n9054_), .Y(u2__abc_52155_new_n9056_));
OR2X2 OR2X2_1472 ( .A(u2__abc_52155_new_n9057_), .B(u2__abc_52155_new_n4032_), .Y(u2__abc_52155_new_n9058_));
OR2X2 OR2X2_1473 ( .A(u2__abc_52155_new_n9061_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9062_));
OR2X2 OR2X2_1474 ( .A(u2__abc_52155_new_n9060_), .B(u2__abc_52155_new_n9062_), .Y(u2__abc_52155_new_n9063_));
OR2X2 OR2X2_1475 ( .A(u2__abc_52155_new_n9067_), .B(u2__abc_52155_new_n9053_), .Y(u2__abc_52155_new_n9068_));
OR2X2 OR2X2_1476 ( .A(u2__abc_52155_new_n4021_), .B(u2__abc_52155_new_n4030_), .Y(u2__abc_52155_new_n9072_));
OR2X2 OR2X2_1477 ( .A(u2__abc_52155_new_n9075_), .B(u2__abc_52155_new_n9074_), .Y(u2__abc_52155_new_n9076_));
OR2X2 OR2X2_1478 ( .A(u2__abc_52155_new_n9076_), .B(u2__abc_52155_new_n9071_), .Y(u2__abc_52155_new_n9079_));
OR2X2 OR2X2_1479 ( .A(u2__abc_52155_new_n9082_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9083_));
OR2X2 OR2X2_148 ( .A(_abc_73687_new_n753_), .B(\a[73] ), .Y(_abc_73687_new_n1050_));
OR2X2 OR2X2_1480 ( .A(u2__abc_52155_new_n9081_), .B(u2__abc_52155_new_n9083_), .Y(u2__abc_52155_new_n9084_));
OR2X2 OR2X2_1481 ( .A(u2__abc_52155_new_n9088_), .B(u2__abc_52155_new_n9070_), .Y(u2__abc_52155_new_n9089_));
OR2X2 OR2X2_1482 ( .A(u2__abc_52155_new_n9093_), .B(u2__abc_52155_new_n4043_), .Y(u2__abc_52155_new_n9094_));
OR2X2 OR2X2_1483 ( .A(u2__abc_52155_new_n9096_), .B(u2__abc_52155_new_n9095_), .Y(u2__abc_52155_new_n9097_));
OR2X2 OR2X2_1484 ( .A(u2__abc_52155_new_n9100_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9101_));
OR2X2 OR2X2_1485 ( .A(u2__abc_52155_new_n9099_), .B(u2__abc_52155_new_n9101_), .Y(u2__abc_52155_new_n9102_));
OR2X2 OR2X2_1486 ( .A(u2__abc_52155_new_n9106_), .B(u2__abc_52155_new_n9091_), .Y(u2__abc_52155_new_n9107_));
OR2X2 OR2X2_1487 ( .A(u2__abc_52155_new_n9092_), .B(u2__abc_52155_new_n4042_), .Y(u2__abc_52155_new_n9112_));
OR2X2 OR2X2_1488 ( .A(u2__abc_52155_new_n9116_), .B(u2__abc_52155_new_n9115_), .Y(u2__abc_52155_new_n9117_));
OR2X2 OR2X2_1489 ( .A(u2__abc_52155_new_n9117_), .B(u2__abc_52155_new_n4075_), .Y(u2__abc_52155_new_n9120_));
OR2X2 OR2X2_149 ( .A(aNan), .B(sqrto_150_), .Y(_abc_73687_new_n1052_));
OR2X2 OR2X2_1490 ( .A(u2__abc_52155_new_n9123_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9124_));
OR2X2 OR2X2_1491 ( .A(u2__abc_52155_new_n9122_), .B(u2__abc_52155_new_n9124_), .Y(u2__abc_52155_new_n9125_));
OR2X2 OR2X2_1492 ( .A(u2__abc_52155_new_n9129_), .B(u2__abc_52155_new_n9109_), .Y(u2__abc_52155_new_n9130_));
OR2X2 OR2X2_1493 ( .A(u2__abc_52155_new_n9134_), .B(u2__abc_52155_new_n4068_), .Y(u2__abc_52155_new_n9137_));
OR2X2 OR2X2_1494 ( .A(u2__abc_52155_new_n9140_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9141_));
OR2X2 OR2X2_1495 ( .A(u2__abc_52155_new_n9139_), .B(u2__abc_52155_new_n9141_), .Y(u2__abc_52155_new_n9142_));
OR2X2 OR2X2_1496 ( .A(u2__abc_52155_new_n9146_), .B(u2__abc_52155_new_n9132_), .Y(u2__abc_52155_new_n9147_));
OR2X2 OR2X2_1497 ( .A(u2__abc_52155_new_n9151_), .B(u2__abc_52155_new_n4053_), .Y(u2__abc_52155_new_n9154_));
OR2X2 OR2X2_1498 ( .A(u2__abc_52155_new_n9157_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9158_));
OR2X2 OR2X2_1499 ( .A(u2__abc_52155_new_n9156_), .B(u2__abc_52155_new_n9158_), .Y(u2__abc_52155_new_n9159_));
OR2X2 OR2X2_15 ( .A(aNan), .B(sqrto_83_), .Y(_abc_73687_new_n851_));
OR2X2 OR2X2_150 ( .A(_abc_73687_new_n753_), .B(\a[74] ), .Y(_abc_73687_new_n1053_));
OR2X2 OR2X2_1500 ( .A(u2__abc_52155_new_n9163_), .B(u2__abc_52155_new_n9149_), .Y(u2__abc_52155_new_n9164_));
OR2X2 OR2X2_1501 ( .A(u2__abc_52155_new_n9168_), .B(u2__abc_52155_new_n9167_), .Y(u2__abc_52155_new_n9169_));
OR2X2 OR2X2_1502 ( .A(u2__abc_52155_new_n9170_), .B(u2__abc_52155_new_n4060_), .Y(u2__abc_52155_new_n9171_));
OR2X2 OR2X2_1503 ( .A(u2__abc_52155_new_n9174_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9175_));
OR2X2 OR2X2_1504 ( .A(u2__abc_52155_new_n9173_), .B(u2__abc_52155_new_n9175_), .Y(u2__abc_52155_new_n9176_));
OR2X2 OR2X2_1505 ( .A(u2__abc_52155_new_n9180_), .B(u2__abc_52155_new_n9166_), .Y(u2__abc_52155_new_n9181_));
OR2X2 OR2X2_1506 ( .A(u2__abc_52155_new_n9186_), .B(u2__abc_52155_new_n4055_), .Y(u2__abc_52155_new_n9187_));
OR2X2 OR2X2_1507 ( .A(u2__abc_52155_new_n4063_), .B(u2__abc_52155_new_n4070_), .Y(u2__abc_52155_new_n9188_));
OR2X2 OR2X2_1508 ( .A(u2__abc_52155_new_n9190_), .B(u2__abc_52155_new_n9187_), .Y(u2__abc_52155_new_n9191_));
OR2X2 OR2X2_1509 ( .A(u2__abc_52155_new_n9185_), .B(u2__abc_52155_new_n9191_), .Y(u2__abc_52155_new_n9192_));
OR2X2 OR2X2_151 ( .A(aNan), .B(sqrto_151_), .Y(_abc_73687_new_n1055_));
OR2X2 OR2X2_1510 ( .A(u2__abc_52155_new_n9184_), .B(u2__abc_52155_new_n9192_), .Y(u2__abc_52155_new_n9193_));
OR2X2 OR2X2_1511 ( .A(u2__abc_52155_new_n9194_), .B(u2__abc_52155_new_n9193_), .Y(u2__abc_52155_new_n9195_));
OR2X2 OR2X2_1512 ( .A(u2__abc_52155_new_n9195_), .B(u2__abc_52155_new_n3964_), .Y(u2__abc_52155_new_n9196_));
OR2X2 OR2X2_1513 ( .A(u2__abc_52155_new_n9199_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n9200_));
OR2X2 OR2X2_1514 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_78_), .Y(u2__abc_52155_new_n9201_));
OR2X2 OR2X2_1515 ( .A(u2__abc_52155_new_n9202_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9203_));
OR2X2 OR2X2_1516 ( .A(u2__abc_52155_new_n9207_), .B(u2__abc_52155_new_n9183_), .Y(u2__abc_52155_new_n9208_));
OR2X2 OR2X2_1517 ( .A(u2__abc_52155_new_n9212_), .B(u2__abc_52155_new_n9211_), .Y(u2__abc_52155_new_n9213_));
OR2X2 OR2X2_1518 ( .A(u2__abc_52155_new_n9214_), .B(u2__abc_52155_new_n3971_), .Y(u2__abc_52155_new_n9215_));
OR2X2 OR2X2_1519 ( .A(u2__abc_52155_new_n9218_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9219_));
OR2X2 OR2X2_152 ( .A(_abc_73687_new_n753_), .B(\a[75] ), .Y(_abc_73687_new_n1056_));
OR2X2 OR2X2_1520 ( .A(u2__abc_52155_new_n9217_), .B(u2__abc_52155_new_n9219_), .Y(u2__abc_52155_new_n9220_));
OR2X2 OR2X2_1521 ( .A(u2__abc_52155_new_n9224_), .B(u2__abc_52155_new_n9210_), .Y(u2__abc_52155_new_n9225_));
OR2X2 OR2X2_1522 ( .A(u2__abc_52155_new_n3960_), .B(u2__abc_52155_new_n3969_), .Y(u2__abc_52155_new_n9229_));
OR2X2 OR2X2_1523 ( .A(u2__abc_52155_new_n9232_), .B(u2__abc_52155_new_n9231_), .Y(u2__abc_52155_new_n9233_));
OR2X2 OR2X2_1524 ( .A(u2__abc_52155_new_n9233_), .B(u2__abc_52155_new_n9228_), .Y(u2__abc_52155_new_n9236_));
OR2X2 OR2X2_1525 ( .A(u2__abc_52155_new_n9239_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9240_));
OR2X2 OR2X2_1526 ( .A(u2__abc_52155_new_n9238_), .B(u2__abc_52155_new_n9240_), .Y(u2__abc_52155_new_n9241_));
OR2X2 OR2X2_1527 ( .A(u2__abc_52155_new_n9245_), .B(u2__abc_52155_new_n9227_), .Y(u2__abc_52155_new_n9246_));
OR2X2 OR2X2_1528 ( .A(u2__abc_52155_new_n9250_), .B(u2__abc_52155_new_n3982_), .Y(u2__abc_52155_new_n9251_));
OR2X2 OR2X2_1529 ( .A(u2__abc_52155_new_n9253_), .B(u2__abc_52155_new_n9252_), .Y(u2__abc_52155_new_n9254_));
OR2X2 OR2X2_153 ( .A(aNan), .B(sqrto_152_), .Y(_abc_73687_new_n1058_));
OR2X2 OR2X2_1530 ( .A(u2__abc_52155_new_n9257_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9258_));
OR2X2 OR2X2_1531 ( .A(u2__abc_52155_new_n9256_), .B(u2__abc_52155_new_n9258_), .Y(u2__abc_52155_new_n9259_));
OR2X2 OR2X2_1532 ( .A(u2__abc_52155_new_n9263_), .B(u2__abc_52155_new_n9248_), .Y(u2__abc_52155_new_n9264_));
OR2X2 OR2X2_1533 ( .A(u2__abc_52155_new_n9249_), .B(u2__abc_52155_new_n3981_), .Y(u2__abc_52155_new_n9269_));
OR2X2 OR2X2_1534 ( .A(u2__abc_52155_new_n9273_), .B(u2__abc_52155_new_n9272_), .Y(u2__abc_52155_new_n9274_));
OR2X2 OR2X2_1535 ( .A(u2__abc_52155_new_n9274_), .B(u2__abc_52155_new_n4014_), .Y(u2__abc_52155_new_n9277_));
OR2X2 OR2X2_1536 ( .A(u2__abc_52155_new_n9280_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9281_));
OR2X2 OR2X2_1537 ( .A(u2__abc_52155_new_n9279_), .B(u2__abc_52155_new_n9281_), .Y(u2__abc_52155_new_n9282_));
OR2X2 OR2X2_1538 ( .A(u2__abc_52155_new_n9286_), .B(u2__abc_52155_new_n9266_), .Y(u2__abc_52155_new_n9287_));
OR2X2 OR2X2_1539 ( .A(u2__abc_52155_new_n9294_), .B(u2__abc_52155_new_n9291_), .Y(u2__abc_52155_new_n9295_));
OR2X2 OR2X2_154 ( .A(_abc_73687_new_n753_), .B(\a[76] ), .Y(_abc_73687_new_n1059_));
OR2X2 OR2X2_1540 ( .A(u2__abc_52155_new_n9297_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9298_));
OR2X2 OR2X2_1541 ( .A(u2__abc_52155_new_n9296_), .B(u2__abc_52155_new_n9298_), .Y(u2__abc_52155_new_n9299_));
OR2X2 OR2X2_1542 ( .A(u2__abc_52155_new_n9303_), .B(u2__abc_52155_new_n9289_), .Y(u2__abc_52155_new_n9304_));
OR2X2 OR2X2_1543 ( .A(u2__abc_52155_new_n9308_), .B(u2__abc_52155_new_n4005_), .Y(u2__abc_52155_new_n9309_));
OR2X2 OR2X2_1544 ( .A(u2__abc_52155_new_n9310_), .B(u2__abc_52155_new_n3992_), .Y(u2__abc_52155_new_n9313_));
OR2X2 OR2X2_1545 ( .A(u2__abc_52155_new_n9316_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9317_));
OR2X2 OR2X2_1546 ( .A(u2__abc_52155_new_n9315_), .B(u2__abc_52155_new_n9317_), .Y(u2__abc_52155_new_n9318_));
OR2X2 OR2X2_1547 ( .A(u2__abc_52155_new_n9322_), .B(u2__abc_52155_new_n9306_), .Y(u2__abc_52155_new_n9323_));
OR2X2 OR2X2_1548 ( .A(u2__abc_52155_new_n9327_), .B(u2__abc_52155_new_n9326_), .Y(u2__abc_52155_new_n9328_));
OR2X2 OR2X2_1549 ( .A(u2__abc_52155_new_n9329_), .B(u2__abc_52155_new_n3999_), .Y(u2__abc_52155_new_n9330_));
OR2X2 OR2X2_155 ( .A(aNan), .B(sqrto_153_), .Y(_abc_73687_new_n1061_));
OR2X2 OR2X2_1550 ( .A(u2__abc_52155_new_n9333_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9334_));
OR2X2 OR2X2_1551 ( .A(u2__abc_52155_new_n9332_), .B(u2__abc_52155_new_n9334_), .Y(u2__abc_52155_new_n9335_));
OR2X2 OR2X2_1552 ( .A(u2__abc_52155_new_n9339_), .B(u2__abc_52155_new_n9325_), .Y(u2__abc_52155_new_n9340_));
OR2X2 OR2X2_1553 ( .A(u2__abc_52155_new_n9345_), .B(u2__abc_52155_new_n3997_), .Y(u2__abc_52155_new_n9346_));
OR2X2 OR2X2_1554 ( .A(u2__abc_52155_new_n9307_), .B(u2__abc_52155_new_n4005_), .Y(u2__abc_52155_new_n9347_));
OR2X2 OR2X2_1555 ( .A(u2__abc_52155_new_n9354_), .B(u2__abc_52155_new_n9353_), .Y(u2__abc_52155_new_n9355_));
OR2X2 OR2X2_1556 ( .A(u2__abc_52155_new_n9355_), .B(u2__abc_52155_new_n3954_), .Y(u2__abc_52155_new_n9358_));
OR2X2 OR2X2_1557 ( .A(u2__abc_52155_new_n9361_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9362_));
OR2X2 OR2X2_1558 ( .A(u2__abc_52155_new_n9360_), .B(u2__abc_52155_new_n9362_), .Y(u2__abc_52155_new_n9363_));
OR2X2 OR2X2_1559 ( .A(u2__abc_52155_new_n9367_), .B(u2__abc_52155_new_n9342_), .Y(u2__abc_52155_new_n9368_));
OR2X2 OR2X2_156 ( .A(_abc_73687_new_n753_), .B(\a[77] ), .Y(_abc_73687_new_n1062_));
OR2X2 OR2X2_1560 ( .A(u2__abc_52155_new_n9372_), .B(u2__abc_52155_new_n3947_), .Y(u2__abc_52155_new_n9373_));
OR2X2 OR2X2_1561 ( .A(u2__abc_52155_new_n9371_), .B(u2__abc_52155_new_n9374_), .Y(u2__abc_52155_new_n9375_));
OR2X2 OR2X2_1562 ( .A(u2__abc_52155_new_n9378_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9379_));
OR2X2 OR2X2_1563 ( .A(u2__abc_52155_new_n9377_), .B(u2__abc_52155_new_n9379_), .Y(u2__abc_52155_new_n9380_));
OR2X2 OR2X2_1564 ( .A(u2__abc_52155_new_n9384_), .B(u2__abc_52155_new_n9370_), .Y(u2__abc_52155_new_n9385_));
OR2X2 OR2X2_1565 ( .A(u2__abc_52155_new_n9388_), .B(u2__abc_52155_new_n3945_), .Y(u2__abc_52155_new_n9389_));
OR2X2 OR2X2_1566 ( .A(u2__abc_52155_new_n9391_), .B(u2__abc_52155_new_n9390_), .Y(u2__abc_52155_new_n9392_));
OR2X2 OR2X2_1567 ( .A(u2__abc_52155_new_n9392_), .B(u2__abc_52155_new_n3932_), .Y(u2__abc_52155_new_n9395_));
OR2X2 OR2X2_1568 ( .A(u2__abc_52155_new_n9398_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9399_));
OR2X2 OR2X2_1569 ( .A(u2__abc_52155_new_n9397_), .B(u2__abc_52155_new_n9399_), .Y(u2__abc_52155_new_n9400_));
OR2X2 OR2X2_157 ( .A(aNan), .B(sqrto_154_), .Y(_abc_73687_new_n1064_));
OR2X2 OR2X2_1570 ( .A(u2__abc_52155_new_n9404_), .B(u2__abc_52155_new_n9387_), .Y(u2__abc_52155_new_n9405_));
OR2X2 OR2X2_1571 ( .A(u2__abc_52155_new_n9409_), .B(u2__abc_52155_new_n9408_), .Y(u2__abc_52155_new_n9410_));
OR2X2 OR2X2_1572 ( .A(u2__abc_52155_new_n9411_), .B(u2__abc_52155_new_n3939_), .Y(u2__abc_52155_new_n9412_));
OR2X2 OR2X2_1573 ( .A(u2__abc_52155_new_n9415_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9416_));
OR2X2 OR2X2_1574 ( .A(u2__abc_52155_new_n9414_), .B(u2__abc_52155_new_n9416_), .Y(u2__abc_52155_new_n9417_));
OR2X2 OR2X2_1575 ( .A(u2__abc_52155_new_n9421_), .B(u2__abc_52155_new_n9407_), .Y(u2__abc_52155_new_n9422_));
OR2X2 OR2X2_1576 ( .A(u2__abc_52155_new_n9426_), .B(u2__abc_52155_new_n3937_), .Y(u2__abc_52155_new_n9427_));
OR2X2 OR2X2_1577 ( .A(u2__abc_52155_new_n9428_), .B(u2__abc_52155_new_n3923_), .Y(u2__abc_52155_new_n9431_));
OR2X2 OR2X2_1578 ( .A(u2__abc_52155_new_n9434_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9435_));
OR2X2 OR2X2_1579 ( .A(u2__abc_52155_new_n9433_), .B(u2__abc_52155_new_n9435_), .Y(u2__abc_52155_new_n9436_));
OR2X2 OR2X2_158 ( .A(_abc_73687_new_n753_), .B(\a[78] ), .Y(_abc_73687_new_n1065_));
OR2X2 OR2X2_1580 ( .A(u2__abc_52155_new_n9440_), .B(u2__abc_52155_new_n9424_), .Y(u2__abc_52155_new_n9441_));
OR2X2 OR2X2_1581 ( .A(u2__abc_52155_new_n9448_), .B(u2__abc_52155_new_n9445_), .Y(u2__abc_52155_new_n9449_));
OR2X2 OR2X2_1582 ( .A(u2__abc_52155_new_n9451_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9452_));
OR2X2 OR2X2_1583 ( .A(u2__abc_52155_new_n9450_), .B(u2__abc_52155_new_n9452_), .Y(u2__abc_52155_new_n9453_));
OR2X2 OR2X2_1584 ( .A(u2__abc_52155_new_n9457_), .B(u2__abc_52155_new_n9443_), .Y(u2__abc_52155_new_n9458_));
OR2X2 OR2X2_1585 ( .A(u2__abc_52155_new_n9462_), .B(u2__abc_52155_new_n3914_), .Y(u2__abc_52155_new_n9463_));
OR2X2 OR2X2_1586 ( .A(u2__abc_52155_new_n9464_), .B(u2__abc_52155_new_n3901_), .Y(u2__abc_52155_new_n9467_));
OR2X2 OR2X2_1587 ( .A(u2__abc_52155_new_n9470_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9471_));
OR2X2 OR2X2_1588 ( .A(u2__abc_52155_new_n9469_), .B(u2__abc_52155_new_n9471_), .Y(u2__abc_52155_new_n9472_));
OR2X2 OR2X2_1589 ( .A(u2__abc_52155_new_n9476_), .B(u2__abc_52155_new_n9460_), .Y(u2__abc_52155_new_n9477_));
OR2X2 OR2X2_159 ( .A(aNan), .B(sqrto_155_), .Y(_abc_73687_new_n1067_));
OR2X2 OR2X2_1590 ( .A(u2__abc_52155_new_n9484_), .B(u2__abc_52155_new_n9481_), .Y(u2__abc_52155_new_n9485_));
OR2X2 OR2X2_1591 ( .A(u2__abc_52155_new_n9487_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9488_));
OR2X2 OR2X2_1592 ( .A(u2__abc_52155_new_n9486_), .B(u2__abc_52155_new_n9488_), .Y(u2__abc_52155_new_n9489_));
OR2X2 OR2X2_1593 ( .A(u2__abc_52155_new_n9493_), .B(u2__abc_52155_new_n9479_), .Y(u2__abc_52155_new_n9494_));
OR2X2 OR2X2_1594 ( .A(u2__abc_52155_new_n9425_), .B(u2__abc_52155_new_n3937_), .Y(u2__abc_52155_new_n9501_));
OR2X2 OR2X2_1595 ( .A(u2__abc_52155_new_n9461_), .B(u2__abc_52155_new_n3914_), .Y(u2__abc_52155_new_n9508_));
OR2X2 OR2X2_1596 ( .A(u2__abc_52155_new_n9512_), .B(u2__abc_52155_new_n3906_), .Y(u2__abc_52155_new_n9513_));
OR2X2 OR2X2_1597 ( .A(u2__abc_52155_new_n9519_), .B(u2__abc_52155_new_n9518_), .Y(u2__abc_52155_new_n9520_));
OR2X2 OR2X2_1598 ( .A(u2__abc_52155_new_n9520_), .B(u2__abc_52155_new_n3858_), .Y(u2__abc_52155_new_n9521_));
OR2X2 OR2X2_1599 ( .A(u2__abc_52155_new_n9524_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n9525_));
OR2X2 OR2X2_16 ( .A(_abc_73687_new_n753_), .B(\a[7] ), .Y(_abc_73687_new_n852_));
OR2X2 OR2X2_160 ( .A(_abc_73687_new_n753_), .B(\a[79] ), .Y(_abc_73687_new_n1068_));
OR2X2 OR2X2_1600 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_94_), .Y(u2__abc_52155_new_n9526_));
OR2X2 OR2X2_1601 ( .A(u2__abc_52155_new_n9527_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9528_));
OR2X2 OR2X2_1602 ( .A(u2__abc_52155_new_n9532_), .B(u2__abc_52155_new_n9496_), .Y(u2__abc_52155_new_n9533_));
OR2X2 OR2X2_1603 ( .A(u2__abc_52155_new_n9540_), .B(u2__abc_52155_new_n9537_), .Y(u2__abc_52155_new_n9541_));
OR2X2 OR2X2_1604 ( .A(u2__abc_52155_new_n9543_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9544_));
OR2X2 OR2X2_1605 ( .A(u2__abc_52155_new_n9542_), .B(u2__abc_52155_new_n9544_), .Y(u2__abc_52155_new_n9545_));
OR2X2 OR2X2_1606 ( .A(u2__abc_52155_new_n9549_), .B(u2__abc_52155_new_n9535_), .Y(u2__abc_52155_new_n9550_));
OR2X2 OR2X2_1607 ( .A(u2__abc_52155_new_n9555_), .B(u2__abc_52155_new_n3849_), .Y(u2__abc_52155_new_n9556_));
OR2X2 OR2X2_1608 ( .A(u2__abc_52155_new_n9557_), .B(u2__abc_52155_new_n9553_), .Y(u2__abc_52155_new_n9560_));
OR2X2 OR2X2_1609 ( .A(u2__abc_52155_new_n9563_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9564_));
OR2X2 OR2X2_161 ( .A(aNan), .B(sqrto_156_), .Y(_abc_73687_new_n1070_));
OR2X2 OR2X2_1610 ( .A(u2__abc_52155_new_n9562_), .B(u2__abc_52155_new_n9564_), .Y(u2__abc_52155_new_n9565_));
OR2X2 OR2X2_1611 ( .A(u2__abc_52155_new_n9569_), .B(u2__abc_52155_new_n9552_), .Y(u2__abc_52155_new_n9570_));
OR2X2 OR2X2_1612 ( .A(u2__abc_52155_new_n9574_), .B(u2__abc_52155_new_n3842_), .Y(u2__abc_52155_new_n9575_));
OR2X2 OR2X2_1613 ( .A(u2__abc_52155_new_n9577_), .B(u2__abc_52155_new_n9576_), .Y(u2__abc_52155_new_n9578_));
OR2X2 OR2X2_1614 ( .A(u2__abc_52155_new_n9581_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9582_));
OR2X2 OR2X2_1615 ( .A(u2__abc_52155_new_n9580_), .B(u2__abc_52155_new_n9582_), .Y(u2__abc_52155_new_n9583_));
OR2X2 OR2X2_1616 ( .A(u2__abc_52155_new_n9587_), .B(u2__abc_52155_new_n9572_), .Y(u2__abc_52155_new_n9588_));
OR2X2 OR2X2_1617 ( .A(u2__abc_52155_new_n9554_), .B(u2__abc_52155_new_n3849_), .Y(u2__abc_52155_new_n9591_));
OR2X2 OR2X2_1618 ( .A(u2__abc_52155_new_n9591_), .B(u2__abc_52155_new_n3843_), .Y(u2__abc_52155_new_n9592_));
OR2X2 OR2X2_1619 ( .A(u2__abc_52155_new_n9573_), .B(u2__abc_52155_new_n3841_), .Y(u2__abc_52155_new_n9593_));
OR2X2 OR2X2_162 ( .A(_abc_73687_new_n753_), .B(\a[80] ), .Y(_abc_73687_new_n1071_));
OR2X2 OR2X2_1620 ( .A(u2__abc_52155_new_n9597_), .B(u2__abc_52155_new_n9596_), .Y(u2__abc_52155_new_n9598_));
OR2X2 OR2X2_1621 ( .A(u2__abc_52155_new_n9598_), .B(u2__abc_52155_new_n3889_), .Y(u2__abc_52155_new_n9601_));
OR2X2 OR2X2_1622 ( .A(u2__abc_52155_new_n9604_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9605_));
OR2X2 OR2X2_1623 ( .A(u2__abc_52155_new_n9603_), .B(u2__abc_52155_new_n9605_), .Y(u2__abc_52155_new_n9606_));
OR2X2 OR2X2_1624 ( .A(u2__abc_52155_new_n9610_), .B(u2__abc_52155_new_n9590_), .Y(u2__abc_52155_new_n9611_));
OR2X2 OR2X2_1625 ( .A(u2__abc_52155_new_n9618_), .B(u2__abc_52155_new_n9615_), .Y(u2__abc_52155_new_n9619_));
OR2X2 OR2X2_1626 ( .A(u2__abc_52155_new_n9621_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9622_));
OR2X2 OR2X2_1627 ( .A(u2__abc_52155_new_n9620_), .B(u2__abc_52155_new_n9622_), .Y(u2__abc_52155_new_n9623_));
OR2X2 OR2X2_1628 ( .A(u2__abc_52155_new_n9627_), .B(u2__abc_52155_new_n9613_), .Y(u2__abc_52155_new_n9628_));
OR2X2 OR2X2_1629 ( .A(u2__abc_52155_new_n9632_), .B(u2__abc_52155_new_n3880_), .Y(u2__abc_52155_new_n9633_));
OR2X2 OR2X2_163 ( .A(aNan), .B(sqrto_157_), .Y(_abc_73687_new_n1073_));
OR2X2 OR2X2_1630 ( .A(u2__abc_52155_new_n9634_), .B(u2__abc_52155_new_n3867_), .Y(u2__abc_52155_new_n9637_));
OR2X2 OR2X2_1631 ( .A(u2__abc_52155_new_n9640_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9641_));
OR2X2 OR2X2_1632 ( .A(u2__abc_52155_new_n9639_), .B(u2__abc_52155_new_n9641_), .Y(u2__abc_52155_new_n9642_));
OR2X2 OR2X2_1633 ( .A(u2__abc_52155_new_n9646_), .B(u2__abc_52155_new_n9630_), .Y(u2__abc_52155_new_n9647_));
OR2X2 OR2X2_1634 ( .A(u2__abc_52155_new_n9651_), .B(u2__abc_52155_new_n9650_), .Y(u2__abc_52155_new_n9652_));
OR2X2 OR2X2_1635 ( .A(u2__abc_52155_new_n9653_), .B(u2__abc_52155_new_n3874_), .Y(u2__abc_52155_new_n9654_));
OR2X2 OR2X2_1636 ( .A(u2__abc_52155_new_n9657_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9658_));
OR2X2 OR2X2_1637 ( .A(u2__abc_52155_new_n9656_), .B(u2__abc_52155_new_n9658_), .Y(u2__abc_52155_new_n9659_));
OR2X2 OR2X2_1638 ( .A(u2__abc_52155_new_n9663_), .B(u2__abc_52155_new_n9649_), .Y(u2__abc_52155_new_n9664_));
OR2X2 OR2X2_1639 ( .A(u2__abc_52155_new_n9631_), .B(u2__abc_52155_new_n3880_), .Y(u2__abc_52155_new_n9668_));
OR2X2 OR2X2_164 ( .A(_abc_73687_new_n753_), .B(\a[81] ), .Y(_abc_73687_new_n1074_));
OR2X2 OR2X2_1640 ( .A(u2__abc_52155_new_n9671_), .B(u2__abc_52155_new_n3869_), .Y(u2__abc_52155_new_n9672_));
OR2X2 OR2X2_1641 ( .A(u2__abc_52155_new_n9670_), .B(u2__abc_52155_new_n9672_), .Y(u2__abc_52155_new_n9673_));
OR2X2 OR2X2_1642 ( .A(u2__abc_52155_new_n9667_), .B(u2__abc_52155_new_n9673_), .Y(u2__abc_52155_new_n9674_));
OR2X2 OR2X2_1643 ( .A(u2__abc_52155_new_n9675_), .B(u2__abc_52155_new_n9674_), .Y(u2__abc_52155_new_n9676_));
OR2X2 OR2X2_1644 ( .A(u2__abc_52155_new_n9676_), .B(u2__abc_52155_new_n3798_), .Y(u2__abc_52155_new_n9679_));
OR2X2 OR2X2_1645 ( .A(u2__abc_52155_new_n9682_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9683_));
OR2X2 OR2X2_1646 ( .A(u2__abc_52155_new_n9681_), .B(u2__abc_52155_new_n9683_), .Y(u2__abc_52155_new_n9684_));
OR2X2 OR2X2_1647 ( .A(u2__abc_52155_new_n9688_), .B(u2__abc_52155_new_n9666_), .Y(u2__abc_52155_new_n9689_));
OR2X2 OR2X2_1648 ( .A(u2__abc_52155_new_n9696_), .B(u2__abc_52155_new_n9693_), .Y(u2__abc_52155_new_n9697_));
OR2X2 OR2X2_1649 ( .A(u2__abc_52155_new_n9699_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9700_));
OR2X2 OR2X2_165 ( .A(aNan), .B(sqrto_158_), .Y(_abc_73687_new_n1076_));
OR2X2 OR2X2_1650 ( .A(u2__abc_52155_new_n9698_), .B(u2__abc_52155_new_n9700_), .Y(u2__abc_52155_new_n9701_));
OR2X2 OR2X2_1651 ( .A(u2__abc_52155_new_n9705_), .B(u2__abc_52155_new_n9691_), .Y(u2__abc_52155_new_n9706_));
OR2X2 OR2X2_1652 ( .A(u2__abc_52155_new_n9710_), .B(u2__abc_52155_new_n3789_), .Y(u2__abc_52155_new_n9711_));
OR2X2 OR2X2_1653 ( .A(u2__abc_52155_new_n9712_), .B(u2__abc_52155_new_n3776_), .Y(u2__abc_52155_new_n9715_));
OR2X2 OR2X2_1654 ( .A(u2__abc_52155_new_n9718_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9719_));
OR2X2 OR2X2_1655 ( .A(u2__abc_52155_new_n9717_), .B(u2__abc_52155_new_n9719_), .Y(u2__abc_52155_new_n9720_));
OR2X2 OR2X2_1656 ( .A(u2__abc_52155_new_n9724_), .B(u2__abc_52155_new_n9708_), .Y(u2__abc_52155_new_n9725_));
OR2X2 OR2X2_1657 ( .A(u2__abc_52155_new_n9729_), .B(u2__abc_52155_new_n9728_), .Y(u2__abc_52155_new_n9730_));
OR2X2 OR2X2_1658 ( .A(u2__abc_52155_new_n9731_), .B(u2__abc_52155_new_n3783_), .Y(u2__abc_52155_new_n9732_));
OR2X2 OR2X2_1659 ( .A(u2__abc_52155_new_n9735_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9736_));
OR2X2 OR2X2_166 ( .A(_abc_73687_new_n753_), .B(\a[82] ), .Y(_abc_73687_new_n1077_));
OR2X2 OR2X2_1660 ( .A(u2__abc_52155_new_n9734_), .B(u2__abc_52155_new_n9736_), .Y(u2__abc_52155_new_n9737_));
OR2X2 OR2X2_1661 ( .A(u2__abc_52155_new_n9741_), .B(u2__abc_52155_new_n9727_), .Y(u2__abc_52155_new_n9742_));
OR2X2 OR2X2_1662 ( .A(u2__abc_52155_new_n9709_), .B(u2__abc_52155_new_n3789_), .Y(u2__abc_52155_new_n9745_));
OR2X2 OR2X2_1663 ( .A(u2__abc_52155_new_n9748_), .B(u2__abc_52155_new_n3778_), .Y(u2__abc_52155_new_n9749_));
OR2X2 OR2X2_1664 ( .A(u2__abc_52155_new_n9747_), .B(u2__abc_52155_new_n9749_), .Y(u2__abc_52155_new_n9750_));
OR2X2 OR2X2_1665 ( .A(u2__abc_52155_new_n9751_), .B(u2__abc_52155_new_n9750_), .Y(u2__abc_52155_new_n9752_));
OR2X2 OR2X2_1666 ( .A(u2__abc_52155_new_n9752_), .B(u2__abc_52155_new_n3829_), .Y(u2__abc_52155_new_n9755_));
OR2X2 OR2X2_1667 ( .A(u2__abc_52155_new_n9758_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9759_));
OR2X2 OR2X2_1668 ( .A(u2__abc_52155_new_n9757_), .B(u2__abc_52155_new_n9759_), .Y(u2__abc_52155_new_n9760_));
OR2X2 OR2X2_1669 ( .A(u2__abc_52155_new_n9764_), .B(u2__abc_52155_new_n9744_), .Y(u2__abc_52155_new_n9765_));
OR2X2 OR2X2_167 ( .A(aNan), .B(sqrto_159_), .Y(_abc_73687_new_n1079_));
OR2X2 OR2X2_1670 ( .A(u2__abc_52155_new_n9772_), .B(u2__abc_52155_new_n9769_), .Y(u2__abc_52155_new_n9773_));
OR2X2 OR2X2_1671 ( .A(u2__abc_52155_new_n9775_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9776_));
OR2X2 OR2X2_1672 ( .A(u2__abc_52155_new_n9774_), .B(u2__abc_52155_new_n9776_), .Y(u2__abc_52155_new_n9777_));
OR2X2 OR2X2_1673 ( .A(u2__abc_52155_new_n9781_), .B(u2__abc_52155_new_n9767_), .Y(u2__abc_52155_new_n9782_));
OR2X2 OR2X2_1674 ( .A(u2__abc_52155_new_n9786_), .B(u2__abc_52155_new_n3820_), .Y(u2__abc_52155_new_n9787_));
OR2X2 OR2X2_1675 ( .A(u2__abc_52155_new_n9788_), .B(u2__abc_52155_new_n3807_), .Y(u2__abc_52155_new_n9791_));
OR2X2 OR2X2_1676 ( .A(u2__abc_52155_new_n9794_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9795_));
OR2X2 OR2X2_1677 ( .A(u2__abc_52155_new_n9793_), .B(u2__abc_52155_new_n9795_), .Y(u2__abc_52155_new_n9796_));
OR2X2 OR2X2_1678 ( .A(u2__abc_52155_new_n9800_), .B(u2__abc_52155_new_n9784_), .Y(u2__abc_52155_new_n9801_));
OR2X2 OR2X2_1679 ( .A(u2__abc_52155_new_n9808_), .B(u2__abc_52155_new_n9805_), .Y(u2__abc_52155_new_n9809_));
OR2X2 OR2X2_168 ( .A(_abc_73687_new_n753_), .B(\a[83] ), .Y(_abc_73687_new_n1080_));
OR2X2 OR2X2_1680 ( .A(u2__abc_52155_new_n9811_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9812_));
OR2X2 OR2X2_1681 ( .A(u2__abc_52155_new_n9810_), .B(u2__abc_52155_new_n9812_), .Y(u2__abc_52155_new_n9813_));
OR2X2 OR2X2_1682 ( .A(u2__abc_52155_new_n9817_), .B(u2__abc_52155_new_n9803_), .Y(u2__abc_52155_new_n9818_));
OR2X2 OR2X2_1683 ( .A(u2__abc_52155_new_n9785_), .B(u2__abc_52155_new_n3820_), .Y(u2__abc_52155_new_n9823_));
OR2X2 OR2X2_1684 ( .A(u2__abc_52155_new_n9826_), .B(u2__abc_52155_new_n3809_), .Y(u2__abc_52155_new_n9827_));
OR2X2 OR2X2_1685 ( .A(u2__abc_52155_new_n9825_), .B(u2__abc_52155_new_n9827_), .Y(u2__abc_52155_new_n9828_));
OR2X2 OR2X2_1686 ( .A(u2__abc_52155_new_n9822_), .B(u2__abc_52155_new_n9828_), .Y(u2__abc_52155_new_n9829_));
OR2X2 OR2X2_1687 ( .A(u2__abc_52155_new_n9821_), .B(u2__abc_52155_new_n9829_), .Y(u2__abc_52155_new_n9830_));
OR2X2 OR2X2_1688 ( .A(u2__abc_52155_new_n9831_), .B(u2__abc_52155_new_n9830_), .Y(u2__abc_52155_new_n9832_));
OR2X2 OR2X2_1689 ( .A(u2__abc_52155_new_n9832_), .B(u2__abc_52155_new_n3712_), .Y(u2__abc_52155_new_n9835_));
OR2X2 OR2X2_169 ( .A(aNan), .B(sqrto_160_), .Y(_abc_73687_new_n1082_));
OR2X2 OR2X2_1690 ( .A(u2__abc_52155_new_n9838_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9839_));
OR2X2 OR2X2_1691 ( .A(u2__abc_52155_new_n9837_), .B(u2__abc_52155_new_n9839_), .Y(u2__abc_52155_new_n9840_));
OR2X2 OR2X2_1692 ( .A(u2__abc_52155_new_n9844_), .B(u2__abc_52155_new_n9820_), .Y(u2__abc_52155_new_n9845_));
OR2X2 OR2X2_1693 ( .A(u2__abc_52155_new_n9849_), .B(u2__abc_52155_new_n9848_), .Y(u2__abc_52155_new_n9850_));
OR2X2 OR2X2_1694 ( .A(u2__abc_52155_new_n9851_), .B(u2__abc_52155_new_n3719_), .Y(u2__abc_52155_new_n9852_));
OR2X2 OR2X2_1695 ( .A(u2__abc_52155_new_n9855_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9856_));
OR2X2 OR2X2_1696 ( .A(u2__abc_52155_new_n9854_), .B(u2__abc_52155_new_n9856_), .Y(u2__abc_52155_new_n9857_));
OR2X2 OR2X2_1697 ( .A(u2__abc_52155_new_n9861_), .B(u2__abc_52155_new_n9847_), .Y(u2__abc_52155_new_n9862_));
OR2X2 OR2X2_1698 ( .A(u2__abc_52155_new_n3708_), .B(u2__abc_52155_new_n3717_), .Y(u2__abc_52155_new_n9865_));
OR2X2 OR2X2_1699 ( .A(u2__abc_52155_new_n9868_), .B(u2__abc_52155_new_n9867_), .Y(u2__abc_52155_new_n9869_));
OR2X2 OR2X2_17 ( .A(aNan), .B(sqrto_84_), .Y(_abc_73687_new_n854_));
OR2X2 OR2X2_170 ( .A(_abc_73687_new_n753_), .B(\a[84] ), .Y(_abc_73687_new_n1083_));
OR2X2 OR2X2_1700 ( .A(u2__abc_52155_new_n9869_), .B(u2__abc_52155_new_n3727_), .Y(u2__abc_52155_new_n9872_));
OR2X2 OR2X2_1701 ( .A(u2__abc_52155_new_n9875_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9876_));
OR2X2 OR2X2_1702 ( .A(u2__abc_52155_new_n9874_), .B(u2__abc_52155_new_n9876_), .Y(u2__abc_52155_new_n9877_));
OR2X2 OR2X2_1703 ( .A(u2__abc_52155_new_n9881_), .B(u2__abc_52155_new_n9864_), .Y(u2__abc_52155_new_n9882_));
OR2X2 OR2X2_1704 ( .A(u2__abc_52155_new_n9886_), .B(u2__abc_52155_new_n9885_), .Y(u2__abc_52155_new_n9887_));
OR2X2 OR2X2_1705 ( .A(u2__abc_52155_new_n9888_), .B(u2__abc_52155_new_n3734_), .Y(u2__abc_52155_new_n9889_));
OR2X2 OR2X2_1706 ( .A(u2__abc_52155_new_n9892_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9893_));
OR2X2 OR2X2_1707 ( .A(u2__abc_52155_new_n9891_), .B(u2__abc_52155_new_n9893_), .Y(u2__abc_52155_new_n9894_));
OR2X2 OR2X2_1708 ( .A(u2__abc_52155_new_n9898_), .B(u2__abc_52155_new_n9884_), .Y(u2__abc_52155_new_n9899_));
OR2X2 OR2X2_1709 ( .A(u2__abc_52155_new_n9903_), .B(u2__abc_52155_new_n3729_), .Y(u2__abc_52155_new_n9904_));
OR2X2 OR2X2_171 ( .A(aNan), .B(sqrto_161_), .Y(_abc_73687_new_n1085_));
OR2X2 OR2X2_1710 ( .A(u2__abc_52155_new_n9902_), .B(u2__abc_52155_new_n9904_), .Y(u2__abc_52155_new_n9905_));
OR2X2 OR2X2_1711 ( .A(u2__abc_52155_new_n9906_), .B(u2__abc_52155_new_n9905_), .Y(u2__abc_52155_new_n9907_));
OR2X2 OR2X2_1712 ( .A(u2__abc_52155_new_n9907_), .B(u2__abc_52155_new_n3765_), .Y(u2__abc_52155_new_n9910_));
OR2X2 OR2X2_1713 ( .A(u2__abc_52155_new_n9913_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9914_));
OR2X2 OR2X2_1714 ( .A(u2__abc_52155_new_n9912_), .B(u2__abc_52155_new_n9914_), .Y(u2__abc_52155_new_n9915_));
OR2X2 OR2X2_1715 ( .A(u2__abc_52155_new_n9919_), .B(u2__abc_52155_new_n9901_), .Y(u2__abc_52155_new_n9920_));
OR2X2 OR2X2_1716 ( .A(u2__abc_52155_new_n9924_), .B(u2__abc_52155_new_n3758_), .Y(u2__abc_52155_new_n9927_));
OR2X2 OR2X2_1717 ( .A(u2__abc_52155_new_n9930_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9931_));
OR2X2 OR2X2_1718 ( .A(u2__abc_52155_new_n9929_), .B(u2__abc_52155_new_n9931_), .Y(u2__abc_52155_new_n9932_));
OR2X2 OR2X2_1719 ( .A(u2__abc_52155_new_n9936_), .B(u2__abc_52155_new_n9922_), .Y(u2__abc_52155_new_n9937_));
OR2X2 OR2X2_172 ( .A(_abc_73687_new_n753_), .B(\a[85] ), .Y(_abc_73687_new_n1086_));
OR2X2 OR2X2_1720 ( .A(u2__abc_52155_new_n9941_), .B(u2__abc_52155_new_n3743_), .Y(u2__abc_52155_new_n9944_));
OR2X2 OR2X2_1721 ( .A(u2__abc_52155_new_n9947_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9948_));
OR2X2 OR2X2_1722 ( .A(u2__abc_52155_new_n9946_), .B(u2__abc_52155_new_n9948_), .Y(u2__abc_52155_new_n9949_));
OR2X2 OR2X2_1723 ( .A(u2__abc_52155_new_n9953_), .B(u2__abc_52155_new_n9939_), .Y(u2__abc_52155_new_n9954_));
OR2X2 OR2X2_1724 ( .A(u2__abc_52155_new_n9961_), .B(u2__abc_52155_new_n9958_), .Y(u2__abc_52155_new_n9962_));
OR2X2 OR2X2_1725 ( .A(u2__abc_52155_new_n9964_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9965_));
OR2X2 OR2X2_1726 ( .A(u2__abc_52155_new_n9963_), .B(u2__abc_52155_new_n9965_), .Y(u2__abc_52155_new_n9966_));
OR2X2 OR2X2_1727 ( .A(u2__abc_52155_new_n9970_), .B(u2__abc_52155_new_n9956_), .Y(u2__abc_52155_new_n9971_));
OR2X2 OR2X2_1728 ( .A(u2__abc_52155_new_n3753_), .B(u2__abc_52155_new_n3760_), .Y(u2__abc_52155_new_n9975_));
OR2X2 OR2X2_1729 ( .A(u2__abc_52155_new_n9978_), .B(u2__abc_52155_new_n3745_), .Y(u2__abc_52155_new_n9979_));
OR2X2 OR2X2_173 ( .A(aNan), .B(sqrto_162_), .Y(_abc_73687_new_n1088_));
OR2X2 OR2X2_1730 ( .A(u2__abc_52155_new_n9977_), .B(u2__abc_52155_new_n9979_), .Y(u2__abc_52155_new_n9980_));
OR2X2 OR2X2_1731 ( .A(u2__abc_52155_new_n9974_), .B(u2__abc_52155_new_n9980_), .Y(u2__abc_52155_new_n9981_));
OR2X2 OR2X2_1732 ( .A(u2__abc_52155_new_n9982_), .B(u2__abc_52155_new_n9981_), .Y(u2__abc_52155_new_n9983_));
OR2X2 OR2X2_1733 ( .A(u2__abc_52155_new_n9983_), .B(u2__abc_52155_new_n3649_), .Y(u2__abc_52155_new_n9986_));
OR2X2 OR2X2_1734 ( .A(u2__abc_52155_new_n9989_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n9990_));
OR2X2 OR2X2_1735 ( .A(u2__abc_52155_new_n9988_), .B(u2__abc_52155_new_n9990_), .Y(u2__abc_52155_new_n9991_));
OR2X2 OR2X2_1736 ( .A(u2__abc_52155_new_n9995_), .B(u2__abc_52155_new_n9973_), .Y(u2__abc_52155_new_n9996_));
OR2X2 OR2X2_1737 ( .A(u2__abc_52155_new_n10000_), .B(u2__abc_52155_new_n9999_), .Y(u2__abc_52155_new_n10001_));
OR2X2 OR2X2_1738 ( .A(u2__abc_52155_new_n10002_), .B(u2__abc_52155_new_n3656_), .Y(u2__abc_52155_new_n10003_));
OR2X2 OR2X2_1739 ( .A(u2__abc_52155_new_n10006_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10007_));
OR2X2 OR2X2_174 ( .A(_abc_73687_new_n753_), .B(\a[86] ), .Y(_abc_73687_new_n1089_));
OR2X2 OR2X2_1740 ( .A(u2__abc_52155_new_n10005_), .B(u2__abc_52155_new_n10007_), .Y(u2__abc_52155_new_n10008_));
OR2X2 OR2X2_1741 ( .A(u2__abc_52155_new_n10012_), .B(u2__abc_52155_new_n9998_), .Y(u2__abc_52155_new_n10013_));
OR2X2 OR2X2_1742 ( .A(u2__abc_52155_new_n3645_), .B(u2__abc_52155_new_n3654_), .Y(u2__abc_52155_new_n10016_));
OR2X2 OR2X2_1743 ( .A(u2__abc_52155_new_n10019_), .B(u2__abc_52155_new_n10018_), .Y(u2__abc_52155_new_n10020_));
OR2X2 OR2X2_1744 ( .A(u2__abc_52155_new_n10020_), .B(u2__abc_52155_new_n3664_), .Y(u2__abc_52155_new_n10023_));
OR2X2 OR2X2_1745 ( .A(u2__abc_52155_new_n10026_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10027_));
OR2X2 OR2X2_1746 ( .A(u2__abc_52155_new_n10025_), .B(u2__abc_52155_new_n10027_), .Y(u2__abc_52155_new_n10028_));
OR2X2 OR2X2_1747 ( .A(u2__abc_52155_new_n10032_), .B(u2__abc_52155_new_n10015_), .Y(u2__abc_52155_new_n10033_));
OR2X2 OR2X2_1748 ( .A(u2__abc_52155_new_n10040_), .B(u2__abc_52155_new_n10037_), .Y(u2__abc_52155_new_n10041_));
OR2X2 OR2X2_1749 ( .A(u2__abc_52155_new_n10043_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10044_));
OR2X2 OR2X2_175 ( .A(aNan), .B(sqrto_163_), .Y(_abc_73687_new_n1091_));
OR2X2 OR2X2_1750 ( .A(u2__abc_52155_new_n10042_), .B(u2__abc_52155_new_n10044_), .Y(u2__abc_52155_new_n10045_));
OR2X2 OR2X2_1751 ( .A(u2__abc_52155_new_n10049_), .B(u2__abc_52155_new_n10035_), .Y(u2__abc_52155_new_n10050_));
OR2X2 OR2X2_1752 ( .A(u2__abc_52155_new_n10054_), .B(u2__abc_52155_new_n3666_), .Y(u2__abc_52155_new_n10055_));
OR2X2 OR2X2_1753 ( .A(u2__abc_52155_new_n10053_), .B(u2__abc_52155_new_n10055_), .Y(u2__abc_52155_new_n10056_));
OR2X2 OR2X2_1754 ( .A(u2__abc_52155_new_n10057_), .B(u2__abc_52155_new_n10056_), .Y(u2__abc_52155_new_n10058_));
OR2X2 OR2X2_1755 ( .A(u2__abc_52155_new_n10058_), .B(u2__abc_52155_new_n3702_), .Y(u2__abc_52155_new_n10061_));
OR2X2 OR2X2_1756 ( .A(u2__abc_52155_new_n10064_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10065_));
OR2X2 OR2X2_1757 ( .A(u2__abc_52155_new_n10063_), .B(u2__abc_52155_new_n10065_), .Y(u2__abc_52155_new_n10066_));
OR2X2 OR2X2_1758 ( .A(u2__abc_52155_new_n10070_), .B(u2__abc_52155_new_n10052_), .Y(u2__abc_52155_new_n10071_));
OR2X2 OR2X2_1759 ( .A(u2__abc_52155_new_n10078_), .B(u2__abc_52155_new_n10075_), .Y(u2__abc_52155_new_n10079_));
OR2X2 OR2X2_176 ( .A(_abc_73687_new_n753_), .B(\a[87] ), .Y(_abc_73687_new_n1092_));
OR2X2 OR2X2_1760 ( .A(u2__abc_52155_new_n10081_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10082_));
OR2X2 OR2X2_1761 ( .A(u2__abc_52155_new_n10080_), .B(u2__abc_52155_new_n10082_), .Y(u2__abc_52155_new_n10083_));
OR2X2 OR2X2_1762 ( .A(u2__abc_52155_new_n10087_), .B(u2__abc_52155_new_n10073_), .Y(u2__abc_52155_new_n10088_));
OR2X2 OR2X2_1763 ( .A(u2__abc_52155_new_n10092_), .B(u2__abc_52155_new_n3693_), .Y(u2__abc_52155_new_n10093_));
OR2X2 OR2X2_1764 ( .A(u2__abc_52155_new_n10094_), .B(u2__abc_52155_new_n3680_), .Y(u2__abc_52155_new_n10097_));
OR2X2 OR2X2_1765 ( .A(u2__abc_52155_new_n10100_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10101_));
OR2X2 OR2X2_1766 ( .A(u2__abc_52155_new_n10099_), .B(u2__abc_52155_new_n10101_), .Y(u2__abc_52155_new_n10102_));
OR2X2 OR2X2_1767 ( .A(u2__abc_52155_new_n10107_), .B(u2__abc_52155_new_n10090_), .Y(u2__abc_52155_new_n10108_));
OR2X2 OR2X2_1768 ( .A(u2__abc_52155_new_n10115_), .B(u2__abc_52155_new_n10112_), .Y(u2__abc_52155_new_n10116_));
OR2X2 OR2X2_1769 ( .A(u2__abc_52155_new_n10118_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10119_));
OR2X2 OR2X2_177 ( .A(aNan), .B(sqrto_164_), .Y(_abc_73687_new_n1094_));
OR2X2 OR2X2_1770 ( .A(u2__abc_52155_new_n10117_), .B(u2__abc_52155_new_n10119_), .Y(u2__abc_52155_new_n10120_));
OR2X2 OR2X2_1771 ( .A(u2__abc_52155_new_n10124_), .B(u2__abc_52155_new_n10110_), .Y(u2__abc_52155_new_n10125_));
OR2X2 OR2X2_1772 ( .A(u2__abc_52155_new_n10138_), .B(u2__abc_52155_new_n3682_), .Y(u2__abc_52155_new_n10139_));
OR2X2 OR2X2_1773 ( .A(u2__abc_52155_new_n10091_), .B(u2__abc_52155_new_n3693_), .Y(u2__abc_52155_new_n10140_));
OR2X2 OR2X2_1774 ( .A(u2__abc_52155_new_n10150_), .B(u2__abc_52155_new_n5237_), .Y(u2__abc_52155_new_n10153_));
OR2X2 OR2X2_1775 ( .A(u2__abc_52155_new_n10154_), .B(u2__abc_52155_new_n7623_), .Y(u2__abc_52155_new_n10155_));
OR2X2 OR2X2_1776 ( .A(u2__abc_52155_new_n7622_), .B(u2_remHi_126_), .Y(u2__abc_52155_new_n10156_));
OR2X2 OR2X2_1777 ( .A(u2__abc_52155_new_n10157_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10158_));
OR2X2 OR2X2_1778 ( .A(u2__abc_52155_new_n10162_), .B(u2__abc_52155_new_n10127_), .Y(u2__abc_52155_new_n10163_));
OR2X2 OR2X2_1779 ( .A(u2__abc_52155_new_n10167_), .B(u2__abc_52155_new_n10166_), .Y(u2__abc_52155_new_n10168_));
OR2X2 OR2X2_178 ( .A(_abc_73687_new_n753_), .B(\a[88] ), .Y(_abc_73687_new_n1095_));
OR2X2 OR2X2_1780 ( .A(u2__abc_52155_new_n10169_), .B(u2__abc_52155_new_n5244_), .Y(u2__abc_52155_new_n10170_));
OR2X2 OR2X2_1781 ( .A(u2__abc_52155_new_n10173_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10174_));
OR2X2 OR2X2_1782 ( .A(u2__abc_52155_new_n10172_), .B(u2__abc_52155_new_n10174_), .Y(u2__abc_52155_new_n10175_));
OR2X2 OR2X2_1783 ( .A(u2__abc_52155_new_n10179_), .B(u2__abc_52155_new_n10165_), .Y(u2__abc_52155_new_n10180_));
OR2X2 OR2X2_1784 ( .A(u2__abc_52155_new_n5235_), .B(u2__abc_52155_new_n5242_), .Y(u2__abc_52155_new_n10184_));
OR2X2 OR2X2_1785 ( .A(u2__abc_52155_new_n10187_), .B(u2__abc_52155_new_n10186_), .Y(u2__abc_52155_new_n10188_));
OR2X2 OR2X2_1786 ( .A(u2__abc_52155_new_n10188_), .B(u2__abc_52155_new_n10183_), .Y(u2__abc_52155_new_n10191_));
OR2X2 OR2X2_1787 ( .A(u2__abc_52155_new_n10194_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10195_));
OR2X2 OR2X2_1788 ( .A(u2__abc_52155_new_n10193_), .B(u2__abc_52155_new_n10195_), .Y(u2__abc_52155_new_n10196_));
OR2X2 OR2X2_1789 ( .A(u2__abc_52155_new_n10200_), .B(u2__abc_52155_new_n10182_), .Y(u2__abc_52155_new_n10201_));
OR2X2 OR2X2_179 ( .A(aNan), .B(sqrto_165_), .Y(_abc_73687_new_n1097_));
OR2X2 OR2X2_1790 ( .A(u2__abc_52155_new_n10205_), .B(u2__abc_52155_new_n5255_), .Y(u2__abc_52155_new_n10206_));
OR2X2 OR2X2_1791 ( .A(u2__abc_52155_new_n10208_), .B(u2__abc_52155_new_n10207_), .Y(u2__abc_52155_new_n10209_));
OR2X2 OR2X2_1792 ( .A(u2__abc_52155_new_n10212_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10213_));
OR2X2 OR2X2_1793 ( .A(u2__abc_52155_new_n10211_), .B(u2__abc_52155_new_n10213_), .Y(u2__abc_52155_new_n10214_));
OR2X2 OR2X2_1794 ( .A(u2__abc_52155_new_n10218_), .B(u2__abc_52155_new_n10203_), .Y(u2__abc_52155_new_n10219_));
OR2X2 OR2X2_1795 ( .A(u2__abc_52155_new_n10224_), .B(u2__abc_52155_new_n5252_), .Y(u2__abc_52155_new_n10225_));
OR2X2 OR2X2_1796 ( .A(u2__abc_52155_new_n10223_), .B(u2__abc_52155_new_n10225_), .Y(u2__abc_52155_new_n10226_));
OR2X2 OR2X2_1797 ( .A(u2__abc_52155_new_n10227_), .B(u2__abc_52155_new_n10226_), .Y(u2__abc_52155_new_n10228_));
OR2X2 OR2X2_1798 ( .A(u2__abc_52155_new_n10228_), .B(u2__abc_52155_new_n10222_), .Y(u2__abc_52155_new_n10231_));
OR2X2 OR2X2_1799 ( .A(u2__abc_52155_new_n10234_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10235_));
OR2X2 OR2X2_18 ( .A(_abc_73687_new_n753_), .B(\a[8] ), .Y(_abc_73687_new_n855_));
OR2X2 OR2X2_180 ( .A(_abc_73687_new_n753_), .B(\a[89] ), .Y(_abc_73687_new_n1098_));
OR2X2 OR2X2_1800 ( .A(u2__abc_52155_new_n10233_), .B(u2__abc_52155_new_n10235_), .Y(u2__abc_52155_new_n10236_));
OR2X2 OR2X2_1801 ( .A(u2__abc_52155_new_n10240_), .B(u2__abc_52155_new_n10221_), .Y(u2__abc_52155_new_n10241_));
OR2X2 OR2X2_1802 ( .A(u2__abc_52155_new_n10249_), .B(u2__abc_52155_new_n10247_), .Y(u2__abc_52155_new_n10250_));
OR2X2 OR2X2_1803 ( .A(u2__abc_52155_new_n10252_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10253_));
OR2X2 OR2X2_1804 ( .A(u2__abc_52155_new_n10251_), .B(u2__abc_52155_new_n10253_), .Y(u2__abc_52155_new_n10254_));
OR2X2 OR2X2_1805 ( .A(u2__abc_52155_new_n10258_), .B(u2__abc_52155_new_n10243_), .Y(u2__abc_52155_new_n10259_));
OR2X2 OR2X2_1806 ( .A(u2__abc_52155_new_n5271_), .B(u2__abc_52155_new_n5276_), .Y(u2__abc_52155_new_n10263_));
OR2X2 OR2X2_1807 ( .A(u2__abc_52155_new_n10265_), .B(u2__abc_52155_new_n5273_), .Y(u2__abc_52155_new_n10266_));
OR2X2 OR2X2_1808 ( .A(u2__abc_52155_new_n10267_), .B(u2__abc_52155_new_n10262_), .Y(u2__abc_52155_new_n10270_));
OR2X2 OR2X2_1809 ( .A(u2__abc_52155_new_n10273_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10274_));
OR2X2 OR2X2_181 ( .A(aNan), .B(sqrto_166_), .Y(_abc_73687_new_n1100_));
OR2X2 OR2X2_1810 ( .A(u2__abc_52155_new_n10272_), .B(u2__abc_52155_new_n10274_), .Y(u2__abc_52155_new_n10275_));
OR2X2 OR2X2_1811 ( .A(u2__abc_52155_new_n10279_), .B(u2__abc_52155_new_n10261_), .Y(u2__abc_52155_new_n10280_));
OR2X2 OR2X2_1812 ( .A(u2__abc_52155_new_n10284_), .B(u2__abc_52155_new_n5268_), .Y(u2__abc_52155_new_n10285_));
OR2X2 OR2X2_1813 ( .A(u2__abc_52155_new_n10287_), .B(u2__abc_52155_new_n10286_), .Y(u2__abc_52155_new_n10288_));
OR2X2 OR2X2_1814 ( .A(u2__abc_52155_new_n10291_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10292_));
OR2X2 OR2X2_1815 ( .A(u2__abc_52155_new_n10290_), .B(u2__abc_52155_new_n10292_), .Y(u2__abc_52155_new_n10293_));
OR2X2 OR2X2_1816 ( .A(u2__abc_52155_new_n10297_), .B(u2__abc_52155_new_n10282_), .Y(u2__abc_52155_new_n10298_));
OR2X2 OR2X2_1817 ( .A(u2__abc_52155_new_n10264_), .B(u2__abc_52155_new_n5273_), .Y(u2__abc_52155_new_n10303_));
OR2X2 OR2X2_1818 ( .A(u2__abc_52155_new_n10303_), .B(u2__abc_52155_new_n5269_), .Y(u2__abc_52155_new_n10304_));
OR2X2 OR2X2_1819 ( .A(u2__abc_52155_new_n10283_), .B(u2__abc_52155_new_n5267_), .Y(u2__abc_52155_new_n10305_));
OR2X2 OR2X2_182 ( .A(_abc_73687_new_n753_), .B(\a[90] ), .Y(_abc_73687_new_n1101_));
OR2X2 OR2X2_1820 ( .A(u2__abc_52155_new_n10310_), .B(u2__abc_52155_new_n10309_), .Y(u2__abc_52155_new_n10311_));
OR2X2 OR2X2_1821 ( .A(u2__abc_52155_new_n10311_), .B(u2__abc_52155_new_n5191_), .Y(u2__abc_52155_new_n10314_));
OR2X2 OR2X2_1822 ( .A(u2__abc_52155_new_n10317_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10318_));
OR2X2 OR2X2_1823 ( .A(u2__abc_52155_new_n10316_), .B(u2__abc_52155_new_n10318_), .Y(u2__abc_52155_new_n10319_));
OR2X2 OR2X2_1824 ( .A(u2__abc_52155_new_n10323_), .B(u2__abc_52155_new_n10300_), .Y(u2__abc_52155_new_n10324_));
OR2X2 OR2X2_1825 ( .A(u2__abc_52155_new_n10330_), .B(u2__abc_52155_new_n10331_), .Y(u2__abc_52155_new_n10332_));
OR2X2 OR2X2_1826 ( .A(u2__abc_52155_new_n10334_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10335_));
OR2X2 OR2X2_1827 ( .A(u2__abc_52155_new_n10333_), .B(u2__abc_52155_new_n10335_), .Y(u2__abc_52155_new_n10336_));
OR2X2 OR2X2_1828 ( .A(u2__abc_52155_new_n10340_), .B(u2__abc_52155_new_n10326_), .Y(u2__abc_52155_new_n10341_));
OR2X2 OR2X2_1829 ( .A(u2__abc_52155_new_n10345_), .B(u2__abc_52155_new_n5193_), .Y(u2__abc_52155_new_n10346_));
OR2X2 OR2X2_183 ( .A(aNan), .B(sqrto_167_), .Y(_abc_73687_new_n1103_));
OR2X2 OR2X2_1830 ( .A(u2__abc_52155_new_n10346_), .B(u2__abc_52155_new_n10344_), .Y(u2__abc_52155_new_n10349_));
OR2X2 OR2X2_1831 ( .A(u2__abc_52155_new_n10352_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10353_));
OR2X2 OR2X2_1832 ( .A(u2__abc_52155_new_n10351_), .B(u2__abc_52155_new_n10353_), .Y(u2__abc_52155_new_n10354_));
OR2X2 OR2X2_1833 ( .A(u2__abc_52155_new_n10358_), .B(u2__abc_52155_new_n10343_), .Y(u2__abc_52155_new_n10359_));
OR2X2 OR2X2_1834 ( .A(u2__abc_52155_new_n10363_), .B(u2__abc_52155_new_n5182_), .Y(u2__abc_52155_new_n10364_));
OR2X2 OR2X2_1835 ( .A(u2__abc_52155_new_n10366_), .B(u2__abc_52155_new_n10365_), .Y(u2__abc_52155_new_n10367_));
OR2X2 OR2X2_1836 ( .A(u2__abc_52155_new_n10370_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10371_));
OR2X2 OR2X2_1837 ( .A(u2__abc_52155_new_n10369_), .B(u2__abc_52155_new_n10371_), .Y(u2__abc_52155_new_n10372_));
OR2X2 OR2X2_1838 ( .A(u2__abc_52155_new_n10376_), .B(u2__abc_52155_new_n10361_), .Y(u2__abc_52155_new_n10377_));
OR2X2 OR2X2_1839 ( .A(u2__abc_52155_new_n10380_), .B(u2__abc_52155_new_n5196_), .Y(u2__abc_52155_new_n10381_));
OR2X2 OR2X2_184 ( .A(_abc_73687_new_n753_), .B(\a[91] ), .Y(_abc_73687_new_n1104_));
OR2X2 OR2X2_1840 ( .A(u2__abc_52155_new_n10381_), .B(u2__abc_52155_new_n5183_), .Y(u2__abc_52155_new_n10382_));
OR2X2 OR2X2_1841 ( .A(u2__abc_52155_new_n10362_), .B(u2__abc_52155_new_n5181_), .Y(u2__abc_52155_new_n10383_));
OR2X2 OR2X2_1842 ( .A(u2__abc_52155_new_n10387_), .B(u2__abc_52155_new_n10386_), .Y(u2__abc_52155_new_n10388_));
OR2X2 OR2X2_1843 ( .A(u2__abc_52155_new_n10388_), .B(u2__abc_52155_new_n5229_), .Y(u2__abc_52155_new_n10391_));
OR2X2 OR2X2_1844 ( .A(u2__abc_52155_new_n10394_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10395_));
OR2X2 OR2X2_1845 ( .A(u2__abc_52155_new_n10393_), .B(u2__abc_52155_new_n10395_), .Y(u2__abc_52155_new_n10396_));
OR2X2 OR2X2_1846 ( .A(u2__abc_52155_new_n10400_), .B(u2__abc_52155_new_n10379_), .Y(u2__abc_52155_new_n10401_));
OR2X2 OR2X2_1847 ( .A(u2__abc_52155_new_n10408_), .B(u2__abc_52155_new_n10405_), .Y(u2__abc_52155_new_n10409_));
OR2X2 OR2X2_1848 ( .A(u2__abc_52155_new_n10411_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10412_));
OR2X2 OR2X2_1849 ( .A(u2__abc_52155_new_n10410_), .B(u2__abc_52155_new_n10412_), .Y(u2__abc_52155_new_n10413_));
OR2X2 OR2X2_185 ( .A(aNan), .B(sqrto_168_), .Y(_abc_73687_new_n1106_));
OR2X2 OR2X2_1850 ( .A(u2__abc_52155_new_n10417_), .B(u2__abc_52155_new_n10403_), .Y(u2__abc_52155_new_n10418_));
OR2X2 OR2X2_1851 ( .A(u2__abc_52155_new_n10422_), .B(u2__abc_52155_new_n5220_), .Y(u2__abc_52155_new_n10423_));
OR2X2 OR2X2_1852 ( .A(u2__abc_52155_new_n10424_), .B(u2__abc_52155_new_n5207_), .Y(u2__abc_52155_new_n10427_));
OR2X2 OR2X2_1853 ( .A(u2__abc_52155_new_n10430_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10431_));
OR2X2 OR2X2_1854 ( .A(u2__abc_52155_new_n10429_), .B(u2__abc_52155_new_n10431_), .Y(u2__abc_52155_new_n10432_));
OR2X2 OR2X2_1855 ( .A(u2__abc_52155_new_n10436_), .B(u2__abc_52155_new_n10420_), .Y(u2__abc_52155_new_n10437_));
OR2X2 OR2X2_1856 ( .A(u2__abc_52155_new_n10444_), .B(u2__abc_52155_new_n10441_), .Y(u2__abc_52155_new_n10445_));
OR2X2 OR2X2_1857 ( .A(u2__abc_52155_new_n10447_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10448_));
OR2X2 OR2X2_1858 ( .A(u2__abc_52155_new_n10446_), .B(u2__abc_52155_new_n10448_), .Y(u2__abc_52155_new_n10449_));
OR2X2 OR2X2_1859 ( .A(u2__abc_52155_new_n10453_), .B(u2__abc_52155_new_n10439_), .Y(u2__abc_52155_new_n10454_));
OR2X2 OR2X2_186 ( .A(_abc_73687_new_n753_), .B(\a[92] ), .Y(_abc_73687_new_n1107_));
OR2X2 OR2X2_1860 ( .A(u2__abc_52155_new_n10421_), .B(u2__abc_52155_new_n5220_), .Y(u2__abc_52155_new_n10459_));
OR2X2 OR2X2_1861 ( .A(u2__abc_52155_new_n10462_), .B(u2__abc_52155_new_n5209_), .Y(u2__abc_52155_new_n10463_));
OR2X2 OR2X2_1862 ( .A(u2__abc_52155_new_n10461_), .B(u2__abc_52155_new_n10463_), .Y(u2__abc_52155_new_n10464_));
OR2X2 OR2X2_1863 ( .A(u2__abc_52155_new_n10458_), .B(u2__abc_52155_new_n10464_), .Y(u2__abc_52155_new_n10465_));
OR2X2 OR2X2_1864 ( .A(u2__abc_52155_new_n10457_), .B(u2__abc_52155_new_n10465_), .Y(u2__abc_52155_new_n10466_));
OR2X2 OR2X2_1865 ( .A(u2__abc_52155_new_n10467_), .B(u2__abc_52155_new_n10466_), .Y(u2__abc_52155_new_n10468_));
OR2X2 OR2X2_1866 ( .A(u2__abc_52155_new_n10468_), .B(u2__abc_52155_new_n5168_), .Y(u2__abc_52155_new_n10471_));
OR2X2 OR2X2_1867 ( .A(u2__abc_52155_new_n10474_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10475_));
OR2X2 OR2X2_1868 ( .A(u2__abc_52155_new_n10473_), .B(u2__abc_52155_new_n10475_), .Y(u2__abc_52155_new_n10476_));
OR2X2 OR2X2_1869 ( .A(u2__abc_52155_new_n10480_), .B(u2__abc_52155_new_n10456_), .Y(u2__abc_52155_new_n10481_));
OR2X2 OR2X2_187 ( .A(aNan), .B(sqrto_169_), .Y(_abc_73687_new_n1109_));
OR2X2 OR2X2_1870 ( .A(u2__abc_52155_new_n10487_), .B(u2__abc_52155_new_n10488_), .Y(u2__abc_52155_new_n10489_));
OR2X2 OR2X2_1871 ( .A(u2__abc_52155_new_n10491_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10492_));
OR2X2 OR2X2_1872 ( .A(u2__abc_52155_new_n10490_), .B(u2__abc_52155_new_n10492_), .Y(u2__abc_52155_new_n10493_));
OR2X2 OR2X2_1873 ( .A(u2__abc_52155_new_n10497_), .B(u2__abc_52155_new_n10483_), .Y(u2__abc_52155_new_n10498_));
OR2X2 OR2X2_1874 ( .A(u2__abc_52155_new_n10502_), .B(u2__abc_52155_new_n5156_), .Y(u2__abc_52155_new_n10503_));
OR2X2 OR2X2_1875 ( .A(u2__abc_52155_new_n10503_), .B(u2__abc_52155_new_n10501_), .Y(u2__abc_52155_new_n10506_));
OR2X2 OR2X2_1876 ( .A(u2__abc_52155_new_n10509_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10510_));
OR2X2 OR2X2_1877 ( .A(u2__abc_52155_new_n10508_), .B(u2__abc_52155_new_n10510_), .Y(u2__abc_52155_new_n10511_));
OR2X2 OR2X2_1878 ( .A(u2__abc_52155_new_n10515_), .B(u2__abc_52155_new_n10500_), .Y(u2__abc_52155_new_n10516_));
OR2X2 OR2X2_1879 ( .A(u2__abc_52155_new_n10520_), .B(u2__abc_52155_new_n5152_), .Y(u2__abc_52155_new_n10521_));
OR2X2 OR2X2_188 ( .A(_abc_73687_new_n753_), .B(\a[93] ), .Y(_abc_73687_new_n1110_));
OR2X2 OR2X2_1880 ( .A(u2__abc_52155_new_n10523_), .B(u2__abc_52155_new_n10522_), .Y(u2__abc_52155_new_n10524_));
OR2X2 OR2X2_1881 ( .A(u2__abc_52155_new_n10527_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10528_));
OR2X2 OR2X2_1882 ( .A(u2__abc_52155_new_n10526_), .B(u2__abc_52155_new_n10528_), .Y(u2__abc_52155_new_n10529_));
OR2X2 OR2X2_1883 ( .A(u2__abc_52155_new_n10533_), .B(u2__abc_52155_new_n10518_), .Y(u2__abc_52155_new_n10534_));
OR2X2 OR2X2_1884 ( .A(u2__abc_52155_new_n10538_), .B(u2__abc_52155_new_n5151_), .Y(u2__abc_52155_new_n10539_));
OR2X2 OR2X2_1885 ( .A(u2__abc_52155_new_n10540_), .B(u2__abc_52155_new_n5140_), .Y(u2__abc_52155_new_n10543_));
OR2X2 OR2X2_1886 ( .A(u2__abc_52155_new_n10546_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10547_));
OR2X2 OR2X2_1887 ( .A(u2__abc_52155_new_n10545_), .B(u2__abc_52155_new_n10547_), .Y(u2__abc_52155_new_n10548_));
OR2X2 OR2X2_1888 ( .A(u2__abc_52155_new_n10552_), .B(u2__abc_52155_new_n10536_), .Y(u2__abc_52155_new_n10553_));
OR2X2 OR2X2_1889 ( .A(u2__abc_52155_new_n10557_), .B(u2__abc_52155_new_n5133_), .Y(u2__abc_52155_new_n10560_));
OR2X2 OR2X2_189 ( .A(aNan), .B(sqrto_170_), .Y(_abc_73687_new_n1112_));
OR2X2 OR2X2_1890 ( .A(u2__abc_52155_new_n10563_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10564_));
OR2X2 OR2X2_1891 ( .A(u2__abc_52155_new_n10562_), .B(u2__abc_52155_new_n10564_), .Y(u2__abc_52155_new_n10565_));
OR2X2 OR2X2_1892 ( .A(u2__abc_52155_new_n10569_), .B(u2__abc_52155_new_n10555_), .Y(u2__abc_52155_new_n10570_));
OR2X2 OR2X2_1893 ( .A(u2__abc_52155_new_n10574_), .B(u2__abc_52155_new_n5118_), .Y(u2__abc_52155_new_n10577_));
OR2X2 OR2X2_1894 ( .A(u2__abc_52155_new_n10580_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10581_));
OR2X2 OR2X2_1895 ( .A(u2__abc_52155_new_n10579_), .B(u2__abc_52155_new_n10581_), .Y(u2__abc_52155_new_n10582_));
OR2X2 OR2X2_1896 ( .A(u2__abc_52155_new_n10586_), .B(u2__abc_52155_new_n10572_), .Y(u2__abc_52155_new_n10587_));
OR2X2 OR2X2_1897 ( .A(u2__abc_52155_new_n10594_), .B(u2__abc_52155_new_n10591_), .Y(u2__abc_52155_new_n10595_));
OR2X2 OR2X2_1898 ( .A(u2__abc_52155_new_n10597_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10598_));
OR2X2 OR2X2_1899 ( .A(u2__abc_52155_new_n10596_), .B(u2__abc_52155_new_n10598_), .Y(u2__abc_52155_new_n10599_));
OR2X2 OR2X2_19 ( .A(aNan), .B(sqrto_85_), .Y(_abc_73687_new_n857_));
OR2X2 OR2X2_190 ( .A(_abc_73687_new_n753_), .B(\a[94] ), .Y(_abc_73687_new_n1113_));
OR2X2 OR2X2_1900 ( .A(u2__abc_52155_new_n10603_), .B(u2__abc_52155_new_n10589_), .Y(u2__abc_52155_new_n10604_));
OR2X2 OR2X2_1901 ( .A(u2__abc_52155_new_n10537_), .B(u2__abc_52155_new_n5151_), .Y(u2__abc_52155_new_n10607_));
OR2X2 OR2X2_1902 ( .A(u2__abc_52155_new_n10608_), .B(u2__abc_52155_new_n5159_), .Y(u2__abc_52155_new_n10609_));
OR2X2 OR2X2_1903 ( .A(u2__abc_52155_new_n10609_), .B(u2__abc_52155_new_n5153_), .Y(u2__abc_52155_new_n10610_));
OR2X2 OR2X2_1904 ( .A(u2__abc_52155_new_n10611_), .B(u2__abc_52155_new_n5138_), .Y(u2__abc_52155_new_n10612_));
OR2X2 OR2X2_1905 ( .A(u2__abc_52155_new_n5116_), .B(u2__abc_52155_new_n5131_), .Y(u2__abc_52155_new_n10615_));
OR2X2 OR2X2_1906 ( .A(u2__abc_52155_new_n10614_), .B(u2__abc_52155_new_n10615_), .Y(u2__abc_52155_new_n10616_));
OR2X2 OR2X2_1907 ( .A(u2__abc_52155_new_n10617_), .B(u2__abc_52155_new_n5123_), .Y(u2__abc_52155_new_n10618_));
OR2X2 OR2X2_1908 ( .A(u2__abc_52155_new_n10621_), .B(u2__abc_52155_new_n10620_), .Y(u2__abc_52155_new_n10622_));
OR2X2 OR2X2_1909 ( .A(u2__abc_52155_new_n10622_), .B(u2__abc_52155_new_n5077_), .Y(u2__abc_52155_new_n10625_));
OR2X2 OR2X2_191 ( .A(aNan), .B(sqrto_171_), .Y(_abc_73687_new_n1115_));
OR2X2 OR2X2_1910 ( .A(u2__abc_52155_new_n10628_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10629_));
OR2X2 OR2X2_1911 ( .A(u2__abc_52155_new_n10627_), .B(u2__abc_52155_new_n10629_), .Y(u2__abc_52155_new_n10630_));
OR2X2 OR2X2_1912 ( .A(u2__abc_52155_new_n10634_), .B(u2__abc_52155_new_n10606_), .Y(u2__abc_52155_new_n10635_));
OR2X2 OR2X2_1913 ( .A(u2__abc_52155_new_n10642_), .B(u2__abc_52155_new_n10639_), .Y(u2__abc_52155_new_n10643_));
OR2X2 OR2X2_1914 ( .A(u2__abc_52155_new_n10645_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10646_));
OR2X2 OR2X2_1915 ( .A(u2__abc_52155_new_n10644_), .B(u2__abc_52155_new_n10646_), .Y(u2__abc_52155_new_n10647_));
OR2X2 OR2X2_1916 ( .A(u2__abc_52155_new_n10651_), .B(u2__abc_52155_new_n10637_), .Y(u2__abc_52155_new_n10652_));
OR2X2 OR2X2_1917 ( .A(u2__abc_52155_new_n10656_), .B(u2__abc_52155_new_n5068_), .Y(u2__abc_52155_new_n10657_));
OR2X2 OR2X2_1918 ( .A(u2__abc_52155_new_n10658_), .B(u2__abc_52155_new_n5055_), .Y(u2__abc_52155_new_n10661_));
OR2X2 OR2X2_1919 ( .A(u2__abc_52155_new_n10664_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10665_));
OR2X2 OR2X2_192 ( .A(_abc_73687_new_n753_), .B(\a[95] ), .Y(_abc_73687_new_n1116_));
OR2X2 OR2X2_1920 ( .A(u2__abc_52155_new_n10663_), .B(u2__abc_52155_new_n10665_), .Y(u2__abc_52155_new_n10666_));
OR2X2 OR2X2_1921 ( .A(u2__abc_52155_new_n10670_), .B(u2__abc_52155_new_n10654_), .Y(u2__abc_52155_new_n10671_));
OR2X2 OR2X2_1922 ( .A(u2__abc_52155_new_n10678_), .B(u2__abc_52155_new_n10675_), .Y(u2__abc_52155_new_n10679_));
OR2X2 OR2X2_1923 ( .A(u2__abc_52155_new_n10681_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10682_));
OR2X2 OR2X2_1924 ( .A(u2__abc_52155_new_n10680_), .B(u2__abc_52155_new_n10682_), .Y(u2__abc_52155_new_n10683_));
OR2X2 OR2X2_1925 ( .A(u2__abc_52155_new_n10687_), .B(u2__abc_52155_new_n10673_), .Y(u2__abc_52155_new_n10688_));
OR2X2 OR2X2_1926 ( .A(u2__abc_52155_new_n10655_), .B(u2__abc_52155_new_n5068_), .Y(u2__abc_52155_new_n10691_));
OR2X2 OR2X2_1927 ( .A(u2__abc_52155_new_n10694_), .B(u2__abc_52155_new_n5057_), .Y(u2__abc_52155_new_n10695_));
OR2X2 OR2X2_1928 ( .A(u2__abc_52155_new_n10693_), .B(u2__abc_52155_new_n10695_), .Y(u2__abc_52155_new_n10696_));
OR2X2 OR2X2_1929 ( .A(u2__abc_52155_new_n10697_), .B(u2__abc_52155_new_n10696_), .Y(u2__abc_52155_new_n10698_));
OR2X2 OR2X2_193 ( .A(aNan), .B(sqrto_172_), .Y(_abc_73687_new_n1118_));
OR2X2 OR2X2_1930 ( .A(u2__abc_52155_new_n10698_), .B(u2__abc_52155_new_n5108_), .Y(u2__abc_52155_new_n10701_));
OR2X2 OR2X2_1931 ( .A(u2__abc_52155_new_n10704_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10705_));
OR2X2 OR2X2_1932 ( .A(u2__abc_52155_new_n10703_), .B(u2__abc_52155_new_n10705_), .Y(u2__abc_52155_new_n10706_));
OR2X2 OR2X2_1933 ( .A(u2__abc_52155_new_n10710_), .B(u2__abc_52155_new_n10690_), .Y(u2__abc_52155_new_n10711_));
OR2X2 OR2X2_1934 ( .A(u2__abc_52155_new_n10718_), .B(u2__abc_52155_new_n10715_), .Y(u2__abc_52155_new_n10719_));
OR2X2 OR2X2_1935 ( .A(u2__abc_52155_new_n10721_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10722_));
OR2X2 OR2X2_1936 ( .A(u2__abc_52155_new_n10720_), .B(u2__abc_52155_new_n10722_), .Y(u2__abc_52155_new_n10723_));
OR2X2 OR2X2_1937 ( .A(u2__abc_52155_new_n10727_), .B(u2__abc_52155_new_n10713_), .Y(u2__abc_52155_new_n10728_));
OR2X2 OR2X2_1938 ( .A(u2__abc_52155_new_n10732_), .B(u2__abc_52155_new_n5099_), .Y(u2__abc_52155_new_n10733_));
OR2X2 OR2X2_1939 ( .A(u2__abc_52155_new_n10734_), .B(u2__abc_52155_new_n5086_), .Y(u2__abc_52155_new_n10737_));
OR2X2 OR2X2_194 ( .A(_abc_73687_new_n753_), .B(\a[96] ), .Y(_abc_73687_new_n1119_));
OR2X2 OR2X2_1940 ( .A(u2__abc_52155_new_n10740_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10741_));
OR2X2 OR2X2_1941 ( .A(u2__abc_52155_new_n10739_), .B(u2__abc_52155_new_n10741_), .Y(u2__abc_52155_new_n10742_));
OR2X2 OR2X2_1942 ( .A(u2__abc_52155_new_n10746_), .B(u2__abc_52155_new_n10730_), .Y(u2__abc_52155_new_n10747_));
OR2X2 OR2X2_1943 ( .A(u2__abc_52155_new_n10754_), .B(u2__abc_52155_new_n10751_), .Y(u2__abc_52155_new_n10755_));
OR2X2 OR2X2_1944 ( .A(u2__abc_52155_new_n10757_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10758_));
OR2X2 OR2X2_1945 ( .A(u2__abc_52155_new_n10756_), .B(u2__abc_52155_new_n10758_), .Y(u2__abc_52155_new_n10759_));
OR2X2 OR2X2_1946 ( .A(u2__abc_52155_new_n10763_), .B(u2__abc_52155_new_n10749_), .Y(u2__abc_52155_new_n10764_));
OR2X2 OR2X2_1947 ( .A(u2__abc_52155_new_n10731_), .B(u2__abc_52155_new_n5099_), .Y(u2__abc_52155_new_n10770_));
OR2X2 OR2X2_1948 ( .A(u2__abc_52155_new_n10773_), .B(u2__abc_52155_new_n5088_), .Y(u2__abc_52155_new_n10774_));
OR2X2 OR2X2_1949 ( .A(u2__abc_52155_new_n10772_), .B(u2__abc_52155_new_n10774_), .Y(u2__abc_52155_new_n10775_));
OR2X2 OR2X2_195 ( .A(aNan), .B(sqrto_173_), .Y(_abc_73687_new_n1121_));
OR2X2 OR2X2_1950 ( .A(u2__abc_52155_new_n10769_), .B(u2__abc_52155_new_n10775_), .Y(u2__abc_52155_new_n10776_));
OR2X2 OR2X2_1951 ( .A(u2__abc_52155_new_n10768_), .B(u2__abc_52155_new_n10776_), .Y(u2__abc_52155_new_n10777_));
OR2X2 OR2X2_1952 ( .A(u2__abc_52155_new_n10777_), .B(u2__abc_52155_new_n10767_), .Y(u2__abc_52155_new_n10778_));
OR2X2 OR2X2_1953 ( .A(u2__abc_52155_new_n10779_), .B(u2__abc_52155_new_n10778_), .Y(u2__abc_52155_new_n10780_));
OR2X2 OR2X2_1954 ( .A(u2__abc_52155_new_n10780_), .B(u2__abc_52155_new_n5012_), .Y(u2__abc_52155_new_n10783_));
OR2X2 OR2X2_1955 ( .A(u2__abc_52155_new_n10786_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10787_));
OR2X2 OR2X2_1956 ( .A(u2__abc_52155_new_n10785_), .B(u2__abc_52155_new_n10787_), .Y(u2__abc_52155_new_n10788_));
OR2X2 OR2X2_1957 ( .A(u2__abc_52155_new_n10792_), .B(u2__abc_52155_new_n10766_), .Y(u2__abc_52155_new_n10793_));
OR2X2 OR2X2_1958 ( .A(u2__abc_52155_new_n10800_), .B(u2__abc_52155_new_n10797_), .Y(u2__abc_52155_new_n10801_));
OR2X2 OR2X2_1959 ( .A(u2__abc_52155_new_n10803_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10804_));
OR2X2 OR2X2_196 ( .A(_abc_73687_new_n753_), .B(\a[97] ), .Y(_abc_73687_new_n1122_));
OR2X2 OR2X2_1960 ( .A(u2__abc_52155_new_n10802_), .B(u2__abc_52155_new_n10804_), .Y(u2__abc_52155_new_n10805_));
OR2X2 OR2X2_1961 ( .A(u2__abc_52155_new_n10809_), .B(u2__abc_52155_new_n10795_), .Y(u2__abc_52155_new_n10810_));
OR2X2 OR2X2_1962 ( .A(u2__abc_52155_new_n10815_), .B(u2__abc_52155_new_n5003_), .Y(u2__abc_52155_new_n10816_));
OR2X2 OR2X2_1963 ( .A(u2__abc_52155_new_n10817_), .B(u2__abc_52155_new_n10813_), .Y(u2__abc_52155_new_n10820_));
OR2X2 OR2X2_1964 ( .A(u2__abc_52155_new_n10823_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10824_));
OR2X2 OR2X2_1965 ( .A(u2__abc_52155_new_n10822_), .B(u2__abc_52155_new_n10824_), .Y(u2__abc_52155_new_n10825_));
OR2X2 OR2X2_1966 ( .A(u2__abc_52155_new_n10829_), .B(u2__abc_52155_new_n10812_), .Y(u2__abc_52155_new_n10830_));
OR2X2 OR2X2_1967 ( .A(u2__abc_52155_new_n10834_), .B(u2__abc_52155_new_n4996_), .Y(u2__abc_52155_new_n10835_));
OR2X2 OR2X2_1968 ( .A(u2__abc_52155_new_n10837_), .B(u2__abc_52155_new_n10836_), .Y(u2__abc_52155_new_n10838_));
OR2X2 OR2X2_1969 ( .A(u2__abc_52155_new_n10841_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10842_));
OR2X2 OR2X2_197 ( .A(aNan), .B(sqrto_174_), .Y(_abc_73687_new_n1124_));
OR2X2 OR2X2_1970 ( .A(u2__abc_52155_new_n10840_), .B(u2__abc_52155_new_n10842_), .Y(u2__abc_52155_new_n10843_));
OR2X2 OR2X2_1971 ( .A(u2__abc_52155_new_n10847_), .B(u2__abc_52155_new_n10832_), .Y(u2__abc_52155_new_n10848_));
OR2X2 OR2X2_1972 ( .A(u2__abc_52155_new_n10814_), .B(u2__abc_52155_new_n5003_), .Y(u2__abc_52155_new_n10851_));
OR2X2 OR2X2_1973 ( .A(u2__abc_52155_new_n10851_), .B(u2__abc_52155_new_n4997_), .Y(u2__abc_52155_new_n10852_));
OR2X2 OR2X2_1974 ( .A(u2__abc_52155_new_n10833_), .B(u2__abc_52155_new_n4995_), .Y(u2__abc_52155_new_n10853_));
OR2X2 OR2X2_1975 ( .A(u2__abc_52155_new_n10857_), .B(u2__abc_52155_new_n10856_), .Y(u2__abc_52155_new_n10858_));
OR2X2 OR2X2_1976 ( .A(u2__abc_52155_new_n10858_), .B(u2__abc_52155_new_n5043_), .Y(u2__abc_52155_new_n10861_));
OR2X2 OR2X2_1977 ( .A(u2__abc_52155_new_n10864_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10865_));
OR2X2 OR2X2_1978 ( .A(u2__abc_52155_new_n10863_), .B(u2__abc_52155_new_n10865_), .Y(u2__abc_52155_new_n10866_));
OR2X2 OR2X2_1979 ( .A(u2__abc_52155_new_n10870_), .B(u2__abc_52155_new_n10850_), .Y(u2__abc_52155_new_n10871_));
OR2X2 OR2X2_198 ( .A(_abc_73687_new_n753_), .B(\a[98] ), .Y(_abc_73687_new_n1125_));
OR2X2 OR2X2_1980 ( .A(u2__abc_52155_new_n10875_), .B(u2__abc_52155_new_n5036_), .Y(u2__abc_52155_new_n10878_));
OR2X2 OR2X2_1981 ( .A(u2__abc_52155_new_n10881_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10882_));
OR2X2 OR2X2_1982 ( .A(u2__abc_52155_new_n10880_), .B(u2__abc_52155_new_n10882_), .Y(u2__abc_52155_new_n10883_));
OR2X2 OR2X2_1983 ( .A(u2__abc_52155_new_n10887_), .B(u2__abc_52155_new_n10873_), .Y(u2__abc_52155_new_n10888_));
OR2X2 OR2X2_1984 ( .A(u2__abc_52155_new_n10892_), .B(u2__abc_52155_new_n5021_), .Y(u2__abc_52155_new_n10895_));
OR2X2 OR2X2_1985 ( .A(u2__abc_52155_new_n10898_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10899_));
OR2X2 OR2X2_1986 ( .A(u2__abc_52155_new_n10897_), .B(u2__abc_52155_new_n10899_), .Y(u2__abc_52155_new_n10900_));
OR2X2 OR2X2_1987 ( .A(u2__abc_52155_new_n10904_), .B(u2__abc_52155_new_n10890_), .Y(u2__abc_52155_new_n10905_));
OR2X2 OR2X2_1988 ( .A(u2__abc_52155_new_n10912_), .B(u2__abc_52155_new_n10909_), .Y(u2__abc_52155_new_n10913_));
OR2X2 OR2X2_1989 ( .A(u2__abc_52155_new_n10915_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10916_));
OR2X2 OR2X2_199 ( .A(aNan), .B(sqrto_175_), .Y(_abc_73687_new_n1127_));
OR2X2 OR2X2_1990 ( .A(u2__abc_52155_new_n10914_), .B(u2__abc_52155_new_n10916_), .Y(u2__abc_52155_new_n10917_));
OR2X2 OR2X2_1991 ( .A(u2__abc_52155_new_n10921_), .B(u2__abc_52155_new_n10907_), .Y(u2__abc_52155_new_n10922_));
OR2X2 OR2X2_1992 ( .A(u2__abc_52155_new_n5031_), .B(u2__abc_52155_new_n5038_), .Y(u2__abc_52155_new_n10926_));
OR2X2 OR2X2_1993 ( .A(u2__abc_52155_new_n10929_), .B(u2__abc_52155_new_n5023_), .Y(u2__abc_52155_new_n10930_));
OR2X2 OR2X2_1994 ( .A(u2__abc_52155_new_n10928_), .B(u2__abc_52155_new_n10930_), .Y(u2__abc_52155_new_n10931_));
OR2X2 OR2X2_1995 ( .A(u2__abc_52155_new_n10925_), .B(u2__abc_52155_new_n10931_), .Y(u2__abc_52155_new_n10932_));
OR2X2 OR2X2_1996 ( .A(u2__abc_52155_new_n10933_), .B(u2__abc_52155_new_n10932_), .Y(u2__abc_52155_new_n10934_));
OR2X2 OR2X2_1997 ( .A(u2__abc_52155_new_n10934_), .B(u2__abc_52155_new_n4983_), .Y(u2__abc_52155_new_n10937_));
OR2X2 OR2X2_1998 ( .A(u2__abc_52155_new_n10940_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10941_));
OR2X2 OR2X2_1999 ( .A(u2__abc_52155_new_n10939_), .B(u2__abc_52155_new_n10941_), .Y(u2__abc_52155_new_n10942_));
OR2X2 OR2X2_2 ( .A(_abc_73687_new_n753_), .B(\a[0] ), .Y(_abc_73687_new_n831_));
OR2X2 OR2X2_20 ( .A(_abc_73687_new_n753_), .B(\a[9] ), .Y(_abc_73687_new_n858_));
OR2X2 OR2X2_200 ( .A(_abc_73687_new_n753_), .B(\a[99] ), .Y(_abc_73687_new_n1128_));
OR2X2 OR2X2_2000 ( .A(u2__abc_52155_new_n10946_), .B(u2__abc_52155_new_n10924_), .Y(u2__abc_52155_new_n10947_));
OR2X2 OR2X2_2001 ( .A(u2__abc_52155_new_n10953_), .B(u2__abc_52155_new_n10954_), .Y(u2__abc_52155_new_n10955_));
OR2X2 OR2X2_2002 ( .A(u2__abc_52155_new_n10957_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10958_));
OR2X2 OR2X2_2003 ( .A(u2__abc_52155_new_n10956_), .B(u2__abc_52155_new_n10958_), .Y(u2__abc_52155_new_n10959_));
OR2X2 OR2X2_2004 ( .A(u2__abc_52155_new_n10963_), .B(u2__abc_52155_new_n10949_), .Y(u2__abc_52155_new_n10964_));
OR2X2 OR2X2_2005 ( .A(u2__abc_52155_new_n10967_), .B(u2__abc_52155_new_n4974_), .Y(u2__abc_52155_new_n10968_));
OR2X2 OR2X2_2006 ( .A(u2__abc_52155_new_n10970_), .B(u2__abc_52155_new_n10969_), .Y(u2__abc_52155_new_n10971_));
OR2X2 OR2X2_2007 ( .A(u2__abc_52155_new_n10971_), .B(u2__abc_52155_new_n4961_), .Y(u2__abc_52155_new_n10974_));
OR2X2 OR2X2_2008 ( .A(u2__abc_52155_new_n10977_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10978_));
OR2X2 OR2X2_2009 ( .A(u2__abc_52155_new_n10976_), .B(u2__abc_52155_new_n10978_), .Y(u2__abc_52155_new_n10979_));
OR2X2 OR2X2_201 ( .A(aNan), .B(sqrto_176_), .Y(_abc_73687_new_n1130_));
OR2X2 OR2X2_2010 ( .A(u2__abc_52155_new_n10983_), .B(u2__abc_52155_new_n10966_), .Y(u2__abc_52155_new_n10984_));
OR2X2 OR2X2_2011 ( .A(u2__abc_52155_new_n10991_), .B(u2__abc_52155_new_n10988_), .Y(u2__abc_52155_new_n10992_));
OR2X2 OR2X2_2012 ( .A(u2__abc_52155_new_n10994_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n10995_));
OR2X2 OR2X2_2013 ( .A(u2__abc_52155_new_n10993_), .B(u2__abc_52155_new_n10995_), .Y(u2__abc_52155_new_n10996_));
OR2X2 OR2X2_2014 ( .A(u2__abc_52155_new_n11000_), .B(u2__abc_52155_new_n10986_), .Y(u2__abc_52155_new_n11001_));
OR2X2 OR2X2_2015 ( .A(u2__abc_52155_new_n11005_), .B(u2__abc_52155_new_n4966_), .Y(u2__abc_52155_new_n11006_));
OR2X2 OR2X2_2016 ( .A(u2__abc_52155_new_n11007_), .B(u2__abc_52155_new_n4952_), .Y(u2__abc_52155_new_n11010_));
OR2X2 OR2X2_2017 ( .A(u2__abc_52155_new_n11013_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11014_));
OR2X2 OR2X2_2018 ( .A(u2__abc_52155_new_n11012_), .B(u2__abc_52155_new_n11014_), .Y(u2__abc_52155_new_n11015_));
OR2X2 OR2X2_2019 ( .A(u2__abc_52155_new_n11019_), .B(u2__abc_52155_new_n11003_), .Y(u2__abc_52155_new_n11020_));
OR2X2 OR2X2_202 ( .A(_abc_73687_new_n753_), .B(\a[100] ), .Y(_abc_73687_new_n1131_));
OR2X2 OR2X2_2020 ( .A(u2__abc_52155_new_n11027_), .B(u2__abc_52155_new_n11024_), .Y(u2__abc_52155_new_n11028_));
OR2X2 OR2X2_2021 ( .A(u2__abc_52155_new_n11030_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11031_));
OR2X2 OR2X2_2022 ( .A(u2__abc_52155_new_n11029_), .B(u2__abc_52155_new_n11031_), .Y(u2__abc_52155_new_n11032_));
OR2X2 OR2X2_2023 ( .A(u2__abc_52155_new_n11036_), .B(u2__abc_52155_new_n11022_), .Y(u2__abc_52155_new_n11037_));
OR2X2 OR2X2_2024 ( .A(u2__abc_52155_new_n11041_), .B(u2__abc_52155_new_n4943_), .Y(u2__abc_52155_new_n11042_));
OR2X2 OR2X2_2025 ( .A(u2__abc_52155_new_n11043_), .B(u2__abc_52155_new_n4930_), .Y(u2__abc_52155_new_n11046_));
OR2X2 OR2X2_2026 ( .A(u2__abc_52155_new_n11049_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11050_));
OR2X2 OR2X2_2027 ( .A(u2__abc_52155_new_n11048_), .B(u2__abc_52155_new_n11050_), .Y(u2__abc_52155_new_n11051_));
OR2X2 OR2X2_2028 ( .A(u2__abc_52155_new_n11055_), .B(u2__abc_52155_new_n11039_), .Y(u2__abc_52155_new_n11056_));
OR2X2 OR2X2_2029 ( .A(u2__abc_52155_new_n11063_), .B(u2__abc_52155_new_n11060_), .Y(u2__abc_52155_new_n11064_));
OR2X2 OR2X2_203 ( .A(aNan), .B(sqrto_177_), .Y(_abc_73687_new_n1133_));
OR2X2 OR2X2_2030 ( .A(u2__abc_52155_new_n11066_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11067_));
OR2X2 OR2X2_2031 ( .A(u2__abc_52155_new_n11065_), .B(u2__abc_52155_new_n11067_), .Y(u2__abc_52155_new_n11068_));
OR2X2 OR2X2_2032 ( .A(u2__abc_52155_new_n11072_), .B(u2__abc_52155_new_n11058_), .Y(u2__abc_52155_new_n11073_));
OR2X2 OR2X2_2033 ( .A(u2__abc_52155_new_n11004_), .B(u2__abc_52155_new_n4966_), .Y(u2__abc_52155_new_n11078_));
OR2X2 OR2X2_2034 ( .A(u2__abc_52155_new_n11040_), .B(u2__abc_52155_new_n4943_), .Y(u2__abc_52155_new_n11085_));
OR2X2 OR2X2_2035 ( .A(u2__abc_52155_new_n11089_), .B(u2__abc_52155_new_n4935_), .Y(u2__abc_52155_new_n11090_));
OR2X2 OR2X2_2036 ( .A(u2__abc_52155_new_n11095_), .B(u2__abc_52155_new_n11094_), .Y(u2__abc_52155_new_n11096_));
OR2X2 OR2X2_2037 ( .A(u2__abc_52155_new_n11096_), .B(u2__abc_52155_new_n4912_), .Y(u2__abc_52155_new_n11099_));
OR2X2 OR2X2_2038 ( .A(u2__abc_52155_new_n11102_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11103_));
OR2X2 OR2X2_2039 ( .A(u2__abc_52155_new_n11101_), .B(u2__abc_52155_new_n11103_), .Y(u2__abc_52155_new_n11104_));
OR2X2 OR2X2_204 ( .A(_abc_73687_new_n753_), .B(\a[101] ), .Y(_abc_73687_new_n1134_));
OR2X2 OR2X2_2040 ( .A(u2__abc_52155_new_n11108_), .B(u2__abc_52155_new_n11075_), .Y(u2__abc_52155_new_n11109_));
OR2X2 OR2X2_2041 ( .A(u2__abc_52155_new_n11113_), .B(u2__abc_52155_new_n11112_), .Y(u2__abc_52155_new_n11114_));
OR2X2 OR2X2_2042 ( .A(u2__abc_52155_new_n11115_), .B(u2__abc_52155_new_n4919_), .Y(u2__abc_52155_new_n11116_));
OR2X2 OR2X2_2043 ( .A(u2__abc_52155_new_n11119_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11120_));
OR2X2 OR2X2_2044 ( .A(u2__abc_52155_new_n11118_), .B(u2__abc_52155_new_n11120_), .Y(u2__abc_52155_new_n11121_));
OR2X2 OR2X2_2045 ( .A(u2__abc_52155_new_n11125_), .B(u2__abc_52155_new_n11111_), .Y(u2__abc_52155_new_n11126_));
OR2X2 OR2X2_2046 ( .A(u2__abc_52155_new_n4908_), .B(u2__abc_52155_new_n4917_), .Y(u2__abc_52155_new_n11129_));
OR2X2 OR2X2_2047 ( .A(u2__abc_52155_new_n11132_), .B(u2__abc_52155_new_n11131_), .Y(u2__abc_52155_new_n11133_));
OR2X2 OR2X2_2048 ( .A(u2__abc_52155_new_n11133_), .B(u2__abc_52155_new_n4897_), .Y(u2__abc_52155_new_n11136_));
OR2X2 OR2X2_2049 ( .A(u2__abc_52155_new_n11139_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11140_));
OR2X2 OR2X2_205 ( .A(aNan), .B(sqrto_178_), .Y(_abc_73687_new_n1136_));
OR2X2 OR2X2_2050 ( .A(u2__abc_52155_new_n11138_), .B(u2__abc_52155_new_n11140_), .Y(u2__abc_52155_new_n11141_));
OR2X2 OR2X2_2051 ( .A(u2__abc_52155_new_n11145_), .B(u2__abc_52155_new_n11128_), .Y(u2__abc_52155_new_n11146_));
OR2X2 OR2X2_2052 ( .A(u2__abc_52155_new_n11153_), .B(u2__abc_52155_new_n11150_), .Y(u2__abc_52155_new_n11154_));
OR2X2 OR2X2_2053 ( .A(u2__abc_52155_new_n11156_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11157_));
OR2X2 OR2X2_2054 ( .A(u2__abc_52155_new_n11155_), .B(u2__abc_52155_new_n11157_), .Y(u2__abc_52155_new_n11158_));
OR2X2 OR2X2_2055 ( .A(u2__abc_52155_new_n11162_), .B(u2__abc_52155_new_n11148_), .Y(u2__abc_52155_new_n11163_));
OR2X2 OR2X2_2056 ( .A(u2__abc_52155_new_n11167_), .B(u2__abc_52155_new_n4902_), .Y(u2__abc_52155_new_n11168_));
OR2X2 OR2X2_2057 ( .A(u2__abc_52155_new_n11169_), .B(u2__abc_52155_new_n4888_), .Y(u2__abc_52155_new_n11172_));
OR2X2 OR2X2_2058 ( .A(u2__abc_52155_new_n11175_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11176_));
OR2X2 OR2X2_2059 ( .A(u2__abc_52155_new_n11174_), .B(u2__abc_52155_new_n11176_), .Y(u2__abc_52155_new_n11177_));
OR2X2 OR2X2_206 ( .A(_abc_73687_new_n753_), .B(\a[102] ), .Y(_abc_73687_new_n1137_));
OR2X2 OR2X2_2060 ( .A(u2__abc_52155_new_n11181_), .B(u2__abc_52155_new_n11165_), .Y(u2__abc_52155_new_n11182_));
OR2X2 OR2X2_2061 ( .A(u2__abc_52155_new_n11189_), .B(u2__abc_52155_new_n11186_), .Y(u2__abc_52155_new_n11190_));
OR2X2 OR2X2_2062 ( .A(u2__abc_52155_new_n11192_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11193_));
OR2X2 OR2X2_2063 ( .A(u2__abc_52155_new_n11191_), .B(u2__abc_52155_new_n11193_), .Y(u2__abc_52155_new_n11194_));
OR2X2 OR2X2_2064 ( .A(u2__abc_52155_new_n11198_), .B(u2__abc_52155_new_n11184_), .Y(u2__abc_52155_new_n11199_));
OR2X2 OR2X2_2065 ( .A(u2__abc_52155_new_n11203_), .B(u2__abc_52155_new_n4879_), .Y(u2__abc_52155_new_n11204_));
OR2X2 OR2X2_2066 ( .A(u2__abc_52155_new_n11205_), .B(u2__abc_52155_new_n4866_), .Y(u2__abc_52155_new_n11208_));
OR2X2 OR2X2_2067 ( .A(u2__abc_52155_new_n11211_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11212_));
OR2X2 OR2X2_2068 ( .A(u2__abc_52155_new_n11210_), .B(u2__abc_52155_new_n11212_), .Y(u2__abc_52155_new_n11213_));
OR2X2 OR2X2_2069 ( .A(u2__abc_52155_new_n11217_), .B(u2__abc_52155_new_n11201_), .Y(u2__abc_52155_new_n11218_));
OR2X2 OR2X2_207 ( .A(aNan), .B(sqrto_179_), .Y(_abc_73687_new_n1139_));
OR2X2 OR2X2_2070 ( .A(u2__abc_52155_new_n11225_), .B(u2__abc_52155_new_n11222_), .Y(u2__abc_52155_new_n11226_));
OR2X2 OR2X2_2071 ( .A(u2__abc_52155_new_n11228_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11229_));
OR2X2 OR2X2_2072 ( .A(u2__abc_52155_new_n11227_), .B(u2__abc_52155_new_n11229_), .Y(u2__abc_52155_new_n11230_));
OR2X2 OR2X2_2073 ( .A(u2__abc_52155_new_n11234_), .B(u2__abc_52155_new_n11220_), .Y(u2__abc_52155_new_n11235_));
OR2X2 OR2X2_2074 ( .A(u2__abc_52155_new_n11166_), .B(u2__abc_52155_new_n4902_), .Y(u2__abc_52155_new_n11238_));
OR2X2 OR2X2_2075 ( .A(u2__abc_52155_new_n11202_), .B(u2__abc_52155_new_n4879_), .Y(u2__abc_52155_new_n11244_));
OR2X2 OR2X2_2076 ( .A(u2__abc_52155_new_n11247_), .B(u2__abc_52155_new_n4868_), .Y(u2__abc_52155_new_n11248_));
OR2X2 OR2X2_2077 ( .A(u2__abc_52155_new_n11246_), .B(u2__abc_52155_new_n11248_), .Y(u2__abc_52155_new_n11249_));
OR2X2 OR2X2_2078 ( .A(u2__abc_52155_new_n11243_), .B(u2__abc_52155_new_n11249_), .Y(u2__abc_52155_new_n11250_));
OR2X2 OR2X2_2079 ( .A(u2__abc_52155_new_n11251_), .B(u2__abc_52155_new_n11250_), .Y(u2__abc_52155_new_n11252_));
OR2X2 OR2X2_208 ( .A(_abc_73687_new_n753_), .B(\a[103] ), .Y(_abc_73687_new_n1140_));
OR2X2 OR2X2_2080 ( .A(u2__abc_52155_new_n11252_), .B(u2__abc_52155_new_n4803_), .Y(u2__abc_52155_new_n11255_));
OR2X2 OR2X2_2081 ( .A(u2__abc_52155_new_n11258_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11259_));
OR2X2 OR2X2_2082 ( .A(u2__abc_52155_new_n11257_), .B(u2__abc_52155_new_n11259_), .Y(u2__abc_52155_new_n11260_));
OR2X2 OR2X2_2083 ( .A(u2__abc_52155_new_n11264_), .B(u2__abc_52155_new_n11237_), .Y(u2__abc_52155_new_n11265_));
OR2X2 OR2X2_2084 ( .A(u2__abc_52155_new_n11272_), .B(u2__abc_52155_new_n11269_), .Y(u2__abc_52155_new_n11273_));
OR2X2 OR2X2_2085 ( .A(u2__abc_52155_new_n11275_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11276_));
OR2X2 OR2X2_2086 ( .A(u2__abc_52155_new_n11274_), .B(u2__abc_52155_new_n11276_), .Y(u2__abc_52155_new_n11277_));
OR2X2 OR2X2_2087 ( .A(u2__abc_52155_new_n11281_), .B(u2__abc_52155_new_n11267_), .Y(u2__abc_52155_new_n11282_));
OR2X2 OR2X2_2088 ( .A(u2__abc_52155_new_n4799_), .B(u2__abc_52155_new_n4808_), .Y(u2__abc_52155_new_n11285_));
OR2X2 OR2X2_2089 ( .A(u2__abc_52155_new_n11288_), .B(u2__abc_52155_new_n11287_), .Y(u2__abc_52155_new_n11289_));
OR2X2 OR2X2_209 ( .A(aNan), .B(sqrto_180_), .Y(_abc_73687_new_n1142_));
OR2X2 OR2X2_2090 ( .A(u2__abc_52155_new_n11289_), .B(u2__abc_52155_new_n4818_), .Y(u2__abc_52155_new_n11292_));
OR2X2 OR2X2_2091 ( .A(u2__abc_52155_new_n11295_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11296_));
OR2X2 OR2X2_2092 ( .A(u2__abc_52155_new_n11294_), .B(u2__abc_52155_new_n11296_), .Y(u2__abc_52155_new_n11297_));
OR2X2 OR2X2_2093 ( .A(u2__abc_52155_new_n11301_), .B(u2__abc_52155_new_n11284_), .Y(u2__abc_52155_new_n11302_));
OR2X2 OR2X2_2094 ( .A(u2__abc_52155_new_n11309_), .B(u2__abc_52155_new_n11306_), .Y(u2__abc_52155_new_n11310_));
OR2X2 OR2X2_2095 ( .A(u2__abc_52155_new_n11312_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11313_));
OR2X2 OR2X2_2096 ( .A(u2__abc_52155_new_n11311_), .B(u2__abc_52155_new_n11313_), .Y(u2__abc_52155_new_n11314_));
OR2X2 OR2X2_2097 ( .A(u2__abc_52155_new_n11318_), .B(u2__abc_52155_new_n11304_), .Y(u2__abc_52155_new_n11319_));
OR2X2 OR2X2_2098 ( .A(u2__abc_52155_new_n11323_), .B(u2__abc_52155_new_n4820_), .Y(u2__abc_52155_new_n11324_));
OR2X2 OR2X2_2099 ( .A(u2__abc_52155_new_n11322_), .B(u2__abc_52155_new_n11324_), .Y(u2__abc_52155_new_n11325_));
OR2X2 OR2X2_21 ( .A(aNan), .B(sqrto_86_), .Y(_abc_73687_new_n860_));
OR2X2 OR2X2_210 ( .A(_abc_73687_new_n753_), .B(\a[104] ), .Y(_abc_73687_new_n1143_));
OR2X2 OR2X2_2100 ( .A(u2__abc_52155_new_n11326_), .B(u2__abc_52155_new_n11325_), .Y(u2__abc_52155_new_n11327_));
OR2X2 OR2X2_2101 ( .A(u2__abc_52155_new_n11327_), .B(u2__abc_52155_new_n4856_), .Y(u2__abc_52155_new_n11330_));
OR2X2 OR2X2_2102 ( .A(u2__abc_52155_new_n11333_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11334_));
OR2X2 OR2X2_2103 ( .A(u2__abc_52155_new_n11332_), .B(u2__abc_52155_new_n11334_), .Y(u2__abc_52155_new_n11335_));
OR2X2 OR2X2_2104 ( .A(u2__abc_52155_new_n11339_), .B(u2__abc_52155_new_n11321_), .Y(u2__abc_52155_new_n11340_));
OR2X2 OR2X2_2105 ( .A(u2__abc_52155_new_n11347_), .B(u2__abc_52155_new_n11344_), .Y(u2__abc_52155_new_n11348_));
OR2X2 OR2X2_2106 ( .A(u2__abc_52155_new_n11350_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11351_));
OR2X2 OR2X2_2107 ( .A(u2__abc_52155_new_n11349_), .B(u2__abc_52155_new_n11351_), .Y(u2__abc_52155_new_n11352_));
OR2X2 OR2X2_2108 ( .A(u2__abc_52155_new_n11356_), .B(u2__abc_52155_new_n11342_), .Y(u2__abc_52155_new_n11357_));
OR2X2 OR2X2_2109 ( .A(u2__abc_52155_new_n11361_), .B(u2__abc_52155_new_n4847_), .Y(u2__abc_52155_new_n11362_));
OR2X2 OR2X2_211 ( .A(aNan), .B(sqrto_181_), .Y(_abc_73687_new_n1145_));
OR2X2 OR2X2_2110 ( .A(u2__abc_52155_new_n11363_), .B(u2__abc_52155_new_n4834_), .Y(u2__abc_52155_new_n11366_));
OR2X2 OR2X2_2111 ( .A(u2__abc_52155_new_n11369_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11370_));
OR2X2 OR2X2_2112 ( .A(u2__abc_52155_new_n11368_), .B(u2__abc_52155_new_n11370_), .Y(u2__abc_52155_new_n11371_));
OR2X2 OR2X2_2113 ( .A(u2__abc_52155_new_n11375_), .B(u2__abc_52155_new_n11359_), .Y(u2__abc_52155_new_n11376_));
OR2X2 OR2X2_2114 ( .A(u2__abc_52155_new_n11383_), .B(u2__abc_52155_new_n11380_), .Y(u2__abc_52155_new_n11384_));
OR2X2 OR2X2_2115 ( .A(u2__abc_52155_new_n11386_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11387_));
OR2X2 OR2X2_2116 ( .A(u2__abc_52155_new_n11385_), .B(u2__abc_52155_new_n11387_), .Y(u2__abc_52155_new_n11388_));
OR2X2 OR2X2_2117 ( .A(u2__abc_52155_new_n11392_), .B(u2__abc_52155_new_n11378_), .Y(u2__abc_52155_new_n11393_));
OR2X2 OR2X2_2118 ( .A(u2__abc_52155_new_n11360_), .B(u2__abc_52155_new_n4847_), .Y(u2__abc_52155_new_n11400_));
OR2X2 OR2X2_2119 ( .A(u2__abc_52155_new_n11403_), .B(u2__abc_52155_new_n4836_), .Y(u2__abc_52155_new_n11404_));
OR2X2 OR2X2_212 ( .A(_abc_73687_new_n753_), .B(\a[105] ), .Y(_abc_73687_new_n1146_));
OR2X2 OR2X2_2120 ( .A(u2__abc_52155_new_n11402_), .B(u2__abc_52155_new_n11404_), .Y(u2__abc_52155_new_n11405_));
OR2X2 OR2X2_2121 ( .A(u2__abc_52155_new_n11399_), .B(u2__abc_52155_new_n11405_), .Y(u2__abc_52155_new_n11406_));
OR2X2 OR2X2_2122 ( .A(u2__abc_52155_new_n11398_), .B(u2__abc_52155_new_n11406_), .Y(u2__abc_52155_new_n11407_));
OR2X2 OR2X2_2123 ( .A(u2__abc_52155_new_n11397_), .B(u2__abc_52155_new_n11407_), .Y(u2__abc_52155_new_n11408_));
OR2X2 OR2X2_2124 ( .A(u2__abc_52155_new_n11396_), .B(u2__abc_52155_new_n11408_), .Y(u2__abc_52155_new_n11409_));
OR2X2 OR2X2_2125 ( .A(u2__abc_52155_new_n11410_), .B(u2__abc_52155_new_n11409_), .Y(u2__abc_52155_new_n11411_));
OR2X2 OR2X2_2126 ( .A(u2__abc_52155_new_n11411_), .B(u2__abc_52155_new_n4783_), .Y(u2__abc_52155_new_n11414_));
OR2X2 OR2X2_2127 ( .A(u2__abc_52155_new_n11417_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11418_));
OR2X2 OR2X2_2128 ( .A(u2__abc_52155_new_n11416_), .B(u2__abc_52155_new_n11418_), .Y(u2__abc_52155_new_n11419_));
OR2X2 OR2X2_2129 ( .A(u2__abc_52155_new_n11423_), .B(u2__abc_52155_new_n11395_), .Y(u2__abc_52155_new_n11424_));
OR2X2 OR2X2_213 ( .A(aNan), .B(sqrto_182_), .Y(_abc_73687_new_n1148_));
OR2X2 OR2X2_2130 ( .A(u2__abc_52155_new_n11430_), .B(u2__abc_52155_new_n11431_), .Y(u2__abc_52155_new_n11432_));
OR2X2 OR2X2_2131 ( .A(u2__abc_52155_new_n11434_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11435_));
OR2X2 OR2X2_2132 ( .A(u2__abc_52155_new_n11433_), .B(u2__abc_52155_new_n11435_), .Y(u2__abc_52155_new_n11436_));
OR2X2 OR2X2_2133 ( .A(u2__abc_52155_new_n11440_), .B(u2__abc_52155_new_n11426_), .Y(u2__abc_52155_new_n11441_));
OR2X2 OR2X2_2134 ( .A(u2__abc_52155_new_n11445_), .B(u2__abc_52155_new_n4785_), .Y(u2__abc_52155_new_n11446_));
OR2X2 OR2X2_2135 ( .A(u2__abc_52155_new_n11446_), .B(u2__abc_52155_new_n11444_), .Y(u2__abc_52155_new_n11449_));
OR2X2 OR2X2_2136 ( .A(u2__abc_52155_new_n11452_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11453_));
OR2X2 OR2X2_2137 ( .A(u2__abc_52155_new_n11451_), .B(u2__abc_52155_new_n11453_), .Y(u2__abc_52155_new_n11454_));
OR2X2 OR2X2_2138 ( .A(u2__abc_52155_new_n11458_), .B(u2__abc_52155_new_n11443_), .Y(u2__abc_52155_new_n11459_));
OR2X2 OR2X2_2139 ( .A(u2__abc_52155_new_n11463_), .B(u2__abc_52155_new_n4774_), .Y(u2__abc_52155_new_n11464_));
OR2X2 OR2X2_214 ( .A(_abc_73687_new_n753_), .B(\a[106] ), .Y(_abc_73687_new_n1149_));
OR2X2 OR2X2_2140 ( .A(u2__abc_52155_new_n11466_), .B(u2__abc_52155_new_n11465_), .Y(u2__abc_52155_new_n11467_));
OR2X2 OR2X2_2141 ( .A(u2__abc_52155_new_n11470_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11471_));
OR2X2 OR2X2_2142 ( .A(u2__abc_52155_new_n11469_), .B(u2__abc_52155_new_n11471_), .Y(u2__abc_52155_new_n11472_));
OR2X2 OR2X2_2143 ( .A(u2__abc_52155_new_n11476_), .B(u2__abc_52155_new_n11461_), .Y(u2__abc_52155_new_n11477_));
OR2X2 OR2X2_2144 ( .A(u2__abc_52155_new_n11480_), .B(u2__abc_52155_new_n4788_), .Y(u2__abc_52155_new_n11481_));
OR2X2 OR2X2_2145 ( .A(u2__abc_52155_new_n11481_), .B(u2__abc_52155_new_n4775_), .Y(u2__abc_52155_new_n11482_));
OR2X2 OR2X2_2146 ( .A(u2__abc_52155_new_n11462_), .B(u2__abc_52155_new_n4773_), .Y(u2__abc_52155_new_n11483_));
OR2X2 OR2X2_2147 ( .A(u2__abc_52155_new_n11487_), .B(u2__abc_52155_new_n11486_), .Y(u2__abc_52155_new_n11488_));
OR2X2 OR2X2_2148 ( .A(u2__abc_52155_new_n11488_), .B(u2__abc_52155_new_n4762_), .Y(u2__abc_52155_new_n11491_));
OR2X2 OR2X2_2149 ( .A(u2__abc_52155_new_n11494_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11495_));
OR2X2 OR2X2_215 ( .A(aNan), .B(sqrto_183_), .Y(_abc_73687_new_n1151_));
OR2X2 OR2X2_2150 ( .A(u2__abc_52155_new_n11493_), .B(u2__abc_52155_new_n11495_), .Y(u2__abc_52155_new_n11496_));
OR2X2 OR2X2_2151 ( .A(u2__abc_52155_new_n11500_), .B(u2__abc_52155_new_n11479_), .Y(u2__abc_52155_new_n11501_));
OR2X2 OR2X2_2152 ( .A(u2__abc_52155_new_n11505_), .B(u2__abc_52155_new_n4755_), .Y(u2__abc_52155_new_n11508_));
OR2X2 OR2X2_2153 ( .A(u2__abc_52155_new_n11511_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11512_));
OR2X2 OR2X2_2154 ( .A(u2__abc_52155_new_n11510_), .B(u2__abc_52155_new_n11512_), .Y(u2__abc_52155_new_n11513_));
OR2X2 OR2X2_2155 ( .A(u2__abc_52155_new_n11517_), .B(u2__abc_52155_new_n11503_), .Y(u2__abc_52155_new_n11518_));
OR2X2 OR2X2_2156 ( .A(u2__abc_52155_new_n11522_), .B(u2__abc_52155_new_n4740_), .Y(u2__abc_52155_new_n11525_));
OR2X2 OR2X2_2157 ( .A(u2__abc_52155_new_n11528_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11529_));
OR2X2 OR2X2_2158 ( .A(u2__abc_52155_new_n11527_), .B(u2__abc_52155_new_n11529_), .Y(u2__abc_52155_new_n11530_));
OR2X2 OR2X2_2159 ( .A(u2__abc_52155_new_n11534_), .B(u2__abc_52155_new_n11520_), .Y(u2__abc_52155_new_n11535_));
OR2X2 OR2X2_216 ( .A(_abc_73687_new_n753_), .B(\a[107] ), .Y(_abc_73687_new_n1152_));
OR2X2 OR2X2_2160 ( .A(u2__abc_52155_new_n11542_), .B(u2__abc_52155_new_n11539_), .Y(u2__abc_52155_new_n11543_));
OR2X2 OR2X2_2161 ( .A(u2__abc_52155_new_n11545_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11546_));
OR2X2 OR2X2_2162 ( .A(u2__abc_52155_new_n11544_), .B(u2__abc_52155_new_n11546_), .Y(u2__abc_52155_new_n11547_));
OR2X2 OR2X2_2163 ( .A(u2__abc_52155_new_n11551_), .B(u2__abc_52155_new_n11537_), .Y(u2__abc_52155_new_n11552_));
OR2X2 OR2X2_2164 ( .A(u2__abc_52155_new_n4750_), .B(u2__abc_52155_new_n4757_), .Y(u2__abc_52155_new_n11556_));
OR2X2 OR2X2_2165 ( .A(u2__abc_52155_new_n11559_), .B(u2__abc_52155_new_n4742_), .Y(u2__abc_52155_new_n11560_));
OR2X2 OR2X2_2166 ( .A(u2__abc_52155_new_n11558_), .B(u2__abc_52155_new_n11560_), .Y(u2__abc_52155_new_n11561_));
OR2X2 OR2X2_2167 ( .A(u2__abc_52155_new_n11555_), .B(u2__abc_52155_new_n11561_), .Y(u2__abc_52155_new_n11562_));
OR2X2 OR2X2_2168 ( .A(u2__abc_52155_new_n11563_), .B(u2__abc_52155_new_n11562_), .Y(u2__abc_52155_new_n11564_));
OR2X2 OR2X2_2169 ( .A(u2__abc_52155_new_n11564_), .B(u2__abc_52155_new_n4699_), .Y(u2__abc_52155_new_n11567_));
OR2X2 OR2X2_217 ( .A(aNan), .B(sqrto_184_), .Y(_abc_73687_new_n1154_));
OR2X2 OR2X2_2170 ( .A(u2__abc_52155_new_n11570_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11571_));
OR2X2 OR2X2_2171 ( .A(u2__abc_52155_new_n11569_), .B(u2__abc_52155_new_n11571_), .Y(u2__abc_52155_new_n11572_));
OR2X2 OR2X2_2172 ( .A(u2__abc_52155_new_n11576_), .B(u2__abc_52155_new_n11554_), .Y(u2__abc_52155_new_n11577_));
OR2X2 OR2X2_2173 ( .A(u2__abc_52155_new_n11584_), .B(u2__abc_52155_new_n11581_), .Y(u2__abc_52155_new_n11585_));
OR2X2 OR2X2_2174 ( .A(u2__abc_52155_new_n11587_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11588_));
OR2X2 OR2X2_2175 ( .A(u2__abc_52155_new_n11586_), .B(u2__abc_52155_new_n11588_), .Y(u2__abc_52155_new_n11589_));
OR2X2 OR2X2_2176 ( .A(u2__abc_52155_new_n11593_), .B(u2__abc_52155_new_n11579_), .Y(u2__abc_52155_new_n11594_));
OR2X2 OR2X2_2177 ( .A(u2__abc_52155_new_n11598_), .B(u2__abc_52155_new_n4690_), .Y(u2__abc_52155_new_n11599_));
OR2X2 OR2X2_2178 ( .A(u2__abc_52155_new_n11600_), .B(u2__abc_52155_new_n4677_), .Y(u2__abc_52155_new_n11603_));
OR2X2 OR2X2_2179 ( .A(u2__abc_52155_new_n11606_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11607_));
OR2X2 OR2X2_218 ( .A(_abc_73687_new_n753_), .B(\a[108] ), .Y(_abc_73687_new_n1155_));
OR2X2 OR2X2_2180 ( .A(u2__abc_52155_new_n11605_), .B(u2__abc_52155_new_n11607_), .Y(u2__abc_52155_new_n11608_));
OR2X2 OR2X2_2181 ( .A(u2__abc_52155_new_n11612_), .B(u2__abc_52155_new_n11596_), .Y(u2__abc_52155_new_n11613_));
OR2X2 OR2X2_2182 ( .A(u2__abc_52155_new_n11620_), .B(u2__abc_52155_new_n11617_), .Y(u2__abc_52155_new_n11621_));
OR2X2 OR2X2_2183 ( .A(u2__abc_52155_new_n11623_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11624_));
OR2X2 OR2X2_2184 ( .A(u2__abc_52155_new_n11622_), .B(u2__abc_52155_new_n11624_), .Y(u2__abc_52155_new_n11625_));
OR2X2 OR2X2_2185 ( .A(u2__abc_52155_new_n11629_), .B(u2__abc_52155_new_n11615_), .Y(u2__abc_52155_new_n11630_));
OR2X2 OR2X2_2186 ( .A(u2__abc_52155_new_n11597_), .B(u2__abc_52155_new_n4690_), .Y(u2__abc_52155_new_n11633_));
OR2X2 OR2X2_2187 ( .A(u2__abc_52155_new_n11636_), .B(u2__abc_52155_new_n4679_), .Y(u2__abc_52155_new_n11637_));
OR2X2 OR2X2_2188 ( .A(u2__abc_52155_new_n11635_), .B(u2__abc_52155_new_n11637_), .Y(u2__abc_52155_new_n11638_));
OR2X2 OR2X2_2189 ( .A(u2__abc_52155_new_n11639_), .B(u2__abc_52155_new_n11638_), .Y(u2__abc_52155_new_n11640_));
OR2X2 OR2X2_219 ( .A(aNan), .B(sqrto_185_), .Y(_abc_73687_new_n1157_));
OR2X2 OR2X2_2190 ( .A(u2__abc_52155_new_n11640_), .B(u2__abc_52155_new_n4730_), .Y(u2__abc_52155_new_n11643_));
OR2X2 OR2X2_2191 ( .A(u2__abc_52155_new_n11646_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11647_));
OR2X2 OR2X2_2192 ( .A(u2__abc_52155_new_n11645_), .B(u2__abc_52155_new_n11647_), .Y(u2__abc_52155_new_n11648_));
OR2X2 OR2X2_2193 ( .A(u2__abc_52155_new_n11652_), .B(u2__abc_52155_new_n11632_), .Y(u2__abc_52155_new_n11653_));
OR2X2 OR2X2_2194 ( .A(u2__abc_52155_new_n11660_), .B(u2__abc_52155_new_n11657_), .Y(u2__abc_52155_new_n11661_));
OR2X2 OR2X2_2195 ( .A(u2__abc_52155_new_n11663_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11664_));
OR2X2 OR2X2_2196 ( .A(u2__abc_52155_new_n11662_), .B(u2__abc_52155_new_n11664_), .Y(u2__abc_52155_new_n11665_));
OR2X2 OR2X2_2197 ( .A(u2__abc_52155_new_n11669_), .B(u2__abc_52155_new_n11655_), .Y(u2__abc_52155_new_n11670_));
OR2X2 OR2X2_2198 ( .A(u2__abc_52155_new_n11674_), .B(u2__abc_52155_new_n4721_), .Y(u2__abc_52155_new_n11675_));
OR2X2 OR2X2_2199 ( .A(u2__abc_52155_new_n11676_), .B(u2__abc_52155_new_n4708_), .Y(u2__abc_52155_new_n11679_));
OR2X2 OR2X2_22 ( .A(_abc_73687_new_n753_), .B(\a[10] ), .Y(_abc_73687_new_n861_));
OR2X2 OR2X2_220 ( .A(_abc_73687_new_n753_), .B(\a[109] ), .Y(_abc_73687_new_n1158_));
OR2X2 OR2X2_2200 ( .A(u2__abc_52155_new_n11682_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11683_));
OR2X2 OR2X2_2201 ( .A(u2__abc_52155_new_n11681_), .B(u2__abc_52155_new_n11683_), .Y(u2__abc_52155_new_n11684_));
OR2X2 OR2X2_2202 ( .A(u2__abc_52155_new_n11688_), .B(u2__abc_52155_new_n11672_), .Y(u2__abc_52155_new_n11689_));
OR2X2 OR2X2_2203 ( .A(u2__abc_52155_new_n11696_), .B(u2__abc_52155_new_n11693_), .Y(u2__abc_52155_new_n11697_));
OR2X2 OR2X2_2204 ( .A(u2__abc_52155_new_n11699_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11700_));
OR2X2 OR2X2_2205 ( .A(u2__abc_52155_new_n11698_), .B(u2__abc_52155_new_n11700_), .Y(u2__abc_52155_new_n11701_));
OR2X2 OR2X2_2206 ( .A(u2__abc_52155_new_n11705_), .B(u2__abc_52155_new_n11691_), .Y(u2__abc_52155_new_n11706_));
OR2X2 OR2X2_2207 ( .A(u2__abc_52155_new_n11673_), .B(u2__abc_52155_new_n4721_), .Y(u2__abc_52155_new_n11711_));
OR2X2 OR2X2_2208 ( .A(u2__abc_52155_new_n11714_), .B(u2__abc_52155_new_n4710_), .Y(u2__abc_52155_new_n11715_));
OR2X2 OR2X2_2209 ( .A(u2__abc_52155_new_n11713_), .B(u2__abc_52155_new_n11715_), .Y(u2__abc_52155_new_n11716_));
OR2X2 OR2X2_221 ( .A(aNan), .B(sqrto_186_), .Y(_abc_73687_new_n1160_));
OR2X2 OR2X2_2210 ( .A(u2__abc_52155_new_n11710_), .B(u2__abc_52155_new_n11716_), .Y(u2__abc_52155_new_n11717_));
OR2X2 OR2X2_2211 ( .A(u2__abc_52155_new_n11709_), .B(u2__abc_52155_new_n11717_), .Y(u2__abc_52155_new_n11718_));
OR2X2 OR2X2_2212 ( .A(u2__abc_52155_new_n11719_), .B(u2__abc_52155_new_n11718_), .Y(u2__abc_52155_new_n11720_));
OR2X2 OR2X2_2213 ( .A(u2__abc_52155_new_n11720_), .B(u2__abc_52155_new_n4628_), .Y(u2__abc_52155_new_n11723_));
OR2X2 OR2X2_2214 ( .A(u2__abc_52155_new_n11726_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11727_));
OR2X2 OR2X2_2215 ( .A(u2__abc_52155_new_n11725_), .B(u2__abc_52155_new_n11727_), .Y(u2__abc_52155_new_n11728_));
OR2X2 OR2X2_2216 ( .A(u2__abc_52155_new_n11732_), .B(u2__abc_52155_new_n11708_), .Y(u2__abc_52155_new_n11733_));
OR2X2 OR2X2_2217 ( .A(u2__abc_52155_new_n11739_), .B(u2__abc_52155_new_n11740_), .Y(u2__abc_52155_new_n11741_));
OR2X2 OR2X2_2218 ( .A(u2__abc_52155_new_n11743_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11744_));
OR2X2 OR2X2_2219 ( .A(u2__abc_52155_new_n11742_), .B(u2__abc_52155_new_n11744_), .Y(u2__abc_52155_new_n11745_));
OR2X2 OR2X2_222 ( .A(_abc_73687_new_n753_), .B(\a[110] ), .Y(_abc_73687_new_n1161_));
OR2X2 OR2X2_2220 ( .A(u2__abc_52155_new_n11749_), .B(u2__abc_52155_new_n11735_), .Y(u2__abc_52155_new_n11750_));
OR2X2 OR2X2_2221 ( .A(u2__abc_52155_new_n11753_), .B(u2__abc_52155_new_n4633_), .Y(u2__abc_52155_new_n11754_));
OR2X2 OR2X2_2222 ( .A(u2__abc_52155_new_n11756_), .B(u2__abc_52155_new_n11755_), .Y(u2__abc_52155_new_n11757_));
OR2X2 OR2X2_2223 ( .A(u2__abc_52155_new_n11757_), .B(u2__abc_52155_new_n4613_), .Y(u2__abc_52155_new_n11760_));
OR2X2 OR2X2_2224 ( .A(u2__abc_52155_new_n11763_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11764_));
OR2X2 OR2X2_2225 ( .A(u2__abc_52155_new_n11762_), .B(u2__abc_52155_new_n11764_), .Y(u2__abc_52155_new_n11765_));
OR2X2 OR2X2_2226 ( .A(u2__abc_52155_new_n11769_), .B(u2__abc_52155_new_n11752_), .Y(u2__abc_52155_new_n11770_));
OR2X2 OR2X2_2227 ( .A(u2__abc_52155_new_n11777_), .B(u2__abc_52155_new_n11774_), .Y(u2__abc_52155_new_n11778_));
OR2X2 OR2X2_2228 ( .A(u2__abc_52155_new_n11780_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11781_));
OR2X2 OR2X2_2229 ( .A(u2__abc_52155_new_n11779_), .B(u2__abc_52155_new_n11781_), .Y(u2__abc_52155_new_n11782_));
OR2X2 OR2X2_223 ( .A(aNan), .B(sqrto_187_), .Y(_abc_73687_new_n1163_));
OR2X2 OR2X2_2230 ( .A(u2__abc_52155_new_n11786_), .B(u2__abc_52155_new_n11772_), .Y(u2__abc_52155_new_n11787_));
OR2X2 OR2X2_2231 ( .A(u2__abc_52155_new_n11791_), .B(u2__abc_52155_new_n4615_), .Y(u2__abc_52155_new_n11792_));
OR2X2 OR2X2_2232 ( .A(u2__abc_52155_new_n11790_), .B(u2__abc_52155_new_n11792_), .Y(u2__abc_52155_new_n11793_));
OR2X2 OR2X2_2233 ( .A(u2__abc_52155_new_n11794_), .B(u2__abc_52155_new_n11793_), .Y(u2__abc_52155_new_n11795_));
OR2X2 OR2X2_2234 ( .A(u2__abc_52155_new_n11795_), .B(u2__abc_52155_new_n4666_), .Y(u2__abc_52155_new_n11798_));
OR2X2 OR2X2_2235 ( .A(u2__abc_52155_new_n11801_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11802_));
OR2X2 OR2X2_2236 ( .A(u2__abc_52155_new_n11800_), .B(u2__abc_52155_new_n11802_), .Y(u2__abc_52155_new_n11803_));
OR2X2 OR2X2_2237 ( .A(u2__abc_52155_new_n11807_), .B(u2__abc_52155_new_n11789_), .Y(u2__abc_52155_new_n11808_));
OR2X2 OR2X2_2238 ( .A(u2__abc_52155_new_n11812_), .B(u2__abc_52155_new_n4659_), .Y(u2__abc_52155_new_n11815_));
OR2X2 OR2X2_2239 ( .A(u2__abc_52155_new_n11818_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11819_));
OR2X2 OR2X2_224 ( .A(_abc_73687_new_n753_), .B(\a[111] ), .Y(_abc_73687_new_n1164_));
OR2X2 OR2X2_2240 ( .A(u2__abc_52155_new_n11817_), .B(u2__abc_52155_new_n11819_), .Y(u2__abc_52155_new_n11820_));
OR2X2 OR2X2_2241 ( .A(u2__abc_52155_new_n11824_), .B(u2__abc_52155_new_n11810_), .Y(u2__abc_52155_new_n11825_));
OR2X2 OR2X2_2242 ( .A(u2__abc_52155_new_n11829_), .B(u2__abc_52155_new_n4644_), .Y(u2__abc_52155_new_n11832_));
OR2X2 OR2X2_2243 ( .A(u2__abc_52155_new_n11835_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11836_));
OR2X2 OR2X2_2244 ( .A(u2__abc_52155_new_n11834_), .B(u2__abc_52155_new_n11836_), .Y(u2__abc_52155_new_n11837_));
OR2X2 OR2X2_2245 ( .A(u2__abc_52155_new_n11841_), .B(u2__abc_52155_new_n11827_), .Y(u2__abc_52155_new_n11842_));
OR2X2 OR2X2_2246 ( .A(u2__abc_52155_new_n11849_), .B(u2__abc_52155_new_n11846_), .Y(u2__abc_52155_new_n11850_));
OR2X2 OR2X2_2247 ( .A(u2__abc_52155_new_n11852_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11853_));
OR2X2 OR2X2_2248 ( .A(u2__abc_52155_new_n11851_), .B(u2__abc_52155_new_n11853_), .Y(u2__abc_52155_new_n11854_));
OR2X2 OR2X2_2249 ( .A(u2__abc_52155_new_n11858_), .B(u2__abc_52155_new_n11844_), .Y(u2__abc_52155_new_n11859_));
OR2X2 OR2X2_225 ( .A(aNan), .B(sqrto_188_), .Y(\o[224] ));
OR2X2 OR2X2_2250 ( .A(u2__abc_52155_new_n4654_), .B(u2__abc_52155_new_n4661_), .Y(u2__abc_52155_new_n11863_));
OR2X2 OR2X2_2251 ( .A(u2__abc_52155_new_n11866_), .B(u2__abc_52155_new_n4646_), .Y(u2__abc_52155_new_n11867_));
OR2X2 OR2X2_2252 ( .A(u2__abc_52155_new_n11865_), .B(u2__abc_52155_new_n11867_), .Y(u2__abc_52155_new_n11868_));
OR2X2 OR2X2_2253 ( .A(u2__abc_52155_new_n11862_), .B(u2__abc_52155_new_n11868_), .Y(u2__abc_52155_new_n11869_));
OR2X2 OR2X2_2254 ( .A(u2__abc_52155_new_n11870_), .B(u2__abc_52155_new_n11869_), .Y(u2__abc_52155_new_n11871_));
OR2X2 OR2X2_2255 ( .A(u2__abc_52155_new_n11871_), .B(u2__abc_52155_new_n4565_), .Y(u2__abc_52155_new_n11874_));
OR2X2 OR2X2_2256 ( .A(u2__abc_52155_new_n11877_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11878_));
OR2X2 OR2X2_2257 ( .A(u2__abc_52155_new_n11876_), .B(u2__abc_52155_new_n11878_), .Y(u2__abc_52155_new_n11879_));
OR2X2 OR2X2_2258 ( .A(u2__abc_52155_new_n11883_), .B(u2__abc_52155_new_n11861_), .Y(u2__abc_52155_new_n11884_));
OR2X2 OR2X2_2259 ( .A(u2__abc_52155_new_n11890_), .B(u2__abc_52155_new_n11891_), .Y(u2__abc_52155_new_n11892_));
OR2X2 OR2X2_226 ( .A(\a[112] ), .B(\a[0] ), .Y(_abc_73687_new_n1169_));
OR2X2 OR2X2_2260 ( .A(u2__abc_52155_new_n11894_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11895_));
OR2X2 OR2X2_2261 ( .A(u2__abc_52155_new_n11893_), .B(u2__abc_52155_new_n11895_), .Y(u2__abc_52155_new_n11896_));
OR2X2 OR2X2_2262 ( .A(u2__abc_52155_new_n11900_), .B(u2__abc_52155_new_n11886_), .Y(u2__abc_52155_new_n11901_));
OR2X2 OR2X2_2263 ( .A(u2__abc_52155_new_n11904_), .B(u2__abc_52155_new_n4570_), .Y(u2__abc_52155_new_n11905_));
OR2X2 OR2X2_2264 ( .A(u2__abc_52155_new_n11907_), .B(u2__abc_52155_new_n11906_), .Y(u2__abc_52155_new_n11908_));
OR2X2 OR2X2_2265 ( .A(u2__abc_52155_new_n11908_), .B(u2__abc_52155_new_n4550_), .Y(u2__abc_52155_new_n11911_));
OR2X2 OR2X2_2266 ( .A(u2__abc_52155_new_n11914_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11915_));
OR2X2 OR2X2_2267 ( .A(u2__abc_52155_new_n11913_), .B(u2__abc_52155_new_n11915_), .Y(u2__abc_52155_new_n11916_));
OR2X2 OR2X2_2268 ( .A(u2__abc_52155_new_n11920_), .B(u2__abc_52155_new_n11903_), .Y(u2__abc_52155_new_n11921_));
OR2X2 OR2X2_2269 ( .A(u2__abc_52155_new_n11928_), .B(u2__abc_52155_new_n11925_), .Y(u2__abc_52155_new_n11929_));
OR2X2 OR2X2_227 ( .A(_abc_73687_new_n1170_), .B(\a[1] ), .Y(_abc_73687_new_n1171_));
OR2X2 OR2X2_2270 ( .A(u2__abc_52155_new_n11931_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11932_));
OR2X2 OR2X2_2271 ( .A(u2__abc_52155_new_n11930_), .B(u2__abc_52155_new_n11932_), .Y(u2__abc_52155_new_n11933_));
OR2X2 OR2X2_2272 ( .A(u2__abc_52155_new_n11937_), .B(u2__abc_52155_new_n11923_), .Y(u2__abc_52155_new_n11938_));
OR2X2 OR2X2_2273 ( .A(u2__abc_52155_new_n11942_), .B(u2__abc_52155_new_n4552_), .Y(u2__abc_52155_new_n11943_));
OR2X2 OR2X2_2274 ( .A(u2__abc_52155_new_n11941_), .B(u2__abc_52155_new_n11943_), .Y(u2__abc_52155_new_n11944_));
OR2X2 OR2X2_2275 ( .A(u2__abc_52155_new_n11945_), .B(u2__abc_52155_new_n11944_), .Y(u2__abc_52155_new_n11946_));
OR2X2 OR2X2_2276 ( .A(u2__abc_52155_new_n11946_), .B(u2__abc_52155_new_n4603_), .Y(u2__abc_52155_new_n11949_));
OR2X2 OR2X2_2277 ( .A(u2__abc_52155_new_n11952_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11953_));
OR2X2 OR2X2_2278 ( .A(u2__abc_52155_new_n11951_), .B(u2__abc_52155_new_n11953_), .Y(u2__abc_52155_new_n11954_));
OR2X2 OR2X2_2279 ( .A(u2__abc_52155_new_n11958_), .B(u2__abc_52155_new_n11940_), .Y(u2__abc_52155_new_n11959_));
OR2X2 OR2X2_228 ( .A(\a[112] ), .B(\a[1] ), .Y(_abc_73687_new_n1173_));
OR2X2 OR2X2_2280 ( .A(u2__abc_52155_new_n11966_), .B(u2__abc_52155_new_n11963_), .Y(u2__abc_52155_new_n11967_));
OR2X2 OR2X2_2281 ( .A(u2__abc_52155_new_n11969_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11970_));
OR2X2 OR2X2_2282 ( .A(u2__abc_52155_new_n11968_), .B(u2__abc_52155_new_n11970_), .Y(u2__abc_52155_new_n11971_));
OR2X2 OR2X2_2283 ( .A(u2__abc_52155_new_n11975_), .B(u2__abc_52155_new_n11961_), .Y(u2__abc_52155_new_n11976_));
OR2X2 OR2X2_2284 ( .A(u2__abc_52155_new_n11980_), .B(u2__abc_52155_new_n4594_), .Y(u2__abc_52155_new_n11981_));
OR2X2 OR2X2_2285 ( .A(u2__abc_52155_new_n11982_), .B(u2__abc_52155_new_n4581_), .Y(u2__abc_52155_new_n11985_));
OR2X2 OR2X2_2286 ( .A(u2__abc_52155_new_n11988_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n11989_));
OR2X2 OR2X2_2287 ( .A(u2__abc_52155_new_n11987_), .B(u2__abc_52155_new_n11989_), .Y(u2__abc_52155_new_n11990_));
OR2X2 OR2X2_2288 ( .A(u2__abc_52155_new_n11994_), .B(u2__abc_52155_new_n11978_), .Y(u2__abc_52155_new_n11995_));
OR2X2 OR2X2_2289 ( .A(u2__abc_52155_new_n12002_), .B(u2__abc_52155_new_n11999_), .Y(u2__abc_52155_new_n12003_));
OR2X2 OR2X2_229 ( .A(_abc_73687_new_n1170_), .B(\a[2] ), .Y(_abc_73687_new_n1174_));
OR2X2 OR2X2_2290 ( .A(u2__abc_52155_new_n12005_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12006_));
OR2X2 OR2X2_2291 ( .A(u2__abc_52155_new_n12004_), .B(u2__abc_52155_new_n12006_), .Y(u2__abc_52155_new_n12007_));
OR2X2 OR2X2_2292 ( .A(u2__abc_52155_new_n12011_), .B(u2__abc_52155_new_n11997_), .Y(u2__abc_52155_new_n12012_));
OR2X2 OR2X2_2293 ( .A(u2__abc_52155_new_n12021_), .B(u2__abc_52155_new_n4586_), .Y(u2__abc_52155_new_n12022_));
OR2X2 OR2X2_2294 ( .A(u2__abc_52155_new_n11979_), .B(u2__abc_52155_new_n4594_), .Y(u2__abc_52155_new_n12023_));
OR2X2 OR2X2_2295 ( .A(u2__abc_52155_new_n12032_), .B(u2__abc_52155_new_n12031_), .Y(u2__abc_52155_new_n12033_));
OR2X2 OR2X2_2296 ( .A(u2__abc_52155_new_n12033_), .B(u2__abc_52155_new_n4507_), .Y(u2__abc_52155_new_n12036_));
OR2X2 OR2X2_2297 ( .A(u2__abc_52155_new_n12039_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12040_));
OR2X2 OR2X2_2298 ( .A(u2__abc_52155_new_n12038_), .B(u2__abc_52155_new_n12040_), .Y(u2__abc_52155_new_n12041_));
OR2X2 OR2X2_2299 ( .A(u2__abc_52155_new_n12045_), .B(u2__abc_52155_new_n12014_), .Y(u2__abc_52155_new_n12046_));
OR2X2 OR2X2_23 ( .A(aNan), .B(sqrto_87_), .Y(_abc_73687_new_n863_));
OR2X2 OR2X2_230 ( .A(\a[112] ), .B(\a[2] ), .Y(_abc_73687_new_n1176_));
OR2X2 OR2X2_2300 ( .A(u2__abc_52155_new_n12053_), .B(u2__abc_52155_new_n12050_), .Y(u2__abc_52155_new_n12054_));
OR2X2 OR2X2_2301 ( .A(u2__abc_52155_new_n12056_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12057_));
OR2X2 OR2X2_2302 ( .A(u2__abc_52155_new_n12055_), .B(u2__abc_52155_new_n12057_), .Y(u2__abc_52155_new_n12058_));
OR2X2 OR2X2_2303 ( .A(u2__abc_52155_new_n12062_), .B(u2__abc_52155_new_n12048_), .Y(u2__abc_52155_new_n12063_));
OR2X2 OR2X2_2304 ( .A(u2__abc_52155_new_n12067_), .B(u2__abc_52155_new_n4498_), .Y(u2__abc_52155_new_n12068_));
OR2X2 OR2X2_2305 ( .A(u2__abc_52155_new_n12069_), .B(u2__abc_52155_new_n4485_), .Y(u2__abc_52155_new_n12072_));
OR2X2 OR2X2_2306 ( .A(u2__abc_52155_new_n12075_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12076_));
OR2X2 OR2X2_2307 ( .A(u2__abc_52155_new_n12074_), .B(u2__abc_52155_new_n12076_), .Y(u2__abc_52155_new_n12077_));
OR2X2 OR2X2_2308 ( .A(u2__abc_52155_new_n12081_), .B(u2__abc_52155_new_n12065_), .Y(u2__abc_52155_new_n12082_));
OR2X2 OR2X2_2309 ( .A(u2__abc_52155_new_n12089_), .B(u2__abc_52155_new_n12086_), .Y(u2__abc_52155_new_n12090_));
OR2X2 OR2X2_231 ( .A(_abc_73687_new_n1170_), .B(\a[3] ), .Y(_abc_73687_new_n1177_));
OR2X2 OR2X2_2310 ( .A(u2__abc_52155_new_n12092_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12093_));
OR2X2 OR2X2_2311 ( .A(u2__abc_52155_new_n12091_), .B(u2__abc_52155_new_n12093_), .Y(u2__abc_52155_new_n12094_));
OR2X2 OR2X2_2312 ( .A(u2__abc_52155_new_n12098_), .B(u2__abc_52155_new_n12084_), .Y(u2__abc_52155_new_n12099_));
OR2X2 OR2X2_2313 ( .A(u2__abc_52155_new_n12102_), .B(u2__abc_52155_new_n4490_), .Y(u2__abc_52155_new_n12103_));
OR2X2 OR2X2_2314 ( .A(u2__abc_52155_new_n12066_), .B(u2__abc_52155_new_n4498_), .Y(u2__abc_52155_new_n12104_));
OR2X2 OR2X2_2315 ( .A(u2__abc_52155_new_n12110_), .B(u2__abc_52155_new_n12109_), .Y(u2__abc_52155_new_n12111_));
OR2X2 OR2X2_2316 ( .A(u2__abc_52155_new_n12111_), .B(u2__abc_52155_new_n4538_), .Y(u2__abc_52155_new_n12114_));
OR2X2 OR2X2_2317 ( .A(u2__abc_52155_new_n12117_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12118_));
OR2X2 OR2X2_2318 ( .A(u2__abc_52155_new_n12116_), .B(u2__abc_52155_new_n12118_), .Y(u2__abc_52155_new_n12119_));
OR2X2 OR2X2_2319 ( .A(u2__abc_52155_new_n12123_), .B(u2__abc_52155_new_n12101_), .Y(u2__abc_52155_new_n12124_));
OR2X2 OR2X2_232 ( .A(\a[112] ), .B(\a[3] ), .Y(_abc_73687_new_n1179_));
OR2X2 OR2X2_2320 ( .A(u2__abc_52155_new_n12131_), .B(u2__abc_52155_new_n12128_), .Y(u2__abc_52155_new_n12132_));
OR2X2 OR2X2_2321 ( .A(u2__abc_52155_new_n12134_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12135_));
OR2X2 OR2X2_2322 ( .A(u2__abc_52155_new_n12133_), .B(u2__abc_52155_new_n12135_), .Y(u2__abc_52155_new_n12136_));
OR2X2 OR2X2_2323 ( .A(u2__abc_52155_new_n12140_), .B(u2__abc_52155_new_n12126_), .Y(u2__abc_52155_new_n12141_));
OR2X2 OR2X2_2324 ( .A(u2__abc_52155_new_n12145_), .B(u2__abc_52155_new_n4529_), .Y(u2__abc_52155_new_n12146_));
OR2X2 OR2X2_2325 ( .A(u2__abc_52155_new_n12147_), .B(u2__abc_52155_new_n4516_), .Y(u2__abc_52155_new_n12150_));
OR2X2 OR2X2_2326 ( .A(u2__abc_52155_new_n12153_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12154_));
OR2X2 OR2X2_2327 ( .A(u2__abc_52155_new_n12152_), .B(u2__abc_52155_new_n12154_), .Y(u2__abc_52155_new_n12155_));
OR2X2 OR2X2_2328 ( .A(u2__abc_52155_new_n12159_), .B(u2__abc_52155_new_n12143_), .Y(u2__abc_52155_new_n12160_));
OR2X2 OR2X2_2329 ( .A(u2__abc_52155_new_n12167_), .B(u2__abc_52155_new_n12164_), .Y(u2__abc_52155_new_n12168_));
OR2X2 OR2X2_233 ( .A(_abc_73687_new_n1170_), .B(\a[4] ), .Y(_abc_73687_new_n1180_));
OR2X2 OR2X2_2330 ( .A(u2__abc_52155_new_n12170_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12171_));
OR2X2 OR2X2_2331 ( .A(u2__abc_52155_new_n12169_), .B(u2__abc_52155_new_n12171_), .Y(u2__abc_52155_new_n12172_));
OR2X2 OR2X2_2332 ( .A(u2__abc_52155_new_n12176_), .B(u2__abc_52155_new_n12162_), .Y(u2__abc_52155_new_n12177_));
OR2X2 OR2X2_2333 ( .A(u2__abc_52155_new_n12144_), .B(u2__abc_52155_new_n4529_), .Y(u2__abc_52155_new_n12181_));
OR2X2 OR2X2_2334 ( .A(u2__abc_52155_new_n12184_), .B(u2__abc_52155_new_n4518_), .Y(u2__abc_52155_new_n12185_));
OR2X2 OR2X2_2335 ( .A(u2__abc_52155_new_n12183_), .B(u2__abc_52155_new_n12185_), .Y(u2__abc_52155_new_n12186_));
OR2X2 OR2X2_2336 ( .A(u2__abc_52155_new_n12180_), .B(u2__abc_52155_new_n12186_), .Y(u2__abc_52155_new_n12187_));
OR2X2 OR2X2_2337 ( .A(u2__abc_52155_new_n12188_), .B(u2__abc_52155_new_n12187_), .Y(u2__abc_52155_new_n12189_));
OR2X2 OR2X2_2338 ( .A(u2__abc_52155_new_n12189_), .B(u2__abc_52155_new_n4475_), .Y(u2__abc_52155_new_n12192_));
OR2X2 OR2X2_2339 ( .A(u2__abc_52155_new_n12195_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12196_));
OR2X2 OR2X2_234 ( .A(\a[112] ), .B(\a[4] ), .Y(_abc_73687_new_n1182_));
OR2X2 OR2X2_2340 ( .A(u2__abc_52155_new_n12194_), .B(u2__abc_52155_new_n12196_), .Y(u2__abc_52155_new_n12197_));
OR2X2 OR2X2_2341 ( .A(u2__abc_52155_new_n12201_), .B(u2__abc_52155_new_n12179_), .Y(u2__abc_52155_new_n12202_));
OR2X2 OR2X2_2342 ( .A(u2__abc_52155_new_n12208_), .B(u2__abc_52155_new_n12209_), .Y(u2__abc_52155_new_n12210_));
OR2X2 OR2X2_2343 ( .A(u2__abc_52155_new_n12212_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12213_));
OR2X2 OR2X2_2344 ( .A(u2__abc_52155_new_n12211_), .B(u2__abc_52155_new_n12213_), .Y(u2__abc_52155_new_n12214_));
OR2X2 OR2X2_2345 ( .A(u2__abc_52155_new_n12218_), .B(u2__abc_52155_new_n12204_), .Y(u2__abc_52155_new_n12219_));
OR2X2 OR2X2_2346 ( .A(u2__abc_52155_new_n12222_), .B(u2__abc_52155_new_n4466_), .Y(u2__abc_52155_new_n12223_));
OR2X2 OR2X2_2347 ( .A(u2__abc_52155_new_n12225_), .B(u2__abc_52155_new_n12224_), .Y(u2__abc_52155_new_n12226_));
OR2X2 OR2X2_2348 ( .A(u2__abc_52155_new_n12226_), .B(u2__abc_52155_new_n4453_), .Y(u2__abc_52155_new_n12229_));
OR2X2 OR2X2_2349 ( .A(u2__abc_52155_new_n12232_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12233_));
OR2X2 OR2X2_235 ( .A(_abc_73687_new_n1170_), .B(\a[5] ), .Y(_abc_73687_new_n1183_));
OR2X2 OR2X2_2350 ( .A(u2__abc_52155_new_n12231_), .B(u2__abc_52155_new_n12233_), .Y(u2__abc_52155_new_n12234_));
OR2X2 OR2X2_2351 ( .A(u2__abc_52155_new_n12238_), .B(u2__abc_52155_new_n12221_), .Y(u2__abc_52155_new_n12239_));
OR2X2 OR2X2_2352 ( .A(u2__abc_52155_new_n12246_), .B(u2__abc_52155_new_n12243_), .Y(u2__abc_52155_new_n12247_));
OR2X2 OR2X2_2353 ( .A(u2__abc_52155_new_n12249_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12250_));
OR2X2 OR2X2_2354 ( .A(u2__abc_52155_new_n12248_), .B(u2__abc_52155_new_n12250_), .Y(u2__abc_52155_new_n12251_));
OR2X2 OR2X2_2355 ( .A(u2__abc_52155_new_n12255_), .B(u2__abc_52155_new_n12241_), .Y(u2__abc_52155_new_n12256_));
OR2X2 OR2X2_2356 ( .A(u2__abc_52155_new_n12260_), .B(u2__abc_52155_new_n4458_), .Y(u2__abc_52155_new_n12261_));
OR2X2 OR2X2_2357 ( .A(u2__abc_52155_new_n12262_), .B(u2__abc_52155_new_n4444_), .Y(u2__abc_52155_new_n12265_));
OR2X2 OR2X2_2358 ( .A(u2__abc_52155_new_n12268_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12269_));
OR2X2 OR2X2_2359 ( .A(u2__abc_52155_new_n12267_), .B(u2__abc_52155_new_n12269_), .Y(u2__abc_52155_new_n12270_));
OR2X2 OR2X2_236 ( .A(\a[112] ), .B(\a[5] ), .Y(_abc_73687_new_n1185_));
OR2X2 OR2X2_2360 ( .A(u2__abc_52155_new_n12274_), .B(u2__abc_52155_new_n12258_), .Y(u2__abc_52155_new_n12275_));
OR2X2 OR2X2_2361 ( .A(u2__abc_52155_new_n12282_), .B(u2__abc_52155_new_n12279_), .Y(u2__abc_52155_new_n12283_));
OR2X2 OR2X2_2362 ( .A(u2__abc_52155_new_n12285_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12286_));
OR2X2 OR2X2_2363 ( .A(u2__abc_52155_new_n12284_), .B(u2__abc_52155_new_n12286_), .Y(u2__abc_52155_new_n12287_));
OR2X2 OR2X2_2364 ( .A(u2__abc_52155_new_n12291_), .B(u2__abc_52155_new_n12277_), .Y(u2__abc_52155_new_n12292_));
OR2X2 OR2X2_2365 ( .A(u2__abc_52155_new_n12296_), .B(u2__abc_52155_new_n4435_), .Y(u2__abc_52155_new_n12297_));
OR2X2 OR2X2_2366 ( .A(u2__abc_52155_new_n12298_), .B(u2__abc_52155_new_n4422_), .Y(u2__abc_52155_new_n12301_));
OR2X2 OR2X2_2367 ( .A(u2__abc_52155_new_n12304_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12305_));
OR2X2 OR2X2_2368 ( .A(u2__abc_52155_new_n12303_), .B(u2__abc_52155_new_n12305_), .Y(u2__abc_52155_new_n12306_));
OR2X2 OR2X2_2369 ( .A(u2__abc_52155_new_n12310_), .B(u2__abc_52155_new_n12294_), .Y(u2__abc_52155_new_n12311_));
OR2X2 OR2X2_237 ( .A(_abc_73687_new_n1170_), .B(\a[6] ), .Y(_abc_73687_new_n1186_));
OR2X2 OR2X2_2370 ( .A(u2__abc_52155_new_n12318_), .B(u2__abc_52155_new_n12315_), .Y(u2__abc_52155_new_n12319_));
OR2X2 OR2X2_2371 ( .A(u2__abc_52155_new_n12321_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12322_));
OR2X2 OR2X2_2372 ( .A(u2__abc_52155_new_n12320_), .B(u2__abc_52155_new_n12322_), .Y(u2__abc_52155_new_n12323_));
OR2X2 OR2X2_2373 ( .A(u2__abc_52155_new_n12327_), .B(u2__abc_52155_new_n12313_), .Y(u2__abc_52155_new_n12328_));
OR2X2 OR2X2_2374 ( .A(u2__abc_52155_new_n12259_), .B(u2__abc_52155_new_n4458_), .Y(u2__abc_52155_new_n12333_));
OR2X2 OR2X2_2375 ( .A(u2__abc_52155_new_n12340_), .B(u2__abc_52155_new_n4427_), .Y(u2__abc_52155_new_n12341_));
OR2X2 OR2X2_2376 ( .A(u2__abc_52155_new_n12295_), .B(u2__abc_52155_new_n4435_), .Y(u2__abc_52155_new_n12342_));
OR2X2 OR2X2_2377 ( .A(u2__abc_52155_new_n12350_), .B(u2__abc_52155_new_n12349_), .Y(u2__abc_52155_new_n12351_));
OR2X2 OR2X2_2378 ( .A(u2__abc_52155_new_n12351_), .B(u2__abc_52155_new_n4358_), .Y(u2__abc_52155_new_n12354_));
OR2X2 OR2X2_2379 ( .A(u2__abc_52155_new_n12357_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12358_));
OR2X2 OR2X2_238 ( .A(\a[112] ), .B(\a[6] ), .Y(_abc_73687_new_n1188_));
OR2X2 OR2X2_2380 ( .A(u2__abc_52155_new_n12356_), .B(u2__abc_52155_new_n12358_), .Y(u2__abc_52155_new_n12359_));
OR2X2 OR2X2_2381 ( .A(u2__abc_52155_new_n12363_), .B(u2__abc_52155_new_n12330_), .Y(u2__abc_52155_new_n12364_));
OR2X2 OR2X2_2382 ( .A(u2__abc_52155_new_n12371_), .B(u2__abc_52155_new_n12368_), .Y(u2__abc_52155_new_n12372_));
OR2X2 OR2X2_2383 ( .A(u2__abc_52155_new_n12374_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12375_));
OR2X2 OR2X2_2384 ( .A(u2__abc_52155_new_n12373_), .B(u2__abc_52155_new_n12375_), .Y(u2__abc_52155_new_n12376_));
OR2X2 OR2X2_2385 ( .A(u2__abc_52155_new_n12380_), .B(u2__abc_52155_new_n12366_), .Y(u2__abc_52155_new_n12381_));
OR2X2 OR2X2_2386 ( .A(u2__abc_52155_new_n4354_), .B(u2__abc_52155_new_n4363_), .Y(u2__abc_52155_new_n12384_));
OR2X2 OR2X2_2387 ( .A(u2__abc_52155_new_n12387_), .B(u2__abc_52155_new_n12386_), .Y(u2__abc_52155_new_n12388_));
OR2X2 OR2X2_2388 ( .A(u2__abc_52155_new_n12388_), .B(u2__abc_52155_new_n4373_), .Y(u2__abc_52155_new_n12391_));
OR2X2 OR2X2_2389 ( .A(u2__abc_52155_new_n12394_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12395_));
OR2X2 OR2X2_239 ( .A(_abc_73687_new_n1170_), .B(\a[7] ), .Y(_abc_73687_new_n1189_));
OR2X2 OR2X2_2390 ( .A(u2__abc_52155_new_n12393_), .B(u2__abc_52155_new_n12395_), .Y(u2__abc_52155_new_n12396_));
OR2X2 OR2X2_2391 ( .A(u2__abc_52155_new_n12400_), .B(u2__abc_52155_new_n12383_), .Y(u2__abc_52155_new_n12401_));
OR2X2 OR2X2_2392 ( .A(u2__abc_52155_new_n12408_), .B(u2__abc_52155_new_n12405_), .Y(u2__abc_52155_new_n12409_));
OR2X2 OR2X2_2393 ( .A(u2__abc_52155_new_n12411_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12412_));
OR2X2 OR2X2_2394 ( .A(u2__abc_52155_new_n12410_), .B(u2__abc_52155_new_n12412_), .Y(u2__abc_52155_new_n12413_));
OR2X2 OR2X2_2395 ( .A(u2__abc_52155_new_n12417_), .B(u2__abc_52155_new_n12403_), .Y(u2__abc_52155_new_n12418_));
OR2X2 OR2X2_2396 ( .A(u2__abc_52155_new_n12422_), .B(u2__abc_52155_new_n4375_), .Y(u2__abc_52155_new_n12423_));
OR2X2 OR2X2_2397 ( .A(u2__abc_52155_new_n12421_), .B(u2__abc_52155_new_n12423_), .Y(u2__abc_52155_new_n12424_));
OR2X2 OR2X2_2398 ( .A(u2__abc_52155_new_n12425_), .B(u2__abc_52155_new_n12424_), .Y(u2__abc_52155_new_n12426_));
OR2X2 OR2X2_2399 ( .A(u2__abc_52155_new_n12426_), .B(u2__abc_52155_new_n4411_), .Y(u2__abc_52155_new_n12429_));
OR2X2 OR2X2_24 ( .A(_abc_73687_new_n753_), .B(\a[11] ), .Y(_abc_73687_new_n864_));
OR2X2 OR2X2_240 ( .A(\a[112] ), .B(\a[7] ), .Y(_abc_73687_new_n1191_));
OR2X2 OR2X2_2400 ( .A(u2__abc_52155_new_n12432_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12433_));
OR2X2 OR2X2_2401 ( .A(u2__abc_52155_new_n12431_), .B(u2__abc_52155_new_n12433_), .Y(u2__abc_52155_new_n12434_));
OR2X2 OR2X2_2402 ( .A(u2__abc_52155_new_n12438_), .B(u2__abc_52155_new_n12420_), .Y(u2__abc_52155_new_n12439_));
OR2X2 OR2X2_2403 ( .A(u2__abc_52155_new_n12443_), .B(u2__abc_52155_new_n4404_), .Y(u2__abc_52155_new_n12446_));
OR2X2 OR2X2_2404 ( .A(u2__abc_52155_new_n12449_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12450_));
OR2X2 OR2X2_2405 ( .A(u2__abc_52155_new_n12448_), .B(u2__abc_52155_new_n12450_), .Y(u2__abc_52155_new_n12451_));
OR2X2 OR2X2_2406 ( .A(u2__abc_52155_new_n12455_), .B(u2__abc_52155_new_n12441_), .Y(u2__abc_52155_new_n12456_));
OR2X2 OR2X2_2407 ( .A(u2__abc_52155_new_n12460_), .B(u2__abc_52155_new_n4389_), .Y(u2__abc_52155_new_n12463_));
OR2X2 OR2X2_2408 ( .A(u2__abc_52155_new_n12466_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12467_));
OR2X2 OR2X2_2409 ( .A(u2__abc_52155_new_n12465_), .B(u2__abc_52155_new_n12467_), .Y(u2__abc_52155_new_n12468_));
OR2X2 OR2X2_241 ( .A(_abc_73687_new_n1170_), .B(\a[8] ), .Y(_abc_73687_new_n1192_));
OR2X2 OR2X2_2410 ( .A(u2__abc_52155_new_n12472_), .B(u2__abc_52155_new_n12458_), .Y(u2__abc_52155_new_n12473_));
OR2X2 OR2X2_2411 ( .A(u2__abc_52155_new_n12480_), .B(u2__abc_52155_new_n12477_), .Y(u2__abc_52155_new_n12481_));
OR2X2 OR2X2_2412 ( .A(u2__abc_52155_new_n12483_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12484_));
OR2X2 OR2X2_2413 ( .A(u2__abc_52155_new_n12482_), .B(u2__abc_52155_new_n12484_), .Y(u2__abc_52155_new_n12485_));
OR2X2 OR2X2_2414 ( .A(u2__abc_52155_new_n12489_), .B(u2__abc_52155_new_n12475_), .Y(u2__abc_52155_new_n12490_));
OR2X2 OR2X2_2415 ( .A(u2__abc_52155_new_n4399_), .B(u2__abc_52155_new_n4406_), .Y(u2__abc_52155_new_n12494_));
OR2X2 OR2X2_2416 ( .A(u2__abc_52155_new_n12497_), .B(u2__abc_52155_new_n4391_), .Y(u2__abc_52155_new_n12498_));
OR2X2 OR2X2_2417 ( .A(u2__abc_52155_new_n12496_), .B(u2__abc_52155_new_n12498_), .Y(u2__abc_52155_new_n12499_));
OR2X2 OR2X2_2418 ( .A(u2__abc_52155_new_n12493_), .B(u2__abc_52155_new_n12499_), .Y(u2__abc_52155_new_n12500_));
OR2X2 OR2X2_2419 ( .A(u2__abc_52155_new_n12501_), .B(u2__abc_52155_new_n12500_), .Y(u2__abc_52155_new_n12502_));
OR2X2 OR2X2_242 ( .A(\a[112] ), .B(\a[8] ), .Y(_abc_73687_new_n1194_));
OR2X2 OR2X2_2420 ( .A(u2__abc_52155_new_n12502_), .B(u2__abc_52155_new_n4295_), .Y(u2__abc_52155_new_n12505_));
OR2X2 OR2X2_2421 ( .A(u2__abc_52155_new_n12508_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12509_));
OR2X2 OR2X2_2422 ( .A(u2__abc_52155_new_n12507_), .B(u2__abc_52155_new_n12509_), .Y(u2__abc_52155_new_n12510_));
OR2X2 OR2X2_2423 ( .A(u2__abc_52155_new_n12514_), .B(u2__abc_52155_new_n12492_), .Y(u2__abc_52155_new_n12515_));
OR2X2 OR2X2_2424 ( .A(u2__abc_52155_new_n12522_), .B(u2__abc_52155_new_n12519_), .Y(u2__abc_52155_new_n12523_));
OR2X2 OR2X2_2425 ( .A(u2__abc_52155_new_n12525_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12526_));
OR2X2 OR2X2_2426 ( .A(u2__abc_52155_new_n12524_), .B(u2__abc_52155_new_n12526_), .Y(u2__abc_52155_new_n12527_));
OR2X2 OR2X2_2427 ( .A(u2__abc_52155_new_n12531_), .B(u2__abc_52155_new_n12517_), .Y(u2__abc_52155_new_n12532_));
OR2X2 OR2X2_2428 ( .A(u2__abc_52155_new_n4291_), .B(u2__abc_52155_new_n4300_), .Y(u2__abc_52155_new_n12535_));
OR2X2 OR2X2_2429 ( .A(u2__abc_52155_new_n12538_), .B(u2__abc_52155_new_n12537_), .Y(u2__abc_52155_new_n12539_));
OR2X2 OR2X2_243 ( .A(_abc_73687_new_n1170_), .B(\a[9] ), .Y(_abc_73687_new_n1195_));
OR2X2 OR2X2_2430 ( .A(u2__abc_52155_new_n12539_), .B(u2__abc_52155_new_n4310_), .Y(u2__abc_52155_new_n12542_));
OR2X2 OR2X2_2431 ( .A(u2__abc_52155_new_n12545_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12546_));
OR2X2 OR2X2_2432 ( .A(u2__abc_52155_new_n12544_), .B(u2__abc_52155_new_n12546_), .Y(u2__abc_52155_new_n12547_));
OR2X2 OR2X2_2433 ( .A(u2__abc_52155_new_n12551_), .B(u2__abc_52155_new_n12534_), .Y(u2__abc_52155_new_n12552_));
OR2X2 OR2X2_2434 ( .A(u2__abc_52155_new_n12559_), .B(u2__abc_52155_new_n12556_), .Y(u2__abc_52155_new_n12560_));
OR2X2 OR2X2_2435 ( .A(u2__abc_52155_new_n12562_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12563_));
OR2X2 OR2X2_2436 ( .A(u2__abc_52155_new_n12561_), .B(u2__abc_52155_new_n12563_), .Y(u2__abc_52155_new_n12564_));
OR2X2 OR2X2_2437 ( .A(u2__abc_52155_new_n12568_), .B(u2__abc_52155_new_n12554_), .Y(u2__abc_52155_new_n12569_));
OR2X2 OR2X2_2438 ( .A(u2__abc_52155_new_n12573_), .B(u2__abc_52155_new_n4312_), .Y(u2__abc_52155_new_n12574_));
OR2X2 OR2X2_2439 ( .A(u2__abc_52155_new_n12572_), .B(u2__abc_52155_new_n12574_), .Y(u2__abc_52155_new_n12575_));
OR2X2 OR2X2_244 ( .A(\a[112] ), .B(\a[9] ), .Y(_abc_73687_new_n1197_));
OR2X2 OR2X2_2440 ( .A(u2__abc_52155_new_n12576_), .B(u2__abc_52155_new_n12575_), .Y(u2__abc_52155_new_n12577_));
OR2X2 OR2X2_2441 ( .A(u2__abc_52155_new_n12577_), .B(u2__abc_52155_new_n4348_), .Y(u2__abc_52155_new_n12580_));
OR2X2 OR2X2_2442 ( .A(u2__abc_52155_new_n12583_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12584_));
OR2X2 OR2X2_2443 ( .A(u2__abc_52155_new_n12582_), .B(u2__abc_52155_new_n12584_), .Y(u2__abc_52155_new_n12585_));
OR2X2 OR2X2_2444 ( .A(u2__abc_52155_new_n12589_), .B(u2__abc_52155_new_n12571_), .Y(u2__abc_52155_new_n12590_));
OR2X2 OR2X2_2445 ( .A(u2__abc_52155_new_n12597_), .B(u2__abc_52155_new_n12594_), .Y(u2__abc_52155_new_n12598_));
OR2X2 OR2X2_2446 ( .A(u2__abc_52155_new_n12600_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12601_));
OR2X2 OR2X2_2447 ( .A(u2__abc_52155_new_n12599_), .B(u2__abc_52155_new_n12601_), .Y(u2__abc_52155_new_n12602_));
OR2X2 OR2X2_2448 ( .A(u2__abc_52155_new_n12606_), .B(u2__abc_52155_new_n12592_), .Y(u2__abc_52155_new_n12607_));
OR2X2 OR2X2_2449 ( .A(u2__abc_52155_new_n12611_), .B(u2__abc_52155_new_n4339_), .Y(u2__abc_52155_new_n12612_));
OR2X2 OR2X2_245 ( .A(_abc_73687_new_n1170_), .B(\a[10] ), .Y(_abc_73687_new_n1198_));
OR2X2 OR2X2_2450 ( .A(u2__abc_52155_new_n12613_), .B(u2__abc_52155_new_n4326_), .Y(u2__abc_52155_new_n12616_));
OR2X2 OR2X2_2451 ( .A(u2__abc_52155_new_n12619_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12620_));
OR2X2 OR2X2_2452 ( .A(u2__abc_52155_new_n12618_), .B(u2__abc_52155_new_n12620_), .Y(u2__abc_52155_new_n12621_));
OR2X2 OR2X2_2453 ( .A(u2__abc_52155_new_n12625_), .B(u2__abc_52155_new_n12609_), .Y(u2__abc_52155_new_n12626_));
OR2X2 OR2X2_2454 ( .A(u2__abc_52155_new_n12633_), .B(u2__abc_52155_new_n12630_), .Y(u2__abc_52155_new_n12634_));
OR2X2 OR2X2_2455 ( .A(u2__abc_52155_new_n12636_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12637_));
OR2X2 OR2X2_2456 ( .A(u2__abc_52155_new_n12635_), .B(u2__abc_52155_new_n12637_), .Y(u2__abc_52155_new_n12638_));
OR2X2 OR2X2_2457 ( .A(u2__abc_52155_new_n12642_), .B(u2__abc_52155_new_n12628_), .Y(u2__abc_52155_new_n12643_));
OR2X2 OR2X2_2458 ( .A(u2__abc_52155_new_n12610_), .B(u2__abc_52155_new_n4339_), .Y(u2__abc_52155_new_n12652_));
OR2X2 OR2X2_2459 ( .A(u2__abc_52155_new_n12655_), .B(u2__abc_52155_new_n4331_), .Y(u2__abc_52155_new_n12656_));
OR2X2 OR2X2_246 ( .A(\a[112] ), .B(\a[10] ), .Y(_abc_73687_new_n1200_));
OR2X2 OR2X2_2460 ( .A(u2__abc_52155_new_n12654_), .B(u2__abc_52155_new_n12656_), .Y(u2__abc_52155_new_n12657_));
OR2X2 OR2X2_2461 ( .A(u2__abc_52155_new_n12651_), .B(u2__abc_52155_new_n12657_), .Y(u2__abc_52155_new_n12658_));
OR2X2 OR2X2_2462 ( .A(u2__abc_52155_new_n12650_), .B(u2__abc_52155_new_n12658_), .Y(u2__abc_52155_new_n12659_));
OR2X2 OR2X2_2463 ( .A(u2__abc_52155_new_n12649_), .B(u2__abc_52155_new_n12659_), .Y(u2__abc_52155_new_n12660_));
OR2X2 OR2X2_2464 ( .A(u2__abc_52155_new_n12660_), .B(u2__abc_52155_new_n12648_), .Y(u2__abc_52155_new_n12661_));
OR2X2 OR2X2_2465 ( .A(u2__abc_52155_new_n12647_), .B(u2__abc_52155_new_n12661_), .Y(u2__abc_52155_new_n12662_));
OR2X2 OR2X2_2466 ( .A(u2__abc_52155_new_n12646_), .B(u2__abc_52155_new_n12662_), .Y(u2__abc_52155_new_n12663_));
OR2X2 OR2X2_2467 ( .A(u2__abc_52155_new_n12663_), .B(u2__abc_52155_new_n6545_), .Y(u2__abc_52155_new_n12666_));
OR2X2 OR2X2_2468 ( .A(u2__abc_52155_new_n12669_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12670_));
OR2X2 OR2X2_2469 ( .A(u2__abc_52155_new_n12668_), .B(u2__abc_52155_new_n12670_), .Y(u2__abc_52155_new_n12671_));
OR2X2 OR2X2_247 ( .A(_abc_73687_new_n1170_), .B(\a[11] ), .Y(_abc_73687_new_n1201_));
OR2X2 OR2X2_2470 ( .A(u2__abc_52155_new_n12675_), .B(u2__abc_52155_new_n12645_), .Y(u2__abc_52155_new_n12676_));
OR2X2 OR2X2_2471 ( .A(u2__abc_52155_new_n12680_), .B(u2__abc_52155_new_n12679_), .Y(u2__abc_52155_new_n12681_));
OR2X2 OR2X2_2472 ( .A(u2__abc_52155_new_n12682_), .B(u2__abc_52155_new_n6552_), .Y(u2__abc_52155_new_n12683_));
OR2X2 OR2X2_2473 ( .A(u2__abc_52155_new_n12686_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12687_));
OR2X2 OR2X2_2474 ( .A(u2__abc_52155_new_n12685_), .B(u2__abc_52155_new_n12687_), .Y(u2__abc_52155_new_n12688_));
OR2X2 OR2X2_2475 ( .A(u2__abc_52155_new_n12692_), .B(u2__abc_52155_new_n12678_), .Y(u2__abc_52155_new_n12693_));
OR2X2 OR2X2_2476 ( .A(u2__abc_52155_new_n12696_), .B(u2__abc_52155_new_n6547_), .Y(u2__abc_52155_new_n12697_));
OR2X2 OR2X2_2477 ( .A(u2__abc_52155_new_n12699_), .B(u2__abc_52155_new_n12698_), .Y(u2__abc_52155_new_n12700_));
OR2X2 OR2X2_2478 ( .A(u2__abc_52155_new_n12700_), .B(u2__abc_52155_new_n6560_), .Y(u2__abc_52155_new_n12703_));
OR2X2 OR2X2_2479 ( .A(u2__abc_52155_new_n12706_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12707_));
OR2X2 OR2X2_248 ( .A(\a[112] ), .B(\a[11] ), .Y(_abc_73687_new_n1203_));
OR2X2 OR2X2_2480 ( .A(u2__abc_52155_new_n12705_), .B(u2__abc_52155_new_n12707_), .Y(u2__abc_52155_new_n12708_));
OR2X2 OR2X2_2481 ( .A(u2__abc_52155_new_n12712_), .B(u2__abc_52155_new_n12695_), .Y(u2__abc_52155_new_n12713_));
OR2X2 OR2X2_2482 ( .A(u2__abc_52155_new_n12717_), .B(u2__abc_52155_new_n12716_), .Y(u2__abc_52155_new_n12718_));
OR2X2 OR2X2_2483 ( .A(u2__abc_52155_new_n12719_), .B(u2__abc_52155_new_n6567_), .Y(u2__abc_52155_new_n12720_));
OR2X2 OR2X2_2484 ( .A(u2__abc_52155_new_n12723_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12724_));
OR2X2 OR2X2_2485 ( .A(u2__abc_52155_new_n12722_), .B(u2__abc_52155_new_n12724_), .Y(u2__abc_52155_new_n12725_));
OR2X2 OR2X2_2486 ( .A(u2__abc_52155_new_n12729_), .B(u2__abc_52155_new_n12715_), .Y(u2__abc_52155_new_n12730_));
OR2X2 OR2X2_2487 ( .A(u2__abc_52155_new_n12734_), .B(u2__abc_52155_new_n6562_), .Y(u2__abc_52155_new_n12735_));
OR2X2 OR2X2_2488 ( .A(u2__abc_52155_new_n12733_), .B(u2__abc_52155_new_n12735_), .Y(u2__abc_52155_new_n12736_));
OR2X2 OR2X2_2489 ( .A(u2__abc_52155_new_n12737_), .B(u2__abc_52155_new_n12736_), .Y(u2__abc_52155_new_n12738_));
OR2X2 OR2X2_249 ( .A(_abc_73687_new_n1170_), .B(\a[12] ), .Y(_abc_73687_new_n1204_));
OR2X2 OR2X2_2490 ( .A(u2__abc_52155_new_n12738_), .B(u2__abc_52155_new_n6591_), .Y(u2__abc_52155_new_n12741_));
OR2X2 OR2X2_2491 ( .A(u2__abc_52155_new_n12744_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12745_));
OR2X2 OR2X2_2492 ( .A(u2__abc_52155_new_n12743_), .B(u2__abc_52155_new_n12745_), .Y(u2__abc_52155_new_n12746_));
OR2X2 OR2X2_2493 ( .A(u2__abc_52155_new_n12750_), .B(u2__abc_52155_new_n12732_), .Y(u2__abc_52155_new_n12751_));
OR2X2 OR2X2_2494 ( .A(u2__abc_52155_new_n12758_), .B(u2__abc_52155_new_n12755_), .Y(u2__abc_52155_new_n12759_));
OR2X2 OR2X2_2495 ( .A(u2__abc_52155_new_n12761_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12762_));
OR2X2 OR2X2_2496 ( .A(u2__abc_52155_new_n12760_), .B(u2__abc_52155_new_n12762_), .Y(u2__abc_52155_new_n12763_));
OR2X2 OR2X2_2497 ( .A(u2__abc_52155_new_n12767_), .B(u2__abc_52155_new_n12753_), .Y(u2__abc_52155_new_n12768_));
OR2X2 OR2X2_2498 ( .A(u2__abc_52155_new_n12772_), .B(u2__abc_52155_new_n6596_), .Y(u2__abc_52155_new_n12773_));
OR2X2 OR2X2_2499 ( .A(u2__abc_52155_new_n12774_), .B(u2__abc_52155_new_n6576_), .Y(u2__abc_52155_new_n12777_));
OR2X2 OR2X2_25 ( .A(aNan), .B(sqrto_88_), .Y(_abc_73687_new_n866_));
OR2X2 OR2X2_250 ( .A(\a[112] ), .B(\a[12] ), .Y(_abc_73687_new_n1206_));
OR2X2 OR2X2_2500 ( .A(u2__abc_52155_new_n12780_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12781_));
OR2X2 OR2X2_2501 ( .A(u2__abc_52155_new_n12779_), .B(u2__abc_52155_new_n12781_), .Y(u2__abc_52155_new_n12782_));
OR2X2 OR2X2_2502 ( .A(u2__abc_52155_new_n12786_), .B(u2__abc_52155_new_n12770_), .Y(u2__abc_52155_new_n12787_));
OR2X2 OR2X2_2503 ( .A(u2__abc_52155_new_n12791_), .B(u2__abc_52155_new_n12790_), .Y(u2__abc_52155_new_n12792_));
OR2X2 OR2X2_2504 ( .A(u2__abc_52155_new_n12793_), .B(u2__abc_52155_new_n6583_), .Y(u2__abc_52155_new_n12794_));
OR2X2 OR2X2_2505 ( .A(u2__abc_52155_new_n12797_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12798_));
OR2X2 OR2X2_2506 ( .A(u2__abc_52155_new_n12796_), .B(u2__abc_52155_new_n12798_), .Y(u2__abc_52155_new_n12799_));
OR2X2 OR2X2_2507 ( .A(u2__abc_52155_new_n12803_), .B(u2__abc_52155_new_n12789_), .Y(u2__abc_52155_new_n12804_));
OR2X2 OR2X2_2508 ( .A(u2__abc_52155_new_n12771_), .B(u2__abc_52155_new_n6596_), .Y(u2__abc_52155_new_n12809_));
OR2X2 OR2X2_2509 ( .A(u2__abc_52155_new_n6641_), .B(u2__abc_52155_new_n12809_), .Y(u2__abc_52155_new_n12810_));
OR2X2 OR2X2_251 ( .A(_abc_73687_new_n1170_), .B(\a[13] ), .Y(_abc_73687_new_n1207_));
OR2X2 OR2X2_2510 ( .A(u2__abc_52155_new_n6571_), .B(u2__abc_52155_new_n6578_), .Y(u2__abc_52155_new_n12811_));
OR2X2 OR2X2_2511 ( .A(u2__abc_52155_new_n12817_), .B(u2__abc_52155_new_n12816_), .Y(u2__abc_52155_new_n12818_));
OR2X2 OR2X2_2512 ( .A(u2__abc_52155_new_n12818_), .B(u2__abc_52155_new_n6528_), .Y(u2__abc_52155_new_n12821_));
OR2X2 OR2X2_2513 ( .A(u2__abc_52155_new_n12824_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12825_));
OR2X2 OR2X2_2514 ( .A(u2__abc_52155_new_n12823_), .B(u2__abc_52155_new_n12825_), .Y(u2__abc_52155_new_n12826_));
OR2X2 OR2X2_2515 ( .A(u2__abc_52155_new_n12830_), .B(u2__abc_52155_new_n12806_), .Y(u2__abc_52155_new_n12831_));
OR2X2 OR2X2_2516 ( .A(u2__abc_52155_new_n12835_), .B(u2__abc_52155_new_n12834_), .Y(u2__abc_52155_new_n12836_));
OR2X2 OR2X2_2517 ( .A(u2__abc_52155_new_n12837_), .B(u2__abc_52155_new_n6535_), .Y(u2__abc_52155_new_n12838_));
OR2X2 OR2X2_2518 ( .A(u2__abc_52155_new_n12841_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12842_));
OR2X2 OR2X2_2519 ( .A(u2__abc_52155_new_n12840_), .B(u2__abc_52155_new_n12842_), .Y(u2__abc_52155_new_n12843_));
OR2X2 OR2X2_252 ( .A(\a[112] ), .B(\a[13] ), .Y(_abc_73687_new_n1209_));
OR2X2 OR2X2_2520 ( .A(u2__abc_52155_new_n12847_), .B(u2__abc_52155_new_n12833_), .Y(u2__abc_52155_new_n12848_));
OR2X2 OR2X2_2521 ( .A(u2__abc_52155_new_n12851_), .B(u2__abc_52155_new_n6530_), .Y(u2__abc_52155_new_n12852_));
OR2X2 OR2X2_2522 ( .A(u2__abc_52155_new_n12854_), .B(u2__abc_52155_new_n12853_), .Y(u2__abc_52155_new_n12855_));
OR2X2 OR2X2_2523 ( .A(u2__abc_52155_new_n12855_), .B(u2__abc_52155_new_n6513_), .Y(u2__abc_52155_new_n12858_));
OR2X2 OR2X2_2524 ( .A(u2__abc_52155_new_n12861_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12862_));
OR2X2 OR2X2_2525 ( .A(u2__abc_52155_new_n12860_), .B(u2__abc_52155_new_n12862_), .Y(u2__abc_52155_new_n12863_));
OR2X2 OR2X2_2526 ( .A(u2__abc_52155_new_n12867_), .B(u2__abc_52155_new_n12850_), .Y(u2__abc_52155_new_n12868_));
OR2X2 OR2X2_2527 ( .A(u2__abc_52155_new_n12872_), .B(u2__abc_52155_new_n12871_), .Y(u2__abc_52155_new_n12873_));
OR2X2 OR2X2_2528 ( .A(u2__abc_52155_new_n12874_), .B(u2__abc_52155_new_n6520_), .Y(u2__abc_52155_new_n12875_));
OR2X2 OR2X2_2529 ( .A(u2__abc_52155_new_n12878_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12879_));
OR2X2 OR2X2_253 ( .A(_abc_73687_new_n1170_), .B(\a[14] ), .Y(_abc_73687_new_n1210_));
OR2X2 OR2X2_2530 ( .A(u2__abc_52155_new_n12877_), .B(u2__abc_52155_new_n12879_), .Y(u2__abc_52155_new_n12880_));
OR2X2 OR2X2_2531 ( .A(u2__abc_52155_new_n12884_), .B(u2__abc_52155_new_n12870_), .Y(u2__abc_52155_new_n12885_));
OR2X2 OR2X2_2532 ( .A(u2__abc_52155_new_n12889_), .B(u2__abc_52155_new_n6518_), .Y(u2__abc_52155_new_n12890_));
OR2X2 OR2X2_2533 ( .A(u2__abc_52155_new_n12891_), .B(u2__abc_52155_new_n6497_), .Y(u2__abc_52155_new_n12894_));
OR2X2 OR2X2_2534 ( .A(u2__abc_52155_new_n12897_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12898_));
OR2X2 OR2X2_2535 ( .A(u2__abc_52155_new_n12896_), .B(u2__abc_52155_new_n12898_), .Y(u2__abc_52155_new_n12899_));
OR2X2 OR2X2_2536 ( .A(u2__abc_52155_new_n12903_), .B(u2__abc_52155_new_n12887_), .Y(u2__abc_52155_new_n12904_));
OR2X2 OR2X2_2537 ( .A(u2__abc_52155_new_n12911_), .B(u2__abc_52155_new_n12908_), .Y(u2__abc_52155_new_n12912_));
OR2X2 OR2X2_2538 ( .A(u2__abc_52155_new_n12914_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12915_));
OR2X2 OR2X2_2539 ( .A(u2__abc_52155_new_n12913_), .B(u2__abc_52155_new_n12915_), .Y(u2__abc_52155_new_n12916_));
OR2X2 OR2X2_254 ( .A(\a[112] ), .B(\a[14] ), .Y(_abc_73687_new_n1212_));
OR2X2 OR2X2_2540 ( .A(u2__abc_52155_new_n12920_), .B(u2__abc_52155_new_n12906_), .Y(u2__abc_52155_new_n12921_));
OR2X2 OR2X2_2541 ( .A(u2__abc_52155_new_n12925_), .B(u2__abc_52155_new_n6502_), .Y(u2__abc_52155_new_n12926_));
OR2X2 OR2X2_2542 ( .A(u2__abc_52155_new_n12927_), .B(u2__abc_52155_new_n6482_), .Y(u2__abc_52155_new_n12930_));
OR2X2 OR2X2_2543 ( .A(u2__abc_52155_new_n12933_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12934_));
OR2X2 OR2X2_2544 ( .A(u2__abc_52155_new_n12932_), .B(u2__abc_52155_new_n12934_), .Y(u2__abc_52155_new_n12935_));
OR2X2 OR2X2_2545 ( .A(u2__abc_52155_new_n12939_), .B(u2__abc_52155_new_n12923_), .Y(u2__abc_52155_new_n12940_));
OR2X2 OR2X2_2546 ( .A(u2__abc_52155_new_n12944_), .B(u2__abc_52155_new_n12943_), .Y(u2__abc_52155_new_n12945_));
OR2X2 OR2X2_2547 ( .A(u2__abc_52155_new_n12946_), .B(u2__abc_52155_new_n6489_), .Y(u2__abc_52155_new_n12947_));
OR2X2 OR2X2_2548 ( .A(u2__abc_52155_new_n12950_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12951_));
OR2X2 OR2X2_2549 ( .A(u2__abc_52155_new_n12949_), .B(u2__abc_52155_new_n12951_), .Y(u2__abc_52155_new_n12952_));
OR2X2 OR2X2_255 ( .A(_abc_73687_new_n1170_), .B(\a[15] ), .Y(_abc_73687_new_n1213_));
OR2X2 OR2X2_2550 ( .A(u2__abc_52155_new_n12956_), .B(u2__abc_52155_new_n12942_), .Y(u2__abc_52155_new_n12957_));
OR2X2 OR2X2_2551 ( .A(u2__abc_52155_new_n12888_), .B(u2__abc_52155_new_n6518_), .Y(u2__abc_52155_new_n12962_));
OR2X2 OR2X2_2552 ( .A(u2__abc_52155_new_n12965_), .B(u2__abc_52155_new_n6651_), .Y(u2__abc_52155_new_n12966_));
OR2X2 OR2X2_2553 ( .A(u2__abc_52155_new_n12967_), .B(u2__abc_52155_new_n6484_), .Y(u2__abc_52155_new_n12968_));
OR2X2 OR2X2_2554 ( .A(u2__abc_52155_new_n12924_), .B(u2__abc_52155_new_n6502_), .Y(u2__abc_52155_new_n12969_));
OR2X2 OR2X2_2555 ( .A(u2__abc_52155_new_n6663_), .B(u2__abc_52155_new_n12969_), .Y(u2__abc_52155_new_n12970_));
OR2X2 OR2X2_2556 ( .A(u2__abc_52155_new_n12975_), .B(u2__abc_52155_new_n12974_), .Y(u2__abc_52155_new_n12976_));
OR2X2 OR2X2_2557 ( .A(u2__abc_52155_new_n12976_), .B(u2__abc_52155_new_n6433_), .Y(u2__abc_52155_new_n12979_));
OR2X2 OR2X2_2558 ( .A(u2__abc_52155_new_n12982_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n12983_));
OR2X2 OR2X2_2559 ( .A(u2__abc_52155_new_n12981_), .B(u2__abc_52155_new_n12983_), .Y(u2__abc_52155_new_n12984_));
OR2X2 OR2X2_256 ( .A(\a[112] ), .B(\a[15] ), .Y(_abc_73687_new_n1215_));
OR2X2 OR2X2_2560 ( .A(u2__abc_52155_new_n12988_), .B(u2__abc_52155_new_n12959_), .Y(u2__abc_52155_new_n12989_));
OR2X2 OR2X2_2561 ( .A(u2__abc_52155_new_n12996_), .B(u2__abc_52155_new_n12993_), .Y(u2__abc_52155_new_n12997_));
OR2X2 OR2X2_2562 ( .A(u2__abc_52155_new_n12999_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13000_));
OR2X2 OR2X2_2563 ( .A(u2__abc_52155_new_n12998_), .B(u2__abc_52155_new_n13000_), .Y(u2__abc_52155_new_n13001_));
OR2X2 OR2X2_2564 ( .A(u2__abc_52155_new_n13005_), .B(u2__abc_52155_new_n12991_), .Y(u2__abc_52155_new_n13006_));
OR2X2 OR2X2_2565 ( .A(u2__abc_52155_new_n13010_), .B(u2__abc_52155_new_n6438_), .Y(u2__abc_52155_new_n13011_));
OR2X2 OR2X2_2566 ( .A(u2__abc_52155_new_n13012_), .B(u2__abc_52155_new_n6418_), .Y(u2__abc_52155_new_n13015_));
OR2X2 OR2X2_2567 ( .A(u2__abc_52155_new_n13018_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13019_));
OR2X2 OR2X2_2568 ( .A(u2__abc_52155_new_n13017_), .B(u2__abc_52155_new_n13019_), .Y(u2__abc_52155_new_n13020_));
OR2X2 OR2X2_2569 ( .A(u2__abc_52155_new_n13024_), .B(u2__abc_52155_new_n13008_), .Y(u2__abc_52155_new_n13025_));
OR2X2 OR2X2_257 ( .A(_abc_73687_new_n1170_), .B(\a[16] ), .Y(_abc_73687_new_n1216_));
OR2X2 OR2X2_2570 ( .A(u2__abc_52155_new_n13029_), .B(u2__abc_52155_new_n13028_), .Y(u2__abc_52155_new_n13030_));
OR2X2 OR2X2_2571 ( .A(u2__abc_52155_new_n13031_), .B(u2__abc_52155_new_n6425_), .Y(u2__abc_52155_new_n13032_));
OR2X2 OR2X2_2572 ( .A(u2__abc_52155_new_n13035_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13036_));
OR2X2 OR2X2_2573 ( .A(u2__abc_52155_new_n13034_), .B(u2__abc_52155_new_n13036_), .Y(u2__abc_52155_new_n13037_));
OR2X2 OR2X2_2574 ( .A(u2__abc_52155_new_n13041_), .B(u2__abc_52155_new_n13027_), .Y(u2__abc_52155_new_n13042_));
OR2X2 OR2X2_2575 ( .A(u2__abc_52155_new_n6413_), .B(u2__abc_52155_new_n6420_), .Y(u2__abc_52155_new_n13045_));
OR2X2 OR2X2_2576 ( .A(u2__abc_52155_new_n13009_), .B(u2__abc_52155_new_n6438_), .Y(u2__abc_52155_new_n13048_));
OR2X2 OR2X2_2577 ( .A(u2__abc_52155_new_n6614_), .B(u2__abc_52155_new_n13048_), .Y(u2__abc_52155_new_n13049_));
OR2X2 OR2X2_2578 ( .A(u2__abc_52155_new_n13052_), .B(u2__abc_52155_new_n13051_), .Y(u2__abc_52155_new_n13053_));
OR2X2 OR2X2_2579 ( .A(u2__abc_52155_new_n13053_), .B(u2__abc_52155_new_n6464_), .Y(u2__abc_52155_new_n13056_));
OR2X2 OR2X2_258 ( .A(\a[112] ), .B(\a[16] ), .Y(_abc_73687_new_n1218_));
OR2X2 OR2X2_2580 ( .A(u2__abc_52155_new_n13059_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13060_));
OR2X2 OR2X2_2581 ( .A(u2__abc_52155_new_n13058_), .B(u2__abc_52155_new_n13060_), .Y(u2__abc_52155_new_n13061_));
OR2X2 OR2X2_2582 ( .A(u2__abc_52155_new_n13065_), .B(u2__abc_52155_new_n13044_), .Y(u2__abc_52155_new_n13066_));
OR2X2 OR2X2_2583 ( .A(u2__abc_52155_new_n13073_), .B(u2__abc_52155_new_n13070_), .Y(u2__abc_52155_new_n13074_));
OR2X2 OR2X2_2584 ( .A(u2__abc_52155_new_n13076_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13077_));
OR2X2 OR2X2_2585 ( .A(u2__abc_52155_new_n13075_), .B(u2__abc_52155_new_n13077_), .Y(u2__abc_52155_new_n13078_));
OR2X2 OR2X2_2586 ( .A(u2__abc_52155_new_n13082_), .B(u2__abc_52155_new_n13068_), .Y(u2__abc_52155_new_n13083_));
OR2X2 OR2X2_2587 ( .A(u2__abc_52155_new_n13087_), .B(u2__abc_52155_new_n6469_), .Y(u2__abc_52155_new_n13088_));
OR2X2 OR2X2_2588 ( .A(u2__abc_52155_new_n13089_), .B(u2__abc_52155_new_n6449_), .Y(u2__abc_52155_new_n13092_));
OR2X2 OR2X2_2589 ( .A(u2__abc_52155_new_n13095_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13096_));
OR2X2 OR2X2_259 ( .A(_abc_73687_new_n1170_), .B(\a[17] ), .Y(_abc_73687_new_n1219_));
OR2X2 OR2X2_2590 ( .A(u2__abc_52155_new_n13094_), .B(u2__abc_52155_new_n13096_), .Y(u2__abc_52155_new_n13097_));
OR2X2 OR2X2_2591 ( .A(u2__abc_52155_new_n13101_), .B(u2__abc_52155_new_n13085_), .Y(u2__abc_52155_new_n13102_));
OR2X2 OR2X2_2592 ( .A(u2__abc_52155_new_n13106_), .B(u2__abc_52155_new_n13105_), .Y(u2__abc_52155_new_n13107_));
OR2X2 OR2X2_2593 ( .A(u2__abc_52155_new_n13108_), .B(u2__abc_52155_new_n6456_), .Y(u2__abc_52155_new_n13109_));
OR2X2 OR2X2_2594 ( .A(u2__abc_52155_new_n13112_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13113_));
OR2X2 OR2X2_2595 ( .A(u2__abc_52155_new_n13111_), .B(u2__abc_52155_new_n13113_), .Y(u2__abc_52155_new_n13114_));
OR2X2 OR2X2_2596 ( .A(u2__abc_52155_new_n13118_), .B(u2__abc_52155_new_n13104_), .Y(u2__abc_52155_new_n13119_));
OR2X2 OR2X2_2597 ( .A(u2__abc_52155_new_n13086_), .B(u2__abc_52155_new_n6469_), .Y(u2__abc_52155_new_n13124_));
OR2X2 OR2X2_2598 ( .A(u2__abc_52155_new_n6624_), .B(u2__abc_52155_new_n13124_), .Y(u2__abc_52155_new_n13125_));
OR2X2 OR2X2_2599 ( .A(u2__abc_52155_new_n13126_), .B(u2__abc_52155_new_n6454_), .Y(u2__abc_52155_new_n13127_));
OR2X2 OR2X2_26 ( .A(_abc_73687_new_n753_), .B(\a[12] ), .Y(_abc_73687_new_n867_));
OR2X2 OR2X2_260 ( .A(\a[112] ), .B(\a[17] ), .Y(_abc_73687_new_n1221_));
OR2X2 OR2X2_2600 ( .A(u2__abc_52155_new_n13131_), .B(u2__abc_52155_new_n13130_), .Y(u2__abc_52155_new_n13132_));
OR2X2 OR2X2_2601 ( .A(u2__abc_52155_new_n13132_), .B(u2__abc_52155_new_n6370_), .Y(u2__abc_52155_new_n13135_));
OR2X2 OR2X2_2602 ( .A(u2__abc_52155_new_n13138_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13139_));
OR2X2 OR2X2_2603 ( .A(u2__abc_52155_new_n13137_), .B(u2__abc_52155_new_n13139_), .Y(u2__abc_52155_new_n13140_));
OR2X2 OR2X2_2604 ( .A(u2__abc_52155_new_n13144_), .B(u2__abc_52155_new_n13121_), .Y(u2__abc_52155_new_n13145_));
OR2X2 OR2X2_2605 ( .A(u2__abc_52155_new_n13152_), .B(u2__abc_52155_new_n13149_), .Y(u2__abc_52155_new_n13153_));
OR2X2 OR2X2_2606 ( .A(u2__abc_52155_new_n13155_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13156_));
OR2X2 OR2X2_2607 ( .A(u2__abc_52155_new_n13154_), .B(u2__abc_52155_new_n13156_), .Y(u2__abc_52155_new_n13157_));
OR2X2 OR2X2_2608 ( .A(u2__abc_52155_new_n13161_), .B(u2__abc_52155_new_n13147_), .Y(u2__abc_52155_new_n13162_));
OR2X2 OR2X2_2609 ( .A(u2__abc_52155_new_n13166_), .B(u2__abc_52155_new_n6375_), .Y(u2__abc_52155_new_n13167_));
OR2X2 OR2X2_261 ( .A(_abc_73687_new_n1170_), .B(\a[18] ), .Y(_abc_73687_new_n1222_));
OR2X2 OR2X2_2610 ( .A(u2__abc_52155_new_n13168_), .B(u2__abc_52155_new_n6355_), .Y(u2__abc_52155_new_n13171_));
OR2X2 OR2X2_2611 ( .A(u2__abc_52155_new_n13174_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13175_));
OR2X2 OR2X2_2612 ( .A(u2__abc_52155_new_n13173_), .B(u2__abc_52155_new_n13175_), .Y(u2__abc_52155_new_n13176_));
OR2X2 OR2X2_2613 ( .A(u2__abc_52155_new_n13180_), .B(u2__abc_52155_new_n13164_), .Y(u2__abc_52155_new_n13181_));
OR2X2 OR2X2_2614 ( .A(u2__abc_52155_new_n13185_), .B(u2__abc_52155_new_n13184_), .Y(u2__abc_52155_new_n13186_));
OR2X2 OR2X2_2615 ( .A(u2__abc_52155_new_n13187_), .B(u2__abc_52155_new_n6362_), .Y(u2__abc_52155_new_n13188_));
OR2X2 OR2X2_2616 ( .A(u2__abc_52155_new_n13191_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13192_));
OR2X2 OR2X2_2617 ( .A(u2__abc_52155_new_n13190_), .B(u2__abc_52155_new_n13192_), .Y(u2__abc_52155_new_n13193_));
OR2X2 OR2X2_2618 ( .A(u2__abc_52155_new_n13197_), .B(u2__abc_52155_new_n13183_), .Y(u2__abc_52155_new_n13198_));
OR2X2 OR2X2_2619 ( .A(u2__abc_52155_new_n13165_), .B(u2__abc_52155_new_n6375_), .Y(u2__abc_52155_new_n13201_));
OR2X2 OR2X2_262 ( .A(\a[112] ), .B(\a[18] ), .Y(_abc_73687_new_n1224_));
OR2X2 OR2X2_2620 ( .A(u2__abc_52155_new_n6672_), .B(u2__abc_52155_new_n13201_), .Y(u2__abc_52155_new_n13202_));
OR2X2 OR2X2_2621 ( .A(u2__abc_52155_new_n13203_), .B(u2__abc_52155_new_n6357_), .Y(u2__abc_52155_new_n13204_));
OR2X2 OR2X2_2622 ( .A(u2__abc_52155_new_n13208_), .B(u2__abc_52155_new_n13207_), .Y(u2__abc_52155_new_n13209_));
OR2X2 OR2X2_2623 ( .A(u2__abc_52155_new_n13209_), .B(u2__abc_52155_new_n6401_), .Y(u2__abc_52155_new_n13212_));
OR2X2 OR2X2_2624 ( .A(u2__abc_52155_new_n13215_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13216_));
OR2X2 OR2X2_2625 ( .A(u2__abc_52155_new_n13214_), .B(u2__abc_52155_new_n13216_), .Y(u2__abc_52155_new_n13217_));
OR2X2 OR2X2_2626 ( .A(u2__abc_52155_new_n13221_), .B(u2__abc_52155_new_n13200_), .Y(u2__abc_52155_new_n13222_));
OR2X2 OR2X2_2627 ( .A(u2__abc_52155_new_n13229_), .B(u2__abc_52155_new_n13226_), .Y(u2__abc_52155_new_n13230_));
OR2X2 OR2X2_2628 ( .A(u2__abc_52155_new_n13232_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13233_));
OR2X2 OR2X2_2629 ( .A(u2__abc_52155_new_n13231_), .B(u2__abc_52155_new_n13233_), .Y(u2__abc_52155_new_n13234_));
OR2X2 OR2X2_263 ( .A(_abc_73687_new_n1170_), .B(\a[19] ), .Y(_abc_73687_new_n1225_));
OR2X2 OR2X2_2630 ( .A(u2__abc_52155_new_n13238_), .B(u2__abc_52155_new_n13224_), .Y(u2__abc_52155_new_n13239_));
OR2X2 OR2X2_2631 ( .A(u2__abc_52155_new_n13243_), .B(u2__abc_52155_new_n6406_), .Y(u2__abc_52155_new_n13244_));
OR2X2 OR2X2_2632 ( .A(u2__abc_52155_new_n13245_), .B(u2__abc_52155_new_n6386_), .Y(u2__abc_52155_new_n13248_));
OR2X2 OR2X2_2633 ( .A(u2__abc_52155_new_n13251_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13252_));
OR2X2 OR2X2_2634 ( .A(u2__abc_52155_new_n13250_), .B(u2__abc_52155_new_n13252_), .Y(u2__abc_52155_new_n13253_));
OR2X2 OR2X2_2635 ( .A(u2__abc_52155_new_n13257_), .B(u2__abc_52155_new_n13241_), .Y(u2__abc_52155_new_n13258_));
OR2X2 OR2X2_2636 ( .A(u2__abc_52155_new_n13262_), .B(u2__abc_52155_new_n13261_), .Y(u2__abc_52155_new_n13263_));
OR2X2 OR2X2_2637 ( .A(u2__abc_52155_new_n13264_), .B(u2__abc_52155_new_n6393_), .Y(u2__abc_52155_new_n13265_));
OR2X2 OR2X2_2638 ( .A(u2__abc_52155_new_n13268_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13269_));
OR2X2 OR2X2_2639 ( .A(u2__abc_52155_new_n13267_), .B(u2__abc_52155_new_n13269_), .Y(u2__abc_52155_new_n13270_));
OR2X2 OR2X2_264 ( .A(\a[112] ), .B(\a[19] ), .Y(_abc_73687_new_n1227_));
OR2X2 OR2X2_2640 ( .A(u2__abc_52155_new_n13274_), .B(u2__abc_52155_new_n13260_), .Y(u2__abc_52155_new_n13275_));
OR2X2 OR2X2_2641 ( .A(u2__abc_52155_new_n13242_), .B(u2__abc_52155_new_n6406_), .Y(u2__abc_52155_new_n13284_));
OR2X2 OR2X2_2642 ( .A(u2__abc_52155_new_n6681_), .B(u2__abc_52155_new_n13284_), .Y(u2__abc_52155_new_n13285_));
OR2X2 OR2X2_2643 ( .A(u2__abc_52155_new_n13286_), .B(u2__abc_52155_new_n6388_), .Y(u2__abc_52155_new_n13287_));
OR2X2 OR2X2_2644 ( .A(u2__abc_52155_new_n13294_), .B(u2__abc_52155_new_n13293_), .Y(u2__abc_52155_new_n13295_));
OR2X2 OR2X2_2645 ( .A(u2__abc_52155_new_n13295_), .B(u2__abc_52155_new_n6305_), .Y(u2__abc_52155_new_n13298_));
OR2X2 OR2X2_2646 ( .A(u2__abc_52155_new_n13301_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13302_));
OR2X2 OR2X2_2647 ( .A(u2__abc_52155_new_n13300_), .B(u2__abc_52155_new_n13302_), .Y(u2__abc_52155_new_n13303_));
OR2X2 OR2X2_2648 ( .A(u2__abc_52155_new_n13307_), .B(u2__abc_52155_new_n13277_), .Y(u2__abc_52155_new_n13308_));
OR2X2 OR2X2_2649 ( .A(u2__abc_52155_new_n13315_), .B(u2__abc_52155_new_n13312_), .Y(u2__abc_52155_new_n13316_));
OR2X2 OR2X2_265 ( .A(_abc_73687_new_n1170_), .B(\a[20] ), .Y(_abc_73687_new_n1228_));
OR2X2 OR2X2_2650 ( .A(u2__abc_52155_new_n13318_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13319_));
OR2X2 OR2X2_2651 ( .A(u2__abc_52155_new_n13317_), .B(u2__abc_52155_new_n13319_), .Y(u2__abc_52155_new_n13320_));
OR2X2 OR2X2_2652 ( .A(u2__abc_52155_new_n13324_), .B(u2__abc_52155_new_n13310_), .Y(u2__abc_52155_new_n13325_));
OR2X2 OR2X2_2653 ( .A(u2__abc_52155_new_n13329_), .B(u2__abc_52155_new_n6310_), .Y(u2__abc_52155_new_n13330_));
OR2X2 OR2X2_2654 ( .A(u2__abc_52155_new_n13331_), .B(u2__abc_52155_new_n6290_), .Y(u2__abc_52155_new_n13334_));
OR2X2 OR2X2_2655 ( .A(u2__abc_52155_new_n13337_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13338_));
OR2X2 OR2X2_2656 ( .A(u2__abc_52155_new_n13336_), .B(u2__abc_52155_new_n13338_), .Y(u2__abc_52155_new_n13339_));
OR2X2 OR2X2_2657 ( .A(u2__abc_52155_new_n13343_), .B(u2__abc_52155_new_n13327_), .Y(u2__abc_52155_new_n13344_));
OR2X2 OR2X2_2658 ( .A(u2__abc_52155_new_n13348_), .B(u2__abc_52155_new_n13347_), .Y(u2__abc_52155_new_n13349_));
OR2X2 OR2X2_2659 ( .A(u2__abc_52155_new_n13350_), .B(u2__abc_52155_new_n6297_), .Y(u2__abc_52155_new_n13351_));
OR2X2 OR2X2_266 ( .A(\a[112] ), .B(\a[20] ), .Y(_abc_73687_new_n1230_));
OR2X2 OR2X2_2660 ( .A(u2__abc_52155_new_n13354_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13355_));
OR2X2 OR2X2_2661 ( .A(u2__abc_52155_new_n13353_), .B(u2__abc_52155_new_n13355_), .Y(u2__abc_52155_new_n13356_));
OR2X2 OR2X2_2662 ( .A(u2__abc_52155_new_n13360_), .B(u2__abc_52155_new_n13346_), .Y(u2__abc_52155_new_n13361_));
OR2X2 OR2X2_2663 ( .A(u2__abc_52155_new_n13328_), .B(u2__abc_52155_new_n6310_), .Y(u2__abc_52155_new_n13364_));
OR2X2 OR2X2_2664 ( .A(u2__abc_52155_new_n6729_), .B(u2__abc_52155_new_n13364_), .Y(u2__abc_52155_new_n13365_));
OR2X2 OR2X2_2665 ( .A(u2__abc_52155_new_n13366_), .B(u2__abc_52155_new_n6292_), .Y(u2__abc_52155_new_n13367_));
OR2X2 OR2X2_2666 ( .A(u2__abc_52155_new_n13371_), .B(u2__abc_52155_new_n13370_), .Y(u2__abc_52155_new_n13372_));
OR2X2 OR2X2_2667 ( .A(u2__abc_52155_new_n13372_), .B(u2__abc_52155_new_n6336_), .Y(u2__abc_52155_new_n13375_));
OR2X2 OR2X2_2668 ( .A(u2__abc_52155_new_n13378_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13379_));
OR2X2 OR2X2_2669 ( .A(u2__abc_52155_new_n13377_), .B(u2__abc_52155_new_n13379_), .Y(u2__abc_52155_new_n13380_));
OR2X2 OR2X2_267 ( .A(_abc_73687_new_n1170_), .B(\a[21] ), .Y(_abc_73687_new_n1231_));
OR2X2 OR2X2_2670 ( .A(u2__abc_52155_new_n13384_), .B(u2__abc_52155_new_n13363_), .Y(u2__abc_52155_new_n13385_));
OR2X2 OR2X2_2671 ( .A(u2__abc_52155_new_n13392_), .B(u2__abc_52155_new_n13389_), .Y(u2__abc_52155_new_n13393_));
OR2X2 OR2X2_2672 ( .A(u2__abc_52155_new_n13395_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13396_));
OR2X2 OR2X2_2673 ( .A(u2__abc_52155_new_n13394_), .B(u2__abc_52155_new_n13396_), .Y(u2__abc_52155_new_n13397_));
OR2X2 OR2X2_2674 ( .A(u2__abc_52155_new_n13401_), .B(u2__abc_52155_new_n13387_), .Y(u2__abc_52155_new_n13402_));
OR2X2 OR2X2_2675 ( .A(u2__abc_52155_new_n13406_), .B(u2__abc_52155_new_n6341_), .Y(u2__abc_52155_new_n13407_));
OR2X2 OR2X2_2676 ( .A(u2__abc_52155_new_n13408_), .B(u2__abc_52155_new_n6321_), .Y(u2__abc_52155_new_n13411_));
OR2X2 OR2X2_2677 ( .A(u2__abc_52155_new_n13414_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13415_));
OR2X2 OR2X2_2678 ( .A(u2__abc_52155_new_n13413_), .B(u2__abc_52155_new_n13415_), .Y(u2__abc_52155_new_n13416_));
OR2X2 OR2X2_2679 ( .A(u2__abc_52155_new_n13420_), .B(u2__abc_52155_new_n13404_), .Y(u2__abc_52155_new_n13421_));
OR2X2 OR2X2_268 ( .A(\a[112] ), .B(\a[21] ), .Y(_abc_73687_new_n1233_));
OR2X2 OR2X2_2680 ( .A(u2__abc_52155_new_n13425_), .B(u2__abc_52155_new_n13424_), .Y(u2__abc_52155_new_n13426_));
OR2X2 OR2X2_2681 ( .A(u2__abc_52155_new_n13427_), .B(u2__abc_52155_new_n6328_), .Y(u2__abc_52155_new_n13428_));
OR2X2 OR2X2_2682 ( .A(u2__abc_52155_new_n13431_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13432_));
OR2X2 OR2X2_2683 ( .A(u2__abc_52155_new_n13430_), .B(u2__abc_52155_new_n13432_), .Y(u2__abc_52155_new_n13433_));
OR2X2 OR2X2_2684 ( .A(u2__abc_52155_new_n13437_), .B(u2__abc_52155_new_n13423_), .Y(u2__abc_52155_new_n13438_));
OR2X2 OR2X2_2685 ( .A(u2__abc_52155_new_n13405_), .B(u2__abc_52155_new_n6341_), .Y(u2__abc_52155_new_n13443_));
OR2X2 OR2X2_2686 ( .A(u2__abc_52155_new_n6735_), .B(u2__abc_52155_new_n13443_), .Y(u2__abc_52155_new_n13444_));
OR2X2 OR2X2_2687 ( .A(u2__abc_52155_new_n13445_), .B(u2__abc_52155_new_n6326_), .Y(u2__abc_52155_new_n13446_));
OR2X2 OR2X2_2688 ( .A(u2__abc_52155_new_n13450_), .B(u2__abc_52155_new_n13449_), .Y(u2__abc_52155_new_n13451_));
OR2X2 OR2X2_2689 ( .A(u2__abc_52155_new_n13451_), .B(u2__abc_52155_new_n6227_), .Y(u2__abc_52155_new_n13454_));
OR2X2 OR2X2_269 ( .A(_abc_73687_new_n1170_), .B(\a[22] ), .Y(_abc_73687_new_n1234_));
OR2X2 OR2X2_2690 ( .A(u2__abc_52155_new_n13457_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13458_));
OR2X2 OR2X2_2691 ( .A(u2__abc_52155_new_n13456_), .B(u2__abc_52155_new_n13458_), .Y(u2__abc_52155_new_n13459_));
OR2X2 OR2X2_2692 ( .A(u2__abc_52155_new_n13463_), .B(u2__abc_52155_new_n13440_), .Y(u2__abc_52155_new_n13464_));
OR2X2 OR2X2_2693 ( .A(u2__abc_52155_new_n13468_), .B(u2__abc_52155_new_n13467_), .Y(u2__abc_52155_new_n13469_));
OR2X2 OR2X2_2694 ( .A(u2__abc_52155_new_n13470_), .B(u2__abc_52155_new_n6234_), .Y(u2__abc_52155_new_n13471_));
OR2X2 OR2X2_2695 ( .A(u2__abc_52155_new_n13474_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13475_));
OR2X2 OR2X2_2696 ( .A(u2__abc_52155_new_n13473_), .B(u2__abc_52155_new_n13475_), .Y(u2__abc_52155_new_n13476_));
OR2X2 OR2X2_2697 ( .A(u2__abc_52155_new_n13480_), .B(u2__abc_52155_new_n13466_), .Y(u2__abc_52155_new_n13481_));
OR2X2 OR2X2_2698 ( .A(u2__abc_52155_new_n13484_), .B(u2__abc_52155_new_n6229_), .Y(u2__abc_52155_new_n13485_));
OR2X2 OR2X2_2699 ( .A(u2__abc_52155_new_n13487_), .B(u2__abc_52155_new_n13486_), .Y(u2__abc_52155_new_n13488_));
OR2X2 OR2X2_27 ( .A(aNan), .B(sqrto_89_), .Y(_abc_73687_new_n869_));
OR2X2 OR2X2_270 ( .A(\a[112] ), .B(\a[22] ), .Y(_abc_73687_new_n1236_));
OR2X2 OR2X2_2700 ( .A(u2__abc_52155_new_n13488_), .B(u2__abc_52155_new_n6242_), .Y(u2__abc_52155_new_n13491_));
OR2X2 OR2X2_2701 ( .A(u2__abc_52155_new_n13494_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13495_));
OR2X2 OR2X2_2702 ( .A(u2__abc_52155_new_n13493_), .B(u2__abc_52155_new_n13495_), .Y(u2__abc_52155_new_n13496_));
OR2X2 OR2X2_2703 ( .A(u2__abc_52155_new_n13500_), .B(u2__abc_52155_new_n13483_), .Y(u2__abc_52155_new_n13501_));
OR2X2 OR2X2_2704 ( .A(u2__abc_52155_new_n13505_), .B(u2__abc_52155_new_n13504_), .Y(u2__abc_52155_new_n13506_));
OR2X2 OR2X2_2705 ( .A(u2__abc_52155_new_n13507_), .B(u2__abc_52155_new_n6249_), .Y(u2__abc_52155_new_n13508_));
OR2X2 OR2X2_2706 ( .A(u2__abc_52155_new_n13511_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13512_));
OR2X2 OR2X2_2707 ( .A(u2__abc_52155_new_n13510_), .B(u2__abc_52155_new_n13512_), .Y(u2__abc_52155_new_n13513_));
OR2X2 OR2X2_2708 ( .A(u2__abc_52155_new_n13517_), .B(u2__abc_52155_new_n13503_), .Y(u2__abc_52155_new_n13518_));
OR2X2 OR2X2_2709 ( .A(u2__abc_52155_new_n13522_), .B(u2__abc_52155_new_n6244_), .Y(u2__abc_52155_new_n13523_));
OR2X2 OR2X2_271 ( .A(_abc_73687_new_n1170_), .B(\a[23] ), .Y(_abc_73687_new_n1237_));
OR2X2 OR2X2_2710 ( .A(u2__abc_52155_new_n13521_), .B(u2__abc_52155_new_n13523_), .Y(u2__abc_52155_new_n13524_));
OR2X2 OR2X2_2711 ( .A(u2__abc_52155_new_n13525_), .B(u2__abc_52155_new_n13524_), .Y(u2__abc_52155_new_n13526_));
OR2X2 OR2X2_2712 ( .A(u2__abc_52155_new_n13526_), .B(u2__abc_52155_new_n6273_), .Y(u2__abc_52155_new_n13529_));
OR2X2 OR2X2_2713 ( .A(u2__abc_52155_new_n13532_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13533_));
OR2X2 OR2X2_2714 ( .A(u2__abc_52155_new_n13531_), .B(u2__abc_52155_new_n13533_), .Y(u2__abc_52155_new_n13534_));
OR2X2 OR2X2_2715 ( .A(u2__abc_52155_new_n13538_), .B(u2__abc_52155_new_n13520_), .Y(u2__abc_52155_new_n13539_));
OR2X2 OR2X2_2716 ( .A(u2__abc_52155_new_n13546_), .B(u2__abc_52155_new_n13543_), .Y(u2__abc_52155_new_n13547_));
OR2X2 OR2X2_2717 ( .A(u2__abc_52155_new_n13549_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13550_));
OR2X2 OR2X2_2718 ( .A(u2__abc_52155_new_n13548_), .B(u2__abc_52155_new_n13550_), .Y(u2__abc_52155_new_n13551_));
OR2X2 OR2X2_2719 ( .A(u2__abc_52155_new_n13555_), .B(u2__abc_52155_new_n13541_), .Y(u2__abc_52155_new_n13556_));
OR2X2 OR2X2_272 ( .A(\a[112] ), .B(\a[23] ), .Y(_abc_73687_new_n1239_));
OR2X2 OR2X2_2720 ( .A(u2__abc_52155_new_n13560_), .B(u2__abc_52155_new_n6278_), .Y(u2__abc_52155_new_n13561_));
OR2X2 OR2X2_2721 ( .A(u2__abc_52155_new_n13562_), .B(u2__abc_52155_new_n6258_), .Y(u2__abc_52155_new_n13565_));
OR2X2 OR2X2_2722 ( .A(u2__abc_52155_new_n13568_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13569_));
OR2X2 OR2X2_2723 ( .A(u2__abc_52155_new_n13567_), .B(u2__abc_52155_new_n13569_), .Y(u2__abc_52155_new_n13570_));
OR2X2 OR2X2_2724 ( .A(u2__abc_52155_new_n13574_), .B(u2__abc_52155_new_n13558_), .Y(u2__abc_52155_new_n13575_));
OR2X2 OR2X2_2725 ( .A(u2__abc_52155_new_n13579_), .B(u2__abc_52155_new_n13578_), .Y(u2__abc_52155_new_n13580_));
OR2X2 OR2X2_2726 ( .A(u2__abc_52155_new_n13581_), .B(u2__abc_52155_new_n6265_), .Y(u2__abc_52155_new_n13582_));
OR2X2 OR2X2_2727 ( .A(u2__abc_52155_new_n13585_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13586_));
OR2X2 OR2X2_2728 ( .A(u2__abc_52155_new_n13584_), .B(u2__abc_52155_new_n13586_), .Y(u2__abc_52155_new_n13587_));
OR2X2 OR2X2_2729 ( .A(u2__abc_52155_new_n13591_), .B(u2__abc_52155_new_n13577_), .Y(u2__abc_52155_new_n13592_));
OR2X2 OR2X2_273 ( .A(_abc_73687_new_n1170_), .B(\a[24] ), .Y(_abc_73687_new_n1240_));
OR2X2 OR2X2_2730 ( .A(u2__abc_52155_new_n13559_), .B(u2__abc_52155_new_n6278_), .Y(u2__abc_52155_new_n13599_));
OR2X2 OR2X2_2731 ( .A(u2__abc_52155_new_n6755_), .B(u2__abc_52155_new_n13599_), .Y(u2__abc_52155_new_n13600_));
OR2X2 OR2X2_2732 ( .A(u2__abc_52155_new_n13601_), .B(u2__abc_52155_new_n6260_), .Y(u2__abc_52155_new_n13602_));
OR2X2 OR2X2_2733 ( .A(u2__abc_52155_new_n13608_), .B(u2__abc_52155_new_n13607_), .Y(u2__abc_52155_new_n13609_));
OR2X2 OR2X2_2734 ( .A(u2__abc_52155_new_n13609_), .B(u2__abc_52155_new_n6163_), .Y(u2__abc_52155_new_n13612_));
OR2X2 OR2X2_2735 ( .A(u2__abc_52155_new_n13615_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13616_));
OR2X2 OR2X2_2736 ( .A(u2__abc_52155_new_n13614_), .B(u2__abc_52155_new_n13616_), .Y(u2__abc_52155_new_n13617_));
OR2X2 OR2X2_2737 ( .A(u2__abc_52155_new_n13621_), .B(u2__abc_52155_new_n13594_), .Y(u2__abc_52155_new_n13622_));
OR2X2 OR2X2_2738 ( .A(u2__abc_52155_new_n13626_), .B(u2__abc_52155_new_n13625_), .Y(u2__abc_52155_new_n13627_));
OR2X2 OR2X2_2739 ( .A(u2__abc_52155_new_n13628_), .B(u2__abc_52155_new_n6170_), .Y(u2__abc_52155_new_n13629_));
OR2X2 OR2X2_274 ( .A(\a[112] ), .B(\a[24] ), .Y(_abc_73687_new_n1242_));
OR2X2 OR2X2_2740 ( .A(u2__abc_52155_new_n13632_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13633_));
OR2X2 OR2X2_2741 ( .A(u2__abc_52155_new_n13631_), .B(u2__abc_52155_new_n13633_), .Y(u2__abc_52155_new_n13634_));
OR2X2 OR2X2_2742 ( .A(u2__abc_52155_new_n13638_), .B(u2__abc_52155_new_n13624_), .Y(u2__abc_52155_new_n13639_));
OR2X2 OR2X2_2743 ( .A(u2__abc_52155_new_n13642_), .B(u2__abc_52155_new_n6165_), .Y(u2__abc_52155_new_n13643_));
OR2X2 OR2X2_2744 ( .A(u2__abc_52155_new_n13645_), .B(u2__abc_52155_new_n13644_), .Y(u2__abc_52155_new_n13646_));
OR2X2 OR2X2_2745 ( .A(u2__abc_52155_new_n13646_), .B(u2__abc_52155_new_n6178_), .Y(u2__abc_52155_new_n13649_));
OR2X2 OR2X2_2746 ( .A(u2__abc_52155_new_n13652_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13653_));
OR2X2 OR2X2_2747 ( .A(u2__abc_52155_new_n13651_), .B(u2__abc_52155_new_n13653_), .Y(u2__abc_52155_new_n13654_));
OR2X2 OR2X2_2748 ( .A(u2__abc_52155_new_n13658_), .B(u2__abc_52155_new_n13641_), .Y(u2__abc_52155_new_n13659_));
OR2X2 OR2X2_2749 ( .A(u2__abc_52155_new_n13663_), .B(u2__abc_52155_new_n13662_), .Y(u2__abc_52155_new_n13664_));
OR2X2 OR2X2_275 ( .A(_abc_73687_new_n1170_), .B(\a[25] ), .Y(_abc_73687_new_n1243_));
OR2X2 OR2X2_2750 ( .A(u2__abc_52155_new_n13665_), .B(u2__abc_52155_new_n6185_), .Y(u2__abc_52155_new_n13666_));
OR2X2 OR2X2_2751 ( .A(u2__abc_52155_new_n13669_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13670_));
OR2X2 OR2X2_2752 ( .A(u2__abc_52155_new_n13668_), .B(u2__abc_52155_new_n13670_), .Y(u2__abc_52155_new_n13671_));
OR2X2 OR2X2_2753 ( .A(u2__abc_52155_new_n13675_), .B(u2__abc_52155_new_n13661_), .Y(u2__abc_52155_new_n13676_));
OR2X2 OR2X2_2754 ( .A(u2__abc_52155_new_n13680_), .B(u2__abc_52155_new_n6180_), .Y(u2__abc_52155_new_n13681_));
OR2X2 OR2X2_2755 ( .A(u2__abc_52155_new_n13679_), .B(u2__abc_52155_new_n13681_), .Y(u2__abc_52155_new_n13682_));
OR2X2 OR2X2_2756 ( .A(u2__abc_52155_new_n13683_), .B(u2__abc_52155_new_n13682_), .Y(u2__abc_52155_new_n13684_));
OR2X2 OR2X2_2757 ( .A(u2__abc_52155_new_n13684_), .B(u2__abc_52155_new_n6216_), .Y(u2__abc_52155_new_n13687_));
OR2X2 OR2X2_2758 ( .A(u2__abc_52155_new_n13690_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13691_));
OR2X2 OR2X2_2759 ( .A(u2__abc_52155_new_n13689_), .B(u2__abc_52155_new_n13691_), .Y(u2__abc_52155_new_n13692_));
OR2X2 OR2X2_276 ( .A(\a[112] ), .B(\a[25] ), .Y(_abc_73687_new_n1245_));
OR2X2 OR2X2_2760 ( .A(u2__abc_52155_new_n13696_), .B(u2__abc_52155_new_n13678_), .Y(u2__abc_52155_new_n13697_));
OR2X2 OR2X2_2761 ( .A(u2__abc_52155_new_n13701_), .B(u2__abc_52155_new_n6209_), .Y(u2__abc_52155_new_n13704_));
OR2X2 OR2X2_2762 ( .A(u2__abc_52155_new_n13707_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13708_));
OR2X2 OR2X2_2763 ( .A(u2__abc_52155_new_n13706_), .B(u2__abc_52155_new_n13708_), .Y(u2__abc_52155_new_n13709_));
OR2X2 OR2X2_2764 ( .A(u2__abc_52155_new_n13713_), .B(u2__abc_52155_new_n13699_), .Y(u2__abc_52155_new_n13714_));
OR2X2 OR2X2_2765 ( .A(u2__abc_52155_new_n13718_), .B(u2__abc_52155_new_n6194_), .Y(u2__abc_52155_new_n13721_));
OR2X2 OR2X2_2766 ( .A(u2__abc_52155_new_n13724_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13725_));
OR2X2 OR2X2_2767 ( .A(u2__abc_52155_new_n13723_), .B(u2__abc_52155_new_n13725_), .Y(u2__abc_52155_new_n13726_));
OR2X2 OR2X2_2768 ( .A(u2__abc_52155_new_n13730_), .B(u2__abc_52155_new_n13716_), .Y(u2__abc_52155_new_n13731_));
OR2X2 OR2X2_2769 ( .A(u2__abc_52155_new_n13735_), .B(u2__abc_52155_new_n13734_), .Y(u2__abc_52155_new_n13736_));
OR2X2 OR2X2_277 ( .A(_abc_73687_new_n1170_), .B(\a[26] ), .Y(_abc_73687_new_n1246_));
OR2X2 OR2X2_2770 ( .A(u2__abc_52155_new_n13737_), .B(u2__abc_52155_new_n6201_), .Y(u2__abc_52155_new_n13738_));
OR2X2 OR2X2_2771 ( .A(u2__abc_52155_new_n13741_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13742_));
OR2X2 OR2X2_2772 ( .A(u2__abc_52155_new_n13740_), .B(u2__abc_52155_new_n13742_), .Y(u2__abc_52155_new_n13743_));
OR2X2 OR2X2_2773 ( .A(u2__abc_52155_new_n13747_), .B(u2__abc_52155_new_n13733_), .Y(u2__abc_52155_new_n13748_));
OR2X2 OR2X2_2774 ( .A(u2__abc_52155_new_n13752_), .B(u2__abc_52155_new_n6204_), .Y(u2__abc_52155_new_n13753_));
OR2X2 OR2X2_2775 ( .A(u2__abc_52155_new_n13755_), .B(u2__abc_52155_new_n6196_), .Y(u2__abc_52155_new_n13756_));
OR2X2 OR2X2_2776 ( .A(u2__abc_52155_new_n13754_), .B(u2__abc_52155_new_n13756_), .Y(u2__abc_52155_new_n13757_));
OR2X2 OR2X2_2777 ( .A(u2__abc_52155_new_n13751_), .B(u2__abc_52155_new_n13757_), .Y(u2__abc_52155_new_n13758_));
OR2X2 OR2X2_2778 ( .A(u2__abc_52155_new_n13759_), .B(u2__abc_52155_new_n13758_), .Y(u2__abc_52155_new_n13760_));
OR2X2 OR2X2_2779 ( .A(u2__abc_52155_new_n13760_), .B(u2__abc_52155_new_n6115_), .Y(u2__abc_52155_new_n13763_));
OR2X2 OR2X2_278 ( .A(\a[112] ), .B(\a[26] ), .Y(_abc_73687_new_n1248_));
OR2X2 OR2X2_2780 ( .A(u2__abc_52155_new_n13766_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13767_));
OR2X2 OR2X2_2781 ( .A(u2__abc_52155_new_n13765_), .B(u2__abc_52155_new_n13767_), .Y(u2__abc_52155_new_n13768_));
OR2X2 OR2X2_2782 ( .A(u2__abc_52155_new_n13772_), .B(u2__abc_52155_new_n13750_), .Y(u2__abc_52155_new_n13773_));
OR2X2 OR2X2_2783 ( .A(u2__abc_52155_new_n13780_), .B(u2__abc_52155_new_n13777_), .Y(u2__abc_52155_new_n13781_));
OR2X2 OR2X2_2784 ( .A(u2__abc_52155_new_n13783_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13784_));
OR2X2 OR2X2_2785 ( .A(u2__abc_52155_new_n13782_), .B(u2__abc_52155_new_n13784_), .Y(u2__abc_52155_new_n13785_));
OR2X2 OR2X2_2786 ( .A(u2__abc_52155_new_n13789_), .B(u2__abc_52155_new_n13775_), .Y(u2__abc_52155_new_n13790_));
OR2X2 OR2X2_2787 ( .A(u2__abc_52155_new_n13794_), .B(u2__abc_52155_new_n6120_), .Y(u2__abc_52155_new_n13795_));
OR2X2 OR2X2_2788 ( .A(u2__abc_52155_new_n13796_), .B(u2__abc_52155_new_n6100_), .Y(u2__abc_52155_new_n13799_));
OR2X2 OR2X2_2789 ( .A(u2__abc_52155_new_n13802_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13803_));
OR2X2 OR2X2_279 ( .A(_abc_73687_new_n1170_), .B(\a[27] ), .Y(_abc_73687_new_n1249_));
OR2X2 OR2X2_2790 ( .A(u2__abc_52155_new_n13801_), .B(u2__abc_52155_new_n13803_), .Y(u2__abc_52155_new_n13804_));
OR2X2 OR2X2_2791 ( .A(u2__abc_52155_new_n13808_), .B(u2__abc_52155_new_n13792_), .Y(u2__abc_52155_new_n13809_));
OR2X2 OR2X2_2792 ( .A(u2__abc_52155_new_n13813_), .B(u2__abc_52155_new_n13812_), .Y(u2__abc_52155_new_n13814_));
OR2X2 OR2X2_2793 ( .A(u2__abc_52155_new_n13815_), .B(u2__abc_52155_new_n6107_), .Y(u2__abc_52155_new_n13816_));
OR2X2 OR2X2_2794 ( .A(u2__abc_52155_new_n13819_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13820_));
OR2X2 OR2X2_2795 ( .A(u2__abc_52155_new_n13818_), .B(u2__abc_52155_new_n13820_), .Y(u2__abc_52155_new_n13821_));
OR2X2 OR2X2_2796 ( .A(u2__abc_52155_new_n13825_), .B(u2__abc_52155_new_n13811_), .Y(u2__abc_52155_new_n13826_));
OR2X2 OR2X2_2797 ( .A(u2__abc_52155_new_n13793_), .B(u2__abc_52155_new_n6120_), .Y(u2__abc_52155_new_n13830_));
OR2X2 OR2X2_2798 ( .A(u2__abc_52155_new_n13829_), .B(u2__abc_52155_new_n13830_), .Y(u2__abc_52155_new_n13831_));
OR2X2 OR2X2_2799 ( .A(u2__abc_52155_new_n13832_), .B(u2__abc_52155_new_n6102_), .Y(u2__abc_52155_new_n13833_));
OR2X2 OR2X2_28 ( .A(_abc_73687_new_n753_), .B(\a[13] ), .Y(_abc_73687_new_n870_));
OR2X2 OR2X2_280 ( .A(\a[112] ), .B(\a[27] ), .Y(_abc_73687_new_n1251_));
OR2X2 OR2X2_2800 ( .A(u2__abc_52155_new_n13837_), .B(u2__abc_52155_new_n13836_), .Y(u2__abc_52155_new_n13838_));
OR2X2 OR2X2_2801 ( .A(u2__abc_52155_new_n13838_), .B(u2__abc_52155_new_n6146_), .Y(u2__abc_52155_new_n13841_));
OR2X2 OR2X2_2802 ( .A(u2__abc_52155_new_n13844_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13845_));
OR2X2 OR2X2_2803 ( .A(u2__abc_52155_new_n13843_), .B(u2__abc_52155_new_n13845_), .Y(u2__abc_52155_new_n13846_));
OR2X2 OR2X2_2804 ( .A(u2__abc_52155_new_n13850_), .B(u2__abc_52155_new_n13828_), .Y(u2__abc_52155_new_n13851_));
OR2X2 OR2X2_2805 ( .A(u2__abc_52155_new_n13858_), .B(u2__abc_52155_new_n13855_), .Y(u2__abc_52155_new_n13859_));
OR2X2 OR2X2_2806 ( .A(u2__abc_52155_new_n13861_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13862_));
OR2X2 OR2X2_2807 ( .A(u2__abc_52155_new_n13860_), .B(u2__abc_52155_new_n13862_), .Y(u2__abc_52155_new_n13863_));
OR2X2 OR2X2_2808 ( .A(u2__abc_52155_new_n13867_), .B(u2__abc_52155_new_n13853_), .Y(u2__abc_52155_new_n13868_));
OR2X2 OR2X2_2809 ( .A(u2__abc_52155_new_n13872_), .B(u2__abc_52155_new_n6151_), .Y(u2__abc_52155_new_n13873_));
OR2X2 OR2X2_281 ( .A(_abc_73687_new_n1170_), .B(\a[28] ), .Y(_abc_73687_new_n1252_));
OR2X2 OR2X2_2810 ( .A(u2__abc_52155_new_n13874_), .B(u2__abc_52155_new_n6131_), .Y(u2__abc_52155_new_n13877_));
OR2X2 OR2X2_2811 ( .A(u2__abc_52155_new_n13880_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13881_));
OR2X2 OR2X2_2812 ( .A(u2__abc_52155_new_n13879_), .B(u2__abc_52155_new_n13881_), .Y(u2__abc_52155_new_n13882_));
OR2X2 OR2X2_2813 ( .A(u2__abc_52155_new_n13886_), .B(u2__abc_52155_new_n13870_), .Y(u2__abc_52155_new_n13887_));
OR2X2 OR2X2_2814 ( .A(u2__abc_52155_new_n13891_), .B(u2__abc_52155_new_n13890_), .Y(u2__abc_52155_new_n13892_));
OR2X2 OR2X2_2815 ( .A(u2__abc_52155_new_n13893_), .B(u2__abc_52155_new_n6138_), .Y(u2__abc_52155_new_n13894_));
OR2X2 OR2X2_2816 ( .A(u2__abc_52155_new_n13897_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13898_));
OR2X2 OR2X2_2817 ( .A(u2__abc_52155_new_n13896_), .B(u2__abc_52155_new_n13898_), .Y(u2__abc_52155_new_n13899_));
OR2X2 OR2X2_2818 ( .A(u2__abc_52155_new_n13903_), .B(u2__abc_52155_new_n13889_), .Y(u2__abc_52155_new_n13904_));
OR2X2 OR2X2_2819 ( .A(u2__abc_52155_new_n13871_), .B(u2__abc_52155_new_n6151_), .Y(u2__abc_52155_new_n13916_));
OR2X2 OR2X2_282 ( .A(\a[112] ), .B(\a[28] ), .Y(_abc_73687_new_n1254_));
OR2X2 OR2X2_2820 ( .A(u2__abc_52155_new_n13915_), .B(u2__abc_52155_new_n13916_), .Y(u2__abc_52155_new_n13917_));
OR2X2 OR2X2_2821 ( .A(u2__abc_52155_new_n13918_), .B(u2__abc_52155_new_n6133_), .Y(u2__abc_52155_new_n13919_));
OR2X2 OR2X2_2822 ( .A(u2__abc_52155_new_n13927_), .B(u2__abc_52155_new_n13926_), .Y(u2__abc_52155_new_n13928_));
OR2X2 OR2X2_2823 ( .A(u2__abc_52155_new_n13928_), .B(u2__abc_52155_new_n6065_), .Y(u2__abc_52155_new_n13931_));
OR2X2 OR2X2_2824 ( .A(u2__abc_52155_new_n13934_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13935_));
OR2X2 OR2X2_2825 ( .A(u2__abc_52155_new_n13933_), .B(u2__abc_52155_new_n13935_), .Y(u2__abc_52155_new_n13936_));
OR2X2 OR2X2_2826 ( .A(u2__abc_52155_new_n13940_), .B(u2__abc_52155_new_n13906_), .Y(u2__abc_52155_new_n13941_));
OR2X2 OR2X2_2827 ( .A(u2__abc_52155_new_n13945_), .B(u2__abc_52155_new_n13944_), .Y(u2__abc_52155_new_n13946_));
OR2X2 OR2X2_2828 ( .A(u2__abc_52155_new_n13947_), .B(u2__abc_52155_new_n6072_), .Y(u2__abc_52155_new_n13948_));
OR2X2 OR2X2_2829 ( .A(u2__abc_52155_new_n13951_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13952_));
OR2X2 OR2X2_283 ( .A(_abc_73687_new_n1170_), .B(\a[29] ), .Y(_abc_73687_new_n1255_));
OR2X2 OR2X2_2830 ( .A(u2__abc_52155_new_n13950_), .B(u2__abc_52155_new_n13952_), .Y(u2__abc_52155_new_n13953_));
OR2X2 OR2X2_2831 ( .A(u2__abc_52155_new_n13957_), .B(u2__abc_52155_new_n13943_), .Y(u2__abc_52155_new_n13958_));
OR2X2 OR2X2_2832 ( .A(u2__abc_52155_new_n13961_), .B(u2__abc_52155_new_n6067_), .Y(u2__abc_52155_new_n13962_));
OR2X2 OR2X2_2833 ( .A(u2__abc_52155_new_n13964_), .B(u2__abc_52155_new_n13963_), .Y(u2__abc_52155_new_n13965_));
OR2X2 OR2X2_2834 ( .A(u2__abc_52155_new_n13965_), .B(u2__abc_52155_new_n6080_), .Y(u2__abc_52155_new_n13968_));
OR2X2 OR2X2_2835 ( .A(u2__abc_52155_new_n13971_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13972_));
OR2X2 OR2X2_2836 ( .A(u2__abc_52155_new_n13970_), .B(u2__abc_52155_new_n13972_), .Y(u2__abc_52155_new_n13973_));
OR2X2 OR2X2_2837 ( .A(u2__abc_52155_new_n13977_), .B(u2__abc_52155_new_n13960_), .Y(u2__abc_52155_new_n13978_));
OR2X2 OR2X2_2838 ( .A(u2__abc_52155_new_n13982_), .B(u2__abc_52155_new_n13981_), .Y(u2__abc_52155_new_n13983_));
OR2X2 OR2X2_2839 ( .A(u2__abc_52155_new_n13984_), .B(u2__abc_52155_new_n6087_), .Y(u2__abc_52155_new_n13985_));
OR2X2 OR2X2_284 ( .A(\a[112] ), .B(\a[29] ), .Y(_abc_73687_new_n1257_));
OR2X2 OR2X2_2840 ( .A(u2__abc_52155_new_n13988_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n13989_));
OR2X2 OR2X2_2841 ( .A(u2__abc_52155_new_n13987_), .B(u2__abc_52155_new_n13989_), .Y(u2__abc_52155_new_n13990_));
OR2X2 OR2X2_2842 ( .A(u2__abc_52155_new_n13994_), .B(u2__abc_52155_new_n13980_), .Y(u2__abc_52155_new_n13995_));
OR2X2 OR2X2_2843 ( .A(u2__abc_52155_new_n13999_), .B(u2__abc_52155_new_n6082_), .Y(u2__abc_52155_new_n14000_));
OR2X2 OR2X2_2844 ( .A(u2__abc_52155_new_n13998_), .B(u2__abc_52155_new_n14000_), .Y(u2__abc_52155_new_n14001_));
OR2X2 OR2X2_2845 ( .A(u2__abc_52155_new_n14002_), .B(u2__abc_52155_new_n14001_), .Y(u2__abc_52155_new_n14003_));
OR2X2 OR2X2_2846 ( .A(u2__abc_52155_new_n14003_), .B(u2__abc_52155_new_n6049_), .Y(u2__abc_52155_new_n14006_));
OR2X2 OR2X2_2847 ( .A(u2__abc_52155_new_n14009_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14010_));
OR2X2 OR2X2_2848 ( .A(u2__abc_52155_new_n14008_), .B(u2__abc_52155_new_n14010_), .Y(u2__abc_52155_new_n14011_));
OR2X2 OR2X2_2849 ( .A(u2__abc_52155_new_n14015_), .B(u2__abc_52155_new_n13997_), .Y(u2__abc_52155_new_n14016_));
OR2X2 OR2X2_285 ( .A(_abc_73687_new_n1170_), .B(\a[30] ), .Y(_abc_73687_new_n1258_));
OR2X2 OR2X2_2850 ( .A(u2__abc_52155_new_n14023_), .B(u2__abc_52155_new_n14020_), .Y(u2__abc_52155_new_n14024_));
OR2X2 OR2X2_2851 ( .A(u2__abc_52155_new_n14026_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14027_));
OR2X2 OR2X2_2852 ( .A(u2__abc_52155_new_n14025_), .B(u2__abc_52155_new_n14027_), .Y(u2__abc_52155_new_n14028_));
OR2X2 OR2X2_2853 ( .A(u2__abc_52155_new_n14032_), .B(u2__abc_52155_new_n14018_), .Y(u2__abc_52155_new_n14033_));
OR2X2 OR2X2_2854 ( .A(u2__abc_52155_new_n14037_), .B(u2__abc_52155_new_n6054_), .Y(u2__abc_52155_new_n14038_));
OR2X2 OR2X2_2855 ( .A(u2__abc_52155_new_n14039_), .B(u2__abc_52155_new_n6034_), .Y(u2__abc_52155_new_n14042_));
OR2X2 OR2X2_2856 ( .A(u2__abc_52155_new_n14045_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14046_));
OR2X2 OR2X2_2857 ( .A(u2__abc_52155_new_n14044_), .B(u2__abc_52155_new_n14046_), .Y(u2__abc_52155_new_n14047_));
OR2X2 OR2X2_2858 ( .A(u2__abc_52155_new_n14051_), .B(u2__abc_52155_new_n14035_), .Y(u2__abc_52155_new_n14052_));
OR2X2 OR2X2_2859 ( .A(u2__abc_52155_new_n14056_), .B(u2__abc_52155_new_n14055_), .Y(u2__abc_52155_new_n14057_));
OR2X2 OR2X2_286 ( .A(\a[112] ), .B(\a[30] ), .Y(_abc_73687_new_n1260_));
OR2X2 OR2X2_2860 ( .A(u2__abc_52155_new_n14058_), .B(u2__abc_52155_new_n6041_), .Y(u2__abc_52155_new_n14059_));
OR2X2 OR2X2_2861 ( .A(u2__abc_52155_new_n14062_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14063_));
OR2X2 OR2X2_2862 ( .A(u2__abc_52155_new_n14061_), .B(u2__abc_52155_new_n14063_), .Y(u2__abc_52155_new_n14064_));
OR2X2 OR2X2_2863 ( .A(u2__abc_52155_new_n14068_), .B(u2__abc_52155_new_n14054_), .Y(u2__abc_52155_new_n14069_));
OR2X2 OR2X2_2864 ( .A(u2__abc_52155_new_n14036_), .B(u2__abc_52155_new_n6054_), .Y(u2__abc_52155_new_n14074_));
OR2X2 OR2X2_2865 ( .A(u2__abc_52155_new_n6784_), .B(u2__abc_52155_new_n14074_), .Y(u2__abc_52155_new_n14075_));
OR2X2 OR2X2_2866 ( .A(u2__abc_52155_new_n14076_), .B(u2__abc_52155_new_n6036_), .Y(u2__abc_52155_new_n14077_));
OR2X2 OR2X2_2867 ( .A(u2__abc_52155_new_n14081_), .B(u2__abc_52155_new_n14080_), .Y(u2__abc_52155_new_n14082_));
OR2X2 OR2X2_2868 ( .A(u2__abc_52155_new_n14082_), .B(u2__abc_52155_new_n5971_), .Y(u2__abc_52155_new_n14085_));
OR2X2 OR2X2_2869 ( .A(u2__abc_52155_new_n14088_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14089_));
OR2X2 OR2X2_287 ( .A(_abc_73687_new_n1170_), .B(\a[31] ), .Y(_abc_73687_new_n1261_));
OR2X2 OR2X2_2870 ( .A(u2__abc_52155_new_n14087_), .B(u2__abc_52155_new_n14089_), .Y(u2__abc_52155_new_n14090_));
OR2X2 OR2X2_2871 ( .A(u2__abc_52155_new_n14094_), .B(u2__abc_52155_new_n14071_), .Y(u2__abc_52155_new_n14095_));
OR2X2 OR2X2_2872 ( .A(u2__abc_52155_new_n14099_), .B(u2__abc_52155_new_n14098_), .Y(u2__abc_52155_new_n14100_));
OR2X2 OR2X2_2873 ( .A(u2__abc_52155_new_n14101_), .B(u2__abc_52155_new_n5978_), .Y(u2__abc_52155_new_n14102_));
OR2X2 OR2X2_2874 ( .A(u2__abc_52155_new_n14105_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14106_));
OR2X2 OR2X2_2875 ( .A(u2__abc_52155_new_n14104_), .B(u2__abc_52155_new_n14106_), .Y(u2__abc_52155_new_n14107_));
OR2X2 OR2X2_2876 ( .A(u2__abc_52155_new_n14111_), .B(u2__abc_52155_new_n14097_), .Y(u2__abc_52155_new_n14112_));
OR2X2 OR2X2_2877 ( .A(u2__abc_52155_new_n14115_), .B(u2__abc_52155_new_n5973_), .Y(u2__abc_52155_new_n14116_));
OR2X2 OR2X2_2878 ( .A(u2__abc_52155_new_n14118_), .B(u2__abc_52155_new_n14117_), .Y(u2__abc_52155_new_n14119_));
OR2X2 OR2X2_2879 ( .A(u2__abc_52155_new_n14119_), .B(u2__abc_52155_new_n5986_), .Y(u2__abc_52155_new_n14122_));
OR2X2 OR2X2_288 ( .A(\a[112] ), .B(\a[31] ), .Y(_abc_73687_new_n1263_));
OR2X2 OR2X2_2880 ( .A(u2__abc_52155_new_n14125_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14126_));
OR2X2 OR2X2_2881 ( .A(u2__abc_52155_new_n14124_), .B(u2__abc_52155_new_n14126_), .Y(u2__abc_52155_new_n14127_));
OR2X2 OR2X2_2882 ( .A(u2__abc_52155_new_n14131_), .B(u2__abc_52155_new_n14114_), .Y(u2__abc_52155_new_n14132_));
OR2X2 OR2X2_2883 ( .A(u2__abc_52155_new_n14136_), .B(u2__abc_52155_new_n14135_), .Y(u2__abc_52155_new_n14137_));
OR2X2 OR2X2_2884 ( .A(u2__abc_52155_new_n14138_), .B(u2__abc_52155_new_n5993_), .Y(u2__abc_52155_new_n14139_));
OR2X2 OR2X2_2885 ( .A(u2__abc_52155_new_n14142_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14143_));
OR2X2 OR2X2_2886 ( .A(u2__abc_52155_new_n14141_), .B(u2__abc_52155_new_n14143_), .Y(u2__abc_52155_new_n14144_));
OR2X2 OR2X2_2887 ( .A(u2__abc_52155_new_n14148_), .B(u2__abc_52155_new_n14134_), .Y(u2__abc_52155_new_n14149_));
OR2X2 OR2X2_2888 ( .A(u2__abc_52155_new_n14153_), .B(u2__abc_52155_new_n5988_), .Y(u2__abc_52155_new_n14154_));
OR2X2 OR2X2_2889 ( .A(u2__abc_52155_new_n14152_), .B(u2__abc_52155_new_n14154_), .Y(u2__abc_52155_new_n14155_));
OR2X2 OR2X2_289 ( .A(_abc_73687_new_n1170_), .B(\a[32] ), .Y(_abc_73687_new_n1264_));
OR2X2 OR2X2_2890 ( .A(u2__abc_52155_new_n14156_), .B(u2__abc_52155_new_n14155_), .Y(u2__abc_52155_new_n14157_));
OR2X2 OR2X2_2891 ( .A(u2__abc_52155_new_n14157_), .B(u2__abc_52155_new_n6017_), .Y(u2__abc_52155_new_n14160_));
OR2X2 OR2X2_2892 ( .A(u2__abc_52155_new_n14163_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14164_));
OR2X2 OR2X2_2893 ( .A(u2__abc_52155_new_n14162_), .B(u2__abc_52155_new_n14164_), .Y(u2__abc_52155_new_n14165_));
OR2X2 OR2X2_2894 ( .A(u2__abc_52155_new_n14169_), .B(u2__abc_52155_new_n14151_), .Y(u2__abc_52155_new_n14170_));
OR2X2 OR2X2_2895 ( .A(u2__abc_52155_new_n14177_), .B(u2__abc_52155_new_n14174_), .Y(u2__abc_52155_new_n14178_));
OR2X2 OR2X2_2896 ( .A(u2__abc_52155_new_n14180_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14181_));
OR2X2 OR2X2_2897 ( .A(u2__abc_52155_new_n14179_), .B(u2__abc_52155_new_n14181_), .Y(u2__abc_52155_new_n14182_));
OR2X2 OR2X2_2898 ( .A(u2__abc_52155_new_n14186_), .B(u2__abc_52155_new_n14172_), .Y(u2__abc_52155_new_n14187_));
OR2X2 OR2X2_2899 ( .A(u2__abc_52155_new_n14191_), .B(u2__abc_52155_new_n6022_), .Y(u2__abc_52155_new_n14192_));
OR2X2 OR2X2_29 ( .A(aNan), .B(sqrto_90_), .Y(_abc_73687_new_n872_));
OR2X2 OR2X2_290 ( .A(\a[112] ), .B(\a[32] ), .Y(_abc_73687_new_n1266_));
OR2X2 OR2X2_2900 ( .A(u2__abc_52155_new_n14193_), .B(u2__abc_52155_new_n6002_), .Y(u2__abc_52155_new_n14196_));
OR2X2 OR2X2_2901 ( .A(u2__abc_52155_new_n14199_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14200_));
OR2X2 OR2X2_2902 ( .A(u2__abc_52155_new_n14198_), .B(u2__abc_52155_new_n14200_), .Y(u2__abc_52155_new_n14201_));
OR2X2 OR2X2_2903 ( .A(u2__abc_52155_new_n14205_), .B(u2__abc_52155_new_n14189_), .Y(u2__abc_52155_new_n14206_));
OR2X2 OR2X2_2904 ( .A(u2__abc_52155_new_n14210_), .B(u2__abc_52155_new_n14209_), .Y(u2__abc_52155_new_n14211_));
OR2X2 OR2X2_2905 ( .A(u2__abc_52155_new_n14212_), .B(u2__abc_52155_new_n6009_), .Y(u2__abc_52155_new_n14213_));
OR2X2 OR2X2_2906 ( .A(u2__abc_52155_new_n14216_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14217_));
OR2X2 OR2X2_2907 ( .A(u2__abc_52155_new_n14215_), .B(u2__abc_52155_new_n14217_), .Y(u2__abc_52155_new_n14218_));
OR2X2 OR2X2_2908 ( .A(u2__abc_52155_new_n14222_), .B(u2__abc_52155_new_n14208_), .Y(u2__abc_52155_new_n14223_));
OR2X2 OR2X2_2909 ( .A(u2__abc_52155_new_n14190_), .B(u2__abc_52155_new_n6022_), .Y(u2__abc_52155_new_n14230_));
OR2X2 OR2X2_291 ( .A(_abc_73687_new_n1170_), .B(\a[33] ), .Y(_abc_73687_new_n1267_));
OR2X2 OR2X2_2910 ( .A(u2__abc_52155_new_n6801_), .B(u2__abc_52155_new_n14230_), .Y(u2__abc_52155_new_n14231_));
OR2X2 OR2X2_2911 ( .A(u2__abc_52155_new_n14232_), .B(u2__abc_52155_new_n6004_), .Y(u2__abc_52155_new_n14233_));
OR2X2 OR2X2_2912 ( .A(u2__abc_52155_new_n14239_), .B(u2__abc_52155_new_n14238_), .Y(u2__abc_52155_new_n14240_));
OR2X2 OR2X2_2913 ( .A(u2__abc_52155_new_n14240_), .B(u2__abc_52155_new_n5922_), .Y(u2__abc_52155_new_n14243_));
OR2X2 OR2X2_2914 ( .A(u2__abc_52155_new_n14246_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14247_));
OR2X2 OR2X2_2915 ( .A(u2__abc_52155_new_n14245_), .B(u2__abc_52155_new_n14247_), .Y(u2__abc_52155_new_n14248_));
OR2X2 OR2X2_2916 ( .A(u2__abc_52155_new_n14252_), .B(u2__abc_52155_new_n14225_), .Y(u2__abc_52155_new_n14253_));
OR2X2 OR2X2_2917 ( .A(u2__abc_52155_new_n14260_), .B(u2__abc_52155_new_n14257_), .Y(u2__abc_52155_new_n14261_));
OR2X2 OR2X2_2918 ( .A(u2__abc_52155_new_n14263_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14264_));
OR2X2 OR2X2_2919 ( .A(u2__abc_52155_new_n14262_), .B(u2__abc_52155_new_n14264_), .Y(u2__abc_52155_new_n14265_));
OR2X2 OR2X2_292 ( .A(\a[112] ), .B(\a[33] ), .Y(_abc_73687_new_n1269_));
OR2X2 OR2X2_2920 ( .A(u2__abc_52155_new_n14269_), .B(u2__abc_52155_new_n14255_), .Y(u2__abc_52155_new_n14270_));
OR2X2 OR2X2_2921 ( .A(u2__abc_52155_new_n14274_), .B(u2__abc_52155_new_n5927_), .Y(u2__abc_52155_new_n14275_));
OR2X2 OR2X2_2922 ( .A(u2__abc_52155_new_n14276_), .B(u2__abc_52155_new_n5907_), .Y(u2__abc_52155_new_n14279_));
OR2X2 OR2X2_2923 ( .A(u2__abc_52155_new_n14282_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14283_));
OR2X2 OR2X2_2924 ( .A(u2__abc_52155_new_n14281_), .B(u2__abc_52155_new_n14283_), .Y(u2__abc_52155_new_n14284_));
OR2X2 OR2X2_2925 ( .A(u2__abc_52155_new_n14288_), .B(u2__abc_52155_new_n14272_), .Y(u2__abc_52155_new_n14289_));
OR2X2 OR2X2_2926 ( .A(u2__abc_52155_new_n14293_), .B(u2__abc_52155_new_n14292_), .Y(u2__abc_52155_new_n14294_));
OR2X2 OR2X2_2927 ( .A(u2__abc_52155_new_n14295_), .B(u2__abc_52155_new_n5914_), .Y(u2__abc_52155_new_n14296_));
OR2X2 OR2X2_2928 ( .A(u2__abc_52155_new_n14299_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14300_));
OR2X2 OR2X2_2929 ( .A(u2__abc_52155_new_n14298_), .B(u2__abc_52155_new_n14300_), .Y(u2__abc_52155_new_n14301_));
OR2X2 OR2X2_293 ( .A(_abc_73687_new_n1170_), .B(\a[34] ), .Y(_abc_73687_new_n1270_));
OR2X2 OR2X2_2930 ( .A(u2__abc_52155_new_n14305_), .B(u2__abc_52155_new_n14291_), .Y(u2__abc_52155_new_n14306_));
OR2X2 OR2X2_2931 ( .A(u2__abc_52155_new_n14273_), .B(u2__abc_52155_new_n5927_), .Y(u2__abc_52155_new_n14309_));
OR2X2 OR2X2_2932 ( .A(u2__abc_52155_new_n6837_), .B(u2__abc_52155_new_n14309_), .Y(u2__abc_52155_new_n14310_));
OR2X2 OR2X2_2933 ( .A(u2__abc_52155_new_n14311_), .B(u2__abc_52155_new_n5909_), .Y(u2__abc_52155_new_n14312_));
OR2X2 OR2X2_2934 ( .A(u2__abc_52155_new_n14316_), .B(u2__abc_52155_new_n14315_), .Y(u2__abc_52155_new_n14317_));
OR2X2 OR2X2_2935 ( .A(u2__abc_52155_new_n14317_), .B(u2__abc_52155_new_n5953_), .Y(u2__abc_52155_new_n14320_));
OR2X2 OR2X2_2936 ( .A(u2__abc_52155_new_n14323_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14324_));
OR2X2 OR2X2_2937 ( .A(u2__abc_52155_new_n14322_), .B(u2__abc_52155_new_n14324_), .Y(u2__abc_52155_new_n14325_));
OR2X2 OR2X2_2938 ( .A(u2__abc_52155_new_n14329_), .B(u2__abc_52155_new_n14308_), .Y(u2__abc_52155_new_n14330_));
OR2X2 OR2X2_2939 ( .A(u2__abc_52155_new_n14337_), .B(u2__abc_52155_new_n14334_), .Y(u2__abc_52155_new_n14338_));
OR2X2 OR2X2_294 ( .A(\a[112] ), .B(\a[34] ), .Y(_abc_73687_new_n1272_));
OR2X2 OR2X2_2940 ( .A(u2__abc_52155_new_n14340_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14341_));
OR2X2 OR2X2_2941 ( .A(u2__abc_52155_new_n14339_), .B(u2__abc_52155_new_n14341_), .Y(u2__abc_52155_new_n14342_));
OR2X2 OR2X2_2942 ( .A(u2__abc_52155_new_n14346_), .B(u2__abc_52155_new_n14332_), .Y(u2__abc_52155_new_n14347_));
OR2X2 OR2X2_2943 ( .A(u2__abc_52155_new_n14351_), .B(u2__abc_52155_new_n5958_), .Y(u2__abc_52155_new_n14352_));
OR2X2 OR2X2_2944 ( .A(u2__abc_52155_new_n14353_), .B(u2__abc_52155_new_n5938_), .Y(u2__abc_52155_new_n14356_));
OR2X2 OR2X2_2945 ( .A(u2__abc_52155_new_n14359_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14360_));
OR2X2 OR2X2_2946 ( .A(u2__abc_52155_new_n14358_), .B(u2__abc_52155_new_n14360_), .Y(u2__abc_52155_new_n14361_));
OR2X2 OR2X2_2947 ( .A(u2__abc_52155_new_n14365_), .B(u2__abc_52155_new_n14349_), .Y(u2__abc_52155_new_n14366_));
OR2X2 OR2X2_2948 ( .A(u2__abc_52155_new_n14370_), .B(u2__abc_52155_new_n14369_), .Y(u2__abc_52155_new_n14371_));
OR2X2 OR2X2_2949 ( .A(u2__abc_52155_new_n14372_), .B(u2__abc_52155_new_n5945_), .Y(u2__abc_52155_new_n14373_));
OR2X2 OR2X2_295 ( .A(_abc_73687_new_n1170_), .B(\a[35] ), .Y(_abc_73687_new_n1273_));
OR2X2 OR2X2_2950 ( .A(u2__abc_52155_new_n14376_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14377_));
OR2X2 OR2X2_2951 ( .A(u2__abc_52155_new_n14375_), .B(u2__abc_52155_new_n14377_), .Y(u2__abc_52155_new_n14378_));
OR2X2 OR2X2_2952 ( .A(u2__abc_52155_new_n14382_), .B(u2__abc_52155_new_n14368_), .Y(u2__abc_52155_new_n14383_));
OR2X2 OR2X2_2953 ( .A(u2__abc_52155_new_n14350_), .B(u2__abc_52155_new_n5958_), .Y(u2__abc_52155_new_n14388_));
OR2X2 OR2X2_2954 ( .A(u2__abc_52155_new_n6844_), .B(u2__abc_52155_new_n14388_), .Y(u2__abc_52155_new_n14389_));
OR2X2 OR2X2_2955 ( .A(u2__abc_52155_new_n14390_), .B(u2__abc_52155_new_n5940_), .Y(u2__abc_52155_new_n14391_));
OR2X2 OR2X2_2956 ( .A(u2__abc_52155_new_n14396_), .B(u2__abc_52155_new_n14395_), .Y(u2__abc_52155_new_n14397_));
OR2X2 OR2X2_2957 ( .A(u2__abc_52155_new_n14397_), .B(u2__abc_52155_new_n5859_), .Y(u2__abc_52155_new_n14400_));
OR2X2 OR2X2_2958 ( .A(u2__abc_52155_new_n14403_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14404_));
OR2X2 OR2X2_2959 ( .A(u2__abc_52155_new_n14402_), .B(u2__abc_52155_new_n14404_), .Y(u2__abc_52155_new_n14405_));
OR2X2 OR2X2_296 ( .A(\a[112] ), .B(\a[35] ), .Y(_abc_73687_new_n1275_));
OR2X2 OR2X2_2960 ( .A(u2__abc_52155_new_n14409_), .B(u2__abc_52155_new_n14385_), .Y(u2__abc_52155_new_n14410_));
OR2X2 OR2X2_2961 ( .A(u2__abc_52155_new_n14417_), .B(u2__abc_52155_new_n14414_), .Y(u2__abc_52155_new_n14418_));
OR2X2 OR2X2_2962 ( .A(u2__abc_52155_new_n14420_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14421_));
OR2X2 OR2X2_2963 ( .A(u2__abc_52155_new_n14419_), .B(u2__abc_52155_new_n14421_), .Y(u2__abc_52155_new_n14422_));
OR2X2 OR2X2_2964 ( .A(u2__abc_52155_new_n14426_), .B(u2__abc_52155_new_n14412_), .Y(u2__abc_52155_new_n14427_));
OR2X2 OR2X2_2965 ( .A(u2__abc_52155_new_n14431_), .B(u2__abc_52155_new_n5864_), .Y(u2__abc_52155_new_n14432_));
OR2X2 OR2X2_2966 ( .A(u2__abc_52155_new_n14433_), .B(u2__abc_52155_new_n5844_), .Y(u2__abc_52155_new_n14436_));
OR2X2 OR2X2_2967 ( .A(u2__abc_52155_new_n14439_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14440_));
OR2X2 OR2X2_2968 ( .A(u2__abc_52155_new_n14438_), .B(u2__abc_52155_new_n14440_), .Y(u2__abc_52155_new_n14441_));
OR2X2 OR2X2_2969 ( .A(u2__abc_52155_new_n14445_), .B(u2__abc_52155_new_n14429_), .Y(u2__abc_52155_new_n14446_));
OR2X2 OR2X2_297 ( .A(_abc_73687_new_n1170_), .B(\a[36] ), .Y(_abc_73687_new_n1276_));
OR2X2 OR2X2_2970 ( .A(u2__abc_52155_new_n14450_), .B(u2__abc_52155_new_n14449_), .Y(u2__abc_52155_new_n14451_));
OR2X2 OR2X2_2971 ( .A(u2__abc_52155_new_n14452_), .B(u2__abc_52155_new_n5851_), .Y(u2__abc_52155_new_n14453_));
OR2X2 OR2X2_2972 ( .A(u2__abc_52155_new_n14456_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14457_));
OR2X2 OR2X2_2973 ( .A(u2__abc_52155_new_n14455_), .B(u2__abc_52155_new_n14457_), .Y(u2__abc_52155_new_n14458_));
OR2X2 OR2X2_2974 ( .A(u2__abc_52155_new_n14462_), .B(u2__abc_52155_new_n14448_), .Y(u2__abc_52155_new_n14463_));
OR2X2 OR2X2_2975 ( .A(u2__abc_52155_new_n14430_), .B(u2__abc_52155_new_n5864_), .Y(u2__abc_52155_new_n14466_));
OR2X2 OR2X2_2976 ( .A(u2__abc_52155_new_n6812_), .B(u2__abc_52155_new_n14466_), .Y(u2__abc_52155_new_n14467_));
OR2X2 OR2X2_2977 ( .A(u2__abc_52155_new_n14468_), .B(u2__abc_52155_new_n5846_), .Y(u2__abc_52155_new_n14469_));
OR2X2 OR2X2_2978 ( .A(u2__abc_52155_new_n14473_), .B(u2__abc_52155_new_n14472_), .Y(u2__abc_52155_new_n14474_));
OR2X2 OR2X2_2979 ( .A(u2__abc_52155_new_n14474_), .B(u2__abc_52155_new_n5890_), .Y(u2__abc_52155_new_n14477_));
OR2X2 OR2X2_298 ( .A(\a[112] ), .B(\a[36] ), .Y(_abc_73687_new_n1278_));
OR2X2 OR2X2_2980 ( .A(u2__abc_52155_new_n14480_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14481_));
OR2X2 OR2X2_2981 ( .A(u2__abc_52155_new_n14479_), .B(u2__abc_52155_new_n14481_), .Y(u2__abc_52155_new_n14482_));
OR2X2 OR2X2_2982 ( .A(u2__abc_52155_new_n14486_), .B(u2__abc_52155_new_n14465_), .Y(u2__abc_52155_new_n14487_));
OR2X2 OR2X2_2983 ( .A(u2__abc_52155_new_n14494_), .B(u2__abc_52155_new_n14491_), .Y(u2__abc_52155_new_n14495_));
OR2X2 OR2X2_2984 ( .A(u2__abc_52155_new_n14497_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14498_));
OR2X2 OR2X2_2985 ( .A(u2__abc_52155_new_n14496_), .B(u2__abc_52155_new_n14498_), .Y(u2__abc_52155_new_n14499_));
OR2X2 OR2X2_2986 ( .A(u2__abc_52155_new_n14503_), .B(u2__abc_52155_new_n14489_), .Y(u2__abc_52155_new_n14504_));
OR2X2 OR2X2_2987 ( .A(u2__abc_52155_new_n14508_), .B(u2__abc_52155_new_n5895_), .Y(u2__abc_52155_new_n14509_));
OR2X2 OR2X2_2988 ( .A(u2__abc_52155_new_n14510_), .B(u2__abc_52155_new_n5875_), .Y(u2__abc_52155_new_n14513_));
OR2X2 OR2X2_2989 ( .A(u2__abc_52155_new_n14516_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14517_));
OR2X2 OR2X2_299 ( .A(_abc_73687_new_n1170_), .B(\a[37] ), .Y(_abc_73687_new_n1279_));
OR2X2 OR2X2_2990 ( .A(u2__abc_52155_new_n14515_), .B(u2__abc_52155_new_n14517_), .Y(u2__abc_52155_new_n14518_));
OR2X2 OR2X2_2991 ( .A(u2__abc_52155_new_n14522_), .B(u2__abc_52155_new_n14506_), .Y(u2__abc_52155_new_n14523_));
OR2X2 OR2X2_2992 ( .A(u2__abc_52155_new_n14527_), .B(u2__abc_52155_new_n14526_), .Y(u2__abc_52155_new_n14528_));
OR2X2 OR2X2_2993 ( .A(u2__abc_52155_new_n14529_), .B(u2__abc_52155_new_n5882_), .Y(u2__abc_52155_new_n14530_));
OR2X2 OR2X2_2994 ( .A(u2__abc_52155_new_n14533_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14534_));
OR2X2 OR2X2_2995 ( .A(u2__abc_52155_new_n14532_), .B(u2__abc_52155_new_n14534_), .Y(u2__abc_52155_new_n14535_));
OR2X2 OR2X2_2996 ( .A(u2__abc_52155_new_n14539_), .B(u2__abc_52155_new_n14525_), .Y(u2__abc_52155_new_n14540_));
OR2X2 OR2X2_2997 ( .A(u2__abc_52155_new_n14507_), .B(u2__abc_52155_new_n5895_), .Y(u2__abc_52155_new_n14549_));
OR2X2 OR2X2_2998 ( .A(u2__abc_52155_new_n6821_), .B(u2__abc_52155_new_n14549_), .Y(u2__abc_52155_new_n14550_));
OR2X2 OR2X2_2999 ( .A(u2__abc_52155_new_n14551_), .B(u2__abc_52155_new_n5877_), .Y(u2__abc_52155_new_n14552_));
OR2X2 OR2X2_3 ( .A(aNan), .B(sqrto_77_), .Y(_abc_73687_new_n833_));
OR2X2 OR2X2_30 ( .A(_abc_73687_new_n753_), .B(\a[14] ), .Y(_abc_73687_new_n873_));
OR2X2 OR2X2_300 ( .A(\a[112] ), .B(\a[37] ), .Y(_abc_73687_new_n1281_));
OR2X2 OR2X2_3000 ( .A(u2__abc_52155_new_n14559_), .B(u2__abc_52155_new_n14558_), .Y(u2__abc_52155_new_n14560_));
OR2X2 OR2X2_3001 ( .A(u2__abc_52155_new_n14560_), .B(u2__abc_52155_new_n5794_), .Y(u2__abc_52155_new_n14563_));
OR2X2 OR2X2_3002 ( .A(u2__abc_52155_new_n14566_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14567_));
OR2X2 OR2X2_3003 ( .A(u2__abc_52155_new_n14565_), .B(u2__abc_52155_new_n14567_), .Y(u2__abc_52155_new_n14568_));
OR2X2 OR2X2_3004 ( .A(u2__abc_52155_new_n14572_), .B(u2__abc_52155_new_n14542_), .Y(u2__abc_52155_new_n14573_));
OR2X2 OR2X2_3005 ( .A(u2__abc_52155_new_n14580_), .B(u2__abc_52155_new_n14577_), .Y(u2__abc_52155_new_n14581_));
OR2X2 OR2X2_3006 ( .A(u2__abc_52155_new_n14583_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14584_));
OR2X2 OR2X2_3007 ( .A(u2__abc_52155_new_n14582_), .B(u2__abc_52155_new_n14584_), .Y(u2__abc_52155_new_n14585_));
OR2X2 OR2X2_3008 ( .A(u2__abc_52155_new_n14589_), .B(u2__abc_52155_new_n14575_), .Y(u2__abc_52155_new_n14590_));
OR2X2 OR2X2_3009 ( .A(u2__abc_52155_new_n14594_), .B(u2__abc_52155_new_n5799_), .Y(u2__abc_52155_new_n14595_));
OR2X2 OR2X2_301 ( .A(_abc_73687_new_n1170_), .B(\a[38] ), .Y(_abc_73687_new_n1282_));
OR2X2 OR2X2_3010 ( .A(u2__abc_52155_new_n14596_), .B(u2__abc_52155_new_n5779_), .Y(u2__abc_52155_new_n14599_));
OR2X2 OR2X2_3011 ( .A(u2__abc_52155_new_n14602_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14603_));
OR2X2 OR2X2_3012 ( .A(u2__abc_52155_new_n14601_), .B(u2__abc_52155_new_n14603_), .Y(u2__abc_52155_new_n14604_));
OR2X2 OR2X2_3013 ( .A(u2__abc_52155_new_n14608_), .B(u2__abc_52155_new_n14592_), .Y(u2__abc_52155_new_n14609_));
OR2X2 OR2X2_3014 ( .A(u2__abc_52155_new_n14613_), .B(u2__abc_52155_new_n14612_), .Y(u2__abc_52155_new_n14614_));
OR2X2 OR2X2_3015 ( .A(u2__abc_52155_new_n14615_), .B(u2__abc_52155_new_n5786_), .Y(u2__abc_52155_new_n14616_));
OR2X2 OR2X2_3016 ( .A(u2__abc_52155_new_n14619_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14620_));
OR2X2 OR2X2_3017 ( .A(u2__abc_52155_new_n14618_), .B(u2__abc_52155_new_n14620_), .Y(u2__abc_52155_new_n14621_));
OR2X2 OR2X2_3018 ( .A(u2__abc_52155_new_n14625_), .B(u2__abc_52155_new_n14611_), .Y(u2__abc_52155_new_n14626_));
OR2X2 OR2X2_3019 ( .A(u2__abc_52155_new_n14593_), .B(u2__abc_52155_new_n5799_), .Y(u2__abc_52155_new_n14629_));
OR2X2 OR2X2_302 ( .A(\a[112] ), .B(\a[38] ), .Y(_abc_73687_new_n1284_));
OR2X2 OR2X2_3020 ( .A(u2__abc_52155_new_n6889_), .B(u2__abc_52155_new_n14629_), .Y(u2__abc_52155_new_n14630_));
OR2X2 OR2X2_3021 ( .A(u2__abc_52155_new_n14631_), .B(u2__abc_52155_new_n5781_), .Y(u2__abc_52155_new_n14632_));
OR2X2 OR2X2_3022 ( .A(u2__abc_52155_new_n14636_), .B(u2__abc_52155_new_n14635_), .Y(u2__abc_52155_new_n14637_));
OR2X2 OR2X2_3023 ( .A(u2__abc_52155_new_n14637_), .B(u2__abc_52155_new_n5825_), .Y(u2__abc_52155_new_n14640_));
OR2X2 OR2X2_3024 ( .A(u2__abc_52155_new_n14643_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14644_));
OR2X2 OR2X2_3025 ( .A(u2__abc_52155_new_n14642_), .B(u2__abc_52155_new_n14644_), .Y(u2__abc_52155_new_n14645_));
OR2X2 OR2X2_3026 ( .A(u2__abc_52155_new_n14649_), .B(u2__abc_52155_new_n14628_), .Y(u2__abc_52155_new_n14650_));
OR2X2 OR2X2_3027 ( .A(u2__abc_52155_new_n14657_), .B(u2__abc_52155_new_n14654_), .Y(u2__abc_52155_new_n14658_));
OR2X2 OR2X2_3028 ( .A(u2__abc_52155_new_n14660_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14661_));
OR2X2 OR2X2_3029 ( .A(u2__abc_52155_new_n14659_), .B(u2__abc_52155_new_n14661_), .Y(u2__abc_52155_new_n14662_));
OR2X2 OR2X2_303 ( .A(_abc_73687_new_n1170_), .B(\a[39] ), .Y(_abc_73687_new_n1285_));
OR2X2 OR2X2_3030 ( .A(u2__abc_52155_new_n14666_), .B(u2__abc_52155_new_n14652_), .Y(u2__abc_52155_new_n14667_));
OR2X2 OR2X2_3031 ( .A(u2__abc_52155_new_n14671_), .B(u2__abc_52155_new_n5830_), .Y(u2__abc_52155_new_n14672_));
OR2X2 OR2X2_3032 ( .A(u2__abc_52155_new_n14673_), .B(u2__abc_52155_new_n5810_), .Y(u2__abc_52155_new_n14676_));
OR2X2 OR2X2_3033 ( .A(u2__abc_52155_new_n14679_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14680_));
OR2X2 OR2X2_3034 ( .A(u2__abc_52155_new_n14678_), .B(u2__abc_52155_new_n14680_), .Y(u2__abc_52155_new_n14681_));
OR2X2 OR2X2_3035 ( .A(u2__abc_52155_new_n14685_), .B(u2__abc_52155_new_n14669_), .Y(u2__abc_52155_new_n14686_));
OR2X2 OR2X2_3036 ( .A(u2__abc_52155_new_n14690_), .B(u2__abc_52155_new_n14689_), .Y(u2__abc_52155_new_n14691_));
OR2X2 OR2X2_3037 ( .A(u2__abc_52155_new_n14692_), .B(u2__abc_52155_new_n5817_), .Y(u2__abc_52155_new_n14693_));
OR2X2 OR2X2_3038 ( .A(u2__abc_52155_new_n14696_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14697_));
OR2X2 OR2X2_3039 ( .A(u2__abc_52155_new_n14695_), .B(u2__abc_52155_new_n14697_), .Y(u2__abc_52155_new_n14698_));
OR2X2 OR2X2_304 ( .A(\a[112] ), .B(\a[39] ), .Y(_abc_73687_new_n1287_));
OR2X2 OR2X2_3040 ( .A(u2__abc_52155_new_n14702_), .B(u2__abc_52155_new_n14688_), .Y(u2__abc_52155_new_n14703_));
OR2X2 OR2X2_3041 ( .A(u2__abc_52155_new_n14670_), .B(u2__abc_52155_new_n5830_), .Y(u2__abc_52155_new_n14709_));
OR2X2 OR2X2_3042 ( .A(u2__abc_52155_new_n14708_), .B(u2__abc_52155_new_n14709_), .Y(u2__abc_52155_new_n14710_));
OR2X2 OR2X2_3043 ( .A(u2__abc_52155_new_n14711_), .B(u2__abc_52155_new_n5815_), .Y(u2__abc_52155_new_n14712_));
OR2X2 OR2X2_3044 ( .A(u2__abc_52155_new_n14716_), .B(u2__abc_52155_new_n14715_), .Y(u2__abc_52155_new_n14717_));
OR2X2 OR2X2_3045 ( .A(u2__abc_52155_new_n14717_), .B(u2__abc_52155_new_n5716_), .Y(u2__abc_52155_new_n14720_));
OR2X2 OR2X2_3046 ( .A(u2__abc_52155_new_n14723_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14724_));
OR2X2 OR2X2_3047 ( .A(u2__abc_52155_new_n14722_), .B(u2__abc_52155_new_n14724_), .Y(u2__abc_52155_new_n14725_));
OR2X2 OR2X2_3048 ( .A(u2__abc_52155_new_n14729_), .B(u2__abc_52155_new_n14705_), .Y(u2__abc_52155_new_n14730_));
OR2X2 OR2X2_3049 ( .A(u2__abc_52155_new_n14734_), .B(u2__abc_52155_new_n14733_), .Y(u2__abc_52155_new_n14735_));
OR2X2 OR2X2_305 ( .A(_abc_73687_new_n1170_), .B(\a[40] ), .Y(_abc_73687_new_n1288_));
OR2X2 OR2X2_3050 ( .A(u2__abc_52155_new_n14736_), .B(u2__abc_52155_new_n5723_), .Y(u2__abc_52155_new_n14737_));
OR2X2 OR2X2_3051 ( .A(u2__abc_52155_new_n14740_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14741_));
OR2X2 OR2X2_3052 ( .A(u2__abc_52155_new_n14739_), .B(u2__abc_52155_new_n14741_), .Y(u2__abc_52155_new_n14742_));
OR2X2 OR2X2_3053 ( .A(u2__abc_52155_new_n14746_), .B(u2__abc_52155_new_n14732_), .Y(u2__abc_52155_new_n14747_));
OR2X2 OR2X2_3054 ( .A(u2__abc_52155_new_n14750_), .B(u2__abc_52155_new_n5718_), .Y(u2__abc_52155_new_n14751_));
OR2X2 OR2X2_3055 ( .A(u2__abc_52155_new_n14753_), .B(u2__abc_52155_new_n14752_), .Y(u2__abc_52155_new_n14754_));
OR2X2 OR2X2_3056 ( .A(u2__abc_52155_new_n14754_), .B(u2__abc_52155_new_n5731_), .Y(u2__abc_52155_new_n14757_));
OR2X2 OR2X2_3057 ( .A(u2__abc_52155_new_n14760_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14761_));
OR2X2 OR2X2_3058 ( .A(u2__abc_52155_new_n14759_), .B(u2__abc_52155_new_n14761_), .Y(u2__abc_52155_new_n14762_));
OR2X2 OR2X2_3059 ( .A(u2__abc_52155_new_n14766_), .B(u2__abc_52155_new_n14749_), .Y(u2__abc_52155_new_n14767_));
OR2X2 OR2X2_306 ( .A(\a[112] ), .B(\a[40] ), .Y(_abc_73687_new_n1290_));
OR2X2 OR2X2_3060 ( .A(u2__abc_52155_new_n14771_), .B(u2__abc_52155_new_n14770_), .Y(u2__abc_52155_new_n14772_));
OR2X2 OR2X2_3061 ( .A(u2__abc_52155_new_n14773_), .B(u2__abc_52155_new_n5738_), .Y(u2__abc_52155_new_n14774_));
OR2X2 OR2X2_3062 ( .A(u2__abc_52155_new_n14777_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14778_));
OR2X2 OR2X2_3063 ( .A(u2__abc_52155_new_n14776_), .B(u2__abc_52155_new_n14778_), .Y(u2__abc_52155_new_n14779_));
OR2X2 OR2X2_3064 ( .A(u2__abc_52155_new_n14783_), .B(u2__abc_52155_new_n14769_), .Y(u2__abc_52155_new_n14784_));
OR2X2 OR2X2_3065 ( .A(u2__abc_52155_new_n14788_), .B(u2__abc_52155_new_n5733_), .Y(u2__abc_52155_new_n14789_));
OR2X2 OR2X2_3066 ( .A(u2__abc_52155_new_n14787_), .B(u2__abc_52155_new_n14789_), .Y(u2__abc_52155_new_n14790_));
OR2X2 OR2X2_3067 ( .A(u2__abc_52155_new_n14791_), .B(u2__abc_52155_new_n14790_), .Y(u2__abc_52155_new_n14792_));
OR2X2 OR2X2_3068 ( .A(u2__abc_52155_new_n14792_), .B(u2__abc_52155_new_n5762_), .Y(u2__abc_52155_new_n14795_));
OR2X2 OR2X2_3069 ( .A(u2__abc_52155_new_n14798_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14799_));
OR2X2 OR2X2_307 ( .A(_abc_73687_new_n1170_), .B(\a[41] ), .Y(_abc_73687_new_n1291_));
OR2X2 OR2X2_3070 ( .A(u2__abc_52155_new_n14797_), .B(u2__abc_52155_new_n14799_), .Y(u2__abc_52155_new_n14800_));
OR2X2 OR2X2_3071 ( .A(u2__abc_52155_new_n14804_), .B(u2__abc_52155_new_n14786_), .Y(u2__abc_52155_new_n14805_));
OR2X2 OR2X2_3072 ( .A(u2__abc_52155_new_n14812_), .B(u2__abc_52155_new_n14809_), .Y(u2__abc_52155_new_n14813_));
OR2X2 OR2X2_3073 ( .A(u2__abc_52155_new_n14815_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14816_));
OR2X2 OR2X2_3074 ( .A(u2__abc_52155_new_n14814_), .B(u2__abc_52155_new_n14816_), .Y(u2__abc_52155_new_n14817_));
OR2X2 OR2X2_3075 ( .A(u2__abc_52155_new_n14821_), .B(u2__abc_52155_new_n14807_), .Y(u2__abc_52155_new_n14822_));
OR2X2 OR2X2_3076 ( .A(u2__abc_52155_new_n14826_), .B(u2__abc_52155_new_n5767_), .Y(u2__abc_52155_new_n14827_));
OR2X2 OR2X2_3077 ( .A(u2__abc_52155_new_n14828_), .B(u2__abc_52155_new_n5747_), .Y(u2__abc_52155_new_n14831_));
OR2X2 OR2X2_3078 ( .A(u2__abc_52155_new_n14834_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14835_));
OR2X2 OR2X2_3079 ( .A(u2__abc_52155_new_n14833_), .B(u2__abc_52155_new_n14835_), .Y(u2__abc_52155_new_n14836_));
OR2X2 OR2X2_308 ( .A(\a[112] ), .B(\a[41] ), .Y(_abc_73687_new_n1293_));
OR2X2 OR2X2_3080 ( .A(u2__abc_52155_new_n14840_), .B(u2__abc_52155_new_n14824_), .Y(u2__abc_52155_new_n14841_));
OR2X2 OR2X2_3081 ( .A(u2__abc_52155_new_n14845_), .B(u2__abc_52155_new_n14844_), .Y(u2__abc_52155_new_n14846_));
OR2X2 OR2X2_3082 ( .A(u2__abc_52155_new_n14847_), .B(u2__abc_52155_new_n5754_), .Y(u2__abc_52155_new_n14848_));
OR2X2 OR2X2_3083 ( .A(u2__abc_52155_new_n14851_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14852_));
OR2X2 OR2X2_3084 ( .A(u2__abc_52155_new_n14850_), .B(u2__abc_52155_new_n14852_), .Y(u2__abc_52155_new_n14853_));
OR2X2 OR2X2_3085 ( .A(u2__abc_52155_new_n14857_), .B(u2__abc_52155_new_n14843_), .Y(u2__abc_52155_new_n14858_));
OR2X2 OR2X2_3086 ( .A(u2__abc_52155_new_n14825_), .B(u2__abc_52155_new_n5767_), .Y(u2__abc_52155_new_n14866_));
OR2X2 OR2X2_3087 ( .A(u2__abc_52155_new_n14865_), .B(u2__abc_52155_new_n14866_), .Y(u2__abc_52155_new_n14867_));
OR2X2 OR2X2_3088 ( .A(u2__abc_52155_new_n14868_), .B(u2__abc_52155_new_n5749_), .Y(u2__abc_52155_new_n14869_));
OR2X2 OR2X2_3089 ( .A(u2__abc_52155_new_n14875_), .B(u2__abc_52155_new_n14874_), .Y(u2__abc_52155_new_n14876_));
OR2X2 OR2X2_309 ( .A(_abc_73687_new_n1170_), .B(\a[42] ), .Y(_abc_73687_new_n1294_));
OR2X2 OR2X2_3090 ( .A(u2__abc_52155_new_n14876_), .B(u2__abc_52155_new_n5667_), .Y(u2__abc_52155_new_n14879_));
OR2X2 OR2X2_3091 ( .A(u2__abc_52155_new_n14882_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14883_));
OR2X2 OR2X2_3092 ( .A(u2__abc_52155_new_n14881_), .B(u2__abc_52155_new_n14883_), .Y(u2__abc_52155_new_n14884_));
OR2X2 OR2X2_3093 ( .A(u2__abc_52155_new_n14888_), .B(u2__abc_52155_new_n14860_), .Y(u2__abc_52155_new_n14889_));
OR2X2 OR2X2_3094 ( .A(u2__abc_52155_new_n14896_), .B(u2__abc_52155_new_n14893_), .Y(u2__abc_52155_new_n14897_));
OR2X2 OR2X2_3095 ( .A(u2__abc_52155_new_n14899_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14900_));
OR2X2 OR2X2_3096 ( .A(u2__abc_52155_new_n14898_), .B(u2__abc_52155_new_n14900_), .Y(u2__abc_52155_new_n14901_));
OR2X2 OR2X2_3097 ( .A(u2__abc_52155_new_n14905_), .B(u2__abc_52155_new_n14891_), .Y(u2__abc_52155_new_n14906_));
OR2X2 OR2X2_3098 ( .A(u2__abc_52155_new_n14910_), .B(u2__abc_52155_new_n5672_), .Y(u2__abc_52155_new_n14911_));
OR2X2 OR2X2_3099 ( .A(u2__abc_52155_new_n14912_), .B(u2__abc_52155_new_n5652_), .Y(u2__abc_52155_new_n14915_));
OR2X2 OR2X2_31 ( .A(aNan), .B(sqrto_91_), .Y(_abc_73687_new_n875_));
OR2X2 OR2X2_310 ( .A(\a[112] ), .B(\a[42] ), .Y(_abc_73687_new_n1296_));
OR2X2 OR2X2_3100 ( .A(u2__abc_52155_new_n14918_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14919_));
OR2X2 OR2X2_3101 ( .A(u2__abc_52155_new_n14917_), .B(u2__abc_52155_new_n14919_), .Y(u2__abc_52155_new_n14920_));
OR2X2 OR2X2_3102 ( .A(u2__abc_52155_new_n14924_), .B(u2__abc_52155_new_n14908_), .Y(u2__abc_52155_new_n14925_));
OR2X2 OR2X2_3103 ( .A(u2__abc_52155_new_n14929_), .B(u2__abc_52155_new_n14928_), .Y(u2__abc_52155_new_n14930_));
OR2X2 OR2X2_3104 ( .A(u2__abc_52155_new_n14931_), .B(u2__abc_52155_new_n5659_), .Y(u2__abc_52155_new_n14932_));
OR2X2 OR2X2_3105 ( .A(u2__abc_52155_new_n14935_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14936_));
OR2X2 OR2X2_3106 ( .A(u2__abc_52155_new_n14934_), .B(u2__abc_52155_new_n14936_), .Y(u2__abc_52155_new_n14937_));
OR2X2 OR2X2_3107 ( .A(u2__abc_52155_new_n14941_), .B(u2__abc_52155_new_n14927_), .Y(u2__abc_52155_new_n14942_));
OR2X2 OR2X2_3108 ( .A(u2__abc_52155_new_n5647_), .B(u2__abc_52155_new_n5654_), .Y(u2__abc_52155_new_n14945_));
OR2X2 OR2X2_3109 ( .A(u2__abc_52155_new_n14909_), .B(u2__abc_52155_new_n5672_), .Y(u2__abc_52155_new_n14948_));
OR2X2 OR2X2_311 ( .A(_abc_73687_new_n1170_), .B(\a[43] ), .Y(_abc_73687_new_n1297_));
OR2X2 OR2X2_3110 ( .A(u2__abc_52155_new_n6858_), .B(u2__abc_52155_new_n14948_), .Y(u2__abc_52155_new_n14949_));
OR2X2 OR2X2_3111 ( .A(u2__abc_52155_new_n14952_), .B(u2__abc_52155_new_n14951_), .Y(u2__abc_52155_new_n14953_));
OR2X2 OR2X2_3112 ( .A(u2__abc_52155_new_n14953_), .B(u2__abc_52155_new_n5705_), .Y(u2__abc_52155_new_n14956_));
OR2X2 OR2X2_3113 ( .A(u2__abc_52155_new_n14959_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14960_));
OR2X2 OR2X2_3114 ( .A(u2__abc_52155_new_n14958_), .B(u2__abc_52155_new_n14960_), .Y(u2__abc_52155_new_n14961_));
OR2X2 OR2X2_3115 ( .A(u2__abc_52155_new_n14965_), .B(u2__abc_52155_new_n14944_), .Y(u2__abc_52155_new_n14966_));
OR2X2 OR2X2_3116 ( .A(u2__abc_52155_new_n14970_), .B(u2__abc_52155_new_n5698_), .Y(u2__abc_52155_new_n14973_));
OR2X2 OR2X2_3117 ( .A(u2__abc_52155_new_n14976_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14977_));
OR2X2 OR2X2_3118 ( .A(u2__abc_52155_new_n14975_), .B(u2__abc_52155_new_n14977_), .Y(u2__abc_52155_new_n14978_));
OR2X2 OR2X2_3119 ( .A(u2__abc_52155_new_n14982_), .B(u2__abc_52155_new_n14968_), .Y(u2__abc_52155_new_n14983_));
OR2X2 OR2X2_312 ( .A(\a[112] ), .B(\a[43] ), .Y(_abc_73687_new_n1299_));
OR2X2 OR2X2_3120 ( .A(u2__abc_52155_new_n14987_), .B(u2__abc_52155_new_n5683_), .Y(u2__abc_52155_new_n14990_));
OR2X2 OR2X2_3121 ( .A(u2__abc_52155_new_n14993_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n14994_));
OR2X2 OR2X2_3122 ( .A(u2__abc_52155_new_n14992_), .B(u2__abc_52155_new_n14994_), .Y(u2__abc_52155_new_n14995_));
OR2X2 OR2X2_3123 ( .A(u2__abc_52155_new_n14999_), .B(u2__abc_52155_new_n14985_), .Y(u2__abc_52155_new_n15000_));
OR2X2 OR2X2_3124 ( .A(u2__abc_52155_new_n15004_), .B(u2__abc_52155_new_n15003_), .Y(u2__abc_52155_new_n15005_));
OR2X2 OR2X2_3125 ( .A(u2__abc_52155_new_n15006_), .B(u2__abc_52155_new_n5690_), .Y(u2__abc_52155_new_n15007_));
OR2X2 OR2X2_3126 ( .A(u2__abc_52155_new_n15010_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15011_));
OR2X2 OR2X2_3127 ( .A(u2__abc_52155_new_n15009_), .B(u2__abc_52155_new_n15011_), .Y(u2__abc_52155_new_n15012_));
OR2X2 OR2X2_3128 ( .A(u2__abc_52155_new_n15016_), .B(u2__abc_52155_new_n15002_), .Y(u2__abc_52155_new_n15017_));
OR2X2 OR2X2_3129 ( .A(u2__abc_52155_new_n15021_), .B(u2__abc_52155_new_n5693_), .Y(u2__abc_52155_new_n15022_));
OR2X2 OR2X2_313 ( .A(_abc_73687_new_n1170_), .B(\a[44] ), .Y(_abc_73687_new_n1300_));
OR2X2 OR2X2_3130 ( .A(u2__abc_52155_new_n15024_), .B(u2__abc_52155_new_n5685_), .Y(u2__abc_52155_new_n15025_));
OR2X2 OR2X2_3131 ( .A(u2__abc_52155_new_n15023_), .B(u2__abc_52155_new_n15025_), .Y(u2__abc_52155_new_n15026_));
OR2X2 OR2X2_3132 ( .A(u2__abc_52155_new_n15020_), .B(u2__abc_52155_new_n15026_), .Y(u2__abc_52155_new_n15027_));
OR2X2 OR2X2_3133 ( .A(u2__abc_52155_new_n15028_), .B(u2__abc_52155_new_n15027_), .Y(u2__abc_52155_new_n15029_));
OR2X2 OR2X2_3134 ( .A(u2__abc_52155_new_n15029_), .B(u2__abc_52155_new_n5620_), .Y(u2__abc_52155_new_n15032_));
OR2X2 OR2X2_3135 ( .A(u2__abc_52155_new_n15035_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15036_));
OR2X2 OR2X2_3136 ( .A(u2__abc_52155_new_n15034_), .B(u2__abc_52155_new_n15036_), .Y(u2__abc_52155_new_n15037_));
OR2X2 OR2X2_3137 ( .A(u2__abc_52155_new_n15041_), .B(u2__abc_52155_new_n15019_), .Y(u2__abc_52155_new_n15042_));
OR2X2 OR2X2_3138 ( .A(u2__abc_52155_new_n15046_), .B(u2__abc_52155_new_n15045_), .Y(u2__abc_52155_new_n15047_));
OR2X2 OR2X2_3139 ( .A(u2__abc_52155_new_n15048_), .B(u2__abc_52155_new_n5627_), .Y(u2__abc_52155_new_n15049_));
OR2X2 OR2X2_314 ( .A(\a[112] ), .B(\a[44] ), .Y(_abc_73687_new_n1302_));
OR2X2 OR2X2_3140 ( .A(u2__abc_52155_new_n15052_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15053_));
OR2X2 OR2X2_3141 ( .A(u2__abc_52155_new_n15051_), .B(u2__abc_52155_new_n15053_), .Y(u2__abc_52155_new_n15054_));
OR2X2 OR2X2_3142 ( .A(u2__abc_52155_new_n15058_), .B(u2__abc_52155_new_n15044_), .Y(u2__abc_52155_new_n15059_));
OR2X2 OR2X2_3143 ( .A(u2__abc_52155_new_n15062_), .B(u2__abc_52155_new_n5622_), .Y(u2__abc_52155_new_n15063_));
OR2X2 OR2X2_3144 ( .A(u2__abc_52155_new_n15065_), .B(u2__abc_52155_new_n15064_), .Y(u2__abc_52155_new_n15066_));
OR2X2 OR2X2_3145 ( .A(u2__abc_52155_new_n15066_), .B(u2__abc_52155_new_n5635_), .Y(u2__abc_52155_new_n15069_));
OR2X2 OR2X2_3146 ( .A(u2__abc_52155_new_n15072_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15073_));
OR2X2 OR2X2_3147 ( .A(u2__abc_52155_new_n15071_), .B(u2__abc_52155_new_n15073_), .Y(u2__abc_52155_new_n15074_));
OR2X2 OR2X2_3148 ( .A(u2__abc_52155_new_n15078_), .B(u2__abc_52155_new_n15061_), .Y(u2__abc_52155_new_n15079_));
OR2X2 OR2X2_3149 ( .A(u2__abc_52155_new_n15083_), .B(u2__abc_52155_new_n15082_), .Y(u2__abc_52155_new_n15084_));
OR2X2 OR2X2_315 ( .A(_abc_73687_new_n1170_), .B(\a[45] ), .Y(_abc_73687_new_n1303_));
OR2X2 OR2X2_3150 ( .A(u2__abc_52155_new_n15085_), .B(u2__abc_52155_new_n5642_), .Y(u2__abc_52155_new_n15086_));
OR2X2 OR2X2_3151 ( .A(u2__abc_52155_new_n15089_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15090_));
OR2X2 OR2X2_3152 ( .A(u2__abc_52155_new_n15088_), .B(u2__abc_52155_new_n15090_), .Y(u2__abc_52155_new_n15091_));
OR2X2 OR2X2_3153 ( .A(u2__abc_52155_new_n15095_), .B(u2__abc_52155_new_n15081_), .Y(u2__abc_52155_new_n15096_));
OR2X2 OR2X2_3154 ( .A(u2__abc_52155_new_n15099_), .B(u2__abc_52155_new_n5637_), .Y(u2__abc_52155_new_n15100_));
OR2X2 OR2X2_3155 ( .A(u2__abc_52155_new_n15101_), .B(u2__abc_52155_new_n15100_), .Y(u2__abc_52155_new_n15102_));
OR2X2 OR2X2_3156 ( .A(u2__abc_52155_new_n15102_), .B(u2__abc_52155_new_n5604_), .Y(u2__abc_52155_new_n15105_));
OR2X2 OR2X2_3157 ( .A(u2__abc_52155_new_n15108_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15109_));
OR2X2 OR2X2_3158 ( .A(u2__abc_52155_new_n15107_), .B(u2__abc_52155_new_n15109_), .Y(u2__abc_52155_new_n15110_));
OR2X2 OR2X2_3159 ( .A(u2__abc_52155_new_n15114_), .B(u2__abc_52155_new_n15098_), .Y(u2__abc_52155_new_n15115_));
OR2X2 OR2X2_316 ( .A(\a[112] ), .B(\a[45] ), .Y(_abc_73687_new_n1305_));
OR2X2 OR2X2_3160 ( .A(u2__abc_52155_new_n15122_), .B(u2__abc_52155_new_n15119_), .Y(u2__abc_52155_new_n15123_));
OR2X2 OR2X2_3161 ( .A(u2__abc_52155_new_n15125_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15126_));
OR2X2 OR2X2_3162 ( .A(u2__abc_52155_new_n15124_), .B(u2__abc_52155_new_n15126_), .Y(u2__abc_52155_new_n15127_));
OR2X2 OR2X2_3163 ( .A(u2__abc_52155_new_n15131_), .B(u2__abc_52155_new_n15117_), .Y(u2__abc_52155_new_n15132_));
OR2X2 OR2X2_3164 ( .A(u2__abc_52155_new_n15136_), .B(u2__abc_52155_new_n5609_), .Y(u2__abc_52155_new_n15137_));
OR2X2 OR2X2_3165 ( .A(u2__abc_52155_new_n15138_), .B(u2__abc_52155_new_n5589_), .Y(u2__abc_52155_new_n15141_));
OR2X2 OR2X2_3166 ( .A(u2__abc_52155_new_n15144_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15145_));
OR2X2 OR2X2_3167 ( .A(u2__abc_52155_new_n15143_), .B(u2__abc_52155_new_n15145_), .Y(u2__abc_52155_new_n15146_));
OR2X2 OR2X2_3168 ( .A(u2__abc_52155_new_n15150_), .B(u2__abc_52155_new_n15134_), .Y(u2__abc_52155_new_n15151_));
OR2X2 OR2X2_3169 ( .A(u2__abc_52155_new_n15155_), .B(u2__abc_52155_new_n15154_), .Y(u2__abc_52155_new_n15156_));
OR2X2 OR2X2_317 ( .A(_abc_73687_new_n1170_), .B(\a[46] ), .Y(_abc_73687_new_n1306_));
OR2X2 OR2X2_3170 ( .A(u2__abc_52155_new_n15157_), .B(u2__abc_52155_new_n5596_), .Y(u2__abc_52155_new_n15158_));
OR2X2 OR2X2_3171 ( .A(u2__abc_52155_new_n15161_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15162_));
OR2X2 OR2X2_3172 ( .A(u2__abc_52155_new_n15160_), .B(u2__abc_52155_new_n15162_), .Y(u2__abc_52155_new_n15163_));
OR2X2 OR2X2_3173 ( .A(u2__abc_52155_new_n15167_), .B(u2__abc_52155_new_n15153_), .Y(u2__abc_52155_new_n15168_));
OR2X2 OR2X2_3174 ( .A(u2__abc_52155_new_n15181_), .B(u2__abc_52155_new_n15100_), .Y(u2__abc_52155_new_n15182_));
OR2X2 OR2X2_3175 ( .A(u2__abc_52155_new_n15135_), .B(u2__abc_52155_new_n5609_), .Y(u2__abc_52155_new_n15185_));
OR2X2 OR2X2_3176 ( .A(u2__abc_52155_new_n6913_), .B(u2__abc_52155_new_n15185_), .Y(u2__abc_52155_new_n15186_));
OR2X2 OR2X2_3177 ( .A(u2__abc_52155_new_n15187_), .B(u2__abc_52155_new_n5594_), .Y(u2__abc_52155_new_n15188_));
OR2X2 OR2X2_3178 ( .A(u2__abc_52155_new_n15197_), .B(u2__abc_52155_new_n7241_), .Y(u2__abc_52155_new_n15200_));
OR2X2 OR2X2_3179 ( .A(u2__abc_52155_new_n15203_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15204_));
OR2X2 OR2X2_318 ( .A(\a[112] ), .B(\a[46] ), .Y(_abc_73687_new_n1308_));
OR2X2 OR2X2_3180 ( .A(u2__abc_52155_new_n15202_), .B(u2__abc_52155_new_n15204_), .Y(u2__abc_52155_new_n15205_));
OR2X2 OR2X2_3181 ( .A(u2__abc_52155_new_n15209_), .B(u2__abc_52155_new_n15170_), .Y(u2__abc_52155_new_n15210_));
OR2X2 OR2X2_3182 ( .A(u2__abc_52155_new_n15214_), .B(u2__abc_52155_new_n15213_), .Y(u2__abc_52155_new_n15215_));
OR2X2 OR2X2_3183 ( .A(u2__abc_52155_new_n15216_), .B(u2__abc_52155_new_n7234_), .Y(u2__abc_52155_new_n15217_));
OR2X2 OR2X2_3184 ( .A(u2__abc_52155_new_n15220_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15221_));
OR2X2 OR2X2_3185 ( .A(u2__abc_52155_new_n15219_), .B(u2__abc_52155_new_n15221_), .Y(u2__abc_52155_new_n15222_));
OR2X2 OR2X2_3186 ( .A(u2__abc_52155_new_n15226_), .B(u2__abc_52155_new_n15212_), .Y(u2__abc_52155_new_n15227_));
OR2X2 OR2X2_3187 ( .A(u2__abc_52155_new_n15231_), .B(u2__abc_52155_new_n7229_), .Y(u2__abc_52155_new_n15232_));
OR2X2 OR2X2_3188 ( .A(u2__abc_52155_new_n15233_), .B(u2__abc_52155_new_n7219_), .Y(u2__abc_52155_new_n15236_));
OR2X2 OR2X2_3189 ( .A(u2__abc_52155_new_n15239_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15240_));
OR2X2 OR2X2_319 ( .A(_abc_73687_new_n1170_), .B(\a[47] ), .Y(_abc_73687_new_n1309_));
OR2X2 OR2X2_3190 ( .A(u2__abc_52155_new_n15238_), .B(u2__abc_52155_new_n15240_), .Y(u2__abc_52155_new_n15241_));
OR2X2 OR2X2_3191 ( .A(u2__abc_52155_new_n15245_), .B(u2__abc_52155_new_n15229_), .Y(u2__abc_52155_new_n15246_));
OR2X2 OR2X2_3192 ( .A(u2__abc_52155_new_n15250_), .B(u2__abc_52155_new_n15249_), .Y(u2__abc_52155_new_n15251_));
OR2X2 OR2X2_3193 ( .A(u2__abc_52155_new_n15252_), .B(u2__abc_52155_new_n7226_), .Y(u2__abc_52155_new_n15253_));
OR2X2 OR2X2_3194 ( .A(u2__abc_52155_new_n15256_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15257_));
OR2X2 OR2X2_3195 ( .A(u2__abc_52155_new_n15255_), .B(u2__abc_52155_new_n15257_), .Y(u2__abc_52155_new_n15258_));
OR2X2 OR2X2_3196 ( .A(u2__abc_52155_new_n15262_), .B(u2__abc_52155_new_n15248_), .Y(u2__abc_52155_new_n15263_));
OR2X2 OR2X2_3197 ( .A(u2__abc_52155_new_n15230_), .B(u2__abc_52155_new_n7229_), .Y(u2__abc_52155_new_n15266_));
OR2X2 OR2X2_3198 ( .A(u2__abc_52155_new_n15269_), .B(u2__abc_52155_new_n7224_), .Y(u2__abc_52155_new_n15270_));
OR2X2 OR2X2_3199 ( .A(u2__abc_52155_new_n15268_), .B(u2__abc_52155_new_n15270_), .Y(u2__abc_52155_new_n15271_));
OR2X2 OR2X2_32 ( .A(_abc_73687_new_n753_), .B(\a[15] ), .Y(_abc_73687_new_n876_));
OR2X2 OR2X2_320 ( .A(\a[112] ), .B(\a[47] ), .Y(_abc_73687_new_n1311_));
OR2X2 OR2X2_3200 ( .A(u2__abc_52155_new_n15272_), .B(u2__abc_52155_new_n15271_), .Y(u2__abc_52155_new_n15273_));
OR2X2 OR2X2_3201 ( .A(u2__abc_52155_new_n15273_), .B(u2__abc_52155_new_n7210_), .Y(u2__abc_52155_new_n15276_));
OR2X2 OR2X2_3202 ( .A(u2__abc_52155_new_n15279_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15280_));
OR2X2 OR2X2_3203 ( .A(u2__abc_52155_new_n15278_), .B(u2__abc_52155_new_n15280_), .Y(u2__abc_52155_new_n15281_));
OR2X2 OR2X2_3204 ( .A(u2__abc_52155_new_n15285_), .B(u2__abc_52155_new_n15265_), .Y(u2__abc_52155_new_n15286_));
OR2X2 OR2X2_3205 ( .A(u2__abc_52155_new_n15293_), .B(u2__abc_52155_new_n15290_), .Y(u2__abc_52155_new_n15294_));
OR2X2 OR2X2_3206 ( .A(u2__abc_52155_new_n15296_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15297_));
OR2X2 OR2X2_3207 ( .A(u2__abc_52155_new_n15295_), .B(u2__abc_52155_new_n15297_), .Y(u2__abc_52155_new_n15298_));
OR2X2 OR2X2_3208 ( .A(u2__abc_52155_new_n15302_), .B(u2__abc_52155_new_n15288_), .Y(u2__abc_52155_new_n15303_));
OR2X2 OR2X2_3209 ( .A(u2__abc_52155_new_n15307_), .B(u2__abc_52155_new_n7198_), .Y(u2__abc_52155_new_n15308_));
OR2X2 OR2X2_321 ( .A(_abc_73687_new_n1170_), .B(\a[48] ), .Y(_abc_73687_new_n1312_));
OR2X2 OR2X2_3210 ( .A(u2__abc_52155_new_n15309_), .B(u2__abc_52155_new_n7188_), .Y(u2__abc_52155_new_n15312_));
OR2X2 OR2X2_3211 ( .A(u2__abc_52155_new_n15315_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15316_));
OR2X2 OR2X2_3212 ( .A(u2__abc_52155_new_n15314_), .B(u2__abc_52155_new_n15316_), .Y(u2__abc_52155_new_n15317_));
OR2X2 OR2X2_3213 ( .A(u2__abc_52155_new_n15321_), .B(u2__abc_52155_new_n15305_), .Y(u2__abc_52155_new_n15322_));
OR2X2 OR2X2_3214 ( .A(u2__abc_52155_new_n15326_), .B(u2__abc_52155_new_n15325_), .Y(u2__abc_52155_new_n15327_));
OR2X2 OR2X2_3215 ( .A(u2__abc_52155_new_n15328_), .B(u2__abc_52155_new_n7195_), .Y(u2__abc_52155_new_n15329_));
OR2X2 OR2X2_3216 ( .A(u2__abc_52155_new_n15332_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15333_));
OR2X2 OR2X2_3217 ( .A(u2__abc_52155_new_n15331_), .B(u2__abc_52155_new_n15333_), .Y(u2__abc_52155_new_n15334_));
OR2X2 OR2X2_3218 ( .A(u2__abc_52155_new_n15338_), .B(u2__abc_52155_new_n15324_), .Y(u2__abc_52155_new_n15339_));
OR2X2 OR2X2_3219 ( .A(u2__abc_52155_new_n15306_), .B(u2__abc_52155_new_n7198_), .Y(u2__abc_52155_new_n15343_));
OR2X2 OR2X2_322 ( .A(\a[112] ), .B(\a[48] ), .Y(_abc_73687_new_n1314_));
OR2X2 OR2X2_3220 ( .A(u2__abc_52155_new_n15346_), .B(u2__abc_52155_new_n7190_), .Y(u2__abc_52155_new_n15347_));
OR2X2 OR2X2_3221 ( .A(u2__abc_52155_new_n15345_), .B(u2__abc_52155_new_n15347_), .Y(u2__abc_52155_new_n15348_));
OR2X2 OR2X2_3222 ( .A(u2__abc_52155_new_n15342_), .B(u2__abc_52155_new_n15348_), .Y(u2__abc_52155_new_n15349_));
OR2X2 OR2X2_3223 ( .A(u2__abc_52155_new_n15350_), .B(u2__abc_52155_new_n15349_), .Y(u2__abc_52155_new_n15351_));
OR2X2 OR2X2_3224 ( .A(u2__abc_52155_new_n15351_), .B(u2__abc_52155_new_n7393_), .Y(u2__abc_52155_new_n15354_));
OR2X2 OR2X2_3225 ( .A(u2__abc_52155_new_n15357_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15358_));
OR2X2 OR2X2_3226 ( .A(u2__abc_52155_new_n15356_), .B(u2__abc_52155_new_n15358_), .Y(u2__abc_52155_new_n15359_));
OR2X2 OR2X2_3227 ( .A(u2__abc_52155_new_n15363_), .B(u2__abc_52155_new_n15341_), .Y(u2__abc_52155_new_n15364_));
OR2X2 OR2X2_3228 ( .A(u2__abc_52155_new_n15370_), .B(u2__abc_52155_new_n15371_), .Y(u2__abc_52155_new_n15372_));
OR2X2 OR2X2_3229 ( .A(u2__abc_52155_new_n15374_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15375_));
OR2X2 OR2X2_323 ( .A(_abc_73687_new_n1170_), .B(\a[49] ), .Y(_abc_73687_new_n1315_));
OR2X2 OR2X2_3230 ( .A(u2__abc_52155_new_n15373_), .B(u2__abc_52155_new_n15375_), .Y(u2__abc_52155_new_n15376_));
OR2X2 OR2X2_3231 ( .A(u2__abc_52155_new_n15380_), .B(u2__abc_52155_new_n15366_), .Y(u2__abc_52155_new_n15381_));
OR2X2 OR2X2_3232 ( .A(u2__abc_52155_new_n15384_), .B(u2__abc_52155_new_n7398_), .Y(u2__abc_52155_new_n15385_));
OR2X2 OR2X2_3233 ( .A(u2__abc_52155_new_n15385_), .B(u2__abc_52155_new_n7378_), .Y(u2__abc_52155_new_n15388_));
OR2X2 OR2X2_3234 ( .A(u2__abc_52155_new_n15391_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15392_));
OR2X2 OR2X2_3235 ( .A(u2__abc_52155_new_n15390_), .B(u2__abc_52155_new_n15392_), .Y(u2__abc_52155_new_n15393_));
OR2X2 OR2X2_3236 ( .A(u2__abc_52155_new_n15397_), .B(u2__abc_52155_new_n15383_), .Y(u2__abc_52155_new_n15398_));
OR2X2 OR2X2_3237 ( .A(u2__abc_52155_new_n15402_), .B(u2__abc_52155_new_n15401_), .Y(u2__abc_52155_new_n15403_));
OR2X2 OR2X2_3238 ( .A(u2__abc_52155_new_n15404_), .B(u2__abc_52155_new_n7385_), .Y(u2__abc_52155_new_n15405_));
OR2X2 OR2X2_3239 ( .A(u2__abc_52155_new_n15408_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15409_));
OR2X2 OR2X2_324 ( .A(\a[112] ), .B(\a[49] ), .Y(_abc_73687_new_n1317_));
OR2X2 OR2X2_3240 ( .A(u2__abc_52155_new_n15407_), .B(u2__abc_52155_new_n15409_), .Y(u2__abc_52155_new_n15410_));
OR2X2 OR2X2_3241 ( .A(u2__abc_52155_new_n15414_), .B(u2__abc_52155_new_n15400_), .Y(u2__abc_52155_new_n15415_));
OR2X2 OR2X2_3242 ( .A(u2__abc_52155_new_n15418_), .B(u2__abc_52155_new_n7395_), .Y(u2__abc_52155_new_n15419_));
OR2X2 OR2X2_3243 ( .A(u2__abc_52155_new_n15422_), .B(u2__abc_52155_new_n7383_), .Y(u2__abc_52155_new_n15423_));
OR2X2 OR2X2_3244 ( .A(u2__abc_52155_new_n15421_), .B(u2__abc_52155_new_n15423_), .Y(u2__abc_52155_new_n15424_));
OR2X2 OR2X2_3245 ( .A(u2__abc_52155_new_n15425_), .B(u2__abc_52155_new_n15424_), .Y(u2__abc_52155_new_n15426_));
OR2X2 OR2X2_3246 ( .A(u2__abc_52155_new_n15426_), .B(u2__abc_52155_new_n7431_), .Y(u2__abc_52155_new_n15429_));
OR2X2 OR2X2_3247 ( .A(u2__abc_52155_new_n15432_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15433_));
OR2X2 OR2X2_3248 ( .A(u2__abc_52155_new_n15431_), .B(u2__abc_52155_new_n15433_), .Y(u2__abc_52155_new_n15434_));
OR2X2 OR2X2_3249 ( .A(u2__abc_52155_new_n15438_), .B(u2__abc_52155_new_n15417_), .Y(u2__abc_52155_new_n15439_));
OR2X2 OR2X2_325 ( .A(_abc_73687_new_n1170_), .B(\a[50] ), .Y(_abc_73687_new_n1318_));
OR2X2 OR2X2_3250 ( .A(u2__abc_52155_new_n15446_), .B(u2__abc_52155_new_n15443_), .Y(u2__abc_52155_new_n15447_));
OR2X2 OR2X2_3251 ( .A(u2__abc_52155_new_n15449_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15450_));
OR2X2 OR2X2_3252 ( .A(u2__abc_52155_new_n15448_), .B(u2__abc_52155_new_n15450_), .Y(u2__abc_52155_new_n15451_));
OR2X2 OR2X2_3253 ( .A(u2__abc_52155_new_n15455_), .B(u2__abc_52155_new_n15441_), .Y(u2__abc_52155_new_n15456_));
OR2X2 OR2X2_3254 ( .A(u2__abc_52155_new_n15460_), .B(u2__abc_52155_new_n7419_), .Y(u2__abc_52155_new_n15461_));
OR2X2 OR2X2_3255 ( .A(u2__abc_52155_new_n15462_), .B(u2__abc_52155_new_n7409_), .Y(u2__abc_52155_new_n15465_));
OR2X2 OR2X2_3256 ( .A(u2__abc_52155_new_n15468_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15469_));
OR2X2 OR2X2_3257 ( .A(u2__abc_52155_new_n15467_), .B(u2__abc_52155_new_n15469_), .Y(u2__abc_52155_new_n15470_));
OR2X2 OR2X2_3258 ( .A(u2__abc_52155_new_n15474_), .B(u2__abc_52155_new_n15458_), .Y(u2__abc_52155_new_n15475_));
OR2X2 OR2X2_3259 ( .A(u2__abc_52155_new_n15479_), .B(u2__abc_52155_new_n15478_), .Y(u2__abc_52155_new_n15480_));
OR2X2 OR2X2_326 ( .A(\a[112] ), .B(\a[50] ), .Y(_abc_73687_new_n1320_));
OR2X2 OR2X2_3260 ( .A(u2__abc_52155_new_n15481_), .B(u2__abc_52155_new_n7416_), .Y(u2__abc_52155_new_n15482_));
OR2X2 OR2X2_3261 ( .A(u2__abc_52155_new_n15485_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15486_));
OR2X2 OR2X2_3262 ( .A(u2__abc_52155_new_n15484_), .B(u2__abc_52155_new_n15486_), .Y(u2__abc_52155_new_n15487_));
OR2X2 OR2X2_3263 ( .A(u2__abc_52155_new_n15491_), .B(u2__abc_52155_new_n15477_), .Y(u2__abc_52155_new_n15492_));
OR2X2 OR2X2_3264 ( .A(u2__abc_52155_new_n15459_), .B(u2__abc_52155_new_n7419_), .Y(u2__abc_52155_new_n15496_));
OR2X2 OR2X2_3265 ( .A(u2__abc_52155_new_n15499_), .B(u2__abc_52155_new_n7411_), .Y(u2__abc_52155_new_n15500_));
OR2X2 OR2X2_3266 ( .A(u2__abc_52155_new_n15498_), .B(u2__abc_52155_new_n15500_), .Y(u2__abc_52155_new_n15501_));
OR2X2 OR2X2_3267 ( .A(u2__abc_52155_new_n15495_), .B(u2__abc_52155_new_n15501_), .Y(u2__abc_52155_new_n15502_));
OR2X2 OR2X2_3268 ( .A(u2__abc_52155_new_n15503_), .B(u2__abc_52155_new_n15502_), .Y(u2__abc_52155_new_n15504_));
OR2X2 OR2X2_3269 ( .A(u2__abc_52155_new_n15504_), .B(u2__abc_52155_new_n7314_), .Y(u2__abc_52155_new_n15507_));
OR2X2 OR2X2_327 ( .A(_abc_73687_new_n1170_), .B(\a[51] ), .Y(_abc_73687_new_n1321_));
OR2X2 OR2X2_3270 ( .A(u2__abc_52155_new_n15510_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15511_));
OR2X2 OR2X2_3271 ( .A(u2__abc_52155_new_n15509_), .B(u2__abc_52155_new_n15511_), .Y(u2__abc_52155_new_n15512_));
OR2X2 OR2X2_3272 ( .A(u2__abc_52155_new_n15516_), .B(u2__abc_52155_new_n15494_), .Y(u2__abc_52155_new_n15517_));
OR2X2 OR2X2_3273 ( .A(u2__abc_52155_new_n15521_), .B(u2__abc_52155_new_n15520_), .Y(u2__abc_52155_new_n15522_));
OR2X2 OR2X2_3274 ( .A(u2__abc_52155_new_n15523_), .B(u2__abc_52155_new_n7321_), .Y(u2__abc_52155_new_n15524_));
OR2X2 OR2X2_3275 ( .A(u2__abc_52155_new_n15527_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15528_));
OR2X2 OR2X2_3276 ( .A(u2__abc_52155_new_n15526_), .B(u2__abc_52155_new_n15528_), .Y(u2__abc_52155_new_n15529_));
OR2X2 OR2X2_3277 ( .A(u2__abc_52155_new_n15533_), .B(u2__abc_52155_new_n15519_), .Y(u2__abc_52155_new_n15534_));
OR2X2 OR2X2_3278 ( .A(u2__abc_52155_new_n7310_), .B(u2__abc_52155_new_n7316_), .Y(u2__abc_52155_new_n15537_));
OR2X2 OR2X2_3279 ( .A(u2__abc_52155_new_n15540_), .B(u2__abc_52155_new_n15539_), .Y(u2__abc_52155_new_n15541_));
OR2X2 OR2X2_328 ( .A(\a[112] ), .B(\a[51] ), .Y(_abc_73687_new_n1323_));
OR2X2 OR2X2_3280 ( .A(u2__abc_52155_new_n15541_), .B(u2__abc_52155_new_n7329_), .Y(u2__abc_52155_new_n15544_));
OR2X2 OR2X2_3281 ( .A(u2__abc_52155_new_n15547_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15548_));
OR2X2 OR2X2_3282 ( .A(u2__abc_52155_new_n15546_), .B(u2__abc_52155_new_n15548_), .Y(u2__abc_52155_new_n15549_));
OR2X2 OR2X2_3283 ( .A(u2__abc_52155_new_n15553_), .B(u2__abc_52155_new_n15536_), .Y(u2__abc_52155_new_n15554_));
OR2X2 OR2X2_3284 ( .A(u2__abc_52155_new_n15558_), .B(u2__abc_52155_new_n15557_), .Y(u2__abc_52155_new_n15559_));
OR2X2 OR2X2_3285 ( .A(u2__abc_52155_new_n15560_), .B(u2__abc_52155_new_n7336_), .Y(u2__abc_52155_new_n15561_));
OR2X2 OR2X2_3286 ( .A(u2__abc_52155_new_n15564_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15565_));
OR2X2 OR2X2_3287 ( .A(u2__abc_52155_new_n15563_), .B(u2__abc_52155_new_n15565_), .Y(u2__abc_52155_new_n15566_));
OR2X2 OR2X2_3288 ( .A(u2__abc_52155_new_n15570_), .B(u2__abc_52155_new_n15556_), .Y(u2__abc_52155_new_n15571_));
OR2X2 OR2X2_3289 ( .A(u2__abc_52155_new_n15575_), .B(u2__abc_52155_new_n7334_), .Y(u2__abc_52155_new_n15576_));
OR2X2 OR2X2_329 ( .A(_abc_73687_new_n1170_), .B(\a[52] ), .Y(_abc_73687_new_n1324_));
OR2X2 OR2X2_3290 ( .A(u2__abc_52155_new_n15574_), .B(u2__abc_52155_new_n15576_), .Y(u2__abc_52155_new_n15577_));
OR2X2 OR2X2_3291 ( .A(u2__abc_52155_new_n15578_), .B(u2__abc_52155_new_n15577_), .Y(u2__abc_52155_new_n15579_));
OR2X2 OR2X2_3292 ( .A(u2__abc_52155_new_n15579_), .B(u2__abc_52155_new_n7367_), .Y(u2__abc_52155_new_n15582_));
OR2X2 OR2X2_3293 ( .A(u2__abc_52155_new_n15585_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15586_));
OR2X2 OR2X2_3294 ( .A(u2__abc_52155_new_n15584_), .B(u2__abc_52155_new_n15586_), .Y(u2__abc_52155_new_n15587_));
OR2X2 OR2X2_3295 ( .A(u2__abc_52155_new_n15591_), .B(u2__abc_52155_new_n15573_), .Y(u2__abc_52155_new_n15592_));
OR2X2 OR2X2_3296 ( .A(u2__abc_52155_new_n15599_), .B(u2__abc_52155_new_n15596_), .Y(u2__abc_52155_new_n15600_));
OR2X2 OR2X2_3297 ( .A(u2__abc_52155_new_n15602_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15603_));
OR2X2 OR2X2_3298 ( .A(u2__abc_52155_new_n15601_), .B(u2__abc_52155_new_n15603_), .Y(u2__abc_52155_new_n15604_));
OR2X2 OR2X2_3299 ( .A(u2__abc_52155_new_n15608_), .B(u2__abc_52155_new_n15594_), .Y(u2__abc_52155_new_n15609_));
OR2X2 OR2X2_33 ( .A(aNan), .B(sqrto_92_), .Y(_abc_73687_new_n878_));
OR2X2 OR2X2_330 ( .A(\a[112] ), .B(\a[52] ), .Y(_abc_73687_new_n1326_));
OR2X2 OR2X2_3300 ( .A(u2__abc_52155_new_n15613_), .B(u2__abc_52155_new_n7355_), .Y(u2__abc_52155_new_n15614_));
OR2X2 OR2X2_3301 ( .A(u2__abc_52155_new_n15615_), .B(u2__abc_52155_new_n7345_), .Y(u2__abc_52155_new_n15618_));
OR2X2 OR2X2_3302 ( .A(u2__abc_52155_new_n15621_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15622_));
OR2X2 OR2X2_3303 ( .A(u2__abc_52155_new_n15620_), .B(u2__abc_52155_new_n15622_), .Y(u2__abc_52155_new_n15623_));
OR2X2 OR2X2_3304 ( .A(u2__abc_52155_new_n15627_), .B(u2__abc_52155_new_n15611_), .Y(u2__abc_52155_new_n15628_));
OR2X2 OR2X2_3305 ( .A(u2__abc_52155_new_n15632_), .B(u2__abc_52155_new_n15631_), .Y(u2__abc_52155_new_n15633_));
OR2X2 OR2X2_3306 ( .A(u2__abc_52155_new_n15634_), .B(u2__abc_52155_new_n7352_), .Y(u2__abc_52155_new_n15635_));
OR2X2 OR2X2_3307 ( .A(u2__abc_52155_new_n15638_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15639_));
OR2X2 OR2X2_3308 ( .A(u2__abc_52155_new_n15637_), .B(u2__abc_52155_new_n15639_), .Y(u2__abc_52155_new_n15640_));
OR2X2 OR2X2_3309 ( .A(u2__abc_52155_new_n15644_), .B(u2__abc_52155_new_n15630_), .Y(u2__abc_52155_new_n15645_));
OR2X2 OR2X2_331 ( .A(_abc_73687_new_n1170_), .B(\a[53] ), .Y(_abc_73687_new_n1327_));
OR2X2 OR2X2_3310 ( .A(u2__abc_52155_new_n15612_), .B(u2__abc_52155_new_n7355_), .Y(u2__abc_52155_new_n15649_));
OR2X2 OR2X2_3311 ( .A(u2__abc_52155_new_n15652_), .B(u2__abc_52155_new_n7347_), .Y(u2__abc_52155_new_n15653_));
OR2X2 OR2X2_3312 ( .A(u2__abc_52155_new_n15651_), .B(u2__abc_52155_new_n15653_), .Y(u2__abc_52155_new_n15654_));
OR2X2 OR2X2_3313 ( .A(u2__abc_52155_new_n15648_), .B(u2__abc_52155_new_n15654_), .Y(u2__abc_52155_new_n15655_));
OR2X2 OR2X2_3314 ( .A(u2__abc_52155_new_n15656_), .B(u2__abc_52155_new_n15655_), .Y(u2__abc_52155_new_n15657_));
OR2X2 OR2X2_3315 ( .A(u2__abc_52155_new_n15657_), .B(u2__abc_52155_new_n7273_), .Y(u2__abc_52155_new_n15660_));
OR2X2 OR2X2_3316 ( .A(u2__abc_52155_new_n15663_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15664_));
OR2X2 OR2X2_3317 ( .A(u2__abc_52155_new_n15662_), .B(u2__abc_52155_new_n15664_), .Y(u2__abc_52155_new_n15665_));
OR2X2 OR2X2_3318 ( .A(u2__abc_52155_new_n15669_), .B(u2__abc_52155_new_n15647_), .Y(u2__abc_52155_new_n15670_));
OR2X2 OR2X2_3319 ( .A(u2__abc_52155_new_n15677_), .B(u2__abc_52155_new_n15674_), .Y(u2__abc_52155_new_n15678_));
OR2X2 OR2X2_332 ( .A(\a[112] ), .B(\a[53] ), .Y(_abc_73687_new_n1329_));
OR2X2 OR2X2_3320 ( .A(u2__abc_52155_new_n15680_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15681_));
OR2X2 OR2X2_3321 ( .A(u2__abc_52155_new_n15679_), .B(u2__abc_52155_new_n15681_), .Y(u2__abc_52155_new_n15682_));
OR2X2 OR2X2_3322 ( .A(u2__abc_52155_new_n15686_), .B(u2__abc_52155_new_n15672_), .Y(u2__abc_52155_new_n15687_));
OR2X2 OR2X2_3323 ( .A(u2__abc_52155_new_n15691_), .B(u2__abc_52155_new_n7261_), .Y(u2__abc_52155_new_n15692_));
OR2X2 OR2X2_3324 ( .A(u2__abc_52155_new_n15693_), .B(u2__abc_52155_new_n7251_), .Y(u2__abc_52155_new_n15696_));
OR2X2 OR2X2_3325 ( .A(u2__abc_52155_new_n15699_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15700_));
OR2X2 OR2X2_3326 ( .A(u2__abc_52155_new_n15698_), .B(u2__abc_52155_new_n15700_), .Y(u2__abc_52155_new_n15701_));
OR2X2 OR2X2_3327 ( .A(u2__abc_52155_new_n15705_), .B(u2__abc_52155_new_n15689_), .Y(u2__abc_52155_new_n15706_));
OR2X2 OR2X2_3328 ( .A(u2__abc_52155_new_n15710_), .B(u2__abc_52155_new_n15709_), .Y(u2__abc_52155_new_n15711_));
OR2X2 OR2X2_3329 ( .A(u2__abc_52155_new_n15712_), .B(u2__abc_52155_new_n7258_), .Y(u2__abc_52155_new_n15713_));
OR2X2 OR2X2_333 ( .A(_abc_73687_new_n1170_), .B(\a[54] ), .Y(_abc_73687_new_n1330_));
OR2X2 OR2X2_3330 ( .A(u2__abc_52155_new_n15716_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15717_));
OR2X2 OR2X2_3331 ( .A(u2__abc_52155_new_n15715_), .B(u2__abc_52155_new_n15717_), .Y(u2__abc_52155_new_n15718_));
OR2X2 OR2X2_3332 ( .A(u2__abc_52155_new_n15722_), .B(u2__abc_52155_new_n15708_), .Y(u2__abc_52155_new_n15723_));
OR2X2 OR2X2_3333 ( .A(u2__abc_52155_new_n15690_), .B(u2__abc_52155_new_n7261_), .Y(u2__abc_52155_new_n15726_));
OR2X2 OR2X2_3334 ( .A(u2__abc_52155_new_n15729_), .B(u2__abc_52155_new_n7256_), .Y(u2__abc_52155_new_n15730_));
OR2X2 OR2X2_3335 ( .A(u2__abc_52155_new_n15728_), .B(u2__abc_52155_new_n15730_), .Y(u2__abc_52155_new_n15731_));
OR2X2 OR2X2_3336 ( .A(u2__abc_52155_new_n15732_), .B(u2__abc_52155_new_n15731_), .Y(u2__abc_52155_new_n15733_));
OR2X2 OR2X2_3337 ( .A(u2__abc_52155_new_n15733_), .B(u2__abc_52155_new_n7304_), .Y(u2__abc_52155_new_n15736_));
OR2X2 OR2X2_3338 ( .A(u2__abc_52155_new_n15739_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15740_));
OR2X2 OR2X2_3339 ( .A(u2__abc_52155_new_n15738_), .B(u2__abc_52155_new_n15740_), .Y(u2__abc_52155_new_n15741_));
OR2X2 OR2X2_334 ( .A(\a[112] ), .B(\a[54] ), .Y(_abc_73687_new_n1332_));
OR2X2 OR2X2_3340 ( .A(u2__abc_52155_new_n15745_), .B(u2__abc_52155_new_n15725_), .Y(u2__abc_52155_new_n15746_));
OR2X2 OR2X2_3341 ( .A(u2__abc_52155_new_n15753_), .B(u2__abc_52155_new_n15750_), .Y(u2__abc_52155_new_n15754_));
OR2X2 OR2X2_3342 ( .A(u2__abc_52155_new_n15756_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15757_));
OR2X2 OR2X2_3343 ( .A(u2__abc_52155_new_n15755_), .B(u2__abc_52155_new_n15757_), .Y(u2__abc_52155_new_n15758_));
OR2X2 OR2X2_3344 ( .A(u2__abc_52155_new_n15762_), .B(u2__abc_52155_new_n15748_), .Y(u2__abc_52155_new_n15763_));
OR2X2 OR2X2_3345 ( .A(u2__abc_52155_new_n15767_), .B(u2__abc_52155_new_n7292_), .Y(u2__abc_52155_new_n15768_));
OR2X2 OR2X2_3346 ( .A(u2__abc_52155_new_n15769_), .B(u2__abc_52155_new_n7282_), .Y(u2__abc_52155_new_n15772_));
OR2X2 OR2X2_3347 ( .A(u2__abc_52155_new_n15775_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15776_));
OR2X2 OR2X2_3348 ( .A(u2__abc_52155_new_n15774_), .B(u2__abc_52155_new_n15776_), .Y(u2__abc_52155_new_n15777_));
OR2X2 OR2X2_3349 ( .A(u2__abc_52155_new_n15781_), .B(u2__abc_52155_new_n15765_), .Y(u2__abc_52155_new_n15782_));
OR2X2 OR2X2_335 ( .A(_abc_73687_new_n1170_), .B(\a[55] ), .Y(_abc_73687_new_n1333_));
OR2X2 OR2X2_3350 ( .A(u2__abc_52155_new_n15786_), .B(u2__abc_52155_new_n15785_), .Y(u2__abc_52155_new_n15787_));
OR2X2 OR2X2_3351 ( .A(u2__abc_52155_new_n15788_), .B(u2__abc_52155_new_n7289_), .Y(u2__abc_52155_new_n15789_));
OR2X2 OR2X2_3352 ( .A(u2__abc_52155_new_n15792_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15793_));
OR2X2 OR2X2_3353 ( .A(u2__abc_52155_new_n15791_), .B(u2__abc_52155_new_n15793_), .Y(u2__abc_52155_new_n15794_));
OR2X2 OR2X2_3354 ( .A(u2__abc_52155_new_n15798_), .B(u2__abc_52155_new_n15784_), .Y(u2__abc_52155_new_n15799_));
OR2X2 OR2X2_3355 ( .A(u2__abc_52155_new_n15766_), .B(u2__abc_52155_new_n7292_), .Y(u2__abc_52155_new_n15804_));
OR2X2 OR2X2_3356 ( .A(u2__abc_52155_new_n15807_), .B(u2__abc_52155_new_n7284_), .Y(u2__abc_52155_new_n15808_));
OR2X2 OR2X2_3357 ( .A(u2__abc_52155_new_n15806_), .B(u2__abc_52155_new_n15808_), .Y(u2__abc_52155_new_n15809_));
OR2X2 OR2X2_3358 ( .A(u2__abc_52155_new_n15803_), .B(u2__abc_52155_new_n15809_), .Y(u2__abc_52155_new_n15810_));
OR2X2 OR2X2_3359 ( .A(u2__abc_52155_new_n15811_), .B(u2__abc_52155_new_n15810_), .Y(u2__abc_52155_new_n15812_));
OR2X2 OR2X2_336 ( .A(\a[112] ), .B(\a[55] ), .Y(_abc_73687_new_n1335_));
OR2X2 OR2X2_3360 ( .A(u2__abc_52155_new_n15814_), .B(u2__abc_52155_new_n15813_), .Y(u2__abc_52155_new_n15815_));
OR2X2 OR2X2_3361 ( .A(u2__abc_52155_new_n15815_), .B(u2__abc_52155_new_n15812_), .Y(u2__abc_52155_new_n15816_));
OR2X2 OR2X2_3362 ( .A(u2__abc_52155_new_n15802_), .B(u2__abc_52155_new_n15816_), .Y(u2__abc_52155_new_n15817_));
OR2X2 OR2X2_3363 ( .A(u2__abc_52155_new_n15817_), .B(u2__abc_52155_new_n7176_), .Y(u2__abc_52155_new_n15820_));
OR2X2 OR2X2_3364 ( .A(u2__abc_52155_new_n15823_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15824_));
OR2X2 OR2X2_3365 ( .A(u2__abc_52155_new_n15822_), .B(u2__abc_52155_new_n15824_), .Y(u2__abc_52155_new_n15825_));
OR2X2 OR2X2_3366 ( .A(u2__abc_52155_new_n15829_), .B(u2__abc_52155_new_n15801_), .Y(u2__abc_52155_new_n15830_));
OR2X2 OR2X2_3367 ( .A(u2__abc_52155_new_n15837_), .B(u2__abc_52155_new_n15834_), .Y(u2__abc_52155_new_n15838_));
OR2X2 OR2X2_3368 ( .A(u2__abc_52155_new_n15840_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15841_));
OR2X2 OR2X2_3369 ( .A(u2__abc_52155_new_n15839_), .B(u2__abc_52155_new_n15841_), .Y(u2__abc_52155_new_n15842_));
OR2X2 OR2X2_337 ( .A(_abc_73687_new_n1170_), .B(\a[56] ), .Y(_abc_73687_new_n1336_));
OR2X2 OR2X2_3370 ( .A(u2__abc_52155_new_n15846_), .B(u2__abc_52155_new_n15832_), .Y(u2__abc_52155_new_n15847_));
OR2X2 OR2X2_3371 ( .A(u2__abc_52155_new_n15851_), .B(u2__abc_52155_new_n7164_), .Y(u2__abc_52155_new_n15852_));
OR2X2 OR2X2_3372 ( .A(u2__abc_52155_new_n15853_), .B(u2__abc_52155_new_n7154_), .Y(u2__abc_52155_new_n15856_));
OR2X2 OR2X2_3373 ( .A(u2__abc_52155_new_n15859_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15860_));
OR2X2 OR2X2_3374 ( .A(u2__abc_52155_new_n15858_), .B(u2__abc_52155_new_n15860_), .Y(u2__abc_52155_new_n15861_));
OR2X2 OR2X2_3375 ( .A(u2__abc_52155_new_n15865_), .B(u2__abc_52155_new_n15849_), .Y(u2__abc_52155_new_n15866_));
OR2X2 OR2X2_3376 ( .A(u2__abc_52155_new_n15870_), .B(u2__abc_52155_new_n15869_), .Y(u2__abc_52155_new_n15871_));
OR2X2 OR2X2_3377 ( .A(u2__abc_52155_new_n15872_), .B(u2__abc_52155_new_n7161_), .Y(u2__abc_52155_new_n15873_));
OR2X2 OR2X2_3378 ( .A(u2__abc_52155_new_n15876_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15877_));
OR2X2 OR2X2_3379 ( .A(u2__abc_52155_new_n15875_), .B(u2__abc_52155_new_n15877_), .Y(u2__abc_52155_new_n15878_));
OR2X2 OR2X2_338 ( .A(\a[112] ), .B(\a[56] ), .Y(_abc_73687_new_n1338_));
OR2X2 OR2X2_3380 ( .A(u2__abc_52155_new_n15882_), .B(u2__abc_52155_new_n15868_), .Y(u2__abc_52155_new_n15883_));
OR2X2 OR2X2_3381 ( .A(u2__abc_52155_new_n15850_), .B(u2__abc_52155_new_n7164_), .Y(u2__abc_52155_new_n15886_));
OR2X2 OR2X2_3382 ( .A(u2__abc_52155_new_n15889_), .B(u2__abc_52155_new_n7159_), .Y(u2__abc_52155_new_n15890_));
OR2X2 OR2X2_3383 ( .A(u2__abc_52155_new_n15888_), .B(u2__abc_52155_new_n15890_), .Y(u2__abc_52155_new_n15891_));
OR2X2 OR2X2_3384 ( .A(u2__abc_52155_new_n15892_), .B(u2__abc_52155_new_n15891_), .Y(u2__abc_52155_new_n15893_));
OR2X2 OR2X2_3385 ( .A(u2__abc_52155_new_n15893_), .B(u2__abc_52155_new_n7145_), .Y(u2__abc_52155_new_n15896_));
OR2X2 OR2X2_3386 ( .A(u2__abc_52155_new_n15899_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15900_));
OR2X2 OR2X2_3387 ( .A(u2__abc_52155_new_n15898_), .B(u2__abc_52155_new_n15900_), .Y(u2__abc_52155_new_n15901_));
OR2X2 OR2X2_3388 ( .A(u2__abc_52155_new_n15905_), .B(u2__abc_52155_new_n15885_), .Y(u2__abc_52155_new_n15906_));
OR2X2 OR2X2_3389 ( .A(u2__abc_52155_new_n15913_), .B(u2__abc_52155_new_n15910_), .Y(u2__abc_52155_new_n15914_));
OR2X2 OR2X2_339 ( .A(_abc_73687_new_n1170_), .B(\a[57] ), .Y(_abc_73687_new_n1339_));
OR2X2 OR2X2_3390 ( .A(u2__abc_52155_new_n15916_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15917_));
OR2X2 OR2X2_3391 ( .A(u2__abc_52155_new_n15915_), .B(u2__abc_52155_new_n15917_), .Y(u2__abc_52155_new_n15918_));
OR2X2 OR2X2_3392 ( .A(u2__abc_52155_new_n15922_), .B(u2__abc_52155_new_n15908_), .Y(u2__abc_52155_new_n15923_));
OR2X2 OR2X2_3393 ( .A(u2__abc_52155_new_n15927_), .B(u2__abc_52155_new_n7133_), .Y(u2__abc_52155_new_n15928_));
OR2X2 OR2X2_3394 ( .A(u2__abc_52155_new_n15929_), .B(u2__abc_52155_new_n7123_), .Y(u2__abc_52155_new_n15932_));
OR2X2 OR2X2_3395 ( .A(u2__abc_52155_new_n15935_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15936_));
OR2X2 OR2X2_3396 ( .A(u2__abc_52155_new_n15934_), .B(u2__abc_52155_new_n15936_), .Y(u2__abc_52155_new_n15937_));
OR2X2 OR2X2_3397 ( .A(u2__abc_52155_new_n15941_), .B(u2__abc_52155_new_n15925_), .Y(u2__abc_52155_new_n15942_));
OR2X2 OR2X2_3398 ( .A(u2__abc_52155_new_n15946_), .B(u2__abc_52155_new_n15945_), .Y(u2__abc_52155_new_n15947_));
OR2X2 OR2X2_3399 ( .A(u2__abc_52155_new_n15948_), .B(u2__abc_52155_new_n7130_), .Y(u2__abc_52155_new_n15949_));
OR2X2 OR2X2_34 ( .A(_abc_73687_new_n753_), .B(\a[16] ), .Y(_abc_73687_new_n879_));
OR2X2 OR2X2_340 ( .A(\a[112] ), .B(\a[57] ), .Y(_abc_73687_new_n1341_));
OR2X2 OR2X2_3400 ( .A(u2__abc_52155_new_n15952_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15953_));
OR2X2 OR2X2_3401 ( .A(u2__abc_52155_new_n15951_), .B(u2__abc_52155_new_n15953_), .Y(u2__abc_52155_new_n15954_));
OR2X2 OR2X2_3402 ( .A(u2__abc_52155_new_n15958_), .B(u2__abc_52155_new_n15944_), .Y(u2__abc_52155_new_n15959_));
OR2X2 OR2X2_3403 ( .A(u2__abc_52155_new_n15926_), .B(u2__abc_52155_new_n7133_), .Y(u2__abc_52155_new_n15963_));
OR2X2 OR2X2_3404 ( .A(u2__abc_52155_new_n15966_), .B(u2__abc_52155_new_n7125_), .Y(u2__abc_52155_new_n15967_));
OR2X2 OR2X2_3405 ( .A(u2__abc_52155_new_n15965_), .B(u2__abc_52155_new_n15967_), .Y(u2__abc_52155_new_n15968_));
OR2X2 OR2X2_3406 ( .A(u2__abc_52155_new_n15962_), .B(u2__abc_52155_new_n15968_), .Y(u2__abc_52155_new_n15969_));
OR2X2 OR2X2_3407 ( .A(u2__abc_52155_new_n15970_), .B(u2__abc_52155_new_n15969_), .Y(u2__abc_52155_new_n15971_));
OR2X2 OR2X2_3408 ( .A(u2__abc_52155_new_n15971_), .B(u2__abc_52155_new_n7075_), .Y(u2__abc_52155_new_n15974_));
OR2X2 OR2X2_3409 ( .A(u2__abc_52155_new_n15977_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15978_));
OR2X2 OR2X2_341 ( .A(_abc_73687_new_n1170_), .B(\a[58] ), .Y(_abc_73687_new_n1342_));
OR2X2 OR2X2_3410 ( .A(u2__abc_52155_new_n15976_), .B(u2__abc_52155_new_n15978_), .Y(u2__abc_52155_new_n15979_));
OR2X2 OR2X2_3411 ( .A(u2__abc_52155_new_n15983_), .B(u2__abc_52155_new_n15961_), .Y(u2__abc_52155_new_n15984_));
OR2X2 OR2X2_3412 ( .A(u2__abc_52155_new_n15990_), .B(u2__abc_52155_new_n15991_), .Y(u2__abc_52155_new_n15992_));
OR2X2 OR2X2_3413 ( .A(u2__abc_52155_new_n15994_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n15995_));
OR2X2 OR2X2_3414 ( .A(u2__abc_52155_new_n15993_), .B(u2__abc_52155_new_n15995_), .Y(u2__abc_52155_new_n15996_));
OR2X2 OR2X2_3415 ( .A(u2__abc_52155_new_n16000_), .B(u2__abc_52155_new_n15986_), .Y(u2__abc_52155_new_n16001_));
OR2X2 OR2X2_3416 ( .A(u2__abc_52155_new_n16004_), .B(u2__abc_52155_new_n7080_), .Y(u2__abc_52155_new_n16005_));
OR2X2 OR2X2_3417 ( .A(u2__abc_52155_new_n16005_), .B(u2__abc_52155_new_n7060_), .Y(u2__abc_52155_new_n16008_));
OR2X2 OR2X2_3418 ( .A(u2__abc_52155_new_n16011_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16012_));
OR2X2 OR2X2_3419 ( .A(u2__abc_52155_new_n16010_), .B(u2__abc_52155_new_n16012_), .Y(u2__abc_52155_new_n16013_));
OR2X2 OR2X2_342 ( .A(\a[112] ), .B(\a[58] ), .Y(_abc_73687_new_n1344_));
OR2X2 OR2X2_3420 ( .A(u2__abc_52155_new_n16017_), .B(u2__abc_52155_new_n16003_), .Y(u2__abc_52155_new_n16018_));
OR2X2 OR2X2_3421 ( .A(u2__abc_52155_new_n16022_), .B(u2__abc_52155_new_n16021_), .Y(u2__abc_52155_new_n16023_));
OR2X2 OR2X2_3422 ( .A(u2__abc_52155_new_n16024_), .B(u2__abc_52155_new_n7067_), .Y(u2__abc_52155_new_n16025_));
OR2X2 OR2X2_3423 ( .A(u2__abc_52155_new_n16028_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16029_));
OR2X2 OR2X2_3424 ( .A(u2__abc_52155_new_n16027_), .B(u2__abc_52155_new_n16029_), .Y(u2__abc_52155_new_n16030_));
OR2X2 OR2X2_3425 ( .A(u2__abc_52155_new_n16034_), .B(u2__abc_52155_new_n16020_), .Y(u2__abc_52155_new_n16035_));
OR2X2 OR2X2_3426 ( .A(u2__abc_52155_new_n16038_), .B(u2__abc_52155_new_n7077_), .Y(u2__abc_52155_new_n16039_));
OR2X2 OR2X2_3427 ( .A(u2__abc_52155_new_n16042_), .B(u2__abc_52155_new_n7065_), .Y(u2__abc_52155_new_n16043_));
OR2X2 OR2X2_3428 ( .A(u2__abc_52155_new_n16041_), .B(u2__abc_52155_new_n16043_), .Y(u2__abc_52155_new_n16044_));
OR2X2 OR2X2_3429 ( .A(u2__abc_52155_new_n16045_), .B(u2__abc_52155_new_n16044_), .Y(u2__abc_52155_new_n16046_));
OR2X2 OR2X2_343 ( .A(_abc_73687_new_n1170_), .B(\a[59] ), .Y(_abc_73687_new_n1345_));
OR2X2 OR2X2_3430 ( .A(u2__abc_52155_new_n16046_), .B(u2__abc_52155_new_n7113_), .Y(u2__abc_52155_new_n16049_));
OR2X2 OR2X2_3431 ( .A(u2__abc_52155_new_n16052_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16053_));
OR2X2 OR2X2_3432 ( .A(u2__abc_52155_new_n16051_), .B(u2__abc_52155_new_n16053_), .Y(u2__abc_52155_new_n16054_));
OR2X2 OR2X2_3433 ( .A(u2__abc_52155_new_n16058_), .B(u2__abc_52155_new_n16037_), .Y(u2__abc_52155_new_n16059_));
OR2X2 OR2X2_3434 ( .A(u2__abc_52155_new_n16066_), .B(u2__abc_52155_new_n16063_), .Y(u2__abc_52155_new_n16067_));
OR2X2 OR2X2_3435 ( .A(u2__abc_52155_new_n16069_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16070_));
OR2X2 OR2X2_3436 ( .A(u2__abc_52155_new_n16068_), .B(u2__abc_52155_new_n16070_), .Y(u2__abc_52155_new_n16071_));
OR2X2 OR2X2_3437 ( .A(u2__abc_52155_new_n16075_), .B(u2__abc_52155_new_n16061_), .Y(u2__abc_52155_new_n16076_));
OR2X2 OR2X2_3438 ( .A(u2__abc_52155_new_n16080_), .B(u2__abc_52155_new_n7101_), .Y(u2__abc_52155_new_n16081_));
OR2X2 OR2X2_3439 ( .A(u2__abc_52155_new_n16082_), .B(u2__abc_52155_new_n7091_), .Y(u2__abc_52155_new_n16085_));
OR2X2 OR2X2_344 ( .A(\a[112] ), .B(\a[59] ), .Y(_abc_73687_new_n1347_));
OR2X2 OR2X2_3440 ( .A(u2__abc_52155_new_n16088_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16089_));
OR2X2 OR2X2_3441 ( .A(u2__abc_52155_new_n16087_), .B(u2__abc_52155_new_n16089_), .Y(u2__abc_52155_new_n16090_));
OR2X2 OR2X2_3442 ( .A(u2__abc_52155_new_n16094_), .B(u2__abc_52155_new_n16078_), .Y(u2__abc_52155_new_n16095_));
OR2X2 OR2X2_3443 ( .A(u2__abc_52155_new_n16099_), .B(u2__abc_52155_new_n16098_), .Y(u2__abc_52155_new_n16100_));
OR2X2 OR2X2_3444 ( .A(u2__abc_52155_new_n16101_), .B(u2__abc_52155_new_n7098_), .Y(u2__abc_52155_new_n16102_));
OR2X2 OR2X2_3445 ( .A(u2__abc_52155_new_n16105_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16106_));
OR2X2 OR2X2_3446 ( .A(u2__abc_52155_new_n16104_), .B(u2__abc_52155_new_n16106_), .Y(u2__abc_52155_new_n16107_));
OR2X2 OR2X2_3447 ( .A(u2__abc_52155_new_n16111_), .B(u2__abc_52155_new_n16097_), .Y(u2__abc_52155_new_n16112_));
OR2X2 OR2X2_3448 ( .A(u2__abc_52155_new_n16079_), .B(u2__abc_52155_new_n7101_), .Y(u2__abc_52155_new_n16117_));
OR2X2 OR2X2_3449 ( .A(u2__abc_52155_new_n16120_), .B(u2__abc_52155_new_n7093_), .Y(u2__abc_52155_new_n16121_));
OR2X2 OR2X2_345 ( .A(_abc_73687_new_n1170_), .B(\a[60] ), .Y(_abc_73687_new_n1348_));
OR2X2 OR2X2_3450 ( .A(u2__abc_52155_new_n16119_), .B(u2__abc_52155_new_n16121_), .Y(u2__abc_52155_new_n16122_));
OR2X2 OR2X2_3451 ( .A(u2__abc_52155_new_n16116_), .B(u2__abc_52155_new_n16122_), .Y(u2__abc_52155_new_n16123_));
OR2X2 OR2X2_3452 ( .A(u2__abc_52155_new_n16115_), .B(u2__abc_52155_new_n16123_), .Y(u2__abc_52155_new_n16124_));
OR2X2 OR2X2_3453 ( .A(u2__abc_52155_new_n16125_), .B(u2__abc_52155_new_n16124_), .Y(u2__abc_52155_new_n16126_));
OR2X2 OR2X2_3454 ( .A(u2__abc_52155_new_n16126_), .B(u2__abc_52155_new_n7027_), .Y(u2__abc_52155_new_n16129_));
OR2X2 OR2X2_3455 ( .A(u2__abc_52155_new_n16132_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16133_));
OR2X2 OR2X2_3456 ( .A(u2__abc_52155_new_n16131_), .B(u2__abc_52155_new_n16133_), .Y(u2__abc_52155_new_n16134_));
OR2X2 OR2X2_3457 ( .A(u2__abc_52155_new_n16138_), .B(u2__abc_52155_new_n16114_), .Y(u2__abc_52155_new_n16139_));
OR2X2 OR2X2_3458 ( .A(u2__abc_52155_new_n16143_), .B(u2__abc_52155_new_n16142_), .Y(u2__abc_52155_new_n16144_));
OR2X2 OR2X2_3459 ( .A(u2__abc_52155_new_n16145_), .B(u2__abc_52155_new_n7034_), .Y(u2__abc_52155_new_n16146_));
OR2X2 OR2X2_346 ( .A(\a[112] ), .B(\a[60] ), .Y(_abc_73687_new_n1350_));
OR2X2 OR2X2_3460 ( .A(u2__abc_52155_new_n16149_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16150_));
OR2X2 OR2X2_3461 ( .A(u2__abc_52155_new_n16148_), .B(u2__abc_52155_new_n16150_), .Y(u2__abc_52155_new_n16151_));
OR2X2 OR2X2_3462 ( .A(u2__abc_52155_new_n16155_), .B(u2__abc_52155_new_n16141_), .Y(u2__abc_52155_new_n16156_));
OR2X2 OR2X2_3463 ( .A(u2__abc_52155_new_n7023_), .B(u2__abc_52155_new_n7029_), .Y(u2__abc_52155_new_n16159_));
OR2X2 OR2X2_3464 ( .A(u2__abc_52155_new_n16162_), .B(u2__abc_52155_new_n16161_), .Y(u2__abc_52155_new_n16163_));
OR2X2 OR2X2_3465 ( .A(u2__abc_52155_new_n16163_), .B(u2__abc_52155_new_n7042_), .Y(u2__abc_52155_new_n16166_));
OR2X2 OR2X2_3466 ( .A(u2__abc_52155_new_n16169_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16170_));
OR2X2 OR2X2_3467 ( .A(u2__abc_52155_new_n16168_), .B(u2__abc_52155_new_n16170_), .Y(u2__abc_52155_new_n16171_));
OR2X2 OR2X2_3468 ( .A(u2__abc_52155_new_n16175_), .B(u2__abc_52155_new_n16158_), .Y(u2__abc_52155_new_n16176_));
OR2X2 OR2X2_3469 ( .A(u2__abc_52155_new_n16180_), .B(u2__abc_52155_new_n16179_), .Y(u2__abc_52155_new_n16181_));
OR2X2 OR2X2_347 ( .A(_abc_73687_new_n1170_), .B(\a[61] ), .Y(_abc_73687_new_n1351_));
OR2X2 OR2X2_3470 ( .A(u2__abc_52155_new_n16182_), .B(u2__abc_52155_new_n7049_), .Y(u2__abc_52155_new_n16183_));
OR2X2 OR2X2_3471 ( .A(u2__abc_52155_new_n16186_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16187_));
OR2X2 OR2X2_3472 ( .A(u2__abc_52155_new_n16185_), .B(u2__abc_52155_new_n16187_), .Y(u2__abc_52155_new_n16188_));
OR2X2 OR2X2_3473 ( .A(u2__abc_52155_new_n16192_), .B(u2__abc_52155_new_n16178_), .Y(u2__abc_52155_new_n16193_));
OR2X2 OR2X2_3474 ( .A(u2__abc_52155_new_n16197_), .B(u2__abc_52155_new_n7044_), .Y(u2__abc_52155_new_n16198_));
OR2X2 OR2X2_3475 ( .A(u2__abc_52155_new_n16199_), .B(u2__abc_52155_new_n7018_), .Y(u2__abc_52155_new_n16202_));
OR2X2 OR2X2_3476 ( .A(u2__abc_52155_new_n16205_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16206_));
OR2X2 OR2X2_3477 ( .A(u2__abc_52155_new_n16204_), .B(u2__abc_52155_new_n16206_), .Y(u2__abc_52155_new_n16207_));
OR2X2 OR2X2_3478 ( .A(u2__abc_52155_new_n16211_), .B(u2__abc_52155_new_n16195_), .Y(u2__abc_52155_new_n16212_));
OR2X2 OR2X2_3479 ( .A(u2__abc_52155_new_n16216_), .B(u2__abc_52155_new_n7011_), .Y(u2__abc_52155_new_n16219_));
OR2X2 OR2X2_348 ( .A(\a[112] ), .B(\a[61] ), .Y(_abc_73687_new_n1353_));
OR2X2 OR2X2_3480 ( .A(u2__abc_52155_new_n16222_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16223_));
OR2X2 OR2X2_3481 ( .A(u2__abc_52155_new_n16221_), .B(u2__abc_52155_new_n16223_), .Y(u2__abc_52155_new_n16224_));
OR2X2 OR2X2_3482 ( .A(u2__abc_52155_new_n16228_), .B(u2__abc_52155_new_n16214_), .Y(u2__abc_52155_new_n16229_));
OR2X2 OR2X2_3483 ( .A(u2__abc_52155_new_n16233_), .B(u2__abc_52155_new_n6996_), .Y(u2__abc_52155_new_n16236_));
OR2X2 OR2X2_3484 ( .A(u2__abc_52155_new_n16239_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16240_));
OR2X2 OR2X2_3485 ( .A(u2__abc_52155_new_n16238_), .B(u2__abc_52155_new_n16240_), .Y(u2__abc_52155_new_n16241_));
OR2X2 OR2X2_3486 ( .A(u2__abc_52155_new_n16245_), .B(u2__abc_52155_new_n16231_), .Y(u2__abc_52155_new_n16246_));
OR2X2 OR2X2_3487 ( .A(u2__abc_52155_new_n16250_), .B(u2__abc_52155_new_n16249_), .Y(u2__abc_52155_new_n16251_));
OR2X2 OR2X2_3488 ( .A(u2__abc_52155_new_n16252_), .B(u2__abc_52155_new_n7003_), .Y(u2__abc_52155_new_n16253_));
OR2X2 OR2X2_3489 ( .A(u2__abc_52155_new_n16256_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16257_));
OR2X2 OR2X2_349 ( .A(_abc_73687_new_n1170_), .B(\a[62] ), .Y(_abc_73687_new_n1354_));
OR2X2 OR2X2_3490 ( .A(u2__abc_52155_new_n16255_), .B(u2__abc_52155_new_n16257_), .Y(u2__abc_52155_new_n16258_));
OR2X2 OR2X2_3491 ( .A(u2__abc_52155_new_n16262_), .B(u2__abc_52155_new_n16248_), .Y(u2__abc_52155_new_n16263_));
OR2X2 OR2X2_3492 ( .A(u2__abc_52155_new_n16196_), .B(u2__abc_52155_new_n7044_), .Y(u2__abc_52155_new_n16266_));
OR2X2 OR2X2_3493 ( .A(u2__abc_52155_new_n16272_), .B(u2__abc_52155_new_n7006_), .Y(u2__abc_52155_new_n16273_));
OR2X2 OR2X2_3494 ( .A(u2__abc_52155_new_n16276_), .B(u2__abc_52155_new_n6998_), .Y(u2__abc_52155_new_n16277_));
OR2X2 OR2X2_3495 ( .A(u2__abc_52155_new_n16275_), .B(u2__abc_52155_new_n16277_), .Y(u2__abc_52155_new_n16278_));
OR2X2 OR2X2_3496 ( .A(u2__abc_52155_new_n16271_), .B(u2__abc_52155_new_n16278_), .Y(u2__abc_52155_new_n16279_));
OR2X2 OR2X2_3497 ( .A(u2__abc_52155_new_n16280_), .B(u2__abc_52155_new_n16279_), .Y(u2__abc_52155_new_n16281_));
OR2X2 OR2X2_3498 ( .A(u2__abc_52155_new_n16281_), .B(u2__abc_52155_new_n6964_), .Y(u2__abc_52155_new_n16284_));
OR2X2 OR2X2_3499 ( .A(u2__abc_52155_new_n16287_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16288_));
OR2X2 OR2X2_35 ( .A(aNan), .B(sqrto_93_), .Y(_abc_73687_new_n881_));
OR2X2 OR2X2_350 ( .A(\a[112] ), .B(\a[62] ), .Y(_abc_73687_new_n1356_));
OR2X2 OR2X2_3500 ( .A(u2__abc_52155_new_n16286_), .B(u2__abc_52155_new_n16288_), .Y(u2__abc_52155_new_n16289_));
OR2X2 OR2X2_3501 ( .A(u2__abc_52155_new_n16293_), .B(u2__abc_52155_new_n16265_), .Y(u2__abc_52155_new_n16294_));
OR2X2 OR2X2_3502 ( .A(u2__abc_52155_new_n16298_), .B(u2__abc_52155_new_n16297_), .Y(u2__abc_52155_new_n16299_));
OR2X2 OR2X2_3503 ( .A(u2__abc_52155_new_n16300_), .B(u2__abc_52155_new_n6971_), .Y(u2__abc_52155_new_n16301_));
OR2X2 OR2X2_3504 ( .A(u2__abc_52155_new_n16304_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16305_));
OR2X2 OR2X2_3505 ( .A(u2__abc_52155_new_n16303_), .B(u2__abc_52155_new_n16305_), .Y(u2__abc_52155_new_n16306_));
OR2X2 OR2X2_3506 ( .A(u2__abc_52155_new_n16310_), .B(u2__abc_52155_new_n16296_), .Y(u2__abc_52155_new_n16311_));
OR2X2 OR2X2_3507 ( .A(u2__abc_52155_new_n6960_), .B(u2__abc_52155_new_n6966_), .Y(u2__abc_52155_new_n16314_));
OR2X2 OR2X2_3508 ( .A(u2__abc_52155_new_n16317_), .B(u2__abc_52155_new_n16316_), .Y(u2__abc_52155_new_n16318_));
OR2X2 OR2X2_3509 ( .A(u2__abc_52155_new_n16318_), .B(u2__abc_52155_new_n6979_), .Y(u2__abc_52155_new_n16321_));
OR2X2 OR2X2_351 ( .A(_abc_73687_new_n1170_), .B(\a[63] ), .Y(_abc_73687_new_n1357_));
OR2X2 OR2X2_3510 ( .A(u2__abc_52155_new_n16324_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16325_));
OR2X2 OR2X2_3511 ( .A(u2__abc_52155_new_n16323_), .B(u2__abc_52155_new_n16325_), .Y(u2__abc_52155_new_n16326_));
OR2X2 OR2X2_3512 ( .A(u2__abc_52155_new_n16330_), .B(u2__abc_52155_new_n16313_), .Y(u2__abc_52155_new_n16331_));
OR2X2 OR2X2_3513 ( .A(u2__abc_52155_new_n16335_), .B(u2__abc_52155_new_n16334_), .Y(u2__abc_52155_new_n16336_));
OR2X2 OR2X2_3514 ( .A(u2__abc_52155_new_n16337_), .B(u2__abc_52155_new_n6986_), .Y(u2__abc_52155_new_n16338_));
OR2X2 OR2X2_3515 ( .A(u2__abc_52155_new_n16341_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16342_));
OR2X2 OR2X2_3516 ( .A(u2__abc_52155_new_n16340_), .B(u2__abc_52155_new_n16342_), .Y(u2__abc_52155_new_n16343_));
OR2X2 OR2X2_3517 ( .A(u2__abc_52155_new_n16347_), .B(u2__abc_52155_new_n16333_), .Y(u2__abc_52155_new_n16348_));
OR2X2 OR2X2_3518 ( .A(u2__abc_52155_new_n16352_), .B(u2__abc_52155_new_n6984_), .Y(u2__abc_52155_new_n16353_));
OR2X2 OR2X2_3519 ( .A(u2__abc_52155_new_n16351_), .B(u2__abc_52155_new_n16353_), .Y(u2__abc_52155_new_n16354_));
OR2X2 OR2X2_352 ( .A(\a[112] ), .B(\a[63] ), .Y(_abc_73687_new_n1359_));
OR2X2 OR2X2_3520 ( .A(u2__abc_52155_new_n16355_), .B(u2__abc_52155_new_n16354_), .Y(u2__abc_52155_new_n16356_));
OR2X2 OR2X2_3521 ( .A(u2__abc_52155_new_n16356_), .B(u2__abc_52155_new_n6955_), .Y(u2__abc_52155_new_n16359_));
OR2X2 OR2X2_3522 ( .A(u2__abc_52155_new_n16362_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16363_));
OR2X2 OR2X2_3523 ( .A(u2__abc_52155_new_n16361_), .B(u2__abc_52155_new_n16363_), .Y(u2__abc_52155_new_n16364_));
OR2X2 OR2X2_3524 ( .A(u2__abc_52155_new_n16368_), .B(u2__abc_52155_new_n16350_), .Y(u2__abc_52155_new_n16369_));
OR2X2 OR2X2_3525 ( .A(u2__abc_52155_new_n16376_), .B(u2__abc_52155_new_n16373_), .Y(u2__abc_52155_new_n16377_));
OR2X2 OR2X2_3526 ( .A(u2__abc_52155_new_n16379_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16380_));
OR2X2 OR2X2_3527 ( .A(u2__abc_52155_new_n16378_), .B(u2__abc_52155_new_n16380_), .Y(u2__abc_52155_new_n16381_));
OR2X2 OR2X2_3528 ( .A(u2__abc_52155_new_n16385_), .B(u2__abc_52155_new_n16371_), .Y(u2__abc_52155_new_n16386_));
OR2X2 OR2X2_3529 ( .A(u2__abc_52155_new_n16390_), .B(u2__abc_52155_new_n6943_), .Y(u2__abc_52155_new_n16391_));
OR2X2 OR2X2_353 ( .A(_abc_73687_new_n1170_), .B(\a[64] ), .Y(_abc_73687_new_n1360_));
OR2X2 OR2X2_3530 ( .A(u2__abc_52155_new_n16392_), .B(u2__abc_52155_new_n6933_), .Y(u2__abc_52155_new_n16395_));
OR2X2 OR2X2_3531 ( .A(u2__abc_52155_new_n16398_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16399_));
OR2X2 OR2X2_3532 ( .A(u2__abc_52155_new_n16397_), .B(u2__abc_52155_new_n16399_), .Y(u2__abc_52155_new_n16400_));
OR2X2 OR2X2_3533 ( .A(u2__abc_52155_new_n16404_), .B(u2__abc_52155_new_n16388_), .Y(u2__abc_52155_new_n16405_));
OR2X2 OR2X2_3534 ( .A(u2__abc_52155_new_n16409_), .B(u2__abc_52155_new_n16408_), .Y(u2__abc_52155_new_n16410_));
OR2X2 OR2X2_3535 ( .A(u2__abc_52155_new_n16411_), .B(u2__abc_52155_new_n6940_), .Y(u2__abc_52155_new_n16412_));
OR2X2 OR2X2_3536 ( .A(u2__abc_52155_new_n16415_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16416_));
OR2X2 OR2X2_3537 ( .A(u2__abc_52155_new_n16414_), .B(u2__abc_52155_new_n16416_), .Y(u2__abc_52155_new_n16417_));
OR2X2 OR2X2_3538 ( .A(u2__abc_52155_new_n16421_), .B(u2__abc_52155_new_n16407_), .Y(u2__abc_52155_new_n16422_));
OR2X2 OR2X2_3539 ( .A(u2__abc_52155_new_n16429_), .B(u2__abc_52155_new_n6938_), .Y(u2__abc_52155_new_n16430_));
OR2X2 OR2X2_354 ( .A(\a[112] ), .B(\a[64] ), .Y(_abc_73687_new_n1362_));
OR2X2 OR2X2_3540 ( .A(u2__abc_52155_new_n16389_), .B(u2__abc_52155_new_n6943_), .Y(u2__abc_52155_new_n16431_));
OR2X2 OR2X2_3541 ( .A(u2__abc_52155_new_n16433_), .B(u2__abc_52155_new_n16430_), .Y(u2__abc_52155_new_n16434_));
OR2X2 OR2X2_3542 ( .A(u2__abc_52155_new_n16428_), .B(u2__abc_52155_new_n16434_), .Y(u2__abc_52155_new_n16435_));
OR2X2 OR2X2_3543 ( .A(u2__abc_52155_new_n16427_), .B(u2__abc_52155_new_n16435_), .Y(u2__abc_52155_new_n16436_));
OR2X2 OR2X2_3544 ( .A(u2__abc_52155_new_n16436_), .B(u2__abc_52155_new_n16426_), .Y(u2__abc_52155_new_n16437_));
OR2X2 OR2X2_3545 ( .A(u2__abc_52155_new_n16425_), .B(u2__abc_52155_new_n16437_), .Y(u2__abc_52155_new_n16438_));
OR2X2 OR2X2_3546 ( .A(u2__abc_52155_new_n16438_), .B(u2__abc_52155_new_n3031_), .Y(u2__abc_52155_new_n16441_));
OR2X2 OR2X2_3547 ( .A(u2__abc_52155_new_n16444_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16445_));
OR2X2 OR2X2_3548 ( .A(u2__abc_52155_new_n16443_), .B(u2__abc_52155_new_n16445_), .Y(u2__abc_52155_new_n16446_));
OR2X2 OR2X2_3549 ( .A(u2__abc_52155_new_n16450_), .B(u2__abc_52155_new_n16424_), .Y(u2__abc_52155_new_n16451_));
OR2X2 OR2X2_355 ( .A(_abc_73687_new_n1170_), .B(\a[65] ), .Y(_abc_73687_new_n1363_));
OR2X2 OR2X2_3550 ( .A(u2__abc_52155_new_n16455_), .B(u2__abc_52155_new_n16454_), .Y(u2__abc_52155_new_n16456_));
OR2X2 OR2X2_3551 ( .A(u2__abc_52155_new_n16457_), .B(u2__abc_52155_new_n3024_), .Y(u2__abc_52155_new_n16458_));
OR2X2 OR2X2_3552 ( .A(u2__abc_52155_new_n16461_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n16462_));
OR2X2 OR2X2_3553 ( .A(u2__abc_52155_new_n16460_), .B(u2__abc_52155_new_n16462_), .Y(u2__abc_52155_new_n16463_));
OR2X2 OR2X2_3554 ( .A(u2__abc_52155_new_n16467_), .B(u2__abc_52155_new_n16453_), .Y(u2__abc_52155_new_n16468_));
OR2X2 OR2X2_3555 ( .A(u2__abc_52155_new_n16473_), .B(u2_cnt_0_), .Y(u2__abc_52155_new_n16474_));
OR2X2 OR2X2_3556 ( .A(u2__abc_52155_new_n2989_), .B(u2__abc_52155_new_n2971_), .Y(u2__abc_52155_new_n16475_));
OR2X2 OR2X2_3557 ( .A(u2__abc_52155_new_n2972_), .B(u2__abc_52155_new_n16479_), .Y(u2__abc_52155_new_n16480_));
OR2X2 OR2X2_3558 ( .A(u2__abc_52155_new_n16481_), .B(u2__abc_52155_new_n16477_), .Y(u2__0cnt_7_0__1_));
OR2X2 OR2X2_3559 ( .A(u2__abc_52155_new_n2980_), .B(u2_cnt_2_), .Y(u2__abc_52155_new_n16483_));
OR2X2 OR2X2_356 ( .A(\a[112] ), .B(\a[65] ), .Y(_abc_73687_new_n1365_));
OR2X2 OR2X2_3560 ( .A(u2__abc_52155_new_n16484_), .B(u2_cnt_2_), .Y(u2__abc_52155_new_n16487_));
OR2X2 OR2X2_3561 ( .A(u2__abc_52155_new_n16489_), .B(u2__abc_52155_new_n2983_), .Y(u2__abc_52155_new_n16490_));
OR2X2 OR2X2_3562 ( .A(u2__abc_52155_new_n16492_), .B(u2_cnt_3_), .Y(u2__abc_52155_new_n16495_));
OR2X2 OR2X2_3563 ( .A(u2__abc_52155_new_n16493_), .B(u2_cnt_4_), .Y(u2__abc_52155_new_n16502_));
OR2X2 OR2X2_3564 ( .A(u2__abc_52155_new_n16500_), .B(u2_cnt_5_), .Y(u2__abc_52155_new_n16507_));
OR2X2 OR2X2_3565 ( .A(u2__abc_52155_new_n16505_), .B(u2_cnt_6_), .Y(u2__abc_52155_new_n16510_));
OR2X2 OR2X2_3566 ( .A(u2__abc_52155_new_n16514_), .B(rst), .Y(u2__0cnt_7_0__6_));
OR2X2 OR2X2_3567 ( .A(u2__abc_52155_new_n16511_), .B(u2_cnt_7_), .Y(u2__abc_52155_new_n16518_));
OR2X2 OR2X2_3568 ( .A(u2__abc_52155_new_n16520_), .B(rst), .Y(u2__0cnt_7_0__7_));
OR2X2 OR2X2_3569 ( .A(u2__abc_52155_new_n2994_), .B(u2__abc_52155_new_n3002_), .Y(u2__abc_52155_new_n16522_));
OR2X2 OR2X2_357 ( .A(_abc_73687_new_n1170_), .B(\a[66] ), .Y(_abc_73687_new_n1366_));
OR2X2 OR2X2_3570 ( .A(u2__abc_52155_new_n16527_), .B(u2__abc_52155_new_n16529_), .Y(u2__abc_52155_new_n16530_));
OR2X2 OR2X2_3571 ( .A(u2__abc_52155_new_n16532_), .B(u2__abc_52155_new_n16534_), .Y(u2__abc_52155_new_n16535_));
OR2X2 OR2X2_3572 ( .A(u2__abc_52155_new_n16537_), .B(u2__abc_52155_new_n16539_), .Y(u2__abc_52155_new_n16540_));
OR2X2 OR2X2_3573 ( .A(u2__abc_52155_new_n16542_), .B(u2__abc_52155_new_n16544_), .Y(u2__abc_52155_new_n16545_));
OR2X2 OR2X2_3574 ( .A(u2__abc_52155_new_n16547_), .B(u2__abc_52155_new_n16549_), .Y(u2__abc_52155_new_n16550_));
OR2X2 OR2X2_3575 ( .A(u2__abc_52155_new_n16552_), .B(u2__abc_52155_new_n16554_), .Y(u2__abc_52155_new_n16555_));
OR2X2 OR2X2_3576 ( .A(u2__abc_52155_new_n16557_), .B(u2__abc_52155_new_n16559_), .Y(u2__abc_52155_new_n16560_));
OR2X2 OR2X2_3577 ( .A(u2__abc_52155_new_n16562_), .B(u2__abc_52155_new_n16564_), .Y(u2__abc_52155_new_n16565_));
OR2X2 OR2X2_3578 ( .A(u2__abc_52155_new_n16567_), .B(u2__abc_52155_new_n16569_), .Y(u2__abc_52155_new_n16570_));
OR2X2 OR2X2_3579 ( .A(u2__abc_52155_new_n16572_), .B(u2__abc_52155_new_n16574_), .Y(u2__abc_52155_new_n16575_));
OR2X2 OR2X2_358 ( .A(\a[112] ), .B(\a[66] ), .Y(_abc_73687_new_n1368_));
OR2X2 OR2X2_3580 ( .A(u2__abc_52155_new_n16577_), .B(u2__abc_52155_new_n16579_), .Y(u2__abc_52155_new_n16580_));
OR2X2 OR2X2_3581 ( .A(u2__abc_52155_new_n16582_), .B(u2__abc_52155_new_n16584_), .Y(u2__abc_52155_new_n16585_));
OR2X2 OR2X2_3582 ( .A(u2__abc_52155_new_n16587_), .B(u2__abc_52155_new_n16589_), .Y(u2__abc_52155_new_n16590_));
OR2X2 OR2X2_3583 ( .A(u2__abc_52155_new_n16592_), .B(u2__abc_52155_new_n16594_), .Y(u2__abc_52155_new_n16595_));
OR2X2 OR2X2_3584 ( .A(u2__abc_52155_new_n16597_), .B(u2__abc_52155_new_n16599_), .Y(u2__abc_52155_new_n16600_));
OR2X2 OR2X2_3585 ( .A(u2__abc_52155_new_n16602_), .B(u2__abc_52155_new_n16604_), .Y(u2__abc_52155_new_n16605_));
OR2X2 OR2X2_3586 ( .A(u2__abc_52155_new_n16607_), .B(u2__abc_52155_new_n16609_), .Y(u2__abc_52155_new_n16610_));
OR2X2 OR2X2_3587 ( .A(u2__abc_52155_new_n16612_), .B(u2__abc_52155_new_n16614_), .Y(u2__abc_52155_new_n16615_));
OR2X2 OR2X2_3588 ( .A(u2__abc_52155_new_n16617_), .B(u2__abc_52155_new_n16619_), .Y(u2__abc_52155_new_n16620_));
OR2X2 OR2X2_3589 ( .A(u2__abc_52155_new_n16622_), .B(u2__abc_52155_new_n16624_), .Y(u2__abc_52155_new_n16625_));
OR2X2 OR2X2_359 ( .A(_abc_73687_new_n1170_), .B(\a[67] ), .Y(_abc_73687_new_n1369_));
OR2X2 OR2X2_3590 ( .A(u2__abc_52155_new_n16627_), .B(u2__abc_52155_new_n16629_), .Y(u2__abc_52155_new_n16630_));
OR2X2 OR2X2_3591 ( .A(u2__abc_52155_new_n16632_), .B(u2__abc_52155_new_n16634_), .Y(u2__abc_52155_new_n16635_));
OR2X2 OR2X2_3592 ( .A(u2__abc_52155_new_n16637_), .B(u2__abc_52155_new_n16639_), .Y(u2__abc_52155_new_n16640_));
OR2X2 OR2X2_3593 ( .A(u2__abc_52155_new_n16642_), .B(u2__abc_52155_new_n16644_), .Y(u2__abc_52155_new_n16645_));
OR2X2 OR2X2_3594 ( .A(u2__abc_52155_new_n16647_), .B(u2__abc_52155_new_n16649_), .Y(u2__abc_52155_new_n16650_));
OR2X2 OR2X2_3595 ( .A(u2__abc_52155_new_n16652_), .B(u2__abc_52155_new_n16654_), .Y(u2__abc_52155_new_n16655_));
OR2X2 OR2X2_3596 ( .A(u2__abc_52155_new_n16657_), .B(u2__abc_52155_new_n16659_), .Y(u2__abc_52155_new_n16660_));
OR2X2 OR2X2_3597 ( .A(u2__abc_52155_new_n16662_), .B(u2__abc_52155_new_n16664_), .Y(u2__abc_52155_new_n16665_));
OR2X2 OR2X2_3598 ( .A(u2__abc_52155_new_n16667_), .B(u2__abc_52155_new_n16669_), .Y(u2__abc_52155_new_n16670_));
OR2X2 OR2X2_3599 ( .A(u2__abc_52155_new_n16672_), .B(u2__abc_52155_new_n16674_), .Y(u2__abc_52155_new_n16675_));
OR2X2 OR2X2_36 ( .A(_abc_73687_new_n753_), .B(\a[17] ), .Y(_abc_73687_new_n882_));
OR2X2 OR2X2_360 ( .A(\a[112] ), .B(\a[67] ), .Y(_abc_73687_new_n1371_));
OR2X2 OR2X2_3600 ( .A(u2__abc_52155_new_n2994_), .B(u2__abc_52155_new_n2985_), .Y(u2__abc_52155_new_n16678_));
OR2X2 OR2X2_3601 ( .A(u2__abc_52155_new_n16679_), .B(u2__abc_52155_new_n16677_), .Y(u2__abc_52155_new_n16680_));
OR2X2 OR2X2_3602 ( .A(u2__abc_52155_new_n16684_), .B(u2__abc_52155_new_n16682_), .Y(u2__abc_52155_new_n16685_));
OR2X2 OR2X2_3603 ( .A(u2__abc_52155_new_n16681_), .B(u2__abc_52155_new_n16686_), .Y(u2__0remLo_451_0__32_));
OR2X2 OR2X2_3604 ( .A(u2__abc_52155_new_n16689_), .B(u2__abc_52155_new_n16690_), .Y(u2__abc_52155_new_n16691_));
OR2X2 OR2X2_3605 ( .A(u2__abc_52155_new_n16688_), .B(u2__abc_52155_new_n16692_), .Y(u2__0remLo_451_0__33_));
OR2X2 OR2X2_3606 ( .A(u2__abc_52155_new_n16694_), .B(u2__abc_52155_new_n16695_), .Y(u2__abc_52155_new_n16696_));
OR2X2 OR2X2_3607 ( .A(u2__abc_52155_new_n16698_), .B(u2__abc_52155_new_n16699_), .Y(u2__abc_52155_new_n16700_));
OR2X2 OR2X2_3608 ( .A(u2__abc_52155_new_n16697_), .B(u2__abc_52155_new_n16701_), .Y(u2__0remLo_451_0__34_));
OR2X2 OR2X2_3609 ( .A(u2__abc_52155_new_n16704_), .B(u2__abc_52155_new_n16705_), .Y(u2__abc_52155_new_n16706_));
OR2X2 OR2X2_361 ( .A(_abc_73687_new_n1170_), .B(\a[68] ), .Y(_abc_73687_new_n1372_));
OR2X2 OR2X2_3610 ( .A(u2__abc_52155_new_n16703_), .B(u2__abc_52155_new_n16707_), .Y(u2__0remLo_451_0__35_));
OR2X2 OR2X2_3611 ( .A(u2__abc_52155_new_n16710_), .B(u2__abc_52155_new_n16711_), .Y(u2__abc_52155_new_n16712_));
OR2X2 OR2X2_3612 ( .A(u2__abc_52155_new_n16709_), .B(u2__abc_52155_new_n16713_), .Y(u2__0remLo_451_0__36_));
OR2X2 OR2X2_3613 ( .A(u2__abc_52155_new_n16716_), .B(u2__abc_52155_new_n16717_), .Y(u2__abc_52155_new_n16718_));
OR2X2 OR2X2_3614 ( .A(u2__abc_52155_new_n16715_), .B(u2__abc_52155_new_n16719_), .Y(u2__0remLo_451_0__37_));
OR2X2 OR2X2_3615 ( .A(u2__abc_52155_new_n16723_), .B(u2__abc_52155_new_n16722_), .Y(u2__abc_52155_new_n16724_));
OR2X2 OR2X2_3616 ( .A(u2__abc_52155_new_n16721_), .B(u2__abc_52155_new_n16725_), .Y(u2__0remLo_451_0__38_));
OR2X2 OR2X2_3617 ( .A(u2__abc_52155_new_n16728_), .B(u2__abc_52155_new_n16729_), .Y(u2__abc_52155_new_n16730_));
OR2X2 OR2X2_3618 ( .A(u2__abc_52155_new_n16727_), .B(u2__abc_52155_new_n16731_), .Y(u2__0remLo_451_0__39_));
OR2X2 OR2X2_3619 ( .A(u2__abc_52155_new_n16734_), .B(u2__abc_52155_new_n16735_), .Y(u2__abc_52155_new_n16736_));
OR2X2 OR2X2_362 ( .A(\a[112] ), .B(\a[68] ), .Y(_abc_73687_new_n1374_));
OR2X2 OR2X2_3620 ( .A(u2__abc_52155_new_n16733_), .B(u2__abc_52155_new_n16737_), .Y(u2__0remLo_451_0__40_));
OR2X2 OR2X2_3621 ( .A(u2__abc_52155_new_n16740_), .B(u2__abc_52155_new_n16741_), .Y(u2__abc_52155_new_n16742_));
OR2X2 OR2X2_3622 ( .A(u2__abc_52155_new_n16739_), .B(u2__abc_52155_new_n16743_), .Y(u2__0remLo_451_0__41_));
OR2X2 OR2X2_3623 ( .A(u2__abc_52155_new_n16747_), .B(u2__abc_52155_new_n16746_), .Y(u2__abc_52155_new_n16748_));
OR2X2 OR2X2_3624 ( .A(u2__abc_52155_new_n16745_), .B(u2__abc_52155_new_n16749_), .Y(u2__0remLo_451_0__42_));
OR2X2 OR2X2_3625 ( .A(u2__abc_52155_new_n16752_), .B(u2__abc_52155_new_n16753_), .Y(u2__abc_52155_new_n16754_));
OR2X2 OR2X2_3626 ( .A(u2__abc_52155_new_n16751_), .B(u2__abc_52155_new_n16755_), .Y(u2__0remLo_451_0__43_));
OR2X2 OR2X2_3627 ( .A(u2__abc_52155_new_n16758_), .B(u2__abc_52155_new_n16759_), .Y(u2__abc_52155_new_n16760_));
OR2X2 OR2X2_3628 ( .A(u2__abc_52155_new_n16757_), .B(u2__abc_52155_new_n16761_), .Y(u2__0remLo_451_0__44_));
OR2X2 OR2X2_3629 ( .A(u2__abc_52155_new_n16764_), .B(u2__abc_52155_new_n16765_), .Y(u2__abc_52155_new_n16766_));
OR2X2 OR2X2_363 ( .A(_abc_73687_new_n1170_), .B(\a[69] ), .Y(_abc_73687_new_n1375_));
OR2X2 OR2X2_3630 ( .A(u2__abc_52155_new_n16763_), .B(u2__abc_52155_new_n16767_), .Y(u2__0remLo_451_0__45_));
OR2X2 OR2X2_3631 ( .A(u2__abc_52155_new_n16769_), .B(u2__abc_52155_new_n16770_), .Y(u2__abc_52155_new_n16771_));
OR2X2 OR2X2_3632 ( .A(u2__abc_52155_new_n16773_), .B(u2__abc_52155_new_n16774_), .Y(u2__abc_52155_new_n16775_));
OR2X2 OR2X2_3633 ( .A(u2__abc_52155_new_n16772_), .B(u2__abc_52155_new_n16776_), .Y(u2__0remLo_451_0__46_));
OR2X2 OR2X2_3634 ( .A(u2__abc_52155_new_n16780_), .B(u2__abc_52155_new_n16779_), .Y(u2__abc_52155_new_n16781_));
OR2X2 OR2X2_3635 ( .A(u2__abc_52155_new_n16778_), .B(u2__abc_52155_new_n16782_), .Y(u2__0remLo_451_0__47_));
OR2X2 OR2X2_3636 ( .A(u2__abc_52155_new_n16785_), .B(u2__abc_52155_new_n16786_), .Y(u2__abc_52155_new_n16787_));
OR2X2 OR2X2_3637 ( .A(u2__abc_52155_new_n16784_), .B(u2__abc_52155_new_n16788_), .Y(u2__0remLo_451_0__48_));
OR2X2 OR2X2_3638 ( .A(u2__abc_52155_new_n16791_), .B(u2__abc_52155_new_n16792_), .Y(u2__abc_52155_new_n16793_));
OR2X2 OR2X2_3639 ( .A(u2__abc_52155_new_n16790_), .B(u2__abc_52155_new_n16794_), .Y(u2__0remLo_451_0__49_));
OR2X2 OR2X2_364 ( .A(\a[112] ), .B(\a[69] ), .Y(_abc_73687_new_n1377_));
OR2X2 OR2X2_3640 ( .A(u2__abc_52155_new_n16797_), .B(u2__abc_52155_new_n16798_), .Y(u2__abc_52155_new_n16799_));
OR2X2 OR2X2_3641 ( .A(u2__abc_52155_new_n16796_), .B(u2__abc_52155_new_n16800_), .Y(u2__0remLo_451_0__50_));
OR2X2 OR2X2_3642 ( .A(u2__abc_52155_new_n16804_), .B(u2__abc_52155_new_n16803_), .Y(u2__abc_52155_new_n16805_));
OR2X2 OR2X2_3643 ( .A(u2__abc_52155_new_n16802_), .B(u2__abc_52155_new_n16806_), .Y(u2__0remLo_451_0__51_));
OR2X2 OR2X2_3644 ( .A(u2__abc_52155_new_n16809_), .B(u2__abc_52155_new_n16810_), .Y(u2__abc_52155_new_n16811_));
OR2X2 OR2X2_3645 ( .A(u2__abc_52155_new_n16808_), .B(u2__abc_52155_new_n16812_), .Y(u2__0remLo_451_0__52_));
OR2X2 OR2X2_3646 ( .A(u2__abc_52155_new_n16815_), .B(u2__abc_52155_new_n16816_), .Y(u2__abc_52155_new_n16817_));
OR2X2 OR2X2_3647 ( .A(u2__abc_52155_new_n16814_), .B(u2__abc_52155_new_n16818_), .Y(u2__0remLo_451_0__53_));
OR2X2 OR2X2_3648 ( .A(u2__abc_52155_new_n16821_), .B(u2__abc_52155_new_n16822_), .Y(u2__abc_52155_new_n16823_));
OR2X2 OR2X2_3649 ( .A(u2__abc_52155_new_n16820_), .B(u2__abc_52155_new_n16824_), .Y(u2__0remLo_451_0__54_));
OR2X2 OR2X2_365 ( .A(_abc_73687_new_n1170_), .B(\a[70] ), .Y(_abc_73687_new_n1378_));
OR2X2 OR2X2_3650 ( .A(u2__abc_52155_new_n16827_), .B(u2__abc_52155_new_n16828_), .Y(u2__abc_52155_new_n16829_));
OR2X2 OR2X2_3651 ( .A(u2__abc_52155_new_n16826_), .B(u2__abc_52155_new_n16830_), .Y(u2__0remLo_451_0__55_));
OR2X2 OR2X2_3652 ( .A(u2__abc_52155_new_n16833_), .B(u2__abc_52155_new_n16834_), .Y(u2__abc_52155_new_n16835_));
OR2X2 OR2X2_3653 ( .A(u2__abc_52155_new_n16832_), .B(u2__abc_52155_new_n16836_), .Y(u2__0remLo_451_0__56_));
OR2X2 OR2X2_3654 ( .A(u2__abc_52155_new_n16840_), .B(u2__abc_52155_new_n16839_), .Y(u2__abc_52155_new_n16841_));
OR2X2 OR2X2_3655 ( .A(u2__abc_52155_new_n16838_), .B(u2__abc_52155_new_n16842_), .Y(u2__0remLo_451_0__57_));
OR2X2 OR2X2_3656 ( .A(u2__abc_52155_new_n16846_), .B(u2__abc_52155_new_n16845_), .Y(u2__abc_52155_new_n16847_));
OR2X2 OR2X2_3657 ( .A(u2__abc_52155_new_n16844_), .B(u2__abc_52155_new_n16848_), .Y(u2__0remLo_451_0__58_));
OR2X2 OR2X2_3658 ( .A(u2__abc_52155_new_n16851_), .B(u2__abc_52155_new_n16852_), .Y(u2__abc_52155_new_n16853_));
OR2X2 OR2X2_3659 ( .A(u2__abc_52155_new_n16850_), .B(u2__abc_52155_new_n16854_), .Y(u2__0remLo_451_0__59_));
OR2X2 OR2X2_366 ( .A(\a[112] ), .B(\a[70] ), .Y(_abc_73687_new_n1380_));
OR2X2 OR2X2_3660 ( .A(u2__abc_52155_new_n16857_), .B(u2__abc_52155_new_n16858_), .Y(u2__abc_52155_new_n16859_));
OR2X2 OR2X2_3661 ( .A(u2__abc_52155_new_n16856_), .B(u2__abc_52155_new_n16860_), .Y(u2__0remLo_451_0__60_));
OR2X2 OR2X2_3662 ( .A(u2__abc_52155_new_n16862_), .B(u2__abc_52155_new_n16863_), .Y(u2__abc_52155_new_n16864_));
OR2X2 OR2X2_3663 ( .A(u2__abc_52155_new_n16866_), .B(u2__abc_52155_new_n16867_), .Y(u2__abc_52155_new_n16868_));
OR2X2 OR2X2_3664 ( .A(u2__abc_52155_new_n16865_), .B(u2__abc_52155_new_n16869_), .Y(u2__0remLo_451_0__61_));
OR2X2 OR2X2_3665 ( .A(u2__abc_52155_new_n16872_), .B(u2__abc_52155_new_n16873_), .Y(u2__abc_52155_new_n16874_));
OR2X2 OR2X2_3666 ( .A(u2__abc_52155_new_n16871_), .B(u2__abc_52155_new_n16875_), .Y(u2__0remLo_451_0__62_));
OR2X2 OR2X2_3667 ( .A(u2__abc_52155_new_n16879_), .B(u2__abc_52155_new_n16878_), .Y(u2__abc_52155_new_n16880_));
OR2X2 OR2X2_3668 ( .A(u2__abc_52155_new_n16877_), .B(u2__abc_52155_new_n16881_), .Y(u2__0remLo_451_0__63_));
OR2X2 OR2X2_3669 ( .A(u2__abc_52155_new_n16885_), .B(u2__abc_52155_new_n16884_), .Y(u2__abc_52155_new_n16886_));
OR2X2 OR2X2_367 ( .A(_abc_73687_new_n1170_), .B(\a[71] ), .Y(_abc_73687_new_n1381_));
OR2X2 OR2X2_3670 ( .A(u2__abc_52155_new_n16883_), .B(u2__abc_52155_new_n16887_), .Y(u2__0remLo_451_0__64_));
OR2X2 OR2X2_3671 ( .A(u2__abc_52155_new_n16889_), .B(u2__abc_52155_new_n16890_), .Y(u2__abc_52155_new_n16891_));
OR2X2 OR2X2_3672 ( .A(u2__abc_52155_new_n16893_), .B(u2__abc_52155_new_n16894_), .Y(u2__abc_52155_new_n16895_));
OR2X2 OR2X2_3673 ( .A(u2__abc_52155_new_n16892_), .B(u2__abc_52155_new_n16896_), .Y(u2__0remLo_451_0__65_));
OR2X2 OR2X2_3674 ( .A(u2__abc_52155_new_n16900_), .B(u2__abc_52155_new_n16899_), .Y(u2__abc_52155_new_n16901_));
OR2X2 OR2X2_3675 ( .A(u2__abc_52155_new_n16898_), .B(u2__abc_52155_new_n16902_), .Y(u2__0remLo_451_0__66_));
OR2X2 OR2X2_3676 ( .A(u2__abc_52155_new_n16905_), .B(u2__abc_52155_new_n16906_), .Y(u2__abc_52155_new_n16907_));
OR2X2 OR2X2_3677 ( .A(u2__abc_52155_new_n16904_), .B(u2__abc_52155_new_n16908_), .Y(u2__0remLo_451_0__67_));
OR2X2 OR2X2_3678 ( .A(u2__abc_52155_new_n16911_), .B(u2__abc_52155_new_n16912_), .Y(u2__abc_52155_new_n16913_));
OR2X2 OR2X2_3679 ( .A(u2__abc_52155_new_n16910_), .B(u2__abc_52155_new_n16914_), .Y(u2__0remLo_451_0__68_));
OR2X2 OR2X2_368 ( .A(\a[112] ), .B(\a[71] ), .Y(_abc_73687_new_n1383_));
OR2X2 OR2X2_3680 ( .A(u2__abc_52155_new_n16917_), .B(u2__abc_52155_new_n16918_), .Y(u2__abc_52155_new_n16919_));
OR2X2 OR2X2_3681 ( .A(u2__abc_52155_new_n16916_), .B(u2__abc_52155_new_n16920_), .Y(u2__0remLo_451_0__69_));
OR2X2 OR2X2_3682 ( .A(u2__abc_52155_new_n16924_), .B(u2__abc_52155_new_n16923_), .Y(u2__abc_52155_new_n16925_));
OR2X2 OR2X2_3683 ( .A(u2__abc_52155_new_n16922_), .B(u2__abc_52155_new_n16926_), .Y(u2__0remLo_451_0__70_));
OR2X2 OR2X2_3684 ( .A(u2__abc_52155_new_n16929_), .B(u2__abc_52155_new_n16930_), .Y(u2__abc_52155_new_n16931_));
OR2X2 OR2X2_3685 ( .A(u2__abc_52155_new_n16928_), .B(u2__abc_52155_new_n16932_), .Y(u2__0remLo_451_0__71_));
OR2X2 OR2X2_3686 ( .A(u2__abc_52155_new_n16935_), .B(u2__abc_52155_new_n16936_), .Y(u2__abc_52155_new_n16937_));
OR2X2 OR2X2_3687 ( .A(u2__abc_52155_new_n16934_), .B(u2__abc_52155_new_n16938_), .Y(u2__0remLo_451_0__72_));
OR2X2 OR2X2_3688 ( .A(u2__abc_52155_new_n16941_), .B(u2__abc_52155_new_n16942_), .Y(u2__abc_52155_new_n16943_));
OR2X2 OR2X2_3689 ( .A(u2__abc_52155_new_n16940_), .B(u2__abc_52155_new_n16944_), .Y(u2__0remLo_451_0__73_));
OR2X2 OR2X2_369 ( .A(_abc_73687_new_n1170_), .B(\a[72] ), .Y(_abc_73687_new_n1384_));
OR2X2 OR2X2_3690 ( .A(u2__abc_52155_new_n16946_), .B(u2__abc_52155_new_n16947_), .Y(u2__abc_52155_new_n16948_));
OR2X2 OR2X2_3691 ( .A(u2__abc_52155_new_n16950_), .B(u2__abc_52155_new_n16951_), .Y(u2__abc_52155_new_n16952_));
OR2X2 OR2X2_3692 ( .A(u2__abc_52155_new_n16949_), .B(u2__abc_52155_new_n16953_), .Y(u2__0remLo_451_0__74_));
OR2X2 OR2X2_3693 ( .A(u2__abc_52155_new_n16956_), .B(u2__abc_52155_new_n16957_), .Y(u2__abc_52155_new_n16958_));
OR2X2 OR2X2_3694 ( .A(u2__abc_52155_new_n16955_), .B(u2__abc_52155_new_n16959_), .Y(u2__0remLo_451_0__75_));
OR2X2 OR2X2_3695 ( .A(u2__abc_52155_new_n16962_), .B(u2__abc_52155_new_n16963_), .Y(u2__abc_52155_new_n16964_));
OR2X2 OR2X2_3696 ( .A(u2__abc_52155_new_n16961_), .B(u2__abc_52155_new_n16965_), .Y(u2__0remLo_451_0__76_));
OR2X2 OR2X2_3697 ( .A(u2__abc_52155_new_n16968_), .B(u2__abc_52155_new_n16969_), .Y(u2__abc_52155_new_n16970_));
OR2X2 OR2X2_3698 ( .A(u2__abc_52155_new_n16967_), .B(u2__abc_52155_new_n16971_), .Y(u2__0remLo_451_0__77_));
OR2X2 OR2X2_3699 ( .A(u2__abc_52155_new_n16974_), .B(u2__abc_52155_new_n16975_), .Y(u2__abc_52155_new_n16976_));
OR2X2 OR2X2_37 ( .A(aNan), .B(sqrto_94_), .Y(_abc_73687_new_n884_));
OR2X2 OR2X2_370 ( .A(\a[112] ), .B(\a[72] ), .Y(_abc_73687_new_n1386_));
OR2X2 OR2X2_3700 ( .A(u2__abc_52155_new_n16973_), .B(u2__abc_52155_new_n16977_), .Y(u2__0remLo_451_0__78_));
OR2X2 OR2X2_3701 ( .A(u2__abc_52155_new_n16981_), .B(u2__abc_52155_new_n16980_), .Y(u2__abc_52155_new_n16982_));
OR2X2 OR2X2_3702 ( .A(u2__abc_52155_new_n16979_), .B(u2__abc_52155_new_n16983_), .Y(u2__0remLo_451_0__79_));
OR2X2 OR2X2_3703 ( .A(u2__abc_52155_new_n16985_), .B(u2__abc_52155_new_n16986_), .Y(u2__abc_52155_new_n16987_));
OR2X2 OR2X2_3704 ( .A(u2__abc_52155_new_n16989_), .B(u2__abc_52155_new_n16990_), .Y(u2__abc_52155_new_n16991_));
OR2X2 OR2X2_3705 ( .A(u2__abc_52155_new_n16988_), .B(u2__abc_52155_new_n16992_), .Y(u2__0remLo_451_0__80_));
OR2X2 OR2X2_3706 ( .A(u2__abc_52155_new_n16995_), .B(u2__abc_52155_new_n16996_), .Y(u2__abc_52155_new_n16997_));
OR2X2 OR2X2_3707 ( .A(u2__abc_52155_new_n16994_), .B(u2__abc_52155_new_n16998_), .Y(u2__0remLo_451_0__81_));
OR2X2 OR2X2_3708 ( .A(u2__abc_52155_new_n17001_), .B(u2__abc_52155_new_n17002_), .Y(u2__abc_52155_new_n17003_));
OR2X2 OR2X2_3709 ( .A(u2__abc_52155_new_n17000_), .B(u2__abc_52155_new_n17004_), .Y(u2__0remLo_451_0__82_));
OR2X2 OR2X2_371 ( .A(_abc_73687_new_n1170_), .B(\a[73] ), .Y(_abc_73687_new_n1387_));
OR2X2 OR2X2_3710 ( .A(u2__abc_52155_new_n17008_), .B(u2__abc_52155_new_n17007_), .Y(u2__abc_52155_new_n17009_));
OR2X2 OR2X2_3711 ( .A(u2__abc_52155_new_n17006_), .B(u2__abc_52155_new_n17010_), .Y(u2__0remLo_451_0__83_));
OR2X2 OR2X2_3712 ( .A(u2__abc_52155_new_n17013_), .B(u2__abc_52155_new_n17014_), .Y(u2__abc_52155_new_n17015_));
OR2X2 OR2X2_3713 ( .A(u2__abc_52155_new_n17012_), .B(u2__abc_52155_new_n17016_), .Y(u2__0remLo_451_0__84_));
OR2X2 OR2X2_3714 ( .A(u2__abc_52155_new_n17019_), .B(u2__abc_52155_new_n17020_), .Y(u2__abc_52155_new_n17021_));
OR2X2 OR2X2_3715 ( .A(u2__abc_52155_new_n17018_), .B(u2__abc_52155_new_n17022_), .Y(u2__0remLo_451_0__85_));
OR2X2 OR2X2_3716 ( .A(u2__abc_52155_new_n17025_), .B(u2__abc_52155_new_n17026_), .Y(u2__abc_52155_new_n17027_));
OR2X2 OR2X2_3717 ( .A(u2__abc_52155_new_n17024_), .B(u2__abc_52155_new_n17028_), .Y(u2__0remLo_451_0__86_));
OR2X2 OR2X2_3718 ( .A(u2__abc_52155_new_n17031_), .B(u2__abc_52155_new_n17032_), .Y(u2__abc_52155_new_n17033_));
OR2X2 OR2X2_3719 ( .A(u2__abc_52155_new_n17030_), .B(u2__abc_52155_new_n17034_), .Y(u2__0remLo_451_0__87_));
OR2X2 OR2X2_372 ( .A(\a[112] ), .B(\a[73] ), .Y(_abc_73687_new_n1389_));
OR2X2 OR2X2_3720 ( .A(u2__abc_52155_new_n17037_), .B(u2__abc_52155_new_n17038_), .Y(u2__abc_52155_new_n17039_));
OR2X2 OR2X2_3721 ( .A(u2__abc_52155_new_n17036_), .B(u2__abc_52155_new_n17040_), .Y(u2__0remLo_451_0__88_));
OR2X2 OR2X2_3722 ( .A(u2__abc_52155_new_n17044_), .B(u2__abc_52155_new_n17043_), .Y(u2__abc_52155_new_n17045_));
OR2X2 OR2X2_3723 ( .A(u2__abc_52155_new_n17042_), .B(u2__abc_52155_new_n17046_), .Y(u2__0remLo_451_0__89_));
OR2X2 OR2X2_3724 ( .A(u2__abc_52155_new_n17049_), .B(u2__abc_52155_new_n17050_), .Y(u2__abc_52155_new_n17051_));
OR2X2 OR2X2_3725 ( .A(u2__abc_52155_new_n17048_), .B(u2__abc_52155_new_n17052_), .Y(u2__0remLo_451_0__90_));
OR2X2 OR2X2_3726 ( .A(u2__abc_52155_new_n17055_), .B(u2__abc_52155_new_n17056_), .Y(u2__abc_52155_new_n17057_));
OR2X2 OR2X2_3727 ( .A(u2__abc_52155_new_n17054_), .B(u2__abc_52155_new_n17058_), .Y(u2__0remLo_451_0__91_));
OR2X2 OR2X2_3728 ( .A(u2__abc_52155_new_n17061_), .B(u2__abc_52155_new_n17062_), .Y(u2__abc_52155_new_n17063_));
OR2X2 OR2X2_3729 ( .A(u2__abc_52155_new_n17060_), .B(u2__abc_52155_new_n17064_), .Y(u2__0remLo_451_0__92_));
OR2X2 OR2X2_373 ( .A(_abc_73687_new_n1170_), .B(\a[74] ), .Y(_abc_73687_new_n1390_));
OR2X2 OR2X2_3730 ( .A(u2__abc_52155_new_n17068_), .B(u2__abc_52155_new_n17067_), .Y(u2__abc_52155_new_n17069_));
OR2X2 OR2X2_3731 ( .A(u2__abc_52155_new_n17066_), .B(u2__abc_52155_new_n17070_), .Y(u2__0remLo_451_0__93_));
OR2X2 OR2X2_3732 ( .A(u2__abc_52155_new_n17073_), .B(u2__abc_52155_new_n17074_), .Y(u2__abc_52155_new_n17075_));
OR2X2 OR2X2_3733 ( .A(u2__abc_52155_new_n17072_), .B(u2__abc_52155_new_n17076_), .Y(u2__0remLo_451_0__94_));
OR2X2 OR2X2_3734 ( .A(u2__abc_52155_new_n17080_), .B(u2__abc_52155_new_n17079_), .Y(u2__abc_52155_new_n17081_));
OR2X2 OR2X2_3735 ( .A(u2__abc_52155_new_n17078_), .B(u2__abc_52155_new_n17082_), .Y(u2__0remLo_451_0__95_));
OR2X2 OR2X2_3736 ( .A(u2__abc_52155_new_n17088_), .B(u2__abc_52155_new_n17086_), .Y(u2__abc_52155_new_n17089_));
OR2X2 OR2X2_3737 ( .A(u2__abc_52155_new_n17084_), .B(u2__abc_52155_new_n17089_), .Y(u2__0remLo_451_0__96_));
OR2X2 OR2X2_3738 ( .A(u2__abc_52155_new_n17091_), .B(u2__abc_52155_new_n17092_), .Y(u2__abc_52155_new_n17093_));
OR2X2 OR2X2_3739 ( .A(u2__abc_52155_new_n17095_), .B(u2__abc_52155_new_n17096_), .Y(u2__abc_52155_new_n17097_));
OR2X2 OR2X2_374 ( .A(\a[112] ), .B(\a[74] ), .Y(_abc_73687_new_n1392_));
OR2X2 OR2X2_3740 ( .A(u2__abc_52155_new_n17094_), .B(u2__abc_52155_new_n17098_), .Y(u2__0remLo_451_0__97_));
OR2X2 OR2X2_3741 ( .A(u2__abc_52155_new_n17103_), .B(u2__abc_52155_new_n17101_), .Y(u2__abc_52155_new_n17104_));
OR2X2 OR2X2_3742 ( .A(u2__abc_52155_new_n17100_), .B(u2__abc_52155_new_n17104_), .Y(u2__0remLo_451_0__98_));
OR2X2 OR2X2_3743 ( .A(u2__abc_52155_new_n17107_), .B(u2__abc_52155_new_n17108_), .Y(u2__abc_52155_new_n17109_));
OR2X2 OR2X2_3744 ( .A(u2__abc_52155_new_n17106_), .B(u2__abc_52155_new_n17110_), .Y(u2__0remLo_451_0__99_));
OR2X2 OR2X2_3745 ( .A(u2__abc_52155_new_n17113_), .B(u2__abc_52155_new_n17114_), .Y(u2__abc_52155_new_n17115_));
OR2X2 OR2X2_3746 ( .A(u2__abc_52155_new_n17112_), .B(u2__abc_52155_new_n17116_), .Y(u2__0remLo_451_0__100_));
OR2X2 OR2X2_3747 ( .A(u2__abc_52155_new_n17119_), .B(u2__abc_52155_new_n17120_), .Y(u2__abc_52155_new_n17121_));
OR2X2 OR2X2_3748 ( .A(u2__abc_52155_new_n17118_), .B(u2__abc_52155_new_n17122_), .Y(u2__0remLo_451_0__101_));
OR2X2 OR2X2_3749 ( .A(u2__abc_52155_new_n17126_), .B(u2__abc_52155_new_n17125_), .Y(u2__abc_52155_new_n17127_));
OR2X2 OR2X2_375 ( .A(_abc_73687_new_n1170_), .B(\a[75] ), .Y(_abc_73687_new_n1393_));
OR2X2 OR2X2_3750 ( .A(u2__abc_52155_new_n17124_), .B(u2__abc_52155_new_n17128_), .Y(u2__0remLo_451_0__102_));
OR2X2 OR2X2_3751 ( .A(u2__abc_52155_new_n17131_), .B(u2__abc_52155_new_n17132_), .Y(u2__abc_52155_new_n17133_));
OR2X2 OR2X2_3752 ( .A(u2__abc_52155_new_n17130_), .B(u2__abc_52155_new_n17134_), .Y(u2__0remLo_451_0__103_));
OR2X2 OR2X2_3753 ( .A(u2__abc_52155_new_n17137_), .B(u2__abc_52155_new_n17138_), .Y(u2__abc_52155_new_n17139_));
OR2X2 OR2X2_3754 ( .A(u2__abc_52155_new_n17136_), .B(u2__abc_52155_new_n17140_), .Y(u2__0remLo_451_0__104_));
OR2X2 OR2X2_3755 ( .A(u2__abc_52155_new_n17143_), .B(u2__abc_52155_new_n17144_), .Y(u2__abc_52155_new_n17145_));
OR2X2 OR2X2_3756 ( .A(u2__abc_52155_new_n17142_), .B(u2__abc_52155_new_n17146_), .Y(u2__0remLo_451_0__105_));
OR2X2 OR2X2_3757 ( .A(u2__abc_52155_new_n17150_), .B(u2__abc_52155_new_n17149_), .Y(u2__abc_52155_new_n17151_));
OR2X2 OR2X2_3758 ( .A(u2__abc_52155_new_n17148_), .B(u2__abc_52155_new_n17152_), .Y(u2__0remLo_451_0__106_));
OR2X2 OR2X2_3759 ( .A(u2__abc_52155_new_n17155_), .B(u2__abc_52155_new_n17156_), .Y(u2__abc_52155_new_n17157_));
OR2X2 OR2X2_376 ( .A(\a[112] ), .B(\a[75] ), .Y(_abc_73687_new_n1395_));
OR2X2 OR2X2_3760 ( .A(u2__abc_52155_new_n17154_), .B(u2__abc_52155_new_n17158_), .Y(u2__0remLo_451_0__107_));
OR2X2 OR2X2_3761 ( .A(u2__abc_52155_new_n17161_), .B(u2__abc_52155_new_n17162_), .Y(u2__abc_52155_new_n17163_));
OR2X2 OR2X2_3762 ( .A(u2__abc_52155_new_n17160_), .B(u2__abc_52155_new_n17164_), .Y(u2__0remLo_451_0__108_));
OR2X2 OR2X2_3763 ( .A(u2__abc_52155_new_n17167_), .B(u2__abc_52155_new_n17168_), .Y(u2__abc_52155_new_n17169_));
OR2X2 OR2X2_3764 ( .A(u2__abc_52155_new_n17166_), .B(u2__abc_52155_new_n17170_), .Y(u2__0remLo_451_0__109_));
OR2X2 OR2X2_3765 ( .A(u2__abc_52155_new_n17172_), .B(u2__abc_52155_new_n17173_), .Y(u2__abc_52155_new_n17174_));
OR2X2 OR2X2_3766 ( .A(u2__abc_52155_new_n17176_), .B(u2__abc_52155_new_n17177_), .Y(u2__abc_52155_new_n17178_));
OR2X2 OR2X2_3767 ( .A(u2__abc_52155_new_n17175_), .B(u2__abc_52155_new_n17179_), .Y(u2__0remLo_451_0__110_));
OR2X2 OR2X2_3768 ( .A(u2__abc_52155_new_n17182_), .B(u2__abc_52155_new_n17183_), .Y(u2__abc_52155_new_n17184_));
OR2X2 OR2X2_3769 ( .A(u2__abc_52155_new_n17181_), .B(u2__abc_52155_new_n17185_), .Y(u2__0remLo_451_0__111_));
OR2X2 OR2X2_377 ( .A(_abc_73687_new_n1170_), .B(\a[76] ), .Y(_abc_73687_new_n1396_));
OR2X2 OR2X2_3770 ( .A(u2__abc_52155_new_n17188_), .B(u2__abc_52155_new_n17189_), .Y(u2__abc_52155_new_n17190_));
OR2X2 OR2X2_3771 ( .A(u2__abc_52155_new_n17187_), .B(u2__abc_52155_new_n17191_), .Y(u2__0remLo_451_0__112_));
OR2X2 OR2X2_3772 ( .A(u2__abc_52155_new_n17194_), .B(u2__abc_52155_new_n17195_), .Y(u2__abc_52155_new_n17196_));
OR2X2 OR2X2_3773 ( .A(u2__abc_52155_new_n17193_), .B(u2__abc_52155_new_n17197_), .Y(u2__0remLo_451_0__113_));
OR2X2 OR2X2_3774 ( .A(u2__abc_52155_new_n17199_), .B(u2__abc_52155_new_n17200_), .Y(u2__abc_52155_new_n17201_));
OR2X2 OR2X2_3775 ( .A(u2__abc_52155_new_n17203_), .B(u2__abc_52155_new_n17204_), .Y(u2__abc_52155_new_n17205_));
OR2X2 OR2X2_3776 ( .A(u2__abc_52155_new_n17202_), .B(u2__abc_52155_new_n17206_), .Y(u2__0remLo_451_0__114_));
OR2X2 OR2X2_3777 ( .A(u2__abc_52155_new_n17210_), .B(u2__abc_52155_new_n17209_), .Y(u2__abc_52155_new_n17211_));
OR2X2 OR2X2_3778 ( .A(u2__abc_52155_new_n17208_), .B(u2__abc_52155_new_n17212_), .Y(u2__0remLo_451_0__115_));
OR2X2 OR2X2_3779 ( .A(u2__abc_52155_new_n17215_), .B(u2__abc_52155_new_n17216_), .Y(u2__abc_52155_new_n17217_));
OR2X2 OR2X2_378 ( .A(\a[112] ), .B(\a[76] ), .Y(_abc_73687_new_n1398_));
OR2X2 OR2X2_3780 ( .A(u2__abc_52155_new_n17214_), .B(u2__abc_52155_new_n17218_), .Y(u2__0remLo_451_0__116_));
OR2X2 OR2X2_3781 ( .A(u2__abc_52155_new_n17221_), .B(u2__abc_52155_new_n17222_), .Y(u2__abc_52155_new_n17223_));
OR2X2 OR2X2_3782 ( .A(u2__abc_52155_new_n17220_), .B(u2__abc_52155_new_n17224_), .Y(u2__0remLo_451_0__117_));
OR2X2 OR2X2_3783 ( .A(u2__abc_52155_new_n17227_), .B(u2__abc_52155_new_n17228_), .Y(u2__abc_52155_new_n17229_));
OR2X2 OR2X2_3784 ( .A(u2__abc_52155_new_n17226_), .B(u2__abc_52155_new_n17230_), .Y(u2__0remLo_451_0__118_));
OR2X2 OR2X2_3785 ( .A(u2__abc_52155_new_n17233_), .B(u2__abc_52155_new_n17234_), .Y(u2__abc_52155_new_n17235_));
OR2X2 OR2X2_3786 ( .A(u2__abc_52155_new_n17232_), .B(u2__abc_52155_new_n17236_), .Y(u2__0remLo_451_0__119_));
OR2X2 OR2X2_3787 ( .A(u2__abc_52155_new_n17239_), .B(u2__abc_52155_new_n17240_), .Y(u2__abc_52155_new_n17241_));
OR2X2 OR2X2_3788 ( .A(u2__abc_52155_new_n17238_), .B(u2__abc_52155_new_n17242_), .Y(u2__0remLo_451_0__120_));
OR2X2 OR2X2_3789 ( .A(u2__abc_52155_new_n17246_), .B(u2__abc_52155_new_n17245_), .Y(u2__abc_52155_new_n17247_));
OR2X2 OR2X2_379 ( .A(_abc_73687_new_n1170_), .B(\a[77] ), .Y(_abc_73687_new_n1399_));
OR2X2 OR2X2_3790 ( .A(u2__abc_52155_new_n17244_), .B(u2__abc_52155_new_n17248_), .Y(u2__0remLo_451_0__121_));
OR2X2 OR2X2_3791 ( .A(u2__abc_52155_new_n17251_), .B(u2__abc_52155_new_n17252_), .Y(u2__abc_52155_new_n17253_));
OR2X2 OR2X2_3792 ( .A(u2__abc_52155_new_n17250_), .B(u2__abc_52155_new_n17254_), .Y(u2__0remLo_451_0__122_));
OR2X2 OR2X2_3793 ( .A(u2__abc_52155_new_n17257_), .B(u2__abc_52155_new_n17258_), .Y(u2__abc_52155_new_n17259_));
OR2X2 OR2X2_3794 ( .A(u2__abc_52155_new_n17256_), .B(u2__abc_52155_new_n17260_), .Y(u2__0remLo_451_0__123_));
OR2X2 OR2X2_3795 ( .A(u2__abc_52155_new_n17263_), .B(u2__abc_52155_new_n17264_), .Y(u2__abc_52155_new_n17265_));
OR2X2 OR2X2_3796 ( .A(u2__abc_52155_new_n17262_), .B(u2__abc_52155_new_n17266_), .Y(u2__0remLo_451_0__124_));
OR2X2 OR2X2_3797 ( .A(u2__abc_52155_new_n17270_), .B(u2__abc_52155_new_n17269_), .Y(u2__abc_52155_new_n17271_));
OR2X2 OR2X2_3798 ( .A(u2__abc_52155_new_n17268_), .B(u2__abc_52155_new_n17272_), .Y(u2__0remLo_451_0__125_));
OR2X2 OR2X2_3799 ( .A(u2__abc_52155_new_n17275_), .B(u2__abc_52155_new_n17276_), .Y(u2__abc_52155_new_n17277_));
OR2X2 OR2X2_38 ( .A(_abc_73687_new_n753_), .B(\a[18] ), .Y(_abc_73687_new_n885_));
OR2X2 OR2X2_380 ( .A(\a[112] ), .B(\a[77] ), .Y(_abc_73687_new_n1401_));
OR2X2 OR2X2_3800 ( .A(u2__abc_52155_new_n17274_), .B(u2__abc_52155_new_n17278_), .Y(u2__0remLo_451_0__126_));
OR2X2 OR2X2_3801 ( .A(u2__abc_52155_new_n17282_), .B(u2__abc_52155_new_n17281_), .Y(u2__abc_52155_new_n17283_));
OR2X2 OR2X2_3802 ( .A(u2__abc_52155_new_n17280_), .B(u2__abc_52155_new_n17284_), .Y(u2__0remLo_451_0__127_));
OR2X2 OR2X2_3803 ( .A(u2__abc_52155_new_n17288_), .B(u2__abc_52155_new_n17287_), .Y(u2__abc_52155_new_n17289_));
OR2X2 OR2X2_3804 ( .A(u2__abc_52155_new_n17286_), .B(u2__abc_52155_new_n17290_), .Y(u2__0remLo_451_0__128_));
OR2X2 OR2X2_3805 ( .A(u2__abc_52155_new_n17292_), .B(u2__abc_52155_new_n17293_), .Y(u2__abc_52155_new_n17294_));
OR2X2 OR2X2_3806 ( .A(u2__abc_52155_new_n17296_), .B(u2__abc_52155_new_n17297_), .Y(u2__abc_52155_new_n17298_));
OR2X2 OR2X2_3807 ( .A(u2__abc_52155_new_n17295_), .B(u2__abc_52155_new_n17299_), .Y(u2__0remLo_451_0__129_));
OR2X2 OR2X2_3808 ( .A(u2__abc_52155_new_n17303_), .B(u2__abc_52155_new_n17302_), .Y(u2__abc_52155_new_n17304_));
OR2X2 OR2X2_3809 ( .A(u2__abc_52155_new_n17301_), .B(u2__abc_52155_new_n17305_), .Y(u2__0remLo_451_0__130_));
OR2X2 OR2X2_381 ( .A(_abc_73687_new_n1170_), .B(\a[78] ), .Y(_abc_73687_new_n1402_));
OR2X2 OR2X2_3810 ( .A(u2__abc_52155_new_n17308_), .B(u2__abc_52155_new_n17309_), .Y(u2__abc_52155_new_n17310_));
OR2X2 OR2X2_3811 ( .A(u2__abc_52155_new_n17307_), .B(u2__abc_52155_new_n17311_), .Y(u2__0remLo_451_0__131_));
OR2X2 OR2X2_3812 ( .A(u2__abc_52155_new_n17314_), .B(u2__abc_52155_new_n17315_), .Y(u2__abc_52155_new_n17316_));
OR2X2 OR2X2_3813 ( .A(u2__abc_52155_new_n17313_), .B(u2__abc_52155_new_n17317_), .Y(u2__0remLo_451_0__132_));
OR2X2 OR2X2_3814 ( .A(u2__abc_52155_new_n17322_), .B(u2__abc_52155_new_n17320_), .Y(u2__abc_52155_new_n17323_));
OR2X2 OR2X2_3815 ( .A(u2__abc_52155_new_n17319_), .B(u2__abc_52155_new_n17323_), .Y(u2__0remLo_451_0__133_));
OR2X2 OR2X2_3816 ( .A(u2__abc_52155_new_n17327_), .B(u2__abc_52155_new_n17326_), .Y(u2__abc_52155_new_n17328_));
OR2X2 OR2X2_3817 ( .A(u2__abc_52155_new_n17325_), .B(u2__abc_52155_new_n17329_), .Y(u2__0remLo_451_0__134_));
OR2X2 OR2X2_3818 ( .A(u2__abc_52155_new_n17332_), .B(u2__abc_52155_new_n17333_), .Y(u2__abc_52155_new_n17334_));
OR2X2 OR2X2_3819 ( .A(u2__abc_52155_new_n17331_), .B(u2__abc_52155_new_n17335_), .Y(u2__0remLo_451_0__135_));
OR2X2 OR2X2_382 ( .A(\a[112] ), .B(\a[78] ), .Y(_abc_73687_new_n1404_));
OR2X2 OR2X2_3820 ( .A(u2__abc_52155_new_n17338_), .B(u2__abc_52155_new_n17339_), .Y(u2__abc_52155_new_n17340_));
OR2X2 OR2X2_3821 ( .A(u2__abc_52155_new_n17337_), .B(u2__abc_52155_new_n17341_), .Y(u2__0remLo_451_0__136_));
OR2X2 OR2X2_3822 ( .A(u2__abc_52155_new_n17344_), .B(u2__abc_52155_new_n17345_), .Y(u2__abc_52155_new_n17346_));
OR2X2 OR2X2_3823 ( .A(u2__abc_52155_new_n17343_), .B(u2__abc_52155_new_n17347_), .Y(u2__0remLo_451_0__137_));
OR2X2 OR2X2_3824 ( .A(u2__abc_52155_new_n17351_), .B(u2__abc_52155_new_n17350_), .Y(u2__abc_52155_new_n17352_));
OR2X2 OR2X2_3825 ( .A(u2__abc_52155_new_n17349_), .B(u2__abc_52155_new_n17353_), .Y(u2__0remLo_451_0__138_));
OR2X2 OR2X2_3826 ( .A(u2__abc_52155_new_n17356_), .B(u2__abc_52155_new_n17357_), .Y(u2__abc_52155_new_n17358_));
OR2X2 OR2X2_3827 ( .A(u2__abc_52155_new_n17355_), .B(u2__abc_52155_new_n17359_), .Y(u2__0remLo_451_0__139_));
OR2X2 OR2X2_3828 ( .A(u2__abc_52155_new_n17362_), .B(u2__abc_52155_new_n17363_), .Y(u2__abc_52155_new_n17364_));
OR2X2 OR2X2_3829 ( .A(u2__abc_52155_new_n17361_), .B(u2__abc_52155_new_n17365_), .Y(u2__0remLo_451_0__140_));
OR2X2 OR2X2_383 ( .A(_abc_73687_new_n1170_), .B(\a[79] ), .Y(_abc_73687_new_n1405_));
OR2X2 OR2X2_3830 ( .A(u2__abc_52155_new_n17368_), .B(u2__abc_52155_new_n17369_), .Y(u2__abc_52155_new_n17370_));
OR2X2 OR2X2_3831 ( .A(u2__abc_52155_new_n17367_), .B(u2__abc_52155_new_n17371_), .Y(u2__0remLo_451_0__141_));
OR2X2 OR2X2_3832 ( .A(u2__abc_52155_new_n17373_), .B(u2__abc_52155_new_n17374_), .Y(u2__abc_52155_new_n17375_));
OR2X2 OR2X2_3833 ( .A(u2__abc_52155_new_n17377_), .B(u2__abc_52155_new_n17378_), .Y(u2__abc_52155_new_n17379_));
OR2X2 OR2X2_3834 ( .A(u2__abc_52155_new_n17376_), .B(u2__abc_52155_new_n17380_), .Y(u2__0remLo_451_0__142_));
OR2X2 OR2X2_3835 ( .A(u2__abc_52155_new_n17384_), .B(u2__abc_52155_new_n17383_), .Y(u2__abc_52155_new_n17385_));
OR2X2 OR2X2_3836 ( .A(u2__abc_52155_new_n17382_), .B(u2__abc_52155_new_n17386_), .Y(u2__0remLo_451_0__143_));
OR2X2 OR2X2_3837 ( .A(u2__abc_52155_new_n17389_), .B(u2__abc_52155_new_n17390_), .Y(u2__abc_52155_new_n17391_));
OR2X2 OR2X2_3838 ( .A(u2__abc_52155_new_n17388_), .B(u2__abc_52155_new_n17392_), .Y(u2__0remLo_451_0__144_));
OR2X2 OR2X2_3839 ( .A(u2__abc_52155_new_n17395_), .B(u2__abc_52155_new_n17396_), .Y(u2__abc_52155_new_n17397_));
OR2X2 OR2X2_384 ( .A(\a[112] ), .B(\a[79] ), .Y(_abc_73687_new_n1407_));
OR2X2 OR2X2_3840 ( .A(u2__abc_52155_new_n17394_), .B(u2__abc_52155_new_n17398_), .Y(u2__0remLo_451_0__145_));
OR2X2 OR2X2_3841 ( .A(u2__abc_52155_new_n17401_), .B(u2__abc_52155_new_n17402_), .Y(u2__abc_52155_new_n17403_));
OR2X2 OR2X2_3842 ( .A(u2__abc_52155_new_n17400_), .B(u2__abc_52155_new_n17404_), .Y(u2__0remLo_451_0__146_));
OR2X2 OR2X2_3843 ( .A(u2__abc_52155_new_n17408_), .B(u2__abc_52155_new_n17407_), .Y(u2__abc_52155_new_n17409_));
OR2X2 OR2X2_3844 ( .A(u2__abc_52155_new_n17406_), .B(u2__abc_52155_new_n17410_), .Y(u2__0remLo_451_0__147_));
OR2X2 OR2X2_3845 ( .A(u2__abc_52155_new_n17413_), .B(u2__abc_52155_new_n17414_), .Y(u2__abc_52155_new_n17415_));
OR2X2 OR2X2_3846 ( .A(u2__abc_52155_new_n17412_), .B(u2__abc_52155_new_n17416_), .Y(u2__0remLo_451_0__148_));
OR2X2 OR2X2_3847 ( .A(u2__abc_52155_new_n17419_), .B(u2__abc_52155_new_n17420_), .Y(u2__abc_52155_new_n17421_));
OR2X2 OR2X2_3848 ( .A(u2__abc_52155_new_n17418_), .B(u2__abc_52155_new_n17422_), .Y(u2__0remLo_451_0__149_));
OR2X2 OR2X2_3849 ( .A(u2__abc_52155_new_n17425_), .B(u2__abc_52155_new_n17426_), .Y(u2__abc_52155_new_n17427_));
OR2X2 OR2X2_385 ( .A(_abc_73687_new_n1170_), .B(\a[80] ), .Y(_abc_73687_new_n1408_));
OR2X2 OR2X2_3850 ( .A(u2__abc_52155_new_n17424_), .B(u2__abc_52155_new_n17428_), .Y(u2__0remLo_451_0__150_));
OR2X2 OR2X2_3851 ( .A(u2__abc_52155_new_n17431_), .B(u2__abc_52155_new_n17432_), .Y(u2__abc_52155_new_n17433_));
OR2X2 OR2X2_3852 ( .A(u2__abc_52155_new_n17430_), .B(u2__abc_52155_new_n17434_), .Y(u2__0remLo_451_0__151_));
OR2X2 OR2X2_3853 ( .A(u2__abc_52155_new_n17437_), .B(u2__abc_52155_new_n17438_), .Y(u2__abc_52155_new_n17439_));
OR2X2 OR2X2_3854 ( .A(u2__abc_52155_new_n17436_), .B(u2__abc_52155_new_n17440_), .Y(u2__0remLo_451_0__152_));
OR2X2 OR2X2_3855 ( .A(u2__abc_52155_new_n17444_), .B(u2__abc_52155_new_n17443_), .Y(u2__abc_52155_new_n17445_));
OR2X2 OR2X2_3856 ( .A(u2__abc_52155_new_n17442_), .B(u2__abc_52155_new_n17446_), .Y(u2__0remLo_451_0__153_));
OR2X2 OR2X2_3857 ( .A(u2__abc_52155_new_n17450_), .B(u2__abc_52155_new_n17449_), .Y(u2__abc_52155_new_n17451_));
OR2X2 OR2X2_3858 ( .A(u2__abc_52155_new_n17448_), .B(u2__abc_52155_new_n17452_), .Y(u2__0remLo_451_0__154_));
OR2X2 OR2X2_3859 ( .A(u2__abc_52155_new_n17455_), .B(u2__abc_52155_new_n17456_), .Y(u2__abc_52155_new_n17457_));
OR2X2 OR2X2_386 ( .A(\a[112] ), .B(\a[80] ), .Y(_abc_73687_new_n1410_));
OR2X2 OR2X2_3860 ( .A(u2__abc_52155_new_n17454_), .B(u2__abc_52155_new_n17458_), .Y(u2__0remLo_451_0__155_));
OR2X2 OR2X2_3861 ( .A(u2__abc_52155_new_n17461_), .B(u2__abc_52155_new_n17462_), .Y(u2__abc_52155_new_n17463_));
OR2X2 OR2X2_3862 ( .A(u2__abc_52155_new_n17460_), .B(u2__abc_52155_new_n17464_), .Y(u2__0remLo_451_0__156_));
OR2X2 OR2X2_3863 ( .A(u2__abc_52155_new_n17467_), .B(u2__abc_52155_new_n17468_), .Y(u2__abc_52155_new_n17469_));
OR2X2 OR2X2_3864 ( .A(u2__abc_52155_new_n17466_), .B(u2__abc_52155_new_n17470_), .Y(u2__0remLo_451_0__157_));
OR2X2 OR2X2_3865 ( .A(u2__abc_52155_new_n17473_), .B(u2__abc_52155_new_n17474_), .Y(u2__abc_52155_new_n17475_));
OR2X2 OR2X2_3866 ( .A(u2__abc_52155_new_n17472_), .B(u2__abc_52155_new_n17476_), .Y(u2__0remLo_451_0__158_));
OR2X2 OR2X2_3867 ( .A(u2__abc_52155_new_n17479_), .B(u2__abc_52155_new_n17480_), .Y(u2__abc_52155_new_n17481_));
OR2X2 OR2X2_3868 ( .A(u2__abc_52155_new_n17478_), .B(u2__abc_52155_new_n17482_), .Y(u2__0remLo_451_0__159_));
OR2X2 OR2X2_3869 ( .A(u2__abc_52155_new_n17484_), .B(u2__abc_52155_new_n17485_), .Y(u2__abc_52155_new_n17486_));
OR2X2 OR2X2_387 ( .A(_abc_73687_new_n1170_), .B(\a[81] ), .Y(_abc_73687_new_n1411_));
OR2X2 OR2X2_3870 ( .A(u2__abc_52155_new_n17488_), .B(u2__abc_52155_new_n17489_), .Y(u2__abc_52155_new_n17490_));
OR2X2 OR2X2_3871 ( .A(u2__abc_52155_new_n17487_), .B(u2__abc_52155_new_n17491_), .Y(u2__0remLo_451_0__160_));
OR2X2 OR2X2_3872 ( .A(u2__abc_52155_new_n17493_), .B(u2__abc_52155_new_n17494_), .Y(u2__abc_52155_new_n17495_));
OR2X2 OR2X2_3873 ( .A(u2__abc_52155_new_n17497_), .B(u2__abc_52155_new_n17498_), .Y(u2__abc_52155_new_n17499_));
OR2X2 OR2X2_3874 ( .A(u2__abc_52155_new_n17496_), .B(u2__abc_52155_new_n17500_), .Y(u2__0remLo_451_0__161_));
OR2X2 OR2X2_3875 ( .A(u2__abc_52155_new_n17503_), .B(u2__abc_52155_new_n17504_), .Y(u2__abc_52155_new_n17505_));
OR2X2 OR2X2_3876 ( .A(u2__abc_52155_new_n17502_), .B(u2__abc_52155_new_n17506_), .Y(u2__0remLo_451_0__162_));
OR2X2 OR2X2_3877 ( .A(u2__abc_52155_new_n17509_), .B(u2__abc_52155_new_n17510_), .Y(u2__abc_52155_new_n17511_));
OR2X2 OR2X2_3878 ( .A(u2__abc_52155_new_n17508_), .B(u2__abc_52155_new_n17512_), .Y(u2__0remLo_451_0__163_));
OR2X2 OR2X2_3879 ( .A(u2__abc_52155_new_n17515_), .B(u2__abc_52155_new_n17516_), .Y(u2__abc_52155_new_n17517_));
OR2X2 OR2X2_388 ( .A(\a[112] ), .B(\a[81] ), .Y(_abc_73687_new_n1413_));
OR2X2 OR2X2_3880 ( .A(u2__abc_52155_new_n17514_), .B(u2__abc_52155_new_n17518_), .Y(u2__0remLo_451_0__164_));
OR2X2 OR2X2_3881 ( .A(u2__abc_52155_new_n17521_), .B(u2__abc_52155_new_n17522_), .Y(u2__abc_52155_new_n17523_));
OR2X2 OR2X2_3882 ( .A(u2__abc_52155_new_n17520_), .B(u2__abc_52155_new_n17524_), .Y(u2__0remLo_451_0__165_));
OR2X2 OR2X2_3883 ( .A(u2__abc_52155_new_n17528_), .B(u2__abc_52155_new_n17527_), .Y(u2__abc_52155_new_n17529_));
OR2X2 OR2X2_3884 ( .A(u2__abc_52155_new_n17526_), .B(u2__abc_52155_new_n17530_), .Y(u2__0remLo_451_0__166_));
OR2X2 OR2X2_3885 ( .A(u2__abc_52155_new_n17533_), .B(u2__abc_52155_new_n17534_), .Y(u2__abc_52155_new_n17535_));
OR2X2 OR2X2_3886 ( .A(u2__abc_52155_new_n17532_), .B(u2__abc_52155_new_n17536_), .Y(u2__0remLo_451_0__167_));
OR2X2 OR2X2_3887 ( .A(u2__abc_52155_new_n17539_), .B(u2__abc_52155_new_n17540_), .Y(u2__abc_52155_new_n17541_));
OR2X2 OR2X2_3888 ( .A(u2__abc_52155_new_n17538_), .B(u2__abc_52155_new_n17542_), .Y(u2__0remLo_451_0__168_));
OR2X2 OR2X2_3889 ( .A(u2__abc_52155_new_n17545_), .B(u2__abc_52155_new_n17546_), .Y(u2__abc_52155_new_n17547_));
OR2X2 OR2X2_389 ( .A(_abc_73687_new_n1170_), .B(\a[82] ), .Y(_abc_73687_new_n1414_));
OR2X2 OR2X2_3890 ( .A(u2__abc_52155_new_n17544_), .B(u2__abc_52155_new_n17548_), .Y(u2__0remLo_451_0__169_));
OR2X2 OR2X2_3891 ( .A(u2__abc_52155_new_n17552_), .B(u2__abc_52155_new_n17551_), .Y(u2__abc_52155_new_n17553_));
OR2X2 OR2X2_3892 ( .A(u2__abc_52155_new_n17550_), .B(u2__abc_52155_new_n17554_), .Y(u2__0remLo_451_0__170_));
OR2X2 OR2X2_3893 ( .A(u2__abc_52155_new_n17557_), .B(u2__abc_52155_new_n17558_), .Y(u2__abc_52155_new_n17559_));
OR2X2 OR2X2_3894 ( .A(u2__abc_52155_new_n17556_), .B(u2__abc_52155_new_n17560_), .Y(u2__0remLo_451_0__171_));
OR2X2 OR2X2_3895 ( .A(u2__abc_52155_new_n17563_), .B(u2__abc_52155_new_n17564_), .Y(u2__abc_52155_new_n17565_));
OR2X2 OR2X2_3896 ( .A(u2__abc_52155_new_n17562_), .B(u2__abc_52155_new_n17566_), .Y(u2__0remLo_451_0__172_));
OR2X2 OR2X2_3897 ( .A(u2__abc_52155_new_n17569_), .B(u2__abc_52155_new_n17570_), .Y(u2__abc_52155_new_n17571_));
OR2X2 OR2X2_3898 ( .A(u2__abc_52155_new_n17568_), .B(u2__abc_52155_new_n17572_), .Y(u2__0remLo_451_0__173_));
OR2X2 OR2X2_3899 ( .A(u2__abc_52155_new_n17577_), .B(u2__abc_52155_new_n17575_), .Y(u2__abc_52155_new_n17578_));
OR2X2 OR2X2_39 ( .A(aNan), .B(sqrto_95_), .Y(_abc_73687_new_n887_));
OR2X2 OR2X2_390 ( .A(\a[112] ), .B(\a[82] ), .Y(_abc_73687_new_n1416_));
OR2X2 OR2X2_3900 ( .A(u2__abc_52155_new_n17574_), .B(u2__abc_52155_new_n17578_), .Y(u2__0remLo_451_0__174_));
OR2X2 OR2X2_3901 ( .A(u2__abc_52155_new_n17581_), .B(u2__abc_52155_new_n17582_), .Y(u2__abc_52155_new_n17583_));
OR2X2 OR2X2_3902 ( .A(u2__abc_52155_new_n17580_), .B(u2__abc_52155_new_n17584_), .Y(u2__0remLo_451_0__175_));
OR2X2 OR2X2_3903 ( .A(u2__abc_52155_new_n17587_), .B(u2__abc_52155_new_n17588_), .Y(u2__abc_52155_new_n17589_));
OR2X2 OR2X2_3904 ( .A(u2__abc_52155_new_n17586_), .B(u2__abc_52155_new_n17590_), .Y(u2__0remLo_451_0__176_));
OR2X2 OR2X2_3905 ( .A(u2__abc_52155_new_n17593_), .B(u2__abc_52155_new_n17594_), .Y(u2__abc_52155_new_n17595_));
OR2X2 OR2X2_3906 ( .A(u2__abc_52155_new_n17592_), .B(u2__abc_52155_new_n17596_), .Y(u2__0remLo_451_0__177_));
OR2X2 OR2X2_3907 ( .A(u2__abc_52155_new_n17599_), .B(u2__abc_52155_new_n17600_), .Y(u2__abc_52155_new_n17601_));
OR2X2 OR2X2_3908 ( .A(u2__abc_52155_new_n17598_), .B(u2__abc_52155_new_n17602_), .Y(u2__0remLo_451_0__178_));
OR2X2 OR2X2_3909 ( .A(u2__abc_52155_new_n17605_), .B(u2__abc_52155_new_n17606_), .Y(u2__abc_52155_new_n17607_));
OR2X2 OR2X2_391 ( .A(_abc_73687_new_n1170_), .B(\a[83] ), .Y(_abc_73687_new_n1417_));
OR2X2 OR2X2_3910 ( .A(u2__abc_52155_new_n17604_), .B(u2__abc_52155_new_n17608_), .Y(u2__0remLo_451_0__179_));
OR2X2 OR2X2_3911 ( .A(u2__abc_52155_new_n17611_), .B(u2__abc_52155_new_n17612_), .Y(u2__abc_52155_new_n17613_));
OR2X2 OR2X2_3912 ( .A(u2__abc_52155_new_n17610_), .B(u2__abc_52155_new_n17614_), .Y(u2__0remLo_451_0__180_));
OR2X2 OR2X2_3913 ( .A(u2__abc_52155_new_n17617_), .B(u2__abc_52155_new_n17618_), .Y(u2__abc_52155_new_n17619_));
OR2X2 OR2X2_3914 ( .A(u2__abc_52155_new_n17616_), .B(u2__abc_52155_new_n17620_), .Y(u2__0remLo_451_0__181_));
OR2X2 OR2X2_3915 ( .A(u2__abc_52155_new_n17623_), .B(u2__abc_52155_new_n17624_), .Y(u2__abc_52155_new_n17625_));
OR2X2 OR2X2_3916 ( .A(u2__abc_52155_new_n17622_), .B(u2__abc_52155_new_n17626_), .Y(u2__0remLo_451_0__182_));
OR2X2 OR2X2_3917 ( .A(u2__abc_52155_new_n17629_), .B(u2__abc_52155_new_n17630_), .Y(u2__abc_52155_new_n17631_));
OR2X2 OR2X2_3918 ( .A(u2__abc_52155_new_n17628_), .B(u2__abc_52155_new_n17632_), .Y(u2__0remLo_451_0__183_));
OR2X2 OR2X2_3919 ( .A(u2__abc_52155_new_n17635_), .B(u2__abc_52155_new_n17636_), .Y(u2__abc_52155_new_n17637_));
OR2X2 OR2X2_392 ( .A(\a[112] ), .B(\a[83] ), .Y(_abc_73687_new_n1419_));
OR2X2 OR2X2_3920 ( .A(u2__abc_52155_new_n17634_), .B(u2__abc_52155_new_n17638_), .Y(u2__0remLo_451_0__184_));
OR2X2 OR2X2_3921 ( .A(u2__abc_52155_new_n17642_), .B(u2__abc_52155_new_n17641_), .Y(u2__abc_52155_new_n17643_));
OR2X2 OR2X2_3922 ( .A(u2__abc_52155_new_n17640_), .B(u2__abc_52155_new_n17644_), .Y(u2__0remLo_451_0__185_));
OR2X2 OR2X2_3923 ( .A(u2__abc_52155_new_n17648_), .B(u2__abc_52155_new_n17647_), .Y(u2__abc_52155_new_n17649_));
OR2X2 OR2X2_3924 ( .A(u2__abc_52155_new_n17646_), .B(u2__abc_52155_new_n17650_), .Y(u2__0remLo_451_0__186_));
OR2X2 OR2X2_3925 ( .A(u2__abc_52155_new_n17653_), .B(u2__abc_52155_new_n17654_), .Y(u2__abc_52155_new_n17655_));
OR2X2 OR2X2_3926 ( .A(u2__abc_52155_new_n17652_), .B(u2__abc_52155_new_n17656_), .Y(u2__0remLo_451_0__187_));
OR2X2 OR2X2_3927 ( .A(u2__abc_52155_new_n17659_), .B(u2__abc_52155_new_n17660_), .Y(u2__abc_52155_new_n17661_));
OR2X2 OR2X2_3928 ( .A(u2__abc_52155_new_n17658_), .B(u2__abc_52155_new_n17662_), .Y(u2__0remLo_451_0__188_));
OR2X2 OR2X2_3929 ( .A(u2__abc_52155_new_n17666_), .B(u2__abc_52155_new_n17665_), .Y(u2__abc_52155_new_n17667_));
OR2X2 OR2X2_393 ( .A(_abc_73687_new_n1170_), .B(\a[84] ), .Y(_abc_73687_new_n1420_));
OR2X2 OR2X2_3930 ( .A(u2__abc_52155_new_n17664_), .B(u2__abc_52155_new_n17668_), .Y(u2__0remLo_451_0__189_));
OR2X2 OR2X2_3931 ( .A(u2__abc_52155_new_n17671_), .B(u2__abc_52155_new_n17672_), .Y(u2__abc_52155_new_n17673_));
OR2X2 OR2X2_3932 ( .A(u2__abc_52155_new_n17670_), .B(u2__abc_52155_new_n17674_), .Y(u2__0remLo_451_0__190_));
OR2X2 OR2X2_3933 ( .A(u2__abc_52155_new_n17678_), .B(u2__abc_52155_new_n17677_), .Y(u2__abc_52155_new_n17679_));
OR2X2 OR2X2_3934 ( .A(u2__abc_52155_new_n17676_), .B(u2__abc_52155_new_n17680_), .Y(u2__0remLo_451_0__191_));
OR2X2 OR2X2_3935 ( .A(u2__abc_52155_new_n17684_), .B(u2__abc_52155_new_n17683_), .Y(u2__abc_52155_new_n17685_));
OR2X2 OR2X2_3936 ( .A(u2__abc_52155_new_n17682_), .B(u2__abc_52155_new_n17686_), .Y(u2__0remLo_451_0__192_));
OR2X2 OR2X2_3937 ( .A(u2__abc_52155_new_n17688_), .B(u2__abc_52155_new_n17689_), .Y(u2__abc_52155_new_n17690_));
OR2X2 OR2X2_3938 ( .A(u2__abc_52155_new_n17692_), .B(u2__abc_52155_new_n17693_), .Y(u2__abc_52155_new_n17694_));
OR2X2 OR2X2_3939 ( .A(u2__abc_52155_new_n17691_), .B(u2__abc_52155_new_n17695_), .Y(u2__0remLo_451_0__193_));
OR2X2 OR2X2_394 ( .A(\a[112] ), .B(\a[84] ), .Y(_abc_73687_new_n1422_));
OR2X2 OR2X2_3940 ( .A(u2__abc_52155_new_n17698_), .B(u2__abc_52155_new_n17699_), .Y(u2__abc_52155_new_n17700_));
OR2X2 OR2X2_3941 ( .A(u2__abc_52155_new_n17697_), .B(u2__abc_52155_new_n17701_), .Y(u2__0remLo_451_0__194_));
OR2X2 OR2X2_3942 ( .A(u2__abc_52155_new_n17704_), .B(u2__abc_52155_new_n17705_), .Y(u2__abc_52155_new_n17706_));
OR2X2 OR2X2_3943 ( .A(u2__abc_52155_new_n17703_), .B(u2__abc_52155_new_n17707_), .Y(u2__0remLo_451_0__195_));
OR2X2 OR2X2_3944 ( .A(u2__abc_52155_new_n17710_), .B(u2__abc_52155_new_n17711_), .Y(u2__abc_52155_new_n17712_));
OR2X2 OR2X2_3945 ( .A(u2__abc_52155_new_n17709_), .B(u2__abc_52155_new_n17713_), .Y(u2__0remLo_451_0__196_));
OR2X2 OR2X2_3946 ( .A(u2__abc_52155_new_n17716_), .B(u2__abc_52155_new_n17717_), .Y(u2__abc_52155_new_n17718_));
OR2X2 OR2X2_3947 ( .A(u2__abc_52155_new_n17715_), .B(u2__abc_52155_new_n17719_), .Y(u2__0remLo_451_0__197_));
OR2X2 OR2X2_3948 ( .A(u2__abc_52155_new_n17723_), .B(u2__abc_52155_new_n17722_), .Y(u2__abc_52155_new_n17724_));
OR2X2 OR2X2_3949 ( .A(u2__abc_52155_new_n17721_), .B(u2__abc_52155_new_n17725_), .Y(u2__0remLo_451_0__198_));
OR2X2 OR2X2_395 ( .A(_abc_73687_new_n1170_), .B(\a[85] ), .Y(_abc_73687_new_n1423_));
OR2X2 OR2X2_3950 ( .A(u2__abc_52155_new_n17728_), .B(u2__abc_52155_new_n17729_), .Y(u2__abc_52155_new_n17730_));
OR2X2 OR2X2_3951 ( .A(u2__abc_52155_new_n17727_), .B(u2__abc_52155_new_n17731_), .Y(u2__0remLo_451_0__199_));
OR2X2 OR2X2_3952 ( .A(u2__abc_52155_new_n17734_), .B(u2__abc_52155_new_n17735_), .Y(u2__abc_52155_new_n17736_));
OR2X2 OR2X2_3953 ( .A(u2__abc_52155_new_n17733_), .B(u2__abc_52155_new_n17737_), .Y(u2__0remLo_451_0__200_));
OR2X2 OR2X2_3954 ( .A(u2__abc_52155_new_n17740_), .B(u2__abc_52155_new_n17741_), .Y(u2__abc_52155_new_n17742_));
OR2X2 OR2X2_3955 ( .A(u2__abc_52155_new_n17739_), .B(u2__abc_52155_new_n17743_), .Y(u2__0remLo_451_0__201_));
OR2X2 OR2X2_3956 ( .A(u2__abc_52155_new_n17745_), .B(u2__abc_52155_new_n17746_), .Y(u2__abc_52155_new_n17747_));
OR2X2 OR2X2_3957 ( .A(u2__abc_52155_new_n17749_), .B(u2__abc_52155_new_n17750_), .Y(u2__abc_52155_new_n17751_));
OR2X2 OR2X2_3958 ( .A(u2__abc_52155_new_n17748_), .B(u2__abc_52155_new_n17752_), .Y(u2__0remLo_451_0__202_));
OR2X2 OR2X2_3959 ( .A(u2__abc_52155_new_n17755_), .B(u2__abc_52155_new_n17756_), .Y(u2__abc_52155_new_n17757_));
OR2X2 OR2X2_396 ( .A(\a[112] ), .B(\a[85] ), .Y(_abc_73687_new_n1425_));
OR2X2 OR2X2_3960 ( .A(u2__abc_52155_new_n17754_), .B(u2__abc_52155_new_n17758_), .Y(u2__0remLo_451_0__203_));
OR2X2 OR2X2_3961 ( .A(u2__abc_52155_new_n17761_), .B(u2__abc_52155_new_n17762_), .Y(u2__abc_52155_new_n17763_));
OR2X2 OR2X2_3962 ( .A(u2__abc_52155_new_n17760_), .B(u2__abc_52155_new_n17764_), .Y(u2__0remLo_451_0__204_));
OR2X2 OR2X2_3963 ( .A(u2__abc_52155_new_n17767_), .B(u2__abc_52155_new_n17768_), .Y(u2__abc_52155_new_n17769_));
OR2X2 OR2X2_3964 ( .A(u2__abc_52155_new_n17766_), .B(u2__abc_52155_new_n17770_), .Y(u2__0remLo_451_0__205_));
OR2X2 OR2X2_3965 ( .A(u2__abc_52155_new_n17775_), .B(u2__abc_52155_new_n17773_), .Y(u2__abc_52155_new_n17776_));
OR2X2 OR2X2_3966 ( .A(u2__abc_52155_new_n17772_), .B(u2__abc_52155_new_n17776_), .Y(u2__0remLo_451_0__206_));
OR2X2 OR2X2_3967 ( .A(u2__abc_52155_new_n17780_), .B(u2__abc_52155_new_n17779_), .Y(u2__abc_52155_new_n17781_));
OR2X2 OR2X2_3968 ( .A(u2__abc_52155_new_n17778_), .B(u2__abc_52155_new_n17782_), .Y(u2__0remLo_451_0__207_));
OR2X2 OR2X2_3969 ( .A(u2__abc_52155_new_n17785_), .B(u2__abc_52155_new_n17786_), .Y(u2__abc_52155_new_n17787_));
OR2X2 OR2X2_397 ( .A(_abc_73687_new_n1170_), .B(\a[86] ), .Y(_abc_73687_new_n1426_));
OR2X2 OR2X2_3970 ( .A(u2__abc_52155_new_n17784_), .B(u2__abc_52155_new_n17788_), .Y(u2__0remLo_451_0__208_));
OR2X2 OR2X2_3971 ( .A(u2__abc_52155_new_n17791_), .B(u2__abc_52155_new_n17792_), .Y(u2__abc_52155_new_n17793_));
OR2X2 OR2X2_3972 ( .A(u2__abc_52155_new_n17790_), .B(u2__abc_52155_new_n17794_), .Y(u2__0remLo_451_0__209_));
OR2X2 OR2X2_3973 ( .A(u2__abc_52155_new_n17797_), .B(u2__abc_52155_new_n17798_), .Y(u2__abc_52155_new_n17799_));
OR2X2 OR2X2_3974 ( .A(u2__abc_52155_new_n17796_), .B(u2__abc_52155_new_n17800_), .Y(u2__0remLo_451_0__210_));
OR2X2 OR2X2_3975 ( .A(u2__abc_52155_new_n17804_), .B(u2__abc_52155_new_n17803_), .Y(u2__abc_52155_new_n17805_));
OR2X2 OR2X2_3976 ( .A(u2__abc_52155_new_n17802_), .B(u2__abc_52155_new_n17806_), .Y(u2__0remLo_451_0__211_));
OR2X2 OR2X2_3977 ( .A(u2__abc_52155_new_n17809_), .B(u2__abc_52155_new_n17810_), .Y(u2__abc_52155_new_n17811_));
OR2X2 OR2X2_3978 ( .A(u2__abc_52155_new_n17808_), .B(u2__abc_52155_new_n17812_), .Y(u2__0remLo_451_0__212_));
OR2X2 OR2X2_3979 ( .A(u2__abc_52155_new_n17815_), .B(u2__abc_52155_new_n17816_), .Y(u2__abc_52155_new_n17817_));
OR2X2 OR2X2_398 ( .A(\a[112] ), .B(\a[86] ), .Y(_abc_73687_new_n1428_));
OR2X2 OR2X2_3980 ( .A(u2__abc_52155_new_n17814_), .B(u2__abc_52155_new_n17818_), .Y(u2__0remLo_451_0__213_));
OR2X2 OR2X2_3981 ( .A(u2__abc_52155_new_n17821_), .B(u2__abc_52155_new_n17822_), .Y(u2__abc_52155_new_n17823_));
OR2X2 OR2X2_3982 ( .A(u2__abc_52155_new_n17820_), .B(u2__abc_52155_new_n17824_), .Y(u2__0remLo_451_0__214_));
OR2X2 OR2X2_3983 ( .A(u2__abc_52155_new_n17827_), .B(u2__abc_52155_new_n17828_), .Y(u2__abc_52155_new_n17829_));
OR2X2 OR2X2_3984 ( .A(u2__abc_52155_new_n17826_), .B(u2__abc_52155_new_n17830_), .Y(u2__0remLo_451_0__215_));
OR2X2 OR2X2_3985 ( .A(u2__abc_52155_new_n17833_), .B(u2__abc_52155_new_n17834_), .Y(u2__abc_52155_new_n17835_));
OR2X2 OR2X2_3986 ( .A(u2__abc_52155_new_n17832_), .B(u2__abc_52155_new_n17836_), .Y(u2__0remLo_451_0__216_));
OR2X2 OR2X2_3987 ( .A(u2__abc_52155_new_n17840_), .B(u2__abc_52155_new_n17839_), .Y(u2__abc_52155_new_n17841_));
OR2X2 OR2X2_3988 ( .A(u2__abc_52155_new_n17838_), .B(u2__abc_52155_new_n17842_), .Y(u2__0remLo_451_0__217_));
OR2X2 OR2X2_3989 ( .A(u2__abc_52155_new_n17846_), .B(u2__abc_52155_new_n17845_), .Y(u2__abc_52155_new_n17847_));
OR2X2 OR2X2_399 ( .A(_abc_73687_new_n1170_), .B(\a[87] ), .Y(_abc_73687_new_n1429_));
OR2X2 OR2X2_3990 ( .A(u2__abc_52155_new_n17844_), .B(u2__abc_52155_new_n17848_), .Y(u2__0remLo_451_0__218_));
OR2X2 OR2X2_3991 ( .A(u2__abc_52155_new_n17851_), .B(u2__abc_52155_new_n17852_), .Y(u2__abc_52155_new_n17853_));
OR2X2 OR2X2_3992 ( .A(u2__abc_52155_new_n17850_), .B(u2__abc_52155_new_n17854_), .Y(u2__0remLo_451_0__219_));
OR2X2 OR2X2_3993 ( .A(u2__abc_52155_new_n17857_), .B(u2__abc_52155_new_n17858_), .Y(u2__abc_52155_new_n17859_));
OR2X2 OR2X2_3994 ( .A(u2__abc_52155_new_n17856_), .B(u2__abc_52155_new_n17860_), .Y(u2__0remLo_451_0__220_));
OR2X2 OR2X2_3995 ( .A(u2__abc_52155_new_n17863_), .B(u2__abc_52155_new_n17864_), .Y(u2__abc_52155_new_n17865_));
OR2X2 OR2X2_3996 ( .A(u2__abc_52155_new_n17862_), .B(u2__abc_52155_new_n17866_), .Y(u2__0remLo_451_0__221_));
OR2X2 OR2X2_3997 ( .A(u2__abc_52155_new_n17869_), .B(u2__abc_52155_new_n17870_), .Y(u2__abc_52155_new_n17871_));
OR2X2 OR2X2_3998 ( .A(u2__abc_52155_new_n17868_), .B(u2__abc_52155_new_n17872_), .Y(u2__0remLo_451_0__222_));
OR2X2 OR2X2_3999 ( .A(u2__abc_52155_new_n17876_), .B(u2__abc_52155_new_n17875_), .Y(u2__abc_52155_new_n17877_));
OR2X2 OR2X2_4 ( .A(_abc_73687_new_n753_), .B(\a[1] ), .Y(_abc_73687_new_n834_));
OR2X2 OR2X2_40 ( .A(_abc_73687_new_n753_), .B(\a[19] ), .Y(_abc_73687_new_n888_));
OR2X2 OR2X2_400 ( .A(\a[112] ), .B(\a[87] ), .Y(_abc_73687_new_n1431_));
OR2X2 OR2X2_4000 ( .A(u2__abc_52155_new_n17874_), .B(u2__abc_52155_new_n17878_), .Y(u2__0remLo_451_0__223_));
OR2X2 OR2X2_4001 ( .A(u2__abc_52155_new_n17881_), .B(u2__abc_52155_new_n17882_), .Y(u2__abc_52155_new_n17883_));
OR2X2 OR2X2_4002 ( .A(u2__abc_52155_new_n17880_), .B(u2__abc_52155_new_n17884_), .Y(u2__0remLo_451_0__224_));
OR2X2 OR2X2_4003 ( .A(u2__abc_52155_new_n17886_), .B(u2__abc_52155_new_n17887_), .Y(u2__abc_52155_new_n17888_));
OR2X2 OR2X2_4004 ( .A(u2__abc_52155_new_n17890_), .B(u2__abc_52155_new_n17891_), .Y(u2__abc_52155_new_n17892_));
OR2X2 OR2X2_4005 ( .A(u2__abc_52155_new_n17889_), .B(u2__abc_52155_new_n17893_), .Y(u2__0remLo_451_0__225_));
OR2X2 OR2X2_4006 ( .A(u2__abc_52155_new_n17895_), .B(u2__abc_52155_new_n17896_), .Y(u2__abc_52155_new_n17897_));
OR2X2 OR2X2_4007 ( .A(u2__abc_52155_new_n17899_), .B(u2__abc_52155_new_n17900_), .Y(u2__abc_52155_new_n17901_));
OR2X2 OR2X2_4008 ( .A(u2__abc_52155_new_n17898_), .B(u2__abc_52155_new_n17902_), .Y(u2__0remLo_451_0__226_));
OR2X2 OR2X2_4009 ( .A(u2__abc_52155_new_n17905_), .B(u2__abc_52155_new_n17906_), .Y(u2__abc_52155_new_n17907_));
OR2X2 OR2X2_401 ( .A(_abc_73687_new_n1170_), .B(\a[88] ), .Y(_abc_73687_new_n1432_));
OR2X2 OR2X2_4010 ( .A(u2__abc_52155_new_n17904_), .B(u2__abc_52155_new_n17908_), .Y(u2__0remLo_451_0__227_));
OR2X2 OR2X2_4011 ( .A(u2__abc_52155_new_n17911_), .B(u2__abc_52155_new_n17912_), .Y(u2__abc_52155_new_n17913_));
OR2X2 OR2X2_4012 ( .A(u2__abc_52155_new_n17910_), .B(u2__abc_52155_new_n17914_), .Y(u2__0remLo_451_0__228_));
OR2X2 OR2X2_4013 ( .A(u2__abc_52155_new_n17917_), .B(u2__abc_52155_new_n17918_), .Y(u2__abc_52155_new_n17919_));
OR2X2 OR2X2_4014 ( .A(u2__abc_52155_new_n17916_), .B(u2__abc_52155_new_n17920_), .Y(u2__0remLo_451_0__229_));
OR2X2 OR2X2_4015 ( .A(u2__abc_52155_new_n17923_), .B(u2__abc_52155_new_n17924_), .Y(u2__abc_52155_new_n17925_));
OR2X2 OR2X2_4016 ( .A(u2__abc_52155_new_n17922_), .B(u2__abc_52155_new_n17926_), .Y(u2__0remLo_451_0__230_));
OR2X2 OR2X2_4017 ( .A(u2__abc_52155_new_n17929_), .B(u2__abc_52155_new_n17930_), .Y(u2__abc_52155_new_n17931_));
OR2X2 OR2X2_4018 ( .A(u2__abc_52155_new_n17928_), .B(u2__abc_52155_new_n17932_), .Y(u2__0remLo_451_0__231_));
OR2X2 OR2X2_4019 ( .A(u2__abc_52155_new_n17935_), .B(u2__abc_52155_new_n17936_), .Y(u2__abc_52155_new_n17937_));
OR2X2 OR2X2_402 ( .A(\a[112] ), .B(\a[88] ), .Y(_abc_73687_new_n1434_));
OR2X2 OR2X2_4020 ( .A(u2__abc_52155_new_n17934_), .B(u2__abc_52155_new_n17938_), .Y(u2__0remLo_451_0__232_));
OR2X2 OR2X2_4021 ( .A(u2__abc_52155_new_n17941_), .B(u2__abc_52155_new_n17942_), .Y(u2__abc_52155_new_n17943_));
OR2X2 OR2X2_4022 ( .A(u2__abc_52155_new_n17940_), .B(u2__abc_52155_new_n17944_), .Y(u2__0remLo_451_0__233_));
OR2X2 OR2X2_4023 ( .A(u2__abc_52155_new_n17949_), .B(u2__abc_52155_new_n17947_), .Y(u2__abc_52155_new_n17950_));
OR2X2 OR2X2_4024 ( .A(u2__abc_52155_new_n17946_), .B(u2__abc_52155_new_n17950_), .Y(u2__0remLo_451_0__234_));
OR2X2 OR2X2_4025 ( .A(u2__abc_52155_new_n17953_), .B(u2__abc_52155_new_n17954_), .Y(u2__abc_52155_new_n17955_));
OR2X2 OR2X2_4026 ( .A(u2__abc_52155_new_n17952_), .B(u2__abc_52155_new_n17956_), .Y(u2__0remLo_451_0__235_));
OR2X2 OR2X2_4027 ( .A(u2__abc_52155_new_n17959_), .B(u2__abc_52155_new_n17960_), .Y(u2__abc_52155_new_n17961_));
OR2X2 OR2X2_4028 ( .A(u2__abc_52155_new_n17958_), .B(u2__abc_52155_new_n17962_), .Y(u2__0remLo_451_0__236_));
OR2X2 OR2X2_4029 ( .A(u2__abc_52155_new_n17965_), .B(u2__abc_52155_new_n17966_), .Y(u2__abc_52155_new_n17967_));
OR2X2 OR2X2_403 ( .A(_abc_73687_new_n1170_), .B(\a[89] ), .Y(_abc_73687_new_n1435_));
OR2X2 OR2X2_4030 ( .A(u2__abc_52155_new_n17964_), .B(u2__abc_52155_new_n17968_), .Y(u2__0remLo_451_0__237_));
OR2X2 OR2X2_4031 ( .A(u2__abc_52155_new_n17971_), .B(u2__abc_52155_new_n17972_), .Y(u2__abc_52155_new_n17973_));
OR2X2 OR2X2_4032 ( .A(u2__abc_52155_new_n17970_), .B(u2__abc_52155_new_n17974_), .Y(u2__0remLo_451_0__238_));
OR2X2 OR2X2_4033 ( .A(u2__abc_52155_new_n17978_), .B(u2__abc_52155_new_n17977_), .Y(u2__abc_52155_new_n17979_));
OR2X2 OR2X2_4034 ( .A(u2__abc_52155_new_n17976_), .B(u2__abc_52155_new_n17980_), .Y(u2__0remLo_451_0__239_));
OR2X2 OR2X2_4035 ( .A(u2__abc_52155_new_n17982_), .B(u2__abc_52155_new_n17983_), .Y(u2__abc_52155_new_n17984_));
OR2X2 OR2X2_4036 ( .A(u2__abc_52155_new_n17986_), .B(u2__abc_52155_new_n17987_), .Y(u2__abc_52155_new_n17988_));
OR2X2 OR2X2_4037 ( .A(u2__abc_52155_new_n17985_), .B(u2__abc_52155_new_n17989_), .Y(u2__0remLo_451_0__240_));
OR2X2 OR2X2_4038 ( .A(u2__abc_52155_new_n17992_), .B(u2__abc_52155_new_n17993_), .Y(u2__abc_52155_new_n17994_));
OR2X2 OR2X2_4039 ( .A(u2__abc_52155_new_n17991_), .B(u2__abc_52155_new_n17995_), .Y(u2__0remLo_451_0__241_));
OR2X2 OR2X2_404 ( .A(\a[112] ), .B(\a[89] ), .Y(_abc_73687_new_n1437_));
OR2X2 OR2X2_4040 ( .A(u2__abc_52155_new_n17998_), .B(u2__abc_52155_new_n17999_), .Y(u2__abc_52155_new_n18000_));
OR2X2 OR2X2_4041 ( .A(u2__abc_52155_new_n17997_), .B(u2__abc_52155_new_n18001_), .Y(u2__0remLo_451_0__242_));
OR2X2 OR2X2_4042 ( .A(u2__abc_52155_new_n18005_), .B(u2__abc_52155_new_n18004_), .Y(u2__abc_52155_new_n18006_));
OR2X2 OR2X2_4043 ( .A(u2__abc_52155_new_n18003_), .B(u2__abc_52155_new_n18007_), .Y(u2__0remLo_451_0__243_));
OR2X2 OR2X2_4044 ( .A(u2__abc_52155_new_n18010_), .B(u2__abc_52155_new_n18011_), .Y(u2__abc_52155_new_n18012_));
OR2X2 OR2X2_4045 ( .A(u2__abc_52155_new_n18009_), .B(u2__abc_52155_new_n18013_), .Y(u2__0remLo_451_0__244_));
OR2X2 OR2X2_4046 ( .A(u2__abc_52155_new_n18016_), .B(u2__abc_52155_new_n18017_), .Y(u2__abc_52155_new_n18018_));
OR2X2 OR2X2_4047 ( .A(u2__abc_52155_new_n18015_), .B(u2__abc_52155_new_n18019_), .Y(u2__0remLo_451_0__245_));
OR2X2 OR2X2_4048 ( .A(u2__abc_52155_new_n18022_), .B(u2__abc_52155_new_n18023_), .Y(u2__abc_52155_new_n18024_));
OR2X2 OR2X2_4049 ( .A(u2__abc_52155_new_n18021_), .B(u2__abc_52155_new_n18025_), .Y(u2__0remLo_451_0__246_));
OR2X2 OR2X2_405 ( .A(_abc_73687_new_n1170_), .B(\a[90] ), .Y(_abc_73687_new_n1438_));
OR2X2 OR2X2_4050 ( .A(u2__abc_52155_new_n18028_), .B(u2__abc_52155_new_n18029_), .Y(u2__abc_52155_new_n18030_));
OR2X2 OR2X2_4051 ( .A(u2__abc_52155_new_n18027_), .B(u2__abc_52155_new_n18031_), .Y(u2__0remLo_451_0__247_));
OR2X2 OR2X2_4052 ( .A(u2__abc_52155_new_n18034_), .B(u2__abc_52155_new_n18035_), .Y(u2__abc_52155_new_n18036_));
OR2X2 OR2X2_4053 ( .A(u2__abc_52155_new_n18033_), .B(u2__abc_52155_new_n18037_), .Y(u2__0remLo_451_0__248_));
OR2X2 OR2X2_4054 ( .A(u2__abc_52155_new_n18041_), .B(u2__abc_52155_new_n18040_), .Y(u2__abc_52155_new_n18042_));
OR2X2 OR2X2_4055 ( .A(u2__abc_52155_new_n18039_), .B(u2__abc_52155_new_n18043_), .Y(u2__0remLo_451_0__249_));
OR2X2 OR2X2_4056 ( .A(u2__abc_52155_new_n18047_), .B(u2__abc_52155_new_n18046_), .Y(u2__abc_52155_new_n18048_));
OR2X2 OR2X2_4057 ( .A(u2__abc_52155_new_n18045_), .B(u2__abc_52155_new_n18049_), .Y(u2__0remLo_451_0__250_));
OR2X2 OR2X2_4058 ( .A(u2__abc_52155_new_n18052_), .B(u2__abc_52155_new_n18053_), .Y(u2__abc_52155_new_n18054_));
OR2X2 OR2X2_4059 ( .A(u2__abc_52155_new_n18051_), .B(u2__abc_52155_new_n18055_), .Y(u2__0remLo_451_0__251_));
OR2X2 OR2X2_406 ( .A(\a[112] ), .B(\a[90] ), .Y(_abc_73687_new_n1440_));
OR2X2 OR2X2_4060 ( .A(u2__abc_52155_new_n18058_), .B(u2__abc_52155_new_n18059_), .Y(u2__abc_52155_new_n18060_));
OR2X2 OR2X2_4061 ( .A(u2__abc_52155_new_n18057_), .B(u2__abc_52155_new_n18061_), .Y(u2__0remLo_451_0__252_));
OR2X2 OR2X2_4062 ( .A(u2__abc_52155_new_n18065_), .B(u2__abc_52155_new_n18064_), .Y(u2__abc_52155_new_n18066_));
OR2X2 OR2X2_4063 ( .A(u2__abc_52155_new_n18063_), .B(u2__abc_52155_new_n18067_), .Y(u2__0remLo_451_0__253_));
OR2X2 OR2X2_4064 ( .A(u2__abc_52155_new_n18070_), .B(u2__abc_52155_new_n18071_), .Y(u2__abc_52155_new_n18072_));
OR2X2 OR2X2_4065 ( .A(u2__abc_52155_new_n18069_), .B(u2__abc_52155_new_n18073_), .Y(u2__0remLo_451_0__254_));
OR2X2 OR2X2_4066 ( .A(u2__abc_52155_new_n18077_), .B(u2__abc_52155_new_n18076_), .Y(u2__abc_52155_new_n18078_));
OR2X2 OR2X2_4067 ( .A(u2__abc_52155_new_n18075_), .B(u2__abc_52155_new_n18079_), .Y(u2__0remLo_451_0__255_));
OR2X2 OR2X2_4068 ( .A(u2__abc_52155_new_n18084_), .B(u2__abc_52155_new_n18082_), .Y(u2__abc_52155_new_n18085_));
OR2X2 OR2X2_4069 ( .A(u2__abc_52155_new_n18081_), .B(u2__abc_52155_new_n18085_), .Y(u2__0remLo_451_0__256_));
OR2X2 OR2X2_407 ( .A(_abc_73687_new_n1170_), .B(\a[91] ), .Y(_abc_73687_new_n1441_));
OR2X2 OR2X2_4070 ( .A(u2__abc_52155_new_n18087_), .B(u2__abc_52155_new_n18088_), .Y(u2__abc_52155_new_n18089_));
OR2X2 OR2X2_4071 ( .A(u2__abc_52155_new_n18091_), .B(u2__abc_52155_new_n18092_), .Y(u2__abc_52155_new_n18093_));
OR2X2 OR2X2_4072 ( .A(u2__abc_52155_new_n18090_), .B(u2__abc_52155_new_n18094_), .Y(u2__0remLo_451_0__257_));
OR2X2 OR2X2_4073 ( .A(u2__abc_52155_new_n18096_), .B(u2__abc_52155_new_n18098_), .Y(u2__abc_52155_new_n18099_));
OR2X2 OR2X2_4074 ( .A(u2__abc_52155_new_n18101_), .B(u2__abc_52155_new_n18103_), .Y(u2__abc_52155_new_n18104_));
OR2X2 OR2X2_4075 ( .A(u2__abc_52155_new_n18106_), .B(u2__abc_52155_new_n18108_), .Y(u2__abc_52155_new_n18109_));
OR2X2 OR2X2_4076 ( .A(u2__abc_52155_new_n18111_), .B(u2__abc_52155_new_n18113_), .Y(u2__abc_52155_new_n18114_));
OR2X2 OR2X2_4077 ( .A(u2__abc_52155_new_n18116_), .B(u2__abc_52155_new_n18118_), .Y(u2__abc_52155_new_n18119_));
OR2X2 OR2X2_4078 ( .A(u2__abc_52155_new_n18121_), .B(u2__abc_52155_new_n18123_), .Y(u2__abc_52155_new_n18124_));
OR2X2 OR2X2_4079 ( .A(u2__abc_52155_new_n18126_), .B(u2__abc_52155_new_n18128_), .Y(u2__abc_52155_new_n18129_));
OR2X2 OR2X2_408 ( .A(\a[112] ), .B(\a[91] ), .Y(_abc_73687_new_n1443_));
OR2X2 OR2X2_4080 ( .A(u2__abc_52155_new_n18131_), .B(u2__abc_52155_new_n18133_), .Y(u2__abc_52155_new_n18134_));
OR2X2 OR2X2_4081 ( .A(u2__abc_52155_new_n18136_), .B(u2__abc_52155_new_n18138_), .Y(u2__abc_52155_new_n18139_));
OR2X2 OR2X2_4082 ( .A(u2__abc_52155_new_n18141_), .B(u2__abc_52155_new_n18143_), .Y(u2__abc_52155_new_n18144_));
OR2X2 OR2X2_4083 ( .A(u2__abc_52155_new_n18146_), .B(u2__abc_52155_new_n18148_), .Y(u2__abc_52155_new_n18149_));
OR2X2 OR2X2_4084 ( .A(u2__abc_52155_new_n18151_), .B(u2__abc_52155_new_n18153_), .Y(u2__abc_52155_new_n18154_));
OR2X2 OR2X2_4085 ( .A(u2__abc_52155_new_n18156_), .B(u2__abc_52155_new_n18158_), .Y(u2__abc_52155_new_n18159_));
OR2X2 OR2X2_4086 ( .A(u2__abc_52155_new_n18161_), .B(u2__abc_52155_new_n18163_), .Y(u2__abc_52155_new_n18164_));
OR2X2 OR2X2_4087 ( .A(u2__abc_52155_new_n18166_), .B(u2__abc_52155_new_n18168_), .Y(u2__abc_52155_new_n18169_));
OR2X2 OR2X2_4088 ( .A(u2__abc_52155_new_n18171_), .B(u2__abc_52155_new_n18173_), .Y(u2__abc_52155_new_n18174_));
OR2X2 OR2X2_4089 ( .A(u2__abc_52155_new_n18176_), .B(u2__abc_52155_new_n18178_), .Y(u2__abc_52155_new_n18179_));
OR2X2 OR2X2_409 ( .A(_abc_73687_new_n1170_), .B(\a[92] ), .Y(_abc_73687_new_n1444_));
OR2X2 OR2X2_4090 ( .A(u2__abc_52155_new_n18181_), .B(u2__abc_52155_new_n18183_), .Y(u2__abc_52155_new_n18184_));
OR2X2 OR2X2_4091 ( .A(u2__abc_52155_new_n18186_), .B(u2__abc_52155_new_n18188_), .Y(u2__abc_52155_new_n18189_));
OR2X2 OR2X2_4092 ( .A(u2__abc_52155_new_n18191_), .B(u2__abc_52155_new_n18193_), .Y(u2__abc_52155_new_n18194_));
OR2X2 OR2X2_4093 ( .A(u2__abc_52155_new_n18196_), .B(u2__abc_52155_new_n18198_), .Y(u2__abc_52155_new_n18199_));
OR2X2 OR2X2_4094 ( .A(u2__abc_52155_new_n18201_), .B(u2__abc_52155_new_n18203_), .Y(u2__abc_52155_new_n18204_));
OR2X2 OR2X2_4095 ( .A(u2__abc_52155_new_n18206_), .B(u2__abc_52155_new_n18208_), .Y(u2__abc_52155_new_n18209_));
OR2X2 OR2X2_4096 ( .A(u2__abc_52155_new_n18211_), .B(u2__abc_52155_new_n18213_), .Y(u2__abc_52155_new_n18214_));
OR2X2 OR2X2_4097 ( .A(u2__abc_52155_new_n18216_), .B(u2__abc_52155_new_n18218_), .Y(u2__abc_52155_new_n18219_));
OR2X2 OR2X2_4098 ( .A(u2__abc_52155_new_n18221_), .B(u2__abc_52155_new_n18223_), .Y(u2__abc_52155_new_n18224_));
OR2X2 OR2X2_4099 ( .A(u2__abc_52155_new_n18226_), .B(u2__abc_52155_new_n18228_), .Y(u2__abc_52155_new_n18229_));
OR2X2 OR2X2_41 ( .A(aNan), .B(sqrto_96_), .Y(_abc_73687_new_n890_));
OR2X2 OR2X2_410 ( .A(\a[112] ), .B(\a[92] ), .Y(_abc_73687_new_n1446_));
OR2X2 OR2X2_4100 ( .A(u2__abc_52155_new_n18231_), .B(u2__abc_52155_new_n18233_), .Y(u2__abc_52155_new_n18234_));
OR2X2 OR2X2_4101 ( .A(u2__abc_52155_new_n18236_), .B(u2__abc_52155_new_n18238_), .Y(u2__abc_52155_new_n18239_));
OR2X2 OR2X2_4102 ( .A(u2__abc_52155_new_n18241_), .B(u2__abc_52155_new_n18243_), .Y(u2__abc_52155_new_n18244_));
OR2X2 OR2X2_4103 ( .A(u2__abc_52155_new_n18246_), .B(u2__abc_52155_new_n18248_), .Y(u2__abc_52155_new_n18249_));
OR2X2 OR2X2_4104 ( .A(u2__abc_52155_new_n18251_), .B(u2__abc_52155_new_n18253_), .Y(u2__abc_52155_new_n18254_));
OR2X2 OR2X2_4105 ( .A(u2__abc_52155_new_n18256_), .B(u2__abc_52155_new_n18258_), .Y(u2__abc_52155_new_n18259_));
OR2X2 OR2X2_4106 ( .A(u2__abc_52155_new_n18261_), .B(u2__abc_52155_new_n18263_), .Y(u2__abc_52155_new_n18264_));
OR2X2 OR2X2_4107 ( .A(u2__abc_52155_new_n18266_), .B(u2__abc_52155_new_n18268_), .Y(u2__abc_52155_new_n18269_));
OR2X2 OR2X2_4108 ( .A(u2__abc_52155_new_n18271_), .B(u2__abc_52155_new_n18273_), .Y(u2__abc_52155_new_n18274_));
OR2X2 OR2X2_4109 ( .A(u2__abc_52155_new_n18276_), .B(u2__abc_52155_new_n18278_), .Y(u2__abc_52155_new_n18279_));
OR2X2 OR2X2_411 ( .A(_abc_73687_new_n1170_), .B(\a[93] ), .Y(_abc_73687_new_n1447_));
OR2X2 OR2X2_4110 ( .A(u2__abc_52155_new_n18281_), .B(u2__abc_52155_new_n18283_), .Y(u2__abc_52155_new_n18284_));
OR2X2 OR2X2_4111 ( .A(u2__abc_52155_new_n18286_), .B(u2__abc_52155_new_n18288_), .Y(u2__abc_52155_new_n18289_));
OR2X2 OR2X2_4112 ( .A(u2__abc_52155_new_n18291_), .B(u2__abc_52155_new_n18293_), .Y(u2__abc_52155_new_n18294_));
OR2X2 OR2X2_4113 ( .A(u2__abc_52155_new_n18296_), .B(u2__abc_52155_new_n18298_), .Y(u2__abc_52155_new_n18299_));
OR2X2 OR2X2_4114 ( .A(u2__abc_52155_new_n18301_), .B(u2__abc_52155_new_n18303_), .Y(u2__abc_52155_new_n18304_));
OR2X2 OR2X2_4115 ( .A(u2__abc_52155_new_n18306_), .B(u2__abc_52155_new_n18308_), .Y(u2__abc_52155_new_n18309_));
OR2X2 OR2X2_4116 ( .A(u2__abc_52155_new_n18311_), .B(u2__abc_52155_new_n18313_), .Y(u2__abc_52155_new_n18314_));
OR2X2 OR2X2_4117 ( .A(u2__abc_52155_new_n18316_), .B(u2__abc_52155_new_n18318_), .Y(u2__abc_52155_new_n18319_));
OR2X2 OR2X2_4118 ( .A(u2__abc_52155_new_n18321_), .B(u2__abc_52155_new_n18323_), .Y(u2__abc_52155_new_n18324_));
OR2X2 OR2X2_4119 ( .A(u2__abc_52155_new_n18326_), .B(u2__abc_52155_new_n18328_), .Y(u2__abc_52155_new_n18329_));
OR2X2 OR2X2_412 ( .A(\a[112] ), .B(\a[93] ), .Y(_abc_73687_new_n1449_));
OR2X2 OR2X2_4120 ( .A(u2__abc_52155_new_n18331_), .B(u2__abc_52155_new_n18333_), .Y(u2__abc_52155_new_n18334_));
OR2X2 OR2X2_4121 ( .A(u2__abc_52155_new_n18336_), .B(u2__abc_52155_new_n18338_), .Y(u2__abc_52155_new_n18339_));
OR2X2 OR2X2_4122 ( .A(u2__abc_52155_new_n18341_), .B(u2__abc_52155_new_n18343_), .Y(u2__abc_52155_new_n18344_));
OR2X2 OR2X2_4123 ( .A(u2__abc_52155_new_n18346_), .B(u2__abc_52155_new_n18348_), .Y(u2__abc_52155_new_n18349_));
OR2X2 OR2X2_4124 ( .A(u2__abc_52155_new_n18351_), .B(u2__abc_52155_new_n18353_), .Y(u2__abc_52155_new_n18354_));
OR2X2 OR2X2_4125 ( .A(u2__abc_52155_new_n18356_), .B(u2__abc_52155_new_n18358_), .Y(u2__abc_52155_new_n18359_));
OR2X2 OR2X2_4126 ( .A(u2__abc_52155_new_n18361_), .B(u2__abc_52155_new_n18363_), .Y(u2__abc_52155_new_n18364_));
OR2X2 OR2X2_4127 ( .A(u2__abc_52155_new_n18366_), .B(u2__abc_52155_new_n18368_), .Y(u2__abc_52155_new_n18369_));
OR2X2 OR2X2_4128 ( .A(u2__abc_52155_new_n18371_), .B(u2__abc_52155_new_n18373_), .Y(u2__abc_52155_new_n18374_));
OR2X2 OR2X2_4129 ( .A(u2__abc_52155_new_n18376_), .B(u2__abc_52155_new_n18378_), .Y(u2__abc_52155_new_n18379_));
OR2X2 OR2X2_413 ( .A(_abc_73687_new_n1170_), .B(\a[94] ), .Y(_abc_73687_new_n1450_));
OR2X2 OR2X2_4130 ( .A(u2__abc_52155_new_n18381_), .B(u2__abc_52155_new_n18383_), .Y(u2__abc_52155_new_n18384_));
OR2X2 OR2X2_4131 ( .A(u2__abc_52155_new_n18386_), .B(u2__abc_52155_new_n18388_), .Y(u2__abc_52155_new_n18389_));
OR2X2 OR2X2_4132 ( .A(u2__abc_52155_new_n18391_), .B(u2__abc_52155_new_n18393_), .Y(u2__abc_52155_new_n18394_));
OR2X2 OR2X2_4133 ( .A(u2__abc_52155_new_n18396_), .B(u2__abc_52155_new_n18398_), .Y(u2__abc_52155_new_n18399_));
OR2X2 OR2X2_4134 ( .A(u2__abc_52155_new_n18401_), .B(u2__abc_52155_new_n18403_), .Y(u2__abc_52155_new_n18404_));
OR2X2 OR2X2_4135 ( .A(u2__abc_52155_new_n18406_), .B(u2__abc_52155_new_n18408_), .Y(u2__abc_52155_new_n18409_));
OR2X2 OR2X2_4136 ( .A(u2__abc_52155_new_n18411_), .B(u2__abc_52155_new_n18413_), .Y(u2__abc_52155_new_n18414_));
OR2X2 OR2X2_4137 ( .A(u2__abc_52155_new_n18416_), .B(u2__abc_52155_new_n18418_), .Y(u2__abc_52155_new_n18419_));
OR2X2 OR2X2_4138 ( .A(u2__abc_52155_new_n18421_), .B(u2__abc_52155_new_n18423_), .Y(u2__abc_52155_new_n18424_));
OR2X2 OR2X2_4139 ( .A(u2__abc_52155_new_n18426_), .B(u2__abc_52155_new_n18428_), .Y(u2__abc_52155_new_n18429_));
OR2X2 OR2X2_414 ( .A(\a[112] ), .B(\a[94] ), .Y(_abc_73687_new_n1452_));
OR2X2 OR2X2_4140 ( .A(u2__abc_52155_new_n18431_), .B(u2__abc_52155_new_n18433_), .Y(u2__abc_52155_new_n18434_));
OR2X2 OR2X2_4141 ( .A(u2__abc_52155_new_n18436_), .B(u2__abc_52155_new_n18438_), .Y(u2__abc_52155_new_n18439_));
OR2X2 OR2X2_4142 ( .A(u2__abc_52155_new_n18441_), .B(u2__abc_52155_new_n18443_), .Y(u2__abc_52155_new_n18444_));
OR2X2 OR2X2_4143 ( .A(u2__abc_52155_new_n18446_), .B(u2__abc_52155_new_n18448_), .Y(u2__abc_52155_new_n18449_));
OR2X2 OR2X2_4144 ( .A(u2__abc_52155_new_n18451_), .B(u2__abc_52155_new_n18453_), .Y(u2__abc_52155_new_n18454_));
OR2X2 OR2X2_4145 ( .A(u2__abc_52155_new_n18456_), .B(u2__abc_52155_new_n18458_), .Y(u2__abc_52155_new_n18459_));
OR2X2 OR2X2_4146 ( .A(u2__abc_52155_new_n18461_), .B(u2__abc_52155_new_n18463_), .Y(u2__abc_52155_new_n18464_));
OR2X2 OR2X2_4147 ( .A(u2__abc_52155_new_n18466_), .B(u2__abc_52155_new_n18468_), .Y(u2__abc_52155_new_n18469_));
OR2X2 OR2X2_4148 ( .A(u2__abc_52155_new_n18471_), .B(u2__abc_52155_new_n18473_), .Y(u2__abc_52155_new_n18474_));
OR2X2 OR2X2_4149 ( .A(u2__abc_52155_new_n18476_), .B(u2__abc_52155_new_n18478_), .Y(u2__abc_52155_new_n18479_));
OR2X2 OR2X2_415 ( .A(_abc_73687_new_n1170_), .B(\a[95] ), .Y(_abc_73687_new_n1453_));
OR2X2 OR2X2_4150 ( .A(u2__abc_52155_new_n18481_), .B(u2__abc_52155_new_n18483_), .Y(u2__abc_52155_new_n18484_));
OR2X2 OR2X2_4151 ( .A(u2__abc_52155_new_n18486_), .B(u2__abc_52155_new_n18488_), .Y(u2__abc_52155_new_n18489_));
OR2X2 OR2X2_4152 ( .A(u2__abc_52155_new_n18491_), .B(u2__abc_52155_new_n18493_), .Y(u2__abc_52155_new_n18494_));
OR2X2 OR2X2_4153 ( .A(u2__abc_52155_new_n18496_), .B(u2__abc_52155_new_n18498_), .Y(u2__abc_52155_new_n18499_));
OR2X2 OR2X2_4154 ( .A(u2__abc_52155_new_n18501_), .B(u2__abc_52155_new_n18503_), .Y(u2__abc_52155_new_n18504_));
OR2X2 OR2X2_4155 ( .A(u2__abc_52155_new_n18506_), .B(u2__abc_52155_new_n18508_), .Y(u2__abc_52155_new_n18509_));
OR2X2 OR2X2_4156 ( .A(u2__abc_52155_new_n18511_), .B(u2__abc_52155_new_n18513_), .Y(u2__abc_52155_new_n18514_));
OR2X2 OR2X2_4157 ( .A(u2__abc_52155_new_n18516_), .B(u2__abc_52155_new_n18518_), .Y(u2__abc_52155_new_n18519_));
OR2X2 OR2X2_4158 ( .A(u2__abc_52155_new_n18521_), .B(u2__abc_52155_new_n18523_), .Y(u2__abc_52155_new_n18524_));
OR2X2 OR2X2_4159 ( .A(u2__abc_52155_new_n18526_), .B(u2__abc_52155_new_n18528_), .Y(u2__abc_52155_new_n18529_));
OR2X2 OR2X2_416 ( .A(\a[112] ), .B(\a[95] ), .Y(_abc_73687_new_n1455_));
OR2X2 OR2X2_4160 ( .A(u2__abc_52155_new_n18531_), .B(u2__abc_52155_new_n18533_), .Y(u2__abc_52155_new_n18534_));
OR2X2 OR2X2_4161 ( .A(u2__abc_52155_new_n18536_), .B(u2__abc_52155_new_n18538_), .Y(u2__abc_52155_new_n18539_));
OR2X2 OR2X2_4162 ( .A(u2__abc_52155_new_n18541_), .B(u2__abc_52155_new_n18543_), .Y(u2__abc_52155_new_n18544_));
OR2X2 OR2X2_4163 ( .A(u2__abc_52155_new_n18546_), .B(u2__abc_52155_new_n18548_), .Y(u2__abc_52155_new_n18549_));
OR2X2 OR2X2_4164 ( .A(u2__abc_52155_new_n18551_), .B(u2__abc_52155_new_n18553_), .Y(u2__abc_52155_new_n18554_));
OR2X2 OR2X2_4165 ( .A(u2__abc_52155_new_n18556_), .B(u2__abc_52155_new_n18558_), .Y(u2__abc_52155_new_n18559_));
OR2X2 OR2X2_4166 ( .A(u2__abc_52155_new_n18561_), .B(u2__abc_52155_new_n18563_), .Y(u2__abc_52155_new_n18564_));
OR2X2 OR2X2_4167 ( .A(u2__abc_52155_new_n18566_), .B(u2__abc_52155_new_n18568_), .Y(u2__abc_52155_new_n18569_));
OR2X2 OR2X2_4168 ( .A(u2__abc_52155_new_n18571_), .B(u2__abc_52155_new_n18573_), .Y(u2__abc_52155_new_n18574_));
OR2X2 OR2X2_4169 ( .A(u2__abc_52155_new_n18576_), .B(u2__abc_52155_new_n18578_), .Y(u2__abc_52155_new_n18579_));
OR2X2 OR2X2_417 ( .A(_abc_73687_new_n1170_), .B(\a[96] ), .Y(_abc_73687_new_n1456_));
OR2X2 OR2X2_4170 ( .A(u2__abc_52155_new_n18581_), .B(u2__abc_52155_new_n18583_), .Y(u2__abc_52155_new_n18584_));
OR2X2 OR2X2_4171 ( .A(u2__abc_52155_new_n18586_), .B(u2__abc_52155_new_n18588_), .Y(u2__abc_52155_new_n18589_));
OR2X2 OR2X2_4172 ( .A(u2__abc_52155_new_n18591_), .B(u2__abc_52155_new_n18593_), .Y(u2__abc_52155_new_n18594_));
OR2X2 OR2X2_4173 ( .A(u2__abc_52155_new_n18596_), .B(u2__abc_52155_new_n18598_), .Y(u2__abc_52155_new_n18599_));
OR2X2 OR2X2_4174 ( .A(u2__abc_52155_new_n18601_), .B(u2__abc_52155_new_n18603_), .Y(u2__abc_52155_new_n18604_));
OR2X2 OR2X2_4175 ( .A(u2__abc_52155_new_n18606_), .B(u2__abc_52155_new_n18608_), .Y(u2__abc_52155_new_n18609_));
OR2X2 OR2X2_4176 ( .A(u2__abc_52155_new_n18611_), .B(u2__abc_52155_new_n18613_), .Y(u2__abc_52155_new_n18614_));
OR2X2 OR2X2_4177 ( .A(u2__abc_52155_new_n18616_), .B(u2__abc_52155_new_n18618_), .Y(u2__abc_52155_new_n18619_));
OR2X2 OR2X2_4178 ( .A(u2__abc_52155_new_n18621_), .B(u2__abc_52155_new_n18623_), .Y(u2__abc_52155_new_n18624_));
OR2X2 OR2X2_4179 ( .A(u2__abc_52155_new_n18626_), .B(u2__abc_52155_new_n18628_), .Y(u2__abc_52155_new_n18629_));
OR2X2 OR2X2_418 ( .A(\a[112] ), .B(\a[96] ), .Y(_abc_73687_new_n1458_));
OR2X2 OR2X2_4180 ( .A(u2__abc_52155_new_n18631_), .B(u2__abc_52155_new_n18633_), .Y(u2__abc_52155_new_n18634_));
OR2X2 OR2X2_4181 ( .A(u2__abc_52155_new_n18636_), .B(u2__abc_52155_new_n18638_), .Y(u2__abc_52155_new_n18639_));
OR2X2 OR2X2_4182 ( .A(u2__abc_52155_new_n18641_), .B(u2__abc_52155_new_n18643_), .Y(u2__abc_52155_new_n18644_));
OR2X2 OR2X2_4183 ( .A(u2__abc_52155_new_n18646_), .B(u2__abc_52155_new_n18648_), .Y(u2__abc_52155_new_n18649_));
OR2X2 OR2X2_4184 ( .A(u2__abc_52155_new_n18651_), .B(u2__abc_52155_new_n18653_), .Y(u2__abc_52155_new_n18654_));
OR2X2 OR2X2_4185 ( .A(u2__abc_52155_new_n18656_), .B(u2__abc_52155_new_n18658_), .Y(u2__abc_52155_new_n18659_));
OR2X2 OR2X2_4186 ( .A(u2__abc_52155_new_n18661_), .B(u2__abc_52155_new_n18663_), .Y(u2__abc_52155_new_n18664_));
OR2X2 OR2X2_4187 ( .A(u2__abc_52155_new_n18666_), .B(u2__abc_52155_new_n18668_), .Y(u2__abc_52155_new_n18669_));
OR2X2 OR2X2_4188 ( .A(u2__abc_52155_new_n18671_), .B(u2__abc_52155_new_n18673_), .Y(u2__abc_52155_new_n18674_));
OR2X2 OR2X2_4189 ( .A(u2__abc_52155_new_n18676_), .B(u2__abc_52155_new_n18678_), .Y(u2__abc_52155_new_n18679_));
OR2X2 OR2X2_419 ( .A(_abc_73687_new_n1170_), .B(\a[97] ), .Y(_abc_73687_new_n1459_));
OR2X2 OR2X2_4190 ( .A(u2__abc_52155_new_n18681_), .B(u2__abc_52155_new_n18683_), .Y(u2__abc_52155_new_n18684_));
OR2X2 OR2X2_4191 ( .A(u2__abc_52155_new_n18686_), .B(u2__abc_52155_new_n18688_), .Y(u2__abc_52155_new_n18689_));
OR2X2 OR2X2_4192 ( .A(u2__abc_52155_new_n18691_), .B(u2__abc_52155_new_n18693_), .Y(u2__abc_52155_new_n18694_));
OR2X2 OR2X2_4193 ( .A(u2__abc_52155_new_n18696_), .B(u2__abc_52155_new_n18698_), .Y(u2__abc_52155_new_n18699_));
OR2X2 OR2X2_4194 ( .A(u2__abc_52155_new_n18701_), .B(u2__abc_52155_new_n18703_), .Y(u2__abc_52155_new_n18704_));
OR2X2 OR2X2_4195 ( .A(u2__abc_52155_new_n18706_), .B(u2__abc_52155_new_n18708_), .Y(u2__abc_52155_new_n18709_));
OR2X2 OR2X2_4196 ( .A(u2__abc_52155_new_n18711_), .B(u2__abc_52155_new_n18713_), .Y(u2__abc_52155_new_n18714_));
OR2X2 OR2X2_4197 ( .A(u2__abc_52155_new_n18716_), .B(u2__abc_52155_new_n18718_), .Y(u2__abc_52155_new_n18719_));
OR2X2 OR2X2_4198 ( .A(u2__abc_52155_new_n18721_), .B(u2__abc_52155_new_n18723_), .Y(u2__abc_52155_new_n18724_));
OR2X2 OR2X2_4199 ( .A(u2__abc_52155_new_n18726_), .B(u2__abc_52155_new_n18728_), .Y(u2__abc_52155_new_n18729_));
OR2X2 OR2X2_42 ( .A(_abc_73687_new_n753_), .B(\a[20] ), .Y(_abc_73687_new_n891_));
OR2X2 OR2X2_420 ( .A(\a[112] ), .B(\a[97] ), .Y(_abc_73687_new_n1461_));
OR2X2 OR2X2_4200 ( .A(u2__abc_52155_new_n18731_), .B(u2__abc_52155_new_n18733_), .Y(u2__abc_52155_new_n18734_));
OR2X2 OR2X2_4201 ( .A(u2__abc_52155_new_n18736_), .B(u2__abc_52155_new_n18738_), .Y(u2__abc_52155_new_n18739_));
OR2X2 OR2X2_4202 ( .A(u2__abc_52155_new_n18741_), .B(u2__abc_52155_new_n18743_), .Y(u2__abc_52155_new_n18744_));
OR2X2 OR2X2_4203 ( .A(u2__abc_52155_new_n18746_), .B(u2__abc_52155_new_n18748_), .Y(u2__abc_52155_new_n18749_));
OR2X2 OR2X2_4204 ( .A(u2__abc_52155_new_n18751_), .B(u2__abc_52155_new_n18753_), .Y(u2__abc_52155_new_n18754_));
OR2X2 OR2X2_4205 ( .A(u2__abc_52155_new_n18756_), .B(u2__abc_52155_new_n18758_), .Y(u2__abc_52155_new_n18759_));
OR2X2 OR2X2_4206 ( .A(u2__abc_52155_new_n18761_), .B(u2__abc_52155_new_n18763_), .Y(u2__abc_52155_new_n18764_));
OR2X2 OR2X2_4207 ( .A(u2__abc_52155_new_n18766_), .B(u2__abc_52155_new_n18768_), .Y(u2__abc_52155_new_n18769_));
OR2X2 OR2X2_4208 ( .A(u2__abc_52155_new_n18771_), .B(u2__abc_52155_new_n18773_), .Y(u2__abc_52155_new_n18774_));
OR2X2 OR2X2_4209 ( .A(u2__abc_52155_new_n18776_), .B(u2__abc_52155_new_n18778_), .Y(u2__abc_52155_new_n18779_));
OR2X2 OR2X2_421 ( .A(_abc_73687_new_n1170_), .B(\a[98] ), .Y(_abc_73687_new_n1462_));
OR2X2 OR2X2_4210 ( .A(u2__abc_52155_new_n18781_), .B(u2__abc_52155_new_n18783_), .Y(u2__abc_52155_new_n18784_));
OR2X2 OR2X2_4211 ( .A(u2__abc_52155_new_n18786_), .B(u2__abc_52155_new_n18788_), .Y(u2__abc_52155_new_n18789_));
OR2X2 OR2X2_4212 ( .A(u2__abc_52155_new_n18791_), .B(u2__abc_52155_new_n18793_), .Y(u2__abc_52155_new_n18794_));
OR2X2 OR2X2_4213 ( .A(u2__abc_52155_new_n18796_), .B(u2__abc_52155_new_n18798_), .Y(u2__abc_52155_new_n18799_));
OR2X2 OR2X2_4214 ( .A(u2__abc_52155_new_n18801_), .B(u2__abc_52155_new_n18803_), .Y(u2__abc_52155_new_n18804_));
OR2X2 OR2X2_4215 ( .A(u2__abc_52155_new_n18806_), .B(u2__abc_52155_new_n18808_), .Y(u2__abc_52155_new_n18809_));
OR2X2 OR2X2_4216 ( .A(u2__abc_52155_new_n18811_), .B(u2__abc_52155_new_n18813_), .Y(u2__abc_52155_new_n18814_));
OR2X2 OR2X2_4217 ( .A(u2__abc_52155_new_n18816_), .B(u2__abc_52155_new_n18818_), .Y(u2__abc_52155_new_n18819_));
OR2X2 OR2X2_4218 ( .A(u2__abc_52155_new_n18821_), .B(u2__abc_52155_new_n18823_), .Y(u2__abc_52155_new_n18824_));
OR2X2 OR2X2_4219 ( .A(u2__abc_52155_new_n18826_), .B(u2__abc_52155_new_n18828_), .Y(u2__abc_52155_new_n18829_));
OR2X2 OR2X2_422 ( .A(\a[112] ), .B(\a[98] ), .Y(_abc_73687_new_n1464_));
OR2X2 OR2X2_4220 ( .A(u2__abc_52155_new_n18831_), .B(u2__abc_52155_new_n18833_), .Y(u2__abc_52155_new_n18834_));
OR2X2 OR2X2_4221 ( .A(u2__abc_52155_new_n18836_), .B(u2__abc_52155_new_n18838_), .Y(u2__abc_52155_new_n18839_));
OR2X2 OR2X2_4222 ( .A(u2__abc_52155_new_n18841_), .B(u2__abc_52155_new_n18843_), .Y(u2__abc_52155_new_n18844_));
OR2X2 OR2X2_4223 ( .A(u2__abc_52155_new_n18846_), .B(u2__abc_52155_new_n18848_), .Y(u2__abc_52155_new_n18849_));
OR2X2 OR2X2_4224 ( .A(u2__abc_52155_new_n18851_), .B(u2__abc_52155_new_n18853_), .Y(u2__abc_52155_new_n18854_));
OR2X2 OR2X2_4225 ( .A(u2__abc_52155_new_n18856_), .B(u2__abc_52155_new_n18858_), .Y(u2__abc_52155_new_n18859_));
OR2X2 OR2X2_4226 ( .A(u2__abc_52155_new_n18861_), .B(u2__abc_52155_new_n18863_), .Y(u2__abc_52155_new_n18864_));
OR2X2 OR2X2_4227 ( .A(u2__abc_52155_new_n18866_), .B(u2__abc_52155_new_n18868_), .Y(u2__abc_52155_new_n18869_));
OR2X2 OR2X2_4228 ( .A(u2__abc_52155_new_n18871_), .B(u2__abc_52155_new_n18873_), .Y(u2__abc_52155_new_n18874_));
OR2X2 OR2X2_4229 ( .A(u2__abc_52155_new_n18876_), .B(u2__abc_52155_new_n18878_), .Y(u2__abc_52155_new_n18879_));
OR2X2 OR2X2_423 ( .A(_abc_73687_new_n1170_), .B(\a[99] ), .Y(_abc_73687_new_n1465_));
OR2X2 OR2X2_4230 ( .A(u2__abc_52155_new_n18881_), .B(u2__abc_52155_new_n18883_), .Y(u2__abc_52155_new_n18884_));
OR2X2 OR2X2_4231 ( .A(u2__abc_52155_new_n18886_), .B(u2__abc_52155_new_n18888_), .Y(u2__abc_52155_new_n18889_));
OR2X2 OR2X2_4232 ( .A(u2__abc_52155_new_n18891_), .B(u2__abc_52155_new_n18893_), .Y(u2__abc_52155_new_n18894_));
OR2X2 OR2X2_4233 ( .A(u2__abc_52155_new_n18896_), .B(u2__abc_52155_new_n18898_), .Y(u2__abc_52155_new_n18899_));
OR2X2 OR2X2_4234 ( .A(u2__abc_52155_new_n18901_), .B(u2__abc_52155_new_n18903_), .Y(u2__abc_52155_new_n18904_));
OR2X2 OR2X2_4235 ( .A(u2__abc_52155_new_n18906_), .B(u2__abc_52155_new_n18908_), .Y(u2__abc_52155_new_n18909_));
OR2X2 OR2X2_4236 ( .A(u2__abc_52155_new_n18911_), .B(u2__abc_52155_new_n18913_), .Y(u2__abc_52155_new_n18914_));
OR2X2 OR2X2_4237 ( .A(u2__abc_52155_new_n18916_), .B(u2__abc_52155_new_n18918_), .Y(u2__abc_52155_new_n18919_));
OR2X2 OR2X2_4238 ( .A(u2__abc_52155_new_n18921_), .B(u2__abc_52155_new_n18923_), .Y(u2__abc_52155_new_n18924_));
OR2X2 OR2X2_4239 ( .A(u2__abc_52155_new_n18926_), .B(u2__abc_52155_new_n18928_), .Y(u2__abc_52155_new_n18929_));
OR2X2 OR2X2_424 ( .A(\a[112] ), .B(\a[99] ), .Y(_abc_73687_new_n1467_));
OR2X2 OR2X2_4240 ( .A(u2__abc_52155_new_n18931_), .B(u2__abc_52155_new_n18933_), .Y(u2__abc_52155_new_n18934_));
OR2X2 OR2X2_4241 ( .A(u2__abc_52155_new_n18936_), .B(u2__abc_52155_new_n18938_), .Y(u2__abc_52155_new_n18939_));
OR2X2 OR2X2_4242 ( .A(u2__abc_52155_new_n18941_), .B(u2__abc_52155_new_n18943_), .Y(u2__abc_52155_new_n18944_));
OR2X2 OR2X2_4243 ( .A(u2__abc_52155_new_n18946_), .B(u2__abc_52155_new_n18948_), .Y(u2__abc_52155_new_n18949_));
OR2X2 OR2X2_4244 ( .A(u2__abc_52155_new_n18951_), .B(u2__abc_52155_new_n18953_), .Y(u2__abc_52155_new_n18954_));
OR2X2 OR2X2_4245 ( .A(u2__abc_52155_new_n18956_), .B(u2__abc_52155_new_n18958_), .Y(u2__abc_52155_new_n18959_));
OR2X2 OR2X2_4246 ( .A(u2__abc_52155_new_n18961_), .B(u2__abc_52155_new_n18963_), .Y(u2__abc_52155_new_n18964_));
OR2X2 OR2X2_4247 ( .A(u2__abc_52155_new_n18966_), .B(u2__abc_52155_new_n18968_), .Y(u2__abc_52155_new_n18969_));
OR2X2 OR2X2_4248 ( .A(u2__abc_52155_new_n18971_), .B(u2__abc_52155_new_n18973_), .Y(u2__abc_52155_new_n18974_));
OR2X2 OR2X2_4249 ( .A(u2__abc_52155_new_n18976_), .B(u2__abc_52155_new_n18978_), .Y(u2__abc_52155_new_n18979_));
OR2X2 OR2X2_425 ( .A(_abc_73687_new_n1170_), .B(\a[100] ), .Y(_abc_73687_new_n1468_));
OR2X2 OR2X2_4250 ( .A(u2__abc_52155_new_n18981_), .B(u2__abc_52155_new_n18983_), .Y(u2__abc_52155_new_n18984_));
OR2X2 OR2X2_4251 ( .A(u2__abc_52155_new_n18986_), .B(u2__abc_52155_new_n18988_), .Y(u2__abc_52155_new_n18989_));
OR2X2 OR2X2_4252 ( .A(u2__abc_52155_new_n18991_), .B(u2__abc_52155_new_n18993_), .Y(u2__abc_52155_new_n18994_));
OR2X2 OR2X2_4253 ( .A(u2__abc_52155_new_n18996_), .B(u2__abc_52155_new_n18998_), .Y(u2__abc_52155_new_n18999_));
OR2X2 OR2X2_4254 ( .A(u2__abc_52155_new_n19001_), .B(u2__abc_52155_new_n19003_), .Y(u2__abc_52155_new_n19004_));
OR2X2 OR2X2_4255 ( .A(u2__abc_52155_new_n19006_), .B(u2__abc_52155_new_n19008_), .Y(u2__abc_52155_new_n19009_));
OR2X2 OR2X2_4256 ( .A(u2__abc_52155_new_n19011_), .B(u2__abc_52155_new_n19013_), .Y(u2__abc_52155_new_n19014_));
OR2X2 OR2X2_4257 ( .A(u2__abc_52155_new_n19016_), .B(u2__abc_52155_new_n19018_), .Y(u2__abc_52155_new_n19019_));
OR2X2 OR2X2_4258 ( .A(u2__abc_52155_new_n19021_), .B(u2__abc_52155_new_n19023_), .Y(u2__abc_52155_new_n19024_));
OR2X2 OR2X2_4259 ( .A(u2__abc_52155_new_n19026_), .B(u2__abc_52155_new_n19028_), .Y(u2__abc_52155_new_n19029_));
OR2X2 OR2X2_426 ( .A(\a[112] ), .B(\a[100] ), .Y(_abc_73687_new_n1470_));
OR2X2 OR2X2_4260 ( .A(u2__abc_52155_new_n19031_), .B(u2__abc_52155_new_n19033_), .Y(u2__abc_52155_new_n19034_));
OR2X2 OR2X2_4261 ( .A(u2__abc_52155_new_n19036_), .B(u2__abc_52155_new_n19038_), .Y(u2__abc_52155_new_n19039_));
OR2X2 OR2X2_4262 ( .A(u2__abc_52155_new_n19041_), .B(u2__abc_52155_new_n19043_), .Y(u2__abc_52155_new_n19044_));
OR2X2 OR2X2_4263 ( .A(u2__abc_52155_new_n19046_), .B(u2__abc_52155_new_n19048_), .Y(u2__abc_52155_new_n19049_));
OR2X2 OR2X2_4264 ( .A(u2__abc_52155_new_n19051_), .B(u2__abc_52155_new_n19053_), .Y(u2__abc_52155_new_n19054_));
OR2X2 OR2X2_4265 ( .A(u2__abc_52155_new_n19056_), .B(u2__abc_52155_new_n19058_), .Y(u2__abc_52155_new_n19059_));
OR2X2 OR2X2_4266 ( .A(u2__abc_52155_new_n19061_), .B(u2__abc_52155_new_n19063_), .Y(u2__abc_52155_new_n19064_));
OR2X2 OR2X2_4267 ( .A(u2__abc_52155_new_n7622_), .B(u2_root_0_), .Y(u2__abc_52155_new_n19071_));
OR2X2 OR2X2_4268 ( .A(u2__abc_52155_new_n19072_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19073_));
OR2X2 OR2X2_4269 ( .A(u2__abc_52155_new_n19077_), .B(u2__abc_52155_new_n19068_), .Y(u2__abc_52155_new_n19078_));
OR2X2 OR2X2_427 ( .A(_abc_73687_new_n1170_), .B(\a[101] ), .Y(_abc_73687_new_n1471_));
OR2X2 OR2X2_4270 ( .A(u2__abc_52155_new_n19069_), .B(sqrto_0_), .Y(u2__abc_52155_new_n19083_));
OR2X2 OR2X2_4271 ( .A(u2__abc_52155_new_n19084_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19085_));
OR2X2 OR2X2_4272 ( .A(u2__abc_52155_new_n19089_), .B(u2__abc_52155_new_n19080_), .Y(u2__abc_52155_new_n19090_));
OR2X2 OR2X2_4273 ( .A(u2__abc_52155_new_n19081_), .B(sqrto_1_), .Y(u2__abc_52155_new_n19093_));
OR2X2 OR2X2_4274 ( .A(u2__abc_52155_new_n19096_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19097_));
OR2X2 OR2X2_4275 ( .A(u2__abc_52155_new_n19101_), .B(u2__abc_52155_new_n19092_), .Y(u2__abc_52155_new_n19102_));
OR2X2 OR2X2_4276 ( .A(u2__abc_52155_new_n19094_), .B(sqrto_2_), .Y(u2__abc_52155_new_n19105_));
OR2X2 OR2X2_4277 ( .A(u2__abc_52155_new_n19108_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19109_));
OR2X2 OR2X2_4278 ( .A(u2__abc_52155_new_n19113_), .B(u2__abc_52155_new_n19104_), .Y(u2__abc_52155_new_n19114_));
OR2X2 OR2X2_4279 ( .A(u2__abc_52155_new_n19106_), .B(sqrto_3_), .Y(u2__abc_52155_new_n19117_));
OR2X2 OR2X2_428 ( .A(\a[112] ), .B(\a[101] ), .Y(_abc_73687_new_n1473_));
OR2X2 OR2X2_4280 ( .A(u2__abc_52155_new_n19120_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19121_));
OR2X2 OR2X2_4281 ( .A(u2__abc_52155_new_n19125_), .B(u2__abc_52155_new_n19116_), .Y(u2__abc_52155_new_n19126_));
OR2X2 OR2X2_4282 ( .A(u2__abc_52155_new_n19118_), .B(sqrto_4_), .Y(u2__abc_52155_new_n19129_));
OR2X2 OR2X2_4283 ( .A(u2__abc_52155_new_n19132_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19133_));
OR2X2 OR2X2_4284 ( .A(u2__abc_52155_new_n19137_), .B(u2__abc_52155_new_n19128_), .Y(u2__abc_52155_new_n19138_));
OR2X2 OR2X2_4285 ( .A(u2__abc_52155_new_n19130_), .B(sqrto_5_), .Y(u2__abc_52155_new_n19141_));
OR2X2 OR2X2_4286 ( .A(u2__abc_52155_new_n19144_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19145_));
OR2X2 OR2X2_4287 ( .A(u2__abc_52155_new_n19149_), .B(u2__abc_52155_new_n19140_), .Y(u2__abc_52155_new_n19150_));
OR2X2 OR2X2_4288 ( .A(u2__abc_52155_new_n19142_), .B(sqrto_6_), .Y(u2__abc_52155_new_n19153_));
OR2X2 OR2X2_4289 ( .A(u2__abc_52155_new_n19156_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19157_));
OR2X2 OR2X2_429 ( .A(_abc_73687_new_n1170_), .B(\a[102] ), .Y(_abc_73687_new_n1474_));
OR2X2 OR2X2_4290 ( .A(u2__abc_52155_new_n19161_), .B(u2__abc_52155_new_n19152_), .Y(u2__abc_52155_new_n19162_));
OR2X2 OR2X2_4291 ( .A(u2__abc_52155_new_n19154_), .B(sqrto_7_), .Y(u2__abc_52155_new_n19165_));
OR2X2 OR2X2_4292 ( .A(u2__abc_52155_new_n19168_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19169_));
OR2X2 OR2X2_4293 ( .A(u2__abc_52155_new_n19173_), .B(u2__abc_52155_new_n19164_), .Y(u2__abc_52155_new_n19174_));
OR2X2 OR2X2_4294 ( .A(u2__abc_52155_new_n19166_), .B(sqrto_8_), .Y(u2__abc_52155_new_n19177_));
OR2X2 OR2X2_4295 ( .A(u2__abc_52155_new_n19180_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19181_));
OR2X2 OR2X2_4296 ( .A(u2__abc_52155_new_n19185_), .B(u2__abc_52155_new_n19176_), .Y(u2__abc_52155_new_n19186_));
OR2X2 OR2X2_4297 ( .A(u2__abc_52155_new_n19178_), .B(sqrto_9_), .Y(u2__abc_52155_new_n19189_));
OR2X2 OR2X2_4298 ( .A(u2__abc_52155_new_n19192_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19193_));
OR2X2 OR2X2_4299 ( .A(u2__abc_52155_new_n19197_), .B(u2__abc_52155_new_n19188_), .Y(u2__abc_52155_new_n19198_));
OR2X2 OR2X2_43 ( .A(aNan), .B(sqrto_97_), .Y(_abc_73687_new_n893_));
OR2X2 OR2X2_430 ( .A(\a[112] ), .B(\a[102] ), .Y(_abc_73687_new_n1476_));
OR2X2 OR2X2_4300 ( .A(u2__abc_52155_new_n19190_), .B(sqrto_10_), .Y(u2__abc_52155_new_n19201_));
OR2X2 OR2X2_4301 ( .A(u2__abc_52155_new_n19204_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19205_));
OR2X2 OR2X2_4302 ( .A(u2__abc_52155_new_n19209_), .B(u2__abc_52155_new_n19200_), .Y(u2__abc_52155_new_n19210_));
OR2X2 OR2X2_4303 ( .A(u2__abc_52155_new_n19202_), .B(sqrto_11_), .Y(u2__abc_52155_new_n19213_));
OR2X2 OR2X2_4304 ( .A(u2__abc_52155_new_n19216_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19217_));
OR2X2 OR2X2_4305 ( .A(u2__abc_52155_new_n19221_), .B(u2__abc_52155_new_n19212_), .Y(u2__abc_52155_new_n19222_));
OR2X2 OR2X2_4306 ( .A(u2__abc_52155_new_n19214_), .B(sqrto_12_), .Y(u2__abc_52155_new_n19225_));
OR2X2 OR2X2_4307 ( .A(u2__abc_52155_new_n19228_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19229_));
OR2X2 OR2X2_4308 ( .A(u2__abc_52155_new_n19233_), .B(u2__abc_52155_new_n19224_), .Y(u2__abc_52155_new_n19234_));
OR2X2 OR2X2_4309 ( .A(u2__abc_52155_new_n19226_), .B(sqrto_13_), .Y(u2__abc_52155_new_n19237_));
OR2X2 OR2X2_431 ( .A(_abc_73687_new_n1170_), .B(\a[103] ), .Y(_abc_73687_new_n1477_));
OR2X2 OR2X2_4310 ( .A(u2__abc_52155_new_n19240_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19241_));
OR2X2 OR2X2_4311 ( .A(u2__abc_52155_new_n19245_), .B(u2__abc_52155_new_n19236_), .Y(u2__abc_52155_new_n19246_));
OR2X2 OR2X2_4312 ( .A(u2__abc_52155_new_n19238_), .B(sqrto_14_), .Y(u2__abc_52155_new_n19249_));
OR2X2 OR2X2_4313 ( .A(u2__abc_52155_new_n19252_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19253_));
OR2X2 OR2X2_4314 ( .A(u2__abc_52155_new_n19257_), .B(u2__abc_52155_new_n19248_), .Y(u2__abc_52155_new_n19258_));
OR2X2 OR2X2_4315 ( .A(u2__abc_52155_new_n19250_), .B(sqrto_15_), .Y(u2__abc_52155_new_n19261_));
OR2X2 OR2X2_4316 ( .A(u2__abc_52155_new_n19264_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19265_));
OR2X2 OR2X2_4317 ( .A(u2__abc_52155_new_n19269_), .B(u2__abc_52155_new_n19260_), .Y(u2__abc_52155_new_n19270_));
OR2X2 OR2X2_4318 ( .A(u2__abc_52155_new_n19262_), .B(sqrto_16_), .Y(u2__abc_52155_new_n19273_));
OR2X2 OR2X2_4319 ( .A(u2__abc_52155_new_n19276_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19277_));
OR2X2 OR2X2_432 ( .A(\a[112] ), .B(\a[103] ), .Y(_abc_73687_new_n1479_));
OR2X2 OR2X2_4320 ( .A(u2__abc_52155_new_n19281_), .B(u2__abc_52155_new_n19272_), .Y(u2__abc_52155_new_n19282_));
OR2X2 OR2X2_4321 ( .A(u2__abc_52155_new_n19274_), .B(sqrto_17_), .Y(u2__abc_52155_new_n19285_));
OR2X2 OR2X2_4322 ( .A(u2__abc_52155_new_n19288_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19289_));
OR2X2 OR2X2_4323 ( .A(u2__abc_52155_new_n19293_), .B(u2__abc_52155_new_n19284_), .Y(u2__abc_52155_new_n19294_));
OR2X2 OR2X2_4324 ( .A(u2__abc_52155_new_n19286_), .B(sqrto_18_), .Y(u2__abc_52155_new_n19297_));
OR2X2 OR2X2_4325 ( .A(u2__abc_52155_new_n19300_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19301_));
OR2X2 OR2X2_4326 ( .A(u2__abc_52155_new_n19305_), .B(u2__abc_52155_new_n19296_), .Y(u2__abc_52155_new_n19306_));
OR2X2 OR2X2_4327 ( .A(u2__abc_52155_new_n19298_), .B(sqrto_19_), .Y(u2__abc_52155_new_n19309_));
OR2X2 OR2X2_4328 ( .A(u2__abc_52155_new_n19312_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19313_));
OR2X2 OR2X2_4329 ( .A(u2__abc_52155_new_n19317_), .B(u2__abc_52155_new_n19308_), .Y(u2__abc_52155_new_n19318_));
OR2X2 OR2X2_433 ( .A(_abc_73687_new_n1170_), .B(\a[104] ), .Y(_abc_73687_new_n1480_));
OR2X2 OR2X2_4330 ( .A(u2__abc_52155_new_n19310_), .B(sqrto_20_), .Y(u2__abc_52155_new_n19321_));
OR2X2 OR2X2_4331 ( .A(u2__abc_52155_new_n19324_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19325_));
OR2X2 OR2X2_4332 ( .A(u2__abc_52155_new_n19329_), .B(u2__abc_52155_new_n19320_), .Y(u2__abc_52155_new_n19330_));
OR2X2 OR2X2_4333 ( .A(u2__abc_52155_new_n19322_), .B(sqrto_21_), .Y(u2__abc_52155_new_n19333_));
OR2X2 OR2X2_4334 ( .A(u2__abc_52155_new_n19336_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19337_));
OR2X2 OR2X2_4335 ( .A(u2__abc_52155_new_n19341_), .B(u2__abc_52155_new_n19332_), .Y(u2__abc_52155_new_n19342_));
OR2X2 OR2X2_4336 ( .A(u2__abc_52155_new_n19334_), .B(sqrto_22_), .Y(u2__abc_52155_new_n19345_));
OR2X2 OR2X2_4337 ( .A(u2__abc_52155_new_n19348_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19349_));
OR2X2 OR2X2_4338 ( .A(u2__abc_52155_new_n19353_), .B(u2__abc_52155_new_n19344_), .Y(u2__abc_52155_new_n19354_));
OR2X2 OR2X2_4339 ( .A(u2__abc_52155_new_n19346_), .B(sqrto_23_), .Y(u2__abc_52155_new_n19357_));
OR2X2 OR2X2_434 ( .A(\a[112] ), .B(\a[104] ), .Y(_abc_73687_new_n1482_));
OR2X2 OR2X2_4340 ( .A(u2__abc_52155_new_n19360_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19361_));
OR2X2 OR2X2_4341 ( .A(u2__abc_52155_new_n19365_), .B(u2__abc_52155_new_n19356_), .Y(u2__abc_52155_new_n19366_));
OR2X2 OR2X2_4342 ( .A(u2__abc_52155_new_n19358_), .B(sqrto_24_), .Y(u2__abc_52155_new_n19369_));
OR2X2 OR2X2_4343 ( .A(u2__abc_52155_new_n19372_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19373_));
OR2X2 OR2X2_4344 ( .A(u2__abc_52155_new_n19377_), .B(u2__abc_52155_new_n19368_), .Y(u2__abc_52155_new_n19378_));
OR2X2 OR2X2_4345 ( .A(u2__abc_52155_new_n19370_), .B(sqrto_25_), .Y(u2__abc_52155_new_n19381_));
OR2X2 OR2X2_4346 ( .A(u2__abc_52155_new_n19384_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19385_));
OR2X2 OR2X2_4347 ( .A(u2__abc_52155_new_n19389_), .B(u2__abc_52155_new_n19380_), .Y(u2__abc_52155_new_n19390_));
OR2X2 OR2X2_4348 ( .A(u2__abc_52155_new_n19382_), .B(sqrto_26_), .Y(u2__abc_52155_new_n19393_));
OR2X2 OR2X2_4349 ( .A(u2__abc_52155_new_n19396_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19397_));
OR2X2 OR2X2_435 ( .A(_abc_73687_new_n1170_), .B(\a[105] ), .Y(_abc_73687_new_n1483_));
OR2X2 OR2X2_4350 ( .A(u2__abc_52155_new_n19401_), .B(u2__abc_52155_new_n19392_), .Y(u2__abc_52155_new_n19402_));
OR2X2 OR2X2_4351 ( .A(u2__abc_52155_new_n19394_), .B(sqrto_27_), .Y(u2__abc_52155_new_n19405_));
OR2X2 OR2X2_4352 ( .A(u2__abc_52155_new_n19408_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19409_));
OR2X2 OR2X2_4353 ( .A(u2__abc_52155_new_n19413_), .B(u2__abc_52155_new_n19404_), .Y(u2__abc_52155_new_n19414_));
OR2X2 OR2X2_4354 ( .A(u2__abc_52155_new_n19406_), .B(sqrto_28_), .Y(u2__abc_52155_new_n19417_));
OR2X2 OR2X2_4355 ( .A(u2__abc_52155_new_n19420_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19421_));
OR2X2 OR2X2_4356 ( .A(u2__abc_52155_new_n19425_), .B(u2__abc_52155_new_n19416_), .Y(u2__abc_52155_new_n19426_));
OR2X2 OR2X2_4357 ( .A(u2__abc_52155_new_n19418_), .B(sqrto_29_), .Y(u2__abc_52155_new_n19429_));
OR2X2 OR2X2_4358 ( .A(u2__abc_52155_new_n19432_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19433_));
OR2X2 OR2X2_4359 ( .A(u2__abc_52155_new_n19437_), .B(u2__abc_52155_new_n19428_), .Y(u2__abc_52155_new_n19438_));
OR2X2 OR2X2_436 ( .A(\a[112] ), .B(\a[105] ), .Y(_abc_73687_new_n1485_));
OR2X2 OR2X2_4360 ( .A(u2__abc_52155_new_n19430_), .B(sqrto_30_), .Y(u2__abc_52155_new_n19441_));
OR2X2 OR2X2_4361 ( .A(u2__abc_52155_new_n19444_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19445_));
OR2X2 OR2X2_4362 ( .A(u2__abc_52155_new_n19449_), .B(u2__abc_52155_new_n19440_), .Y(u2__abc_52155_new_n19450_));
OR2X2 OR2X2_4363 ( .A(u2__abc_52155_new_n19442_), .B(sqrto_31_), .Y(u2__abc_52155_new_n19453_));
OR2X2 OR2X2_4364 ( .A(u2__abc_52155_new_n19456_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19457_));
OR2X2 OR2X2_4365 ( .A(u2__abc_52155_new_n19461_), .B(u2__abc_52155_new_n19452_), .Y(u2__abc_52155_new_n19462_));
OR2X2 OR2X2_4366 ( .A(u2__abc_52155_new_n19454_), .B(sqrto_32_), .Y(u2__abc_52155_new_n19465_));
OR2X2 OR2X2_4367 ( .A(u2__abc_52155_new_n19468_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19469_));
OR2X2 OR2X2_4368 ( .A(u2__abc_52155_new_n19473_), .B(u2__abc_52155_new_n19464_), .Y(u2__abc_52155_new_n19474_));
OR2X2 OR2X2_4369 ( .A(u2__abc_52155_new_n19466_), .B(sqrto_33_), .Y(u2__abc_52155_new_n19477_));
OR2X2 OR2X2_437 ( .A(_abc_73687_new_n1170_), .B(\a[106] ), .Y(_abc_73687_new_n1486_));
OR2X2 OR2X2_4370 ( .A(u2__abc_52155_new_n19480_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19481_));
OR2X2 OR2X2_4371 ( .A(u2__abc_52155_new_n19485_), .B(u2__abc_52155_new_n19476_), .Y(u2__abc_52155_new_n19486_));
OR2X2 OR2X2_4372 ( .A(u2__abc_52155_new_n19478_), .B(sqrto_34_), .Y(u2__abc_52155_new_n19489_));
OR2X2 OR2X2_4373 ( .A(u2__abc_52155_new_n19492_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19493_));
OR2X2 OR2X2_4374 ( .A(u2__abc_52155_new_n19497_), .B(u2__abc_52155_new_n19488_), .Y(u2__abc_52155_new_n19498_));
OR2X2 OR2X2_4375 ( .A(u2__abc_52155_new_n19490_), .B(sqrto_35_), .Y(u2__abc_52155_new_n19501_));
OR2X2 OR2X2_4376 ( .A(u2__abc_52155_new_n19504_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19505_));
OR2X2 OR2X2_4377 ( .A(u2__abc_52155_new_n19509_), .B(u2__abc_52155_new_n19500_), .Y(u2__abc_52155_new_n19510_));
OR2X2 OR2X2_4378 ( .A(u2__abc_52155_new_n19502_), .B(sqrto_36_), .Y(u2__abc_52155_new_n19513_));
OR2X2 OR2X2_4379 ( .A(u2__abc_52155_new_n19516_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19517_));
OR2X2 OR2X2_438 ( .A(\a[112] ), .B(\a[106] ), .Y(_abc_73687_new_n1488_));
OR2X2 OR2X2_4380 ( .A(u2__abc_52155_new_n19521_), .B(u2__abc_52155_new_n19512_), .Y(u2__abc_52155_new_n19522_));
OR2X2 OR2X2_4381 ( .A(u2__abc_52155_new_n19514_), .B(sqrto_37_), .Y(u2__abc_52155_new_n19525_));
OR2X2 OR2X2_4382 ( .A(u2__abc_52155_new_n19528_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19529_));
OR2X2 OR2X2_4383 ( .A(u2__abc_52155_new_n19533_), .B(u2__abc_52155_new_n19524_), .Y(u2__abc_52155_new_n19534_));
OR2X2 OR2X2_4384 ( .A(u2__abc_52155_new_n19526_), .B(sqrto_38_), .Y(u2__abc_52155_new_n19537_));
OR2X2 OR2X2_4385 ( .A(u2__abc_52155_new_n19540_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19541_));
OR2X2 OR2X2_4386 ( .A(u2__abc_52155_new_n19545_), .B(u2__abc_52155_new_n19536_), .Y(u2__abc_52155_new_n19546_));
OR2X2 OR2X2_4387 ( .A(u2__abc_52155_new_n19538_), .B(sqrto_39_), .Y(u2__abc_52155_new_n19549_));
OR2X2 OR2X2_4388 ( .A(u2__abc_52155_new_n19552_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19553_));
OR2X2 OR2X2_4389 ( .A(u2__abc_52155_new_n19557_), .B(u2__abc_52155_new_n19548_), .Y(u2__abc_52155_new_n19558_));
OR2X2 OR2X2_439 ( .A(_abc_73687_new_n1170_), .B(\a[107] ), .Y(_abc_73687_new_n1489_));
OR2X2 OR2X2_4390 ( .A(u2__abc_52155_new_n19550_), .B(sqrto_40_), .Y(u2__abc_52155_new_n19561_));
OR2X2 OR2X2_4391 ( .A(u2__abc_52155_new_n19564_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19565_));
OR2X2 OR2X2_4392 ( .A(u2__abc_52155_new_n19569_), .B(u2__abc_52155_new_n19560_), .Y(u2__abc_52155_new_n19570_));
OR2X2 OR2X2_4393 ( .A(u2__abc_52155_new_n19562_), .B(sqrto_41_), .Y(u2__abc_52155_new_n19573_));
OR2X2 OR2X2_4394 ( .A(u2__abc_52155_new_n19576_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19577_));
OR2X2 OR2X2_4395 ( .A(u2__abc_52155_new_n19581_), .B(u2__abc_52155_new_n19572_), .Y(u2__abc_52155_new_n19582_));
OR2X2 OR2X2_4396 ( .A(u2__abc_52155_new_n19574_), .B(sqrto_42_), .Y(u2__abc_52155_new_n19585_));
OR2X2 OR2X2_4397 ( .A(u2__abc_52155_new_n19588_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19589_));
OR2X2 OR2X2_4398 ( .A(u2__abc_52155_new_n19593_), .B(u2__abc_52155_new_n19584_), .Y(u2__abc_52155_new_n19594_));
OR2X2 OR2X2_4399 ( .A(u2__abc_52155_new_n19586_), .B(sqrto_43_), .Y(u2__abc_52155_new_n19597_));
OR2X2 OR2X2_44 ( .A(_abc_73687_new_n753_), .B(\a[21] ), .Y(_abc_73687_new_n894_));
OR2X2 OR2X2_440 ( .A(\a[112] ), .B(\a[107] ), .Y(_abc_73687_new_n1491_));
OR2X2 OR2X2_4400 ( .A(u2__abc_52155_new_n19600_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19601_));
OR2X2 OR2X2_4401 ( .A(u2__abc_52155_new_n19605_), .B(u2__abc_52155_new_n19596_), .Y(u2__abc_52155_new_n19606_));
OR2X2 OR2X2_4402 ( .A(u2__abc_52155_new_n19598_), .B(sqrto_44_), .Y(u2__abc_52155_new_n19609_));
OR2X2 OR2X2_4403 ( .A(u2__abc_52155_new_n19612_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19613_));
OR2X2 OR2X2_4404 ( .A(u2__abc_52155_new_n19617_), .B(u2__abc_52155_new_n19608_), .Y(u2__abc_52155_new_n19618_));
OR2X2 OR2X2_4405 ( .A(u2__abc_52155_new_n19610_), .B(sqrto_45_), .Y(u2__abc_52155_new_n19621_));
OR2X2 OR2X2_4406 ( .A(u2__abc_52155_new_n19624_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19625_));
OR2X2 OR2X2_4407 ( .A(u2__abc_52155_new_n19629_), .B(u2__abc_52155_new_n19620_), .Y(u2__abc_52155_new_n19630_));
OR2X2 OR2X2_4408 ( .A(u2__abc_52155_new_n19622_), .B(sqrto_46_), .Y(u2__abc_52155_new_n19633_));
OR2X2 OR2X2_4409 ( .A(u2__abc_52155_new_n19636_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19637_));
OR2X2 OR2X2_441 ( .A(_abc_73687_new_n1170_), .B(\a[108] ), .Y(_abc_73687_new_n1492_));
OR2X2 OR2X2_4410 ( .A(u2__abc_52155_new_n19641_), .B(u2__abc_52155_new_n19632_), .Y(u2__abc_52155_new_n19642_));
OR2X2 OR2X2_4411 ( .A(u2__abc_52155_new_n19634_), .B(sqrto_47_), .Y(u2__abc_52155_new_n19645_));
OR2X2 OR2X2_4412 ( .A(u2__abc_52155_new_n19648_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19649_));
OR2X2 OR2X2_4413 ( .A(u2__abc_52155_new_n19653_), .B(u2__abc_52155_new_n19644_), .Y(u2__abc_52155_new_n19654_));
OR2X2 OR2X2_4414 ( .A(u2__abc_52155_new_n19646_), .B(sqrto_48_), .Y(u2__abc_52155_new_n19657_));
OR2X2 OR2X2_4415 ( .A(u2__abc_52155_new_n19660_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19661_));
OR2X2 OR2X2_4416 ( .A(u2__abc_52155_new_n19665_), .B(u2__abc_52155_new_n19656_), .Y(u2__abc_52155_new_n19666_));
OR2X2 OR2X2_4417 ( .A(u2__abc_52155_new_n19658_), .B(sqrto_49_), .Y(u2__abc_52155_new_n19669_));
OR2X2 OR2X2_4418 ( .A(u2__abc_52155_new_n19672_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19673_));
OR2X2 OR2X2_4419 ( .A(u2__abc_52155_new_n19677_), .B(u2__abc_52155_new_n19668_), .Y(u2__abc_52155_new_n19678_));
OR2X2 OR2X2_442 ( .A(\a[112] ), .B(\a[108] ), .Y(_abc_73687_new_n1494_));
OR2X2 OR2X2_4420 ( .A(u2__abc_52155_new_n19670_), .B(sqrto_50_), .Y(u2__abc_52155_new_n19681_));
OR2X2 OR2X2_4421 ( .A(u2__abc_52155_new_n19684_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19685_));
OR2X2 OR2X2_4422 ( .A(u2__abc_52155_new_n19689_), .B(u2__abc_52155_new_n19680_), .Y(u2__abc_52155_new_n19690_));
OR2X2 OR2X2_4423 ( .A(u2__abc_52155_new_n19682_), .B(sqrto_51_), .Y(u2__abc_52155_new_n19693_));
OR2X2 OR2X2_4424 ( .A(u2__abc_52155_new_n19696_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19697_));
OR2X2 OR2X2_4425 ( .A(u2__abc_52155_new_n19701_), .B(u2__abc_52155_new_n19692_), .Y(u2__abc_52155_new_n19702_));
OR2X2 OR2X2_4426 ( .A(u2__abc_52155_new_n19694_), .B(sqrto_52_), .Y(u2__abc_52155_new_n19705_));
OR2X2 OR2X2_4427 ( .A(u2__abc_52155_new_n19708_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19709_));
OR2X2 OR2X2_4428 ( .A(u2__abc_52155_new_n19713_), .B(u2__abc_52155_new_n19704_), .Y(u2__abc_52155_new_n19714_));
OR2X2 OR2X2_4429 ( .A(u2__abc_52155_new_n19706_), .B(sqrto_53_), .Y(u2__abc_52155_new_n19717_));
OR2X2 OR2X2_443 ( .A(_abc_73687_new_n1170_), .B(\a[109] ), .Y(_abc_73687_new_n1495_));
OR2X2 OR2X2_4430 ( .A(u2__abc_52155_new_n19720_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19721_));
OR2X2 OR2X2_4431 ( .A(u2__abc_52155_new_n19725_), .B(u2__abc_52155_new_n19716_), .Y(u2__abc_52155_new_n19726_));
OR2X2 OR2X2_4432 ( .A(u2__abc_52155_new_n19718_), .B(sqrto_54_), .Y(u2__abc_52155_new_n19729_));
OR2X2 OR2X2_4433 ( .A(u2__abc_52155_new_n19732_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19733_));
OR2X2 OR2X2_4434 ( .A(u2__abc_52155_new_n19737_), .B(u2__abc_52155_new_n19728_), .Y(u2__abc_52155_new_n19738_));
OR2X2 OR2X2_4435 ( .A(u2__abc_52155_new_n19730_), .B(sqrto_55_), .Y(u2__abc_52155_new_n19741_));
OR2X2 OR2X2_4436 ( .A(u2__abc_52155_new_n19744_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19745_));
OR2X2 OR2X2_4437 ( .A(u2__abc_52155_new_n19749_), .B(u2__abc_52155_new_n19740_), .Y(u2__abc_52155_new_n19750_));
OR2X2 OR2X2_4438 ( .A(u2__abc_52155_new_n19742_), .B(sqrto_56_), .Y(u2__abc_52155_new_n19753_));
OR2X2 OR2X2_4439 ( .A(u2__abc_52155_new_n19756_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19757_));
OR2X2 OR2X2_444 ( .A(\a[112] ), .B(\a[109] ), .Y(_abc_73687_new_n1497_));
OR2X2 OR2X2_4440 ( .A(u2__abc_52155_new_n19761_), .B(u2__abc_52155_new_n19752_), .Y(u2__abc_52155_new_n19762_));
OR2X2 OR2X2_4441 ( .A(u2__abc_52155_new_n19754_), .B(sqrto_57_), .Y(u2__abc_52155_new_n19765_));
OR2X2 OR2X2_4442 ( .A(u2__abc_52155_new_n19768_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19769_));
OR2X2 OR2X2_4443 ( .A(u2__abc_52155_new_n19773_), .B(u2__abc_52155_new_n19764_), .Y(u2__abc_52155_new_n19774_));
OR2X2 OR2X2_4444 ( .A(u2__abc_52155_new_n19766_), .B(sqrto_58_), .Y(u2__abc_52155_new_n19777_));
OR2X2 OR2X2_4445 ( .A(u2__abc_52155_new_n19780_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19781_));
OR2X2 OR2X2_4446 ( .A(u2__abc_52155_new_n19785_), .B(u2__abc_52155_new_n19776_), .Y(u2__abc_52155_new_n19786_));
OR2X2 OR2X2_4447 ( .A(u2__abc_52155_new_n19778_), .B(sqrto_59_), .Y(u2__abc_52155_new_n19789_));
OR2X2 OR2X2_4448 ( .A(u2__abc_52155_new_n19792_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19793_));
OR2X2 OR2X2_4449 ( .A(u2__abc_52155_new_n19797_), .B(u2__abc_52155_new_n19788_), .Y(u2__abc_52155_new_n19798_));
OR2X2 OR2X2_445 ( .A(_abc_73687_new_n1170_), .B(\a[110] ), .Y(_abc_73687_new_n1498_));
OR2X2 OR2X2_4450 ( .A(u2__abc_52155_new_n19790_), .B(sqrto_60_), .Y(u2__abc_52155_new_n19801_));
OR2X2 OR2X2_4451 ( .A(u2__abc_52155_new_n19804_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19805_));
OR2X2 OR2X2_4452 ( .A(u2__abc_52155_new_n19809_), .B(u2__abc_52155_new_n19800_), .Y(u2__abc_52155_new_n19810_));
OR2X2 OR2X2_4453 ( .A(u2__abc_52155_new_n19802_), .B(sqrto_61_), .Y(u2__abc_52155_new_n19813_));
OR2X2 OR2X2_4454 ( .A(u2__abc_52155_new_n19816_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19817_));
OR2X2 OR2X2_4455 ( .A(u2__abc_52155_new_n19821_), .B(u2__abc_52155_new_n19812_), .Y(u2__abc_52155_new_n19822_));
OR2X2 OR2X2_4456 ( .A(u2__abc_52155_new_n19814_), .B(sqrto_62_), .Y(u2__abc_52155_new_n19825_));
OR2X2 OR2X2_4457 ( .A(u2__abc_52155_new_n19828_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19829_));
OR2X2 OR2X2_4458 ( .A(u2__abc_52155_new_n19833_), .B(u2__abc_52155_new_n19824_), .Y(u2__abc_52155_new_n19834_));
OR2X2 OR2X2_4459 ( .A(u2__abc_52155_new_n19826_), .B(sqrto_63_), .Y(u2__abc_52155_new_n19837_));
OR2X2 OR2X2_446 ( .A(\a[112] ), .B(\a[110] ), .Y(_abc_73687_new_n1500_));
OR2X2 OR2X2_4460 ( .A(u2__abc_52155_new_n19840_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19841_));
OR2X2 OR2X2_4461 ( .A(u2__abc_52155_new_n19845_), .B(u2__abc_52155_new_n19836_), .Y(u2__abc_52155_new_n19846_));
OR2X2 OR2X2_4462 ( .A(u2__abc_52155_new_n19838_), .B(sqrto_64_), .Y(u2__abc_52155_new_n19849_));
OR2X2 OR2X2_4463 ( .A(u2__abc_52155_new_n19852_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19853_));
OR2X2 OR2X2_4464 ( .A(u2__abc_52155_new_n19857_), .B(u2__abc_52155_new_n19848_), .Y(u2__abc_52155_new_n19858_));
OR2X2 OR2X2_4465 ( .A(u2__abc_52155_new_n19850_), .B(sqrto_65_), .Y(u2__abc_52155_new_n19861_));
OR2X2 OR2X2_4466 ( .A(u2__abc_52155_new_n19864_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19865_));
OR2X2 OR2X2_4467 ( .A(u2__abc_52155_new_n19869_), .B(u2__abc_52155_new_n19860_), .Y(u2__abc_52155_new_n19870_));
OR2X2 OR2X2_4468 ( .A(u2__abc_52155_new_n19862_), .B(sqrto_66_), .Y(u2__abc_52155_new_n19873_));
OR2X2 OR2X2_4469 ( .A(u2__abc_52155_new_n19876_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19877_));
OR2X2 OR2X2_447 ( .A(_abc_73687_new_n1170_), .B(\a[111] ), .Y(_abc_73687_new_n1501_));
OR2X2 OR2X2_4470 ( .A(u2__abc_52155_new_n19881_), .B(u2__abc_52155_new_n19872_), .Y(u2__abc_52155_new_n19882_));
OR2X2 OR2X2_4471 ( .A(u2__abc_52155_new_n19874_), .B(sqrto_67_), .Y(u2__abc_52155_new_n19885_));
OR2X2 OR2X2_4472 ( .A(u2__abc_52155_new_n19888_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19889_));
OR2X2 OR2X2_4473 ( .A(u2__abc_52155_new_n19893_), .B(u2__abc_52155_new_n19884_), .Y(u2__abc_52155_new_n19894_));
OR2X2 OR2X2_4474 ( .A(u2__abc_52155_new_n19886_), .B(sqrto_68_), .Y(u2__abc_52155_new_n19897_));
OR2X2 OR2X2_4475 ( .A(u2__abc_52155_new_n19900_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19901_));
OR2X2 OR2X2_4476 ( .A(u2__abc_52155_new_n19905_), .B(u2__abc_52155_new_n19896_), .Y(u2__abc_52155_new_n19906_));
OR2X2 OR2X2_4477 ( .A(u2__abc_52155_new_n19898_), .B(sqrto_69_), .Y(u2__abc_52155_new_n19909_));
OR2X2 OR2X2_4478 ( .A(u2__abc_52155_new_n19912_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19913_));
OR2X2 OR2X2_4479 ( .A(u2__abc_52155_new_n19917_), .B(u2__abc_52155_new_n19908_), .Y(u2__abc_52155_new_n19918_));
OR2X2 OR2X2_448 ( .A(\a[112] ), .B(\a[111] ), .Y(_abc_73687_new_n1503_));
OR2X2 OR2X2_4480 ( .A(u2__abc_52155_new_n19910_), .B(sqrto_70_), .Y(u2__abc_52155_new_n19921_));
OR2X2 OR2X2_4481 ( .A(u2__abc_52155_new_n19924_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19925_));
OR2X2 OR2X2_4482 ( .A(u2__abc_52155_new_n19929_), .B(u2__abc_52155_new_n19920_), .Y(u2__abc_52155_new_n19930_));
OR2X2 OR2X2_4483 ( .A(u2__abc_52155_new_n19922_), .B(sqrto_71_), .Y(u2__abc_52155_new_n19933_));
OR2X2 OR2X2_4484 ( .A(u2__abc_52155_new_n19936_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19937_));
OR2X2 OR2X2_4485 ( .A(u2__abc_52155_new_n19941_), .B(u2__abc_52155_new_n19932_), .Y(u2__abc_52155_new_n19942_));
OR2X2 OR2X2_4486 ( .A(u2__abc_52155_new_n19934_), .B(sqrto_72_), .Y(u2__abc_52155_new_n19945_));
OR2X2 OR2X2_4487 ( .A(u2__abc_52155_new_n19948_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19949_));
OR2X2 OR2X2_4488 ( .A(u2__abc_52155_new_n19953_), .B(u2__abc_52155_new_n19944_), .Y(u2__abc_52155_new_n19954_));
OR2X2 OR2X2_4489 ( .A(u2__abc_52155_new_n19946_), .B(sqrto_73_), .Y(u2__abc_52155_new_n19957_));
OR2X2 OR2X2_449 ( .A(_abc_73687_new_n1170_), .B(fracta_112_), .Y(_abc_73687_new_n1504_));
OR2X2 OR2X2_4490 ( .A(u2__abc_52155_new_n19960_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19961_));
OR2X2 OR2X2_4491 ( .A(u2__abc_52155_new_n19965_), .B(u2__abc_52155_new_n19956_), .Y(u2__abc_52155_new_n19966_));
OR2X2 OR2X2_4492 ( .A(u2__abc_52155_new_n19958_), .B(sqrto_74_), .Y(u2__abc_52155_new_n19969_));
OR2X2 OR2X2_4493 ( .A(u2__abc_52155_new_n19972_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19973_));
OR2X2 OR2X2_4494 ( .A(u2__abc_52155_new_n19977_), .B(u2__abc_52155_new_n19968_), .Y(u2__abc_52155_new_n19978_));
OR2X2 OR2X2_4495 ( .A(u2__abc_52155_new_n19970_), .B(sqrto_75_), .Y(u2__abc_52155_new_n19981_));
OR2X2 OR2X2_4496 ( .A(u2__abc_52155_new_n19984_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19985_));
OR2X2 OR2X2_4497 ( .A(u2__abc_52155_new_n19989_), .B(u2__abc_52155_new_n19980_), .Y(u2__abc_52155_new_n19990_));
OR2X2 OR2X2_4498 ( .A(u2__abc_52155_new_n19982_), .B(sqrto_76_), .Y(u2__abc_52155_new_n19993_));
OR2X2 OR2X2_4499 ( .A(u2__abc_52155_new_n19996_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n19997_));
OR2X2 OR2X2_45 ( .A(aNan), .B(sqrto_98_), .Y(_abc_73687_new_n896_));
OR2X2 OR2X2_450 ( .A(_abc_73687_new_n1509_), .B(_abc_73687_new_n1507_), .Y(_abc_73687_new_n1510_));
OR2X2 OR2X2_4500 ( .A(u2__abc_52155_new_n20001_), .B(u2__abc_52155_new_n19992_), .Y(u2__abc_52155_new_n20002_));
OR2X2 OR2X2_4501 ( .A(u2__abc_52155_new_n19994_), .B(sqrto_77_), .Y(u2__abc_52155_new_n20005_));
OR2X2 OR2X2_4502 ( .A(u2__abc_52155_new_n20008_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20009_));
OR2X2 OR2X2_4503 ( .A(u2__abc_52155_new_n20013_), .B(u2__abc_52155_new_n20004_), .Y(u2__abc_52155_new_n20014_));
OR2X2 OR2X2_4504 ( .A(u2__abc_52155_new_n20006_), .B(sqrto_78_), .Y(u2__abc_52155_new_n20017_));
OR2X2 OR2X2_4505 ( .A(u2__abc_52155_new_n20020_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20021_));
OR2X2 OR2X2_4506 ( .A(u2__abc_52155_new_n20025_), .B(u2__abc_52155_new_n20016_), .Y(u2__abc_52155_new_n20026_));
OR2X2 OR2X2_4507 ( .A(u2__abc_52155_new_n20018_), .B(sqrto_79_), .Y(u2__abc_52155_new_n20031_));
OR2X2 OR2X2_4508 ( .A(u2__abc_52155_new_n20032_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20033_));
OR2X2 OR2X2_4509 ( .A(u2__abc_52155_new_n20037_), .B(u2__abc_52155_new_n20028_), .Y(u2__abc_52155_new_n20038_));
OR2X2 OR2X2_451 ( .A(_abc_73687_new_n1511_), .B(_abc_73687_new_n1512_), .Y(\o[226] ));
OR2X2 OR2X2_4510 ( .A(u2__abc_52155_new_n20029_), .B(sqrto_80_), .Y(u2__abc_52155_new_n20041_));
OR2X2 OR2X2_4511 ( .A(u2__abc_52155_new_n20044_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20045_));
OR2X2 OR2X2_4512 ( .A(u2__abc_52155_new_n20049_), .B(u2__abc_52155_new_n20040_), .Y(u2__abc_52155_new_n20050_));
OR2X2 OR2X2_4513 ( .A(u2__abc_52155_new_n20042_), .B(sqrto_81_), .Y(u2__abc_52155_new_n20053_));
OR2X2 OR2X2_4514 ( .A(u2__abc_52155_new_n20056_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20057_));
OR2X2 OR2X2_4515 ( .A(u2__abc_52155_new_n20061_), .B(u2__abc_52155_new_n20052_), .Y(u2__abc_52155_new_n20062_));
OR2X2 OR2X2_4516 ( .A(u2__abc_52155_new_n20054_), .B(sqrto_82_), .Y(u2__abc_52155_new_n20065_));
OR2X2 OR2X2_4517 ( .A(u2__abc_52155_new_n20068_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20069_));
OR2X2 OR2X2_4518 ( .A(u2__abc_52155_new_n20073_), .B(u2__abc_52155_new_n20064_), .Y(u2__abc_52155_new_n20074_));
OR2X2 OR2X2_4519 ( .A(u2__abc_52155_new_n20066_), .B(sqrto_83_), .Y(u2__abc_52155_new_n20077_));
OR2X2 OR2X2_452 ( .A(aNan), .B(\a[114] ), .Y(_abc_73687_new_n1514_));
OR2X2 OR2X2_4520 ( .A(u2__abc_52155_new_n20080_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20081_));
OR2X2 OR2X2_4521 ( .A(u2__abc_52155_new_n20085_), .B(u2__abc_52155_new_n20076_), .Y(u2__abc_52155_new_n20086_));
OR2X2 OR2X2_4522 ( .A(u2__abc_52155_new_n20078_), .B(sqrto_84_), .Y(u2__abc_52155_new_n20089_));
OR2X2 OR2X2_4523 ( .A(u2__abc_52155_new_n20092_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20093_));
OR2X2 OR2X2_4524 ( .A(u2__abc_52155_new_n20097_), .B(u2__abc_52155_new_n20088_), .Y(u2__abc_52155_new_n20098_));
OR2X2 OR2X2_4525 ( .A(u2__abc_52155_new_n20090_), .B(sqrto_85_), .Y(u2__abc_52155_new_n20101_));
OR2X2 OR2X2_4526 ( .A(u2__abc_52155_new_n20104_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20105_));
OR2X2 OR2X2_4527 ( .A(u2__abc_52155_new_n20109_), .B(u2__abc_52155_new_n20100_), .Y(u2__abc_52155_new_n20110_));
OR2X2 OR2X2_4528 ( .A(u2__abc_52155_new_n20102_), .B(sqrto_86_), .Y(u2__abc_52155_new_n20113_));
OR2X2 OR2X2_4529 ( .A(u2__abc_52155_new_n20116_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20117_));
OR2X2 OR2X2_453 ( .A(_abc_73687_new_n1509_), .B(_abc_73687_new_n1514_), .Y(_abc_73687_new_n1515_));
OR2X2 OR2X2_4530 ( .A(u2__abc_52155_new_n20121_), .B(u2__abc_52155_new_n20112_), .Y(u2__abc_52155_new_n20122_));
OR2X2 OR2X2_4531 ( .A(u2__abc_52155_new_n20114_), .B(sqrto_87_), .Y(u2__abc_52155_new_n20127_));
OR2X2 OR2X2_4532 ( .A(u2__abc_52155_new_n20128_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20129_));
OR2X2 OR2X2_4533 ( .A(u2__abc_52155_new_n20133_), .B(u2__abc_52155_new_n20124_), .Y(u2__abc_52155_new_n20134_));
OR2X2 OR2X2_4534 ( .A(u2__abc_52155_new_n20125_), .B(sqrto_88_), .Y(u2__abc_52155_new_n20137_));
OR2X2 OR2X2_4535 ( .A(u2__abc_52155_new_n20140_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20141_));
OR2X2 OR2X2_4536 ( .A(u2__abc_52155_new_n20145_), .B(u2__abc_52155_new_n20136_), .Y(u2__abc_52155_new_n20146_));
OR2X2 OR2X2_4537 ( .A(u2__abc_52155_new_n20138_), .B(sqrto_89_), .Y(u2__abc_52155_new_n20149_));
OR2X2 OR2X2_4538 ( .A(u2__abc_52155_new_n20152_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20153_));
OR2X2 OR2X2_4539 ( .A(u2__abc_52155_new_n20157_), .B(u2__abc_52155_new_n20148_), .Y(u2__abc_52155_new_n20158_));
OR2X2 OR2X2_454 ( .A(_abc_73687_new_n1516_), .B(\a[112] ), .Y(_abc_73687_new_n1517_));
OR2X2 OR2X2_4540 ( .A(u2__abc_52155_new_n20150_), .B(sqrto_90_), .Y(u2__abc_52155_new_n20161_));
OR2X2 OR2X2_4541 ( .A(u2__abc_52155_new_n20164_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20165_));
OR2X2 OR2X2_4542 ( .A(u2__abc_52155_new_n20169_), .B(u2__abc_52155_new_n20160_), .Y(u2__abc_52155_new_n20170_));
OR2X2 OR2X2_4543 ( .A(u2__abc_52155_new_n20162_), .B(sqrto_91_), .Y(u2__abc_52155_new_n20175_));
OR2X2 OR2X2_4544 ( .A(u2__abc_52155_new_n20176_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20177_));
OR2X2 OR2X2_4545 ( .A(u2__abc_52155_new_n20181_), .B(u2__abc_52155_new_n20172_), .Y(u2__abc_52155_new_n20182_));
OR2X2 OR2X2_4546 ( .A(u2__abc_52155_new_n20173_), .B(sqrto_92_), .Y(u2__abc_52155_new_n20185_));
OR2X2 OR2X2_4547 ( .A(u2__abc_52155_new_n20188_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20189_));
OR2X2 OR2X2_4548 ( .A(u2__abc_52155_new_n20193_), .B(u2__abc_52155_new_n20184_), .Y(u2__abc_52155_new_n20194_));
OR2X2 OR2X2_4549 ( .A(u2__abc_52155_new_n20186_), .B(sqrto_93_), .Y(u2__abc_52155_new_n20199_));
OR2X2 OR2X2_455 ( .A(_abc_73687_new_n1518_), .B(\a[113] ), .Y(_abc_73687_new_n1519_));
OR2X2 OR2X2_4550 ( .A(u2__abc_52155_new_n20200_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20201_));
OR2X2 OR2X2_4551 ( .A(u2__abc_52155_new_n20205_), .B(u2__abc_52155_new_n20196_), .Y(u2__abc_52155_new_n20206_));
OR2X2 OR2X2_4552 ( .A(u2__abc_52155_new_n20197_), .B(sqrto_94_), .Y(u2__abc_52155_new_n20209_));
OR2X2 OR2X2_4553 ( .A(u2__abc_52155_new_n20212_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20213_));
OR2X2 OR2X2_4554 ( .A(u2__abc_52155_new_n20217_), .B(u2__abc_52155_new_n20208_), .Y(u2__abc_52155_new_n20218_));
OR2X2 OR2X2_4555 ( .A(u2__abc_52155_new_n20210_), .B(sqrto_95_), .Y(u2__abc_52155_new_n20221_));
OR2X2 OR2X2_4556 ( .A(u2__abc_52155_new_n20224_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20225_));
OR2X2 OR2X2_4557 ( .A(u2__abc_52155_new_n20229_), .B(u2__abc_52155_new_n20220_), .Y(u2__abc_52155_new_n20230_));
OR2X2 OR2X2_4558 ( .A(u2__abc_52155_new_n20222_), .B(sqrto_96_), .Y(u2__abc_52155_new_n20233_));
OR2X2 OR2X2_4559 ( .A(u2__abc_52155_new_n20236_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20237_));
OR2X2 OR2X2_456 ( .A(_abc_73687_new_n1525_), .B(\a[114] ), .Y(_abc_73687_new_n1526_));
OR2X2 OR2X2_4560 ( .A(u2__abc_52155_new_n20241_), .B(u2__abc_52155_new_n20232_), .Y(u2__abc_52155_new_n20242_));
OR2X2 OR2X2_4561 ( .A(u2__abc_52155_new_n20234_), .B(sqrto_97_), .Y(u2__abc_52155_new_n20245_));
OR2X2 OR2X2_4562 ( .A(u2__abc_52155_new_n20248_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20249_));
OR2X2 OR2X2_4563 ( .A(u2__abc_52155_new_n20253_), .B(u2__abc_52155_new_n20244_), .Y(u2__abc_52155_new_n20254_));
OR2X2 OR2X2_4564 ( .A(u2__abc_52155_new_n20246_), .B(sqrto_98_), .Y(u2__abc_52155_new_n20257_));
OR2X2 OR2X2_4565 ( .A(u2__abc_52155_new_n20260_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20261_));
OR2X2 OR2X2_4566 ( .A(u2__abc_52155_new_n20265_), .B(u2__abc_52155_new_n20256_), .Y(u2__abc_52155_new_n20266_));
OR2X2 OR2X2_4567 ( .A(u2__abc_52155_new_n20258_), .B(sqrto_99_), .Y(u2__abc_52155_new_n20269_));
OR2X2 OR2X2_4568 ( .A(u2__abc_52155_new_n20272_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20273_));
OR2X2 OR2X2_4569 ( .A(u2__abc_52155_new_n20277_), .B(u2__abc_52155_new_n20268_), .Y(u2__abc_52155_new_n20278_));
OR2X2 OR2X2_457 ( .A(_abc_73687_new_n1527_), .B(_abc_73687_new_n1523_), .Y(_abc_73687_new_n1528_));
OR2X2 OR2X2_4570 ( .A(u2__abc_52155_new_n20270_), .B(sqrto_100_), .Y(u2__abc_52155_new_n20281_));
OR2X2 OR2X2_4571 ( .A(u2__abc_52155_new_n20284_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20285_));
OR2X2 OR2X2_4572 ( .A(u2__abc_52155_new_n20289_), .B(u2__abc_52155_new_n20280_), .Y(u2__abc_52155_new_n20290_));
OR2X2 OR2X2_4573 ( .A(u2__abc_52155_new_n20282_), .B(sqrto_101_), .Y(u2__abc_52155_new_n20293_));
OR2X2 OR2X2_4574 ( .A(u2__abc_52155_new_n20296_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20297_));
OR2X2 OR2X2_4575 ( .A(u2__abc_52155_new_n20301_), .B(u2__abc_52155_new_n20292_), .Y(u2__abc_52155_new_n20302_));
OR2X2 OR2X2_4576 ( .A(u2__abc_52155_new_n20294_), .B(sqrto_102_), .Y(u2__abc_52155_new_n20305_));
OR2X2 OR2X2_4577 ( .A(u2__abc_52155_new_n20308_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20309_));
OR2X2 OR2X2_4578 ( .A(u2__abc_52155_new_n20313_), .B(u2__abc_52155_new_n20304_), .Y(u2__abc_52155_new_n20314_));
OR2X2 OR2X2_4579 ( .A(u2__abc_52155_new_n20306_), .B(sqrto_103_), .Y(u2__abc_52155_new_n20319_));
OR2X2 OR2X2_458 ( .A(_abc_73687_new_n1526_), .B(_abc_73687_new_n1522_), .Y(_abc_73687_new_n1529_));
OR2X2 OR2X2_4580 ( .A(u2__abc_52155_new_n20320_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20321_));
OR2X2 OR2X2_4581 ( .A(u2__abc_52155_new_n20325_), .B(u2__abc_52155_new_n20316_), .Y(u2__abc_52155_new_n20326_));
OR2X2 OR2X2_4582 ( .A(u2__abc_52155_new_n20317_), .B(sqrto_104_), .Y(u2__abc_52155_new_n20329_));
OR2X2 OR2X2_4583 ( .A(u2__abc_52155_new_n20332_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20333_));
OR2X2 OR2X2_4584 ( .A(u2__abc_52155_new_n20337_), .B(u2__abc_52155_new_n20328_), .Y(u2__abc_52155_new_n20338_));
OR2X2 OR2X2_4585 ( .A(u2__abc_52155_new_n20330_), .B(sqrto_105_), .Y(u2__abc_52155_new_n20341_));
OR2X2 OR2X2_4586 ( .A(u2__abc_52155_new_n20344_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20345_));
OR2X2 OR2X2_4587 ( .A(u2__abc_52155_new_n20349_), .B(u2__abc_52155_new_n20340_), .Y(u2__abc_52155_new_n20350_));
OR2X2 OR2X2_4588 ( .A(u2__abc_52155_new_n20342_), .B(sqrto_106_), .Y(u2__abc_52155_new_n20353_));
OR2X2 OR2X2_4589 ( .A(u2__abc_52155_new_n20356_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20357_));
OR2X2 OR2X2_459 ( .A(_abc_73687_new_n1534_), .B(_abc_73687_new_n1532_), .Y(_abc_73687_new_n1535_));
OR2X2 OR2X2_4590 ( .A(u2__abc_52155_new_n20361_), .B(u2__abc_52155_new_n20352_), .Y(u2__abc_52155_new_n20362_));
OR2X2 OR2X2_4591 ( .A(u2__abc_52155_new_n20354_), .B(sqrto_107_), .Y(u2__abc_52155_new_n20367_));
OR2X2 OR2X2_4592 ( .A(u2__abc_52155_new_n20368_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20369_));
OR2X2 OR2X2_4593 ( .A(u2__abc_52155_new_n20373_), .B(u2__abc_52155_new_n20364_), .Y(u2__abc_52155_new_n20374_));
OR2X2 OR2X2_4594 ( .A(u2__abc_52155_new_n20365_), .B(sqrto_108_), .Y(u2__abc_52155_new_n20377_));
OR2X2 OR2X2_4595 ( .A(u2__abc_52155_new_n20380_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20381_));
OR2X2 OR2X2_4596 ( .A(u2__abc_52155_new_n20385_), .B(u2__abc_52155_new_n20376_), .Y(u2__abc_52155_new_n20386_));
OR2X2 OR2X2_4597 ( .A(u2__abc_52155_new_n20378_), .B(sqrto_109_), .Y(u2__abc_52155_new_n20391_));
OR2X2 OR2X2_4598 ( .A(u2__abc_52155_new_n20392_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20393_));
OR2X2 OR2X2_4599 ( .A(u2__abc_52155_new_n20397_), .B(u2__abc_52155_new_n20388_), .Y(u2__abc_52155_new_n20398_));
OR2X2 OR2X2_46 ( .A(_abc_73687_new_n753_), .B(\a[22] ), .Y(_abc_73687_new_n897_));
OR2X2 OR2X2_460 ( .A(_abc_73687_new_n1539_), .B(_abc_73687_new_n1536_), .Y(_abc_73687_new_n1540_));
OR2X2 OR2X2_4600 ( .A(u2__abc_52155_new_n20389_), .B(sqrto_110_), .Y(u2__abc_52155_new_n20401_));
OR2X2 OR2X2_4601 ( .A(u2__abc_52155_new_n20404_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20405_));
OR2X2 OR2X2_4602 ( .A(u2__abc_52155_new_n20409_), .B(u2__abc_52155_new_n20400_), .Y(u2__abc_52155_new_n20410_));
OR2X2 OR2X2_4603 ( .A(u2__abc_52155_new_n20402_), .B(sqrto_111_), .Y(u2__abc_52155_new_n20413_));
OR2X2 OR2X2_4604 ( .A(u2__abc_52155_new_n20416_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20417_));
OR2X2 OR2X2_4605 ( .A(u2__abc_52155_new_n20421_), .B(u2__abc_52155_new_n20412_), .Y(u2__abc_52155_new_n20422_));
OR2X2 OR2X2_4606 ( .A(u2__abc_52155_new_n20414_), .B(sqrto_112_), .Y(u2__abc_52155_new_n20425_));
OR2X2 OR2X2_4607 ( .A(u2__abc_52155_new_n20428_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20429_));
OR2X2 OR2X2_4608 ( .A(u2__abc_52155_new_n20433_), .B(u2__abc_52155_new_n20424_), .Y(u2__abc_52155_new_n20434_));
OR2X2 OR2X2_4609 ( .A(u2__abc_52155_new_n20426_), .B(sqrto_113_), .Y(u2__abc_52155_new_n20437_));
OR2X2 OR2X2_461 ( .A(_abc_73687_new_n1541_), .B(_abc_73687_new_n1543_), .Y(_abc_73687_new_n1544_));
OR2X2 OR2X2_4610 ( .A(u2__abc_52155_new_n20440_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20441_));
OR2X2 OR2X2_4611 ( .A(u2__abc_52155_new_n20445_), .B(u2__abc_52155_new_n20436_), .Y(u2__abc_52155_new_n20446_));
OR2X2 OR2X2_4612 ( .A(u2__abc_52155_new_n20438_), .B(sqrto_114_), .Y(u2__abc_52155_new_n20449_));
OR2X2 OR2X2_4613 ( .A(u2__abc_52155_new_n20452_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20453_));
OR2X2 OR2X2_4614 ( .A(u2__abc_52155_new_n20457_), .B(u2__abc_52155_new_n20448_), .Y(u2__abc_52155_new_n20458_));
OR2X2 OR2X2_4615 ( .A(u2__abc_52155_new_n20450_), .B(sqrto_115_), .Y(u2__abc_52155_new_n20463_));
OR2X2 OR2X2_4616 ( .A(u2__abc_52155_new_n20464_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20465_));
OR2X2 OR2X2_4617 ( .A(u2__abc_52155_new_n20469_), .B(u2__abc_52155_new_n20460_), .Y(u2__abc_52155_new_n20470_));
OR2X2 OR2X2_4618 ( .A(u2__abc_52155_new_n20461_), .B(sqrto_116_), .Y(u2__abc_52155_new_n20473_));
OR2X2 OR2X2_4619 ( .A(u2__abc_52155_new_n20476_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20477_));
OR2X2 OR2X2_462 ( .A(_abc_73687_new_n1545_), .B(_abc_73687_new_n1546_), .Y(\o[229] ));
OR2X2 OR2X2_4620 ( .A(u2__abc_52155_new_n20481_), .B(u2__abc_52155_new_n20472_), .Y(u2__abc_52155_new_n20482_));
OR2X2 OR2X2_4621 ( .A(u2__abc_52155_new_n20474_), .B(sqrto_117_), .Y(u2__abc_52155_new_n20487_));
OR2X2 OR2X2_4622 ( .A(u2__abc_52155_new_n20488_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20489_));
OR2X2 OR2X2_4623 ( .A(u2__abc_52155_new_n20493_), .B(u2__abc_52155_new_n20484_), .Y(u2__abc_52155_new_n20494_));
OR2X2 OR2X2_4624 ( .A(u2__abc_52155_new_n20485_), .B(sqrto_118_), .Y(u2__abc_52155_new_n20497_));
OR2X2 OR2X2_4625 ( .A(u2__abc_52155_new_n20500_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20501_));
OR2X2 OR2X2_4626 ( .A(u2__abc_52155_new_n20505_), .B(u2__abc_52155_new_n20496_), .Y(u2__abc_52155_new_n20506_));
OR2X2 OR2X2_4627 ( .A(u2__abc_52155_new_n20498_), .B(sqrto_119_), .Y(u2__abc_52155_new_n20509_));
OR2X2 OR2X2_4628 ( .A(u2__abc_52155_new_n20512_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20513_));
OR2X2 OR2X2_4629 ( .A(u2__abc_52155_new_n20517_), .B(u2__abc_52155_new_n20508_), .Y(u2__abc_52155_new_n20518_));
OR2X2 OR2X2_463 ( .A(_abc_73687_new_n1550_), .B(_abc_73687_new_n1551_), .Y(_abc_73687_new_n1552_));
OR2X2 OR2X2_4630 ( .A(u2__abc_52155_new_n20510_), .B(sqrto_120_), .Y(u2__abc_52155_new_n20521_));
OR2X2 OR2X2_4631 ( .A(u2__abc_52155_new_n20524_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20525_));
OR2X2 OR2X2_4632 ( .A(u2__abc_52155_new_n20529_), .B(u2__abc_52155_new_n20520_), .Y(u2__abc_52155_new_n20530_));
OR2X2 OR2X2_4633 ( .A(u2__abc_52155_new_n20522_), .B(sqrto_121_), .Y(u2__abc_52155_new_n20535_));
OR2X2 OR2X2_4634 ( .A(u2__abc_52155_new_n20536_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20537_));
OR2X2 OR2X2_4635 ( .A(u2__abc_52155_new_n20541_), .B(u2__abc_52155_new_n20532_), .Y(u2__abc_52155_new_n20542_));
OR2X2 OR2X2_4636 ( .A(u2__abc_52155_new_n20533_), .B(sqrto_122_), .Y(u2__abc_52155_new_n20545_));
OR2X2 OR2X2_4637 ( .A(u2__abc_52155_new_n20548_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20549_));
OR2X2 OR2X2_4638 ( .A(u2__abc_52155_new_n20553_), .B(u2__abc_52155_new_n20544_), .Y(u2__abc_52155_new_n20554_));
OR2X2 OR2X2_4639 ( .A(u2__abc_52155_new_n20546_), .B(sqrto_123_), .Y(u2__abc_52155_new_n20557_));
OR2X2 OR2X2_464 ( .A(_abc_73687_new_n1556_), .B(_abc_73687_new_n1553_), .Y(_abc_73687_new_n1557_));
OR2X2 OR2X2_4640 ( .A(u2__abc_52155_new_n20560_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20561_));
OR2X2 OR2X2_4641 ( .A(u2__abc_52155_new_n20565_), .B(u2__abc_52155_new_n20556_), .Y(u2__abc_52155_new_n20566_));
OR2X2 OR2X2_4642 ( .A(u2__abc_52155_new_n20558_), .B(sqrto_124_), .Y(u2__abc_52155_new_n20569_));
OR2X2 OR2X2_4643 ( .A(u2__abc_52155_new_n20572_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20573_));
OR2X2 OR2X2_4644 ( .A(u2__abc_52155_new_n20577_), .B(u2__abc_52155_new_n20568_), .Y(u2__abc_52155_new_n20578_));
OR2X2 OR2X2_4645 ( .A(u2__abc_52155_new_n20570_), .B(sqrto_125_), .Y(u2__abc_52155_new_n20583_));
OR2X2 OR2X2_4646 ( .A(u2__abc_52155_new_n20584_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20585_));
OR2X2 OR2X2_4647 ( .A(u2__abc_52155_new_n20589_), .B(u2__abc_52155_new_n20580_), .Y(u2__abc_52155_new_n20590_));
OR2X2 OR2X2_4648 ( .A(u2__abc_52155_new_n20581_), .B(sqrto_126_), .Y(u2__abc_52155_new_n20593_));
OR2X2 OR2X2_4649 ( .A(u2__abc_52155_new_n20596_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20597_));
OR2X2 OR2X2_465 ( .A(_abc_73687_new_n1557_), .B(aNan), .Y(_abc_73687_new_n1558_));
OR2X2 OR2X2_4650 ( .A(u2__abc_52155_new_n20601_), .B(u2__abc_52155_new_n20592_), .Y(u2__abc_52155_new_n20602_));
OR2X2 OR2X2_4651 ( .A(u2__abc_52155_new_n20594_), .B(sqrto_127_), .Y(u2__abc_52155_new_n20605_));
OR2X2 OR2X2_4652 ( .A(u2__abc_52155_new_n20608_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20609_));
OR2X2 OR2X2_4653 ( .A(u2__abc_52155_new_n20613_), .B(u2__abc_52155_new_n20604_), .Y(u2__abc_52155_new_n20614_));
OR2X2 OR2X2_4654 ( .A(u2__abc_52155_new_n20606_), .B(sqrto_128_), .Y(u2__abc_52155_new_n20617_));
OR2X2 OR2X2_4655 ( .A(u2__abc_52155_new_n20620_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20621_));
OR2X2 OR2X2_4656 ( .A(u2__abc_52155_new_n20625_), .B(u2__abc_52155_new_n20616_), .Y(u2__abc_52155_new_n20626_));
OR2X2 OR2X2_4657 ( .A(u2__abc_52155_new_n20618_), .B(sqrto_129_), .Y(u2__abc_52155_new_n20629_));
OR2X2 OR2X2_4658 ( .A(u2__abc_52155_new_n20632_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20633_));
OR2X2 OR2X2_4659 ( .A(u2__abc_52155_new_n20637_), .B(u2__abc_52155_new_n20628_), .Y(u2__abc_52155_new_n20638_));
OR2X2 OR2X2_466 ( .A(_abc_73687_new_n753_), .B(\a[116] ), .Y(_abc_73687_new_n1559_));
OR2X2 OR2X2_4660 ( .A(u2__abc_52155_new_n20630_), .B(sqrto_130_), .Y(u2__abc_52155_new_n20641_));
OR2X2 OR2X2_4661 ( .A(u2__abc_52155_new_n20644_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20645_));
OR2X2 OR2X2_4662 ( .A(u2__abc_52155_new_n20649_), .B(u2__abc_52155_new_n20640_), .Y(u2__abc_52155_new_n20650_));
OR2X2 OR2X2_4663 ( .A(u2__abc_52155_new_n20642_), .B(sqrto_131_), .Y(u2__abc_52155_new_n20653_));
OR2X2 OR2X2_4664 ( .A(u2__abc_52155_new_n20656_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20657_));
OR2X2 OR2X2_4665 ( .A(u2__abc_52155_new_n20661_), .B(u2__abc_52155_new_n20652_), .Y(u2__abc_52155_new_n20662_));
OR2X2 OR2X2_4666 ( .A(u2__abc_52155_new_n20654_), .B(sqrto_132_), .Y(u2__abc_52155_new_n20665_));
OR2X2 OR2X2_4667 ( .A(u2__abc_52155_new_n20668_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20669_));
OR2X2 OR2X2_4668 ( .A(u2__abc_52155_new_n20673_), .B(u2__abc_52155_new_n20664_), .Y(u2__abc_52155_new_n20674_));
OR2X2 OR2X2_4669 ( .A(u2__abc_52155_new_n20666_), .B(sqrto_133_), .Y(u2__abc_52155_new_n20677_));
OR2X2 OR2X2_467 ( .A(_abc_73687_new_n1565_), .B(_abc_73687_new_n1562_), .Y(_abc_73687_new_n1566_));
OR2X2 OR2X2_4670 ( .A(u2__abc_52155_new_n20680_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20681_));
OR2X2 OR2X2_4671 ( .A(u2__abc_52155_new_n20685_), .B(u2__abc_52155_new_n20676_), .Y(u2__abc_52155_new_n20686_));
OR2X2 OR2X2_4672 ( .A(u2__abc_52155_new_n20678_), .B(sqrto_134_), .Y(u2__abc_52155_new_n20689_));
OR2X2 OR2X2_4673 ( .A(u2__abc_52155_new_n20692_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20693_));
OR2X2 OR2X2_4674 ( .A(u2__abc_52155_new_n20697_), .B(u2__abc_52155_new_n20688_), .Y(u2__abc_52155_new_n20698_));
OR2X2 OR2X2_4675 ( .A(u2__abc_52155_new_n20690_), .B(sqrto_135_), .Y(u2__abc_52155_new_n20703_));
OR2X2 OR2X2_4676 ( .A(u2__abc_52155_new_n20704_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20705_));
OR2X2 OR2X2_4677 ( .A(u2__abc_52155_new_n20709_), .B(u2__abc_52155_new_n20700_), .Y(u2__abc_52155_new_n20710_));
OR2X2 OR2X2_4678 ( .A(u2__abc_52155_new_n20701_), .B(sqrto_136_), .Y(u2__abc_52155_new_n20713_));
OR2X2 OR2X2_4679 ( .A(u2__abc_52155_new_n20716_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20717_));
OR2X2 OR2X2_468 ( .A(_abc_73687_new_n1570_), .B(_abc_73687_new_n1567_), .Y(_abc_73687_new_n1571_));
OR2X2 OR2X2_4680 ( .A(u2__abc_52155_new_n20721_), .B(u2__abc_52155_new_n20712_), .Y(u2__abc_52155_new_n20722_));
OR2X2 OR2X2_4681 ( .A(u2__abc_52155_new_n20714_), .B(sqrto_137_), .Y(u2__abc_52155_new_n20725_));
OR2X2 OR2X2_4682 ( .A(u2__abc_52155_new_n20728_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20729_));
OR2X2 OR2X2_4683 ( .A(u2__abc_52155_new_n20733_), .B(u2__abc_52155_new_n20724_), .Y(u2__abc_52155_new_n20734_));
OR2X2 OR2X2_4684 ( .A(u2__abc_52155_new_n20726_), .B(sqrto_138_), .Y(u2__abc_52155_new_n20737_));
OR2X2 OR2X2_4685 ( .A(u2__abc_52155_new_n20740_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20741_));
OR2X2 OR2X2_4686 ( .A(u2__abc_52155_new_n20745_), .B(u2__abc_52155_new_n20736_), .Y(u2__abc_52155_new_n20746_));
OR2X2 OR2X2_4687 ( .A(u2__abc_52155_new_n20738_), .B(sqrto_139_), .Y(u2__abc_52155_new_n20751_));
OR2X2 OR2X2_4688 ( .A(u2__abc_52155_new_n20752_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20753_));
OR2X2 OR2X2_4689 ( .A(u2__abc_52155_new_n20757_), .B(u2__abc_52155_new_n20748_), .Y(u2__abc_52155_new_n20758_));
OR2X2 OR2X2_469 ( .A(_abc_73687_new_n1572_), .B(_abc_73687_new_n1561_), .Y(\o[231] ));
OR2X2 OR2X2_4690 ( .A(u2__abc_52155_new_n20749_), .B(sqrto_140_), .Y(u2__abc_52155_new_n20761_));
OR2X2 OR2X2_4691 ( .A(u2__abc_52155_new_n20764_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20765_));
OR2X2 OR2X2_4692 ( .A(u2__abc_52155_new_n20769_), .B(u2__abc_52155_new_n20760_), .Y(u2__abc_52155_new_n20770_));
OR2X2 OR2X2_4693 ( .A(u2__abc_52155_new_n20762_), .B(sqrto_141_), .Y(u2__abc_52155_new_n20775_));
OR2X2 OR2X2_4694 ( .A(u2__abc_52155_new_n20776_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20777_));
OR2X2 OR2X2_4695 ( .A(u2__abc_52155_new_n20781_), .B(u2__abc_52155_new_n20772_), .Y(u2__abc_52155_new_n20782_));
OR2X2 OR2X2_4696 ( .A(u2__abc_52155_new_n20773_), .B(sqrto_142_), .Y(u2__abc_52155_new_n20785_));
OR2X2 OR2X2_4697 ( .A(u2__abc_52155_new_n20788_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20789_));
OR2X2 OR2X2_4698 ( .A(u2__abc_52155_new_n20793_), .B(u2__abc_52155_new_n20784_), .Y(u2__abc_52155_new_n20794_));
OR2X2 OR2X2_4699 ( .A(u2__abc_52155_new_n20786_), .B(sqrto_143_), .Y(u2__abc_52155_new_n20797_));
OR2X2 OR2X2_47 ( .A(aNan), .B(sqrto_99_), .Y(_abc_73687_new_n899_));
OR2X2 OR2X2_470 ( .A(_abc_73687_new_n1577_), .B(_abc_73687_new_n1578_), .Y(_abc_73687_new_n1579_));
OR2X2 OR2X2_4700 ( .A(u2__abc_52155_new_n20800_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20801_));
OR2X2 OR2X2_4701 ( .A(u2__abc_52155_new_n20805_), .B(u2__abc_52155_new_n20796_), .Y(u2__abc_52155_new_n20806_));
OR2X2 OR2X2_4702 ( .A(u2__abc_52155_new_n20798_), .B(sqrto_144_), .Y(u2__abc_52155_new_n20809_));
OR2X2 OR2X2_4703 ( .A(u2__abc_52155_new_n20812_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20813_));
OR2X2 OR2X2_4704 ( .A(u2__abc_52155_new_n20817_), .B(u2__abc_52155_new_n20808_), .Y(u2__abc_52155_new_n20818_));
OR2X2 OR2X2_4705 ( .A(u2__abc_52155_new_n20810_), .B(sqrto_145_), .Y(u2__abc_52155_new_n20821_));
OR2X2 OR2X2_4706 ( .A(u2__abc_52155_new_n20824_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20825_));
OR2X2 OR2X2_4707 ( .A(u2__abc_52155_new_n20829_), .B(u2__abc_52155_new_n20820_), .Y(u2__abc_52155_new_n20830_));
OR2X2 OR2X2_4708 ( .A(u2__abc_52155_new_n20822_), .B(sqrto_146_), .Y(u2__abc_52155_new_n20833_));
OR2X2 OR2X2_4709 ( .A(u2__abc_52155_new_n20836_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20837_));
OR2X2 OR2X2_471 ( .A(_abc_73687_new_n1581_), .B(_abc_73687_new_n1582_), .Y(_abc_73687_new_n1583_));
OR2X2 OR2X2_4710 ( .A(u2__abc_52155_new_n20841_), .B(u2__abc_52155_new_n20832_), .Y(u2__abc_52155_new_n20842_));
OR2X2 OR2X2_4711 ( .A(u2__abc_52155_new_n20834_), .B(sqrto_147_), .Y(u2__abc_52155_new_n20847_));
OR2X2 OR2X2_4712 ( .A(u2__abc_52155_new_n20848_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20849_));
OR2X2 OR2X2_4713 ( .A(u2__abc_52155_new_n20853_), .B(u2__abc_52155_new_n20844_), .Y(u2__abc_52155_new_n20854_));
OR2X2 OR2X2_4714 ( .A(u2__abc_52155_new_n20845_), .B(sqrto_148_), .Y(u2__abc_52155_new_n20857_));
OR2X2 OR2X2_4715 ( .A(u2__abc_52155_new_n20860_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20861_));
OR2X2 OR2X2_4716 ( .A(u2__abc_52155_new_n20865_), .B(u2__abc_52155_new_n20856_), .Y(u2__abc_52155_new_n20866_));
OR2X2 OR2X2_4717 ( .A(u2__abc_52155_new_n20858_), .B(sqrto_149_), .Y(u2__abc_52155_new_n20871_));
OR2X2 OR2X2_4718 ( .A(u2__abc_52155_new_n20872_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20873_));
OR2X2 OR2X2_4719 ( .A(u2__abc_52155_new_n20877_), .B(u2__abc_52155_new_n20868_), .Y(u2__abc_52155_new_n20878_));
OR2X2 OR2X2_472 ( .A(_abc_73687_new_n1584_), .B(_abc_73687_new_n1585_), .Y(\o[232] ));
OR2X2 OR2X2_4720 ( .A(u2__abc_52155_new_n20869_), .B(sqrto_150_), .Y(u2__abc_52155_new_n20881_));
OR2X2 OR2X2_4721 ( .A(u2__abc_52155_new_n20884_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20885_));
OR2X2 OR2X2_4722 ( .A(u2__abc_52155_new_n20889_), .B(u2__abc_52155_new_n20880_), .Y(u2__abc_52155_new_n20890_));
OR2X2 OR2X2_4723 ( .A(u2__abc_52155_new_n20882_), .B(sqrto_151_), .Y(u2__abc_52155_new_n20893_));
OR2X2 OR2X2_4724 ( .A(u2__abc_52155_new_n20896_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20897_));
OR2X2 OR2X2_4725 ( .A(u2__abc_52155_new_n20901_), .B(u2__abc_52155_new_n20892_), .Y(u2__abc_52155_new_n20902_));
OR2X2 OR2X2_4726 ( .A(u2__abc_52155_new_n20894_), .B(sqrto_152_), .Y(u2__abc_52155_new_n20905_));
OR2X2 OR2X2_4727 ( .A(u2__abc_52155_new_n20908_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20909_));
OR2X2 OR2X2_4728 ( .A(u2__abc_52155_new_n20913_), .B(u2__abc_52155_new_n20904_), .Y(u2__abc_52155_new_n20914_));
OR2X2 OR2X2_4729 ( .A(u2__abc_52155_new_n20906_), .B(sqrto_153_), .Y(u2__abc_52155_new_n20919_));
OR2X2 OR2X2_473 ( .A(_abc_73687_new_n1591_), .B(_abc_73687_new_n1588_), .Y(_abc_73687_new_n1592_));
OR2X2 OR2X2_4730 ( .A(u2__abc_52155_new_n20920_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20921_));
OR2X2 OR2X2_4731 ( .A(u2__abc_52155_new_n20925_), .B(u2__abc_52155_new_n20916_), .Y(u2__abc_52155_new_n20926_));
OR2X2 OR2X2_4732 ( .A(u2__abc_52155_new_n20917_), .B(sqrto_154_), .Y(u2__abc_52155_new_n20929_));
OR2X2 OR2X2_4733 ( .A(u2__abc_52155_new_n20932_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20933_));
OR2X2 OR2X2_4734 ( .A(u2__abc_52155_new_n20937_), .B(u2__abc_52155_new_n20928_), .Y(u2__abc_52155_new_n20938_));
OR2X2 OR2X2_4735 ( .A(u2__abc_52155_new_n20930_), .B(sqrto_155_), .Y(u2__abc_52155_new_n20941_));
OR2X2 OR2X2_4736 ( .A(u2__abc_52155_new_n20944_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20945_));
OR2X2 OR2X2_4737 ( .A(u2__abc_52155_new_n20949_), .B(u2__abc_52155_new_n20940_), .Y(u2__abc_52155_new_n20950_));
OR2X2 OR2X2_4738 ( .A(u2__abc_52155_new_n20942_), .B(sqrto_156_), .Y(u2__abc_52155_new_n20953_));
OR2X2 OR2X2_4739 ( .A(u2__abc_52155_new_n20956_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20957_));
OR2X2 OR2X2_474 ( .A(_abc_73687_new_n1596_), .B(_abc_73687_new_n1593_), .Y(_abc_73687_new_n1597_));
OR2X2 OR2X2_4740 ( .A(u2__abc_52155_new_n20961_), .B(u2__abc_52155_new_n20952_), .Y(u2__abc_52155_new_n20962_));
OR2X2 OR2X2_4741 ( .A(u2__abc_52155_new_n20954_), .B(sqrto_157_), .Y(u2__abc_52155_new_n20967_));
OR2X2 OR2X2_4742 ( .A(u2__abc_52155_new_n20968_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20969_));
OR2X2 OR2X2_4743 ( .A(u2__abc_52155_new_n20973_), .B(u2__abc_52155_new_n20964_), .Y(u2__abc_52155_new_n20974_));
OR2X2 OR2X2_4744 ( .A(u2__abc_52155_new_n20965_), .B(sqrto_158_), .Y(u2__abc_52155_new_n20977_));
OR2X2 OR2X2_4745 ( .A(u2__abc_52155_new_n20980_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20981_));
OR2X2 OR2X2_4746 ( .A(u2__abc_52155_new_n20985_), .B(u2__abc_52155_new_n20976_), .Y(u2__abc_52155_new_n20986_));
OR2X2 OR2X2_4747 ( .A(u2__abc_52155_new_n20978_), .B(sqrto_159_), .Y(u2__abc_52155_new_n20989_));
OR2X2 OR2X2_4748 ( .A(u2__abc_52155_new_n20992_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n20993_));
OR2X2 OR2X2_4749 ( .A(u2__abc_52155_new_n20997_), .B(u2__abc_52155_new_n20988_), .Y(u2__abc_52155_new_n20998_));
OR2X2 OR2X2_475 ( .A(_abc_73687_new_n1598_), .B(_abc_73687_new_n1587_), .Y(\o[233] ));
OR2X2 OR2X2_4750 ( .A(u2__abc_52155_new_n20990_), .B(sqrto_160_), .Y(u2__abc_52155_new_n21001_));
OR2X2 OR2X2_4751 ( .A(u2__abc_52155_new_n21004_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21005_));
OR2X2 OR2X2_4752 ( .A(u2__abc_52155_new_n21009_), .B(u2__abc_52155_new_n21000_), .Y(u2__abc_52155_new_n21010_));
OR2X2 OR2X2_4753 ( .A(u2__abc_52155_new_n21002_), .B(sqrto_161_), .Y(u2__abc_52155_new_n21013_));
OR2X2 OR2X2_4754 ( .A(u2__abc_52155_new_n21016_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21017_));
OR2X2 OR2X2_4755 ( .A(u2__abc_52155_new_n21021_), .B(u2__abc_52155_new_n21012_), .Y(u2__abc_52155_new_n21022_));
OR2X2 OR2X2_4756 ( .A(u2__abc_52155_new_n21014_), .B(sqrto_162_), .Y(u2__abc_52155_new_n21025_));
OR2X2 OR2X2_4757 ( .A(u2__abc_52155_new_n21028_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21029_));
OR2X2 OR2X2_4758 ( .A(u2__abc_52155_new_n21033_), .B(u2__abc_52155_new_n21024_), .Y(u2__abc_52155_new_n21034_));
OR2X2 OR2X2_4759 ( .A(u2__abc_52155_new_n21026_), .B(sqrto_163_), .Y(u2__abc_52155_new_n21039_));
OR2X2 OR2X2_476 ( .A(_abc_73687_new_n1603_), .B(_abc_73687_new_n1600_), .Y(_abc_73687_new_n1604_));
OR2X2 OR2X2_4760 ( .A(u2__abc_52155_new_n21040_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21041_));
OR2X2 OR2X2_4761 ( .A(u2__abc_52155_new_n21045_), .B(u2__abc_52155_new_n21036_), .Y(u2__abc_52155_new_n21046_));
OR2X2 OR2X2_4762 ( .A(u2__abc_52155_new_n21037_), .B(sqrto_164_), .Y(u2__abc_52155_new_n21049_));
OR2X2 OR2X2_4763 ( .A(u2__abc_52155_new_n21052_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21053_));
OR2X2 OR2X2_4764 ( .A(u2__abc_52155_new_n21057_), .B(u2__abc_52155_new_n21048_), .Y(u2__abc_52155_new_n21058_));
OR2X2 OR2X2_4765 ( .A(u2__abc_52155_new_n21050_), .B(sqrto_165_), .Y(u2__abc_52155_new_n21063_));
OR2X2 OR2X2_4766 ( .A(u2__abc_52155_new_n21064_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21065_));
OR2X2 OR2X2_4767 ( .A(u2__abc_52155_new_n21069_), .B(u2__abc_52155_new_n21060_), .Y(u2__abc_52155_new_n21070_));
OR2X2 OR2X2_4768 ( .A(u2__abc_52155_new_n21061_), .B(sqrto_166_), .Y(u2__abc_52155_new_n21073_));
OR2X2 OR2X2_4769 ( .A(u2__abc_52155_new_n21076_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21077_));
OR2X2 OR2X2_477 ( .A(_abc_73687_new_n1608_), .B(_abc_73687_new_n1605_), .Y(_abc_73687_new_n1609_));
OR2X2 OR2X2_4770 ( .A(u2__abc_52155_new_n21081_), .B(u2__abc_52155_new_n21072_), .Y(u2__abc_52155_new_n21082_));
OR2X2 OR2X2_4771 ( .A(u2__abc_52155_new_n21074_), .B(sqrto_167_), .Y(u2__abc_52155_new_n21085_));
OR2X2 OR2X2_4772 ( .A(u2__abc_52155_new_n21088_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21089_));
OR2X2 OR2X2_4773 ( .A(u2__abc_52155_new_n21093_), .B(u2__abc_52155_new_n21084_), .Y(u2__abc_52155_new_n21094_));
OR2X2 OR2X2_4774 ( .A(u2__abc_52155_new_n21086_), .B(sqrto_168_), .Y(u2__abc_52155_new_n21097_));
OR2X2 OR2X2_4775 ( .A(u2__abc_52155_new_n21100_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21101_));
OR2X2 OR2X2_4776 ( .A(u2__abc_52155_new_n21105_), .B(u2__abc_52155_new_n21096_), .Y(u2__abc_52155_new_n21106_));
OR2X2 OR2X2_4777 ( .A(u2__abc_52155_new_n21098_), .B(sqrto_169_), .Y(u2__abc_52155_new_n21111_));
OR2X2 OR2X2_4778 ( .A(u2__abc_52155_new_n21112_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21113_));
OR2X2 OR2X2_4779 ( .A(u2__abc_52155_new_n21117_), .B(u2__abc_52155_new_n21108_), .Y(u2__abc_52155_new_n21118_));
OR2X2 OR2X2_478 ( .A(_abc_73687_new_n1610_), .B(_abc_73687_new_n1611_), .Y(\o[234] ));
OR2X2 OR2X2_4780 ( .A(u2__abc_52155_new_n21109_), .B(sqrto_170_), .Y(u2__abc_52155_new_n21121_));
OR2X2 OR2X2_4781 ( .A(u2__abc_52155_new_n21124_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21125_));
OR2X2 OR2X2_4782 ( .A(u2__abc_52155_new_n21129_), .B(u2__abc_52155_new_n21120_), .Y(u2__abc_52155_new_n21130_));
OR2X2 OR2X2_4783 ( .A(u2__abc_52155_new_n21122_), .B(sqrto_171_), .Y(u2__abc_52155_new_n21133_));
OR2X2 OR2X2_4784 ( .A(u2__abc_52155_new_n21136_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21137_));
OR2X2 OR2X2_4785 ( .A(u2__abc_52155_new_n21141_), .B(u2__abc_52155_new_n21132_), .Y(u2__abc_52155_new_n21142_));
OR2X2 OR2X2_4786 ( .A(u2__abc_52155_new_n21134_), .B(sqrto_172_), .Y(u2__abc_52155_new_n21145_));
OR2X2 OR2X2_4787 ( .A(u2__abc_52155_new_n21148_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21149_));
OR2X2 OR2X2_4788 ( .A(u2__abc_52155_new_n21153_), .B(u2__abc_52155_new_n21144_), .Y(u2__abc_52155_new_n21154_));
OR2X2 OR2X2_4789 ( .A(u2__abc_52155_new_n21146_), .B(sqrto_173_), .Y(u2__abc_52155_new_n21159_));
OR2X2 OR2X2_479 ( .A(_abc_73687_new_n1617_), .B(_abc_73687_new_n1614_), .Y(_abc_73687_new_n1618_));
OR2X2 OR2X2_4790 ( .A(u2__abc_52155_new_n21160_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21161_));
OR2X2 OR2X2_4791 ( .A(u2__abc_52155_new_n21165_), .B(u2__abc_52155_new_n21156_), .Y(u2__abc_52155_new_n21166_));
OR2X2 OR2X2_4792 ( .A(u2__abc_52155_new_n21157_), .B(sqrto_174_), .Y(u2__abc_52155_new_n21169_));
OR2X2 OR2X2_4793 ( .A(u2__abc_52155_new_n21172_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21173_));
OR2X2 OR2X2_4794 ( .A(u2__abc_52155_new_n21177_), .B(u2__abc_52155_new_n21168_), .Y(u2__abc_52155_new_n21178_));
OR2X2 OR2X2_4795 ( .A(u2__abc_52155_new_n21170_), .B(sqrto_175_), .Y(u2__abc_52155_new_n21181_));
OR2X2 OR2X2_4796 ( .A(u2__abc_52155_new_n21184_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21185_));
OR2X2 OR2X2_4797 ( .A(u2__abc_52155_new_n21189_), .B(u2__abc_52155_new_n21180_), .Y(u2__abc_52155_new_n21190_));
OR2X2 OR2X2_4798 ( .A(u2__abc_52155_new_n21182_), .B(sqrto_176_), .Y(u2__abc_52155_new_n21193_));
OR2X2 OR2X2_4799 ( .A(u2__abc_52155_new_n21196_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21197_));
OR2X2 OR2X2_48 ( .A(_abc_73687_new_n753_), .B(\a[23] ), .Y(_abc_73687_new_n900_));
OR2X2 OR2X2_480 ( .A(_abc_73687_new_n1622_), .B(_abc_73687_new_n1619_), .Y(_abc_73687_new_n1623_));
OR2X2 OR2X2_4800 ( .A(u2__abc_52155_new_n21201_), .B(u2__abc_52155_new_n21192_), .Y(u2__abc_52155_new_n21202_));
OR2X2 OR2X2_4801 ( .A(u2__abc_52155_new_n21194_), .B(sqrto_177_), .Y(u2__abc_52155_new_n21207_));
OR2X2 OR2X2_4802 ( .A(u2__abc_52155_new_n21208_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21209_));
OR2X2 OR2X2_4803 ( .A(u2__abc_52155_new_n21213_), .B(u2__abc_52155_new_n21204_), .Y(u2__abc_52155_new_n21214_));
OR2X2 OR2X2_4804 ( .A(u2__abc_52155_new_n21205_), .B(sqrto_178_), .Y(u2__abc_52155_new_n21217_));
OR2X2 OR2X2_4805 ( .A(u2__abc_52155_new_n21220_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21221_));
OR2X2 OR2X2_4806 ( .A(u2__abc_52155_new_n21225_), .B(u2__abc_52155_new_n21216_), .Y(u2__abc_52155_new_n21226_));
OR2X2 OR2X2_4807 ( .A(u2__abc_52155_new_n21218_), .B(sqrto_179_), .Y(u2__abc_52155_new_n21229_));
OR2X2 OR2X2_4808 ( .A(u2__abc_52155_new_n21232_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21233_));
OR2X2 OR2X2_4809 ( .A(u2__abc_52155_new_n21237_), .B(u2__abc_52155_new_n21228_), .Y(u2__abc_52155_new_n21238_));
OR2X2 OR2X2_481 ( .A(_abc_73687_new_n1624_), .B(_abc_73687_new_n1613_), .Y(\o[235] ));
OR2X2 OR2X2_4810 ( .A(u2__abc_52155_new_n21230_), .B(sqrto_180_), .Y(u2__abc_52155_new_n21241_));
OR2X2 OR2X2_4811 ( .A(u2__abc_52155_new_n21244_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21245_));
OR2X2 OR2X2_4812 ( .A(u2__abc_52155_new_n21249_), .B(u2__abc_52155_new_n21240_), .Y(u2__abc_52155_new_n21250_));
OR2X2 OR2X2_4813 ( .A(u2__abc_52155_new_n21242_), .B(sqrto_181_), .Y(u2__abc_52155_new_n21255_));
OR2X2 OR2X2_4814 ( .A(u2__abc_52155_new_n21256_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21257_));
OR2X2 OR2X2_4815 ( .A(u2__abc_52155_new_n21261_), .B(u2__abc_52155_new_n21252_), .Y(u2__abc_52155_new_n21262_));
OR2X2 OR2X2_4816 ( .A(u2__abc_52155_new_n21253_), .B(sqrto_182_), .Y(u2__abc_52155_new_n21265_));
OR2X2 OR2X2_4817 ( .A(u2__abc_52155_new_n21268_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21269_));
OR2X2 OR2X2_4818 ( .A(u2__abc_52155_new_n21273_), .B(u2__abc_52155_new_n21264_), .Y(u2__abc_52155_new_n21274_));
OR2X2 OR2X2_4819 ( .A(u2__abc_52155_new_n21266_), .B(sqrto_183_), .Y(u2__abc_52155_new_n21277_));
OR2X2 OR2X2_482 ( .A(_abc_73687_new_n1632_), .B(_abc_73687_new_n1633_), .Y(_abc_73687_new_n1634_));
OR2X2 OR2X2_4820 ( .A(u2__abc_52155_new_n21280_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21281_));
OR2X2 OR2X2_4821 ( .A(u2__abc_52155_new_n21285_), .B(u2__abc_52155_new_n21276_), .Y(u2__abc_52155_new_n21286_));
OR2X2 OR2X2_4822 ( .A(u2__abc_52155_new_n21278_), .B(sqrto_184_), .Y(u2__abc_52155_new_n21289_));
OR2X2 OR2X2_4823 ( .A(u2__abc_52155_new_n21292_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21293_));
OR2X2 OR2X2_4824 ( .A(u2__abc_52155_new_n21297_), .B(u2__abc_52155_new_n21288_), .Y(u2__abc_52155_new_n21298_));
OR2X2 OR2X2_4825 ( .A(u2__abc_52155_new_n21290_), .B(sqrto_185_), .Y(u2__abc_52155_new_n21303_));
OR2X2 OR2X2_4826 ( .A(u2__abc_52155_new_n21304_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21305_));
OR2X2 OR2X2_4827 ( .A(u2__abc_52155_new_n21309_), .B(u2__abc_52155_new_n21300_), .Y(u2__abc_52155_new_n21310_));
OR2X2 OR2X2_4828 ( .A(u2__abc_52155_new_n21301_), .B(sqrto_186_), .Y(u2__abc_52155_new_n21313_));
OR2X2 OR2X2_4829 ( .A(u2__abc_52155_new_n21316_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21317_));
OR2X2 OR2X2_483 ( .A(_abc_73687_new_n1636_), .B(_abc_73687_new_n1637_), .Y(_abc_73687_new_n1638_));
OR2X2 OR2X2_4830 ( .A(u2__abc_52155_new_n21321_), .B(u2__abc_52155_new_n21312_), .Y(u2__abc_52155_new_n21322_));
OR2X2 OR2X2_4831 ( .A(u2__abc_52155_new_n21314_), .B(sqrto_187_), .Y(u2__abc_52155_new_n21325_));
OR2X2 OR2X2_4832 ( .A(u2__abc_52155_new_n21328_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21329_));
OR2X2 OR2X2_4833 ( .A(u2__abc_52155_new_n21333_), .B(u2__abc_52155_new_n21324_), .Y(u2__abc_52155_new_n21334_));
OR2X2 OR2X2_4834 ( .A(u2__abc_52155_new_n21326_), .B(sqrto_188_), .Y(u2__abc_52155_new_n21337_));
OR2X2 OR2X2_4835 ( .A(u2__abc_52155_new_n21340_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21341_));
OR2X2 OR2X2_4836 ( .A(u2__abc_52155_new_n21345_), .B(u2__abc_52155_new_n21336_), .Y(u2__abc_52155_new_n21346_));
OR2X2 OR2X2_4837 ( .A(u2__abc_52155_new_n21338_), .B(sqrto_189_), .Y(u2__abc_52155_new_n21351_));
OR2X2 OR2X2_4838 ( .A(u2__abc_52155_new_n21352_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21353_));
OR2X2 OR2X2_4839 ( .A(u2__abc_52155_new_n21357_), .B(u2__abc_52155_new_n21348_), .Y(u2__abc_52155_new_n21358_));
OR2X2 OR2X2_484 ( .A(_abc_73687_new_n1639_), .B(_abc_73687_new_n1640_), .Y(\o[236] ));
OR2X2 OR2X2_4840 ( .A(u2__abc_52155_new_n21349_), .B(sqrto_190_), .Y(u2__abc_52155_new_n21361_));
OR2X2 OR2X2_4841 ( .A(u2__abc_52155_new_n21364_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21365_));
OR2X2 OR2X2_4842 ( .A(u2__abc_52155_new_n21369_), .B(u2__abc_52155_new_n21360_), .Y(u2__abc_52155_new_n21370_));
OR2X2 OR2X2_4843 ( .A(u2__abc_52155_new_n21362_), .B(sqrto_191_), .Y(u2__abc_52155_new_n21375_));
OR2X2 OR2X2_4844 ( .A(u2__abc_52155_new_n21376_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21377_));
OR2X2 OR2X2_4845 ( .A(u2__abc_52155_new_n21381_), .B(u2__abc_52155_new_n21372_), .Y(u2__abc_52155_new_n21382_));
OR2X2 OR2X2_4846 ( .A(u2__abc_52155_new_n21373_), .B(sqrto_192_), .Y(u2__abc_52155_new_n21385_));
OR2X2 OR2X2_4847 ( .A(u2__abc_52155_new_n21388_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21389_));
OR2X2 OR2X2_4848 ( .A(u2__abc_52155_new_n21393_), .B(u2__abc_52155_new_n21384_), .Y(u2__abc_52155_new_n21394_));
OR2X2 OR2X2_4849 ( .A(u2__abc_52155_new_n21386_), .B(sqrto_193_), .Y(u2__abc_52155_new_n21397_));
OR2X2 OR2X2_485 ( .A(_abc_73687_new_n1633_), .B(_abc_73687_new_n1643_), .Y(_abc_73687_new_n1646_));
OR2X2 OR2X2_4850 ( .A(u2__abc_52155_new_n21400_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21401_));
OR2X2 OR2X2_4851 ( .A(u2__abc_52155_new_n21405_), .B(u2__abc_52155_new_n21396_), .Y(u2__abc_52155_new_n21406_));
OR2X2 OR2X2_4852 ( .A(u2__abc_52155_new_n21398_), .B(sqrto_194_), .Y(u2__abc_52155_new_n21409_));
OR2X2 OR2X2_4853 ( .A(u2__abc_52155_new_n21412_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21413_));
OR2X2 OR2X2_4854 ( .A(u2__abc_52155_new_n21417_), .B(u2__abc_52155_new_n21408_), .Y(u2__abc_52155_new_n21418_));
OR2X2 OR2X2_4855 ( .A(u2__abc_52155_new_n21410_), .B(sqrto_195_), .Y(u2__abc_52155_new_n21423_));
OR2X2 OR2X2_4856 ( .A(u2__abc_52155_new_n21424_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21425_));
OR2X2 OR2X2_4857 ( .A(u2__abc_52155_new_n21429_), .B(u2__abc_52155_new_n21420_), .Y(u2__abc_52155_new_n21430_));
OR2X2 OR2X2_4858 ( .A(u2__abc_52155_new_n21421_), .B(sqrto_196_), .Y(u2__abc_52155_new_n21433_));
OR2X2 OR2X2_4859 ( .A(u2__abc_52155_new_n21436_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21437_));
OR2X2 OR2X2_486 ( .A(_abc_73687_new_n1651_), .B(_abc_73687_new_n1648_), .Y(_abc_73687_new_n1652_));
OR2X2 OR2X2_4860 ( .A(u2__abc_52155_new_n21441_), .B(u2__abc_52155_new_n21432_), .Y(u2__abc_52155_new_n21442_));
OR2X2 OR2X2_4861 ( .A(u2__abc_52155_new_n21434_), .B(sqrto_197_), .Y(u2__abc_52155_new_n21447_));
OR2X2 OR2X2_4862 ( .A(u2__abc_52155_new_n21448_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21449_));
OR2X2 OR2X2_4863 ( .A(u2__abc_52155_new_n21453_), .B(u2__abc_52155_new_n21444_), .Y(u2__abc_52155_new_n21454_));
OR2X2 OR2X2_4864 ( .A(u2__abc_52155_new_n21445_), .B(sqrto_198_), .Y(u2__abc_52155_new_n21457_));
OR2X2 OR2X2_4865 ( .A(u2__abc_52155_new_n21460_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21461_));
OR2X2 OR2X2_4866 ( .A(u2__abc_52155_new_n21465_), .B(u2__abc_52155_new_n21456_), .Y(u2__abc_52155_new_n21466_));
OR2X2 OR2X2_4867 ( .A(u2__abc_52155_new_n21458_), .B(sqrto_199_), .Y(u2__abc_52155_new_n21469_));
OR2X2 OR2X2_4868 ( .A(u2__abc_52155_new_n21472_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21473_));
OR2X2 OR2X2_4869 ( .A(u2__abc_52155_new_n21477_), .B(u2__abc_52155_new_n21468_), .Y(u2__abc_52155_new_n21478_));
OR2X2 OR2X2_487 ( .A(_abc_73687_new_n1653_), .B(_abc_73687_new_n1642_), .Y(\o[237] ));
OR2X2 OR2X2_4870 ( .A(u2__abc_52155_new_n21470_), .B(sqrto_200_), .Y(u2__abc_52155_new_n21481_));
OR2X2 OR2X2_4871 ( .A(u2__abc_52155_new_n21484_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21485_));
OR2X2 OR2X2_4872 ( .A(u2__abc_52155_new_n21489_), .B(u2__abc_52155_new_n21480_), .Y(u2__abc_52155_new_n21490_));
OR2X2 OR2X2_4873 ( .A(u2__abc_52155_new_n21482_), .B(sqrto_201_), .Y(u2__abc_52155_new_n21495_));
OR2X2 OR2X2_4874 ( .A(u2__abc_52155_new_n21496_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21497_));
OR2X2 OR2X2_4875 ( .A(u2__abc_52155_new_n21501_), .B(u2__abc_52155_new_n21492_), .Y(u2__abc_52155_new_n21502_));
OR2X2 OR2X2_4876 ( .A(u2__abc_52155_new_n21493_), .B(sqrto_202_), .Y(u2__abc_52155_new_n21505_));
OR2X2 OR2X2_4877 ( .A(u2__abc_52155_new_n21508_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21509_));
OR2X2 OR2X2_4878 ( .A(u2__abc_52155_new_n21513_), .B(u2__abc_52155_new_n21504_), .Y(u2__abc_52155_new_n21514_));
OR2X2 OR2X2_4879 ( .A(u2__abc_52155_new_n21506_), .B(sqrto_203_), .Y(u2__abc_52155_new_n21517_));
OR2X2 OR2X2_488 ( .A(_abc_73687_new_n1659_), .B(_abc_73687_new_n1660_), .Y(_abc_73687_new_n1661_));
OR2X2 OR2X2_4880 ( .A(u2__abc_52155_new_n21520_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21521_));
OR2X2 OR2X2_4881 ( .A(u2__abc_52155_new_n21525_), .B(u2__abc_52155_new_n21516_), .Y(u2__abc_52155_new_n21526_));
OR2X2 OR2X2_4882 ( .A(u2__abc_52155_new_n21518_), .B(sqrto_204_), .Y(u2__abc_52155_new_n21529_));
OR2X2 OR2X2_4883 ( .A(u2__abc_52155_new_n21532_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21533_));
OR2X2 OR2X2_4884 ( .A(u2__abc_52155_new_n21537_), .B(u2__abc_52155_new_n21528_), .Y(u2__abc_52155_new_n21538_));
OR2X2 OR2X2_4885 ( .A(u2__abc_52155_new_n21530_), .B(sqrto_205_), .Y(u2__abc_52155_new_n21543_));
OR2X2 OR2X2_4886 ( .A(u2__abc_52155_new_n21544_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21545_));
OR2X2 OR2X2_4887 ( .A(u2__abc_52155_new_n21549_), .B(u2__abc_52155_new_n21540_), .Y(u2__abc_52155_new_n21550_));
OR2X2 OR2X2_4888 ( .A(u2__abc_52155_new_n21541_), .B(sqrto_206_), .Y(u2__abc_52155_new_n21553_));
OR2X2 OR2X2_4889 ( .A(u2__abc_52155_new_n21556_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21557_));
OR2X2 OR2X2_489 ( .A(_abc_73687_new_n1663_), .B(_abc_73687_new_n1664_), .Y(_abc_73687_new_n1665_));
OR2X2 OR2X2_4890 ( .A(u2__abc_52155_new_n21561_), .B(u2__abc_52155_new_n21552_), .Y(u2__abc_52155_new_n21562_));
OR2X2 OR2X2_4891 ( .A(u2__abc_52155_new_n21554_), .B(sqrto_207_), .Y(u2__abc_52155_new_n21565_));
OR2X2 OR2X2_4892 ( .A(u2__abc_52155_new_n21568_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21569_));
OR2X2 OR2X2_4893 ( .A(u2__abc_52155_new_n21573_), .B(u2__abc_52155_new_n21564_), .Y(u2__abc_52155_new_n21574_));
OR2X2 OR2X2_4894 ( .A(u2__abc_52155_new_n21566_), .B(sqrto_208_), .Y(u2__abc_52155_new_n21577_));
OR2X2 OR2X2_4895 ( .A(u2__abc_52155_new_n21580_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21581_));
OR2X2 OR2X2_4896 ( .A(u2__abc_52155_new_n21585_), .B(u2__abc_52155_new_n21576_), .Y(u2__abc_52155_new_n21586_));
OR2X2 OR2X2_4897 ( .A(u2__abc_52155_new_n21578_), .B(sqrto_209_), .Y(u2__abc_52155_new_n21591_));
OR2X2 OR2X2_4898 ( .A(u2__abc_52155_new_n21592_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21593_));
OR2X2 OR2X2_4899 ( .A(u2__abc_52155_new_n21597_), .B(u2__abc_52155_new_n21588_), .Y(u2__abc_52155_new_n21598_));
OR2X2 OR2X2_49 ( .A(aNan), .B(sqrto_100_), .Y(_abc_73687_new_n902_));
OR2X2 OR2X2_490 ( .A(_abc_73687_new_n1666_), .B(_abc_73687_new_n1667_), .Y(\o[238] ));
OR2X2 OR2X2_4900 ( .A(u2__abc_52155_new_n21589_), .B(sqrto_210_), .Y(u2__abc_52155_new_n21601_));
OR2X2 OR2X2_4901 ( .A(u2__abc_52155_new_n21604_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21605_));
OR2X2 OR2X2_4902 ( .A(u2__abc_52155_new_n21609_), .B(u2__abc_52155_new_n21600_), .Y(u2__abc_52155_new_n21610_));
OR2X2 OR2X2_4903 ( .A(u2__abc_52155_new_n21602_), .B(sqrto_211_), .Y(u2__abc_52155_new_n21613_));
OR2X2 OR2X2_4904 ( .A(u2__abc_52155_new_n21616_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21617_));
OR2X2 OR2X2_4905 ( .A(u2__abc_52155_new_n21621_), .B(u2__abc_52155_new_n21612_), .Y(u2__abc_52155_new_n21622_));
OR2X2 OR2X2_4906 ( .A(u2__abc_52155_new_n21614_), .B(sqrto_212_), .Y(u2__abc_52155_new_n21625_));
OR2X2 OR2X2_4907 ( .A(u2__abc_52155_new_n21628_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21629_));
OR2X2 OR2X2_4908 ( .A(u2__abc_52155_new_n21633_), .B(u2__abc_52155_new_n21624_), .Y(u2__abc_52155_new_n21634_));
OR2X2 OR2X2_4909 ( .A(u2__abc_52155_new_n21626_), .B(sqrto_213_), .Y(u2__abc_52155_new_n21639_));
OR2X2 OR2X2_491 ( .A(_abc_73687_new_n753_), .B(\a[125] ), .Y(_abc_73687_new_n1669_));
OR2X2 OR2X2_4910 ( .A(u2__abc_52155_new_n21640_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21641_));
OR2X2 OR2X2_4911 ( .A(u2__abc_52155_new_n21645_), .B(u2__abc_52155_new_n21636_), .Y(u2__abc_52155_new_n21646_));
OR2X2 OR2X2_4912 ( .A(u2__abc_52155_new_n21637_), .B(sqrto_214_), .Y(u2__abc_52155_new_n21649_));
OR2X2 OR2X2_4913 ( .A(u2__abc_52155_new_n21652_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21653_));
OR2X2 OR2X2_4914 ( .A(u2__abc_52155_new_n21657_), .B(u2__abc_52155_new_n21648_), .Y(u2__abc_52155_new_n21658_));
OR2X2 OR2X2_4915 ( .A(u2__abc_52155_new_n21650_), .B(sqrto_215_), .Y(u2__abc_52155_new_n21661_));
OR2X2 OR2X2_4916 ( .A(u2__abc_52155_new_n21664_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21665_));
OR2X2 OR2X2_4917 ( .A(u2__abc_52155_new_n21669_), .B(u2__abc_52155_new_n21660_), .Y(u2__abc_52155_new_n21670_));
OR2X2 OR2X2_4918 ( .A(u2__abc_52155_new_n21662_), .B(sqrto_216_), .Y(u2__abc_52155_new_n21673_));
OR2X2 OR2X2_4919 ( .A(u2__abc_52155_new_n21676_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21677_));
OR2X2 OR2X2_492 ( .A(_abc_73687_new_n1660_), .B(_abc_73687_new_n1670_), .Y(_abc_73687_new_n1671_));
OR2X2 OR2X2_4920 ( .A(u2__abc_52155_new_n21681_), .B(u2__abc_52155_new_n21672_), .Y(u2__abc_52155_new_n21682_));
OR2X2 OR2X2_4921 ( .A(u2__abc_52155_new_n21674_), .B(sqrto_217_), .Y(u2__abc_52155_new_n21687_));
OR2X2 OR2X2_4922 ( .A(u2__abc_52155_new_n21688_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21689_));
OR2X2 OR2X2_4923 ( .A(u2__abc_52155_new_n21693_), .B(u2__abc_52155_new_n21684_), .Y(u2__abc_52155_new_n21694_));
OR2X2 OR2X2_4924 ( .A(u2__abc_52155_new_n21685_), .B(sqrto_218_), .Y(u2__abc_52155_new_n21697_));
OR2X2 OR2X2_4925 ( .A(u2__abc_52155_new_n21700_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21701_));
OR2X2 OR2X2_4926 ( .A(u2__abc_52155_new_n21705_), .B(u2__abc_52155_new_n21696_), .Y(u2__abc_52155_new_n21706_));
OR2X2 OR2X2_4927 ( .A(u2__abc_52155_new_n21698_), .B(sqrto_219_), .Y(u2__abc_52155_new_n21709_));
OR2X2 OR2X2_4928 ( .A(u2__abc_52155_new_n21712_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21713_));
OR2X2 OR2X2_4929 ( .A(u2__abc_52155_new_n21717_), .B(u2__abc_52155_new_n21708_), .Y(u2__abc_52155_new_n21718_));
OR2X2 OR2X2_493 ( .A(_abc_73687_new_n1664_), .B(_abc_73687_new_n1674_), .Y(_abc_73687_new_n1675_));
OR2X2 OR2X2_4930 ( .A(u2__abc_52155_new_n21710_), .B(sqrto_220_), .Y(u2__abc_52155_new_n21721_));
OR2X2 OR2X2_4931 ( .A(u2__abc_52155_new_n21724_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21725_));
OR2X2 OR2X2_4932 ( .A(u2__abc_52155_new_n21729_), .B(u2__abc_52155_new_n21720_), .Y(u2__abc_52155_new_n21730_));
OR2X2 OR2X2_4933 ( .A(u2__abc_52155_new_n21722_), .B(sqrto_221_), .Y(u2__abc_52155_new_n21735_));
OR2X2 OR2X2_4934 ( .A(u2__abc_52155_new_n21736_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21737_));
OR2X2 OR2X2_4935 ( .A(u2__abc_52155_new_n21741_), .B(u2__abc_52155_new_n21732_), .Y(u2__abc_52155_new_n21742_));
OR2X2 OR2X2_4936 ( .A(u2__abc_52155_new_n21733_), .B(sqrto_222_), .Y(u2__abc_52155_new_n21745_));
OR2X2 OR2X2_4937 ( .A(u2__abc_52155_new_n21748_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21749_));
OR2X2 OR2X2_4938 ( .A(u2__abc_52155_new_n21753_), .B(u2__abc_52155_new_n21744_), .Y(u2__abc_52155_new_n21754_));
OR2X2 OR2X2_4939 ( .A(u2__abc_52155_new_n21746_), .B(sqrto_223_), .Y(u2__abc_52155_new_n21759_));
OR2X2 OR2X2_494 ( .A(_abc_73687_new_n1678_), .B(aNan), .Y(_abc_73687_new_n1679_));
OR2X2 OR2X2_4940 ( .A(u2__abc_52155_new_n21760_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21761_));
OR2X2 OR2X2_4941 ( .A(u2__abc_52155_new_n21765_), .B(u2__abc_52155_new_n21756_), .Y(u2__abc_52155_new_n21766_));
OR2X2 OR2X2_4942 ( .A(u2__abc_52155_new_n21757_), .B(sqrto_224_), .Y(u2__abc_52155_new_n21769_));
OR2X2 OR2X2_4943 ( .A(u2__abc_52155_new_n21772_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21773_));
OR2X2 OR2X2_4944 ( .A(u2__abc_52155_new_n21777_), .B(u2__abc_52155_new_n21768_), .Y(u2__abc_52155_new_n21778_));
OR2X2 OR2X2_4945 ( .A(u2__abc_52155_new_n21770_), .B(sqrto_225_), .Y(u2__abc_52155_new_n21783_));
OR2X2 OR2X2_4946 ( .A(u2__abc_52155_new_n21784_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21785_));
OR2X2 OR2X2_4947 ( .A(u2__abc_52155_new_n21789_), .B(u2__abc_52155_new_n21780_), .Y(u2__abc_52155_new_n21790_));
OR2X2 OR2X2_4948 ( .A(u2__abc_52155_new_n21781_), .B(u2_o_226_), .Y(u2__abc_52155_new_n21793_));
OR2X2 OR2X2_4949 ( .A(u2__abc_52155_new_n21796_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21797_));
OR2X2 OR2X2_495 ( .A(_abc_73687_new_n1683_), .B(aNan), .Y(_abc_73687_new_n1684_));
OR2X2 OR2X2_4950 ( .A(u2__abc_52155_new_n21801_), .B(u2__abc_52155_new_n21792_), .Y(u2__abc_52155_new_n21802_));
OR2X2 OR2X2_4951 ( .A(u2__abc_52155_new_n21794_), .B(u2_o_227_), .Y(u2__abc_52155_new_n21805_));
OR2X2 OR2X2_4952 ( .A(u2__abc_52155_new_n21808_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21809_));
OR2X2 OR2X2_4953 ( .A(u2__abc_52155_new_n21813_), .B(u2__abc_52155_new_n21804_), .Y(u2__abc_52155_new_n21814_));
OR2X2 OR2X2_4954 ( .A(u2__abc_52155_new_n21806_), .B(u2_o_228_), .Y(u2__abc_52155_new_n21817_));
OR2X2 OR2X2_4955 ( .A(u2__abc_52155_new_n21820_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21821_));
OR2X2 OR2X2_4956 ( .A(u2__abc_52155_new_n21825_), .B(u2__abc_52155_new_n21816_), .Y(u2__abc_52155_new_n21826_));
OR2X2 OR2X2_4957 ( .A(u2__abc_52155_new_n21818_), .B(u2_o_229_), .Y(u2__abc_52155_new_n21831_));
OR2X2 OR2X2_4958 ( .A(u2__abc_52155_new_n21832_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21833_));
OR2X2 OR2X2_4959 ( .A(u2__abc_52155_new_n21837_), .B(u2__abc_52155_new_n21828_), .Y(u2__abc_52155_new_n21838_));
OR2X2 OR2X2_496 ( .A(_abc_73687_new_n1687_), .B(_abc_73687_new_n1685_), .Y(\o[240] ));
OR2X2 OR2X2_4960 ( .A(u2__abc_52155_new_n21829_), .B(u2_o_230_), .Y(u2__abc_52155_new_n21841_));
OR2X2 OR2X2_4961 ( .A(u2__abc_52155_new_n21844_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21845_));
OR2X2 OR2X2_4962 ( .A(u2__abc_52155_new_n21849_), .B(u2__abc_52155_new_n21840_), .Y(u2__abc_52155_new_n21850_));
OR2X2 OR2X2_4963 ( .A(u2__abc_52155_new_n21842_), .B(u2_o_231_), .Y(u2__abc_52155_new_n21853_));
OR2X2 OR2X2_4964 ( .A(u2__abc_52155_new_n21856_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21857_));
OR2X2 OR2X2_4965 ( .A(u2__abc_52155_new_n21861_), .B(u2__abc_52155_new_n21852_), .Y(u2__abc_52155_new_n21862_));
OR2X2 OR2X2_4966 ( .A(u2__abc_52155_new_n21854_), .B(u2_o_232_), .Y(u2__abc_52155_new_n21865_));
OR2X2 OR2X2_4967 ( .A(u2__abc_52155_new_n21868_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21869_));
OR2X2 OR2X2_4968 ( .A(u2__abc_52155_new_n21873_), .B(u2__abc_52155_new_n21864_), .Y(u2__abc_52155_new_n21874_));
OR2X2 OR2X2_4969 ( .A(u2__abc_52155_new_n21866_), .B(u2_o_233_), .Y(u2__abc_52155_new_n21879_));
OR2X2 OR2X2_497 ( .A(\a[121] ), .B(\a[122] ), .Y(u1__abc_51895_new_n137_));
OR2X2 OR2X2_4970 ( .A(u2__abc_52155_new_n21880_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21881_));
OR2X2 OR2X2_4971 ( .A(u2__abc_52155_new_n21885_), .B(u2__abc_52155_new_n21876_), .Y(u2__abc_52155_new_n21886_));
OR2X2 OR2X2_4972 ( .A(u2__abc_52155_new_n21877_), .B(u2_o_234_), .Y(u2__abc_52155_new_n21889_));
OR2X2 OR2X2_4973 ( .A(u2__abc_52155_new_n21892_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21893_));
OR2X2 OR2X2_4974 ( .A(u2__abc_52155_new_n21897_), .B(u2__abc_52155_new_n21888_), .Y(u2__abc_52155_new_n21898_));
OR2X2 OR2X2_4975 ( .A(u2__abc_52155_new_n21890_), .B(u2_o_235_), .Y(u2__abc_52155_new_n21901_));
OR2X2 OR2X2_4976 ( .A(u2__abc_52155_new_n21904_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21905_));
OR2X2 OR2X2_4977 ( .A(u2__abc_52155_new_n21909_), .B(u2__abc_52155_new_n21900_), .Y(u2__abc_52155_new_n21910_));
OR2X2 OR2X2_4978 ( .A(u2__abc_52155_new_n21902_), .B(u2_o_236_), .Y(u2__abc_52155_new_n21913_));
OR2X2 OR2X2_4979 ( .A(u2__abc_52155_new_n21916_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21917_));
OR2X2 OR2X2_498 ( .A(\a[119] ), .B(\a[120] ), .Y(u1__abc_51895_new_n138_));
OR2X2 OR2X2_4980 ( .A(u2__abc_52155_new_n21921_), .B(u2__abc_52155_new_n21912_), .Y(u2__abc_52155_new_n21922_));
OR2X2 OR2X2_4981 ( .A(u2__abc_52155_new_n21914_), .B(u2_o_237_), .Y(u2__abc_52155_new_n21927_));
OR2X2 OR2X2_4982 ( .A(u2__abc_52155_new_n21928_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21929_));
OR2X2 OR2X2_4983 ( .A(u2__abc_52155_new_n21933_), .B(u2__abc_52155_new_n21924_), .Y(u2__abc_52155_new_n21934_));
OR2X2 OR2X2_4984 ( .A(u2__abc_52155_new_n21925_), .B(u2_o_238_), .Y(u2__abc_52155_new_n21937_));
OR2X2 OR2X2_4985 ( .A(u2__abc_52155_new_n21940_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21941_));
OR2X2 OR2X2_4986 ( .A(u2__abc_52155_new_n21945_), .B(u2__abc_52155_new_n21936_), .Y(u2__abc_52155_new_n21946_));
OR2X2 OR2X2_4987 ( .A(u2__abc_52155_new_n21938_), .B(u2_o_239_), .Y(u2__abc_52155_new_n21951_));
OR2X2 OR2X2_4988 ( .A(u2__abc_52155_new_n21952_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21953_));
OR2X2 OR2X2_4989 ( .A(u2__abc_52155_new_n21957_), .B(u2__abc_52155_new_n21948_), .Y(u2__abc_52155_new_n21958_));
OR2X2 OR2X2_499 ( .A(u1__abc_51895_new_n137_), .B(u1__abc_51895_new_n138_), .Y(u1__abc_51895_new_n139_));
OR2X2 OR2X2_4990 ( .A(u2__abc_52155_new_n21949_), .B(u2_o_240_), .Y(u2__abc_52155_new_n21961_));
OR2X2 OR2X2_4991 ( .A(u2__abc_52155_new_n21964_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21965_));
OR2X2 OR2X2_4992 ( .A(u2__abc_52155_new_n21969_), .B(u2__abc_52155_new_n21960_), .Y(u2__abc_52155_new_n21970_));
OR2X2 OR2X2_4993 ( .A(u2__abc_52155_new_n21962_), .B(u2_o_241_), .Y(u2__abc_52155_new_n21975_));
OR2X2 OR2X2_4994 ( .A(u2__abc_52155_new_n21976_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21977_));
OR2X2 OR2X2_4995 ( .A(u2__abc_52155_new_n21981_), .B(u2__abc_52155_new_n21972_), .Y(u2__abc_52155_new_n21982_));
OR2X2 OR2X2_4996 ( .A(u2__abc_52155_new_n21973_), .B(u2_o_242_), .Y(u2__abc_52155_new_n21985_));
OR2X2 OR2X2_4997 ( .A(u2__abc_52155_new_n21988_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n21989_));
OR2X2 OR2X2_4998 ( .A(u2__abc_52155_new_n21993_), .B(u2__abc_52155_new_n21984_), .Y(u2__abc_52155_new_n21994_));
OR2X2 OR2X2_4999 ( .A(u2__abc_52155_new_n21986_), .B(u2_o_243_), .Y(u2__abc_52155_new_n21997_));
OR2X2 OR2X2_5 ( .A(aNan), .B(sqrto_78_), .Y(_abc_73687_new_n836_));
OR2X2 OR2X2_50 ( .A(_abc_73687_new_n753_), .B(\a[24] ), .Y(_abc_73687_new_n903_));
OR2X2 OR2X2_500 ( .A(\a[125] ), .B(\a[126] ), .Y(u1__abc_51895_new_n140_));
OR2X2 OR2X2_5000 ( .A(u2__abc_52155_new_n22000_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22001_));
OR2X2 OR2X2_5001 ( .A(u2__abc_52155_new_n22005_), .B(u2__abc_52155_new_n21996_), .Y(u2__abc_52155_new_n22006_));
OR2X2 OR2X2_5002 ( .A(u2__abc_52155_new_n21998_), .B(u2_o_244_), .Y(u2__abc_52155_new_n22009_));
OR2X2 OR2X2_5003 ( .A(u2__abc_52155_new_n22012_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22013_));
OR2X2 OR2X2_5004 ( .A(u2__abc_52155_new_n22017_), .B(u2__abc_52155_new_n22008_), .Y(u2__abc_52155_new_n22018_));
OR2X2 OR2X2_5005 ( .A(u2__abc_52155_new_n22010_), .B(u2_o_245_), .Y(u2__abc_52155_new_n22023_));
OR2X2 OR2X2_5006 ( .A(u2__abc_52155_new_n22024_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22025_));
OR2X2 OR2X2_5007 ( .A(u2__abc_52155_new_n22029_), .B(u2__abc_52155_new_n22020_), .Y(u2__abc_52155_new_n22030_));
OR2X2 OR2X2_5008 ( .A(u2__abc_52155_new_n22021_), .B(u2_o_246_), .Y(u2__abc_52155_new_n22033_));
OR2X2 OR2X2_5009 ( .A(u2__abc_52155_new_n22036_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22037_));
OR2X2 OR2X2_501 ( .A(\a[123] ), .B(\a[124] ), .Y(u1__abc_51895_new_n141_));
OR2X2 OR2X2_5010 ( .A(u2__abc_52155_new_n22041_), .B(u2__abc_52155_new_n22032_), .Y(u2__abc_52155_new_n22042_));
OR2X2 OR2X2_5011 ( .A(u2__abc_52155_new_n22034_), .B(u2_o_247_), .Y(u2__abc_52155_new_n22047_));
OR2X2 OR2X2_5012 ( .A(u2__abc_52155_new_n22048_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22049_));
OR2X2 OR2X2_5013 ( .A(u2__abc_52155_new_n22053_), .B(u2__abc_52155_new_n22044_), .Y(u2__abc_52155_new_n22054_));
OR2X2 OR2X2_5014 ( .A(u2__abc_52155_new_n22045_), .B(u2_o_248_), .Y(u2__abc_52155_new_n22057_));
OR2X2 OR2X2_5015 ( .A(u2__abc_52155_new_n22060_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22061_));
OR2X2 OR2X2_5016 ( .A(u2__abc_52155_new_n22065_), .B(u2__abc_52155_new_n22056_), .Y(u2__abc_52155_new_n22066_));
OR2X2 OR2X2_5017 ( .A(u2__abc_52155_new_n22058_), .B(u2_o_249_), .Y(u2__abc_52155_new_n22071_));
OR2X2 OR2X2_5018 ( .A(u2__abc_52155_new_n22072_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22073_));
OR2X2 OR2X2_5019 ( .A(u2__abc_52155_new_n22077_), .B(u2__abc_52155_new_n22068_), .Y(u2__abc_52155_new_n22078_));
OR2X2 OR2X2_502 ( .A(u1__abc_51895_new_n140_), .B(u1__abc_51895_new_n141_), .Y(u1__abc_51895_new_n142_));
OR2X2 OR2X2_5020 ( .A(u2__abc_52155_new_n22069_), .B(u2_o_250_), .Y(u2__abc_52155_new_n22081_));
OR2X2 OR2X2_5021 ( .A(u2__abc_52155_new_n22084_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22085_));
OR2X2 OR2X2_5022 ( .A(u2__abc_52155_new_n22089_), .B(u2__abc_52155_new_n22080_), .Y(u2__abc_52155_new_n22090_));
OR2X2 OR2X2_5023 ( .A(u2__abc_52155_new_n22082_), .B(u2_o_251_), .Y(u2__abc_52155_new_n22095_));
OR2X2 OR2X2_5024 ( .A(u2__abc_52155_new_n22096_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22097_));
OR2X2 OR2X2_5025 ( .A(u2__abc_52155_new_n22101_), .B(u2__abc_52155_new_n22092_), .Y(u2__abc_52155_new_n22102_));
OR2X2 OR2X2_5026 ( .A(u2__abc_52155_new_n22093_), .B(u2_o_252_), .Y(u2__abc_52155_new_n22105_));
OR2X2 OR2X2_5027 ( .A(u2__abc_52155_new_n22108_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22109_));
OR2X2 OR2X2_5028 ( .A(u2__abc_52155_new_n22113_), .B(u2__abc_52155_new_n22104_), .Y(u2__abc_52155_new_n22114_));
OR2X2 OR2X2_5029 ( .A(u2__abc_52155_new_n22106_), .B(u2_o_253_), .Y(u2__abc_52155_new_n22119_));
OR2X2 OR2X2_503 ( .A(u1__abc_51895_new_n139_), .B(u1__abc_51895_new_n142_), .Y(u1__abc_51895_new_n143_));
OR2X2 OR2X2_5030 ( .A(u2__abc_52155_new_n22120_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22121_));
OR2X2 OR2X2_5031 ( .A(u2__abc_52155_new_n22125_), .B(u2__abc_52155_new_n22116_), .Y(u2__abc_52155_new_n22126_));
OR2X2 OR2X2_5032 ( .A(u2__abc_52155_new_n22117_), .B(u2_o_254_), .Y(u2__abc_52155_new_n22129_));
OR2X2 OR2X2_5033 ( .A(u2__abc_52155_new_n22132_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22133_));
OR2X2 OR2X2_5034 ( .A(u2__abc_52155_new_n22137_), .B(u2__abc_52155_new_n22128_), .Y(u2__abc_52155_new_n22138_));
OR2X2 OR2X2_5035 ( .A(u2__abc_52155_new_n22130_), .B(u2_o_255_), .Y(u2__abc_52155_new_n22143_));
OR2X2 OR2X2_5036 ( .A(u2__abc_52155_new_n22144_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22145_));
OR2X2 OR2X2_5037 ( .A(u2__abc_52155_new_n22149_), .B(u2__abc_52155_new_n22140_), .Y(u2__abc_52155_new_n22150_));
OR2X2 OR2X2_5038 ( .A(u2__abc_52155_new_n22141_), .B(u2_o_256_), .Y(u2__abc_52155_new_n22153_));
OR2X2 OR2X2_5039 ( .A(u2__abc_52155_new_n22156_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22157_));
OR2X2 OR2X2_504 ( .A(\a[113] ), .B(\a[114] ), .Y(u1__abc_51895_new_n144_));
OR2X2 OR2X2_5040 ( .A(u2__abc_52155_new_n22161_), .B(u2__abc_52155_new_n22152_), .Y(u2__abc_52155_new_n22162_));
OR2X2 OR2X2_5041 ( .A(u2__abc_52155_new_n22154_), .B(u2_o_257_), .Y(u2__abc_52155_new_n22165_));
OR2X2 OR2X2_5042 ( .A(u2__abc_52155_new_n22168_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22169_));
OR2X2 OR2X2_5043 ( .A(u2__abc_52155_new_n22173_), .B(u2__abc_52155_new_n22164_), .Y(u2__abc_52155_new_n22174_));
OR2X2 OR2X2_5044 ( .A(u2__abc_52155_new_n22166_), .B(u2_o_258_), .Y(u2__abc_52155_new_n22177_));
OR2X2 OR2X2_5045 ( .A(u2__abc_52155_new_n22180_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22181_));
OR2X2 OR2X2_5046 ( .A(u2__abc_52155_new_n22185_), .B(u2__abc_52155_new_n22176_), .Y(u2__abc_52155_new_n22186_));
OR2X2 OR2X2_5047 ( .A(u2__abc_52155_new_n22178_), .B(u2_o_259_), .Y(u2__abc_52155_new_n22191_));
OR2X2 OR2X2_5048 ( .A(u2__abc_52155_new_n22192_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22193_));
OR2X2 OR2X2_5049 ( .A(u2__abc_52155_new_n22197_), .B(u2__abc_52155_new_n22188_), .Y(u2__abc_52155_new_n22198_));
OR2X2 OR2X2_505 ( .A(u1__abc_51895_new_n144_), .B(\a[112] ), .Y(u1__abc_51895_new_n145_));
OR2X2 OR2X2_5050 ( .A(u2__abc_52155_new_n22189_), .B(u2_o_260_), .Y(u2__abc_52155_new_n22201_));
OR2X2 OR2X2_5051 ( .A(u2__abc_52155_new_n22204_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22205_));
OR2X2 OR2X2_5052 ( .A(u2__abc_52155_new_n22209_), .B(u2__abc_52155_new_n22200_), .Y(u2__abc_52155_new_n22210_));
OR2X2 OR2X2_5053 ( .A(u2__abc_52155_new_n22202_), .B(u2_o_261_), .Y(u2__abc_52155_new_n22215_));
OR2X2 OR2X2_5054 ( .A(u2__abc_52155_new_n22216_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22217_));
OR2X2 OR2X2_5055 ( .A(u2__abc_52155_new_n22221_), .B(u2__abc_52155_new_n22212_), .Y(u2__abc_52155_new_n22222_));
OR2X2 OR2X2_5056 ( .A(u2__abc_52155_new_n22213_), .B(u2_o_262_), .Y(u2__abc_52155_new_n22225_));
OR2X2 OR2X2_5057 ( .A(u2__abc_52155_new_n22228_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22229_));
OR2X2 OR2X2_5058 ( .A(u2__abc_52155_new_n22233_), .B(u2__abc_52155_new_n22224_), .Y(u2__abc_52155_new_n22234_));
OR2X2 OR2X2_5059 ( .A(u2__abc_52155_new_n22226_), .B(u2_o_263_), .Y(u2__abc_52155_new_n22237_));
OR2X2 OR2X2_506 ( .A(\a[117] ), .B(\a[118] ), .Y(u1__abc_51895_new_n146_));
OR2X2 OR2X2_5060 ( .A(u2__abc_52155_new_n22240_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22241_));
OR2X2 OR2X2_5061 ( .A(u2__abc_52155_new_n22245_), .B(u2__abc_52155_new_n22236_), .Y(u2__abc_52155_new_n22246_));
OR2X2 OR2X2_5062 ( .A(u2__abc_52155_new_n22238_), .B(u2_o_264_), .Y(u2__abc_52155_new_n22249_));
OR2X2 OR2X2_5063 ( .A(u2__abc_52155_new_n22252_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22253_));
OR2X2 OR2X2_5064 ( .A(u2__abc_52155_new_n22257_), .B(u2__abc_52155_new_n22248_), .Y(u2__abc_52155_new_n22258_));
OR2X2 OR2X2_5065 ( .A(u2__abc_52155_new_n22250_), .B(u2_o_265_), .Y(u2__abc_52155_new_n22263_));
OR2X2 OR2X2_5066 ( .A(u2__abc_52155_new_n22264_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22265_));
OR2X2 OR2X2_5067 ( .A(u2__abc_52155_new_n22269_), .B(u2__abc_52155_new_n22260_), .Y(u2__abc_52155_new_n22270_));
OR2X2 OR2X2_5068 ( .A(u2__abc_52155_new_n22261_), .B(u2_o_266_), .Y(u2__abc_52155_new_n22273_));
OR2X2 OR2X2_5069 ( .A(u2__abc_52155_new_n22276_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22277_));
OR2X2 OR2X2_507 ( .A(\a[115] ), .B(\a[116] ), .Y(u1__abc_51895_new_n147_));
OR2X2 OR2X2_5070 ( .A(u2__abc_52155_new_n22281_), .B(u2__abc_52155_new_n22272_), .Y(u2__abc_52155_new_n22282_));
OR2X2 OR2X2_5071 ( .A(u2__abc_52155_new_n22274_), .B(u2_o_267_), .Y(u2__abc_52155_new_n22285_));
OR2X2 OR2X2_5072 ( .A(u2__abc_52155_new_n22288_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22289_));
OR2X2 OR2X2_5073 ( .A(u2__abc_52155_new_n22293_), .B(u2__abc_52155_new_n22284_), .Y(u2__abc_52155_new_n22294_));
OR2X2 OR2X2_5074 ( .A(u2__abc_52155_new_n22286_), .B(u2_o_268_), .Y(u2__abc_52155_new_n22297_));
OR2X2 OR2X2_5075 ( .A(u2__abc_52155_new_n22300_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22301_));
OR2X2 OR2X2_5076 ( .A(u2__abc_52155_new_n22305_), .B(u2__abc_52155_new_n22296_), .Y(u2__abc_52155_new_n22306_));
OR2X2 OR2X2_5077 ( .A(u2__abc_52155_new_n22298_), .B(u2_o_269_), .Y(u2__abc_52155_new_n22311_));
OR2X2 OR2X2_5078 ( .A(u2__abc_52155_new_n22312_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22313_));
OR2X2 OR2X2_5079 ( .A(u2__abc_52155_new_n22317_), .B(u2__abc_52155_new_n22308_), .Y(u2__abc_52155_new_n22318_));
OR2X2 OR2X2_508 ( .A(u1__abc_51895_new_n146_), .B(u1__abc_51895_new_n147_), .Y(u1__abc_51895_new_n148_));
OR2X2 OR2X2_5080 ( .A(u2__abc_52155_new_n22309_), .B(u2_o_270_), .Y(u2__abc_52155_new_n22321_));
OR2X2 OR2X2_5081 ( .A(u2__abc_52155_new_n22324_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22325_));
OR2X2 OR2X2_5082 ( .A(u2__abc_52155_new_n22329_), .B(u2__abc_52155_new_n22320_), .Y(u2__abc_52155_new_n22330_));
OR2X2 OR2X2_5083 ( .A(u2__abc_52155_new_n22322_), .B(u2_o_271_), .Y(u2__abc_52155_new_n22333_));
OR2X2 OR2X2_5084 ( .A(u2__abc_52155_new_n22336_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22337_));
OR2X2 OR2X2_5085 ( .A(u2__abc_52155_new_n22341_), .B(u2__abc_52155_new_n22332_), .Y(u2__abc_52155_new_n22342_));
OR2X2 OR2X2_5086 ( .A(u2__abc_52155_new_n22334_), .B(u2_o_272_), .Y(u2__abc_52155_new_n22345_));
OR2X2 OR2X2_5087 ( .A(u2__abc_52155_new_n22348_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22349_));
OR2X2 OR2X2_5088 ( .A(u2__abc_52155_new_n22353_), .B(u2__abc_52155_new_n22344_), .Y(u2__abc_52155_new_n22354_));
OR2X2 OR2X2_5089 ( .A(u2__abc_52155_new_n22346_), .B(u2_o_273_), .Y(u2__abc_52155_new_n22359_));
OR2X2 OR2X2_509 ( .A(u1__abc_51895_new_n148_), .B(u1__abc_51895_new_n145_), .Y(u1__abc_51895_new_n149_));
OR2X2 OR2X2_5090 ( .A(u2__abc_52155_new_n22360_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22361_));
OR2X2 OR2X2_5091 ( .A(u2__abc_52155_new_n22365_), .B(u2__abc_52155_new_n22356_), .Y(u2__abc_52155_new_n22366_));
OR2X2 OR2X2_5092 ( .A(u2__abc_52155_new_n22357_), .B(u2_o_274_), .Y(u2__abc_52155_new_n22369_));
OR2X2 OR2X2_5093 ( .A(u2__abc_52155_new_n22372_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22373_));
OR2X2 OR2X2_5094 ( .A(u2__abc_52155_new_n22377_), .B(u2__abc_52155_new_n22368_), .Y(u2__abc_52155_new_n22378_));
OR2X2 OR2X2_5095 ( .A(u2__abc_52155_new_n22370_), .B(u2_o_275_), .Y(u2__abc_52155_new_n22381_));
OR2X2 OR2X2_5096 ( .A(u2__abc_52155_new_n22384_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22385_));
OR2X2 OR2X2_5097 ( .A(u2__abc_52155_new_n22389_), .B(u2__abc_52155_new_n22380_), .Y(u2__abc_52155_new_n22390_));
OR2X2 OR2X2_5098 ( .A(u2__abc_52155_new_n22382_), .B(u2_o_276_), .Y(u2__abc_52155_new_n22393_));
OR2X2 OR2X2_5099 ( .A(u2__abc_52155_new_n22396_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22397_));
OR2X2 OR2X2_51 ( .A(aNan), .B(sqrto_101_), .Y(_abc_73687_new_n905_));
OR2X2 OR2X2_510 ( .A(u1__abc_51895_new_n143_), .B(u1__abc_51895_new_n149_), .Y(fracta_112_));
OR2X2 OR2X2_5100 ( .A(u2__abc_52155_new_n22401_), .B(u2__abc_52155_new_n22392_), .Y(u2__abc_52155_new_n22402_));
OR2X2 OR2X2_5101 ( .A(u2__abc_52155_new_n22394_), .B(u2_o_277_), .Y(u2__abc_52155_new_n22407_));
OR2X2 OR2X2_5102 ( .A(u2__abc_52155_new_n22408_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22409_));
OR2X2 OR2X2_5103 ( .A(u2__abc_52155_new_n22413_), .B(u2__abc_52155_new_n22404_), .Y(u2__abc_52155_new_n22414_));
OR2X2 OR2X2_5104 ( .A(u2__abc_52155_new_n22405_), .B(u2_o_278_), .Y(u2__abc_52155_new_n22417_));
OR2X2 OR2X2_5105 ( .A(u2__abc_52155_new_n22420_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22421_));
OR2X2 OR2X2_5106 ( .A(u2__abc_52155_new_n22425_), .B(u2__abc_52155_new_n22416_), .Y(u2__abc_52155_new_n22426_));
OR2X2 OR2X2_5107 ( .A(u2__abc_52155_new_n22418_), .B(u2_o_279_), .Y(u2__abc_52155_new_n22429_));
OR2X2 OR2X2_5108 ( .A(u2__abc_52155_new_n22432_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22433_));
OR2X2 OR2X2_5109 ( .A(u2__abc_52155_new_n22437_), .B(u2__abc_52155_new_n22428_), .Y(u2__abc_52155_new_n22438_));
OR2X2 OR2X2_511 ( .A(u2_cnt_3_), .B(u2_cnt_2_), .Y(u2__abc_52155_new_n2969_));
OR2X2 OR2X2_5110 ( .A(u2__abc_52155_new_n22430_), .B(u2_o_280_), .Y(u2__abc_52155_new_n22441_));
OR2X2 OR2X2_5111 ( .A(u2__abc_52155_new_n22444_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22445_));
OR2X2 OR2X2_5112 ( .A(u2__abc_52155_new_n22449_), .B(u2__abc_52155_new_n22440_), .Y(u2__abc_52155_new_n22450_));
OR2X2 OR2X2_5113 ( .A(u2__abc_52155_new_n22442_), .B(u2_o_281_), .Y(u2__abc_52155_new_n22455_));
OR2X2 OR2X2_5114 ( .A(u2__abc_52155_new_n22456_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22457_));
OR2X2 OR2X2_5115 ( .A(u2__abc_52155_new_n22461_), .B(u2__abc_52155_new_n22452_), .Y(u2__abc_52155_new_n22462_));
OR2X2 OR2X2_5116 ( .A(u2__abc_52155_new_n22453_), .B(u2_o_282_), .Y(u2__abc_52155_new_n22465_));
OR2X2 OR2X2_5117 ( .A(u2__abc_52155_new_n22468_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22469_));
OR2X2 OR2X2_5118 ( .A(u2__abc_52155_new_n22473_), .B(u2__abc_52155_new_n22464_), .Y(u2__abc_52155_new_n22474_));
OR2X2 OR2X2_5119 ( .A(u2__abc_52155_new_n22466_), .B(u2_o_283_), .Y(u2__abc_52155_new_n22477_));
OR2X2 OR2X2_512 ( .A(u2__abc_52155_new_n2977_), .B(u2__abc_52155_new_n2964_), .Y(u2__abc_52155_new_n2978_));
OR2X2 OR2X2_5120 ( .A(u2__abc_52155_new_n22480_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22481_));
OR2X2 OR2X2_5121 ( .A(u2__abc_52155_new_n22485_), .B(u2__abc_52155_new_n22476_), .Y(u2__abc_52155_new_n22486_));
OR2X2 OR2X2_5122 ( .A(u2__abc_52155_new_n22478_), .B(u2_o_284_), .Y(u2__abc_52155_new_n22489_));
OR2X2 OR2X2_5123 ( .A(u2__abc_52155_new_n22492_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22493_));
OR2X2 OR2X2_5124 ( .A(u2__abc_52155_new_n22497_), .B(u2__abc_52155_new_n22488_), .Y(u2__abc_52155_new_n22498_));
OR2X2 OR2X2_5125 ( .A(u2__abc_52155_new_n22490_), .B(u2_o_285_), .Y(u2__abc_52155_new_n22503_));
OR2X2 OR2X2_5126 ( .A(u2__abc_52155_new_n22504_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22505_));
OR2X2 OR2X2_5127 ( .A(u2__abc_52155_new_n22509_), .B(u2__abc_52155_new_n22500_), .Y(u2__abc_52155_new_n22510_));
OR2X2 OR2X2_5128 ( .A(u2__abc_52155_new_n22501_), .B(u2_o_286_), .Y(u2__abc_52155_new_n22513_));
OR2X2 OR2X2_5129 ( .A(u2__abc_52155_new_n22516_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22517_));
OR2X2 OR2X2_513 ( .A(rst), .B(ce), .Y(u2__abc_52155_new_n2980_));
OR2X2 OR2X2_5130 ( .A(u2__abc_52155_new_n22521_), .B(u2__abc_52155_new_n22512_), .Y(u2__abc_52155_new_n22522_));
OR2X2 OR2X2_5131 ( .A(u2__abc_52155_new_n22514_), .B(u2_o_287_), .Y(u2__abc_52155_new_n22527_));
OR2X2 OR2X2_5132 ( .A(u2__abc_52155_new_n22528_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22529_));
OR2X2 OR2X2_5133 ( .A(u2__abc_52155_new_n22533_), .B(u2__abc_52155_new_n22524_), .Y(u2__abc_52155_new_n22534_));
OR2X2 OR2X2_5134 ( .A(u2__abc_52155_new_n22525_), .B(u2_o_288_), .Y(u2__abc_52155_new_n22537_));
OR2X2 OR2X2_5135 ( .A(u2__abc_52155_new_n22540_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22541_));
OR2X2 OR2X2_5136 ( .A(u2__abc_52155_new_n22545_), .B(u2__abc_52155_new_n22536_), .Y(u2__abc_52155_new_n22546_));
OR2X2 OR2X2_5137 ( .A(u2__abc_52155_new_n22538_), .B(u2_o_289_), .Y(u2__abc_52155_new_n22551_));
OR2X2 OR2X2_5138 ( .A(u2__abc_52155_new_n22552_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22553_));
OR2X2 OR2X2_5139 ( .A(u2__abc_52155_new_n22557_), .B(u2__abc_52155_new_n22548_), .Y(u2__abc_52155_new_n22558_));
OR2X2 OR2X2_514 ( .A(u2__abc_52155_new_n2980_), .B(u2_state_0_), .Y(u2__abc_52155_new_n2981_));
OR2X2 OR2X2_5140 ( .A(u2__abc_52155_new_n22549_), .B(u2_o_290_), .Y(u2__abc_52155_new_n22561_));
OR2X2 OR2X2_5141 ( .A(u2__abc_52155_new_n22564_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22565_));
OR2X2 OR2X2_5142 ( .A(u2__abc_52155_new_n22569_), .B(u2__abc_52155_new_n22560_), .Y(u2__abc_52155_new_n22570_));
OR2X2 OR2X2_5143 ( .A(u2__abc_52155_new_n22562_), .B(u2_o_291_), .Y(u2__abc_52155_new_n22573_));
OR2X2 OR2X2_5144 ( .A(u2__abc_52155_new_n22576_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22577_));
OR2X2 OR2X2_5145 ( .A(u2__abc_52155_new_n22581_), .B(u2__abc_52155_new_n22572_), .Y(u2__abc_52155_new_n22582_));
OR2X2 OR2X2_5146 ( .A(u2__abc_52155_new_n22574_), .B(u2_o_292_), .Y(u2__abc_52155_new_n22585_));
OR2X2 OR2X2_5147 ( .A(u2__abc_52155_new_n22588_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22589_));
OR2X2 OR2X2_5148 ( .A(u2__abc_52155_new_n22593_), .B(u2__abc_52155_new_n22584_), .Y(u2__abc_52155_new_n22594_));
OR2X2 OR2X2_5149 ( .A(u2__abc_52155_new_n22586_), .B(u2_o_293_), .Y(u2__abc_52155_new_n22599_));
OR2X2 OR2X2_515 ( .A(u2__abc_52155_new_n2985_), .B(done), .Y(u2__abc_52155_new_n2986_));
OR2X2 OR2X2_5150 ( .A(u2__abc_52155_new_n22600_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22601_));
OR2X2 OR2X2_5151 ( .A(u2__abc_52155_new_n22605_), .B(u2__abc_52155_new_n22596_), .Y(u2__abc_52155_new_n22606_));
OR2X2 OR2X2_5152 ( .A(u2__abc_52155_new_n22597_), .B(u2_o_294_), .Y(u2__abc_52155_new_n22609_));
OR2X2 OR2X2_5153 ( .A(u2__abc_52155_new_n22612_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22613_));
OR2X2 OR2X2_5154 ( .A(u2__abc_52155_new_n22617_), .B(u2__abc_52155_new_n22608_), .Y(u2__abc_52155_new_n22618_));
OR2X2 OR2X2_5155 ( .A(u2__abc_52155_new_n22610_), .B(u2_o_295_), .Y(u2__abc_52155_new_n22621_));
OR2X2 OR2X2_5156 ( .A(u2__abc_52155_new_n22624_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22625_));
OR2X2 OR2X2_5157 ( .A(u2__abc_52155_new_n22629_), .B(u2__abc_52155_new_n22620_), .Y(u2__abc_52155_new_n22630_));
OR2X2 OR2X2_5158 ( .A(u2__abc_52155_new_n22622_), .B(u2_o_296_), .Y(u2__abc_52155_new_n22633_));
OR2X2 OR2X2_5159 ( .A(u2__abc_52155_new_n22636_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22637_));
OR2X2 OR2X2_516 ( .A(u2__abc_52155_new_n2986_), .B(u2__abc_52155_new_n2983_), .Y(u2__abc_52155_new_n2987_));
OR2X2 OR2X2_5160 ( .A(u2__abc_52155_new_n22641_), .B(u2__abc_52155_new_n22632_), .Y(u2__abc_52155_new_n22642_));
OR2X2 OR2X2_5161 ( .A(u2__abc_52155_new_n22634_), .B(u2_o_297_), .Y(u2__abc_52155_new_n22647_));
OR2X2 OR2X2_5162 ( .A(u2__abc_52155_new_n22648_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22649_));
OR2X2 OR2X2_5163 ( .A(u2__abc_52155_new_n22653_), .B(u2__abc_52155_new_n22644_), .Y(u2__abc_52155_new_n22654_));
OR2X2 OR2X2_5164 ( .A(u2__abc_52155_new_n22645_), .B(u2_o_298_), .Y(u2__abc_52155_new_n22657_));
OR2X2 OR2X2_5165 ( .A(u2__abc_52155_new_n22660_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22661_));
OR2X2 OR2X2_5166 ( .A(u2__abc_52155_new_n22665_), .B(u2__abc_52155_new_n22656_), .Y(u2__abc_52155_new_n22666_));
OR2X2 OR2X2_5167 ( .A(u2__abc_52155_new_n22658_), .B(u2_o_299_), .Y(u2__abc_52155_new_n22669_));
OR2X2 OR2X2_5168 ( .A(u2__abc_52155_new_n22672_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22673_));
OR2X2 OR2X2_5169 ( .A(u2__abc_52155_new_n22677_), .B(u2__abc_52155_new_n22668_), .Y(u2__abc_52155_new_n22678_));
OR2X2 OR2X2_517 ( .A(u2__abc_52155_new_n2995_), .B(u2__abc_52155_new_n2990_), .Y(u2__abc_34132_auto_fsm_map_cc_170_map_fsm_175_1_));
OR2X2 OR2X2_5170 ( .A(u2__abc_52155_new_n22670_), .B(u2_o_300_), .Y(u2__abc_52155_new_n22681_));
OR2X2 OR2X2_5171 ( .A(u2__abc_52155_new_n22684_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22685_));
OR2X2 OR2X2_5172 ( .A(u2__abc_52155_new_n22689_), .B(u2__abc_52155_new_n22680_), .Y(u2__abc_52155_new_n22690_));
OR2X2 OR2X2_5173 ( .A(u2__abc_52155_new_n22682_), .B(u2_o_301_), .Y(u2__abc_52155_new_n22695_));
OR2X2 OR2X2_5174 ( .A(u2__abc_52155_new_n22696_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22697_));
OR2X2 OR2X2_5175 ( .A(u2__abc_52155_new_n22701_), .B(u2__abc_52155_new_n22692_), .Y(u2__abc_52155_new_n22702_));
OR2X2 OR2X2_5176 ( .A(u2__abc_52155_new_n22693_), .B(u2_o_302_), .Y(u2__abc_52155_new_n22705_));
OR2X2 OR2X2_5177 ( .A(u2__abc_52155_new_n22708_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22709_));
OR2X2 OR2X2_5178 ( .A(u2__abc_52155_new_n22713_), .B(u2__abc_52155_new_n22704_), .Y(u2__abc_52155_new_n22714_));
OR2X2 OR2X2_5179 ( .A(u2__abc_52155_new_n22706_), .B(u2_o_303_), .Y(u2__abc_52155_new_n22719_));
OR2X2 OR2X2_518 ( .A(u2__abc_52155_new_n3001_), .B(u2__abc_52155_new_n2985_), .Y(u2__abc_52155_new_n3002_));
OR2X2 OR2X2_5180 ( .A(u2__abc_52155_new_n22720_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22721_));
OR2X2 OR2X2_5181 ( .A(u2__abc_52155_new_n22725_), .B(u2__abc_52155_new_n22716_), .Y(u2__abc_52155_new_n22726_));
OR2X2 OR2X2_5182 ( .A(u2__abc_52155_new_n22717_), .B(u2_o_304_), .Y(u2__abc_52155_new_n22729_));
OR2X2 OR2X2_5183 ( .A(u2__abc_52155_new_n22732_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22733_));
OR2X2 OR2X2_5184 ( .A(u2__abc_52155_new_n22737_), .B(u2__abc_52155_new_n22728_), .Y(u2__abc_52155_new_n22738_));
OR2X2 OR2X2_5185 ( .A(u2__abc_52155_new_n22730_), .B(u2_o_305_), .Y(u2__abc_52155_new_n22743_));
OR2X2 OR2X2_5186 ( .A(u2__abc_52155_new_n22744_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22745_));
OR2X2 OR2X2_5187 ( .A(u2__abc_52155_new_n22749_), .B(u2__abc_52155_new_n22740_), .Y(u2__abc_52155_new_n22750_));
OR2X2 OR2X2_5188 ( .A(u2__abc_52155_new_n22741_), .B(u2_o_306_), .Y(u2__abc_52155_new_n22753_));
OR2X2 OR2X2_5189 ( .A(u2__abc_52155_new_n22756_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22757_));
OR2X2 OR2X2_519 ( .A(u2__abc_52155_new_n3012_), .B(u2__abc_52155_new_n3014_), .Y(u2__abc_52155_new_n3015_));
OR2X2 OR2X2_5190 ( .A(u2__abc_52155_new_n22761_), .B(u2__abc_52155_new_n22752_), .Y(u2__abc_52155_new_n22762_));
OR2X2 OR2X2_5191 ( .A(u2__abc_52155_new_n22754_), .B(u2_o_307_), .Y(u2__abc_52155_new_n22765_));
OR2X2 OR2X2_5192 ( .A(u2__abc_52155_new_n22768_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22769_));
OR2X2 OR2X2_5193 ( .A(u2__abc_52155_new_n22773_), .B(u2__abc_52155_new_n22764_), .Y(u2__abc_52155_new_n22774_));
OR2X2 OR2X2_5194 ( .A(u2__abc_52155_new_n22766_), .B(u2_o_308_), .Y(u2__abc_52155_new_n22777_));
OR2X2 OR2X2_5195 ( .A(u2__abc_52155_new_n22780_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22781_));
OR2X2 OR2X2_5196 ( .A(u2__abc_52155_new_n22785_), .B(u2__abc_52155_new_n22776_), .Y(u2__abc_52155_new_n22786_));
OR2X2 OR2X2_5197 ( .A(u2__abc_52155_new_n22778_), .B(u2_o_309_), .Y(u2__abc_52155_new_n22791_));
OR2X2 OR2X2_5198 ( .A(u2__abc_52155_new_n22792_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22793_));
OR2X2 OR2X2_5199 ( .A(u2__abc_52155_new_n22797_), .B(u2__abc_52155_new_n22788_), .Y(u2__abc_52155_new_n22798_));
OR2X2 OR2X2_52 ( .A(_abc_73687_new_n753_), .B(\a[25] ), .Y(_abc_73687_new_n906_));
OR2X2 OR2X2_520 ( .A(u2__abc_52155_new_n3036_), .B(u2__abc_52155_new_n3038_), .Y(u2__abc_52155_new_n3039_));
OR2X2 OR2X2_5200 ( .A(u2__abc_52155_new_n22789_), .B(u2_o_310_), .Y(u2__abc_52155_new_n22801_));
OR2X2 OR2X2_5201 ( .A(u2__abc_52155_new_n22804_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22805_));
OR2X2 OR2X2_5202 ( .A(u2__abc_52155_new_n22809_), .B(u2__abc_52155_new_n22800_), .Y(u2__abc_52155_new_n22810_));
OR2X2 OR2X2_5203 ( .A(u2__abc_52155_new_n22802_), .B(u2_o_311_), .Y(u2__abc_52155_new_n22815_));
OR2X2 OR2X2_5204 ( .A(u2__abc_52155_new_n22816_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22817_));
OR2X2 OR2X2_5205 ( .A(u2__abc_52155_new_n22821_), .B(u2__abc_52155_new_n22812_), .Y(u2__abc_52155_new_n22822_));
OR2X2 OR2X2_5206 ( .A(u2__abc_52155_new_n22813_), .B(u2_o_312_), .Y(u2__abc_52155_new_n22825_));
OR2X2 OR2X2_5207 ( .A(u2__abc_52155_new_n22828_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22829_));
OR2X2 OR2X2_5208 ( .A(u2__abc_52155_new_n22833_), .B(u2__abc_52155_new_n22824_), .Y(u2__abc_52155_new_n22834_));
OR2X2 OR2X2_5209 ( .A(u2__abc_52155_new_n22826_), .B(u2_o_313_), .Y(u2__abc_52155_new_n22839_));
OR2X2 OR2X2_521 ( .A(u2__abc_52155_new_n3042_), .B(u2__abc_52155_new_n3044_), .Y(u2__abc_52155_new_n3045_));
OR2X2 OR2X2_5210 ( .A(u2__abc_52155_new_n22840_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22841_));
OR2X2 OR2X2_5211 ( .A(u2__abc_52155_new_n22845_), .B(u2__abc_52155_new_n22836_), .Y(u2__abc_52155_new_n22846_));
OR2X2 OR2X2_5212 ( .A(u2__abc_52155_new_n22837_), .B(u2_o_314_), .Y(u2__abc_52155_new_n22849_));
OR2X2 OR2X2_5213 ( .A(u2__abc_52155_new_n22852_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22853_));
OR2X2 OR2X2_5214 ( .A(u2__abc_52155_new_n22857_), .B(u2__abc_52155_new_n22848_), .Y(u2__abc_52155_new_n22858_));
OR2X2 OR2X2_5215 ( .A(u2__abc_52155_new_n22850_), .B(u2_o_315_), .Y(u2__abc_52155_new_n22863_));
OR2X2 OR2X2_5216 ( .A(u2__abc_52155_new_n22864_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22865_));
OR2X2 OR2X2_5217 ( .A(u2__abc_52155_new_n22869_), .B(u2__abc_52155_new_n22860_), .Y(u2__abc_52155_new_n22870_));
OR2X2 OR2X2_5218 ( .A(u2__abc_52155_new_n22861_), .B(u2_o_316_), .Y(u2__abc_52155_new_n22873_));
OR2X2 OR2X2_5219 ( .A(u2__abc_52155_new_n22876_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22877_));
OR2X2 OR2X2_522 ( .A(u2__abc_52155_new_n3056_), .B(u2__abc_52155_new_n3058_), .Y(u2__abc_52155_new_n3059_));
OR2X2 OR2X2_5220 ( .A(u2__abc_52155_new_n22881_), .B(u2__abc_52155_new_n22872_), .Y(u2__abc_52155_new_n22882_));
OR2X2 OR2X2_5221 ( .A(u2__abc_52155_new_n22874_), .B(u2_o_317_), .Y(u2__abc_52155_new_n22887_));
OR2X2 OR2X2_5222 ( .A(u2__abc_52155_new_n22888_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22889_));
OR2X2 OR2X2_5223 ( .A(u2__abc_52155_new_n22893_), .B(u2__abc_52155_new_n22884_), .Y(u2__abc_52155_new_n22894_));
OR2X2 OR2X2_5224 ( .A(u2__abc_52155_new_n22885_), .B(u2_o_318_), .Y(u2__abc_52155_new_n22897_));
OR2X2 OR2X2_5225 ( .A(u2__abc_52155_new_n22900_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22901_));
OR2X2 OR2X2_5226 ( .A(u2__abc_52155_new_n22905_), .B(u2__abc_52155_new_n22896_), .Y(u2__abc_52155_new_n22906_));
OR2X2 OR2X2_5227 ( .A(u2__abc_52155_new_n22898_), .B(u2_o_319_), .Y(u2__abc_52155_new_n22911_));
OR2X2 OR2X2_5228 ( .A(u2__abc_52155_new_n22912_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22913_));
OR2X2 OR2X2_5229 ( .A(u2__abc_52155_new_n22917_), .B(u2__abc_52155_new_n22908_), .Y(u2__abc_52155_new_n22918_));
OR2X2 OR2X2_523 ( .A(u2__abc_52155_new_n3064_), .B(u2__abc_52155_new_n3066_), .Y(u2__abc_52155_new_n3067_));
OR2X2 OR2X2_5230 ( .A(u2__abc_52155_new_n22909_), .B(u2_o_320_), .Y(u2__abc_52155_new_n22921_));
OR2X2 OR2X2_5231 ( .A(u2__abc_52155_new_n22924_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22925_));
OR2X2 OR2X2_5232 ( .A(u2__abc_52155_new_n22929_), .B(u2__abc_52155_new_n22920_), .Y(u2__abc_52155_new_n22930_));
OR2X2 OR2X2_5233 ( .A(u2__abc_52155_new_n22922_), .B(u2_o_321_), .Y(u2__abc_52155_new_n22935_));
OR2X2 OR2X2_5234 ( .A(u2__abc_52155_new_n22936_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22937_));
OR2X2 OR2X2_5235 ( .A(u2__abc_52155_new_n22941_), .B(u2__abc_52155_new_n22932_), .Y(u2__abc_52155_new_n22942_));
OR2X2 OR2X2_5236 ( .A(u2__abc_52155_new_n22933_), .B(u2_o_322_), .Y(u2__abc_52155_new_n22945_));
OR2X2 OR2X2_5237 ( .A(u2__abc_52155_new_n22948_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22949_));
OR2X2 OR2X2_5238 ( .A(u2__abc_52155_new_n22953_), .B(u2__abc_52155_new_n22944_), .Y(u2__abc_52155_new_n22954_));
OR2X2 OR2X2_5239 ( .A(u2__abc_52155_new_n22946_), .B(u2_o_323_), .Y(u2__abc_52155_new_n22957_));
OR2X2 OR2X2_524 ( .A(u2__abc_52155_new_n3077_), .B(u2_remHi_7_), .Y(u2__abc_52155_new_n3080_));
OR2X2 OR2X2_5240 ( .A(u2__abc_52155_new_n22960_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22961_));
OR2X2 OR2X2_5241 ( .A(u2__abc_52155_new_n22965_), .B(u2__abc_52155_new_n22956_), .Y(u2__abc_52155_new_n22966_));
OR2X2 OR2X2_5242 ( .A(u2__abc_52155_new_n22958_), .B(u2_o_324_), .Y(u2__abc_52155_new_n22969_));
OR2X2 OR2X2_5243 ( .A(u2__abc_52155_new_n22972_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22973_));
OR2X2 OR2X2_5244 ( .A(u2__abc_52155_new_n22977_), .B(u2__abc_52155_new_n22968_), .Y(u2__abc_52155_new_n22978_));
OR2X2 OR2X2_5245 ( .A(u2__abc_52155_new_n22970_), .B(u2_o_325_), .Y(u2__abc_52155_new_n22983_));
OR2X2 OR2X2_5246 ( .A(u2__abc_52155_new_n22984_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22985_));
OR2X2 OR2X2_5247 ( .A(u2__abc_52155_new_n22989_), .B(u2__abc_52155_new_n22980_), .Y(u2__abc_52155_new_n22990_));
OR2X2 OR2X2_5248 ( .A(u2__abc_52155_new_n22981_), .B(u2_o_326_), .Y(u2__abc_52155_new_n22993_));
OR2X2 OR2X2_5249 ( .A(u2__abc_52155_new_n22996_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n22997_));
OR2X2 OR2X2_525 ( .A(u2__abc_52155_new_n3082_), .B(sqrto_6_), .Y(u2__abc_52155_new_n3083_));
OR2X2 OR2X2_5250 ( .A(u2__abc_52155_new_n23001_), .B(u2__abc_52155_new_n22992_), .Y(u2__abc_52155_new_n23002_));
OR2X2 OR2X2_5251 ( .A(u2__abc_52155_new_n22994_), .B(u2_o_327_), .Y(u2__abc_52155_new_n23005_));
OR2X2 OR2X2_5252 ( .A(u2__abc_52155_new_n23008_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23009_));
OR2X2 OR2X2_5253 ( .A(u2__abc_52155_new_n23013_), .B(u2__abc_52155_new_n23004_), .Y(u2__abc_52155_new_n23014_));
OR2X2 OR2X2_5254 ( .A(u2__abc_52155_new_n23006_), .B(u2_o_328_), .Y(u2__abc_52155_new_n23017_));
OR2X2 OR2X2_5255 ( .A(u2__abc_52155_new_n23020_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23021_));
OR2X2 OR2X2_5256 ( .A(u2__abc_52155_new_n23025_), .B(u2__abc_52155_new_n23016_), .Y(u2__abc_52155_new_n23026_));
OR2X2 OR2X2_5257 ( .A(u2__abc_52155_new_n23018_), .B(u2_o_329_), .Y(u2__abc_52155_new_n23031_));
OR2X2 OR2X2_5258 ( .A(u2__abc_52155_new_n23032_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23033_));
OR2X2 OR2X2_5259 ( .A(u2__abc_52155_new_n23037_), .B(u2__abc_52155_new_n23028_), .Y(u2__abc_52155_new_n23038_));
OR2X2 OR2X2_526 ( .A(u2__abc_52155_new_n3084_), .B(u2_remHi_6_), .Y(u2__abc_52155_new_n3085_));
OR2X2 OR2X2_5260 ( .A(u2__abc_52155_new_n23029_), .B(u2_o_330_), .Y(u2__abc_52155_new_n23041_));
OR2X2 OR2X2_5261 ( .A(u2__abc_52155_new_n23044_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23045_));
OR2X2 OR2X2_5262 ( .A(u2__abc_52155_new_n23049_), .B(u2__abc_52155_new_n23040_), .Y(u2__abc_52155_new_n23050_));
OR2X2 OR2X2_5263 ( .A(u2__abc_52155_new_n23042_), .B(u2_o_331_), .Y(u2__abc_52155_new_n23053_));
OR2X2 OR2X2_5264 ( .A(u2__abc_52155_new_n23056_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23057_));
OR2X2 OR2X2_5265 ( .A(u2__abc_52155_new_n23061_), .B(u2__abc_52155_new_n23052_), .Y(u2__abc_52155_new_n23062_));
OR2X2 OR2X2_5266 ( .A(u2__abc_52155_new_n23054_), .B(u2_o_332_), .Y(u2__abc_52155_new_n23065_));
OR2X2 OR2X2_5267 ( .A(u2__abc_52155_new_n23068_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23069_));
OR2X2 OR2X2_5268 ( .A(u2__abc_52155_new_n23073_), .B(u2__abc_52155_new_n23064_), .Y(u2__abc_52155_new_n23074_));
OR2X2 OR2X2_5269 ( .A(u2__abc_52155_new_n23066_), .B(u2_o_333_), .Y(u2__abc_52155_new_n23079_));
OR2X2 OR2X2_527 ( .A(u2__abc_52155_new_n3092_), .B(u2__abc_52155_new_n3094_), .Y(u2__abc_52155_new_n3095_));
OR2X2 OR2X2_5270 ( .A(u2__abc_52155_new_n23080_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23081_));
OR2X2 OR2X2_5271 ( .A(u2__abc_52155_new_n23085_), .B(u2__abc_52155_new_n23076_), .Y(u2__abc_52155_new_n23086_));
OR2X2 OR2X2_5272 ( .A(u2__abc_52155_new_n23077_), .B(u2_o_334_), .Y(u2__abc_52155_new_n23089_));
OR2X2 OR2X2_5273 ( .A(u2__abc_52155_new_n23092_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23093_));
OR2X2 OR2X2_5274 ( .A(u2__abc_52155_new_n23097_), .B(u2__abc_52155_new_n23088_), .Y(u2__abc_52155_new_n23098_));
OR2X2 OR2X2_5275 ( .A(u2__abc_52155_new_n23090_), .B(u2_o_335_), .Y(u2__abc_52155_new_n23103_));
OR2X2 OR2X2_5276 ( .A(u2__abc_52155_new_n23104_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23105_));
OR2X2 OR2X2_5277 ( .A(u2__abc_52155_new_n23109_), .B(u2__abc_52155_new_n23100_), .Y(u2__abc_52155_new_n23110_));
OR2X2 OR2X2_5278 ( .A(u2__abc_52155_new_n23101_), .B(u2_o_336_), .Y(u2__abc_52155_new_n23113_));
OR2X2 OR2X2_5279 ( .A(u2__abc_52155_new_n23116_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23117_));
OR2X2 OR2X2_528 ( .A(u2__abc_52155_new_n3097_), .B(u2__abc_52155_new_n3099_), .Y(u2__abc_52155_new_n3100_));
OR2X2 OR2X2_5280 ( .A(u2__abc_52155_new_n23121_), .B(u2__abc_52155_new_n23112_), .Y(u2__abc_52155_new_n23122_));
OR2X2 OR2X2_5281 ( .A(u2__abc_52155_new_n23114_), .B(u2_o_337_), .Y(u2__abc_52155_new_n23127_));
OR2X2 OR2X2_5282 ( .A(u2__abc_52155_new_n23128_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23129_));
OR2X2 OR2X2_5283 ( .A(u2__abc_52155_new_n23133_), .B(u2__abc_52155_new_n23124_), .Y(u2__abc_52155_new_n23134_));
OR2X2 OR2X2_5284 ( .A(u2__abc_52155_new_n23125_), .B(u2_o_338_), .Y(u2__abc_52155_new_n23137_));
OR2X2 OR2X2_5285 ( .A(u2__abc_52155_new_n23140_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23141_));
OR2X2 OR2X2_5286 ( .A(u2__abc_52155_new_n23145_), .B(u2__abc_52155_new_n23136_), .Y(u2__abc_52155_new_n23146_));
OR2X2 OR2X2_5287 ( .A(u2__abc_52155_new_n23138_), .B(u2_o_339_), .Y(u2__abc_52155_new_n23149_));
OR2X2 OR2X2_5288 ( .A(u2__abc_52155_new_n23152_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23153_));
OR2X2 OR2X2_5289 ( .A(u2__abc_52155_new_n23157_), .B(u2__abc_52155_new_n23148_), .Y(u2__abc_52155_new_n23158_));
OR2X2 OR2X2_529 ( .A(u2__abc_52155_new_n3095_), .B(u2__abc_52155_new_n3100_), .Y(u2__abc_52155_new_n3101_));
OR2X2 OR2X2_5290 ( .A(u2__abc_52155_new_n23150_), .B(u2_o_340_), .Y(u2__abc_52155_new_n23161_));
OR2X2 OR2X2_5291 ( .A(u2__abc_52155_new_n23164_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23165_));
OR2X2 OR2X2_5292 ( .A(u2__abc_52155_new_n23169_), .B(u2__abc_52155_new_n23160_), .Y(u2__abc_52155_new_n23170_));
OR2X2 OR2X2_5293 ( .A(u2__abc_52155_new_n23162_), .B(u2_o_341_), .Y(u2__abc_52155_new_n23175_));
OR2X2 OR2X2_5294 ( .A(u2__abc_52155_new_n23176_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23177_));
OR2X2 OR2X2_5295 ( .A(u2__abc_52155_new_n23181_), .B(u2__abc_52155_new_n23172_), .Y(u2__abc_52155_new_n23182_));
OR2X2 OR2X2_5296 ( .A(u2__abc_52155_new_n23173_), .B(u2_o_342_), .Y(u2__abc_52155_new_n23185_));
OR2X2 OR2X2_5297 ( .A(u2__abc_52155_new_n23188_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23189_));
OR2X2 OR2X2_5298 ( .A(u2__abc_52155_new_n23193_), .B(u2__abc_52155_new_n23184_), .Y(u2__abc_52155_new_n23194_));
OR2X2 OR2X2_5299 ( .A(u2__abc_52155_new_n23186_), .B(u2_o_343_), .Y(u2__abc_52155_new_n23199_));
OR2X2 OR2X2_53 ( .A(aNan), .B(sqrto_102_), .Y(_abc_73687_new_n908_));
OR2X2 OR2X2_530 ( .A(u2__abc_52155_new_n3103_), .B(u2__abc_52155_new_n3105_), .Y(u2__abc_52155_new_n3106_));
OR2X2 OR2X2_5300 ( .A(u2__abc_52155_new_n23200_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23201_));
OR2X2 OR2X2_5301 ( .A(u2__abc_52155_new_n23205_), .B(u2__abc_52155_new_n23196_), .Y(u2__abc_52155_new_n23206_));
OR2X2 OR2X2_5302 ( .A(u2__abc_52155_new_n23197_), .B(u2_o_344_), .Y(u2__abc_52155_new_n23209_));
OR2X2 OR2X2_5303 ( .A(u2__abc_52155_new_n23212_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23213_));
OR2X2 OR2X2_5304 ( .A(u2__abc_52155_new_n23217_), .B(u2__abc_52155_new_n23208_), .Y(u2__abc_52155_new_n23218_));
OR2X2 OR2X2_5305 ( .A(u2__abc_52155_new_n23210_), .B(u2_o_345_), .Y(u2__abc_52155_new_n23223_));
OR2X2 OR2X2_5306 ( .A(u2__abc_52155_new_n23224_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23225_));
OR2X2 OR2X2_5307 ( .A(u2__abc_52155_new_n23229_), .B(u2__abc_52155_new_n23220_), .Y(u2__abc_52155_new_n23230_));
OR2X2 OR2X2_5308 ( .A(u2__abc_52155_new_n23221_), .B(u2_o_346_), .Y(u2__abc_52155_new_n23233_));
OR2X2 OR2X2_5309 ( .A(u2__abc_52155_new_n23236_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23237_));
OR2X2 OR2X2_531 ( .A(u2__abc_52155_new_n3108_), .B(u2__abc_52155_new_n3110_), .Y(u2__abc_52155_new_n3111_));
OR2X2 OR2X2_5310 ( .A(u2__abc_52155_new_n23241_), .B(u2__abc_52155_new_n23232_), .Y(u2__abc_52155_new_n23242_));
OR2X2 OR2X2_5311 ( .A(u2__abc_52155_new_n23234_), .B(u2_o_347_), .Y(u2__abc_52155_new_n23247_));
OR2X2 OR2X2_5312 ( .A(u2__abc_52155_new_n23248_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23249_));
OR2X2 OR2X2_5313 ( .A(u2__abc_52155_new_n23253_), .B(u2__abc_52155_new_n23244_), .Y(u2__abc_52155_new_n23254_));
OR2X2 OR2X2_5314 ( .A(u2__abc_52155_new_n23245_), .B(u2_o_348_), .Y(u2__abc_52155_new_n23257_));
OR2X2 OR2X2_5315 ( .A(u2__abc_52155_new_n23260_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23261_));
OR2X2 OR2X2_5316 ( .A(u2__abc_52155_new_n23265_), .B(u2__abc_52155_new_n23256_), .Y(u2__abc_52155_new_n23266_));
OR2X2 OR2X2_5317 ( .A(u2__abc_52155_new_n23258_), .B(u2_o_349_), .Y(u2__abc_52155_new_n23271_));
OR2X2 OR2X2_5318 ( .A(u2__abc_52155_new_n23272_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23273_));
OR2X2 OR2X2_5319 ( .A(u2__abc_52155_new_n23277_), .B(u2__abc_52155_new_n23268_), .Y(u2__abc_52155_new_n23278_));
OR2X2 OR2X2_532 ( .A(u2__abc_52155_new_n3106_), .B(u2__abc_52155_new_n3111_), .Y(u2__abc_52155_new_n3112_));
OR2X2 OR2X2_5320 ( .A(u2__abc_52155_new_n23269_), .B(u2_o_350_), .Y(u2__abc_52155_new_n23281_));
OR2X2 OR2X2_5321 ( .A(u2__abc_52155_new_n23284_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23285_));
OR2X2 OR2X2_5322 ( .A(u2__abc_52155_new_n23289_), .B(u2__abc_52155_new_n23280_), .Y(u2__abc_52155_new_n23290_));
OR2X2 OR2X2_5323 ( .A(u2__abc_52155_new_n23282_), .B(u2_o_351_), .Y(u2__abc_52155_new_n23295_));
OR2X2 OR2X2_5324 ( .A(u2__abc_52155_new_n23296_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23297_));
OR2X2 OR2X2_5325 ( .A(u2__abc_52155_new_n23301_), .B(u2__abc_52155_new_n23292_), .Y(u2__abc_52155_new_n23302_));
OR2X2 OR2X2_5326 ( .A(u2__abc_52155_new_n23293_), .B(u2_o_352_), .Y(u2__abc_52155_new_n23305_));
OR2X2 OR2X2_5327 ( .A(u2__abc_52155_new_n23308_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23309_));
OR2X2 OR2X2_5328 ( .A(u2__abc_52155_new_n23313_), .B(u2__abc_52155_new_n23304_), .Y(u2__abc_52155_new_n23314_));
OR2X2 OR2X2_5329 ( .A(u2__abc_52155_new_n23306_), .B(u2_o_353_), .Y(u2__abc_52155_new_n23319_));
OR2X2 OR2X2_533 ( .A(u2__abc_52155_new_n3101_), .B(u2__abc_52155_new_n3112_), .Y(u2__abc_52155_new_n3113_));
OR2X2 OR2X2_5330 ( .A(u2__abc_52155_new_n23320_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23321_));
OR2X2 OR2X2_5331 ( .A(u2__abc_52155_new_n23325_), .B(u2__abc_52155_new_n23316_), .Y(u2__abc_52155_new_n23326_));
OR2X2 OR2X2_5332 ( .A(u2__abc_52155_new_n23317_), .B(u2_o_354_), .Y(u2__abc_52155_new_n23329_));
OR2X2 OR2X2_5333 ( .A(u2__abc_52155_new_n23332_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23333_));
OR2X2 OR2X2_5334 ( .A(u2__abc_52155_new_n23337_), .B(u2__abc_52155_new_n23328_), .Y(u2__abc_52155_new_n23338_));
OR2X2 OR2X2_5335 ( .A(u2__abc_52155_new_n23330_), .B(u2_o_355_), .Y(u2__abc_52155_new_n23341_));
OR2X2 OR2X2_5336 ( .A(u2__abc_52155_new_n23344_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23345_));
OR2X2 OR2X2_5337 ( .A(u2__abc_52155_new_n23349_), .B(u2__abc_52155_new_n23340_), .Y(u2__abc_52155_new_n23350_));
OR2X2 OR2X2_5338 ( .A(u2__abc_52155_new_n23342_), .B(u2_o_356_), .Y(u2__abc_52155_new_n23353_));
OR2X2 OR2X2_5339 ( .A(u2__abc_52155_new_n23356_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23357_));
OR2X2 OR2X2_534 ( .A(u2__abc_52155_new_n3115_), .B(u2__abc_52155_new_n3117_), .Y(u2__abc_52155_new_n3118_));
OR2X2 OR2X2_5340 ( .A(u2__abc_52155_new_n23361_), .B(u2__abc_52155_new_n23352_), .Y(u2__abc_52155_new_n23362_));
OR2X2 OR2X2_5341 ( .A(u2__abc_52155_new_n23354_), .B(u2_o_357_), .Y(u2__abc_52155_new_n23367_));
OR2X2 OR2X2_5342 ( .A(u2__abc_52155_new_n23368_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23369_));
OR2X2 OR2X2_5343 ( .A(u2__abc_52155_new_n23373_), .B(u2__abc_52155_new_n23364_), .Y(u2__abc_52155_new_n23374_));
OR2X2 OR2X2_5344 ( .A(u2__abc_52155_new_n23365_), .B(u2_o_358_), .Y(u2__abc_52155_new_n23377_));
OR2X2 OR2X2_5345 ( .A(u2__abc_52155_new_n23380_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23381_));
OR2X2 OR2X2_5346 ( .A(u2__abc_52155_new_n23385_), .B(u2__abc_52155_new_n23376_), .Y(u2__abc_52155_new_n23386_));
OR2X2 OR2X2_5347 ( .A(u2__abc_52155_new_n23378_), .B(u2_o_359_), .Y(u2__abc_52155_new_n23391_));
OR2X2 OR2X2_5348 ( .A(u2__abc_52155_new_n23392_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23393_));
OR2X2 OR2X2_5349 ( .A(u2__abc_52155_new_n23397_), .B(u2__abc_52155_new_n23388_), .Y(u2__abc_52155_new_n23398_));
OR2X2 OR2X2_535 ( .A(u2__abc_52155_new_n3120_), .B(u2__abc_52155_new_n3122_), .Y(u2__abc_52155_new_n3123_));
OR2X2 OR2X2_5350 ( .A(u2__abc_52155_new_n23389_), .B(u2_o_360_), .Y(u2__abc_52155_new_n23401_));
OR2X2 OR2X2_5351 ( .A(u2__abc_52155_new_n23404_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23405_));
OR2X2 OR2X2_5352 ( .A(u2__abc_52155_new_n23409_), .B(u2__abc_52155_new_n23400_), .Y(u2__abc_52155_new_n23410_));
OR2X2 OR2X2_5353 ( .A(u2__abc_52155_new_n23402_), .B(u2_o_361_), .Y(u2__abc_52155_new_n23415_));
OR2X2 OR2X2_5354 ( .A(u2__abc_52155_new_n23416_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23417_));
OR2X2 OR2X2_5355 ( .A(u2__abc_52155_new_n23421_), .B(u2__abc_52155_new_n23412_), .Y(u2__abc_52155_new_n23422_));
OR2X2 OR2X2_5356 ( .A(u2__abc_52155_new_n23413_), .B(u2_o_362_), .Y(u2__abc_52155_new_n23425_));
OR2X2 OR2X2_5357 ( .A(u2__abc_52155_new_n23428_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23429_));
OR2X2 OR2X2_5358 ( .A(u2__abc_52155_new_n23433_), .B(u2__abc_52155_new_n23424_), .Y(u2__abc_52155_new_n23434_));
OR2X2 OR2X2_5359 ( .A(u2__abc_52155_new_n23426_), .B(u2_o_363_), .Y(u2__abc_52155_new_n23439_));
OR2X2 OR2X2_536 ( .A(u2__abc_52155_new_n3118_), .B(u2__abc_52155_new_n3123_), .Y(u2__abc_52155_new_n3124_));
OR2X2 OR2X2_5360 ( .A(u2__abc_52155_new_n23440_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23441_));
OR2X2 OR2X2_5361 ( .A(u2__abc_52155_new_n23445_), .B(u2__abc_52155_new_n23436_), .Y(u2__abc_52155_new_n23446_));
OR2X2 OR2X2_5362 ( .A(u2__abc_52155_new_n23437_), .B(u2_o_364_), .Y(u2__abc_52155_new_n23449_));
OR2X2 OR2X2_5363 ( .A(u2__abc_52155_new_n23452_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23453_));
OR2X2 OR2X2_5364 ( .A(u2__abc_52155_new_n23457_), .B(u2__abc_52155_new_n23448_), .Y(u2__abc_52155_new_n23458_));
OR2X2 OR2X2_5365 ( .A(u2__abc_52155_new_n23450_), .B(u2_o_365_), .Y(u2__abc_52155_new_n23463_));
OR2X2 OR2X2_5366 ( .A(u2__abc_52155_new_n23464_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23465_));
OR2X2 OR2X2_5367 ( .A(u2__abc_52155_new_n23469_), .B(u2__abc_52155_new_n23460_), .Y(u2__abc_52155_new_n23470_));
OR2X2 OR2X2_5368 ( .A(u2__abc_52155_new_n23461_), .B(u2_o_366_), .Y(u2__abc_52155_new_n23473_));
OR2X2 OR2X2_5369 ( .A(u2__abc_52155_new_n23476_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23477_));
OR2X2 OR2X2_537 ( .A(u2__abc_52155_new_n3124_), .B(u2__abc_52155_new_n3126_), .Y(u2__abc_52155_new_n3127_));
OR2X2 OR2X2_5370 ( .A(u2__abc_52155_new_n23481_), .B(u2__abc_52155_new_n23472_), .Y(u2__abc_52155_new_n23482_));
OR2X2 OR2X2_5371 ( .A(u2__abc_52155_new_n23474_), .B(u2_o_367_), .Y(u2__abc_52155_new_n23487_));
OR2X2 OR2X2_5372 ( .A(u2__abc_52155_new_n23488_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23489_));
OR2X2 OR2X2_5373 ( .A(u2__abc_52155_new_n23493_), .B(u2__abc_52155_new_n23484_), .Y(u2__abc_52155_new_n23494_));
OR2X2 OR2X2_5374 ( .A(u2__abc_52155_new_n23485_), .B(u2_o_368_), .Y(u2__abc_52155_new_n23497_));
OR2X2 OR2X2_5375 ( .A(u2__abc_52155_new_n23500_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23501_));
OR2X2 OR2X2_5376 ( .A(u2__abc_52155_new_n23505_), .B(u2__abc_52155_new_n23496_), .Y(u2__abc_52155_new_n23506_));
OR2X2 OR2X2_5377 ( .A(u2__abc_52155_new_n23498_), .B(u2_o_369_), .Y(u2__abc_52155_new_n23511_));
OR2X2 OR2X2_5378 ( .A(u2__abc_52155_new_n23512_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23513_));
OR2X2 OR2X2_5379 ( .A(u2__abc_52155_new_n23517_), .B(u2__abc_52155_new_n23508_), .Y(u2__abc_52155_new_n23518_));
OR2X2 OR2X2_538 ( .A(u2__abc_52155_new_n3129_), .B(u2__abc_52155_new_n3122_), .Y(u2__abc_52155_new_n3130_));
OR2X2 OR2X2_5380 ( .A(u2__abc_52155_new_n23509_), .B(u2_o_370_), .Y(u2__abc_52155_new_n23521_));
OR2X2 OR2X2_5381 ( .A(u2__abc_52155_new_n23524_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23525_));
OR2X2 OR2X2_5382 ( .A(u2__abc_52155_new_n23529_), .B(u2__abc_52155_new_n23520_), .Y(u2__abc_52155_new_n23530_));
OR2X2 OR2X2_5383 ( .A(u2__abc_52155_new_n23522_), .B(u2_o_371_), .Y(u2__abc_52155_new_n23535_));
OR2X2 OR2X2_5384 ( .A(u2__abc_52155_new_n23536_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23537_));
OR2X2 OR2X2_5385 ( .A(u2__abc_52155_new_n23541_), .B(u2__abc_52155_new_n23532_), .Y(u2__abc_52155_new_n23542_));
OR2X2 OR2X2_5386 ( .A(u2__abc_52155_new_n23533_), .B(u2_o_372_), .Y(u2__abc_52155_new_n23545_));
OR2X2 OR2X2_5387 ( .A(u2__abc_52155_new_n23548_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23549_));
OR2X2 OR2X2_5388 ( .A(u2__abc_52155_new_n23553_), .B(u2__abc_52155_new_n23544_), .Y(u2__abc_52155_new_n23554_));
OR2X2 OR2X2_5389 ( .A(u2__abc_52155_new_n23546_), .B(u2_o_373_), .Y(u2__abc_52155_new_n23559_));
OR2X2 OR2X2_539 ( .A(u2__abc_52155_new_n3132_), .B(u2__abc_52155_new_n3113_), .Y(u2__abc_52155_new_n3133_));
OR2X2 OR2X2_5390 ( .A(u2__abc_52155_new_n23560_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23561_));
OR2X2 OR2X2_5391 ( .A(u2__abc_52155_new_n23565_), .B(u2__abc_52155_new_n23556_), .Y(u2__abc_52155_new_n23566_));
OR2X2 OR2X2_5392 ( .A(u2__abc_52155_new_n23557_), .B(u2_o_374_), .Y(u2__abc_52155_new_n23569_));
OR2X2 OR2X2_5393 ( .A(u2__abc_52155_new_n23572_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23573_));
OR2X2 OR2X2_5394 ( .A(u2__abc_52155_new_n23577_), .B(u2__abc_52155_new_n23568_), .Y(u2__abc_52155_new_n23578_));
OR2X2 OR2X2_5395 ( .A(u2__abc_52155_new_n23570_), .B(u2_o_375_), .Y(u2__abc_52155_new_n23583_));
OR2X2 OR2X2_5396 ( .A(u2__abc_52155_new_n23584_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23585_));
OR2X2 OR2X2_5397 ( .A(u2__abc_52155_new_n23589_), .B(u2__abc_52155_new_n23580_), .Y(u2__abc_52155_new_n23590_));
OR2X2 OR2X2_5398 ( .A(u2__abc_52155_new_n23581_), .B(u2_o_376_), .Y(u2__abc_52155_new_n23593_));
OR2X2 OR2X2_5399 ( .A(u2__abc_52155_new_n23596_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23597_));
OR2X2 OR2X2_54 ( .A(_abc_73687_new_n753_), .B(\a[26] ), .Y(_abc_73687_new_n909_));
OR2X2 OR2X2_540 ( .A(u2__abc_52155_new_n3135_), .B(u2__abc_52155_new_n3103_), .Y(u2__abc_52155_new_n3136_));
OR2X2 OR2X2_5400 ( .A(u2__abc_52155_new_n23601_), .B(u2__abc_52155_new_n23592_), .Y(u2__abc_52155_new_n23602_));
OR2X2 OR2X2_5401 ( .A(u2__abc_52155_new_n23594_), .B(u2_o_377_), .Y(u2__abc_52155_new_n23607_));
OR2X2 OR2X2_5402 ( .A(u2__abc_52155_new_n23608_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23609_));
OR2X2 OR2X2_5403 ( .A(u2__abc_52155_new_n23613_), .B(u2__abc_52155_new_n23604_), .Y(u2__abc_52155_new_n23614_));
OR2X2 OR2X2_5404 ( .A(u2__abc_52155_new_n23605_), .B(u2_o_378_), .Y(u2__abc_52155_new_n23617_));
OR2X2 OR2X2_5405 ( .A(u2__abc_52155_new_n23620_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23621_));
OR2X2 OR2X2_5406 ( .A(u2__abc_52155_new_n23625_), .B(u2__abc_52155_new_n23616_), .Y(u2__abc_52155_new_n23626_));
OR2X2 OR2X2_5407 ( .A(u2__abc_52155_new_n23618_), .B(u2_o_379_), .Y(u2__abc_52155_new_n23631_));
OR2X2 OR2X2_5408 ( .A(u2__abc_52155_new_n23632_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23633_));
OR2X2 OR2X2_5409 ( .A(u2__abc_52155_new_n23637_), .B(u2__abc_52155_new_n23628_), .Y(u2__abc_52155_new_n23638_));
OR2X2 OR2X2_541 ( .A(u2__abc_52155_new_n3137_), .B(u2__abc_52155_new_n3101_), .Y(u2__abc_52155_new_n3138_));
OR2X2 OR2X2_5410 ( .A(u2__abc_52155_new_n23629_), .B(u2_o_380_), .Y(u2__abc_52155_new_n23641_));
OR2X2 OR2X2_5411 ( .A(u2__abc_52155_new_n23644_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23645_));
OR2X2 OR2X2_5412 ( .A(u2__abc_52155_new_n23649_), .B(u2__abc_52155_new_n23640_), .Y(u2__abc_52155_new_n23650_));
OR2X2 OR2X2_5413 ( .A(u2__abc_52155_new_n23642_), .B(u2_o_381_), .Y(u2__abc_52155_new_n23655_));
OR2X2 OR2X2_5414 ( .A(u2__abc_52155_new_n23656_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23657_));
OR2X2 OR2X2_5415 ( .A(u2__abc_52155_new_n23661_), .B(u2__abc_52155_new_n23652_), .Y(u2__abc_52155_new_n23662_));
OR2X2 OR2X2_5416 ( .A(u2__abc_52155_new_n23653_), .B(u2_o_382_), .Y(u2__abc_52155_new_n23665_));
OR2X2 OR2X2_5417 ( .A(u2__abc_52155_new_n23668_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23669_));
OR2X2 OR2X2_5418 ( .A(u2__abc_52155_new_n23673_), .B(u2__abc_52155_new_n23664_), .Y(u2__abc_52155_new_n23674_));
OR2X2 OR2X2_5419 ( .A(u2__abc_52155_new_n23666_), .B(u2_o_383_), .Y(u2__abc_52155_new_n23679_));
OR2X2 OR2X2_542 ( .A(u2__abc_52155_new_n3140_), .B(u2__abc_52155_new_n3099_), .Y(u2__abc_52155_new_n3141_));
OR2X2 OR2X2_5420 ( .A(u2__abc_52155_new_n23680_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23681_));
OR2X2 OR2X2_5421 ( .A(u2__abc_52155_new_n23685_), .B(u2__abc_52155_new_n23676_), .Y(u2__abc_52155_new_n23686_));
OR2X2 OR2X2_5422 ( .A(u2__abc_52155_new_n23677_), .B(u2_o_384_), .Y(u2__abc_52155_new_n23689_));
OR2X2 OR2X2_5423 ( .A(u2__abc_52155_new_n23692_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23693_));
OR2X2 OR2X2_5424 ( .A(u2__abc_52155_new_n23697_), .B(u2__abc_52155_new_n23688_), .Y(u2__abc_52155_new_n23698_));
OR2X2 OR2X2_5425 ( .A(u2__abc_52155_new_n23690_), .B(u2_o_385_), .Y(u2__abc_52155_new_n23703_));
OR2X2 OR2X2_5426 ( .A(u2__abc_52155_new_n23704_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23705_));
OR2X2 OR2X2_5427 ( .A(u2__abc_52155_new_n23709_), .B(u2__abc_52155_new_n23700_), .Y(u2__abc_52155_new_n23710_));
OR2X2 OR2X2_5428 ( .A(u2__abc_52155_new_n23701_), .B(u2_o_386_), .Y(u2__abc_52155_new_n23713_));
OR2X2 OR2X2_5429 ( .A(u2__abc_52155_new_n23716_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23717_));
OR2X2 OR2X2_543 ( .A(u2__abc_52155_new_n3144_), .B(u2__abc_52155_new_n3090_), .Y(u2__abc_52155_new_n3145_));
OR2X2 OR2X2_5430 ( .A(u2__abc_52155_new_n23721_), .B(u2__abc_52155_new_n23712_), .Y(u2__abc_52155_new_n23722_));
OR2X2 OR2X2_5431 ( .A(u2__abc_52155_new_n23714_), .B(u2_o_387_), .Y(u2__abc_52155_new_n23725_));
OR2X2 OR2X2_5432 ( .A(u2__abc_52155_new_n23728_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23729_));
OR2X2 OR2X2_5433 ( .A(u2__abc_52155_new_n23733_), .B(u2__abc_52155_new_n23724_), .Y(u2__abc_52155_new_n23734_));
OR2X2 OR2X2_5434 ( .A(u2__abc_52155_new_n23726_), .B(u2_o_388_), .Y(u2__abc_52155_new_n23737_));
OR2X2 OR2X2_5435 ( .A(u2__abc_52155_new_n23740_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23741_));
OR2X2 OR2X2_5436 ( .A(u2__abc_52155_new_n23745_), .B(u2__abc_52155_new_n23736_), .Y(u2__abc_52155_new_n23746_));
OR2X2 OR2X2_5437 ( .A(u2__abc_52155_new_n23738_), .B(u2_o_389_), .Y(u2__abc_52155_new_n23751_));
OR2X2 OR2X2_5438 ( .A(u2__abc_52155_new_n23752_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23753_));
OR2X2 OR2X2_5439 ( .A(u2__abc_52155_new_n23757_), .B(u2__abc_52155_new_n23748_), .Y(u2__abc_52155_new_n23758_));
OR2X2 OR2X2_544 ( .A(u2__abc_52155_new_n3085_), .B(u2__abc_52155_new_n3078_), .Y(u2__abc_52155_new_n3148_));
OR2X2 OR2X2_5440 ( .A(u2__abc_52155_new_n23749_), .B(u2_o_390_), .Y(u2__abc_52155_new_n23761_));
OR2X2 OR2X2_5441 ( .A(u2__abc_52155_new_n23764_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23765_));
OR2X2 OR2X2_5442 ( .A(u2__abc_52155_new_n23769_), .B(u2__abc_52155_new_n23760_), .Y(u2__abc_52155_new_n23770_));
OR2X2 OR2X2_5443 ( .A(u2__abc_52155_new_n23762_), .B(u2_o_391_), .Y(u2__abc_52155_new_n23773_));
OR2X2 OR2X2_5444 ( .A(u2__abc_52155_new_n23776_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23777_));
OR2X2 OR2X2_5445 ( .A(u2__abc_52155_new_n23781_), .B(u2__abc_52155_new_n23772_), .Y(u2__abc_52155_new_n23782_));
OR2X2 OR2X2_5446 ( .A(u2__abc_52155_new_n23774_), .B(u2_o_392_), .Y(u2__abc_52155_new_n23785_));
OR2X2 OR2X2_5447 ( .A(u2__abc_52155_new_n23788_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23789_));
OR2X2 OR2X2_5448 ( .A(u2__abc_52155_new_n23793_), .B(u2__abc_52155_new_n23784_), .Y(u2__abc_52155_new_n23794_));
OR2X2 OR2X2_5449 ( .A(u2__abc_52155_new_n23786_), .B(u2_o_393_), .Y(u2__abc_52155_new_n23799_));
OR2X2 OR2X2_545 ( .A(u2__abc_52155_new_n3147_), .B(u2__abc_52155_new_n3149_), .Y(u2__abc_52155_new_n3150_));
OR2X2 OR2X2_5450 ( .A(u2__abc_52155_new_n23800_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23801_));
OR2X2 OR2X2_5451 ( .A(u2__abc_52155_new_n23805_), .B(u2__abc_52155_new_n23796_), .Y(u2__abc_52155_new_n23806_));
OR2X2 OR2X2_5452 ( .A(u2__abc_52155_new_n23797_), .B(u2_o_394_), .Y(u2__abc_52155_new_n23809_));
OR2X2 OR2X2_5453 ( .A(u2__abc_52155_new_n23812_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23813_));
OR2X2 OR2X2_5454 ( .A(u2__abc_52155_new_n23817_), .B(u2__abc_52155_new_n23808_), .Y(u2__abc_52155_new_n23818_));
OR2X2 OR2X2_5455 ( .A(u2__abc_52155_new_n23810_), .B(u2_o_395_), .Y(u2__abc_52155_new_n23821_));
OR2X2 OR2X2_5456 ( .A(u2__abc_52155_new_n23824_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23825_));
OR2X2 OR2X2_5457 ( .A(u2__abc_52155_new_n23829_), .B(u2__abc_52155_new_n23820_), .Y(u2__abc_52155_new_n23830_));
OR2X2 OR2X2_5458 ( .A(u2__abc_52155_new_n23822_), .B(u2_o_396_), .Y(u2__abc_52155_new_n23833_));
OR2X2 OR2X2_5459 ( .A(u2__abc_52155_new_n23836_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23837_));
OR2X2 OR2X2_546 ( .A(u2__abc_52155_new_n3154_), .B(u2__abc_52155_new_n3146_), .Y(u2__abc_52155_new_n3155_));
OR2X2 OR2X2_5460 ( .A(u2__abc_52155_new_n23841_), .B(u2__abc_52155_new_n23832_), .Y(u2__abc_52155_new_n23842_));
OR2X2 OR2X2_5461 ( .A(u2__abc_52155_new_n23834_), .B(u2_o_397_), .Y(u2__abc_52155_new_n23847_));
OR2X2 OR2X2_5462 ( .A(u2__abc_52155_new_n23848_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23849_));
OR2X2 OR2X2_5463 ( .A(u2__abc_52155_new_n23853_), .B(u2__abc_52155_new_n23844_), .Y(u2__abc_52155_new_n23854_));
OR2X2 OR2X2_5464 ( .A(u2__abc_52155_new_n23845_), .B(u2_o_398_), .Y(u2__abc_52155_new_n23857_));
OR2X2 OR2X2_5465 ( .A(u2__abc_52155_new_n23860_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23861_));
OR2X2 OR2X2_5466 ( .A(u2__abc_52155_new_n23865_), .B(u2__abc_52155_new_n23856_), .Y(u2__abc_52155_new_n23866_));
OR2X2 OR2X2_5467 ( .A(u2__abc_52155_new_n23858_), .B(u2_o_399_), .Y(u2__abc_52155_new_n23871_));
OR2X2 OR2X2_5468 ( .A(u2__abc_52155_new_n23872_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23873_));
OR2X2 OR2X2_5469 ( .A(u2__abc_52155_new_n23877_), .B(u2__abc_52155_new_n23868_), .Y(u2__abc_52155_new_n23878_));
OR2X2 OR2X2_547 ( .A(u2__abc_52155_new_n3156_), .B(u2__abc_52155_new_n3042_), .Y(u2__abc_52155_new_n3157_));
OR2X2 OR2X2_5470 ( .A(u2__abc_52155_new_n23869_), .B(u2_o_400_), .Y(u2__abc_52155_new_n23881_));
OR2X2 OR2X2_5471 ( .A(u2__abc_52155_new_n23884_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23885_));
OR2X2 OR2X2_5472 ( .A(u2__abc_52155_new_n23889_), .B(u2__abc_52155_new_n23880_), .Y(u2__abc_52155_new_n23890_));
OR2X2 OR2X2_5473 ( .A(u2__abc_52155_new_n23882_), .B(u2_o_401_), .Y(u2__abc_52155_new_n23895_));
OR2X2 OR2X2_5474 ( .A(u2__abc_52155_new_n23896_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23897_));
OR2X2 OR2X2_5475 ( .A(u2__abc_52155_new_n23901_), .B(u2__abc_52155_new_n23892_), .Y(u2__abc_52155_new_n23902_));
OR2X2 OR2X2_5476 ( .A(u2__abc_52155_new_n23893_), .B(u2_o_402_), .Y(u2__abc_52155_new_n23905_));
OR2X2 OR2X2_5477 ( .A(u2__abc_52155_new_n23908_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23909_));
OR2X2 OR2X2_5478 ( .A(u2__abc_52155_new_n23913_), .B(u2__abc_52155_new_n23904_), .Y(u2__abc_52155_new_n23914_));
OR2X2 OR2X2_5479 ( .A(u2__abc_52155_new_n23906_), .B(u2_o_403_), .Y(u2__abc_52155_new_n23917_));
OR2X2 OR2X2_548 ( .A(u2__abc_52155_new_n3159_), .B(u2__abc_52155_new_n3162_), .Y(u2__abc_52155_new_n3163_));
OR2X2 OR2X2_5480 ( .A(u2__abc_52155_new_n23920_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23921_));
OR2X2 OR2X2_5481 ( .A(u2__abc_52155_new_n23925_), .B(u2__abc_52155_new_n23916_), .Y(u2__abc_52155_new_n23926_));
OR2X2 OR2X2_5482 ( .A(u2__abc_52155_new_n23918_), .B(u2_o_404_), .Y(u2__abc_52155_new_n23929_));
OR2X2 OR2X2_5483 ( .A(u2__abc_52155_new_n23932_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23933_));
OR2X2 OR2X2_5484 ( .A(u2__abc_52155_new_n23937_), .B(u2__abc_52155_new_n23928_), .Y(u2__abc_52155_new_n23938_));
OR2X2 OR2X2_5485 ( .A(u2__abc_52155_new_n23930_), .B(u2_o_405_), .Y(u2__abc_52155_new_n23943_));
OR2X2 OR2X2_5486 ( .A(u2__abc_52155_new_n23944_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23945_));
OR2X2 OR2X2_5487 ( .A(u2__abc_52155_new_n23949_), .B(u2__abc_52155_new_n23940_), .Y(u2__abc_52155_new_n23950_));
OR2X2 OR2X2_5488 ( .A(u2__abc_52155_new_n23941_), .B(u2_o_406_), .Y(u2__abc_52155_new_n23953_));
OR2X2 OR2X2_5489 ( .A(u2__abc_52155_new_n23956_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23957_));
OR2X2 OR2X2_549 ( .A(u2__abc_52155_new_n3168_), .B(u2__abc_52155_new_n3170_), .Y(u2__abc_52155_new_n3171_));
OR2X2 OR2X2_5490 ( .A(u2__abc_52155_new_n23961_), .B(u2__abc_52155_new_n23952_), .Y(u2__abc_52155_new_n23962_));
OR2X2 OR2X2_5491 ( .A(u2__abc_52155_new_n23954_), .B(u2_o_407_), .Y(u2__abc_52155_new_n23967_));
OR2X2 OR2X2_5492 ( .A(u2__abc_52155_new_n23968_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23969_));
OR2X2 OR2X2_5493 ( .A(u2__abc_52155_new_n23973_), .B(u2__abc_52155_new_n23964_), .Y(u2__abc_52155_new_n23974_));
OR2X2 OR2X2_5494 ( .A(u2__abc_52155_new_n23965_), .B(u2_o_408_), .Y(u2__abc_52155_new_n23977_));
OR2X2 OR2X2_5495 ( .A(u2__abc_52155_new_n23980_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23981_));
OR2X2 OR2X2_5496 ( .A(u2__abc_52155_new_n23985_), .B(u2__abc_52155_new_n23976_), .Y(u2__abc_52155_new_n23986_));
OR2X2 OR2X2_5497 ( .A(u2__abc_52155_new_n23978_), .B(u2_o_409_), .Y(u2__abc_52155_new_n23991_));
OR2X2 OR2X2_5498 ( .A(u2__abc_52155_new_n23992_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n23993_));
OR2X2 OR2X2_5499 ( .A(u2__abc_52155_new_n23997_), .B(u2__abc_52155_new_n23988_), .Y(u2__abc_52155_new_n23998_));
OR2X2 OR2X2_55 ( .A(aNan), .B(sqrto_103_), .Y(_abc_73687_new_n911_));
OR2X2 OR2X2_550 ( .A(u2__abc_52155_new_n3173_), .B(u2__abc_52155_new_n3175_), .Y(u2__abc_52155_new_n3176_));
OR2X2 OR2X2_5500 ( .A(u2__abc_52155_new_n23989_), .B(u2_o_410_), .Y(u2__abc_52155_new_n24001_));
OR2X2 OR2X2_5501 ( .A(u2__abc_52155_new_n24004_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24005_));
OR2X2 OR2X2_5502 ( .A(u2__abc_52155_new_n24009_), .B(u2__abc_52155_new_n24000_), .Y(u2__abc_52155_new_n24010_));
OR2X2 OR2X2_5503 ( .A(u2__abc_52155_new_n24002_), .B(u2_o_411_), .Y(u2__abc_52155_new_n24015_));
OR2X2 OR2X2_5504 ( .A(u2__abc_52155_new_n24016_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24017_));
OR2X2 OR2X2_5505 ( .A(u2__abc_52155_new_n24021_), .B(u2__abc_52155_new_n24012_), .Y(u2__abc_52155_new_n24022_));
OR2X2 OR2X2_5506 ( .A(u2__abc_52155_new_n24013_), .B(u2_o_412_), .Y(u2__abc_52155_new_n24025_));
OR2X2 OR2X2_5507 ( .A(u2__abc_52155_new_n24028_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24029_));
OR2X2 OR2X2_5508 ( .A(u2__abc_52155_new_n24033_), .B(u2__abc_52155_new_n24024_), .Y(u2__abc_52155_new_n24034_));
OR2X2 OR2X2_5509 ( .A(u2__abc_52155_new_n24026_), .B(u2_o_413_), .Y(u2__abc_52155_new_n24039_));
OR2X2 OR2X2_551 ( .A(u2__abc_52155_new_n3171_), .B(u2__abc_52155_new_n3176_), .Y(u2__abc_52155_new_n3177_));
OR2X2 OR2X2_5510 ( .A(u2__abc_52155_new_n24040_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24041_));
OR2X2 OR2X2_5511 ( .A(u2__abc_52155_new_n24045_), .B(u2__abc_52155_new_n24036_), .Y(u2__abc_52155_new_n24046_));
OR2X2 OR2X2_5512 ( .A(u2__abc_52155_new_n24037_), .B(u2_o_414_), .Y(u2__abc_52155_new_n24049_));
OR2X2 OR2X2_5513 ( .A(u2__abc_52155_new_n24052_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24053_));
OR2X2 OR2X2_5514 ( .A(u2__abc_52155_new_n24057_), .B(u2__abc_52155_new_n24048_), .Y(u2__abc_52155_new_n24058_));
OR2X2 OR2X2_5515 ( .A(u2__abc_52155_new_n24050_), .B(u2_o_415_), .Y(u2__abc_52155_new_n24063_));
OR2X2 OR2X2_5516 ( .A(u2__abc_52155_new_n24064_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24065_));
OR2X2 OR2X2_5517 ( .A(u2__abc_52155_new_n24069_), .B(u2__abc_52155_new_n24060_), .Y(u2__abc_52155_new_n24070_));
OR2X2 OR2X2_5518 ( .A(u2__abc_52155_new_n24061_), .B(u2_o_416_), .Y(u2__abc_52155_new_n24073_));
OR2X2 OR2X2_5519 ( .A(u2__abc_52155_new_n24076_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24077_));
OR2X2 OR2X2_552 ( .A(u2__abc_52155_new_n3228_), .B(u2__abc_52155_new_n3230_), .Y(u2__abc_52155_new_n3231_));
OR2X2 OR2X2_5520 ( .A(u2__abc_52155_new_n24081_), .B(u2__abc_52155_new_n24072_), .Y(u2__abc_52155_new_n24082_));
OR2X2 OR2X2_5521 ( .A(u2__abc_52155_new_n24074_), .B(u2_o_417_), .Y(u2__abc_52155_new_n24087_));
OR2X2 OR2X2_5522 ( .A(u2__abc_52155_new_n24088_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24089_));
OR2X2 OR2X2_5523 ( .A(u2__abc_52155_new_n24093_), .B(u2__abc_52155_new_n24084_), .Y(u2__abc_52155_new_n24094_));
OR2X2 OR2X2_5524 ( .A(u2__abc_52155_new_n24085_), .B(u2_o_418_), .Y(u2__abc_52155_new_n24097_));
OR2X2 OR2X2_5525 ( .A(u2__abc_52155_new_n24100_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24101_));
OR2X2 OR2X2_5526 ( .A(u2__abc_52155_new_n24105_), .B(u2__abc_52155_new_n24096_), .Y(u2__abc_52155_new_n24106_));
OR2X2 OR2X2_5527 ( .A(u2__abc_52155_new_n24098_), .B(u2_o_419_), .Y(u2__abc_52155_new_n24109_));
OR2X2 OR2X2_5528 ( .A(u2__abc_52155_new_n24112_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24113_));
OR2X2 OR2X2_5529 ( .A(u2__abc_52155_new_n24117_), .B(u2__abc_52155_new_n24108_), .Y(u2__abc_52155_new_n24118_));
OR2X2 OR2X2_553 ( .A(u2__abc_52155_new_n3233_), .B(u2__abc_52155_new_n3235_), .Y(u2__abc_52155_new_n3236_));
OR2X2 OR2X2_5530 ( .A(u2__abc_52155_new_n24110_), .B(u2_o_420_), .Y(u2__abc_52155_new_n24121_));
OR2X2 OR2X2_5531 ( .A(u2__abc_52155_new_n24124_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24125_));
OR2X2 OR2X2_5532 ( .A(u2__abc_52155_new_n24129_), .B(u2__abc_52155_new_n24120_), .Y(u2__abc_52155_new_n24130_));
OR2X2 OR2X2_5533 ( .A(u2__abc_52155_new_n24122_), .B(u2_o_421_), .Y(u2__abc_52155_new_n24135_));
OR2X2 OR2X2_5534 ( .A(u2__abc_52155_new_n24136_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24137_));
OR2X2 OR2X2_5535 ( .A(u2__abc_52155_new_n24141_), .B(u2__abc_52155_new_n24132_), .Y(u2__abc_52155_new_n24142_));
OR2X2 OR2X2_5536 ( .A(u2__abc_52155_new_n24133_), .B(u2_o_422_), .Y(u2__abc_52155_new_n24145_));
OR2X2 OR2X2_5537 ( .A(u2__abc_52155_new_n24148_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24149_));
OR2X2 OR2X2_5538 ( .A(u2__abc_52155_new_n24153_), .B(u2__abc_52155_new_n24144_), .Y(u2__abc_52155_new_n24154_));
OR2X2 OR2X2_5539 ( .A(u2__abc_52155_new_n24146_), .B(u2_o_423_), .Y(u2__abc_52155_new_n24159_));
OR2X2 OR2X2_554 ( .A(u2__abc_52155_new_n3231_), .B(u2__abc_52155_new_n3236_), .Y(u2__abc_52155_new_n3237_));
OR2X2 OR2X2_5540 ( .A(u2__abc_52155_new_n24160_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24161_));
OR2X2 OR2X2_5541 ( .A(u2__abc_52155_new_n24165_), .B(u2__abc_52155_new_n24156_), .Y(u2__abc_52155_new_n24166_));
OR2X2 OR2X2_5542 ( .A(u2__abc_52155_new_n24157_), .B(u2_o_424_), .Y(u2__abc_52155_new_n24169_));
OR2X2 OR2X2_5543 ( .A(u2__abc_52155_new_n24172_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24173_));
OR2X2 OR2X2_5544 ( .A(u2__abc_52155_new_n24177_), .B(u2__abc_52155_new_n24168_), .Y(u2__abc_52155_new_n24178_));
OR2X2 OR2X2_5545 ( .A(u2__abc_52155_new_n24170_), .B(u2_o_425_), .Y(u2__abc_52155_new_n24183_));
OR2X2 OR2X2_5546 ( .A(u2__abc_52155_new_n24184_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24185_));
OR2X2 OR2X2_5547 ( .A(u2__abc_52155_new_n24189_), .B(u2__abc_52155_new_n24180_), .Y(u2__abc_52155_new_n24190_));
OR2X2 OR2X2_5548 ( .A(u2__abc_52155_new_n24181_), .B(u2_o_426_), .Y(u2__abc_52155_new_n24193_));
OR2X2 OR2X2_5549 ( .A(u2__abc_52155_new_n24196_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24197_));
OR2X2 OR2X2_555 ( .A(u2__abc_52155_new_n3239_), .B(u2_remHi_14_), .Y(u2__abc_52155_new_n3242_));
OR2X2 OR2X2_5550 ( .A(u2__abc_52155_new_n24201_), .B(u2__abc_52155_new_n24192_), .Y(u2__abc_52155_new_n24202_));
OR2X2 OR2X2_5551 ( .A(u2__abc_52155_new_n24194_), .B(u2_o_427_), .Y(u2__abc_52155_new_n24207_));
OR2X2 OR2X2_5552 ( .A(u2__abc_52155_new_n24208_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24209_));
OR2X2 OR2X2_5553 ( .A(u2__abc_52155_new_n24213_), .B(u2__abc_52155_new_n24204_), .Y(u2__abc_52155_new_n24214_));
OR2X2 OR2X2_5554 ( .A(u2__abc_52155_new_n24205_), .B(u2_o_428_), .Y(u2__abc_52155_new_n24217_));
OR2X2 OR2X2_5555 ( .A(u2__abc_52155_new_n24220_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24221_));
OR2X2 OR2X2_5556 ( .A(u2__abc_52155_new_n24225_), .B(u2__abc_52155_new_n24216_), .Y(u2__abc_52155_new_n24226_));
OR2X2 OR2X2_5557 ( .A(u2__abc_52155_new_n24218_), .B(u2_o_429_), .Y(u2__abc_52155_new_n24231_));
OR2X2 OR2X2_5558 ( .A(u2__abc_52155_new_n24232_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24233_));
OR2X2 OR2X2_5559 ( .A(u2__abc_52155_new_n24237_), .B(u2__abc_52155_new_n24228_), .Y(u2__abc_52155_new_n24238_));
OR2X2 OR2X2_556 ( .A(u2__abc_52155_new_n3254_), .B(u2__abc_52155_new_n3256_), .Y(u2__abc_52155_new_n3257_));
OR2X2 OR2X2_5560 ( .A(u2__abc_52155_new_n24229_), .B(u2_o_430_), .Y(u2__abc_52155_new_n24241_));
OR2X2 OR2X2_5561 ( .A(u2__abc_52155_new_n24244_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24245_));
OR2X2 OR2X2_5562 ( .A(u2__abc_52155_new_n24249_), .B(u2__abc_52155_new_n24240_), .Y(u2__abc_52155_new_n24250_));
OR2X2 OR2X2_5563 ( .A(u2__abc_52155_new_n24242_), .B(u2_o_431_), .Y(u2__abc_52155_new_n24255_));
OR2X2 OR2X2_5564 ( .A(u2__abc_52155_new_n24256_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24257_));
OR2X2 OR2X2_5565 ( .A(u2__abc_52155_new_n24261_), .B(u2__abc_52155_new_n24252_), .Y(u2__abc_52155_new_n24262_));
OR2X2 OR2X2_5566 ( .A(u2__abc_52155_new_n24253_), .B(u2_o_432_), .Y(u2__abc_52155_new_n24265_));
OR2X2 OR2X2_5567 ( .A(u2__abc_52155_new_n24268_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24269_));
OR2X2 OR2X2_5568 ( .A(u2__abc_52155_new_n24273_), .B(u2__abc_52155_new_n24264_), .Y(u2__abc_52155_new_n24274_));
OR2X2 OR2X2_5569 ( .A(u2__abc_52155_new_n24266_), .B(u2_o_433_), .Y(u2__abc_52155_new_n24279_));
OR2X2 OR2X2_557 ( .A(u2__abc_52155_new_n3259_), .B(u2__abc_52155_new_n3261_), .Y(u2__abc_52155_new_n3262_));
OR2X2 OR2X2_5570 ( .A(u2__abc_52155_new_n24280_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24281_));
OR2X2 OR2X2_5571 ( .A(u2__abc_52155_new_n24285_), .B(u2__abc_52155_new_n24276_), .Y(u2__abc_52155_new_n24286_));
OR2X2 OR2X2_5572 ( .A(u2__abc_52155_new_n24277_), .B(u2_o_434_), .Y(u2__abc_52155_new_n24289_));
OR2X2 OR2X2_5573 ( .A(u2__abc_52155_new_n24292_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24293_));
OR2X2 OR2X2_5574 ( .A(u2__abc_52155_new_n24297_), .B(u2__abc_52155_new_n24288_), .Y(u2__abc_52155_new_n24298_));
OR2X2 OR2X2_5575 ( .A(u2__abc_52155_new_n24290_), .B(u2_o_435_), .Y(u2__abc_52155_new_n24303_));
OR2X2 OR2X2_5576 ( .A(u2__abc_52155_new_n24304_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24305_));
OR2X2 OR2X2_5577 ( .A(u2__abc_52155_new_n24309_), .B(u2__abc_52155_new_n24300_), .Y(u2__abc_52155_new_n24310_));
OR2X2 OR2X2_5578 ( .A(u2__abc_52155_new_n24301_), .B(u2_o_436_), .Y(u2__abc_52155_new_n24313_));
OR2X2 OR2X2_5579 ( .A(u2__abc_52155_new_n24316_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24317_));
OR2X2 OR2X2_558 ( .A(u2__abc_52155_new_n3257_), .B(u2__abc_52155_new_n3262_), .Y(u2__abc_52155_new_n3263_));
OR2X2 OR2X2_5580 ( .A(u2__abc_52155_new_n24321_), .B(u2__abc_52155_new_n24312_), .Y(u2__abc_52155_new_n24322_));
OR2X2 OR2X2_5581 ( .A(u2__abc_52155_new_n24314_), .B(u2_o_437_), .Y(u2__abc_52155_new_n24327_));
OR2X2 OR2X2_5582 ( .A(u2__abc_52155_new_n24328_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24329_));
OR2X2 OR2X2_5583 ( .A(u2__abc_52155_new_n24333_), .B(u2__abc_52155_new_n24324_), .Y(u2__abc_52155_new_n24334_));
OR2X2 OR2X2_5584 ( .A(u2__abc_52155_new_n24325_), .B(u2_o_438_), .Y(u2__abc_52155_new_n24337_));
OR2X2 OR2X2_5585 ( .A(u2__abc_52155_new_n24340_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24341_));
OR2X2 OR2X2_5586 ( .A(u2__abc_52155_new_n24345_), .B(u2__abc_52155_new_n24336_), .Y(u2__abc_52155_new_n24346_));
OR2X2 OR2X2_5587 ( .A(u2__abc_52155_new_n24338_), .B(u2_o_439_), .Y(u2__abc_52155_new_n24351_));
OR2X2 OR2X2_5588 ( .A(u2__abc_52155_new_n24352_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24353_));
OR2X2 OR2X2_5589 ( .A(u2__abc_52155_new_n24357_), .B(u2__abc_52155_new_n24348_), .Y(u2__abc_52155_new_n24358_));
OR2X2 OR2X2_559 ( .A(u2__abc_52155_new_n3265_), .B(u2__abc_52155_new_n3267_), .Y(u2__abc_52155_new_n3268_));
OR2X2 OR2X2_5590 ( .A(u2__abc_52155_new_n24349_), .B(u2_o_440_), .Y(u2__abc_52155_new_n24361_));
OR2X2 OR2X2_5591 ( .A(u2__abc_52155_new_n24364_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24365_));
OR2X2 OR2X2_5592 ( .A(u2__abc_52155_new_n24369_), .B(u2__abc_52155_new_n24360_), .Y(u2__abc_52155_new_n24370_));
OR2X2 OR2X2_5593 ( .A(u2__abc_52155_new_n24362_), .B(u2_o_441_), .Y(u2__abc_52155_new_n24375_));
OR2X2 OR2X2_5594 ( .A(u2__abc_52155_new_n24376_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24377_));
OR2X2 OR2X2_5595 ( .A(u2__abc_52155_new_n24381_), .B(u2__abc_52155_new_n24372_), .Y(u2__abc_52155_new_n24382_));
OR2X2 OR2X2_5596 ( .A(u2__abc_52155_new_n24373_), .B(u2_o_442_), .Y(u2__abc_52155_new_n24385_));
OR2X2 OR2X2_5597 ( .A(u2__abc_52155_new_n24388_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24389_));
OR2X2 OR2X2_5598 ( .A(u2__abc_52155_new_n24393_), .B(u2__abc_52155_new_n24384_), .Y(u2__abc_52155_new_n24394_));
OR2X2 OR2X2_5599 ( .A(u2__abc_52155_new_n24386_), .B(u2_o_443_), .Y(u2__abc_52155_new_n24399_));
OR2X2 OR2X2_56 ( .A(_abc_73687_new_n753_), .B(\a[27] ), .Y(_abc_73687_new_n912_));
OR2X2 OR2X2_560 ( .A(u2__abc_52155_new_n3270_), .B(u2__abc_52155_new_n3272_), .Y(u2__abc_52155_new_n3273_));
OR2X2 OR2X2_5600 ( .A(u2__abc_52155_new_n24400_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24401_));
OR2X2 OR2X2_5601 ( .A(u2__abc_52155_new_n24405_), .B(u2__abc_52155_new_n24396_), .Y(u2__abc_52155_new_n24406_));
OR2X2 OR2X2_5602 ( .A(u2__abc_52155_new_n24397_), .B(u2_o_444_), .Y(u2__abc_52155_new_n24409_));
OR2X2 OR2X2_5603 ( .A(u2__abc_52155_new_n24412_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24413_));
OR2X2 OR2X2_5604 ( .A(u2__abc_52155_new_n24417_), .B(u2__abc_52155_new_n24408_), .Y(u2__abc_52155_new_n24418_));
OR2X2 OR2X2_5605 ( .A(u2__abc_52155_new_n24410_), .B(u2_o_445_), .Y(u2__abc_52155_new_n24423_));
OR2X2 OR2X2_5606 ( .A(u2__abc_52155_new_n24424_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24425_));
OR2X2 OR2X2_5607 ( .A(u2__abc_52155_new_n24429_), .B(u2__abc_52155_new_n24420_), .Y(u2__abc_52155_new_n24430_));
OR2X2 OR2X2_5608 ( .A(u2__abc_52155_new_n24421_), .B(u2_o_446_), .Y(u2__abc_52155_new_n24433_));
OR2X2 OR2X2_5609 ( .A(u2__abc_52155_new_n24436_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24437_));
OR2X2 OR2X2_561 ( .A(u2__abc_52155_new_n3268_), .B(u2__abc_52155_new_n3273_), .Y(u2__abc_52155_new_n3274_));
OR2X2 OR2X2_5610 ( .A(u2__abc_52155_new_n24441_), .B(u2__abc_52155_new_n24432_), .Y(u2__abc_52155_new_n24442_));
OR2X2 OR2X2_5611 ( .A(u2__abc_52155_new_n24434_), .B(u2_o_447_), .Y(u2__abc_52155_new_n24445_));
OR2X2 OR2X2_5612 ( .A(u2__abc_52155_new_n24448_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24449_));
OR2X2 OR2X2_5613 ( .A(u2__abc_52155_new_n24453_), .B(u2__abc_52155_new_n24444_), .Y(u2__abc_52155_new_n24454_));
OR2X2 OR2X2_5614 ( .A(u2__abc_52155_new_n24446_), .B(u2_o_448_), .Y(u2__abc_52155_new_n24457_));
OR2X2 OR2X2_5615 ( .A(u2__abc_52155_new_n24460_), .B(u2__abc_52155_new_n2974_), .Y(u2__abc_52155_new_n24461_));
OR2X2 OR2X2_5616 ( .A(u2__abc_52155_new_n24465_), .B(u2__abc_52155_new_n24456_), .Y(u2__abc_52155_new_n24466_));
OR2X2 OR2X2_562 ( .A(u2__abc_52155_new_n3263_), .B(u2__abc_52155_new_n3274_), .Y(u2__abc_52155_new_n3275_));
OR2X2 OR2X2_563 ( .A(u2__abc_52155_new_n3166_), .B(u2__abc_52155_new_n3279_), .Y(u2__abc_52155_new_n3280_));
OR2X2 OR2X2_564 ( .A(u2__abc_52155_new_n3242_), .B(u2__abc_52155_new_n3245_), .Y(u2__abc_52155_new_n3282_));
OR2X2 OR2X2_565 ( .A(u2__abc_52155_new_n3237_), .B(u2__abc_52155_new_n3283_), .Y(u2__abc_52155_new_n3284_));
OR2X2 OR2X2_566 ( .A(u2__abc_52155_new_n3286_), .B(u2__abc_52155_new_n3233_), .Y(u2__abc_52155_new_n3287_));
OR2X2 OR2X2_567 ( .A(u2__abc_52155_new_n3289_), .B(u2__abc_52155_new_n3275_), .Y(u2__abc_52155_new_n3290_));
OR2X2 OR2X2_568 ( .A(u2__abc_52155_new_n3292_), .B(u2__abc_52155_new_n3265_), .Y(u2__abc_52155_new_n3293_));
OR2X2 OR2X2_569 ( .A(u2__abc_52155_new_n3294_), .B(u2__abc_52155_new_n3263_), .Y(u2__abc_52155_new_n3295_));
OR2X2 OR2X2_57 ( .A(aNan), .B(sqrto_104_), .Y(_abc_73687_new_n914_));
OR2X2 OR2X2_570 ( .A(u2__abc_52155_new_n3297_), .B(u2__abc_52155_new_n3261_), .Y(u2__abc_52155_new_n3298_));
OR2X2 OR2X2_571 ( .A(u2__abc_52155_new_n3301_), .B(u2__abc_52155_new_n3281_), .Y(u2__abc_52155_new_n3302_));
OR2X2 OR2X2_572 ( .A(u2__abc_52155_new_n3191_), .B(u2__abc_52155_new_n3180_), .Y(u2__abc_52155_new_n3304_));
OR2X2 OR2X2_573 ( .A(u2__abc_52155_new_n3305_), .B(u2__abc_52155_new_n3177_), .Y(u2__abc_52155_new_n3306_));
OR2X2 OR2X2_574 ( .A(u2__abc_52155_new_n3308_), .B(u2__abc_52155_new_n3175_), .Y(u2__abc_52155_new_n3309_));
OR2X2 OR2X2_575 ( .A(u2__abc_52155_new_n3311_), .B(u2__abc_52155_new_n3303_), .Y(u2__abc_52155_new_n3312_));
OR2X2 OR2X2_576 ( .A(u2__abc_52155_new_n3313_), .B(u2__abc_52155_new_n3203_), .Y(u2__abc_52155_new_n3314_));
OR2X2 OR2X2_577 ( .A(u2__abc_52155_new_n3315_), .B(u2__abc_52155_new_n3214_), .Y(u2__abc_52155_new_n3316_));
OR2X2 OR2X2_578 ( .A(u2__abc_52155_new_n3317_), .B(u2__abc_52155_new_n3314_), .Y(u2__abc_52155_new_n3318_));
OR2X2 OR2X2_579 ( .A(u2__abc_52155_new_n3387_), .B(u2__abc_52155_new_n3389_), .Y(u2__abc_52155_new_n3390_));
OR2X2 OR2X2_58 ( .A(_abc_73687_new_n753_), .B(\a[28] ), .Y(_abc_73687_new_n915_));
OR2X2 OR2X2_580 ( .A(u2__abc_52155_new_n3392_), .B(u2__abc_52155_new_n3394_), .Y(u2__abc_52155_new_n3395_));
OR2X2 OR2X2_581 ( .A(u2__abc_52155_new_n3390_), .B(u2__abc_52155_new_n3395_), .Y(u2__abc_52155_new_n3396_));
OR2X2 OR2X2_582 ( .A(u2__abc_52155_new_n3448_), .B(u2__abc_52155_new_n3450_), .Y(u2__abc_52155_new_n3451_));
OR2X2 OR2X2_583 ( .A(u2__abc_52155_new_n3453_), .B(u2__abc_52155_new_n3455_), .Y(u2__abc_52155_new_n3456_));
OR2X2 OR2X2_584 ( .A(u2__abc_52155_new_n3451_), .B(u2__abc_52155_new_n3456_), .Y(u2__abc_52155_new_n3457_));
OR2X2 OR2X2_585 ( .A(u2__abc_52155_new_n3508_), .B(u2__abc_52155_new_n3510_), .Y(u2__abc_52155_new_n3511_));
OR2X2 OR2X2_586 ( .A(u2__abc_52155_new_n3513_), .B(u2__abc_52155_new_n3515_), .Y(u2__abc_52155_new_n3516_));
OR2X2 OR2X2_587 ( .A(u2__abc_52155_new_n3511_), .B(u2__abc_52155_new_n3516_), .Y(u2__abc_52155_new_n3517_));
OR2X2 OR2X2_588 ( .A(u2__abc_52155_new_n3519_), .B(u2_remHi_30_), .Y(u2__abc_52155_new_n3522_));
OR2X2 OR2X2_589 ( .A(u2__abc_52155_new_n3534_), .B(u2__abc_52155_new_n3536_), .Y(u2__abc_52155_new_n3537_));
OR2X2 OR2X2_59 ( .A(aNan), .B(sqrto_105_), .Y(_abc_73687_new_n917_));
OR2X2 OR2X2_590 ( .A(u2__abc_52155_new_n3539_), .B(u2__abc_52155_new_n3541_), .Y(u2__abc_52155_new_n3542_));
OR2X2 OR2X2_591 ( .A(u2__abc_52155_new_n3537_), .B(u2__abc_52155_new_n3542_), .Y(u2__abc_52155_new_n3543_));
OR2X2 OR2X2_592 ( .A(u2__abc_52155_new_n3545_), .B(u2__abc_52155_new_n3547_), .Y(u2__abc_52155_new_n3548_));
OR2X2 OR2X2_593 ( .A(u2__abc_52155_new_n3550_), .B(u2__abc_52155_new_n3552_), .Y(u2__abc_52155_new_n3553_));
OR2X2 OR2X2_594 ( .A(u2__abc_52155_new_n3548_), .B(u2__abc_52155_new_n3553_), .Y(u2__abc_52155_new_n3554_));
OR2X2 OR2X2_595 ( .A(u2__abc_52155_new_n3543_), .B(u2__abc_52155_new_n3554_), .Y(u2__abc_52155_new_n3555_));
OR2X2 OR2X2_596 ( .A(u2__abc_52155_new_n3322_), .B(u2__abc_52155_new_n3560_), .Y(u2__abc_52155_new_n3561_));
OR2X2 OR2X2_597 ( .A(u2__abc_52155_new_n3522_), .B(u2__abc_52155_new_n3525_), .Y(u2__abc_52155_new_n3564_));
OR2X2 OR2X2_598 ( .A(u2__abc_52155_new_n3517_), .B(u2__abc_52155_new_n3565_), .Y(u2__abc_52155_new_n3566_));
OR2X2 OR2X2_599 ( .A(u2__abc_52155_new_n3568_), .B(u2__abc_52155_new_n3513_), .Y(u2__abc_52155_new_n3569_));
OR2X2 OR2X2_6 ( .A(_abc_73687_new_n753_), .B(\a[2] ), .Y(_abc_73687_new_n837_));
OR2X2 OR2X2_60 ( .A(_abc_73687_new_n753_), .B(\a[29] ), .Y(_abc_73687_new_n918_));
OR2X2 OR2X2_600 ( .A(u2__abc_52155_new_n3571_), .B(u2__abc_52155_new_n3555_), .Y(u2__abc_52155_new_n3572_));
OR2X2 OR2X2_601 ( .A(u2__abc_52155_new_n3574_), .B(u2__abc_52155_new_n3545_), .Y(u2__abc_52155_new_n3575_));
OR2X2 OR2X2_602 ( .A(u2__abc_52155_new_n3576_), .B(u2__abc_52155_new_n3543_), .Y(u2__abc_52155_new_n3577_));
OR2X2 OR2X2_603 ( .A(u2__abc_52155_new_n3579_), .B(u2__abc_52155_new_n3541_), .Y(u2__abc_52155_new_n3580_));
OR2X2 OR2X2_604 ( .A(u2__abc_52155_new_n3583_), .B(u2__abc_52155_new_n3563_), .Y(u2__abc_52155_new_n3584_));
OR2X2 OR2X2_605 ( .A(u2__abc_52155_new_n3464_), .B(u2__abc_52155_new_n3467_), .Y(u2__abc_52155_new_n3586_));
OR2X2 OR2X2_606 ( .A(u2__abc_52155_new_n3587_), .B(u2__abc_52155_new_n3457_), .Y(u2__abc_52155_new_n3588_));
OR2X2 OR2X2_607 ( .A(u2__abc_52155_new_n3590_), .B(u2__abc_52155_new_n3455_), .Y(u2__abc_52155_new_n3591_));
OR2X2 OR2X2_608 ( .A(u2__abc_52155_new_n3593_), .B(u2__abc_52155_new_n3585_), .Y(u2__abc_52155_new_n3594_));
OR2X2 OR2X2_609 ( .A(u2__abc_52155_new_n3595_), .B(u2__abc_52155_new_n3494_), .Y(u2__abc_52155_new_n3596_));
OR2X2 OR2X2_61 ( .A(aNan), .B(sqrto_106_), .Y(_abc_73687_new_n920_));
OR2X2 OR2X2_610 ( .A(u2__abc_52155_new_n3598_), .B(u2__abc_52155_new_n3486_), .Y(u2__abc_52155_new_n3599_));
OR2X2 OR2X2_611 ( .A(u2__abc_52155_new_n3597_), .B(u2__abc_52155_new_n3599_), .Y(u2__abc_52155_new_n3600_));
OR2X2 OR2X2_612 ( .A(u2__abc_52155_new_n3603_), .B(u2__abc_52155_new_n3562_), .Y(u2__abc_52155_new_n3604_));
OR2X2 OR2X2_613 ( .A(u2__abc_52155_new_n3410_), .B(u2__abc_52155_new_n3399_), .Y(u2__abc_52155_new_n3607_));
OR2X2 OR2X2_614 ( .A(u2__abc_52155_new_n3608_), .B(u2__abc_52155_new_n3396_), .Y(u2__abc_52155_new_n3609_));
OR2X2 OR2X2_615 ( .A(u2__abc_52155_new_n3611_), .B(u2__abc_52155_new_n3394_), .Y(u2__abc_52155_new_n3612_));
OR2X2 OR2X2_616 ( .A(u2__abc_52155_new_n3614_), .B(u2__abc_52155_new_n3606_), .Y(u2__abc_52155_new_n3615_));
OR2X2 OR2X2_617 ( .A(u2__abc_52155_new_n3616_), .B(u2__abc_52155_new_n3433_), .Y(u2__abc_52155_new_n3617_));
OR2X2 OR2X2_618 ( .A(u2__abc_52155_new_n3619_), .B(u2__abc_52155_new_n3425_), .Y(u2__abc_52155_new_n3620_));
OR2X2 OR2X2_619 ( .A(u2__abc_52155_new_n3618_), .B(u2__abc_52155_new_n3620_), .Y(u2__abc_52155_new_n3621_));
OR2X2 OR2X2_62 ( .A(_abc_73687_new_n753_), .B(\a[30] ), .Y(_abc_73687_new_n921_));
OR2X2 OR2X2_620 ( .A(u2__abc_52155_new_n3623_), .B(u2__abc_52155_new_n3605_), .Y(u2__abc_52155_new_n3624_));
OR2X2 OR2X2_621 ( .A(u2__abc_52155_new_n3625_), .B(u2__abc_52155_new_n3349_), .Y(u2__abc_52155_new_n3626_));
OR2X2 OR2X2_622 ( .A(u2__abc_52155_new_n3628_), .B(u2__abc_52155_new_n3334_), .Y(u2__abc_52155_new_n3629_));
OR2X2 OR2X2_623 ( .A(u2__abc_52155_new_n3627_), .B(u2__abc_52155_new_n3629_), .Y(u2__abc_52155_new_n3630_));
OR2X2 OR2X2_624 ( .A(u2__abc_52155_new_n3632_), .B(u2__abc_52155_new_n3373_), .Y(u2__abc_52155_new_n3633_));
OR2X2 OR2X2_625 ( .A(u2__abc_52155_new_n3635_), .B(u2__abc_52155_new_n3362_), .Y(u2__abc_52155_new_n3636_));
OR2X2 OR2X2_626 ( .A(u2__abc_52155_new_n3634_), .B(u2__abc_52155_new_n3636_), .Y(u2__abc_52155_new_n3637_));
OR2X2 OR2X2_627 ( .A(u2__abc_52155_new_n3631_), .B(u2__abc_52155_new_n3637_), .Y(u2__abc_52155_new_n3638_));
OR2X2 OR2X2_628 ( .A(u2__abc_52155_new_n3834_), .B(u2__abc_52155_new_n3836_), .Y(u2__abc_52155_new_n3837_));
OR2X2 OR2X2_629 ( .A(u2__abc_52155_new_n3839_), .B(u2__abc_52155_new_n3841_), .Y(u2__abc_52155_new_n3842_));
OR2X2 OR2X2_63 ( .A(aNan), .B(sqrto_107_), .Y(_abc_73687_new_n923_));
OR2X2 OR2X2_630 ( .A(u2__abc_52155_new_n3837_), .B(u2__abc_52155_new_n3842_), .Y(u2__abc_52155_new_n3843_));
OR2X2 OR2X2_631 ( .A(u2__abc_52155_new_n3974_), .B(u2__abc_52155_new_n3976_), .Y(u2__abc_52155_new_n3977_));
OR2X2 OR2X2_632 ( .A(u2__abc_52155_new_n3979_), .B(u2__abc_52155_new_n3981_), .Y(u2__abc_52155_new_n3982_));
OR2X2 OR2X2_633 ( .A(u2__abc_52155_new_n3977_), .B(u2__abc_52155_new_n3982_), .Y(u2__abc_52155_new_n3983_));
OR2X2 OR2X2_634 ( .A(u2__abc_52155_new_n4035_), .B(u2__abc_52155_new_n4037_), .Y(u2__abc_52155_new_n4038_));
OR2X2 OR2X2_635 ( .A(u2__abc_52155_new_n4040_), .B(u2__abc_52155_new_n4042_), .Y(u2__abc_52155_new_n4043_));
OR2X2 OR2X2_636 ( .A(u2__abc_52155_new_n4038_), .B(u2__abc_52155_new_n4043_), .Y(u2__abc_52155_new_n4044_));
OR2X2 OR2X2_637 ( .A(u2__abc_52155_new_n4079_), .B(u2_remHi_62_), .Y(u2__abc_52155_new_n4082_));
OR2X2 OR2X2_638 ( .A(u2__abc_52155_new_n4093_), .B(u2__abc_52155_new_n4095_), .Y(u2__abc_52155_new_n4096_));
OR2X2 OR2X2_639 ( .A(u2__abc_52155_new_n4098_), .B(u2__abc_52155_new_n4100_), .Y(u2__abc_52155_new_n4101_));
OR2X2 OR2X2_64 ( .A(_abc_73687_new_n753_), .B(\a[31] ), .Y(_abc_73687_new_n924_));
OR2X2 OR2X2_640 ( .A(u2__abc_52155_new_n4096_), .B(u2__abc_52155_new_n4101_), .Y(u2__abc_52155_new_n4102_));
OR2X2 OR2X2_641 ( .A(u2__abc_52155_new_n4106_), .B(u2__abc_52155_new_n4108_), .Y(u2__abc_52155_new_n4109_));
OR2X2 OR2X2_642 ( .A(u2__abc_52155_new_n4111_), .B(u2__abc_52155_new_n4113_), .Y(u2__abc_52155_new_n4114_));
OR2X2 OR2X2_643 ( .A(u2__abc_52155_new_n4109_), .B(u2__abc_52155_new_n4114_), .Y(u2__abc_52155_new_n4115_));
OR2X2 OR2X2_644 ( .A(u2__abc_52155_new_n4117_), .B(u2__abc_52155_new_n4119_), .Y(u2__abc_52155_new_n4120_));
OR2X2 OR2X2_645 ( .A(u2__abc_52155_new_n4122_), .B(u2__abc_52155_new_n4124_), .Y(u2__abc_52155_new_n4125_));
OR2X2 OR2X2_646 ( .A(u2__abc_52155_new_n4120_), .B(u2__abc_52155_new_n4125_), .Y(u2__abc_52155_new_n4126_));
OR2X2 OR2X2_647 ( .A(u2__abc_52155_new_n4115_), .B(u2__abc_52155_new_n4126_), .Y(u2__abc_52155_new_n4127_));
OR2X2 OR2X2_648 ( .A(u2__abc_52155_new_n3642_), .B(u2__abc_52155_new_n4133_), .Y(u2__abc_52155_new_n4134_));
OR2X2 OR2X2_649 ( .A(u2__abc_52155_new_n4082_), .B(u2__abc_52155_new_n4085_), .Y(u2__abc_52155_new_n4138_));
OR2X2 OR2X2_65 ( .A(aNan), .B(sqrto_108_), .Y(_abc_73687_new_n926_));
OR2X2 OR2X2_650 ( .A(u2__abc_52155_new_n4102_), .B(u2__abc_52155_new_n4139_), .Y(u2__abc_52155_new_n4140_));
OR2X2 OR2X2_651 ( .A(u2__abc_52155_new_n4142_), .B(u2__abc_52155_new_n4098_), .Y(u2__abc_52155_new_n4143_));
OR2X2 OR2X2_652 ( .A(u2__abc_52155_new_n4145_), .B(u2__abc_52155_new_n4127_), .Y(u2__abc_52155_new_n4146_));
OR2X2 OR2X2_653 ( .A(u2__abc_52155_new_n4148_), .B(u2__abc_52155_new_n4117_), .Y(u2__abc_52155_new_n4149_));
OR2X2 OR2X2_654 ( .A(u2__abc_52155_new_n4150_), .B(u2__abc_52155_new_n4115_), .Y(u2__abc_52155_new_n4151_));
OR2X2 OR2X2_655 ( .A(u2__abc_52155_new_n4153_), .B(u2__abc_52155_new_n4113_), .Y(u2__abc_52155_new_n4154_));
OR2X2 OR2X2_656 ( .A(u2__abc_52155_new_n4157_), .B(u2__abc_52155_new_n4137_), .Y(u2__abc_52155_new_n4158_));
OR2X2 OR2X2_657 ( .A(u2__abc_52155_new_n4024_), .B(u2__abc_52155_new_n4027_), .Y(u2__abc_52155_new_n4160_));
OR2X2 OR2X2_658 ( .A(u2__abc_52155_new_n4161_), .B(u2__abc_52155_new_n4044_), .Y(u2__abc_52155_new_n4162_));
OR2X2 OR2X2_659 ( .A(u2__abc_52155_new_n4164_), .B(u2__abc_52155_new_n4042_), .Y(u2__abc_52155_new_n4165_));
OR2X2 OR2X2_66 ( .A(_abc_73687_new_n753_), .B(\a[32] ), .Y(_abc_73687_new_n927_));
OR2X2 OR2X2_660 ( .A(u2__abc_52155_new_n4167_), .B(u2__abc_52155_new_n4159_), .Y(u2__abc_52155_new_n4168_));
OR2X2 OR2X2_661 ( .A(u2__abc_52155_new_n4169_), .B(u2__abc_52155_new_n4066_), .Y(u2__abc_52155_new_n4170_));
OR2X2 OR2X2_662 ( .A(u2__abc_52155_new_n4172_), .B(u2__abc_52155_new_n4058_), .Y(u2__abc_52155_new_n4173_));
OR2X2 OR2X2_663 ( .A(u2__abc_52155_new_n4171_), .B(u2__abc_52155_new_n4173_), .Y(u2__abc_52155_new_n4174_));
OR2X2 OR2X2_664 ( .A(u2__abc_52155_new_n4177_), .B(u2__abc_52155_new_n4136_), .Y(u2__abc_52155_new_n4178_));
OR2X2 OR2X2_665 ( .A(u2__abc_52155_new_n3963_), .B(u2__abc_52155_new_n3966_), .Y(u2__abc_52155_new_n4181_));
OR2X2 OR2X2_666 ( .A(u2__abc_52155_new_n4182_), .B(u2__abc_52155_new_n3983_), .Y(u2__abc_52155_new_n4183_));
OR2X2 OR2X2_667 ( .A(u2__abc_52155_new_n4185_), .B(u2__abc_52155_new_n3981_), .Y(u2__abc_52155_new_n4186_));
OR2X2 OR2X2_668 ( .A(u2__abc_52155_new_n4188_), .B(u2__abc_52155_new_n4180_), .Y(u2__abc_52155_new_n4189_));
OR2X2 OR2X2_669 ( .A(u2__abc_52155_new_n4190_), .B(u2__abc_52155_new_n4005_), .Y(u2__abc_52155_new_n4191_));
OR2X2 OR2X2_67 ( .A(aNan), .B(sqrto_109_), .Y(_abc_73687_new_n929_));
OR2X2 OR2X2_670 ( .A(u2__abc_52155_new_n4193_), .B(u2__abc_52155_new_n3997_), .Y(u2__abc_52155_new_n4194_));
OR2X2 OR2X2_671 ( .A(u2__abc_52155_new_n4192_), .B(u2__abc_52155_new_n4194_), .Y(u2__abc_52155_new_n4195_));
OR2X2 OR2X2_672 ( .A(u2__abc_52155_new_n4197_), .B(u2__abc_52155_new_n4179_), .Y(u2__abc_52155_new_n4198_));
OR2X2 OR2X2_673 ( .A(u2__abc_52155_new_n4199_), .B(u2__abc_52155_new_n3945_), .Y(u2__abc_52155_new_n4200_));
OR2X2 OR2X2_674 ( .A(u2__abc_52155_new_n4202_), .B(u2__abc_52155_new_n3937_), .Y(u2__abc_52155_new_n4203_));
OR2X2 OR2X2_675 ( .A(u2__abc_52155_new_n4201_), .B(u2__abc_52155_new_n4203_), .Y(u2__abc_52155_new_n4204_));
OR2X2 OR2X2_676 ( .A(u2__abc_52155_new_n4206_), .B(u2__abc_52155_new_n3914_), .Y(u2__abc_52155_new_n4207_));
OR2X2 OR2X2_677 ( .A(u2__abc_52155_new_n4209_), .B(u2__abc_52155_new_n3906_), .Y(u2__abc_52155_new_n4210_));
OR2X2 OR2X2_678 ( .A(u2__abc_52155_new_n4208_), .B(u2__abc_52155_new_n4210_), .Y(u2__abc_52155_new_n4211_));
OR2X2 OR2X2_679 ( .A(u2__abc_52155_new_n4205_), .B(u2__abc_52155_new_n4211_), .Y(u2__abc_52155_new_n4212_));
OR2X2 OR2X2_68 ( .A(_abc_73687_new_n753_), .B(\a[33] ), .Y(_abc_73687_new_n930_));
OR2X2 OR2X2_680 ( .A(u2__abc_52155_new_n4215_), .B(u2__abc_52155_new_n4135_), .Y(u2__abc_52155_new_n4216_));
OR2X2 OR2X2_681 ( .A(u2__abc_52155_new_n3857_), .B(u2__abc_52155_new_n3846_), .Y(u2__abc_52155_new_n4220_));
OR2X2 OR2X2_682 ( .A(u2__abc_52155_new_n4221_), .B(u2__abc_52155_new_n3843_), .Y(u2__abc_52155_new_n4222_));
OR2X2 OR2X2_683 ( .A(u2__abc_52155_new_n4224_), .B(u2__abc_52155_new_n3841_), .Y(u2__abc_52155_new_n4225_));
OR2X2 OR2X2_684 ( .A(u2__abc_52155_new_n4227_), .B(u2__abc_52155_new_n4219_), .Y(u2__abc_52155_new_n4228_));
OR2X2 OR2X2_685 ( .A(u2__abc_52155_new_n4229_), .B(u2__abc_52155_new_n3880_), .Y(u2__abc_52155_new_n4230_));
OR2X2 OR2X2_686 ( .A(u2__abc_52155_new_n4232_), .B(u2__abc_52155_new_n3872_), .Y(u2__abc_52155_new_n4233_));
OR2X2 OR2X2_687 ( .A(u2__abc_52155_new_n4231_), .B(u2__abc_52155_new_n4233_), .Y(u2__abc_52155_new_n4234_));
OR2X2 OR2X2_688 ( .A(u2__abc_52155_new_n4236_), .B(u2__abc_52155_new_n4218_), .Y(u2__abc_52155_new_n4237_));
OR2X2 OR2X2_689 ( .A(u2__abc_52155_new_n4238_), .B(u2__abc_52155_new_n3789_), .Y(u2__abc_52155_new_n4239_));
OR2X2 OR2X2_69 ( .A(aNan), .B(sqrto_110_), .Y(_abc_73687_new_n932_));
OR2X2 OR2X2_690 ( .A(u2__abc_52155_new_n4241_), .B(u2__abc_52155_new_n3781_), .Y(u2__abc_52155_new_n4242_));
OR2X2 OR2X2_691 ( .A(u2__abc_52155_new_n4240_), .B(u2__abc_52155_new_n4242_), .Y(u2__abc_52155_new_n4243_));
OR2X2 OR2X2_692 ( .A(u2__abc_52155_new_n4245_), .B(u2__abc_52155_new_n3820_), .Y(u2__abc_52155_new_n4246_));
OR2X2 OR2X2_693 ( .A(u2__abc_52155_new_n4248_), .B(u2__abc_52155_new_n3812_), .Y(u2__abc_52155_new_n4249_));
OR2X2 OR2X2_694 ( .A(u2__abc_52155_new_n4247_), .B(u2__abc_52155_new_n4249_), .Y(u2__abc_52155_new_n4250_));
OR2X2 OR2X2_695 ( .A(u2__abc_52155_new_n4244_), .B(u2__abc_52155_new_n4250_), .Y(u2__abc_52155_new_n4251_));
OR2X2 OR2X2_696 ( .A(u2__abc_52155_new_n4253_), .B(u2__abc_52155_new_n4217_), .Y(u2__abc_52155_new_n4254_));
OR2X2 OR2X2_697 ( .A(u2__abc_52155_new_n4255_), .B(u2__abc_52155_new_n3654_), .Y(u2__abc_52155_new_n4256_));
OR2X2 OR2X2_698 ( .A(u2__abc_52155_new_n4258_), .B(u2__abc_52155_new_n3669_), .Y(u2__abc_52155_new_n4259_));
OR2X2 OR2X2_699 ( .A(u2__abc_52155_new_n4257_), .B(u2__abc_52155_new_n4259_), .Y(u2__abc_52155_new_n4260_));
OR2X2 OR2X2_7 ( .A(aNan), .B(sqrto_79_), .Y(_abc_73687_new_n839_));
OR2X2 OR2X2_70 ( .A(_abc_73687_new_n753_), .B(\a[34] ), .Y(_abc_73687_new_n933_));
OR2X2 OR2X2_700 ( .A(u2__abc_52155_new_n4262_), .B(u2__abc_52155_new_n3682_), .Y(u2__abc_52155_new_n4263_));
OR2X2 OR2X2_701 ( .A(u2__abc_52155_new_n4264_), .B(u2__abc_52155_new_n3693_), .Y(u2__abc_52155_new_n4265_));
OR2X2 OR2X2_702 ( .A(u2__abc_52155_new_n4266_), .B(u2__abc_52155_new_n4263_), .Y(u2__abc_52155_new_n4267_));
OR2X2 OR2X2_703 ( .A(u2__abc_52155_new_n4261_), .B(u2__abc_52155_new_n4267_), .Y(u2__abc_52155_new_n4268_));
OR2X2 OR2X2_704 ( .A(u2__abc_52155_new_n4269_), .B(u2__abc_52155_new_n3717_), .Y(u2__abc_52155_new_n4270_));
OR2X2 OR2X2_705 ( .A(u2__abc_52155_new_n4272_), .B(u2__abc_52155_new_n3732_), .Y(u2__abc_52155_new_n4273_));
OR2X2 OR2X2_706 ( .A(u2__abc_52155_new_n4271_), .B(u2__abc_52155_new_n4273_), .Y(u2__abc_52155_new_n4274_));
OR2X2 OR2X2_707 ( .A(u2__abc_52155_new_n4276_), .B(u2__abc_52155_new_n3748_), .Y(u2__abc_52155_new_n4277_));
OR2X2 OR2X2_708 ( .A(u2__abc_52155_new_n4278_), .B(u2__abc_52155_new_n3756_), .Y(u2__abc_52155_new_n4279_));
OR2X2 OR2X2_709 ( .A(u2__abc_52155_new_n4280_), .B(u2__abc_52155_new_n4277_), .Y(u2__abc_52155_new_n4281_));
OR2X2 OR2X2_71 ( .A(aNan), .B(sqrto_111_), .Y(_abc_73687_new_n935_));
OR2X2 OR2X2_710 ( .A(u2__abc_52155_new_n4275_), .B(u2__abc_52155_new_n4281_), .Y(u2__abc_52155_new_n4282_));
OR2X2 OR2X2_711 ( .A(u2__abc_52155_new_n4283_), .B(u2__abc_52155_new_n4268_), .Y(u2__abc_52155_new_n4284_));
OR2X2 OR2X2_712 ( .A(u2__abc_52155_new_n4766_), .B(u2__abc_52155_new_n4768_), .Y(u2__abc_52155_new_n4769_));
OR2X2 OR2X2_713 ( .A(u2__abc_52155_new_n4771_), .B(u2__abc_52155_new_n4773_), .Y(u2__abc_52155_new_n4774_));
OR2X2 OR2X2_714 ( .A(u2__abc_52155_new_n4769_), .B(u2__abc_52155_new_n4774_), .Y(u2__abc_52155_new_n4775_));
OR2X2 OR2X2_715 ( .A(u2__abc_52155_new_n4988_), .B(u2__abc_52155_new_n4990_), .Y(u2__abc_52155_new_n4991_));
OR2X2 OR2X2_716 ( .A(u2__abc_52155_new_n4993_), .B(u2__abc_52155_new_n4995_), .Y(u2__abc_52155_new_n4996_));
OR2X2 OR2X2_717 ( .A(u2__abc_52155_new_n4991_), .B(u2__abc_52155_new_n4996_), .Y(u2__abc_52155_new_n4997_));
OR2X2 OR2X2_718 ( .A(u2__abc_52155_new_n5144_), .B(u2__abc_52155_new_n5146_), .Y(u2__abc_52155_new_n5147_));
OR2X2 OR2X2_719 ( .A(u2__abc_52155_new_n5149_), .B(u2__abc_52155_new_n5151_), .Y(u2__abc_52155_new_n5152_));
OR2X2 OR2X2_72 ( .A(_abc_73687_new_n753_), .B(\a[35] ), .Y(_abc_73687_new_n936_));
OR2X2 OR2X2_720 ( .A(u2__abc_52155_new_n5147_), .B(u2__abc_52155_new_n5152_), .Y(u2__abc_52155_new_n5153_));
OR2X2 OR2X2_721 ( .A(u2__abc_52155_new_n5174_), .B(u2__abc_52155_new_n5176_), .Y(u2__abc_52155_new_n5177_));
OR2X2 OR2X2_722 ( .A(u2__abc_52155_new_n5179_), .B(u2__abc_52155_new_n5181_), .Y(u2__abc_52155_new_n5182_));
OR2X2 OR2X2_723 ( .A(u2__abc_52155_new_n5177_), .B(u2__abc_52155_new_n5182_), .Y(u2__abc_52155_new_n5183_));
OR2X2 OR2X2_724 ( .A(u2__abc_52155_new_n5233_), .B(u2_remHi_126_), .Y(u2__abc_52155_new_n5236_));
OR2X2 OR2X2_725 ( .A(u2__abc_52155_new_n5247_), .B(u2__abc_52155_new_n5249_), .Y(u2__abc_52155_new_n5250_));
OR2X2 OR2X2_726 ( .A(u2__abc_52155_new_n5252_), .B(u2__abc_52155_new_n5254_), .Y(u2__abc_52155_new_n5255_));
OR2X2 OR2X2_727 ( .A(u2__abc_52155_new_n5250_), .B(u2__abc_52155_new_n5255_), .Y(u2__abc_52155_new_n5256_));
OR2X2 OR2X2_728 ( .A(u2__abc_52155_new_n5260_), .B(u2__abc_52155_new_n5262_), .Y(u2__abc_52155_new_n5263_));
OR2X2 OR2X2_729 ( .A(u2__abc_52155_new_n5265_), .B(u2__abc_52155_new_n5267_), .Y(u2__abc_52155_new_n5268_));
OR2X2 OR2X2_73 ( .A(aNan), .B(sqrto_112_), .Y(_abc_73687_new_n938_));
OR2X2 OR2X2_730 ( .A(u2__abc_52155_new_n5263_), .B(u2__abc_52155_new_n5268_), .Y(u2__abc_52155_new_n5269_));
OR2X2 OR2X2_731 ( .A(u2__abc_52155_new_n5271_), .B(u2__abc_52155_new_n5273_), .Y(u2__abc_52155_new_n5274_));
OR2X2 OR2X2_732 ( .A(u2__abc_52155_new_n5276_), .B(u2__abc_52155_new_n5278_), .Y(u2__abc_52155_new_n5279_));
OR2X2 OR2X2_733 ( .A(u2__abc_52155_new_n5274_), .B(u2__abc_52155_new_n5279_), .Y(u2__abc_52155_new_n5280_));
OR2X2 OR2X2_734 ( .A(u2__abc_52155_new_n5269_), .B(u2__abc_52155_new_n5280_), .Y(u2__abc_52155_new_n5281_));
OR2X2 OR2X2_735 ( .A(u2__abc_52155_new_n4288_), .B(u2__abc_52155_new_n5288_), .Y(u2__abc_52155_new_n5289_));
OR2X2 OR2X2_736 ( .A(u2__abc_52155_new_n5236_), .B(u2__abc_52155_new_n5239_), .Y(u2__abc_52155_new_n5294_));
OR2X2 OR2X2_737 ( .A(u2__abc_52155_new_n5256_), .B(u2__abc_52155_new_n5295_), .Y(u2__abc_52155_new_n5296_));
OR2X2 OR2X2_738 ( .A(u2__abc_52155_new_n5298_), .B(u2__abc_52155_new_n5252_), .Y(u2__abc_52155_new_n5299_));
OR2X2 OR2X2_739 ( .A(u2__abc_52155_new_n5301_), .B(u2__abc_52155_new_n5281_), .Y(u2__abc_52155_new_n5302_));
OR2X2 OR2X2_74 ( .A(_abc_73687_new_n753_), .B(\a[36] ), .Y(_abc_73687_new_n939_));
OR2X2 OR2X2_740 ( .A(u2__abc_52155_new_n5304_), .B(u2__abc_52155_new_n5271_), .Y(u2__abc_52155_new_n5305_));
OR2X2 OR2X2_741 ( .A(u2__abc_52155_new_n5306_), .B(u2__abc_52155_new_n5269_), .Y(u2__abc_52155_new_n5307_));
OR2X2 OR2X2_742 ( .A(u2__abc_52155_new_n5309_), .B(u2__abc_52155_new_n5267_), .Y(u2__abc_52155_new_n5310_));
OR2X2 OR2X2_743 ( .A(u2__abc_52155_new_n5313_), .B(u2__abc_52155_new_n5293_), .Y(u2__abc_52155_new_n5314_));
OR2X2 OR2X2_744 ( .A(u2__abc_52155_new_n5190_), .B(u2__abc_52155_new_n5193_), .Y(u2__abc_52155_new_n5316_));
OR2X2 OR2X2_745 ( .A(u2__abc_52155_new_n5317_), .B(u2__abc_52155_new_n5183_), .Y(u2__abc_52155_new_n5318_));
OR2X2 OR2X2_746 ( .A(u2__abc_52155_new_n5320_), .B(u2__abc_52155_new_n5181_), .Y(u2__abc_52155_new_n5321_));
OR2X2 OR2X2_747 ( .A(u2__abc_52155_new_n5323_), .B(u2__abc_52155_new_n5315_), .Y(u2__abc_52155_new_n5324_));
OR2X2 OR2X2_748 ( .A(u2__abc_52155_new_n5325_), .B(u2__abc_52155_new_n5220_), .Y(u2__abc_52155_new_n5326_));
OR2X2 OR2X2_749 ( .A(u2__abc_52155_new_n5328_), .B(u2__abc_52155_new_n5212_), .Y(u2__abc_52155_new_n5329_));
OR2X2 OR2X2_75 ( .A(aNan), .B(sqrto_113_), .Y(_abc_73687_new_n941_));
OR2X2 OR2X2_750 ( .A(u2__abc_52155_new_n5327_), .B(u2__abc_52155_new_n5329_), .Y(u2__abc_52155_new_n5330_));
OR2X2 OR2X2_751 ( .A(u2__abc_52155_new_n5333_), .B(u2__abc_52155_new_n5292_), .Y(u2__abc_52155_new_n5334_));
OR2X2 OR2X2_752 ( .A(u2__abc_52155_new_n5167_), .B(u2__abc_52155_new_n5156_), .Y(u2__abc_52155_new_n5337_));
OR2X2 OR2X2_753 ( .A(u2__abc_52155_new_n5338_), .B(u2__abc_52155_new_n5153_), .Y(u2__abc_52155_new_n5339_));
OR2X2 OR2X2_754 ( .A(u2__abc_52155_new_n5341_), .B(u2__abc_52155_new_n5151_), .Y(u2__abc_52155_new_n5342_));
OR2X2 OR2X2_755 ( .A(u2__abc_52155_new_n5344_), .B(u2__abc_52155_new_n5336_), .Y(u2__abc_52155_new_n5345_));
OR2X2 OR2X2_756 ( .A(u2__abc_52155_new_n5346_), .B(u2__abc_52155_new_n5131_), .Y(u2__abc_52155_new_n5347_));
OR2X2 OR2X2_757 ( .A(u2__abc_52155_new_n5349_), .B(u2__abc_52155_new_n5123_), .Y(u2__abc_52155_new_n5350_));
OR2X2 OR2X2_758 ( .A(u2__abc_52155_new_n5348_), .B(u2__abc_52155_new_n5350_), .Y(u2__abc_52155_new_n5351_));
OR2X2 OR2X2_759 ( .A(u2__abc_52155_new_n5353_), .B(u2__abc_52155_new_n5335_), .Y(u2__abc_52155_new_n5354_));
OR2X2 OR2X2_76 ( .A(_abc_73687_new_n753_), .B(\a[37] ), .Y(_abc_73687_new_n942_));
OR2X2 OR2X2_760 ( .A(u2__abc_52155_new_n5355_), .B(u2__abc_52155_new_n5068_), .Y(u2__abc_52155_new_n5356_));
OR2X2 OR2X2_761 ( .A(u2__abc_52155_new_n5358_), .B(u2__abc_52155_new_n5060_), .Y(u2__abc_52155_new_n5359_));
OR2X2 OR2X2_762 ( .A(u2__abc_52155_new_n5357_), .B(u2__abc_52155_new_n5359_), .Y(u2__abc_52155_new_n5360_));
OR2X2 OR2X2_763 ( .A(u2__abc_52155_new_n5362_), .B(u2__abc_52155_new_n5099_), .Y(u2__abc_52155_new_n5363_));
OR2X2 OR2X2_764 ( .A(u2__abc_52155_new_n5365_), .B(u2__abc_52155_new_n5091_), .Y(u2__abc_52155_new_n5366_));
OR2X2 OR2X2_765 ( .A(u2__abc_52155_new_n5364_), .B(u2__abc_52155_new_n5366_), .Y(u2__abc_52155_new_n5367_));
OR2X2 OR2X2_766 ( .A(u2__abc_52155_new_n5361_), .B(u2__abc_52155_new_n5367_), .Y(u2__abc_52155_new_n5368_));
OR2X2 OR2X2_767 ( .A(u2__abc_52155_new_n5371_), .B(u2__abc_52155_new_n5291_), .Y(u2__abc_52155_new_n5372_));
OR2X2 OR2X2_768 ( .A(u2__abc_52155_new_n5011_), .B(u2__abc_52155_new_n5000_), .Y(u2__abc_52155_new_n5376_));
OR2X2 OR2X2_769 ( .A(u2__abc_52155_new_n5377_), .B(u2__abc_52155_new_n4997_), .Y(u2__abc_52155_new_n5378_));
OR2X2 OR2X2_77 ( .A(aNan), .B(sqrto_114_), .Y(_abc_73687_new_n944_));
OR2X2 OR2X2_770 ( .A(u2__abc_52155_new_n5380_), .B(u2__abc_52155_new_n4995_), .Y(u2__abc_52155_new_n5381_));
OR2X2 OR2X2_771 ( .A(u2__abc_52155_new_n5383_), .B(u2__abc_52155_new_n5375_), .Y(u2__abc_52155_new_n5384_));
OR2X2 OR2X2_772 ( .A(u2__abc_52155_new_n5385_), .B(u2__abc_52155_new_n5034_), .Y(u2__abc_52155_new_n5386_));
OR2X2 OR2X2_773 ( .A(u2__abc_52155_new_n5388_), .B(u2__abc_52155_new_n5026_), .Y(u2__abc_52155_new_n5389_));
OR2X2 OR2X2_774 ( .A(u2__abc_52155_new_n5387_), .B(u2__abc_52155_new_n5389_), .Y(u2__abc_52155_new_n5390_));
OR2X2 OR2X2_775 ( .A(u2__abc_52155_new_n5392_), .B(u2__abc_52155_new_n5374_), .Y(u2__abc_52155_new_n5393_));
OR2X2 OR2X2_776 ( .A(u2__abc_52155_new_n5394_), .B(u2__abc_52155_new_n4974_), .Y(u2__abc_52155_new_n5395_));
OR2X2 OR2X2_777 ( .A(u2__abc_52155_new_n5397_), .B(u2__abc_52155_new_n4966_), .Y(u2__abc_52155_new_n5398_));
OR2X2 OR2X2_778 ( .A(u2__abc_52155_new_n5396_), .B(u2__abc_52155_new_n5398_), .Y(u2__abc_52155_new_n5399_));
OR2X2 OR2X2_779 ( .A(u2__abc_52155_new_n5401_), .B(u2__abc_52155_new_n4943_), .Y(u2__abc_52155_new_n5402_));
OR2X2 OR2X2_78 ( .A(_abc_73687_new_n753_), .B(\a[38] ), .Y(_abc_73687_new_n945_));
OR2X2 OR2X2_780 ( .A(u2__abc_52155_new_n5404_), .B(u2__abc_52155_new_n4935_), .Y(u2__abc_52155_new_n5405_));
OR2X2 OR2X2_781 ( .A(u2__abc_52155_new_n5403_), .B(u2__abc_52155_new_n5405_), .Y(u2__abc_52155_new_n5406_));
OR2X2 OR2X2_782 ( .A(u2__abc_52155_new_n5400_), .B(u2__abc_52155_new_n5406_), .Y(u2__abc_52155_new_n5407_));
OR2X2 OR2X2_783 ( .A(u2__abc_52155_new_n5409_), .B(u2__abc_52155_new_n5373_), .Y(u2__abc_52155_new_n5410_));
OR2X2 OR2X2_784 ( .A(u2__abc_52155_new_n5411_), .B(u2__abc_52155_new_n4917_), .Y(u2__abc_52155_new_n5412_));
OR2X2 OR2X2_785 ( .A(u2__abc_52155_new_n5414_), .B(u2__abc_52155_new_n4902_), .Y(u2__abc_52155_new_n5415_));
OR2X2 OR2X2_786 ( .A(u2__abc_52155_new_n5413_), .B(u2__abc_52155_new_n5415_), .Y(u2__abc_52155_new_n5416_));
OR2X2 OR2X2_787 ( .A(u2__abc_52155_new_n5418_), .B(u2__abc_52155_new_n4871_), .Y(u2__abc_52155_new_n5419_));
OR2X2 OR2X2_788 ( .A(u2__abc_52155_new_n5420_), .B(u2__abc_52155_new_n4879_), .Y(u2__abc_52155_new_n5421_));
OR2X2 OR2X2_789 ( .A(u2__abc_52155_new_n5422_), .B(u2__abc_52155_new_n5419_), .Y(u2__abc_52155_new_n5423_));
OR2X2 OR2X2_79 ( .A(aNan), .B(sqrto_115_), .Y(_abc_73687_new_n947_));
OR2X2 OR2X2_790 ( .A(u2__abc_52155_new_n5417_), .B(u2__abc_52155_new_n5423_), .Y(u2__abc_52155_new_n5424_));
OR2X2 OR2X2_791 ( .A(u2__abc_52155_new_n5426_), .B(u2__abc_52155_new_n4808_), .Y(u2__abc_52155_new_n5427_));
OR2X2 OR2X2_792 ( .A(u2__abc_52155_new_n5429_), .B(u2__abc_52155_new_n4823_), .Y(u2__abc_52155_new_n5430_));
OR2X2 OR2X2_793 ( .A(u2__abc_52155_new_n5428_), .B(u2__abc_52155_new_n5430_), .Y(u2__abc_52155_new_n5431_));
OR2X2 OR2X2_794 ( .A(u2__abc_52155_new_n5433_), .B(u2__abc_52155_new_n4847_), .Y(u2__abc_52155_new_n5434_));
OR2X2 OR2X2_795 ( .A(u2__abc_52155_new_n5436_), .B(u2__abc_52155_new_n4839_), .Y(u2__abc_52155_new_n5437_));
OR2X2 OR2X2_796 ( .A(u2__abc_52155_new_n5435_), .B(u2__abc_52155_new_n5437_), .Y(u2__abc_52155_new_n5438_));
OR2X2 OR2X2_797 ( .A(u2__abc_52155_new_n5432_), .B(u2__abc_52155_new_n5438_), .Y(u2__abc_52155_new_n5439_));
OR2X2 OR2X2_798 ( .A(u2__abc_52155_new_n5425_), .B(u2__abc_52155_new_n5439_), .Y(u2__abc_52155_new_n5440_));
OR2X2 OR2X2_799 ( .A(u2__abc_52155_new_n5443_), .B(u2__abc_52155_new_n5290_), .Y(u2__abc_52155_new_n5444_));
OR2X2 OR2X2_8 ( .A(_abc_73687_new_n753_), .B(\a[3] ), .Y(_abc_73687_new_n840_));
OR2X2 OR2X2_80 ( .A(_abc_73687_new_n753_), .B(\a[39] ), .Y(_abc_73687_new_n948_));
OR2X2 OR2X2_800 ( .A(u2__abc_52155_new_n4782_), .B(u2__abc_52155_new_n4785_), .Y(u2__abc_52155_new_n5449_));
OR2X2 OR2X2_801 ( .A(u2__abc_52155_new_n5450_), .B(u2__abc_52155_new_n4775_), .Y(u2__abc_52155_new_n5451_));
OR2X2 OR2X2_802 ( .A(u2__abc_52155_new_n5453_), .B(u2__abc_52155_new_n4773_), .Y(u2__abc_52155_new_n5454_));
OR2X2 OR2X2_803 ( .A(u2__abc_52155_new_n5456_), .B(u2__abc_52155_new_n5448_), .Y(u2__abc_52155_new_n5457_));
OR2X2 OR2X2_804 ( .A(u2__abc_52155_new_n5458_), .B(u2__abc_52155_new_n4753_), .Y(u2__abc_52155_new_n5459_));
OR2X2 OR2X2_805 ( .A(u2__abc_52155_new_n5461_), .B(u2__abc_52155_new_n4745_), .Y(u2__abc_52155_new_n5462_));
OR2X2 OR2X2_806 ( .A(u2__abc_52155_new_n5460_), .B(u2__abc_52155_new_n5462_), .Y(u2__abc_52155_new_n5463_));
OR2X2 OR2X2_807 ( .A(u2__abc_52155_new_n5465_), .B(u2__abc_52155_new_n5447_), .Y(u2__abc_52155_new_n5466_));
OR2X2 OR2X2_808 ( .A(u2__abc_52155_new_n5467_), .B(u2__abc_52155_new_n4690_), .Y(u2__abc_52155_new_n5468_));
OR2X2 OR2X2_809 ( .A(u2__abc_52155_new_n5470_), .B(u2__abc_52155_new_n4682_), .Y(u2__abc_52155_new_n5471_));
OR2X2 OR2X2_81 ( .A(aNan), .B(sqrto_116_), .Y(_abc_73687_new_n950_));
OR2X2 OR2X2_810 ( .A(u2__abc_52155_new_n5469_), .B(u2__abc_52155_new_n5471_), .Y(u2__abc_52155_new_n5472_));
OR2X2 OR2X2_811 ( .A(u2__abc_52155_new_n5474_), .B(u2__abc_52155_new_n4721_), .Y(u2__abc_52155_new_n5475_));
OR2X2 OR2X2_812 ( .A(u2__abc_52155_new_n5477_), .B(u2__abc_52155_new_n4713_), .Y(u2__abc_52155_new_n5478_));
OR2X2 OR2X2_813 ( .A(u2__abc_52155_new_n5476_), .B(u2__abc_52155_new_n5478_), .Y(u2__abc_52155_new_n5479_));
OR2X2 OR2X2_814 ( .A(u2__abc_52155_new_n5473_), .B(u2__abc_52155_new_n5479_), .Y(u2__abc_52155_new_n5480_));
OR2X2 OR2X2_815 ( .A(u2__abc_52155_new_n5482_), .B(u2__abc_52155_new_n5446_), .Y(u2__abc_52155_new_n5483_));
OR2X2 OR2X2_816 ( .A(u2__abc_52155_new_n5484_), .B(u2__abc_52155_new_n4633_), .Y(u2__abc_52155_new_n5485_));
OR2X2 OR2X2_817 ( .A(u2__abc_52155_new_n5487_), .B(u2__abc_52155_new_n4618_), .Y(u2__abc_52155_new_n5488_));
OR2X2 OR2X2_818 ( .A(u2__abc_52155_new_n5486_), .B(u2__abc_52155_new_n5488_), .Y(u2__abc_52155_new_n5489_));
OR2X2 OR2X2_819 ( .A(u2__abc_52155_new_n5491_), .B(u2__abc_52155_new_n4657_), .Y(u2__abc_52155_new_n5492_));
OR2X2 OR2X2_82 ( .A(_abc_73687_new_n753_), .B(\a[40] ), .Y(_abc_73687_new_n951_));
OR2X2 OR2X2_820 ( .A(u2__abc_52155_new_n5494_), .B(u2__abc_52155_new_n4649_), .Y(u2__abc_52155_new_n5495_));
OR2X2 OR2X2_821 ( .A(u2__abc_52155_new_n5493_), .B(u2__abc_52155_new_n5495_), .Y(u2__abc_52155_new_n5496_));
OR2X2 OR2X2_822 ( .A(u2__abc_52155_new_n5490_), .B(u2__abc_52155_new_n5496_), .Y(u2__abc_52155_new_n5497_));
OR2X2 OR2X2_823 ( .A(u2__abc_52155_new_n5499_), .B(u2__abc_52155_new_n4570_), .Y(u2__abc_52155_new_n5500_));
OR2X2 OR2X2_824 ( .A(u2__abc_52155_new_n5502_), .B(u2__abc_52155_new_n4555_), .Y(u2__abc_52155_new_n5503_));
OR2X2 OR2X2_825 ( .A(u2__abc_52155_new_n5501_), .B(u2__abc_52155_new_n5503_), .Y(u2__abc_52155_new_n5504_));
OR2X2 OR2X2_826 ( .A(u2__abc_52155_new_n5506_), .B(u2__abc_52155_new_n4586_), .Y(u2__abc_52155_new_n5507_));
OR2X2 OR2X2_827 ( .A(u2__abc_52155_new_n5508_), .B(u2__abc_52155_new_n4594_), .Y(u2__abc_52155_new_n5509_));
OR2X2 OR2X2_828 ( .A(u2__abc_52155_new_n5510_), .B(u2__abc_52155_new_n5507_), .Y(u2__abc_52155_new_n5511_));
OR2X2 OR2X2_829 ( .A(u2__abc_52155_new_n5505_), .B(u2__abc_52155_new_n5511_), .Y(u2__abc_52155_new_n5512_));
OR2X2 OR2X2_83 ( .A(aNan), .B(sqrto_117_), .Y(_abc_73687_new_n953_));
OR2X2 OR2X2_830 ( .A(u2__abc_52155_new_n5498_), .B(u2__abc_52155_new_n5512_), .Y(u2__abc_52155_new_n5513_));
OR2X2 OR2X2_831 ( .A(u2__abc_52155_new_n5515_), .B(u2__abc_52155_new_n5445_), .Y(u2__abc_52155_new_n5516_));
OR2X2 OR2X2_832 ( .A(u2__abc_52155_new_n5517_), .B(u2__abc_52155_new_n4498_), .Y(u2__abc_52155_new_n5518_));
OR2X2 OR2X2_833 ( .A(u2__abc_52155_new_n5520_), .B(u2__abc_52155_new_n4490_), .Y(u2__abc_52155_new_n5521_));
OR2X2 OR2X2_834 ( .A(u2__abc_52155_new_n5519_), .B(u2__abc_52155_new_n5521_), .Y(u2__abc_52155_new_n5522_));
OR2X2 OR2X2_835 ( .A(u2__abc_52155_new_n5524_), .B(u2__abc_52155_new_n4529_), .Y(u2__abc_52155_new_n5525_));
OR2X2 OR2X2_836 ( .A(u2__abc_52155_new_n5527_), .B(u2__abc_52155_new_n4521_), .Y(u2__abc_52155_new_n5528_));
OR2X2 OR2X2_837 ( .A(u2__abc_52155_new_n5526_), .B(u2__abc_52155_new_n5528_), .Y(u2__abc_52155_new_n5529_));
OR2X2 OR2X2_838 ( .A(u2__abc_52155_new_n5523_), .B(u2__abc_52155_new_n5529_), .Y(u2__abc_52155_new_n5530_));
OR2X2 OR2X2_839 ( .A(u2__abc_52155_new_n5532_), .B(u2__abc_52155_new_n4466_), .Y(u2__abc_52155_new_n5533_));
OR2X2 OR2X2_84 ( .A(_abc_73687_new_n753_), .B(\a[41] ), .Y(_abc_73687_new_n954_));
OR2X2 OR2X2_840 ( .A(u2__abc_52155_new_n5535_), .B(u2__abc_52155_new_n4458_), .Y(u2__abc_52155_new_n5536_));
OR2X2 OR2X2_841 ( .A(u2__abc_52155_new_n5534_), .B(u2__abc_52155_new_n5536_), .Y(u2__abc_52155_new_n5537_));
OR2X2 OR2X2_842 ( .A(u2__abc_52155_new_n5539_), .B(u2__abc_52155_new_n4435_), .Y(u2__abc_52155_new_n5540_));
OR2X2 OR2X2_843 ( .A(u2__abc_52155_new_n5542_), .B(u2__abc_52155_new_n4427_), .Y(u2__abc_52155_new_n5543_));
OR2X2 OR2X2_844 ( .A(u2__abc_52155_new_n5541_), .B(u2__abc_52155_new_n5543_), .Y(u2__abc_52155_new_n5544_));
OR2X2 OR2X2_845 ( .A(u2__abc_52155_new_n5538_), .B(u2__abc_52155_new_n5544_), .Y(u2__abc_52155_new_n5545_));
OR2X2 OR2X2_846 ( .A(u2__abc_52155_new_n5531_), .B(u2__abc_52155_new_n5545_), .Y(u2__abc_52155_new_n5546_));
OR2X2 OR2X2_847 ( .A(u2__abc_52155_new_n5548_), .B(u2__abc_52155_new_n4300_), .Y(u2__abc_52155_new_n5549_));
OR2X2 OR2X2_848 ( .A(u2__abc_52155_new_n5551_), .B(u2__abc_52155_new_n4315_), .Y(u2__abc_52155_new_n5552_));
OR2X2 OR2X2_849 ( .A(u2__abc_52155_new_n5550_), .B(u2__abc_52155_new_n5552_), .Y(u2__abc_52155_new_n5553_));
OR2X2 OR2X2_85 ( .A(aNan), .B(sqrto_118_), .Y(_abc_73687_new_n956_));
OR2X2 OR2X2_850 ( .A(u2__abc_52155_new_n5555_), .B(u2__abc_52155_new_n4328_), .Y(u2__abc_52155_new_n5556_));
OR2X2 OR2X2_851 ( .A(u2__abc_52155_new_n5557_), .B(u2__abc_52155_new_n4339_), .Y(u2__abc_52155_new_n5558_));
OR2X2 OR2X2_852 ( .A(u2__abc_52155_new_n5559_), .B(u2__abc_52155_new_n5556_), .Y(u2__abc_52155_new_n5560_));
OR2X2 OR2X2_853 ( .A(u2__abc_52155_new_n5554_), .B(u2__abc_52155_new_n5560_), .Y(u2__abc_52155_new_n5561_));
OR2X2 OR2X2_854 ( .A(u2__abc_52155_new_n5562_), .B(u2__abc_52155_new_n4363_), .Y(u2__abc_52155_new_n5563_));
OR2X2 OR2X2_855 ( .A(u2__abc_52155_new_n5565_), .B(u2__abc_52155_new_n4378_), .Y(u2__abc_52155_new_n5566_));
OR2X2 OR2X2_856 ( .A(u2__abc_52155_new_n5564_), .B(u2__abc_52155_new_n5566_), .Y(u2__abc_52155_new_n5567_));
OR2X2 OR2X2_857 ( .A(u2__abc_52155_new_n5569_), .B(u2__abc_52155_new_n4394_), .Y(u2__abc_52155_new_n5570_));
OR2X2 OR2X2_858 ( .A(u2__abc_52155_new_n5571_), .B(u2__abc_52155_new_n4402_), .Y(u2__abc_52155_new_n5572_));
OR2X2 OR2X2_859 ( .A(u2__abc_52155_new_n5573_), .B(u2__abc_52155_new_n5570_), .Y(u2__abc_52155_new_n5574_));
OR2X2 OR2X2_86 ( .A(_abc_73687_new_n753_), .B(\a[42] ), .Y(_abc_73687_new_n957_));
OR2X2 OR2X2_860 ( .A(u2__abc_52155_new_n5568_), .B(u2__abc_52155_new_n5574_), .Y(u2__abc_52155_new_n5575_));
OR2X2 OR2X2_861 ( .A(u2__abc_52155_new_n5576_), .B(u2__abc_52155_new_n5561_), .Y(u2__abc_52155_new_n5577_));
OR2X2 OR2X2_862 ( .A(u2__abc_52155_new_n5547_), .B(u2__abc_52155_new_n5577_), .Y(u2__abc_52155_new_n5578_));
OR2X2 OR2X2_863 ( .A(u2__abc_52155_new_n5582_), .B(u2__abc_52155_new_n6606_), .Y(u2__abc_52155_new_n6607_));
OR2X2 OR2X2_864 ( .A(u2__abc_52155_new_n6611_), .B(u2__abc_52155_new_n6451_), .Y(u2__abc_52155_new_n6612_));
OR2X2 OR2X2_865 ( .A(u2__abc_52155_new_n6615_), .B(u2__abc_52155_new_n6435_), .Y(u2__abc_52155_new_n6616_));
OR2X2 OR2X2_866 ( .A(u2__abc_52155_new_n6614_), .B(u2__abc_52155_new_n6616_), .Y(u2__abc_52155_new_n6617_));
OR2X2 OR2X2_867 ( .A(u2__abc_52155_new_n6618_), .B(u2__abc_52155_new_n6423_), .Y(u2__abc_52155_new_n6619_));
OR2X2 OR2X2_868 ( .A(u2__abc_52155_new_n6621_), .B(u2__abc_52155_new_n6459_), .Y(u2__abc_52155_new_n6622_));
OR2X2 OR2X2_869 ( .A(u2__abc_52155_new_n6624_), .B(u2__abc_52155_new_n6466_), .Y(u2__abc_52155_new_n6625_));
OR2X2 OR2X2_87 ( .A(aNan), .B(sqrto_119_), .Y(_abc_73687_new_n959_));
OR2X2 OR2X2_870 ( .A(u2__abc_52155_new_n6623_), .B(u2__abc_52155_new_n6625_), .Y(u2__abc_52155_new_n6626_));
OR2X2 OR2X2_871 ( .A(u2__abc_52155_new_n6627_), .B(u2__abc_52155_new_n6610_), .Y(u2__abc_52155_new_n6628_));
OR2X2 OR2X2_872 ( .A(u2__abc_52155_new_n6633_), .B(u2__abc_52155_new_n6550_), .Y(u2__abc_52155_new_n6634_));
OR2X2 OR2X2_873 ( .A(u2__abc_52155_new_n6632_), .B(u2__abc_52155_new_n6634_), .Y(u2__abc_52155_new_n6635_));
OR2X2 OR2X2_874 ( .A(u2__abc_52155_new_n6636_), .B(u2__abc_52155_new_n6565_), .Y(u2__abc_52155_new_n6637_));
OR2X2 OR2X2_875 ( .A(u2__abc_52155_new_n6639_), .B(u2__abc_52155_new_n6631_), .Y(u2__abc_52155_new_n6640_));
OR2X2 OR2X2_876 ( .A(u2__abc_52155_new_n6642_), .B(u2__abc_52155_new_n6593_), .Y(u2__abc_52155_new_n6643_));
OR2X2 OR2X2_877 ( .A(u2__abc_52155_new_n6641_), .B(u2__abc_52155_new_n6643_), .Y(u2__abc_52155_new_n6644_));
OR2X2 OR2X2_878 ( .A(u2__abc_52155_new_n6645_), .B(u2__abc_52155_new_n6581_), .Y(u2__abc_52155_new_n6646_));
OR2X2 OR2X2_879 ( .A(u2__abc_52155_new_n6649_), .B(u2__abc_52155_new_n6630_), .Y(u2__abc_52155_new_n6650_));
OR2X2 OR2X2_88 ( .A(_abc_73687_new_n753_), .B(\a[43] ), .Y(_abc_73687_new_n960_));
OR2X2 OR2X2_880 ( .A(u2__abc_52155_new_n6653_), .B(u2__abc_52155_new_n6533_), .Y(u2__abc_52155_new_n6654_));
OR2X2 OR2X2_881 ( .A(u2__abc_52155_new_n6652_), .B(u2__abc_52155_new_n6654_), .Y(u2__abc_52155_new_n6655_));
OR2X2 OR2X2_882 ( .A(u2__abc_52155_new_n6656_), .B(u2__abc_52155_new_n6518_), .Y(u2__abc_52155_new_n6657_));
OR2X2 OR2X2_883 ( .A(u2__abc_52155_new_n6659_), .B(u2__abc_52155_new_n6651_), .Y(u2__abc_52155_new_n6660_));
OR2X2 OR2X2_884 ( .A(u2__abc_52155_new_n6661_), .B(u2__abc_52155_new_n6487_), .Y(u2__abc_52155_new_n6662_));
OR2X2 OR2X2_885 ( .A(u2__abc_52155_new_n6664_), .B(u2__abc_52155_new_n6499_), .Y(u2__abc_52155_new_n6665_));
OR2X2 OR2X2_886 ( .A(u2__abc_52155_new_n6663_), .B(u2__abc_52155_new_n6665_), .Y(u2__abc_52155_new_n6666_));
OR2X2 OR2X2_887 ( .A(u2__abc_52155_new_n6669_), .B(u2__abc_52155_new_n6629_), .Y(u2__abc_52155_new_n6670_));
OR2X2 OR2X2_888 ( .A(u2__abc_52155_new_n6673_), .B(u2__abc_52155_new_n6372_), .Y(u2__abc_52155_new_n6674_));
OR2X2 OR2X2_889 ( .A(u2__abc_52155_new_n6672_), .B(u2__abc_52155_new_n6674_), .Y(u2__abc_52155_new_n6675_));
OR2X2 OR2X2_89 ( .A(aNan), .B(sqrto_120_), .Y(_abc_73687_new_n962_));
OR2X2 OR2X2_890 ( .A(u2__abc_52155_new_n6676_), .B(u2__abc_52155_new_n6360_), .Y(u2__abc_52155_new_n6677_));
OR2X2 OR2X2_891 ( .A(u2__abc_52155_new_n6679_), .B(u2__abc_52155_new_n6671_), .Y(u2__abc_52155_new_n6680_));
OR2X2 OR2X2_892 ( .A(u2__abc_52155_new_n6682_), .B(u2__abc_52155_new_n6403_), .Y(u2__abc_52155_new_n6683_));
OR2X2 OR2X2_893 ( .A(u2__abc_52155_new_n6681_), .B(u2__abc_52155_new_n6683_), .Y(u2__abc_52155_new_n6684_));
OR2X2 OR2X2_894 ( .A(u2__abc_52155_new_n6685_), .B(u2__abc_52155_new_n6388_), .Y(u2__abc_52155_new_n6686_));
OR2X2 OR2X2_895 ( .A(u2__abc_52155_new_n6690_), .B(u2__abc_52155_new_n6609_), .Y(u2__abc_52155_new_n6691_));
OR2X2 OR2X2_896 ( .A(u2__abc_52155_new_n6695_), .B(u2__abc_52155_new_n6168_), .Y(u2__abc_52155_new_n6696_));
OR2X2 OR2X2_897 ( .A(u2__abc_52155_new_n6694_), .B(u2__abc_52155_new_n6696_), .Y(u2__abc_52155_new_n6697_));
OR2X2 OR2X2_898 ( .A(u2__abc_52155_new_n6698_), .B(u2__abc_52155_new_n6183_), .Y(u2__abc_52155_new_n6699_));
OR2X2 OR2X2_899 ( .A(u2__abc_52155_new_n6701_), .B(u2__abc_52155_new_n6211_), .Y(u2__abc_52155_new_n6702_));
OR2X2 OR2X2_9 ( .A(aNan), .B(sqrto_80_), .Y(_abc_73687_new_n842_));
OR2X2 OR2X2_90 ( .A(_abc_73687_new_n753_), .B(\a[44] ), .Y(_abc_73687_new_n963_));
OR2X2 OR2X2_900 ( .A(u2__abc_52155_new_n6189_), .B(u2__abc_52155_new_n6204_), .Y(u2__abc_52155_new_n6704_));
OR2X2 OR2X2_901 ( .A(u2__abc_52155_new_n6703_), .B(u2__abc_52155_new_n6704_), .Y(u2__abc_52155_new_n6705_));
OR2X2 OR2X2_902 ( .A(u2__abc_52155_new_n6706_), .B(u2__abc_52155_new_n6196_), .Y(u2__abc_52155_new_n6707_));
OR2X2 OR2X2_903 ( .A(u2__abc_52155_new_n6708_), .B(u2__abc_52155_new_n6692_), .Y(u2__abc_52155_new_n6709_));
OR2X2 OR2X2_904 ( .A(u2__abc_52155_new_n6095_), .B(u2__abc_52155_new_n6117_), .Y(u2__abc_52155_new_n6712_));
OR2X2 OR2X2_905 ( .A(u2__abc_52155_new_n6711_), .B(u2__abc_52155_new_n6712_), .Y(u2__abc_52155_new_n6713_));
OR2X2 OR2X2_906 ( .A(u2__abc_52155_new_n6714_), .B(u2__abc_52155_new_n6102_), .Y(u2__abc_52155_new_n6715_));
OR2X2 OR2X2_907 ( .A(u2__abc_52155_new_n6716_), .B(u2__abc_52155_new_n6141_), .Y(u2__abc_52155_new_n6717_));
OR2X2 OR2X2_908 ( .A(u2__abc_52155_new_n6126_), .B(u2__abc_52155_new_n6148_), .Y(u2__abc_52155_new_n6719_));
OR2X2 OR2X2_909 ( .A(u2__abc_52155_new_n6718_), .B(u2__abc_52155_new_n6719_), .Y(u2__abc_52155_new_n6720_));
OR2X2 OR2X2_91 ( .A(aNan), .B(sqrto_121_), .Y(_abc_73687_new_n965_));
OR2X2 OR2X2_910 ( .A(u2__abc_52155_new_n6721_), .B(u2__abc_52155_new_n6133_), .Y(u2__abc_52155_new_n6722_));
OR2X2 OR2X2_911 ( .A(u2__abc_52155_new_n6727_), .B(u2__abc_52155_new_n6292_), .Y(u2__abc_52155_new_n6728_));
OR2X2 OR2X2_912 ( .A(u2__abc_52155_new_n6730_), .B(u2__abc_52155_new_n6307_), .Y(u2__abc_52155_new_n6731_));
OR2X2 OR2X2_913 ( .A(u2__abc_52155_new_n6729_), .B(u2__abc_52155_new_n6731_), .Y(u2__abc_52155_new_n6732_));
OR2X2 OR2X2_914 ( .A(u2__abc_52155_new_n6733_), .B(u2__abc_52155_new_n6726_), .Y(u2__abc_52155_new_n6734_));
OR2X2 OR2X2_915 ( .A(u2__abc_52155_new_n6736_), .B(u2__abc_52155_new_n6338_), .Y(u2__abc_52155_new_n6737_));
OR2X2 OR2X2_916 ( .A(u2__abc_52155_new_n6735_), .B(u2__abc_52155_new_n6737_), .Y(u2__abc_52155_new_n6738_));
OR2X2 OR2X2_917 ( .A(u2__abc_52155_new_n6739_), .B(u2__abc_52155_new_n6326_), .Y(u2__abc_52155_new_n6740_));
OR2X2 OR2X2_918 ( .A(u2__abc_52155_new_n6743_), .B(u2__abc_52155_new_n6725_), .Y(u2__abc_52155_new_n6744_));
OR2X2 OR2X2_919 ( .A(u2__abc_52155_new_n6747_), .B(u2__abc_52155_new_n6232_), .Y(u2__abc_52155_new_n6748_));
OR2X2 OR2X2_92 ( .A(_abc_73687_new_n753_), .B(\a[45] ), .Y(_abc_73687_new_n966_));
OR2X2 OR2X2_920 ( .A(u2__abc_52155_new_n6746_), .B(u2__abc_52155_new_n6748_), .Y(u2__abc_52155_new_n6749_));
OR2X2 OR2X2_921 ( .A(u2__abc_52155_new_n6750_), .B(u2__abc_52155_new_n6247_), .Y(u2__abc_52155_new_n6751_));
OR2X2 OR2X2_922 ( .A(u2__abc_52155_new_n6753_), .B(u2__abc_52155_new_n6745_), .Y(u2__abc_52155_new_n6754_));
OR2X2 OR2X2_923 ( .A(u2__abc_52155_new_n6756_), .B(u2__abc_52155_new_n6275_), .Y(u2__abc_52155_new_n6757_));
OR2X2 OR2X2_924 ( .A(u2__abc_52155_new_n6755_), .B(u2__abc_52155_new_n6757_), .Y(u2__abc_52155_new_n6758_));
OR2X2 OR2X2_925 ( .A(u2__abc_52155_new_n6759_), .B(u2__abc_52155_new_n6263_), .Y(u2__abc_52155_new_n6760_));
OR2X2 OR2X2_926 ( .A(u2__abc_52155_new_n6764_), .B(u2__abc_52155_new_n6724_), .Y(u2__abc_52155_new_n6765_));
OR2X2 OR2X2_927 ( .A(u2__abc_52155_new_n6768_), .B(u2__abc_52155_new_n6608_), .Y(u2__abc_52155_new_n6769_));
OR2X2 OR2X2_928 ( .A(u2__abc_52155_new_n6775_), .B(u2__abc_52155_new_n6070_), .Y(u2__abc_52155_new_n6776_));
OR2X2 OR2X2_929 ( .A(u2__abc_52155_new_n6774_), .B(u2__abc_52155_new_n6776_), .Y(u2__abc_52155_new_n6777_));
OR2X2 OR2X2_93 ( .A(aNan), .B(sqrto_122_), .Y(_abc_73687_new_n968_));
OR2X2 OR2X2_930 ( .A(u2__abc_52155_new_n6079_), .B(u2__abc_52155_new_n6082_), .Y(u2__abc_52155_new_n6778_));
OR2X2 OR2X2_931 ( .A(u2__abc_52155_new_n6780_), .B(u2__abc_52155_new_n6773_), .Y(u2__abc_52155_new_n6781_));
OR2X2 OR2X2_932 ( .A(u2__abc_52155_new_n6782_), .B(u2__abc_52155_new_n6039_), .Y(u2__abc_52155_new_n6783_));
OR2X2 OR2X2_933 ( .A(u2__abc_52155_new_n6785_), .B(u2__abc_52155_new_n6051_), .Y(u2__abc_52155_new_n6786_));
OR2X2 OR2X2_934 ( .A(u2__abc_52155_new_n6784_), .B(u2__abc_52155_new_n6786_), .Y(u2__abc_52155_new_n6787_));
OR2X2 OR2X2_935 ( .A(u2__abc_52155_new_n6789_), .B(u2__abc_52155_new_n6772_), .Y(u2__abc_52155_new_n6790_));
OR2X2 OR2X2_936 ( .A(u2__abc_52155_new_n6793_), .B(u2__abc_52155_new_n5976_), .Y(u2__abc_52155_new_n6794_));
OR2X2 OR2X2_937 ( .A(u2__abc_52155_new_n6792_), .B(u2__abc_52155_new_n6794_), .Y(u2__abc_52155_new_n6795_));
OR2X2 OR2X2_938 ( .A(u2__abc_52155_new_n6796_), .B(u2__abc_52155_new_n5991_), .Y(u2__abc_52155_new_n6797_));
OR2X2 OR2X2_939 ( .A(u2__abc_52155_new_n6799_), .B(u2__abc_52155_new_n6791_), .Y(u2__abc_52155_new_n6800_));
OR2X2 OR2X2_94 ( .A(_abc_73687_new_n753_), .B(\a[46] ), .Y(_abc_73687_new_n969_));
OR2X2 OR2X2_940 ( .A(u2__abc_52155_new_n6802_), .B(u2__abc_52155_new_n6019_), .Y(u2__abc_52155_new_n6803_));
OR2X2 OR2X2_941 ( .A(u2__abc_52155_new_n6801_), .B(u2__abc_52155_new_n6803_), .Y(u2__abc_52155_new_n6804_));
OR2X2 OR2X2_942 ( .A(u2__abc_52155_new_n6805_), .B(u2__abc_52155_new_n6004_), .Y(u2__abc_52155_new_n6806_));
OR2X2 OR2X2_943 ( .A(u2__abc_52155_new_n6809_), .B(u2__abc_52155_new_n6771_), .Y(u2__abc_52155_new_n6810_));
OR2X2 OR2X2_944 ( .A(u2__abc_52155_new_n6813_), .B(u2__abc_52155_new_n5861_), .Y(u2__abc_52155_new_n6814_));
OR2X2 OR2X2_945 ( .A(u2__abc_52155_new_n6812_), .B(u2__abc_52155_new_n6814_), .Y(u2__abc_52155_new_n6815_));
OR2X2 OR2X2_946 ( .A(u2__abc_52155_new_n6816_), .B(u2__abc_52155_new_n5849_), .Y(u2__abc_52155_new_n6817_));
OR2X2 OR2X2_947 ( .A(u2__abc_52155_new_n6819_), .B(u2__abc_52155_new_n6811_), .Y(u2__abc_52155_new_n6820_));
OR2X2 OR2X2_948 ( .A(u2__abc_52155_new_n6822_), .B(u2__abc_52155_new_n5892_), .Y(u2__abc_52155_new_n6823_));
OR2X2 OR2X2_949 ( .A(u2__abc_52155_new_n6821_), .B(u2__abc_52155_new_n6823_), .Y(u2__abc_52155_new_n6824_));
OR2X2 OR2X2_95 ( .A(aNan), .B(sqrto_123_), .Y(_abc_73687_new_n971_));
OR2X2 OR2X2_950 ( .A(u2__abc_52155_new_n6825_), .B(u2__abc_52155_new_n5880_), .Y(u2__abc_52155_new_n6826_));
OR2X2 OR2X2_951 ( .A(u2__abc_52155_new_n6831_), .B(u2__abc_52155_new_n5943_), .Y(u2__abc_52155_new_n6832_));
OR2X2 OR2X2_952 ( .A(u2__abc_52155_new_n6835_), .B(u2__abc_52155_new_n5909_), .Y(u2__abc_52155_new_n6836_));
OR2X2 OR2X2_953 ( .A(u2__abc_52155_new_n6838_), .B(u2__abc_52155_new_n5924_), .Y(u2__abc_52155_new_n6839_));
OR2X2 OR2X2_954 ( .A(u2__abc_52155_new_n6837_), .B(u2__abc_52155_new_n6839_), .Y(u2__abc_52155_new_n6840_));
OR2X2 OR2X2_955 ( .A(u2__abc_52155_new_n6841_), .B(u2__abc_52155_new_n5948_), .Y(u2__abc_52155_new_n6842_));
OR2X2 OR2X2_956 ( .A(u2__abc_52155_new_n6844_), .B(u2__abc_52155_new_n5955_), .Y(u2__abc_52155_new_n6845_));
OR2X2 OR2X2_957 ( .A(u2__abc_52155_new_n6843_), .B(u2__abc_52155_new_n6845_), .Y(u2__abc_52155_new_n6846_));
OR2X2 OR2X2_958 ( .A(u2__abc_52155_new_n6847_), .B(u2__abc_52155_new_n6830_), .Y(u2__abc_52155_new_n6848_));
OR2X2 OR2X2_959 ( .A(u2__abc_52155_new_n6850_), .B(u2__abc_52155_new_n6770_), .Y(u2__abc_52155_new_n6851_));
OR2X2 OR2X2_96 ( .A(_abc_73687_new_n753_), .B(\a[47] ), .Y(_abc_73687_new_n972_));
OR2X2 OR2X2_960 ( .A(u2__abc_52155_new_n6853_), .B(u2__abc_52155_new_n5693_), .Y(u2__abc_52155_new_n6854_));
OR2X2 OR2X2_961 ( .A(u2__abc_52155_new_n6856_), .B(u2__abc_52155_new_n5654_), .Y(u2__abc_52155_new_n6857_));
OR2X2 OR2X2_962 ( .A(u2__abc_52155_new_n6859_), .B(u2__abc_52155_new_n5669_), .Y(u2__abc_52155_new_n6860_));
OR2X2 OR2X2_963 ( .A(u2__abc_52155_new_n6858_), .B(u2__abc_52155_new_n6860_), .Y(u2__abc_52155_new_n6861_));
OR2X2 OR2X2_964 ( .A(u2__abc_52155_new_n6862_), .B(u2__abc_52155_new_n6855_), .Y(u2__abc_52155_new_n6863_));
OR2X2 OR2X2_965 ( .A(u2__abc_52155_new_n6864_), .B(u2__abc_52155_new_n5678_), .Y(u2__abc_52155_new_n6865_));
OR2X2 OR2X2_966 ( .A(u2__abc_52155_new_n6866_), .B(u2__abc_52155_new_n5685_), .Y(u2__abc_52155_new_n6867_));
OR2X2 OR2X2_967 ( .A(u2__abc_52155_new_n6868_), .B(u2__abc_52155_new_n6852_), .Y(u2__abc_52155_new_n6869_));
OR2X2 OR2X2_968 ( .A(u2__abc_52155_new_n5721_), .B(u2__abc_52155_new_n5726_), .Y(u2__abc_52155_new_n6874_));
OR2X2 OR2X2_969 ( .A(u2__abc_52155_new_n6873_), .B(u2__abc_52155_new_n6874_), .Y(u2__abc_52155_new_n6875_));
OR2X2 OR2X2_97 ( .A(aNan), .B(sqrto_124_), .Y(_abc_73687_new_n974_));
OR2X2 OR2X2_970 ( .A(u2__abc_52155_new_n5733_), .B(u2__abc_52155_new_n5757_), .Y(u2__abc_52155_new_n6877_));
OR2X2 OR2X2_971 ( .A(u2__abc_52155_new_n6876_), .B(u2__abc_52155_new_n6877_), .Y(u2__abc_52155_new_n6878_));
OR2X2 OR2X2_972 ( .A(u2__abc_52155_new_n5742_), .B(u2__abc_52155_new_n5764_), .Y(u2__abc_52155_new_n6880_));
OR2X2 OR2X2_973 ( .A(u2__abc_52155_new_n6879_), .B(u2__abc_52155_new_n6880_), .Y(u2__abc_52155_new_n6881_));
OR2X2 OR2X2_974 ( .A(u2__abc_52155_new_n6882_), .B(u2__abc_52155_new_n5749_), .Y(u2__abc_52155_new_n6883_));
OR2X2 OR2X2_975 ( .A(u2__abc_52155_new_n6887_), .B(u2__abc_52155_new_n5781_), .Y(u2__abc_52155_new_n6888_));
OR2X2 OR2X2_976 ( .A(u2__abc_52155_new_n6890_), .B(u2__abc_52155_new_n5796_), .Y(u2__abc_52155_new_n6891_));
OR2X2 OR2X2_977 ( .A(u2__abc_52155_new_n6889_), .B(u2__abc_52155_new_n6891_), .Y(u2__abc_52155_new_n6892_));
OR2X2 OR2X2_978 ( .A(u2__abc_52155_new_n6893_), .B(u2__abc_52155_new_n5820_), .Y(u2__abc_52155_new_n6894_));
OR2X2 OR2X2_979 ( .A(u2__abc_52155_new_n5805_), .B(u2__abc_52155_new_n5827_), .Y(u2__abc_52155_new_n6896_));
OR2X2 OR2X2_98 ( .A(_abc_73687_new_n753_), .B(\a[48] ), .Y(_abc_73687_new_n975_));
OR2X2 OR2X2_980 ( .A(u2__abc_52155_new_n6895_), .B(u2__abc_52155_new_n6896_), .Y(u2__abc_52155_new_n6897_));
OR2X2 OR2X2_981 ( .A(u2__abc_52155_new_n6898_), .B(u2__abc_52155_new_n6900_), .Y(u2__abc_52155_new_n6901_));
OR2X2 OR2X2_982 ( .A(u2__abc_52155_new_n6902_), .B(u2__abc_52155_new_n6870_), .Y(u2__abc_52155_new_n6903_));
OR2X2 OR2X2_983 ( .A(u2__abc_52155_new_n6905_), .B(u2__abc_52155_new_n5637_), .Y(u2__abc_52155_new_n6906_));
OR2X2 OR2X2_984 ( .A(u2__abc_52155_new_n6908_), .B(u2__abc_52155_new_n5625_), .Y(u2__abc_52155_new_n6909_));
OR2X2 OR2X2_985 ( .A(u2__abc_52155_new_n6907_), .B(u2__abc_52155_new_n6909_), .Y(u2__abc_52155_new_n6910_));
OR2X2 OR2X2_986 ( .A(u2__abc_52155_new_n6911_), .B(u2__abc_52155_new_n6904_), .Y(u2__abc_52155_new_n6912_));
OR2X2 OR2X2_987 ( .A(u2__abc_52155_new_n6914_), .B(u2__abc_52155_new_n5606_), .Y(u2__abc_52155_new_n6915_));
OR2X2 OR2X2_988 ( .A(u2__abc_52155_new_n6913_), .B(u2__abc_52155_new_n6915_), .Y(u2__abc_52155_new_n6916_));
OR2X2 OR2X2_989 ( .A(u2__abc_52155_new_n6917_), .B(u2__abc_52155_new_n5591_), .Y(u2__abc_52155_new_n6918_));
OR2X2 OR2X2_99 ( .A(aNan), .B(sqrto_125_), .Y(_abc_73687_new_n977_));
OR2X2 OR2X2_990 ( .A(u2__abc_52155_new_n6926_), .B(u2__abc_52155_new_n7438_), .Y(u2__abc_52155_new_n7439_));
OR2X2 OR2X2_991 ( .A(u2__abc_52155_new_n7440_), .B(u2__abc_52155_new_n7229_), .Y(u2__abc_52155_new_n7441_));
OR2X2 OR2X2_992 ( .A(u2__abc_52155_new_n7443_), .B(u2__abc_52155_new_n7221_), .Y(u2__abc_52155_new_n7444_));
OR2X2 OR2X2_993 ( .A(u2__abc_52155_new_n7442_), .B(u2__abc_52155_new_n7444_), .Y(u2__abc_52155_new_n7445_));
OR2X2 OR2X2_994 ( .A(u2__abc_52155_new_n7447_), .B(u2__abc_52155_new_n7198_), .Y(u2__abc_52155_new_n7448_));
OR2X2 OR2X2_995 ( .A(u2__abc_52155_new_n7450_), .B(u2__abc_52155_new_n7193_), .Y(u2__abc_52155_new_n7451_));
OR2X2 OR2X2_996 ( .A(u2__abc_52155_new_n7449_), .B(u2__abc_52155_new_n7451_), .Y(u2__abc_52155_new_n7452_));
OR2X2 OR2X2_997 ( .A(u2__abc_52155_new_n7446_), .B(u2__abc_52155_new_n7452_), .Y(u2__abc_52155_new_n7453_));
OR2X2 OR2X2_998 ( .A(u2__abc_52155_new_n7455_), .B(u2__abc_52155_new_n7419_), .Y(u2__abc_52155_new_n7456_));
OR2X2 OR2X2_999 ( .A(u2__abc_52155_new_n7458_), .B(u2__abc_52155_new_n7414_), .Y(u2__abc_52155_new_n7459_));

assign \o[0]  = 1'h0;
assign \o[1]  = 1'h0;
assign \o[2]  = 1'h0;
assign \o[3]  = 1'h0;
assign \o[4]  = 1'h0;
assign \o[5]  = 1'h0;
assign \o[6]  = 1'h0;
assign \o[7]  = 1'h0;
assign \o[8]  = 1'h0;
assign \o[9]  = 1'h0;
assign \o[10]  = 1'h0;
assign \o[11]  = 1'h0;
assign \o[12]  = 1'h0;
assign \o[13]  = 1'h0;
assign \o[14]  = 1'h0;
assign \o[15]  = 1'h0;
assign \o[16]  = 1'h0;
assign \o[17]  = 1'h0;
assign \o[18]  = 1'h0;
assign \o[19]  = 1'h0;
assign \o[20]  = 1'h0;
assign \o[21]  = 1'h0;
assign \o[22]  = 1'h0;
assign \o[23]  = 1'h0;
assign \o[24]  = 1'h0;
assign \o[25]  = 1'h0;
assign \o[26]  = 1'h0;
assign \o[27]  = 1'h0;
assign \o[28]  = 1'h0;
assign \o[29]  = 1'h0;
assign \o[30]  = 1'h0;
assign \o[31]  = 1'h0;
assign \o[32]  = 1'h0;
assign \o[33]  = 1'h0;
assign \o[34]  = 1'h0;
assign \o[35]  = 1'h0;

endmodule