module FSM(clk, reset, \codif[0] , \codif[1] , \codif[2] , \codif[3] , \codif[4] , \codif[5] , \codif[6] , \codif[7] , \codif[8] , \codif[9] , \codif[10] , \codif[11] , busy_mem, done_mem, aligned_mem, done_exec, is_exec, \W_R_mem[0] , \W_R_mem[1] , \wordsize_mem[0] , \wordsize_mem[1] , sign_mem, en_mem, enable_exec, enable_exec_mem, trap, enable_pc);

output \W_R_mem[0] ;
output \W_R_mem[1] ;
wire _0W_R_mem_1_0__0_; 
wire _0W_R_mem_1_0__1_; 
wire _0en_mem_0_0_; 
wire _0enable_exec_0_0_; 
wire _0enable_exec_mem_0_0_; 
wire _0enable_pc_aux_0_0_; 
wire _0enable_pc_fsm_0_0_; 
wire _0trap_0_0_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_0_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_1_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_2_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_3_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_4_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_5_; 
wire _abc_801_auto_fsm_map_cc_170_map_fsm_238_6_; 
wire _abc_934_new_n100_; 
wire _abc_934_new_n101_; 
wire _abc_934_new_n102_; 
wire _abc_934_new_n103_; 
wire _abc_934_new_n105_; 
wire _abc_934_new_n106_; 
wire _abc_934_new_n107_; 
wire _abc_934_new_n108_; 
wire _abc_934_new_n110_; 
wire _abc_934_new_n111_; 
wire _abc_934_new_n114_; 
wire _abc_934_new_n116_; 
wire _abc_934_new_n117_; 
wire _abc_934_new_n118_; 
wire _abc_934_new_n119_; 
wire _abc_934_new_n120_; 
wire _abc_934_new_n121_; 
wire _abc_934_new_n122_; 
wire _abc_934_new_n123_; 
wire _abc_934_new_n124_; 
wire _abc_934_new_n125_; 
wire _abc_934_new_n126_; 
wire _abc_934_new_n127_; 
wire _abc_934_new_n128_; 
wire _abc_934_new_n129_; 
wire _abc_934_new_n130_; 
wire _abc_934_new_n131_; 
wire _abc_934_new_n132_; 
wire _abc_934_new_n134_; 
wire _abc_934_new_n135_; 
wire _abc_934_new_n136_; 
wire _abc_934_new_n137_; 
wire _abc_934_new_n138_; 
wire _abc_934_new_n139_; 
wire _abc_934_new_n140_; 
wire _abc_934_new_n141_; 
wire _abc_934_new_n142_; 
wire _abc_934_new_n143_; 
wire _abc_934_new_n144_; 
wire _abc_934_new_n145_; 
wire _abc_934_new_n146_; 
wire _abc_934_new_n149_; 
wire _abc_934_new_n150_; 
wire _abc_934_new_n151_; 
wire _abc_934_new_n152_; 
wire _abc_934_new_n153_; 
wire _abc_934_new_n154_; 
wire _abc_934_new_n155_; 
wire _abc_934_new_n156_; 
wire _abc_934_new_n157_; 
wire _abc_934_new_n158_; 
wire _abc_934_new_n160_; 
wire _abc_934_new_n162_; 
wire _abc_934_new_n163_; 
wire _abc_934_new_n164_; 
wire _abc_934_new_n165_; 
wire _abc_934_new_n166_; 
wire _abc_934_new_n167_; 
wire _abc_934_new_n168_; 
wire _abc_934_new_n169_; 
wire _abc_934_new_n170_; 
wire _abc_934_new_n171_; 
wire _abc_934_new_n173_; 
wire _abc_934_new_n174_; 
wire _abc_934_new_n175_; 
wire _abc_934_new_n176_; 
wire _abc_934_new_n178_; 
wire _abc_934_new_n179_; 
wire _abc_934_new_n180_; 
wire _abc_934_new_n181_; 
wire _abc_934_new_n182_; 
wire _abc_934_new_n49_; 
wire _abc_934_new_n50_; 
wire _abc_934_new_n51_; 
wire _abc_934_new_n52_; 
wire _abc_934_new_n53_; 
wire _abc_934_new_n54_; 
wire _abc_934_new_n55_; 
wire _abc_934_new_n56_; 
wire _abc_934_new_n57_; 
wire _abc_934_new_n58_; 
wire _abc_934_new_n59_; 
wire _abc_934_new_n60_; 
wire _abc_934_new_n61_; 
wire _abc_934_new_n62_; 
wire _abc_934_new_n63_; 
wire _abc_934_new_n64_; 
wire _abc_934_new_n65_; 
wire _abc_934_new_n66_; 
wire _abc_934_new_n67_; 
wire _abc_934_new_n68_; 
wire _abc_934_new_n69_; 
wire _abc_934_new_n70_; 
wire _abc_934_new_n71_; 
wire _abc_934_new_n72_; 
wire _abc_934_new_n73_; 
wire _abc_934_new_n74_; 
wire _abc_934_new_n75_; 
wire _abc_934_new_n76_; 
wire _abc_934_new_n77_; 
wire _abc_934_new_n78_; 
wire _abc_934_new_n80_; 
wire _abc_934_new_n81_; 
wire _abc_934_new_n82_; 
wire _abc_934_new_n83_; 
wire _abc_934_new_n84_; 
wire _abc_934_new_n86_; 
wire _abc_934_new_n87_; 
wire _abc_934_new_n88_; 
wire _abc_934_new_n89_; 
wire _abc_934_new_n91_; 
wire _abc_934_new_n92_; 
wire _abc_934_new_n93_; 
wire _abc_934_new_n94_; 
wire _abc_934_new_n95_; 
wire _abc_934_new_n96_; 
wire _abc_934_new_n97_; 
wire _abc_934_new_n98_; 
wire _abc_934_new_n99_; 
wire _auto_iopadmap_cc_368_execute_1071_0_; 
wire _auto_iopadmap_cc_368_execute_1071_1_; 
wire _auto_iopadmap_cc_368_execute_1074; 
wire _auto_iopadmap_cc_368_execute_1076; 
wire _auto_iopadmap_cc_368_execute_1078; 
wire _auto_iopadmap_cc_368_execute_1080; 
wire _auto_iopadmap_cc_368_execute_1082; 
wire _auto_iopadmap_cc_368_execute_1084; 
input aligned_mem;
input busy_mem;
input clk;
input \codif[0] ;
input \codif[10] ;
input \codif[11] ;
input \codif[1] ;
input \codif[2] ;
input \codif[3] ;
input \codif[4] ;
input \codif[5] ;
input \codif[6] ;
input \codif[7] ;
input \codif[8] ;
input \codif[9] ;
input done_exec;
input done_mem;
output en_mem;
output enable_exec;
output enable_exec_mem;
output enable_pc;
wire enable_pc_aux; 
wire enable_pc_fsm; 
input is_exec;
input reset;
output sign_mem;
wire state_0_; 
wire state_1_; 
wire state_2_; 
wire state_3_; 
wire state_4_; 
wire state_5_; 
wire state_6_; 
output trap;
output \wordsize_mem[0] ;
output \wordsize_mem[1] ;
AND2X2 AND2X2_1 ( .A(_abc_934_new_n114_), .B(enable_pc_fsm), .Y(_auto_iopadmap_cc_368_execute_1080));
AND2X2 AND2X2_10 ( .A(_auto_iopadmap_cc_368_execute_1074), .B(done_mem), .Y(_abc_934_new_n134_));
AND2X2 AND2X2_11 ( .A(_abc_934_new_n136_), .B(_abc_934_new_n135_), .Y(_abc_934_new_n137_));
AND2X2 AND2X2_12 ( .A(_abc_934_new_n116_), .B(_abc_934_new_n86_), .Y(_abc_934_new_n139_));
AND2X2 AND2X2_13 ( .A(_abc_934_new_n119_), .B(_abc_934_new_n140_), .Y(_abc_934_new_n141_));
AND2X2 AND2X2_14 ( .A(_abc_934_new_n141_), .B(_abc_934_new_n138_), .Y(_abc_934_new_n142_));
AND2X2 AND2X2_15 ( .A(_abc_934_new_n143_), .B(_auto_iopadmap_cc_368_execute_1071_1_), .Y(_abc_934_new_n144_));
AND2X2 AND2X2_16 ( .A(_abc_934_new_n119_), .B(_abc_934_new_n95_), .Y(_abc_934_new_n145_));
AND2X2 AND2X2_17 ( .A(_abc_934_new_n146_), .B(reset), .Y(_0W_R_mem_1_0__1_));
AND2X2 AND2X2_18 ( .A(_abc_934_new_n150_), .B(_abc_934_new_n151_), .Y(_abc_934_new_n152_));
AND2X2 AND2X2_19 ( .A(_abc_934_new_n153_), .B(enable_pc_fsm), .Y(_abc_934_new_n154_));
AND2X2 AND2X2_2 ( .A(_abc_934_new_n118_), .B(aligned_mem), .Y(_abc_934_new_n119_));
AND2X2 AND2X2_20 ( .A(_abc_934_new_n155_), .B(aligned_mem), .Y(_abc_934_new_n156_));
AND2X2 AND2X2_21 ( .A(_abc_934_new_n157_), .B(reset), .Y(_abc_934_new_n158_));
AND2X2 AND2X2_22 ( .A(_abc_934_new_n158_), .B(_abc_934_new_n149_), .Y(_0enable_pc_fsm_0_0_));
AND2X2 AND2X2_23 ( .A(_abc_934_new_n160_), .B(reset), .Y(_0trap_0_0_));
AND2X2 AND2X2_24 ( .A(_abc_934_new_n106_), .B(_abc_934_new_n125_), .Y(_abc_934_new_n162_));
AND2X2 AND2X2_25 ( .A(_abc_934_new_n163_), .B(_abc_934_new_n86_), .Y(_abc_934_new_n164_));
AND2X2 AND2X2_26 ( .A(_abc_934_new_n165_), .B(_abc_934_new_n166_), .Y(_abc_934_new_n167_));
AND2X2 AND2X2_27 ( .A(reset), .B(_auto_iopadmap_cc_368_execute_1078), .Y(_abc_934_new_n170_));
AND2X2 AND2X2_28 ( .A(_abc_934_new_n169_), .B(_abc_934_new_n170_), .Y(_abc_934_new_n171_));
AND2X2 AND2X2_29 ( .A(_abc_934_new_n153_), .B(_auto_iopadmap_cc_368_execute_1076), .Y(_abc_934_new_n174_));
AND2X2 AND2X2_3 ( .A(_abc_934_new_n120_), .B(_auto_iopadmap_cc_368_execute_1071_0_), .Y(_abc_934_new_n121_));
AND2X2 AND2X2_30 ( .A(_abc_934_new_n175_), .B(reset), .Y(_abc_934_new_n176_));
AND2X2 AND2X2_31 ( .A(_abc_934_new_n176_), .B(_abc_934_new_n173_), .Y(_0enable_exec_0_0_));
AND2X2 AND2X2_32 ( .A(_abc_934_new_n94_), .B(aligned_mem), .Y(_abc_934_new_n178_));
AND2X2 AND2X2_33 ( .A(_abc_934_new_n178_), .B(_abc_934_new_n117_), .Y(_abc_934_new_n179_));
AND2X2 AND2X2_34 ( .A(_abc_934_new_n180_), .B(_auto_iopadmap_cc_368_execute_1074), .Y(_abc_934_new_n181_));
AND2X2 AND2X2_35 ( .A(_abc_934_new_n182_), .B(reset), .Y(_0en_mem_0_0_));
AND2X2 AND2X2_36 ( .A(reset), .B(enable_pc_fsm), .Y(_0enable_pc_aux_0_0_));
AND2X2 AND2X2_37 ( .A(reset), .B(aligned_mem), .Y(_abc_934_new_n49_));
AND2X2 AND2X2_38 ( .A(\codif[0] ), .B(\codif[1] ), .Y(_abc_934_new_n50_));
AND2X2 AND2X2_39 ( .A(_abc_934_new_n56_), .B(state_2_), .Y(_abc_934_new_n57_));
AND2X2 AND2X2_4 ( .A(_abc_934_new_n86_), .B(_auto_iopadmap_cc_368_execute_1071_0_), .Y(_abc_934_new_n122_));
AND2X2 AND2X2_40 ( .A(_abc_934_new_n55_), .B(_abc_934_new_n57_), .Y(_abc_934_new_n58_));
AND2X2 AND2X2_41 ( .A(\codif[4] ), .B(\codif[5] ), .Y(_abc_934_new_n59_));
AND2X2 AND2X2_42 ( .A(\codif[6] ), .B(\codif[7] ), .Y(_abc_934_new_n60_));
AND2X2 AND2X2_43 ( .A(_abc_934_new_n59_), .B(_abc_934_new_n60_), .Y(_abc_934_new_n61_));
AND2X2 AND2X2_44 ( .A(\codif[2] ), .B(\codif[3] ), .Y(_abc_934_new_n62_));
AND2X2 AND2X2_45 ( .A(_abc_934_new_n50_), .B(_abc_934_new_n62_), .Y(_abc_934_new_n63_));
AND2X2 AND2X2_46 ( .A(\codif[10] ), .B(\codif[11] ), .Y(_abc_934_new_n64_));
AND2X2 AND2X2_47 ( .A(\codif[8] ), .B(\codif[9] ), .Y(_abc_934_new_n65_));
AND2X2 AND2X2_48 ( .A(_abc_934_new_n64_), .B(_abc_934_new_n65_), .Y(_abc_934_new_n66_));
AND2X2 AND2X2_49 ( .A(_abc_934_new_n63_), .B(_abc_934_new_n66_), .Y(_abc_934_new_n67_));
AND2X2 AND2X2_5 ( .A(_abc_934_new_n122_), .B(_abc_934_new_n116_), .Y(_abc_934_new_n123_));
AND2X2 AND2X2_50 ( .A(_abc_934_new_n67_), .B(_abc_934_new_n61_), .Y(_abc_934_new_n68_));
AND2X2 AND2X2_51 ( .A(_abc_934_new_n75_), .B(_abc_934_new_n69_), .Y(_abc_934_new_n76_));
AND2X2 AND2X2_52 ( .A(_abc_934_new_n76_), .B(state_4_), .Y(_abc_934_new_n77_));
AND2X2 AND2X2_53 ( .A(_abc_934_new_n78_), .B(_abc_934_new_n49_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_2_));
AND2X2 AND2X2_54 ( .A(_abc_934_new_n82_), .B(state_4_), .Y(_abc_934_new_n83_));
AND2X2 AND2X2_55 ( .A(_abc_934_new_n84_), .B(reset), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_1_));
AND2X2 AND2X2_56 ( .A(_abc_934_new_n49_), .B(_abc_934_new_n86_), .Y(_abc_934_new_n87_));
AND2X2 AND2X2_57 ( .A(state_6_), .B(_auto_iopadmap_cc_368_execute_1074), .Y(_abc_934_new_n88_));
AND2X2 AND2X2_58 ( .A(_abc_934_new_n89_), .B(_abc_934_new_n87_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_3_));
AND2X2 AND2X2_59 ( .A(_abc_934_new_n49_), .B(state_2_), .Y(_abc_934_new_n91_));
AND2X2 AND2X2_6 ( .A(_abc_934_new_n126_), .B(state_6_), .Y(_abc_934_new_n127_));
AND2X2 AND2X2_60 ( .A(_abc_934_new_n91_), .B(done_exec), .Y(_abc_934_new_n92_));
AND2X2 AND2X2_61 ( .A(_abc_934_new_n55_), .B(_abc_934_new_n92_), .Y(_abc_934_new_n93_));
AND2X2 AND2X2_62 ( .A(_abc_934_new_n94_), .B(state_0_), .Y(_abc_934_new_n95_));
AND2X2 AND2X2_63 ( .A(_abc_934_new_n88_), .B(done_mem), .Y(_abc_934_new_n96_));
AND2X2 AND2X2_64 ( .A(_abc_934_new_n97_), .B(aligned_mem), .Y(_abc_934_new_n98_));
AND2X2 AND2X2_65 ( .A(_abc_934_new_n49_), .B(done_mem), .Y(_abc_934_new_n100_));
AND2X2 AND2X2_66 ( .A(_abc_934_new_n100_), .B(state_3_), .Y(_abc_934_new_n101_));
AND2X2 AND2X2_67 ( .A(_abc_934_new_n94_), .B(state_6_), .Y(_abc_934_new_n105_));
AND2X2 AND2X2_68 ( .A(_abc_934_new_n105_), .B(_abc_934_new_n49_), .Y(_abc_934_new_n106_));
AND2X2 AND2X2_69 ( .A(_abc_934_new_n107_), .B(_abc_934_new_n91_), .Y(_abc_934_new_n108_));
AND2X2 AND2X2_7 ( .A(_abc_934_new_n128_), .B(_abc_934_new_n124_), .Y(_abc_934_new_n129_));
AND2X2 AND2X2_70 ( .A(_auto_iopadmap_cc_368_execute_1074), .B(state_0_), .Y(_abc_934_new_n110_));
AND2X2 AND2X2_71 ( .A(_abc_934_new_n111_), .B(_abc_934_new_n100_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_4_));
AND2X2 AND2X2_72 ( .A(_abc_934_new_n111_), .B(_abc_934_new_n87_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_5_));
AND2X2 AND2X2_8 ( .A(_abc_934_new_n130_), .B(aligned_mem), .Y(_abc_934_new_n131_));
AND2X2 AND2X2_9 ( .A(_abc_934_new_n132_), .B(reset), .Y(_0W_R_mem_1_0__0_));
BUFX2 BUFX2_1 ( .A(_auto_iopadmap_cc_368_execute_1071_0_), .Y(\W_R_mem[0] ));
BUFX2 BUFX2_10 ( .A(\codif[8] ), .Y(\wordsize_mem[1] ));
BUFX2 BUFX2_2 ( .A(_auto_iopadmap_cc_368_execute_1071_1_), .Y(\W_R_mem[1] ));
BUFX2 BUFX2_3 ( .A(_auto_iopadmap_cc_368_execute_1074), .Y(en_mem));
BUFX2 BUFX2_4 ( .A(_auto_iopadmap_cc_368_execute_1076), .Y(enable_exec));
BUFX2 BUFX2_5 ( .A(_auto_iopadmap_cc_368_execute_1078), .Y(enable_exec_mem));
BUFX2 BUFX2_6 ( .A(_auto_iopadmap_cc_368_execute_1080), .Y(enable_pc));
BUFX2 BUFX2_7 ( .A(_auto_iopadmap_cc_368_execute_1082), .Y(sign_mem));
BUFX2 BUFX2_8 ( .A(_auto_iopadmap_cc_368_execute_1084), .Y(trap));
BUFX2 BUFX2_9 ( .A(\codif[7] ), .Y(\wordsize_mem[0] ));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_0_), .Q(state_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(_0en_mem_0_0_), .Q(_auto_iopadmap_cc_368_execute_1074));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(_0enable_exec_0_0_), .Q(_auto_iopadmap_cc_368_execute_1076));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(_0enable_exec_mem_0_0_), .Q(_auto_iopadmap_cc_368_execute_1078));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(_0trap_0_0_), .Q(_auto_iopadmap_cc_368_execute_1084));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(_0enable_pc_fsm_0_0_), .Q(enable_pc_fsm));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(_0enable_pc_aux_0_0_), .Q(enable_pc_aux));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_1_), .Q(state_1_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_2_), .Q(state_2_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_3_), .Q(state_3_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_4_), .Q(state_4_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_5_), .Q(state_5_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(_abc_801_auto_fsm_map_cc_170_map_fsm_238_6_), .Q(state_6_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(_0W_R_mem_1_0__0_), .Q(_auto_iopadmap_cc_368_execute_1071_0_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(_0W_R_mem_1_0__1_), .Q(_auto_iopadmap_cc_368_execute_1071_1_));
INVX1 INVX1_1 ( .A(enable_pc_aux), .Y(_abc_934_new_n114_));
INVX1 INVX1_10 ( .A(state_4_), .Y(_abc_934_new_n151_));
INVX1 INVX1_11 ( .A(state_3_), .Y(_abc_934_new_n165_));
INVX1 INVX1_12 ( .A(state_6_), .Y(_abc_934_new_n166_));
INVX1 INVX1_13 ( .A(_abc_934_new_n141_), .Y(_abc_934_new_n180_));
INVX1 INVX1_14 ( .A(_abc_934_new_n50_), .Y(_abc_934_new_n51_));
INVX1 INVX1_15 ( .A(done_exec), .Y(_abc_934_new_n56_));
INVX1 INVX1_16 ( .A(_abc_934_new_n68_), .Y(_abc_934_new_n69_));
INVX1 INVX1_17 ( .A(_abc_934_new_n61_), .Y(_abc_934_new_n73_));
INVX1 INVX1_18 ( .A(aligned_mem), .Y(_abc_934_new_n80_));
INVX1 INVX1_19 ( .A(_abc_934_new_n76_), .Y(_abc_934_new_n82_));
INVX1 INVX1_2 ( .A(_abc_934_new_n119_), .Y(_abc_934_new_n120_));
INVX1 INVX1_20 ( .A(done_mem), .Y(_abc_934_new_n86_));
INVX1 INVX1_21 ( .A(_auto_iopadmap_cc_368_execute_1074), .Y(_abc_934_new_n94_));
INVX1 INVX1_22 ( .A(reset), .Y(_abc_934_new_n99_));
INVX1 INVX1_23 ( .A(_abc_934_new_n55_), .Y(_abc_934_new_n107_));
INVX1 INVX1_3 ( .A(\codif[5] ), .Y(_abc_934_new_n125_));
INVX1 INVX1_4 ( .A(state_0_), .Y(_abc_934_new_n135_));
INVX1 INVX1_5 ( .A(_abc_934_new_n88_), .Y(_abc_934_new_n136_));
INVX1 INVX1_6 ( .A(_abc_934_new_n139_), .Y(_abc_934_new_n140_));
INVX1 INVX1_7 ( .A(_abc_934_new_n142_), .Y(_abc_934_new_n143_));
INVX1 INVX1_8 ( .A(\codif[9] ), .Y(_auto_iopadmap_cc_368_execute_1082));
INVX1 INVX1_9 ( .A(state_2_), .Y(_abc_934_new_n150_));
OR2X2 OR2X2_1 ( .A(state_3_), .B(state_5_), .Y(_abc_934_new_n116_));
OR2X2 OR2X2_10 ( .A(_abc_934_new_n144_), .B(_abc_934_new_n145_), .Y(_abc_934_new_n146_));
OR2X2 OR2X2_11 ( .A(_abc_934_new_n77_), .B(enable_pc_fsm), .Y(_abc_934_new_n149_));
OR2X2 OR2X2_12 ( .A(_abc_934_new_n152_), .B(_abc_934_new_n80_), .Y(_abc_934_new_n153_));
OR2X2 OR2X2_13 ( .A(_abc_934_new_n58_), .B(state_4_), .Y(_abc_934_new_n155_));
OR2X2 OR2X2_14 ( .A(_abc_934_new_n156_), .B(_abc_934_new_n154_), .Y(_abc_934_new_n157_));
OR2X2 OR2X2_15 ( .A(_abc_934_new_n81_), .B(_auto_iopadmap_cc_368_execute_1084), .Y(_abc_934_new_n160_));
OR2X2 OR2X2_16 ( .A(_abc_934_new_n127_), .B(state_3_), .Y(_abc_934_new_n163_));
OR2X2 OR2X2_17 ( .A(_abc_934_new_n167_), .B(_abc_934_new_n80_), .Y(_abc_934_new_n168_));
OR2X2 OR2X2_18 ( .A(_abc_934_new_n164_), .B(_abc_934_new_n168_), .Y(_abc_934_new_n169_));
OR2X2 OR2X2_19 ( .A(_abc_934_new_n171_), .B(_abc_934_new_n162_), .Y(_0enable_exec_mem_0_0_));
OR2X2 OR2X2_2 ( .A(state_6_), .B(state_0_), .Y(_abc_934_new_n117_));
OR2X2 OR2X2_20 ( .A(_abc_934_new_n77_), .B(_auto_iopadmap_cc_368_execute_1076), .Y(_abc_934_new_n173_));
OR2X2 OR2X2_21 ( .A(_abc_934_new_n156_), .B(_abc_934_new_n174_), .Y(_abc_934_new_n175_));
OR2X2 OR2X2_22 ( .A(_abc_934_new_n181_), .B(_abc_934_new_n179_), .Y(_abc_934_new_n182_));
OR2X2 OR2X2_23 ( .A(\codif[2] ), .B(\codif[3] ), .Y(_abc_934_new_n52_));
OR2X2 OR2X2_24 ( .A(_abc_934_new_n51_), .B(_abc_934_new_n52_), .Y(_abc_934_new_n53_));
OR2X2 OR2X2_25 ( .A(\codif[4] ), .B(\codif[6] ), .Y(_abc_934_new_n54_));
OR2X2 OR2X2_26 ( .A(_abc_934_new_n53_), .B(_abc_934_new_n54_), .Y(_abc_934_new_n55_));
OR2X2 OR2X2_27 ( .A(\codif[10] ), .B(\codif[11] ), .Y(_abc_934_new_n70_));
OR2X2 OR2X2_28 ( .A(\codif[8] ), .B(\codif[9] ), .Y(_abc_934_new_n71_));
OR2X2 OR2X2_29 ( .A(_abc_934_new_n70_), .B(_abc_934_new_n71_), .Y(_abc_934_new_n72_));
OR2X2 OR2X2_3 ( .A(_abc_934_new_n116_), .B(_abc_934_new_n117_), .Y(_abc_934_new_n118_));
OR2X2 OR2X2_30 ( .A(_abc_934_new_n53_), .B(_abc_934_new_n73_), .Y(_abc_934_new_n74_));
OR2X2 OR2X2_31 ( .A(_abc_934_new_n74_), .B(_abc_934_new_n72_), .Y(_abc_934_new_n75_));
OR2X2 OR2X2_32 ( .A(_abc_934_new_n77_), .B(_abc_934_new_n58_), .Y(_abc_934_new_n78_));
OR2X2 OR2X2_33 ( .A(_abc_934_new_n80_), .B(state_1_), .Y(_abc_934_new_n81_));
OR2X2 OR2X2_34 ( .A(_abc_934_new_n83_), .B(_abc_934_new_n81_), .Y(_abc_934_new_n84_));
OR2X2 OR2X2_35 ( .A(_abc_934_new_n88_), .B(state_3_), .Y(_abc_934_new_n89_));
OR2X2 OR2X2_36 ( .A(_abc_934_new_n96_), .B(_abc_934_new_n95_), .Y(_abc_934_new_n97_));
OR2X2 OR2X2_37 ( .A(_abc_934_new_n101_), .B(_abc_934_new_n99_), .Y(_abc_934_new_n102_));
OR2X2 OR2X2_38 ( .A(_abc_934_new_n98_), .B(_abc_934_new_n102_), .Y(_abc_934_new_n103_));
OR2X2 OR2X2_39 ( .A(_abc_934_new_n103_), .B(_abc_934_new_n93_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_0_));
OR2X2 OR2X2_4 ( .A(_abc_934_new_n122_), .B(_abc_934_new_n94_), .Y(_abc_934_new_n124_));
OR2X2 OR2X2_40 ( .A(_abc_934_new_n108_), .B(_abc_934_new_n106_), .Y(_abc_801_auto_fsm_map_cc_170_map_fsm_238_6_));
OR2X2 OR2X2_41 ( .A(_abc_934_new_n110_), .B(state_5_), .Y(_abc_934_new_n111_));
OR2X2 OR2X2_5 ( .A(_abc_934_new_n125_), .B(_auto_iopadmap_cc_368_execute_1074), .Y(_abc_934_new_n126_));
OR2X2 OR2X2_6 ( .A(_abc_934_new_n127_), .B(state_0_), .Y(_abc_934_new_n128_));
OR2X2 OR2X2_7 ( .A(_abc_934_new_n129_), .B(_abc_934_new_n123_), .Y(_abc_934_new_n130_));
OR2X2 OR2X2_8 ( .A(_abc_934_new_n131_), .B(_abc_934_new_n121_), .Y(_abc_934_new_n132_));
OR2X2 OR2X2_9 ( .A(_abc_934_new_n137_), .B(_abc_934_new_n134_), .Y(_abc_934_new_n138_));


endmodule