module b09_reset(clock, RESET_G, nRESET_G, X, Y_REG);

wire D_IN_REG_0_; 
wire D_IN_REG_1_; 
wire D_IN_REG_2_; 
wire D_IN_REG_3_; 
wire D_IN_REG_4_; 
wire D_IN_REG_5_; 
wire D_IN_REG_6_; 
wire D_IN_REG_7_; 
wire D_IN_REG_8_; 
wire D_OUT_REG_0_; 
wire D_OUT_REG_1_; 
wire D_OUT_REG_2_; 
wire D_OUT_REG_3_; 
wire D_OUT_REG_4_; 
wire D_OUT_REG_5_; 
wire D_OUT_REG_6_; 
wire D_OUT_REG_7_; 
wire OLD_REG_0_; 
wire OLD_REG_1_; 
wire OLD_REG_2_; 
wire OLD_REG_3_; 
wire OLD_REG_4_; 
wire OLD_REG_5_; 
wire OLD_REG_6_; 
wire OLD_REG_7_; 
input RESET_G;
wire STATO_REG_0_; 
wire STATO_REG_1_; 
input X;
output Y_REG;
wire _abc_898_new_n100_; 
wire _abc_898_new_n102_; 
wire _abc_898_new_n104_; 
wire _abc_898_new_n106_; 
wire _abc_898_new_n108_; 
wire _abc_898_new_n110_; 
wire _abc_898_new_n112_; 
wire _abc_898_new_n114_; 
wire _abc_898_new_n115_; 
wire _abc_898_new_n116_; 
wire _abc_898_new_n117_; 
wire _abc_898_new_n118_; 
wire _abc_898_new_n119_; 
wire _abc_898_new_n120_; 
wire _abc_898_new_n121_; 
wire _abc_898_new_n122_; 
wire _abc_898_new_n123_; 
wire _abc_898_new_n124_; 
wire _abc_898_new_n125_; 
wire _abc_898_new_n126_; 
wire _abc_898_new_n127_; 
wire _abc_898_new_n128_; 
wire _abc_898_new_n129_; 
wire _abc_898_new_n130_; 
wire _abc_898_new_n132_; 
wire _abc_898_new_n133_; 
wire _abc_898_new_n135_; 
wire _abc_898_new_n136_; 
wire _abc_898_new_n138_; 
wire _abc_898_new_n139_; 
wire _abc_898_new_n141_; 
wire _abc_898_new_n142_; 
wire _abc_898_new_n144_; 
wire _abc_898_new_n145_; 
wire _abc_898_new_n147_; 
wire _abc_898_new_n148_; 
wire _abc_898_new_n150_; 
wire _abc_898_new_n151_; 
wire _abc_898_new_n153_; 
wire _abc_898_new_n154_; 
wire _abc_898_new_n156_; 
wire _abc_898_new_n157_; 
wire _abc_898_new_n158_; 
wire _abc_898_new_n159_; 
wire _abc_898_new_n160_; 
wire _abc_898_new_n161_; 
wire _abc_898_new_n162_; 
wire _abc_898_new_n164_; 
wire _abc_898_new_n165_; 
wire _abc_898_new_n166_; 
wire _abc_898_new_n167_; 
wire _abc_898_new_n168_; 
wire _abc_898_new_n170_; 
wire _abc_898_new_n171_; 
wire _abc_898_new_n172_; 
wire _abc_898_new_n173_; 
wire _abc_898_new_n174_; 
wire _abc_898_new_n176_; 
wire _abc_898_new_n177_; 
wire _abc_898_new_n178_; 
wire _abc_898_new_n179_; 
wire _abc_898_new_n180_; 
wire _abc_898_new_n182_; 
wire _abc_898_new_n183_; 
wire _abc_898_new_n184_; 
wire _abc_898_new_n185_; 
wire _abc_898_new_n186_; 
wire _abc_898_new_n188_; 
wire _abc_898_new_n189_; 
wire _abc_898_new_n190_; 
wire _abc_898_new_n191_; 
wire _abc_898_new_n192_; 
wire _abc_898_new_n194_; 
wire _abc_898_new_n195_; 
wire _abc_898_new_n196_; 
wire _abc_898_new_n198_; 
wire _abc_898_new_n199_; 
wire _abc_898_new_n200_; 
wire _abc_898_new_n201_; 
wire _abc_898_new_n202_; 
wire _abc_898_new_n59_; 
wire _abc_898_new_n60_; 
wire _abc_898_new_n61_; 
wire _abc_898_new_n62_; 
wire _abc_898_new_n64_; 
wire _abc_898_new_n65_; 
wire _abc_898_new_n66_; 
wire _abc_898_new_n67_; 
wire _abc_898_new_n68_; 
wire _abc_898_new_n69_; 
wire _abc_898_new_n70_; 
wire _abc_898_new_n71_; 
wire _abc_898_new_n72_; 
wire _abc_898_new_n73_; 
wire _abc_898_new_n74_; 
wire _abc_898_new_n75_; 
wire _abc_898_new_n76_; 
wire _abc_898_new_n77_; 
wire _abc_898_new_n78_; 
wire _abc_898_new_n79_; 
wire _abc_898_new_n80_; 
wire _abc_898_new_n81_; 
wire _abc_898_new_n82_; 
wire _abc_898_new_n83_; 
wire _abc_898_new_n84_; 
wire _abc_898_new_n85_; 
wire _abc_898_new_n86_; 
wire _abc_898_new_n87_; 
wire _abc_898_new_n89_; 
wire _abc_898_new_n90_; 
wire _abc_898_new_n91_; 
wire _abc_898_new_n92_; 
wire _abc_898_new_n93_; 
wire _abc_898_new_n94_; 
wire _abc_898_new_n96_; 
wire _abc_898_new_n97_; 
wire _abc_898_new_n98_; 
wire _auto_iopadmap_cc_368_execute_1044; 
input clock;
wire clock_bF_buf0; 
wire clock_bF_buf1; 
wire clock_bF_buf2; 
wire clock_bF_buf3; 
wire clock_bF_buf4; 
wire n10; 
wire n104; 
wire n109; 
wire n114; 
wire n119; 
wire n124; 
wire n129; 
wire n134; 
wire n139; 
wire n144; 
wire n15; 
wire n20; 
wire n25; 
wire n30; 
wire n35; 
wire n40; 
wire n45; 
wire n50; 
wire n55; 
wire n60; 
wire n65; 
wire n70; 
wire n75; 
wire n80; 
wire n85; 
wire n90; 
wire n95; 
wire n99; 
input nRESET_G;
wire nRESET_G_bF_buf0; 
wire nRESET_G_bF_buf1; 
wire nRESET_G_bF_buf2; 
wire nRESET_G_bF_buf3; 
AOI21X1 AOI21X1_1 ( .A(_abc_898_new_n93_), .B(_abc_898_new_n158_), .C(_abc_898_new_n161_), .Y(_abc_898_new_n162_));
AOI21X1 AOI21X1_10 ( .A(_abc_898_new_n93_), .B(_abc_898_new_n92_), .C(_abc_898_new_n61_), .Y(_abc_898_new_n94_));
AOI21X1 AOI21X1_11 ( .A(_abc_898_new_n60_), .B(_abc_898_new_n82_), .C(_abc_898_new_n92_), .Y(_abc_898_new_n97_));
AOI21X1 AOI21X1_12 ( .A(D_OUT_REG_0_), .B(_abc_898_new_n127_), .C(_abc_898_new_n129_), .Y(_abc_898_new_n130_));
AOI21X1 AOI21X1_2 ( .A(_abc_898_new_n93_), .B(_abc_898_new_n165_), .C(_abc_898_new_n167_), .Y(_abc_898_new_n168_));
AOI21X1 AOI21X1_3 ( .A(_abc_898_new_n93_), .B(_abc_898_new_n171_), .C(_abc_898_new_n173_), .Y(_abc_898_new_n174_));
AOI21X1 AOI21X1_4 ( .A(_abc_898_new_n93_), .B(_abc_898_new_n177_), .C(_abc_898_new_n179_), .Y(_abc_898_new_n180_));
AOI21X1 AOI21X1_5 ( .A(_abc_898_new_n93_), .B(_abc_898_new_n183_), .C(_abc_898_new_n185_), .Y(_abc_898_new_n186_));
AOI21X1 AOI21X1_6 ( .A(_abc_898_new_n93_), .B(_abc_898_new_n189_), .C(_abc_898_new_n191_), .Y(_abc_898_new_n192_));
AOI21X1 AOI21X1_7 ( .A(_abc_898_new_n93_), .B(_abc_898_new_n195_), .C(_abc_898_new_n61_), .Y(_abc_898_new_n196_));
AOI21X1 AOI21X1_8 ( .A(_abc_898_new_n93_), .B(_abc_898_new_n199_), .C(_abc_898_new_n201_), .Y(_abc_898_new_n202_));
AOI21X1 AOI21X1_9 ( .A(_abc_898_new_n86_), .B(_abc_898_new_n60_), .C(_abc_898_new_n61_), .Y(_abc_898_new_n87_));
AOI22X1 AOI22X1_1 ( .A(_abc_898_new_n121_), .B(_abc_898_new_n74_), .C(_abc_898_new_n77_), .D(_abc_898_new_n122_), .Y(_abc_898_new_n123_));
BUFX2 BUFX2_1 ( .A(nRESET_G), .Y(nRESET_G_bF_buf3));
BUFX2 BUFX2_2 ( .A(nRESET_G), .Y(nRESET_G_bF_buf2));
BUFX2 BUFX2_3 ( .A(nRESET_G), .Y(nRESET_G_bF_buf1));
BUFX2 BUFX2_4 ( .A(nRESET_G), .Y(nRESET_G_bF_buf0));
BUFX2 BUFX2_5 ( .A(_auto_iopadmap_cc_368_execute_1044), .Y(Y_REG));
BUFX4 BUFX4_1 ( .A(clock), .Y(clock_bF_buf4));
BUFX4 BUFX4_2 ( .A(clock), .Y(clock_bF_buf3));
BUFX4 BUFX4_3 ( .A(clock), .Y(clock_bF_buf2));
BUFX4 BUFX4_4 ( .A(clock), .Y(clock_bF_buf1));
BUFX4 BUFX4_5 ( .A(clock), .Y(clock_bF_buf0));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock_bF_buf4), .D(n25), .Q(D_OUT_REG_5_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock_bF_buf0), .D(n50), .Q(D_OUT_REG_0_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock_bF_buf4), .D(n55), .Q(OLD_REG_7_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock_bF_buf3), .D(n60), .Q(OLD_REG_6_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock_bF_buf2), .D(n65), .Q(OLD_REG_5_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock_bF_buf1), .D(n70), .Q(OLD_REG_4_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock_bF_buf0), .D(n75), .Q(OLD_REG_3_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock_bF_buf4), .D(n80), .Q(OLD_REG_2_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock_bF_buf3), .D(n85), .Q(OLD_REG_1_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock_bF_buf2), .D(n90), .Q(OLD_REG_0_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock_bF_buf1), .D(n99), .Q(STATO_REG_1_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock_bF_buf3), .D(n15), .Q(D_OUT_REG_7_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock_bF_buf0), .D(n104), .Q(STATO_REG_0_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock_bF_buf4), .D(n109), .Q(D_IN_REG_8_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock_bF_buf3), .D(n114), .Q(D_IN_REG_7_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock_bF_buf2), .D(n119), .Q(D_IN_REG_6_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock_bF_buf1), .D(n124), .Q(D_IN_REG_5_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock_bF_buf0), .D(n129), .Q(D_IN_REG_4_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock_bF_buf4), .D(n134), .Q(D_IN_REG_3_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock_bF_buf3), .D(n139), .Q(D_IN_REG_2_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock_bF_buf2), .D(n144), .Q(D_IN_REG_1_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock_bF_buf2), .D(n10), .Q(D_IN_REG_0_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock_bF_buf1), .D(n20), .Q(D_OUT_REG_6_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock_bF_buf0), .D(n95), .Q(_auto_iopadmap_cc_368_execute_1044));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock_bF_buf4), .D(n30), .Q(D_OUT_REG_4_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock_bF_buf3), .D(n35), .Q(D_OUT_REG_3_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock_bF_buf2), .D(n40), .Q(D_OUT_REG_2_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock_bF_buf1), .D(n45), .Q(D_OUT_REG_1_));
INVX1 INVX1_1 ( .A(_abc_898_new_n136_), .Y(_abc_898_new_n165_));
INVX1 INVX1_10 ( .A(D_OUT_REG_6_), .Y(_abc_898_new_n190_));
INVX1 INVX1_11 ( .A(_abc_898_new_n154_), .Y(_abc_898_new_n195_));
INVX1 INVX1_12 ( .A(_abc_898_new_n151_), .Y(_abc_898_new_n199_));
INVX1 INVX1_13 ( .A(D_OUT_REG_7_), .Y(_abc_898_new_n200_));
INVX1 INVX1_14 ( .A(D_IN_REG_0_), .Y(_abc_898_new_n59_));
INVX1 INVX1_15 ( .A(_abc_898_new_n74_), .Y(_abc_898_new_n75_));
INVX1 INVX1_16 ( .A(_abc_898_new_n77_), .Y(_abc_898_new_n78_));
INVX1 INVX1_17 ( .A(D_IN_REG_1_), .Y(_abc_898_new_n96_));
INVX1 INVX1_18 ( .A(D_IN_REG_2_), .Y(_abc_898_new_n100_));
INVX1 INVX1_19 ( .A(D_IN_REG_3_), .Y(_abc_898_new_n102_));
INVX1 INVX1_2 ( .A(D_OUT_REG_2_), .Y(_abc_898_new_n166_));
INVX1 INVX1_20 ( .A(D_IN_REG_4_), .Y(_abc_898_new_n104_));
INVX1 INVX1_21 ( .A(D_IN_REG_5_), .Y(_abc_898_new_n106_));
INVX1 INVX1_22 ( .A(D_IN_REG_6_), .Y(_abc_898_new_n108_));
INVX1 INVX1_23 ( .A(D_IN_REG_7_), .Y(_abc_898_new_n110_));
INVX1 INVX1_24 ( .A(D_IN_REG_8_), .Y(_abc_898_new_n112_));
INVX1 INVX1_25 ( .A(_abc_898_new_n76_), .Y(_abc_898_new_n121_));
INVX1 INVX1_26 ( .A(_abc_898_new_n79_), .Y(_abc_898_new_n122_));
INVX1 INVX1_27 ( .A(_abc_898_new_n133_), .Y(_abc_898_new_n158_));
INVX1 INVX1_28 ( .A(D_OUT_REG_1_), .Y(_abc_898_new_n159_));
INVX1 INVX1_3 ( .A(_abc_898_new_n139_), .Y(_abc_898_new_n171_));
INVX1 INVX1_4 ( .A(D_OUT_REG_3_), .Y(_abc_898_new_n172_));
INVX1 INVX1_5 ( .A(_abc_898_new_n142_), .Y(_abc_898_new_n177_));
INVX1 INVX1_6 ( .A(D_OUT_REG_4_), .Y(_abc_898_new_n178_));
INVX1 INVX1_7 ( .A(_abc_898_new_n145_), .Y(_abc_898_new_n183_));
INVX1 INVX1_8 ( .A(D_OUT_REG_5_), .Y(_abc_898_new_n184_));
INVX1 INVX1_9 ( .A(_abc_898_new_n148_), .Y(_abc_898_new_n189_));
INVX2 INVX2_1 ( .A(nRESET_G_bF_buf0), .Y(_abc_898_new_n61_));
INVX2 INVX2_2 ( .A(STATO_REG_1_), .Y(_abc_898_new_n82_));
INVX4 INVX4_1 ( .A(_abc_898_new_n127_), .Y(_abc_898_new_n160_));
INVX4 INVX4_2 ( .A(STATO_REG_0_), .Y(_abc_898_new_n60_));
MUX2X1 MUX2X1_1 ( .A(_abc_898_new_n82_), .B(_abc_898_new_n60_), .S(D_IN_REG_0_), .Y(_abc_898_new_n156_));
NAND2X1 NAND2X1_1 ( .A(_abc_898_new_n157_), .B(_abc_898_new_n162_), .Y(n50));
NAND2X1 NAND2X1_10 ( .A(_abc_898_new_n67_), .B(_abc_898_new_n68_), .Y(_abc_898_new_n69_));
NAND2X1 NAND2X1_11 ( .A(_abc_898_new_n71_), .B(_abc_898_new_n72_), .Y(_abc_898_new_n73_));
NAND2X1 NAND2X1_12 ( .A(OLD_REG_0_), .B(D_IN_REG_1_), .Y(_abc_898_new_n74_));
NAND2X1 NAND2X1_13 ( .A(OLD_REG_1_), .B(D_IN_REG_2_), .Y(_abc_898_new_n77_));
NAND2X1 NAND2X1_14 ( .A(STATO_REG_0_), .B(_abc_898_new_n59_), .Y(_abc_898_new_n85_));
NAND2X1 NAND2X1_15 ( .A(STATO_REG_1_), .B(_abc_898_new_n59_), .Y(_abc_898_new_n86_));
NAND2X1 NAND2X1_16 ( .A(_abc_898_new_n91_), .B(_abc_898_new_n94_), .Y(n109));
NAND2X1 NAND2X1_17 ( .A(nRESET_G_bF_buf3), .B(_abc_898_new_n97_), .Y(_abc_898_new_n98_));
NAND2X1 NAND2X1_18 ( .A(_abc_898_new_n116_), .B(_abc_898_new_n119_), .Y(_abc_898_new_n120_));
NAND2X1 NAND2X1_19 ( .A(STATO_REG_1_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n126_));
NAND2X1 NAND2X1_2 ( .A(_abc_898_new_n164_), .B(_abc_898_new_n168_), .Y(n45));
NAND2X1 NAND2X1_20 ( .A(nRESET_G_bF_buf2), .B(_abc_898_new_n128_), .Y(_abc_898_new_n129_));
NAND2X1 NAND2X1_21 ( .A(_abc_898_new_n130_), .B(_abc_898_new_n125_), .Y(n95));
NAND2X1 NAND2X1_22 ( .A(OLD_REG_0_), .B(_abc_898_new_n97_), .Y(_abc_898_new_n132_));
NAND2X1 NAND2X1_23 ( .A(D_IN_REG_1_), .B(_abc_898_new_n92_), .Y(_abc_898_new_n133_));
NAND2X1 NAND2X1_24 ( .A(OLD_REG_1_), .B(_abc_898_new_n97_), .Y(_abc_898_new_n135_));
NAND2X1 NAND2X1_25 ( .A(D_IN_REG_2_), .B(_abc_898_new_n92_), .Y(_abc_898_new_n136_));
NAND2X1 NAND2X1_26 ( .A(OLD_REG_2_), .B(_abc_898_new_n97_), .Y(_abc_898_new_n138_));
NAND2X1 NAND2X1_27 ( .A(D_IN_REG_3_), .B(_abc_898_new_n92_), .Y(_abc_898_new_n139_));
NAND2X1 NAND2X1_28 ( .A(OLD_REG_3_), .B(_abc_898_new_n97_), .Y(_abc_898_new_n141_));
NAND2X1 NAND2X1_29 ( .A(D_IN_REG_4_), .B(_abc_898_new_n92_), .Y(_abc_898_new_n142_));
NAND2X1 NAND2X1_3 ( .A(_abc_898_new_n170_), .B(_abc_898_new_n174_), .Y(n40));
NAND2X1 NAND2X1_30 ( .A(OLD_REG_4_), .B(_abc_898_new_n97_), .Y(_abc_898_new_n144_));
NAND2X1 NAND2X1_31 ( .A(D_IN_REG_5_), .B(_abc_898_new_n92_), .Y(_abc_898_new_n145_));
NAND2X1 NAND2X1_32 ( .A(OLD_REG_5_), .B(_abc_898_new_n97_), .Y(_abc_898_new_n147_));
NAND2X1 NAND2X1_33 ( .A(D_IN_REG_6_), .B(_abc_898_new_n92_), .Y(_abc_898_new_n148_));
NAND2X1 NAND2X1_34 ( .A(OLD_REG_6_), .B(_abc_898_new_n97_), .Y(_abc_898_new_n150_));
NAND2X1 NAND2X1_35 ( .A(D_IN_REG_7_), .B(_abc_898_new_n92_), .Y(_abc_898_new_n151_));
NAND2X1 NAND2X1_36 ( .A(OLD_REG_7_), .B(_abc_898_new_n97_), .Y(_abc_898_new_n153_));
NAND2X1 NAND2X1_37 ( .A(D_IN_REG_8_), .B(_abc_898_new_n92_), .Y(_abc_898_new_n154_));
NAND2X1 NAND2X1_4 ( .A(_abc_898_new_n176_), .B(_abc_898_new_n180_), .Y(n35));
NAND2X1 NAND2X1_5 ( .A(_abc_898_new_n182_), .B(_abc_898_new_n186_), .Y(n30));
NAND2X1 NAND2X1_6 ( .A(_abc_898_new_n188_), .B(_abc_898_new_n192_), .Y(n25));
NAND2X1 NAND2X1_7 ( .A(_abc_898_new_n194_), .B(_abc_898_new_n196_), .Y(n15));
NAND2X1 NAND2X1_8 ( .A(_abc_898_new_n198_), .B(_abc_898_new_n202_), .Y(n20));
NAND2X1 NAND2X1_9 ( .A(_abc_898_new_n64_), .B(_abc_898_new_n65_), .Y(_abc_898_new_n66_));
NAND3X1 NAND3X1_1 ( .A(D_OUT_REG_1_), .B(_abc_898_new_n156_), .C(_abc_898_new_n125_), .Y(_abc_898_new_n164_));
NAND3X1 NAND3X1_10 ( .A(STATO_REG_1_), .B(_abc_898_new_n81_), .C(_abc_898_new_n70_), .Y(_abc_898_new_n93_));
NAND3X1 NAND3X1_11 ( .A(_abc_898_new_n71_), .B(_abc_898_new_n72_), .C(_abc_898_new_n123_), .Y(_abc_898_new_n124_));
NAND3X1 NAND3X1_12 ( .A(nRESET_G_bF_buf1), .B(_abc_898_new_n133_), .C(_abc_898_new_n132_), .Y(n90));
NAND3X1 NAND3X1_13 ( .A(nRESET_G_bF_buf0), .B(_abc_898_new_n136_), .C(_abc_898_new_n135_), .Y(n85));
NAND3X1 NAND3X1_14 ( .A(nRESET_G_bF_buf3), .B(_abc_898_new_n139_), .C(_abc_898_new_n138_), .Y(n80));
NAND3X1 NAND3X1_15 ( .A(nRESET_G_bF_buf2), .B(_abc_898_new_n142_), .C(_abc_898_new_n141_), .Y(n75));
NAND3X1 NAND3X1_16 ( .A(nRESET_G_bF_buf1), .B(_abc_898_new_n145_), .C(_abc_898_new_n144_), .Y(n70));
NAND3X1 NAND3X1_17 ( .A(nRESET_G_bF_buf0), .B(_abc_898_new_n148_), .C(_abc_898_new_n147_), .Y(n65));
NAND3X1 NAND3X1_18 ( .A(nRESET_G_bF_buf3), .B(_abc_898_new_n151_), .C(_abc_898_new_n150_), .Y(n60));
NAND3X1 NAND3X1_19 ( .A(nRESET_G_bF_buf2), .B(_abc_898_new_n154_), .C(_abc_898_new_n153_), .Y(n55));
NAND3X1 NAND3X1_2 ( .A(D_OUT_REG_2_), .B(_abc_898_new_n156_), .C(_abc_898_new_n125_), .Y(_abc_898_new_n170_));
NAND3X1 NAND3X1_20 ( .A(D_OUT_REG_0_), .B(_abc_898_new_n156_), .C(_abc_898_new_n125_), .Y(_abc_898_new_n157_));
NAND3X1 NAND3X1_3 ( .A(D_OUT_REG_3_), .B(_abc_898_new_n156_), .C(_abc_898_new_n125_), .Y(_abc_898_new_n176_));
NAND3X1 NAND3X1_4 ( .A(D_OUT_REG_4_), .B(_abc_898_new_n156_), .C(_abc_898_new_n125_), .Y(_abc_898_new_n182_));
NAND3X1 NAND3X1_5 ( .A(D_OUT_REG_5_), .B(_abc_898_new_n156_), .C(_abc_898_new_n125_), .Y(_abc_898_new_n188_));
NAND3X1 NAND3X1_6 ( .A(D_OUT_REG_7_), .B(_abc_898_new_n156_), .C(_abc_898_new_n125_), .Y(_abc_898_new_n194_));
NAND3X1 NAND3X1_7 ( .A(D_OUT_REG_6_), .B(_abc_898_new_n156_), .C(_abc_898_new_n125_), .Y(_abc_898_new_n198_));
NAND3X1 NAND3X1_8 ( .A(_abc_898_new_n83_), .B(_abc_898_new_n81_), .C(_abc_898_new_n70_), .Y(_abc_898_new_n84_));
NAND3X1 NAND3X1_9 ( .A(_abc_898_new_n85_), .B(_abc_898_new_n87_), .C(_abc_898_new_n84_), .Y(n104));
NOR2X1 NOR2X1_1 ( .A(STATO_REG_1_), .B(_abc_898_new_n61_), .Y(_abc_898_new_n62_));
NOR2X1 NOR2X1_10 ( .A(_abc_898_new_n100_), .B(_abc_898_new_n98_), .Y(n144));
NOR2X1 NOR2X1_11 ( .A(_abc_898_new_n102_), .B(_abc_898_new_n98_), .Y(n139));
NOR2X1 NOR2X1_12 ( .A(_abc_898_new_n104_), .B(_abc_898_new_n98_), .Y(n134));
NOR2X1 NOR2X1_13 ( .A(_abc_898_new_n106_), .B(_abc_898_new_n98_), .Y(n129));
NOR2X1 NOR2X1_14 ( .A(_abc_898_new_n108_), .B(_abc_898_new_n98_), .Y(n124));
NOR2X1 NOR2X1_15 ( .A(_abc_898_new_n110_), .B(_abc_898_new_n98_), .Y(n119));
NOR2X1 NOR2X1_16 ( .A(_abc_898_new_n112_), .B(_abc_898_new_n98_), .Y(n114));
NOR2X1 NOR2X1_17 ( .A(_abc_898_new_n114_), .B(_abc_898_new_n115_), .Y(_abc_898_new_n116_));
NOR2X1 NOR2X1_18 ( .A(_abc_898_new_n117_), .B(_abc_898_new_n118_), .Y(_abc_898_new_n119_));
NOR2X1 NOR2X1_19 ( .A(D_IN_REG_0_), .B(_abc_898_new_n126_), .Y(_abc_898_new_n127_));
NOR2X1 NOR2X1_2 ( .A(_abc_898_new_n66_), .B(_abc_898_new_n69_), .Y(_abc_898_new_n70_));
NOR2X1 NOR2X1_3 ( .A(OLD_REG_0_), .B(D_IN_REG_1_), .Y(_abc_898_new_n76_));
NOR2X1 NOR2X1_4 ( .A(OLD_REG_1_), .B(D_IN_REG_2_), .Y(_abc_898_new_n79_));
NOR2X1 NOR2X1_5 ( .A(_abc_898_new_n80_), .B(_abc_898_new_n73_), .Y(_abc_898_new_n81_));
NOR2X1 NOR2X1_6 ( .A(_abc_898_new_n60_), .B(_abc_898_new_n82_), .Y(_abc_898_new_n83_));
NOR2X1 NOR2X1_7 ( .A(STATO_REG_1_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n89_));
NOR2X1 NOR2X1_8 ( .A(_abc_898_new_n59_), .B(_abc_898_new_n60_), .Y(_abc_898_new_n92_));
NOR2X1 NOR2X1_9 ( .A(_abc_898_new_n96_), .B(_abc_898_new_n98_), .Y(n10));
OAI21X1 OAI21X1_1 ( .A(_abc_898_new_n159_), .B(_abc_898_new_n160_), .C(nRESET_G_bF_buf3), .Y(_abc_898_new_n161_));
OAI21X1 OAI21X1_10 ( .A(_abc_898_new_n89_), .B(_abc_898_new_n90_), .C(X), .Y(_abc_898_new_n91_));
OAI21X1 OAI21X1_11 ( .A(_abc_898_new_n124_), .B(_abc_898_new_n120_), .C(_abc_898_new_n92_), .Y(_abc_898_new_n125_));
OAI21X1 OAI21X1_12 ( .A(D_IN_REG_0_), .B(_auto_iopadmap_cc_368_execute_1044), .C(_abc_898_new_n89_), .Y(_abc_898_new_n128_));
OAI21X1 OAI21X1_2 ( .A(_abc_898_new_n166_), .B(_abc_898_new_n160_), .C(nRESET_G_bF_buf2), .Y(_abc_898_new_n167_));
OAI21X1 OAI21X1_3 ( .A(_abc_898_new_n172_), .B(_abc_898_new_n160_), .C(nRESET_G_bF_buf1), .Y(_abc_898_new_n173_));
OAI21X1 OAI21X1_4 ( .A(_abc_898_new_n178_), .B(_abc_898_new_n160_), .C(nRESET_G_bF_buf0), .Y(_abc_898_new_n179_));
OAI21X1 OAI21X1_5 ( .A(_abc_898_new_n184_), .B(_abc_898_new_n160_), .C(nRESET_G_bF_buf3), .Y(_abc_898_new_n185_));
OAI21X1 OAI21X1_6 ( .A(_abc_898_new_n190_), .B(_abc_898_new_n160_), .C(nRESET_G_bF_buf2), .Y(_abc_898_new_n191_));
OAI21X1 OAI21X1_7 ( .A(_abc_898_new_n200_), .B(_abc_898_new_n160_), .C(nRESET_G_bF_buf1), .Y(_abc_898_new_n201_));
OAI21X1 OAI21X1_8 ( .A(_abc_898_new_n59_), .B(_abc_898_new_n60_), .C(_abc_898_new_n62_), .Y(n99));
OAI21X1 OAI21X1_9 ( .A(STATO_REG_0_), .B(_abc_898_new_n82_), .C(_abc_898_new_n86_), .Y(_abc_898_new_n90_));
OAI22X1 OAI22X1_1 ( .A(_abc_898_new_n76_), .B(_abc_898_new_n75_), .C(_abc_898_new_n78_), .D(_abc_898_new_n79_), .Y(_abc_898_new_n80_));
XNOR2X1 XNOR2X1_1 ( .A(OLD_REG_7_), .B(D_IN_REG_8_), .Y(_abc_898_new_n64_));
XNOR2X1 XNOR2X1_2 ( .A(D_IN_REG_7_), .B(OLD_REG_6_), .Y(_abc_898_new_n65_));
XNOR2X1 XNOR2X1_3 ( .A(OLD_REG_2_), .B(D_IN_REG_3_), .Y(_abc_898_new_n67_));
XNOR2X1 XNOR2X1_4 ( .A(D_IN_REG_4_), .B(OLD_REG_3_), .Y(_abc_898_new_n68_));
XNOR2X1 XNOR2X1_5 ( .A(OLD_REG_4_), .B(D_IN_REG_5_), .Y(_abc_898_new_n71_));
XNOR2X1 XNOR2X1_6 ( .A(D_IN_REG_6_), .B(OLD_REG_5_), .Y(_abc_898_new_n72_));
XOR2X1 XOR2X1_1 ( .A(OLD_REG_7_), .B(D_IN_REG_8_), .Y(_abc_898_new_n114_));
XOR2X1 XOR2X1_2 ( .A(D_IN_REG_7_), .B(OLD_REG_6_), .Y(_abc_898_new_n115_));
XOR2X1 XOR2X1_3 ( .A(OLD_REG_2_), .B(D_IN_REG_3_), .Y(_abc_898_new_n117_));
XOR2X1 XOR2X1_4 ( .A(D_IN_REG_4_), .B(OLD_REG_3_), .Y(_abc_898_new_n118_));


endmodule