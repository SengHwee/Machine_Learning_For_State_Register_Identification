module cpu8080(\data[0] , \data[1] , \data[2] , \data[3] , \data[4] , \data[5] , \data[6] , \data[7] , intr, waitr, reset, clock, \addr[0] , \addr[1] , \addr[2] , \addr[3] , \addr[4] , \addr[5] , \addr[6] , \addr[7] , \addr[8] , \addr[9] , \addr[10] , \addr[11] , \addr[12] , \addr[13] , \addr[14] , \addr[15] , readmem, writemem, readio, writeio, inta);

wire _0addr_15_0__0_; 
wire _0addr_15_0__10_; 
wire _0addr_15_0__11_; 
wire _0addr_15_0__12_; 
wire _0addr_15_0__13_; 
wire _0addr_15_0__14_; 
wire _0addr_15_0__15_; 
wire _0addr_15_0__1_; 
wire _0addr_15_0__2_; 
wire _0addr_15_0__3_; 
wire _0addr_15_0__4_; 
wire _0addr_15_0__5_; 
wire _0addr_15_0__6_; 
wire _0addr_15_0__7_; 
wire _0addr_15_0__8_; 
wire _0addr_15_0__9_; 
wire _0alucin_0_0_; 
wire _0aluopra_7_0__0_; 
wire _0aluopra_7_0__1_; 
wire _0aluopra_7_0__2_; 
wire _0aluopra_7_0__3_; 
wire _0aluopra_7_0__4_; 
wire _0aluopra_7_0__5_; 
wire _0aluopra_7_0__6_; 
wire _0aluopra_7_0__7_; 
wire _0aluoprb_7_0__0_; 
wire _0aluoprb_7_0__1_; 
wire _0aluoprb_7_0__2_; 
wire _0aluoprb_7_0__3_; 
wire _0aluoprb_7_0__4_; 
wire _0aluoprb_7_0__5_; 
wire _0aluoprb_7_0__6_; 
wire _0aluoprb_7_0__7_; 
wire _0alusel_2_0__0_; 
wire _0alusel_2_0__1_; 
wire _0alusel_2_0__2_; 
wire _0auxcar_0_0_; 
wire _0carry_0_0_; 
wire _0datao_7_0__0_; 
wire _0datao_7_0__1_; 
wire _0datao_7_0__2_; 
wire _0datao_7_0__3_; 
wire _0datao_7_0__4_; 
wire _0datao_7_0__5_; 
wire _0datao_7_0__6_; 
wire _0datao_7_0__7_; 
wire _0ei_0_0_; 
wire _0eienb_0_0_; 
wire _0inta_0_0_; 
wire _0intcyc_0_0_; 
wire _0opcode_7_0__0_; 
wire _0opcode_7_0__1_; 
wire _0opcode_7_0__2_; 
wire _0opcode_7_0__3_; 
wire _0opcode_7_0__4_; 
wire _0opcode_7_0__5_; 
wire _0opcode_7_0__6_; 
wire _0opcode_7_0__7_; 
wire _0parity_0_0_; 
wire _0pc_15_0__0_; 
wire _0pc_15_0__10_; 
wire _0pc_15_0__11_; 
wire _0pc_15_0__12_; 
wire _0pc_15_0__13_; 
wire _0pc_15_0__14_; 
wire _0pc_15_0__15_; 
wire _0pc_15_0__1_; 
wire _0pc_15_0__2_; 
wire _0pc_15_0__3_; 
wire _0pc_15_0__4_; 
wire _0pc_15_0__5_; 
wire _0pc_15_0__6_; 
wire _0pc_15_0__7_; 
wire _0pc_15_0__8_; 
wire _0pc_15_0__9_; 
wire _0popdes_1_0__0_; 
wire _0popdes_1_0__1_; 
wire _0raddrhold_15_0__0_; 
wire _0raddrhold_15_0__10_; 
wire _0raddrhold_15_0__11_; 
wire _0raddrhold_15_0__12_; 
wire _0raddrhold_15_0__13_; 
wire _0raddrhold_15_0__14_; 
wire _0raddrhold_15_0__15_; 
wire _0raddrhold_15_0__1_; 
wire _0raddrhold_15_0__2_; 
wire _0raddrhold_15_0__3_; 
wire _0raddrhold_15_0__4_; 
wire _0raddrhold_15_0__5_; 
wire _0raddrhold_15_0__6_; 
wire _0raddrhold_15_0__7_; 
wire _0raddrhold_15_0__8_; 
wire _0raddrhold_15_0__9_; 
wire _0rdatahold2_7_0__0_; 
wire _0rdatahold2_7_0__1_; 
wire _0rdatahold2_7_0__2_; 
wire _0rdatahold2_7_0__3_; 
wire _0rdatahold2_7_0__4_; 
wire _0rdatahold2_7_0__5_; 
wire _0rdatahold2_7_0__6_; 
wire _0rdatahold2_7_0__7_; 
wire _0rdatahold_7_0__0_; 
wire _0rdatahold_7_0__1_; 
wire _0rdatahold_7_0__2_; 
wire _0rdatahold_7_0__3_; 
wire _0rdatahold_7_0__4_; 
wire _0rdatahold_7_0__5_; 
wire _0rdatahold_7_0__6_; 
wire _0rdatahold_7_0__7_; 
wire _0readio_0_0_; 
wire _0readmem_0_0_; 
wire _0regd_2_0__0_; 
wire _0regd_2_0__1_; 
wire _0regd_2_0__2_; 
wire _0sign_0_0_; 
wire _0sp_15_0__0_; 
wire _0sp_15_0__10_; 
wire _0sp_15_0__11_; 
wire _0sp_15_0__12_; 
wire _0sp_15_0__13_; 
wire _0sp_15_0__14_; 
wire _0sp_15_0__15_; 
wire _0sp_15_0__1_; 
wire _0sp_15_0__2_; 
wire _0sp_15_0__3_; 
wire _0sp_15_0__4_; 
wire _0sp_15_0__5_; 
wire _0sp_15_0__6_; 
wire _0sp_15_0__7_; 
wire _0sp_15_0__8_; 
wire _0sp_15_0__9_; 
wire _0statesel_5_0__0_; 
wire _0statesel_5_0__1_; 
wire _0statesel_5_0__2_; 
wire _0statesel_5_0__3_; 
wire _0statesel_5_0__4_; 
wire _0statesel_5_0__5_; 
wire _0waddrhold_15_0__0_; 
wire _0waddrhold_15_0__10_; 
wire _0waddrhold_15_0__11_; 
wire _0waddrhold_15_0__12_; 
wire _0waddrhold_15_0__13_; 
wire _0waddrhold_15_0__14_; 
wire _0waddrhold_15_0__15_; 
wire _0waddrhold_15_0__1_; 
wire _0waddrhold_15_0__2_; 
wire _0waddrhold_15_0__3_; 
wire _0waddrhold_15_0__4_; 
wire _0waddrhold_15_0__5_; 
wire _0waddrhold_15_0__6_; 
wire _0waddrhold_15_0__7_; 
wire _0waddrhold_15_0__8_; 
wire _0waddrhold_15_0__9_; 
wire _0wdatahold2_7_0__0_; 
wire _0wdatahold2_7_0__1_; 
wire _0wdatahold2_7_0__2_; 
wire _0wdatahold2_7_0__3_; 
wire _0wdatahold2_7_0__4_; 
wire _0wdatahold2_7_0__5_; 
wire _0wdatahold2_7_0__6_; 
wire _0wdatahold2_7_0__7_; 
wire _0wdatahold_7_0__0_; 
wire _0wdatahold_7_0__1_; 
wire _0wdatahold_7_0__2_; 
wire _0wdatahold_7_0__3_; 
wire _0wdatahold_7_0__4_; 
wire _0wdatahold_7_0__5_; 
wire _0wdatahold_7_0__6_; 
wire _0wdatahold_7_0__7_; 
wire _0writeio_0_0_; 
wire _0writemem_0_0_; 
wire _0zero_0_0_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_0_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_1_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_2_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_3_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_4_; 
wire _abc_36060_auto_fsm_map_cc_170_map_fsm_12881_5_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_0_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_1_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_2_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_3_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_4_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_5_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_6_; 
wire _abc_36060_memoryregfil_wrmux_0__0__0__y_15937_7_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_0_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_1_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_2_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_3_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_4_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_5_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_6_; 
wire _abc_36060_memoryregfil_wrmux_1__1__0__y_16001_7_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_0_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_1_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_2_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_3_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_4_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_5_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_6_; 
wire _abc_36060_memoryregfil_wrmux_2__1__0__y_16043_7_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_0_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_1_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_2_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_3_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_4_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_5_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_6_; 
wire _abc_36060_memoryregfil_wrmux_3__2__0__y_16089_7_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_0_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_1_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_2_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_3_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_4_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_5_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_6_; 
wire _abc_36060_memoryregfil_wrmux_4__4__0__y_16147_7_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_0_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_1_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_2_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_3_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_4_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_5_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_6_; 
wire _abc_36060_memoryregfil_wrmux_5__3__0__y_16171_7_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_0_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_1_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_2_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_3_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_4_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_5_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_6_; 
wire _abc_36060_memoryregfil_wrmux_6__0__0__y_16185_7_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_0_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_1_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_2_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_3_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_4_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_5_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_6_; 
wire _abc_36060_memoryregfil_wrmux_7__4__0__y_16247_7_; 
wire _abc_41356_new_n1000_; 
wire _abc_41356_new_n1001_; 
wire _abc_41356_new_n1002_; 
wire _abc_41356_new_n1003_; 
wire _abc_41356_new_n1004_; 
wire _abc_41356_new_n1005_; 
wire _abc_41356_new_n1006_; 
wire _abc_41356_new_n1007_; 
wire _abc_41356_new_n1008_; 
wire _abc_41356_new_n1009_; 
wire _abc_41356_new_n1010_; 
wire _abc_41356_new_n1011_; 
wire _abc_41356_new_n1012_; 
wire _abc_41356_new_n1013_; 
wire _abc_41356_new_n1014_; 
wire _abc_41356_new_n1015_; 
wire _abc_41356_new_n1016_; 
wire _abc_41356_new_n1017_; 
wire _abc_41356_new_n1018_; 
wire _abc_41356_new_n1019_; 
wire _abc_41356_new_n1020_; 
wire _abc_41356_new_n1021_; 
wire _abc_41356_new_n1022_; 
wire _abc_41356_new_n1023_; 
wire _abc_41356_new_n1024_; 
wire _abc_41356_new_n1025_; 
wire _abc_41356_new_n1026_; 
wire _abc_41356_new_n1027_; 
wire _abc_41356_new_n1028_; 
wire _abc_41356_new_n1029_; 
wire _abc_41356_new_n1030_; 
wire _abc_41356_new_n1031_; 
wire _abc_41356_new_n1032_; 
wire _abc_41356_new_n1033_; 
wire _abc_41356_new_n1034_; 
wire _abc_41356_new_n1035_; 
wire _abc_41356_new_n1036_; 
wire _abc_41356_new_n1037_; 
wire _abc_41356_new_n1038_; 
wire _abc_41356_new_n1039_; 
wire _abc_41356_new_n1040_; 
wire _abc_41356_new_n1041_; 
wire _abc_41356_new_n1042_; 
wire _abc_41356_new_n1043_; 
wire _abc_41356_new_n1044_; 
wire _abc_41356_new_n1045_; 
wire _abc_41356_new_n1046_; 
wire _abc_41356_new_n1047_; 
wire _abc_41356_new_n1048_; 
wire _abc_41356_new_n1049_; 
wire _abc_41356_new_n1050_; 
wire _abc_41356_new_n1052_; 
wire _abc_41356_new_n1053_; 
wire _abc_41356_new_n1054_; 
wire _abc_41356_new_n1055_; 
wire _abc_41356_new_n1056_; 
wire _abc_41356_new_n1057_; 
wire _abc_41356_new_n1058_; 
wire _abc_41356_new_n1059_; 
wire _abc_41356_new_n1060_; 
wire _abc_41356_new_n1061_; 
wire _abc_41356_new_n1062_; 
wire _abc_41356_new_n1063_; 
wire _abc_41356_new_n1064_; 
wire _abc_41356_new_n1065_; 
wire _abc_41356_new_n1066_; 
wire _abc_41356_new_n1067_; 
wire _abc_41356_new_n1068_; 
wire _abc_41356_new_n1069_; 
wire _abc_41356_new_n1070_; 
wire _abc_41356_new_n1071_; 
wire _abc_41356_new_n1072_; 
wire _abc_41356_new_n1073_; 
wire _abc_41356_new_n1074_; 
wire _abc_41356_new_n1075_; 
wire _abc_41356_new_n1076_; 
wire _abc_41356_new_n1077_; 
wire _abc_41356_new_n1078_; 
wire _abc_41356_new_n1079_; 
wire _abc_41356_new_n1080_; 
wire _abc_41356_new_n1081_; 
wire _abc_41356_new_n1082_; 
wire _abc_41356_new_n1083_; 
wire _abc_41356_new_n1084_; 
wire _abc_41356_new_n1085_; 
wire _abc_41356_new_n1086_; 
wire _abc_41356_new_n1087_; 
wire _abc_41356_new_n1088_; 
wire _abc_41356_new_n1089_; 
wire _abc_41356_new_n1090_; 
wire _abc_41356_new_n1091_; 
wire _abc_41356_new_n1092_; 
wire _abc_41356_new_n1093_; 
wire _abc_41356_new_n1094_; 
wire _abc_41356_new_n1095_; 
wire _abc_41356_new_n1096_; 
wire _abc_41356_new_n1097_; 
wire _abc_41356_new_n1098_; 
wire _abc_41356_new_n1099_; 
wire _abc_41356_new_n1100_; 
wire _abc_41356_new_n1101_; 
wire _abc_41356_new_n1102_; 
wire _abc_41356_new_n1103_; 
wire _abc_41356_new_n1104_; 
wire _abc_41356_new_n1105_; 
wire _abc_41356_new_n1106_; 
wire _abc_41356_new_n1107_; 
wire _abc_41356_new_n1108_; 
wire _abc_41356_new_n1109_; 
wire _abc_41356_new_n1110_; 
wire _abc_41356_new_n1111_; 
wire _abc_41356_new_n1112_; 
wire _abc_41356_new_n1113_; 
wire _abc_41356_new_n1114_; 
wire _abc_41356_new_n1115_; 
wire _abc_41356_new_n1116_; 
wire _abc_41356_new_n1117_; 
wire _abc_41356_new_n1118_; 
wire _abc_41356_new_n1119_; 
wire _abc_41356_new_n1120_; 
wire _abc_41356_new_n1121_; 
wire _abc_41356_new_n1122_; 
wire _abc_41356_new_n1123_; 
wire _abc_41356_new_n1124_; 
wire _abc_41356_new_n1125_; 
wire _abc_41356_new_n1126_; 
wire _abc_41356_new_n1127_; 
wire _abc_41356_new_n1128_; 
wire _abc_41356_new_n1129_; 
wire _abc_41356_new_n1130_; 
wire _abc_41356_new_n1131_; 
wire _abc_41356_new_n1132_; 
wire _abc_41356_new_n1134_; 
wire _abc_41356_new_n1135_; 
wire _abc_41356_new_n1136_; 
wire _abc_41356_new_n1137_; 
wire _abc_41356_new_n1138_; 
wire _abc_41356_new_n1139_; 
wire _abc_41356_new_n1140_; 
wire _abc_41356_new_n1141_; 
wire _abc_41356_new_n1142_; 
wire _abc_41356_new_n1143_; 
wire _abc_41356_new_n1144_; 
wire _abc_41356_new_n1145_; 
wire _abc_41356_new_n1146_; 
wire _abc_41356_new_n1147_; 
wire _abc_41356_new_n1148_; 
wire _abc_41356_new_n1149_; 
wire _abc_41356_new_n1150_; 
wire _abc_41356_new_n1151_; 
wire _abc_41356_new_n1152_; 
wire _abc_41356_new_n1153_; 
wire _abc_41356_new_n1154_; 
wire _abc_41356_new_n1155_; 
wire _abc_41356_new_n1156_; 
wire _abc_41356_new_n1157_; 
wire _abc_41356_new_n1158_; 
wire _abc_41356_new_n1159_; 
wire _abc_41356_new_n1160_; 
wire _abc_41356_new_n1161_; 
wire _abc_41356_new_n1162_; 
wire _abc_41356_new_n1163_; 
wire _abc_41356_new_n1164_; 
wire _abc_41356_new_n1165_; 
wire _abc_41356_new_n1166_; 
wire _abc_41356_new_n1167_; 
wire _abc_41356_new_n1168_; 
wire _abc_41356_new_n1169_; 
wire _abc_41356_new_n1170_; 
wire _abc_41356_new_n1171_; 
wire _abc_41356_new_n1172_; 
wire _abc_41356_new_n1173_; 
wire _abc_41356_new_n1174_; 
wire _abc_41356_new_n1175_; 
wire _abc_41356_new_n1176_; 
wire _abc_41356_new_n1177_; 
wire _abc_41356_new_n1178_; 
wire _abc_41356_new_n1179_; 
wire _abc_41356_new_n1180_; 
wire _abc_41356_new_n1181_; 
wire _abc_41356_new_n1182_; 
wire _abc_41356_new_n1183_; 
wire _abc_41356_new_n1184_; 
wire _abc_41356_new_n1185_; 
wire _abc_41356_new_n1186_; 
wire _abc_41356_new_n1187_; 
wire _abc_41356_new_n1188_; 
wire _abc_41356_new_n1189_; 
wire _abc_41356_new_n1190_; 
wire _abc_41356_new_n1191_; 
wire _abc_41356_new_n1192_; 
wire _abc_41356_new_n1193_; 
wire _abc_41356_new_n1194_; 
wire _abc_41356_new_n1195_; 
wire _abc_41356_new_n1196_; 
wire _abc_41356_new_n1197_; 
wire _abc_41356_new_n1198_; 
wire _abc_41356_new_n1199_; 
wire _abc_41356_new_n1200_; 
wire _abc_41356_new_n1201_; 
wire _abc_41356_new_n1202_; 
wire _abc_41356_new_n1203_; 
wire _abc_41356_new_n1204_; 
wire _abc_41356_new_n1205_; 
wire _abc_41356_new_n1207_; 
wire _abc_41356_new_n1208_; 
wire _abc_41356_new_n1209_; 
wire _abc_41356_new_n1210_; 
wire _abc_41356_new_n1211_; 
wire _abc_41356_new_n1212_; 
wire _abc_41356_new_n1213_; 
wire _abc_41356_new_n1214_; 
wire _abc_41356_new_n1215_; 
wire _abc_41356_new_n1216_; 
wire _abc_41356_new_n1217_; 
wire _abc_41356_new_n1218_; 
wire _abc_41356_new_n1219_; 
wire _abc_41356_new_n1220_; 
wire _abc_41356_new_n1221_; 
wire _abc_41356_new_n1222_; 
wire _abc_41356_new_n1223_; 
wire _abc_41356_new_n1224_; 
wire _abc_41356_new_n1225_; 
wire _abc_41356_new_n1226_; 
wire _abc_41356_new_n1227_; 
wire _abc_41356_new_n1228_; 
wire _abc_41356_new_n1229_; 
wire _abc_41356_new_n1230_; 
wire _abc_41356_new_n1231_; 
wire _abc_41356_new_n1232_; 
wire _abc_41356_new_n1233_; 
wire _abc_41356_new_n1234_; 
wire _abc_41356_new_n1235_; 
wire _abc_41356_new_n1236_; 
wire _abc_41356_new_n1237_; 
wire _abc_41356_new_n1238_; 
wire _abc_41356_new_n1239_; 
wire _abc_41356_new_n1240_; 
wire _abc_41356_new_n1241_; 
wire _abc_41356_new_n1242_; 
wire _abc_41356_new_n1243_; 
wire _abc_41356_new_n1244_; 
wire _abc_41356_new_n1245_; 
wire _abc_41356_new_n1246_; 
wire _abc_41356_new_n1247_; 
wire _abc_41356_new_n1248_; 
wire _abc_41356_new_n1249_; 
wire _abc_41356_new_n1250_; 
wire _abc_41356_new_n1251_; 
wire _abc_41356_new_n1252_; 
wire _abc_41356_new_n1253_; 
wire _abc_41356_new_n1254_; 
wire _abc_41356_new_n1255_; 
wire _abc_41356_new_n1256_; 
wire _abc_41356_new_n1257_; 
wire _abc_41356_new_n1258_; 
wire _abc_41356_new_n1259_; 
wire _abc_41356_new_n1260_; 
wire _abc_41356_new_n1261_; 
wire _abc_41356_new_n1262_; 
wire _abc_41356_new_n1263_; 
wire _abc_41356_new_n1264_; 
wire _abc_41356_new_n1265_; 
wire _abc_41356_new_n1266_; 
wire _abc_41356_new_n1267_; 
wire _abc_41356_new_n1268_; 
wire _abc_41356_new_n1269_; 
wire _abc_41356_new_n1270_; 
wire _abc_41356_new_n1271_; 
wire _abc_41356_new_n1272_; 
wire _abc_41356_new_n1273_; 
wire _abc_41356_new_n1274_; 
wire _abc_41356_new_n1275_; 
wire _abc_41356_new_n1276_; 
wire _abc_41356_new_n1277_; 
wire _abc_41356_new_n1278_; 
wire _abc_41356_new_n1279_; 
wire _abc_41356_new_n1280_; 
wire _abc_41356_new_n1281_; 
wire _abc_41356_new_n1282_; 
wire _abc_41356_new_n1283_; 
wire _abc_41356_new_n1284_; 
wire _abc_41356_new_n1285_; 
wire _abc_41356_new_n1286_; 
wire _abc_41356_new_n1287_; 
wire _abc_41356_new_n1288_; 
wire _abc_41356_new_n1289_; 
wire _abc_41356_new_n1290_; 
wire _abc_41356_new_n1291_; 
wire _abc_41356_new_n1292_; 
wire _abc_41356_new_n1293_; 
wire _abc_41356_new_n1294_; 
wire _abc_41356_new_n1295_; 
wire _abc_41356_new_n1296_; 
wire _abc_41356_new_n1297_; 
wire _abc_41356_new_n1298_; 
wire _abc_41356_new_n1299_; 
wire _abc_41356_new_n1300_; 
wire _abc_41356_new_n1301_; 
wire _abc_41356_new_n1302_; 
wire _abc_41356_new_n1303_; 
wire _abc_41356_new_n1304_; 
wire _abc_41356_new_n1305_; 
wire _abc_41356_new_n1306_; 
wire _abc_41356_new_n1307_; 
wire _abc_41356_new_n1308_; 
wire _abc_41356_new_n1309_; 
wire _abc_41356_new_n1310_; 
wire _abc_41356_new_n1311_; 
wire _abc_41356_new_n1312_; 
wire _abc_41356_new_n1313_; 
wire _abc_41356_new_n1314_; 
wire _abc_41356_new_n1315_; 
wire _abc_41356_new_n1316_; 
wire _abc_41356_new_n1317_; 
wire _abc_41356_new_n1318_; 
wire _abc_41356_new_n1319_; 
wire _abc_41356_new_n1320_; 
wire _abc_41356_new_n1321_; 
wire _abc_41356_new_n1322_; 
wire _abc_41356_new_n1323_; 
wire _abc_41356_new_n1324_; 
wire _abc_41356_new_n1325_; 
wire _abc_41356_new_n1326_; 
wire _abc_41356_new_n1327_; 
wire _abc_41356_new_n1328_; 
wire _abc_41356_new_n1329_; 
wire _abc_41356_new_n1330_; 
wire _abc_41356_new_n1331_; 
wire _abc_41356_new_n1332_; 
wire _abc_41356_new_n1333_; 
wire _abc_41356_new_n1334_; 
wire _abc_41356_new_n1335_; 
wire _abc_41356_new_n1336_; 
wire _abc_41356_new_n1337_; 
wire _abc_41356_new_n1338_; 
wire _abc_41356_new_n1339_; 
wire _abc_41356_new_n1340_; 
wire _abc_41356_new_n1341_; 
wire _abc_41356_new_n1342_; 
wire _abc_41356_new_n1343_; 
wire _abc_41356_new_n1344_; 
wire _abc_41356_new_n1345_; 
wire _abc_41356_new_n1346_; 
wire _abc_41356_new_n1347_; 
wire _abc_41356_new_n1348_; 
wire _abc_41356_new_n1349_; 
wire _abc_41356_new_n1350_; 
wire _abc_41356_new_n1351_; 
wire _abc_41356_new_n1352_; 
wire _abc_41356_new_n1353_; 
wire _abc_41356_new_n1354_; 
wire _abc_41356_new_n1355_; 
wire _abc_41356_new_n1356_; 
wire _abc_41356_new_n1357_; 
wire _abc_41356_new_n1358_; 
wire _abc_41356_new_n1359_; 
wire _abc_41356_new_n1360_; 
wire _abc_41356_new_n1361_; 
wire _abc_41356_new_n1362_; 
wire _abc_41356_new_n1363_; 
wire _abc_41356_new_n1364_; 
wire _abc_41356_new_n1365_; 
wire _abc_41356_new_n1366_; 
wire _abc_41356_new_n1367_; 
wire _abc_41356_new_n1368_; 
wire _abc_41356_new_n1369_; 
wire _abc_41356_new_n1370_; 
wire _abc_41356_new_n1371_; 
wire _abc_41356_new_n1372_; 
wire _abc_41356_new_n1373_; 
wire _abc_41356_new_n1374_; 
wire _abc_41356_new_n1375_; 
wire _abc_41356_new_n1376_; 
wire _abc_41356_new_n1377_; 
wire _abc_41356_new_n1378_; 
wire _abc_41356_new_n1379_; 
wire _abc_41356_new_n1380_; 
wire _abc_41356_new_n1381_; 
wire _abc_41356_new_n1382_; 
wire _abc_41356_new_n1383_; 
wire _abc_41356_new_n1384_; 
wire _abc_41356_new_n1385_; 
wire _abc_41356_new_n1386_; 
wire _abc_41356_new_n1387_; 
wire _abc_41356_new_n1388_; 
wire _abc_41356_new_n1389_; 
wire _abc_41356_new_n1390_; 
wire _abc_41356_new_n1391_; 
wire _abc_41356_new_n1392_; 
wire _abc_41356_new_n1393_; 
wire _abc_41356_new_n1394_; 
wire _abc_41356_new_n1395_; 
wire _abc_41356_new_n1396_; 
wire _abc_41356_new_n1397_; 
wire _abc_41356_new_n1398_; 
wire _abc_41356_new_n1399_; 
wire _abc_41356_new_n1400_; 
wire _abc_41356_new_n1401_; 
wire _abc_41356_new_n1402_; 
wire _abc_41356_new_n1403_; 
wire _abc_41356_new_n1404_; 
wire _abc_41356_new_n1405_; 
wire _abc_41356_new_n1406_; 
wire _abc_41356_new_n1407_; 
wire _abc_41356_new_n1408_; 
wire _abc_41356_new_n1409_; 
wire _abc_41356_new_n1410_; 
wire _abc_41356_new_n1411_; 
wire _abc_41356_new_n1412_; 
wire _abc_41356_new_n1413_; 
wire _abc_41356_new_n1414_; 
wire _abc_41356_new_n1415_; 
wire _abc_41356_new_n1416_; 
wire _abc_41356_new_n1417_; 
wire _abc_41356_new_n1418_; 
wire _abc_41356_new_n1419_; 
wire _abc_41356_new_n1420_; 
wire _abc_41356_new_n1421_; 
wire _abc_41356_new_n1422_; 
wire _abc_41356_new_n1423_; 
wire _abc_41356_new_n1424_; 
wire _abc_41356_new_n1425_; 
wire _abc_41356_new_n1426_; 
wire _abc_41356_new_n1427_; 
wire _abc_41356_new_n1428_; 
wire _abc_41356_new_n1429_; 
wire _abc_41356_new_n1430_; 
wire _abc_41356_new_n1431_; 
wire _abc_41356_new_n1432_; 
wire _abc_41356_new_n1433_; 
wire _abc_41356_new_n1434_; 
wire _abc_41356_new_n1435_; 
wire _abc_41356_new_n1436_; 
wire _abc_41356_new_n1437_; 
wire _abc_41356_new_n1438_; 
wire _abc_41356_new_n1439_; 
wire _abc_41356_new_n1440_; 
wire _abc_41356_new_n1441_; 
wire _abc_41356_new_n1442_; 
wire _abc_41356_new_n1443_; 
wire _abc_41356_new_n1444_; 
wire _abc_41356_new_n1445_; 
wire _abc_41356_new_n1446_; 
wire _abc_41356_new_n1447_; 
wire _abc_41356_new_n1448_; 
wire _abc_41356_new_n1449_; 
wire _abc_41356_new_n1450_; 
wire _abc_41356_new_n1451_; 
wire _abc_41356_new_n1452_; 
wire _abc_41356_new_n1453_; 
wire _abc_41356_new_n1454_; 
wire _abc_41356_new_n1455_; 
wire _abc_41356_new_n1456_; 
wire _abc_41356_new_n1457_; 
wire _abc_41356_new_n1458_; 
wire _abc_41356_new_n1459_; 
wire _abc_41356_new_n1460_; 
wire _abc_41356_new_n1461_; 
wire _abc_41356_new_n1462_; 
wire _abc_41356_new_n1463_; 
wire _abc_41356_new_n1464_; 
wire _abc_41356_new_n1465_; 
wire _abc_41356_new_n1466_; 
wire _abc_41356_new_n1467_; 
wire _abc_41356_new_n1468_; 
wire _abc_41356_new_n1469_; 
wire _abc_41356_new_n1470_; 
wire _abc_41356_new_n1471_; 
wire _abc_41356_new_n1472_; 
wire _abc_41356_new_n1473_; 
wire _abc_41356_new_n1474_; 
wire _abc_41356_new_n1475_; 
wire _abc_41356_new_n1476_; 
wire _abc_41356_new_n1477_; 
wire _abc_41356_new_n1478_; 
wire _abc_41356_new_n1479_; 
wire _abc_41356_new_n1480_; 
wire _abc_41356_new_n1481_; 
wire _abc_41356_new_n1482_; 
wire _abc_41356_new_n1483_; 
wire _abc_41356_new_n1484_; 
wire _abc_41356_new_n1485_; 
wire _abc_41356_new_n1486_; 
wire _abc_41356_new_n1487_; 
wire _abc_41356_new_n1488_; 
wire _abc_41356_new_n1489_; 
wire _abc_41356_new_n1490_; 
wire _abc_41356_new_n1491_; 
wire _abc_41356_new_n1492_; 
wire _abc_41356_new_n1493_; 
wire _abc_41356_new_n1494_; 
wire _abc_41356_new_n1496_; 
wire _abc_41356_new_n1497_; 
wire _abc_41356_new_n1498_; 
wire _abc_41356_new_n1499_; 
wire _abc_41356_new_n1500_; 
wire _abc_41356_new_n1501_; 
wire _abc_41356_new_n1502_; 
wire _abc_41356_new_n1503_; 
wire _abc_41356_new_n1504_; 
wire _abc_41356_new_n1505_; 
wire _abc_41356_new_n1506_; 
wire _abc_41356_new_n1507_; 
wire _abc_41356_new_n1508_; 
wire _abc_41356_new_n1509_; 
wire _abc_41356_new_n1510_; 
wire _abc_41356_new_n1511_; 
wire _abc_41356_new_n1512_; 
wire _abc_41356_new_n1513_; 
wire _abc_41356_new_n1514_; 
wire _abc_41356_new_n1515_; 
wire _abc_41356_new_n1516_; 
wire _abc_41356_new_n1517_; 
wire _abc_41356_new_n1518_; 
wire _abc_41356_new_n1519_; 
wire _abc_41356_new_n1520_; 
wire _abc_41356_new_n1521_; 
wire _abc_41356_new_n1522_; 
wire _abc_41356_new_n1523_; 
wire _abc_41356_new_n1524_; 
wire _abc_41356_new_n1525_; 
wire _abc_41356_new_n1526_; 
wire _abc_41356_new_n1527_; 
wire _abc_41356_new_n1528_; 
wire _abc_41356_new_n1529_; 
wire _abc_41356_new_n1530_; 
wire _abc_41356_new_n1531_; 
wire _abc_41356_new_n1532_; 
wire _abc_41356_new_n1533_; 
wire _abc_41356_new_n1534_; 
wire _abc_41356_new_n1535_; 
wire _abc_41356_new_n1536_; 
wire _abc_41356_new_n1537_; 
wire _abc_41356_new_n1538_; 
wire _abc_41356_new_n1539_; 
wire _abc_41356_new_n1540_; 
wire _abc_41356_new_n1541_; 
wire _abc_41356_new_n1542_; 
wire _abc_41356_new_n1543_; 
wire _abc_41356_new_n1544_; 
wire _abc_41356_new_n1545_; 
wire _abc_41356_new_n1546_; 
wire _abc_41356_new_n1547_; 
wire _abc_41356_new_n1548_; 
wire _abc_41356_new_n1549_; 
wire _abc_41356_new_n1550_; 
wire _abc_41356_new_n1551_; 
wire _abc_41356_new_n1552_; 
wire _abc_41356_new_n1553_; 
wire _abc_41356_new_n1554_; 
wire _abc_41356_new_n1555_; 
wire _abc_41356_new_n1556_; 
wire _abc_41356_new_n1557_; 
wire _abc_41356_new_n1558_; 
wire _abc_41356_new_n1559_; 
wire _abc_41356_new_n1560_; 
wire _abc_41356_new_n1561_; 
wire _abc_41356_new_n1562_; 
wire _abc_41356_new_n1563_; 
wire _abc_41356_new_n1564_; 
wire _abc_41356_new_n1565_; 
wire _abc_41356_new_n1566_; 
wire _abc_41356_new_n1567_; 
wire _abc_41356_new_n1568_; 
wire _abc_41356_new_n1569_; 
wire _abc_41356_new_n1570_; 
wire _abc_41356_new_n1572_; 
wire _abc_41356_new_n1573_; 
wire _abc_41356_new_n1574_; 
wire _abc_41356_new_n1575_; 
wire _abc_41356_new_n1576_; 
wire _abc_41356_new_n1577_; 
wire _abc_41356_new_n1578_; 
wire _abc_41356_new_n1579_; 
wire _abc_41356_new_n1580_; 
wire _abc_41356_new_n1581_; 
wire _abc_41356_new_n1582_; 
wire _abc_41356_new_n1583_; 
wire _abc_41356_new_n1584_; 
wire _abc_41356_new_n1585_; 
wire _abc_41356_new_n1586_; 
wire _abc_41356_new_n1587_; 
wire _abc_41356_new_n1588_; 
wire _abc_41356_new_n1589_; 
wire _abc_41356_new_n1590_; 
wire _abc_41356_new_n1591_; 
wire _abc_41356_new_n1592_; 
wire _abc_41356_new_n1593_; 
wire _abc_41356_new_n1594_; 
wire _abc_41356_new_n1595_; 
wire _abc_41356_new_n1596_; 
wire _abc_41356_new_n1597_; 
wire _abc_41356_new_n1598_; 
wire _abc_41356_new_n1599_; 
wire _abc_41356_new_n1600_; 
wire _abc_41356_new_n1601_; 
wire _abc_41356_new_n1602_; 
wire _abc_41356_new_n1603_; 
wire _abc_41356_new_n1604_; 
wire _abc_41356_new_n1605_; 
wire _abc_41356_new_n1606_; 
wire _abc_41356_new_n1607_; 
wire _abc_41356_new_n1608_; 
wire _abc_41356_new_n1609_; 
wire _abc_41356_new_n1610_; 
wire _abc_41356_new_n1611_; 
wire _abc_41356_new_n1612_; 
wire _abc_41356_new_n1613_; 
wire _abc_41356_new_n1614_; 
wire _abc_41356_new_n1615_; 
wire _abc_41356_new_n1616_; 
wire _abc_41356_new_n1617_; 
wire _abc_41356_new_n1618_; 
wire _abc_41356_new_n1619_; 
wire _abc_41356_new_n1620_; 
wire _abc_41356_new_n1621_; 
wire _abc_41356_new_n1622_; 
wire _abc_41356_new_n1623_; 
wire _abc_41356_new_n1624_; 
wire _abc_41356_new_n1625_; 
wire _abc_41356_new_n1626_; 
wire _abc_41356_new_n1627_; 
wire _abc_41356_new_n1628_; 
wire _abc_41356_new_n1629_; 
wire _abc_41356_new_n1630_; 
wire _abc_41356_new_n1631_; 
wire _abc_41356_new_n1632_; 
wire _abc_41356_new_n1633_; 
wire _abc_41356_new_n1634_; 
wire _abc_41356_new_n1635_; 
wire _abc_41356_new_n1636_; 
wire _abc_41356_new_n1637_; 
wire _abc_41356_new_n1638_; 
wire _abc_41356_new_n1639_; 
wire _abc_41356_new_n1640_; 
wire _abc_41356_new_n1641_; 
wire _abc_41356_new_n1643_; 
wire _abc_41356_new_n1644_; 
wire _abc_41356_new_n1645_; 
wire _abc_41356_new_n1646_; 
wire _abc_41356_new_n1647_; 
wire _abc_41356_new_n1648_; 
wire _abc_41356_new_n1649_; 
wire _abc_41356_new_n1650_; 
wire _abc_41356_new_n1651_; 
wire _abc_41356_new_n1652_; 
wire _abc_41356_new_n1653_; 
wire _abc_41356_new_n1654_; 
wire _abc_41356_new_n1655_; 
wire _abc_41356_new_n1656_; 
wire _abc_41356_new_n1657_; 
wire _abc_41356_new_n1658_; 
wire _abc_41356_new_n1659_; 
wire _abc_41356_new_n1660_; 
wire _abc_41356_new_n1661_; 
wire _abc_41356_new_n1662_; 
wire _abc_41356_new_n1663_; 
wire _abc_41356_new_n1664_; 
wire _abc_41356_new_n1665_; 
wire _abc_41356_new_n1666_; 
wire _abc_41356_new_n1667_; 
wire _abc_41356_new_n1668_; 
wire _abc_41356_new_n1669_; 
wire _abc_41356_new_n1670_; 
wire _abc_41356_new_n1671_; 
wire _abc_41356_new_n1672_; 
wire _abc_41356_new_n1673_; 
wire _abc_41356_new_n1674_; 
wire _abc_41356_new_n1675_; 
wire _abc_41356_new_n1676_; 
wire _abc_41356_new_n1677_; 
wire _abc_41356_new_n1678_; 
wire _abc_41356_new_n1679_; 
wire _abc_41356_new_n1680_; 
wire _abc_41356_new_n1681_; 
wire _abc_41356_new_n1682_; 
wire _abc_41356_new_n1683_; 
wire _abc_41356_new_n1684_; 
wire _abc_41356_new_n1685_; 
wire _abc_41356_new_n1686_; 
wire _abc_41356_new_n1687_; 
wire _abc_41356_new_n1688_; 
wire _abc_41356_new_n1689_; 
wire _abc_41356_new_n1690_; 
wire _abc_41356_new_n1691_; 
wire _abc_41356_new_n1692_; 
wire _abc_41356_new_n1693_; 
wire _abc_41356_new_n1694_; 
wire _abc_41356_new_n1695_; 
wire _abc_41356_new_n1696_; 
wire _abc_41356_new_n1697_; 
wire _abc_41356_new_n1698_; 
wire _abc_41356_new_n1699_; 
wire _abc_41356_new_n1700_; 
wire _abc_41356_new_n1701_; 
wire _abc_41356_new_n1702_; 
wire _abc_41356_new_n1703_; 
wire _abc_41356_new_n1704_; 
wire _abc_41356_new_n1705_; 
wire _abc_41356_new_n1706_; 
wire _abc_41356_new_n1707_; 
wire _abc_41356_new_n1708_; 
wire _abc_41356_new_n1709_; 
wire _abc_41356_new_n1710_; 
wire _abc_41356_new_n1711_; 
wire _abc_41356_new_n1712_; 
wire _abc_41356_new_n1713_; 
wire _abc_41356_new_n1715_; 
wire _abc_41356_new_n1716_; 
wire _abc_41356_new_n1717_; 
wire _abc_41356_new_n1718_; 
wire _abc_41356_new_n1719_; 
wire _abc_41356_new_n1720_; 
wire _abc_41356_new_n1721_; 
wire _abc_41356_new_n1722_; 
wire _abc_41356_new_n1723_; 
wire _abc_41356_new_n1724_; 
wire _abc_41356_new_n1725_; 
wire _abc_41356_new_n1726_; 
wire _abc_41356_new_n1727_; 
wire _abc_41356_new_n1728_; 
wire _abc_41356_new_n1729_; 
wire _abc_41356_new_n1730_; 
wire _abc_41356_new_n1731_; 
wire _abc_41356_new_n1732_; 
wire _abc_41356_new_n1733_; 
wire _abc_41356_new_n1734_; 
wire _abc_41356_new_n1735_; 
wire _abc_41356_new_n1736_; 
wire _abc_41356_new_n1737_; 
wire _abc_41356_new_n1738_; 
wire _abc_41356_new_n1739_; 
wire _abc_41356_new_n1740_; 
wire _abc_41356_new_n1741_; 
wire _abc_41356_new_n1742_; 
wire _abc_41356_new_n1743_; 
wire _abc_41356_new_n1744_; 
wire _abc_41356_new_n1745_; 
wire _abc_41356_new_n1746_; 
wire _abc_41356_new_n1747_; 
wire _abc_41356_new_n1748_; 
wire _abc_41356_new_n1749_; 
wire _abc_41356_new_n1750_; 
wire _abc_41356_new_n1751_; 
wire _abc_41356_new_n1752_; 
wire _abc_41356_new_n1753_; 
wire _abc_41356_new_n1754_; 
wire _abc_41356_new_n1755_; 
wire _abc_41356_new_n1756_; 
wire _abc_41356_new_n1757_; 
wire _abc_41356_new_n1758_; 
wire _abc_41356_new_n1759_; 
wire _abc_41356_new_n1760_; 
wire _abc_41356_new_n1761_; 
wire _abc_41356_new_n1762_; 
wire _abc_41356_new_n1763_; 
wire _abc_41356_new_n1764_; 
wire _abc_41356_new_n1765_; 
wire _abc_41356_new_n1766_; 
wire _abc_41356_new_n1767_; 
wire _abc_41356_new_n1768_; 
wire _abc_41356_new_n1769_; 
wire _abc_41356_new_n1770_; 
wire _abc_41356_new_n1771_; 
wire _abc_41356_new_n1772_; 
wire _abc_41356_new_n1773_; 
wire _abc_41356_new_n1774_; 
wire _abc_41356_new_n1775_; 
wire _abc_41356_new_n1776_; 
wire _abc_41356_new_n1777_; 
wire _abc_41356_new_n1778_; 
wire _abc_41356_new_n1779_; 
wire _abc_41356_new_n1780_; 
wire _abc_41356_new_n1781_; 
wire _abc_41356_new_n1782_; 
wire _abc_41356_new_n1783_; 
wire _abc_41356_new_n1784_; 
wire _abc_41356_new_n1785_; 
wire _abc_41356_new_n1786_; 
wire _abc_41356_new_n1787_; 
wire _abc_41356_new_n1788_; 
wire _abc_41356_new_n1789_; 
wire _abc_41356_new_n1790_; 
wire _abc_41356_new_n1791_; 
wire _abc_41356_new_n1792_; 
wire _abc_41356_new_n1793_; 
wire _abc_41356_new_n1794_; 
wire _abc_41356_new_n1795_; 
wire _abc_41356_new_n1796_; 
wire _abc_41356_new_n1797_; 
wire _abc_41356_new_n1798_; 
wire _abc_41356_new_n1799_; 
wire _abc_41356_new_n1800_; 
wire _abc_41356_new_n1801_; 
wire _abc_41356_new_n1802_; 
wire _abc_41356_new_n1803_; 
wire _abc_41356_new_n1804_; 
wire _abc_41356_new_n1805_; 
wire _abc_41356_new_n1806_; 
wire _abc_41356_new_n1807_; 
wire _abc_41356_new_n1808_; 
wire _abc_41356_new_n1809_; 
wire _abc_41356_new_n1811_; 
wire _abc_41356_new_n1812_; 
wire _abc_41356_new_n1813_; 
wire _abc_41356_new_n1814_; 
wire _abc_41356_new_n1815_; 
wire _abc_41356_new_n1816_; 
wire _abc_41356_new_n1817_; 
wire _abc_41356_new_n1818_; 
wire _abc_41356_new_n1819_; 
wire _abc_41356_new_n1820_; 
wire _abc_41356_new_n1821_; 
wire _abc_41356_new_n1822_; 
wire _abc_41356_new_n1823_; 
wire _abc_41356_new_n1824_; 
wire _abc_41356_new_n1825_; 
wire _abc_41356_new_n1826_; 
wire _abc_41356_new_n1827_; 
wire _abc_41356_new_n1828_; 
wire _abc_41356_new_n1829_; 
wire _abc_41356_new_n1830_; 
wire _abc_41356_new_n1831_; 
wire _abc_41356_new_n1832_; 
wire _abc_41356_new_n1833_; 
wire _abc_41356_new_n1834_; 
wire _abc_41356_new_n1835_; 
wire _abc_41356_new_n1836_; 
wire _abc_41356_new_n1837_; 
wire _abc_41356_new_n1838_; 
wire _abc_41356_new_n1839_; 
wire _abc_41356_new_n1840_; 
wire _abc_41356_new_n1841_; 
wire _abc_41356_new_n1842_; 
wire _abc_41356_new_n1843_; 
wire _abc_41356_new_n1844_; 
wire _abc_41356_new_n1845_; 
wire _abc_41356_new_n1846_; 
wire _abc_41356_new_n1847_; 
wire _abc_41356_new_n1848_; 
wire _abc_41356_new_n1849_; 
wire _abc_41356_new_n1850_; 
wire _abc_41356_new_n1851_; 
wire _abc_41356_new_n1852_; 
wire _abc_41356_new_n1853_; 
wire _abc_41356_new_n1854_; 
wire _abc_41356_new_n1855_; 
wire _abc_41356_new_n1856_; 
wire _abc_41356_new_n1857_; 
wire _abc_41356_new_n1858_; 
wire _abc_41356_new_n1859_; 
wire _abc_41356_new_n1860_; 
wire _abc_41356_new_n1861_; 
wire _abc_41356_new_n1862_; 
wire _abc_41356_new_n1863_; 
wire _abc_41356_new_n1864_; 
wire _abc_41356_new_n1865_; 
wire _abc_41356_new_n1866_; 
wire _abc_41356_new_n1867_; 
wire _abc_41356_new_n1868_; 
wire _abc_41356_new_n1869_; 
wire _abc_41356_new_n1870_; 
wire _abc_41356_new_n1871_; 
wire _abc_41356_new_n1872_; 
wire _abc_41356_new_n1873_; 
wire _abc_41356_new_n1874_; 
wire _abc_41356_new_n1875_; 
wire _abc_41356_new_n1876_; 
wire _abc_41356_new_n1877_; 
wire _abc_41356_new_n1878_; 
wire _abc_41356_new_n1879_; 
wire _abc_41356_new_n1880_; 
wire _abc_41356_new_n1881_; 
wire _abc_41356_new_n1882_; 
wire _abc_41356_new_n1883_; 
wire _abc_41356_new_n1885_; 
wire _abc_41356_new_n1886_; 
wire _abc_41356_new_n1887_; 
wire _abc_41356_new_n1888_; 
wire _abc_41356_new_n1889_; 
wire _abc_41356_new_n1890_; 
wire _abc_41356_new_n1891_; 
wire _abc_41356_new_n1892_; 
wire _abc_41356_new_n1893_; 
wire _abc_41356_new_n1894_; 
wire _abc_41356_new_n1895_; 
wire _abc_41356_new_n1896_; 
wire _abc_41356_new_n1897_; 
wire _abc_41356_new_n1898_; 
wire _abc_41356_new_n1899_; 
wire _abc_41356_new_n1900_; 
wire _abc_41356_new_n1901_; 
wire _abc_41356_new_n1902_; 
wire _abc_41356_new_n1903_; 
wire _abc_41356_new_n1904_; 
wire _abc_41356_new_n1905_; 
wire _abc_41356_new_n1906_; 
wire _abc_41356_new_n1907_; 
wire _abc_41356_new_n1908_; 
wire _abc_41356_new_n1909_; 
wire _abc_41356_new_n1910_; 
wire _abc_41356_new_n1911_; 
wire _abc_41356_new_n1912_; 
wire _abc_41356_new_n1913_; 
wire _abc_41356_new_n1914_; 
wire _abc_41356_new_n1915_; 
wire _abc_41356_new_n1916_; 
wire _abc_41356_new_n1917_; 
wire _abc_41356_new_n1918_; 
wire _abc_41356_new_n1919_; 
wire _abc_41356_new_n1920_; 
wire _abc_41356_new_n1921_; 
wire _abc_41356_new_n1922_; 
wire _abc_41356_new_n1923_; 
wire _abc_41356_new_n1924_; 
wire _abc_41356_new_n1925_; 
wire _abc_41356_new_n1926_; 
wire _abc_41356_new_n1927_; 
wire _abc_41356_new_n1928_; 
wire _abc_41356_new_n1929_; 
wire _abc_41356_new_n1930_; 
wire _abc_41356_new_n1931_; 
wire _abc_41356_new_n1932_; 
wire _abc_41356_new_n1933_; 
wire _abc_41356_new_n1934_; 
wire _abc_41356_new_n1935_; 
wire _abc_41356_new_n1936_; 
wire _abc_41356_new_n1937_; 
wire _abc_41356_new_n1938_; 
wire _abc_41356_new_n1939_; 
wire _abc_41356_new_n1940_; 
wire _abc_41356_new_n1941_; 
wire _abc_41356_new_n1942_; 
wire _abc_41356_new_n1943_; 
wire _abc_41356_new_n1944_; 
wire _abc_41356_new_n1945_; 
wire _abc_41356_new_n1946_; 
wire _abc_41356_new_n1947_; 
wire _abc_41356_new_n1948_; 
wire _abc_41356_new_n1949_; 
wire _abc_41356_new_n1950_; 
wire _abc_41356_new_n1952_; 
wire _abc_41356_new_n1953_; 
wire _abc_41356_new_n1954_; 
wire _abc_41356_new_n1955_; 
wire _abc_41356_new_n1956_; 
wire _abc_41356_new_n1957_; 
wire _abc_41356_new_n1958_; 
wire _abc_41356_new_n1959_; 
wire _abc_41356_new_n1960_; 
wire _abc_41356_new_n1961_; 
wire _abc_41356_new_n1962_; 
wire _abc_41356_new_n1963_; 
wire _abc_41356_new_n1964_; 
wire _abc_41356_new_n1965_; 
wire _abc_41356_new_n1966_; 
wire _abc_41356_new_n1967_; 
wire _abc_41356_new_n1968_; 
wire _abc_41356_new_n1969_; 
wire _abc_41356_new_n1970_; 
wire _abc_41356_new_n1971_; 
wire _abc_41356_new_n1972_; 
wire _abc_41356_new_n1973_; 
wire _abc_41356_new_n1974_; 
wire _abc_41356_new_n1975_; 
wire _abc_41356_new_n1976_; 
wire _abc_41356_new_n1977_; 
wire _abc_41356_new_n1978_; 
wire _abc_41356_new_n1979_; 
wire _abc_41356_new_n1980_; 
wire _abc_41356_new_n1981_; 
wire _abc_41356_new_n1982_; 
wire _abc_41356_new_n1983_; 
wire _abc_41356_new_n1984_; 
wire _abc_41356_new_n1985_; 
wire _abc_41356_new_n1986_; 
wire _abc_41356_new_n1987_; 
wire _abc_41356_new_n1988_; 
wire _abc_41356_new_n1989_; 
wire _abc_41356_new_n1990_; 
wire _abc_41356_new_n1991_; 
wire _abc_41356_new_n1992_; 
wire _abc_41356_new_n1993_; 
wire _abc_41356_new_n1994_; 
wire _abc_41356_new_n1995_; 
wire _abc_41356_new_n1996_; 
wire _abc_41356_new_n1997_; 
wire _abc_41356_new_n1998_; 
wire _abc_41356_new_n1999_; 
wire _abc_41356_new_n2000_; 
wire _abc_41356_new_n2001_; 
wire _abc_41356_new_n2002_; 
wire _abc_41356_new_n2003_; 
wire _abc_41356_new_n2004_; 
wire _abc_41356_new_n2005_; 
wire _abc_41356_new_n2006_; 
wire _abc_41356_new_n2007_; 
wire _abc_41356_new_n2008_; 
wire _abc_41356_new_n2009_; 
wire _abc_41356_new_n2010_; 
wire _abc_41356_new_n2011_; 
wire _abc_41356_new_n2012_; 
wire _abc_41356_new_n2013_; 
wire _abc_41356_new_n2014_; 
wire _abc_41356_new_n2015_; 
wire _abc_41356_new_n2016_; 
wire _abc_41356_new_n2017_; 
wire _abc_41356_new_n2018_; 
wire _abc_41356_new_n2020_; 
wire _abc_41356_new_n2021_; 
wire _abc_41356_new_n2022_; 
wire _abc_41356_new_n2023_; 
wire _abc_41356_new_n2024_; 
wire _abc_41356_new_n2025_; 
wire _abc_41356_new_n2026_; 
wire _abc_41356_new_n2027_; 
wire _abc_41356_new_n2028_; 
wire _abc_41356_new_n2029_; 
wire _abc_41356_new_n2030_; 
wire _abc_41356_new_n2031_; 
wire _abc_41356_new_n2032_; 
wire _abc_41356_new_n2033_; 
wire _abc_41356_new_n2034_; 
wire _abc_41356_new_n2035_; 
wire _abc_41356_new_n2036_; 
wire _abc_41356_new_n2037_; 
wire _abc_41356_new_n2038_; 
wire _abc_41356_new_n2039_; 
wire _abc_41356_new_n2040_; 
wire _abc_41356_new_n2041_; 
wire _abc_41356_new_n2042_; 
wire _abc_41356_new_n2043_; 
wire _abc_41356_new_n2044_; 
wire _abc_41356_new_n2045_; 
wire _abc_41356_new_n2046_; 
wire _abc_41356_new_n2047_; 
wire _abc_41356_new_n2048_; 
wire _abc_41356_new_n2049_; 
wire _abc_41356_new_n2050_; 
wire _abc_41356_new_n2051_; 
wire _abc_41356_new_n2052_; 
wire _abc_41356_new_n2053_; 
wire _abc_41356_new_n2054_; 
wire _abc_41356_new_n2055_; 
wire _abc_41356_new_n2056_; 
wire _abc_41356_new_n2057_; 
wire _abc_41356_new_n2058_; 
wire _abc_41356_new_n2059_; 
wire _abc_41356_new_n2060_; 
wire _abc_41356_new_n2061_; 
wire _abc_41356_new_n2062_; 
wire _abc_41356_new_n2063_; 
wire _abc_41356_new_n2064_; 
wire _abc_41356_new_n2065_; 
wire _abc_41356_new_n2066_; 
wire _abc_41356_new_n2067_; 
wire _abc_41356_new_n2068_; 
wire _abc_41356_new_n2069_; 
wire _abc_41356_new_n2070_; 
wire _abc_41356_new_n2071_; 
wire _abc_41356_new_n2072_; 
wire _abc_41356_new_n2073_; 
wire _abc_41356_new_n2074_; 
wire _abc_41356_new_n2075_; 
wire _abc_41356_new_n2076_; 
wire _abc_41356_new_n2077_; 
wire _abc_41356_new_n2078_; 
wire _abc_41356_new_n2079_; 
wire _abc_41356_new_n2080_; 
wire _abc_41356_new_n2081_; 
wire _abc_41356_new_n2082_; 
wire _abc_41356_new_n2083_; 
wire _abc_41356_new_n2084_; 
wire _abc_41356_new_n2085_; 
wire _abc_41356_new_n2086_; 
wire _abc_41356_new_n2087_; 
wire _abc_41356_new_n2088_; 
wire _abc_41356_new_n2089_; 
wire _abc_41356_new_n2090_; 
wire _abc_41356_new_n2091_; 
wire _abc_41356_new_n2092_; 
wire _abc_41356_new_n2093_; 
wire _abc_41356_new_n2094_; 
wire _abc_41356_new_n2095_; 
wire _abc_41356_new_n2096_; 
wire _abc_41356_new_n2097_; 
wire _abc_41356_new_n2098_; 
wire _abc_41356_new_n2099_; 
wire _abc_41356_new_n2100_; 
wire _abc_41356_new_n2101_; 
wire _abc_41356_new_n2103_; 
wire _abc_41356_new_n2104_; 
wire _abc_41356_new_n2105_; 
wire _abc_41356_new_n2106_; 
wire _abc_41356_new_n2107_; 
wire _abc_41356_new_n2108_; 
wire _abc_41356_new_n2109_; 
wire _abc_41356_new_n2110_; 
wire _abc_41356_new_n2111_; 
wire _abc_41356_new_n2112_; 
wire _abc_41356_new_n2113_; 
wire _abc_41356_new_n2114_; 
wire _abc_41356_new_n2115_; 
wire _abc_41356_new_n2116_; 
wire _abc_41356_new_n2117_; 
wire _abc_41356_new_n2118_; 
wire _abc_41356_new_n2119_; 
wire _abc_41356_new_n2120_; 
wire _abc_41356_new_n2121_; 
wire _abc_41356_new_n2122_; 
wire _abc_41356_new_n2123_; 
wire _abc_41356_new_n2124_; 
wire _abc_41356_new_n2125_; 
wire _abc_41356_new_n2126_; 
wire _abc_41356_new_n2127_; 
wire _abc_41356_new_n2128_; 
wire _abc_41356_new_n2129_; 
wire _abc_41356_new_n2130_; 
wire _abc_41356_new_n2131_; 
wire _abc_41356_new_n2132_; 
wire _abc_41356_new_n2133_; 
wire _abc_41356_new_n2134_; 
wire _abc_41356_new_n2135_; 
wire _abc_41356_new_n2136_; 
wire _abc_41356_new_n2137_; 
wire _abc_41356_new_n2138_; 
wire _abc_41356_new_n2139_; 
wire _abc_41356_new_n2140_; 
wire _abc_41356_new_n2141_; 
wire _abc_41356_new_n2143_; 
wire _abc_41356_new_n2144_; 
wire _abc_41356_new_n2145_; 
wire _abc_41356_new_n2146_; 
wire _abc_41356_new_n2147_; 
wire _abc_41356_new_n2148_; 
wire _abc_41356_new_n2149_; 
wire _abc_41356_new_n2150_; 
wire _abc_41356_new_n2151_; 
wire _abc_41356_new_n2152_; 
wire _abc_41356_new_n2153_; 
wire _abc_41356_new_n2154_; 
wire _abc_41356_new_n2155_; 
wire _abc_41356_new_n2156_; 
wire _abc_41356_new_n2157_; 
wire _abc_41356_new_n2158_; 
wire _abc_41356_new_n2159_; 
wire _abc_41356_new_n2160_; 
wire _abc_41356_new_n2161_; 
wire _abc_41356_new_n2162_; 
wire _abc_41356_new_n2163_; 
wire _abc_41356_new_n2164_; 
wire _abc_41356_new_n2165_; 
wire _abc_41356_new_n2166_; 
wire _abc_41356_new_n2167_; 
wire _abc_41356_new_n2168_; 
wire _abc_41356_new_n2169_; 
wire _abc_41356_new_n2170_; 
wire _abc_41356_new_n2171_; 
wire _abc_41356_new_n2172_; 
wire _abc_41356_new_n2173_; 
wire _abc_41356_new_n2174_; 
wire _abc_41356_new_n2175_; 
wire _abc_41356_new_n2176_; 
wire _abc_41356_new_n2177_; 
wire _abc_41356_new_n2178_; 
wire _abc_41356_new_n2179_; 
wire _abc_41356_new_n2180_; 
wire _abc_41356_new_n2181_; 
wire _abc_41356_new_n2183_; 
wire _abc_41356_new_n2184_; 
wire _abc_41356_new_n2185_; 
wire _abc_41356_new_n2186_; 
wire _abc_41356_new_n2187_; 
wire _abc_41356_new_n2188_; 
wire _abc_41356_new_n2189_; 
wire _abc_41356_new_n2190_; 
wire _abc_41356_new_n2191_; 
wire _abc_41356_new_n2192_; 
wire _abc_41356_new_n2193_; 
wire _abc_41356_new_n2194_; 
wire _abc_41356_new_n2195_; 
wire _abc_41356_new_n2196_; 
wire _abc_41356_new_n2197_; 
wire _abc_41356_new_n2198_; 
wire _abc_41356_new_n2199_; 
wire _abc_41356_new_n2200_; 
wire _abc_41356_new_n2201_; 
wire _abc_41356_new_n2202_; 
wire _abc_41356_new_n2203_; 
wire _abc_41356_new_n2204_; 
wire _abc_41356_new_n2205_; 
wire _abc_41356_new_n2206_; 
wire _abc_41356_new_n2207_; 
wire _abc_41356_new_n2208_; 
wire _abc_41356_new_n2209_; 
wire _abc_41356_new_n2210_; 
wire _abc_41356_new_n2211_; 
wire _abc_41356_new_n2212_; 
wire _abc_41356_new_n2213_; 
wire _abc_41356_new_n2214_; 
wire _abc_41356_new_n2215_; 
wire _abc_41356_new_n2216_; 
wire _abc_41356_new_n2217_; 
wire _abc_41356_new_n2218_; 
wire _abc_41356_new_n2219_; 
wire _abc_41356_new_n2221_; 
wire _abc_41356_new_n2222_; 
wire _abc_41356_new_n2223_; 
wire _abc_41356_new_n2224_; 
wire _abc_41356_new_n2225_; 
wire _abc_41356_new_n2226_; 
wire _abc_41356_new_n2227_; 
wire _abc_41356_new_n2228_; 
wire _abc_41356_new_n2229_; 
wire _abc_41356_new_n2230_; 
wire _abc_41356_new_n2231_; 
wire _abc_41356_new_n2232_; 
wire _abc_41356_new_n2233_; 
wire _abc_41356_new_n2234_; 
wire _abc_41356_new_n2235_; 
wire _abc_41356_new_n2236_; 
wire _abc_41356_new_n2237_; 
wire _abc_41356_new_n2238_; 
wire _abc_41356_new_n2239_; 
wire _abc_41356_new_n2240_; 
wire _abc_41356_new_n2241_; 
wire _abc_41356_new_n2242_; 
wire _abc_41356_new_n2243_; 
wire _abc_41356_new_n2244_; 
wire _abc_41356_new_n2245_; 
wire _abc_41356_new_n2246_; 
wire _abc_41356_new_n2247_; 
wire _abc_41356_new_n2248_; 
wire _abc_41356_new_n2249_; 
wire _abc_41356_new_n2250_; 
wire _abc_41356_new_n2251_; 
wire _abc_41356_new_n2252_; 
wire _abc_41356_new_n2253_; 
wire _abc_41356_new_n2254_; 
wire _abc_41356_new_n2255_; 
wire _abc_41356_new_n2256_; 
wire _abc_41356_new_n2257_; 
wire _abc_41356_new_n2258_; 
wire _abc_41356_new_n2259_; 
wire _abc_41356_new_n2261_; 
wire _abc_41356_new_n2262_; 
wire _abc_41356_new_n2263_; 
wire _abc_41356_new_n2264_; 
wire _abc_41356_new_n2265_; 
wire _abc_41356_new_n2266_; 
wire _abc_41356_new_n2267_; 
wire _abc_41356_new_n2268_; 
wire _abc_41356_new_n2269_; 
wire _abc_41356_new_n2270_; 
wire _abc_41356_new_n2271_; 
wire _abc_41356_new_n2272_; 
wire _abc_41356_new_n2273_; 
wire _abc_41356_new_n2274_; 
wire _abc_41356_new_n2275_; 
wire _abc_41356_new_n2276_; 
wire _abc_41356_new_n2277_; 
wire _abc_41356_new_n2278_; 
wire _abc_41356_new_n2279_; 
wire _abc_41356_new_n2280_; 
wire _abc_41356_new_n2281_; 
wire _abc_41356_new_n2282_; 
wire _abc_41356_new_n2283_; 
wire _abc_41356_new_n2284_; 
wire _abc_41356_new_n2285_; 
wire _abc_41356_new_n2286_; 
wire _abc_41356_new_n2287_; 
wire _abc_41356_new_n2288_; 
wire _abc_41356_new_n2289_; 
wire _abc_41356_new_n2290_; 
wire _abc_41356_new_n2291_; 
wire _abc_41356_new_n2292_; 
wire _abc_41356_new_n2293_; 
wire _abc_41356_new_n2294_; 
wire _abc_41356_new_n2295_; 
wire _abc_41356_new_n2296_; 
wire _abc_41356_new_n2297_; 
wire _abc_41356_new_n2299_; 
wire _abc_41356_new_n2300_; 
wire _abc_41356_new_n2301_; 
wire _abc_41356_new_n2302_; 
wire _abc_41356_new_n2303_; 
wire _abc_41356_new_n2304_; 
wire _abc_41356_new_n2305_; 
wire _abc_41356_new_n2306_; 
wire _abc_41356_new_n2307_; 
wire _abc_41356_new_n2308_; 
wire _abc_41356_new_n2309_; 
wire _abc_41356_new_n2310_; 
wire _abc_41356_new_n2311_; 
wire _abc_41356_new_n2312_; 
wire _abc_41356_new_n2313_; 
wire _abc_41356_new_n2314_; 
wire _abc_41356_new_n2315_; 
wire _abc_41356_new_n2316_; 
wire _abc_41356_new_n2317_; 
wire _abc_41356_new_n2318_; 
wire _abc_41356_new_n2319_; 
wire _abc_41356_new_n2320_; 
wire _abc_41356_new_n2321_; 
wire _abc_41356_new_n2322_; 
wire _abc_41356_new_n2323_; 
wire _abc_41356_new_n2324_; 
wire _abc_41356_new_n2325_; 
wire _abc_41356_new_n2326_; 
wire _abc_41356_new_n2327_; 
wire _abc_41356_new_n2328_; 
wire _abc_41356_new_n2329_; 
wire _abc_41356_new_n2330_; 
wire _abc_41356_new_n2331_; 
wire _abc_41356_new_n2332_; 
wire _abc_41356_new_n2333_; 
wire _abc_41356_new_n2334_; 
wire _abc_41356_new_n2335_; 
wire _abc_41356_new_n2337_; 
wire _abc_41356_new_n2338_; 
wire _abc_41356_new_n2339_; 
wire _abc_41356_new_n2340_; 
wire _abc_41356_new_n2341_; 
wire _abc_41356_new_n2342_; 
wire _abc_41356_new_n2343_; 
wire _abc_41356_new_n2344_; 
wire _abc_41356_new_n2345_; 
wire _abc_41356_new_n2346_; 
wire _abc_41356_new_n2347_; 
wire _abc_41356_new_n2348_; 
wire _abc_41356_new_n2349_; 
wire _abc_41356_new_n2350_; 
wire _abc_41356_new_n2351_; 
wire _abc_41356_new_n2352_; 
wire _abc_41356_new_n2353_; 
wire _abc_41356_new_n2354_; 
wire _abc_41356_new_n2355_; 
wire _abc_41356_new_n2356_; 
wire _abc_41356_new_n2357_; 
wire _abc_41356_new_n2358_; 
wire _abc_41356_new_n2359_; 
wire _abc_41356_new_n2360_; 
wire _abc_41356_new_n2361_; 
wire _abc_41356_new_n2362_; 
wire _abc_41356_new_n2363_; 
wire _abc_41356_new_n2364_; 
wire _abc_41356_new_n2365_; 
wire _abc_41356_new_n2366_; 
wire _abc_41356_new_n2367_; 
wire _abc_41356_new_n2368_; 
wire _abc_41356_new_n2369_; 
wire _abc_41356_new_n2370_; 
wire _abc_41356_new_n2371_; 
wire _abc_41356_new_n2372_; 
wire _abc_41356_new_n2373_; 
wire _abc_41356_new_n2375_; 
wire _abc_41356_new_n2376_; 
wire _abc_41356_new_n2377_; 
wire _abc_41356_new_n2378_; 
wire _abc_41356_new_n2379_; 
wire _abc_41356_new_n2380_; 
wire _abc_41356_new_n2381_; 
wire _abc_41356_new_n2382_; 
wire _abc_41356_new_n2383_; 
wire _abc_41356_new_n2384_; 
wire _abc_41356_new_n2385_; 
wire _abc_41356_new_n2386_; 
wire _abc_41356_new_n2387_; 
wire _abc_41356_new_n2388_; 
wire _abc_41356_new_n2389_; 
wire _abc_41356_new_n2390_; 
wire _abc_41356_new_n2391_; 
wire _abc_41356_new_n2392_; 
wire _abc_41356_new_n2393_; 
wire _abc_41356_new_n2394_; 
wire _abc_41356_new_n2395_; 
wire _abc_41356_new_n2396_; 
wire _abc_41356_new_n2397_; 
wire _abc_41356_new_n2398_; 
wire _abc_41356_new_n2399_; 
wire _abc_41356_new_n2400_; 
wire _abc_41356_new_n2401_; 
wire _abc_41356_new_n2403_; 
wire _abc_41356_new_n2404_; 
wire _abc_41356_new_n2405_; 
wire _abc_41356_new_n2406_; 
wire _abc_41356_new_n2407_; 
wire _abc_41356_new_n2408_; 
wire _abc_41356_new_n2409_; 
wire _abc_41356_new_n2410_; 
wire _abc_41356_new_n2411_; 
wire _abc_41356_new_n2412_; 
wire _abc_41356_new_n2413_; 
wire _abc_41356_new_n2414_; 
wire _abc_41356_new_n2415_; 
wire _abc_41356_new_n2416_; 
wire _abc_41356_new_n2417_; 
wire _abc_41356_new_n2418_; 
wire _abc_41356_new_n2419_; 
wire _abc_41356_new_n2420_; 
wire _abc_41356_new_n2421_; 
wire _abc_41356_new_n2422_; 
wire _abc_41356_new_n2423_; 
wire _abc_41356_new_n2424_; 
wire _abc_41356_new_n2425_; 
wire _abc_41356_new_n2426_; 
wire _abc_41356_new_n2428_; 
wire _abc_41356_new_n2429_; 
wire _abc_41356_new_n2430_; 
wire _abc_41356_new_n2431_; 
wire _abc_41356_new_n2432_; 
wire _abc_41356_new_n2433_; 
wire _abc_41356_new_n2434_; 
wire _abc_41356_new_n2435_; 
wire _abc_41356_new_n2436_; 
wire _abc_41356_new_n2437_; 
wire _abc_41356_new_n2438_; 
wire _abc_41356_new_n2439_; 
wire _abc_41356_new_n2440_; 
wire _abc_41356_new_n2441_; 
wire _abc_41356_new_n2442_; 
wire _abc_41356_new_n2443_; 
wire _abc_41356_new_n2444_; 
wire _abc_41356_new_n2445_; 
wire _abc_41356_new_n2446_; 
wire _abc_41356_new_n2448_; 
wire _abc_41356_new_n2449_; 
wire _abc_41356_new_n2450_; 
wire _abc_41356_new_n2451_; 
wire _abc_41356_new_n2452_; 
wire _abc_41356_new_n2453_; 
wire _abc_41356_new_n2454_; 
wire _abc_41356_new_n2455_; 
wire _abc_41356_new_n2456_; 
wire _abc_41356_new_n2457_; 
wire _abc_41356_new_n2458_; 
wire _abc_41356_new_n2459_; 
wire _abc_41356_new_n2460_; 
wire _abc_41356_new_n2461_; 
wire _abc_41356_new_n2462_; 
wire _abc_41356_new_n2463_; 
wire _abc_41356_new_n2464_; 
wire _abc_41356_new_n2465_; 
wire _abc_41356_new_n2466_; 
wire _abc_41356_new_n2468_; 
wire _abc_41356_new_n2469_; 
wire _abc_41356_new_n2470_; 
wire _abc_41356_new_n2471_; 
wire _abc_41356_new_n2472_; 
wire _abc_41356_new_n2473_; 
wire _abc_41356_new_n2474_; 
wire _abc_41356_new_n2475_; 
wire _abc_41356_new_n2476_; 
wire _abc_41356_new_n2477_; 
wire _abc_41356_new_n2478_; 
wire _abc_41356_new_n2479_; 
wire _abc_41356_new_n2480_; 
wire _abc_41356_new_n2481_; 
wire _abc_41356_new_n2482_; 
wire _abc_41356_new_n2483_; 
wire _abc_41356_new_n2484_; 
wire _abc_41356_new_n2485_; 
wire _abc_41356_new_n2486_; 
wire _abc_41356_new_n2487_; 
wire _abc_41356_new_n2489_; 
wire _abc_41356_new_n2490_; 
wire _abc_41356_new_n2491_; 
wire _abc_41356_new_n2492_; 
wire _abc_41356_new_n2493_; 
wire _abc_41356_new_n2494_; 
wire _abc_41356_new_n2495_; 
wire _abc_41356_new_n2496_; 
wire _abc_41356_new_n2497_; 
wire _abc_41356_new_n2498_; 
wire _abc_41356_new_n2499_; 
wire _abc_41356_new_n2500_; 
wire _abc_41356_new_n2501_; 
wire _abc_41356_new_n2502_; 
wire _abc_41356_new_n2503_; 
wire _abc_41356_new_n2504_; 
wire _abc_41356_new_n2505_; 
wire _abc_41356_new_n2506_; 
wire _abc_41356_new_n2507_; 
wire _abc_41356_new_n2509_; 
wire _abc_41356_new_n2510_; 
wire _abc_41356_new_n2511_; 
wire _abc_41356_new_n2512_; 
wire _abc_41356_new_n2513_; 
wire _abc_41356_new_n2514_; 
wire _abc_41356_new_n2515_; 
wire _abc_41356_new_n2516_; 
wire _abc_41356_new_n2517_; 
wire _abc_41356_new_n2518_; 
wire _abc_41356_new_n2519_; 
wire _abc_41356_new_n2520_; 
wire _abc_41356_new_n2521_; 
wire _abc_41356_new_n2522_; 
wire _abc_41356_new_n2523_; 
wire _abc_41356_new_n2524_; 
wire _abc_41356_new_n2525_; 
wire _abc_41356_new_n2526_; 
wire _abc_41356_new_n2527_; 
wire _abc_41356_new_n2529_; 
wire _abc_41356_new_n2530_; 
wire _abc_41356_new_n2531_; 
wire _abc_41356_new_n2532_; 
wire _abc_41356_new_n2533_; 
wire _abc_41356_new_n2534_; 
wire _abc_41356_new_n2535_; 
wire _abc_41356_new_n2536_; 
wire _abc_41356_new_n2537_; 
wire _abc_41356_new_n2538_; 
wire _abc_41356_new_n2539_; 
wire _abc_41356_new_n2540_; 
wire _abc_41356_new_n2541_; 
wire _abc_41356_new_n2542_; 
wire _abc_41356_new_n2543_; 
wire _abc_41356_new_n2544_; 
wire _abc_41356_new_n2545_; 
wire _abc_41356_new_n2546_; 
wire _abc_41356_new_n2547_; 
wire _abc_41356_new_n2549_; 
wire _abc_41356_new_n2550_; 
wire _abc_41356_new_n2551_; 
wire _abc_41356_new_n2552_; 
wire _abc_41356_new_n2553_; 
wire _abc_41356_new_n2554_; 
wire _abc_41356_new_n2555_; 
wire _abc_41356_new_n2556_; 
wire _abc_41356_new_n2557_; 
wire _abc_41356_new_n2558_; 
wire _abc_41356_new_n2559_; 
wire _abc_41356_new_n2560_; 
wire _abc_41356_new_n2561_; 
wire _abc_41356_new_n2563_; 
wire _abc_41356_new_n2564_; 
wire _abc_41356_new_n2565_; 
wire _abc_41356_new_n2566_; 
wire _abc_41356_new_n2567_; 
wire _abc_41356_new_n2568_; 
wire _abc_41356_new_n2569_; 
wire _abc_41356_new_n2570_; 
wire _abc_41356_new_n2571_; 
wire _abc_41356_new_n2572_; 
wire _abc_41356_new_n2573_; 
wire _abc_41356_new_n2574_; 
wire _abc_41356_new_n2576_; 
wire _abc_41356_new_n2577_; 
wire _abc_41356_new_n2578_; 
wire _abc_41356_new_n2579_; 
wire _abc_41356_new_n2580_; 
wire _abc_41356_new_n2581_; 
wire _abc_41356_new_n2582_; 
wire _abc_41356_new_n2583_; 
wire _abc_41356_new_n2584_; 
wire _abc_41356_new_n2585_; 
wire _abc_41356_new_n2586_; 
wire _abc_41356_new_n2587_; 
wire _abc_41356_new_n2588_; 
wire _abc_41356_new_n2589_; 
wire _abc_41356_new_n2590_; 
wire _abc_41356_new_n2592_; 
wire _abc_41356_new_n2593_; 
wire _abc_41356_new_n2594_; 
wire _abc_41356_new_n2595_; 
wire _abc_41356_new_n2596_; 
wire _abc_41356_new_n2597_; 
wire _abc_41356_new_n2598_; 
wire _abc_41356_new_n2599_; 
wire _abc_41356_new_n2600_; 
wire _abc_41356_new_n2601_; 
wire _abc_41356_new_n2602_; 
wire _abc_41356_new_n2603_; 
wire _abc_41356_new_n2604_; 
wire _abc_41356_new_n2605_; 
wire _abc_41356_new_n2606_; 
wire _abc_41356_new_n2608_; 
wire _abc_41356_new_n2609_; 
wire _abc_41356_new_n2610_; 
wire _abc_41356_new_n2611_; 
wire _abc_41356_new_n2612_; 
wire _abc_41356_new_n2613_; 
wire _abc_41356_new_n2614_; 
wire _abc_41356_new_n2615_; 
wire _abc_41356_new_n2616_; 
wire _abc_41356_new_n2617_; 
wire _abc_41356_new_n2618_; 
wire _abc_41356_new_n2619_; 
wire _abc_41356_new_n2620_; 
wire _abc_41356_new_n2621_; 
wire _abc_41356_new_n2622_; 
wire _abc_41356_new_n2624_; 
wire _abc_41356_new_n2625_; 
wire _abc_41356_new_n2626_; 
wire _abc_41356_new_n2627_; 
wire _abc_41356_new_n2628_; 
wire _abc_41356_new_n2629_; 
wire _abc_41356_new_n2630_; 
wire _abc_41356_new_n2631_; 
wire _abc_41356_new_n2632_; 
wire _abc_41356_new_n2633_; 
wire _abc_41356_new_n2634_; 
wire _abc_41356_new_n2635_; 
wire _abc_41356_new_n2636_; 
wire _abc_41356_new_n2637_; 
wire _abc_41356_new_n2638_; 
wire _abc_41356_new_n2640_; 
wire _abc_41356_new_n2641_; 
wire _abc_41356_new_n2642_; 
wire _abc_41356_new_n2643_; 
wire _abc_41356_new_n2644_; 
wire _abc_41356_new_n2645_; 
wire _abc_41356_new_n2646_; 
wire _abc_41356_new_n2647_; 
wire _abc_41356_new_n2648_; 
wire _abc_41356_new_n2649_; 
wire _abc_41356_new_n2650_; 
wire _abc_41356_new_n2651_; 
wire _abc_41356_new_n2652_; 
wire _abc_41356_new_n2653_; 
wire _abc_41356_new_n2654_; 
wire _abc_41356_new_n2656_; 
wire _abc_41356_new_n2657_; 
wire _abc_41356_new_n2658_; 
wire _abc_41356_new_n2659_; 
wire _abc_41356_new_n2660_; 
wire _abc_41356_new_n2661_; 
wire _abc_41356_new_n2662_; 
wire _abc_41356_new_n2663_; 
wire _abc_41356_new_n2664_; 
wire _abc_41356_new_n2665_; 
wire _abc_41356_new_n2666_; 
wire _abc_41356_new_n2667_; 
wire _abc_41356_new_n2668_; 
wire _abc_41356_new_n2669_; 
wire _abc_41356_new_n2671_; 
wire _abc_41356_new_n2672_; 
wire _abc_41356_new_n2673_; 
wire _abc_41356_new_n2674_; 
wire _abc_41356_new_n2676_; 
wire _abc_41356_new_n2677_; 
wire _abc_41356_new_n2679_; 
wire _abc_41356_new_n2680_; 
wire _abc_41356_new_n2682_; 
wire _abc_41356_new_n2683_; 
wire _abc_41356_new_n2685_; 
wire _abc_41356_new_n2686_; 
wire _abc_41356_new_n2688_; 
wire _abc_41356_new_n2689_; 
wire _abc_41356_new_n2691_; 
wire _abc_41356_new_n2692_; 
wire _abc_41356_new_n2694_; 
wire _abc_41356_new_n2695_; 
wire _abc_41356_new_n2697_; 
wire _abc_41356_new_n2698_; 
wire _abc_41356_new_n2699_; 
wire _abc_41356_new_n2700_; 
wire _abc_41356_new_n2701_; 
wire _abc_41356_new_n2702_; 
wire _abc_41356_new_n2703_; 
wire _abc_41356_new_n2704_; 
wire _abc_41356_new_n2705_; 
wire _abc_41356_new_n2706_; 
wire _abc_41356_new_n2707_; 
wire _abc_41356_new_n2708_; 
wire _abc_41356_new_n2709_; 
wire _abc_41356_new_n2710_; 
wire _abc_41356_new_n2711_; 
wire _abc_41356_new_n2712_; 
wire _abc_41356_new_n2713_; 
wire _abc_41356_new_n2714_; 
wire _abc_41356_new_n2715_; 
wire _abc_41356_new_n2716_; 
wire _abc_41356_new_n2717_; 
wire _abc_41356_new_n2719_; 
wire _abc_41356_new_n2720_; 
wire _abc_41356_new_n2721_; 
wire _abc_41356_new_n2722_; 
wire _abc_41356_new_n2723_; 
wire _abc_41356_new_n2724_; 
wire _abc_41356_new_n2725_; 
wire _abc_41356_new_n2726_; 
wire _abc_41356_new_n2727_; 
wire _abc_41356_new_n2728_; 
wire _abc_41356_new_n2729_; 
wire _abc_41356_new_n2730_; 
wire _abc_41356_new_n2731_; 
wire _abc_41356_new_n2732_; 
wire _abc_41356_new_n2733_; 
wire _abc_41356_new_n2734_; 
wire _abc_41356_new_n2735_; 
wire _abc_41356_new_n2736_; 
wire _abc_41356_new_n2737_; 
wire _abc_41356_new_n2739_; 
wire _abc_41356_new_n2740_; 
wire _abc_41356_new_n2741_; 
wire _abc_41356_new_n2742_; 
wire _abc_41356_new_n2743_; 
wire _abc_41356_new_n2744_; 
wire _abc_41356_new_n2745_; 
wire _abc_41356_new_n2746_; 
wire _abc_41356_new_n2747_; 
wire _abc_41356_new_n2748_; 
wire _abc_41356_new_n2749_; 
wire _abc_41356_new_n2750_; 
wire _abc_41356_new_n2751_; 
wire _abc_41356_new_n2752_; 
wire _abc_41356_new_n2753_; 
wire _abc_41356_new_n2754_; 
wire _abc_41356_new_n2755_; 
wire _abc_41356_new_n2756_; 
wire _abc_41356_new_n2757_; 
wire _abc_41356_new_n2759_; 
wire _abc_41356_new_n2760_; 
wire _abc_41356_new_n2761_; 
wire _abc_41356_new_n2762_; 
wire _abc_41356_new_n2763_; 
wire _abc_41356_new_n2764_; 
wire _abc_41356_new_n2765_; 
wire _abc_41356_new_n2766_; 
wire _abc_41356_new_n2767_; 
wire _abc_41356_new_n2768_; 
wire _abc_41356_new_n2769_; 
wire _abc_41356_new_n2770_; 
wire _abc_41356_new_n2771_; 
wire _abc_41356_new_n2772_; 
wire _abc_41356_new_n2773_; 
wire _abc_41356_new_n2774_; 
wire _abc_41356_new_n2775_; 
wire _abc_41356_new_n2776_; 
wire _abc_41356_new_n2777_; 
wire _abc_41356_new_n2778_; 
wire _abc_41356_new_n2779_; 
wire _abc_41356_new_n2781_; 
wire _abc_41356_new_n2782_; 
wire _abc_41356_new_n2783_; 
wire _abc_41356_new_n2784_; 
wire _abc_41356_new_n2785_; 
wire _abc_41356_new_n2786_; 
wire _abc_41356_new_n2787_; 
wire _abc_41356_new_n2788_; 
wire _abc_41356_new_n2789_; 
wire _abc_41356_new_n2790_; 
wire _abc_41356_new_n2791_; 
wire _abc_41356_new_n2792_; 
wire _abc_41356_new_n2793_; 
wire _abc_41356_new_n2794_; 
wire _abc_41356_new_n2795_; 
wire _abc_41356_new_n2796_; 
wire _abc_41356_new_n2797_; 
wire _abc_41356_new_n2798_; 
wire _abc_41356_new_n2799_; 
wire _abc_41356_new_n2800_; 
wire _abc_41356_new_n2801_; 
wire _abc_41356_new_n2803_; 
wire _abc_41356_new_n2804_; 
wire _abc_41356_new_n2805_; 
wire _abc_41356_new_n2806_; 
wire _abc_41356_new_n2807_; 
wire _abc_41356_new_n2808_; 
wire _abc_41356_new_n2809_; 
wire _abc_41356_new_n2810_; 
wire _abc_41356_new_n2811_; 
wire _abc_41356_new_n2812_; 
wire _abc_41356_new_n2813_; 
wire _abc_41356_new_n2814_; 
wire _abc_41356_new_n2815_; 
wire _abc_41356_new_n2816_; 
wire _abc_41356_new_n2817_; 
wire _abc_41356_new_n2818_; 
wire _abc_41356_new_n2819_; 
wire _abc_41356_new_n2820_; 
wire _abc_41356_new_n2821_; 
wire _abc_41356_new_n2822_; 
wire _abc_41356_new_n2823_; 
wire _abc_41356_new_n2825_; 
wire _abc_41356_new_n2826_; 
wire _abc_41356_new_n2827_; 
wire _abc_41356_new_n2828_; 
wire _abc_41356_new_n2829_; 
wire _abc_41356_new_n2830_; 
wire _abc_41356_new_n2831_; 
wire _abc_41356_new_n2832_; 
wire _abc_41356_new_n2833_; 
wire _abc_41356_new_n2834_; 
wire _abc_41356_new_n2835_; 
wire _abc_41356_new_n2836_; 
wire _abc_41356_new_n2837_; 
wire _abc_41356_new_n2838_; 
wire _abc_41356_new_n2839_; 
wire _abc_41356_new_n2840_; 
wire _abc_41356_new_n2841_; 
wire _abc_41356_new_n2842_; 
wire _abc_41356_new_n2843_; 
wire _abc_41356_new_n2844_; 
wire _abc_41356_new_n2845_; 
wire _abc_41356_new_n2847_; 
wire _abc_41356_new_n2848_; 
wire _abc_41356_new_n2849_; 
wire _abc_41356_new_n2850_; 
wire _abc_41356_new_n2851_; 
wire _abc_41356_new_n2852_; 
wire _abc_41356_new_n2853_; 
wire _abc_41356_new_n2854_; 
wire _abc_41356_new_n2855_; 
wire _abc_41356_new_n2856_; 
wire _abc_41356_new_n2857_; 
wire _abc_41356_new_n2858_; 
wire _abc_41356_new_n2859_; 
wire _abc_41356_new_n2860_; 
wire _abc_41356_new_n2861_; 
wire _abc_41356_new_n2862_; 
wire _abc_41356_new_n2863_; 
wire _abc_41356_new_n2864_; 
wire _abc_41356_new_n2865_; 
wire _abc_41356_new_n2866_; 
wire _abc_41356_new_n2867_; 
wire _abc_41356_new_n2868_; 
wire _abc_41356_new_n2869_; 
wire _abc_41356_new_n2870_; 
wire _abc_41356_new_n2871_; 
wire _abc_41356_new_n2872_; 
wire _abc_41356_new_n2874_; 
wire _abc_41356_new_n2875_; 
wire _abc_41356_new_n2876_; 
wire _abc_41356_new_n2877_; 
wire _abc_41356_new_n2878_; 
wire _abc_41356_new_n2879_; 
wire _abc_41356_new_n2880_; 
wire _abc_41356_new_n2881_; 
wire _abc_41356_new_n2882_; 
wire _abc_41356_new_n2883_; 
wire _abc_41356_new_n2884_; 
wire _abc_41356_new_n2885_; 
wire _abc_41356_new_n2886_; 
wire _abc_41356_new_n2887_; 
wire _abc_41356_new_n2888_; 
wire _abc_41356_new_n2889_; 
wire _abc_41356_new_n2890_; 
wire _abc_41356_new_n2891_; 
wire _abc_41356_new_n2892_; 
wire _abc_41356_new_n2893_; 
wire _abc_41356_new_n2895_; 
wire _abc_41356_new_n2896_; 
wire _abc_41356_new_n2897_; 
wire _abc_41356_new_n2898_; 
wire _abc_41356_new_n2899_; 
wire _abc_41356_new_n2900_; 
wire _abc_41356_new_n2901_; 
wire _abc_41356_new_n2902_; 
wire _abc_41356_new_n2903_; 
wire _abc_41356_new_n2904_; 
wire _abc_41356_new_n2905_; 
wire _abc_41356_new_n2906_; 
wire _abc_41356_new_n2907_; 
wire _abc_41356_new_n2909_; 
wire _abc_41356_new_n2910_; 
wire _abc_41356_new_n2911_; 
wire _abc_41356_new_n2912_; 
wire _abc_41356_new_n2913_; 
wire _abc_41356_new_n2914_; 
wire _abc_41356_new_n2915_; 
wire _abc_41356_new_n2916_; 
wire _abc_41356_new_n2917_; 
wire _abc_41356_new_n2919_; 
wire _abc_41356_new_n2920_; 
wire _abc_41356_new_n2921_; 
wire _abc_41356_new_n2922_; 
wire _abc_41356_new_n2924_; 
wire _abc_41356_new_n2925_; 
wire _abc_41356_new_n2926_; 
wire _abc_41356_new_n2927_; 
wire _abc_41356_new_n2928_; 
wire _abc_41356_new_n2929_; 
wire _abc_41356_new_n2930_; 
wire _abc_41356_new_n2931_; 
wire _abc_41356_new_n2932_; 
wire _abc_41356_new_n2933_; 
wire _abc_41356_new_n2934_; 
wire _abc_41356_new_n2935_; 
wire _abc_41356_new_n2936_; 
wire _abc_41356_new_n2937_; 
wire _abc_41356_new_n2938_; 
wire _abc_41356_new_n2939_; 
wire _abc_41356_new_n2940_; 
wire _abc_41356_new_n2941_; 
wire _abc_41356_new_n2942_; 
wire _abc_41356_new_n2944_; 
wire _abc_41356_new_n2945_; 
wire _abc_41356_new_n2946_; 
wire _abc_41356_new_n2947_; 
wire _abc_41356_new_n2948_; 
wire _abc_41356_new_n2949_; 
wire _abc_41356_new_n2950_; 
wire _abc_41356_new_n2952_; 
wire _abc_41356_new_n2953_; 
wire _abc_41356_new_n2954_; 
wire _abc_41356_new_n2955_; 
wire _abc_41356_new_n2957_; 
wire _abc_41356_new_n2958_; 
wire _abc_41356_new_n2959_; 
wire _abc_41356_new_n2960_; 
wire _abc_41356_new_n2961_; 
wire _abc_41356_new_n2962_; 
wire _abc_41356_new_n2963_; 
wire _abc_41356_new_n2965_; 
wire _abc_41356_new_n2966_; 
wire _abc_41356_new_n2967_; 
wire _abc_41356_new_n2968_; 
wire _abc_41356_new_n2970_; 
wire _abc_41356_new_n2971_; 
wire _abc_41356_new_n2972_; 
wire _abc_41356_new_n2973_; 
wire _abc_41356_new_n2975_; 
wire _abc_41356_new_n2976_; 
wire _abc_41356_new_n2977_; 
wire _abc_41356_new_n2978_; 
wire _abc_41356_new_n2979_; 
wire _abc_41356_new_n2980_; 
wire _abc_41356_new_n2981_; 
wire _abc_41356_new_n2983_; 
wire _abc_41356_new_n2984_; 
wire _abc_41356_new_n2985_; 
wire _abc_41356_new_n2986_; 
wire _abc_41356_new_n2988_; 
wire _abc_41356_new_n2989_; 
wire _abc_41356_new_n2990_; 
wire _abc_41356_new_n2991_; 
wire _abc_41356_new_n2992_; 
wire _abc_41356_new_n2993_; 
wire _abc_41356_new_n2994_; 
wire _abc_41356_new_n2995_; 
wire _abc_41356_new_n2996_; 
wire _abc_41356_new_n2997_; 
wire _abc_41356_new_n2998_; 
wire _abc_41356_new_n2999_; 
wire _abc_41356_new_n3000_; 
wire _abc_41356_new_n3001_; 
wire _abc_41356_new_n3002_; 
wire _abc_41356_new_n3003_; 
wire _abc_41356_new_n3004_; 
wire _abc_41356_new_n3005_; 
wire _abc_41356_new_n3006_; 
wire _abc_41356_new_n3007_; 
wire _abc_41356_new_n3008_; 
wire _abc_41356_new_n3009_; 
wire _abc_41356_new_n3010_; 
wire _abc_41356_new_n3011_; 
wire _abc_41356_new_n3012_; 
wire _abc_41356_new_n3013_; 
wire _abc_41356_new_n3014_; 
wire _abc_41356_new_n3015_; 
wire _abc_41356_new_n3016_; 
wire _abc_41356_new_n3017_; 
wire _abc_41356_new_n3018_; 
wire _abc_41356_new_n3019_; 
wire _abc_41356_new_n3020_; 
wire _abc_41356_new_n3021_; 
wire _abc_41356_new_n3022_; 
wire _abc_41356_new_n3023_; 
wire _abc_41356_new_n3025_; 
wire _abc_41356_new_n3026_; 
wire _abc_41356_new_n3027_; 
wire _abc_41356_new_n3028_; 
wire _abc_41356_new_n3029_; 
wire _abc_41356_new_n3030_; 
wire _abc_41356_new_n3031_; 
wire _abc_41356_new_n3032_; 
wire _abc_41356_new_n3033_; 
wire _abc_41356_new_n3034_; 
wire _abc_41356_new_n3035_; 
wire _abc_41356_new_n3036_; 
wire _abc_41356_new_n3037_; 
wire _abc_41356_new_n3038_; 
wire _abc_41356_new_n3039_; 
wire _abc_41356_new_n3040_; 
wire _abc_41356_new_n3041_; 
wire _abc_41356_new_n3042_; 
wire _abc_41356_new_n3043_; 
wire _abc_41356_new_n3044_; 
wire _abc_41356_new_n3045_; 
wire _abc_41356_new_n3046_; 
wire _abc_41356_new_n3047_; 
wire _abc_41356_new_n3048_; 
wire _abc_41356_new_n3050_; 
wire _abc_41356_new_n3051_; 
wire _abc_41356_new_n3052_; 
wire _abc_41356_new_n3053_; 
wire _abc_41356_new_n3054_; 
wire _abc_41356_new_n3055_; 
wire _abc_41356_new_n3056_; 
wire _abc_41356_new_n3057_; 
wire _abc_41356_new_n3058_; 
wire _abc_41356_new_n3059_; 
wire _abc_41356_new_n3060_; 
wire _abc_41356_new_n3061_; 
wire _abc_41356_new_n3062_; 
wire _abc_41356_new_n3063_; 
wire _abc_41356_new_n3064_; 
wire _abc_41356_new_n3065_; 
wire _abc_41356_new_n3066_; 
wire _abc_41356_new_n3067_; 
wire _abc_41356_new_n3068_; 
wire _abc_41356_new_n3069_; 
wire _abc_41356_new_n3070_; 
wire _abc_41356_new_n3071_; 
wire _abc_41356_new_n3072_; 
wire _abc_41356_new_n3073_; 
wire _abc_41356_new_n3075_; 
wire _abc_41356_new_n3076_; 
wire _abc_41356_new_n3077_; 
wire _abc_41356_new_n3078_; 
wire _abc_41356_new_n3079_; 
wire _abc_41356_new_n3080_; 
wire _abc_41356_new_n3081_; 
wire _abc_41356_new_n3082_; 
wire _abc_41356_new_n3083_; 
wire _abc_41356_new_n3084_; 
wire _abc_41356_new_n3085_; 
wire _abc_41356_new_n3086_; 
wire _abc_41356_new_n3087_; 
wire _abc_41356_new_n3088_; 
wire _abc_41356_new_n3089_; 
wire _abc_41356_new_n3090_; 
wire _abc_41356_new_n3091_; 
wire _abc_41356_new_n3092_; 
wire _abc_41356_new_n3093_; 
wire _abc_41356_new_n3094_; 
wire _abc_41356_new_n3095_; 
wire _abc_41356_new_n3096_; 
wire _abc_41356_new_n3097_; 
wire _abc_41356_new_n3098_; 
wire _abc_41356_new_n3100_; 
wire _abc_41356_new_n3101_; 
wire _abc_41356_new_n3102_; 
wire _abc_41356_new_n3103_; 
wire _abc_41356_new_n3104_; 
wire _abc_41356_new_n3105_; 
wire _abc_41356_new_n3106_; 
wire _abc_41356_new_n3107_; 
wire _abc_41356_new_n3108_; 
wire _abc_41356_new_n3109_; 
wire _abc_41356_new_n3110_; 
wire _abc_41356_new_n3111_; 
wire _abc_41356_new_n3112_; 
wire _abc_41356_new_n3113_; 
wire _abc_41356_new_n3114_; 
wire _abc_41356_new_n3115_; 
wire _abc_41356_new_n3116_; 
wire _abc_41356_new_n3117_; 
wire _abc_41356_new_n3118_; 
wire _abc_41356_new_n3119_; 
wire _abc_41356_new_n3120_; 
wire _abc_41356_new_n3121_; 
wire _abc_41356_new_n3122_; 
wire _abc_41356_new_n3123_; 
wire _abc_41356_new_n3125_; 
wire _abc_41356_new_n3126_; 
wire _abc_41356_new_n3127_; 
wire _abc_41356_new_n3128_; 
wire _abc_41356_new_n3129_; 
wire _abc_41356_new_n3130_; 
wire _abc_41356_new_n3131_; 
wire _abc_41356_new_n3132_; 
wire _abc_41356_new_n3133_; 
wire _abc_41356_new_n3134_; 
wire _abc_41356_new_n3135_; 
wire _abc_41356_new_n3136_; 
wire _abc_41356_new_n3137_; 
wire _abc_41356_new_n3138_; 
wire _abc_41356_new_n3139_; 
wire _abc_41356_new_n3140_; 
wire _abc_41356_new_n3141_; 
wire _abc_41356_new_n3142_; 
wire _abc_41356_new_n3143_; 
wire _abc_41356_new_n3144_; 
wire _abc_41356_new_n3145_; 
wire _abc_41356_new_n3146_; 
wire _abc_41356_new_n3147_; 
wire _abc_41356_new_n3148_; 
wire _abc_41356_new_n3150_; 
wire _abc_41356_new_n3151_; 
wire _abc_41356_new_n3152_; 
wire _abc_41356_new_n3153_; 
wire _abc_41356_new_n3154_; 
wire _abc_41356_new_n3155_; 
wire _abc_41356_new_n3156_; 
wire _abc_41356_new_n3157_; 
wire _abc_41356_new_n3158_; 
wire _abc_41356_new_n3159_; 
wire _abc_41356_new_n3160_; 
wire _abc_41356_new_n3161_; 
wire _abc_41356_new_n3162_; 
wire _abc_41356_new_n3163_; 
wire _abc_41356_new_n3164_; 
wire _abc_41356_new_n3165_; 
wire _abc_41356_new_n3166_; 
wire _abc_41356_new_n3167_; 
wire _abc_41356_new_n3168_; 
wire _abc_41356_new_n3169_; 
wire _abc_41356_new_n3170_; 
wire _abc_41356_new_n3171_; 
wire _abc_41356_new_n3172_; 
wire _abc_41356_new_n3173_; 
wire _abc_41356_new_n3175_; 
wire _abc_41356_new_n3176_; 
wire _abc_41356_new_n3177_; 
wire _abc_41356_new_n3178_; 
wire _abc_41356_new_n3179_; 
wire _abc_41356_new_n3180_; 
wire _abc_41356_new_n3181_; 
wire _abc_41356_new_n3182_; 
wire _abc_41356_new_n3183_; 
wire _abc_41356_new_n3184_; 
wire _abc_41356_new_n3185_; 
wire _abc_41356_new_n3186_; 
wire _abc_41356_new_n3187_; 
wire _abc_41356_new_n3188_; 
wire _abc_41356_new_n3189_; 
wire _abc_41356_new_n3190_; 
wire _abc_41356_new_n3191_; 
wire _abc_41356_new_n3192_; 
wire _abc_41356_new_n3193_; 
wire _abc_41356_new_n3194_; 
wire _abc_41356_new_n3195_; 
wire _abc_41356_new_n3196_; 
wire _abc_41356_new_n3197_; 
wire _abc_41356_new_n3198_; 
wire _abc_41356_new_n3200_; 
wire _abc_41356_new_n3201_; 
wire _abc_41356_new_n3202_; 
wire _abc_41356_new_n3203_; 
wire _abc_41356_new_n3204_; 
wire _abc_41356_new_n3205_; 
wire _abc_41356_new_n3206_; 
wire _abc_41356_new_n3207_; 
wire _abc_41356_new_n3209_; 
wire _abc_41356_new_n3210_; 
wire _abc_41356_new_n3211_; 
wire _abc_41356_new_n3212_; 
wire _abc_41356_new_n3213_; 
wire _abc_41356_new_n3214_; 
wire _abc_41356_new_n3215_; 
wire _abc_41356_new_n3216_; 
wire _abc_41356_new_n3217_; 
wire _abc_41356_new_n3218_; 
wire _abc_41356_new_n3219_; 
wire _abc_41356_new_n3220_; 
wire _abc_41356_new_n3221_; 
wire _abc_41356_new_n3222_; 
wire _abc_41356_new_n3223_; 
wire _abc_41356_new_n3224_; 
wire _abc_41356_new_n3226_; 
wire _abc_41356_new_n3227_; 
wire _abc_41356_new_n3228_; 
wire _abc_41356_new_n3229_; 
wire _abc_41356_new_n3230_; 
wire _abc_41356_new_n3231_; 
wire _abc_41356_new_n3232_; 
wire _abc_41356_new_n3233_; 
wire _abc_41356_new_n3235_; 
wire _abc_41356_new_n3236_; 
wire _abc_41356_new_n3237_; 
wire _abc_41356_new_n3238_; 
wire _abc_41356_new_n3239_; 
wire _abc_41356_new_n3240_; 
wire _abc_41356_new_n3241_; 
wire _abc_41356_new_n3242_; 
wire _abc_41356_new_n3243_; 
wire _abc_41356_new_n3244_; 
wire _abc_41356_new_n3245_; 
wire _abc_41356_new_n3246_; 
wire _abc_41356_new_n3248_; 
wire _abc_41356_new_n3249_; 
wire _abc_41356_new_n3250_; 
wire _abc_41356_new_n3251_; 
wire _abc_41356_new_n3252_; 
wire _abc_41356_new_n3253_; 
wire _abc_41356_new_n3254_; 
wire _abc_41356_new_n3255_; 
wire _abc_41356_new_n3256_; 
wire _abc_41356_new_n3257_; 
wire _abc_41356_new_n3258_; 
wire _abc_41356_new_n3259_; 
wire _abc_41356_new_n3260_; 
wire _abc_41356_new_n3261_; 
wire _abc_41356_new_n3262_; 
wire _abc_41356_new_n3263_; 
wire _abc_41356_new_n3265_; 
wire _abc_41356_new_n3266_; 
wire _abc_41356_new_n3267_; 
wire _abc_41356_new_n3268_; 
wire _abc_41356_new_n3269_; 
wire _abc_41356_new_n3270_; 
wire _abc_41356_new_n3271_; 
wire _abc_41356_new_n3272_; 
wire _abc_41356_new_n3273_; 
wire _abc_41356_new_n3274_; 
wire _abc_41356_new_n3275_; 
wire _abc_41356_new_n3276_; 
wire _abc_41356_new_n3277_; 
wire _abc_41356_new_n3278_; 
wire _abc_41356_new_n3279_; 
wire _abc_41356_new_n3280_; 
wire _abc_41356_new_n3281_; 
wire _abc_41356_new_n3282_; 
wire _abc_41356_new_n3283_; 
wire _abc_41356_new_n3284_; 
wire _abc_41356_new_n3285_; 
wire _abc_41356_new_n3286_; 
wire _abc_41356_new_n3287_; 
wire _abc_41356_new_n3288_; 
wire _abc_41356_new_n3289_; 
wire _abc_41356_new_n3290_; 
wire _abc_41356_new_n3291_; 
wire _abc_41356_new_n3292_; 
wire _abc_41356_new_n3293_; 
wire _abc_41356_new_n3294_; 
wire _abc_41356_new_n3295_; 
wire _abc_41356_new_n3296_; 
wire _abc_41356_new_n3297_; 
wire _abc_41356_new_n3298_; 
wire _abc_41356_new_n3299_; 
wire _abc_41356_new_n3300_; 
wire _abc_41356_new_n3301_; 
wire _abc_41356_new_n3302_; 
wire _abc_41356_new_n3303_; 
wire _abc_41356_new_n3304_; 
wire _abc_41356_new_n3305_; 
wire _abc_41356_new_n3306_; 
wire _abc_41356_new_n3307_; 
wire _abc_41356_new_n3308_; 
wire _abc_41356_new_n3309_; 
wire _abc_41356_new_n3310_; 
wire _abc_41356_new_n3311_; 
wire _abc_41356_new_n3312_; 
wire _abc_41356_new_n3313_; 
wire _abc_41356_new_n3314_; 
wire _abc_41356_new_n3315_; 
wire _abc_41356_new_n3317_; 
wire _abc_41356_new_n3318_; 
wire _abc_41356_new_n3319_; 
wire _abc_41356_new_n3320_; 
wire _abc_41356_new_n3321_; 
wire _abc_41356_new_n3322_; 
wire _abc_41356_new_n3324_; 
wire _abc_41356_new_n3325_; 
wire _abc_41356_new_n3327_; 
wire _abc_41356_new_n3328_; 
wire _abc_41356_new_n3330_; 
wire _abc_41356_new_n3331_; 
wire _abc_41356_new_n3333_; 
wire _abc_41356_new_n3334_; 
wire _abc_41356_new_n3336_; 
wire _abc_41356_new_n3337_; 
wire _abc_41356_new_n3339_; 
wire _abc_41356_new_n3340_; 
wire _abc_41356_new_n3342_; 
wire _abc_41356_new_n3343_; 
wire _abc_41356_new_n3345_; 
wire _abc_41356_new_n3346_; 
wire _abc_41356_new_n3347_; 
wire _abc_41356_new_n3348_; 
wire _abc_41356_new_n3349_; 
wire _abc_41356_new_n3350_; 
wire _abc_41356_new_n3351_; 
wire _abc_41356_new_n3353_; 
wire _abc_41356_new_n3354_; 
wire _abc_41356_new_n3355_; 
wire _abc_41356_new_n3356_; 
wire _abc_41356_new_n3357_; 
wire _abc_41356_new_n3358_; 
wire _abc_41356_new_n3359_; 
wire _abc_41356_new_n3360_; 
wire _abc_41356_new_n3361_; 
wire _abc_41356_new_n3362_; 
wire _abc_41356_new_n3363_; 
wire _abc_41356_new_n3364_; 
wire _abc_41356_new_n3365_; 
wire _abc_41356_new_n3366_; 
wire _abc_41356_new_n3367_; 
wire _abc_41356_new_n3368_; 
wire _abc_41356_new_n3369_; 
wire _abc_41356_new_n3370_; 
wire _abc_41356_new_n3371_; 
wire _abc_41356_new_n3372_; 
wire _abc_41356_new_n3373_; 
wire _abc_41356_new_n3374_; 
wire _abc_41356_new_n3375_; 
wire _abc_41356_new_n3376_; 
wire _abc_41356_new_n3377_; 
wire _abc_41356_new_n3378_; 
wire _abc_41356_new_n3379_; 
wire _abc_41356_new_n3380_; 
wire _abc_41356_new_n3381_; 
wire _abc_41356_new_n3382_; 
wire _abc_41356_new_n3383_; 
wire _abc_41356_new_n3384_; 
wire _abc_41356_new_n3385_; 
wire _abc_41356_new_n3386_; 
wire _abc_41356_new_n3387_; 
wire _abc_41356_new_n3388_; 
wire _abc_41356_new_n3389_; 
wire _abc_41356_new_n3390_; 
wire _abc_41356_new_n3391_; 
wire _abc_41356_new_n3392_; 
wire _abc_41356_new_n3393_; 
wire _abc_41356_new_n3394_; 
wire _abc_41356_new_n3395_; 
wire _abc_41356_new_n3396_; 
wire _abc_41356_new_n3397_; 
wire _abc_41356_new_n3398_; 
wire _abc_41356_new_n3399_; 
wire _abc_41356_new_n3400_; 
wire _abc_41356_new_n3401_; 
wire _abc_41356_new_n3402_; 
wire _abc_41356_new_n3403_; 
wire _abc_41356_new_n3404_; 
wire _abc_41356_new_n3405_; 
wire _abc_41356_new_n3406_; 
wire _abc_41356_new_n3407_; 
wire _abc_41356_new_n3408_; 
wire _abc_41356_new_n3409_; 
wire _abc_41356_new_n3410_; 
wire _abc_41356_new_n3411_; 
wire _abc_41356_new_n3412_; 
wire _abc_41356_new_n3413_; 
wire _abc_41356_new_n3414_; 
wire _abc_41356_new_n3415_; 
wire _abc_41356_new_n3416_; 
wire _abc_41356_new_n3417_; 
wire _abc_41356_new_n3418_; 
wire _abc_41356_new_n3419_; 
wire _abc_41356_new_n3420_; 
wire _abc_41356_new_n3421_; 
wire _abc_41356_new_n3422_; 
wire _abc_41356_new_n3423_; 
wire _abc_41356_new_n3424_; 
wire _abc_41356_new_n3425_; 
wire _abc_41356_new_n3426_; 
wire _abc_41356_new_n3427_; 
wire _abc_41356_new_n3428_; 
wire _abc_41356_new_n3429_; 
wire _abc_41356_new_n3430_; 
wire _abc_41356_new_n3431_; 
wire _abc_41356_new_n3432_; 
wire _abc_41356_new_n3433_; 
wire _abc_41356_new_n3434_; 
wire _abc_41356_new_n3435_; 
wire _abc_41356_new_n3436_; 
wire _abc_41356_new_n3437_; 
wire _abc_41356_new_n3438_; 
wire _abc_41356_new_n3439_; 
wire _abc_41356_new_n3440_; 
wire _abc_41356_new_n3441_; 
wire _abc_41356_new_n3442_; 
wire _abc_41356_new_n3443_; 
wire _abc_41356_new_n3444_; 
wire _abc_41356_new_n3445_; 
wire _abc_41356_new_n3446_; 
wire _abc_41356_new_n3447_; 
wire _abc_41356_new_n3448_; 
wire _abc_41356_new_n3449_; 
wire _abc_41356_new_n3450_; 
wire _abc_41356_new_n3451_; 
wire _abc_41356_new_n3452_; 
wire _abc_41356_new_n3453_; 
wire _abc_41356_new_n3454_; 
wire _abc_41356_new_n3455_; 
wire _abc_41356_new_n3456_; 
wire _abc_41356_new_n3458_; 
wire _abc_41356_new_n3459_; 
wire _abc_41356_new_n3460_; 
wire _abc_41356_new_n3461_; 
wire _abc_41356_new_n3462_; 
wire _abc_41356_new_n3463_; 
wire _abc_41356_new_n3464_; 
wire _abc_41356_new_n3465_; 
wire _abc_41356_new_n3466_; 
wire _abc_41356_new_n3467_; 
wire _abc_41356_new_n3468_; 
wire _abc_41356_new_n3469_; 
wire _abc_41356_new_n3470_; 
wire _abc_41356_new_n3471_; 
wire _abc_41356_new_n3472_; 
wire _abc_41356_new_n3473_; 
wire _abc_41356_new_n3474_; 
wire _abc_41356_new_n3475_; 
wire _abc_41356_new_n3476_; 
wire _abc_41356_new_n3477_; 
wire _abc_41356_new_n3478_; 
wire _abc_41356_new_n3479_; 
wire _abc_41356_new_n3480_; 
wire _abc_41356_new_n3481_; 
wire _abc_41356_new_n3482_; 
wire _abc_41356_new_n3483_; 
wire _abc_41356_new_n3484_; 
wire _abc_41356_new_n3485_; 
wire _abc_41356_new_n3486_; 
wire _abc_41356_new_n3487_; 
wire _abc_41356_new_n3488_; 
wire _abc_41356_new_n3489_; 
wire _abc_41356_new_n3490_; 
wire _abc_41356_new_n3491_; 
wire _abc_41356_new_n3492_; 
wire _abc_41356_new_n3494_; 
wire _abc_41356_new_n3495_; 
wire _abc_41356_new_n3496_; 
wire _abc_41356_new_n3497_; 
wire _abc_41356_new_n3498_; 
wire _abc_41356_new_n3499_; 
wire _abc_41356_new_n3500_; 
wire _abc_41356_new_n3501_; 
wire _abc_41356_new_n3502_; 
wire _abc_41356_new_n3503_; 
wire _abc_41356_new_n3504_; 
wire _abc_41356_new_n3505_; 
wire _abc_41356_new_n3506_; 
wire _abc_41356_new_n3507_; 
wire _abc_41356_new_n3508_; 
wire _abc_41356_new_n3509_; 
wire _abc_41356_new_n3510_; 
wire _abc_41356_new_n3511_; 
wire _abc_41356_new_n3512_; 
wire _abc_41356_new_n3513_; 
wire _abc_41356_new_n3514_; 
wire _abc_41356_new_n3515_; 
wire _abc_41356_new_n3516_; 
wire _abc_41356_new_n3517_; 
wire _abc_41356_new_n3518_; 
wire _abc_41356_new_n3519_; 
wire _abc_41356_new_n3520_; 
wire _abc_41356_new_n3521_; 
wire _abc_41356_new_n3522_; 
wire _abc_41356_new_n3523_; 
wire _abc_41356_new_n3524_; 
wire _abc_41356_new_n3525_; 
wire _abc_41356_new_n3526_; 
wire _abc_41356_new_n3527_; 
wire _abc_41356_new_n3528_; 
wire _abc_41356_new_n3529_; 
wire _abc_41356_new_n3531_; 
wire _abc_41356_new_n3532_; 
wire _abc_41356_new_n3533_; 
wire _abc_41356_new_n3534_; 
wire _abc_41356_new_n3535_; 
wire _abc_41356_new_n3536_; 
wire _abc_41356_new_n3537_; 
wire _abc_41356_new_n3538_; 
wire _abc_41356_new_n3539_; 
wire _abc_41356_new_n3540_; 
wire _abc_41356_new_n3541_; 
wire _abc_41356_new_n3542_; 
wire _abc_41356_new_n3543_; 
wire _abc_41356_new_n3544_; 
wire _abc_41356_new_n3545_; 
wire _abc_41356_new_n3546_; 
wire _abc_41356_new_n3547_; 
wire _abc_41356_new_n3548_; 
wire _abc_41356_new_n3549_; 
wire _abc_41356_new_n3550_; 
wire _abc_41356_new_n3551_; 
wire _abc_41356_new_n3552_; 
wire _abc_41356_new_n3553_; 
wire _abc_41356_new_n3554_; 
wire _abc_41356_new_n3555_; 
wire _abc_41356_new_n3556_; 
wire _abc_41356_new_n3557_; 
wire _abc_41356_new_n3558_; 
wire _abc_41356_new_n3559_; 
wire _abc_41356_new_n3560_; 
wire _abc_41356_new_n3561_; 
wire _abc_41356_new_n3562_; 
wire _abc_41356_new_n3563_; 
wire _abc_41356_new_n3565_; 
wire _abc_41356_new_n3566_; 
wire _abc_41356_new_n3567_; 
wire _abc_41356_new_n3568_; 
wire _abc_41356_new_n3569_; 
wire _abc_41356_new_n3570_; 
wire _abc_41356_new_n3571_; 
wire _abc_41356_new_n3572_; 
wire _abc_41356_new_n3573_; 
wire _abc_41356_new_n3574_; 
wire _abc_41356_new_n3575_; 
wire _abc_41356_new_n3576_; 
wire _abc_41356_new_n3577_; 
wire _abc_41356_new_n3578_; 
wire _abc_41356_new_n3579_; 
wire _abc_41356_new_n3580_; 
wire _abc_41356_new_n3581_; 
wire _abc_41356_new_n3582_; 
wire _abc_41356_new_n3583_; 
wire _abc_41356_new_n3584_; 
wire _abc_41356_new_n3585_; 
wire _abc_41356_new_n3586_; 
wire _abc_41356_new_n3587_; 
wire _abc_41356_new_n3588_; 
wire _abc_41356_new_n3589_; 
wire _abc_41356_new_n3590_; 
wire _abc_41356_new_n3591_; 
wire _abc_41356_new_n3593_; 
wire _abc_41356_new_n3594_; 
wire _abc_41356_new_n3595_; 
wire _abc_41356_new_n3596_; 
wire _abc_41356_new_n3597_; 
wire _abc_41356_new_n3598_; 
wire _abc_41356_new_n3599_; 
wire _abc_41356_new_n3600_; 
wire _abc_41356_new_n3601_; 
wire _abc_41356_new_n3602_; 
wire _abc_41356_new_n3603_; 
wire _abc_41356_new_n3604_; 
wire _abc_41356_new_n3605_; 
wire _abc_41356_new_n3606_; 
wire _abc_41356_new_n3607_; 
wire _abc_41356_new_n3608_; 
wire _abc_41356_new_n3609_; 
wire _abc_41356_new_n3610_; 
wire _abc_41356_new_n3611_; 
wire _abc_41356_new_n3612_; 
wire _abc_41356_new_n3613_; 
wire _abc_41356_new_n3615_; 
wire _abc_41356_new_n3616_; 
wire _abc_41356_new_n3617_; 
wire _abc_41356_new_n3618_; 
wire _abc_41356_new_n3620_; 
wire _abc_41356_new_n3621_; 
wire _abc_41356_new_n3623_; 
wire _abc_41356_new_n3624_; 
wire _abc_41356_new_n3625_; 
wire _abc_41356_new_n3626_; 
wire _abc_41356_new_n3628_; 
wire _abc_41356_new_n3629_; 
wire _abc_41356_new_n3630_; 
wire _abc_41356_new_n3631_; 
wire _abc_41356_new_n3633_; 
wire _abc_41356_new_n3634_; 
wire _abc_41356_new_n3635_; 
wire _abc_41356_new_n3637_; 
wire _abc_41356_new_n3638_; 
wire _abc_41356_new_n3639_; 
wire _abc_41356_new_n3641_; 
wire _abc_41356_new_n3642_; 
wire _abc_41356_new_n3643_; 
wire _abc_41356_new_n3644_; 
wire _abc_41356_new_n3646_; 
wire _abc_41356_new_n3647_; 
wire _abc_41356_new_n3648_; 
wire _abc_41356_new_n3650_; 
wire _abc_41356_new_n3651_; 
wire _abc_41356_new_n3652_; 
wire _abc_41356_new_n3654_; 
wire _abc_41356_new_n3655_; 
wire _abc_41356_new_n3656_; 
wire _abc_41356_new_n3658_; 
wire _abc_41356_new_n3659_; 
wire _abc_41356_new_n3660_; 
wire _abc_41356_new_n3661_; 
wire _abc_41356_new_n3663_; 
wire _abc_41356_new_n3664_; 
wire _abc_41356_new_n3665_; 
wire _abc_41356_new_n3666_; 
wire _abc_41356_new_n3668_; 
wire _abc_41356_new_n3669_; 
wire _abc_41356_new_n3670_; 
wire _abc_41356_new_n3671_; 
wire _abc_41356_new_n3673_; 
wire _abc_41356_new_n3674_; 
wire _abc_41356_new_n3675_; 
wire _abc_41356_new_n3676_; 
wire _abc_41356_new_n3678_; 
wire _abc_41356_new_n3679_; 
wire _abc_41356_new_n3680_; 
wire _abc_41356_new_n3681_; 
wire _abc_41356_new_n3683_; 
wire _abc_41356_new_n3684_; 
wire _abc_41356_new_n3685_; 
wire _abc_41356_new_n3686_; 
wire _abc_41356_new_n3688_; 
wire _abc_41356_new_n3689_; 
wire _abc_41356_new_n3690_; 
wire _abc_41356_new_n3691_; 
wire _abc_41356_new_n3693_; 
wire _abc_41356_new_n3694_; 
wire _abc_41356_new_n3695_; 
wire _abc_41356_new_n3696_; 
wire _abc_41356_new_n3698_; 
wire _abc_41356_new_n3699_; 
wire _abc_41356_new_n3700_; 
wire _abc_41356_new_n3701_; 
wire _abc_41356_new_n3702_; 
wire _abc_41356_new_n3703_; 
wire _abc_41356_new_n3704_; 
wire _abc_41356_new_n3705_; 
wire _abc_41356_new_n3706_; 
wire _abc_41356_new_n3707_; 
wire _abc_41356_new_n3708_; 
wire _abc_41356_new_n3709_; 
wire _abc_41356_new_n3710_; 
wire _abc_41356_new_n3711_; 
wire _abc_41356_new_n3712_; 
wire _abc_41356_new_n3713_; 
wire _abc_41356_new_n3714_; 
wire _abc_41356_new_n3715_; 
wire _abc_41356_new_n3716_; 
wire _abc_41356_new_n3717_; 
wire _abc_41356_new_n3718_; 
wire _abc_41356_new_n3719_; 
wire _abc_41356_new_n3720_; 
wire _abc_41356_new_n3721_; 
wire _abc_41356_new_n3722_; 
wire _abc_41356_new_n3723_; 
wire _abc_41356_new_n3724_; 
wire _abc_41356_new_n3725_; 
wire _abc_41356_new_n3726_; 
wire _abc_41356_new_n3727_; 
wire _abc_41356_new_n3728_; 
wire _abc_41356_new_n3729_; 
wire _abc_41356_new_n3730_; 
wire _abc_41356_new_n3731_; 
wire _abc_41356_new_n3732_; 
wire _abc_41356_new_n3733_; 
wire _abc_41356_new_n3734_; 
wire _abc_41356_new_n3735_; 
wire _abc_41356_new_n3736_; 
wire _abc_41356_new_n3737_; 
wire _abc_41356_new_n3738_; 
wire _abc_41356_new_n3739_; 
wire _abc_41356_new_n3740_; 
wire _abc_41356_new_n3741_; 
wire _abc_41356_new_n3742_; 
wire _abc_41356_new_n3743_; 
wire _abc_41356_new_n3744_; 
wire _abc_41356_new_n3745_; 
wire _abc_41356_new_n3746_; 
wire _abc_41356_new_n3747_; 
wire _abc_41356_new_n3748_; 
wire _abc_41356_new_n3749_; 
wire _abc_41356_new_n3750_; 
wire _abc_41356_new_n3751_; 
wire _abc_41356_new_n3752_; 
wire _abc_41356_new_n3753_; 
wire _abc_41356_new_n3755_; 
wire _abc_41356_new_n3756_; 
wire _abc_41356_new_n3757_; 
wire _abc_41356_new_n3758_; 
wire _abc_41356_new_n3759_; 
wire _abc_41356_new_n3760_; 
wire _abc_41356_new_n3761_; 
wire _abc_41356_new_n3762_; 
wire _abc_41356_new_n3763_; 
wire _abc_41356_new_n3764_; 
wire _abc_41356_new_n3765_; 
wire _abc_41356_new_n3766_; 
wire _abc_41356_new_n3767_; 
wire _abc_41356_new_n3768_; 
wire _abc_41356_new_n3769_; 
wire _abc_41356_new_n3770_; 
wire _abc_41356_new_n3771_; 
wire _abc_41356_new_n3772_; 
wire _abc_41356_new_n3773_; 
wire _abc_41356_new_n3774_; 
wire _abc_41356_new_n3775_; 
wire _abc_41356_new_n3776_; 
wire _abc_41356_new_n3777_; 
wire _abc_41356_new_n3778_; 
wire _abc_41356_new_n3779_; 
wire _abc_41356_new_n3780_; 
wire _abc_41356_new_n3781_; 
wire _abc_41356_new_n3782_; 
wire _abc_41356_new_n3783_; 
wire _abc_41356_new_n3784_; 
wire _abc_41356_new_n3785_; 
wire _abc_41356_new_n3786_; 
wire _abc_41356_new_n3787_; 
wire _abc_41356_new_n3788_; 
wire _abc_41356_new_n3789_; 
wire _abc_41356_new_n3790_; 
wire _abc_41356_new_n3791_; 
wire _abc_41356_new_n3792_; 
wire _abc_41356_new_n3793_; 
wire _abc_41356_new_n3794_; 
wire _abc_41356_new_n3795_; 
wire _abc_41356_new_n3796_; 
wire _abc_41356_new_n3797_; 
wire _abc_41356_new_n3798_; 
wire _abc_41356_new_n3799_; 
wire _abc_41356_new_n3800_; 
wire _abc_41356_new_n3801_; 
wire _abc_41356_new_n3802_; 
wire _abc_41356_new_n3803_; 
wire _abc_41356_new_n3804_; 
wire _abc_41356_new_n3805_; 
wire _abc_41356_new_n3806_; 
wire _abc_41356_new_n3808_; 
wire _abc_41356_new_n3809_; 
wire _abc_41356_new_n3810_; 
wire _abc_41356_new_n3811_; 
wire _abc_41356_new_n3812_; 
wire _abc_41356_new_n3813_; 
wire _abc_41356_new_n3814_; 
wire _abc_41356_new_n3815_; 
wire _abc_41356_new_n3816_; 
wire _abc_41356_new_n3817_; 
wire _abc_41356_new_n3818_; 
wire _abc_41356_new_n3819_; 
wire _abc_41356_new_n3820_; 
wire _abc_41356_new_n3821_; 
wire _abc_41356_new_n3822_; 
wire _abc_41356_new_n3823_; 
wire _abc_41356_new_n3824_; 
wire _abc_41356_new_n3825_; 
wire _abc_41356_new_n3826_; 
wire _abc_41356_new_n3827_; 
wire _abc_41356_new_n3828_; 
wire _abc_41356_new_n3829_; 
wire _abc_41356_new_n3830_; 
wire _abc_41356_new_n3831_; 
wire _abc_41356_new_n3832_; 
wire _abc_41356_new_n3833_; 
wire _abc_41356_new_n3834_; 
wire _abc_41356_new_n3835_; 
wire _abc_41356_new_n3836_; 
wire _abc_41356_new_n3837_; 
wire _abc_41356_new_n3838_; 
wire _abc_41356_new_n3839_; 
wire _abc_41356_new_n3840_; 
wire _abc_41356_new_n3841_; 
wire _abc_41356_new_n3842_; 
wire _abc_41356_new_n3843_; 
wire _abc_41356_new_n3844_; 
wire _abc_41356_new_n3845_; 
wire _abc_41356_new_n3846_; 
wire _abc_41356_new_n3847_; 
wire _abc_41356_new_n3848_; 
wire _abc_41356_new_n3849_; 
wire _abc_41356_new_n3850_; 
wire _abc_41356_new_n3851_; 
wire _abc_41356_new_n3852_; 
wire _abc_41356_new_n3853_; 
wire _abc_41356_new_n3854_; 
wire _abc_41356_new_n3855_; 
wire _abc_41356_new_n3856_; 
wire _abc_41356_new_n3857_; 
wire _abc_41356_new_n3858_; 
wire _abc_41356_new_n3859_; 
wire _abc_41356_new_n3860_; 
wire _abc_41356_new_n3861_; 
wire _abc_41356_new_n3863_; 
wire _abc_41356_new_n3864_; 
wire _abc_41356_new_n3865_; 
wire _abc_41356_new_n3866_; 
wire _abc_41356_new_n3867_; 
wire _abc_41356_new_n3868_; 
wire _abc_41356_new_n3869_; 
wire _abc_41356_new_n3870_; 
wire _abc_41356_new_n3871_; 
wire _abc_41356_new_n3872_; 
wire _abc_41356_new_n3873_; 
wire _abc_41356_new_n3874_; 
wire _abc_41356_new_n3875_; 
wire _abc_41356_new_n3876_; 
wire _abc_41356_new_n3877_; 
wire _abc_41356_new_n3878_; 
wire _abc_41356_new_n3879_; 
wire _abc_41356_new_n3880_; 
wire _abc_41356_new_n3881_; 
wire _abc_41356_new_n3882_; 
wire _abc_41356_new_n3883_; 
wire _abc_41356_new_n3884_; 
wire _abc_41356_new_n3885_; 
wire _abc_41356_new_n3886_; 
wire _abc_41356_new_n3887_; 
wire _abc_41356_new_n3888_; 
wire _abc_41356_new_n3889_; 
wire _abc_41356_new_n3890_; 
wire _abc_41356_new_n3891_; 
wire _abc_41356_new_n3892_; 
wire _abc_41356_new_n3893_; 
wire _abc_41356_new_n3894_; 
wire _abc_41356_new_n3895_; 
wire _abc_41356_new_n3896_; 
wire _abc_41356_new_n3897_; 
wire _abc_41356_new_n3898_; 
wire _abc_41356_new_n3899_; 
wire _abc_41356_new_n3900_; 
wire _abc_41356_new_n3901_; 
wire _abc_41356_new_n3902_; 
wire _abc_41356_new_n3903_; 
wire _abc_41356_new_n3904_; 
wire _abc_41356_new_n3905_; 
wire _abc_41356_new_n3906_; 
wire _abc_41356_new_n3907_; 
wire _abc_41356_new_n3908_; 
wire _abc_41356_new_n3909_; 
wire _abc_41356_new_n3910_; 
wire _abc_41356_new_n3912_; 
wire _abc_41356_new_n3913_; 
wire _abc_41356_new_n3914_; 
wire _abc_41356_new_n3915_; 
wire _abc_41356_new_n3916_; 
wire _abc_41356_new_n3917_; 
wire _abc_41356_new_n3918_; 
wire _abc_41356_new_n3919_; 
wire _abc_41356_new_n3920_; 
wire _abc_41356_new_n3921_; 
wire _abc_41356_new_n3922_; 
wire _abc_41356_new_n3923_; 
wire _abc_41356_new_n3924_; 
wire _abc_41356_new_n3925_; 
wire _abc_41356_new_n3926_; 
wire _abc_41356_new_n3927_; 
wire _abc_41356_new_n3928_; 
wire _abc_41356_new_n3929_; 
wire _abc_41356_new_n3930_; 
wire _abc_41356_new_n3931_; 
wire _abc_41356_new_n3932_; 
wire _abc_41356_new_n3933_; 
wire _abc_41356_new_n3934_; 
wire _abc_41356_new_n3935_; 
wire _abc_41356_new_n3936_; 
wire _abc_41356_new_n3937_; 
wire _abc_41356_new_n3938_; 
wire _abc_41356_new_n3939_; 
wire _abc_41356_new_n3940_; 
wire _abc_41356_new_n3941_; 
wire _abc_41356_new_n3942_; 
wire _abc_41356_new_n3943_; 
wire _abc_41356_new_n3944_; 
wire _abc_41356_new_n3945_; 
wire _abc_41356_new_n3946_; 
wire _abc_41356_new_n3947_; 
wire _abc_41356_new_n3948_; 
wire _abc_41356_new_n3949_; 
wire _abc_41356_new_n3950_; 
wire _abc_41356_new_n3951_; 
wire _abc_41356_new_n3952_; 
wire _abc_41356_new_n3953_; 
wire _abc_41356_new_n3954_; 
wire _abc_41356_new_n3955_; 
wire _abc_41356_new_n3956_; 
wire _abc_41356_new_n3957_; 
wire _abc_41356_new_n3958_; 
wire _abc_41356_new_n3959_; 
wire _abc_41356_new_n3960_; 
wire _abc_41356_new_n3961_; 
wire _abc_41356_new_n3962_; 
wire _abc_41356_new_n3963_; 
wire _abc_41356_new_n3965_; 
wire _abc_41356_new_n3966_; 
wire _abc_41356_new_n3967_; 
wire _abc_41356_new_n3968_; 
wire _abc_41356_new_n3969_; 
wire _abc_41356_new_n3970_; 
wire _abc_41356_new_n3971_; 
wire _abc_41356_new_n3972_; 
wire _abc_41356_new_n3973_; 
wire _abc_41356_new_n3974_; 
wire _abc_41356_new_n3975_; 
wire _abc_41356_new_n3976_; 
wire _abc_41356_new_n3977_; 
wire _abc_41356_new_n3978_; 
wire _abc_41356_new_n3979_; 
wire _abc_41356_new_n3980_; 
wire _abc_41356_new_n3981_; 
wire _abc_41356_new_n3982_; 
wire _abc_41356_new_n3983_; 
wire _abc_41356_new_n3984_; 
wire _abc_41356_new_n3985_; 
wire _abc_41356_new_n3986_; 
wire _abc_41356_new_n3987_; 
wire _abc_41356_new_n3988_; 
wire _abc_41356_new_n3989_; 
wire _abc_41356_new_n3990_; 
wire _abc_41356_new_n3991_; 
wire _abc_41356_new_n3992_; 
wire _abc_41356_new_n3993_; 
wire _abc_41356_new_n3994_; 
wire _abc_41356_new_n3995_; 
wire _abc_41356_new_n3996_; 
wire _abc_41356_new_n3997_; 
wire _abc_41356_new_n3998_; 
wire _abc_41356_new_n3999_; 
wire _abc_41356_new_n4000_; 
wire _abc_41356_new_n4001_; 
wire _abc_41356_new_n4002_; 
wire _abc_41356_new_n4003_; 
wire _abc_41356_new_n4004_; 
wire _abc_41356_new_n4005_; 
wire _abc_41356_new_n4006_; 
wire _abc_41356_new_n4007_; 
wire _abc_41356_new_n4008_; 
wire _abc_41356_new_n4009_; 
wire _abc_41356_new_n4010_; 
wire _abc_41356_new_n4011_; 
wire _abc_41356_new_n4012_; 
wire _abc_41356_new_n4013_; 
wire _abc_41356_new_n4014_; 
wire _abc_41356_new_n4015_; 
wire _abc_41356_new_n4017_; 
wire _abc_41356_new_n4018_; 
wire _abc_41356_new_n4019_; 
wire _abc_41356_new_n4020_; 
wire _abc_41356_new_n4021_; 
wire _abc_41356_new_n4022_; 
wire _abc_41356_new_n4023_; 
wire _abc_41356_new_n4024_; 
wire _abc_41356_new_n4025_; 
wire _abc_41356_new_n4026_; 
wire _abc_41356_new_n4027_; 
wire _abc_41356_new_n4028_; 
wire _abc_41356_new_n4029_; 
wire _abc_41356_new_n4030_; 
wire _abc_41356_new_n4031_; 
wire _abc_41356_new_n4032_; 
wire _abc_41356_new_n4033_; 
wire _abc_41356_new_n4034_; 
wire _abc_41356_new_n4035_; 
wire _abc_41356_new_n4036_; 
wire _abc_41356_new_n4037_; 
wire _abc_41356_new_n4038_; 
wire _abc_41356_new_n4039_; 
wire _abc_41356_new_n4040_; 
wire _abc_41356_new_n4041_; 
wire _abc_41356_new_n4042_; 
wire _abc_41356_new_n4043_; 
wire _abc_41356_new_n4044_; 
wire _abc_41356_new_n4045_; 
wire _abc_41356_new_n4046_; 
wire _abc_41356_new_n4047_; 
wire _abc_41356_new_n4048_; 
wire _abc_41356_new_n4049_; 
wire _abc_41356_new_n4050_; 
wire _abc_41356_new_n4051_; 
wire _abc_41356_new_n4052_; 
wire _abc_41356_new_n4053_; 
wire _abc_41356_new_n4054_; 
wire _abc_41356_new_n4055_; 
wire _abc_41356_new_n4056_; 
wire _abc_41356_new_n4057_; 
wire _abc_41356_new_n4058_; 
wire _abc_41356_new_n4059_; 
wire _abc_41356_new_n4060_; 
wire _abc_41356_new_n4061_; 
wire _abc_41356_new_n4062_; 
wire _abc_41356_new_n4063_; 
wire _abc_41356_new_n4064_; 
wire _abc_41356_new_n4065_; 
wire _abc_41356_new_n4066_; 
wire _abc_41356_new_n4068_; 
wire _abc_41356_new_n4069_; 
wire _abc_41356_new_n4070_; 
wire _abc_41356_new_n4071_; 
wire _abc_41356_new_n4072_; 
wire _abc_41356_new_n4073_; 
wire _abc_41356_new_n4074_; 
wire _abc_41356_new_n4075_; 
wire _abc_41356_new_n4076_; 
wire _abc_41356_new_n4077_; 
wire _abc_41356_new_n4078_; 
wire _abc_41356_new_n4079_; 
wire _abc_41356_new_n4080_; 
wire _abc_41356_new_n4081_; 
wire _abc_41356_new_n4082_; 
wire _abc_41356_new_n4083_; 
wire _abc_41356_new_n4084_; 
wire _abc_41356_new_n4085_; 
wire _abc_41356_new_n4086_; 
wire _abc_41356_new_n4087_; 
wire _abc_41356_new_n4088_; 
wire _abc_41356_new_n4089_; 
wire _abc_41356_new_n4090_; 
wire _abc_41356_new_n4091_; 
wire _abc_41356_new_n4092_; 
wire _abc_41356_new_n4093_; 
wire _abc_41356_new_n4094_; 
wire _abc_41356_new_n4095_; 
wire _abc_41356_new_n4096_; 
wire _abc_41356_new_n4097_; 
wire _abc_41356_new_n4098_; 
wire _abc_41356_new_n4099_; 
wire _abc_41356_new_n4100_; 
wire _abc_41356_new_n4101_; 
wire _abc_41356_new_n4102_; 
wire _abc_41356_new_n4103_; 
wire _abc_41356_new_n4104_; 
wire _abc_41356_new_n4105_; 
wire _abc_41356_new_n4106_; 
wire _abc_41356_new_n4107_; 
wire _abc_41356_new_n4108_; 
wire _abc_41356_new_n4109_; 
wire _abc_41356_new_n4110_; 
wire _abc_41356_new_n4111_; 
wire _abc_41356_new_n4112_; 
wire _abc_41356_new_n4113_; 
wire _abc_41356_new_n4114_; 
wire _abc_41356_new_n4115_; 
wire _abc_41356_new_n4117_; 
wire _abc_41356_new_n4118_; 
wire _abc_41356_new_n4119_; 
wire _abc_41356_new_n4120_; 
wire _abc_41356_new_n4121_; 
wire _abc_41356_new_n4122_; 
wire _abc_41356_new_n4123_; 
wire _abc_41356_new_n4124_; 
wire _abc_41356_new_n4125_; 
wire _abc_41356_new_n4126_; 
wire _abc_41356_new_n4127_; 
wire _abc_41356_new_n4128_; 
wire _abc_41356_new_n4129_; 
wire _abc_41356_new_n4130_; 
wire _abc_41356_new_n4131_; 
wire _abc_41356_new_n4132_; 
wire _abc_41356_new_n4133_; 
wire _abc_41356_new_n4134_; 
wire _abc_41356_new_n4135_; 
wire _abc_41356_new_n4136_; 
wire _abc_41356_new_n4137_; 
wire _abc_41356_new_n4138_; 
wire _abc_41356_new_n4139_; 
wire _abc_41356_new_n4140_; 
wire _abc_41356_new_n4141_; 
wire _abc_41356_new_n4142_; 
wire _abc_41356_new_n4143_; 
wire _abc_41356_new_n4144_; 
wire _abc_41356_new_n4145_; 
wire _abc_41356_new_n4146_; 
wire _abc_41356_new_n4147_; 
wire _abc_41356_new_n4148_; 
wire _abc_41356_new_n4149_; 
wire _abc_41356_new_n4150_; 
wire _abc_41356_new_n4151_; 
wire _abc_41356_new_n4152_; 
wire _abc_41356_new_n4153_; 
wire _abc_41356_new_n4154_; 
wire _abc_41356_new_n4155_; 
wire _abc_41356_new_n4156_; 
wire _abc_41356_new_n4157_; 
wire _abc_41356_new_n4158_; 
wire _abc_41356_new_n4159_; 
wire _abc_41356_new_n4160_; 
wire _abc_41356_new_n4161_; 
wire _abc_41356_new_n4162_; 
wire _abc_41356_new_n4163_; 
wire _abc_41356_new_n4164_; 
wire _abc_41356_new_n4165_; 
wire _abc_41356_new_n4166_; 
wire _abc_41356_new_n4167_; 
wire _abc_41356_new_n4168_; 
wire _abc_41356_new_n4169_; 
wire _abc_41356_new_n4170_; 
wire _abc_41356_new_n4171_; 
wire _abc_41356_new_n4172_; 
wire _abc_41356_new_n4173_; 
wire _abc_41356_new_n4174_; 
wire _abc_41356_new_n4175_; 
wire _abc_41356_new_n4176_; 
wire _abc_41356_new_n4177_; 
wire _abc_41356_new_n4178_; 
wire _abc_41356_new_n4179_; 
wire _abc_41356_new_n4180_; 
wire _abc_41356_new_n4181_; 
wire _abc_41356_new_n4182_; 
wire _abc_41356_new_n4183_; 
wire _abc_41356_new_n4184_; 
wire _abc_41356_new_n4185_; 
wire _abc_41356_new_n4186_; 
wire _abc_41356_new_n4187_; 
wire _abc_41356_new_n4188_; 
wire _abc_41356_new_n4189_; 
wire _abc_41356_new_n4190_; 
wire _abc_41356_new_n4191_; 
wire _abc_41356_new_n4192_; 
wire _abc_41356_new_n4193_; 
wire _abc_41356_new_n4194_; 
wire _abc_41356_new_n4195_; 
wire _abc_41356_new_n4196_; 
wire _abc_41356_new_n4197_; 
wire _abc_41356_new_n4198_; 
wire _abc_41356_new_n4199_; 
wire _abc_41356_new_n4200_; 
wire _abc_41356_new_n4202_; 
wire _abc_41356_new_n4203_; 
wire _abc_41356_new_n4204_; 
wire _abc_41356_new_n4205_; 
wire _abc_41356_new_n4206_; 
wire _abc_41356_new_n4207_; 
wire _abc_41356_new_n4208_; 
wire _abc_41356_new_n4209_; 
wire _abc_41356_new_n4210_; 
wire _abc_41356_new_n4211_; 
wire _abc_41356_new_n4212_; 
wire _abc_41356_new_n4213_; 
wire _abc_41356_new_n4214_; 
wire _abc_41356_new_n4215_; 
wire _abc_41356_new_n4216_; 
wire _abc_41356_new_n4217_; 
wire _abc_41356_new_n4218_; 
wire _abc_41356_new_n4219_; 
wire _abc_41356_new_n4220_; 
wire _abc_41356_new_n4221_; 
wire _abc_41356_new_n4222_; 
wire _abc_41356_new_n4223_; 
wire _abc_41356_new_n4224_; 
wire _abc_41356_new_n4225_; 
wire _abc_41356_new_n4226_; 
wire _abc_41356_new_n4227_; 
wire _abc_41356_new_n4228_; 
wire _abc_41356_new_n4229_; 
wire _abc_41356_new_n4230_; 
wire _abc_41356_new_n4231_; 
wire _abc_41356_new_n4232_; 
wire _abc_41356_new_n4233_; 
wire _abc_41356_new_n4234_; 
wire _abc_41356_new_n4235_; 
wire _abc_41356_new_n4236_; 
wire _abc_41356_new_n4237_; 
wire _abc_41356_new_n4238_; 
wire _abc_41356_new_n4239_; 
wire _abc_41356_new_n4240_; 
wire _abc_41356_new_n4241_; 
wire _abc_41356_new_n4242_; 
wire _abc_41356_new_n4243_; 
wire _abc_41356_new_n4245_; 
wire _abc_41356_new_n4246_; 
wire _abc_41356_new_n4247_; 
wire _abc_41356_new_n4248_; 
wire _abc_41356_new_n4249_; 
wire _abc_41356_new_n4250_; 
wire _abc_41356_new_n4251_; 
wire _abc_41356_new_n4252_; 
wire _abc_41356_new_n4253_; 
wire _abc_41356_new_n4254_; 
wire _abc_41356_new_n4255_; 
wire _abc_41356_new_n4256_; 
wire _abc_41356_new_n4257_; 
wire _abc_41356_new_n4258_; 
wire _abc_41356_new_n4259_; 
wire _abc_41356_new_n4260_; 
wire _abc_41356_new_n4261_; 
wire _abc_41356_new_n4262_; 
wire _abc_41356_new_n4263_; 
wire _abc_41356_new_n4264_; 
wire _abc_41356_new_n4265_; 
wire _abc_41356_new_n4266_; 
wire _abc_41356_new_n4267_; 
wire _abc_41356_new_n4268_; 
wire _abc_41356_new_n4269_; 
wire _abc_41356_new_n4270_; 
wire _abc_41356_new_n4271_; 
wire _abc_41356_new_n4272_; 
wire _abc_41356_new_n4273_; 
wire _abc_41356_new_n4274_; 
wire _abc_41356_new_n4275_; 
wire _abc_41356_new_n4276_; 
wire _abc_41356_new_n4277_; 
wire _abc_41356_new_n4278_; 
wire _abc_41356_new_n4279_; 
wire _abc_41356_new_n4280_; 
wire _abc_41356_new_n4281_; 
wire _abc_41356_new_n4282_; 
wire _abc_41356_new_n4283_; 
wire _abc_41356_new_n4284_; 
wire _abc_41356_new_n4285_; 
wire _abc_41356_new_n4286_; 
wire _abc_41356_new_n4288_; 
wire _abc_41356_new_n4289_; 
wire _abc_41356_new_n4290_; 
wire _abc_41356_new_n4291_; 
wire _abc_41356_new_n4292_; 
wire _abc_41356_new_n4293_; 
wire _abc_41356_new_n4294_; 
wire _abc_41356_new_n4295_; 
wire _abc_41356_new_n4296_; 
wire _abc_41356_new_n4297_; 
wire _abc_41356_new_n4298_; 
wire _abc_41356_new_n4299_; 
wire _abc_41356_new_n4300_; 
wire _abc_41356_new_n4301_; 
wire _abc_41356_new_n4302_; 
wire _abc_41356_new_n4303_; 
wire _abc_41356_new_n4304_; 
wire _abc_41356_new_n4305_; 
wire _abc_41356_new_n4306_; 
wire _abc_41356_new_n4307_; 
wire _abc_41356_new_n4308_; 
wire _abc_41356_new_n4309_; 
wire _abc_41356_new_n4310_; 
wire _abc_41356_new_n4311_; 
wire _abc_41356_new_n4312_; 
wire _abc_41356_new_n4313_; 
wire _abc_41356_new_n4314_; 
wire _abc_41356_new_n4315_; 
wire _abc_41356_new_n4316_; 
wire _abc_41356_new_n4317_; 
wire _abc_41356_new_n4318_; 
wire _abc_41356_new_n4319_; 
wire _abc_41356_new_n4320_; 
wire _abc_41356_new_n4321_; 
wire _abc_41356_new_n4322_; 
wire _abc_41356_new_n4323_; 
wire _abc_41356_new_n4324_; 
wire _abc_41356_new_n4325_; 
wire _abc_41356_new_n4326_; 
wire _abc_41356_new_n4327_; 
wire _abc_41356_new_n4328_; 
wire _abc_41356_new_n4329_; 
wire _abc_41356_new_n4331_; 
wire _abc_41356_new_n4332_; 
wire _abc_41356_new_n4333_; 
wire _abc_41356_new_n4334_; 
wire _abc_41356_new_n4335_; 
wire _abc_41356_new_n4336_; 
wire _abc_41356_new_n4337_; 
wire _abc_41356_new_n4338_; 
wire _abc_41356_new_n4339_; 
wire _abc_41356_new_n4340_; 
wire _abc_41356_new_n4341_; 
wire _abc_41356_new_n4342_; 
wire _abc_41356_new_n4343_; 
wire _abc_41356_new_n4344_; 
wire _abc_41356_new_n4345_; 
wire _abc_41356_new_n4346_; 
wire _abc_41356_new_n4347_; 
wire _abc_41356_new_n4348_; 
wire _abc_41356_new_n4349_; 
wire _abc_41356_new_n4350_; 
wire _abc_41356_new_n4351_; 
wire _abc_41356_new_n4352_; 
wire _abc_41356_new_n4353_; 
wire _abc_41356_new_n4354_; 
wire _abc_41356_new_n4355_; 
wire _abc_41356_new_n4356_; 
wire _abc_41356_new_n4357_; 
wire _abc_41356_new_n4358_; 
wire _abc_41356_new_n4359_; 
wire _abc_41356_new_n4360_; 
wire _abc_41356_new_n4361_; 
wire _abc_41356_new_n4362_; 
wire _abc_41356_new_n4363_; 
wire _abc_41356_new_n4364_; 
wire _abc_41356_new_n4365_; 
wire _abc_41356_new_n4366_; 
wire _abc_41356_new_n4367_; 
wire _abc_41356_new_n4368_; 
wire _abc_41356_new_n4369_; 
wire _abc_41356_new_n4370_; 
wire _abc_41356_new_n4371_; 
wire _abc_41356_new_n4372_; 
wire _abc_41356_new_n4374_; 
wire _abc_41356_new_n4375_; 
wire _abc_41356_new_n4376_; 
wire _abc_41356_new_n4377_; 
wire _abc_41356_new_n4378_; 
wire _abc_41356_new_n4379_; 
wire _abc_41356_new_n4380_; 
wire _abc_41356_new_n4381_; 
wire _abc_41356_new_n4382_; 
wire _abc_41356_new_n4383_; 
wire _abc_41356_new_n4384_; 
wire _abc_41356_new_n4385_; 
wire _abc_41356_new_n4386_; 
wire _abc_41356_new_n4387_; 
wire _abc_41356_new_n4388_; 
wire _abc_41356_new_n4389_; 
wire _abc_41356_new_n4390_; 
wire _abc_41356_new_n4391_; 
wire _abc_41356_new_n4392_; 
wire _abc_41356_new_n4393_; 
wire _abc_41356_new_n4394_; 
wire _abc_41356_new_n4395_; 
wire _abc_41356_new_n4396_; 
wire _abc_41356_new_n4397_; 
wire _abc_41356_new_n4398_; 
wire _abc_41356_new_n4399_; 
wire _abc_41356_new_n4400_; 
wire _abc_41356_new_n4401_; 
wire _abc_41356_new_n4402_; 
wire _abc_41356_new_n4403_; 
wire _abc_41356_new_n4404_; 
wire _abc_41356_new_n4405_; 
wire _abc_41356_new_n4406_; 
wire _abc_41356_new_n4407_; 
wire _abc_41356_new_n4408_; 
wire _abc_41356_new_n4409_; 
wire _abc_41356_new_n4410_; 
wire _abc_41356_new_n4411_; 
wire _abc_41356_new_n4412_; 
wire _abc_41356_new_n4413_; 
wire _abc_41356_new_n4414_; 
wire _abc_41356_new_n4415_; 
wire _abc_41356_new_n4417_; 
wire _abc_41356_new_n4418_; 
wire _abc_41356_new_n4419_; 
wire _abc_41356_new_n4420_; 
wire _abc_41356_new_n4421_; 
wire _abc_41356_new_n4422_; 
wire _abc_41356_new_n4423_; 
wire _abc_41356_new_n4424_; 
wire _abc_41356_new_n4425_; 
wire _abc_41356_new_n4426_; 
wire _abc_41356_new_n4427_; 
wire _abc_41356_new_n4428_; 
wire _abc_41356_new_n4429_; 
wire _abc_41356_new_n4430_; 
wire _abc_41356_new_n4431_; 
wire _abc_41356_new_n4432_; 
wire _abc_41356_new_n4433_; 
wire _abc_41356_new_n4434_; 
wire _abc_41356_new_n4435_; 
wire _abc_41356_new_n4436_; 
wire _abc_41356_new_n4437_; 
wire _abc_41356_new_n4438_; 
wire _abc_41356_new_n4439_; 
wire _abc_41356_new_n4440_; 
wire _abc_41356_new_n4441_; 
wire _abc_41356_new_n4442_; 
wire _abc_41356_new_n4443_; 
wire _abc_41356_new_n4444_; 
wire _abc_41356_new_n4445_; 
wire _abc_41356_new_n4446_; 
wire _abc_41356_new_n4447_; 
wire _abc_41356_new_n4448_; 
wire _abc_41356_new_n4449_; 
wire _abc_41356_new_n4450_; 
wire _abc_41356_new_n4451_; 
wire _abc_41356_new_n4452_; 
wire _abc_41356_new_n4453_; 
wire _abc_41356_new_n4454_; 
wire _abc_41356_new_n4455_; 
wire _abc_41356_new_n4456_; 
wire _abc_41356_new_n4457_; 
wire _abc_41356_new_n4459_; 
wire _abc_41356_new_n4460_; 
wire _abc_41356_new_n4461_; 
wire _abc_41356_new_n4462_; 
wire _abc_41356_new_n4463_; 
wire _abc_41356_new_n4464_; 
wire _abc_41356_new_n4465_; 
wire _abc_41356_new_n4466_; 
wire _abc_41356_new_n4467_; 
wire _abc_41356_new_n4468_; 
wire _abc_41356_new_n4469_; 
wire _abc_41356_new_n4470_; 
wire _abc_41356_new_n4471_; 
wire _abc_41356_new_n4472_; 
wire _abc_41356_new_n4473_; 
wire _abc_41356_new_n4474_; 
wire _abc_41356_new_n4475_; 
wire _abc_41356_new_n4476_; 
wire _abc_41356_new_n4477_; 
wire _abc_41356_new_n4478_; 
wire _abc_41356_new_n4479_; 
wire _abc_41356_new_n4480_; 
wire _abc_41356_new_n4481_; 
wire _abc_41356_new_n4482_; 
wire _abc_41356_new_n4483_; 
wire _abc_41356_new_n4484_; 
wire _abc_41356_new_n4485_; 
wire _abc_41356_new_n4486_; 
wire _abc_41356_new_n4487_; 
wire _abc_41356_new_n4488_; 
wire _abc_41356_new_n4489_; 
wire _abc_41356_new_n4490_; 
wire _abc_41356_new_n4491_; 
wire _abc_41356_new_n4492_; 
wire _abc_41356_new_n4493_; 
wire _abc_41356_new_n4494_; 
wire _abc_41356_new_n4495_; 
wire _abc_41356_new_n4496_; 
wire _abc_41356_new_n4497_; 
wire _abc_41356_new_n4498_; 
wire _abc_41356_new_n4499_; 
wire _abc_41356_new_n4500_; 
wire _abc_41356_new_n4502_; 
wire _abc_41356_new_n4503_; 
wire _abc_41356_new_n4504_; 
wire _abc_41356_new_n4505_; 
wire _abc_41356_new_n4506_; 
wire _abc_41356_new_n4507_; 
wire _abc_41356_new_n4508_; 
wire _abc_41356_new_n4509_; 
wire _abc_41356_new_n4510_; 
wire _abc_41356_new_n4511_; 
wire _abc_41356_new_n4512_; 
wire _abc_41356_new_n4513_; 
wire _abc_41356_new_n4514_; 
wire _abc_41356_new_n4515_; 
wire _abc_41356_new_n4516_; 
wire _abc_41356_new_n4517_; 
wire _abc_41356_new_n4518_; 
wire _abc_41356_new_n4519_; 
wire _abc_41356_new_n4520_; 
wire _abc_41356_new_n4521_; 
wire _abc_41356_new_n4522_; 
wire _abc_41356_new_n4523_; 
wire _abc_41356_new_n4524_; 
wire _abc_41356_new_n4525_; 
wire _abc_41356_new_n4526_; 
wire _abc_41356_new_n4527_; 
wire _abc_41356_new_n4528_; 
wire _abc_41356_new_n4529_; 
wire _abc_41356_new_n4530_; 
wire _abc_41356_new_n4531_; 
wire _abc_41356_new_n4532_; 
wire _abc_41356_new_n4533_; 
wire _abc_41356_new_n4534_; 
wire _abc_41356_new_n4535_; 
wire _abc_41356_new_n4536_; 
wire _abc_41356_new_n4537_; 
wire _abc_41356_new_n4538_; 
wire _abc_41356_new_n4539_; 
wire _abc_41356_new_n4540_; 
wire _abc_41356_new_n4541_; 
wire _abc_41356_new_n4543_; 
wire _abc_41356_new_n4544_; 
wire _abc_41356_new_n4545_; 
wire _abc_41356_new_n4546_; 
wire _abc_41356_new_n4547_; 
wire _abc_41356_new_n4548_; 
wire _abc_41356_new_n4549_; 
wire _abc_41356_new_n4550_; 
wire _abc_41356_new_n4551_; 
wire _abc_41356_new_n4552_; 
wire _abc_41356_new_n4553_; 
wire _abc_41356_new_n4554_; 
wire _abc_41356_new_n4555_; 
wire _abc_41356_new_n4556_; 
wire _abc_41356_new_n4557_; 
wire _abc_41356_new_n4558_; 
wire _abc_41356_new_n4559_; 
wire _abc_41356_new_n4560_; 
wire _abc_41356_new_n4561_; 
wire _abc_41356_new_n4562_; 
wire _abc_41356_new_n4563_; 
wire _abc_41356_new_n4564_; 
wire _abc_41356_new_n4565_; 
wire _abc_41356_new_n4566_; 
wire _abc_41356_new_n4567_; 
wire _abc_41356_new_n4568_; 
wire _abc_41356_new_n4569_; 
wire _abc_41356_new_n4570_; 
wire _abc_41356_new_n4571_; 
wire _abc_41356_new_n4572_; 
wire _abc_41356_new_n4573_; 
wire _abc_41356_new_n4574_; 
wire _abc_41356_new_n4575_; 
wire _abc_41356_new_n4576_; 
wire _abc_41356_new_n4577_; 
wire _abc_41356_new_n4578_; 
wire _abc_41356_new_n4579_; 
wire _abc_41356_new_n4580_; 
wire _abc_41356_new_n4581_; 
wire _abc_41356_new_n4582_; 
wire _abc_41356_new_n4584_; 
wire _abc_41356_new_n4585_; 
wire _abc_41356_new_n4586_; 
wire _abc_41356_new_n4587_; 
wire _abc_41356_new_n4588_; 
wire _abc_41356_new_n4589_; 
wire _abc_41356_new_n4590_; 
wire _abc_41356_new_n4591_; 
wire _abc_41356_new_n4592_; 
wire _abc_41356_new_n4593_; 
wire _abc_41356_new_n4594_; 
wire _abc_41356_new_n4595_; 
wire _abc_41356_new_n4596_; 
wire _abc_41356_new_n4597_; 
wire _abc_41356_new_n4598_; 
wire _abc_41356_new_n4599_; 
wire _abc_41356_new_n4600_; 
wire _abc_41356_new_n4601_; 
wire _abc_41356_new_n4602_; 
wire _abc_41356_new_n4603_; 
wire _abc_41356_new_n4604_; 
wire _abc_41356_new_n4605_; 
wire _abc_41356_new_n4606_; 
wire _abc_41356_new_n4607_; 
wire _abc_41356_new_n4608_; 
wire _abc_41356_new_n4609_; 
wire _abc_41356_new_n4610_; 
wire _abc_41356_new_n4611_; 
wire _abc_41356_new_n4612_; 
wire _abc_41356_new_n4613_; 
wire _abc_41356_new_n4614_; 
wire _abc_41356_new_n4615_; 
wire _abc_41356_new_n4616_; 
wire _abc_41356_new_n4617_; 
wire _abc_41356_new_n4618_; 
wire _abc_41356_new_n4619_; 
wire _abc_41356_new_n4620_; 
wire _abc_41356_new_n4621_; 
wire _abc_41356_new_n4622_; 
wire _abc_41356_new_n4623_; 
wire _abc_41356_new_n4625_; 
wire _abc_41356_new_n4626_; 
wire _abc_41356_new_n4627_; 
wire _abc_41356_new_n4628_; 
wire _abc_41356_new_n4629_; 
wire _abc_41356_new_n4630_; 
wire _abc_41356_new_n4631_; 
wire _abc_41356_new_n4632_; 
wire _abc_41356_new_n4633_; 
wire _abc_41356_new_n4634_; 
wire _abc_41356_new_n4635_; 
wire _abc_41356_new_n4636_; 
wire _abc_41356_new_n4637_; 
wire _abc_41356_new_n4638_; 
wire _abc_41356_new_n4639_; 
wire _abc_41356_new_n4640_; 
wire _abc_41356_new_n4641_; 
wire _abc_41356_new_n4642_; 
wire _abc_41356_new_n4643_; 
wire _abc_41356_new_n4644_; 
wire _abc_41356_new_n4645_; 
wire _abc_41356_new_n4646_; 
wire _abc_41356_new_n4647_; 
wire _abc_41356_new_n4648_; 
wire _abc_41356_new_n4649_; 
wire _abc_41356_new_n4650_; 
wire _abc_41356_new_n4651_; 
wire _abc_41356_new_n4652_; 
wire _abc_41356_new_n4653_; 
wire _abc_41356_new_n4654_; 
wire _abc_41356_new_n4655_; 
wire _abc_41356_new_n4656_; 
wire _abc_41356_new_n4657_; 
wire _abc_41356_new_n4658_; 
wire _abc_41356_new_n4659_; 
wire _abc_41356_new_n4660_; 
wire _abc_41356_new_n4661_; 
wire _abc_41356_new_n4662_; 
wire _abc_41356_new_n4663_; 
wire _abc_41356_new_n4665_; 
wire _abc_41356_new_n4666_; 
wire _abc_41356_new_n4667_; 
wire _abc_41356_new_n4668_; 
wire _abc_41356_new_n4669_; 
wire _abc_41356_new_n4670_; 
wire _abc_41356_new_n4671_; 
wire _abc_41356_new_n4672_; 
wire _abc_41356_new_n4673_; 
wire _abc_41356_new_n4674_; 
wire _abc_41356_new_n4675_; 
wire _abc_41356_new_n4676_; 
wire _abc_41356_new_n4677_; 
wire _abc_41356_new_n4678_; 
wire _abc_41356_new_n4679_; 
wire _abc_41356_new_n4680_; 
wire _abc_41356_new_n4681_; 
wire _abc_41356_new_n4682_; 
wire _abc_41356_new_n4683_; 
wire _abc_41356_new_n4684_; 
wire _abc_41356_new_n4685_; 
wire _abc_41356_new_n4686_; 
wire _abc_41356_new_n4687_; 
wire _abc_41356_new_n4688_; 
wire _abc_41356_new_n4689_; 
wire _abc_41356_new_n4690_; 
wire _abc_41356_new_n4691_; 
wire _abc_41356_new_n4692_; 
wire _abc_41356_new_n4693_; 
wire _abc_41356_new_n4694_; 
wire _abc_41356_new_n4695_; 
wire _abc_41356_new_n4696_; 
wire _abc_41356_new_n4697_; 
wire _abc_41356_new_n4698_; 
wire _abc_41356_new_n4699_; 
wire _abc_41356_new_n4700_; 
wire _abc_41356_new_n4702_; 
wire _abc_41356_new_n4703_; 
wire _abc_41356_new_n4704_; 
wire _abc_41356_new_n4705_; 
wire _abc_41356_new_n4706_; 
wire _abc_41356_new_n4707_; 
wire _abc_41356_new_n4708_; 
wire _abc_41356_new_n4709_; 
wire _abc_41356_new_n4710_; 
wire _abc_41356_new_n4711_; 
wire _abc_41356_new_n4712_; 
wire _abc_41356_new_n4713_; 
wire _abc_41356_new_n4714_; 
wire _abc_41356_new_n4715_; 
wire _abc_41356_new_n4716_; 
wire _abc_41356_new_n4717_; 
wire _abc_41356_new_n4718_; 
wire _abc_41356_new_n4719_; 
wire _abc_41356_new_n4720_; 
wire _abc_41356_new_n4721_; 
wire _abc_41356_new_n4722_; 
wire _abc_41356_new_n4723_; 
wire _abc_41356_new_n4724_; 
wire _abc_41356_new_n4725_; 
wire _abc_41356_new_n4726_; 
wire _abc_41356_new_n4727_; 
wire _abc_41356_new_n4728_; 
wire _abc_41356_new_n4729_; 
wire _abc_41356_new_n4730_; 
wire _abc_41356_new_n4731_; 
wire _abc_41356_new_n4732_; 
wire _abc_41356_new_n4733_; 
wire _abc_41356_new_n4734_; 
wire _abc_41356_new_n4735_; 
wire _abc_41356_new_n4736_; 
wire _abc_41356_new_n4737_; 
wire _abc_41356_new_n4739_; 
wire _abc_41356_new_n4740_; 
wire _abc_41356_new_n4741_; 
wire _abc_41356_new_n4742_; 
wire _abc_41356_new_n4743_; 
wire _abc_41356_new_n4744_; 
wire _abc_41356_new_n4745_; 
wire _abc_41356_new_n4746_; 
wire _abc_41356_new_n4747_; 
wire _abc_41356_new_n4748_; 
wire _abc_41356_new_n4749_; 
wire _abc_41356_new_n4750_; 
wire _abc_41356_new_n4751_; 
wire _abc_41356_new_n4752_; 
wire _abc_41356_new_n4753_; 
wire _abc_41356_new_n4754_; 
wire _abc_41356_new_n4755_; 
wire _abc_41356_new_n4756_; 
wire _abc_41356_new_n4757_; 
wire _abc_41356_new_n4758_; 
wire _abc_41356_new_n4759_; 
wire _abc_41356_new_n4760_; 
wire _abc_41356_new_n4761_; 
wire _abc_41356_new_n4762_; 
wire _abc_41356_new_n4763_; 
wire _abc_41356_new_n4764_; 
wire _abc_41356_new_n4765_; 
wire _abc_41356_new_n4766_; 
wire _abc_41356_new_n4767_; 
wire _abc_41356_new_n4768_; 
wire _abc_41356_new_n4769_; 
wire _abc_41356_new_n4770_; 
wire _abc_41356_new_n4771_; 
wire _abc_41356_new_n4772_; 
wire _abc_41356_new_n4773_; 
wire _abc_41356_new_n4774_; 
wire _abc_41356_new_n4775_; 
wire _abc_41356_new_n4776_; 
wire _abc_41356_new_n4778_; 
wire _abc_41356_new_n4779_; 
wire _abc_41356_new_n4780_; 
wire _abc_41356_new_n4781_; 
wire _abc_41356_new_n4782_; 
wire _abc_41356_new_n4783_; 
wire _abc_41356_new_n4784_; 
wire _abc_41356_new_n4785_; 
wire _abc_41356_new_n4786_; 
wire _abc_41356_new_n4787_; 
wire _abc_41356_new_n4788_; 
wire _abc_41356_new_n4789_; 
wire _abc_41356_new_n4790_; 
wire _abc_41356_new_n4791_; 
wire _abc_41356_new_n4792_; 
wire _abc_41356_new_n4793_; 
wire _abc_41356_new_n4794_; 
wire _abc_41356_new_n4795_; 
wire _abc_41356_new_n4796_; 
wire _abc_41356_new_n4797_; 
wire _abc_41356_new_n4798_; 
wire _abc_41356_new_n4799_; 
wire _abc_41356_new_n4800_; 
wire _abc_41356_new_n4801_; 
wire _abc_41356_new_n4802_; 
wire _abc_41356_new_n4803_; 
wire _abc_41356_new_n4804_; 
wire _abc_41356_new_n4805_; 
wire _abc_41356_new_n4806_; 
wire _abc_41356_new_n4807_; 
wire _abc_41356_new_n4808_; 
wire _abc_41356_new_n4809_; 
wire _abc_41356_new_n4810_; 
wire _abc_41356_new_n4811_; 
wire _abc_41356_new_n4812_; 
wire _abc_41356_new_n4813_; 
wire _abc_41356_new_n4814_; 
wire _abc_41356_new_n4815_; 
wire _abc_41356_new_n4816_; 
wire _abc_41356_new_n4817_; 
wire _abc_41356_new_n4819_; 
wire _abc_41356_new_n4820_; 
wire _abc_41356_new_n4821_; 
wire _abc_41356_new_n4822_; 
wire _abc_41356_new_n4823_; 
wire _abc_41356_new_n4824_; 
wire _abc_41356_new_n4825_; 
wire _abc_41356_new_n4826_; 
wire _abc_41356_new_n4827_; 
wire _abc_41356_new_n4828_; 
wire _abc_41356_new_n4829_; 
wire _abc_41356_new_n4830_; 
wire _abc_41356_new_n4831_; 
wire _abc_41356_new_n4832_; 
wire _abc_41356_new_n4833_; 
wire _abc_41356_new_n4834_; 
wire _abc_41356_new_n4835_; 
wire _abc_41356_new_n4836_; 
wire _abc_41356_new_n4837_; 
wire _abc_41356_new_n4838_; 
wire _abc_41356_new_n4839_; 
wire _abc_41356_new_n4840_; 
wire _abc_41356_new_n4841_; 
wire _abc_41356_new_n4842_; 
wire _abc_41356_new_n4843_; 
wire _abc_41356_new_n4844_; 
wire _abc_41356_new_n4845_; 
wire _abc_41356_new_n4846_; 
wire _abc_41356_new_n4847_; 
wire _abc_41356_new_n4848_; 
wire _abc_41356_new_n4849_; 
wire _abc_41356_new_n4850_; 
wire _abc_41356_new_n4851_; 
wire _abc_41356_new_n4852_; 
wire _abc_41356_new_n4853_; 
wire _abc_41356_new_n4854_; 
wire _abc_41356_new_n4856_; 
wire _abc_41356_new_n4857_; 
wire _abc_41356_new_n4858_; 
wire _abc_41356_new_n4859_; 
wire _abc_41356_new_n4860_; 
wire _abc_41356_new_n4861_; 
wire _abc_41356_new_n4862_; 
wire _abc_41356_new_n4863_; 
wire _abc_41356_new_n4864_; 
wire _abc_41356_new_n4865_; 
wire _abc_41356_new_n4866_; 
wire _abc_41356_new_n4867_; 
wire _abc_41356_new_n4868_; 
wire _abc_41356_new_n4869_; 
wire _abc_41356_new_n4870_; 
wire _abc_41356_new_n4871_; 
wire _abc_41356_new_n4872_; 
wire _abc_41356_new_n4873_; 
wire _abc_41356_new_n4874_; 
wire _abc_41356_new_n4875_; 
wire _abc_41356_new_n4876_; 
wire _abc_41356_new_n4877_; 
wire _abc_41356_new_n4878_; 
wire _abc_41356_new_n4879_; 
wire _abc_41356_new_n4880_; 
wire _abc_41356_new_n4881_; 
wire _abc_41356_new_n4882_; 
wire _abc_41356_new_n4883_; 
wire _abc_41356_new_n4884_; 
wire _abc_41356_new_n4885_; 
wire _abc_41356_new_n4886_; 
wire _abc_41356_new_n4887_; 
wire _abc_41356_new_n4888_; 
wire _abc_41356_new_n4889_; 
wire _abc_41356_new_n4890_; 
wire _abc_41356_new_n4891_; 
wire _abc_41356_new_n4893_; 
wire _abc_41356_new_n4894_; 
wire _abc_41356_new_n4895_; 
wire _abc_41356_new_n4896_; 
wire _abc_41356_new_n4897_; 
wire _abc_41356_new_n4898_; 
wire _abc_41356_new_n4899_; 
wire _abc_41356_new_n4900_; 
wire _abc_41356_new_n4901_; 
wire _abc_41356_new_n4902_; 
wire _abc_41356_new_n4903_; 
wire _abc_41356_new_n4904_; 
wire _abc_41356_new_n4905_; 
wire _abc_41356_new_n4906_; 
wire _abc_41356_new_n4907_; 
wire _abc_41356_new_n4908_; 
wire _abc_41356_new_n4909_; 
wire _abc_41356_new_n4910_; 
wire _abc_41356_new_n4911_; 
wire _abc_41356_new_n4912_; 
wire _abc_41356_new_n4913_; 
wire _abc_41356_new_n4914_; 
wire _abc_41356_new_n4915_; 
wire _abc_41356_new_n4916_; 
wire _abc_41356_new_n4917_; 
wire _abc_41356_new_n4918_; 
wire _abc_41356_new_n4919_; 
wire _abc_41356_new_n4920_; 
wire _abc_41356_new_n4921_; 
wire _abc_41356_new_n4922_; 
wire _abc_41356_new_n4923_; 
wire _abc_41356_new_n4924_; 
wire _abc_41356_new_n4925_; 
wire _abc_41356_new_n4926_; 
wire _abc_41356_new_n4927_; 
wire _abc_41356_new_n4929_; 
wire _abc_41356_new_n4930_; 
wire _abc_41356_new_n4931_; 
wire _abc_41356_new_n4932_; 
wire _abc_41356_new_n4933_; 
wire _abc_41356_new_n4934_; 
wire _abc_41356_new_n4935_; 
wire _abc_41356_new_n4936_; 
wire _abc_41356_new_n4937_; 
wire _abc_41356_new_n4938_; 
wire _abc_41356_new_n4939_; 
wire _abc_41356_new_n4940_; 
wire _abc_41356_new_n4941_; 
wire _abc_41356_new_n4942_; 
wire _abc_41356_new_n4943_; 
wire _abc_41356_new_n4944_; 
wire _abc_41356_new_n4945_; 
wire _abc_41356_new_n4946_; 
wire _abc_41356_new_n4947_; 
wire _abc_41356_new_n4948_; 
wire _abc_41356_new_n4949_; 
wire _abc_41356_new_n4950_; 
wire _abc_41356_new_n4951_; 
wire _abc_41356_new_n4952_; 
wire _abc_41356_new_n4953_; 
wire _abc_41356_new_n4954_; 
wire _abc_41356_new_n4955_; 
wire _abc_41356_new_n4956_; 
wire _abc_41356_new_n4957_; 
wire _abc_41356_new_n4958_; 
wire _abc_41356_new_n4959_; 
wire _abc_41356_new_n4960_; 
wire _abc_41356_new_n4961_; 
wire _abc_41356_new_n4962_; 
wire _abc_41356_new_n4963_; 
wire _abc_41356_new_n4964_; 
wire _abc_41356_new_n4966_; 
wire _abc_41356_new_n4967_; 
wire _abc_41356_new_n4968_; 
wire _abc_41356_new_n4969_; 
wire _abc_41356_new_n4970_; 
wire _abc_41356_new_n4971_; 
wire _abc_41356_new_n4972_; 
wire _abc_41356_new_n4973_; 
wire _abc_41356_new_n4974_; 
wire _abc_41356_new_n4975_; 
wire _abc_41356_new_n4976_; 
wire _abc_41356_new_n4977_; 
wire _abc_41356_new_n4978_; 
wire _abc_41356_new_n4979_; 
wire _abc_41356_new_n4980_; 
wire _abc_41356_new_n4981_; 
wire _abc_41356_new_n4982_; 
wire _abc_41356_new_n4983_; 
wire _abc_41356_new_n4984_; 
wire _abc_41356_new_n4985_; 
wire _abc_41356_new_n4986_; 
wire _abc_41356_new_n4987_; 
wire _abc_41356_new_n4988_; 
wire _abc_41356_new_n4989_; 
wire _abc_41356_new_n4990_; 
wire _abc_41356_new_n4991_; 
wire _abc_41356_new_n4992_; 
wire _abc_41356_new_n4993_; 
wire _abc_41356_new_n4994_; 
wire _abc_41356_new_n4995_; 
wire _abc_41356_new_n4996_; 
wire _abc_41356_new_n4997_; 
wire _abc_41356_new_n4998_; 
wire _abc_41356_new_n4999_; 
wire _abc_41356_new_n5000_; 
wire _abc_41356_new_n5001_; 
wire _abc_41356_new_n5002_; 
wire _abc_41356_new_n5004_; 
wire _abc_41356_new_n5005_; 
wire _abc_41356_new_n5006_; 
wire _abc_41356_new_n5007_; 
wire _abc_41356_new_n5008_; 
wire _abc_41356_new_n5009_; 
wire _abc_41356_new_n5010_; 
wire _abc_41356_new_n5011_; 
wire _abc_41356_new_n5012_; 
wire _abc_41356_new_n5013_; 
wire _abc_41356_new_n5014_; 
wire _abc_41356_new_n5015_; 
wire _abc_41356_new_n5016_; 
wire _abc_41356_new_n5017_; 
wire _abc_41356_new_n5018_; 
wire _abc_41356_new_n5019_; 
wire _abc_41356_new_n501_; 
wire _abc_41356_new_n5020_; 
wire _abc_41356_new_n5021_; 
wire _abc_41356_new_n5022_; 
wire _abc_41356_new_n5023_; 
wire _abc_41356_new_n5024_; 
wire _abc_41356_new_n5025_; 
wire _abc_41356_new_n5026_; 
wire _abc_41356_new_n5027_; 
wire _abc_41356_new_n5028_; 
wire _abc_41356_new_n5029_; 
wire _abc_41356_new_n502_; 
wire _abc_41356_new_n5030_; 
wire _abc_41356_new_n5031_; 
wire _abc_41356_new_n5032_; 
wire _abc_41356_new_n5033_; 
wire _abc_41356_new_n5034_; 
wire _abc_41356_new_n5035_; 
wire _abc_41356_new_n5036_; 
wire _abc_41356_new_n5037_; 
wire _abc_41356_new_n5038_; 
wire _abc_41356_new_n5039_; 
wire _abc_41356_new_n503_; 
wire _abc_41356_new_n5041_; 
wire _abc_41356_new_n5042_; 
wire _abc_41356_new_n5043_; 
wire _abc_41356_new_n5044_; 
wire _abc_41356_new_n5045_; 
wire _abc_41356_new_n5046_; 
wire _abc_41356_new_n5047_; 
wire _abc_41356_new_n5048_; 
wire _abc_41356_new_n5049_; 
wire _abc_41356_new_n504_; 
wire _abc_41356_new_n5050_; 
wire _abc_41356_new_n5051_; 
wire _abc_41356_new_n5052_; 
wire _abc_41356_new_n5053_; 
wire _abc_41356_new_n5054_; 
wire _abc_41356_new_n5055_; 
wire _abc_41356_new_n5056_; 
wire _abc_41356_new_n5057_; 
wire _abc_41356_new_n5058_; 
wire _abc_41356_new_n5059_; 
wire _abc_41356_new_n505_; 
wire _abc_41356_new_n5060_; 
wire _abc_41356_new_n5061_; 
wire _abc_41356_new_n5062_; 
wire _abc_41356_new_n5063_; 
wire _abc_41356_new_n5064_; 
wire _abc_41356_new_n5065_; 
wire _abc_41356_new_n5066_; 
wire _abc_41356_new_n5067_; 
wire _abc_41356_new_n5068_; 
wire _abc_41356_new_n5069_; 
wire _abc_41356_new_n506_; 
wire _abc_41356_new_n5070_; 
wire _abc_41356_new_n5071_; 
wire _abc_41356_new_n5072_; 
wire _abc_41356_new_n5073_; 
wire _abc_41356_new_n5074_; 
wire _abc_41356_new_n5075_; 
wire _abc_41356_new_n5076_; 
wire _abc_41356_new_n5078_; 
wire _abc_41356_new_n5079_; 
wire _abc_41356_new_n507_; 
wire _abc_41356_new_n5080_; 
wire _abc_41356_new_n5081_; 
wire _abc_41356_new_n5082_; 
wire _abc_41356_new_n5083_; 
wire _abc_41356_new_n5084_; 
wire _abc_41356_new_n5085_; 
wire _abc_41356_new_n5086_; 
wire _abc_41356_new_n5087_; 
wire _abc_41356_new_n5088_; 
wire _abc_41356_new_n5089_; 
wire _abc_41356_new_n508_; 
wire _abc_41356_new_n5090_; 
wire _abc_41356_new_n5091_; 
wire _abc_41356_new_n5092_; 
wire _abc_41356_new_n5093_; 
wire _abc_41356_new_n5094_; 
wire _abc_41356_new_n5095_; 
wire _abc_41356_new_n5096_; 
wire _abc_41356_new_n5097_; 
wire _abc_41356_new_n5098_; 
wire _abc_41356_new_n5099_; 
wire _abc_41356_new_n509_; 
wire _abc_41356_new_n5100_; 
wire _abc_41356_new_n5101_; 
wire _abc_41356_new_n5102_; 
wire _abc_41356_new_n5103_; 
wire _abc_41356_new_n5104_; 
wire _abc_41356_new_n5105_; 
wire _abc_41356_new_n5106_; 
wire _abc_41356_new_n5107_; 
wire _abc_41356_new_n5108_; 
wire _abc_41356_new_n5109_; 
wire _abc_41356_new_n510_; 
wire _abc_41356_new_n5110_; 
wire _abc_41356_new_n5111_; 
wire _abc_41356_new_n5112_; 
wire _abc_41356_new_n5113_; 
wire _abc_41356_new_n5115_; 
wire _abc_41356_new_n5116_; 
wire _abc_41356_new_n5117_; 
wire _abc_41356_new_n5118_; 
wire _abc_41356_new_n5119_; 
wire _abc_41356_new_n511_; 
wire _abc_41356_new_n5120_; 
wire _abc_41356_new_n5121_; 
wire _abc_41356_new_n5122_; 
wire _abc_41356_new_n5123_; 
wire _abc_41356_new_n5124_; 
wire _abc_41356_new_n5125_; 
wire _abc_41356_new_n5126_; 
wire _abc_41356_new_n5127_; 
wire _abc_41356_new_n5128_; 
wire _abc_41356_new_n5129_; 
wire _abc_41356_new_n512_; 
wire _abc_41356_new_n5130_; 
wire _abc_41356_new_n5131_; 
wire _abc_41356_new_n5132_; 
wire _abc_41356_new_n5133_; 
wire _abc_41356_new_n5134_; 
wire _abc_41356_new_n5135_; 
wire _abc_41356_new_n5136_; 
wire _abc_41356_new_n5137_; 
wire _abc_41356_new_n5138_; 
wire _abc_41356_new_n5139_; 
wire _abc_41356_new_n513_; 
wire _abc_41356_new_n5140_; 
wire _abc_41356_new_n5141_; 
wire _abc_41356_new_n5142_; 
wire _abc_41356_new_n5143_; 
wire _abc_41356_new_n5144_; 
wire _abc_41356_new_n5145_; 
wire _abc_41356_new_n5146_; 
wire _abc_41356_new_n5147_; 
wire _abc_41356_new_n5148_; 
wire _abc_41356_new_n5149_; 
wire _abc_41356_new_n514_; 
wire _abc_41356_new_n5150_; 
wire _abc_41356_new_n5152_; 
wire _abc_41356_new_n5153_; 
wire _abc_41356_new_n5154_; 
wire _abc_41356_new_n5155_; 
wire _abc_41356_new_n5156_; 
wire _abc_41356_new_n5157_; 
wire _abc_41356_new_n5158_; 
wire _abc_41356_new_n5159_; 
wire _abc_41356_new_n515_; 
wire _abc_41356_new_n5160_; 
wire _abc_41356_new_n5161_; 
wire _abc_41356_new_n5162_; 
wire _abc_41356_new_n5163_; 
wire _abc_41356_new_n5164_; 
wire _abc_41356_new_n5165_; 
wire _abc_41356_new_n5166_; 
wire _abc_41356_new_n5167_; 
wire _abc_41356_new_n5168_; 
wire _abc_41356_new_n5169_; 
wire _abc_41356_new_n516_; 
wire _abc_41356_new_n5170_; 
wire _abc_41356_new_n5171_; 
wire _abc_41356_new_n5172_; 
wire _abc_41356_new_n5173_; 
wire _abc_41356_new_n5174_; 
wire _abc_41356_new_n5175_; 
wire _abc_41356_new_n5176_; 
wire _abc_41356_new_n5177_; 
wire _abc_41356_new_n5178_; 
wire _abc_41356_new_n5179_; 
wire _abc_41356_new_n517_; 
wire _abc_41356_new_n5180_; 
wire _abc_41356_new_n5181_; 
wire _abc_41356_new_n5182_; 
wire _abc_41356_new_n5183_; 
wire _abc_41356_new_n5184_; 
wire _abc_41356_new_n5185_; 
wire _abc_41356_new_n5186_; 
wire _abc_41356_new_n5187_; 
wire _abc_41356_new_n5189_; 
wire _abc_41356_new_n518_; 
wire _abc_41356_new_n5190_; 
wire _abc_41356_new_n5191_; 
wire _abc_41356_new_n5192_; 
wire _abc_41356_new_n5193_; 
wire _abc_41356_new_n5194_; 
wire _abc_41356_new_n5195_; 
wire _abc_41356_new_n5196_; 
wire _abc_41356_new_n5197_; 
wire _abc_41356_new_n5198_; 
wire _abc_41356_new_n5199_; 
wire _abc_41356_new_n519_; 
wire _abc_41356_new_n5200_; 
wire _abc_41356_new_n5201_; 
wire _abc_41356_new_n5202_; 
wire _abc_41356_new_n5203_; 
wire _abc_41356_new_n5204_; 
wire _abc_41356_new_n5205_; 
wire _abc_41356_new_n5206_; 
wire _abc_41356_new_n5207_; 
wire _abc_41356_new_n5208_; 
wire _abc_41356_new_n5209_; 
wire _abc_41356_new_n520_; 
wire _abc_41356_new_n5210_; 
wire _abc_41356_new_n5211_; 
wire _abc_41356_new_n5212_; 
wire _abc_41356_new_n5213_; 
wire _abc_41356_new_n5214_; 
wire _abc_41356_new_n5215_; 
wire _abc_41356_new_n5216_; 
wire _abc_41356_new_n5217_; 
wire _abc_41356_new_n5218_; 
wire _abc_41356_new_n5219_; 
wire _abc_41356_new_n521_; 
wire _abc_41356_new_n5220_; 
wire _abc_41356_new_n5221_; 
wire _abc_41356_new_n5222_; 
wire _abc_41356_new_n5223_; 
wire _abc_41356_new_n5224_; 
wire _abc_41356_new_n5226_; 
wire _abc_41356_new_n5227_; 
wire _abc_41356_new_n5228_; 
wire _abc_41356_new_n5229_; 
wire _abc_41356_new_n522_; 
wire _abc_41356_new_n5230_; 
wire _abc_41356_new_n5231_; 
wire _abc_41356_new_n5232_; 
wire _abc_41356_new_n5233_; 
wire _abc_41356_new_n5234_; 
wire _abc_41356_new_n5235_; 
wire _abc_41356_new_n5236_; 
wire _abc_41356_new_n5237_; 
wire _abc_41356_new_n5238_; 
wire _abc_41356_new_n5239_; 
wire _abc_41356_new_n523_; 
wire _abc_41356_new_n5240_; 
wire _abc_41356_new_n5241_; 
wire _abc_41356_new_n5242_; 
wire _abc_41356_new_n5243_; 
wire _abc_41356_new_n5244_; 
wire _abc_41356_new_n5245_; 
wire _abc_41356_new_n5246_; 
wire _abc_41356_new_n5247_; 
wire _abc_41356_new_n5248_; 
wire _abc_41356_new_n5249_; 
wire _abc_41356_new_n524_; 
wire _abc_41356_new_n5250_; 
wire _abc_41356_new_n5251_; 
wire _abc_41356_new_n5252_; 
wire _abc_41356_new_n5253_; 
wire _abc_41356_new_n5254_; 
wire _abc_41356_new_n5255_; 
wire _abc_41356_new_n5256_; 
wire _abc_41356_new_n5257_; 
wire _abc_41356_new_n5258_; 
wire _abc_41356_new_n5259_; 
wire _abc_41356_new_n525_; 
wire _abc_41356_new_n5260_; 
wire _abc_41356_new_n5261_; 
wire _abc_41356_new_n5263_; 
wire _abc_41356_new_n5264_; 
wire _abc_41356_new_n5265_; 
wire _abc_41356_new_n5266_; 
wire _abc_41356_new_n5267_; 
wire _abc_41356_new_n5268_; 
wire _abc_41356_new_n5269_; 
wire _abc_41356_new_n526_; 
wire _abc_41356_new_n5270_; 
wire _abc_41356_new_n5271_; 
wire _abc_41356_new_n5272_; 
wire _abc_41356_new_n5273_; 
wire _abc_41356_new_n5274_; 
wire _abc_41356_new_n5275_; 
wire _abc_41356_new_n5276_; 
wire _abc_41356_new_n5277_; 
wire _abc_41356_new_n5278_; 
wire _abc_41356_new_n5279_; 
wire _abc_41356_new_n527_; 
wire _abc_41356_new_n5280_; 
wire _abc_41356_new_n5281_; 
wire _abc_41356_new_n5282_; 
wire _abc_41356_new_n5283_; 
wire _abc_41356_new_n5284_; 
wire _abc_41356_new_n5285_; 
wire _abc_41356_new_n5286_; 
wire _abc_41356_new_n5287_; 
wire _abc_41356_new_n5288_; 
wire _abc_41356_new_n5289_; 
wire _abc_41356_new_n528_; 
wire _abc_41356_new_n5290_; 
wire _abc_41356_new_n5291_; 
wire _abc_41356_new_n5292_; 
wire _abc_41356_new_n5293_; 
wire _abc_41356_new_n5294_; 
wire _abc_41356_new_n5295_; 
wire _abc_41356_new_n5296_; 
wire _abc_41356_new_n5297_; 
wire _abc_41356_new_n5298_; 
wire _abc_41356_new_n5299_; 
wire _abc_41356_new_n529_; 
wire _abc_41356_new_n5301_; 
wire _abc_41356_new_n5302_; 
wire _abc_41356_new_n5303_; 
wire _abc_41356_new_n5304_; 
wire _abc_41356_new_n5305_; 
wire _abc_41356_new_n5306_; 
wire _abc_41356_new_n5307_; 
wire _abc_41356_new_n5308_; 
wire _abc_41356_new_n5309_; 
wire _abc_41356_new_n530_; 
wire _abc_41356_new_n5310_; 
wire _abc_41356_new_n5311_; 
wire _abc_41356_new_n5312_; 
wire _abc_41356_new_n5313_; 
wire _abc_41356_new_n5314_; 
wire _abc_41356_new_n5315_; 
wire _abc_41356_new_n5316_; 
wire _abc_41356_new_n5317_; 
wire _abc_41356_new_n5318_; 
wire _abc_41356_new_n5319_; 
wire _abc_41356_new_n531_; 
wire _abc_41356_new_n5320_; 
wire _abc_41356_new_n5321_; 
wire _abc_41356_new_n5322_; 
wire _abc_41356_new_n5323_; 
wire _abc_41356_new_n5324_; 
wire _abc_41356_new_n5325_; 
wire _abc_41356_new_n5326_; 
wire _abc_41356_new_n5327_; 
wire _abc_41356_new_n5328_; 
wire _abc_41356_new_n5329_; 
wire _abc_41356_new_n532_; 
wire _abc_41356_new_n5330_; 
wire _abc_41356_new_n5331_; 
wire _abc_41356_new_n5332_; 
wire _abc_41356_new_n5333_; 
wire _abc_41356_new_n5334_; 
wire _abc_41356_new_n5335_; 
wire _abc_41356_new_n5336_; 
wire _abc_41356_new_n5338_; 
wire _abc_41356_new_n5339_; 
wire _abc_41356_new_n533_; 
wire _abc_41356_new_n5340_; 
wire _abc_41356_new_n5341_; 
wire _abc_41356_new_n5342_; 
wire _abc_41356_new_n5343_; 
wire _abc_41356_new_n5344_; 
wire _abc_41356_new_n5345_; 
wire _abc_41356_new_n5346_; 
wire _abc_41356_new_n5347_; 
wire _abc_41356_new_n5348_; 
wire _abc_41356_new_n5349_; 
wire _abc_41356_new_n534_; 
wire _abc_41356_new_n5350_; 
wire _abc_41356_new_n5351_; 
wire _abc_41356_new_n5352_; 
wire _abc_41356_new_n5353_; 
wire _abc_41356_new_n5354_; 
wire _abc_41356_new_n5355_; 
wire _abc_41356_new_n5356_; 
wire _abc_41356_new_n5357_; 
wire _abc_41356_new_n5358_; 
wire _abc_41356_new_n5359_; 
wire _abc_41356_new_n535_; 
wire _abc_41356_new_n5360_; 
wire _abc_41356_new_n5361_; 
wire _abc_41356_new_n5362_; 
wire _abc_41356_new_n5363_; 
wire _abc_41356_new_n5364_; 
wire _abc_41356_new_n5365_; 
wire _abc_41356_new_n5366_; 
wire _abc_41356_new_n5367_; 
wire _abc_41356_new_n5368_; 
wire _abc_41356_new_n5369_; 
wire _abc_41356_new_n536_; 
wire _abc_41356_new_n5370_; 
wire _abc_41356_new_n5371_; 
wire _abc_41356_new_n5372_; 
wire _abc_41356_new_n5373_; 
wire _abc_41356_new_n5375_; 
wire _abc_41356_new_n5376_; 
wire _abc_41356_new_n5377_; 
wire _abc_41356_new_n5378_; 
wire _abc_41356_new_n5379_; 
wire _abc_41356_new_n537_; 
wire _abc_41356_new_n5380_; 
wire _abc_41356_new_n5381_; 
wire _abc_41356_new_n5382_; 
wire _abc_41356_new_n5383_; 
wire _abc_41356_new_n5384_; 
wire _abc_41356_new_n5385_; 
wire _abc_41356_new_n5386_; 
wire _abc_41356_new_n5387_; 
wire _abc_41356_new_n5388_; 
wire _abc_41356_new_n5389_; 
wire _abc_41356_new_n538_; 
wire _abc_41356_new_n5390_; 
wire _abc_41356_new_n5391_; 
wire _abc_41356_new_n5392_; 
wire _abc_41356_new_n5393_; 
wire _abc_41356_new_n5394_; 
wire _abc_41356_new_n5395_; 
wire _abc_41356_new_n5396_; 
wire _abc_41356_new_n5397_; 
wire _abc_41356_new_n5398_; 
wire _abc_41356_new_n5399_; 
wire _abc_41356_new_n539_; 
wire _abc_41356_new_n5400_; 
wire _abc_41356_new_n5401_; 
wire _abc_41356_new_n5402_; 
wire _abc_41356_new_n5403_; 
wire _abc_41356_new_n5404_; 
wire _abc_41356_new_n5405_; 
wire _abc_41356_new_n5406_; 
wire _abc_41356_new_n5407_; 
wire _abc_41356_new_n5408_; 
wire _abc_41356_new_n5409_; 
wire _abc_41356_new_n540_; 
wire _abc_41356_new_n5410_; 
wire _abc_41356_new_n5412_; 
wire _abc_41356_new_n5413_; 
wire _abc_41356_new_n5414_; 
wire _abc_41356_new_n5415_; 
wire _abc_41356_new_n5416_; 
wire _abc_41356_new_n5417_; 
wire _abc_41356_new_n5418_; 
wire _abc_41356_new_n5419_; 
wire _abc_41356_new_n541_; 
wire _abc_41356_new_n5421_; 
wire _abc_41356_new_n5422_; 
wire _abc_41356_new_n5423_; 
wire _abc_41356_new_n5424_; 
wire _abc_41356_new_n5426_; 
wire _abc_41356_new_n5427_; 
wire _abc_41356_new_n5428_; 
wire _abc_41356_new_n5429_; 
wire _abc_41356_new_n542_; 
wire _abc_41356_new_n5431_; 
wire _abc_41356_new_n5432_; 
wire _abc_41356_new_n5433_; 
wire _abc_41356_new_n5434_; 
wire _abc_41356_new_n5436_; 
wire _abc_41356_new_n5437_; 
wire _abc_41356_new_n5438_; 
wire _abc_41356_new_n5439_; 
wire _abc_41356_new_n543_; 
wire _abc_41356_new_n5441_; 
wire _abc_41356_new_n5442_; 
wire _abc_41356_new_n5443_; 
wire _abc_41356_new_n5444_; 
wire _abc_41356_new_n5446_; 
wire _abc_41356_new_n5447_; 
wire _abc_41356_new_n5448_; 
wire _abc_41356_new_n5449_; 
wire _abc_41356_new_n544_; 
wire _abc_41356_new_n5451_; 
wire _abc_41356_new_n5452_; 
wire _abc_41356_new_n5453_; 
wire _abc_41356_new_n5454_; 
wire _abc_41356_new_n5456_; 
wire _abc_41356_new_n5457_; 
wire _abc_41356_new_n5458_; 
wire _abc_41356_new_n5459_; 
wire _abc_41356_new_n545_; 
wire _abc_41356_new_n5460_; 
wire _abc_41356_new_n5461_; 
wire _abc_41356_new_n5462_; 
wire _abc_41356_new_n5463_; 
wire _abc_41356_new_n5464_; 
wire _abc_41356_new_n5465_; 
wire _abc_41356_new_n5466_; 
wire _abc_41356_new_n5467_; 
wire _abc_41356_new_n5468_; 
wire _abc_41356_new_n5469_; 
wire _abc_41356_new_n546_; 
wire _abc_41356_new_n5470_; 
wire _abc_41356_new_n5471_; 
wire _abc_41356_new_n5473_; 
wire _abc_41356_new_n5474_; 
wire _abc_41356_new_n5475_; 
wire _abc_41356_new_n5476_; 
wire _abc_41356_new_n5477_; 
wire _abc_41356_new_n5478_; 
wire _abc_41356_new_n5479_; 
wire _abc_41356_new_n547_; 
wire _abc_41356_new_n5480_; 
wire _abc_41356_new_n5481_; 
wire _abc_41356_new_n5482_; 
wire _abc_41356_new_n5484_; 
wire _abc_41356_new_n5485_; 
wire _abc_41356_new_n5486_; 
wire _abc_41356_new_n5487_; 
wire _abc_41356_new_n5488_; 
wire _abc_41356_new_n5489_; 
wire _abc_41356_new_n548_; 
wire _abc_41356_new_n5490_; 
wire _abc_41356_new_n5491_; 
wire _abc_41356_new_n5492_; 
wire _abc_41356_new_n5493_; 
wire _abc_41356_new_n5495_; 
wire _abc_41356_new_n5496_; 
wire _abc_41356_new_n5497_; 
wire _abc_41356_new_n5498_; 
wire _abc_41356_new_n5499_; 
wire _abc_41356_new_n549_; 
wire _abc_41356_new_n5500_; 
wire _abc_41356_new_n5501_; 
wire _abc_41356_new_n5502_; 
wire _abc_41356_new_n5503_; 
wire _abc_41356_new_n5504_; 
wire _abc_41356_new_n5505_; 
wire _abc_41356_new_n5506_; 
wire _abc_41356_new_n5507_; 
wire _abc_41356_new_n5508_; 
wire _abc_41356_new_n5509_; 
wire _abc_41356_new_n550_; 
wire _abc_41356_new_n5510_; 
wire _abc_41356_new_n5511_; 
wire _abc_41356_new_n5512_; 
wire _abc_41356_new_n5513_; 
wire _abc_41356_new_n5514_; 
wire _abc_41356_new_n5515_; 
wire _abc_41356_new_n5516_; 
wire _abc_41356_new_n5517_; 
wire _abc_41356_new_n5518_; 
wire _abc_41356_new_n5519_; 
wire _abc_41356_new_n551_; 
wire _abc_41356_new_n5520_; 
wire _abc_41356_new_n5521_; 
wire _abc_41356_new_n5523_; 
wire _abc_41356_new_n5524_; 
wire _abc_41356_new_n5525_; 
wire _abc_41356_new_n5526_; 
wire _abc_41356_new_n5527_; 
wire _abc_41356_new_n5528_; 
wire _abc_41356_new_n5529_; 
wire _abc_41356_new_n552_; 
wire _abc_41356_new_n5530_; 
wire _abc_41356_new_n5531_; 
wire _abc_41356_new_n5532_; 
wire _abc_41356_new_n5533_; 
wire _abc_41356_new_n5534_; 
wire _abc_41356_new_n5535_; 
wire _abc_41356_new_n5536_; 
wire _abc_41356_new_n5537_; 
wire _abc_41356_new_n5538_; 
wire _abc_41356_new_n5539_; 
wire _abc_41356_new_n553_; 
wire _abc_41356_new_n5540_; 
wire _abc_41356_new_n5541_; 
wire _abc_41356_new_n5542_; 
wire _abc_41356_new_n5543_; 
wire _abc_41356_new_n5544_; 
wire _abc_41356_new_n5545_; 
wire _abc_41356_new_n5546_; 
wire _abc_41356_new_n5547_; 
wire _abc_41356_new_n5548_; 
wire _abc_41356_new_n5549_; 
wire _abc_41356_new_n554_; 
wire _abc_41356_new_n5550_; 
wire _abc_41356_new_n5551_; 
wire _abc_41356_new_n5552_; 
wire _abc_41356_new_n5553_; 
wire _abc_41356_new_n5554_; 
wire _abc_41356_new_n5555_; 
wire _abc_41356_new_n5557_; 
wire _abc_41356_new_n5558_; 
wire _abc_41356_new_n5559_; 
wire _abc_41356_new_n555_; 
wire _abc_41356_new_n5560_; 
wire _abc_41356_new_n5561_; 
wire _abc_41356_new_n5562_; 
wire _abc_41356_new_n5563_; 
wire _abc_41356_new_n5564_; 
wire _abc_41356_new_n5565_; 
wire _abc_41356_new_n5566_; 
wire _abc_41356_new_n5567_; 
wire _abc_41356_new_n5568_; 
wire _abc_41356_new_n5569_; 
wire _abc_41356_new_n556_; 
wire _abc_41356_new_n5570_; 
wire _abc_41356_new_n5571_; 
wire _abc_41356_new_n5572_; 
wire _abc_41356_new_n5573_; 
wire _abc_41356_new_n5574_; 
wire _abc_41356_new_n5575_; 
wire _abc_41356_new_n5576_; 
wire _abc_41356_new_n5577_; 
wire _abc_41356_new_n5578_; 
wire _abc_41356_new_n5579_; 
wire _abc_41356_new_n557_; 
wire _abc_41356_new_n5580_; 
wire _abc_41356_new_n5581_; 
wire _abc_41356_new_n5582_; 
wire _abc_41356_new_n5583_; 
wire _abc_41356_new_n5584_; 
wire _abc_41356_new_n5585_; 
wire _abc_41356_new_n5586_; 
wire _abc_41356_new_n5587_; 
wire _abc_41356_new_n5588_; 
wire _abc_41356_new_n5589_; 
wire _abc_41356_new_n558_; 
wire _abc_41356_new_n5590_; 
wire _abc_41356_new_n5591_; 
wire _abc_41356_new_n5592_; 
wire _abc_41356_new_n5593_; 
wire _abc_41356_new_n5594_; 
wire _abc_41356_new_n5595_; 
wire _abc_41356_new_n5596_; 
wire _abc_41356_new_n5597_; 
wire _abc_41356_new_n5598_; 
wire _abc_41356_new_n5599_; 
wire _abc_41356_new_n559_; 
wire _abc_41356_new_n5600_; 
wire _abc_41356_new_n5602_; 
wire _abc_41356_new_n5603_; 
wire _abc_41356_new_n5604_; 
wire _abc_41356_new_n5605_; 
wire _abc_41356_new_n5606_; 
wire _abc_41356_new_n5607_; 
wire _abc_41356_new_n5608_; 
wire _abc_41356_new_n5609_; 
wire _abc_41356_new_n560_; 
wire _abc_41356_new_n5610_; 
wire _abc_41356_new_n5611_; 
wire _abc_41356_new_n5612_; 
wire _abc_41356_new_n5613_; 
wire _abc_41356_new_n5614_; 
wire _abc_41356_new_n5615_; 
wire _abc_41356_new_n5616_; 
wire _abc_41356_new_n5617_; 
wire _abc_41356_new_n5618_; 
wire _abc_41356_new_n5619_; 
wire _abc_41356_new_n561_; 
wire _abc_41356_new_n5620_; 
wire _abc_41356_new_n5621_; 
wire _abc_41356_new_n5622_; 
wire _abc_41356_new_n5623_; 
wire _abc_41356_new_n5624_; 
wire _abc_41356_new_n5625_; 
wire _abc_41356_new_n5626_; 
wire _abc_41356_new_n5627_; 
wire _abc_41356_new_n5628_; 
wire _abc_41356_new_n5629_; 
wire _abc_41356_new_n562_; 
wire _abc_41356_new_n5630_; 
wire _abc_41356_new_n5631_; 
wire _abc_41356_new_n5632_; 
wire _abc_41356_new_n5633_; 
wire _abc_41356_new_n5634_; 
wire _abc_41356_new_n5635_; 
wire _abc_41356_new_n5636_; 
wire _abc_41356_new_n5637_; 
wire _abc_41356_new_n5638_; 
wire _abc_41356_new_n5639_; 
wire _abc_41356_new_n563_; 
wire _abc_41356_new_n5640_; 
wire _abc_41356_new_n5641_; 
wire _abc_41356_new_n5642_; 
wire _abc_41356_new_n5643_; 
wire _abc_41356_new_n5644_; 
wire _abc_41356_new_n5645_; 
wire _abc_41356_new_n5646_; 
wire _abc_41356_new_n5647_; 
wire _abc_41356_new_n5649_; 
wire _abc_41356_new_n564_; 
wire _abc_41356_new_n5650_; 
wire _abc_41356_new_n5651_; 
wire _abc_41356_new_n5652_; 
wire _abc_41356_new_n5653_; 
wire _abc_41356_new_n5654_; 
wire _abc_41356_new_n5655_; 
wire _abc_41356_new_n5656_; 
wire _abc_41356_new_n5657_; 
wire _abc_41356_new_n5658_; 
wire _abc_41356_new_n5659_; 
wire _abc_41356_new_n565_; 
wire _abc_41356_new_n5660_; 
wire _abc_41356_new_n5661_; 
wire _abc_41356_new_n5662_; 
wire _abc_41356_new_n5663_; 
wire _abc_41356_new_n5664_; 
wire _abc_41356_new_n5665_; 
wire _abc_41356_new_n5666_; 
wire _abc_41356_new_n5667_; 
wire _abc_41356_new_n5668_; 
wire _abc_41356_new_n5669_; 
wire _abc_41356_new_n566_; 
wire _abc_41356_new_n5670_; 
wire _abc_41356_new_n5671_; 
wire _abc_41356_new_n5672_; 
wire _abc_41356_new_n5673_; 
wire _abc_41356_new_n5674_; 
wire _abc_41356_new_n5675_; 
wire _abc_41356_new_n5676_; 
wire _abc_41356_new_n5677_; 
wire _abc_41356_new_n5678_; 
wire _abc_41356_new_n5679_; 
wire _abc_41356_new_n567_; 
wire _abc_41356_new_n5680_; 
wire _abc_41356_new_n5681_; 
wire _abc_41356_new_n5682_; 
wire _abc_41356_new_n5683_; 
wire _abc_41356_new_n5684_; 
wire _abc_41356_new_n5685_; 
wire _abc_41356_new_n5686_; 
wire _abc_41356_new_n5687_; 
wire _abc_41356_new_n5688_; 
wire _abc_41356_new_n5689_; 
wire _abc_41356_new_n568_; 
wire _abc_41356_new_n5690_; 
wire _abc_41356_new_n5691_; 
wire _abc_41356_new_n5693_; 
wire _abc_41356_new_n5694_; 
wire _abc_41356_new_n5695_; 
wire _abc_41356_new_n5696_; 
wire _abc_41356_new_n5697_; 
wire _abc_41356_new_n5698_; 
wire _abc_41356_new_n5699_; 
wire _abc_41356_new_n569_; 
wire _abc_41356_new_n5700_; 
wire _abc_41356_new_n5701_; 
wire _abc_41356_new_n5702_; 
wire _abc_41356_new_n5703_; 
wire _abc_41356_new_n5704_; 
wire _abc_41356_new_n5705_; 
wire _abc_41356_new_n5706_; 
wire _abc_41356_new_n5707_; 
wire _abc_41356_new_n5708_; 
wire _abc_41356_new_n5709_; 
wire _abc_41356_new_n570_; 
wire _abc_41356_new_n5710_; 
wire _abc_41356_new_n5711_; 
wire _abc_41356_new_n5712_; 
wire _abc_41356_new_n5713_; 
wire _abc_41356_new_n5714_; 
wire _abc_41356_new_n5715_; 
wire _abc_41356_new_n5716_; 
wire _abc_41356_new_n5717_; 
wire _abc_41356_new_n5718_; 
wire _abc_41356_new_n5719_; 
wire _abc_41356_new_n571_; 
wire _abc_41356_new_n5720_; 
wire _abc_41356_new_n5721_; 
wire _abc_41356_new_n5722_; 
wire _abc_41356_new_n5723_; 
wire _abc_41356_new_n5724_; 
wire _abc_41356_new_n5725_; 
wire _abc_41356_new_n5726_; 
wire _abc_41356_new_n5727_; 
wire _abc_41356_new_n5728_; 
wire _abc_41356_new_n5729_; 
wire _abc_41356_new_n572_; 
wire _abc_41356_new_n5730_; 
wire _abc_41356_new_n5731_; 
wire _abc_41356_new_n5732_; 
wire _abc_41356_new_n5733_; 
wire _abc_41356_new_n5734_; 
wire _abc_41356_new_n5735_; 
wire _abc_41356_new_n5736_; 
wire _abc_41356_new_n5737_; 
wire _abc_41356_new_n5738_; 
wire _abc_41356_new_n5739_; 
wire _abc_41356_new_n573_; 
wire _abc_41356_new_n5740_; 
wire _abc_41356_new_n5742_; 
wire _abc_41356_new_n5743_; 
wire _abc_41356_new_n5744_; 
wire _abc_41356_new_n5745_; 
wire _abc_41356_new_n5746_; 
wire _abc_41356_new_n5747_; 
wire _abc_41356_new_n5748_; 
wire _abc_41356_new_n5749_; 
wire _abc_41356_new_n574_; 
wire _abc_41356_new_n5750_; 
wire _abc_41356_new_n5751_; 
wire _abc_41356_new_n5752_; 
wire _abc_41356_new_n5753_; 
wire _abc_41356_new_n5754_; 
wire _abc_41356_new_n5755_; 
wire _abc_41356_new_n5756_; 
wire _abc_41356_new_n5757_; 
wire _abc_41356_new_n5758_; 
wire _abc_41356_new_n5759_; 
wire _abc_41356_new_n575_; 
wire _abc_41356_new_n5760_; 
wire _abc_41356_new_n5761_; 
wire _abc_41356_new_n5762_; 
wire _abc_41356_new_n5763_; 
wire _abc_41356_new_n5764_; 
wire _abc_41356_new_n5765_; 
wire _abc_41356_new_n5766_; 
wire _abc_41356_new_n5767_; 
wire _abc_41356_new_n5768_; 
wire _abc_41356_new_n5769_; 
wire _abc_41356_new_n576_; 
wire _abc_41356_new_n5770_; 
wire _abc_41356_new_n5771_; 
wire _abc_41356_new_n5772_; 
wire _abc_41356_new_n5773_; 
wire _abc_41356_new_n5774_; 
wire _abc_41356_new_n5775_; 
wire _abc_41356_new_n5776_; 
wire _abc_41356_new_n5777_; 
wire _abc_41356_new_n5778_; 
wire _abc_41356_new_n5779_; 
wire _abc_41356_new_n577_; 
wire _abc_41356_new_n5780_; 
wire _abc_41356_new_n5781_; 
wire _abc_41356_new_n5782_; 
wire _abc_41356_new_n5783_; 
wire _abc_41356_new_n5784_; 
wire _abc_41356_new_n5785_; 
wire _abc_41356_new_n5786_; 
wire _abc_41356_new_n5787_; 
wire _abc_41356_new_n5788_; 
wire _abc_41356_new_n578_; 
wire _abc_41356_new_n5790_; 
wire _abc_41356_new_n5791_; 
wire _abc_41356_new_n5792_; 
wire _abc_41356_new_n5793_; 
wire _abc_41356_new_n5794_; 
wire _abc_41356_new_n5795_; 
wire _abc_41356_new_n5796_; 
wire _abc_41356_new_n5797_; 
wire _abc_41356_new_n5798_; 
wire _abc_41356_new_n5799_; 
wire _abc_41356_new_n579_; 
wire _abc_41356_new_n5800_; 
wire _abc_41356_new_n5801_; 
wire _abc_41356_new_n5802_; 
wire _abc_41356_new_n5803_; 
wire _abc_41356_new_n5804_; 
wire _abc_41356_new_n5805_; 
wire _abc_41356_new_n5806_; 
wire _abc_41356_new_n5807_; 
wire _abc_41356_new_n5808_; 
wire _abc_41356_new_n5809_; 
wire _abc_41356_new_n580_; 
wire _abc_41356_new_n5810_; 
wire _abc_41356_new_n5811_; 
wire _abc_41356_new_n5812_; 
wire _abc_41356_new_n5813_; 
wire _abc_41356_new_n5814_; 
wire _abc_41356_new_n5815_; 
wire _abc_41356_new_n5816_; 
wire _abc_41356_new_n5817_; 
wire _abc_41356_new_n5818_; 
wire _abc_41356_new_n5819_; 
wire _abc_41356_new_n581_; 
wire _abc_41356_new_n5820_; 
wire _abc_41356_new_n5821_; 
wire _abc_41356_new_n5822_; 
wire _abc_41356_new_n5823_; 
wire _abc_41356_new_n5824_; 
wire _abc_41356_new_n5825_; 
wire _abc_41356_new_n5826_; 
wire _abc_41356_new_n5827_; 
wire _abc_41356_new_n5828_; 
wire _abc_41356_new_n5829_; 
wire _abc_41356_new_n582_; 
wire _abc_41356_new_n5830_; 
wire _abc_41356_new_n5831_; 
wire _abc_41356_new_n5832_; 
wire _abc_41356_new_n5833_; 
wire _abc_41356_new_n5834_; 
wire _abc_41356_new_n5835_; 
wire _abc_41356_new_n5836_; 
wire _abc_41356_new_n5838_; 
wire _abc_41356_new_n5839_; 
wire _abc_41356_new_n583_; 
wire _abc_41356_new_n5840_; 
wire _abc_41356_new_n5841_; 
wire _abc_41356_new_n5842_; 
wire _abc_41356_new_n5843_; 
wire _abc_41356_new_n5844_; 
wire _abc_41356_new_n5845_; 
wire _abc_41356_new_n5846_; 
wire _abc_41356_new_n5847_; 
wire _abc_41356_new_n5848_; 
wire _abc_41356_new_n5849_; 
wire _abc_41356_new_n584_; 
wire _abc_41356_new_n5850_; 
wire _abc_41356_new_n5851_; 
wire _abc_41356_new_n5852_; 
wire _abc_41356_new_n5853_; 
wire _abc_41356_new_n5854_; 
wire _abc_41356_new_n5855_; 
wire _abc_41356_new_n5856_; 
wire _abc_41356_new_n5857_; 
wire _abc_41356_new_n5858_; 
wire _abc_41356_new_n5859_; 
wire _abc_41356_new_n585_; 
wire _abc_41356_new_n5860_; 
wire _abc_41356_new_n5861_; 
wire _abc_41356_new_n5862_; 
wire _abc_41356_new_n5863_; 
wire _abc_41356_new_n5864_; 
wire _abc_41356_new_n5865_; 
wire _abc_41356_new_n5866_; 
wire _abc_41356_new_n5867_; 
wire _abc_41356_new_n5868_; 
wire _abc_41356_new_n5869_; 
wire _abc_41356_new_n586_; 
wire _abc_41356_new_n5870_; 
wire _abc_41356_new_n5871_; 
wire _abc_41356_new_n5873_; 
wire _abc_41356_new_n5874_; 
wire _abc_41356_new_n5875_; 
wire _abc_41356_new_n5876_; 
wire _abc_41356_new_n5877_; 
wire _abc_41356_new_n5878_; 
wire _abc_41356_new_n5879_; 
wire _abc_41356_new_n587_; 
wire _abc_41356_new_n5880_; 
wire _abc_41356_new_n5881_; 
wire _abc_41356_new_n5882_; 
wire _abc_41356_new_n5883_; 
wire _abc_41356_new_n5884_; 
wire _abc_41356_new_n5885_; 
wire _abc_41356_new_n5886_; 
wire _abc_41356_new_n5887_; 
wire _abc_41356_new_n5888_; 
wire _abc_41356_new_n5889_; 
wire _abc_41356_new_n588_; 
wire _abc_41356_new_n5890_; 
wire _abc_41356_new_n5891_; 
wire _abc_41356_new_n5892_; 
wire _abc_41356_new_n5893_; 
wire _abc_41356_new_n5894_; 
wire _abc_41356_new_n5895_; 
wire _abc_41356_new_n5896_; 
wire _abc_41356_new_n5897_; 
wire _abc_41356_new_n5898_; 
wire _abc_41356_new_n5899_; 
wire _abc_41356_new_n589_; 
wire _abc_41356_new_n5900_; 
wire _abc_41356_new_n5901_; 
wire _abc_41356_new_n5902_; 
wire _abc_41356_new_n5903_; 
wire _abc_41356_new_n5904_; 
wire _abc_41356_new_n5905_; 
wire _abc_41356_new_n5906_; 
wire _abc_41356_new_n5908_; 
wire _abc_41356_new_n5909_; 
wire _abc_41356_new_n590_; 
wire _abc_41356_new_n5910_; 
wire _abc_41356_new_n5911_; 
wire _abc_41356_new_n5912_; 
wire _abc_41356_new_n5913_; 
wire _abc_41356_new_n5914_; 
wire _abc_41356_new_n5915_; 
wire _abc_41356_new_n5916_; 
wire _abc_41356_new_n5917_; 
wire _abc_41356_new_n5918_; 
wire _abc_41356_new_n5919_; 
wire _abc_41356_new_n591_; 
wire _abc_41356_new_n5920_; 
wire _abc_41356_new_n5921_; 
wire _abc_41356_new_n5922_; 
wire _abc_41356_new_n5923_; 
wire _abc_41356_new_n5924_; 
wire _abc_41356_new_n5925_; 
wire _abc_41356_new_n5926_; 
wire _abc_41356_new_n5927_; 
wire _abc_41356_new_n5928_; 
wire _abc_41356_new_n5929_; 
wire _abc_41356_new_n592_; 
wire _abc_41356_new_n5930_; 
wire _abc_41356_new_n5931_; 
wire _abc_41356_new_n5932_; 
wire _abc_41356_new_n5933_; 
wire _abc_41356_new_n5934_; 
wire _abc_41356_new_n5935_; 
wire _abc_41356_new_n5936_; 
wire _abc_41356_new_n5937_; 
wire _abc_41356_new_n5938_; 
wire _abc_41356_new_n5939_; 
wire _abc_41356_new_n593_; 
wire _abc_41356_new_n5940_; 
wire _abc_41356_new_n5941_; 
wire _abc_41356_new_n5943_; 
wire _abc_41356_new_n5944_; 
wire _abc_41356_new_n5945_; 
wire _abc_41356_new_n5946_; 
wire _abc_41356_new_n5947_; 
wire _abc_41356_new_n5948_; 
wire _abc_41356_new_n5949_; 
wire _abc_41356_new_n594_; 
wire _abc_41356_new_n5950_; 
wire _abc_41356_new_n5951_; 
wire _abc_41356_new_n5952_; 
wire _abc_41356_new_n5953_; 
wire _abc_41356_new_n5954_; 
wire _abc_41356_new_n5955_; 
wire _abc_41356_new_n5956_; 
wire _abc_41356_new_n5957_; 
wire _abc_41356_new_n5958_; 
wire _abc_41356_new_n5959_; 
wire _abc_41356_new_n595_; 
wire _abc_41356_new_n5960_; 
wire _abc_41356_new_n5961_; 
wire _abc_41356_new_n5962_; 
wire _abc_41356_new_n5963_; 
wire _abc_41356_new_n5964_; 
wire _abc_41356_new_n5965_; 
wire _abc_41356_new_n5966_; 
wire _abc_41356_new_n5967_; 
wire _abc_41356_new_n5968_; 
wire _abc_41356_new_n5969_; 
wire _abc_41356_new_n596_; 
wire _abc_41356_new_n5970_; 
wire _abc_41356_new_n5971_; 
wire _abc_41356_new_n5972_; 
wire _abc_41356_new_n5973_; 
wire _abc_41356_new_n5974_; 
wire _abc_41356_new_n5975_; 
wire _abc_41356_new_n5976_; 
wire _abc_41356_new_n5977_; 
wire _abc_41356_new_n5978_; 
wire _abc_41356_new_n5979_; 
wire _abc_41356_new_n597_; 
wire _abc_41356_new_n5981_; 
wire _abc_41356_new_n5982_; 
wire _abc_41356_new_n5983_; 
wire _abc_41356_new_n5984_; 
wire _abc_41356_new_n5985_; 
wire _abc_41356_new_n5986_; 
wire _abc_41356_new_n5987_; 
wire _abc_41356_new_n5988_; 
wire _abc_41356_new_n5989_; 
wire _abc_41356_new_n598_; 
wire _abc_41356_new_n5990_; 
wire _abc_41356_new_n5991_; 
wire _abc_41356_new_n5992_; 
wire _abc_41356_new_n5993_; 
wire _abc_41356_new_n5994_; 
wire _abc_41356_new_n5995_; 
wire _abc_41356_new_n5996_; 
wire _abc_41356_new_n5997_; 
wire _abc_41356_new_n5998_; 
wire _abc_41356_new_n5999_; 
wire _abc_41356_new_n599_; 
wire _abc_41356_new_n6000_; 
wire _abc_41356_new_n6001_; 
wire _abc_41356_new_n6002_; 
wire _abc_41356_new_n6003_; 
wire _abc_41356_new_n6004_; 
wire _abc_41356_new_n6005_; 
wire _abc_41356_new_n6006_; 
wire _abc_41356_new_n6007_; 
wire _abc_41356_new_n6008_; 
wire _abc_41356_new_n6009_; 
wire _abc_41356_new_n600_; 
wire _abc_41356_new_n6010_; 
wire _abc_41356_new_n6011_; 
wire _abc_41356_new_n6012_; 
wire _abc_41356_new_n6013_; 
wire _abc_41356_new_n6014_; 
wire _abc_41356_new_n6015_; 
wire _abc_41356_new_n6016_; 
wire _abc_41356_new_n6017_; 
wire _abc_41356_new_n6018_; 
wire _abc_41356_new_n6019_; 
wire _abc_41356_new_n601_; 
wire _abc_41356_new_n6021_; 
wire _abc_41356_new_n6022_; 
wire _abc_41356_new_n6023_; 
wire _abc_41356_new_n6024_; 
wire _abc_41356_new_n6025_; 
wire _abc_41356_new_n6026_; 
wire _abc_41356_new_n6027_; 
wire _abc_41356_new_n6028_; 
wire _abc_41356_new_n6029_; 
wire _abc_41356_new_n602_; 
wire _abc_41356_new_n6030_; 
wire _abc_41356_new_n6031_; 
wire _abc_41356_new_n6032_; 
wire _abc_41356_new_n6033_; 
wire _abc_41356_new_n6034_; 
wire _abc_41356_new_n6035_; 
wire _abc_41356_new_n6036_; 
wire _abc_41356_new_n6037_; 
wire _abc_41356_new_n6038_; 
wire _abc_41356_new_n6039_; 
wire _abc_41356_new_n603_; 
wire _abc_41356_new_n6040_; 
wire _abc_41356_new_n6041_; 
wire _abc_41356_new_n6042_; 
wire _abc_41356_new_n6043_; 
wire _abc_41356_new_n6044_; 
wire _abc_41356_new_n6045_; 
wire _abc_41356_new_n6046_; 
wire _abc_41356_new_n6047_; 
wire _abc_41356_new_n6048_; 
wire _abc_41356_new_n6049_; 
wire _abc_41356_new_n604_; 
wire _abc_41356_new_n6050_; 
wire _abc_41356_new_n6051_; 
wire _abc_41356_new_n6052_; 
wire _abc_41356_new_n6053_; 
wire _abc_41356_new_n6054_; 
wire _abc_41356_new_n6055_; 
wire _abc_41356_new_n6056_; 
wire _abc_41356_new_n6057_; 
wire _abc_41356_new_n6059_; 
wire _abc_41356_new_n605_; 
wire _abc_41356_new_n6060_; 
wire _abc_41356_new_n6061_; 
wire _abc_41356_new_n6062_; 
wire _abc_41356_new_n6063_; 
wire _abc_41356_new_n6064_; 
wire _abc_41356_new_n6065_; 
wire _abc_41356_new_n6066_; 
wire _abc_41356_new_n6067_; 
wire _abc_41356_new_n6068_; 
wire _abc_41356_new_n6069_; 
wire _abc_41356_new_n606_; 
wire _abc_41356_new_n6070_; 
wire _abc_41356_new_n6071_; 
wire _abc_41356_new_n6072_; 
wire _abc_41356_new_n6073_; 
wire _abc_41356_new_n6074_; 
wire _abc_41356_new_n6075_; 
wire _abc_41356_new_n6076_; 
wire _abc_41356_new_n6077_; 
wire _abc_41356_new_n6078_; 
wire _abc_41356_new_n6079_; 
wire _abc_41356_new_n607_; 
wire _abc_41356_new_n6080_; 
wire _abc_41356_new_n6081_; 
wire _abc_41356_new_n6082_; 
wire _abc_41356_new_n6083_; 
wire _abc_41356_new_n6084_; 
wire _abc_41356_new_n6085_; 
wire _abc_41356_new_n6086_; 
wire _abc_41356_new_n6087_; 
wire _abc_41356_new_n6088_; 
wire _abc_41356_new_n6089_; 
wire _abc_41356_new_n608_; 
wire _abc_41356_new_n6090_; 
wire _abc_41356_new_n6091_; 
wire _abc_41356_new_n6092_; 
wire _abc_41356_new_n6093_; 
wire _abc_41356_new_n6095_; 
wire _abc_41356_new_n6096_; 
wire _abc_41356_new_n6097_; 
wire _abc_41356_new_n6098_; 
wire _abc_41356_new_n6099_; 
wire _abc_41356_new_n609_; 
wire _abc_41356_new_n6100_; 
wire _abc_41356_new_n6101_; 
wire _abc_41356_new_n6102_; 
wire _abc_41356_new_n6103_; 
wire _abc_41356_new_n6104_; 
wire _abc_41356_new_n6105_; 
wire _abc_41356_new_n6106_; 
wire _abc_41356_new_n6107_; 
wire _abc_41356_new_n6108_; 
wire _abc_41356_new_n6109_; 
wire _abc_41356_new_n610_; 
wire _abc_41356_new_n6110_; 
wire _abc_41356_new_n6111_; 
wire _abc_41356_new_n6112_; 
wire _abc_41356_new_n6113_; 
wire _abc_41356_new_n6114_; 
wire _abc_41356_new_n6115_; 
wire _abc_41356_new_n6116_; 
wire _abc_41356_new_n6117_; 
wire _abc_41356_new_n6118_; 
wire _abc_41356_new_n6119_; 
wire _abc_41356_new_n611_; 
wire _abc_41356_new_n6120_; 
wire _abc_41356_new_n6121_; 
wire _abc_41356_new_n6122_; 
wire _abc_41356_new_n6123_; 
wire _abc_41356_new_n6124_; 
wire _abc_41356_new_n6125_; 
wire _abc_41356_new_n6126_; 
wire _abc_41356_new_n6127_; 
wire _abc_41356_new_n6128_; 
wire _abc_41356_new_n6129_; 
wire _abc_41356_new_n612_; 
wire _abc_41356_new_n6130_; 
wire _abc_41356_new_n6131_; 
wire _abc_41356_new_n6132_; 
wire _abc_41356_new_n6134_; 
wire _abc_41356_new_n6135_; 
wire _abc_41356_new_n6136_; 
wire _abc_41356_new_n6137_; 
wire _abc_41356_new_n6138_; 
wire _abc_41356_new_n6139_; 
wire _abc_41356_new_n613_; 
wire _abc_41356_new_n6140_; 
wire _abc_41356_new_n6141_; 
wire _abc_41356_new_n6142_; 
wire _abc_41356_new_n6143_; 
wire _abc_41356_new_n6144_; 
wire _abc_41356_new_n6145_; 
wire _abc_41356_new_n6146_; 
wire _abc_41356_new_n6147_; 
wire _abc_41356_new_n6148_; 
wire _abc_41356_new_n6149_; 
wire _abc_41356_new_n614_; 
wire _abc_41356_new_n6150_; 
wire _abc_41356_new_n6151_; 
wire _abc_41356_new_n6152_; 
wire _abc_41356_new_n6153_; 
wire _abc_41356_new_n6154_; 
wire _abc_41356_new_n6155_; 
wire _abc_41356_new_n6156_; 
wire _abc_41356_new_n6157_; 
wire _abc_41356_new_n6158_; 
wire _abc_41356_new_n6159_; 
wire _abc_41356_new_n615_; 
wire _abc_41356_new_n6160_; 
wire _abc_41356_new_n6161_; 
wire _abc_41356_new_n6162_; 
wire _abc_41356_new_n6163_; 
wire _abc_41356_new_n6164_; 
wire _abc_41356_new_n6165_; 
wire _abc_41356_new_n6166_; 
wire _abc_41356_new_n6167_; 
wire _abc_41356_new_n6168_; 
wire _abc_41356_new_n6169_; 
wire _abc_41356_new_n616_; 
wire _abc_41356_new_n6170_; 
wire _abc_41356_new_n6171_; 
wire _abc_41356_new_n6173_; 
wire _abc_41356_new_n6174_; 
wire _abc_41356_new_n6175_; 
wire _abc_41356_new_n6176_; 
wire _abc_41356_new_n6177_; 
wire _abc_41356_new_n6178_; 
wire _abc_41356_new_n6179_; 
wire _abc_41356_new_n617_; 
wire _abc_41356_new_n6180_; 
wire _abc_41356_new_n6181_; 
wire _abc_41356_new_n6182_; 
wire _abc_41356_new_n6183_; 
wire _abc_41356_new_n6184_; 
wire _abc_41356_new_n6185_; 
wire _abc_41356_new_n6186_; 
wire _abc_41356_new_n6187_; 
wire _abc_41356_new_n6188_; 
wire _abc_41356_new_n6189_; 
wire _abc_41356_new_n618_; 
wire _abc_41356_new_n6190_; 
wire _abc_41356_new_n6191_; 
wire _abc_41356_new_n6192_; 
wire _abc_41356_new_n6193_; 
wire _abc_41356_new_n6194_; 
wire _abc_41356_new_n6195_; 
wire _abc_41356_new_n6196_; 
wire _abc_41356_new_n6197_; 
wire _abc_41356_new_n6198_; 
wire _abc_41356_new_n6199_; 
wire _abc_41356_new_n619_; 
wire _abc_41356_new_n6200_; 
wire _abc_41356_new_n6201_; 
wire _abc_41356_new_n6202_; 
wire _abc_41356_new_n6203_; 
wire _abc_41356_new_n6204_; 
wire _abc_41356_new_n6205_; 
wire _abc_41356_new_n6206_; 
wire _abc_41356_new_n6207_; 
wire _abc_41356_new_n6208_; 
wire _abc_41356_new_n6209_; 
wire _abc_41356_new_n620_; 
wire _abc_41356_new_n6210_; 
wire _abc_41356_new_n6212_; 
wire _abc_41356_new_n6213_; 
wire _abc_41356_new_n6214_; 
wire _abc_41356_new_n6215_; 
wire _abc_41356_new_n6216_; 
wire _abc_41356_new_n6217_; 
wire _abc_41356_new_n6218_; 
wire _abc_41356_new_n6219_; 
wire _abc_41356_new_n621_; 
wire _abc_41356_new_n6220_; 
wire _abc_41356_new_n6221_; 
wire _abc_41356_new_n6222_; 
wire _abc_41356_new_n6223_; 
wire _abc_41356_new_n6224_; 
wire _abc_41356_new_n6225_; 
wire _abc_41356_new_n6226_; 
wire _abc_41356_new_n6227_; 
wire _abc_41356_new_n6228_; 
wire _abc_41356_new_n6229_; 
wire _abc_41356_new_n622_; 
wire _abc_41356_new_n6230_; 
wire _abc_41356_new_n6231_; 
wire _abc_41356_new_n6232_; 
wire _abc_41356_new_n6233_; 
wire _abc_41356_new_n6234_; 
wire _abc_41356_new_n6235_; 
wire _abc_41356_new_n6236_; 
wire _abc_41356_new_n6237_; 
wire _abc_41356_new_n6238_; 
wire _abc_41356_new_n6239_; 
wire _abc_41356_new_n623_; 
wire _abc_41356_new_n6240_; 
wire _abc_41356_new_n6241_; 
wire _abc_41356_new_n6242_; 
wire _abc_41356_new_n6243_; 
wire _abc_41356_new_n6244_; 
wire _abc_41356_new_n6245_; 
wire _abc_41356_new_n6247_; 
wire _abc_41356_new_n6248_; 
wire _abc_41356_new_n6249_; 
wire _abc_41356_new_n624_; 
wire _abc_41356_new_n6250_; 
wire _abc_41356_new_n6251_; 
wire _abc_41356_new_n6252_; 
wire _abc_41356_new_n6253_; 
wire _abc_41356_new_n6254_; 
wire _abc_41356_new_n6255_; 
wire _abc_41356_new_n6256_; 
wire _abc_41356_new_n6257_; 
wire _abc_41356_new_n6258_; 
wire _abc_41356_new_n6259_; 
wire _abc_41356_new_n625_; 
wire _abc_41356_new_n6260_; 
wire _abc_41356_new_n6261_; 
wire _abc_41356_new_n6262_; 
wire _abc_41356_new_n6263_; 
wire _abc_41356_new_n6264_; 
wire _abc_41356_new_n6265_; 
wire _abc_41356_new_n6266_; 
wire _abc_41356_new_n6267_; 
wire _abc_41356_new_n6268_; 
wire _abc_41356_new_n6269_; 
wire _abc_41356_new_n626_; 
wire _abc_41356_new_n6270_; 
wire _abc_41356_new_n6271_; 
wire _abc_41356_new_n6272_; 
wire _abc_41356_new_n6273_; 
wire _abc_41356_new_n6274_; 
wire _abc_41356_new_n6275_; 
wire _abc_41356_new_n6276_; 
wire _abc_41356_new_n6277_; 
wire _abc_41356_new_n6278_; 
wire _abc_41356_new_n6279_; 
wire _abc_41356_new_n627_; 
wire _abc_41356_new_n6280_; 
wire _abc_41356_new_n6281_; 
wire _abc_41356_new_n6282_; 
wire _abc_41356_new_n6283_; 
wire _abc_41356_new_n6284_; 
wire _abc_41356_new_n6285_; 
wire _abc_41356_new_n6287_; 
wire _abc_41356_new_n6288_; 
wire _abc_41356_new_n6289_; 
wire _abc_41356_new_n628_; 
wire _abc_41356_new_n6290_; 
wire _abc_41356_new_n6291_; 
wire _abc_41356_new_n6292_; 
wire _abc_41356_new_n6293_; 
wire _abc_41356_new_n6294_; 
wire _abc_41356_new_n6295_; 
wire _abc_41356_new_n6296_; 
wire _abc_41356_new_n6297_; 
wire _abc_41356_new_n6298_; 
wire _abc_41356_new_n6299_; 
wire _abc_41356_new_n629_; 
wire _abc_41356_new_n6300_; 
wire _abc_41356_new_n6301_; 
wire _abc_41356_new_n6302_; 
wire _abc_41356_new_n6303_; 
wire _abc_41356_new_n6304_; 
wire _abc_41356_new_n6305_; 
wire _abc_41356_new_n6306_; 
wire _abc_41356_new_n6307_; 
wire _abc_41356_new_n6308_; 
wire _abc_41356_new_n6309_; 
wire _abc_41356_new_n630_; 
wire _abc_41356_new_n6310_; 
wire _abc_41356_new_n6311_; 
wire _abc_41356_new_n6312_; 
wire _abc_41356_new_n6313_; 
wire _abc_41356_new_n6314_; 
wire _abc_41356_new_n6315_; 
wire _abc_41356_new_n6316_; 
wire _abc_41356_new_n6317_; 
wire _abc_41356_new_n6318_; 
wire _abc_41356_new_n6319_; 
wire _abc_41356_new_n631_; 
wire _abc_41356_new_n6320_; 
wire _abc_41356_new_n6322_; 
wire _abc_41356_new_n6323_; 
wire _abc_41356_new_n6324_; 
wire _abc_41356_new_n6325_; 
wire _abc_41356_new_n6326_; 
wire _abc_41356_new_n6327_; 
wire _abc_41356_new_n6328_; 
wire _abc_41356_new_n6329_; 
wire _abc_41356_new_n632_; 
wire _abc_41356_new_n6330_; 
wire _abc_41356_new_n6331_; 
wire _abc_41356_new_n6332_; 
wire _abc_41356_new_n6333_; 
wire _abc_41356_new_n6334_; 
wire _abc_41356_new_n6335_; 
wire _abc_41356_new_n6336_; 
wire _abc_41356_new_n6337_; 
wire _abc_41356_new_n6338_; 
wire _abc_41356_new_n6339_; 
wire _abc_41356_new_n633_; 
wire _abc_41356_new_n6340_; 
wire _abc_41356_new_n6341_; 
wire _abc_41356_new_n6342_; 
wire _abc_41356_new_n6343_; 
wire _abc_41356_new_n6344_; 
wire _abc_41356_new_n6345_; 
wire _abc_41356_new_n6346_; 
wire _abc_41356_new_n6347_; 
wire _abc_41356_new_n6348_; 
wire _abc_41356_new_n6349_; 
wire _abc_41356_new_n634_; 
wire _abc_41356_new_n6350_; 
wire _abc_41356_new_n6351_; 
wire _abc_41356_new_n6352_; 
wire _abc_41356_new_n6353_; 
wire _abc_41356_new_n6354_; 
wire _abc_41356_new_n6355_; 
wire _abc_41356_new_n6356_; 
wire _abc_41356_new_n6357_; 
wire _abc_41356_new_n6358_; 
wire _abc_41356_new_n6359_; 
wire _abc_41356_new_n635_; 
wire _abc_41356_new_n6361_; 
wire _abc_41356_new_n6362_; 
wire _abc_41356_new_n6363_; 
wire _abc_41356_new_n6364_; 
wire _abc_41356_new_n6365_; 
wire _abc_41356_new_n6366_; 
wire _abc_41356_new_n6367_; 
wire _abc_41356_new_n6368_; 
wire _abc_41356_new_n6369_; 
wire _abc_41356_new_n636_; 
wire _abc_41356_new_n6370_; 
wire _abc_41356_new_n6371_; 
wire _abc_41356_new_n6372_; 
wire _abc_41356_new_n6373_; 
wire _abc_41356_new_n6374_; 
wire _abc_41356_new_n6375_; 
wire _abc_41356_new_n6376_; 
wire _abc_41356_new_n6377_; 
wire _abc_41356_new_n6378_; 
wire _abc_41356_new_n6379_; 
wire _abc_41356_new_n637_; 
wire _abc_41356_new_n6380_; 
wire _abc_41356_new_n6381_; 
wire _abc_41356_new_n6382_; 
wire _abc_41356_new_n6383_; 
wire _abc_41356_new_n6384_; 
wire _abc_41356_new_n6385_; 
wire _abc_41356_new_n6386_; 
wire _abc_41356_new_n6387_; 
wire _abc_41356_new_n6388_; 
wire _abc_41356_new_n6389_; 
wire _abc_41356_new_n638_; 
wire _abc_41356_new_n6390_; 
wire _abc_41356_new_n6391_; 
wire _abc_41356_new_n6392_; 
wire _abc_41356_new_n6393_; 
wire _abc_41356_new_n6394_; 
wire _abc_41356_new_n6395_; 
wire _abc_41356_new_n6396_; 
wire _abc_41356_new_n6397_; 
wire _abc_41356_new_n6398_; 
wire _abc_41356_new_n639_; 
wire _abc_41356_new_n6400_; 
wire _abc_41356_new_n6401_; 
wire _abc_41356_new_n6402_; 
wire _abc_41356_new_n6403_; 
wire _abc_41356_new_n6404_; 
wire _abc_41356_new_n6405_; 
wire _abc_41356_new_n6406_; 
wire _abc_41356_new_n6407_; 
wire _abc_41356_new_n6408_; 
wire _abc_41356_new_n6409_; 
wire _abc_41356_new_n640_; 
wire _abc_41356_new_n6410_; 
wire _abc_41356_new_n6411_; 
wire _abc_41356_new_n6412_; 
wire _abc_41356_new_n6413_; 
wire _abc_41356_new_n6414_; 
wire _abc_41356_new_n6415_; 
wire _abc_41356_new_n6416_; 
wire _abc_41356_new_n6417_; 
wire _abc_41356_new_n6418_; 
wire _abc_41356_new_n6419_; 
wire _abc_41356_new_n641_; 
wire _abc_41356_new_n6420_; 
wire _abc_41356_new_n6421_; 
wire _abc_41356_new_n6422_; 
wire _abc_41356_new_n6423_; 
wire _abc_41356_new_n6424_; 
wire _abc_41356_new_n6425_; 
wire _abc_41356_new_n6426_; 
wire _abc_41356_new_n6427_; 
wire _abc_41356_new_n6428_; 
wire _abc_41356_new_n6429_; 
wire _abc_41356_new_n642_; 
wire _abc_41356_new_n6430_; 
wire _abc_41356_new_n6431_; 
wire _abc_41356_new_n6432_; 
wire _abc_41356_new_n6433_; 
wire _abc_41356_new_n6434_; 
wire _abc_41356_new_n6436_; 
wire _abc_41356_new_n6437_; 
wire _abc_41356_new_n6438_; 
wire _abc_41356_new_n6439_; 
wire _abc_41356_new_n643_; 
wire _abc_41356_new_n6441_; 
wire _abc_41356_new_n6442_; 
wire _abc_41356_new_n6444_; 
wire _abc_41356_new_n6445_; 
wire _abc_41356_new_n6447_; 
wire _abc_41356_new_n6448_; 
wire _abc_41356_new_n644_; 
wire _abc_41356_new_n6450_; 
wire _abc_41356_new_n6451_; 
wire _abc_41356_new_n6453_; 
wire _abc_41356_new_n6454_; 
wire _abc_41356_new_n6456_; 
wire _abc_41356_new_n6457_; 
wire _abc_41356_new_n6459_; 
wire _abc_41356_new_n645_; 
wire _abc_41356_new_n6460_; 
wire _abc_41356_new_n6462_; 
wire _abc_41356_new_n6463_; 
wire _abc_41356_new_n6464_; 
wire _abc_41356_new_n6465_; 
wire _abc_41356_new_n6466_; 
wire _abc_41356_new_n6467_; 
wire _abc_41356_new_n6468_; 
wire _abc_41356_new_n6469_; 
wire _abc_41356_new_n646_; 
wire _abc_41356_new_n6470_; 
wire _abc_41356_new_n6471_; 
wire _abc_41356_new_n6472_; 
wire _abc_41356_new_n6473_; 
wire _abc_41356_new_n6474_; 
wire _abc_41356_new_n6475_; 
wire _abc_41356_new_n6476_; 
wire _abc_41356_new_n6477_; 
wire _abc_41356_new_n6478_; 
wire _abc_41356_new_n6479_; 
wire _abc_41356_new_n647_; 
wire _abc_41356_new_n6480_; 
wire _abc_41356_new_n6481_; 
wire _abc_41356_new_n6482_; 
wire _abc_41356_new_n6483_; 
wire _abc_41356_new_n6484_; 
wire _abc_41356_new_n6485_; 
wire _abc_41356_new_n6486_; 
wire _abc_41356_new_n6487_; 
wire _abc_41356_new_n6488_; 
wire _abc_41356_new_n6489_; 
wire _abc_41356_new_n648_; 
wire _abc_41356_new_n6490_; 
wire _abc_41356_new_n6491_; 
wire _abc_41356_new_n6492_; 
wire _abc_41356_new_n6493_; 
wire _abc_41356_new_n6494_; 
wire _abc_41356_new_n6495_; 
wire _abc_41356_new_n6496_; 
wire _abc_41356_new_n6497_; 
wire _abc_41356_new_n6498_; 
wire _abc_41356_new_n6499_; 
wire _abc_41356_new_n649_; 
wire _abc_41356_new_n6500_; 
wire _abc_41356_new_n6501_; 
wire _abc_41356_new_n6502_; 
wire _abc_41356_new_n6503_; 
wire _abc_41356_new_n6504_; 
wire _abc_41356_new_n6505_; 
wire _abc_41356_new_n6506_; 
wire _abc_41356_new_n6507_; 
wire _abc_41356_new_n6508_; 
wire _abc_41356_new_n6509_; 
wire _abc_41356_new_n650_; 
wire _abc_41356_new_n6510_; 
wire _abc_41356_new_n6511_; 
wire _abc_41356_new_n6513_; 
wire _abc_41356_new_n6514_; 
wire _abc_41356_new_n6515_; 
wire _abc_41356_new_n6516_; 
wire _abc_41356_new_n6517_; 
wire _abc_41356_new_n6518_; 
wire _abc_41356_new_n6519_; 
wire _abc_41356_new_n651_; 
wire _abc_41356_new_n6520_; 
wire _abc_41356_new_n6521_; 
wire _abc_41356_new_n6522_; 
wire _abc_41356_new_n6523_; 
wire _abc_41356_new_n6524_; 
wire _abc_41356_new_n6525_; 
wire _abc_41356_new_n6526_; 
wire _abc_41356_new_n6527_; 
wire _abc_41356_new_n6528_; 
wire _abc_41356_new_n6529_; 
wire _abc_41356_new_n652_; 
wire _abc_41356_new_n6530_; 
wire _abc_41356_new_n6531_; 
wire _abc_41356_new_n6532_; 
wire _abc_41356_new_n6533_; 
wire _abc_41356_new_n6534_; 
wire _abc_41356_new_n6535_; 
wire _abc_41356_new_n6536_; 
wire _abc_41356_new_n6537_; 
wire _abc_41356_new_n6538_; 
wire _abc_41356_new_n6539_; 
wire _abc_41356_new_n653_; 
wire _abc_41356_new_n6540_; 
wire _abc_41356_new_n6541_; 
wire _abc_41356_new_n6542_; 
wire _abc_41356_new_n6543_; 
wire _abc_41356_new_n6544_; 
wire _abc_41356_new_n6545_; 
wire _abc_41356_new_n6546_; 
wire _abc_41356_new_n6547_; 
wire _abc_41356_new_n6548_; 
wire _abc_41356_new_n6549_; 
wire _abc_41356_new_n654_; 
wire _abc_41356_new_n6550_; 
wire _abc_41356_new_n6551_; 
wire _abc_41356_new_n6552_; 
wire _abc_41356_new_n6553_; 
wire _abc_41356_new_n6554_; 
wire _abc_41356_new_n6555_; 
wire _abc_41356_new_n6556_; 
wire _abc_41356_new_n6557_; 
wire _abc_41356_new_n6558_; 
wire _abc_41356_new_n6559_; 
wire _abc_41356_new_n655_; 
wire _abc_41356_new_n6560_; 
wire _abc_41356_new_n6561_; 
wire _abc_41356_new_n6562_; 
wire _abc_41356_new_n6563_; 
wire _abc_41356_new_n6564_; 
wire _abc_41356_new_n6565_; 
wire _abc_41356_new_n6567_; 
wire _abc_41356_new_n6568_; 
wire _abc_41356_new_n6569_; 
wire _abc_41356_new_n656_; 
wire _abc_41356_new_n6570_; 
wire _abc_41356_new_n6571_; 
wire _abc_41356_new_n6572_; 
wire _abc_41356_new_n6573_; 
wire _abc_41356_new_n6574_; 
wire _abc_41356_new_n6575_; 
wire _abc_41356_new_n6576_; 
wire _abc_41356_new_n6577_; 
wire _abc_41356_new_n6578_; 
wire _abc_41356_new_n6579_; 
wire _abc_41356_new_n657_; 
wire _abc_41356_new_n6580_; 
wire _abc_41356_new_n6581_; 
wire _abc_41356_new_n6582_; 
wire _abc_41356_new_n6583_; 
wire _abc_41356_new_n6584_; 
wire _abc_41356_new_n6585_; 
wire _abc_41356_new_n6586_; 
wire _abc_41356_new_n6587_; 
wire _abc_41356_new_n6588_; 
wire _abc_41356_new_n6589_; 
wire _abc_41356_new_n658_; 
wire _abc_41356_new_n6590_; 
wire _abc_41356_new_n6591_; 
wire _abc_41356_new_n6592_; 
wire _abc_41356_new_n6593_; 
wire _abc_41356_new_n6594_; 
wire _abc_41356_new_n6595_; 
wire _abc_41356_new_n6596_; 
wire _abc_41356_new_n6598_; 
wire _abc_41356_new_n6599_; 
wire _abc_41356_new_n659_; 
wire _abc_41356_new_n6600_; 
wire _abc_41356_new_n6601_; 
wire _abc_41356_new_n6602_; 
wire _abc_41356_new_n6603_; 
wire _abc_41356_new_n6604_; 
wire _abc_41356_new_n6605_; 
wire _abc_41356_new_n6606_; 
wire _abc_41356_new_n6607_; 
wire _abc_41356_new_n6608_; 
wire _abc_41356_new_n6609_; 
wire _abc_41356_new_n660_; 
wire _abc_41356_new_n6610_; 
wire _abc_41356_new_n6611_; 
wire _abc_41356_new_n6612_; 
wire _abc_41356_new_n6613_; 
wire _abc_41356_new_n6614_; 
wire _abc_41356_new_n6615_; 
wire _abc_41356_new_n6616_; 
wire _abc_41356_new_n6617_; 
wire _abc_41356_new_n6618_; 
wire _abc_41356_new_n6619_; 
wire _abc_41356_new_n661_; 
wire _abc_41356_new_n6620_; 
wire _abc_41356_new_n6621_; 
wire _abc_41356_new_n6622_; 
wire _abc_41356_new_n6623_; 
wire _abc_41356_new_n6624_; 
wire _abc_41356_new_n6625_; 
wire _abc_41356_new_n6626_; 
wire _abc_41356_new_n6627_; 
wire _abc_41356_new_n6628_; 
wire _abc_41356_new_n6629_; 
wire _abc_41356_new_n662_; 
wire _abc_41356_new_n6630_; 
wire _abc_41356_new_n6631_; 
wire _abc_41356_new_n6632_; 
wire _abc_41356_new_n6633_; 
wire _abc_41356_new_n6634_; 
wire _abc_41356_new_n6635_; 
wire _abc_41356_new_n6636_; 
wire _abc_41356_new_n6637_; 
wire _abc_41356_new_n6639_; 
wire _abc_41356_new_n663_; 
wire _abc_41356_new_n6640_; 
wire _abc_41356_new_n6641_; 
wire _abc_41356_new_n6642_; 
wire _abc_41356_new_n6643_; 
wire _abc_41356_new_n6644_; 
wire _abc_41356_new_n6645_; 
wire _abc_41356_new_n6646_; 
wire _abc_41356_new_n6647_; 
wire _abc_41356_new_n6648_; 
wire _abc_41356_new_n6649_; 
wire _abc_41356_new_n664_; 
wire _abc_41356_new_n6650_; 
wire _abc_41356_new_n6651_; 
wire _abc_41356_new_n6652_; 
wire _abc_41356_new_n6653_; 
wire _abc_41356_new_n6654_; 
wire _abc_41356_new_n6655_; 
wire _abc_41356_new_n6656_; 
wire _abc_41356_new_n6657_; 
wire _abc_41356_new_n6658_; 
wire _abc_41356_new_n6659_; 
wire _abc_41356_new_n665_; 
wire _abc_41356_new_n6660_; 
wire _abc_41356_new_n6661_; 
wire _abc_41356_new_n6662_; 
wire _abc_41356_new_n6663_; 
wire _abc_41356_new_n6664_; 
wire _abc_41356_new_n6665_; 
wire _abc_41356_new_n6666_; 
wire _abc_41356_new_n6667_; 
wire _abc_41356_new_n6668_; 
wire _abc_41356_new_n6669_; 
wire _abc_41356_new_n666_; 
wire _abc_41356_new_n6670_; 
wire _abc_41356_new_n6671_; 
wire _abc_41356_new_n6673_; 
wire _abc_41356_new_n6674_; 
wire _abc_41356_new_n6675_; 
wire _abc_41356_new_n6676_; 
wire _abc_41356_new_n6677_; 
wire _abc_41356_new_n6678_; 
wire _abc_41356_new_n6679_; 
wire _abc_41356_new_n667_; 
wire _abc_41356_new_n6680_; 
wire _abc_41356_new_n6681_; 
wire _abc_41356_new_n6682_; 
wire _abc_41356_new_n6683_; 
wire _abc_41356_new_n6684_; 
wire _abc_41356_new_n6685_; 
wire _abc_41356_new_n6686_; 
wire _abc_41356_new_n6687_; 
wire _abc_41356_new_n6688_; 
wire _abc_41356_new_n6689_; 
wire _abc_41356_new_n668_; 
wire _abc_41356_new_n6690_; 
wire _abc_41356_new_n6691_; 
wire _abc_41356_new_n6692_; 
wire _abc_41356_new_n6693_; 
wire _abc_41356_new_n6694_; 
wire _abc_41356_new_n6695_; 
wire _abc_41356_new_n6696_; 
wire _abc_41356_new_n6697_; 
wire _abc_41356_new_n6698_; 
wire _abc_41356_new_n6699_; 
wire _abc_41356_new_n669_; 
wire _abc_41356_new_n6700_; 
wire _abc_41356_new_n6701_; 
wire _abc_41356_new_n6702_; 
wire _abc_41356_new_n6703_; 
wire _abc_41356_new_n6704_; 
wire _abc_41356_new_n6705_; 
wire _abc_41356_new_n6706_; 
wire _abc_41356_new_n6707_; 
wire _abc_41356_new_n6708_; 
wire _abc_41356_new_n6709_; 
wire _abc_41356_new_n670_; 
wire _abc_41356_new_n6711_; 
wire _abc_41356_new_n6712_; 
wire _abc_41356_new_n6713_; 
wire _abc_41356_new_n6714_; 
wire _abc_41356_new_n6715_; 
wire _abc_41356_new_n6716_; 
wire _abc_41356_new_n6717_; 
wire _abc_41356_new_n6718_; 
wire _abc_41356_new_n6719_; 
wire _abc_41356_new_n671_; 
wire _abc_41356_new_n6720_; 
wire _abc_41356_new_n6721_; 
wire _abc_41356_new_n6722_; 
wire _abc_41356_new_n6723_; 
wire _abc_41356_new_n6724_; 
wire _abc_41356_new_n6725_; 
wire _abc_41356_new_n6726_; 
wire _abc_41356_new_n6727_; 
wire _abc_41356_new_n6728_; 
wire _abc_41356_new_n6729_; 
wire _abc_41356_new_n672_; 
wire _abc_41356_new_n6730_; 
wire _abc_41356_new_n6731_; 
wire _abc_41356_new_n6732_; 
wire _abc_41356_new_n6733_; 
wire _abc_41356_new_n6734_; 
wire _abc_41356_new_n6735_; 
wire _abc_41356_new_n6736_; 
wire _abc_41356_new_n6737_; 
wire _abc_41356_new_n6738_; 
wire _abc_41356_new_n6739_; 
wire _abc_41356_new_n673_; 
wire _abc_41356_new_n6740_; 
wire _abc_41356_new_n6741_; 
wire _abc_41356_new_n6742_; 
wire _abc_41356_new_n6743_; 
wire _abc_41356_new_n6744_; 
wire _abc_41356_new_n6745_; 
wire _abc_41356_new_n6746_; 
wire _abc_41356_new_n6748_; 
wire _abc_41356_new_n6749_; 
wire _abc_41356_new_n674_; 
wire _abc_41356_new_n6750_; 
wire _abc_41356_new_n6751_; 
wire _abc_41356_new_n6752_; 
wire _abc_41356_new_n6753_; 
wire _abc_41356_new_n6754_; 
wire _abc_41356_new_n6755_; 
wire _abc_41356_new_n6756_; 
wire _abc_41356_new_n6757_; 
wire _abc_41356_new_n6758_; 
wire _abc_41356_new_n6759_; 
wire _abc_41356_new_n675_; 
wire _abc_41356_new_n6760_; 
wire _abc_41356_new_n6761_; 
wire _abc_41356_new_n6762_; 
wire _abc_41356_new_n6763_; 
wire _abc_41356_new_n6764_; 
wire _abc_41356_new_n6765_; 
wire _abc_41356_new_n6766_; 
wire _abc_41356_new_n6767_; 
wire _abc_41356_new_n6768_; 
wire _abc_41356_new_n6769_; 
wire _abc_41356_new_n676_; 
wire _abc_41356_new_n6770_; 
wire _abc_41356_new_n6771_; 
wire _abc_41356_new_n6772_; 
wire _abc_41356_new_n6773_; 
wire _abc_41356_new_n6774_; 
wire _abc_41356_new_n6775_; 
wire _abc_41356_new_n6776_; 
wire _abc_41356_new_n6777_; 
wire _abc_41356_new_n6778_; 
wire _abc_41356_new_n6779_; 
wire _abc_41356_new_n677_; 
wire _abc_41356_new_n6780_; 
wire _abc_41356_new_n6781_; 
wire _abc_41356_new_n6782_; 
wire _abc_41356_new_n6783_; 
wire _abc_41356_new_n6784_; 
wire _abc_41356_new_n6785_; 
wire _abc_41356_new_n6786_; 
wire _abc_41356_new_n6788_; 
wire _abc_41356_new_n6789_; 
wire _abc_41356_new_n678_; 
wire _abc_41356_new_n6790_; 
wire _abc_41356_new_n6791_; 
wire _abc_41356_new_n6792_; 
wire _abc_41356_new_n6793_; 
wire _abc_41356_new_n6794_; 
wire _abc_41356_new_n6795_; 
wire _abc_41356_new_n6796_; 
wire _abc_41356_new_n6797_; 
wire _abc_41356_new_n6798_; 
wire _abc_41356_new_n6799_; 
wire _abc_41356_new_n679_; 
wire _abc_41356_new_n6800_; 
wire _abc_41356_new_n6801_; 
wire _abc_41356_new_n6802_; 
wire _abc_41356_new_n6803_; 
wire _abc_41356_new_n6804_; 
wire _abc_41356_new_n6805_; 
wire _abc_41356_new_n6806_; 
wire _abc_41356_new_n6807_; 
wire _abc_41356_new_n6808_; 
wire _abc_41356_new_n6809_; 
wire _abc_41356_new_n680_; 
wire _abc_41356_new_n6810_; 
wire _abc_41356_new_n6811_; 
wire _abc_41356_new_n6812_; 
wire _abc_41356_new_n6813_; 
wire _abc_41356_new_n6814_; 
wire _abc_41356_new_n6815_; 
wire _abc_41356_new_n6816_; 
wire _abc_41356_new_n6817_; 
wire _abc_41356_new_n6818_; 
wire _abc_41356_new_n6819_; 
wire _abc_41356_new_n681_; 
wire _abc_41356_new_n6820_; 
wire _abc_41356_new_n6822_; 
wire _abc_41356_new_n6823_; 
wire _abc_41356_new_n6824_; 
wire _abc_41356_new_n6825_; 
wire _abc_41356_new_n6826_; 
wire _abc_41356_new_n6827_; 
wire _abc_41356_new_n6828_; 
wire _abc_41356_new_n6829_; 
wire _abc_41356_new_n682_; 
wire _abc_41356_new_n6830_; 
wire _abc_41356_new_n6831_; 
wire _abc_41356_new_n6832_; 
wire _abc_41356_new_n6833_; 
wire _abc_41356_new_n6834_; 
wire _abc_41356_new_n6835_; 
wire _abc_41356_new_n6836_; 
wire _abc_41356_new_n6837_; 
wire _abc_41356_new_n6838_; 
wire _abc_41356_new_n6839_; 
wire _abc_41356_new_n683_; 
wire _abc_41356_new_n6840_; 
wire _abc_41356_new_n6841_; 
wire _abc_41356_new_n6842_; 
wire _abc_41356_new_n6843_; 
wire _abc_41356_new_n6844_; 
wire _abc_41356_new_n6845_; 
wire _abc_41356_new_n6846_; 
wire _abc_41356_new_n6847_; 
wire _abc_41356_new_n6848_; 
wire _abc_41356_new_n6849_; 
wire _abc_41356_new_n684_; 
wire _abc_41356_new_n6850_; 
wire _abc_41356_new_n6851_; 
wire _abc_41356_new_n6852_; 
wire _abc_41356_new_n6853_; 
wire _abc_41356_new_n6854_; 
wire _abc_41356_new_n6855_; 
wire _abc_41356_new_n6856_; 
wire _abc_41356_new_n6857_; 
wire _abc_41356_new_n6858_; 
wire _abc_41356_new_n685_; 
wire _abc_41356_new_n6860_; 
wire _abc_41356_new_n6861_; 
wire _abc_41356_new_n6862_; 
wire _abc_41356_new_n6863_; 
wire _abc_41356_new_n6864_; 
wire _abc_41356_new_n6865_; 
wire _abc_41356_new_n6866_; 
wire _abc_41356_new_n6867_; 
wire _abc_41356_new_n6868_; 
wire _abc_41356_new_n6869_; 
wire _abc_41356_new_n686_; 
wire _abc_41356_new_n6870_; 
wire _abc_41356_new_n6871_; 
wire _abc_41356_new_n6872_; 
wire _abc_41356_new_n6873_; 
wire _abc_41356_new_n6874_; 
wire _abc_41356_new_n6875_; 
wire _abc_41356_new_n6876_; 
wire _abc_41356_new_n6877_; 
wire _abc_41356_new_n6878_; 
wire _abc_41356_new_n6879_; 
wire _abc_41356_new_n687_; 
wire _abc_41356_new_n6880_; 
wire _abc_41356_new_n6881_; 
wire _abc_41356_new_n6882_; 
wire _abc_41356_new_n6883_; 
wire _abc_41356_new_n6884_; 
wire _abc_41356_new_n6885_; 
wire _abc_41356_new_n6886_; 
wire _abc_41356_new_n6887_; 
wire _abc_41356_new_n6888_; 
wire _abc_41356_new_n6889_; 
wire _abc_41356_new_n688_; 
wire _abc_41356_new_n6890_; 
wire _abc_41356_new_n6891_; 
wire _abc_41356_new_n6892_; 
wire _abc_41356_new_n6894_; 
wire _abc_41356_new_n6895_; 
wire _abc_41356_new_n6896_; 
wire _abc_41356_new_n6897_; 
wire _abc_41356_new_n6898_; 
wire _abc_41356_new_n6899_; 
wire _abc_41356_new_n689_; 
wire _abc_41356_new_n6900_; 
wire _abc_41356_new_n6901_; 
wire _abc_41356_new_n6902_; 
wire _abc_41356_new_n6903_; 
wire _abc_41356_new_n6904_; 
wire _abc_41356_new_n6905_; 
wire _abc_41356_new_n6906_; 
wire _abc_41356_new_n6907_; 
wire _abc_41356_new_n6908_; 
wire _abc_41356_new_n6909_; 
wire _abc_41356_new_n690_; 
wire _abc_41356_new_n6910_; 
wire _abc_41356_new_n6911_; 
wire _abc_41356_new_n6912_; 
wire _abc_41356_new_n6913_; 
wire _abc_41356_new_n6914_; 
wire _abc_41356_new_n6915_; 
wire _abc_41356_new_n6916_; 
wire _abc_41356_new_n6917_; 
wire _abc_41356_new_n6918_; 
wire _abc_41356_new_n6919_; 
wire _abc_41356_new_n691_; 
wire _abc_41356_new_n6920_; 
wire _abc_41356_new_n6921_; 
wire _abc_41356_new_n6922_; 
wire _abc_41356_new_n6923_; 
wire _abc_41356_new_n6924_; 
wire _abc_41356_new_n6925_; 
wire _abc_41356_new_n6926_; 
wire _abc_41356_new_n6927_; 
wire _abc_41356_new_n6928_; 
wire _abc_41356_new_n692_; 
wire _abc_41356_new_n6930_; 
wire _abc_41356_new_n6931_; 
wire _abc_41356_new_n6932_; 
wire _abc_41356_new_n6933_; 
wire _abc_41356_new_n6934_; 
wire _abc_41356_new_n6935_; 
wire _abc_41356_new_n6936_; 
wire _abc_41356_new_n6937_; 
wire _abc_41356_new_n6938_; 
wire _abc_41356_new_n6939_; 
wire _abc_41356_new_n693_; 
wire _abc_41356_new_n6940_; 
wire _abc_41356_new_n6941_; 
wire _abc_41356_new_n6942_; 
wire _abc_41356_new_n6943_; 
wire _abc_41356_new_n6944_; 
wire _abc_41356_new_n6945_; 
wire _abc_41356_new_n6946_; 
wire _abc_41356_new_n6947_; 
wire _abc_41356_new_n6948_; 
wire _abc_41356_new_n6949_; 
wire _abc_41356_new_n694_; 
wire _abc_41356_new_n6950_; 
wire _abc_41356_new_n6951_; 
wire _abc_41356_new_n6952_; 
wire _abc_41356_new_n6953_; 
wire _abc_41356_new_n6954_; 
wire _abc_41356_new_n6955_; 
wire _abc_41356_new_n6956_; 
wire _abc_41356_new_n6957_; 
wire _abc_41356_new_n6958_; 
wire _abc_41356_new_n6959_; 
wire _abc_41356_new_n695_; 
wire _abc_41356_new_n6960_; 
wire _abc_41356_new_n6961_; 
wire _abc_41356_new_n6963_; 
wire _abc_41356_new_n6964_; 
wire _abc_41356_new_n6965_; 
wire _abc_41356_new_n6966_; 
wire _abc_41356_new_n6967_; 
wire _abc_41356_new_n6968_; 
wire _abc_41356_new_n6969_; 
wire _abc_41356_new_n696_; 
wire _abc_41356_new_n6970_; 
wire _abc_41356_new_n6971_; 
wire _abc_41356_new_n6972_; 
wire _abc_41356_new_n6973_; 
wire _abc_41356_new_n6974_; 
wire _abc_41356_new_n6975_; 
wire _abc_41356_new_n6976_; 
wire _abc_41356_new_n6977_; 
wire _abc_41356_new_n6978_; 
wire _abc_41356_new_n6979_; 
wire _abc_41356_new_n697_; 
wire _abc_41356_new_n6980_; 
wire _abc_41356_new_n6981_; 
wire _abc_41356_new_n6982_; 
wire _abc_41356_new_n6983_; 
wire _abc_41356_new_n6984_; 
wire _abc_41356_new_n6985_; 
wire _abc_41356_new_n6986_; 
wire _abc_41356_new_n6987_; 
wire _abc_41356_new_n6988_; 
wire _abc_41356_new_n6989_; 
wire _abc_41356_new_n698_; 
wire _abc_41356_new_n6990_; 
wire _abc_41356_new_n6991_; 
wire _abc_41356_new_n6992_; 
wire _abc_41356_new_n6993_; 
wire _abc_41356_new_n6995_; 
wire _abc_41356_new_n6996_; 
wire _abc_41356_new_n6997_; 
wire _abc_41356_new_n6998_; 
wire _abc_41356_new_n6999_; 
wire _abc_41356_new_n699_; 
wire _abc_41356_new_n7000_; 
wire _abc_41356_new_n7001_; 
wire _abc_41356_new_n7002_; 
wire _abc_41356_new_n7003_; 
wire _abc_41356_new_n7004_; 
wire _abc_41356_new_n7005_; 
wire _abc_41356_new_n7006_; 
wire _abc_41356_new_n7007_; 
wire _abc_41356_new_n7008_; 
wire _abc_41356_new_n7009_; 
wire _abc_41356_new_n700_; 
wire _abc_41356_new_n7010_; 
wire _abc_41356_new_n7011_; 
wire _abc_41356_new_n7012_; 
wire _abc_41356_new_n7013_; 
wire _abc_41356_new_n7014_; 
wire _abc_41356_new_n7015_; 
wire _abc_41356_new_n7016_; 
wire _abc_41356_new_n7017_; 
wire _abc_41356_new_n7018_; 
wire _abc_41356_new_n7019_; 
wire _abc_41356_new_n701_; 
wire _abc_41356_new_n7020_; 
wire _abc_41356_new_n7021_; 
wire _abc_41356_new_n7022_; 
wire _abc_41356_new_n7023_; 
wire _abc_41356_new_n7024_; 
wire _abc_41356_new_n7026_; 
wire _abc_41356_new_n7027_; 
wire _abc_41356_new_n7028_; 
wire _abc_41356_new_n7029_; 
wire _abc_41356_new_n702_; 
wire _abc_41356_new_n7030_; 
wire _abc_41356_new_n7031_; 
wire _abc_41356_new_n7032_; 
wire _abc_41356_new_n7033_; 
wire _abc_41356_new_n7034_; 
wire _abc_41356_new_n7035_; 
wire _abc_41356_new_n7036_; 
wire _abc_41356_new_n7037_; 
wire _abc_41356_new_n7038_; 
wire _abc_41356_new_n7039_; 
wire _abc_41356_new_n703_; 
wire _abc_41356_new_n7040_; 
wire _abc_41356_new_n7041_; 
wire _abc_41356_new_n7042_; 
wire _abc_41356_new_n7043_; 
wire _abc_41356_new_n7044_; 
wire _abc_41356_new_n7045_; 
wire _abc_41356_new_n7046_; 
wire _abc_41356_new_n7047_; 
wire _abc_41356_new_n7048_; 
wire _abc_41356_new_n7049_; 
wire _abc_41356_new_n704_; 
wire _abc_41356_new_n7050_; 
wire _abc_41356_new_n7051_; 
wire _abc_41356_new_n7052_; 
wire _abc_41356_new_n7053_; 
wire _abc_41356_new_n7054_; 
wire _abc_41356_new_n7055_; 
wire _abc_41356_new_n7057_; 
wire _abc_41356_new_n7058_; 
wire _abc_41356_new_n7059_; 
wire _abc_41356_new_n705_; 
wire _abc_41356_new_n7060_; 
wire _abc_41356_new_n7061_; 
wire _abc_41356_new_n7062_; 
wire _abc_41356_new_n7064_; 
wire _abc_41356_new_n7065_; 
wire _abc_41356_new_n7066_; 
wire _abc_41356_new_n7067_; 
wire _abc_41356_new_n7068_; 
wire _abc_41356_new_n7069_; 
wire _abc_41356_new_n706_; 
wire _abc_41356_new_n7070_; 
wire _abc_41356_new_n7071_; 
wire _abc_41356_new_n7072_; 
wire _abc_41356_new_n7073_; 
wire _abc_41356_new_n7074_; 
wire _abc_41356_new_n7075_; 
wire _abc_41356_new_n7076_; 
wire _abc_41356_new_n7078_; 
wire _abc_41356_new_n7079_; 
wire _abc_41356_new_n707_; 
wire _abc_41356_new_n7080_; 
wire _abc_41356_new_n7081_; 
wire _abc_41356_new_n7082_; 
wire _abc_41356_new_n7083_; 
wire _abc_41356_new_n7084_; 
wire _abc_41356_new_n7085_; 
wire _abc_41356_new_n7086_; 
wire _abc_41356_new_n7087_; 
wire _abc_41356_new_n7088_; 
wire _abc_41356_new_n7089_; 
wire _abc_41356_new_n708_; 
wire _abc_41356_new_n7090_; 
wire _abc_41356_new_n7091_; 
wire _abc_41356_new_n7092_; 
wire _abc_41356_new_n7093_; 
wire _abc_41356_new_n7095_; 
wire _abc_41356_new_n7096_; 
wire _abc_41356_new_n7097_; 
wire _abc_41356_new_n7098_; 
wire _abc_41356_new_n7099_; 
wire _abc_41356_new_n709_; 
wire _abc_41356_new_n7100_; 
wire _abc_41356_new_n7101_; 
wire _abc_41356_new_n7102_; 
wire _abc_41356_new_n7103_; 
wire _abc_41356_new_n7105_; 
wire _abc_41356_new_n7106_; 
wire _abc_41356_new_n7107_; 
wire _abc_41356_new_n7108_; 
wire _abc_41356_new_n7109_; 
wire _abc_41356_new_n710_; 
wire _abc_41356_new_n7110_; 
wire _abc_41356_new_n7111_; 
wire _abc_41356_new_n7112_; 
wire _abc_41356_new_n7113_; 
wire _abc_41356_new_n7115_; 
wire _abc_41356_new_n7116_; 
wire _abc_41356_new_n7117_; 
wire _abc_41356_new_n7118_; 
wire _abc_41356_new_n7119_; 
wire _abc_41356_new_n711_; 
wire _abc_41356_new_n7120_; 
wire _abc_41356_new_n7121_; 
wire _abc_41356_new_n7122_; 
wire _abc_41356_new_n7123_; 
wire _abc_41356_new_n7125_; 
wire _abc_41356_new_n7126_; 
wire _abc_41356_new_n7127_; 
wire _abc_41356_new_n7128_; 
wire _abc_41356_new_n7129_; 
wire _abc_41356_new_n712_; 
wire _abc_41356_new_n7130_; 
wire _abc_41356_new_n7131_; 
wire _abc_41356_new_n7132_; 
wire _abc_41356_new_n7133_; 
wire _abc_41356_new_n7135_; 
wire _abc_41356_new_n7136_; 
wire _abc_41356_new_n7137_; 
wire _abc_41356_new_n7138_; 
wire _abc_41356_new_n7139_; 
wire _abc_41356_new_n713_; 
wire _abc_41356_new_n7140_; 
wire _abc_41356_new_n7141_; 
wire _abc_41356_new_n7142_; 
wire _abc_41356_new_n7143_; 
wire _abc_41356_new_n7145_; 
wire _abc_41356_new_n7146_; 
wire _abc_41356_new_n7147_; 
wire _abc_41356_new_n7148_; 
wire _abc_41356_new_n7149_; 
wire _abc_41356_new_n714_; 
wire _abc_41356_new_n7150_; 
wire _abc_41356_new_n7151_; 
wire _abc_41356_new_n7152_; 
wire _abc_41356_new_n7153_; 
wire _abc_41356_new_n7155_; 
wire _abc_41356_new_n7156_; 
wire _abc_41356_new_n7157_; 
wire _abc_41356_new_n7158_; 
wire _abc_41356_new_n7159_; 
wire _abc_41356_new_n715_; 
wire _abc_41356_new_n7160_; 
wire _abc_41356_new_n7161_; 
wire _abc_41356_new_n7162_; 
wire _abc_41356_new_n7163_; 
wire _abc_41356_new_n7165_; 
wire _abc_41356_new_n7166_; 
wire _abc_41356_new_n7167_; 
wire _abc_41356_new_n7168_; 
wire _abc_41356_new_n7169_; 
wire _abc_41356_new_n716_; 
wire _abc_41356_new_n7170_; 
wire _abc_41356_new_n7171_; 
wire _abc_41356_new_n7173_; 
wire _abc_41356_new_n7174_; 
wire _abc_41356_new_n7175_; 
wire _abc_41356_new_n7176_; 
wire _abc_41356_new_n7177_; 
wire _abc_41356_new_n7178_; 
wire _abc_41356_new_n7179_; 
wire _abc_41356_new_n717_; 
wire _abc_41356_new_n7180_; 
wire _abc_41356_new_n7182_; 
wire _abc_41356_new_n7183_; 
wire _abc_41356_new_n7184_; 
wire _abc_41356_new_n7185_; 
wire _abc_41356_new_n7186_; 
wire _abc_41356_new_n7187_; 
wire _abc_41356_new_n7188_; 
wire _abc_41356_new_n718_; 
wire _abc_41356_new_n7190_; 
wire _abc_41356_new_n7191_; 
wire _abc_41356_new_n7192_; 
wire _abc_41356_new_n7193_; 
wire _abc_41356_new_n7194_; 
wire _abc_41356_new_n7195_; 
wire _abc_41356_new_n7196_; 
wire _abc_41356_new_n7198_; 
wire _abc_41356_new_n7199_; 
wire _abc_41356_new_n719_; 
wire _abc_41356_new_n7200_; 
wire _abc_41356_new_n7201_; 
wire _abc_41356_new_n7202_; 
wire _abc_41356_new_n7203_; 
wire _abc_41356_new_n7204_; 
wire _abc_41356_new_n7206_; 
wire _abc_41356_new_n7207_; 
wire _abc_41356_new_n7208_; 
wire _abc_41356_new_n7209_; 
wire _abc_41356_new_n720_; 
wire _abc_41356_new_n7210_; 
wire _abc_41356_new_n7211_; 
wire _abc_41356_new_n7212_; 
wire _abc_41356_new_n7214_; 
wire _abc_41356_new_n7215_; 
wire _abc_41356_new_n7216_; 
wire _abc_41356_new_n7217_; 
wire _abc_41356_new_n7218_; 
wire _abc_41356_new_n7219_; 
wire _abc_41356_new_n721_; 
wire _abc_41356_new_n7221_; 
wire _abc_41356_new_n7222_; 
wire _abc_41356_new_n7223_; 
wire _abc_41356_new_n7224_; 
wire _abc_41356_new_n7225_; 
wire _abc_41356_new_n7226_; 
wire _abc_41356_new_n7228_; 
wire _abc_41356_new_n7229_; 
wire _abc_41356_new_n722_; 
wire _abc_41356_new_n7230_; 
wire _abc_41356_new_n7231_; 
wire _abc_41356_new_n7232_; 
wire _abc_41356_new_n7234_; 
wire _abc_41356_new_n7235_; 
wire _abc_41356_new_n7236_; 
wire _abc_41356_new_n7237_; 
wire _abc_41356_new_n7238_; 
wire _abc_41356_new_n7239_; 
wire _abc_41356_new_n723_; 
wire _abc_41356_new_n7240_; 
wire _abc_41356_new_n7241_; 
wire _abc_41356_new_n7243_; 
wire _abc_41356_new_n7244_; 
wire _abc_41356_new_n7245_; 
wire _abc_41356_new_n7246_; 
wire _abc_41356_new_n7247_; 
wire _abc_41356_new_n7248_; 
wire _abc_41356_new_n724_; 
wire _abc_41356_new_n7250_; 
wire _abc_41356_new_n7251_; 
wire _abc_41356_new_n7252_; 
wire _abc_41356_new_n7253_; 
wire _abc_41356_new_n7254_; 
wire _abc_41356_new_n7255_; 
wire _abc_41356_new_n7256_; 
wire _abc_41356_new_n7257_; 
wire _abc_41356_new_n7258_; 
wire _abc_41356_new_n7259_; 
wire _abc_41356_new_n725_; 
wire _abc_41356_new_n7260_; 
wire _abc_41356_new_n7261_; 
wire _abc_41356_new_n7262_; 
wire _abc_41356_new_n7263_; 
wire _abc_41356_new_n7264_; 
wire _abc_41356_new_n7265_; 
wire _abc_41356_new_n7266_; 
wire _abc_41356_new_n7267_; 
wire _abc_41356_new_n7268_; 
wire _abc_41356_new_n7269_; 
wire _abc_41356_new_n726_; 
wire _abc_41356_new_n7270_; 
wire _abc_41356_new_n7271_; 
wire _abc_41356_new_n7272_; 
wire _abc_41356_new_n7273_; 
wire _abc_41356_new_n7274_; 
wire _abc_41356_new_n7275_; 
wire _abc_41356_new_n7276_; 
wire _abc_41356_new_n7277_; 
wire _abc_41356_new_n7278_; 
wire _abc_41356_new_n7279_; 
wire _abc_41356_new_n727_; 
wire _abc_41356_new_n7280_; 
wire _abc_41356_new_n7281_; 
wire _abc_41356_new_n7282_; 
wire _abc_41356_new_n7283_; 
wire _abc_41356_new_n7284_; 
wire _abc_41356_new_n7285_; 
wire _abc_41356_new_n7286_; 
wire _abc_41356_new_n7287_; 
wire _abc_41356_new_n7288_; 
wire _abc_41356_new_n7289_; 
wire _abc_41356_new_n728_; 
wire _abc_41356_new_n7290_; 
wire _abc_41356_new_n7291_; 
wire _abc_41356_new_n7292_; 
wire _abc_41356_new_n7293_; 
wire _abc_41356_new_n7294_; 
wire _abc_41356_new_n7295_; 
wire _abc_41356_new_n7296_; 
wire _abc_41356_new_n7297_; 
wire _abc_41356_new_n7298_; 
wire _abc_41356_new_n7299_; 
wire _abc_41356_new_n729_; 
wire _abc_41356_new_n7300_; 
wire _abc_41356_new_n7301_; 
wire _abc_41356_new_n7302_; 
wire _abc_41356_new_n7303_; 
wire _abc_41356_new_n7304_; 
wire _abc_41356_new_n7305_; 
wire _abc_41356_new_n7306_; 
wire _abc_41356_new_n7307_; 
wire _abc_41356_new_n7308_; 
wire _abc_41356_new_n7309_; 
wire _abc_41356_new_n730_; 
wire _abc_41356_new_n7310_; 
wire _abc_41356_new_n7311_; 
wire _abc_41356_new_n7312_; 
wire _abc_41356_new_n7313_; 
wire _abc_41356_new_n7314_; 
wire _abc_41356_new_n7315_; 
wire _abc_41356_new_n7316_; 
wire _abc_41356_new_n7317_; 
wire _abc_41356_new_n7318_; 
wire _abc_41356_new_n7319_; 
wire _abc_41356_new_n731_; 
wire _abc_41356_new_n7320_; 
wire _abc_41356_new_n7321_; 
wire _abc_41356_new_n7322_; 
wire _abc_41356_new_n7323_; 
wire _abc_41356_new_n7324_; 
wire _abc_41356_new_n7325_; 
wire _abc_41356_new_n7326_; 
wire _abc_41356_new_n7327_; 
wire _abc_41356_new_n7328_; 
wire _abc_41356_new_n7329_; 
wire _abc_41356_new_n732_; 
wire _abc_41356_new_n7330_; 
wire _abc_41356_new_n7331_; 
wire _abc_41356_new_n7332_; 
wire _abc_41356_new_n7333_; 
wire _abc_41356_new_n7334_; 
wire _abc_41356_new_n7335_; 
wire _abc_41356_new_n7336_; 
wire _abc_41356_new_n7337_; 
wire _abc_41356_new_n7338_; 
wire _abc_41356_new_n7339_; 
wire _abc_41356_new_n733_; 
wire _abc_41356_new_n7340_; 
wire _abc_41356_new_n7341_; 
wire _abc_41356_new_n7342_; 
wire _abc_41356_new_n7343_; 
wire _abc_41356_new_n7344_; 
wire _abc_41356_new_n7345_; 
wire _abc_41356_new_n7346_; 
wire _abc_41356_new_n7347_; 
wire _abc_41356_new_n7348_; 
wire _abc_41356_new_n7349_; 
wire _abc_41356_new_n7350_; 
wire _abc_41356_new_n7351_; 
wire _abc_41356_new_n7352_; 
wire _abc_41356_new_n7353_; 
wire _abc_41356_new_n7354_; 
wire _abc_41356_new_n7355_; 
wire _abc_41356_new_n7356_; 
wire _abc_41356_new_n7357_; 
wire _abc_41356_new_n7358_; 
wire _abc_41356_new_n7359_; 
wire _abc_41356_new_n735_; 
wire _abc_41356_new_n7360_; 
wire _abc_41356_new_n7361_; 
wire _abc_41356_new_n7362_; 
wire _abc_41356_new_n7363_; 
wire _abc_41356_new_n7364_; 
wire _abc_41356_new_n7365_; 
wire _abc_41356_new_n7366_; 
wire _abc_41356_new_n7367_; 
wire _abc_41356_new_n7368_; 
wire _abc_41356_new_n7369_; 
wire _abc_41356_new_n736_; 
wire _abc_41356_new_n7370_; 
wire _abc_41356_new_n7371_; 
wire _abc_41356_new_n7372_; 
wire _abc_41356_new_n7373_; 
wire _abc_41356_new_n7374_; 
wire _abc_41356_new_n7375_; 
wire _abc_41356_new_n7376_; 
wire _abc_41356_new_n7377_; 
wire _abc_41356_new_n7378_; 
wire _abc_41356_new_n7379_; 
wire _abc_41356_new_n737_; 
wire _abc_41356_new_n7380_; 
wire _abc_41356_new_n7381_; 
wire _abc_41356_new_n7382_; 
wire _abc_41356_new_n7383_; 
wire _abc_41356_new_n7384_; 
wire _abc_41356_new_n7385_; 
wire _abc_41356_new_n7386_; 
wire _abc_41356_new_n7387_; 
wire _abc_41356_new_n7388_; 
wire _abc_41356_new_n7389_; 
wire _abc_41356_new_n738_; 
wire _abc_41356_new_n7390_; 
wire _abc_41356_new_n7391_; 
wire _abc_41356_new_n7392_; 
wire _abc_41356_new_n7393_; 
wire _abc_41356_new_n7394_; 
wire _abc_41356_new_n7395_; 
wire _abc_41356_new_n7396_; 
wire _abc_41356_new_n7397_; 
wire _abc_41356_new_n7398_; 
wire _abc_41356_new_n7399_; 
wire _abc_41356_new_n739_; 
wire _abc_41356_new_n7400_; 
wire _abc_41356_new_n7401_; 
wire _abc_41356_new_n7402_; 
wire _abc_41356_new_n7403_; 
wire _abc_41356_new_n7404_; 
wire _abc_41356_new_n7405_; 
wire _abc_41356_new_n7406_; 
wire _abc_41356_new_n7407_; 
wire _abc_41356_new_n7408_; 
wire _abc_41356_new_n7409_; 
wire _abc_41356_new_n740_; 
wire _abc_41356_new_n7410_; 
wire _abc_41356_new_n7411_; 
wire _abc_41356_new_n7412_; 
wire _abc_41356_new_n7413_; 
wire _abc_41356_new_n7414_; 
wire _abc_41356_new_n7415_; 
wire _abc_41356_new_n7416_; 
wire _abc_41356_new_n7417_; 
wire _abc_41356_new_n7418_; 
wire _abc_41356_new_n7419_; 
wire _abc_41356_new_n741_; 
wire _abc_41356_new_n7420_; 
wire _abc_41356_new_n7421_; 
wire _abc_41356_new_n7422_; 
wire _abc_41356_new_n7423_; 
wire _abc_41356_new_n7424_; 
wire _abc_41356_new_n7425_; 
wire _abc_41356_new_n7426_; 
wire _abc_41356_new_n7427_; 
wire _abc_41356_new_n7428_; 
wire _abc_41356_new_n7429_; 
wire _abc_41356_new_n742_; 
wire _abc_41356_new_n7430_; 
wire _abc_41356_new_n7431_; 
wire _abc_41356_new_n7432_; 
wire _abc_41356_new_n7433_; 
wire _abc_41356_new_n7434_; 
wire _abc_41356_new_n7435_; 
wire _abc_41356_new_n7436_; 
wire _abc_41356_new_n7437_; 
wire _abc_41356_new_n7438_; 
wire _abc_41356_new_n743_; 
wire _abc_41356_new_n7440_; 
wire _abc_41356_new_n7441_; 
wire _abc_41356_new_n7442_; 
wire _abc_41356_new_n7443_; 
wire _abc_41356_new_n7444_; 
wire _abc_41356_new_n7445_; 
wire _abc_41356_new_n7446_; 
wire _abc_41356_new_n7447_; 
wire _abc_41356_new_n7448_; 
wire _abc_41356_new_n7449_; 
wire _abc_41356_new_n744_; 
wire _abc_41356_new_n7450_; 
wire _abc_41356_new_n7451_; 
wire _abc_41356_new_n7452_; 
wire _abc_41356_new_n7453_; 
wire _abc_41356_new_n7454_; 
wire _abc_41356_new_n7455_; 
wire _abc_41356_new_n7456_; 
wire _abc_41356_new_n7457_; 
wire _abc_41356_new_n7458_; 
wire _abc_41356_new_n7459_; 
wire _abc_41356_new_n745_; 
wire _abc_41356_new_n7460_; 
wire _abc_41356_new_n7461_; 
wire _abc_41356_new_n7462_; 
wire _abc_41356_new_n7463_; 
wire _abc_41356_new_n7464_; 
wire _abc_41356_new_n7465_; 
wire _abc_41356_new_n7466_; 
wire _abc_41356_new_n7467_; 
wire _abc_41356_new_n7468_; 
wire _abc_41356_new_n7469_; 
wire _abc_41356_new_n746_; 
wire _abc_41356_new_n7470_; 
wire _abc_41356_new_n7471_; 
wire _abc_41356_new_n7472_; 
wire _abc_41356_new_n7473_; 
wire _abc_41356_new_n7474_; 
wire _abc_41356_new_n7475_; 
wire _abc_41356_new_n7477_; 
wire _abc_41356_new_n7478_; 
wire _abc_41356_new_n7479_; 
wire _abc_41356_new_n747_; 
wire _abc_41356_new_n7480_; 
wire _abc_41356_new_n7481_; 
wire _abc_41356_new_n7482_; 
wire _abc_41356_new_n7483_; 
wire _abc_41356_new_n7484_; 
wire _abc_41356_new_n7485_; 
wire _abc_41356_new_n7486_; 
wire _abc_41356_new_n7487_; 
wire _abc_41356_new_n7488_; 
wire _abc_41356_new_n7489_; 
wire _abc_41356_new_n748_; 
wire _abc_41356_new_n7490_; 
wire _abc_41356_new_n7491_; 
wire _abc_41356_new_n7492_; 
wire _abc_41356_new_n7493_; 
wire _abc_41356_new_n7494_; 
wire _abc_41356_new_n7495_; 
wire _abc_41356_new_n7496_; 
wire _abc_41356_new_n7497_; 
wire _abc_41356_new_n7498_; 
wire _abc_41356_new_n7499_; 
wire _abc_41356_new_n749_; 
wire _abc_41356_new_n7500_; 
wire _abc_41356_new_n7501_; 
wire _abc_41356_new_n7502_; 
wire _abc_41356_new_n7503_; 
wire _abc_41356_new_n7504_; 
wire _abc_41356_new_n7505_; 
wire _abc_41356_new_n7506_; 
wire _abc_41356_new_n7507_; 
wire _abc_41356_new_n7508_; 
wire _abc_41356_new_n750_; 
wire _abc_41356_new_n7510_; 
wire _abc_41356_new_n7511_; 
wire _abc_41356_new_n7512_; 
wire _abc_41356_new_n7513_; 
wire _abc_41356_new_n7514_; 
wire _abc_41356_new_n7515_; 
wire _abc_41356_new_n7516_; 
wire _abc_41356_new_n7517_; 
wire _abc_41356_new_n7518_; 
wire _abc_41356_new_n7519_; 
wire _abc_41356_new_n751_; 
wire _abc_41356_new_n7520_; 
wire _abc_41356_new_n7521_; 
wire _abc_41356_new_n7522_; 
wire _abc_41356_new_n7523_; 
wire _abc_41356_new_n7524_; 
wire _abc_41356_new_n7525_; 
wire _abc_41356_new_n7527_; 
wire _abc_41356_new_n7528_; 
wire _abc_41356_new_n7529_; 
wire _abc_41356_new_n752_; 
wire _abc_41356_new_n7530_; 
wire _abc_41356_new_n7531_; 
wire _abc_41356_new_n7532_; 
wire _abc_41356_new_n7533_; 
wire _abc_41356_new_n7534_; 
wire _abc_41356_new_n7535_; 
wire _abc_41356_new_n7536_; 
wire _abc_41356_new_n7537_; 
wire _abc_41356_new_n7538_; 
wire _abc_41356_new_n7539_; 
wire _abc_41356_new_n753_; 
wire _abc_41356_new_n7540_; 
wire _abc_41356_new_n7541_; 
wire _abc_41356_new_n7542_; 
wire _abc_41356_new_n7543_; 
wire _abc_41356_new_n7545_; 
wire _abc_41356_new_n7546_; 
wire _abc_41356_new_n7547_; 
wire _abc_41356_new_n7548_; 
wire _abc_41356_new_n7549_; 
wire _abc_41356_new_n754_; 
wire _abc_41356_new_n7550_; 
wire _abc_41356_new_n7551_; 
wire _abc_41356_new_n7552_; 
wire _abc_41356_new_n7554_; 
wire _abc_41356_new_n7555_; 
wire _abc_41356_new_n7556_; 
wire _abc_41356_new_n7557_; 
wire _abc_41356_new_n7558_; 
wire _abc_41356_new_n7559_; 
wire _abc_41356_new_n755_; 
wire _abc_41356_new_n7560_; 
wire _abc_41356_new_n7561_; 
wire _abc_41356_new_n7562_; 
wire _abc_41356_new_n756_; 
wire _abc_41356_new_n757_; 
wire _abc_41356_new_n758_; 
wire _abc_41356_new_n759_; 
wire _abc_41356_new_n760_; 
wire _abc_41356_new_n761_; 
wire _abc_41356_new_n762_; 
wire _abc_41356_new_n763_; 
wire _abc_41356_new_n764_; 
wire _abc_41356_new_n765_; 
wire _abc_41356_new_n766_; 
wire _abc_41356_new_n767_; 
wire _abc_41356_new_n768_; 
wire _abc_41356_new_n769_; 
wire _abc_41356_new_n770_; 
wire _abc_41356_new_n771_; 
wire _abc_41356_new_n772_; 
wire _abc_41356_new_n773_; 
wire _abc_41356_new_n774_; 
wire _abc_41356_new_n775_; 
wire _abc_41356_new_n776_; 
wire _abc_41356_new_n777_; 
wire _abc_41356_new_n778_; 
wire _abc_41356_new_n779_; 
wire _abc_41356_new_n780_; 
wire _abc_41356_new_n781_; 
wire _abc_41356_new_n782_; 
wire _abc_41356_new_n783_; 
wire _abc_41356_new_n784_; 
wire _abc_41356_new_n785_; 
wire _abc_41356_new_n786_; 
wire _abc_41356_new_n787_; 
wire _abc_41356_new_n788_; 
wire _abc_41356_new_n790_; 
wire _abc_41356_new_n791_; 
wire _abc_41356_new_n792_; 
wire _abc_41356_new_n793_; 
wire _abc_41356_new_n794_; 
wire _abc_41356_new_n795_; 
wire _abc_41356_new_n796_; 
wire _abc_41356_new_n797_; 
wire _abc_41356_new_n798_; 
wire _abc_41356_new_n799_; 
wire _abc_41356_new_n800_; 
wire _abc_41356_new_n801_; 
wire _abc_41356_new_n802_; 
wire _abc_41356_new_n803_; 
wire _abc_41356_new_n804_; 
wire _abc_41356_new_n805_; 
wire _abc_41356_new_n806_; 
wire _abc_41356_new_n807_; 
wire _abc_41356_new_n808_; 
wire _abc_41356_new_n809_; 
wire _abc_41356_new_n810_; 
wire _abc_41356_new_n811_; 
wire _abc_41356_new_n812_; 
wire _abc_41356_new_n813_; 
wire _abc_41356_new_n814_; 
wire _abc_41356_new_n815_; 
wire _abc_41356_new_n816_; 
wire _abc_41356_new_n817_; 
wire _abc_41356_new_n818_; 
wire _abc_41356_new_n819_; 
wire _abc_41356_new_n820_; 
wire _abc_41356_new_n821_; 
wire _abc_41356_new_n822_; 
wire _abc_41356_new_n823_; 
wire _abc_41356_new_n824_; 
wire _abc_41356_new_n825_; 
wire _abc_41356_new_n826_; 
wire _abc_41356_new_n827_; 
wire _abc_41356_new_n828_; 
wire _abc_41356_new_n829_; 
wire _abc_41356_new_n830_; 
wire _abc_41356_new_n831_; 
wire _abc_41356_new_n832_; 
wire _abc_41356_new_n833_; 
wire _abc_41356_new_n834_; 
wire _abc_41356_new_n835_; 
wire _abc_41356_new_n836_; 
wire _abc_41356_new_n837_; 
wire _abc_41356_new_n838_; 
wire _abc_41356_new_n839_; 
wire _abc_41356_new_n840_; 
wire _abc_41356_new_n841_; 
wire _abc_41356_new_n842_; 
wire _abc_41356_new_n843_; 
wire _abc_41356_new_n844_; 
wire _abc_41356_new_n845_; 
wire _abc_41356_new_n846_; 
wire _abc_41356_new_n847_; 
wire _abc_41356_new_n848_; 
wire _abc_41356_new_n849_; 
wire _abc_41356_new_n851_; 
wire _abc_41356_new_n852_; 
wire _abc_41356_new_n853_; 
wire _abc_41356_new_n854_; 
wire _abc_41356_new_n855_; 
wire _abc_41356_new_n856_; 
wire _abc_41356_new_n857_; 
wire _abc_41356_new_n858_; 
wire _abc_41356_new_n859_; 
wire _abc_41356_new_n860_; 
wire _abc_41356_new_n861_; 
wire _abc_41356_new_n862_; 
wire _abc_41356_new_n863_; 
wire _abc_41356_new_n864_; 
wire _abc_41356_new_n865_; 
wire _abc_41356_new_n866_; 
wire _abc_41356_new_n867_; 
wire _abc_41356_new_n868_; 
wire _abc_41356_new_n869_; 
wire _abc_41356_new_n870_; 
wire _abc_41356_new_n871_; 
wire _abc_41356_new_n872_; 
wire _abc_41356_new_n873_; 
wire _abc_41356_new_n874_; 
wire _abc_41356_new_n875_; 
wire _abc_41356_new_n876_; 
wire _abc_41356_new_n877_; 
wire _abc_41356_new_n878_; 
wire _abc_41356_new_n879_; 
wire _abc_41356_new_n880_; 
wire _abc_41356_new_n881_; 
wire _abc_41356_new_n882_; 
wire _abc_41356_new_n883_; 
wire _abc_41356_new_n884_; 
wire _abc_41356_new_n885_; 
wire _abc_41356_new_n886_; 
wire _abc_41356_new_n887_; 
wire _abc_41356_new_n888_; 
wire _abc_41356_new_n889_; 
wire _abc_41356_new_n890_; 
wire _abc_41356_new_n891_; 
wire _abc_41356_new_n892_; 
wire _abc_41356_new_n893_; 
wire _abc_41356_new_n894_; 
wire _abc_41356_new_n895_; 
wire _abc_41356_new_n896_; 
wire _abc_41356_new_n897_; 
wire _abc_41356_new_n898_; 
wire _abc_41356_new_n899_; 
wire _abc_41356_new_n900_; 
wire _abc_41356_new_n901_; 
wire _abc_41356_new_n902_; 
wire _abc_41356_new_n903_; 
wire _abc_41356_new_n904_; 
wire _abc_41356_new_n905_; 
wire _abc_41356_new_n906_; 
wire _abc_41356_new_n907_; 
wire _abc_41356_new_n908_; 
wire _abc_41356_new_n909_; 
wire _abc_41356_new_n910_; 
wire _abc_41356_new_n911_; 
wire _abc_41356_new_n912_; 
wire _abc_41356_new_n913_; 
wire _abc_41356_new_n914_; 
wire _abc_41356_new_n915_; 
wire _abc_41356_new_n916_; 
wire _abc_41356_new_n918_; 
wire _abc_41356_new_n919_; 
wire _abc_41356_new_n920_; 
wire _abc_41356_new_n921_; 
wire _abc_41356_new_n922_; 
wire _abc_41356_new_n923_; 
wire _abc_41356_new_n924_; 
wire _abc_41356_new_n925_; 
wire _abc_41356_new_n926_; 
wire _abc_41356_new_n927_; 
wire _abc_41356_new_n928_; 
wire _abc_41356_new_n929_; 
wire _abc_41356_new_n930_; 
wire _abc_41356_new_n931_; 
wire _abc_41356_new_n932_; 
wire _abc_41356_new_n933_; 
wire _abc_41356_new_n934_; 
wire _abc_41356_new_n935_; 
wire _abc_41356_new_n936_; 
wire _abc_41356_new_n937_; 
wire _abc_41356_new_n938_; 
wire _abc_41356_new_n939_; 
wire _abc_41356_new_n940_; 
wire _abc_41356_new_n941_; 
wire _abc_41356_new_n942_; 
wire _abc_41356_new_n943_; 
wire _abc_41356_new_n944_; 
wire _abc_41356_new_n945_; 
wire _abc_41356_new_n946_; 
wire _abc_41356_new_n947_; 
wire _abc_41356_new_n948_; 
wire _abc_41356_new_n949_; 
wire _abc_41356_new_n950_; 
wire _abc_41356_new_n951_; 
wire _abc_41356_new_n952_; 
wire _abc_41356_new_n953_; 
wire _abc_41356_new_n954_; 
wire _abc_41356_new_n955_; 
wire _abc_41356_new_n956_; 
wire _abc_41356_new_n957_; 
wire _abc_41356_new_n958_; 
wire _abc_41356_new_n959_; 
wire _abc_41356_new_n960_; 
wire _abc_41356_new_n961_; 
wire _abc_41356_new_n962_; 
wire _abc_41356_new_n963_; 
wire _abc_41356_new_n964_; 
wire _abc_41356_new_n965_; 
wire _abc_41356_new_n966_; 
wire _abc_41356_new_n967_; 
wire _abc_41356_new_n968_; 
wire _abc_41356_new_n969_; 
wire _abc_41356_new_n970_; 
wire _abc_41356_new_n971_; 
wire _abc_41356_new_n972_; 
wire _abc_41356_new_n973_; 
wire _abc_41356_new_n974_; 
wire _abc_41356_new_n975_; 
wire _abc_41356_new_n976_; 
wire _abc_41356_new_n977_; 
wire _abc_41356_new_n978_; 
wire _abc_41356_new_n979_; 
wire _abc_41356_new_n980_; 
wire _abc_41356_new_n981_; 
wire _abc_41356_new_n982_; 
wire _abc_41356_new_n983_; 
wire _abc_41356_new_n985_; 
wire _abc_41356_new_n986_; 
wire _abc_41356_new_n987_; 
wire _abc_41356_new_n988_; 
wire _abc_41356_new_n989_; 
wire _abc_41356_new_n990_; 
wire _abc_41356_new_n991_; 
wire _abc_41356_new_n992_; 
wire _abc_41356_new_n993_; 
wire _abc_41356_new_n994_; 
wire _abc_41356_new_n995_; 
wire _abc_41356_new_n996_; 
wire _abc_41356_new_n997_; 
wire _abc_41356_new_n998_; 
wire _abc_41356_new_n999_; 
output \addr[0] ;
output \addr[10] ;
output \addr[11] ;
output \addr[12] ;
output \addr[13] ;
output \addr[14] ;
output \addr[15] ;
output \addr[1] ;
output \addr[2] ;
output \addr[3] ;
output \addr[4] ;
output \addr[5] ;
output \addr[6] ;
output \addr[7] ;
output \addr[8] ;
output \addr[9] ;
wire alu__abc_40887_new_n100_; 
wire alu__abc_40887_new_n101_; 
wire alu__abc_40887_new_n102_; 
wire alu__abc_40887_new_n103_; 
wire alu__abc_40887_new_n104_; 
wire alu__abc_40887_new_n105_; 
wire alu__abc_40887_new_n106_; 
wire alu__abc_40887_new_n107_; 
wire alu__abc_40887_new_n108_; 
wire alu__abc_40887_new_n109_; 
wire alu__abc_40887_new_n110_; 
wire alu__abc_40887_new_n111_; 
wire alu__abc_40887_new_n112_; 
wire alu__abc_40887_new_n113_; 
wire alu__abc_40887_new_n114_; 
wire alu__abc_40887_new_n115_; 
wire alu__abc_40887_new_n116_; 
wire alu__abc_40887_new_n117_; 
wire alu__abc_40887_new_n118_; 
wire alu__abc_40887_new_n119_; 
wire alu__abc_40887_new_n120_; 
wire alu__abc_40887_new_n121_; 
wire alu__abc_40887_new_n122_; 
wire alu__abc_40887_new_n123_; 
wire alu__abc_40887_new_n124_; 
wire alu__abc_40887_new_n125_; 
wire alu__abc_40887_new_n126_; 
wire alu__abc_40887_new_n127_; 
wire alu__abc_40887_new_n128_; 
wire alu__abc_40887_new_n129_; 
wire alu__abc_40887_new_n130_; 
wire alu__abc_40887_new_n131_; 
wire alu__abc_40887_new_n132_; 
wire alu__abc_40887_new_n133_; 
wire alu__abc_40887_new_n134_; 
wire alu__abc_40887_new_n135_; 
wire alu__abc_40887_new_n136_; 
wire alu__abc_40887_new_n137_; 
wire alu__abc_40887_new_n138_; 
wire alu__abc_40887_new_n139_; 
wire alu__abc_40887_new_n140_; 
wire alu__abc_40887_new_n141_; 
wire alu__abc_40887_new_n142_; 
wire alu__abc_40887_new_n143_; 
wire alu__abc_40887_new_n144_; 
wire alu__abc_40887_new_n145_; 
wire alu__abc_40887_new_n146_; 
wire alu__abc_40887_new_n147_; 
wire alu__abc_40887_new_n148_; 
wire alu__abc_40887_new_n149_; 
wire alu__abc_40887_new_n150_; 
wire alu__abc_40887_new_n151_; 
wire alu__abc_40887_new_n152_; 
wire alu__abc_40887_new_n153_; 
wire alu__abc_40887_new_n154_; 
wire alu__abc_40887_new_n155_; 
wire alu__abc_40887_new_n156_; 
wire alu__abc_40887_new_n157_; 
wire alu__abc_40887_new_n158_; 
wire alu__abc_40887_new_n159_; 
wire alu__abc_40887_new_n160_; 
wire alu__abc_40887_new_n161_; 
wire alu__abc_40887_new_n162_; 
wire alu__abc_40887_new_n163_; 
wire alu__abc_40887_new_n164_; 
wire alu__abc_40887_new_n165_; 
wire alu__abc_40887_new_n166_; 
wire alu__abc_40887_new_n167_; 
wire alu__abc_40887_new_n168_; 
wire alu__abc_40887_new_n169_; 
wire alu__abc_40887_new_n170_; 
wire alu__abc_40887_new_n171_; 
wire alu__abc_40887_new_n172_; 
wire alu__abc_40887_new_n173_; 
wire alu__abc_40887_new_n174_; 
wire alu__abc_40887_new_n175_; 
wire alu__abc_40887_new_n176_; 
wire alu__abc_40887_new_n177_; 
wire alu__abc_40887_new_n178_; 
wire alu__abc_40887_new_n179_; 
wire alu__abc_40887_new_n180_; 
wire alu__abc_40887_new_n181_; 
wire alu__abc_40887_new_n182_; 
wire alu__abc_40887_new_n183_; 
wire alu__abc_40887_new_n184_; 
wire alu__abc_40887_new_n185_; 
wire alu__abc_40887_new_n186_; 
wire alu__abc_40887_new_n187_; 
wire alu__abc_40887_new_n188_; 
wire alu__abc_40887_new_n189_; 
wire alu__abc_40887_new_n190_; 
wire alu__abc_40887_new_n191_; 
wire alu__abc_40887_new_n192_; 
wire alu__abc_40887_new_n193_; 
wire alu__abc_40887_new_n194_; 
wire alu__abc_40887_new_n195_; 
wire alu__abc_40887_new_n196_; 
wire alu__abc_40887_new_n197_; 
wire alu__abc_40887_new_n198_; 
wire alu__abc_40887_new_n199_; 
wire alu__abc_40887_new_n200_; 
wire alu__abc_40887_new_n201_; 
wire alu__abc_40887_new_n202_; 
wire alu__abc_40887_new_n203_; 
wire alu__abc_40887_new_n204_; 
wire alu__abc_40887_new_n205_; 
wire alu__abc_40887_new_n206_; 
wire alu__abc_40887_new_n207_; 
wire alu__abc_40887_new_n208_; 
wire alu__abc_40887_new_n209_; 
wire alu__abc_40887_new_n210_; 
wire alu__abc_40887_new_n211_; 
wire alu__abc_40887_new_n212_; 
wire alu__abc_40887_new_n213_; 
wire alu__abc_40887_new_n214_; 
wire alu__abc_40887_new_n215_; 
wire alu__abc_40887_new_n216_; 
wire alu__abc_40887_new_n217_; 
wire alu__abc_40887_new_n218_; 
wire alu__abc_40887_new_n219_; 
wire alu__abc_40887_new_n220_; 
wire alu__abc_40887_new_n221_; 
wire alu__abc_40887_new_n222_; 
wire alu__abc_40887_new_n223_; 
wire alu__abc_40887_new_n224_; 
wire alu__abc_40887_new_n225_; 
wire alu__abc_40887_new_n226_; 
wire alu__abc_40887_new_n227_; 
wire alu__abc_40887_new_n228_; 
wire alu__abc_40887_new_n229_; 
wire alu__abc_40887_new_n230_; 
wire alu__abc_40887_new_n231_; 
wire alu__abc_40887_new_n232_; 
wire alu__abc_40887_new_n233_; 
wire alu__abc_40887_new_n234_; 
wire alu__abc_40887_new_n235_; 
wire alu__abc_40887_new_n236_; 
wire alu__abc_40887_new_n237_; 
wire alu__abc_40887_new_n238_; 
wire alu__abc_40887_new_n239_; 
wire alu__abc_40887_new_n240_; 
wire alu__abc_40887_new_n241_; 
wire alu__abc_40887_new_n242_; 
wire alu__abc_40887_new_n243_; 
wire alu__abc_40887_new_n244_; 
wire alu__abc_40887_new_n245_; 
wire alu__abc_40887_new_n246_; 
wire alu__abc_40887_new_n247_; 
wire alu__abc_40887_new_n248_; 
wire alu__abc_40887_new_n249_; 
wire alu__abc_40887_new_n251_; 
wire alu__abc_40887_new_n252_; 
wire alu__abc_40887_new_n253_; 
wire alu__abc_40887_new_n254_; 
wire alu__abc_40887_new_n255_; 
wire alu__abc_40887_new_n256_; 
wire alu__abc_40887_new_n257_; 
wire alu__abc_40887_new_n258_; 
wire alu__abc_40887_new_n259_; 
wire alu__abc_40887_new_n260_; 
wire alu__abc_40887_new_n261_; 
wire alu__abc_40887_new_n262_; 
wire alu__abc_40887_new_n263_; 
wire alu__abc_40887_new_n264_; 
wire alu__abc_40887_new_n265_; 
wire alu__abc_40887_new_n266_; 
wire alu__abc_40887_new_n267_; 
wire alu__abc_40887_new_n268_; 
wire alu__abc_40887_new_n269_; 
wire alu__abc_40887_new_n270_; 
wire alu__abc_40887_new_n271_; 
wire alu__abc_40887_new_n272_; 
wire alu__abc_40887_new_n273_; 
wire alu__abc_40887_new_n274_; 
wire alu__abc_40887_new_n275_; 
wire alu__abc_40887_new_n276_; 
wire alu__abc_40887_new_n277_; 
wire alu__abc_40887_new_n278_; 
wire alu__abc_40887_new_n279_; 
wire alu__abc_40887_new_n280_; 
wire alu__abc_40887_new_n281_; 
wire alu__abc_40887_new_n282_; 
wire alu__abc_40887_new_n283_; 
wire alu__abc_40887_new_n284_; 
wire alu__abc_40887_new_n285_; 
wire alu__abc_40887_new_n286_; 
wire alu__abc_40887_new_n287_; 
wire alu__abc_40887_new_n288_; 
wire alu__abc_40887_new_n289_; 
wire alu__abc_40887_new_n290_; 
wire alu__abc_40887_new_n291_; 
wire alu__abc_40887_new_n292_; 
wire alu__abc_40887_new_n293_; 
wire alu__abc_40887_new_n294_; 
wire alu__abc_40887_new_n295_; 
wire alu__abc_40887_new_n296_; 
wire alu__abc_40887_new_n297_; 
wire alu__abc_40887_new_n298_; 
wire alu__abc_40887_new_n299_; 
wire alu__abc_40887_new_n300_; 
wire alu__abc_40887_new_n301_; 
wire alu__abc_40887_new_n302_; 
wire alu__abc_40887_new_n303_; 
wire alu__abc_40887_new_n304_; 
wire alu__abc_40887_new_n305_; 
wire alu__abc_40887_new_n306_; 
wire alu__abc_40887_new_n307_; 
wire alu__abc_40887_new_n308_; 
wire alu__abc_40887_new_n309_; 
wire alu__abc_40887_new_n310_; 
wire alu__abc_40887_new_n311_; 
wire alu__abc_40887_new_n312_; 
wire alu__abc_40887_new_n313_; 
wire alu__abc_40887_new_n314_; 
wire alu__abc_40887_new_n315_; 
wire alu__abc_40887_new_n316_; 
wire alu__abc_40887_new_n317_; 
wire alu__abc_40887_new_n318_; 
wire alu__abc_40887_new_n319_; 
wire alu__abc_40887_new_n320_; 
wire alu__abc_40887_new_n321_; 
wire alu__abc_40887_new_n322_; 
wire alu__abc_40887_new_n323_; 
wire alu__abc_40887_new_n324_; 
wire alu__abc_40887_new_n325_; 
wire alu__abc_40887_new_n326_; 
wire alu__abc_40887_new_n327_; 
wire alu__abc_40887_new_n328_; 
wire alu__abc_40887_new_n329_; 
wire alu__abc_40887_new_n330_; 
wire alu__abc_40887_new_n331_; 
wire alu__abc_40887_new_n332_; 
wire alu__abc_40887_new_n333_; 
wire alu__abc_40887_new_n334_; 
wire alu__abc_40887_new_n335_; 
wire alu__abc_40887_new_n336_; 
wire alu__abc_40887_new_n337_; 
wire alu__abc_40887_new_n338_; 
wire alu__abc_40887_new_n339_; 
wire alu__abc_40887_new_n33_; 
wire alu__abc_40887_new_n340_; 
wire alu__abc_40887_new_n341_; 
wire alu__abc_40887_new_n342_; 
wire alu__abc_40887_new_n343_; 
wire alu__abc_40887_new_n344_; 
wire alu__abc_40887_new_n345_; 
wire alu__abc_40887_new_n346_; 
wire alu__abc_40887_new_n347_; 
wire alu__abc_40887_new_n348_; 
wire alu__abc_40887_new_n349_; 
wire alu__abc_40887_new_n34_; 
wire alu__abc_40887_new_n350_; 
wire alu__abc_40887_new_n351_; 
wire alu__abc_40887_new_n352_; 
wire alu__abc_40887_new_n353_; 
wire alu__abc_40887_new_n354_; 
wire alu__abc_40887_new_n355_; 
wire alu__abc_40887_new_n356_; 
wire alu__abc_40887_new_n357_; 
wire alu__abc_40887_new_n358_; 
wire alu__abc_40887_new_n359_; 
wire alu__abc_40887_new_n35_; 
wire alu__abc_40887_new_n360_; 
wire alu__abc_40887_new_n361_; 
wire alu__abc_40887_new_n362_; 
wire alu__abc_40887_new_n363_; 
wire alu__abc_40887_new_n364_; 
wire alu__abc_40887_new_n365_; 
wire alu__abc_40887_new_n366_; 
wire alu__abc_40887_new_n367_; 
wire alu__abc_40887_new_n368_; 
wire alu__abc_40887_new_n369_; 
wire alu__abc_40887_new_n36_; 
wire alu__abc_40887_new_n370_; 
wire alu__abc_40887_new_n371_; 
wire alu__abc_40887_new_n372_; 
wire alu__abc_40887_new_n373_; 
wire alu__abc_40887_new_n374_; 
wire alu__abc_40887_new_n375_; 
wire alu__abc_40887_new_n376_; 
wire alu__abc_40887_new_n377_; 
wire alu__abc_40887_new_n378_; 
wire alu__abc_40887_new_n379_; 
wire alu__abc_40887_new_n37_; 
wire alu__abc_40887_new_n380_; 
wire alu__abc_40887_new_n381_; 
wire alu__abc_40887_new_n382_; 
wire alu__abc_40887_new_n383_; 
wire alu__abc_40887_new_n384_; 
wire alu__abc_40887_new_n385_; 
wire alu__abc_40887_new_n386_; 
wire alu__abc_40887_new_n387_; 
wire alu__abc_40887_new_n388_; 
wire alu__abc_40887_new_n389_; 
wire alu__abc_40887_new_n38_; 
wire alu__abc_40887_new_n390_; 
wire alu__abc_40887_new_n391_; 
wire alu__abc_40887_new_n392_; 
wire alu__abc_40887_new_n393_; 
wire alu__abc_40887_new_n394_; 
wire alu__abc_40887_new_n395_; 
wire alu__abc_40887_new_n396_; 
wire alu__abc_40887_new_n397_; 
wire alu__abc_40887_new_n398_; 
wire alu__abc_40887_new_n399_; 
wire alu__abc_40887_new_n39_; 
wire alu__abc_40887_new_n400_; 
wire alu__abc_40887_new_n401_; 
wire alu__abc_40887_new_n402_; 
wire alu__abc_40887_new_n403_; 
wire alu__abc_40887_new_n404_; 
wire alu__abc_40887_new_n405_; 
wire alu__abc_40887_new_n406_; 
wire alu__abc_40887_new_n407_; 
wire alu__abc_40887_new_n408_; 
wire alu__abc_40887_new_n409_; 
wire alu__abc_40887_new_n40_; 
wire alu__abc_40887_new_n410_; 
wire alu__abc_40887_new_n411_; 
wire alu__abc_40887_new_n412_; 
wire alu__abc_40887_new_n413_; 
wire alu__abc_40887_new_n414_; 
wire alu__abc_40887_new_n415_; 
wire alu__abc_40887_new_n416_; 
wire alu__abc_40887_new_n417_; 
wire alu__abc_40887_new_n418_; 
wire alu__abc_40887_new_n419_; 
wire alu__abc_40887_new_n41_; 
wire alu__abc_40887_new_n420_; 
wire alu__abc_40887_new_n421_; 
wire alu__abc_40887_new_n422_; 
wire alu__abc_40887_new_n423_; 
wire alu__abc_40887_new_n424_; 
wire alu__abc_40887_new_n425_; 
wire alu__abc_40887_new_n426_; 
wire alu__abc_40887_new_n427_; 
wire alu__abc_40887_new_n428_; 
wire alu__abc_40887_new_n429_; 
wire alu__abc_40887_new_n42_; 
wire alu__abc_40887_new_n430_; 
wire alu__abc_40887_new_n431_; 
wire alu__abc_40887_new_n432_; 
wire alu__abc_40887_new_n433_; 
wire alu__abc_40887_new_n434_; 
wire alu__abc_40887_new_n435_; 
wire alu__abc_40887_new_n436_; 
wire alu__abc_40887_new_n437_; 
wire alu__abc_40887_new_n438_; 
wire alu__abc_40887_new_n439_; 
wire alu__abc_40887_new_n43_; 
wire alu__abc_40887_new_n440_; 
wire alu__abc_40887_new_n441_; 
wire alu__abc_40887_new_n442_; 
wire alu__abc_40887_new_n443_; 
wire alu__abc_40887_new_n444_; 
wire alu__abc_40887_new_n445_; 
wire alu__abc_40887_new_n446_; 
wire alu__abc_40887_new_n447_; 
wire alu__abc_40887_new_n448_; 
wire alu__abc_40887_new_n449_; 
wire alu__abc_40887_new_n44_; 
wire alu__abc_40887_new_n450_; 
wire alu__abc_40887_new_n451_; 
wire alu__abc_40887_new_n452_; 
wire alu__abc_40887_new_n453_; 
wire alu__abc_40887_new_n454_; 
wire alu__abc_40887_new_n455_; 
wire alu__abc_40887_new_n456_; 
wire alu__abc_40887_new_n457_; 
wire alu__abc_40887_new_n459_; 
wire alu__abc_40887_new_n45_; 
wire alu__abc_40887_new_n460_; 
wire alu__abc_40887_new_n462_; 
wire alu__abc_40887_new_n463_; 
wire alu__abc_40887_new_n464_; 
wire alu__abc_40887_new_n466_; 
wire alu__abc_40887_new_n467_; 
wire alu__abc_40887_new_n469_; 
wire alu__abc_40887_new_n46_; 
wire alu__abc_40887_new_n470_; 
wire alu__abc_40887_new_n472_; 
wire alu__abc_40887_new_n473_; 
wire alu__abc_40887_new_n475_; 
wire alu__abc_40887_new_n476_; 
wire alu__abc_40887_new_n478_; 
wire alu__abc_40887_new_n479_; 
wire alu__abc_40887_new_n47_; 
wire alu__abc_40887_new_n481_; 
wire alu__abc_40887_new_n482_; 
wire alu__abc_40887_new_n484_; 
wire alu__abc_40887_new_n485_; 
wire alu__abc_40887_new_n487_; 
wire alu__abc_40887_new_n488_; 
wire alu__abc_40887_new_n489_; 
wire alu__abc_40887_new_n48_; 
wire alu__abc_40887_new_n490_; 
wire alu__abc_40887_new_n491_; 
wire alu__abc_40887_new_n492_; 
wire alu__abc_40887_new_n493_; 
wire alu__abc_40887_new_n494_; 
wire alu__abc_40887_new_n495_; 
wire alu__abc_40887_new_n496_; 
wire alu__abc_40887_new_n497_; 
wire alu__abc_40887_new_n498_; 
wire alu__abc_40887_new_n499_; 
wire alu__abc_40887_new_n49_; 
wire alu__abc_40887_new_n50_; 
wire alu__abc_40887_new_n51_; 
wire alu__abc_40887_new_n52_; 
wire alu__abc_40887_new_n53_; 
wire alu__abc_40887_new_n54_; 
wire alu__abc_40887_new_n55_; 
wire alu__abc_40887_new_n56_; 
wire alu__abc_40887_new_n57_; 
wire alu__abc_40887_new_n58_; 
wire alu__abc_40887_new_n59_; 
wire alu__abc_40887_new_n60_; 
wire alu__abc_40887_new_n61_; 
wire alu__abc_40887_new_n62_; 
wire alu__abc_40887_new_n63_; 
wire alu__abc_40887_new_n64_; 
wire alu__abc_40887_new_n65_; 
wire alu__abc_40887_new_n66_; 
wire alu__abc_40887_new_n67_; 
wire alu__abc_40887_new_n68_; 
wire alu__abc_40887_new_n69_; 
wire alu__abc_40887_new_n70_; 
wire alu__abc_40887_new_n71_; 
wire alu__abc_40887_new_n72_; 
wire alu__abc_40887_new_n73_; 
wire alu__abc_40887_new_n74_; 
wire alu__abc_40887_new_n75_; 
wire alu__abc_40887_new_n76_; 
wire alu__abc_40887_new_n77_; 
wire alu__abc_40887_new_n78_; 
wire alu__abc_40887_new_n79_; 
wire alu__abc_40887_new_n80_; 
wire alu__abc_40887_new_n81_; 
wire alu__abc_40887_new_n82_; 
wire alu__abc_40887_new_n83_; 
wire alu__abc_40887_new_n84_; 
wire alu__abc_40887_new_n85_; 
wire alu__abc_40887_new_n86_; 
wire alu__abc_40887_new_n87_; 
wire alu__abc_40887_new_n88_; 
wire alu__abc_40887_new_n89_; 
wire alu__abc_40887_new_n90_; 
wire alu__abc_40887_new_n91_; 
wire alu__abc_40887_new_n92_; 
wire alu__abc_40887_new_n93_; 
wire alu__abc_40887_new_n94_; 
wire alu__abc_40887_new_n95_; 
wire alu__abc_40887_new_n96_; 
wire alu__abc_40887_new_n97_; 
wire alu__abc_40887_new_n98_; 
wire alu__abc_40887_new_n99_; 
wire alu_cin; 
wire alu_cout; 
wire alu_opra_0_; 
wire alu_opra_1_; 
wire alu_opra_2_; 
wire alu_opra_3_; 
wire alu_opra_4_; 
wire alu_opra_5_; 
wire alu_opra_6_; 
wire alu_opra_7_; 
wire alu_oprb_0_; 
wire alu_oprb_1_; 
wire alu_oprb_2_; 
wire alu_oprb_3_; 
wire alu_oprb_4_; 
wire alu_oprb_5_; 
wire alu_oprb_6_; 
wire alu_oprb_7_; 
wire alu_parity; 
wire alu_res_0_; 
wire alu_res_1_; 
wire alu_res_2_; 
wire alu_res_3_; 
wire alu_res_4_; 
wire alu_res_5_; 
wire alu_res_6_; 
wire alu_res_7_; 
wire alu_sel_0_; 
wire alu_sel_1_; 
wire alu_sel_2_; 
wire alu_sout; 
wire alu_zout; 
wire auxcar; 
wire carry; 
input clock;
input \data[0] ;
input \data[1] ;
input \data[2] ;
input \data[3] ;
input \data[4] ;
input \data[5] ;
input \data[6] ;
input \data[7] ;
wire ei; 
wire eienb; 
output inta;
wire intcyc; 
input intr;
wire opcode_0_; 
wire opcode_1_; 
wire opcode_2_; 
wire opcode_3_; 
wire opcode_4_; 
wire opcode_5_; 
wire opcode_6_; 
wire opcode_7_; 
wire parity; 
wire pc_0_; 
wire pc_10_; 
wire pc_11_; 
wire pc_12_; 
wire pc_13_; 
wire pc_14_; 
wire pc_15_; 
wire pc_1_; 
wire pc_2_; 
wire pc_3_; 
wire pc_4_; 
wire pc_5_; 
wire pc_6_; 
wire pc_7_; 
wire pc_8_; 
wire pc_9_; 
wire popdes_0_; 
wire popdes_1_; 
wire raddrhold_0_; 
wire raddrhold_10_; 
wire raddrhold_11_; 
wire raddrhold_12_; 
wire raddrhold_13_; 
wire raddrhold_14_; 
wire raddrhold_15_; 
wire raddrhold_1_; 
wire raddrhold_2_; 
wire raddrhold_3_; 
wire raddrhold_4_; 
wire raddrhold_5_; 
wire raddrhold_6_; 
wire raddrhold_7_; 
wire raddrhold_8_; 
wire raddrhold_9_; 
wire rdatahold2_0_; 
wire rdatahold2_1_; 
wire rdatahold2_2_; 
wire rdatahold2_3_; 
wire rdatahold2_4_; 
wire rdatahold2_5_; 
wire rdatahold2_6_; 
wire rdatahold2_7_; 
wire rdatahold_0_; 
wire rdatahold_1_; 
wire rdatahold_2_; 
wire rdatahold_3_; 
wire rdatahold_4_; 
wire rdatahold_5_; 
wire rdatahold_6_; 
wire rdatahold_7_; 
output readio;
output readmem;
wire regd_0_; 
wire regd_1_; 
wire regd_2_; 
wire regfil_0__0_; 
wire regfil_0__1_; 
wire regfil_0__2_; 
wire regfil_0__3_; 
wire regfil_0__4_; 
wire regfil_0__5_; 
wire regfil_0__6_; 
wire regfil_0__7_; 
wire regfil_1__0_; 
wire regfil_1__1_; 
wire regfil_1__2_; 
wire regfil_1__3_; 
wire regfil_1__4_; 
wire regfil_1__5_; 
wire regfil_1__6_; 
wire regfil_1__7_; 
wire regfil_2__0_; 
wire regfil_2__1_; 
wire regfil_2__2_; 
wire regfil_2__3_; 
wire regfil_2__4_; 
wire regfil_2__5_; 
wire regfil_2__6_; 
wire regfil_2__7_; 
wire regfil_3__0_; 
wire regfil_3__1_; 
wire regfil_3__2_; 
wire regfil_3__3_; 
wire regfil_3__4_; 
wire regfil_3__5_; 
wire regfil_3__6_; 
wire regfil_3__7_; 
wire regfil_4__0_; 
wire regfil_4__1_; 
wire regfil_4__2_; 
wire regfil_4__3_; 
wire regfil_4__4_; 
wire regfil_4__5_; 
wire regfil_4__6_; 
wire regfil_4__7_; 
wire regfil_5__0_; 
wire regfil_5__1_; 
wire regfil_5__2_; 
wire regfil_5__3_; 
wire regfil_5__4_; 
wire regfil_5__5_; 
wire regfil_5__6_; 
wire regfil_5__7_; 
wire regfil_6__0_; 
wire regfil_6__1_; 
wire regfil_6__2_; 
wire regfil_6__3_; 
wire regfil_6__4_; 
wire regfil_6__5_; 
wire regfil_6__6_; 
wire regfil_6__7_; 
wire regfil_7__0_; 
wire regfil_7__1_; 
wire regfil_7__2_; 
wire regfil_7__3_; 
wire regfil_7__4_; 
wire regfil_7__5_; 
wire regfil_7__6_; 
wire regfil_7__7_; 
input reset;
wire sign; 
wire sp_0_; 
wire sp_10_; 
wire sp_11_; 
wire sp_12_; 
wire sp_13_; 
wire sp_14_; 
wire sp_15_; 
wire sp_1_; 
wire sp_2_; 
wire sp_3_; 
wire sp_4_; 
wire sp_5_; 
wire sp_6_; 
wire sp_7_; 
wire sp_8_; 
wire sp_9_; 
wire state_0_; 
wire state_1_; 
wire state_2_; 
wire state_3_; 
wire state_4_; 
wire state_5_; 
wire statesel_0_; 
wire statesel_1_; 
wire statesel_2_; 
wire statesel_3_; 
wire statesel_4_; 
wire statesel_5_; 
wire waddrhold_0_; 
wire waddrhold_10_; 
wire waddrhold_11_; 
wire waddrhold_12_; 
wire waddrhold_13_; 
wire waddrhold_14_; 
wire waddrhold_15_; 
wire waddrhold_1_; 
wire waddrhold_2_; 
wire waddrhold_3_; 
wire waddrhold_4_; 
wire waddrhold_5_; 
wire waddrhold_6_; 
wire waddrhold_7_; 
wire waddrhold_8_; 
wire waddrhold_9_; 
input waitr;
wire wdatahold2_0_; 
wire wdatahold2_1_; 
wire wdatahold2_2_; 
wire wdatahold2_3_; 
wire wdatahold2_4_; 
wire wdatahold2_5_; 
wire wdatahold2_6_; 
wire wdatahold2_7_; 
wire wdatahold_0_; 
wire wdatahold_1_; 
wire wdatahold_2_; 
wire wdatahold_3_; 
wire wdatahold_4_; 
wire wdatahold_5_; 
wire wdatahold_6_; 
wire wdatahold_7_; 
output writeio;
output writemem;
wire zero; 
AND2X2 AND2X2_1 ( .A(_abc_41356_new_n501_), .B(state_4_), .Y(_abc_41356_new_n502_));
AND2X2 AND2X2_10 ( .A(_abc_41356_new_n501_), .B(_abc_41356_new_n517_), .Y(_abc_41356_new_n518_));
AND2X2 AND2X2_100 ( .A(_abc_41356_new_n666_), .B(_abc_41356_new_n664_), .Y(_abc_41356_new_n667_));
AND2X2 AND2X2_1000 ( .A(_abc_41356_new_n1235_), .B(regfil_5__2_), .Y(_abc_41356_new_n2444_));
AND2X2 AND2X2_1001 ( .A(_abc_41356_new_n2449_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2450_));
AND2X2 AND2X2_1002 ( .A(_abc_41356_new_n2448_), .B(_abc_41356_new_n2450_), .Y(_abc_41356_new_n2451_));
AND2X2 AND2X2_1003 ( .A(_abc_41356_new_n2393_), .B(rdatahold2_3_), .Y(_abc_41356_new_n2452_));
AND2X2 AND2X2_1004 ( .A(_abc_41356_new_n2433_), .B(_abc_41356_new_n1356_), .Y(_abc_41356_new_n2453_));
AND2X2 AND2X2_1005 ( .A(_abc_41356_new_n2454_), .B(regfil_3__3_), .Y(_abc_41356_new_n2455_));
AND2X2 AND2X2_1006 ( .A(_abc_41356_new_n2412_), .B(_abc_41356_new_n2456_), .Y(_abc_41356_new_n2457_));
AND2X2 AND2X2_1007 ( .A(_abc_41356_new_n2439_), .B(regfil_3__3_), .Y(_abc_41356_new_n2459_));
AND2X2 AND2X2_1008 ( .A(_abc_41356_new_n2460_), .B(_abc_41356_new_n2458_), .Y(_abc_41356_new_n2461_));
AND2X2 AND2X2_1009 ( .A(_abc_41356_new_n2415_), .B(_abc_41356_new_n2461_), .Y(_abc_41356_new_n2462_));
AND2X2 AND2X2_101 ( .A(_abc_41356_new_n604_), .B(_abc_41356_new_n667_), .Y(_abc_41356_new_n668_));
AND2X2 AND2X2_1010 ( .A(_abc_41356_new_n1235_), .B(regfil_5__3_), .Y(_abc_41356_new_n2464_));
AND2X2 AND2X2_1011 ( .A(_abc_41356_new_n2469_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2470_));
AND2X2 AND2X2_1012 ( .A(_abc_41356_new_n2468_), .B(_abc_41356_new_n2470_), .Y(_abc_41356_new_n2471_));
AND2X2 AND2X2_1013 ( .A(_abc_41356_new_n2393_), .B(rdatahold2_4_), .Y(_abc_41356_new_n2472_));
AND2X2 AND2X2_1014 ( .A(_abc_41356_new_n2473_), .B(regfil_3__4_), .Y(_abc_41356_new_n2476_));
AND2X2 AND2X2_1015 ( .A(_abc_41356_new_n2477_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2478_));
AND2X2 AND2X2_1016 ( .A(_abc_41356_new_n2459_), .B(regfil_3__4_), .Y(_abc_41356_new_n2480_));
AND2X2 AND2X2_1017 ( .A(_abc_41356_new_n2481_), .B(_abc_41356_new_n2479_), .Y(_abc_41356_new_n2482_));
AND2X2 AND2X2_1018 ( .A(_abc_41356_new_n2415_), .B(_abc_41356_new_n2482_), .Y(_abc_41356_new_n2483_));
AND2X2 AND2X2_1019 ( .A(_abc_41356_new_n1235_), .B(regfil_5__4_), .Y(_abc_41356_new_n2485_));
AND2X2 AND2X2_102 ( .A(_abc_41356_new_n614_), .B(_abc_41356_new_n534_), .Y(_abc_41356_new_n670_));
AND2X2 AND2X2_1020 ( .A(_abc_41356_new_n2490_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2491_));
AND2X2 AND2X2_1021 ( .A(_abc_41356_new_n2489_), .B(_abc_41356_new_n2491_), .Y(_abc_41356_new_n2492_));
AND2X2 AND2X2_1022 ( .A(_abc_41356_new_n2393_), .B(rdatahold2_5_), .Y(_abc_41356_new_n2493_));
AND2X2 AND2X2_1023 ( .A(_abc_41356_new_n2474_), .B(regfil_3__5_), .Y(_abc_41356_new_n2496_));
AND2X2 AND2X2_1024 ( .A(_abc_41356_new_n2497_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2498_));
AND2X2 AND2X2_1025 ( .A(_abc_41356_new_n2480_), .B(regfil_3__5_), .Y(_abc_41356_new_n2499_));
AND2X2 AND2X2_1026 ( .A(_abc_41356_new_n2500_), .B(_abc_41356_new_n2501_), .Y(_abc_41356_new_n2502_));
AND2X2 AND2X2_1027 ( .A(_abc_41356_new_n2415_), .B(_abc_41356_new_n2502_), .Y(_abc_41356_new_n2503_));
AND2X2 AND2X2_1028 ( .A(_abc_41356_new_n1235_), .B(regfil_5__5_), .Y(_abc_41356_new_n2505_));
AND2X2 AND2X2_1029 ( .A(_abc_41356_new_n2510_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2511_));
AND2X2 AND2X2_103 ( .A(_abc_41356_new_n671_), .B(_abc_41356_new_n669_), .Y(_abc_41356_new_n672_));
AND2X2 AND2X2_1030 ( .A(_abc_41356_new_n2509_), .B(_abc_41356_new_n2511_), .Y(_abc_41356_new_n2512_));
AND2X2 AND2X2_1031 ( .A(_abc_41356_new_n2393_), .B(rdatahold2_6_), .Y(_abc_41356_new_n2513_));
AND2X2 AND2X2_1032 ( .A(_abc_41356_new_n2494_), .B(regfil_3__6_), .Y(_abc_41356_new_n2516_));
AND2X2 AND2X2_1033 ( .A(_abc_41356_new_n2517_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2518_));
AND2X2 AND2X2_1034 ( .A(_abc_41356_new_n2499_), .B(regfil_3__6_), .Y(_abc_41356_new_n2519_));
AND2X2 AND2X2_1035 ( .A(_abc_41356_new_n2415_), .B(_abc_41356_new_n2521_), .Y(_abc_41356_new_n2522_));
AND2X2 AND2X2_1036 ( .A(_abc_41356_new_n2522_), .B(_abc_41356_new_n2520_), .Y(_abc_41356_new_n2523_));
AND2X2 AND2X2_1037 ( .A(_abc_41356_new_n1235_), .B(regfil_5__6_), .Y(_abc_41356_new_n2525_));
AND2X2 AND2X2_1038 ( .A(_abc_41356_new_n2530_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2531_));
AND2X2 AND2X2_1039 ( .A(_abc_41356_new_n2529_), .B(_abc_41356_new_n2531_), .Y(_abc_41356_new_n2532_));
AND2X2 AND2X2_104 ( .A(_abc_41356_new_n668_), .B(_abc_41356_new_n672_), .Y(_abc_41356_new_n673_));
AND2X2 AND2X2_1040 ( .A(_abc_41356_new_n2393_), .B(rdatahold2_7_), .Y(_abc_41356_new_n2533_));
AND2X2 AND2X2_1041 ( .A(_abc_41356_new_n2514_), .B(regfil_3__7_), .Y(_abc_41356_new_n2536_));
AND2X2 AND2X2_1042 ( .A(_abc_41356_new_n2537_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2538_));
AND2X2 AND2X2_1043 ( .A(_abc_41356_new_n2519_), .B(regfil_3__7_), .Y(_abc_41356_new_n2540_));
AND2X2 AND2X2_1044 ( .A(_abc_41356_new_n2541_), .B(_abc_41356_new_n2415_), .Y(_abc_41356_new_n2542_));
AND2X2 AND2X2_1045 ( .A(_abc_41356_new_n2542_), .B(_abc_41356_new_n2539_), .Y(_abc_41356_new_n2543_));
AND2X2 AND2X2_1046 ( .A(_abc_41356_new_n1235_), .B(regfil_5__7_), .Y(_abc_41356_new_n2545_));
AND2X2 AND2X2_1047 ( .A(_abc_41356_new_n2383_), .B(_abc_41356_new_n1208_), .Y(_abc_41356_new_n2549_));
AND2X2 AND2X2_1048 ( .A(_abc_41356_new_n694_), .B(_abc_41356_new_n2549_), .Y(_abc_41356_new_n2550_));
AND2X2 AND2X2_1049 ( .A(_abc_41356_new_n2553_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n2554_));
AND2X2 AND2X2_105 ( .A(_abc_41356_new_n522_), .B(_abc_41356_new_n518_), .Y(_abc_41356_new_n676_));
AND2X2 AND2X2_1050 ( .A(_abc_41356_new_n2552_), .B(_abc_41356_new_n2554_), .Y(_abc_41356_new_n2555_));
AND2X2 AND2X2_1051 ( .A(_abc_41356_new_n2419_), .B(_abc_41356_new_n1224_), .Y(_abc_41356_new_n2556_));
AND2X2 AND2X2_1052 ( .A(_abc_41356_new_n2557_), .B(_abc_41356_new_n647_), .Y(_abc_41356_new_n2558_));
AND2X2 AND2X2_1053 ( .A(_abc_41356_new_n1082_), .B(_abc_41356_new_n2558_), .Y(_abc_41356_new_n2559_));
AND2X2 AND2X2_1054 ( .A(_abc_41356_new_n595_), .B(rdatahold2_0_), .Y(_abc_41356_new_n2560_));
AND2X2 AND2X2_1055 ( .A(_abc_41356_new_n2564_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n2565_));
AND2X2 AND2X2_1056 ( .A(_abc_41356_new_n2563_), .B(_abc_41356_new_n2565_), .Y(_abc_41356_new_n2566_));
AND2X2 AND2X2_1057 ( .A(_abc_41356_new_n2570_), .B(_abc_41356_new_n2557_), .Y(_abc_41356_new_n2571_));
AND2X2 AND2X2_1058 ( .A(_abc_41356_new_n2571_), .B(_abc_41356_new_n2568_), .Y(_abc_41356_new_n2572_));
AND2X2 AND2X2_1059 ( .A(_abc_41356_new_n595_), .B(rdatahold2_1_), .Y(_abc_41356_new_n2573_));
AND2X2 AND2X2_106 ( .A(_abc_41356_new_n623_), .B(opcode_2_), .Y(_abc_41356_new_n677_));
AND2X2 AND2X2_1060 ( .A(_abc_41356_new_n2577_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n2578_));
AND2X2 AND2X2_1061 ( .A(_abc_41356_new_n2576_), .B(_abc_41356_new_n2578_), .Y(_abc_41356_new_n2579_));
AND2X2 AND2X2_1062 ( .A(_abc_41356_new_n2580_), .B(regfil_1__2_), .Y(_abc_41356_new_n2581_));
AND2X2 AND2X2_1063 ( .A(_abc_41356_new_n601_), .B(_abc_41356_new_n2582_), .Y(_abc_41356_new_n2583_));
AND2X2 AND2X2_1064 ( .A(_abc_41356_new_n2584_), .B(_abc_41356_new_n2585_), .Y(_abc_41356_new_n2586_));
AND2X2 AND2X2_1065 ( .A(_abc_41356_new_n581_), .B(_abc_41356_new_n2586_), .Y(_abc_41356_new_n2587_));
AND2X2 AND2X2_1066 ( .A(_abc_41356_new_n595_), .B(rdatahold2_2_), .Y(_abc_41356_new_n2589_));
AND2X2 AND2X2_1067 ( .A(_abc_41356_new_n2593_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n2594_));
AND2X2 AND2X2_1068 ( .A(_abc_41356_new_n2592_), .B(_abc_41356_new_n2594_), .Y(_abc_41356_new_n2595_));
AND2X2 AND2X2_1069 ( .A(_abc_41356_new_n2596_), .B(regfil_1__3_), .Y(_abc_41356_new_n2597_));
AND2X2 AND2X2_107 ( .A(_abc_41356_new_n515_), .B(opcode_6_), .Y(_abc_41356_new_n679_));
AND2X2 AND2X2_1070 ( .A(_abc_41356_new_n601_), .B(_abc_41356_new_n2598_), .Y(_abc_41356_new_n2599_));
AND2X2 AND2X2_1071 ( .A(_abc_41356_new_n2600_), .B(_abc_41356_new_n2601_), .Y(_abc_41356_new_n2602_));
AND2X2 AND2X2_1072 ( .A(_abc_41356_new_n581_), .B(_abc_41356_new_n2602_), .Y(_abc_41356_new_n2603_));
AND2X2 AND2X2_1073 ( .A(_abc_41356_new_n595_), .B(rdatahold2_3_), .Y(_abc_41356_new_n2605_));
AND2X2 AND2X2_1074 ( .A(_abc_41356_new_n2609_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n2610_));
AND2X2 AND2X2_1075 ( .A(_abc_41356_new_n2608_), .B(_abc_41356_new_n2610_), .Y(_abc_41356_new_n2611_));
AND2X2 AND2X2_1076 ( .A(_abc_41356_new_n652_), .B(regfil_1__4_), .Y(_abc_41356_new_n2613_));
AND2X2 AND2X2_1077 ( .A(_abc_41356_new_n2614_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n2615_));
AND2X2 AND2X2_1078 ( .A(_abc_41356_new_n2616_), .B(_abc_41356_new_n2617_), .Y(_abc_41356_new_n2618_));
AND2X2 AND2X2_1079 ( .A(_abc_41356_new_n581_), .B(_abc_41356_new_n2618_), .Y(_abc_41356_new_n2619_));
AND2X2 AND2X2_108 ( .A(_abc_41356_new_n679_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n680_));
AND2X2 AND2X2_1080 ( .A(_abc_41356_new_n595_), .B(rdatahold2_4_), .Y(_abc_41356_new_n2621_));
AND2X2 AND2X2_1081 ( .A(_abc_41356_new_n2625_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n2626_));
AND2X2 AND2X2_1082 ( .A(_abc_41356_new_n2624_), .B(_abc_41356_new_n2626_), .Y(_abc_41356_new_n2627_));
AND2X2 AND2X2_1083 ( .A(_abc_41356_new_n653_), .B(regfil_1__5_), .Y(_abc_41356_new_n2629_));
AND2X2 AND2X2_1084 ( .A(_abc_41356_new_n2630_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n2631_));
AND2X2 AND2X2_1085 ( .A(_abc_41356_new_n2632_), .B(_abc_41356_new_n2633_), .Y(_abc_41356_new_n2634_));
AND2X2 AND2X2_1086 ( .A(_abc_41356_new_n2634_), .B(_abc_41356_new_n581_), .Y(_abc_41356_new_n2635_));
AND2X2 AND2X2_1087 ( .A(_abc_41356_new_n595_), .B(rdatahold2_5_), .Y(_abc_41356_new_n2637_));
AND2X2 AND2X2_1088 ( .A(_abc_41356_new_n2641_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n2642_));
AND2X2 AND2X2_1089 ( .A(_abc_41356_new_n2640_), .B(_abc_41356_new_n2642_), .Y(_abc_41356_new_n2643_));
AND2X2 AND2X2_109 ( .A(opcode_4_), .B(opcode_5_), .Y(_abc_41356_new_n681_));
AND2X2 AND2X2_1090 ( .A(_abc_41356_new_n595_), .B(rdatahold2_6_), .Y(_abc_41356_new_n2644_));
AND2X2 AND2X2_1091 ( .A(_abc_41356_new_n654_), .B(regfil_1__6_), .Y(_abc_41356_new_n2646_));
AND2X2 AND2X2_1092 ( .A(_abc_41356_new_n2647_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n2648_));
AND2X2 AND2X2_1093 ( .A(_abc_41356_new_n2650_), .B(_abc_41356_new_n581_), .Y(_abc_41356_new_n2651_));
AND2X2 AND2X2_1094 ( .A(_abc_41356_new_n2651_), .B(_abc_41356_new_n2649_), .Y(_abc_41356_new_n2652_));
AND2X2 AND2X2_1095 ( .A(_abc_41356_new_n2657_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n2658_));
AND2X2 AND2X2_1096 ( .A(_abc_41356_new_n2656_), .B(_abc_41356_new_n2658_), .Y(_abc_41356_new_n2659_));
AND2X2 AND2X2_1097 ( .A(_abc_41356_new_n595_), .B(rdatahold2_7_), .Y(_abc_41356_new_n2660_));
AND2X2 AND2X2_1098 ( .A(_abc_41356_new_n655_), .B(regfil_1__7_), .Y(_abc_41356_new_n2661_));
AND2X2 AND2X2_1099 ( .A(_abc_41356_new_n2662_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n2663_));
AND2X2 AND2X2_11 ( .A(_abc_41356_new_n518_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n519_));
AND2X2 AND2X2_110 ( .A(_abc_41356_new_n681_), .B(_abc_41356_new_n545_), .Y(_abc_41356_new_n682_));
AND2X2 AND2X2_1100 ( .A(_abc_41356_new_n2665_), .B(_abc_41356_new_n581_), .Y(_abc_41356_new_n2666_));
AND2X2 AND2X2_1101 ( .A(_abc_41356_new_n2666_), .B(_abc_41356_new_n2664_), .Y(_abc_41356_new_n2667_));
AND2X2 AND2X2_1102 ( .A(_abc_41356_new_n1211_), .B(_abc_41356_new_n673_), .Y(_abc_41356_new_n2671_));
AND2X2 AND2X2_1103 ( .A(_abc_41356_new_n2673_), .B(_abc_41356_new_n2674_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_0_));
AND2X2 AND2X2_1104 ( .A(_abc_41356_new_n2676_), .B(_abc_41356_new_n2677_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_1_));
AND2X2 AND2X2_1105 ( .A(_abc_41356_new_n2679_), .B(_abc_41356_new_n2680_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_2_));
AND2X2 AND2X2_1106 ( .A(_abc_41356_new_n2682_), .B(_abc_41356_new_n2683_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_3_));
AND2X2 AND2X2_1107 ( .A(_abc_41356_new_n2685_), .B(_abc_41356_new_n2686_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_4_));
AND2X2 AND2X2_1108 ( .A(_abc_41356_new_n2688_), .B(_abc_41356_new_n2689_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_5_));
AND2X2 AND2X2_1109 ( .A(_abc_41356_new_n2691_), .B(_abc_41356_new_n2692_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_6_));
AND2X2 AND2X2_111 ( .A(_abc_41356_new_n683_), .B(_abc_41356_new_n680_), .Y(_abc_41356_new_n684_));
AND2X2 AND2X2_1110 ( .A(_abc_41356_new_n2694_), .B(_abc_41356_new_n2695_), .Y(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_7_));
AND2X2 AND2X2_1111 ( .A(_abc_41356_new_n1211_), .B(_abc_41356_new_n2384_), .Y(_abc_41356_new_n2697_));
AND2X2 AND2X2_1112 ( .A(_abc_41356_new_n2700_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2701_));
AND2X2 AND2X2_1113 ( .A(_abc_41356_new_n2699_), .B(_abc_41356_new_n2701_), .Y(_abc_41356_new_n2702_));
AND2X2 AND2X2_1114 ( .A(_abc_41356_new_n2393_), .B(rdatahold_0_), .Y(_abc_41356_new_n2703_));
AND2X2 AND2X2_1115 ( .A(_abc_41356_new_n2534_), .B(regfil_2__0_), .Y(_abc_41356_new_n2706_));
AND2X2 AND2X2_1116 ( .A(_abc_41356_new_n2707_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2708_));
AND2X2 AND2X2_1117 ( .A(_abc_41356_new_n2540_), .B(regfil_2__0_), .Y(_abc_41356_new_n2710_));
AND2X2 AND2X2_1118 ( .A(_abc_41356_new_n2711_), .B(_abc_41356_new_n2415_), .Y(_abc_41356_new_n2712_));
AND2X2 AND2X2_1119 ( .A(_abc_41356_new_n2712_), .B(_abc_41356_new_n2709_), .Y(_abc_41356_new_n2713_));
AND2X2 AND2X2_112 ( .A(_abc_41356_new_n684_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n685_));
AND2X2 AND2X2_1120 ( .A(_abc_41356_new_n1235_), .B(regfil_4__0_), .Y(_abc_41356_new_n2715_));
AND2X2 AND2X2_1121 ( .A(_abc_41356_new_n2720_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2721_));
AND2X2 AND2X2_1122 ( .A(_abc_41356_new_n2719_), .B(_abc_41356_new_n2721_), .Y(_abc_41356_new_n2722_));
AND2X2 AND2X2_1123 ( .A(_abc_41356_new_n2393_), .B(rdatahold_1_), .Y(_abc_41356_new_n2723_));
AND2X2 AND2X2_1124 ( .A(_abc_41356_new_n2704_), .B(regfil_2__1_), .Y(_abc_41356_new_n2726_));
AND2X2 AND2X2_1125 ( .A(_abc_41356_new_n2727_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2728_));
AND2X2 AND2X2_1126 ( .A(_abc_41356_new_n2710_), .B(regfil_2__1_), .Y(_abc_41356_new_n2730_));
AND2X2 AND2X2_1127 ( .A(_abc_41356_new_n2731_), .B(_abc_41356_new_n2415_), .Y(_abc_41356_new_n2732_));
AND2X2 AND2X2_1128 ( .A(_abc_41356_new_n2732_), .B(_abc_41356_new_n2729_), .Y(_abc_41356_new_n2733_));
AND2X2 AND2X2_1129 ( .A(_abc_41356_new_n1235_), .B(regfil_4__1_), .Y(_abc_41356_new_n2735_));
AND2X2 AND2X2_113 ( .A(_abc_41356_new_n685_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n686_));
AND2X2 AND2X2_1130 ( .A(_abc_41356_new_n2740_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2741_));
AND2X2 AND2X2_1131 ( .A(_abc_41356_new_n2739_), .B(_abc_41356_new_n2741_), .Y(_abc_41356_new_n2742_));
AND2X2 AND2X2_1132 ( .A(_abc_41356_new_n2393_), .B(rdatahold_2_), .Y(_abc_41356_new_n2743_));
AND2X2 AND2X2_1133 ( .A(_abc_41356_new_n2724_), .B(regfil_2__2_), .Y(_abc_41356_new_n2746_));
AND2X2 AND2X2_1134 ( .A(_abc_41356_new_n2747_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2748_));
AND2X2 AND2X2_1135 ( .A(_abc_41356_new_n2730_), .B(regfil_2__2_), .Y(_abc_41356_new_n2750_));
AND2X2 AND2X2_1136 ( .A(_abc_41356_new_n2751_), .B(_abc_41356_new_n2415_), .Y(_abc_41356_new_n2752_));
AND2X2 AND2X2_1137 ( .A(_abc_41356_new_n2752_), .B(_abc_41356_new_n2749_), .Y(_abc_41356_new_n2753_));
AND2X2 AND2X2_1138 ( .A(_abc_41356_new_n1235_), .B(regfil_4__2_), .Y(_abc_41356_new_n2755_));
AND2X2 AND2X2_1139 ( .A(_abc_41356_new_n2760_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2761_));
AND2X2 AND2X2_114 ( .A(_abc_41356_new_n614_), .B(_abc_41356_new_n545_), .Y(_abc_41356_new_n689_));
AND2X2 AND2X2_1140 ( .A(_abc_41356_new_n2759_), .B(_abc_41356_new_n2761_), .Y(_abc_41356_new_n2762_));
AND2X2 AND2X2_1141 ( .A(_abc_41356_new_n2393_), .B(rdatahold_3_), .Y(_abc_41356_new_n2763_));
AND2X2 AND2X2_1142 ( .A(_abc_41356_new_n2750_), .B(regfil_2__3_), .Y(_abc_41356_new_n2764_));
AND2X2 AND2X2_1143 ( .A(_abc_41356_new_n2766_), .B(_abc_41356_new_n2415_), .Y(_abc_41356_new_n2767_));
AND2X2 AND2X2_1144 ( .A(_abc_41356_new_n2767_), .B(_abc_41356_new_n2765_), .Y(_abc_41356_new_n2768_));
AND2X2 AND2X2_1145 ( .A(_abc_41356_new_n2744_), .B(regfil_2__3_), .Y(_abc_41356_new_n2771_));
AND2X2 AND2X2_1146 ( .A(_abc_41356_new_n2772_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2773_));
AND2X2 AND2X2_1147 ( .A(_abc_41356_new_n2776_), .B(_abc_41356_new_n2422_), .Y(_abc_41356_new_n2777_));
AND2X2 AND2X2_1148 ( .A(_abc_41356_new_n2775_), .B(_abc_41356_new_n2777_), .Y(_abc_41356_new_n2778_));
AND2X2 AND2X2_1149 ( .A(_abc_41356_new_n2782_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2783_));
AND2X2 AND2X2_115 ( .A(_abc_41356_new_n690_), .B(_abc_41356_new_n691_), .Y(_abc_41356_new_n692_));
AND2X2 AND2X2_1150 ( .A(_abc_41356_new_n2781_), .B(_abc_41356_new_n2783_), .Y(_abc_41356_new_n2784_));
AND2X2 AND2X2_1151 ( .A(_abc_41356_new_n2393_), .B(rdatahold_4_), .Y(_abc_41356_new_n2785_));
AND2X2 AND2X2_1152 ( .A(_abc_41356_new_n2764_), .B(regfil_2__4_), .Y(_abc_41356_new_n2786_));
AND2X2 AND2X2_1153 ( .A(_abc_41356_new_n2788_), .B(_abc_41356_new_n2415_), .Y(_abc_41356_new_n2789_));
AND2X2 AND2X2_1154 ( .A(_abc_41356_new_n2789_), .B(_abc_41356_new_n2787_), .Y(_abc_41356_new_n2790_));
AND2X2 AND2X2_1155 ( .A(_abc_41356_new_n2769_), .B(regfil_2__4_), .Y(_abc_41356_new_n2793_));
AND2X2 AND2X2_1156 ( .A(_abc_41356_new_n2794_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2795_));
AND2X2 AND2X2_1157 ( .A(_abc_41356_new_n2798_), .B(_abc_41356_new_n2422_), .Y(_abc_41356_new_n2799_));
AND2X2 AND2X2_1158 ( .A(_abc_41356_new_n2797_), .B(_abc_41356_new_n2799_), .Y(_abc_41356_new_n2800_));
AND2X2 AND2X2_1159 ( .A(_abc_41356_new_n2804_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2805_));
AND2X2 AND2X2_116 ( .A(_abc_41356_new_n604_), .B(_abc_41356_new_n692_), .Y(_abc_41356_new_n693_));
AND2X2 AND2X2_1160 ( .A(_abc_41356_new_n2803_), .B(_abc_41356_new_n2805_), .Y(_abc_41356_new_n2806_));
AND2X2 AND2X2_1161 ( .A(_abc_41356_new_n2393_), .B(rdatahold_5_), .Y(_abc_41356_new_n2807_));
AND2X2 AND2X2_1162 ( .A(_abc_41356_new_n2786_), .B(regfil_2__5_), .Y(_abc_41356_new_n2808_));
AND2X2 AND2X2_1163 ( .A(_abc_41356_new_n2810_), .B(_abc_41356_new_n2415_), .Y(_abc_41356_new_n2811_));
AND2X2 AND2X2_1164 ( .A(_abc_41356_new_n2811_), .B(_abc_41356_new_n2809_), .Y(_abc_41356_new_n2812_));
AND2X2 AND2X2_1165 ( .A(_abc_41356_new_n2791_), .B(regfil_2__5_), .Y(_abc_41356_new_n2815_));
AND2X2 AND2X2_1166 ( .A(_abc_41356_new_n2816_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2817_));
AND2X2 AND2X2_1167 ( .A(_abc_41356_new_n2820_), .B(_abc_41356_new_n2422_), .Y(_abc_41356_new_n2821_));
AND2X2 AND2X2_1168 ( .A(_abc_41356_new_n2819_), .B(_abc_41356_new_n2821_), .Y(_abc_41356_new_n2822_));
AND2X2 AND2X2_1169 ( .A(_abc_41356_new_n2826_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2827_));
AND2X2 AND2X2_117 ( .A(_abc_41356_new_n688_), .B(_abc_41356_new_n693_), .Y(_abc_41356_new_n694_));
AND2X2 AND2X2_1170 ( .A(_abc_41356_new_n2825_), .B(_abc_41356_new_n2827_), .Y(_abc_41356_new_n2828_));
AND2X2 AND2X2_1171 ( .A(_abc_41356_new_n2393_), .B(rdatahold_6_), .Y(_abc_41356_new_n2829_));
AND2X2 AND2X2_1172 ( .A(_abc_41356_new_n2808_), .B(regfil_2__6_), .Y(_abc_41356_new_n2831_));
AND2X2 AND2X2_1173 ( .A(_abc_41356_new_n2832_), .B(_abc_41356_new_n2415_), .Y(_abc_41356_new_n2833_));
AND2X2 AND2X2_1174 ( .A(_abc_41356_new_n2833_), .B(_abc_41356_new_n2830_), .Y(_abc_41356_new_n2834_));
AND2X2 AND2X2_1175 ( .A(_abc_41356_new_n2813_), .B(regfil_2__6_), .Y(_abc_41356_new_n2837_));
AND2X2 AND2X2_1176 ( .A(_abc_41356_new_n2838_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2839_));
AND2X2 AND2X2_1177 ( .A(_abc_41356_new_n2842_), .B(_abc_41356_new_n2422_), .Y(_abc_41356_new_n2843_));
AND2X2 AND2X2_1178 ( .A(_abc_41356_new_n2841_), .B(_abc_41356_new_n2843_), .Y(_abc_41356_new_n2844_));
AND2X2 AND2X2_1179 ( .A(_abc_41356_new_n2847_), .B(_abc_41356_new_n2697_), .Y(_abc_41356_new_n2848_));
AND2X2 AND2X2_118 ( .A(_abc_41356_new_n694_), .B(_abc_41356_new_n673_), .Y(_abc_41356_new_n695_));
AND2X2 AND2X2_1180 ( .A(_abc_41356_new_n2698_), .B(_abc_41356_new_n1996_), .Y(_abc_41356_new_n2849_));
AND2X2 AND2X2_1181 ( .A(_abc_41356_new_n2831_), .B(_abc_41356_new_n2415_), .Y(_abc_41356_new_n2855_));
AND2X2 AND2X2_1182 ( .A(_abc_41356_new_n2836_), .B(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2857_));
AND2X2 AND2X2_1183 ( .A(_abc_41356_new_n2858_), .B(_abc_41356_new_n1996_), .Y(_abc_41356_new_n2859_));
AND2X2 AND2X2_1184 ( .A(_abc_41356_new_n2859_), .B(_abc_41356_new_n2856_), .Y(_abc_41356_new_n2860_));
AND2X2 AND2X2_1185 ( .A(_abc_41356_new_n2863_), .B(regfil_2__7_), .Y(_abc_41356_new_n2864_));
AND2X2 AND2X2_1186 ( .A(_abc_41356_new_n2862_), .B(_abc_41356_new_n2864_), .Y(_abc_41356_new_n2865_));
AND2X2 AND2X2_1187 ( .A(_abc_41356_new_n2866_), .B(_abc_41356_new_n1236_), .Y(_abc_41356_new_n2867_));
AND2X2 AND2X2_1188 ( .A(_abc_41356_new_n1235_), .B(_abc_41356_new_n1961_), .Y(_abc_41356_new_n2868_));
AND2X2 AND2X2_1189 ( .A(_abc_41356_new_n2870_), .B(_abc_41356_new_n2854_), .Y(_abc_41356_new_n2871_));
AND2X2 AND2X2_119 ( .A(_abc_41356_new_n700_), .B(_abc_41356_new_n701_), .Y(_abc_41356_new_n702_));
AND2X2 AND2X2_1190 ( .A(_abc_41356_new_n2871_), .B(_abc_41356_new_n2851_), .Y(_abc_41356_new_n2872_));
AND2X2 AND2X2_1191 ( .A(_abc_41356_new_n615_), .B(opcode_2_), .Y(_abc_41356_new_n2874_));
AND2X2 AND2X2_1192 ( .A(_abc_41356_new_n2875_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n2876_));
AND2X2 AND2X2_1193 ( .A(_abc_41356_new_n523_), .B(_abc_41356_new_n2878_), .Y(_abc_41356_new_n2879_));
AND2X2 AND2X2_1194 ( .A(_abc_41356_new_n2879_), .B(_abc_41356_new_n2877_), .Y(_abc_41356_new_n2880_));
AND2X2 AND2X2_1195 ( .A(_abc_41356_new_n2880_), .B(_abc_41356_new_n2882_), .Y(_abc_41356_new_n2883_));
AND2X2 AND2X2_1196 ( .A(_abc_41356_new_n2884_), .B(alu_sel_0_), .Y(_abc_41356_new_n2885_));
AND2X2 AND2X2_1197 ( .A(_abc_41356_new_n514_), .B(opcode_7_), .Y(_abc_41356_new_n2886_));
AND2X2 AND2X2_1198 ( .A(_abc_41356_new_n677_), .B(opcode_7_), .Y(_abc_41356_new_n2888_));
AND2X2 AND2X2_1199 ( .A(_abc_41356_new_n2889_), .B(_abc_41356_new_n2887_), .Y(_abc_41356_new_n2890_));
AND2X2 AND2X2_12 ( .A(_abc_41356_new_n505_), .B(_abc_41356_new_n520_), .Y(_abc_41356_new_n521_));
AND2X2 AND2X2_120 ( .A(_abc_41356_new_n703_), .B(regfil_7__7_), .Y(_abc_41356_new_n704_));
AND2X2 AND2X2_1200 ( .A(_abc_41356_new_n523_), .B(opcode_3_), .Y(_abc_41356_new_n2892_));
AND2X2 AND2X2_1201 ( .A(_abc_41356_new_n2891_), .B(_abc_41356_new_n2892_), .Y(_abc_41356_new_n2893_));
AND2X2 AND2X2_1202 ( .A(_abc_41356_new_n2896_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2897_));
AND2X2 AND2X2_1203 ( .A(_abc_41356_new_n2897_), .B(_abc_41356_new_n2895_), .Y(_abc_41356_new_n2898_));
AND2X2 AND2X2_1204 ( .A(_abc_41356_new_n2054_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n2900_));
AND2X2 AND2X2_1205 ( .A(_abc_41356_new_n2900_), .B(_abc_41356_new_n2899_), .Y(_abc_41356_new_n2901_));
AND2X2 AND2X2_1206 ( .A(_abc_41356_new_n2886_), .B(opcode_4_), .Y(_abc_41356_new_n2902_));
AND2X2 AND2X2_1207 ( .A(_abc_41356_new_n2904_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2905_));
AND2X2 AND2X2_1208 ( .A(_abc_41356_new_n2906_), .B(alu_sel_1_), .Y(_abc_41356_new_n2907_));
AND2X2 AND2X2_1209 ( .A(_abc_41356_new_n2909_), .B(alu_sel_2_), .Y(_abc_41356_new_n2910_));
AND2X2 AND2X2_121 ( .A(_abc_41356_new_n517_), .B(state_5_), .Y(_abc_41356_new_n706_));
AND2X2 AND2X2_1210 ( .A(_abc_41356_new_n2886_), .B(opcode_5_), .Y(_abc_41356_new_n2911_));
AND2X2 AND2X2_1211 ( .A(_abc_41356_new_n2912_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2913_));
AND2X2 AND2X2_1212 ( .A(_abc_41356_new_n2915_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2916_));
AND2X2 AND2X2_1213 ( .A(_abc_41356_new_n2914_), .B(_abc_41356_new_n2916_), .Y(_abc_41356_new_n2917_));
AND2X2 AND2X2_1214 ( .A(_abc_41356_new_n2891_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2919_));
AND2X2 AND2X2_1215 ( .A(_abc_41356_new_n2922_), .B(_abc_41356_new_n2920_), .Y(_0alucin_0_0_));
AND2X2 AND2X2_1216 ( .A(_abc_41356_new_n713_), .B(_abc_41356_new_n706_), .Y(_abc_41356_new_n2924_));
AND2X2 AND2X2_1217 ( .A(_abc_41356_new_n708_), .B(_abc_41356_new_n506_), .Y(_abc_41356_new_n2926_));
AND2X2 AND2X2_1218 ( .A(_abc_41356_new_n2926_), .B(_abc_41356_new_n706_), .Y(_abc_41356_new_n2927_));
AND2X2 AND2X2_1219 ( .A(_abc_41356_new_n2925_), .B(_abc_41356_new_n2928_), .Y(_abc_41356_new_n2929_));
AND2X2 AND2X2_122 ( .A(_abc_41356_new_n520_), .B(state_1_), .Y(_abc_41356_new_n707_));
AND2X2 AND2X2_1220 ( .A(_abc_41356_new_n2930_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n2931_));
AND2X2 AND2X2_1221 ( .A(_abc_41356_new_n2931_), .B(rdatahold_0_), .Y(_abc_41356_new_n2932_));
AND2X2 AND2X2_1222 ( .A(_abc_41356_new_n2933_), .B(_abc_41356_new_n2020_), .Y(_abc_41356_new_n2934_));
AND2X2 AND2X2_1223 ( .A(_abc_41356_new_n2934_), .B(alu_oprb_0_), .Y(_abc_41356_new_n2935_));
AND2X2 AND2X2_1224 ( .A(_abc_41356_new_n2936_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2937_));
AND2X2 AND2X2_1225 ( .A(_abc_41356_new_n2938_), .B(_abc_41356_new_n2941_), .Y(_abc_41356_new_n2942_));
AND2X2 AND2X2_1226 ( .A(_abc_41356_new_n2939_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2944_));
AND2X2 AND2X2_1227 ( .A(_abc_41356_new_n2945_), .B(alu_oprb_1_), .Y(_abc_41356_new_n2946_));
AND2X2 AND2X2_1228 ( .A(_abc_41356_new_n2931_), .B(rdatahold_1_), .Y(_abc_41356_new_n2947_));
AND2X2 AND2X2_1229 ( .A(_abc_41356_new_n523_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n2948_));
AND2X2 AND2X2_123 ( .A(_abc_41356_new_n503_), .B(_abc_41356_new_n586_), .Y(_abc_41356_new_n708_));
AND2X2 AND2X2_1230 ( .A(_abc_41356_new_n764_), .B(_abc_41356_new_n2948_), .Y(_abc_41356_new_n2949_));
AND2X2 AND2X2_1231 ( .A(_abc_41356_new_n2945_), .B(alu_oprb_2_), .Y(_abc_41356_new_n2952_));
AND2X2 AND2X2_1232 ( .A(_abc_41356_new_n2931_), .B(rdatahold_2_), .Y(_abc_41356_new_n2953_));
AND2X2 AND2X2_1233 ( .A(_abc_41356_new_n817_), .B(_abc_41356_new_n2948_), .Y(_abc_41356_new_n2954_));
AND2X2 AND2X2_1234 ( .A(_abc_41356_new_n878_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n2957_));
AND2X2 AND2X2_1235 ( .A(_abc_41356_new_n2939_), .B(alu_oprb_3_), .Y(_abc_41356_new_n2958_));
AND2X2 AND2X2_1236 ( .A(_abc_41356_new_n2959_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2960_));
AND2X2 AND2X2_1237 ( .A(_abc_41356_new_n2934_), .B(alu_oprb_3_), .Y(_abc_41356_new_n2961_));
AND2X2 AND2X2_1238 ( .A(_abc_41356_new_n2931_), .B(rdatahold_3_), .Y(_abc_41356_new_n2962_));
AND2X2 AND2X2_1239 ( .A(_abc_41356_new_n2945_), .B(alu_oprb_4_), .Y(_abc_41356_new_n2965_));
AND2X2 AND2X2_124 ( .A(_abc_41356_new_n708_), .B(_abc_41356_new_n707_), .Y(_abc_41356_new_n709_));
AND2X2 AND2X2_1240 ( .A(_abc_41356_new_n2931_), .B(rdatahold_4_), .Y(_abc_41356_new_n2966_));
AND2X2 AND2X2_1241 ( .A(_abc_41356_new_n945_), .B(_abc_41356_new_n2948_), .Y(_abc_41356_new_n2967_));
AND2X2 AND2X2_1242 ( .A(_abc_41356_new_n2945_), .B(alu_oprb_5_), .Y(_abc_41356_new_n2970_));
AND2X2 AND2X2_1243 ( .A(_abc_41356_new_n2931_), .B(rdatahold_5_), .Y(_abc_41356_new_n2971_));
AND2X2 AND2X2_1244 ( .A(_abc_41356_new_n1012_), .B(_abc_41356_new_n2948_), .Y(_abc_41356_new_n2972_));
AND2X2 AND2X2_1245 ( .A(_abc_41356_new_n1069_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n2975_));
AND2X2 AND2X2_1246 ( .A(_abc_41356_new_n2939_), .B(alu_oprb_6_), .Y(_abc_41356_new_n2976_));
AND2X2 AND2X2_1247 ( .A(_abc_41356_new_n2977_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2978_));
AND2X2 AND2X2_1248 ( .A(_abc_41356_new_n2931_), .B(rdatahold_6_), .Y(_abc_41356_new_n2979_));
AND2X2 AND2X2_1249 ( .A(_abc_41356_new_n2934_), .B(alu_oprb_6_), .Y(_abc_41356_new_n2980_));
AND2X2 AND2X2_125 ( .A(_abc_41356_new_n709_), .B(_abc_41356_new_n706_), .Y(_abc_41356_new_n710_));
AND2X2 AND2X2_1250 ( .A(_abc_41356_new_n2945_), .B(alu_oprb_7_), .Y(_abc_41356_new_n2983_));
AND2X2 AND2X2_1251 ( .A(_abc_41356_new_n2930_), .B(_abc_41356_new_n1164_), .Y(_abc_41356_new_n2984_));
AND2X2 AND2X2_1252 ( .A(_abc_41356_new_n1161_), .B(_abc_41356_new_n2948_), .Y(_abc_41356_new_n2985_));
AND2X2 AND2X2_1253 ( .A(_abc_41356_new_n2891_), .B(regfil_7__0_), .Y(_abc_41356_new_n2988_));
AND2X2 AND2X2_1254 ( .A(opcode_4_), .B(opcode_3_), .Y(_abc_41356_new_n2989_));
AND2X2 AND2X2_1255 ( .A(_abc_41356_new_n2989_), .B(regfil_7__0_), .Y(_abc_41356_new_n2990_));
AND2X2 AND2X2_1256 ( .A(_abc_41356_new_n534_), .B(opcode_3_), .Y(_abc_41356_new_n2992_));
AND2X2 AND2X2_1257 ( .A(_abc_41356_new_n2992_), .B(regfil_5__0_), .Y(_abc_41356_new_n2993_));
AND2X2 AND2X2_1258 ( .A(_abc_41356_new_n534_), .B(_abc_41356_new_n545_), .Y(_abc_41356_new_n2994_));
AND2X2 AND2X2_1259 ( .A(_abc_41356_new_n2994_), .B(regfil_4__0_), .Y(_abc_41356_new_n2995_));
AND2X2 AND2X2_126 ( .A(_abc_41356_new_n710_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n711_));
AND2X2 AND2X2_1260 ( .A(_abc_41356_new_n545_), .B(opcode_4_), .Y(_abc_41356_new_n2997_));
AND2X2 AND2X2_1261 ( .A(_abc_41356_new_n2997_), .B(regfil_6__0_), .Y(_abc_41356_new_n2998_));
AND2X2 AND2X2_1262 ( .A(_abc_41356_new_n516_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n3001_));
AND2X2 AND2X2_1263 ( .A(_abc_41356_new_n2992_), .B(regfil_1__0_), .Y(_abc_41356_new_n3002_));
AND2X2 AND2X2_1264 ( .A(_abc_41356_new_n2989_), .B(regfil_3__0_), .Y(_abc_41356_new_n3004_));
AND2X2 AND2X2_1265 ( .A(_abc_41356_new_n2994_), .B(regfil_0__0_), .Y(_abc_41356_new_n3005_));
AND2X2 AND2X2_1266 ( .A(_abc_41356_new_n2997_), .B(regfil_2__0_), .Y(_abc_41356_new_n3006_));
AND2X2 AND2X2_1267 ( .A(_abc_41356_new_n3009_), .B(_abc_41356_new_n3001_), .Y(_abc_41356_new_n3010_));
AND2X2 AND2X2_1268 ( .A(_abc_41356_new_n3010_), .B(_abc_41356_new_n3000_), .Y(_abc_41356_new_n3011_));
AND2X2 AND2X2_1269 ( .A(_abc_41356_new_n3012_), .B(_abc_41356_new_n2879_), .Y(_abc_41356_new_n3013_));
AND2X2 AND2X2_127 ( .A(_abc_41356_new_n711_), .B(_abc_41356_new_n705_), .Y(_abc_41356_new_n712_));
AND2X2 AND2X2_1270 ( .A(_abc_41356_new_n507_), .B(_abc_41356_new_n706_), .Y(_abc_41356_new_n3014_));
AND2X2 AND2X2_1271 ( .A(_abc_41356_new_n3014_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3015_));
AND2X2 AND2X2_1272 ( .A(_abc_41356_new_n3015_), .B(rdatahold_0_), .Y(_abc_41356_new_n3016_));
AND2X2 AND2X2_1273 ( .A(_abc_41356_new_n3017_), .B(_abc_41356_new_n2020_), .Y(_abc_41356_new_n3018_));
AND2X2 AND2X2_1274 ( .A(_abc_41356_new_n2939_), .B(_abc_41356_new_n2889_), .Y(_abc_41356_new_n3019_));
AND2X2 AND2X2_1275 ( .A(_abc_41356_new_n3019_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n3020_));
AND2X2 AND2X2_1276 ( .A(_abc_41356_new_n3021_), .B(alu_opra_0_), .Y(_abc_41356_new_n3022_));
AND2X2 AND2X2_1277 ( .A(_abc_41356_new_n2891_), .B(regfil_7__1_), .Y(_abc_41356_new_n3025_));
AND2X2 AND2X2_1278 ( .A(_abc_41356_new_n2989_), .B(regfil_7__1_), .Y(_abc_41356_new_n3026_));
AND2X2 AND2X2_1279 ( .A(_abc_41356_new_n2992_), .B(regfil_5__1_), .Y(_abc_41356_new_n3028_));
AND2X2 AND2X2_128 ( .A(_abc_41356_new_n504_), .B(_abc_41356_new_n707_), .Y(_abc_41356_new_n713_));
AND2X2 AND2X2_1280 ( .A(_abc_41356_new_n2994_), .B(regfil_4__1_), .Y(_abc_41356_new_n3029_));
AND2X2 AND2X2_1281 ( .A(_abc_41356_new_n2997_), .B(regfil_6__1_), .Y(_abc_41356_new_n3031_));
AND2X2 AND2X2_1282 ( .A(_abc_41356_new_n2992_), .B(regfil_1__1_), .Y(_abc_41356_new_n3034_));
AND2X2 AND2X2_1283 ( .A(_abc_41356_new_n2989_), .B(regfil_3__1_), .Y(_abc_41356_new_n3036_));
AND2X2 AND2X2_1284 ( .A(_abc_41356_new_n2994_), .B(regfil_0__1_), .Y(_abc_41356_new_n3037_));
AND2X2 AND2X2_1285 ( .A(_abc_41356_new_n2997_), .B(regfil_2__1_), .Y(_abc_41356_new_n3038_));
AND2X2 AND2X2_1286 ( .A(_abc_41356_new_n3041_), .B(_abc_41356_new_n3001_), .Y(_abc_41356_new_n3042_));
AND2X2 AND2X2_1287 ( .A(_abc_41356_new_n3042_), .B(_abc_41356_new_n3033_), .Y(_abc_41356_new_n3043_));
AND2X2 AND2X2_1288 ( .A(_abc_41356_new_n3044_), .B(_abc_41356_new_n2879_), .Y(_abc_41356_new_n3045_));
AND2X2 AND2X2_1289 ( .A(_abc_41356_new_n3015_), .B(rdatahold_1_), .Y(_abc_41356_new_n3046_));
AND2X2 AND2X2_129 ( .A(_abc_41356_new_n519_), .B(_abc_41356_new_n713_), .Y(_abc_41356_new_n714_));
AND2X2 AND2X2_1290 ( .A(_abc_41356_new_n3021_), .B(alu_opra_1_), .Y(_abc_41356_new_n3047_));
AND2X2 AND2X2_1291 ( .A(_abc_41356_new_n2891_), .B(regfil_7__2_), .Y(_abc_41356_new_n3050_));
AND2X2 AND2X2_1292 ( .A(_abc_41356_new_n2989_), .B(regfil_7__2_), .Y(_abc_41356_new_n3051_));
AND2X2 AND2X2_1293 ( .A(_abc_41356_new_n2992_), .B(regfil_5__2_), .Y(_abc_41356_new_n3053_));
AND2X2 AND2X2_1294 ( .A(_abc_41356_new_n2994_), .B(regfil_4__2_), .Y(_abc_41356_new_n3054_));
AND2X2 AND2X2_1295 ( .A(_abc_41356_new_n2997_), .B(regfil_6__2_), .Y(_abc_41356_new_n3056_));
AND2X2 AND2X2_1296 ( .A(_abc_41356_new_n2992_), .B(regfil_1__2_), .Y(_abc_41356_new_n3059_));
AND2X2 AND2X2_1297 ( .A(_abc_41356_new_n2989_), .B(regfil_3__2_), .Y(_abc_41356_new_n3061_));
AND2X2 AND2X2_1298 ( .A(_abc_41356_new_n2994_), .B(regfil_0__2_), .Y(_abc_41356_new_n3062_));
AND2X2 AND2X2_1299 ( .A(_abc_41356_new_n2997_), .B(regfil_2__2_), .Y(_abc_41356_new_n3063_));
AND2X2 AND2X2_13 ( .A(_abc_41356_new_n521_), .B(_abc_41356_new_n504_), .Y(_abc_41356_new_n522_));
AND2X2 AND2X2_130 ( .A(_abc_41356_new_n588_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n715_));
AND2X2 AND2X2_1300 ( .A(_abc_41356_new_n3066_), .B(_abc_41356_new_n3001_), .Y(_abc_41356_new_n3067_));
AND2X2 AND2X2_1301 ( .A(_abc_41356_new_n3067_), .B(_abc_41356_new_n3058_), .Y(_abc_41356_new_n3068_));
AND2X2 AND2X2_1302 ( .A(_abc_41356_new_n3069_), .B(_abc_41356_new_n2879_), .Y(_abc_41356_new_n3070_));
AND2X2 AND2X2_1303 ( .A(_abc_41356_new_n3015_), .B(rdatahold_2_), .Y(_abc_41356_new_n3071_));
AND2X2 AND2X2_1304 ( .A(_abc_41356_new_n3021_), .B(alu_opra_2_), .Y(_abc_41356_new_n3072_));
AND2X2 AND2X2_1305 ( .A(_abc_41356_new_n2891_), .B(regfil_7__3_), .Y(_abc_41356_new_n3075_));
AND2X2 AND2X2_1306 ( .A(_abc_41356_new_n2989_), .B(regfil_7__3_), .Y(_abc_41356_new_n3076_));
AND2X2 AND2X2_1307 ( .A(_abc_41356_new_n2992_), .B(regfil_5__3_), .Y(_abc_41356_new_n3078_));
AND2X2 AND2X2_1308 ( .A(_abc_41356_new_n2994_), .B(regfil_4__3_), .Y(_abc_41356_new_n3079_));
AND2X2 AND2X2_1309 ( .A(_abc_41356_new_n2997_), .B(regfil_6__3_), .Y(_abc_41356_new_n3081_));
AND2X2 AND2X2_131 ( .A(_abc_41356_new_n509_), .B(_abc_41356_new_n716_), .Y(_abc_41356_new_n717_));
AND2X2 AND2X2_1310 ( .A(_abc_41356_new_n2992_), .B(regfil_1__3_), .Y(_abc_41356_new_n3084_));
AND2X2 AND2X2_1311 ( .A(_abc_41356_new_n2989_), .B(regfil_3__3_), .Y(_abc_41356_new_n3086_));
AND2X2 AND2X2_1312 ( .A(_abc_41356_new_n2994_), .B(regfil_0__3_), .Y(_abc_41356_new_n3087_));
AND2X2 AND2X2_1313 ( .A(_abc_41356_new_n2997_), .B(regfil_2__3_), .Y(_abc_41356_new_n3088_));
AND2X2 AND2X2_1314 ( .A(_abc_41356_new_n3091_), .B(_abc_41356_new_n3001_), .Y(_abc_41356_new_n3092_));
AND2X2 AND2X2_1315 ( .A(_abc_41356_new_n3092_), .B(_abc_41356_new_n3083_), .Y(_abc_41356_new_n3093_));
AND2X2 AND2X2_1316 ( .A(_abc_41356_new_n3094_), .B(_abc_41356_new_n2879_), .Y(_abc_41356_new_n3095_));
AND2X2 AND2X2_1317 ( .A(_abc_41356_new_n3015_), .B(rdatahold_3_), .Y(_abc_41356_new_n3096_));
AND2X2 AND2X2_1318 ( .A(_abc_41356_new_n3021_), .B(alu_opra_3_), .Y(_abc_41356_new_n3097_));
AND2X2 AND2X2_1319 ( .A(_abc_41356_new_n2891_), .B(regfil_7__4_), .Y(_abc_41356_new_n3100_));
AND2X2 AND2X2_132 ( .A(_abc_41356_new_n715_), .B(_abc_41356_new_n717_), .Y(_abc_41356_new_n718_));
AND2X2 AND2X2_1320 ( .A(_abc_41356_new_n2989_), .B(regfil_7__4_), .Y(_abc_41356_new_n3101_));
AND2X2 AND2X2_1321 ( .A(_abc_41356_new_n2992_), .B(regfil_5__4_), .Y(_abc_41356_new_n3103_));
AND2X2 AND2X2_1322 ( .A(_abc_41356_new_n2994_), .B(regfil_4__4_), .Y(_abc_41356_new_n3104_));
AND2X2 AND2X2_1323 ( .A(_abc_41356_new_n2997_), .B(regfil_6__4_), .Y(_abc_41356_new_n3106_));
AND2X2 AND2X2_1324 ( .A(_abc_41356_new_n2992_), .B(regfil_1__4_), .Y(_abc_41356_new_n3109_));
AND2X2 AND2X2_1325 ( .A(_abc_41356_new_n2989_), .B(regfil_3__4_), .Y(_abc_41356_new_n3111_));
AND2X2 AND2X2_1326 ( .A(_abc_41356_new_n2994_), .B(regfil_0__4_), .Y(_abc_41356_new_n3112_));
AND2X2 AND2X2_1327 ( .A(_abc_41356_new_n2997_), .B(regfil_2__4_), .Y(_abc_41356_new_n3113_));
AND2X2 AND2X2_1328 ( .A(_abc_41356_new_n3116_), .B(_abc_41356_new_n3001_), .Y(_abc_41356_new_n3117_));
AND2X2 AND2X2_1329 ( .A(_abc_41356_new_n3117_), .B(_abc_41356_new_n3108_), .Y(_abc_41356_new_n3118_));
AND2X2 AND2X2_133 ( .A(_abc_41356_new_n725_), .B(_abc_41356_new_n724_), .Y(_abc_41356_new_n726_));
AND2X2 AND2X2_1330 ( .A(_abc_41356_new_n3119_), .B(_abc_41356_new_n2879_), .Y(_abc_41356_new_n3120_));
AND2X2 AND2X2_1331 ( .A(_abc_41356_new_n3015_), .B(rdatahold_4_), .Y(_abc_41356_new_n3121_));
AND2X2 AND2X2_1332 ( .A(_abc_41356_new_n3021_), .B(alu_opra_4_), .Y(_abc_41356_new_n3122_));
AND2X2 AND2X2_1333 ( .A(_abc_41356_new_n2891_), .B(regfil_7__5_), .Y(_abc_41356_new_n3125_));
AND2X2 AND2X2_1334 ( .A(_abc_41356_new_n2992_), .B(regfil_1__5_), .Y(_abc_41356_new_n3126_));
AND2X2 AND2X2_1335 ( .A(_abc_41356_new_n2989_), .B(regfil_3__5_), .Y(_abc_41356_new_n3128_));
AND2X2 AND2X2_1336 ( .A(_abc_41356_new_n2994_), .B(regfil_0__5_), .Y(_abc_41356_new_n3129_));
AND2X2 AND2X2_1337 ( .A(_abc_41356_new_n2997_), .B(regfil_2__5_), .Y(_abc_41356_new_n3130_));
AND2X2 AND2X2_1338 ( .A(_abc_41356_new_n2989_), .B(regfil_7__5_), .Y(_abc_41356_new_n3134_));
AND2X2 AND2X2_1339 ( .A(_abc_41356_new_n2992_), .B(regfil_5__5_), .Y(_abc_41356_new_n3136_));
AND2X2 AND2X2_134 ( .A(_abc_41356_new_n697_), .B(_abc_41356_new_n726_), .Y(_abc_41356_new_n727_));
AND2X2 AND2X2_1340 ( .A(_abc_41356_new_n2994_), .B(regfil_4__5_), .Y(_abc_41356_new_n3137_));
AND2X2 AND2X2_1341 ( .A(_abc_41356_new_n2997_), .B(regfil_6__5_), .Y(_abc_41356_new_n3139_));
AND2X2 AND2X2_1342 ( .A(_abc_41356_new_n3141_), .B(_abc_41356_new_n3001_), .Y(_abc_41356_new_n3142_));
AND2X2 AND2X2_1343 ( .A(_abc_41356_new_n3142_), .B(_abc_41356_new_n3133_), .Y(_abc_41356_new_n3143_));
AND2X2 AND2X2_1344 ( .A(_abc_41356_new_n3144_), .B(_abc_41356_new_n2879_), .Y(_abc_41356_new_n3145_));
AND2X2 AND2X2_1345 ( .A(_abc_41356_new_n3015_), .B(rdatahold_5_), .Y(_abc_41356_new_n3146_));
AND2X2 AND2X2_1346 ( .A(_abc_41356_new_n3021_), .B(alu_opra_5_), .Y(_abc_41356_new_n3147_));
AND2X2 AND2X2_1347 ( .A(_abc_41356_new_n2891_), .B(regfil_7__6_), .Y(_abc_41356_new_n3150_));
AND2X2 AND2X2_1348 ( .A(_abc_41356_new_n2992_), .B(regfil_1__6_), .Y(_abc_41356_new_n3151_));
AND2X2 AND2X2_1349 ( .A(_abc_41356_new_n2989_), .B(regfil_3__6_), .Y(_abc_41356_new_n3153_));
AND2X2 AND2X2_135 ( .A(_abc_41356_new_n712_), .B(regfil_7__0_), .Y(_abc_41356_new_n728_));
AND2X2 AND2X2_1350 ( .A(_abc_41356_new_n2994_), .B(regfil_0__6_), .Y(_abc_41356_new_n3154_));
AND2X2 AND2X2_1351 ( .A(_abc_41356_new_n2997_), .B(regfil_2__6_), .Y(_abc_41356_new_n3155_));
AND2X2 AND2X2_1352 ( .A(_abc_41356_new_n2989_), .B(regfil_7__6_), .Y(_abc_41356_new_n3159_));
AND2X2 AND2X2_1353 ( .A(_abc_41356_new_n2992_), .B(regfil_5__6_), .Y(_abc_41356_new_n3161_));
AND2X2 AND2X2_1354 ( .A(_abc_41356_new_n2994_), .B(regfil_4__6_), .Y(_abc_41356_new_n3162_));
AND2X2 AND2X2_1355 ( .A(_abc_41356_new_n2997_), .B(regfil_6__6_), .Y(_abc_41356_new_n3164_));
AND2X2 AND2X2_1356 ( .A(_abc_41356_new_n3166_), .B(_abc_41356_new_n3001_), .Y(_abc_41356_new_n3167_));
AND2X2 AND2X2_1357 ( .A(_abc_41356_new_n3167_), .B(_abc_41356_new_n3158_), .Y(_abc_41356_new_n3168_));
AND2X2 AND2X2_1358 ( .A(_abc_41356_new_n3169_), .B(_abc_41356_new_n2879_), .Y(_abc_41356_new_n3170_));
AND2X2 AND2X2_1359 ( .A(_abc_41356_new_n3015_), .B(rdatahold_6_), .Y(_abc_41356_new_n3171_));
AND2X2 AND2X2_136 ( .A(_abc_41356_new_n714_), .B(alu_res_0_), .Y(_abc_41356_new_n729_));
AND2X2 AND2X2_1360 ( .A(_abc_41356_new_n3021_), .B(alu_opra_6_), .Y(_abc_41356_new_n3172_));
AND2X2 AND2X2_1361 ( .A(_abc_41356_new_n2891_), .B(regfil_7__7_), .Y(_abc_41356_new_n3175_));
AND2X2 AND2X2_1362 ( .A(_abc_41356_new_n2994_), .B(regfil_0__7_), .Y(_abc_41356_new_n3176_));
AND2X2 AND2X2_1363 ( .A(_abc_41356_new_n2992_), .B(regfil_1__7_), .Y(_abc_41356_new_n3177_));
AND2X2 AND2X2_1364 ( .A(_abc_41356_new_n2989_), .B(regfil_3__7_), .Y(_abc_41356_new_n3179_));
AND2X2 AND2X2_1365 ( .A(_abc_41356_new_n2997_), .B(regfil_2__7_), .Y(_abc_41356_new_n3180_));
AND2X2 AND2X2_1366 ( .A(_abc_41356_new_n3182_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3183_));
AND2X2 AND2X2_1367 ( .A(_abc_41356_new_n2992_), .B(regfil_5__7_), .Y(_abc_41356_new_n3184_));
AND2X2 AND2X2_1368 ( .A(_abc_41356_new_n2989_), .B(regfil_7__7_), .Y(_abc_41356_new_n3185_));
AND2X2 AND2X2_1369 ( .A(_abc_41356_new_n2994_), .B(regfil_4__7_), .Y(_abc_41356_new_n3187_));
AND2X2 AND2X2_137 ( .A(_abc_41356_new_n718_), .B(\data[0] ), .Y(_abc_41356_new_n730_));
AND2X2 AND2X2_1370 ( .A(_abc_41356_new_n2997_), .B(regfil_6__7_), .Y(_abc_41356_new_n3188_));
AND2X2 AND2X2_1371 ( .A(_abc_41356_new_n3190_), .B(opcode_5_), .Y(_abc_41356_new_n3191_));
AND2X2 AND2X2_1372 ( .A(_abc_41356_new_n3192_), .B(_abc_41356_new_n3001_), .Y(_abc_41356_new_n3193_));
AND2X2 AND2X2_1373 ( .A(_abc_41356_new_n3194_), .B(_abc_41356_new_n2879_), .Y(_abc_41356_new_n3195_));
AND2X2 AND2X2_1374 ( .A(_abc_41356_new_n3014_), .B(_abc_41356_new_n1164_), .Y(_abc_41356_new_n3196_));
AND2X2 AND2X2_1375 ( .A(_abc_41356_new_n3021_), .B(alu_opra_7_), .Y(_abc_41356_new_n3197_));
AND2X2 AND2X2_1376 ( .A(ei), .B(intr), .Y(_abc_41356_new_n3202_));
AND2X2 AND2X2_1377 ( .A(_abc_41356_new_n2926_), .B(_abc_41356_new_n518_), .Y(_abc_41356_new_n3205_));
AND2X2 AND2X2_1378 ( .A(_abc_41356_new_n3206_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3207_));
AND2X2 AND2X2_1379 ( .A(_abc_41356_new_n3207_), .B(_abc_41356_new_n3204_), .Y(_0intcyc_0_0_));
AND2X2 AND2X2_138 ( .A(_abc_41356_new_n738_), .B(regfil_0__1_), .Y(_abc_41356_new_n739_));
AND2X2 AND2X2_1380 ( .A(_abc_41356_new_n611_), .B(_abc_41356_new_n517_), .Y(_abc_41356_new_n3210_));
AND2X2 AND2X2_1381 ( .A(_abc_41356_new_n713_), .B(_abc_41356_new_n518_), .Y(_abc_41356_new_n3211_));
AND2X2 AND2X2_1382 ( .A(_abc_41356_new_n3213_), .B(_abc_41356_new_n3209_), .Y(_abc_41356_new_n3214_));
AND2X2 AND2X2_1383 ( .A(_abc_41356_new_n3215_), .B(parity), .Y(_abc_41356_new_n3216_));
AND2X2 AND2X2_1384 ( .A(_abc_41356_new_n3212_), .B(alu_parity), .Y(_abc_41356_new_n3217_));
AND2X2 AND2X2_1385 ( .A(_abc_41356_new_n510_), .B(rdatahold2_2_), .Y(_abc_41356_new_n3218_));
AND2X2 AND2X2_1386 ( .A(_abc_41356_new_n3219_), .B(parity), .Y(_abc_41356_new_n3220_));
AND2X2 AND2X2_1387 ( .A(_abc_41356_new_n3221_), .B(_abc_41356_new_n508_), .Y(_abc_41356_new_n3222_));
AND2X2 AND2X2_1388 ( .A(_abc_41356_new_n3223_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3224_));
AND2X2 AND2X2_1389 ( .A(_abc_41356_new_n3215_), .B(zero), .Y(_abc_41356_new_n3226_));
AND2X2 AND2X2_139 ( .A(_abc_41356_new_n740_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n741_));
AND2X2 AND2X2_1390 ( .A(_abc_41356_new_n3212_), .B(alu_zout), .Y(_abc_41356_new_n3227_));
AND2X2 AND2X2_1391 ( .A(_abc_41356_new_n510_), .B(rdatahold2_6_), .Y(_abc_41356_new_n3228_));
AND2X2 AND2X2_1392 ( .A(_abc_41356_new_n3219_), .B(zero), .Y(_abc_41356_new_n3229_));
AND2X2 AND2X2_1393 ( .A(_abc_41356_new_n3230_), .B(_abc_41356_new_n508_), .Y(_abc_41356_new_n3231_));
AND2X2 AND2X2_1394 ( .A(_abc_41356_new_n3232_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3233_));
AND2X2 AND2X2_1395 ( .A(_abc_41356_new_n3215_), .B(sign), .Y(_abc_41356_new_n3235_));
AND2X2 AND2X2_1396 ( .A(_abc_41356_new_n510_), .B(_abc_41356_new_n3236_), .Y(_abc_41356_new_n3237_));
AND2X2 AND2X2_1397 ( .A(_abc_41356_new_n3238_), .B(_abc_41356_new_n3239_), .Y(_abc_41356_new_n3240_));
AND2X2 AND2X2_1398 ( .A(_abc_41356_new_n508_), .B(_abc_41356_new_n3240_), .Y(_abc_41356_new_n3241_));
AND2X2 AND2X2_1399 ( .A(_abc_41356_new_n3210_), .B(alu_res_7_), .Y(_abc_41356_new_n3242_));
AND2X2 AND2X2_14 ( .A(_abc_41356_new_n519_), .B(_abc_41356_new_n522_), .Y(_abc_41356_new_n523_));
AND2X2 AND2X2_140 ( .A(_abc_41356_new_n582_), .B(regfil_0__1_), .Y(_abc_41356_new_n743_));
AND2X2 AND2X2_1400 ( .A(_abc_41356_new_n3211_), .B(alu_sout), .Y(_abc_41356_new_n3243_));
AND2X2 AND2X2_1401 ( .A(_abc_41356_new_n3245_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3246_));
AND2X2 AND2X2_1402 ( .A(_abc_41356_new_n1107_), .B(regfil_7__7_), .Y(_abc_41356_new_n3249_));
AND2X2 AND2X2_1403 ( .A(_abc_41356_new_n3251_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3252_));
AND2X2 AND2X2_1404 ( .A(_abc_41356_new_n3250_), .B(_abc_41356_new_n3252_), .Y(_abc_41356_new_n3253_));
AND2X2 AND2X2_1405 ( .A(_abc_41356_new_n3219_), .B(auxcar), .Y(_abc_41356_new_n3254_));
AND2X2 AND2X2_1406 ( .A(_abc_41356_new_n510_), .B(rdatahold2_4_), .Y(_abc_41356_new_n3255_));
AND2X2 AND2X2_1407 ( .A(_abc_41356_new_n3256_), .B(_abc_41356_new_n508_), .Y(_abc_41356_new_n3257_));
AND2X2 AND2X2_1408 ( .A(_abc_41356_new_n3212_), .B(1'h0), .Y(_abc_41356_new_n3258_));
AND2X2 AND2X2_1409 ( .A(_abc_41356_new_n3260_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3261_));
AND2X2 AND2X2_141 ( .A(_abc_41356_new_n744_), .B(_abc_41356_new_n581_), .Y(_abc_41356_new_n745_));
AND2X2 AND2X2_1410 ( .A(_abc_41356_new_n2020_), .B(auxcar), .Y(_abc_41356_new_n3262_));
AND2X2 AND2X2_1411 ( .A(_abc_41356_new_n3215_), .B(_abc_41356_new_n3262_), .Y(_abc_41356_new_n3263_));
AND2X2 AND2X2_1412 ( .A(_abc_41356_new_n3209_), .B(_abc_41356_new_n3265_), .Y(_abc_41356_new_n3266_));
AND2X2 AND2X2_1413 ( .A(_abc_41356_new_n975_), .B(carry), .Y(_abc_41356_new_n3269_));
AND2X2 AND2X2_1414 ( .A(_abc_41356_new_n3269_), .B(_abc_41356_new_n3268_), .Y(_abc_41356_new_n3270_));
AND2X2 AND2X2_1415 ( .A(_abc_41356_new_n3267_), .B(_abc_41356_new_n3270_), .Y(_abc_41356_new_n3271_));
AND2X2 AND2X2_1416 ( .A(_abc_41356_new_n1985_), .B(_abc_41356_new_n1983_), .Y(_abc_41356_new_n3272_));
AND2X2 AND2X2_1417 ( .A(_abc_41356_new_n3273_), .B(_abc_41356_new_n1481_), .Y(_abc_41356_new_n3274_));
AND2X2 AND2X2_1418 ( .A(_abc_41356_new_n1414_), .B(_abc_41356_new_n3276_), .Y(_abc_41356_new_n3277_));
AND2X2 AND2X2_1419 ( .A(_abc_41356_new_n3275_), .B(_abc_41356_new_n3277_), .Y(_abc_41356_new_n3278_));
AND2X2 AND2X2_142 ( .A(_abc_41356_new_n745_), .B(_abc_41356_new_n742_), .Y(_abc_41356_new_n746_));
AND2X2 AND2X2_1420 ( .A(_abc_41356_new_n528_), .B(_abc_41356_new_n681_), .Y(_abc_41356_new_n3280_));
AND2X2 AND2X2_1421 ( .A(_abc_41356_new_n3280_), .B(_abc_41356_new_n3279_), .Y(_abc_41356_new_n3281_));
AND2X2 AND2X2_1422 ( .A(_abc_41356_new_n1417_), .B(regfil_4__7_), .Y(_abc_41356_new_n3282_));
AND2X2 AND2X2_1423 ( .A(_abc_41356_new_n529_), .B(regfil_7__0_), .Y(_abc_41356_new_n3284_));
AND2X2 AND2X2_1424 ( .A(_abc_41356_new_n554_), .B(regfil_7__7_), .Y(_abc_41356_new_n3285_));
AND2X2 AND2X2_1425 ( .A(_abc_41356_new_n1286_), .B(_abc_41356_new_n3291_), .Y(_abc_41356_new_n3292_));
AND2X2 AND2X2_1426 ( .A(_abc_41356_new_n3290_), .B(_abc_41356_new_n3292_), .Y(_abc_41356_new_n3293_));
AND2X2 AND2X2_1427 ( .A(_abc_41356_new_n3296_), .B(_abc_41356_new_n3295_), .Y(_abc_41356_new_n3297_));
AND2X2 AND2X2_1428 ( .A(_abc_41356_new_n3297_), .B(carry), .Y(_abc_41356_new_n3298_));
AND2X2 AND2X2_1429 ( .A(_abc_41356_new_n547_), .B(_abc_41356_new_n681_), .Y(_abc_41356_new_n3299_));
AND2X2 AND2X2_143 ( .A(_abc_41356_new_n642_), .B(rdatahold_1_), .Y(_abc_41356_new_n747_));
AND2X2 AND2X2_1430 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n3303_), .Y(_abc_41356_new_n3304_));
AND2X2 AND2X2_1431 ( .A(_abc_41356_new_n3302_), .B(_abc_41356_new_n3304_), .Y(_abc_41356_new_n3305_));
AND2X2 AND2X2_1432 ( .A(_abc_41356_new_n3211_), .B(alu_cout), .Y(_abc_41356_new_n3306_));
AND2X2 AND2X2_1433 ( .A(_abc_41356_new_n710_), .B(_abc_41356_new_n704_), .Y(_abc_41356_new_n3307_));
AND2X2 AND2X2_1434 ( .A(_abc_41356_new_n3219_), .B(carry), .Y(_abc_41356_new_n3309_));
AND2X2 AND2X2_1435 ( .A(_abc_41356_new_n510_), .B(rdatahold2_0_), .Y(_abc_41356_new_n3310_));
AND2X2 AND2X2_1436 ( .A(_abc_41356_new_n3311_), .B(_abc_41356_new_n508_), .Y(_abc_41356_new_n3312_));
AND2X2 AND2X2_1437 ( .A(_abc_41356_new_n3314_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3315_));
AND2X2 AND2X2_1438 ( .A(_abc_41356_new_n708_), .B(_abc_41356_new_n610_), .Y(_abc_41356_new_n3317_));
AND2X2 AND2X2_1439 ( .A(_abc_41356_new_n3317_), .B(_abc_41356_new_n518_), .Y(_abc_41356_new_n3318_));
AND2X2 AND2X2_144 ( .A(_abc_41356_new_n619_), .B(regfil_4__1_), .Y(_abc_41356_new_n748_));
AND2X2 AND2X2_1440 ( .A(_abc_41356_new_n3318_), .B(_abc_41356_new_n717_), .Y(_abc_41356_new_n3319_));
AND2X2 AND2X2_1441 ( .A(_abc_41356_new_n3322_), .B(_abc_41356_new_n3320_), .Y(_0opcode_7_0__0_));
AND2X2 AND2X2_1442 ( .A(_abc_41356_new_n3319_), .B(\data[1] ), .Y(_abc_41356_new_n3324_));
AND2X2 AND2X2_1443 ( .A(_abc_41356_new_n3321_), .B(opcode_1_), .Y(_abc_41356_new_n3325_));
AND2X2 AND2X2_1444 ( .A(_abc_41356_new_n3328_), .B(_abc_41356_new_n3327_), .Y(_0opcode_7_0__2_));
AND2X2 AND2X2_1445 ( .A(_abc_41356_new_n3319_), .B(\data[3] ), .Y(_abc_41356_new_n3330_));
AND2X2 AND2X2_1446 ( .A(_abc_41356_new_n3321_), .B(opcode_3_), .Y(_abc_41356_new_n3331_));
AND2X2 AND2X2_1447 ( .A(_abc_41356_new_n3334_), .B(_abc_41356_new_n3333_), .Y(_0opcode_7_0__4_));
AND2X2 AND2X2_1448 ( .A(_abc_41356_new_n3337_), .B(_abc_41356_new_n3336_), .Y(_0opcode_7_0__5_));
AND2X2 AND2X2_1449 ( .A(_abc_41356_new_n3319_), .B(\data[6] ), .Y(_abc_41356_new_n3339_));
AND2X2 AND2X2_145 ( .A(_abc_41356_new_n616_), .B(regfil_5__1_), .Y(_abc_41356_new_n749_));
AND2X2 AND2X2_1450 ( .A(_abc_41356_new_n3321_), .B(opcode_6_), .Y(_abc_41356_new_n3340_));
AND2X2 AND2X2_1451 ( .A(_abc_41356_new_n3319_), .B(\data[7] ), .Y(_abc_41356_new_n3342_));
AND2X2 AND2X2_1452 ( .A(_abc_41356_new_n3321_), .B(opcode_7_), .Y(_abc_41356_new_n3343_));
AND2X2 AND2X2_1453 ( .A(_abc_41356_new_n3345_), .B(eienb), .Y(_abc_41356_new_n3346_));
AND2X2 AND2X2_1454 ( .A(_abc_41356_new_n509_), .B(eienb), .Y(_abc_41356_new_n3348_));
AND2X2 AND2X2_1455 ( .A(_abc_41356_new_n599_), .B(_abc_41356_new_n681_), .Y(_abc_41356_new_n3349_));
AND2X2 AND2X2_1456 ( .A(_abc_41356_new_n3349_), .B(_abc_41356_new_n1233_), .Y(_abc_41356_new_n3350_));
AND2X2 AND2X2_1457 ( .A(_abc_41356_new_n3347_), .B(_abc_41356_new_n3351_), .Y(_0eienb_0_0_));
AND2X2 AND2X2_1458 ( .A(_abc_41356_new_n619_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n3354_));
AND2X2 AND2X2_1459 ( .A(_abc_41356_new_n3353_), .B(_abc_41356_new_n3355_), .Y(_abc_41356_new_n3356_));
AND2X2 AND2X2_146 ( .A(_abc_41356_new_n526_), .B(regfil_7__1_), .Y(_abc_41356_new_n751_));
AND2X2 AND2X2_1460 ( .A(_abc_41356_new_n2064_), .B(_abc_41356_new_n2054_), .Y(_abc_41356_new_n3358_));
AND2X2 AND2X2_1461 ( .A(_abc_41356_new_n3358_), .B(_abc_41356_new_n3357_), .Y(_abc_41356_new_n3359_));
AND2X2 AND2X2_1462 ( .A(_abc_41356_new_n3359_), .B(_abc_41356_new_n3356_), .Y(_abc_41356_new_n3360_));
AND2X2 AND2X2_1463 ( .A(_abc_41356_new_n578_), .B(_abc_41356_new_n616_), .Y(_abc_41356_new_n3361_));
AND2X2 AND2X2_1464 ( .A(_abc_41356_new_n2061_), .B(_abc_41356_new_n2066_), .Y(_abc_41356_new_n3363_));
AND2X2 AND2X2_1465 ( .A(_abc_41356_new_n3363_), .B(_abc_41356_new_n3362_), .Y(_abc_41356_new_n3364_));
AND2X2 AND2X2_1466 ( .A(_abc_41356_new_n2063_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n3365_));
AND2X2 AND2X2_1467 ( .A(_abc_41356_new_n3366_), .B(opcode_5_), .Y(_abc_41356_new_n3367_));
AND2X2 AND2X2_1468 ( .A(_abc_41356_new_n623_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n3368_));
AND2X2 AND2X2_1469 ( .A(_abc_41356_new_n3367_), .B(_abc_41356_new_n3368_), .Y(_abc_41356_new_n3369_));
AND2X2 AND2X2_147 ( .A(_abc_41356_new_n623_), .B(regfil_6__1_), .Y(_abc_41356_new_n752_));
AND2X2 AND2X2_1470 ( .A(_abc_41356_new_n2026_), .B(_abc_41356_new_n1413_), .Y(_abc_41356_new_n3371_));
AND2X2 AND2X2_1471 ( .A(_abc_41356_new_n598_), .B(_abc_41356_new_n623_), .Y(_abc_41356_new_n3372_));
AND2X2 AND2X2_1472 ( .A(_abc_41356_new_n3372_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3373_));
AND2X2 AND2X2_1473 ( .A(_abc_41356_new_n2026_), .B(_abc_41356_new_n576_), .Y(_abc_41356_new_n3377_));
AND2X2 AND2X2_1474 ( .A(_abc_41356_new_n3379_), .B(_abc_41356_new_n3365_), .Y(_abc_41356_new_n3380_));
AND2X2 AND2X2_1475 ( .A(_abc_41356_new_n3380_), .B(_abc_41356_new_n3364_), .Y(_abc_41356_new_n3381_));
AND2X2 AND2X2_1476 ( .A(_abc_41356_new_n3381_), .B(_abc_41356_new_n3360_), .Y(_abc_41356_new_n3382_));
AND2X2 AND2X2_1477 ( .A(_abc_41356_new_n3382_), .B(statesel_0_), .Y(_abc_41356_new_n3383_));
AND2X2 AND2X2_1478 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n1413_), .Y(_abc_41356_new_n3385_));
AND2X2 AND2X2_1479 ( .A(_abc_41356_new_n3389_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3390_));
AND2X2 AND2X2_148 ( .A(_abc_41356_new_n619_), .B(regfil_0__1_), .Y(_abc_41356_new_n756_));
AND2X2 AND2X2_1480 ( .A(_abc_41356_new_n678_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n3391_));
AND2X2 AND2X2_1481 ( .A(_abc_41356_new_n3368_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3393_));
AND2X2 AND2X2_1482 ( .A(_abc_41356_new_n3361_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3394_));
AND2X2 AND2X2_1483 ( .A(_abc_41356_new_n3361_), .B(opcode_5_), .Y(_abc_41356_new_n3395_));
AND2X2 AND2X2_1484 ( .A(_abc_41356_new_n3402_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3403_));
AND2X2 AND2X2_1485 ( .A(_abc_41356_new_n3403_), .B(_abc_41356_new_n3404_), .Y(_abc_41356_new_n3405_));
AND2X2 AND2X2_1486 ( .A(_abc_41356_new_n3406_), .B(statesel_0_), .Y(_abc_41356_new_n3407_));
AND2X2 AND2X2_1487 ( .A(_abc_41356_new_n683_), .B(_abc_41356_new_n677_), .Y(_abc_41356_new_n3408_));
AND2X2 AND2X2_1488 ( .A(_abc_41356_new_n3409_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n3410_));
AND2X2 AND2X2_1489 ( .A(_abc_41356_new_n678_), .B(_abc_41356_new_n682_), .Y(_abc_41356_new_n3411_));
AND2X2 AND2X2_149 ( .A(_abc_41356_new_n616_), .B(regfil_1__1_), .Y(_abc_41356_new_n757_));
AND2X2 AND2X2_1490 ( .A(_abc_41356_new_n3412_), .B(_abc_41356_new_n3410_), .Y(_abc_41356_new_n3413_));
AND2X2 AND2X2_1491 ( .A(_abc_41356_new_n2026_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3414_));
AND2X2 AND2X2_1492 ( .A(_abc_41356_new_n3416_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3417_));
AND2X2 AND2X2_1493 ( .A(_abc_41356_new_n3420_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n3421_));
AND2X2 AND2X2_1494 ( .A(_abc_41356_new_n521_), .B(_abc_41356_new_n708_), .Y(_abc_41356_new_n3423_));
AND2X2 AND2X2_1495 ( .A(_abc_41356_new_n3423_), .B(_abc_41356_new_n706_), .Y(_abc_41356_new_n3424_));
AND2X2 AND2X2_1496 ( .A(_abc_41356_new_n2926_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n3425_));
AND2X2 AND2X2_1497 ( .A(_abc_41356_new_n707_), .B(_abc_41356_new_n605_), .Y(_abc_41356_new_n3426_));
AND2X2 AND2X2_1498 ( .A(_abc_41356_new_n3426_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n3427_));
AND2X2 AND2X2_1499 ( .A(_abc_41356_new_n611_), .B(_abc_41356_new_n706_), .Y(_abc_41356_new_n3430_));
AND2X2 AND2X2_15 ( .A(_abc_41356_new_n523_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n524_));
AND2X2 AND2X2_150 ( .A(_abc_41356_new_n526_), .B(regfil_3__1_), .Y(_abc_41356_new_n759_));
AND2X2 AND2X2_1500 ( .A(_abc_41356_new_n605_), .B(_abc_41356_new_n610_), .Y(_abc_41356_new_n3431_));
AND2X2 AND2X2_1501 ( .A(_abc_41356_new_n3431_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n3432_));
AND2X2 AND2X2_1502 ( .A(_abc_41356_new_n1222_), .B(_abc_41356_new_n518_), .Y(_abc_41356_new_n3434_));
AND2X2 AND2X2_1503 ( .A(_abc_41356_new_n522_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n3440_));
AND2X2 AND2X2_1504 ( .A(_abc_41356_new_n3441_), .B(_abc_41356_new_n3265_), .Y(_abc_41356_new_n3442_));
AND2X2 AND2X2_1505 ( .A(_abc_41356_new_n3439_), .B(_abc_41356_new_n3442_), .Y(_abc_41356_new_n3443_));
AND2X2 AND2X2_1506 ( .A(_abc_41356_new_n509_), .B(waitr), .Y(_abc_41356_new_n3445_));
AND2X2 AND2X2_1507 ( .A(_abc_41356_new_n3440_), .B(_abc_41356_new_n3445_), .Y(_abc_41356_new_n3446_));
AND2X2 AND2X2_1508 ( .A(_abc_41356_new_n3447_), .B(statesel_0_), .Y(_abc_41356_new_n3448_));
AND2X2 AND2X2_1509 ( .A(_abc_41356_new_n3440_), .B(_abc_41356_new_n716_), .Y(_abc_41356_new_n3450_));
AND2X2 AND2X2_151 ( .A(_abc_41356_new_n623_), .B(regfil_2__1_), .Y(_abc_41356_new_n760_));
AND2X2 AND2X2_1510 ( .A(_abc_41356_new_n3454_), .B(_abc_41356_new_n3449_), .Y(_abc_41356_new_n3455_));
AND2X2 AND2X2_1511 ( .A(_abc_41356_new_n3382_), .B(statesel_1_), .Y(_abc_41356_new_n3458_));
AND2X2 AND2X2_1512 ( .A(_abc_41356_new_n3460_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3461_));
AND2X2 AND2X2_1513 ( .A(_abc_41356_new_n683_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n3462_));
AND2X2 AND2X2_1514 ( .A(_abc_41356_new_n3463_), .B(statesel_1_), .Y(_abc_41356_new_n3464_));
AND2X2 AND2X2_1515 ( .A(_abc_41356_new_n3368_), .B(_abc_41356_new_n535_), .Y(_abc_41356_new_n3465_));
AND2X2 AND2X2_1516 ( .A(_abc_41356_new_n3361_), .B(opcode_4_), .Y(_abc_41356_new_n3466_));
AND2X2 AND2X2_1517 ( .A(_abc_41356_new_n3470_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3471_));
AND2X2 AND2X2_1518 ( .A(_abc_41356_new_n3472_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n3473_));
AND2X2 AND2X2_1519 ( .A(_abc_41356_new_n3475_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n3476_));
AND2X2 AND2X2_152 ( .A(_abc_41356_new_n755_), .B(_abc_41356_new_n763_), .Y(_abc_41356_new_n764_));
AND2X2 AND2X2_1520 ( .A(_abc_41356_new_n3476_), .B(_abc_41356_new_n3474_), .Y(_abc_41356_new_n3477_));
AND2X2 AND2X2_1521 ( .A(_abc_41356_new_n3480_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3481_));
AND2X2 AND2X2_1522 ( .A(_abc_41356_new_n3440_), .B(waitr), .Y(_abc_41356_new_n3482_));
AND2X2 AND2X2_1523 ( .A(_abc_41356_new_n3482_), .B(statesel_1_), .Y(_abc_41356_new_n3483_));
AND2X2 AND2X2_1524 ( .A(_abc_41356_new_n3484_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3485_));
AND2X2 AND2X2_1525 ( .A(_abc_41356_new_n3444_), .B(statesel_1_), .Y(_abc_41356_new_n3486_));
AND2X2 AND2X2_1526 ( .A(_abc_41356_new_n3449_), .B(statesel_1_), .Y(_abc_41356_new_n3487_));
AND2X2 AND2X2_1527 ( .A(_abc_41356_new_n3488_), .B(statesel_0_), .Y(_abc_41356_new_n3489_));
AND2X2 AND2X2_1528 ( .A(_abc_41356_new_n3454_), .B(_abc_41356_new_n3490_), .Y(_abc_41356_new_n3491_));
AND2X2 AND2X2_1529 ( .A(_abc_41356_new_n3357_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n3494_));
AND2X2 AND2X2_153 ( .A(_abc_41356_new_n764_), .B(_abc_41356_new_n614_), .Y(_abc_41356_new_n765_));
AND2X2 AND2X2_1530 ( .A(_abc_41356_new_n3382_), .B(statesel_2_), .Y(_abc_41356_new_n3498_));
AND2X2 AND2X2_1531 ( .A(_abc_41356_new_n3499_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3500_));
AND2X2 AND2X2_1532 ( .A(_abc_41356_new_n3402_), .B(_abc_41356_new_n3501_), .Y(_abc_41356_new_n3502_));
AND2X2 AND2X2_1533 ( .A(_abc_41356_new_n3372_), .B(opcode_5_), .Y(_abc_41356_new_n3503_));
AND2X2 AND2X2_1534 ( .A(_abc_41356_new_n3507_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3508_));
AND2X2 AND2X2_1535 ( .A(_abc_41356_new_n3506_), .B(_abc_41356_new_n3508_), .Y(_abc_41356_new_n3509_));
AND2X2 AND2X2_1536 ( .A(_abc_41356_new_n3410_), .B(_abc_41356_new_n3475_), .Y(_abc_41356_new_n3510_));
AND2X2 AND2X2_1537 ( .A(_abc_41356_new_n3511_), .B(statesel_2_), .Y(_abc_41356_new_n3512_));
AND2X2 AND2X2_1538 ( .A(_abc_41356_new_n3514_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3515_));
AND2X2 AND2X2_1539 ( .A(_abc_41356_new_n3482_), .B(statesel_2_), .Y(_abc_41356_new_n3516_));
AND2X2 AND2X2_154 ( .A(_abc_41356_new_n612_), .B(alu_res_1_), .Y(_abc_41356_new_n766_));
AND2X2 AND2X2_1540 ( .A(_abc_41356_new_n3517_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3518_));
AND2X2 AND2X2_1541 ( .A(_abc_41356_new_n3444_), .B(statesel_2_), .Y(_abc_41356_new_n3519_));
AND2X2 AND2X2_1542 ( .A(statesel_0_), .B(statesel_1_), .Y(_abc_41356_new_n3520_));
AND2X2 AND2X2_1543 ( .A(_abc_41356_new_n3520_), .B(statesel_2_), .Y(_abc_41356_new_n3521_));
AND2X2 AND2X2_1544 ( .A(_abc_41356_new_n3438_), .B(_abc_41356_new_n3522_), .Y(_abc_41356_new_n3523_));
AND2X2 AND2X2_1545 ( .A(_abc_41356_new_n3450_), .B(_abc_41356_new_n3522_), .Y(_abc_41356_new_n3524_));
AND2X2 AND2X2_1546 ( .A(_abc_41356_new_n3526_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3527_));
AND2X2 AND2X2_1547 ( .A(_abc_41356_new_n3525_), .B(_abc_41356_new_n3527_), .Y(_abc_41356_new_n3528_));
AND2X2 AND2X2_1548 ( .A(_abc_41356_new_n3444_), .B(statesel_3_), .Y(_abc_41356_new_n3531_));
AND2X2 AND2X2_1549 ( .A(_abc_41356_new_n3382_), .B(statesel_3_), .Y(_abc_41356_new_n3532_));
AND2X2 AND2X2_155 ( .A(_abc_41356_new_n767_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n768_));
AND2X2 AND2X2_1550 ( .A(_abc_41356_new_n3536_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3537_));
AND2X2 AND2X2_1551 ( .A(_abc_41356_new_n3402_), .B(_abc_41356_new_n3540_), .Y(_abc_41356_new_n3541_));
AND2X2 AND2X2_1552 ( .A(_abc_41356_new_n3543_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3544_));
AND2X2 AND2X2_1553 ( .A(_abc_41356_new_n3542_), .B(_abc_41356_new_n3544_), .Y(_abc_41356_new_n3545_));
AND2X2 AND2X2_1554 ( .A(_abc_41356_new_n677_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n3546_));
AND2X2 AND2X2_1555 ( .A(_abc_41356_new_n3548_), .B(_abc_41356_new_n3547_), .Y(_abc_41356_new_n3549_));
AND2X2 AND2X2_1556 ( .A(_abc_41356_new_n3551_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3552_));
AND2X2 AND2X2_1557 ( .A(_abc_41356_new_n3553_), .B(statesel_2_), .Y(_abc_41356_new_n3554_));
AND2X2 AND2X2_1558 ( .A(_abc_41356_new_n3554_), .B(_abc_41356_new_n3520_), .Y(_abc_41356_new_n3555_));
AND2X2 AND2X2_1559 ( .A(_abc_41356_new_n3451_), .B(_abc_41356_new_n3555_), .Y(_abc_41356_new_n3556_));
AND2X2 AND2X2_156 ( .A(_abc_41356_new_n773_), .B(_abc_41356_new_n724_), .Y(_abc_41356_new_n774_));
AND2X2 AND2X2_1560 ( .A(_abc_41356_new_n3440_), .B(_abc_41356_new_n3522_), .Y(_abc_41356_new_n3557_));
AND2X2 AND2X2_1561 ( .A(_abc_41356_new_n3559_), .B(statesel_3_), .Y(_abc_41356_new_n3560_));
AND2X2 AND2X2_1562 ( .A(_abc_41356_new_n3562_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3563_));
AND2X2 AND2X2_1563 ( .A(_abc_41356_new_n3444_), .B(statesel_4_), .Y(_abc_41356_new_n3565_));
AND2X2 AND2X2_1564 ( .A(_abc_41356_new_n3381_), .B(statesel_4_), .Y(_abc_41356_new_n3567_));
AND2X2 AND2X2_1565 ( .A(_abc_41356_new_n3568_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3569_));
AND2X2 AND2X2_1566 ( .A(_abc_41356_new_n3570_), .B(statesel_4_), .Y(_abc_41356_new_n3571_));
AND2X2 AND2X2_1567 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n3572_));
AND2X2 AND2X2_1568 ( .A(_abc_41356_new_n3573_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3574_));
AND2X2 AND2X2_1569 ( .A(_abc_41356_new_n3577_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3578_));
AND2X2 AND2X2_157 ( .A(_abc_41356_new_n772_), .B(_abc_41356_new_n774_), .Y(_abc_41356_new_n775_));
AND2X2 AND2X2_1570 ( .A(_abc_41356_new_n3482_), .B(statesel_4_), .Y(_abc_41356_new_n3579_));
AND2X2 AND2X2_1571 ( .A(statesel_2_), .B(statesel_3_), .Y(_abc_41356_new_n3580_));
AND2X2 AND2X2_1572 ( .A(_abc_41356_new_n3520_), .B(_abc_41356_new_n3580_), .Y(_abc_41356_new_n3581_));
AND2X2 AND2X2_1573 ( .A(_abc_41356_new_n3581_), .B(statesel_4_), .Y(_abc_41356_new_n3583_));
AND2X2 AND2X2_1574 ( .A(_abc_41356_new_n3438_), .B(_abc_41356_new_n3584_), .Y(_abc_41356_new_n3585_));
AND2X2 AND2X2_1575 ( .A(_abc_41356_new_n3450_), .B(_abc_41356_new_n3584_), .Y(_abc_41356_new_n3586_));
AND2X2 AND2X2_1576 ( .A(_abc_41356_new_n3587_), .B(_abc_41356_new_n3582_), .Y(_abc_41356_new_n3588_));
AND2X2 AND2X2_1577 ( .A(_abc_41356_new_n3590_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3591_));
AND2X2 AND2X2_1578 ( .A(_abc_41356_new_n3444_), .B(statesel_5_), .Y(_abc_41356_new_n3593_));
AND2X2 AND2X2_1579 ( .A(_abc_41356_new_n3382_), .B(_abc_41356_new_n3594_), .Y(_abc_41356_new_n3595_));
AND2X2 AND2X2_158 ( .A(_abc_41356_new_n530_), .B(regfil_7__2_), .Y(_abc_41356_new_n776_));
AND2X2 AND2X2_1580 ( .A(_abc_41356_new_n3596_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3597_));
AND2X2 AND2X2_1581 ( .A(_abc_41356_new_n3570_), .B(statesel_5_), .Y(_abc_41356_new_n3598_));
AND2X2 AND2X2_1582 ( .A(_abc_41356_new_n3001_), .B(_abc_41356_new_n682_), .Y(_abc_41356_new_n3599_));
AND2X2 AND2X2_1583 ( .A(_abc_41356_new_n3602_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3603_));
AND2X2 AND2X2_1584 ( .A(_abc_41356_new_n3584_), .B(_abc_41356_new_n3440_), .Y(_abc_41356_new_n3604_));
AND2X2 AND2X2_1585 ( .A(_abc_41356_new_n3606_), .B(statesel_5_), .Y(_abc_41356_new_n3607_));
AND2X2 AND2X2_1586 ( .A(_abc_41356_new_n3594_), .B(statesel_4_), .Y(_abc_41356_new_n3608_));
AND2X2 AND2X2_1587 ( .A(_abc_41356_new_n3581_), .B(_abc_41356_new_n3608_), .Y(_abc_41356_new_n3609_));
AND2X2 AND2X2_1588 ( .A(_abc_41356_new_n3451_), .B(_abc_41356_new_n3609_), .Y(_abc_41356_new_n3610_));
AND2X2 AND2X2_1589 ( .A(_abc_41356_new_n3612_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3613_));
AND2X2 AND2X2_159 ( .A(_abc_41356_new_n555_), .B(regfil_7__0_), .Y(_abc_41356_new_n777_));
AND2X2 AND2X2_1590 ( .A(_abc_41356_new_n1234_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n3615_));
AND2X2 AND2X2_1591 ( .A(_abc_41356_new_n3617_), .B(_abc_41356_new_n3618_), .Y(_0popdes_1_0__0_));
AND2X2 AND2X2_1592 ( .A(_abc_41356_new_n3620_), .B(_abc_41356_new_n3621_), .Y(_0popdes_1_0__1_));
AND2X2 AND2X2_1593 ( .A(_abc_41356_new_n3440_), .B(_abc_41356_new_n717_), .Y(_abc_41356_new_n3623_));
AND2X2 AND2X2_1594 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n564_), .Y(_abc_41356_new_n3625_));
AND2X2 AND2X2_1595 ( .A(_abc_41356_new_n3626_), .B(_abc_41356_new_n3624_), .Y(_0rdatahold2_7_0__0_));
AND2X2 AND2X2_1596 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n3629_), .Y(_abc_41356_new_n3630_));
AND2X2 AND2X2_1597 ( .A(_abc_41356_new_n3631_), .B(_abc_41356_new_n3628_), .Y(_0rdatahold2_7_0__1_));
AND2X2 AND2X2_1598 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n829_), .Y(_abc_41356_new_n3634_));
AND2X2 AND2X2_1599 ( .A(_abc_41356_new_n3635_), .B(_abc_41356_new_n3633_), .Y(_0rdatahold2_7_0__2_));
AND2X2 AND2X2_16 ( .A(opcode_1_), .B(opcode_0_), .Y(_abc_41356_new_n526_));
AND2X2 AND2X2_160 ( .A(_abc_41356_new_n698_), .B(_abc_41356_new_n513_), .Y(_abc_41356_new_n778_));
AND2X2 AND2X2_1600 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n890_), .Y(_abc_41356_new_n3638_));
AND2X2 AND2X2_1601 ( .A(_abc_41356_new_n3639_), .B(_abc_41356_new_n3637_), .Y(_0rdatahold2_7_0__3_));
AND2X2 AND2X2_1602 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n3642_), .Y(_abc_41356_new_n3643_));
AND2X2 AND2X2_1603 ( .A(_abc_41356_new_n3644_), .B(_abc_41356_new_n3641_), .Y(_0rdatahold2_7_0__4_));
AND2X2 AND2X2_1604 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n1024_), .Y(_abc_41356_new_n3647_));
AND2X2 AND2X2_1605 ( .A(_abc_41356_new_n3648_), .B(_abc_41356_new_n3646_), .Y(_0rdatahold2_7_0__5_));
AND2X2 AND2X2_1606 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n1097_), .Y(_abc_41356_new_n3651_));
AND2X2 AND2X2_1607 ( .A(_abc_41356_new_n3652_), .B(_abc_41356_new_n3650_), .Y(_0rdatahold2_7_0__6_));
AND2X2 AND2X2_1608 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n2852_), .Y(_abc_41356_new_n3655_));
AND2X2 AND2X2_1609 ( .A(_abc_41356_new_n3656_), .B(_abc_41356_new_n3654_), .Y(_0rdatahold2_7_0__7_));
AND2X2 AND2X2_161 ( .A(_abc_41356_new_n712_), .B(regfil_7__1_), .Y(_abc_41356_new_n781_));
AND2X2 AND2X2_1610 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n3659_), .Y(_abc_41356_new_n3660_));
AND2X2 AND2X2_1611 ( .A(_abc_41356_new_n3661_), .B(_abc_41356_new_n3658_), .Y(_0rdatahold_7_0__0_));
AND2X2 AND2X2_1612 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n3664_), .Y(_abc_41356_new_n3665_));
AND2X2 AND2X2_1613 ( .A(_abc_41356_new_n3666_), .B(_abc_41356_new_n3663_), .Y(_0rdatahold_7_0__1_));
AND2X2 AND2X2_1614 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n3669_), .Y(_abc_41356_new_n3670_));
AND2X2 AND2X2_1615 ( .A(_abc_41356_new_n3671_), .B(_abc_41356_new_n3668_), .Y(_0rdatahold_7_0__2_));
AND2X2 AND2X2_1616 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n3674_), .Y(_abc_41356_new_n3675_));
AND2X2 AND2X2_1617 ( .A(_abc_41356_new_n3676_), .B(_abc_41356_new_n3673_), .Y(_0rdatahold_7_0__3_));
AND2X2 AND2X2_1618 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n3679_), .Y(_abc_41356_new_n3680_));
AND2X2 AND2X2_1619 ( .A(_abc_41356_new_n3681_), .B(_abc_41356_new_n3678_), .Y(_0rdatahold_7_0__4_));
AND2X2 AND2X2_162 ( .A(_abc_41356_new_n714_), .B(alu_res_1_), .Y(_abc_41356_new_n782_));
AND2X2 AND2X2_1620 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n3684_), .Y(_abc_41356_new_n3685_));
AND2X2 AND2X2_1621 ( .A(_abc_41356_new_n3686_), .B(_abc_41356_new_n3683_), .Y(_0rdatahold_7_0__5_));
AND2X2 AND2X2_1622 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n3689_), .Y(_abc_41356_new_n3690_));
AND2X2 AND2X2_1623 ( .A(_abc_41356_new_n3691_), .B(_abc_41356_new_n3688_), .Y(_0rdatahold_7_0__6_));
AND2X2 AND2X2_1624 ( .A(_abc_41356_new_n3623_), .B(_abc_41356_new_n3694_), .Y(_abc_41356_new_n3695_));
AND2X2 AND2X2_1625 ( .A(_abc_41356_new_n3696_), .B(_abc_41356_new_n3693_), .Y(_0rdatahold_7_0__7_));
AND2X2 AND2X2_1626 ( .A(_abc_41356_new_n3426_), .B(_abc_41356_new_n518_), .Y(_abc_41356_new_n3698_));
AND2X2 AND2X2_1627 ( .A(_abc_41356_new_n3265_), .B(_abc_41356_new_n3699_), .Y(_abc_41356_new_n3700_));
AND2X2 AND2X2_1628 ( .A(_abc_41356_new_n3701_), .B(_abc_41356_new_n3702_), .Y(_abc_41356_new_n3703_));
AND2X2 AND2X2_1629 ( .A(_abc_41356_new_n3703_), .B(_abc_41356_new_n3700_), .Y(_abc_41356_new_n3704_));
AND2X2 AND2X2_163 ( .A(_abc_41356_new_n512_), .B(rdatahold_1_), .Y(_abc_41356_new_n783_));
AND2X2 AND2X2_1630 ( .A(_abc_41356_new_n3705_), .B(wdatahold_0_), .Y(_abc_41356_new_n3706_));
AND2X2 AND2X2_1631 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3707_));
AND2X2 AND2X2_1632 ( .A(_abc_41356_new_n3708_), .B(wdatahold_0_), .Y(_abc_41356_new_n3709_));
AND2X2 AND2X2_1633 ( .A(_abc_41356_new_n535_), .B(regfil_5__0_), .Y(_abc_41356_new_n3711_));
AND2X2 AND2X2_1634 ( .A(_abc_41356_new_n2056_), .B(regfil_7__0_), .Y(_abc_41356_new_n3712_));
AND2X2 AND2X2_1635 ( .A(_abc_41356_new_n3715_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3716_));
AND2X2 AND2X2_1636 ( .A(_abc_41356_new_n3714_), .B(_abc_41356_new_n3716_), .Y(_abc_41356_new_n3717_));
AND2X2 AND2X2_1637 ( .A(_abc_41356_new_n3719_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n3720_));
AND2X2 AND2X2_1638 ( .A(_abc_41356_new_n3718_), .B(_abc_41356_new_n3720_), .Y(_abc_41356_new_n3721_));
AND2X2 AND2X2_1639 ( .A(_abc_41356_new_n3724_), .B(_abc_41356_new_n3723_), .Y(_abc_41356_new_n3725_));
AND2X2 AND2X2_164 ( .A(_abc_41356_new_n718_), .B(\data[1] ), .Y(_abc_41356_new_n784_));
AND2X2 AND2X2_1640 ( .A(pc_0_), .B(intcyc), .Y(_abc_41356_new_n3726_));
AND2X2 AND2X2_1641 ( .A(_abc_41356_new_n3723_), .B(_abc_41356_new_n2049_), .Y(_abc_41356_new_n3727_));
AND2X2 AND2X2_1642 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n3728_), .Y(_abc_41356_new_n3729_));
AND2X2 AND2X2_1643 ( .A(_abc_41356_new_n681_), .B(carry), .Y(_abc_41356_new_n3730_));
AND2X2 AND2X2_1644 ( .A(_abc_41356_new_n3732_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3733_));
AND2X2 AND2X2_1645 ( .A(_abc_41356_new_n3736_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n3737_));
AND2X2 AND2X2_1646 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n3711_), .Y(_abc_41356_new_n3738_));
AND2X2 AND2X2_1647 ( .A(_abc_41356_new_n3739_), .B(_abc_41356_new_n3734_), .Y(_abc_41356_new_n3740_));
AND2X2 AND2X2_1648 ( .A(_abc_41356_new_n3742_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3743_));
AND2X2 AND2X2_1649 ( .A(_abc_41356_new_n3745_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3746_));
AND2X2 AND2X2_165 ( .A(_abc_41356_new_n736_), .B(regfil_0__2_), .Y(_abc_41356_new_n792_));
AND2X2 AND2X2_1650 ( .A(_abc_41356_new_n3430_), .B(alu_res_0_), .Y(_abc_41356_new_n3747_));
AND2X2 AND2X2_1651 ( .A(_abc_41356_new_n3698_), .B(wdatahold2_0_), .Y(_abc_41356_new_n3748_));
AND2X2 AND2X2_1652 ( .A(_abc_41356_new_n3427_), .B(rdatahold_0_), .Y(_abc_41356_new_n3749_));
AND2X2 AND2X2_1653 ( .A(_abc_41356_new_n3752_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3753_));
AND2X2 AND2X2_1654 ( .A(_abc_41356_new_n3705_), .B(wdatahold_1_), .Y(_abc_41356_new_n3755_));
AND2X2 AND2X2_1655 ( .A(_abc_41356_new_n3710_), .B(_abc_41356_new_n514_), .Y(_abc_41356_new_n3756_));
AND2X2 AND2X2_1656 ( .A(_abc_41356_new_n3758_), .B(wdatahold_1_), .Y(_abc_41356_new_n3759_));
AND2X2 AND2X2_1657 ( .A(pc_1_), .B(pc_0_), .Y(_abc_41356_new_n3760_));
AND2X2 AND2X2_1658 ( .A(_abc_41356_new_n3761_), .B(_abc_41356_new_n2033_), .Y(_abc_41356_new_n3762_));
AND2X2 AND2X2_1659 ( .A(_abc_41356_new_n2060_), .B(_abc_41356_new_n3762_), .Y(_abc_41356_new_n3763_));
AND2X2 AND2X2_166 ( .A(_abc_41356_new_n793_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n794_));
AND2X2 AND2X2_1660 ( .A(_abc_41356_new_n3765_), .B(_abc_41356_new_n3766_), .Y(_abc_41356_new_n3767_));
AND2X2 AND2X2_1661 ( .A(_abc_41356_new_n3767_), .B(_abc_41356_new_n2048_), .Y(_abc_41356_new_n3768_));
AND2X2 AND2X2_1662 ( .A(_abc_41356_new_n3764_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n3769_));
AND2X2 AND2X2_1663 ( .A(opcode_5_), .B(regfil_5__1_), .Y(_abc_41356_new_n3771_));
AND2X2 AND2X2_1664 ( .A(_abc_41356_new_n534_), .B(regfil_1__1_), .Y(_abc_41356_new_n3772_));
AND2X2 AND2X2_1665 ( .A(_abc_41356_new_n3772_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3773_));
AND2X2 AND2X2_1666 ( .A(opcode_4_), .B(regfil_3__1_), .Y(_abc_41356_new_n3774_));
AND2X2 AND2X2_1667 ( .A(_abc_41356_new_n3776_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n3777_));
AND2X2 AND2X2_1668 ( .A(_abc_41356_new_n2376_), .B(_abc_41356_new_n2994_), .Y(_abc_41356_new_n3779_));
AND2X2 AND2X2_1669 ( .A(_abc_41356_new_n3778_), .B(_abc_41356_new_n3780_), .Y(_abc_41356_new_n3781_));
AND2X2 AND2X2_167 ( .A(_abc_41356_new_n743_), .B(regfil_0__2_), .Y(_abc_41356_new_n796_));
AND2X2 AND2X2_1670 ( .A(_abc_41356_new_n2096_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3784_));
AND2X2 AND2X2_1671 ( .A(_abc_41356_new_n3784_), .B(_abc_41356_new_n3783_), .Y(_abc_41356_new_n3785_));
AND2X2 AND2X2_1672 ( .A(_abc_41356_new_n2027_), .B(regfil_5__1_), .Y(_abc_41356_new_n3786_));
AND2X2 AND2X2_1673 ( .A(_abc_41356_new_n2056_), .B(regfil_7__1_), .Y(_abc_41356_new_n3787_));
AND2X2 AND2X2_1674 ( .A(_abc_41356_new_n3787_), .B(_abc_41356_new_n2026_), .Y(_abc_41356_new_n3788_));
AND2X2 AND2X2_1675 ( .A(_abc_41356_new_n3789_), .B(_abc_41356_new_n514_), .Y(_abc_41356_new_n3790_));
AND2X2 AND2X2_1676 ( .A(_abc_41356_new_n3411_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n3791_));
AND2X2 AND2X2_1677 ( .A(_abc_41356_new_n764_), .B(_abc_41356_new_n3791_), .Y(_abc_41356_new_n3792_));
AND2X2 AND2X2_1678 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n3797_), .Y(_abc_41356_new_n3798_));
AND2X2 AND2X2_1679 ( .A(_abc_41356_new_n3796_), .B(_abc_41356_new_n3798_), .Y(_abc_41356_new_n3799_));
AND2X2 AND2X2_168 ( .A(_abc_41356_new_n797_), .B(_abc_41356_new_n581_), .Y(_abc_41356_new_n798_));
AND2X2 AND2X2_1680 ( .A(_abc_41356_new_n3430_), .B(alu_res_1_), .Y(_abc_41356_new_n3800_));
AND2X2 AND2X2_1681 ( .A(_abc_41356_new_n3698_), .B(wdatahold2_1_), .Y(_abc_41356_new_n3801_));
AND2X2 AND2X2_1682 ( .A(_abc_41356_new_n3427_), .B(rdatahold_1_), .Y(_abc_41356_new_n3802_));
AND2X2 AND2X2_1683 ( .A(_abc_41356_new_n3805_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3806_));
AND2X2 AND2X2_1684 ( .A(_abc_41356_new_n3705_), .B(wdatahold_2_), .Y(_abc_41356_new_n3808_));
AND2X2 AND2X2_1685 ( .A(_abc_41356_new_n2069_), .B(wdatahold_2_), .Y(_abc_41356_new_n3809_));
AND2X2 AND2X2_1686 ( .A(_abc_41356_new_n2070_), .B(pc_0_), .Y(_abc_41356_new_n3810_));
AND2X2 AND2X2_1687 ( .A(_abc_41356_new_n3761_), .B(_abc_41356_new_n3811_), .Y(_abc_41356_new_n3812_));
AND2X2 AND2X2_1688 ( .A(_abc_41356_new_n2060_), .B(_abc_41356_new_n3814_), .Y(_abc_41356_new_n3815_));
AND2X2 AND2X2_1689 ( .A(_abc_41356_new_n3811_), .B(_abc_41356_new_n3817_), .Y(_abc_41356_new_n3818_));
AND2X2 AND2X2_169 ( .A(_abc_41356_new_n798_), .B(_abc_41356_new_n795_), .Y(_abc_41356_new_n799_));
AND2X2 AND2X2_1690 ( .A(_abc_41356_new_n3818_), .B(_abc_41356_new_n3723_), .Y(_abc_41356_new_n3819_));
AND2X2 AND2X2_1691 ( .A(_abc_41356_new_n3822_), .B(_abc_41356_new_n3816_), .Y(_abc_41356_new_n3823_));
AND2X2 AND2X2_1692 ( .A(_abc_41356_new_n3823_), .B(_abc_41356_new_n2048_), .Y(_abc_41356_new_n3824_));
AND2X2 AND2X2_1693 ( .A(_abc_41356_new_n681_), .B(parity), .Y(_abc_41356_new_n3825_));
AND2X2 AND2X2_1694 ( .A(_abc_41356_new_n535_), .B(regfil_5__2_), .Y(_abc_41356_new_n3826_));
AND2X2 AND2X2_1695 ( .A(_abc_41356_new_n3827_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3828_));
AND2X2 AND2X2_1696 ( .A(_abc_41356_new_n3831_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n3832_));
AND2X2 AND2X2_1697 ( .A(_abc_41356_new_n3830_), .B(_abc_41356_new_n3832_), .Y(_abc_41356_new_n3833_));
AND2X2 AND2X2_1698 ( .A(_abc_41356_new_n3821_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n3834_));
AND2X2 AND2X2_1699 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n3826_), .Y(_abc_41356_new_n3835_));
AND2X2 AND2X2_17 ( .A(opcode_3_), .B(opcode_2_), .Y(_abc_41356_new_n527_));
AND2X2 AND2X2_170 ( .A(_abc_41356_new_n642_), .B(rdatahold_2_), .Y(_abc_41356_new_n800_));
AND2X2 AND2X2_1700 ( .A(_abc_41356_new_n3840_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3841_));
AND2X2 AND2X2_1701 ( .A(_abc_41356_new_n817_), .B(_abc_41356_new_n3791_), .Y(_abc_41356_new_n3842_));
AND2X2 AND2X2_1702 ( .A(_abc_41356_new_n2056_), .B(regfil_7__2_), .Y(_abc_41356_new_n3843_));
AND2X2 AND2X2_1703 ( .A(_abc_41356_new_n3846_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3847_));
AND2X2 AND2X2_1704 ( .A(_abc_41356_new_n3845_), .B(_abc_41356_new_n3847_), .Y(_abc_41356_new_n3848_));
AND2X2 AND2X2_1705 ( .A(_abc_41356_new_n3849_), .B(wdatahold_2_), .Y(_abc_41356_new_n3850_));
AND2X2 AND2X2_1706 ( .A(_abc_41356_new_n3853_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3854_));
AND2X2 AND2X2_1707 ( .A(_abc_41356_new_n3430_), .B(alu_res_2_), .Y(_abc_41356_new_n3855_));
AND2X2 AND2X2_1708 ( .A(_abc_41356_new_n3698_), .B(wdatahold2_2_), .Y(_abc_41356_new_n3856_));
AND2X2 AND2X2_1709 ( .A(_abc_41356_new_n3427_), .B(rdatahold_2_), .Y(_abc_41356_new_n3857_));
AND2X2 AND2X2_171 ( .A(_abc_41356_new_n616_), .B(regfil_1__2_), .Y(_abc_41356_new_n801_));
AND2X2 AND2X2_1710 ( .A(_abc_41356_new_n3860_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3861_));
AND2X2 AND2X2_1711 ( .A(_abc_41356_new_n3705_), .B(wdatahold_3_), .Y(_abc_41356_new_n3863_));
AND2X2 AND2X2_1712 ( .A(_abc_41356_new_n3708_), .B(wdatahold_3_), .Y(_abc_41356_new_n3864_));
AND2X2 AND2X2_1713 ( .A(_abc_41356_new_n535_), .B(regfil_5__3_), .Y(_abc_41356_new_n3865_));
AND2X2 AND2X2_1714 ( .A(_abc_41356_new_n2056_), .B(regfil_7__3_), .Y(_abc_41356_new_n3866_));
AND2X2 AND2X2_1715 ( .A(_abc_41356_new_n3869_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3870_));
AND2X2 AND2X2_1716 ( .A(_abc_41356_new_n3868_), .B(_abc_41356_new_n3870_), .Y(_abc_41356_new_n3871_));
AND2X2 AND2X2_1717 ( .A(_abc_41356_new_n3873_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n3874_));
AND2X2 AND2X2_1718 ( .A(_abc_41356_new_n3872_), .B(_abc_41356_new_n3874_), .Y(_abc_41356_new_n3875_));
AND2X2 AND2X2_1719 ( .A(_abc_41356_new_n3877_), .B(_abc_41356_new_n3878_), .Y(_abc_41356_new_n3879_));
AND2X2 AND2X2_172 ( .A(_abc_41356_new_n619_), .B(regfil_0__2_), .Y(_abc_41356_new_n802_));
AND2X2 AND2X2_1720 ( .A(_abc_41356_new_n2060_), .B(_abc_41356_new_n3879_), .Y(_abc_41356_new_n3880_));
AND2X2 AND2X2_1721 ( .A(_abc_41356_new_n3881_), .B(_abc_41356_new_n3882_), .Y(_abc_41356_new_n3883_));
AND2X2 AND2X2_1722 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n3885_), .Y(_abc_41356_new_n3886_));
AND2X2 AND2X2_1723 ( .A(_abc_41356_new_n3884_), .B(_abc_41356_new_n3886_), .Y(_abc_41356_new_n3887_));
AND2X2 AND2X2_1724 ( .A(_abc_41356_new_n3883_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n3888_));
AND2X2 AND2X2_1725 ( .A(_abc_41356_new_n3889_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3890_));
AND2X2 AND2X2_1726 ( .A(_abc_41356_new_n3892_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n3893_));
AND2X2 AND2X2_1727 ( .A(_abc_41356_new_n3893_), .B(_abc_41356_new_n3891_), .Y(_abc_41356_new_n3894_));
AND2X2 AND2X2_1728 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n3865_), .Y(_abc_41356_new_n3895_));
AND2X2 AND2X2_1729 ( .A(_abc_41356_new_n3899_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3900_));
AND2X2 AND2X2_173 ( .A(_abc_41356_new_n526_), .B(regfil_3__2_), .Y(_abc_41356_new_n804_));
AND2X2 AND2X2_1730 ( .A(_abc_41356_new_n3902_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3903_));
AND2X2 AND2X2_1731 ( .A(_abc_41356_new_n3430_), .B(alu_res_3_), .Y(_abc_41356_new_n3904_));
AND2X2 AND2X2_1732 ( .A(_abc_41356_new_n3698_), .B(wdatahold2_3_), .Y(_abc_41356_new_n3905_));
AND2X2 AND2X2_1733 ( .A(_abc_41356_new_n3427_), .B(rdatahold_3_), .Y(_abc_41356_new_n3906_));
AND2X2 AND2X2_1734 ( .A(_abc_41356_new_n3909_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3910_));
AND2X2 AND2X2_1735 ( .A(_abc_41356_new_n3705_), .B(wdatahold_4_), .Y(_abc_41356_new_n3912_));
AND2X2 AND2X2_1736 ( .A(_abc_41356_new_n3708_), .B(wdatahold_4_), .Y(_abc_41356_new_n3913_));
AND2X2 AND2X2_1737 ( .A(_abc_41356_new_n535_), .B(regfil_5__4_), .Y(_abc_41356_new_n3914_));
AND2X2 AND2X2_1738 ( .A(_abc_41356_new_n2056_), .B(regfil_7__4_), .Y(_abc_41356_new_n3915_));
AND2X2 AND2X2_1739 ( .A(_abc_41356_new_n3918_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3919_));
AND2X2 AND2X2_174 ( .A(_abc_41356_new_n623_), .B(regfil_2__2_), .Y(_abc_41356_new_n805_));
AND2X2 AND2X2_1740 ( .A(_abc_41356_new_n3917_), .B(_abc_41356_new_n3919_), .Y(_abc_41356_new_n3920_));
AND2X2 AND2X2_1741 ( .A(_abc_41356_new_n3922_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n3923_));
AND2X2 AND2X2_1742 ( .A(_abc_41356_new_n3921_), .B(_abc_41356_new_n3923_), .Y(_abc_41356_new_n3924_));
AND2X2 AND2X2_1743 ( .A(_abc_41356_new_n2072_), .B(pc_4_), .Y(_abc_41356_new_n3926_));
AND2X2 AND2X2_1744 ( .A(_abc_41356_new_n3927_), .B(_abc_41356_new_n3928_), .Y(_abc_41356_new_n3929_));
AND2X2 AND2X2_1745 ( .A(_abc_41356_new_n2060_), .B(_abc_41356_new_n3929_), .Y(_abc_41356_new_n3930_));
AND2X2 AND2X2_1746 ( .A(_abc_41356_new_n2035_), .B(pc_4_), .Y(_abc_41356_new_n3931_));
AND2X2 AND2X2_1747 ( .A(_abc_41356_new_n3932_), .B(_abc_41356_new_n3933_), .Y(_abc_41356_new_n3934_));
AND2X2 AND2X2_1748 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n3936_), .Y(_abc_41356_new_n3937_));
AND2X2 AND2X2_1749 ( .A(_abc_41356_new_n3935_), .B(_abc_41356_new_n3937_), .Y(_abc_41356_new_n3938_));
AND2X2 AND2X2_175 ( .A(_abc_41356_new_n616_), .B(regfil_5__2_), .Y(_abc_41356_new_n809_));
AND2X2 AND2X2_1750 ( .A(_abc_41356_new_n3934_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n3939_));
AND2X2 AND2X2_1751 ( .A(_abc_41356_new_n681_), .B(auxcar), .Y(_abc_41356_new_n3940_));
AND2X2 AND2X2_1752 ( .A(_abc_41356_new_n3942_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3943_));
AND2X2 AND2X2_1753 ( .A(_abc_41356_new_n3945_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n3946_));
AND2X2 AND2X2_1754 ( .A(_abc_41356_new_n3944_), .B(_abc_41356_new_n3946_), .Y(_abc_41356_new_n3947_));
AND2X2 AND2X2_1755 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n3914_), .Y(_abc_41356_new_n3948_));
AND2X2 AND2X2_1756 ( .A(_abc_41356_new_n3952_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n3953_));
AND2X2 AND2X2_1757 ( .A(_abc_41356_new_n3955_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3956_));
AND2X2 AND2X2_1758 ( .A(_abc_41356_new_n3430_), .B(alu_res_4_), .Y(_abc_41356_new_n3957_));
AND2X2 AND2X2_1759 ( .A(_abc_41356_new_n3698_), .B(wdatahold2_4_), .Y(_abc_41356_new_n3958_));
AND2X2 AND2X2_176 ( .A(_abc_41356_new_n623_), .B(regfil_6__2_), .Y(_abc_41356_new_n811_));
AND2X2 AND2X2_1760 ( .A(_abc_41356_new_n3427_), .B(rdatahold_4_), .Y(_abc_41356_new_n3959_));
AND2X2 AND2X2_1761 ( .A(_abc_41356_new_n3962_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n3963_));
AND2X2 AND2X2_1762 ( .A(_abc_41356_new_n3705_), .B(wdatahold_5_), .Y(_abc_41356_new_n3965_));
AND2X2 AND2X2_1763 ( .A(_abc_41356_new_n3708_), .B(wdatahold_5_), .Y(_abc_41356_new_n3966_));
AND2X2 AND2X2_1764 ( .A(_abc_41356_new_n535_), .B(regfil_5__5_), .Y(_abc_41356_new_n3967_));
AND2X2 AND2X2_1765 ( .A(_abc_41356_new_n2056_), .B(regfil_7__5_), .Y(_abc_41356_new_n3968_));
AND2X2 AND2X2_1766 ( .A(_abc_41356_new_n3971_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n3972_));
AND2X2 AND2X2_1767 ( .A(_abc_41356_new_n3970_), .B(_abc_41356_new_n3972_), .Y(_abc_41356_new_n3973_));
AND2X2 AND2X2_1768 ( .A(_abc_41356_new_n3975_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n3976_));
AND2X2 AND2X2_1769 ( .A(_abc_41356_new_n3974_), .B(_abc_41356_new_n3976_), .Y(_abc_41356_new_n3977_));
AND2X2 AND2X2_177 ( .A(_abc_41356_new_n619_), .B(regfil_4__2_), .Y(_abc_41356_new_n812_));
AND2X2 AND2X2_1770 ( .A(_abc_41356_new_n2072_), .B(_abc_41356_new_n2036_), .Y(_abc_41356_new_n3979_));
AND2X2 AND2X2_1771 ( .A(_abc_41356_new_n3927_), .B(_abc_41356_new_n3980_), .Y(_abc_41356_new_n3981_));
AND2X2 AND2X2_1772 ( .A(_abc_41356_new_n3983_), .B(_abc_41356_new_n2060_), .Y(_abc_41356_new_n3984_));
AND2X2 AND2X2_1773 ( .A(_abc_41356_new_n2035_), .B(_abc_41356_new_n2036_), .Y(_abc_41356_new_n3985_));
AND2X2 AND2X2_1774 ( .A(_abc_41356_new_n3932_), .B(_abc_41356_new_n3980_), .Y(_abc_41356_new_n3986_));
AND2X2 AND2X2_1775 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n3989_), .Y(_abc_41356_new_n3990_));
AND2X2 AND2X2_1776 ( .A(_abc_41356_new_n3990_), .B(intcyc), .Y(_abc_41356_new_n3991_));
AND2X2 AND2X2_1777 ( .A(_abc_41356_new_n3992_), .B(_abc_41356_new_n3993_), .Y(_abc_41356_new_n3994_));
AND2X2 AND2X2_1778 ( .A(_abc_41356_new_n3995_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3996_));
AND2X2 AND2X2_1779 ( .A(_abc_41356_new_n3998_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n3999_));
AND2X2 AND2X2_178 ( .A(_abc_41356_new_n526_), .B(regfil_7__2_), .Y(_abc_41356_new_n813_));
AND2X2 AND2X2_1780 ( .A(_abc_41356_new_n3999_), .B(_abc_41356_new_n3997_), .Y(_abc_41356_new_n4000_));
AND2X2 AND2X2_1781 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n3967_), .Y(_abc_41356_new_n4001_));
AND2X2 AND2X2_1782 ( .A(_abc_41356_new_n4004_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4005_));
AND2X2 AND2X2_1783 ( .A(_abc_41356_new_n4007_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4008_));
AND2X2 AND2X2_1784 ( .A(_abc_41356_new_n3430_), .B(alu_res_5_), .Y(_abc_41356_new_n4009_));
AND2X2 AND2X2_1785 ( .A(_abc_41356_new_n3698_), .B(wdatahold2_5_), .Y(_abc_41356_new_n4010_));
AND2X2 AND2X2_1786 ( .A(_abc_41356_new_n3427_), .B(rdatahold_5_), .Y(_abc_41356_new_n4011_));
AND2X2 AND2X2_1787 ( .A(_abc_41356_new_n4014_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4015_));
AND2X2 AND2X2_1788 ( .A(_abc_41356_new_n3705_), .B(wdatahold_6_), .Y(_abc_41356_new_n4017_));
AND2X2 AND2X2_1789 ( .A(_abc_41356_new_n4018_), .B(wdatahold_6_), .Y(_abc_41356_new_n4019_));
AND2X2 AND2X2_179 ( .A(_abc_41356_new_n808_), .B(_abc_41356_new_n816_), .Y(_abc_41356_new_n817_));
AND2X2 AND2X2_1790 ( .A(_abc_41356_new_n3979_), .B(pc_6_), .Y(_abc_41356_new_n4020_));
AND2X2 AND2X2_1791 ( .A(_abc_41356_new_n4021_), .B(_abc_41356_new_n4022_), .Y(_abc_41356_new_n4023_));
AND2X2 AND2X2_1792 ( .A(_abc_41356_new_n2060_), .B(_abc_41356_new_n4023_), .Y(_abc_41356_new_n4024_));
AND2X2 AND2X2_1793 ( .A(_abc_41356_new_n3985_), .B(pc_6_), .Y(_abc_41356_new_n4025_));
AND2X2 AND2X2_1794 ( .A(_abc_41356_new_n4026_), .B(_abc_41356_new_n4027_), .Y(_abc_41356_new_n4028_));
AND2X2 AND2X2_1795 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n2049_), .Y(_abc_41356_new_n4029_));
AND2X2 AND2X2_1796 ( .A(_abc_41356_new_n4028_), .B(_abc_41356_new_n4030_), .Y(_abc_41356_new_n4031_));
AND2X2 AND2X2_1797 ( .A(_abc_41356_new_n681_), .B(zero), .Y(_abc_41356_new_n4032_));
AND2X2 AND2X2_1798 ( .A(_abc_41356_new_n535_), .B(regfil_5__6_), .Y(_abc_41356_new_n4033_));
AND2X2 AND2X2_1799 ( .A(_abc_41356_new_n4034_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n4035_));
AND2X2 AND2X2_18 ( .A(_abc_41356_new_n526_), .B(_abc_41356_new_n527_), .Y(_abc_41356_new_n528_));
AND2X2 AND2X2_180 ( .A(_abc_41356_new_n817_), .B(_abc_41356_new_n614_), .Y(_abc_41356_new_n818_));
AND2X2 AND2X2_1800 ( .A(_abc_41356_new_n4038_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n4039_));
AND2X2 AND2X2_1801 ( .A(_abc_41356_new_n4037_), .B(_abc_41356_new_n4039_), .Y(_abc_41356_new_n4040_));
AND2X2 AND2X2_1802 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n4033_), .Y(_abc_41356_new_n4041_));
AND2X2 AND2X2_1803 ( .A(pc_6_), .B(intcyc), .Y(_abc_41356_new_n4042_));
AND2X2 AND2X2_1804 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n4042_), .Y(_abc_41356_new_n4043_));
AND2X2 AND2X2_1805 ( .A(_abc_41356_new_n4047_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4048_));
AND2X2 AND2X2_1806 ( .A(_abc_41356_new_n2056_), .B(regfil_7__6_), .Y(_abc_41356_new_n4049_));
AND2X2 AND2X2_1807 ( .A(_abc_41356_new_n4052_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4053_));
AND2X2 AND2X2_1808 ( .A(_abc_41356_new_n4051_), .B(_abc_41356_new_n4053_), .Y(_abc_41356_new_n4054_));
AND2X2 AND2X2_1809 ( .A(_abc_41356_new_n1069_), .B(_abc_41356_new_n3791_), .Y(_abc_41356_new_n4055_));
AND2X2 AND2X2_181 ( .A(_abc_41356_new_n612_), .B(alu_res_2_), .Y(_abc_41356_new_n819_));
AND2X2 AND2X2_1810 ( .A(_abc_41356_new_n4058_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4059_));
AND2X2 AND2X2_1811 ( .A(_abc_41356_new_n3430_), .B(alu_res_6_), .Y(_abc_41356_new_n4060_));
AND2X2 AND2X2_1812 ( .A(_abc_41356_new_n3698_), .B(wdatahold2_6_), .Y(_abc_41356_new_n4061_));
AND2X2 AND2X2_1813 ( .A(_abc_41356_new_n3427_), .B(rdatahold_6_), .Y(_abc_41356_new_n4062_));
AND2X2 AND2X2_1814 ( .A(_abc_41356_new_n4065_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4066_));
AND2X2 AND2X2_1815 ( .A(_abc_41356_new_n3705_), .B(wdatahold_7_), .Y(_abc_41356_new_n4068_));
AND2X2 AND2X2_1816 ( .A(_abc_41356_new_n4069_), .B(_abc_41356_new_n2042_), .Y(_abc_41356_new_n4070_));
AND2X2 AND2X2_1817 ( .A(_abc_41356_new_n4070_), .B(_abc_41356_new_n4030_), .Y(_abc_41356_new_n4071_));
AND2X2 AND2X2_1818 ( .A(_abc_41356_new_n4021_), .B(_abc_41356_new_n4072_), .Y(_abc_41356_new_n4073_));
AND2X2 AND2X2_1819 ( .A(_abc_41356_new_n4075_), .B(_abc_41356_new_n2060_), .Y(_abc_41356_new_n4076_));
AND2X2 AND2X2_182 ( .A(_abc_41356_new_n820_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n821_));
AND2X2 AND2X2_1820 ( .A(_abc_41356_new_n535_), .B(regfil_5__7_), .Y(_abc_41356_new_n4077_));
AND2X2 AND2X2_1821 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n4077_), .Y(_abc_41356_new_n4078_));
AND2X2 AND2X2_1822 ( .A(_abc_41356_new_n681_), .B(sign), .Y(_abc_41356_new_n4079_));
AND2X2 AND2X2_1823 ( .A(_abc_41356_new_n4081_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n4082_));
AND2X2 AND2X2_1824 ( .A(_abc_41356_new_n4084_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n4085_));
AND2X2 AND2X2_1825 ( .A(_abc_41356_new_n4083_), .B(_abc_41356_new_n4085_), .Y(_abc_41356_new_n4086_));
AND2X2 AND2X2_1826 ( .A(pc_7_), .B(intcyc), .Y(_abc_41356_new_n4087_));
AND2X2 AND2X2_1827 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n4087_), .Y(_abc_41356_new_n4088_));
AND2X2 AND2X2_1828 ( .A(_abc_41356_new_n4092_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4093_));
AND2X2 AND2X2_1829 ( .A(_abc_41356_new_n2056_), .B(regfil_7__7_), .Y(_abc_41356_new_n4094_));
AND2X2 AND2X2_183 ( .A(_abc_41356_new_n826_), .B(_abc_41356_new_n724_), .Y(_abc_41356_new_n827_));
AND2X2 AND2X2_1830 ( .A(_abc_41356_new_n4097_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4098_));
AND2X2 AND2X2_1831 ( .A(_abc_41356_new_n4096_), .B(_abc_41356_new_n4098_), .Y(_abc_41356_new_n4099_));
AND2X2 AND2X2_1832 ( .A(_abc_41356_new_n4101_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n4102_));
AND2X2 AND2X2_1833 ( .A(_abc_41356_new_n4100_), .B(_abc_41356_new_n4102_), .Y(_abc_41356_new_n4103_));
AND2X2 AND2X2_1834 ( .A(_abc_41356_new_n3708_), .B(wdatahold_7_), .Y(_abc_41356_new_n4105_));
AND2X2 AND2X2_1835 ( .A(_abc_41356_new_n4107_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4108_));
AND2X2 AND2X2_1836 ( .A(_abc_41356_new_n3430_), .B(alu_res_7_), .Y(_abc_41356_new_n4109_));
AND2X2 AND2X2_1837 ( .A(_abc_41356_new_n3698_), .B(wdatahold2_7_), .Y(_abc_41356_new_n4110_));
AND2X2 AND2X2_1838 ( .A(_abc_41356_new_n3427_), .B(rdatahold_7_), .Y(_abc_41356_new_n4111_));
AND2X2 AND2X2_1839 ( .A(_abc_41356_new_n4114_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4115_));
AND2X2 AND2X2_184 ( .A(_abc_41356_new_n825_), .B(_abc_41356_new_n827_), .Y(_abc_41356_new_n828_));
AND2X2 AND2X2_1840 ( .A(_abc_41356_new_n709_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n4117_));
AND2X2 AND2X2_1841 ( .A(_abc_41356_new_n4119_), .B(_abc_41356_new_n3265_), .Y(_abc_41356_new_n4120_));
AND2X2 AND2X2_1842 ( .A(_abc_41356_new_n4120_), .B(_abc_41356_new_n4118_), .Y(_abc_41356_new_n4121_));
AND2X2 AND2X2_1843 ( .A(_abc_41356_new_n4122_), .B(raddrhold_0_), .Y(_abc_41356_new_n4123_));
AND2X2 AND2X2_1844 ( .A(_abc_41356_new_n4125_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n4126_));
AND2X2 AND2X2_1845 ( .A(_abc_41356_new_n4129_), .B(_abc_41356_new_n2875_), .Y(_abc_41356_new_n4130_));
AND2X2 AND2X2_1846 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1258_), .Y(_abc_41356_new_n4131_));
AND2X2 AND2X2_1847 ( .A(_abc_41356_new_n4132_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4133_));
AND2X2 AND2X2_1848 ( .A(_abc_41356_new_n4133_), .B(_abc_41356_new_n4134_), .Y(_abc_41356_new_n4135_));
AND2X2 AND2X2_1849 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n3723_), .Y(_abc_41356_new_n4136_));
AND2X2 AND2X2_185 ( .A(_abc_41356_new_n512_), .B(_abc_41356_new_n829_), .Y(_abc_41356_new_n830_));
AND2X2 AND2X2_1850 ( .A(_abc_41356_new_n3732_), .B(_abc_41356_new_n4137_), .Y(_abc_41356_new_n4138_));
AND2X2 AND2X2_1851 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n4138_), .Y(_abc_41356_new_n4139_));
AND2X2 AND2X2_1852 ( .A(_abc_41356_new_n4144_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4145_));
AND2X2 AND2X2_1853 ( .A(_abc_41356_new_n4145_), .B(_abc_41356_new_n4142_), .Y(_abc_41356_new_n4146_));
AND2X2 AND2X2_1854 ( .A(_abc_41356_new_n681_), .B(opcode_3_), .Y(_abc_41356_new_n4147_));
AND2X2 AND2X2_1855 ( .A(_abc_41356_new_n3354_), .B(_abc_41356_new_n4147_), .Y(_abc_41356_new_n4148_));
AND2X2 AND2X2_1856 ( .A(_abc_41356_new_n2063_), .B(_abc_41356_new_n4149_), .Y(_abc_41356_new_n4150_));
AND2X2 AND2X2_1857 ( .A(_abc_41356_new_n4151_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n4152_));
AND2X2 AND2X2_1858 ( .A(_abc_41356_new_n4154_), .B(_abc_41356_new_n4150_), .Y(_abc_41356_new_n4155_));
AND2X2 AND2X2_1859 ( .A(_abc_41356_new_n3353_), .B(_abc_41356_new_n3362_), .Y(_abc_41356_new_n4156_));
AND2X2 AND2X2_186 ( .A(_abc_41356_new_n555_), .B(regfil_7__1_), .Y(_abc_41356_new_n832_));
AND2X2 AND2X2_1860 ( .A(_abc_41356_new_n3354_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n4157_));
AND2X2 AND2X2_1861 ( .A(_abc_41356_new_n4157_), .B(_abc_41356_new_n2994_), .Y(_abc_41356_new_n4158_));
AND2X2 AND2X2_1862 ( .A(_abc_41356_new_n4160_), .B(_abc_41356_new_n4161_), .Y(_abc_41356_new_n4162_));
AND2X2 AND2X2_1863 ( .A(_abc_41356_new_n4163_), .B(_abc_41356_new_n4157_), .Y(_abc_41356_new_n4164_));
AND2X2 AND2X2_1864 ( .A(_abc_41356_new_n4165_), .B(_abc_41356_new_n4159_), .Y(_abc_41356_new_n4166_));
AND2X2 AND2X2_1865 ( .A(_abc_41356_new_n4166_), .B(_abc_41356_new_n4156_), .Y(_abc_41356_new_n4167_));
AND2X2 AND2X2_1866 ( .A(_abc_41356_new_n4167_), .B(_abc_41356_new_n4155_), .Y(_abc_41356_new_n4168_));
AND2X2 AND2X2_1867 ( .A(_abc_41356_new_n3379_), .B(_abc_41356_new_n3358_), .Y(_abc_41356_new_n4169_));
AND2X2 AND2X2_1868 ( .A(_abc_41356_new_n4169_), .B(_abc_41356_new_n3494_), .Y(_abc_41356_new_n4170_));
AND2X2 AND2X2_1869 ( .A(_abc_41356_new_n4170_), .B(_abc_41356_new_n4168_), .Y(_abc_41356_new_n4171_));
AND2X2 AND2X2_187 ( .A(_abc_41356_new_n551_), .B(regfil_7__1_), .Y(_abc_41356_new_n833_));
AND2X2 AND2X2_1870 ( .A(_abc_41356_new_n4171_), .B(raddrhold_0_), .Y(_abc_41356_new_n4172_));
AND2X2 AND2X2_1871 ( .A(_abc_41356_new_n4173_), .B(sp_0_), .Y(_abc_41356_new_n4174_));
AND2X2 AND2X2_1872 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n3723_), .Y(_abc_41356_new_n4176_));
AND2X2 AND2X2_1873 ( .A(_abc_41356_new_n4178_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4179_));
AND2X2 AND2X2_1874 ( .A(_abc_41356_new_n677_), .B(regfil_5__0_), .Y(_abc_41356_new_n4180_));
AND2X2 AND2X2_1875 ( .A(_abc_41356_new_n678_), .B(raddrhold_0_), .Y(_abc_41356_new_n4181_));
AND2X2 AND2X2_1876 ( .A(_abc_41356_new_n677_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n4183_));
AND2X2 AND2X2_1877 ( .A(_abc_41356_new_n4183_), .B(_abc_41356_new_n682_), .Y(_abc_41356_new_n4184_));
AND2X2 AND2X2_1878 ( .A(_abc_41356_new_n4185_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n4186_));
AND2X2 AND2X2_1879 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4182_), .Y(_abc_41356_new_n4187_));
AND2X2 AND2X2_188 ( .A(_abc_41356_new_n834_), .B(_abc_41356_new_n540_), .Y(_abc_41356_new_n835_));
AND2X2 AND2X2_1880 ( .A(_abc_41356_new_n4182_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4188_));
AND2X2 AND2X2_1881 ( .A(_abc_41356_new_n4184_), .B(raddrhold_0_), .Y(_abc_41356_new_n4189_));
AND2X2 AND2X2_1882 ( .A(_abc_41356_new_n4193_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4194_));
AND2X2 AND2X2_1883 ( .A(_abc_41356_new_n3424_), .B(rdatahold2_0_), .Y(_abc_41356_new_n4195_));
AND2X2 AND2X2_1884 ( .A(_abc_41356_new_n4117_), .B(_abc_41356_new_n4196_), .Y(_abc_41356_new_n4197_));
AND2X2 AND2X2_1885 ( .A(_abc_41356_new_n4199_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4200_));
AND2X2 AND2X2_1886 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1259_), .Y(_abc_41356_new_n4202_));
AND2X2 AND2X2_1887 ( .A(_abc_41356_new_n4204_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4205_));
AND2X2 AND2X2_1888 ( .A(_abc_41356_new_n4205_), .B(_abc_41356_new_n4203_), .Y(_abc_41356_new_n4206_));
AND2X2 AND2X2_1889 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n3762_), .Y(_abc_41356_new_n4207_));
AND2X2 AND2X2_189 ( .A(_abc_41356_new_n833_), .B(regfil_7__2_), .Y(_abc_41356_new_n836_));
AND2X2 AND2X2_1890 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n4208_), .Y(_abc_41356_new_n4209_));
AND2X2 AND2X2_1891 ( .A(_abc_41356_new_n4213_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4214_));
AND2X2 AND2X2_1892 ( .A(_abc_41356_new_n4214_), .B(_abc_41356_new_n4212_), .Y(_abc_41356_new_n4215_));
AND2X2 AND2X2_1893 ( .A(_abc_41356_new_n4171_), .B(raddrhold_1_), .Y(_abc_41356_new_n4216_));
AND2X2 AND2X2_1894 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n3762_), .Y(_abc_41356_new_n4217_));
AND2X2 AND2X2_1895 ( .A(_abc_41356_new_n4173_), .B(sp_1_), .Y(_abc_41356_new_n4218_));
AND2X2 AND2X2_1896 ( .A(_abc_41356_new_n4220_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4221_));
AND2X2 AND2X2_1897 ( .A(_abc_41356_new_n677_), .B(regfil_5__1_), .Y(_abc_41356_new_n4222_));
AND2X2 AND2X2_1898 ( .A(_abc_41356_new_n678_), .B(raddrhold_1_), .Y(_abc_41356_new_n4223_));
AND2X2 AND2X2_1899 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4224_), .Y(_abc_41356_new_n4225_));
AND2X2 AND2X2_19 ( .A(_abc_41356_new_n528_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n529_));
AND2X2 AND2X2_190 ( .A(_abc_41356_new_n837_), .B(_abc_41356_new_n698_), .Y(_abc_41356_new_n838_));
AND2X2 AND2X2_1900 ( .A(_abc_41356_new_n4224_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4226_));
AND2X2 AND2X2_1901 ( .A(_abc_41356_new_n4184_), .B(raddrhold_1_), .Y(_abc_41356_new_n4227_));
AND2X2 AND2X2_1902 ( .A(_abc_41356_new_n4231_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4232_));
AND2X2 AND2X2_1903 ( .A(_abc_41356_new_n3424_), .B(rdatahold2_1_), .Y(_abc_41356_new_n4233_));
AND2X2 AND2X2_1904 ( .A(_abc_41356_new_n4234_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4235_));
AND2X2 AND2X2_1905 ( .A(_abc_41356_new_n4122_), .B(raddrhold_1_), .Y(_abc_41356_new_n4236_));
AND2X2 AND2X2_1906 ( .A(raddrhold_0_), .B(raddrhold_1_), .Y(_abc_41356_new_n4238_));
AND2X2 AND2X2_1907 ( .A(_abc_41356_new_n4239_), .B(_abc_41356_new_n4237_), .Y(_abc_41356_new_n4240_));
AND2X2 AND2X2_1908 ( .A(_abc_41356_new_n709_), .B(_abc_41356_new_n607_), .Y(_abc_41356_new_n4241_));
AND2X2 AND2X2_1909 ( .A(_abc_41356_new_n4241_), .B(_abc_41356_new_n4240_), .Y(_abc_41356_new_n4242_));
AND2X2 AND2X2_191 ( .A(_abc_41356_new_n530_), .B(regfil_7__3_), .Y(_abc_41356_new_n840_));
AND2X2 AND2X2_1910 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1257_), .Y(_abc_41356_new_n4245_));
AND2X2 AND2X2_1911 ( .A(_abc_41356_new_n4246_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4247_));
AND2X2 AND2X2_1912 ( .A(_abc_41356_new_n4247_), .B(_abc_41356_new_n4248_), .Y(_abc_41356_new_n4249_));
AND2X2 AND2X2_1913 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n3814_), .Y(_abc_41356_new_n4250_));
AND2X2 AND2X2_1914 ( .A(_abc_41356_new_n3827_), .B(_abc_41356_new_n4251_), .Y(_abc_41356_new_n4252_));
AND2X2 AND2X2_1915 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n4252_), .Y(_abc_41356_new_n4253_));
AND2X2 AND2X2_1916 ( .A(_abc_41356_new_n4257_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4258_));
AND2X2 AND2X2_1917 ( .A(_abc_41356_new_n4258_), .B(_abc_41356_new_n4256_), .Y(_abc_41356_new_n4259_));
AND2X2 AND2X2_1918 ( .A(_abc_41356_new_n4171_), .B(raddrhold_2_), .Y(_abc_41356_new_n4260_));
AND2X2 AND2X2_1919 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n3814_), .Y(_abc_41356_new_n4261_));
AND2X2 AND2X2_192 ( .A(_abc_41356_new_n842_), .B(_abc_41356_new_n831_), .Y(_abc_41356_new_n843_));
AND2X2 AND2X2_1920 ( .A(_abc_41356_new_n4173_), .B(sp_2_), .Y(_abc_41356_new_n4262_));
AND2X2 AND2X2_1921 ( .A(_abc_41356_new_n4264_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4265_));
AND2X2 AND2X2_1922 ( .A(_abc_41356_new_n677_), .B(regfil_5__2_), .Y(_abc_41356_new_n4266_));
AND2X2 AND2X2_1923 ( .A(_abc_41356_new_n678_), .B(raddrhold_2_), .Y(_abc_41356_new_n4267_));
AND2X2 AND2X2_1924 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4268_), .Y(_abc_41356_new_n4269_));
AND2X2 AND2X2_1925 ( .A(_abc_41356_new_n4268_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4270_));
AND2X2 AND2X2_1926 ( .A(_abc_41356_new_n4184_), .B(raddrhold_2_), .Y(_abc_41356_new_n4271_));
AND2X2 AND2X2_1927 ( .A(_abc_41356_new_n4275_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4276_));
AND2X2 AND2X2_1928 ( .A(_abc_41356_new_n3424_), .B(rdatahold2_2_), .Y(_abc_41356_new_n4277_));
AND2X2 AND2X2_1929 ( .A(_abc_41356_new_n4278_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4279_));
AND2X2 AND2X2_193 ( .A(_abc_41356_new_n712_), .B(regfil_7__2_), .Y(_abc_41356_new_n844_));
AND2X2 AND2X2_1930 ( .A(_abc_41356_new_n4122_), .B(raddrhold_2_), .Y(_abc_41356_new_n4280_));
AND2X2 AND2X2_1931 ( .A(_abc_41356_new_n4238_), .B(raddrhold_2_), .Y(_abc_41356_new_n4282_));
AND2X2 AND2X2_1932 ( .A(_abc_41356_new_n4283_), .B(_abc_41356_new_n4281_), .Y(_abc_41356_new_n4284_));
AND2X2 AND2X2_1933 ( .A(_abc_41356_new_n4241_), .B(_abc_41356_new_n4284_), .Y(_abc_41356_new_n4285_));
AND2X2 AND2X2_1934 ( .A(_abc_41356_new_n4122_), .B(raddrhold_3_), .Y(_abc_41356_new_n4288_));
AND2X2 AND2X2_1935 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1256_), .Y(_abc_41356_new_n4289_));
AND2X2 AND2X2_1936 ( .A(_abc_41356_new_n4290_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4291_));
AND2X2 AND2X2_1937 ( .A(_abc_41356_new_n4291_), .B(_abc_41356_new_n4292_), .Y(_abc_41356_new_n4293_));
AND2X2 AND2X2_1938 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n3879_), .Y(_abc_41356_new_n4294_));
AND2X2 AND2X2_1939 ( .A(_abc_41356_new_n3889_), .B(_abc_41356_new_n4295_), .Y(_abc_41356_new_n4296_));
AND2X2 AND2X2_194 ( .A(_abc_41356_new_n714_), .B(alu_res_2_), .Y(_abc_41356_new_n845_));
AND2X2 AND2X2_1940 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n4296_), .Y(_abc_41356_new_n4297_));
AND2X2 AND2X2_1941 ( .A(_abc_41356_new_n4301_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4302_));
AND2X2 AND2X2_1942 ( .A(_abc_41356_new_n4302_), .B(_abc_41356_new_n4300_), .Y(_abc_41356_new_n4303_));
AND2X2 AND2X2_1943 ( .A(_abc_41356_new_n4171_), .B(raddrhold_3_), .Y(_abc_41356_new_n4304_));
AND2X2 AND2X2_1944 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n3879_), .Y(_abc_41356_new_n4305_));
AND2X2 AND2X2_1945 ( .A(_abc_41356_new_n4173_), .B(sp_3_), .Y(_abc_41356_new_n4306_));
AND2X2 AND2X2_1946 ( .A(_abc_41356_new_n4308_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4309_));
AND2X2 AND2X2_1947 ( .A(_abc_41356_new_n677_), .B(regfil_5__3_), .Y(_abc_41356_new_n4310_));
AND2X2 AND2X2_1948 ( .A(_abc_41356_new_n678_), .B(raddrhold_3_), .Y(_abc_41356_new_n4311_));
AND2X2 AND2X2_1949 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4312_), .Y(_abc_41356_new_n4313_));
AND2X2 AND2X2_195 ( .A(_abc_41356_new_n718_), .B(\data[2] ), .Y(_abc_41356_new_n846_));
AND2X2 AND2X2_1950 ( .A(_abc_41356_new_n4312_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4314_));
AND2X2 AND2X2_1951 ( .A(_abc_41356_new_n4184_), .B(raddrhold_3_), .Y(_abc_41356_new_n4315_));
AND2X2 AND2X2_1952 ( .A(_abc_41356_new_n4319_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4320_));
AND2X2 AND2X2_1953 ( .A(_abc_41356_new_n4282_), .B(raddrhold_3_), .Y(_abc_41356_new_n4321_));
AND2X2 AND2X2_1954 ( .A(_abc_41356_new_n4117_), .B(_abc_41356_new_n4323_), .Y(_abc_41356_new_n4324_));
AND2X2 AND2X2_1955 ( .A(_abc_41356_new_n4324_), .B(_abc_41356_new_n4322_), .Y(_abc_41356_new_n4325_));
AND2X2 AND2X2_1956 ( .A(_abc_41356_new_n3424_), .B(rdatahold2_3_), .Y(_abc_41356_new_n4326_));
AND2X2 AND2X2_1957 ( .A(_abc_41356_new_n4328_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4329_));
AND2X2 AND2X2_1958 ( .A(_abc_41356_new_n4122_), .B(raddrhold_4_), .Y(_abc_41356_new_n4331_));
AND2X2 AND2X2_1959 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1255_), .Y(_abc_41356_new_n4332_));
AND2X2 AND2X2_196 ( .A(_abc_41356_new_n790_), .B(regfil_0__3_), .Y(_abc_41356_new_n853_));
AND2X2 AND2X2_1960 ( .A(_abc_41356_new_n4333_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4334_));
AND2X2 AND2X2_1961 ( .A(_abc_41356_new_n4334_), .B(_abc_41356_new_n4335_), .Y(_abc_41356_new_n4336_));
AND2X2 AND2X2_1962 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n3929_), .Y(_abc_41356_new_n4337_));
AND2X2 AND2X2_1963 ( .A(_abc_41356_new_n3942_), .B(_abc_41356_new_n4338_), .Y(_abc_41356_new_n4339_));
AND2X2 AND2X2_1964 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n4339_), .Y(_abc_41356_new_n4340_));
AND2X2 AND2X2_1965 ( .A(_abc_41356_new_n4344_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4345_));
AND2X2 AND2X2_1966 ( .A(_abc_41356_new_n4345_), .B(_abc_41356_new_n4343_), .Y(_abc_41356_new_n4346_));
AND2X2 AND2X2_1967 ( .A(_abc_41356_new_n4171_), .B(raddrhold_4_), .Y(_abc_41356_new_n4347_));
AND2X2 AND2X2_1968 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n3929_), .Y(_abc_41356_new_n4348_));
AND2X2 AND2X2_1969 ( .A(_abc_41356_new_n4173_), .B(sp_4_), .Y(_abc_41356_new_n4349_));
AND2X2 AND2X2_197 ( .A(_abc_41356_new_n854_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n855_));
AND2X2 AND2X2_1970 ( .A(_abc_41356_new_n4351_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4352_));
AND2X2 AND2X2_1971 ( .A(_abc_41356_new_n677_), .B(regfil_5__4_), .Y(_abc_41356_new_n4353_));
AND2X2 AND2X2_1972 ( .A(_abc_41356_new_n678_), .B(raddrhold_4_), .Y(_abc_41356_new_n4354_));
AND2X2 AND2X2_1973 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4355_), .Y(_abc_41356_new_n4356_));
AND2X2 AND2X2_1974 ( .A(_abc_41356_new_n4355_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4357_));
AND2X2 AND2X2_1975 ( .A(_abc_41356_new_n4184_), .B(raddrhold_4_), .Y(_abc_41356_new_n4358_));
AND2X2 AND2X2_1976 ( .A(_abc_41356_new_n4362_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4363_));
AND2X2 AND2X2_1977 ( .A(_abc_41356_new_n4321_), .B(raddrhold_4_), .Y(_abc_41356_new_n4364_));
AND2X2 AND2X2_1978 ( .A(_abc_41356_new_n4366_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4367_));
AND2X2 AND2X2_1979 ( .A(_abc_41356_new_n4367_), .B(_abc_41356_new_n4365_), .Y(_abc_41356_new_n4368_));
AND2X2 AND2X2_198 ( .A(_abc_41356_new_n796_), .B(regfil_0__3_), .Y(_abc_41356_new_n857_));
AND2X2 AND2X2_1980 ( .A(_abc_41356_new_n3424_), .B(rdatahold2_4_), .Y(_abc_41356_new_n4369_));
AND2X2 AND2X2_1981 ( .A(_abc_41356_new_n4371_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4372_));
AND2X2 AND2X2_1982 ( .A(_abc_41356_new_n4122_), .B(raddrhold_5_), .Y(_abc_41356_new_n4374_));
AND2X2 AND2X2_1983 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1254_), .Y(_abc_41356_new_n4375_));
AND2X2 AND2X2_1984 ( .A(_abc_41356_new_n4376_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4377_));
AND2X2 AND2X2_1985 ( .A(_abc_41356_new_n4377_), .B(_abc_41356_new_n4378_), .Y(_abc_41356_new_n4379_));
AND2X2 AND2X2_1986 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n3983_), .Y(_abc_41356_new_n4380_));
AND2X2 AND2X2_1987 ( .A(_abc_41356_new_n3995_), .B(_abc_41356_new_n4381_), .Y(_abc_41356_new_n4382_));
AND2X2 AND2X2_1988 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n4382_), .Y(_abc_41356_new_n4383_));
AND2X2 AND2X2_1989 ( .A(_abc_41356_new_n4387_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4388_));
AND2X2 AND2X2_199 ( .A(_abc_41356_new_n858_), .B(_abc_41356_new_n581_), .Y(_abc_41356_new_n859_));
AND2X2 AND2X2_1990 ( .A(_abc_41356_new_n4388_), .B(_abc_41356_new_n4386_), .Y(_abc_41356_new_n4389_));
AND2X2 AND2X2_1991 ( .A(_abc_41356_new_n4171_), .B(raddrhold_5_), .Y(_abc_41356_new_n4390_));
AND2X2 AND2X2_1992 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n3983_), .Y(_abc_41356_new_n4391_));
AND2X2 AND2X2_1993 ( .A(_abc_41356_new_n4173_), .B(sp_5_), .Y(_abc_41356_new_n4392_));
AND2X2 AND2X2_1994 ( .A(_abc_41356_new_n4394_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4395_));
AND2X2 AND2X2_1995 ( .A(_abc_41356_new_n677_), .B(regfil_5__5_), .Y(_abc_41356_new_n4396_));
AND2X2 AND2X2_1996 ( .A(_abc_41356_new_n678_), .B(raddrhold_5_), .Y(_abc_41356_new_n4397_));
AND2X2 AND2X2_1997 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4398_), .Y(_abc_41356_new_n4399_));
AND2X2 AND2X2_1998 ( .A(_abc_41356_new_n4398_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4400_));
AND2X2 AND2X2_1999 ( .A(_abc_41356_new_n4184_), .B(raddrhold_5_), .Y(_abc_41356_new_n4401_));
AND2X2 AND2X2_2 ( .A(_abc_41356_new_n503_), .B(state_2_), .Y(_abc_41356_new_n504_));
AND2X2 AND2X2_20 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n529_), .Y(_abc_41356_new_n530_));
AND2X2 AND2X2_200 ( .A(_abc_41356_new_n859_), .B(_abc_41356_new_n856_), .Y(_abc_41356_new_n860_));
AND2X2 AND2X2_2000 ( .A(_abc_41356_new_n4405_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4406_));
AND2X2 AND2X2_2001 ( .A(_abc_41356_new_n4364_), .B(raddrhold_5_), .Y(_abc_41356_new_n4407_));
AND2X2 AND2X2_2002 ( .A(_abc_41356_new_n4409_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4410_));
AND2X2 AND2X2_2003 ( .A(_abc_41356_new_n4410_), .B(_abc_41356_new_n4408_), .Y(_abc_41356_new_n4411_));
AND2X2 AND2X2_2004 ( .A(_abc_41356_new_n3424_), .B(rdatahold2_5_), .Y(_abc_41356_new_n4412_));
AND2X2 AND2X2_2005 ( .A(_abc_41356_new_n4414_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4415_));
AND2X2 AND2X2_2006 ( .A(_abc_41356_new_n4122_), .B(raddrhold_6_), .Y(_abc_41356_new_n4417_));
AND2X2 AND2X2_2007 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1253_), .Y(_abc_41356_new_n4418_));
AND2X2 AND2X2_2008 ( .A(_abc_41356_new_n4419_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4420_));
AND2X2 AND2X2_2009 ( .A(_abc_41356_new_n4421_), .B(raddrhold_6_), .Y(_abc_41356_new_n4422_));
AND2X2 AND2X2_201 ( .A(_abc_41356_new_n642_), .B(rdatahold_3_), .Y(_abc_41356_new_n861_));
AND2X2 AND2X2_2010 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n4023_), .Y(_abc_41356_new_n4423_));
AND2X2 AND2X2_2011 ( .A(_abc_41356_new_n4034_), .B(_abc_41356_new_n4424_), .Y(_abc_41356_new_n4425_));
AND2X2 AND2X2_2012 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n4425_), .Y(_abc_41356_new_n4426_));
AND2X2 AND2X2_2013 ( .A(_abc_41356_new_n4420_), .B(_abc_41356_new_n682_), .Y(_abc_41356_new_n4427_));
AND2X2 AND2X2_2014 ( .A(_abc_41356_new_n4430_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4431_));
AND2X2 AND2X2_2015 ( .A(_abc_41356_new_n4171_), .B(raddrhold_6_), .Y(_abc_41356_new_n4432_));
AND2X2 AND2X2_2016 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n4023_), .Y(_abc_41356_new_n4433_));
AND2X2 AND2X2_2017 ( .A(_abc_41356_new_n4173_), .B(sp_6_), .Y(_abc_41356_new_n4434_));
AND2X2 AND2X2_2018 ( .A(_abc_41356_new_n4436_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4437_));
AND2X2 AND2X2_2019 ( .A(_abc_41356_new_n677_), .B(regfil_5__6_), .Y(_abc_41356_new_n4438_));
AND2X2 AND2X2_202 ( .A(_abc_41356_new_n619_), .B(regfil_4__3_), .Y(_abc_41356_new_n862_));
AND2X2 AND2X2_2020 ( .A(_abc_41356_new_n678_), .B(raddrhold_6_), .Y(_abc_41356_new_n4439_));
AND2X2 AND2X2_2021 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4440_), .Y(_abc_41356_new_n4441_));
AND2X2 AND2X2_2022 ( .A(_abc_41356_new_n4440_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4442_));
AND2X2 AND2X2_2023 ( .A(_abc_41356_new_n4184_), .B(raddrhold_6_), .Y(_abc_41356_new_n4443_));
AND2X2 AND2X2_2024 ( .A(_abc_41356_new_n4447_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4448_));
AND2X2 AND2X2_2025 ( .A(_abc_41356_new_n4407_), .B(raddrhold_6_), .Y(_abc_41356_new_n4449_));
AND2X2 AND2X2_2026 ( .A(_abc_41356_new_n4451_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4452_));
AND2X2 AND2X2_2027 ( .A(_abc_41356_new_n4452_), .B(_abc_41356_new_n4450_), .Y(_abc_41356_new_n4453_));
AND2X2 AND2X2_2028 ( .A(_abc_41356_new_n3424_), .B(rdatahold2_6_), .Y(_abc_41356_new_n4454_));
AND2X2 AND2X2_2029 ( .A(_abc_41356_new_n4456_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4457_));
AND2X2 AND2X2_203 ( .A(_abc_41356_new_n616_), .B(regfil_5__3_), .Y(_abc_41356_new_n863_));
AND2X2 AND2X2_2030 ( .A(_abc_41356_new_n4122_), .B(raddrhold_7_), .Y(_abc_41356_new_n4459_));
AND2X2 AND2X2_2031 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1252_), .Y(_abc_41356_new_n4460_));
AND2X2 AND2X2_2032 ( .A(_abc_41356_new_n4461_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4462_));
AND2X2 AND2X2_2033 ( .A(_abc_41356_new_n4462_), .B(_abc_41356_new_n4463_), .Y(_abc_41356_new_n4464_));
AND2X2 AND2X2_2034 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n4075_), .Y(_abc_41356_new_n4465_));
AND2X2 AND2X2_2035 ( .A(_abc_41356_new_n4081_), .B(_abc_41356_new_n4466_), .Y(_abc_41356_new_n4467_));
AND2X2 AND2X2_2036 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n4467_), .Y(_abc_41356_new_n4468_));
AND2X2 AND2X2_2037 ( .A(_abc_41356_new_n4472_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4473_));
AND2X2 AND2X2_2038 ( .A(_abc_41356_new_n4473_), .B(_abc_41356_new_n4471_), .Y(_abc_41356_new_n4474_));
AND2X2 AND2X2_2039 ( .A(_abc_41356_new_n4171_), .B(raddrhold_7_), .Y(_abc_41356_new_n4475_));
AND2X2 AND2X2_204 ( .A(_abc_41356_new_n526_), .B(regfil_7__3_), .Y(_abc_41356_new_n865_));
AND2X2 AND2X2_2040 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n4075_), .Y(_abc_41356_new_n4476_));
AND2X2 AND2X2_2041 ( .A(_abc_41356_new_n4173_), .B(sp_7_), .Y(_abc_41356_new_n4477_));
AND2X2 AND2X2_2042 ( .A(_abc_41356_new_n4479_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4480_));
AND2X2 AND2X2_2043 ( .A(_abc_41356_new_n677_), .B(regfil_5__7_), .Y(_abc_41356_new_n4481_));
AND2X2 AND2X2_2044 ( .A(_abc_41356_new_n678_), .B(raddrhold_7_), .Y(_abc_41356_new_n4482_));
AND2X2 AND2X2_2045 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4483_), .Y(_abc_41356_new_n4484_));
AND2X2 AND2X2_2046 ( .A(_abc_41356_new_n4483_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4485_));
AND2X2 AND2X2_2047 ( .A(_abc_41356_new_n4184_), .B(raddrhold_7_), .Y(_abc_41356_new_n4486_));
AND2X2 AND2X2_2048 ( .A(_abc_41356_new_n4490_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4491_));
AND2X2 AND2X2_2049 ( .A(_abc_41356_new_n4449_), .B(raddrhold_7_), .Y(_abc_41356_new_n4492_));
AND2X2 AND2X2_205 ( .A(_abc_41356_new_n623_), .B(regfil_6__3_), .Y(_abc_41356_new_n866_));
AND2X2 AND2X2_2050 ( .A(_abc_41356_new_n4494_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4495_));
AND2X2 AND2X2_2051 ( .A(_abc_41356_new_n4495_), .B(_abc_41356_new_n4493_), .Y(_abc_41356_new_n4496_));
AND2X2 AND2X2_2052 ( .A(_abc_41356_new_n3424_), .B(rdatahold2_7_), .Y(_abc_41356_new_n4497_));
AND2X2 AND2X2_2053 ( .A(_abc_41356_new_n4499_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4500_));
AND2X2 AND2X2_2054 ( .A(_abc_41356_new_n4122_), .B(raddrhold_8_), .Y(_abc_41356_new_n4502_));
AND2X2 AND2X2_2055 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1251_), .Y(_abc_41356_new_n4503_));
AND2X2 AND2X2_2056 ( .A(_abc_41356_new_n4504_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4505_));
AND2X2 AND2X2_2057 ( .A(_abc_41356_new_n4505_), .B(_abc_41356_new_n4506_), .Y(_abc_41356_new_n4507_));
AND2X2 AND2X2_2058 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n2078_), .Y(_abc_41356_new_n4508_));
AND2X2 AND2X2_2059 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n2086_), .Y(_abc_41356_new_n4509_));
AND2X2 AND2X2_206 ( .A(_abc_41356_new_n619_), .B(regfil_0__3_), .Y(_abc_41356_new_n870_));
AND2X2 AND2X2_2060 ( .A(_abc_41356_new_n4513_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4514_));
AND2X2 AND2X2_2061 ( .A(_abc_41356_new_n4514_), .B(_abc_41356_new_n4512_), .Y(_abc_41356_new_n4515_));
AND2X2 AND2X2_2062 ( .A(_abc_41356_new_n4171_), .B(raddrhold_8_), .Y(_abc_41356_new_n4516_));
AND2X2 AND2X2_2063 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n2078_), .Y(_abc_41356_new_n4517_));
AND2X2 AND2X2_2064 ( .A(_abc_41356_new_n4173_), .B(sp_8_), .Y(_abc_41356_new_n4518_));
AND2X2 AND2X2_2065 ( .A(_abc_41356_new_n4520_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4521_));
AND2X2 AND2X2_2066 ( .A(_abc_41356_new_n677_), .B(regfil_4__0_), .Y(_abc_41356_new_n4522_));
AND2X2 AND2X2_2067 ( .A(_abc_41356_new_n678_), .B(raddrhold_8_), .Y(_abc_41356_new_n4523_));
AND2X2 AND2X2_2068 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4524_), .Y(_abc_41356_new_n4525_));
AND2X2 AND2X2_2069 ( .A(_abc_41356_new_n4524_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4526_));
AND2X2 AND2X2_207 ( .A(_abc_41356_new_n616_), .B(regfil_1__3_), .Y(_abc_41356_new_n871_));
AND2X2 AND2X2_2070 ( .A(_abc_41356_new_n4184_), .B(raddrhold_8_), .Y(_abc_41356_new_n4527_));
AND2X2 AND2X2_2071 ( .A(_abc_41356_new_n4531_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4532_));
AND2X2 AND2X2_2072 ( .A(_abc_41356_new_n4492_), .B(raddrhold_8_), .Y(_abc_41356_new_n4533_));
AND2X2 AND2X2_2073 ( .A(_abc_41356_new_n4535_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4536_));
AND2X2 AND2X2_2074 ( .A(_abc_41356_new_n4536_), .B(_abc_41356_new_n4534_), .Y(_abc_41356_new_n4537_));
AND2X2 AND2X2_2075 ( .A(_abc_41356_new_n3424_), .B(rdatahold_0_), .Y(_abc_41356_new_n4538_));
AND2X2 AND2X2_2076 ( .A(_abc_41356_new_n4540_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4541_));
AND2X2 AND2X2_2077 ( .A(_abc_41356_new_n4122_), .B(raddrhold_9_), .Y(_abc_41356_new_n4543_));
AND2X2 AND2X2_2078 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1504_), .Y(_abc_41356_new_n4544_));
AND2X2 AND2X2_2079 ( .A(_abc_41356_new_n4545_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4546_));
AND2X2 AND2X2_208 ( .A(_abc_41356_new_n526_), .B(regfil_3__3_), .Y(_abc_41356_new_n873_));
AND2X2 AND2X2_2080 ( .A(_abc_41356_new_n4546_), .B(_abc_41356_new_n4547_), .Y(_abc_41356_new_n4548_));
AND2X2 AND2X2_2081 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n2119_), .Y(_abc_41356_new_n4549_));
AND2X2 AND2X2_2082 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n2127_), .Y(_abc_41356_new_n4550_));
AND2X2 AND2X2_2083 ( .A(_abc_41356_new_n4554_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4555_));
AND2X2 AND2X2_2084 ( .A(_abc_41356_new_n4555_), .B(_abc_41356_new_n4553_), .Y(_abc_41356_new_n4556_));
AND2X2 AND2X2_2085 ( .A(_abc_41356_new_n4171_), .B(raddrhold_9_), .Y(_abc_41356_new_n4557_));
AND2X2 AND2X2_2086 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n2119_), .Y(_abc_41356_new_n4558_));
AND2X2 AND2X2_2087 ( .A(_abc_41356_new_n4173_), .B(sp_9_), .Y(_abc_41356_new_n4559_));
AND2X2 AND2X2_2088 ( .A(_abc_41356_new_n4561_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4562_));
AND2X2 AND2X2_2089 ( .A(_abc_41356_new_n677_), .B(regfil_4__1_), .Y(_abc_41356_new_n4563_));
AND2X2 AND2X2_209 ( .A(_abc_41356_new_n623_), .B(regfil_2__3_), .Y(_abc_41356_new_n874_));
AND2X2 AND2X2_2090 ( .A(_abc_41356_new_n678_), .B(raddrhold_9_), .Y(_abc_41356_new_n4564_));
AND2X2 AND2X2_2091 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4565_), .Y(_abc_41356_new_n4566_));
AND2X2 AND2X2_2092 ( .A(_abc_41356_new_n4565_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4567_));
AND2X2 AND2X2_2093 ( .A(_abc_41356_new_n4184_), .B(raddrhold_9_), .Y(_abc_41356_new_n4568_));
AND2X2 AND2X2_2094 ( .A(_abc_41356_new_n4572_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4573_));
AND2X2 AND2X2_2095 ( .A(_abc_41356_new_n4533_), .B(raddrhold_9_), .Y(_abc_41356_new_n4574_));
AND2X2 AND2X2_2096 ( .A(_abc_41356_new_n4576_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4577_));
AND2X2 AND2X2_2097 ( .A(_abc_41356_new_n4577_), .B(_abc_41356_new_n4575_), .Y(_abc_41356_new_n4578_));
AND2X2 AND2X2_2098 ( .A(_abc_41356_new_n3424_), .B(rdatahold_1_), .Y(_abc_41356_new_n4579_));
AND2X2 AND2X2_2099 ( .A(_abc_41356_new_n4581_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4582_));
AND2X2 AND2X2_21 ( .A(_abc_41356_new_n530_), .B(_abc_41356_new_n513_), .Y(_abc_41356_new_n531_));
AND2X2 AND2X2_210 ( .A(_abc_41356_new_n869_), .B(_abc_41356_new_n877_), .Y(_abc_41356_new_n878_));
AND2X2 AND2X2_2100 ( .A(_abc_41356_new_n4122_), .B(raddrhold_10_), .Y(_abc_41356_new_n4584_));
AND2X2 AND2X2_2101 ( .A(_abc_41356_new_n4171_), .B(raddrhold_10_), .Y(_abc_41356_new_n4585_));
AND2X2 AND2X2_2102 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n2160_), .Y(_abc_41356_new_n4586_));
AND2X2 AND2X2_2103 ( .A(_abc_41356_new_n4173_), .B(sp_10_), .Y(_abc_41356_new_n4587_));
AND2X2 AND2X2_2104 ( .A(_abc_41356_new_n4589_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4590_));
AND2X2 AND2X2_2105 ( .A(_abc_41356_new_n2160_), .B(_abc_41356_new_n4127_), .Y(_abc_41356_new_n4591_));
AND2X2 AND2X2_2106 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1580_), .Y(_abc_41356_new_n4592_));
AND2X2 AND2X2_2107 ( .A(_abc_41356_new_n4594_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4595_));
AND2X2 AND2X2_2108 ( .A(_abc_41356_new_n4595_), .B(_abc_41356_new_n4593_), .Y(_abc_41356_new_n4596_));
AND2X2 AND2X2_2109 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n2165_), .Y(_abc_41356_new_n4597_));
AND2X2 AND2X2_211 ( .A(_abc_41356_new_n878_), .B(_abc_41356_new_n614_), .Y(_abc_41356_new_n879_));
AND2X2 AND2X2_2110 ( .A(_abc_41356_new_n4601_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4602_));
AND2X2 AND2X2_2111 ( .A(_abc_41356_new_n4602_), .B(_abc_41356_new_n4600_), .Y(_abc_41356_new_n4603_));
AND2X2 AND2X2_2112 ( .A(_abc_41356_new_n677_), .B(regfil_4__2_), .Y(_abc_41356_new_n4604_));
AND2X2 AND2X2_2113 ( .A(_abc_41356_new_n678_), .B(raddrhold_10_), .Y(_abc_41356_new_n4605_));
AND2X2 AND2X2_2114 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n4606_), .Y(_abc_41356_new_n4607_));
AND2X2 AND2X2_2115 ( .A(_abc_41356_new_n4606_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4608_));
AND2X2 AND2X2_2116 ( .A(_abc_41356_new_n4184_), .B(raddrhold_10_), .Y(_abc_41356_new_n4609_));
AND2X2 AND2X2_2117 ( .A(_abc_41356_new_n4613_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4614_));
AND2X2 AND2X2_2118 ( .A(_abc_41356_new_n3424_), .B(rdatahold_2_), .Y(_abc_41356_new_n4615_));
AND2X2 AND2X2_2119 ( .A(_abc_41356_new_n4574_), .B(raddrhold_10_), .Y(_abc_41356_new_n4617_));
AND2X2 AND2X2_212 ( .A(_abc_41356_new_n612_), .B(alu_res_3_), .Y(_abc_41356_new_n880_));
AND2X2 AND2X2_2120 ( .A(_abc_41356_new_n4618_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4619_));
AND2X2 AND2X2_2121 ( .A(_abc_41356_new_n4619_), .B(_abc_41356_new_n4616_), .Y(_abc_41356_new_n4620_));
AND2X2 AND2X2_2122 ( .A(_abc_41356_new_n4622_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4623_));
AND2X2 AND2X2_2123 ( .A(_abc_41356_new_n4122_), .B(raddrhold_11_), .Y(_abc_41356_new_n4625_));
AND2X2 AND2X2_2124 ( .A(_abc_41356_new_n2199_), .B(_abc_41356_new_n4127_), .Y(_abc_41356_new_n4626_));
AND2X2 AND2X2_2125 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1652_), .Y(_abc_41356_new_n4627_));
AND2X2 AND2X2_2126 ( .A(_abc_41356_new_n4629_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4630_));
AND2X2 AND2X2_2127 ( .A(_abc_41356_new_n4630_), .B(_abc_41356_new_n4628_), .Y(_abc_41356_new_n4631_));
AND2X2 AND2X2_2128 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n2205_), .Y(_abc_41356_new_n4632_));
AND2X2 AND2X2_2129 ( .A(_abc_41356_new_n4143_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4635_));
AND2X2 AND2X2_213 ( .A(_abc_41356_new_n881_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n882_));
AND2X2 AND2X2_2130 ( .A(_abc_41356_new_n4635_), .B(_abc_41356_new_n4634_), .Y(_abc_41356_new_n4636_));
AND2X2 AND2X2_2131 ( .A(_abc_41356_new_n677_), .B(regfil_4__3_), .Y(_abc_41356_new_n4637_));
AND2X2 AND2X2_2132 ( .A(_abc_41356_new_n678_), .B(raddrhold_11_), .Y(_abc_41356_new_n4638_));
AND2X2 AND2X2_2133 ( .A(_abc_41356_new_n4640_), .B(_abc_41356_new_n4639_), .Y(_abc_41356_new_n4641_));
AND2X2 AND2X2_2134 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n2199_), .Y(_abc_41356_new_n4643_));
AND2X2 AND2X2_2135 ( .A(_abc_41356_new_n4173_), .B(sp_11_), .Y(_abc_41356_new_n4644_));
AND2X2 AND2X2_2136 ( .A(_abc_41356_new_n4645_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4646_));
AND2X2 AND2X2_2137 ( .A(_abc_41356_new_n4171_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4647_));
AND2X2 AND2X2_2138 ( .A(_abc_41356_new_n4130_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4648_));
AND2X2 AND2X2_2139 ( .A(_abc_41356_new_n4650_), .B(raddrhold_11_), .Y(_abc_41356_new_n4651_));
AND2X2 AND2X2_214 ( .A(_abc_41356_new_n887_), .B(_abc_41356_new_n724_), .Y(_abc_41356_new_n888_));
AND2X2 AND2X2_2140 ( .A(_abc_41356_new_n4653_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4654_));
AND2X2 AND2X2_2141 ( .A(_abc_41356_new_n3424_), .B(rdatahold_3_), .Y(_abc_41356_new_n4655_));
AND2X2 AND2X2_2142 ( .A(_abc_41356_new_n4617_), .B(raddrhold_11_), .Y(_abc_41356_new_n4657_));
AND2X2 AND2X2_2143 ( .A(_abc_41356_new_n4658_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4659_));
AND2X2 AND2X2_2144 ( .A(_abc_41356_new_n4659_), .B(_abc_41356_new_n4656_), .Y(_abc_41356_new_n4660_));
AND2X2 AND2X2_2145 ( .A(_abc_41356_new_n4662_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4663_));
AND2X2 AND2X2_2146 ( .A(_abc_41356_new_n4122_), .B(raddrhold_12_), .Y(_abc_41356_new_n4665_));
AND2X2 AND2X2_2147 ( .A(_abc_41356_new_n2238_), .B(_abc_41356_new_n4127_), .Y(_abc_41356_new_n4666_));
AND2X2 AND2X2_2148 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1723_), .Y(_abc_41356_new_n4667_));
AND2X2 AND2X2_2149 ( .A(_abc_41356_new_n4669_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4670_));
AND2X2 AND2X2_215 ( .A(_abc_41356_new_n886_), .B(_abc_41356_new_n888_), .Y(_abc_41356_new_n889_));
AND2X2 AND2X2_2150 ( .A(_abc_41356_new_n4670_), .B(_abc_41356_new_n4668_), .Y(_abc_41356_new_n4671_));
AND2X2 AND2X2_2151 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n2243_), .Y(_abc_41356_new_n4672_));
AND2X2 AND2X2_2152 ( .A(_abc_41356_new_n4130_), .B(raddrhold_12_), .Y(_abc_41356_new_n4675_));
AND2X2 AND2X2_2153 ( .A(_abc_41356_new_n4676_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4677_));
AND2X2 AND2X2_2154 ( .A(_abc_41356_new_n4173_), .B(sp_12_), .Y(_abc_41356_new_n4678_));
AND2X2 AND2X2_2155 ( .A(_abc_41356_new_n4175_), .B(_abc_41356_new_n2238_), .Y(_abc_41356_new_n4679_));
AND2X2 AND2X2_2156 ( .A(_abc_41356_new_n4680_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4681_));
AND2X2 AND2X2_2157 ( .A(_abc_41356_new_n677_), .B(regfil_4__4_), .Y(_abc_41356_new_n4682_));
AND2X2 AND2X2_2158 ( .A(_abc_41356_new_n678_), .B(raddrhold_12_), .Y(_abc_41356_new_n4683_));
AND2X2 AND2X2_2159 ( .A(_abc_41356_new_n4640_), .B(_abc_41356_new_n4684_), .Y(_abc_41356_new_n4685_));
AND2X2 AND2X2_216 ( .A(_abc_41356_new_n512_), .B(_abc_41356_new_n890_), .Y(_abc_41356_new_n891_));
AND2X2 AND2X2_2160 ( .A(_abc_41356_new_n4686_), .B(raddrhold_12_), .Y(_abc_41356_new_n4687_));
AND2X2 AND2X2_2161 ( .A(_abc_41356_new_n4690_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4691_));
AND2X2 AND2X2_2162 ( .A(_abc_41356_new_n4657_), .B(raddrhold_12_), .Y(_abc_41356_new_n4692_));
AND2X2 AND2X2_2163 ( .A(_abc_41356_new_n4694_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4695_));
AND2X2 AND2X2_2164 ( .A(_abc_41356_new_n4695_), .B(_abc_41356_new_n4693_), .Y(_abc_41356_new_n4696_));
AND2X2 AND2X2_2165 ( .A(_abc_41356_new_n3424_), .B(rdatahold_4_), .Y(_abc_41356_new_n4697_));
AND2X2 AND2X2_2166 ( .A(_abc_41356_new_n4699_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4700_));
AND2X2 AND2X2_2167 ( .A(_abc_41356_new_n4122_), .B(raddrhold_13_), .Y(_abc_41356_new_n4702_));
AND2X2 AND2X2_2168 ( .A(_abc_41356_new_n2277_), .B(_abc_41356_new_n4127_), .Y(_abc_41356_new_n4703_));
AND2X2 AND2X2_2169 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1819_), .Y(_abc_41356_new_n4704_));
AND2X2 AND2X2_217 ( .A(_abc_41356_new_n530_), .B(_abc_41356_new_n893_), .Y(_abc_41356_new_n894_));
AND2X2 AND2X2_2170 ( .A(_abc_41356_new_n4706_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4707_));
AND2X2 AND2X2_2171 ( .A(_abc_41356_new_n4707_), .B(_abc_41356_new_n4705_), .Y(_abc_41356_new_n4708_));
AND2X2 AND2X2_2172 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n2284_), .Y(_abc_41356_new_n4709_));
AND2X2 AND2X2_2173 ( .A(_abc_41356_new_n4711_), .B(_abc_41356_new_n4635_), .Y(_abc_41356_new_n4712_));
AND2X2 AND2X2_2174 ( .A(_abc_41356_new_n2277_), .B(_abc_41356_new_n4175_), .Y(_abc_41356_new_n4713_));
AND2X2 AND2X2_2175 ( .A(_abc_41356_new_n4173_), .B(sp_13_), .Y(_abc_41356_new_n4714_));
AND2X2 AND2X2_2176 ( .A(_abc_41356_new_n4715_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4716_));
AND2X2 AND2X2_2177 ( .A(_abc_41356_new_n4717_), .B(raddrhold_13_), .Y(_abc_41356_new_n4718_));
AND2X2 AND2X2_2178 ( .A(_abc_41356_new_n4184_), .B(raddrhold_13_), .Y(_abc_41356_new_n4719_));
AND2X2 AND2X2_2179 ( .A(_abc_41356_new_n677_), .B(regfil_4__5_), .Y(_abc_41356_new_n4720_));
AND2X2 AND2X2_218 ( .A(_abc_41356_new_n555_), .B(_abc_41356_new_n540_), .Y(_abc_41356_new_n896_));
AND2X2 AND2X2_2180 ( .A(_abc_41356_new_n678_), .B(raddrhold_13_), .Y(_abc_41356_new_n4721_));
AND2X2 AND2X2_2181 ( .A(_abc_41356_new_n4640_), .B(_abc_41356_new_n4722_), .Y(_abc_41356_new_n4723_));
AND2X2 AND2X2_2182 ( .A(_abc_41356_new_n4727_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4728_));
AND2X2 AND2X2_2183 ( .A(_abc_41356_new_n3424_), .B(rdatahold_5_), .Y(_abc_41356_new_n4729_));
AND2X2 AND2X2_2184 ( .A(_abc_41356_new_n4692_), .B(raddrhold_13_), .Y(_abc_41356_new_n4731_));
AND2X2 AND2X2_2185 ( .A(_abc_41356_new_n4732_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4733_));
AND2X2 AND2X2_2186 ( .A(_abc_41356_new_n4733_), .B(_abc_41356_new_n4730_), .Y(_abc_41356_new_n4734_));
AND2X2 AND2X2_2187 ( .A(_abc_41356_new_n4736_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4737_));
AND2X2 AND2X2_2188 ( .A(_abc_41356_new_n4122_), .B(raddrhold_14_), .Y(_abc_41356_new_n4739_));
AND2X2 AND2X2_2189 ( .A(_abc_41356_new_n2315_), .B(_abc_41356_new_n4127_), .Y(_abc_41356_new_n4740_));
AND2X2 AND2X2_219 ( .A(_abc_41356_new_n537_), .B(_abc_41356_new_n539_), .Y(_abc_41356_new_n898_));
AND2X2 AND2X2_2190 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1893_), .Y(_abc_41356_new_n4741_));
AND2X2 AND2X2_2191 ( .A(_abc_41356_new_n4743_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4744_));
AND2X2 AND2X2_2192 ( .A(_abc_41356_new_n4744_), .B(_abc_41356_new_n4742_), .Y(_abc_41356_new_n4745_));
AND2X2 AND2X2_2193 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n2320_), .Y(_abc_41356_new_n4746_));
AND2X2 AND2X2_2194 ( .A(_abc_41356_new_n4750_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4751_));
AND2X2 AND2X2_2195 ( .A(_abc_41356_new_n4749_), .B(_abc_41356_new_n4751_), .Y(_abc_41356_new_n4752_));
AND2X2 AND2X2_2196 ( .A(_abc_41356_new_n2315_), .B(_abc_41356_new_n4175_), .Y(_abc_41356_new_n4753_));
AND2X2 AND2X2_2197 ( .A(_abc_41356_new_n4171_), .B(raddrhold_14_), .Y(_abc_41356_new_n4754_));
AND2X2 AND2X2_2198 ( .A(_abc_41356_new_n4173_), .B(sp_14_), .Y(_abc_41356_new_n4755_));
AND2X2 AND2X2_2199 ( .A(_abc_41356_new_n4757_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4758_));
AND2X2 AND2X2_22 ( .A(_abc_41356_new_n534_), .B(opcode_5_), .Y(_abc_41356_new_n535_));
AND2X2 AND2X2_220 ( .A(_abc_41356_new_n551_), .B(_abc_41356_new_n542_), .Y(_abc_41356_new_n899_));
AND2X2 AND2X2_2200 ( .A(_abc_41356_new_n4184_), .B(raddrhold_14_), .Y(_abc_41356_new_n4759_));
AND2X2 AND2X2_2201 ( .A(_abc_41356_new_n677_), .B(regfil_4__6_), .Y(_abc_41356_new_n4760_));
AND2X2 AND2X2_2202 ( .A(_abc_41356_new_n678_), .B(raddrhold_14_), .Y(_abc_41356_new_n4761_));
AND2X2 AND2X2_2203 ( .A(_abc_41356_new_n4640_), .B(_abc_41356_new_n4762_), .Y(_abc_41356_new_n4763_));
AND2X2 AND2X2_2204 ( .A(_abc_41356_new_n4766_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4767_));
AND2X2 AND2X2_2205 ( .A(_abc_41356_new_n3424_), .B(rdatahold_6_), .Y(_abc_41356_new_n4768_));
AND2X2 AND2X2_2206 ( .A(_abc_41356_new_n4731_), .B(raddrhold_14_), .Y(_abc_41356_new_n4769_));
AND2X2 AND2X2_2207 ( .A(_abc_41356_new_n4771_), .B(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4772_));
AND2X2 AND2X2_2208 ( .A(_abc_41356_new_n4772_), .B(_abc_41356_new_n4770_), .Y(_abc_41356_new_n4773_));
AND2X2 AND2X2_2209 ( .A(_abc_41356_new_n4775_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4776_));
AND2X2 AND2X2_221 ( .A(_abc_41356_new_n541_), .B(_abc_41356_new_n539_), .Y(_abc_41356_new_n901_));
AND2X2 AND2X2_2210 ( .A(_abc_41356_new_n4122_), .B(raddrhold_15_), .Y(_abc_41356_new_n4778_));
AND2X2 AND2X2_2211 ( .A(_abc_41356_new_n2353_), .B(_abc_41356_new_n4127_), .Y(_abc_41356_new_n4779_));
AND2X2 AND2X2_2212 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n1961_), .Y(_abc_41356_new_n4781_));
AND2X2 AND2X2_2213 ( .A(_abc_41356_new_n4782_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n4783_));
AND2X2 AND2X2_2214 ( .A(_abc_41356_new_n4783_), .B(_abc_41356_new_n4780_), .Y(_abc_41356_new_n4784_));
AND2X2 AND2X2_2215 ( .A(_abc_41356_new_n3373_), .B(_abc_41356_new_n2360_), .Y(_abc_41356_new_n4785_));
AND2X2 AND2X2_2216 ( .A(_abc_41356_new_n4789_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4790_));
AND2X2 AND2X2_2217 ( .A(_abc_41356_new_n4788_), .B(_abc_41356_new_n4790_), .Y(_abc_41356_new_n4791_));
AND2X2 AND2X2_2218 ( .A(_abc_41356_new_n2353_), .B(_abc_41356_new_n4175_), .Y(_abc_41356_new_n4792_));
AND2X2 AND2X2_2219 ( .A(_abc_41356_new_n4171_), .B(raddrhold_15_), .Y(_abc_41356_new_n4793_));
AND2X2 AND2X2_222 ( .A(_abc_41356_new_n551_), .B(_abc_41356_new_n901_), .Y(_abc_41356_new_n902_));
AND2X2 AND2X2_2220 ( .A(_abc_41356_new_n4173_), .B(sp_15_), .Y(_abc_41356_new_n4794_));
AND2X2 AND2X2_2221 ( .A(_abc_41356_new_n4796_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4797_));
AND2X2 AND2X2_2222 ( .A(_abc_41356_new_n4184_), .B(raddrhold_15_), .Y(_abc_41356_new_n4798_));
AND2X2 AND2X2_2223 ( .A(_abc_41356_new_n677_), .B(regfil_4__7_), .Y(_abc_41356_new_n4799_));
AND2X2 AND2X2_2224 ( .A(_abc_41356_new_n678_), .B(raddrhold_15_), .Y(_abc_41356_new_n4800_));
AND2X2 AND2X2_2225 ( .A(_abc_41356_new_n4640_), .B(_abc_41356_new_n4801_), .Y(_abc_41356_new_n4802_));
AND2X2 AND2X2_2226 ( .A(_abc_41356_new_n4805_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n4806_));
AND2X2 AND2X2_2227 ( .A(_abc_41356_new_n4117_), .B(raddrhold_15_), .Y(_abc_41356_new_n4807_));
AND2X2 AND2X2_2228 ( .A(_abc_41356_new_n4770_), .B(_abc_41356_new_n4807_), .Y(_abc_41356_new_n4808_));
AND2X2 AND2X2_2229 ( .A(_abc_41356_new_n3424_), .B(rdatahold_7_), .Y(_abc_41356_new_n4809_));
AND2X2 AND2X2_223 ( .A(_abc_41356_new_n900_), .B(_abc_41356_new_n903_), .Y(_abc_41356_new_n904_));
AND2X2 AND2X2_2230 ( .A(_abc_41356_new_n4117_), .B(raddrhold_14_), .Y(_abc_41356_new_n4811_));
AND2X2 AND2X2_2231 ( .A(_abc_41356_new_n4811_), .B(_abc_41356_new_n4810_), .Y(_abc_41356_new_n4812_));
AND2X2 AND2X2_2232 ( .A(_abc_41356_new_n4731_), .B(_abc_41356_new_n4812_), .Y(_abc_41356_new_n4813_));
AND2X2 AND2X2_2233 ( .A(_abc_41356_new_n4816_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4817_));
AND2X2 AND2X2_2234 ( .A(_abc_41356_new_n4819_), .B(_abc_41356_new_n3700_), .Y(_abc_41356_new_n4820_));
AND2X2 AND2X2_2235 ( .A(_abc_41356_new_n4821_), .B(waddrhold_0_), .Y(_abc_41356_new_n4822_));
AND2X2 AND2X2_2236 ( .A(_abc_41356_new_n4824_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4825_));
AND2X2 AND2X2_2237 ( .A(_abc_41356_new_n4825_), .B(_abc_41356_new_n4823_), .Y(_abc_41356_new_n4826_));
AND2X2 AND2X2_2238 ( .A(_abc_41356_new_n678_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4828_));
AND2X2 AND2X2_2239 ( .A(_abc_41356_new_n4827_), .B(_abc_41356_new_n4828_), .Y(_abc_41356_new_n4829_));
AND2X2 AND2X2_224 ( .A(_abc_41356_new_n905_), .B(_abc_41356_new_n897_), .Y(_abc_41356_new_n906_));
AND2X2 AND2X2_2240 ( .A(_abc_41356_new_n4830_), .B(waddrhold_0_), .Y(_abc_41356_new_n4831_));
AND2X2 AND2X2_2241 ( .A(_abc_41356_new_n4138_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4832_));
AND2X2 AND2X2_2242 ( .A(_abc_41356_new_n4832_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n4833_));
AND2X2 AND2X2_2243 ( .A(_abc_41356_new_n4132_), .B(_abc_41356_new_n4834_), .Y(_abc_41356_new_n4835_));
AND2X2 AND2X2_2244 ( .A(_abc_41356_new_n678_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n4836_));
AND2X2 AND2X2_2245 ( .A(_abc_41356_new_n677_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4837_));
AND2X2 AND2X2_2246 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n4835_), .Y(_abc_41356_new_n4839_));
AND2X2 AND2X2_2247 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n4844_), .Y(_abc_41356_new_n4845_));
AND2X2 AND2X2_2248 ( .A(_abc_41356_new_n4843_), .B(_abc_41356_new_n4845_), .Y(_abc_41356_new_n4846_));
AND2X2 AND2X2_2249 ( .A(_abc_41356_new_n3430_), .B(regfil_5__0_), .Y(_abc_41356_new_n4847_));
AND2X2 AND2X2_225 ( .A(_abc_41356_new_n907_), .B(_abc_41356_new_n895_), .Y(_abc_41356_new_n908_));
AND2X2 AND2X2_2250 ( .A(_abc_41356_new_n3698_), .B(_abc_41356_new_n4848_), .Y(_abc_41356_new_n4849_));
AND2X2 AND2X2_2251 ( .A(_abc_41356_new_n3432_), .B(rdatahold2_0_), .Y(_abc_41356_new_n4850_));
AND2X2 AND2X2_2252 ( .A(_abc_41356_new_n4853_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4854_));
AND2X2 AND2X2_2253 ( .A(_abc_41356_new_n4821_), .B(waddrhold_1_), .Y(_abc_41356_new_n4856_));
AND2X2 AND2X2_2254 ( .A(_abc_41356_new_n4860_), .B(_abc_41356_new_n4857_), .Y(_abc_41356_new_n4861_));
AND2X2 AND2X2_2255 ( .A(_abc_41356_new_n1218_), .B(sp_1_), .Y(_abc_41356_new_n4862_));
AND2X2 AND2X2_2256 ( .A(_abc_41356_new_n4865_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4866_));
AND2X2 AND2X2_2257 ( .A(_abc_41356_new_n4864_), .B(_abc_41356_new_n4866_), .Y(_abc_41356_new_n4867_));
AND2X2 AND2X2_2258 ( .A(_abc_41356_new_n4830_), .B(waddrhold_1_), .Y(_abc_41356_new_n4868_));
AND2X2 AND2X2_2259 ( .A(_abc_41356_new_n4208_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4869_));
AND2X2 AND2X2_226 ( .A(_abc_41356_new_n909_), .B(_abc_41356_new_n892_), .Y(_abc_41356_new_n910_));
AND2X2 AND2X2_2260 ( .A(_abc_41356_new_n4869_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n4870_));
AND2X2 AND2X2_2261 ( .A(_abc_41356_new_n4203_), .B(_abc_41356_new_n4871_), .Y(_abc_41356_new_n4872_));
AND2X2 AND2X2_2262 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n4872_), .Y(_abc_41356_new_n4873_));
AND2X2 AND2X2_2263 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n4878_), .Y(_abc_41356_new_n4879_));
AND2X2 AND2X2_2264 ( .A(_abc_41356_new_n4877_), .B(_abc_41356_new_n4879_), .Y(_abc_41356_new_n4880_));
AND2X2 AND2X2_2265 ( .A(_abc_41356_new_n3430_), .B(regfil_5__1_), .Y(_abc_41356_new_n4881_));
AND2X2 AND2X2_2266 ( .A(_abc_41356_new_n3432_), .B(rdatahold2_1_), .Y(_abc_41356_new_n4882_));
AND2X2 AND2X2_2267 ( .A(waddrhold_0_), .B(waddrhold_1_), .Y(_abc_41356_new_n4883_));
AND2X2 AND2X2_2268 ( .A(_abc_41356_new_n4884_), .B(_abc_41356_new_n4885_), .Y(_abc_41356_new_n4886_));
AND2X2 AND2X2_2269 ( .A(_abc_41356_new_n3698_), .B(_abc_41356_new_n4886_), .Y(_abc_41356_new_n4887_));
AND2X2 AND2X2_227 ( .A(_abc_41356_new_n712_), .B(regfil_7__3_), .Y(_abc_41356_new_n911_));
AND2X2 AND2X2_2270 ( .A(_abc_41356_new_n4890_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4891_));
AND2X2 AND2X2_2271 ( .A(_abc_41356_new_n4821_), .B(waddrhold_2_), .Y(_abc_41356_new_n4893_));
AND2X2 AND2X2_2272 ( .A(_abc_41356_new_n1298_), .B(_abc_41356_new_n4857_), .Y(_abc_41356_new_n4894_));
AND2X2 AND2X2_2273 ( .A(sp_2_), .B(sp_1_), .Y(_abc_41356_new_n4895_));
AND2X2 AND2X2_2274 ( .A(_abc_41356_new_n4860_), .B(_abc_41356_new_n4896_), .Y(_abc_41356_new_n4897_));
AND2X2 AND2X2_2275 ( .A(_abc_41356_new_n1218_), .B(sp_2_), .Y(_abc_41356_new_n4898_));
AND2X2 AND2X2_2276 ( .A(_abc_41356_new_n4901_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4902_));
AND2X2 AND2X2_2277 ( .A(_abc_41356_new_n4900_), .B(_abc_41356_new_n4902_), .Y(_abc_41356_new_n4903_));
AND2X2 AND2X2_2278 ( .A(_abc_41356_new_n4830_), .B(waddrhold_2_), .Y(_abc_41356_new_n4904_));
AND2X2 AND2X2_2279 ( .A(_abc_41356_new_n4252_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4905_));
AND2X2 AND2X2_228 ( .A(_abc_41356_new_n714_), .B(alu_res_3_), .Y(_abc_41356_new_n912_));
AND2X2 AND2X2_2280 ( .A(_abc_41356_new_n4905_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n4906_));
AND2X2 AND2X2_2281 ( .A(_abc_41356_new_n4246_), .B(_abc_41356_new_n4907_), .Y(_abc_41356_new_n4908_));
AND2X2 AND2X2_2282 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n4908_), .Y(_abc_41356_new_n4909_));
AND2X2 AND2X2_2283 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n4914_), .Y(_abc_41356_new_n4915_));
AND2X2 AND2X2_2284 ( .A(_abc_41356_new_n4913_), .B(_abc_41356_new_n4915_), .Y(_abc_41356_new_n4916_));
AND2X2 AND2X2_2285 ( .A(_abc_41356_new_n3430_), .B(regfil_5__2_), .Y(_abc_41356_new_n4917_));
AND2X2 AND2X2_2286 ( .A(_abc_41356_new_n3432_), .B(rdatahold2_2_), .Y(_abc_41356_new_n4918_));
AND2X2 AND2X2_2287 ( .A(_abc_41356_new_n4883_), .B(waddrhold_2_), .Y(_abc_41356_new_n4920_));
AND2X2 AND2X2_2288 ( .A(_abc_41356_new_n4921_), .B(_abc_41356_new_n4919_), .Y(_abc_41356_new_n4922_));
AND2X2 AND2X2_2289 ( .A(_abc_41356_new_n4922_), .B(_abc_41356_new_n3698_), .Y(_abc_41356_new_n4923_));
AND2X2 AND2X2_229 ( .A(_abc_41356_new_n718_), .B(\data[3] ), .Y(_abc_41356_new_n913_));
AND2X2 AND2X2_2290 ( .A(_abc_41356_new_n4926_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4927_));
AND2X2 AND2X2_2291 ( .A(_abc_41356_new_n4821_), .B(waddrhold_3_), .Y(_abc_41356_new_n4929_));
AND2X2 AND2X2_2292 ( .A(_abc_41356_new_n4931_), .B(_abc_41356_new_n4932_), .Y(_abc_41356_new_n4933_));
AND2X2 AND2X2_2293 ( .A(_abc_41356_new_n4860_), .B(_abc_41356_new_n4933_), .Y(_abc_41356_new_n4934_));
AND2X2 AND2X2_2294 ( .A(_abc_41356_new_n1218_), .B(sp_3_), .Y(_abc_41356_new_n4935_));
AND2X2 AND2X2_2295 ( .A(_abc_41356_new_n4938_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4939_));
AND2X2 AND2X2_2296 ( .A(_abc_41356_new_n4937_), .B(_abc_41356_new_n4939_), .Y(_abc_41356_new_n4940_));
AND2X2 AND2X2_2297 ( .A(_abc_41356_new_n4830_), .B(waddrhold_3_), .Y(_abc_41356_new_n4941_));
AND2X2 AND2X2_2298 ( .A(_abc_41356_new_n4296_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4942_));
AND2X2 AND2X2_2299 ( .A(_abc_41356_new_n4942_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n4943_));
AND2X2 AND2X2_23 ( .A(_abc_41356_new_n528_), .B(_abc_41356_new_n535_), .Y(_abc_41356_new_n536_));
AND2X2 AND2X2_230 ( .A(_abc_41356_new_n851_), .B(regfil_0__4_), .Y(_abc_41356_new_n920_));
AND2X2 AND2X2_2300 ( .A(_abc_41356_new_n4290_), .B(_abc_41356_new_n4944_), .Y(_abc_41356_new_n4945_));
AND2X2 AND2X2_2301 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n4945_), .Y(_abc_41356_new_n4946_));
AND2X2 AND2X2_2302 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n4951_), .Y(_abc_41356_new_n4952_));
AND2X2 AND2X2_2303 ( .A(_abc_41356_new_n4950_), .B(_abc_41356_new_n4952_), .Y(_abc_41356_new_n4953_));
AND2X2 AND2X2_2304 ( .A(_abc_41356_new_n3430_), .B(regfil_5__3_), .Y(_abc_41356_new_n4954_));
AND2X2 AND2X2_2305 ( .A(_abc_41356_new_n3432_), .B(rdatahold2_3_), .Y(_abc_41356_new_n4955_));
AND2X2 AND2X2_2306 ( .A(_abc_41356_new_n4920_), .B(waddrhold_3_), .Y(_abc_41356_new_n4956_));
AND2X2 AND2X2_2307 ( .A(_abc_41356_new_n3698_), .B(_abc_41356_new_n4958_), .Y(_abc_41356_new_n4959_));
AND2X2 AND2X2_2308 ( .A(_abc_41356_new_n4959_), .B(_abc_41356_new_n4957_), .Y(_abc_41356_new_n4960_));
AND2X2 AND2X2_2309 ( .A(_abc_41356_new_n4963_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n4964_));
AND2X2 AND2X2_231 ( .A(_abc_41356_new_n921_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n922_));
AND2X2 AND2X2_2310 ( .A(_abc_41356_new_n4821_), .B(waddrhold_4_), .Y(_abc_41356_new_n4966_));
AND2X2 AND2X2_2311 ( .A(_abc_41356_new_n4894_), .B(_abc_41356_new_n1303_), .Y(_abc_41356_new_n4967_));
AND2X2 AND2X2_2312 ( .A(_abc_41356_new_n4967_), .B(_abc_41356_new_n1325_), .Y(_abc_41356_new_n4968_));
AND2X2 AND2X2_2313 ( .A(_abc_41356_new_n4969_), .B(sp_4_), .Y(_abc_41356_new_n4970_));
AND2X2 AND2X2_2314 ( .A(_abc_41356_new_n4860_), .B(_abc_41356_new_n4971_), .Y(_abc_41356_new_n4972_));
AND2X2 AND2X2_2315 ( .A(_abc_41356_new_n1218_), .B(sp_4_), .Y(_abc_41356_new_n4973_));
AND2X2 AND2X2_2316 ( .A(_abc_41356_new_n4976_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n4977_));
AND2X2 AND2X2_2317 ( .A(_abc_41356_new_n4975_), .B(_abc_41356_new_n4977_), .Y(_abc_41356_new_n4978_));
AND2X2 AND2X2_2318 ( .A(_abc_41356_new_n4830_), .B(waddrhold_4_), .Y(_abc_41356_new_n4979_));
AND2X2 AND2X2_2319 ( .A(_abc_41356_new_n4339_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n4980_));
AND2X2 AND2X2_232 ( .A(_abc_41356_new_n857_), .B(regfil_0__4_), .Y(_abc_41356_new_n924_));
AND2X2 AND2X2_2320 ( .A(_abc_41356_new_n4980_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n4981_));
AND2X2 AND2X2_2321 ( .A(_abc_41356_new_n4333_), .B(_abc_41356_new_n4982_), .Y(_abc_41356_new_n4983_));
AND2X2 AND2X2_2322 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n4983_), .Y(_abc_41356_new_n4984_));
AND2X2 AND2X2_2323 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n4989_), .Y(_abc_41356_new_n4990_));
AND2X2 AND2X2_2324 ( .A(_abc_41356_new_n4988_), .B(_abc_41356_new_n4990_), .Y(_abc_41356_new_n4991_));
AND2X2 AND2X2_2325 ( .A(_abc_41356_new_n3432_), .B(rdatahold2_4_), .Y(_abc_41356_new_n4992_));
AND2X2 AND2X2_2326 ( .A(_abc_41356_new_n3430_), .B(regfil_5__4_), .Y(_abc_41356_new_n4993_));
AND2X2 AND2X2_2327 ( .A(_abc_41356_new_n4956_), .B(waddrhold_4_), .Y(_abc_41356_new_n4995_));
AND2X2 AND2X2_2328 ( .A(_abc_41356_new_n4997_), .B(_abc_41356_new_n3698_), .Y(_abc_41356_new_n4998_));
AND2X2 AND2X2_2329 ( .A(_abc_41356_new_n4998_), .B(_abc_41356_new_n4996_), .Y(_abc_41356_new_n4999_));
AND2X2 AND2X2_233 ( .A(_abc_41356_new_n925_), .B(_abc_41356_new_n581_), .Y(_abc_41356_new_n926_));
AND2X2 AND2X2_2330 ( .A(_abc_41356_new_n5001_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5002_));
AND2X2 AND2X2_2331 ( .A(_abc_41356_new_n4821_), .B(waddrhold_5_), .Y(_abc_41356_new_n5004_));
AND2X2 AND2X2_2332 ( .A(_abc_41356_new_n5005_), .B(sp_5_), .Y(_abc_41356_new_n5006_));
AND2X2 AND2X2_2333 ( .A(_abc_41356_new_n4968_), .B(_abc_41356_new_n1331_), .Y(_abc_41356_new_n5007_));
AND2X2 AND2X2_2334 ( .A(_abc_41356_new_n4860_), .B(_abc_41356_new_n5008_), .Y(_abc_41356_new_n5009_));
AND2X2 AND2X2_2335 ( .A(_abc_41356_new_n1218_), .B(sp_5_), .Y(_abc_41356_new_n5010_));
AND2X2 AND2X2_2336 ( .A(_abc_41356_new_n5013_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5014_));
AND2X2 AND2X2_2337 ( .A(_abc_41356_new_n5012_), .B(_abc_41356_new_n5014_), .Y(_abc_41356_new_n5015_));
AND2X2 AND2X2_2338 ( .A(_abc_41356_new_n4830_), .B(waddrhold_5_), .Y(_abc_41356_new_n5016_));
AND2X2 AND2X2_2339 ( .A(_abc_41356_new_n4382_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5017_));
AND2X2 AND2X2_234 ( .A(_abc_41356_new_n926_), .B(_abc_41356_new_n923_), .Y(_abc_41356_new_n927_));
AND2X2 AND2X2_2340 ( .A(_abc_41356_new_n5017_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5018_));
AND2X2 AND2X2_2341 ( .A(_abc_41356_new_n4376_), .B(_abc_41356_new_n5019_), .Y(_abc_41356_new_n5020_));
AND2X2 AND2X2_2342 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5020_), .Y(_abc_41356_new_n5021_));
AND2X2 AND2X2_2343 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5026_), .Y(_abc_41356_new_n5027_));
AND2X2 AND2X2_2344 ( .A(_abc_41356_new_n5025_), .B(_abc_41356_new_n5027_), .Y(_abc_41356_new_n5028_));
AND2X2 AND2X2_2345 ( .A(_abc_41356_new_n3432_), .B(rdatahold2_5_), .Y(_abc_41356_new_n5029_));
AND2X2 AND2X2_2346 ( .A(_abc_41356_new_n3430_), .B(regfil_5__5_), .Y(_abc_41356_new_n5030_));
AND2X2 AND2X2_2347 ( .A(_abc_41356_new_n4995_), .B(waddrhold_5_), .Y(_abc_41356_new_n5032_));
AND2X2 AND2X2_2348 ( .A(_abc_41356_new_n5034_), .B(_abc_41356_new_n3698_), .Y(_abc_41356_new_n5035_));
AND2X2 AND2X2_2349 ( .A(_abc_41356_new_n5035_), .B(_abc_41356_new_n5033_), .Y(_abc_41356_new_n5036_));
AND2X2 AND2X2_235 ( .A(_abc_41356_new_n642_), .B(rdatahold_4_), .Y(_abc_41356_new_n928_));
AND2X2 AND2X2_2350 ( .A(_abc_41356_new_n5038_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5039_));
AND2X2 AND2X2_2351 ( .A(_abc_41356_new_n4821_), .B(waddrhold_6_), .Y(_abc_41356_new_n5041_));
AND2X2 AND2X2_2352 ( .A(_abc_41356_new_n5007_), .B(_abc_41356_new_n1319_), .Y(_abc_41356_new_n5042_));
AND2X2 AND2X2_2353 ( .A(_abc_41356_new_n5043_), .B(sp_6_), .Y(_abc_41356_new_n5044_));
AND2X2 AND2X2_2354 ( .A(_abc_41356_new_n4860_), .B(_abc_41356_new_n5045_), .Y(_abc_41356_new_n5046_));
AND2X2 AND2X2_2355 ( .A(_abc_41356_new_n1218_), .B(sp_6_), .Y(_abc_41356_new_n5047_));
AND2X2 AND2X2_2356 ( .A(_abc_41356_new_n5050_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5051_));
AND2X2 AND2X2_2357 ( .A(_abc_41356_new_n5049_), .B(_abc_41356_new_n5051_), .Y(_abc_41356_new_n5052_));
AND2X2 AND2X2_2358 ( .A(_abc_41356_new_n4830_), .B(waddrhold_6_), .Y(_abc_41356_new_n5053_));
AND2X2 AND2X2_2359 ( .A(_abc_41356_new_n4425_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5054_));
AND2X2 AND2X2_236 ( .A(_abc_41356_new_n616_), .B(regfil_5__4_), .Y(_abc_41356_new_n929_));
AND2X2 AND2X2_2360 ( .A(_abc_41356_new_n5054_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5055_));
AND2X2 AND2X2_2361 ( .A(_abc_41356_new_n4419_), .B(_abc_41356_new_n5056_), .Y(_abc_41356_new_n5057_));
AND2X2 AND2X2_2362 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5057_), .Y(_abc_41356_new_n5058_));
AND2X2 AND2X2_2363 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5063_), .Y(_abc_41356_new_n5064_));
AND2X2 AND2X2_2364 ( .A(_abc_41356_new_n5062_), .B(_abc_41356_new_n5064_), .Y(_abc_41356_new_n5065_));
AND2X2 AND2X2_2365 ( .A(_abc_41356_new_n3432_), .B(rdatahold2_6_), .Y(_abc_41356_new_n5066_));
AND2X2 AND2X2_2366 ( .A(_abc_41356_new_n3430_), .B(regfil_5__6_), .Y(_abc_41356_new_n5067_));
AND2X2 AND2X2_2367 ( .A(_abc_41356_new_n5032_), .B(waddrhold_6_), .Y(_abc_41356_new_n5069_));
AND2X2 AND2X2_2368 ( .A(_abc_41356_new_n5071_), .B(_abc_41356_new_n3698_), .Y(_abc_41356_new_n5072_));
AND2X2 AND2X2_2369 ( .A(_abc_41356_new_n5072_), .B(_abc_41356_new_n5070_), .Y(_abc_41356_new_n5073_));
AND2X2 AND2X2_237 ( .A(_abc_41356_new_n619_), .B(regfil_4__4_), .Y(_abc_41356_new_n930_));
AND2X2 AND2X2_2370 ( .A(_abc_41356_new_n5075_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5076_));
AND2X2 AND2X2_2371 ( .A(_abc_41356_new_n4821_), .B(waddrhold_7_), .Y(_abc_41356_new_n5078_));
AND2X2 AND2X2_2372 ( .A(_abc_41356_new_n5079_), .B(sp_7_), .Y(_abc_41356_new_n5080_));
AND2X2 AND2X2_2373 ( .A(_abc_41356_new_n5042_), .B(_abc_41356_new_n1314_), .Y(_abc_41356_new_n5081_));
AND2X2 AND2X2_2374 ( .A(_abc_41356_new_n4860_), .B(_abc_41356_new_n5082_), .Y(_abc_41356_new_n5083_));
AND2X2 AND2X2_2375 ( .A(_abc_41356_new_n1218_), .B(sp_7_), .Y(_abc_41356_new_n5084_));
AND2X2 AND2X2_2376 ( .A(_abc_41356_new_n5087_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5088_));
AND2X2 AND2X2_2377 ( .A(_abc_41356_new_n5086_), .B(_abc_41356_new_n5088_), .Y(_abc_41356_new_n5089_));
AND2X2 AND2X2_2378 ( .A(_abc_41356_new_n4830_), .B(waddrhold_7_), .Y(_abc_41356_new_n5090_));
AND2X2 AND2X2_2379 ( .A(_abc_41356_new_n4467_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5091_));
AND2X2 AND2X2_238 ( .A(_abc_41356_new_n526_), .B(regfil_7__4_), .Y(_abc_41356_new_n932_));
AND2X2 AND2X2_2380 ( .A(_abc_41356_new_n5091_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5092_));
AND2X2 AND2X2_2381 ( .A(_abc_41356_new_n4461_), .B(_abc_41356_new_n5093_), .Y(_abc_41356_new_n5094_));
AND2X2 AND2X2_2382 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5094_), .Y(_abc_41356_new_n5095_));
AND2X2 AND2X2_2383 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5100_), .Y(_abc_41356_new_n5101_));
AND2X2 AND2X2_2384 ( .A(_abc_41356_new_n5099_), .B(_abc_41356_new_n5101_), .Y(_abc_41356_new_n5102_));
AND2X2 AND2X2_2385 ( .A(_abc_41356_new_n3432_), .B(rdatahold2_7_), .Y(_abc_41356_new_n5103_));
AND2X2 AND2X2_2386 ( .A(_abc_41356_new_n3430_), .B(regfil_5__7_), .Y(_abc_41356_new_n5104_));
AND2X2 AND2X2_2387 ( .A(_abc_41356_new_n5069_), .B(waddrhold_7_), .Y(_abc_41356_new_n5106_));
AND2X2 AND2X2_2388 ( .A(_abc_41356_new_n5108_), .B(_abc_41356_new_n3698_), .Y(_abc_41356_new_n5109_));
AND2X2 AND2X2_2389 ( .A(_abc_41356_new_n5109_), .B(_abc_41356_new_n5107_), .Y(_abc_41356_new_n5110_));
AND2X2 AND2X2_239 ( .A(_abc_41356_new_n623_), .B(regfil_6__4_), .Y(_abc_41356_new_n933_));
AND2X2 AND2X2_2390 ( .A(_abc_41356_new_n5112_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5113_));
AND2X2 AND2X2_2391 ( .A(_abc_41356_new_n4821_), .B(waddrhold_8_), .Y(_abc_41356_new_n5115_));
AND2X2 AND2X2_2392 ( .A(_abc_41356_new_n5081_), .B(_abc_41356_new_n1345_), .Y(_abc_41356_new_n5116_));
AND2X2 AND2X2_2393 ( .A(_abc_41356_new_n5117_), .B(sp_8_), .Y(_abc_41356_new_n5118_));
AND2X2 AND2X2_2394 ( .A(_abc_41356_new_n4860_), .B(_abc_41356_new_n5119_), .Y(_abc_41356_new_n5120_));
AND2X2 AND2X2_2395 ( .A(_abc_41356_new_n1218_), .B(sp_8_), .Y(_abc_41356_new_n5121_));
AND2X2 AND2X2_2396 ( .A(_abc_41356_new_n5124_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5125_));
AND2X2 AND2X2_2397 ( .A(_abc_41356_new_n5123_), .B(_abc_41356_new_n5125_), .Y(_abc_41356_new_n5126_));
AND2X2 AND2X2_2398 ( .A(_abc_41356_new_n4830_), .B(waddrhold_8_), .Y(_abc_41356_new_n5127_));
AND2X2 AND2X2_2399 ( .A(_abc_41356_new_n2086_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5128_));
AND2X2 AND2X2_24 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n536_), .Y(_abc_41356_new_n537_));
AND2X2 AND2X2_240 ( .A(_abc_41356_new_n616_), .B(regfil_1__4_), .Y(_abc_41356_new_n937_));
AND2X2 AND2X2_2400 ( .A(_abc_41356_new_n5128_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5129_));
AND2X2 AND2X2_2401 ( .A(_abc_41356_new_n4504_), .B(_abc_41356_new_n5130_), .Y(_abc_41356_new_n5131_));
AND2X2 AND2X2_2402 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5131_), .Y(_abc_41356_new_n5132_));
AND2X2 AND2X2_2403 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5137_), .Y(_abc_41356_new_n5138_));
AND2X2 AND2X2_2404 ( .A(_abc_41356_new_n5136_), .B(_abc_41356_new_n5138_), .Y(_abc_41356_new_n5139_));
AND2X2 AND2X2_2405 ( .A(_abc_41356_new_n3432_), .B(rdatahold_0_), .Y(_abc_41356_new_n5140_));
AND2X2 AND2X2_2406 ( .A(_abc_41356_new_n3430_), .B(regfil_4__0_), .Y(_abc_41356_new_n5141_));
AND2X2 AND2X2_2407 ( .A(_abc_41356_new_n5106_), .B(waddrhold_8_), .Y(_abc_41356_new_n5143_));
AND2X2 AND2X2_2408 ( .A(_abc_41356_new_n5145_), .B(_abc_41356_new_n3698_), .Y(_abc_41356_new_n5146_));
AND2X2 AND2X2_2409 ( .A(_abc_41356_new_n5146_), .B(_abc_41356_new_n5144_), .Y(_abc_41356_new_n5147_));
AND2X2 AND2X2_241 ( .A(_abc_41356_new_n623_), .B(regfil_2__4_), .Y(_abc_41356_new_n939_));
AND2X2 AND2X2_2410 ( .A(_abc_41356_new_n5149_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5150_));
AND2X2 AND2X2_2411 ( .A(_abc_41356_new_n4821_), .B(waddrhold_9_), .Y(_abc_41356_new_n5152_));
AND2X2 AND2X2_2412 ( .A(_abc_41356_new_n5153_), .B(sp_9_), .Y(_abc_41356_new_n5154_));
AND2X2 AND2X2_2413 ( .A(_abc_41356_new_n5116_), .B(_abc_41356_new_n1515_), .Y(_abc_41356_new_n5155_));
AND2X2 AND2X2_2414 ( .A(_abc_41356_new_n5156_), .B(_abc_41356_new_n4860_), .Y(_abc_41356_new_n5157_));
AND2X2 AND2X2_2415 ( .A(_abc_41356_new_n1218_), .B(sp_9_), .Y(_abc_41356_new_n5158_));
AND2X2 AND2X2_2416 ( .A(_abc_41356_new_n5161_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5162_));
AND2X2 AND2X2_2417 ( .A(_abc_41356_new_n5160_), .B(_abc_41356_new_n5162_), .Y(_abc_41356_new_n5163_));
AND2X2 AND2X2_2418 ( .A(_abc_41356_new_n4830_), .B(waddrhold_9_), .Y(_abc_41356_new_n5164_));
AND2X2 AND2X2_2419 ( .A(_abc_41356_new_n2127_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5165_));
AND2X2 AND2X2_242 ( .A(_abc_41356_new_n619_), .B(regfil_0__4_), .Y(_abc_41356_new_n940_));
AND2X2 AND2X2_2420 ( .A(_abc_41356_new_n5165_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5166_));
AND2X2 AND2X2_2421 ( .A(_abc_41356_new_n4545_), .B(_abc_41356_new_n5167_), .Y(_abc_41356_new_n5168_));
AND2X2 AND2X2_2422 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5168_), .Y(_abc_41356_new_n5169_));
AND2X2 AND2X2_2423 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5174_), .Y(_abc_41356_new_n5175_));
AND2X2 AND2X2_2424 ( .A(_abc_41356_new_n5173_), .B(_abc_41356_new_n5175_), .Y(_abc_41356_new_n5176_));
AND2X2 AND2X2_2425 ( .A(_abc_41356_new_n3432_), .B(rdatahold_1_), .Y(_abc_41356_new_n5177_));
AND2X2 AND2X2_2426 ( .A(_abc_41356_new_n3430_), .B(regfil_4__1_), .Y(_abc_41356_new_n5178_));
AND2X2 AND2X2_2427 ( .A(_abc_41356_new_n5143_), .B(waddrhold_9_), .Y(_abc_41356_new_n5180_));
AND2X2 AND2X2_2428 ( .A(_abc_41356_new_n5182_), .B(_abc_41356_new_n3698_), .Y(_abc_41356_new_n5183_));
AND2X2 AND2X2_2429 ( .A(_abc_41356_new_n5183_), .B(_abc_41356_new_n5181_), .Y(_abc_41356_new_n5184_));
AND2X2 AND2X2_243 ( .A(_abc_41356_new_n526_), .B(regfil_3__4_), .Y(_abc_41356_new_n941_));
AND2X2 AND2X2_2430 ( .A(_abc_41356_new_n5186_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5187_));
AND2X2 AND2X2_2431 ( .A(_abc_41356_new_n4821_), .B(waddrhold_10_), .Y(_abc_41356_new_n5189_));
AND2X2 AND2X2_2432 ( .A(_abc_41356_new_n5155_), .B(_abc_41356_new_n1596_), .Y(_abc_41356_new_n5190_));
AND2X2 AND2X2_2433 ( .A(_abc_41356_new_n5191_), .B(sp_10_), .Y(_abc_41356_new_n5192_));
AND2X2 AND2X2_2434 ( .A(_abc_41356_new_n5193_), .B(_abc_41356_new_n4860_), .Y(_abc_41356_new_n5194_));
AND2X2 AND2X2_2435 ( .A(_abc_41356_new_n1218_), .B(sp_10_), .Y(_abc_41356_new_n5195_));
AND2X2 AND2X2_2436 ( .A(_abc_41356_new_n5198_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5199_));
AND2X2 AND2X2_2437 ( .A(_abc_41356_new_n5197_), .B(_abc_41356_new_n5199_), .Y(_abc_41356_new_n5200_));
AND2X2 AND2X2_2438 ( .A(_abc_41356_new_n4830_), .B(waddrhold_10_), .Y(_abc_41356_new_n5201_));
AND2X2 AND2X2_2439 ( .A(_abc_41356_new_n2165_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5202_));
AND2X2 AND2X2_244 ( .A(_abc_41356_new_n936_), .B(_abc_41356_new_n944_), .Y(_abc_41356_new_n945_));
AND2X2 AND2X2_2440 ( .A(_abc_41356_new_n5202_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5203_));
AND2X2 AND2X2_2441 ( .A(_abc_41356_new_n4593_), .B(_abc_41356_new_n5204_), .Y(_abc_41356_new_n5205_));
AND2X2 AND2X2_2442 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5205_), .Y(_abc_41356_new_n5206_));
AND2X2 AND2X2_2443 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5211_), .Y(_abc_41356_new_n5212_));
AND2X2 AND2X2_2444 ( .A(_abc_41356_new_n5210_), .B(_abc_41356_new_n5212_), .Y(_abc_41356_new_n5213_));
AND2X2 AND2X2_2445 ( .A(_abc_41356_new_n3432_), .B(rdatahold_2_), .Y(_abc_41356_new_n5214_));
AND2X2 AND2X2_2446 ( .A(_abc_41356_new_n3430_), .B(regfil_4__2_), .Y(_abc_41356_new_n5215_));
AND2X2 AND2X2_2447 ( .A(_abc_41356_new_n5180_), .B(waddrhold_10_), .Y(_abc_41356_new_n5217_));
AND2X2 AND2X2_2448 ( .A(_abc_41356_new_n5219_), .B(_abc_41356_new_n3698_), .Y(_abc_41356_new_n5220_));
AND2X2 AND2X2_2449 ( .A(_abc_41356_new_n5220_), .B(_abc_41356_new_n5218_), .Y(_abc_41356_new_n5221_));
AND2X2 AND2X2_245 ( .A(_abc_41356_new_n945_), .B(_abc_41356_new_n614_), .Y(_abc_41356_new_n946_));
AND2X2 AND2X2_2450 ( .A(_abc_41356_new_n5223_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5224_));
AND2X2 AND2X2_2451 ( .A(_abc_41356_new_n4821_), .B(waddrhold_11_), .Y(_abc_41356_new_n5226_));
AND2X2 AND2X2_2452 ( .A(_abc_41356_new_n5227_), .B(sp_11_), .Y(_abc_41356_new_n5228_));
AND2X2 AND2X2_2453 ( .A(_abc_41356_new_n5190_), .B(_abc_41356_new_n1653_), .Y(_abc_41356_new_n5229_));
AND2X2 AND2X2_2454 ( .A(_abc_41356_new_n5230_), .B(_abc_41356_new_n4860_), .Y(_abc_41356_new_n5231_));
AND2X2 AND2X2_2455 ( .A(_abc_41356_new_n1218_), .B(sp_11_), .Y(_abc_41356_new_n5232_));
AND2X2 AND2X2_2456 ( .A(_abc_41356_new_n5235_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5236_));
AND2X2 AND2X2_2457 ( .A(_abc_41356_new_n5234_), .B(_abc_41356_new_n5236_), .Y(_abc_41356_new_n5237_));
AND2X2 AND2X2_2458 ( .A(_abc_41356_new_n4830_), .B(waddrhold_11_), .Y(_abc_41356_new_n5238_));
AND2X2 AND2X2_2459 ( .A(_abc_41356_new_n2205_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5239_));
AND2X2 AND2X2_246 ( .A(_abc_41356_new_n612_), .B(alu_res_4_), .Y(_abc_41356_new_n947_));
AND2X2 AND2X2_2460 ( .A(_abc_41356_new_n5239_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5240_));
AND2X2 AND2X2_2461 ( .A(_abc_41356_new_n4628_), .B(_abc_41356_new_n5241_), .Y(_abc_41356_new_n5242_));
AND2X2 AND2X2_2462 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5242_), .Y(_abc_41356_new_n5243_));
AND2X2 AND2X2_2463 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5248_), .Y(_abc_41356_new_n5249_));
AND2X2 AND2X2_2464 ( .A(_abc_41356_new_n5247_), .B(_abc_41356_new_n5249_), .Y(_abc_41356_new_n5250_));
AND2X2 AND2X2_2465 ( .A(_abc_41356_new_n3432_), .B(rdatahold_3_), .Y(_abc_41356_new_n5251_));
AND2X2 AND2X2_2466 ( .A(_abc_41356_new_n3430_), .B(regfil_4__3_), .Y(_abc_41356_new_n5252_));
AND2X2 AND2X2_2467 ( .A(_abc_41356_new_n5217_), .B(waddrhold_11_), .Y(_abc_41356_new_n5254_));
AND2X2 AND2X2_2468 ( .A(_abc_41356_new_n5256_), .B(_abc_41356_new_n3698_), .Y(_abc_41356_new_n5257_));
AND2X2 AND2X2_2469 ( .A(_abc_41356_new_n5257_), .B(_abc_41356_new_n5255_), .Y(_abc_41356_new_n5258_));
AND2X2 AND2X2_247 ( .A(_abc_41356_new_n948_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n949_));
AND2X2 AND2X2_2470 ( .A(_abc_41356_new_n5260_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5261_));
AND2X2 AND2X2_2471 ( .A(_abc_41356_new_n3432_), .B(rdatahold_4_), .Y(_abc_41356_new_n5263_));
AND2X2 AND2X2_2472 ( .A(_abc_41356_new_n3430_), .B(regfil_4__4_), .Y(_abc_41356_new_n5264_));
AND2X2 AND2X2_2473 ( .A(_abc_41356_new_n5229_), .B(_abc_41356_new_n1738_), .Y(_abc_41356_new_n5266_));
AND2X2 AND2X2_2474 ( .A(_abc_41356_new_n5267_), .B(sp_12_), .Y(_abc_41356_new_n5268_));
AND2X2 AND2X2_2475 ( .A(_abc_41356_new_n5269_), .B(_abc_41356_new_n4860_), .Y(_abc_41356_new_n5270_));
AND2X2 AND2X2_2476 ( .A(_abc_41356_new_n1218_), .B(sp_12_), .Y(_abc_41356_new_n5271_));
AND2X2 AND2X2_2477 ( .A(_abc_41356_new_n5274_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5275_));
AND2X2 AND2X2_2478 ( .A(_abc_41356_new_n5273_), .B(_abc_41356_new_n5275_), .Y(_abc_41356_new_n5276_));
AND2X2 AND2X2_2479 ( .A(_abc_41356_new_n4830_), .B(waddrhold_12_), .Y(_abc_41356_new_n5277_));
AND2X2 AND2X2_248 ( .A(_abc_41356_new_n954_), .B(_abc_41356_new_n724_), .Y(_abc_41356_new_n955_));
AND2X2 AND2X2_2480 ( .A(_abc_41356_new_n4668_), .B(_abc_41356_new_n5278_), .Y(_abc_41356_new_n5279_));
AND2X2 AND2X2_2481 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5279_), .Y(_abc_41356_new_n5280_));
AND2X2 AND2X2_2482 ( .A(_abc_41356_new_n2243_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5281_));
AND2X2 AND2X2_2483 ( .A(_abc_41356_new_n5281_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5282_));
AND2X2 AND2X2_2484 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5287_), .Y(_abc_41356_new_n5288_));
AND2X2 AND2X2_2485 ( .A(_abc_41356_new_n5286_), .B(_abc_41356_new_n5288_), .Y(_abc_41356_new_n5289_));
AND2X2 AND2X2_2486 ( .A(_abc_41356_new_n5290_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5291_));
AND2X2 AND2X2_2487 ( .A(_abc_41356_new_n5254_), .B(waddrhold_12_), .Y(_abc_41356_new_n5292_));
AND2X2 AND2X2_2488 ( .A(_abc_41356_new_n519_), .B(_abc_41356_new_n3426_), .Y(_abc_41356_new_n5295_));
AND2X2 AND2X2_2489 ( .A(_abc_41356_new_n5294_), .B(_abc_41356_new_n5295_), .Y(_abc_41356_new_n5296_));
AND2X2 AND2X2_249 ( .A(_abc_41356_new_n953_), .B(_abc_41356_new_n955_), .Y(_abc_41356_new_n956_));
AND2X2 AND2X2_2490 ( .A(_abc_41356_new_n5296_), .B(_abc_41356_new_n5293_), .Y(_abc_41356_new_n5297_));
AND2X2 AND2X2_2491 ( .A(_abc_41356_new_n4821_), .B(waddrhold_12_), .Y(_abc_41356_new_n5298_));
AND2X2 AND2X2_2492 ( .A(_abc_41356_new_n3432_), .B(rdatahold_5_), .Y(_abc_41356_new_n5301_));
AND2X2 AND2X2_2493 ( .A(_abc_41356_new_n3430_), .B(regfil_4__5_), .Y(_abc_41356_new_n5302_));
AND2X2 AND2X2_2494 ( .A(_abc_41356_new_n5304_), .B(sp_13_), .Y(_abc_41356_new_n5305_));
AND2X2 AND2X2_2495 ( .A(_abc_41356_new_n5266_), .B(_abc_41356_new_n1826_), .Y(_abc_41356_new_n5306_));
AND2X2 AND2X2_2496 ( .A(_abc_41356_new_n5307_), .B(_abc_41356_new_n4860_), .Y(_abc_41356_new_n5308_));
AND2X2 AND2X2_2497 ( .A(_abc_41356_new_n1218_), .B(sp_13_), .Y(_abc_41356_new_n5309_));
AND2X2 AND2X2_2498 ( .A(_abc_41356_new_n5312_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5313_));
AND2X2 AND2X2_2499 ( .A(_abc_41356_new_n5311_), .B(_abc_41356_new_n5313_), .Y(_abc_41356_new_n5314_));
AND2X2 AND2X2_25 ( .A(_abc_41356_new_n537_), .B(_abc_41356_new_n533_), .Y(_abc_41356_new_n538_));
AND2X2 AND2X2_250 ( .A(_abc_41356_new_n555_), .B(regfil_7__3_), .Y(_abc_41356_new_n957_));
AND2X2 AND2X2_2500 ( .A(_abc_41356_new_n4830_), .B(waddrhold_13_), .Y(_abc_41356_new_n5315_));
AND2X2 AND2X2_2501 ( .A(_abc_41356_new_n2284_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5316_));
AND2X2 AND2X2_2502 ( .A(_abc_41356_new_n5316_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5317_));
AND2X2 AND2X2_2503 ( .A(_abc_41356_new_n4705_), .B(_abc_41356_new_n5318_), .Y(_abc_41356_new_n5319_));
AND2X2 AND2X2_2504 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5319_), .Y(_abc_41356_new_n5320_));
AND2X2 AND2X2_2505 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5325_), .Y(_abc_41356_new_n5326_));
AND2X2 AND2X2_2506 ( .A(_abc_41356_new_n5324_), .B(_abc_41356_new_n5326_), .Y(_abc_41356_new_n5327_));
AND2X2 AND2X2_2507 ( .A(_abc_41356_new_n5328_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5329_));
AND2X2 AND2X2_2508 ( .A(_abc_41356_new_n4821_), .B(waddrhold_13_), .Y(_abc_41356_new_n5330_));
AND2X2 AND2X2_2509 ( .A(_abc_41356_new_n5292_), .B(waddrhold_13_), .Y(_abc_41356_new_n5332_));
AND2X2 AND2X2_251 ( .A(_abc_41356_new_n961_), .B(_abc_41356_new_n958_), .Y(_abc_41356_new_n962_));
AND2X2 AND2X2_2510 ( .A(_abc_41356_new_n5333_), .B(_abc_41356_new_n5331_), .Y(_abc_41356_new_n5334_));
AND2X2 AND2X2_2511 ( .A(_abc_41356_new_n5334_), .B(_abc_41356_new_n5295_), .Y(_abc_41356_new_n5335_));
AND2X2 AND2X2_2512 ( .A(_abc_41356_new_n3432_), .B(rdatahold_6_), .Y(_abc_41356_new_n5338_));
AND2X2 AND2X2_2513 ( .A(_abc_41356_new_n3430_), .B(regfil_4__6_), .Y(_abc_41356_new_n5339_));
AND2X2 AND2X2_2514 ( .A(_abc_41356_new_n5306_), .B(_abc_41356_new_n1902_), .Y(_abc_41356_new_n5341_));
AND2X2 AND2X2_2515 ( .A(_abc_41356_new_n5342_), .B(sp_14_), .Y(_abc_41356_new_n5343_));
AND2X2 AND2X2_2516 ( .A(_abc_41356_new_n5344_), .B(_abc_41356_new_n4860_), .Y(_abc_41356_new_n5345_));
AND2X2 AND2X2_2517 ( .A(_abc_41356_new_n1218_), .B(sp_14_), .Y(_abc_41356_new_n5346_));
AND2X2 AND2X2_2518 ( .A(_abc_41356_new_n5349_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5350_));
AND2X2 AND2X2_2519 ( .A(_abc_41356_new_n5348_), .B(_abc_41356_new_n5350_), .Y(_abc_41356_new_n5351_));
AND2X2 AND2X2_252 ( .A(_abc_41356_new_n530_), .B(regfil_7__5_), .Y(_abc_41356_new_n963_));
AND2X2 AND2X2_2520 ( .A(_abc_41356_new_n4830_), .B(waddrhold_14_), .Y(_abc_41356_new_n5352_));
AND2X2 AND2X2_2521 ( .A(_abc_41356_new_n2320_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5353_));
AND2X2 AND2X2_2522 ( .A(_abc_41356_new_n5353_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5354_));
AND2X2 AND2X2_2523 ( .A(_abc_41356_new_n4742_), .B(_abc_41356_new_n5355_), .Y(_abc_41356_new_n5356_));
AND2X2 AND2X2_2524 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5356_), .Y(_abc_41356_new_n5357_));
AND2X2 AND2X2_2525 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5362_), .Y(_abc_41356_new_n5363_));
AND2X2 AND2X2_2526 ( .A(_abc_41356_new_n5361_), .B(_abc_41356_new_n5363_), .Y(_abc_41356_new_n5364_));
AND2X2 AND2X2_2527 ( .A(_abc_41356_new_n5365_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5366_));
AND2X2 AND2X2_2528 ( .A(_abc_41356_new_n4821_), .B(waddrhold_14_), .Y(_abc_41356_new_n5368_));
AND2X2 AND2X2_2529 ( .A(_abc_41356_new_n5332_), .B(waddrhold_14_), .Y(_abc_41356_new_n5369_));
AND2X2 AND2X2_253 ( .A(_abc_41356_new_n967_), .B(_abc_41356_new_n964_), .Y(_abc_41356_new_n968_));
AND2X2 AND2X2_2530 ( .A(_abc_41356_new_n5370_), .B(_abc_41356_new_n5295_), .Y(_abc_41356_new_n5371_));
AND2X2 AND2X2_2531 ( .A(_abc_41356_new_n5372_), .B(_abc_41356_new_n5367_), .Y(_abc_41356_new_n5373_));
AND2X2 AND2X2_2532 ( .A(_abc_41356_new_n3432_), .B(rdatahold_7_), .Y(_abc_41356_new_n5375_));
AND2X2 AND2X2_2533 ( .A(_abc_41356_new_n3430_), .B(regfil_4__7_), .Y(_abc_41356_new_n5376_));
AND2X2 AND2X2_2534 ( .A(_abc_41356_new_n5380_), .B(_abc_41356_new_n5378_), .Y(_abc_41356_new_n5381_));
AND2X2 AND2X2_2535 ( .A(_abc_41356_new_n5381_), .B(_abc_41356_new_n4860_), .Y(_abc_41356_new_n5382_));
AND2X2 AND2X2_2536 ( .A(_abc_41356_new_n1218_), .B(sp_15_), .Y(_abc_41356_new_n5383_));
AND2X2 AND2X2_2537 ( .A(_abc_41356_new_n5386_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n5387_));
AND2X2 AND2X2_2538 ( .A(_abc_41356_new_n5385_), .B(_abc_41356_new_n5387_), .Y(_abc_41356_new_n5388_));
AND2X2 AND2X2_2539 ( .A(_abc_41356_new_n4830_), .B(waddrhold_15_), .Y(_abc_41356_new_n5389_));
AND2X2 AND2X2_254 ( .A(_abc_41356_new_n962_), .B(_abc_41356_new_n968_), .Y(_abc_41356_new_n969_));
AND2X2 AND2X2_2540 ( .A(_abc_41356_new_n2360_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5390_));
AND2X2 AND2X2_2541 ( .A(_abc_41356_new_n5390_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n5391_));
AND2X2 AND2X2_2542 ( .A(_abc_41356_new_n4782_), .B(_abc_41356_new_n5392_), .Y(_abc_41356_new_n5393_));
AND2X2 AND2X2_2543 ( .A(_abc_41356_new_n4838_), .B(_abc_41356_new_n5393_), .Y(_abc_41356_new_n5394_));
AND2X2 AND2X2_2544 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n5399_), .Y(_abc_41356_new_n5400_));
AND2X2 AND2X2_2545 ( .A(_abc_41356_new_n5398_), .B(_abc_41356_new_n5400_), .Y(_abc_41356_new_n5401_));
AND2X2 AND2X2_2546 ( .A(_abc_41356_new_n5402_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5403_));
AND2X2 AND2X2_2547 ( .A(_abc_41356_new_n5369_), .B(waddrhold_15_), .Y(_abc_41356_new_n5404_));
AND2X2 AND2X2_2548 ( .A(_abc_41356_new_n5406_), .B(_abc_41356_new_n5295_), .Y(_abc_41356_new_n5407_));
AND2X2 AND2X2_2549 ( .A(_abc_41356_new_n5407_), .B(_abc_41356_new_n5405_), .Y(_abc_41356_new_n5408_));
AND2X2 AND2X2_255 ( .A(_abc_41356_new_n712_), .B(regfil_7__4_), .Y(_abc_41356_new_n970_));
AND2X2 AND2X2_2550 ( .A(_abc_41356_new_n4821_), .B(waddrhold_15_), .Y(_abc_41356_new_n5409_));
AND2X2 AND2X2_2551 ( .A(_abc_41356_new_n2388_), .B(_abc_41356_new_n607_), .Y(_abc_41356_new_n5413_));
AND2X2 AND2X2_2552 ( .A(_abc_41356_new_n5414_), .B(_abc_41356_new_n5412_), .Y(_abc_41356_new_n5415_));
AND2X2 AND2X2_2553 ( .A(_abc_41356_new_n5415_), .B(\data[0] ), .Y(_abc_41356_new_n5416_));
AND2X2 AND2X2_2554 ( .A(_abc_41356_new_n5295_), .B(wdatahold_0_), .Y(_abc_41356_new_n5417_));
AND2X2 AND2X2_2555 ( .A(_abc_41356_new_n5413_), .B(regfil_7__0_), .Y(_abc_41356_new_n5418_));
AND2X2 AND2X2_2556 ( .A(_abc_41356_new_n5415_), .B(\data[1] ), .Y(_abc_41356_new_n5421_));
AND2X2 AND2X2_2557 ( .A(_abc_41356_new_n5295_), .B(wdatahold_1_), .Y(_abc_41356_new_n5422_));
AND2X2 AND2X2_2558 ( .A(_abc_41356_new_n5413_), .B(regfil_7__1_), .Y(_abc_41356_new_n5423_));
AND2X2 AND2X2_2559 ( .A(_abc_41356_new_n5415_), .B(\data[2] ), .Y(_abc_41356_new_n5426_));
AND2X2 AND2X2_256 ( .A(_abc_41356_new_n718_), .B(\data[4] ), .Y(_abc_41356_new_n972_));
AND2X2 AND2X2_2560 ( .A(_abc_41356_new_n5295_), .B(wdatahold_2_), .Y(_abc_41356_new_n5427_));
AND2X2 AND2X2_2561 ( .A(_abc_41356_new_n5413_), .B(regfil_7__2_), .Y(_abc_41356_new_n5428_));
AND2X2 AND2X2_2562 ( .A(_abc_41356_new_n5415_), .B(\data[3] ), .Y(_abc_41356_new_n5431_));
AND2X2 AND2X2_2563 ( .A(_abc_41356_new_n5295_), .B(wdatahold_3_), .Y(_abc_41356_new_n5432_));
AND2X2 AND2X2_2564 ( .A(_abc_41356_new_n5413_), .B(regfil_7__3_), .Y(_abc_41356_new_n5433_));
AND2X2 AND2X2_2565 ( .A(_abc_41356_new_n5415_), .B(\data[4] ), .Y(_abc_41356_new_n5436_));
AND2X2 AND2X2_2566 ( .A(_abc_41356_new_n5295_), .B(wdatahold_4_), .Y(_abc_41356_new_n5437_));
AND2X2 AND2X2_2567 ( .A(_abc_41356_new_n5413_), .B(regfil_7__4_), .Y(_abc_41356_new_n5438_));
AND2X2 AND2X2_2568 ( .A(_abc_41356_new_n5415_), .B(\data[5] ), .Y(_abc_41356_new_n5441_));
AND2X2 AND2X2_2569 ( .A(_abc_41356_new_n5295_), .B(wdatahold_5_), .Y(_abc_41356_new_n5442_));
AND2X2 AND2X2_257 ( .A(_abc_41356_new_n512_), .B(rdatahold_4_), .Y(_abc_41356_new_n977_));
AND2X2 AND2X2_2570 ( .A(_abc_41356_new_n5413_), .B(regfil_7__5_), .Y(_abc_41356_new_n5443_));
AND2X2 AND2X2_2571 ( .A(_abc_41356_new_n5415_), .B(\data[6] ), .Y(_abc_41356_new_n5446_));
AND2X2 AND2X2_2572 ( .A(_abc_41356_new_n5295_), .B(wdatahold_6_), .Y(_abc_41356_new_n5447_));
AND2X2 AND2X2_2573 ( .A(_abc_41356_new_n5413_), .B(regfil_7__6_), .Y(_abc_41356_new_n5448_));
AND2X2 AND2X2_2574 ( .A(_abc_41356_new_n5415_), .B(\data[7] ), .Y(_abc_41356_new_n5451_));
AND2X2 AND2X2_2575 ( .A(_abc_41356_new_n5295_), .B(wdatahold_7_), .Y(_abc_41356_new_n5452_));
AND2X2 AND2X2_2576 ( .A(_abc_41356_new_n5413_), .B(regfil_7__7_), .Y(_abc_41356_new_n5453_));
AND2X2 AND2X2_2577 ( .A(_abc_41356_new_n5456_), .B(regd_0_), .Y(_abc_41356_new_n5457_));
AND2X2 AND2X2_2578 ( .A(_abc_41356_new_n4185_), .B(_abc_41356_new_n677_), .Y(_abc_41356_new_n5458_));
AND2X2 AND2X2_2579 ( .A(_abc_41356_new_n679_), .B(opcode_3_), .Y(_abc_41356_new_n5460_));
AND2X2 AND2X2_258 ( .A(_abc_41356_new_n978_), .B(_abc_41356_new_n976_), .Y(_abc_41356_new_n979_));
AND2X2 AND2X2_2580 ( .A(_abc_41356_new_n5459_), .B(_abc_41356_new_n5461_), .Y(_abc_41356_new_n5462_));
AND2X2 AND2X2_2581 ( .A(_abc_41356_new_n3372_), .B(_abc_41356_new_n2056_), .Y(_abc_41356_new_n5463_));
AND2X2 AND2X2_2582 ( .A(_abc_41356_new_n5467_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5468_));
AND2X2 AND2X2_2583 ( .A(_abc_41356_new_n5468_), .B(_abc_41356_new_n5465_), .Y(_abc_41356_new_n5469_));
AND2X2 AND2X2_2584 ( .A(_abc_41356_new_n5470_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n5471_));
AND2X2 AND2X2_2585 ( .A(_abc_41356_new_n5456_), .B(regd_1_), .Y(_abc_41356_new_n5473_));
AND2X2 AND2X2_2586 ( .A(_abc_41356_new_n2895_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n5475_));
AND2X2 AND2X2_2587 ( .A(_abc_41356_new_n5474_), .B(_abc_41356_new_n5475_), .Y(_abc_41356_new_n5476_));
AND2X2 AND2X2_2588 ( .A(_abc_41356_new_n5478_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5479_));
AND2X2 AND2X2_2589 ( .A(_abc_41356_new_n5479_), .B(_abc_41356_new_n5477_), .Y(_abc_41356_new_n5480_));
AND2X2 AND2X2_259 ( .A(_abc_41356_new_n979_), .B(_abc_41356_new_n973_), .Y(_abc_41356_new_n980_));
AND2X2 AND2X2_2590 ( .A(_abc_41356_new_n5481_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n5482_));
AND2X2 AND2X2_2591 ( .A(_abc_41356_new_n5456_), .B(regd_2_), .Y(_abc_41356_new_n5484_));
AND2X2 AND2X2_2592 ( .A(_abc_41356_new_n2915_), .B(_abc_41356_new_n679_), .Y(_abc_41356_new_n5486_));
AND2X2 AND2X2_2593 ( .A(_abc_41356_new_n5485_), .B(_abc_41356_new_n5486_), .Y(_abc_41356_new_n5487_));
AND2X2 AND2X2_2594 ( .A(_abc_41356_new_n5489_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5490_));
AND2X2 AND2X2_2595 ( .A(_abc_41356_new_n5490_), .B(_abc_41356_new_n5488_), .Y(_abc_41356_new_n5491_));
AND2X2 AND2X2_2596 ( .A(_abc_41356_new_n5492_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n5493_));
AND2X2 AND2X2_2597 ( .A(_abc_41356_new_n694_), .B(_abc_41356_new_n1209_), .Y(_abc_41356_new_n5495_));
AND2X2 AND2X2_2598 ( .A(_abc_41356_new_n5498_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n5499_));
AND2X2 AND2X2_2599 ( .A(_abc_41356_new_n5497_), .B(_abc_41356_new_n5499_), .Y(_abc_41356_new_n5500_));
AND2X2 AND2X2_26 ( .A(_abc_41356_new_n540_), .B(_abc_41356_new_n513_), .Y(_abc_41356_new_n541_));
AND2X2 AND2X2_260 ( .A(_abc_41356_new_n980_), .B(_abc_41356_new_n971_), .Y(_abc_41356_new_n981_));
AND2X2 AND2X2_2600 ( .A(_abc_41356_new_n1230_), .B(rdatahold2_0_), .Y(_abc_41356_new_n5501_));
AND2X2 AND2X2_2601 ( .A(_abc_41356_new_n5502_), .B(_abc_41356_new_n1248_), .Y(_abc_41356_new_n5503_));
AND2X2 AND2X2_2602 ( .A(_abc_41356_new_n5504_), .B(_abc_41356_new_n5505_), .Y(_abc_41356_new_n5506_));
AND2X2 AND2X2_2603 ( .A(_abc_41356_new_n1287_), .B(_abc_41356_new_n5506_), .Y(_abc_41356_new_n5507_));
AND2X2 AND2X2_2604 ( .A(_abc_41356_new_n5508_), .B(_abc_41356_new_n5509_), .Y(_abc_41356_new_n5510_));
AND2X2 AND2X2_2605 ( .A(_abc_41356_new_n2001_), .B(_abc_41356_new_n5510_), .Y(_abc_41356_new_n5511_));
AND2X2 AND2X2_2606 ( .A(_abc_41356_new_n1422_), .B(_abc_41356_new_n5512_), .Y(_abc_41356_new_n5513_));
AND2X2 AND2X2_2607 ( .A(_abc_41356_new_n1988_), .B(_abc_41356_new_n5513_), .Y(_abc_41356_new_n5514_));
AND2X2 AND2X2_2608 ( .A(_abc_41356_new_n1285_), .B(_abc_41356_new_n1258_), .Y(_abc_41356_new_n5517_));
AND2X2 AND2X2_2609 ( .A(_abc_41356_new_n5519_), .B(_abc_41356_new_n5503_), .Y(_abc_41356_new_n5520_));
AND2X2 AND2X2_261 ( .A(_abc_41356_new_n969_), .B(_abc_41356_new_n981_), .Y(_abc_41356_new_n982_));
AND2X2 AND2X2_2610 ( .A(_abc_41356_new_n1230_), .B(rdatahold2_1_), .Y(_abc_41356_new_n5523_));
AND2X2 AND2X2_2611 ( .A(_abc_41356_new_n5525_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n5526_));
AND2X2 AND2X2_2612 ( .A(_abc_41356_new_n5524_), .B(_abc_41356_new_n5526_), .Y(_abc_41356_new_n5527_));
AND2X2 AND2X2_2613 ( .A(_abc_41356_new_n1216_), .B(_abc_41356_new_n5529_), .Y(_abc_41356_new_n5530_));
AND2X2 AND2X2_2614 ( .A(_abc_41356_new_n1294_), .B(_abc_41356_new_n5532_), .Y(_abc_41356_new_n5533_));
AND2X2 AND2X2_2615 ( .A(_abc_41356_new_n1287_), .B(_abc_41356_new_n5533_), .Y(_abc_41356_new_n5534_));
AND2X2 AND2X2_2616 ( .A(_abc_41356_new_n1418_), .B(regfil_5__0_), .Y(_abc_41356_new_n5536_));
AND2X2 AND2X2_2617 ( .A(_abc_41356_new_n1482_), .B(_abc_41356_new_n1425_), .Y(_abc_41356_new_n5537_));
AND2X2 AND2X2_2618 ( .A(_abc_41356_new_n1665_), .B(_abc_41356_new_n5539_), .Y(_abc_41356_new_n5540_));
AND2X2 AND2X2_2619 ( .A(_abc_41356_new_n5540_), .B(_abc_41356_new_n5537_), .Y(_abc_41356_new_n5541_));
AND2X2 AND2X2_262 ( .A(_abc_41356_new_n918_), .B(regfil_0__5_), .Y(_abc_41356_new_n987_));
AND2X2 AND2X2_2620 ( .A(_abc_41356_new_n5542_), .B(_abc_41356_new_n5543_), .Y(_abc_41356_new_n5544_));
AND2X2 AND2X2_2621 ( .A(_abc_41356_new_n1415_), .B(_abc_41356_new_n5544_), .Y(_abc_41356_new_n5545_));
AND2X2 AND2X2_2622 ( .A(_abc_41356_new_n1219_), .B(_abc_41356_new_n5529_), .Y(_abc_41356_new_n5549_));
AND2X2 AND2X2_2623 ( .A(_abc_41356_new_n5550_), .B(_abc_41356_new_n1217_), .Y(_abc_41356_new_n5551_));
AND2X2 AND2X2_2624 ( .A(_abc_41356_new_n5548_), .B(_abc_41356_new_n5551_), .Y(_abc_41356_new_n5552_));
AND2X2 AND2X2_2625 ( .A(_abc_41356_new_n5553_), .B(_abc_41356_new_n5528_), .Y(_abc_41356_new_n5554_));
AND2X2 AND2X2_2626 ( .A(_abc_41356_new_n5496_), .B(regfil_5__2_), .Y(_abc_41356_new_n5557_));
AND2X2 AND2X2_2627 ( .A(_abc_41356_new_n824_), .B(_abc_41356_new_n5495_), .Y(_abc_41356_new_n5558_));
AND2X2 AND2X2_2628 ( .A(_abc_41356_new_n5559_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n5560_));
AND2X2 AND2X2_2629 ( .A(_abc_41356_new_n1230_), .B(rdatahold2_2_), .Y(_abc_41356_new_n5561_));
AND2X2 AND2X2_263 ( .A(_abc_41356_new_n988_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n989_));
AND2X2 AND2X2_2630 ( .A(_abc_41356_new_n1216_), .B(_abc_41356_new_n5564_), .Y(_abc_41356_new_n5565_));
AND2X2 AND2X2_2631 ( .A(_abc_41356_new_n5565_), .B(_abc_41356_new_n5563_), .Y(_abc_41356_new_n5566_));
AND2X2 AND2X2_2632 ( .A(_abc_41356_new_n5568_), .B(_abc_41356_new_n1257_), .Y(_abc_41356_new_n5569_));
AND2X2 AND2X2_2633 ( .A(_abc_41356_new_n1219_), .B(_abc_41356_new_n5570_), .Y(_abc_41356_new_n5571_));
AND2X2 AND2X2_2634 ( .A(_abc_41356_new_n1296_), .B(_abc_41356_new_n1301_), .Y(_abc_41356_new_n5573_));
AND2X2 AND2X2_2635 ( .A(_abc_41356_new_n5574_), .B(_abc_41356_new_n5575_), .Y(_abc_41356_new_n5576_));
AND2X2 AND2X2_2636 ( .A(_abc_41356_new_n5576_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n5577_));
AND2X2 AND2X2_2637 ( .A(_abc_41356_new_n5578_), .B(_abc_41356_new_n1434_), .Y(_abc_41356_new_n5580_));
AND2X2 AND2X2_2638 ( .A(_abc_41356_new_n5581_), .B(_abc_41356_new_n5579_), .Y(_abc_41356_new_n5582_));
AND2X2 AND2X2_2639 ( .A(_abc_41356_new_n5582_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n5583_));
AND2X2 AND2X2_264 ( .A(_abc_41356_new_n924_), .B(regfil_0__5_), .Y(_abc_41356_new_n991_));
AND2X2 AND2X2_2640 ( .A(_abc_41356_new_n1369_), .B(_abc_41356_new_n1373_), .Y(_abc_41356_new_n5584_));
AND2X2 AND2X2_2641 ( .A(_abc_41356_new_n5585_), .B(_abc_41356_new_n5586_), .Y(_abc_41356_new_n5587_));
AND2X2 AND2X2_2642 ( .A(_abc_41356_new_n5587_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n5588_));
AND2X2 AND2X2_2643 ( .A(_abc_41356_new_n1418_), .B(_abc_41356_new_n1259_), .Y(_abc_41356_new_n5591_));
AND2X2 AND2X2_2644 ( .A(_abc_41356_new_n5590_), .B(_abc_41356_new_n5592_), .Y(_abc_41356_new_n5593_));
AND2X2 AND2X2_2645 ( .A(_abc_41356_new_n5595_), .B(_abc_41356_new_n5572_), .Y(_abc_41356_new_n5596_));
AND2X2 AND2X2_2646 ( .A(_abc_41356_new_n5596_), .B(_abc_41356_new_n5567_), .Y(_abc_41356_new_n5597_));
AND2X2 AND2X2_2647 ( .A(_abc_41356_new_n5598_), .B(_abc_41356_new_n5562_), .Y(_abc_41356_new_n5599_));
AND2X2 AND2X2_2648 ( .A(_abc_41356_new_n5603_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n5604_));
AND2X2 AND2X2_2649 ( .A(_abc_41356_new_n5602_), .B(_abc_41356_new_n5604_), .Y(_abc_41356_new_n5605_));
AND2X2 AND2X2_265 ( .A(_abc_41356_new_n992_), .B(_abc_41356_new_n581_), .Y(_abc_41356_new_n993_));
AND2X2 AND2X2_2650 ( .A(_abc_41356_new_n1230_), .B(rdatahold2_3_), .Y(_abc_41356_new_n5606_));
AND2X2 AND2X2_2651 ( .A(_abc_41356_new_n5563_), .B(regfil_5__3_), .Y(_abc_41356_new_n5608_));
AND2X2 AND2X2_2652 ( .A(_abc_41356_new_n1216_), .B(_abc_41356_new_n5609_), .Y(_abc_41356_new_n5610_));
AND2X2 AND2X2_2653 ( .A(_abc_41356_new_n5574_), .B(_abc_41356_new_n5612_), .Y(_abc_41356_new_n5613_));
AND2X2 AND2X2_2654 ( .A(_abc_41356_new_n5615_), .B(_abc_41356_new_n5616_), .Y(_abc_41356_new_n5617_));
AND2X2 AND2X2_2655 ( .A(_abc_41356_new_n5617_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n5618_));
AND2X2 AND2X2_2656 ( .A(_abc_41356_new_n1418_), .B(regfil_5__2_), .Y(_abc_41356_new_n5620_));
AND2X2 AND2X2_2657 ( .A(_abc_41356_new_n5581_), .B(_abc_41356_new_n5621_), .Y(_abc_41356_new_n5622_));
AND2X2 AND2X2_2658 ( .A(_abc_41356_new_n5624_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n5625_));
AND2X2 AND2X2_2659 ( .A(_abc_41356_new_n5626_), .B(_abc_41356_new_n1665_), .Y(_abc_41356_new_n5627_));
AND2X2 AND2X2_266 ( .A(_abc_41356_new_n993_), .B(_abc_41356_new_n990_), .Y(_abc_41356_new_n994_));
AND2X2 AND2X2_2660 ( .A(_abc_41356_new_n5625_), .B(_abc_41356_new_n5627_), .Y(_abc_41356_new_n5628_));
AND2X2 AND2X2_2661 ( .A(_abc_41356_new_n5585_), .B(_abc_41356_new_n5629_), .Y(_abc_41356_new_n5630_));
AND2X2 AND2X2_2662 ( .A(_abc_41356_new_n5633_), .B(_abc_41356_new_n5631_), .Y(_abc_41356_new_n5634_));
AND2X2 AND2X2_2663 ( .A(_abc_41356_new_n5634_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n5635_));
AND2X2 AND2X2_2664 ( .A(_abc_41356_new_n5639_), .B(_abc_41356_new_n1256_), .Y(_abc_41356_new_n5640_));
AND2X2 AND2X2_2665 ( .A(_abc_41356_new_n1219_), .B(_abc_41356_new_n5641_), .Y(_abc_41356_new_n5642_));
AND2X2 AND2X2_2666 ( .A(_abc_41356_new_n5638_), .B(_abc_41356_new_n5643_), .Y(_abc_41356_new_n5644_));
AND2X2 AND2X2_2667 ( .A(_abc_41356_new_n5645_), .B(_abc_41356_new_n5607_), .Y(_abc_41356_new_n5646_));
AND2X2 AND2X2_2668 ( .A(_abc_41356_new_n5650_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n5651_));
AND2X2 AND2X2_2669 ( .A(_abc_41356_new_n5649_), .B(_abc_41356_new_n5651_), .Y(_abc_41356_new_n5652_));
AND2X2 AND2X2_267 ( .A(_abc_41356_new_n642_), .B(rdatahold_5_), .Y(_abc_41356_new_n995_));
AND2X2 AND2X2_2670 ( .A(_abc_41356_new_n1230_), .B(rdatahold2_4_), .Y(_abc_41356_new_n5653_));
AND2X2 AND2X2_2671 ( .A(_abc_41356_new_n5655_), .B(regfil_5__4_), .Y(_abc_41356_new_n5656_));
AND2X2 AND2X2_2672 ( .A(_abc_41356_new_n5657_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n5658_));
AND2X2 AND2X2_2673 ( .A(_abc_41356_new_n1376_), .B(_abc_41356_new_n1393_), .Y(_abc_41356_new_n5661_));
AND2X2 AND2X2_2674 ( .A(_abc_41356_new_n5662_), .B(_abc_41356_new_n5660_), .Y(_abc_41356_new_n5663_));
AND2X2 AND2X2_2675 ( .A(_abc_41356_new_n5663_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n5664_));
AND2X2 AND2X2_2676 ( .A(_abc_41356_new_n5665_), .B(_abc_41356_new_n1455_), .Y(_abc_41356_new_n5666_));
AND2X2 AND2X2_2677 ( .A(_abc_41356_new_n5667_), .B(_abc_41356_new_n5668_), .Y(_abc_41356_new_n5669_));
AND2X2 AND2X2_2678 ( .A(_abc_41356_new_n5669_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n5670_));
AND2X2 AND2X2_2679 ( .A(_abc_41356_new_n1418_), .B(_abc_41356_new_n1256_), .Y(_abc_41356_new_n5673_));
AND2X2 AND2X2_268 ( .A(_abc_41356_new_n619_), .B(regfil_4__5_), .Y(_abc_41356_new_n996_));
AND2X2 AND2X2_2680 ( .A(_abc_41356_new_n5672_), .B(_abc_41356_new_n5674_), .Y(_abc_41356_new_n5675_));
AND2X2 AND2X2_2681 ( .A(_abc_41356_new_n1311_), .B(_abc_41356_new_n1328_), .Y(_abc_41356_new_n5676_));
AND2X2 AND2X2_2682 ( .A(_abc_41356_new_n5677_), .B(_abc_41356_new_n5678_), .Y(_abc_41356_new_n5679_));
AND2X2 AND2X2_2683 ( .A(_abc_41356_new_n5679_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n5680_));
AND2X2 AND2X2_2684 ( .A(_abc_41356_new_n5683_), .B(_abc_41356_new_n1255_), .Y(_abc_41356_new_n5684_));
AND2X2 AND2X2_2685 ( .A(_abc_41356_new_n5685_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n5686_));
AND2X2 AND2X2_2686 ( .A(_abc_41356_new_n5682_), .B(_abc_41356_new_n5687_), .Y(_abc_41356_new_n5688_));
AND2X2 AND2X2_2687 ( .A(_abc_41356_new_n5689_), .B(_abc_41356_new_n5654_), .Y(_abc_41356_new_n5690_));
AND2X2 AND2X2_2688 ( .A(_abc_41356_new_n5694_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n5695_));
AND2X2 AND2X2_2689 ( .A(_abc_41356_new_n5693_), .B(_abc_41356_new_n5695_), .Y(_abc_41356_new_n5696_));
AND2X2 AND2X2_269 ( .A(_abc_41356_new_n616_), .B(regfil_5__5_), .Y(_abc_41356_new_n997_));
AND2X2 AND2X2_2690 ( .A(_abc_41356_new_n1230_), .B(rdatahold2_5_), .Y(_abc_41356_new_n5697_));
AND2X2 AND2X2_2691 ( .A(_abc_41356_new_n5699_), .B(regfil_5__5_), .Y(_abc_41356_new_n5700_));
AND2X2 AND2X2_2692 ( .A(_abc_41356_new_n5701_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n5702_));
AND2X2 AND2X2_2693 ( .A(_abc_41356_new_n5677_), .B(_abc_41356_new_n5704_), .Y(_abc_41356_new_n5705_));
AND2X2 AND2X2_2694 ( .A(_abc_41356_new_n5709_), .B(_abc_41356_new_n5707_), .Y(_abc_41356_new_n5710_));
AND2X2 AND2X2_2695 ( .A(_abc_41356_new_n5710_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n5711_));
AND2X2 AND2X2_2696 ( .A(_abc_41356_new_n5662_), .B(_abc_41356_new_n1391_), .Y(_abc_41356_new_n5713_));
AND2X2 AND2X2_2697 ( .A(_abc_41356_new_n5715_), .B(_abc_41356_new_n5717_), .Y(_abc_41356_new_n5718_));
AND2X2 AND2X2_2698 ( .A(_abc_41356_new_n5667_), .B(_abc_41356_new_n1453_), .Y(_abc_41356_new_n5720_));
AND2X2 AND2X2_2699 ( .A(_abc_41356_new_n5724_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n5725_));
AND2X2 AND2X2_27 ( .A(_abc_41356_new_n545_), .B(opcode_2_), .Y(_abc_41356_new_n546_));
AND2X2 AND2X2_270 ( .A(_abc_41356_new_n526_), .B(regfil_7__5_), .Y(_abc_41356_new_n999_));
AND2X2 AND2X2_2700 ( .A(_abc_41356_new_n5725_), .B(_abc_41356_new_n5722_), .Y(_abc_41356_new_n5726_));
AND2X2 AND2X2_2701 ( .A(_abc_41356_new_n5727_), .B(_abc_41356_new_n5719_), .Y(_abc_41356_new_n5728_));
AND2X2 AND2X2_2702 ( .A(_abc_41356_new_n1418_), .B(regfil_5__4_), .Y(_abc_41356_new_n5729_));
AND2X2 AND2X2_2703 ( .A(_abc_41356_new_n5732_), .B(_abc_41356_new_n5733_), .Y(_abc_41356_new_n5734_));
AND2X2 AND2X2_2704 ( .A(_abc_41356_new_n5735_), .B(_abc_41356_new_n1217_), .Y(_abc_41356_new_n5736_));
AND2X2 AND2X2_2705 ( .A(_abc_41356_new_n5731_), .B(_abc_41356_new_n5736_), .Y(_abc_41356_new_n5737_));
AND2X2 AND2X2_2706 ( .A(_abc_41356_new_n5738_), .B(_abc_41356_new_n5698_), .Y(_abc_41356_new_n5739_));
AND2X2 AND2X2_2707 ( .A(_abc_41356_new_n1230_), .B(rdatahold2_6_), .Y(_abc_41356_new_n5742_));
AND2X2 AND2X2_2708 ( .A(_abc_41356_new_n5744_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n5745_));
AND2X2 AND2X2_2709 ( .A(_abc_41356_new_n5743_), .B(_abc_41356_new_n5745_), .Y(_abc_41356_new_n5746_));
AND2X2 AND2X2_271 ( .A(_abc_41356_new_n623_), .B(regfil_6__5_), .Y(_abc_41356_new_n1000_));
AND2X2 AND2X2_2710 ( .A(_abc_41356_new_n5748_), .B(regfil_5__6_), .Y(_abc_41356_new_n5749_));
AND2X2 AND2X2_2711 ( .A(_abc_41356_new_n5750_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n5751_));
AND2X2 AND2X2_2712 ( .A(_abc_41356_new_n1376_), .B(_abc_41356_new_n1394_), .Y(_abc_41356_new_n5753_));
AND2X2 AND2X2_2713 ( .A(_abc_41356_new_n5754_), .B(_abc_41356_new_n1384_), .Y(_abc_41356_new_n5755_));
AND2X2 AND2X2_2714 ( .A(_abc_41356_new_n5756_), .B(_abc_41356_new_n5757_), .Y(_abc_41356_new_n5758_));
AND2X2 AND2X2_2715 ( .A(_abc_41356_new_n5758_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n5759_));
AND2X2 AND2X2_2716 ( .A(_abc_41356_new_n5665_), .B(_abc_41356_new_n1460_), .Y(_abc_41356_new_n5760_));
AND2X2 AND2X2_2717 ( .A(_abc_41356_new_n5761_), .B(_abc_41356_new_n1450_), .Y(_abc_41356_new_n5763_));
AND2X2 AND2X2_2718 ( .A(_abc_41356_new_n5764_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n5765_));
AND2X2 AND2X2_2719 ( .A(_abc_41356_new_n5765_), .B(_abc_41356_new_n5762_), .Y(_abc_41356_new_n5766_));
AND2X2 AND2X2_272 ( .A(_abc_41356_new_n619_), .B(regfil_0__5_), .Y(_abc_41356_new_n1004_));
AND2X2 AND2X2_2720 ( .A(_abc_41356_new_n1418_), .B(_abc_41356_new_n1254_), .Y(_abc_41356_new_n5769_));
AND2X2 AND2X2_2721 ( .A(_abc_41356_new_n5768_), .B(_abc_41356_new_n5770_), .Y(_abc_41356_new_n5771_));
AND2X2 AND2X2_2722 ( .A(_abc_41356_new_n1311_), .B(_abc_41356_new_n1335_), .Y(_abc_41356_new_n5772_));
AND2X2 AND2X2_2723 ( .A(_abc_41356_new_n5773_), .B(_abc_41356_new_n1322_), .Y(_abc_41356_new_n5775_));
AND2X2 AND2X2_2724 ( .A(_abc_41356_new_n5776_), .B(_abc_41356_new_n5774_), .Y(_abc_41356_new_n5777_));
AND2X2 AND2X2_2725 ( .A(_abc_41356_new_n5777_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n5778_));
AND2X2 AND2X2_2726 ( .A(_abc_41356_new_n5781_), .B(_abc_41356_new_n5782_), .Y(_abc_41356_new_n5783_));
AND2X2 AND2X2_2727 ( .A(_abc_41356_new_n5780_), .B(_abc_41356_new_n5784_), .Y(_abc_41356_new_n5785_));
AND2X2 AND2X2_2728 ( .A(_abc_41356_new_n5786_), .B(_abc_41356_new_n5747_), .Y(_abc_41356_new_n5787_));
AND2X2 AND2X2_2729 ( .A(_abc_41356_new_n5496_), .B(regfil_5__7_), .Y(_abc_41356_new_n5790_));
AND2X2 AND2X2_273 ( .A(_abc_41356_new_n616_), .B(regfil_1__5_), .Y(_abc_41356_new_n1005_));
AND2X2 AND2X2_2730 ( .A(_abc_41356_new_n1173_), .B(_abc_41356_new_n5495_), .Y(_abc_41356_new_n5791_));
AND2X2 AND2X2_2731 ( .A(_abc_41356_new_n5792_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n5793_));
AND2X2 AND2X2_2732 ( .A(_abc_41356_new_n1230_), .B(rdatahold2_7_), .Y(_abc_41356_new_n5794_));
AND2X2 AND2X2_2733 ( .A(_abc_41356_new_n5796_), .B(_abc_41356_new_n1248_), .Y(_abc_41356_new_n5797_));
AND2X2 AND2X2_2734 ( .A(_abc_41356_new_n5798_), .B(regfil_5__7_), .Y(_abc_41356_new_n5799_));
AND2X2 AND2X2_2735 ( .A(_abc_41356_new_n5800_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n5801_));
AND2X2 AND2X2_2736 ( .A(_abc_41356_new_n5807_), .B(_abc_41356_new_n5804_), .Y(_abc_41356_new_n5808_));
AND2X2 AND2X2_2737 ( .A(_abc_41356_new_n5808_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n5809_));
AND2X2 AND2X2_2738 ( .A(_abc_41356_new_n1418_), .B(regfil_5__6_), .Y(_abc_41356_new_n5811_));
AND2X2 AND2X2_2739 ( .A(_abc_41356_new_n5764_), .B(_abc_41356_new_n1448_), .Y(_abc_41356_new_n5812_));
AND2X2 AND2X2_274 ( .A(_abc_41356_new_n526_), .B(regfil_3__5_), .Y(_abc_41356_new_n1007_));
AND2X2 AND2X2_2740 ( .A(_abc_41356_new_n5814_), .B(_abc_41356_new_n5816_), .Y(_abc_41356_new_n5817_));
AND2X2 AND2X2_2741 ( .A(_abc_41356_new_n5817_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n5818_));
AND2X2 AND2X2_2742 ( .A(_abc_41356_new_n5756_), .B(_abc_41356_new_n1382_), .Y(_abc_41356_new_n5820_));
AND2X2 AND2X2_2743 ( .A(_abc_41356_new_n5820_), .B(_abc_41356_new_n1380_), .Y(_abc_41356_new_n5821_));
AND2X2 AND2X2_2744 ( .A(_abc_41356_new_n5823_), .B(_abc_41356_new_n5822_), .Y(_abc_41356_new_n5824_));
AND2X2 AND2X2_2745 ( .A(_abc_41356_new_n5819_), .B(_abc_41356_new_n5826_), .Y(_abc_41356_new_n5827_));
AND2X2 AND2X2_2746 ( .A(_abc_41356_new_n5831_), .B(_abc_41356_new_n5830_), .Y(_abc_41356_new_n5832_));
AND2X2 AND2X2_2747 ( .A(_abc_41356_new_n5829_), .B(_abc_41356_new_n5833_), .Y(_abc_41356_new_n5834_));
AND2X2 AND2X2_2748 ( .A(_abc_41356_new_n5835_), .B(_abc_41356_new_n5797_), .Y(_abc_41356_new_n5836_));
AND2X2 AND2X2_2749 ( .A(_abc_41356_new_n3317_), .B(_abc_41356_new_n706_), .Y(_abc_41356_new_n5838_));
AND2X2 AND2X2_275 ( .A(_abc_41356_new_n623_), .B(regfil_2__5_), .Y(_abc_41356_new_n1008_));
AND2X2 AND2X2_2750 ( .A(_abc_41356_new_n522_), .B(_abc_41356_new_n706_), .Y(_abc_41356_new_n5839_));
AND2X2 AND2X2_2751 ( .A(_abc_41356_new_n587_), .B(_abc_41356_new_n610_), .Y(_abc_41356_new_n5842_));
AND2X2 AND2X2_2752 ( .A(_abc_41356_new_n5842_), .B(_abc_41356_new_n518_), .Y(_abc_41356_new_n5843_));
AND2X2 AND2X2_2753 ( .A(_abc_41356_new_n3265_), .B(_abc_41356_new_n5844_), .Y(_abc_41356_new_n5845_));
AND2X2 AND2X2_2754 ( .A(_abc_41356_new_n5841_), .B(_abc_41356_new_n5845_), .Y(_abc_41356_new_n5846_));
AND2X2 AND2X2_2755 ( .A(_abc_41356_new_n5847_), .B(sp_0_), .Y(_abc_41356_new_n5848_));
AND2X2 AND2X2_2756 ( .A(_abc_41356_new_n5849_), .B(sp_0_), .Y(_abc_41356_new_n5850_));
AND2X2 AND2X2_2757 ( .A(_abc_41356_new_n1286_), .B(regfil_5__0_), .Y(_abc_41356_new_n5851_));
AND2X2 AND2X2_2758 ( .A(_abc_41356_new_n2376_), .B(_abc_41356_new_n681_), .Y(_abc_41356_new_n5854_));
AND2X2 AND2X2_2759 ( .A(_abc_41356_new_n5855_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5856_));
AND2X2 AND2X2_276 ( .A(_abc_41356_new_n1003_), .B(_abc_41356_new_n1011_), .Y(_abc_41356_new_n1012_));
AND2X2 AND2X2_2760 ( .A(_abc_41356_new_n5857_), .B(_abc_41356_new_n5853_), .Y(_abc_41356_new_n5858_));
AND2X2 AND2X2_2761 ( .A(_abc_41356_new_n5859_), .B(_abc_41356_new_n5852_), .Y(_abc_41356_new_n5860_));
AND2X2 AND2X2_2762 ( .A(_abc_41356_new_n516_), .B(sp_0_), .Y(_abc_41356_new_n5862_));
AND2X2 AND2X2_2763 ( .A(_abc_41356_new_n5854_), .B(_abc_41356_new_n5862_), .Y(_abc_41356_new_n5863_));
AND2X2 AND2X2_2764 ( .A(_abc_41356_new_n5864_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n5865_));
AND2X2 AND2X2_2765 ( .A(_abc_41356_new_n5861_), .B(_abc_41356_new_n5865_), .Y(_abc_41356_new_n5866_));
AND2X2 AND2X2_2766 ( .A(_abc_41356_new_n5843_), .B(rdatahold2_0_), .Y(_abc_41356_new_n5867_));
AND2X2 AND2X2_2767 ( .A(_abc_41356_new_n5840_), .B(sp_0_), .Y(_abc_41356_new_n5868_));
AND2X2 AND2X2_2768 ( .A(_abc_41356_new_n5870_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5871_));
AND2X2 AND2X2_2769 ( .A(_abc_41356_new_n5847_), .B(sp_1_), .Y(_abc_41356_new_n5873_));
AND2X2 AND2X2_277 ( .A(_abc_41356_new_n1012_), .B(_abc_41356_new_n614_), .Y(_abc_41356_new_n1013_));
AND2X2 AND2X2_2770 ( .A(_abc_41356_new_n5849_), .B(_abc_41356_new_n3362_), .Y(_abc_41356_new_n5874_));
AND2X2 AND2X2_2771 ( .A(_abc_41356_new_n3363_), .B(_abc_41356_new_n5874_), .Y(_abc_41356_new_n5875_));
AND2X2 AND2X2_2772 ( .A(_abc_41356_new_n5875_), .B(sp_1_), .Y(_abc_41356_new_n5876_));
AND2X2 AND2X2_2773 ( .A(_abc_41356_new_n1286_), .B(regfil_5__1_), .Y(_abc_41356_new_n5877_));
AND2X2 AND2X2_2774 ( .A(_abc_41356_new_n3384_), .B(_abc_41356_new_n4857_), .Y(_abc_41356_new_n5879_));
AND2X2 AND2X2_2775 ( .A(_abc_41356_new_n4857_), .B(_abc_41356_new_n5883_), .Y(_abc_41356_new_n5884_));
AND2X2 AND2X2_2776 ( .A(sp_1_), .B(sp_0_), .Y(_abc_41356_new_n5886_));
AND2X2 AND2X2_2777 ( .A(_abc_41356_new_n5885_), .B(_abc_41356_new_n5887_), .Y(_abc_41356_new_n5888_));
AND2X2 AND2X2_2778 ( .A(_abc_41356_new_n2376_), .B(_abc_41356_new_n682_), .Y(_abc_41356_new_n5890_));
AND2X2 AND2X2_2779 ( .A(_abc_41356_new_n5888_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n5891_));
AND2X2 AND2X2_278 ( .A(_abc_41356_new_n612_), .B(alu_res_5_), .Y(_abc_41356_new_n1014_));
AND2X2 AND2X2_2780 ( .A(_abc_41356_new_n5893_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n5894_));
AND2X2 AND2X2_2781 ( .A(_abc_41356_new_n5894_), .B(_abc_41356_new_n5892_), .Y(_abc_41356_new_n5895_));
AND2X2 AND2X2_2782 ( .A(_abc_41356_new_n5895_), .B(_abc_41356_new_n5889_), .Y(_abc_41356_new_n5896_));
AND2X2 AND2X2_2783 ( .A(_abc_41356_new_n5898_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n5899_));
AND2X2 AND2X2_2784 ( .A(_abc_41356_new_n5897_), .B(_abc_41356_new_n5899_), .Y(_abc_41356_new_n5900_));
AND2X2 AND2X2_2785 ( .A(_abc_41356_new_n5881_), .B(_abc_41356_new_n5900_), .Y(_abc_41356_new_n5901_));
AND2X2 AND2X2_2786 ( .A(_abc_41356_new_n5843_), .B(rdatahold2_1_), .Y(_abc_41356_new_n5902_));
AND2X2 AND2X2_2787 ( .A(_abc_41356_new_n5840_), .B(_abc_41356_new_n4857_), .Y(_abc_41356_new_n5903_));
AND2X2 AND2X2_2788 ( .A(_abc_41356_new_n5905_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5906_));
AND2X2 AND2X2_2789 ( .A(_abc_41356_new_n5847_), .B(sp_2_), .Y(_abc_41356_new_n5908_));
AND2X2 AND2X2_279 ( .A(_abc_41356_new_n1015_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n1016_));
AND2X2 AND2X2_2790 ( .A(_abc_41356_new_n5875_), .B(sp_2_), .Y(_abc_41356_new_n5909_));
AND2X2 AND2X2_2791 ( .A(_abc_41356_new_n4859_), .B(_abc_41356_new_n4896_), .Y(_abc_41356_new_n5910_));
AND2X2 AND2X2_2792 ( .A(_abc_41356_new_n1286_), .B(regfil_5__2_), .Y(_abc_41356_new_n5911_));
AND2X2 AND2X2_2793 ( .A(_abc_41356_new_n5912_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n5913_));
AND2X2 AND2X2_2794 ( .A(_abc_41356_new_n5855_), .B(sp_2_), .Y(_abc_41356_new_n5919_));
AND2X2 AND2X2_2795 ( .A(_abc_41356_new_n4895_), .B(sp_0_), .Y(_abc_41356_new_n5920_));
AND2X2 AND2X2_2796 ( .A(_abc_41356_new_n5890_), .B(_abc_41356_new_n5921_), .Y(_abc_41356_new_n5922_));
AND2X2 AND2X2_2797 ( .A(_abc_41356_new_n5923_), .B(_abc_41356_new_n5918_), .Y(_abc_41356_new_n5924_));
AND2X2 AND2X2_2798 ( .A(_abc_41356_new_n5884_), .B(_abc_41356_new_n1298_), .Y(_abc_41356_new_n5925_));
AND2X2 AND2X2_2799 ( .A(_abc_41356_new_n5885_), .B(sp_2_), .Y(_abc_41356_new_n5926_));
AND2X2 AND2X2_28 ( .A(_abc_41356_new_n546_), .B(_abc_41356_new_n526_), .Y(_abc_41356_new_n547_));
AND2X2 AND2X2_280 ( .A(_abc_41356_new_n1021_), .B(_abc_41356_new_n724_), .Y(_abc_41356_new_n1022_));
AND2X2 AND2X2_2800 ( .A(_abc_41356_new_n5927_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n5928_));
AND2X2 AND2X2_2801 ( .A(_abc_41356_new_n5931_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n5932_));
AND2X2 AND2X2_2802 ( .A(_abc_41356_new_n5930_), .B(_abc_41356_new_n5932_), .Y(_abc_41356_new_n5933_));
AND2X2 AND2X2_2803 ( .A(_abc_41356_new_n5917_), .B(_abc_41356_new_n5933_), .Y(_abc_41356_new_n5934_));
AND2X2 AND2X2_2804 ( .A(_abc_41356_new_n5839_), .B(_abc_41356_new_n5912_), .Y(_abc_41356_new_n5935_));
AND2X2 AND2X2_2805 ( .A(_abc_41356_new_n5843_), .B(rdatahold2_2_), .Y(_abc_41356_new_n5936_));
AND2X2 AND2X2_2806 ( .A(_abc_41356_new_n5838_), .B(_abc_41356_new_n4896_), .Y(_abc_41356_new_n5937_));
AND2X2 AND2X2_2807 ( .A(_abc_41356_new_n5940_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5941_));
AND2X2 AND2X2_2808 ( .A(_abc_41356_new_n5847_), .B(sp_3_), .Y(_abc_41356_new_n5943_));
AND2X2 AND2X2_2809 ( .A(_abc_41356_new_n5875_), .B(sp_3_), .Y(_abc_41356_new_n5944_));
AND2X2 AND2X2_281 ( .A(_abc_41356_new_n1020_), .B(_abc_41356_new_n1022_), .Y(_abc_41356_new_n1023_));
AND2X2 AND2X2_2810 ( .A(_abc_41356_new_n4859_), .B(_abc_41356_new_n4933_), .Y(_abc_41356_new_n5945_));
AND2X2 AND2X2_2811 ( .A(_abc_41356_new_n4895_), .B(sp_3_), .Y(_abc_41356_new_n5946_));
AND2X2 AND2X2_2812 ( .A(_abc_41356_new_n5947_), .B(_abc_41356_new_n5948_), .Y(_abc_41356_new_n5949_));
AND2X2 AND2X2_2813 ( .A(_abc_41356_new_n5949_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n5950_));
AND2X2 AND2X2_2814 ( .A(_abc_41356_new_n1286_), .B(regfil_5__3_), .Y(_abc_41356_new_n5951_));
AND2X2 AND2X2_2815 ( .A(_abc_41356_new_n5956_), .B(_abc_41356_new_n5957_), .Y(_abc_41356_new_n5958_));
AND2X2 AND2X2_2816 ( .A(_abc_41356_new_n5958_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n5959_));
AND2X2 AND2X2_2817 ( .A(_abc_41356_new_n5855_), .B(sp_3_), .Y(_abc_41356_new_n5960_));
AND2X2 AND2X2_2818 ( .A(_abc_41356_new_n5920_), .B(sp_3_), .Y(_abc_41356_new_n5962_));
AND2X2 AND2X2_2819 ( .A(_abc_41356_new_n5964_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n5965_));
AND2X2 AND2X2_282 ( .A(_abc_41356_new_n512_), .B(_abc_41356_new_n1024_), .Y(_abc_41356_new_n1025_));
AND2X2 AND2X2_2820 ( .A(_abc_41356_new_n5965_), .B(_abc_41356_new_n5963_), .Y(_abc_41356_new_n5966_));
AND2X2 AND2X2_2821 ( .A(_abc_41356_new_n5969_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n5970_));
AND2X2 AND2X2_2822 ( .A(_abc_41356_new_n5968_), .B(_abc_41356_new_n5970_), .Y(_abc_41356_new_n5971_));
AND2X2 AND2X2_2823 ( .A(_abc_41356_new_n5955_), .B(_abc_41356_new_n5971_), .Y(_abc_41356_new_n5972_));
AND2X2 AND2X2_2824 ( .A(_abc_41356_new_n5839_), .B(_abc_41356_new_n5949_), .Y(_abc_41356_new_n5973_));
AND2X2 AND2X2_2825 ( .A(_abc_41356_new_n4933_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n5974_));
AND2X2 AND2X2_2826 ( .A(_abc_41356_new_n5843_), .B(rdatahold2_3_), .Y(_abc_41356_new_n5975_));
AND2X2 AND2X2_2827 ( .A(_abc_41356_new_n5978_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n5979_));
AND2X2 AND2X2_2828 ( .A(_abc_41356_new_n5847_), .B(sp_4_), .Y(_abc_41356_new_n5981_));
AND2X2 AND2X2_2829 ( .A(_abc_41356_new_n5875_), .B(sp_4_), .Y(_abc_41356_new_n5982_));
AND2X2 AND2X2_283 ( .A(_abc_41356_new_n530_), .B(regfil_7__6_), .Y(_abc_41356_new_n1027_));
AND2X2 AND2X2_2830 ( .A(_abc_41356_new_n4859_), .B(_abc_41356_new_n4971_), .Y(_abc_41356_new_n5983_));
AND2X2 AND2X2_2831 ( .A(_abc_41356_new_n5946_), .B(sp_4_), .Y(_abc_41356_new_n5984_));
AND2X2 AND2X2_2832 ( .A(_abc_41356_new_n5985_), .B(_abc_41356_new_n5986_), .Y(_abc_41356_new_n5987_));
AND2X2 AND2X2_2833 ( .A(_abc_41356_new_n5987_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n5988_));
AND2X2 AND2X2_2834 ( .A(_abc_41356_new_n1286_), .B(regfil_5__4_), .Y(_abc_41356_new_n5989_));
AND2X2 AND2X2_2835 ( .A(_abc_41356_new_n5855_), .B(sp_4_), .Y(_abc_41356_new_n5994_));
AND2X2 AND2X2_2836 ( .A(_abc_41356_new_n4967_), .B(_abc_41356_new_n5883_), .Y(_abc_41356_new_n5995_));
AND2X2 AND2X2_2837 ( .A(_abc_41356_new_n5995_), .B(_abc_41356_new_n1325_), .Y(_abc_41356_new_n5996_));
AND2X2 AND2X2_2838 ( .A(_abc_41356_new_n5997_), .B(sp_4_), .Y(_abc_41356_new_n5998_));
AND2X2 AND2X2_2839 ( .A(_abc_41356_new_n5999_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6000_));
AND2X2 AND2X2_284 ( .A(_abc_41356_new_n555_), .B(_abc_41356_new_n893_), .Y(_abc_41356_new_n1030_));
AND2X2 AND2X2_2840 ( .A(_abc_41356_new_n5962_), .B(sp_4_), .Y(_abc_41356_new_n6002_));
AND2X2 AND2X2_2841 ( .A(_abc_41356_new_n6004_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6005_));
AND2X2 AND2X2_2842 ( .A(_abc_41356_new_n6005_), .B(_abc_41356_new_n6003_), .Y(_abc_41356_new_n6006_));
AND2X2 AND2X2_2843 ( .A(_abc_41356_new_n6009_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6010_));
AND2X2 AND2X2_2844 ( .A(_abc_41356_new_n6008_), .B(_abc_41356_new_n6010_), .Y(_abc_41356_new_n6011_));
AND2X2 AND2X2_2845 ( .A(_abc_41356_new_n5993_), .B(_abc_41356_new_n6011_), .Y(_abc_41356_new_n6012_));
AND2X2 AND2X2_2846 ( .A(_abc_41356_new_n5987_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6013_));
AND2X2 AND2X2_2847 ( .A(_abc_41356_new_n5843_), .B(rdatahold2_4_), .Y(_abc_41356_new_n6014_));
AND2X2 AND2X2_2848 ( .A(_abc_41356_new_n4971_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6016_));
AND2X2 AND2X2_2849 ( .A(_abc_41356_new_n6018_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6019_));
AND2X2 AND2X2_285 ( .A(_abc_41356_new_n1031_), .B(_abc_41356_new_n1029_), .Y(_abc_41356_new_n1032_));
AND2X2 AND2X2_2850 ( .A(_abc_41356_new_n5847_), .B(sp_5_), .Y(_abc_41356_new_n6021_));
AND2X2 AND2X2_2851 ( .A(_abc_41356_new_n6022_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6023_));
AND2X2 AND2X2_2852 ( .A(_abc_41356_new_n6024_), .B(sp_5_), .Y(_abc_41356_new_n6025_));
AND2X2 AND2X2_2853 ( .A(_abc_41356_new_n4859_), .B(_abc_41356_new_n5008_), .Y(_abc_41356_new_n6026_));
AND2X2 AND2X2_2854 ( .A(_abc_41356_new_n5984_), .B(sp_5_), .Y(_abc_41356_new_n6027_));
AND2X2 AND2X2_2855 ( .A(_abc_41356_new_n6028_), .B(_abc_41356_new_n6029_), .Y(_abc_41356_new_n6030_));
AND2X2 AND2X2_2856 ( .A(_abc_41356_new_n6030_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6031_));
AND2X2 AND2X2_2857 ( .A(_abc_41356_new_n1286_), .B(regfil_5__5_), .Y(_abc_41356_new_n6032_));
AND2X2 AND2X2_2858 ( .A(_abc_41356_new_n6034_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n6035_));
AND2X2 AND2X2_2859 ( .A(_abc_41356_new_n6002_), .B(sp_5_), .Y(_abc_41356_new_n6036_));
AND2X2 AND2X2_286 ( .A(_abc_41356_new_n543_), .B(regfil_7__4_), .Y(_abc_41356_new_n1033_));
AND2X2 AND2X2_2860 ( .A(_abc_41356_new_n6038_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6039_));
AND2X2 AND2X2_2861 ( .A(_abc_41356_new_n6039_), .B(_abc_41356_new_n6037_), .Y(_abc_41356_new_n6040_));
AND2X2 AND2X2_2862 ( .A(_abc_41356_new_n6043_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6044_));
AND2X2 AND2X2_2863 ( .A(_abc_41356_new_n6044_), .B(_abc_41356_new_n6042_), .Y(_abc_41356_new_n6045_));
AND2X2 AND2X2_2864 ( .A(_abc_41356_new_n6046_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n6047_));
AND2X2 AND2X2_2865 ( .A(_abc_41356_new_n6049_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6050_));
AND2X2 AND2X2_2866 ( .A(_abc_41356_new_n6030_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6051_));
AND2X2 AND2X2_2867 ( .A(_abc_41356_new_n5008_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6052_));
AND2X2 AND2X2_2868 ( .A(_abc_41356_new_n5843_), .B(rdatahold2_5_), .Y(_abc_41356_new_n6053_));
AND2X2 AND2X2_2869 ( .A(_abc_41356_new_n6056_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6057_));
AND2X2 AND2X2_287 ( .A(_abc_41356_new_n551_), .B(_abc_41356_new_n1034_), .Y(_abc_41356_new_n1035_));
AND2X2 AND2X2_2870 ( .A(_abc_41356_new_n5847_), .B(sp_6_), .Y(_abc_41356_new_n6059_));
AND2X2 AND2X2_2871 ( .A(_abc_41356_new_n6024_), .B(sp_6_), .Y(_abc_41356_new_n6060_));
AND2X2 AND2X2_2872 ( .A(_abc_41356_new_n5042_), .B(_abc_41356_new_n5883_), .Y(_abc_41356_new_n6061_));
AND2X2 AND2X2_2873 ( .A(_abc_41356_new_n6062_), .B(sp_6_), .Y(_abc_41356_new_n6063_));
AND2X2 AND2X2_2874 ( .A(_abc_41356_new_n6064_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6065_));
AND2X2 AND2X2_2875 ( .A(_abc_41356_new_n6036_), .B(sp_6_), .Y(_abc_41356_new_n6066_));
AND2X2 AND2X2_2876 ( .A(_abc_41356_new_n6068_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6069_));
AND2X2 AND2X2_2877 ( .A(_abc_41356_new_n6069_), .B(_abc_41356_new_n6067_), .Y(_abc_41356_new_n6070_));
AND2X2 AND2X2_2878 ( .A(_abc_41356_new_n6071_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n6072_));
AND2X2 AND2X2_2879 ( .A(_abc_41356_new_n6073_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6074_));
AND2X2 AND2X2_288 ( .A(_abc_41356_new_n698_), .B(_abc_41356_new_n701_), .Y(_abc_41356_new_n1037_));
AND2X2 AND2X2_2880 ( .A(_abc_41356_new_n6027_), .B(sp_6_), .Y(_abc_41356_new_n6075_));
AND2X2 AND2X2_2881 ( .A(_abc_41356_new_n6076_), .B(_abc_41356_new_n6077_), .Y(_abc_41356_new_n6078_));
AND2X2 AND2X2_2882 ( .A(_abc_41356_new_n6078_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6079_));
AND2X2 AND2X2_2883 ( .A(_abc_41356_new_n5045_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6080_));
AND2X2 AND2X2_2884 ( .A(_abc_41356_new_n5843_), .B(rdatahold2_6_), .Y(_abc_41356_new_n6081_));
AND2X2 AND2X2_2885 ( .A(_abc_41356_new_n4859_), .B(_abc_41356_new_n5045_), .Y(_abc_41356_new_n6084_));
AND2X2 AND2X2_2886 ( .A(_abc_41356_new_n6078_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6085_));
AND2X2 AND2X2_2887 ( .A(_abc_41356_new_n1286_), .B(regfil_5__6_), .Y(_abc_41356_new_n6086_));
AND2X2 AND2X2_2888 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n6089_));
AND2X2 AND2X2_2889 ( .A(_abc_41356_new_n6088_), .B(_abc_41356_new_n6089_), .Y(_abc_41356_new_n6090_));
AND2X2 AND2X2_289 ( .A(_abc_41356_new_n1037_), .B(_abc_41356_new_n1036_), .Y(_abc_41356_new_n1038_));
AND2X2 AND2X2_2890 ( .A(_abc_41356_new_n6092_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6093_));
AND2X2 AND2X2_2891 ( .A(_abc_41356_new_n5847_), .B(sp_7_), .Y(_abc_41356_new_n6095_));
AND2X2 AND2X2_2892 ( .A(_abc_41356_new_n5875_), .B(sp_7_), .Y(_abc_41356_new_n6096_));
AND2X2 AND2X2_2893 ( .A(_abc_41356_new_n4859_), .B(_abc_41356_new_n5082_), .Y(_abc_41356_new_n6097_));
AND2X2 AND2X2_2894 ( .A(_abc_41356_new_n6075_), .B(sp_7_), .Y(_abc_41356_new_n6098_));
AND2X2 AND2X2_2895 ( .A(_abc_41356_new_n6099_), .B(_abc_41356_new_n6100_), .Y(_abc_41356_new_n6101_));
AND2X2 AND2X2_2896 ( .A(_abc_41356_new_n6101_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6102_));
AND2X2 AND2X2_2897 ( .A(_abc_41356_new_n1286_), .B(regfil_5__7_), .Y(_abc_41356_new_n6103_));
AND2X2 AND2X2_2898 ( .A(_abc_41356_new_n6066_), .B(sp_7_), .Y(_abc_41356_new_n6109_));
AND2X2 AND2X2_2899 ( .A(_abc_41356_new_n6110_), .B(_abc_41356_new_n6108_), .Y(_abc_41356_new_n6111_));
AND2X2 AND2X2_29 ( .A(_abc_41356_new_n547_), .B(_abc_41356_new_n535_), .Y(_abc_41356_new_n548_));
AND2X2 AND2X2_290 ( .A(_abc_41356_new_n1035_), .B(regfil_7__5_), .Y(_abc_41356_new_n1039_));
AND2X2 AND2X2_2900 ( .A(_abc_41356_new_n6111_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6112_));
AND2X2 AND2X2_2901 ( .A(_abc_41356_new_n6113_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6114_));
AND2X2 AND2X2_2902 ( .A(_abc_41356_new_n6115_), .B(sp_7_), .Y(_abc_41356_new_n6116_));
AND2X2 AND2X2_2903 ( .A(_abc_41356_new_n5081_), .B(_abc_41356_new_n5883_), .Y(_abc_41356_new_n6117_));
AND2X2 AND2X2_2904 ( .A(_abc_41356_new_n6117_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6118_));
AND2X2 AND2X2_2905 ( .A(_abc_41356_new_n6122_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6123_));
AND2X2 AND2X2_2906 ( .A(_abc_41356_new_n6121_), .B(_abc_41356_new_n6123_), .Y(_abc_41356_new_n6124_));
AND2X2 AND2X2_2907 ( .A(_abc_41356_new_n6124_), .B(_abc_41356_new_n6107_), .Y(_abc_41356_new_n6125_));
AND2X2 AND2X2_2908 ( .A(_abc_41356_new_n6101_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6126_));
AND2X2 AND2X2_2909 ( .A(_abc_41356_new_n5082_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6127_));
AND2X2 AND2X2_291 ( .A(_abc_41356_new_n1041_), .B(_abc_41356_new_n1032_), .Y(_abc_41356_new_n1042_));
AND2X2 AND2X2_2910 ( .A(_abc_41356_new_n5843_), .B(rdatahold2_7_), .Y(_abc_41356_new_n6128_));
AND2X2 AND2X2_2911 ( .A(_abc_41356_new_n6131_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6132_));
AND2X2 AND2X2_2912 ( .A(_abc_41356_new_n5847_), .B(sp_8_), .Y(_abc_41356_new_n6134_));
AND2X2 AND2X2_2913 ( .A(_abc_41356_new_n5875_), .B(sp_8_), .Y(_abc_41356_new_n6135_));
AND2X2 AND2X2_2914 ( .A(_abc_41356_new_n6098_), .B(sp_8_), .Y(_abc_41356_new_n6136_));
AND2X2 AND2X2_2915 ( .A(_abc_41356_new_n6137_), .B(_abc_41356_new_n6138_), .Y(_abc_41356_new_n6139_));
AND2X2 AND2X2_2916 ( .A(_abc_41356_new_n6139_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6140_));
AND2X2 AND2X2_2917 ( .A(_abc_41356_new_n5119_), .B(_abc_41356_new_n4859_), .Y(_abc_41356_new_n6141_));
AND2X2 AND2X2_2918 ( .A(_abc_41356_new_n1286_), .B(regfil_4__0_), .Y(_abc_41356_new_n6142_));
AND2X2 AND2X2_2919 ( .A(_abc_41356_new_n6109_), .B(sp_8_), .Y(_abc_41356_new_n6148_));
AND2X2 AND2X2_292 ( .A(_abc_41356_new_n1043_), .B(_abc_41356_new_n1026_), .Y(_abc_41356_new_n1044_));
AND2X2 AND2X2_2920 ( .A(_abc_41356_new_n6149_), .B(_abc_41356_new_n6147_), .Y(_abc_41356_new_n6150_));
AND2X2 AND2X2_2921 ( .A(_abc_41356_new_n6150_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6151_));
AND2X2 AND2X2_2922 ( .A(_abc_41356_new_n6152_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6153_));
AND2X2 AND2X2_2923 ( .A(_abc_41356_new_n6154_), .B(sp_8_), .Y(_abc_41356_new_n6155_));
AND2X2 AND2X2_2924 ( .A(_abc_41356_new_n6117_), .B(_abc_41356_new_n1345_), .Y(_abc_41356_new_n6156_));
AND2X2 AND2X2_2925 ( .A(_abc_41356_new_n6156_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6157_));
AND2X2 AND2X2_2926 ( .A(_abc_41356_new_n6161_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6162_));
AND2X2 AND2X2_2927 ( .A(_abc_41356_new_n6160_), .B(_abc_41356_new_n6162_), .Y(_abc_41356_new_n6163_));
AND2X2 AND2X2_2928 ( .A(_abc_41356_new_n6163_), .B(_abc_41356_new_n6146_), .Y(_abc_41356_new_n6164_));
AND2X2 AND2X2_2929 ( .A(_abc_41356_new_n6139_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6165_));
AND2X2 AND2X2_293 ( .A(_abc_41356_new_n712_), .B(_abc_41356_new_n701_), .Y(_abc_41356_new_n1045_));
AND2X2 AND2X2_2930 ( .A(_abc_41356_new_n5119_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6166_));
AND2X2 AND2X2_2931 ( .A(_abc_41356_new_n5843_), .B(rdatahold_0_), .Y(_abc_41356_new_n6167_));
AND2X2 AND2X2_2932 ( .A(_abc_41356_new_n6170_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6171_));
AND2X2 AND2X2_2933 ( .A(_abc_41356_new_n5847_), .B(sp_9_), .Y(_abc_41356_new_n6173_));
AND2X2 AND2X2_2934 ( .A(_abc_41356_new_n6148_), .B(sp_9_), .Y(_abc_41356_new_n6175_));
AND2X2 AND2X2_2935 ( .A(_abc_41356_new_n6176_), .B(_abc_41356_new_n6174_), .Y(_abc_41356_new_n6177_));
AND2X2 AND2X2_2936 ( .A(_abc_41356_new_n6177_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6178_));
AND2X2 AND2X2_2937 ( .A(_abc_41356_new_n6180_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6181_));
AND2X2 AND2X2_2938 ( .A(_abc_41356_new_n5854_), .B(sp_9_), .Y(_abc_41356_new_n6182_));
AND2X2 AND2X2_2939 ( .A(_abc_41356_new_n6184_), .B(_abc_41356_new_n6179_), .Y(_abc_41356_new_n6185_));
AND2X2 AND2X2_294 ( .A(_abc_41356_new_n714_), .B(alu_res_5_), .Y(_abc_41356_new_n1046_));
AND2X2 AND2X2_2940 ( .A(_abc_41356_new_n5156_), .B(_abc_41356_new_n4859_), .Y(_abc_41356_new_n6188_));
AND2X2 AND2X2_2941 ( .A(_abc_41356_new_n1286_), .B(regfil_4__1_), .Y(_abc_41356_new_n6189_));
AND2X2 AND2X2_2942 ( .A(_abc_41356_new_n5875_), .B(sp_9_), .Y(_abc_41356_new_n6192_));
AND2X2 AND2X2_2943 ( .A(_abc_41356_new_n6136_), .B(sp_9_), .Y(_abc_41356_new_n6193_));
AND2X2 AND2X2_2944 ( .A(_abc_41356_new_n6194_), .B(_abc_41356_new_n6195_), .Y(_abc_41356_new_n6196_));
AND2X2 AND2X2_2945 ( .A(_abc_41356_new_n6196_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6197_));
AND2X2 AND2X2_2946 ( .A(_abc_41356_new_n6200_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6201_));
AND2X2 AND2X2_2947 ( .A(_abc_41356_new_n6199_), .B(_abc_41356_new_n6201_), .Y(_abc_41356_new_n6202_));
AND2X2 AND2X2_2948 ( .A(_abc_41356_new_n6187_), .B(_abc_41356_new_n6202_), .Y(_abc_41356_new_n6203_));
AND2X2 AND2X2_2949 ( .A(_abc_41356_new_n6196_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6204_));
AND2X2 AND2X2_295 ( .A(_abc_41356_new_n718_), .B(\data[5] ), .Y(_abc_41356_new_n1047_));
AND2X2 AND2X2_2950 ( .A(_abc_41356_new_n5156_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6205_));
AND2X2 AND2X2_2951 ( .A(_abc_41356_new_n5843_), .B(rdatahold_1_), .Y(_abc_41356_new_n6206_));
AND2X2 AND2X2_2952 ( .A(_abc_41356_new_n6209_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6210_));
AND2X2 AND2X2_2953 ( .A(_abc_41356_new_n5847_), .B(sp_10_), .Y(_abc_41356_new_n6212_));
AND2X2 AND2X2_2954 ( .A(_abc_41356_new_n5190_), .B(_abc_41356_new_n5883_), .Y(_abc_41356_new_n6213_));
AND2X2 AND2X2_2955 ( .A(_abc_41356_new_n6214_), .B(sp_10_), .Y(_abc_41356_new_n6215_));
AND2X2 AND2X2_2956 ( .A(_abc_41356_new_n6216_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6217_));
AND2X2 AND2X2_2957 ( .A(_abc_41356_new_n6193_), .B(sp_10_), .Y(_abc_41356_new_n6218_));
AND2X2 AND2X2_2958 ( .A(_abc_41356_new_n6218_), .B(sp_0_), .Y(_abc_41356_new_n6219_));
AND2X2 AND2X2_2959 ( .A(_abc_41356_new_n6221_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6222_));
AND2X2 AND2X2_296 ( .A(_abc_41356_new_n595_), .B(rdatahold_6_), .Y(_abc_41356_new_n1052_));
AND2X2 AND2X2_2960 ( .A(_abc_41356_new_n6222_), .B(_abc_41356_new_n6220_), .Y(_abc_41356_new_n6223_));
AND2X2 AND2X2_2961 ( .A(_abc_41356_new_n6224_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n6225_));
AND2X2 AND2X2_2962 ( .A(_abc_41356_new_n6024_), .B(sp_10_), .Y(_abc_41356_new_n6226_));
AND2X2 AND2X2_2963 ( .A(_abc_41356_new_n6227_), .B(_abc_41356_new_n6228_), .Y(_abc_41356_new_n6229_));
AND2X2 AND2X2_2964 ( .A(_abc_41356_new_n6229_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6230_));
AND2X2 AND2X2_2965 ( .A(_abc_41356_new_n1286_), .B(regfil_4__2_), .Y(_abc_41356_new_n6231_));
AND2X2 AND2X2_2966 ( .A(_abc_41356_new_n5193_), .B(_abc_41356_new_n4859_), .Y(_abc_41356_new_n6232_));
AND2X2 AND2X2_2967 ( .A(_abc_41356_new_n6234_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n6235_));
AND2X2 AND2X2_2968 ( .A(_abc_41356_new_n6237_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6238_));
AND2X2 AND2X2_2969 ( .A(_abc_41356_new_n6229_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6239_));
AND2X2 AND2X2_297 ( .A(_abc_41356_new_n619_), .B(regfil_4__6_), .Y(_abc_41356_new_n1053_));
AND2X2 AND2X2_2970 ( .A(_abc_41356_new_n5843_), .B(rdatahold_2_), .Y(_abc_41356_new_n6240_));
AND2X2 AND2X2_2971 ( .A(_abc_41356_new_n5193_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6241_));
AND2X2 AND2X2_2972 ( .A(_abc_41356_new_n6244_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6245_));
AND2X2 AND2X2_2973 ( .A(_abc_41356_new_n5847_), .B(sp_11_), .Y(_abc_41356_new_n6247_));
AND2X2 AND2X2_2974 ( .A(_abc_41356_new_n5229_), .B(_abc_41356_new_n5883_), .Y(_abc_41356_new_n6248_));
AND2X2 AND2X2_2975 ( .A(_abc_41356_new_n6249_), .B(sp_11_), .Y(_abc_41356_new_n6250_));
AND2X2 AND2X2_2976 ( .A(_abc_41356_new_n6251_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6252_));
AND2X2 AND2X2_2977 ( .A(_abc_41356_new_n5855_), .B(sp_11_), .Y(_abc_41356_new_n6253_));
AND2X2 AND2X2_2978 ( .A(_abc_41356_new_n6175_), .B(sp_10_), .Y(_abc_41356_new_n6257_));
AND2X2 AND2X2_2979 ( .A(_abc_41356_new_n6257_), .B(sp_11_), .Y(_abc_41356_new_n6258_));
AND2X2 AND2X2_298 ( .A(_abc_41356_new_n616_), .B(regfil_5__6_), .Y(_abc_41356_new_n1054_));
AND2X2 AND2X2_2980 ( .A(_abc_41356_new_n6259_), .B(_abc_41356_new_n6256_), .Y(_abc_41356_new_n6260_));
AND2X2 AND2X2_2981 ( .A(_abc_41356_new_n6260_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6261_));
AND2X2 AND2X2_2982 ( .A(_abc_41356_new_n6218_), .B(sp_11_), .Y(_abc_41356_new_n6263_));
AND2X2 AND2X2_2983 ( .A(_abc_41356_new_n6264_), .B(_abc_41356_new_n6265_), .Y(_abc_41356_new_n6266_));
AND2X2 AND2X2_2984 ( .A(_abc_41356_new_n6266_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6267_));
AND2X2 AND2X2_2985 ( .A(_abc_41356_new_n5230_), .B(_abc_41356_new_n4859_), .Y(_abc_41356_new_n6268_));
AND2X2 AND2X2_2986 ( .A(_abc_41356_new_n5875_), .B(sp_11_), .Y(_abc_41356_new_n6269_));
AND2X2 AND2X2_2987 ( .A(_abc_41356_new_n1286_), .B(regfil_4__3_), .Y(_abc_41356_new_n6270_));
AND2X2 AND2X2_2988 ( .A(_abc_41356_new_n6275_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6276_));
AND2X2 AND2X2_2989 ( .A(_abc_41356_new_n6274_), .B(_abc_41356_new_n6276_), .Y(_abc_41356_new_n6277_));
AND2X2 AND2X2_299 ( .A(_abc_41356_new_n526_), .B(regfil_7__6_), .Y(_abc_41356_new_n1056_));
AND2X2 AND2X2_2990 ( .A(_abc_41356_new_n6277_), .B(_abc_41356_new_n6262_), .Y(_abc_41356_new_n6278_));
AND2X2 AND2X2_2991 ( .A(_abc_41356_new_n6266_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6279_));
AND2X2 AND2X2_2992 ( .A(_abc_41356_new_n5230_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6280_));
AND2X2 AND2X2_2993 ( .A(_abc_41356_new_n5843_), .B(rdatahold_3_), .Y(_abc_41356_new_n6281_));
AND2X2 AND2X2_2994 ( .A(_abc_41356_new_n6284_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6285_));
AND2X2 AND2X2_2995 ( .A(_abc_41356_new_n5847_), .B(sp_12_), .Y(_abc_41356_new_n6287_));
AND2X2 AND2X2_2996 ( .A(_abc_41356_new_n6263_), .B(sp_12_), .Y(_abc_41356_new_n6288_));
AND2X2 AND2X2_2997 ( .A(_abc_41356_new_n6289_), .B(_abc_41356_new_n6290_), .Y(_abc_41356_new_n6291_));
AND2X2 AND2X2_2998 ( .A(_abc_41356_new_n6291_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6292_));
AND2X2 AND2X2_2999 ( .A(_abc_41356_new_n1286_), .B(regfil_4__4_), .Y(_abc_41356_new_n6293_));
AND2X2 AND2X2_3 ( .A(_abc_41356_new_n505_), .B(state_0_), .Y(_abc_41356_new_n506_));
AND2X2 AND2X2_30 ( .A(_abc_41356_new_n548_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n549_));
AND2X2 AND2X2_300 ( .A(_abc_41356_new_n623_), .B(regfil_6__6_), .Y(_abc_41356_new_n1057_));
AND2X2 AND2X2_3000 ( .A(_abc_41356_new_n5269_), .B(_abc_41356_new_n4859_), .Y(_abc_41356_new_n6294_));
AND2X2 AND2X2_3001 ( .A(_abc_41356_new_n6296_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n6297_));
AND2X2 AND2X2_3002 ( .A(_abc_41356_new_n6248_), .B(_abc_41356_new_n1738_), .Y(_abc_41356_new_n6298_));
AND2X2 AND2X2_3003 ( .A(_abc_41356_new_n6299_), .B(sp_12_), .Y(_abc_41356_new_n6300_));
AND2X2 AND2X2_3004 ( .A(_abc_41356_new_n6301_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6302_));
AND2X2 AND2X2_3005 ( .A(_abc_41356_new_n6258_), .B(sp_12_), .Y(_abc_41356_new_n6304_));
AND2X2 AND2X2_3006 ( .A(_abc_41356_new_n6305_), .B(_abc_41356_new_n6303_), .Y(_abc_41356_new_n6306_));
AND2X2 AND2X2_3007 ( .A(_abc_41356_new_n6306_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6307_));
AND2X2 AND2X2_3008 ( .A(_abc_41356_new_n6308_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n6309_));
AND2X2 AND2X2_3009 ( .A(_abc_41356_new_n6024_), .B(sp_12_), .Y(_abc_41356_new_n6310_));
AND2X2 AND2X2_301 ( .A(_abc_41356_new_n619_), .B(regfil_0__6_), .Y(_abc_41356_new_n1061_));
AND2X2 AND2X2_3010 ( .A(_abc_41356_new_n6312_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6313_));
AND2X2 AND2X2_3011 ( .A(_abc_41356_new_n6291_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6314_));
AND2X2 AND2X2_3012 ( .A(_abc_41356_new_n5269_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6315_));
AND2X2 AND2X2_3013 ( .A(_abc_41356_new_n5843_), .B(rdatahold_4_), .Y(_abc_41356_new_n6316_));
AND2X2 AND2X2_3014 ( .A(_abc_41356_new_n6319_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6320_));
AND2X2 AND2X2_3015 ( .A(_abc_41356_new_n5847_), .B(sp_13_), .Y(_abc_41356_new_n6322_));
AND2X2 AND2X2_3016 ( .A(_abc_41356_new_n6288_), .B(sp_13_), .Y(_abc_41356_new_n6323_));
AND2X2 AND2X2_3017 ( .A(_abc_41356_new_n6323_), .B(sp_0_), .Y(_abc_41356_new_n6324_));
AND2X2 AND2X2_3018 ( .A(_abc_41356_new_n6326_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6327_));
AND2X2 AND2X2_3019 ( .A(_abc_41356_new_n6327_), .B(_abc_41356_new_n6325_), .Y(_abc_41356_new_n6328_));
AND2X2 AND2X2_302 ( .A(_abc_41356_new_n616_), .B(regfil_1__6_), .Y(_abc_41356_new_n1062_));
AND2X2 AND2X2_3020 ( .A(_abc_41356_new_n6329_), .B(sp_13_), .Y(_abc_41356_new_n6330_));
AND2X2 AND2X2_3021 ( .A(_abc_41356_new_n5306_), .B(_abc_41356_new_n5883_), .Y(_abc_41356_new_n6331_));
AND2X2 AND2X2_3022 ( .A(_abc_41356_new_n6332_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6333_));
AND2X2 AND2X2_3023 ( .A(_abc_41356_new_n5855_), .B(sp_13_), .Y(_abc_41356_new_n6334_));
AND2X2 AND2X2_3024 ( .A(_abc_41356_new_n6338_), .B(_abc_41356_new_n6339_), .Y(_abc_41356_new_n6340_));
AND2X2 AND2X2_3025 ( .A(_abc_41356_new_n6340_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6341_));
AND2X2 AND2X2_3026 ( .A(_abc_41356_new_n5307_), .B(_abc_41356_new_n4859_), .Y(_abc_41356_new_n6342_));
AND2X2 AND2X2_3027 ( .A(_abc_41356_new_n5875_), .B(sp_13_), .Y(_abc_41356_new_n6343_));
AND2X2 AND2X2_3028 ( .A(_abc_41356_new_n1286_), .B(regfil_4__5_), .Y(_abc_41356_new_n6344_));
AND2X2 AND2X2_3029 ( .A(_abc_41356_new_n6349_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6350_));
AND2X2 AND2X2_303 ( .A(_abc_41356_new_n526_), .B(regfil_3__6_), .Y(_abc_41356_new_n1064_));
AND2X2 AND2X2_3030 ( .A(_abc_41356_new_n6348_), .B(_abc_41356_new_n6350_), .Y(_abc_41356_new_n6351_));
AND2X2 AND2X2_3031 ( .A(_abc_41356_new_n6351_), .B(_abc_41356_new_n6337_), .Y(_abc_41356_new_n6352_));
AND2X2 AND2X2_3032 ( .A(_abc_41356_new_n6340_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6353_));
AND2X2 AND2X2_3033 ( .A(_abc_41356_new_n5307_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6354_));
AND2X2 AND2X2_3034 ( .A(_abc_41356_new_n5843_), .B(rdatahold_5_), .Y(_abc_41356_new_n6355_));
AND2X2 AND2X2_3035 ( .A(_abc_41356_new_n6358_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6359_));
AND2X2 AND2X2_3036 ( .A(_abc_41356_new_n5847_), .B(sp_14_), .Y(_abc_41356_new_n6361_));
AND2X2 AND2X2_3037 ( .A(_abc_41356_new_n6323_), .B(sp_14_), .Y(_abc_41356_new_n6362_));
AND2X2 AND2X2_3038 ( .A(_abc_41356_new_n6362_), .B(sp_0_), .Y(_abc_41356_new_n6363_));
AND2X2 AND2X2_3039 ( .A(_abc_41356_new_n6365_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6366_));
AND2X2 AND2X2_304 ( .A(_abc_41356_new_n623_), .B(regfil_2__6_), .Y(_abc_41356_new_n1065_));
AND2X2 AND2X2_3040 ( .A(_abc_41356_new_n6366_), .B(_abc_41356_new_n6364_), .Y(_abc_41356_new_n6367_));
AND2X2 AND2X2_3041 ( .A(_abc_41356_new_n5341_), .B(_abc_41356_new_n5883_), .Y(_abc_41356_new_n6368_));
AND2X2 AND2X2_3042 ( .A(_abc_41356_new_n6369_), .B(sp_14_), .Y(_abc_41356_new_n6370_));
AND2X2 AND2X2_3043 ( .A(_abc_41356_new_n6371_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6372_));
AND2X2 AND2X2_3044 ( .A(_abc_41356_new_n5855_), .B(sp_14_), .Y(_abc_41356_new_n6373_));
AND2X2 AND2X2_3045 ( .A(_abc_41356_new_n6377_), .B(_abc_41356_new_n6378_), .Y(_abc_41356_new_n6379_));
AND2X2 AND2X2_3046 ( .A(_abc_41356_new_n6379_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6380_));
AND2X2 AND2X2_3047 ( .A(_abc_41356_new_n5344_), .B(_abc_41356_new_n4859_), .Y(_abc_41356_new_n6381_));
AND2X2 AND2X2_3048 ( .A(_abc_41356_new_n5875_), .B(sp_14_), .Y(_abc_41356_new_n6382_));
AND2X2 AND2X2_3049 ( .A(_abc_41356_new_n1286_), .B(regfil_4__6_), .Y(_abc_41356_new_n6383_));
AND2X2 AND2X2_305 ( .A(_abc_41356_new_n1060_), .B(_abc_41356_new_n1068_), .Y(_abc_41356_new_n1069_));
AND2X2 AND2X2_3050 ( .A(_abc_41356_new_n6388_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6389_));
AND2X2 AND2X2_3051 ( .A(_abc_41356_new_n6387_), .B(_abc_41356_new_n6389_), .Y(_abc_41356_new_n6390_));
AND2X2 AND2X2_3052 ( .A(_abc_41356_new_n6390_), .B(_abc_41356_new_n6376_), .Y(_abc_41356_new_n6391_));
AND2X2 AND2X2_3053 ( .A(_abc_41356_new_n6379_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6392_));
AND2X2 AND2X2_3054 ( .A(_abc_41356_new_n5344_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6393_));
AND2X2 AND2X2_3055 ( .A(_abc_41356_new_n5843_), .B(rdatahold_6_), .Y(_abc_41356_new_n6394_));
AND2X2 AND2X2_3056 ( .A(_abc_41356_new_n6397_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6398_));
AND2X2 AND2X2_3057 ( .A(_abc_41356_new_n5847_), .B(sp_15_), .Y(_abc_41356_new_n6400_));
AND2X2 AND2X2_3058 ( .A(_abc_41356_new_n6364_), .B(sp_15_), .Y(_abc_41356_new_n6401_));
AND2X2 AND2X2_3059 ( .A(_abc_41356_new_n6363_), .B(_abc_41356_new_n1967_), .Y(_abc_41356_new_n6402_));
AND2X2 AND2X2_306 ( .A(_abc_41356_new_n1069_), .B(_abc_41356_new_n614_), .Y(_abc_41356_new_n1070_));
AND2X2 AND2X2_3060 ( .A(_abc_41356_new_n6403_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6404_));
AND2X2 AND2X2_3061 ( .A(_abc_41356_new_n6406_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6407_));
AND2X2 AND2X2_3062 ( .A(_abc_41356_new_n6407_), .B(_abc_41356_new_n6405_), .Y(_abc_41356_new_n6408_));
AND2X2 AND2X2_3063 ( .A(_abc_41356_new_n5855_), .B(sp_15_), .Y(_abc_41356_new_n6409_));
AND2X2 AND2X2_3064 ( .A(_abc_41356_new_n6377_), .B(sp_15_), .Y(_abc_41356_new_n6413_));
AND2X2 AND2X2_3065 ( .A(_abc_41356_new_n6362_), .B(_abc_41356_new_n1967_), .Y(_abc_41356_new_n6414_));
AND2X2 AND2X2_3066 ( .A(_abc_41356_new_n6415_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n6416_));
AND2X2 AND2X2_3067 ( .A(_abc_41356_new_n5381_), .B(_abc_41356_new_n4859_), .Y(_abc_41356_new_n6417_));
AND2X2 AND2X2_3068 ( .A(_abc_41356_new_n5875_), .B(sp_15_), .Y(_abc_41356_new_n6418_));
AND2X2 AND2X2_3069 ( .A(_abc_41356_new_n1286_), .B(regfil_4__7_), .Y(_abc_41356_new_n6419_));
AND2X2 AND2X2_307 ( .A(_abc_41356_new_n612_), .B(alu_res_6_), .Y(_abc_41356_new_n1071_));
AND2X2 AND2X2_3070 ( .A(_abc_41356_new_n6424_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6425_));
AND2X2 AND2X2_3071 ( .A(_abc_41356_new_n6423_), .B(_abc_41356_new_n6425_), .Y(_abc_41356_new_n6426_));
AND2X2 AND2X2_3072 ( .A(_abc_41356_new_n6412_), .B(_abc_41356_new_n6426_), .Y(_abc_41356_new_n6427_));
AND2X2 AND2X2_3073 ( .A(_abc_41356_new_n6415_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n6428_));
AND2X2 AND2X2_3074 ( .A(_abc_41356_new_n5381_), .B(_abc_41356_new_n5838_), .Y(_abc_41356_new_n6429_));
AND2X2 AND2X2_3075 ( .A(_abc_41356_new_n5843_), .B(rdatahold_7_), .Y(_abc_41356_new_n6430_));
AND2X2 AND2X2_3076 ( .A(_abc_41356_new_n6433_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n6434_));
AND2X2 AND2X2_3077 ( .A(_abc_41356_new_n1211_), .B(_abc_41356_new_n2549_), .Y(_abc_41356_new_n6436_));
AND2X2 AND2X2_3078 ( .A(_abc_41356_new_n6439_), .B(_abc_41356_new_n6437_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_0_));
AND2X2 AND2X2_3079 ( .A(_abc_41356_new_n6442_), .B(_abc_41356_new_n6441_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_1_));
AND2X2 AND2X2_308 ( .A(_abc_41356_new_n608_), .B(rdatahold_6_), .Y(_abc_41356_new_n1072_));
AND2X2 AND2X2_3080 ( .A(_abc_41356_new_n6445_), .B(_abc_41356_new_n6444_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_2_));
AND2X2 AND2X2_3081 ( .A(_abc_41356_new_n6448_), .B(_abc_41356_new_n6447_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_3_));
AND2X2 AND2X2_3082 ( .A(_abc_41356_new_n6451_), .B(_abc_41356_new_n6450_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_4_));
AND2X2 AND2X2_3083 ( .A(_abc_41356_new_n6454_), .B(_abc_41356_new_n6453_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_5_));
AND2X2 AND2X2_3084 ( .A(_abc_41356_new_n6457_), .B(_abc_41356_new_n6456_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_6_));
AND2X2 AND2X2_3085 ( .A(_abc_41356_new_n6460_), .B(_abc_41356_new_n6459_), .Y(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_7_));
AND2X2 AND2X2_3086 ( .A(_abc_41356_new_n6463_), .B(_abc_41356_new_n3723_), .Y(_abc_41356_new_n6464_));
AND2X2 AND2X2_3087 ( .A(_abc_41356_new_n6462_), .B(pc_0_), .Y(_abc_41356_new_n6465_));
AND2X2 AND2X2_3088 ( .A(_abc_41356_new_n6466_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n6467_));
AND2X2 AND2X2_3089 ( .A(_abc_41356_new_n2023_), .B(_abc_41356_new_n3723_), .Y(_abc_41356_new_n6468_));
AND2X2 AND2X2_309 ( .A(_abc_41356_new_n1074_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n1075_));
AND2X2 AND2X2_3090 ( .A(_abc_41356_new_n6469_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6470_));
AND2X2 AND2X2_3091 ( .A(_abc_41356_new_n1237_), .B(_abc_41356_new_n3711_), .Y(_abc_41356_new_n6471_));
AND2X2 AND2X2_3092 ( .A(_abc_41356_new_n599_), .B(_abc_41356_new_n534_), .Y(_abc_41356_new_n6472_));
AND2X2 AND2X2_3093 ( .A(_abc_41356_new_n6473_), .B(_abc_41356_new_n2047_), .Y(_abc_41356_new_n6474_));
AND2X2 AND2X2_3094 ( .A(_abc_41356_new_n6477_), .B(_abc_41356_new_n4166_), .Y(_abc_41356_new_n6478_));
AND2X2 AND2X2_3095 ( .A(_abc_41356_new_n2047_), .B(_abc_41356_new_n681_), .Y(_abc_41356_new_n6479_));
AND2X2 AND2X2_3096 ( .A(_abc_41356_new_n5874_), .B(_abc_41356_new_n5882_), .Y(_abc_41356_new_n6483_));
AND2X2 AND2X2_3097 ( .A(_abc_41356_new_n6482_), .B(_abc_41356_new_n6483_), .Y(_abc_41356_new_n6484_));
AND2X2 AND2X2_3098 ( .A(_abc_41356_new_n6478_), .B(_abc_41356_new_n6484_), .Y(_abc_41356_new_n6485_));
AND2X2 AND2X2_3099 ( .A(_abc_41356_new_n6485_), .B(_abc_41356_new_n4155_), .Y(_abc_41356_new_n6486_));
AND2X2 AND2X2_31 ( .A(_abc_41356_new_n549_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n550_));
AND2X2 AND2X2_310 ( .A(_abc_41356_new_n992_), .B(_abc_41356_new_n1076_), .Y(_abc_41356_new_n1077_));
AND2X2 AND2X2_3100 ( .A(_abc_41356_new_n2054_), .B(_abc_41356_new_n6488_), .Y(_abc_41356_new_n6489_));
AND2X2 AND2X2_3101 ( .A(_abc_41356_new_n6494_), .B(_abc_41356_new_n6489_), .Y(_abc_41356_new_n6495_));
AND2X2 AND2X2_3102 ( .A(_abc_41356_new_n6495_), .B(_abc_41356_new_n3494_), .Y(_abc_41356_new_n6496_));
AND2X2 AND2X2_3103 ( .A(_abc_41356_new_n2061_), .B(_abc_41356_new_n6496_), .Y(_abc_41356_new_n6497_));
AND2X2 AND2X2_3104 ( .A(_abc_41356_new_n6486_), .B(_abc_41356_new_n6497_), .Y(_abc_41356_new_n6498_));
AND2X2 AND2X2_3105 ( .A(_abc_41356_new_n6499_), .B(_abc_41356_new_n6492_), .Y(_abc_41356_new_n6500_));
AND2X2 AND2X2_3106 ( .A(_abc_41356_new_n6501_), .B(_abc_41356_new_n6089_), .Y(_abc_41356_new_n6502_));
AND2X2 AND2X2_3107 ( .A(_abc_41356_new_n606_), .B(_abc_41356_new_n518_), .Y(_abc_41356_new_n6503_));
AND2X2 AND2X2_3108 ( .A(_abc_41356_new_n6505_), .B(_abc_41356_new_n3265_), .Y(_abc_41356_new_n6506_));
AND2X2 AND2X2_3109 ( .A(_abc_41356_new_n6506_), .B(pc_0_), .Y(_abc_41356_new_n6507_));
AND2X2 AND2X2_311 ( .A(_abc_41356_new_n991_), .B(regfil_0__6_), .Y(_abc_41356_new_n1078_));
AND2X2 AND2X2_3110 ( .A(_abc_41356_new_n6504_), .B(rdatahold2_0_), .Y(_abc_41356_new_n6508_));
AND2X2 AND2X2_3111 ( .A(_abc_41356_new_n6511_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__0_));
AND2X2 AND2X2_3112 ( .A(_abc_41356_new_n1237_), .B(_abc_41356_new_n6513_), .Y(_abc_41356_new_n6514_));
AND2X2 AND2X2_3113 ( .A(_abc_41356_new_n2376_), .B(_abc_41356_new_n534_), .Y(_abc_41356_new_n6515_));
AND2X2 AND2X2_3114 ( .A(_abc_41356_new_n4154_), .B(_abc_41356_new_n6519_), .Y(_abc_41356_new_n6520_));
AND2X2 AND2X2_3115 ( .A(_abc_41356_new_n6520_), .B(_abc_41356_new_n6518_), .Y(_abc_41356_new_n6521_));
AND2X2 AND2X2_3116 ( .A(_abc_41356_new_n6530_), .B(_abc_41356_new_n6521_), .Y(_abc_41356_new_n6531_));
AND2X2 AND2X2_3117 ( .A(_abc_41356_new_n6532_), .B(_abc_41356_new_n6533_), .Y(_abc_41356_new_n6534_));
AND2X2 AND2X2_3118 ( .A(_abc_41356_new_n6534_), .B(_abc_41356_new_n5849_), .Y(_abc_41356_new_n6535_));
AND2X2 AND2X2_3119 ( .A(_abc_41356_new_n6535_), .B(_abc_41356_new_n3358_), .Y(_abc_41356_new_n6536_));
AND2X2 AND2X2_312 ( .A(_abc_41356_new_n1079_), .B(_abc_41356_new_n602_), .Y(_abc_41356_new_n1080_));
AND2X2 AND2X2_3120 ( .A(_abc_41356_new_n6531_), .B(_abc_41356_new_n6536_), .Y(_abc_41356_new_n6537_));
AND2X2 AND2X2_3121 ( .A(_abc_41356_new_n6538_), .B(_abc_41356_new_n3762_), .Y(_abc_41356_new_n6539_));
AND2X2 AND2X2_3122 ( .A(_abc_41356_new_n4124_), .B(_abc_41356_new_n3764_), .Y(_abc_41356_new_n6540_));
AND2X2 AND2X2_3123 ( .A(_abc_41356_new_n677_), .B(_abc_41356_new_n3817_), .Y(_abc_41356_new_n6541_));
AND2X2 AND2X2_3124 ( .A(_abc_41356_new_n6545_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n6546_));
AND2X2 AND2X2_3125 ( .A(_abc_41356_new_n6544_), .B(_abc_41356_new_n6546_), .Y(_abc_41356_new_n6547_));
AND2X2 AND2X2_3126 ( .A(_abc_41356_new_n2023_), .B(_abc_41356_new_n3762_), .Y(_abc_41356_new_n6548_));
AND2X2 AND2X2_3127 ( .A(_abc_41356_new_n6498_), .B(pc_1_), .Y(_abc_41356_new_n6549_));
AND2X2 AND2X2_3128 ( .A(_abc_41356_new_n6487_), .B(_abc_41356_new_n3762_), .Y(_abc_41356_new_n6550_));
AND2X2 AND2X2_3129 ( .A(_abc_41356_new_n3495_), .B(_abc_41356_new_n3817_), .Y(_abc_41356_new_n6551_));
AND2X2 AND2X2_313 ( .A(_abc_41356_new_n985_), .B(regfil_0__6_), .Y(_abc_41356_new_n1085_));
AND2X2 AND2X2_3130 ( .A(_abc_41356_new_n1417_), .B(regfil_5__1_), .Y(_abc_41356_new_n6552_));
AND2X2 AND2X2_3131 ( .A(_abc_41356_new_n6490_), .B(_abc_41356_new_n3764_), .Y(_abc_41356_new_n6553_));
AND2X2 AND2X2_3132 ( .A(_abc_41356_new_n6557_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n6558_));
AND2X2 AND2X2_3133 ( .A(_abc_41356_new_n6560_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6561_));
AND2X2 AND2X2_3134 ( .A(_abc_41356_new_n6506_), .B(pc_1_), .Y(_abc_41356_new_n6562_));
AND2X2 AND2X2_3135 ( .A(_abc_41356_new_n6504_), .B(rdatahold2_1_), .Y(_abc_41356_new_n6563_));
AND2X2 AND2X2_3136 ( .A(_abc_41356_new_n6565_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__1_));
AND2X2 AND2X2_3137 ( .A(_abc_41356_new_n6570_), .B(_abc_41356_new_n4149_), .Y(_abc_41356_new_n6571_));
AND2X2 AND2X2_3138 ( .A(_abc_41356_new_n6568_), .B(_abc_41356_new_n6571_), .Y(_abc_41356_new_n6572_));
AND2X2 AND2X2_3139 ( .A(_abc_41356_new_n6567_), .B(_abc_41356_new_n6572_), .Y(_abc_41356_new_n6573_));
AND2X2 AND2X2_314 ( .A(_abc_41356_new_n1087_), .B(_abc_41356_new_n1082_), .Y(_abc_41356_new_n1088_));
AND2X2 AND2X2_3140 ( .A(_abc_41356_new_n4148_), .B(_abc_41356_new_n3811_), .Y(_abc_41356_new_n6574_));
AND2X2 AND2X2_3141 ( .A(_abc_41356_new_n6498_), .B(pc_2_), .Y(_abc_41356_new_n6577_));
AND2X2 AND2X2_3142 ( .A(_abc_41356_new_n6582_), .B(_abc_41356_new_n6581_), .Y(_abc_41356_new_n6583_));
AND2X2 AND2X2_3143 ( .A(_abc_41356_new_n6583_), .B(_abc_41356_new_n6580_), .Y(_abc_41356_new_n6584_));
AND2X2 AND2X2_3144 ( .A(_abc_41356_new_n6579_), .B(_abc_41356_new_n6584_), .Y(_abc_41356_new_n6585_));
AND2X2 AND2X2_3145 ( .A(_abc_41356_new_n6578_), .B(_abc_41356_new_n6585_), .Y(_abc_41356_new_n6586_));
AND2X2 AND2X2_3146 ( .A(_abc_41356_new_n6587_), .B(_abc_41356_new_n6588_), .Y(_abc_41356_new_n6589_));
AND2X2 AND2X2_3147 ( .A(_abc_41356_new_n6589_), .B(_abc_41356_new_n6576_), .Y(_abc_41356_new_n6590_));
AND2X2 AND2X2_3148 ( .A(_abc_41356_new_n6591_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6592_));
AND2X2 AND2X2_3149 ( .A(_abc_41356_new_n6506_), .B(pc_2_), .Y(_abc_41356_new_n6593_));
AND2X2 AND2X2_315 ( .A(_abc_41356_new_n1088_), .B(_abc_41356_new_n1081_), .Y(_abc_41356_new_n1089_));
AND2X2 AND2X2_3150 ( .A(_abc_41356_new_n6504_), .B(rdatahold2_2_), .Y(_abc_41356_new_n6594_));
AND2X2 AND2X2_3151 ( .A(_abc_41356_new_n6596_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__2_));
AND2X2 AND2X2_3152 ( .A(_abc_41356_new_n6603_), .B(_abc_41356_new_n6602_), .Y(_abc_41356_new_n6604_));
AND2X2 AND2X2_3153 ( .A(_abc_41356_new_n6606_), .B(_abc_41356_new_n4149_), .Y(_abc_41356_new_n6607_));
AND2X2 AND2X2_3154 ( .A(_abc_41356_new_n6601_), .B(_abc_41356_new_n6607_), .Y(_abc_41356_new_n6608_));
AND2X2 AND2X2_3155 ( .A(_abc_41356_new_n6599_), .B(_abc_41356_new_n6608_), .Y(_abc_41356_new_n6609_));
AND2X2 AND2X2_3156 ( .A(_abc_41356_new_n4148_), .B(_abc_41356_new_n6602_), .Y(_abc_41356_new_n6610_));
AND2X2 AND2X2_3157 ( .A(_abc_41356_new_n6498_), .B(pc_3_), .Y(_abc_41356_new_n6613_));
AND2X2 AND2X2_3158 ( .A(_abc_41356_new_n6490_), .B(_abc_41356_new_n3883_), .Y(_abc_41356_new_n6616_));
AND2X2 AND2X2_3159 ( .A(_abc_41356_new_n1417_), .B(regfil_5__3_), .Y(_abc_41356_new_n6620_));
AND2X2 AND2X2_316 ( .A(_abc_41356_new_n1092_), .B(_abc_41356_new_n695_), .Y(_abc_41356_new_n1093_));
AND2X2 AND2X2_3160 ( .A(_abc_41356_new_n6621_), .B(_abc_41356_new_n6619_), .Y(_abc_41356_new_n6622_));
AND2X2 AND2X2_3161 ( .A(_abc_41356_new_n6622_), .B(_abc_41356_new_n6618_), .Y(_abc_41356_new_n6623_));
AND2X2 AND2X2_3162 ( .A(_abc_41356_new_n6623_), .B(_abc_41356_new_n6617_), .Y(_abc_41356_new_n6624_));
AND2X2 AND2X2_3163 ( .A(_abc_41356_new_n6615_), .B(_abc_41356_new_n6624_), .Y(_abc_41356_new_n6625_));
AND2X2 AND2X2_3164 ( .A(_abc_41356_new_n6614_), .B(_abc_41356_new_n6625_), .Y(_abc_41356_new_n6626_));
AND2X2 AND2X2_3165 ( .A(_abc_41356_new_n3879_), .B(_abc_41356_new_n2023_), .Y(_abc_41356_new_n6628_));
AND2X2 AND2X2_3166 ( .A(_abc_41356_new_n6627_), .B(_abc_41356_new_n6629_), .Y(_abc_41356_new_n6630_));
AND2X2 AND2X2_3167 ( .A(_abc_41356_new_n6630_), .B(_abc_41356_new_n6612_), .Y(_abc_41356_new_n6631_));
AND2X2 AND2X2_3168 ( .A(_abc_41356_new_n6632_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6633_));
AND2X2 AND2X2_3169 ( .A(_abc_41356_new_n6506_), .B(pc_3_), .Y(_abc_41356_new_n6634_));
AND2X2 AND2X2_317 ( .A(_abc_41356_new_n696_), .B(_abc_41356_new_n700_), .Y(_abc_41356_new_n1094_));
AND2X2 AND2X2_3170 ( .A(_abc_41356_new_n6504_), .B(rdatahold2_3_), .Y(_abc_41356_new_n6635_));
AND2X2 AND2X2_3171 ( .A(_abc_41356_new_n6637_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__3_));
AND2X2 AND2X2_3172 ( .A(_abc_41356_new_n6538_), .B(_abc_41356_new_n3929_), .Y(_abc_41356_new_n6639_));
AND2X2 AND2X2_3173 ( .A(_abc_41356_new_n4124_), .B(_abc_41356_new_n3934_), .Y(_abc_41356_new_n6640_));
AND2X2 AND2X2_3174 ( .A(_abc_41356_new_n2071_), .B(pc_4_), .Y(_abc_41356_new_n6641_));
AND2X2 AND2X2_3175 ( .A(_abc_41356_new_n6642_), .B(_abc_41356_new_n6643_), .Y(_abc_41356_new_n6644_));
AND2X2 AND2X2_3176 ( .A(_abc_41356_new_n6644_), .B(_abc_41356_new_n677_), .Y(_abc_41356_new_n6645_));
AND2X2 AND2X2_3177 ( .A(_abc_41356_new_n6649_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n6650_));
AND2X2 AND2X2_3178 ( .A(_abc_41356_new_n6648_), .B(_abc_41356_new_n6650_), .Y(_abc_41356_new_n6651_));
AND2X2 AND2X2_3179 ( .A(_abc_41356_new_n3929_), .B(_abc_41356_new_n2023_), .Y(_abc_41356_new_n6652_));
AND2X2 AND2X2_318 ( .A(_abc_41356_new_n512_), .B(_abc_41356_new_n1097_), .Y(_abc_41356_new_n1098_));
AND2X2 AND2X2_3180 ( .A(_abc_41356_new_n6653_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6654_));
AND2X2 AND2X2_3181 ( .A(_abc_41356_new_n6498_), .B(pc_4_), .Y(_abc_41356_new_n6655_));
AND2X2 AND2X2_3182 ( .A(_abc_41356_new_n6487_), .B(_abc_41356_new_n3929_), .Y(_abc_41356_new_n6656_));
AND2X2 AND2X2_3183 ( .A(_abc_41356_new_n2059_), .B(opcode_4_), .Y(_abc_41356_new_n6657_));
AND2X2 AND2X2_3184 ( .A(_abc_41356_new_n3934_), .B(_abc_41356_new_n6490_), .Y(_abc_41356_new_n6658_));
AND2X2 AND2X2_3185 ( .A(_abc_41356_new_n3495_), .B(_abc_41356_new_n6644_), .Y(_abc_41356_new_n6659_));
AND2X2 AND2X2_3186 ( .A(_abc_41356_new_n1417_), .B(regfil_5__4_), .Y(_abc_41356_new_n6660_));
AND2X2 AND2X2_3187 ( .A(_abc_41356_new_n6665_), .B(_abc_41356_new_n6089_), .Y(_abc_41356_new_n6666_));
AND2X2 AND2X2_3188 ( .A(_abc_41356_new_n6506_), .B(pc_4_), .Y(_abc_41356_new_n6667_));
AND2X2 AND2X2_3189 ( .A(_abc_41356_new_n6504_), .B(rdatahold2_4_), .Y(_abc_41356_new_n6668_));
AND2X2 AND2X2_319 ( .A(_abc_41356_new_n551_), .B(_abc_41356_new_n700_), .Y(_abc_41356_new_n1100_));
AND2X2 AND2X2_3190 ( .A(_abc_41356_new_n6671_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__4_));
AND2X2 AND2X2_3191 ( .A(_abc_41356_new_n2071_), .B(_abc_41356_new_n2036_), .Y(_abc_41356_new_n6675_));
AND2X2 AND2X2_3192 ( .A(_abc_41356_new_n6642_), .B(_abc_41356_new_n3980_), .Y(_abc_41356_new_n6676_));
AND2X2 AND2X2_3193 ( .A(_abc_41356_new_n6678_), .B(_abc_41356_new_n4149_), .Y(_abc_41356_new_n6679_));
AND2X2 AND2X2_3194 ( .A(_abc_41356_new_n6674_), .B(_abc_41356_new_n6679_), .Y(_abc_41356_new_n6680_));
AND2X2 AND2X2_3195 ( .A(_abc_41356_new_n6673_), .B(_abc_41356_new_n6680_), .Y(_abc_41356_new_n6681_));
AND2X2 AND2X2_3196 ( .A(_abc_41356_new_n4148_), .B(_abc_41356_new_n3980_), .Y(_abc_41356_new_n6682_));
AND2X2 AND2X2_3197 ( .A(_abc_41356_new_n6498_), .B(pc_5_), .Y(_abc_41356_new_n6685_));
AND2X2 AND2X2_3198 ( .A(_abc_41356_new_n3988_), .B(_abc_41356_new_n6490_), .Y(_abc_41356_new_n6688_));
AND2X2 AND2X2_3199 ( .A(_abc_41356_new_n1417_), .B(regfil_5__5_), .Y(_abc_41356_new_n6691_));
AND2X2 AND2X2_32 ( .A(_abc_41356_new_n550_), .B(_abc_41356_new_n544_), .Y(_abc_41356_new_n551_));
AND2X2 AND2X2_320 ( .A(_abc_41356_new_n1101_), .B(_abc_41356_new_n701_), .Y(_abc_41356_new_n1102_));
AND2X2 AND2X2_3200 ( .A(_abc_41356_new_n6693_), .B(_abc_41356_new_n6692_), .Y(_abc_41356_new_n6694_));
AND2X2 AND2X2_3201 ( .A(_abc_41356_new_n6690_), .B(_abc_41356_new_n6694_), .Y(_abc_41356_new_n6695_));
AND2X2 AND2X2_3202 ( .A(_abc_41356_new_n6695_), .B(_abc_41356_new_n6689_), .Y(_abc_41356_new_n6696_));
AND2X2 AND2X2_3203 ( .A(_abc_41356_new_n6687_), .B(_abc_41356_new_n6696_), .Y(_abc_41356_new_n6697_));
AND2X2 AND2X2_3204 ( .A(_abc_41356_new_n6686_), .B(_abc_41356_new_n6697_), .Y(_abc_41356_new_n6698_));
AND2X2 AND2X2_3205 ( .A(_abc_41356_new_n3983_), .B(_abc_41356_new_n2023_), .Y(_abc_41356_new_n6700_));
AND2X2 AND2X2_3206 ( .A(_abc_41356_new_n6699_), .B(_abc_41356_new_n6701_), .Y(_abc_41356_new_n6702_));
AND2X2 AND2X2_3207 ( .A(_abc_41356_new_n6702_), .B(_abc_41356_new_n6684_), .Y(_abc_41356_new_n6703_));
AND2X2 AND2X2_3208 ( .A(_abc_41356_new_n6704_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6705_));
AND2X2 AND2X2_3209 ( .A(_abc_41356_new_n6506_), .B(pc_5_), .Y(_abc_41356_new_n6706_));
AND2X2 AND2X2_321 ( .A(_abc_41356_new_n537_), .B(_abc_41356_new_n700_), .Y(_abc_41356_new_n1104_));
AND2X2 AND2X2_3210 ( .A(_abc_41356_new_n6504_), .B(rdatahold2_5_), .Y(_abc_41356_new_n6707_));
AND2X2 AND2X2_3211 ( .A(_abc_41356_new_n6709_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__5_));
AND2X2 AND2X2_3212 ( .A(_abc_41356_new_n6675_), .B(pc_6_), .Y(_abc_41356_new_n6715_));
AND2X2 AND2X2_3213 ( .A(_abc_41356_new_n6717_), .B(_abc_41356_new_n6716_), .Y(_abc_41356_new_n6718_));
AND2X2 AND2X2_3214 ( .A(_abc_41356_new_n6720_), .B(_abc_41356_new_n4149_), .Y(_abc_41356_new_n6721_));
AND2X2 AND2X2_3215 ( .A(_abc_41356_new_n6714_), .B(_abc_41356_new_n6721_), .Y(_abc_41356_new_n6722_));
AND2X2 AND2X2_3216 ( .A(_abc_41356_new_n6712_), .B(_abc_41356_new_n6722_), .Y(_abc_41356_new_n6723_));
AND2X2 AND2X2_3217 ( .A(_abc_41356_new_n4148_), .B(_abc_41356_new_n6716_), .Y(_abc_41356_new_n6724_));
AND2X2 AND2X2_3218 ( .A(_abc_41356_new_n6498_), .B(pc_6_), .Y(_abc_41356_new_n6727_));
AND2X2 AND2X2_3219 ( .A(_abc_41356_new_n6732_), .B(_abc_41356_new_n6731_), .Y(_abc_41356_new_n6733_));
AND2X2 AND2X2_322 ( .A(regfil_7__6_), .B(regfil_7__5_), .Y(_abc_41356_new_n1106_));
AND2X2 AND2X2_3220 ( .A(_abc_41356_new_n6730_), .B(_abc_41356_new_n6733_), .Y(_abc_41356_new_n6734_));
AND2X2 AND2X2_3221 ( .A(_abc_41356_new_n6729_), .B(_abc_41356_new_n6734_), .Y(_abc_41356_new_n6735_));
AND2X2 AND2X2_3222 ( .A(_abc_41356_new_n6728_), .B(_abc_41356_new_n6735_), .Y(_abc_41356_new_n6736_));
AND2X2 AND2X2_3223 ( .A(_abc_41356_new_n6737_), .B(_abc_41356_new_n6738_), .Y(_abc_41356_new_n6739_));
AND2X2 AND2X2_3224 ( .A(_abc_41356_new_n6739_), .B(_abc_41356_new_n6726_), .Y(_abc_41356_new_n6740_));
AND2X2 AND2X2_3225 ( .A(_abc_41356_new_n6741_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6742_));
AND2X2 AND2X2_3226 ( .A(_abc_41356_new_n6506_), .B(pc_6_), .Y(_abc_41356_new_n6743_));
AND2X2 AND2X2_3227 ( .A(_abc_41356_new_n6504_), .B(rdatahold2_6_), .Y(_abc_41356_new_n6744_));
AND2X2 AND2X2_3228 ( .A(_abc_41356_new_n6746_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__6_));
AND2X2 AND2X2_3229 ( .A(_abc_41356_new_n4070_), .B(_abc_41356_new_n4124_), .Y(_abc_41356_new_n6749_));
AND2X2 AND2X2_323 ( .A(_abc_41356_new_n1033_), .B(_abc_41356_new_n1106_), .Y(_abc_41356_new_n1107_));
AND2X2 AND2X2_3230 ( .A(_abc_41356_new_n6675_), .B(_abc_41356_new_n2037_), .Y(_abc_41356_new_n6751_));
AND2X2 AND2X2_3231 ( .A(_abc_41356_new_n6753_), .B(_abc_41356_new_n6752_), .Y(_abc_41356_new_n6754_));
AND2X2 AND2X2_3232 ( .A(_abc_41356_new_n6754_), .B(_abc_41356_new_n677_), .Y(_abc_41356_new_n6755_));
AND2X2 AND2X2_3233 ( .A(_abc_41356_new_n6756_), .B(_abc_41356_new_n4149_), .Y(_abc_41356_new_n6757_));
AND2X2 AND2X2_3234 ( .A(_abc_41356_new_n6750_), .B(_abc_41356_new_n6757_), .Y(_abc_41356_new_n6758_));
AND2X2 AND2X2_3235 ( .A(_abc_41356_new_n6748_), .B(_abc_41356_new_n6758_), .Y(_abc_41356_new_n6759_));
AND2X2 AND2X2_3236 ( .A(_abc_41356_new_n4148_), .B(_abc_41356_new_n4072_), .Y(_abc_41356_new_n6760_));
AND2X2 AND2X2_3237 ( .A(_abc_41356_new_n6498_), .B(pc_7_), .Y(_abc_41356_new_n6763_));
AND2X2 AND2X2_3238 ( .A(_abc_41356_new_n4070_), .B(_abc_41356_new_n6490_), .Y(_abc_41356_new_n6765_));
AND2X2 AND2X2_3239 ( .A(_abc_41356_new_n1417_), .B(regfil_5__7_), .Y(_abc_41356_new_n6768_));
AND2X2 AND2X2_324 ( .A(_abc_41356_new_n551_), .B(_abc_41356_new_n1108_), .Y(_abc_41356_new_n1109_));
AND2X2 AND2X2_3240 ( .A(_abc_41356_new_n6754_), .B(_abc_41356_new_n3495_), .Y(_abc_41356_new_n6770_));
AND2X2 AND2X2_3241 ( .A(_abc_41356_new_n6771_), .B(_abc_41356_new_n6769_), .Y(_abc_41356_new_n6772_));
AND2X2 AND2X2_3242 ( .A(_abc_41356_new_n6767_), .B(_abc_41356_new_n6772_), .Y(_abc_41356_new_n6773_));
AND2X2 AND2X2_3243 ( .A(_abc_41356_new_n6773_), .B(_abc_41356_new_n6766_), .Y(_abc_41356_new_n6774_));
AND2X2 AND2X2_3244 ( .A(_abc_41356_new_n6774_), .B(_abc_41356_new_n6764_), .Y(_abc_41356_new_n6775_));
AND2X2 AND2X2_3245 ( .A(_abc_41356_new_n4075_), .B(_abc_41356_new_n2023_), .Y(_abc_41356_new_n6777_));
AND2X2 AND2X2_3246 ( .A(_abc_41356_new_n6776_), .B(_abc_41356_new_n6778_), .Y(_abc_41356_new_n6779_));
AND2X2 AND2X2_3247 ( .A(_abc_41356_new_n6779_), .B(_abc_41356_new_n6762_), .Y(_abc_41356_new_n6780_));
AND2X2 AND2X2_3248 ( .A(_abc_41356_new_n6781_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6782_));
AND2X2 AND2X2_3249 ( .A(_abc_41356_new_n6506_), .B(pc_7_), .Y(_abc_41356_new_n6783_));
AND2X2 AND2X2_325 ( .A(_abc_41356_new_n1110_), .B(_abc_41356_new_n1105_), .Y(_abc_41356_new_n1111_));
AND2X2 AND2X2_3250 ( .A(_abc_41356_new_n6504_), .B(rdatahold2_7_), .Y(_abc_41356_new_n6784_));
AND2X2 AND2X2_3251 ( .A(_abc_41356_new_n6786_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__7_));
AND2X2 AND2X2_3252 ( .A(_abc_41356_new_n6752_), .B(_abc_41356_new_n2041_), .Y(_abc_41356_new_n6790_));
AND2X2 AND2X2_3253 ( .A(_abc_41356_new_n6751_), .B(pc_8_), .Y(_abc_41356_new_n6791_));
AND2X2 AND2X2_3254 ( .A(_abc_41356_new_n6793_), .B(_abc_41356_new_n4149_), .Y(_abc_41356_new_n6794_));
AND2X2 AND2X2_3255 ( .A(_abc_41356_new_n6794_), .B(_abc_41356_new_n6789_), .Y(_abc_41356_new_n6795_));
AND2X2 AND2X2_3256 ( .A(_abc_41356_new_n6788_), .B(_abc_41356_new_n6795_), .Y(_abc_41356_new_n6796_));
AND2X2 AND2X2_3257 ( .A(_abc_41356_new_n4148_), .B(_abc_41356_new_n2041_), .Y(_abc_41356_new_n6797_));
AND2X2 AND2X2_3258 ( .A(_abc_41356_new_n6498_), .B(pc_8_), .Y(_abc_41356_new_n6800_));
AND2X2 AND2X2_3259 ( .A(_abc_41356_new_n6802_), .B(_abc_41356_new_n6803_), .Y(_abc_41356_new_n6804_));
AND2X2 AND2X2_326 ( .A(_abc_41356_new_n1035_), .B(_abc_41356_new_n700_), .Y(_abc_41356_new_n1112_));
AND2X2 AND2X2_3260 ( .A(_abc_41356_new_n1417_), .B(regfil_4__0_), .Y(_abc_41356_new_n6806_));
AND2X2 AND2X2_3261 ( .A(_abc_41356_new_n6805_), .B(_abc_41356_new_n6807_), .Y(_abc_41356_new_n6808_));
AND2X2 AND2X2_3262 ( .A(_abc_41356_new_n6808_), .B(_abc_41356_new_n6804_), .Y(_abc_41356_new_n6809_));
AND2X2 AND2X2_3263 ( .A(_abc_41356_new_n6809_), .B(_abc_41356_new_n6801_), .Y(_abc_41356_new_n6810_));
AND2X2 AND2X2_3264 ( .A(_abc_41356_new_n6811_), .B(_abc_41356_new_n6812_), .Y(_abc_41356_new_n6813_));
AND2X2 AND2X2_3265 ( .A(_abc_41356_new_n6813_), .B(_abc_41356_new_n6799_), .Y(_abc_41356_new_n6814_));
AND2X2 AND2X2_3266 ( .A(_abc_41356_new_n6815_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6816_));
AND2X2 AND2X2_3267 ( .A(_abc_41356_new_n6506_), .B(pc_8_), .Y(_abc_41356_new_n6817_));
AND2X2 AND2X2_3268 ( .A(_abc_41356_new_n6504_), .B(rdatahold_0_), .Y(_abc_41356_new_n6818_));
AND2X2 AND2X2_3269 ( .A(_abc_41356_new_n6820_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__8_));
AND2X2 AND2X2_327 ( .A(_abc_41356_new_n1113_), .B(_abc_41356_new_n1103_), .Y(_abc_41356_new_n1114_));
AND2X2 AND2X2_3270 ( .A(_abc_41356_new_n6791_), .B(pc_9_), .Y(_abc_41356_new_n6822_));
AND2X2 AND2X2_3271 ( .A(_abc_41356_new_n6824_), .B(_abc_41356_new_n6823_), .Y(_abc_41356_new_n6825_));
AND2X2 AND2X2_3272 ( .A(_abc_41356_new_n6827_), .B(_abc_41356_new_n4149_), .Y(_abc_41356_new_n6828_));
AND2X2 AND2X2_3273 ( .A(_abc_41356_new_n6832_), .B(_abc_41356_new_n6830_), .Y(_abc_41356_new_n6833_));
AND2X2 AND2X2_3274 ( .A(_abc_41356_new_n6833_), .B(_abc_41356_new_n6828_), .Y(_abc_41356_new_n6834_));
AND2X2 AND2X2_3275 ( .A(_abc_41356_new_n4148_), .B(_abc_41356_new_n6823_), .Y(_abc_41356_new_n6835_));
AND2X2 AND2X2_3276 ( .A(_abc_41356_new_n6498_), .B(pc_9_), .Y(_abc_41356_new_n6838_));
AND2X2 AND2X2_3277 ( .A(_abc_41356_new_n6840_), .B(_abc_41356_new_n6841_), .Y(_abc_41356_new_n6842_));
AND2X2 AND2X2_3278 ( .A(_abc_41356_new_n1417_), .B(regfil_4__1_), .Y(_abc_41356_new_n6844_));
AND2X2 AND2X2_3279 ( .A(_abc_41356_new_n6843_), .B(_abc_41356_new_n6845_), .Y(_abc_41356_new_n6846_));
AND2X2 AND2X2_328 ( .A(_abc_41356_new_n1115_), .B(_abc_41356_new_n1029_), .Y(_abc_41356_new_n1116_));
AND2X2 AND2X2_3280 ( .A(_abc_41356_new_n6846_), .B(_abc_41356_new_n6842_), .Y(_abc_41356_new_n6847_));
AND2X2 AND2X2_3281 ( .A(_abc_41356_new_n6847_), .B(_abc_41356_new_n6839_), .Y(_abc_41356_new_n6848_));
AND2X2 AND2X2_3282 ( .A(_abc_41356_new_n6849_), .B(_abc_41356_new_n6850_), .Y(_abc_41356_new_n6851_));
AND2X2 AND2X2_3283 ( .A(_abc_41356_new_n6837_), .B(_abc_41356_new_n6851_), .Y(_abc_41356_new_n6852_));
AND2X2 AND2X2_3284 ( .A(_abc_41356_new_n6853_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6854_));
AND2X2 AND2X2_3285 ( .A(_abc_41356_new_n6506_), .B(pc_9_), .Y(_abc_41356_new_n6855_));
AND2X2 AND2X2_3286 ( .A(_abc_41356_new_n6504_), .B(rdatahold_1_), .Y(_abc_41356_new_n6856_));
AND2X2 AND2X2_3287 ( .A(_abc_41356_new_n6858_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__9_));
AND2X2 AND2X2_3288 ( .A(_abc_41356_new_n6822_), .B(pc_10_), .Y(_abc_41356_new_n6860_));
AND2X2 AND2X2_3289 ( .A(_abc_41356_new_n6861_), .B(_abc_41356_new_n2149_), .Y(_abc_41356_new_n6862_));
AND2X2 AND2X2_329 ( .A(_abc_41356_new_n530_), .B(_abc_41356_new_n1117_), .Y(_abc_41356_new_n1118_));
AND2X2 AND2X2_3290 ( .A(_abc_41356_new_n6866_), .B(_abc_41356_new_n4149_), .Y(_abc_41356_new_n6867_));
AND2X2 AND2X2_3291 ( .A(_abc_41356_new_n6865_), .B(_abc_41356_new_n6867_), .Y(_abc_41356_new_n6868_));
AND2X2 AND2X2_3292 ( .A(_abc_41356_new_n6868_), .B(_abc_41356_new_n6864_), .Y(_abc_41356_new_n6869_));
AND2X2 AND2X2_3293 ( .A(_abc_41356_new_n4148_), .B(_abc_41356_new_n2149_), .Y(_abc_41356_new_n6870_));
AND2X2 AND2X2_3294 ( .A(_abc_41356_new_n6498_), .B(pc_10_), .Y(_abc_41356_new_n6873_));
AND2X2 AND2X2_3295 ( .A(_abc_41356_new_n6878_), .B(_abc_41356_new_n6877_), .Y(_abc_41356_new_n6879_));
AND2X2 AND2X2_3296 ( .A(_abc_41356_new_n6879_), .B(_abc_41356_new_n6876_), .Y(_abc_41356_new_n6880_));
AND2X2 AND2X2_3297 ( .A(_abc_41356_new_n6880_), .B(_abc_41356_new_n6875_), .Y(_abc_41356_new_n6881_));
AND2X2 AND2X2_3298 ( .A(_abc_41356_new_n6881_), .B(_abc_41356_new_n6874_), .Y(_abc_41356_new_n6882_));
AND2X2 AND2X2_3299 ( .A(_abc_41356_new_n6883_), .B(_abc_41356_new_n6884_), .Y(_abc_41356_new_n6885_));
AND2X2 AND2X2_33 ( .A(_abc_41356_new_n551_), .B(regfil_7__0_), .Y(_abc_41356_new_n552_));
AND2X2 AND2X2_330 ( .A(_abc_41356_new_n1119_), .B(_abc_41356_new_n1099_), .Y(_abc_41356_new_n1120_));
AND2X2 AND2X2_3300 ( .A(_abc_41356_new_n6885_), .B(_abc_41356_new_n6872_), .Y(_abc_41356_new_n6886_));
AND2X2 AND2X2_3301 ( .A(_abc_41356_new_n6887_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6888_));
AND2X2 AND2X2_3302 ( .A(_abc_41356_new_n6506_), .B(pc_10_), .Y(_abc_41356_new_n6889_));
AND2X2 AND2X2_3303 ( .A(_abc_41356_new_n6504_), .B(rdatahold_2_), .Y(_abc_41356_new_n6890_));
AND2X2 AND2X2_3304 ( .A(_abc_41356_new_n6892_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__10_));
AND2X2 AND2X2_3305 ( .A(_abc_41356_new_n6860_), .B(pc_11_), .Y(_abc_41356_new_n6894_));
AND2X2 AND2X2_3306 ( .A(_abc_41356_new_n6895_), .B(_abc_41356_new_n6896_), .Y(_abc_41356_new_n6897_));
AND2X2 AND2X2_3307 ( .A(_abc_41356_new_n6903_), .B(_abc_41356_new_n6901_), .Y(_abc_41356_new_n6904_));
AND2X2 AND2X2_3308 ( .A(_abc_41356_new_n6904_), .B(_abc_41356_new_n6899_), .Y(_abc_41356_new_n6905_));
AND2X2 AND2X2_3309 ( .A(_abc_41356_new_n6905_), .B(_abc_41356_new_n6907_), .Y(_abc_41356_new_n6908_));
AND2X2 AND2X2_331 ( .A(_abc_41356_new_n712_), .B(_abc_41356_new_n1122_), .Y(_abc_41356_new_n1123_));
AND2X2 AND2X2_3310 ( .A(_abc_41356_new_n6909_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n6910_));
AND2X2 AND2X2_3311 ( .A(_abc_41356_new_n2199_), .B(_abc_41356_new_n2023_), .Y(_abc_41356_new_n6911_));
AND2X2 AND2X2_3312 ( .A(_abc_41356_new_n6897_), .B(_abc_41356_new_n3495_), .Y(_abc_41356_new_n6912_));
AND2X2 AND2X2_3313 ( .A(_abc_41356_new_n6498_), .B(pc_11_), .Y(_abc_41356_new_n6913_));
AND2X2 AND2X2_3314 ( .A(_abc_41356_new_n1417_), .B(regfil_4__3_), .Y(_abc_41356_new_n6914_));
AND2X2 AND2X2_3315 ( .A(_abc_41356_new_n2191_), .B(_abc_41356_new_n6490_), .Y(_abc_41356_new_n6916_));
AND2X2 AND2X2_3316 ( .A(_abc_41356_new_n6487_), .B(_abc_41356_new_n2199_), .Y(_abc_41356_new_n6917_));
AND2X2 AND2X2_3317 ( .A(_abc_41356_new_n6920_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n6921_));
AND2X2 AND2X2_3318 ( .A(_abc_41356_new_n6923_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6924_));
AND2X2 AND2X2_3319 ( .A(_abc_41356_new_n6506_), .B(pc_11_), .Y(_abc_41356_new_n6925_));
AND2X2 AND2X2_332 ( .A(_abc_41356_new_n718_), .B(\data[6] ), .Y(_abc_41356_new_n1127_));
AND2X2 AND2X2_3320 ( .A(_abc_41356_new_n6504_), .B(rdatahold_3_), .Y(_abc_41356_new_n6926_));
AND2X2 AND2X2_3321 ( .A(_abc_41356_new_n6928_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__11_));
AND2X2 AND2X2_3322 ( .A(_abc_41356_new_n6895_), .B(_abc_41356_new_n2227_), .Y(_abc_41356_new_n6930_));
AND2X2 AND2X2_3323 ( .A(_abc_41356_new_n6894_), .B(pc_12_), .Y(_abc_41356_new_n6931_));
AND2X2 AND2X2_3324 ( .A(_abc_41356_new_n6935_), .B(_abc_41356_new_n6934_), .Y(_abc_41356_new_n6936_));
AND2X2 AND2X2_3325 ( .A(_abc_41356_new_n6936_), .B(_abc_41356_new_n4149_), .Y(_abc_41356_new_n6937_));
AND2X2 AND2X2_3326 ( .A(_abc_41356_new_n6937_), .B(_abc_41356_new_n6933_), .Y(_abc_41356_new_n6938_));
AND2X2 AND2X2_3327 ( .A(_abc_41356_new_n6940_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n6941_));
AND2X2 AND2X2_3328 ( .A(_abc_41356_new_n6939_), .B(_abc_41356_new_n6941_), .Y(_abc_41356_new_n6942_));
AND2X2 AND2X2_3329 ( .A(_abc_41356_new_n2238_), .B(_abc_41356_new_n2023_), .Y(_abc_41356_new_n6943_));
AND2X2 AND2X2_333 ( .A(_abc_41356_new_n1128_), .B(_abc_41356_new_n1126_), .Y(_abc_41356_new_n1129_));
AND2X2 AND2X2_3330 ( .A(_abc_41356_new_n2230_), .B(_abc_41356_new_n6490_), .Y(_abc_41356_new_n6944_));
AND2X2 AND2X2_3331 ( .A(_abc_41356_new_n6945_), .B(_abc_41356_new_n3495_), .Y(_abc_41356_new_n6946_));
AND2X2 AND2X2_3332 ( .A(_abc_41356_new_n2238_), .B(_abc_41356_new_n6487_), .Y(_abc_41356_new_n6947_));
AND2X2 AND2X2_3333 ( .A(_abc_41356_new_n1237_), .B(_abc_41356_new_n2248_), .Y(_abc_41356_new_n6948_));
AND2X2 AND2X2_3334 ( .A(_abc_41356_new_n6498_), .B(pc_12_), .Y(_abc_41356_new_n6949_));
AND2X2 AND2X2_3335 ( .A(_abc_41356_new_n6953_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n6954_));
AND2X2 AND2X2_3336 ( .A(_abc_41356_new_n6956_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6957_));
AND2X2 AND2X2_3337 ( .A(_abc_41356_new_n6506_), .B(pc_12_), .Y(_abc_41356_new_n6958_));
AND2X2 AND2X2_3338 ( .A(_abc_41356_new_n6504_), .B(rdatahold_4_), .Y(_abc_41356_new_n6959_));
AND2X2 AND2X2_3339 ( .A(_abc_41356_new_n6961_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__12_));
AND2X2 AND2X2_334 ( .A(_abc_41356_new_n1124_), .B(_abc_41356_new_n1129_), .Y(_abc_41356_new_n1130_));
AND2X2 AND2X2_3340 ( .A(_abc_41356_new_n6931_), .B(pc_13_), .Y(_abc_41356_new_n6963_));
AND2X2 AND2X2_3341 ( .A(_abc_41356_new_n6964_), .B(_abc_41356_new_n6965_), .Y(_abc_41356_new_n6966_));
AND2X2 AND2X2_3342 ( .A(_abc_41356_new_n6966_), .B(_abc_41356_new_n677_), .Y(_abc_41356_new_n6967_));
AND2X2 AND2X2_3343 ( .A(_abc_41356_new_n2269_), .B(_abc_41356_new_n4124_), .Y(_abc_41356_new_n6968_));
AND2X2 AND2X2_3344 ( .A(_abc_41356_new_n6538_), .B(_abc_41356_new_n2277_), .Y(_abc_41356_new_n6969_));
AND2X2 AND2X2_3345 ( .A(_abc_41356_new_n6973_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n6974_));
AND2X2 AND2X2_3346 ( .A(_abc_41356_new_n6972_), .B(_abc_41356_new_n6974_), .Y(_abc_41356_new_n6975_));
AND2X2 AND2X2_3347 ( .A(_abc_41356_new_n2277_), .B(_abc_41356_new_n2023_), .Y(_abc_41356_new_n6976_));
AND2X2 AND2X2_3348 ( .A(_abc_41356_new_n6966_), .B(_abc_41356_new_n3495_), .Y(_abc_41356_new_n6977_));
AND2X2 AND2X2_3349 ( .A(_abc_41356_new_n2269_), .B(_abc_41356_new_n6490_), .Y(_abc_41356_new_n6978_));
AND2X2 AND2X2_335 ( .A(_abc_41356_new_n1121_), .B(_abc_41356_new_n1130_), .Y(_abc_41356_new_n1131_));
AND2X2 AND2X2_3350 ( .A(_abc_41356_new_n1417_), .B(regfil_4__5_), .Y(_abc_41356_new_n6979_));
AND2X2 AND2X2_3351 ( .A(_abc_41356_new_n2277_), .B(_abc_41356_new_n6487_), .Y(_abc_41356_new_n6981_));
AND2X2 AND2X2_3352 ( .A(_abc_41356_new_n6498_), .B(pc_13_), .Y(_abc_41356_new_n6982_));
AND2X2 AND2X2_3353 ( .A(_abc_41356_new_n6985_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n6986_));
AND2X2 AND2X2_3354 ( .A(_abc_41356_new_n6988_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n6989_));
AND2X2 AND2X2_3355 ( .A(_abc_41356_new_n6506_), .B(pc_13_), .Y(_abc_41356_new_n6990_));
AND2X2 AND2X2_3356 ( .A(_abc_41356_new_n6504_), .B(rdatahold_5_), .Y(_abc_41356_new_n6991_));
AND2X2 AND2X2_3357 ( .A(_abc_41356_new_n6993_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__13_));
AND2X2 AND2X2_3358 ( .A(_abc_41356_new_n2307_), .B(_abc_41356_new_n4124_), .Y(_abc_41356_new_n6995_));
AND2X2 AND2X2_3359 ( .A(_abc_41356_new_n6963_), .B(pc_14_), .Y(_abc_41356_new_n6996_));
AND2X2 AND2X2_336 ( .A(_abc_41356_new_n1096_), .B(_abc_41356_new_n1131_), .Y(_abc_41356_new_n1132_));
AND2X2 AND2X2_3360 ( .A(_abc_41356_new_n6997_), .B(_abc_41356_new_n6998_), .Y(_abc_41356_new_n6999_));
AND2X2 AND2X2_3361 ( .A(_abc_41356_new_n6999_), .B(_abc_41356_new_n677_), .Y(_abc_41356_new_n7000_));
AND2X2 AND2X2_3362 ( .A(_abc_41356_new_n2315_), .B(_abc_41356_new_n6538_), .Y(_abc_41356_new_n7001_));
AND2X2 AND2X2_3363 ( .A(_abc_41356_new_n7005_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n7006_));
AND2X2 AND2X2_3364 ( .A(_abc_41356_new_n7004_), .B(_abc_41356_new_n7006_), .Y(_abc_41356_new_n7007_));
AND2X2 AND2X2_3365 ( .A(_abc_41356_new_n2315_), .B(_abc_41356_new_n2023_), .Y(_abc_41356_new_n7008_));
AND2X2 AND2X2_3366 ( .A(_abc_41356_new_n2307_), .B(_abc_41356_new_n6490_), .Y(_abc_41356_new_n7009_));
AND2X2 AND2X2_3367 ( .A(_abc_41356_new_n2315_), .B(_abc_41356_new_n6487_), .Y(_abc_41356_new_n7010_));
AND2X2 AND2X2_3368 ( .A(_abc_41356_new_n6999_), .B(_abc_41356_new_n3495_), .Y(_abc_41356_new_n7011_));
AND2X2 AND2X2_3369 ( .A(_abc_41356_new_n6498_), .B(pc_14_), .Y(_abc_41356_new_n7012_));
AND2X2 AND2X2_337 ( .A(_abc_41356_new_n1078_), .B(_abc_41356_new_n1134_), .Y(_abc_41356_new_n1136_));
AND2X2 AND2X2_3370 ( .A(_abc_41356_new_n7016_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n7017_));
AND2X2 AND2X2_3371 ( .A(_abc_41356_new_n7019_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n7020_));
AND2X2 AND2X2_3372 ( .A(_abc_41356_new_n6506_), .B(pc_14_), .Y(_abc_41356_new_n7021_));
AND2X2 AND2X2_3373 ( .A(_abc_41356_new_n6504_), .B(rdatahold_6_), .Y(_abc_41356_new_n7022_));
AND2X2 AND2X2_3374 ( .A(_abc_41356_new_n7024_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__14_));
AND2X2 AND2X2_3375 ( .A(_abc_41356_new_n2345_), .B(_abc_41356_new_n4124_), .Y(_abc_41356_new_n7026_));
AND2X2 AND2X2_3376 ( .A(_abc_41356_new_n6996_), .B(pc_15_), .Y(_abc_41356_new_n7028_));
AND2X2 AND2X2_3377 ( .A(_abc_41356_new_n7029_), .B(_abc_41356_new_n7027_), .Y(_abc_41356_new_n7030_));
AND2X2 AND2X2_3378 ( .A(_abc_41356_new_n7030_), .B(_abc_41356_new_n677_), .Y(_abc_41356_new_n7031_));
AND2X2 AND2X2_3379 ( .A(_abc_41356_new_n2353_), .B(_abc_41356_new_n6538_), .Y(_abc_41356_new_n7032_));
AND2X2 AND2X2_338 ( .A(_abc_41356_new_n1137_), .B(_abc_41356_new_n1135_), .Y(_abc_41356_new_n1138_));
AND2X2 AND2X2_3380 ( .A(_abc_41356_new_n7036_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n7037_));
AND2X2 AND2X2_3381 ( .A(_abc_41356_new_n7035_), .B(_abc_41356_new_n7037_), .Y(_abc_41356_new_n7038_));
AND2X2 AND2X2_3382 ( .A(_abc_41356_new_n2345_), .B(_abc_41356_new_n6490_), .Y(_abc_41356_new_n7039_));
AND2X2 AND2X2_3383 ( .A(_abc_41356_new_n7030_), .B(_abc_41356_new_n3495_), .Y(_abc_41356_new_n7040_));
AND2X2 AND2X2_3384 ( .A(_abc_41356_new_n2353_), .B(_abc_41356_new_n6487_), .Y(_abc_41356_new_n7041_));
AND2X2 AND2X2_3385 ( .A(_abc_41356_new_n6498_), .B(pc_15_), .Y(_abc_41356_new_n7042_));
AND2X2 AND2X2_3386 ( .A(_abc_41356_new_n7046_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n7047_));
AND2X2 AND2X2_3387 ( .A(_abc_41356_new_n2353_), .B(_abc_41356_new_n2023_), .Y(_abc_41356_new_n7048_));
AND2X2 AND2X2_3388 ( .A(_abc_41356_new_n7050_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n7051_));
AND2X2 AND2X2_3389 ( .A(_abc_41356_new_n6506_), .B(pc_15_), .Y(_abc_41356_new_n7052_));
AND2X2 AND2X2_339 ( .A(_abc_41356_new_n1083_), .B(regfil_0__7_), .Y(_abc_41356_new_n1141_));
AND2X2 AND2X2_3390 ( .A(_abc_41356_new_n6504_), .B(rdatahold_7_), .Y(_abc_41356_new_n7053_));
AND2X2 AND2X2_3391 ( .A(_abc_41356_new_n7055_), .B(_abc_41356_new_n509_), .Y(_0pc_15_0__15_));
AND2X2 AND2X2_3392 ( .A(_abc_41356_new_n519_), .B(_abc_41356_new_n3431_), .Y(_abc_41356_new_n7057_));
AND2X2 AND2X2_3393 ( .A(_abc_41356_new_n3423_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n7058_));
AND2X2 AND2X2_3394 ( .A(_abc_41356_new_n509_), .B(writemem), .Y(_abc_41356_new_n7061_));
AND2X2 AND2X2_3395 ( .A(_abc_41356_new_n7060_), .B(_abc_41356_new_n7061_), .Y(_abc_41356_new_n7062_));
AND2X2 AND2X2_3396 ( .A(_abc_41356_new_n3441_), .B(_abc_41356_new_n7064_), .Y(_abc_41356_new_n7065_));
AND2X2 AND2X2_3397 ( .A(_abc_41356_new_n3345_), .B(_abc_41356_new_n4118_), .Y(_abc_41356_new_n7066_));
AND2X2 AND2X2_3398 ( .A(_abc_41356_new_n7068_), .B(waitr), .Y(_abc_41356_new_n7069_));
AND2X2 AND2X2_3399 ( .A(_abc_41356_new_n4117_), .B(_abc_41356_new_n2049_), .Y(_abc_41356_new_n7073_));
AND2X2 AND2X2_34 ( .A(_abc_41356_new_n547_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n554_));
AND2X2 AND2X2_340 ( .A(_abc_41356_new_n1084_), .B(_abc_41356_new_n1134_), .Y(_abc_41356_new_n1142_));
AND2X2 AND2X2_3400 ( .A(_abc_41356_new_n7075_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7076_));
AND2X2 AND2X2_3401 ( .A(_abc_41356_new_n7071_), .B(_abc_41356_new_n7076_), .Y(_0readmem_0_0_));
AND2X2 AND2X2_3402 ( .A(_abc_41356_new_n2388_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n7078_));
AND2X2 AND2X2_3403 ( .A(_abc_41356_new_n713_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n7079_));
AND2X2 AND2X2_3404 ( .A(_abc_41356_new_n7066_), .B(_abc_41356_new_n3699_), .Y(_abc_41356_new_n7082_));
AND2X2 AND2X2_3405 ( .A(_abc_41356_new_n7082_), .B(_abc_41356_new_n7081_), .Y(_abc_41356_new_n7083_));
AND2X2 AND2X2_3406 ( .A(_abc_41356_new_n7084_), .B(\addr[0] ), .Y(_abc_41356_new_n7085_));
AND2X2 AND2X2_3407 ( .A(_abc_41356_new_n7080_), .B(rdatahold_0_), .Y(_abc_41356_new_n7086_));
AND2X2 AND2X2_3408 ( .A(_abc_41356_new_n3698_), .B(waddrhold_0_), .Y(_abc_41356_new_n7087_));
AND2X2 AND2X2_3409 ( .A(_abc_41356_new_n3205_), .B(pc_0_), .Y(_abc_41356_new_n7088_));
AND2X2 AND2X2_341 ( .A(_abc_41356_new_n1143_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n1144_));
AND2X2 AND2X2_3410 ( .A(_abc_41356_new_n4117_), .B(raddrhold_0_), .Y(_abc_41356_new_n7090_));
AND2X2 AND2X2_3411 ( .A(_abc_41356_new_n7092_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7093_));
AND2X2 AND2X2_3412 ( .A(_abc_41356_new_n7084_), .B(\addr[1] ), .Y(_abc_41356_new_n7095_));
AND2X2 AND2X2_3413 ( .A(_abc_41356_new_n7080_), .B(rdatahold_1_), .Y(_abc_41356_new_n7096_));
AND2X2 AND2X2_3414 ( .A(_abc_41356_new_n3698_), .B(waddrhold_1_), .Y(_abc_41356_new_n7097_));
AND2X2 AND2X2_3415 ( .A(_abc_41356_new_n3205_), .B(pc_1_), .Y(_abc_41356_new_n7098_));
AND2X2 AND2X2_3416 ( .A(_abc_41356_new_n4117_), .B(raddrhold_1_), .Y(_abc_41356_new_n7100_));
AND2X2 AND2X2_3417 ( .A(_abc_41356_new_n7102_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7103_));
AND2X2 AND2X2_3418 ( .A(_abc_41356_new_n7084_), .B(\addr[2] ), .Y(_abc_41356_new_n7105_));
AND2X2 AND2X2_3419 ( .A(_abc_41356_new_n7080_), .B(rdatahold_2_), .Y(_abc_41356_new_n7106_));
AND2X2 AND2X2_342 ( .A(_abc_41356_new_n616_), .B(regfil_1__7_), .Y(_abc_41356_new_n1145_));
AND2X2 AND2X2_3420 ( .A(_abc_41356_new_n3698_), .B(waddrhold_2_), .Y(_abc_41356_new_n7107_));
AND2X2 AND2X2_3421 ( .A(_abc_41356_new_n3205_), .B(pc_2_), .Y(_abc_41356_new_n7108_));
AND2X2 AND2X2_3422 ( .A(_abc_41356_new_n4117_), .B(raddrhold_2_), .Y(_abc_41356_new_n7110_));
AND2X2 AND2X2_3423 ( .A(_abc_41356_new_n7112_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7113_));
AND2X2 AND2X2_3424 ( .A(_abc_41356_new_n7084_), .B(\addr[3] ), .Y(_abc_41356_new_n7115_));
AND2X2 AND2X2_3425 ( .A(_abc_41356_new_n7080_), .B(rdatahold_3_), .Y(_abc_41356_new_n7116_));
AND2X2 AND2X2_3426 ( .A(_abc_41356_new_n3698_), .B(waddrhold_3_), .Y(_abc_41356_new_n7117_));
AND2X2 AND2X2_3427 ( .A(_abc_41356_new_n3205_), .B(pc_3_), .Y(_abc_41356_new_n7118_));
AND2X2 AND2X2_3428 ( .A(_abc_41356_new_n4117_), .B(raddrhold_3_), .Y(_abc_41356_new_n7120_));
AND2X2 AND2X2_3429 ( .A(_abc_41356_new_n7122_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7123_));
AND2X2 AND2X2_343 ( .A(_abc_41356_new_n619_), .B(regfil_0__7_), .Y(_abc_41356_new_n1146_));
AND2X2 AND2X2_3430 ( .A(_abc_41356_new_n7084_), .B(\addr[4] ), .Y(_abc_41356_new_n7125_));
AND2X2 AND2X2_3431 ( .A(_abc_41356_new_n7080_), .B(rdatahold_4_), .Y(_abc_41356_new_n7126_));
AND2X2 AND2X2_3432 ( .A(_abc_41356_new_n3698_), .B(waddrhold_4_), .Y(_abc_41356_new_n7127_));
AND2X2 AND2X2_3433 ( .A(_abc_41356_new_n3205_), .B(pc_4_), .Y(_abc_41356_new_n7128_));
AND2X2 AND2X2_3434 ( .A(_abc_41356_new_n4117_), .B(raddrhold_4_), .Y(_abc_41356_new_n7130_));
AND2X2 AND2X2_3435 ( .A(_abc_41356_new_n7132_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7133_));
AND2X2 AND2X2_3436 ( .A(_abc_41356_new_n7084_), .B(\addr[5] ), .Y(_abc_41356_new_n7135_));
AND2X2 AND2X2_3437 ( .A(_abc_41356_new_n7080_), .B(rdatahold_5_), .Y(_abc_41356_new_n7136_));
AND2X2 AND2X2_3438 ( .A(_abc_41356_new_n3698_), .B(waddrhold_5_), .Y(_abc_41356_new_n7137_));
AND2X2 AND2X2_3439 ( .A(_abc_41356_new_n3205_), .B(pc_5_), .Y(_abc_41356_new_n7138_));
AND2X2 AND2X2_344 ( .A(_abc_41356_new_n526_), .B(regfil_3__7_), .Y(_abc_41356_new_n1148_));
AND2X2 AND2X2_3440 ( .A(_abc_41356_new_n4117_), .B(raddrhold_5_), .Y(_abc_41356_new_n7140_));
AND2X2 AND2X2_3441 ( .A(_abc_41356_new_n7142_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7143_));
AND2X2 AND2X2_3442 ( .A(_abc_41356_new_n7084_), .B(\addr[6] ), .Y(_abc_41356_new_n7145_));
AND2X2 AND2X2_3443 ( .A(_abc_41356_new_n7080_), .B(rdatahold_6_), .Y(_abc_41356_new_n7146_));
AND2X2 AND2X2_3444 ( .A(_abc_41356_new_n3698_), .B(waddrhold_6_), .Y(_abc_41356_new_n7147_));
AND2X2 AND2X2_3445 ( .A(_abc_41356_new_n3205_), .B(pc_6_), .Y(_abc_41356_new_n7148_));
AND2X2 AND2X2_3446 ( .A(_abc_41356_new_n4117_), .B(raddrhold_6_), .Y(_abc_41356_new_n7150_));
AND2X2 AND2X2_3447 ( .A(_abc_41356_new_n7152_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7153_));
AND2X2 AND2X2_3448 ( .A(_abc_41356_new_n7084_), .B(\addr[7] ), .Y(_abc_41356_new_n7155_));
AND2X2 AND2X2_3449 ( .A(_abc_41356_new_n7080_), .B(rdatahold_7_), .Y(_abc_41356_new_n7156_));
AND2X2 AND2X2_345 ( .A(_abc_41356_new_n623_), .B(regfil_2__7_), .Y(_abc_41356_new_n1149_));
AND2X2 AND2X2_3450 ( .A(_abc_41356_new_n3698_), .B(waddrhold_7_), .Y(_abc_41356_new_n7157_));
AND2X2 AND2X2_3451 ( .A(_abc_41356_new_n3205_), .B(pc_7_), .Y(_abc_41356_new_n7158_));
AND2X2 AND2X2_3452 ( .A(_abc_41356_new_n4117_), .B(raddrhold_7_), .Y(_abc_41356_new_n7160_));
AND2X2 AND2X2_3453 ( .A(_abc_41356_new_n7162_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7163_));
AND2X2 AND2X2_3454 ( .A(_abc_41356_new_n7084_), .B(\addr[8] ), .Y(_abc_41356_new_n7165_));
AND2X2 AND2X2_3455 ( .A(_abc_41356_new_n4117_), .B(raddrhold_8_), .Y(_abc_41356_new_n7166_));
AND2X2 AND2X2_3456 ( .A(_abc_41356_new_n3698_), .B(waddrhold_8_), .Y(_abc_41356_new_n7167_));
AND2X2 AND2X2_3457 ( .A(_abc_41356_new_n3205_), .B(pc_8_), .Y(_abc_41356_new_n7168_));
AND2X2 AND2X2_3458 ( .A(_abc_41356_new_n7170_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7171_));
AND2X2 AND2X2_3459 ( .A(_abc_41356_new_n7084_), .B(\addr[9] ), .Y(_abc_41356_new_n7173_));
AND2X2 AND2X2_346 ( .A(_abc_41356_new_n616_), .B(regfil_5__7_), .Y(_abc_41356_new_n1153_));
AND2X2 AND2X2_3460 ( .A(_abc_41356_new_n5295_), .B(waddrhold_9_), .Y(_abc_41356_new_n7174_));
AND2X2 AND2X2_3461 ( .A(_abc_41356_new_n519_), .B(_abc_41356_new_n2926_), .Y(_abc_41356_new_n7175_));
AND2X2 AND2X2_3462 ( .A(_abc_41356_new_n7175_), .B(pc_9_), .Y(_abc_41356_new_n7176_));
AND2X2 AND2X2_3463 ( .A(_abc_41356_new_n509_), .B(raddrhold_9_), .Y(_abc_41356_new_n7177_));
AND2X2 AND2X2_3464 ( .A(_abc_41356_new_n4117_), .B(_abc_41356_new_n7177_), .Y(_abc_41356_new_n7178_));
AND2X2 AND2X2_3465 ( .A(_abc_41356_new_n7084_), .B(\addr[10] ), .Y(_abc_41356_new_n7182_));
AND2X2 AND2X2_3466 ( .A(_abc_41356_new_n5295_), .B(waddrhold_10_), .Y(_abc_41356_new_n7183_));
AND2X2 AND2X2_3467 ( .A(_abc_41356_new_n7175_), .B(pc_10_), .Y(_abc_41356_new_n7184_));
AND2X2 AND2X2_3468 ( .A(_abc_41356_new_n509_), .B(raddrhold_10_), .Y(_abc_41356_new_n7185_));
AND2X2 AND2X2_3469 ( .A(_abc_41356_new_n4117_), .B(_abc_41356_new_n7185_), .Y(_abc_41356_new_n7186_));
AND2X2 AND2X2_347 ( .A(_abc_41356_new_n623_), .B(regfil_6__7_), .Y(_abc_41356_new_n1155_));
AND2X2 AND2X2_3470 ( .A(_abc_41356_new_n7084_), .B(\addr[11] ), .Y(_abc_41356_new_n7190_));
AND2X2 AND2X2_3471 ( .A(_abc_41356_new_n5295_), .B(waddrhold_11_), .Y(_abc_41356_new_n7191_));
AND2X2 AND2X2_3472 ( .A(_abc_41356_new_n7175_), .B(pc_11_), .Y(_abc_41356_new_n7192_));
AND2X2 AND2X2_3473 ( .A(_abc_41356_new_n509_), .B(raddrhold_11_), .Y(_abc_41356_new_n7193_));
AND2X2 AND2X2_3474 ( .A(_abc_41356_new_n4117_), .B(_abc_41356_new_n7193_), .Y(_abc_41356_new_n7194_));
AND2X2 AND2X2_3475 ( .A(_abc_41356_new_n7084_), .B(\addr[12] ), .Y(_abc_41356_new_n7198_));
AND2X2 AND2X2_3476 ( .A(_abc_41356_new_n4117_), .B(raddrhold_12_), .Y(_abc_41356_new_n7199_));
AND2X2 AND2X2_3477 ( .A(_abc_41356_new_n3205_), .B(pc_12_), .Y(_abc_41356_new_n7200_));
AND2X2 AND2X2_3478 ( .A(_abc_41356_new_n3698_), .B(waddrhold_12_), .Y(_abc_41356_new_n7201_));
AND2X2 AND2X2_3479 ( .A(_abc_41356_new_n7203_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7204_));
AND2X2 AND2X2_348 ( .A(_abc_41356_new_n619_), .B(regfil_4__7_), .Y(_abc_41356_new_n1156_));
AND2X2 AND2X2_3480 ( .A(_abc_41356_new_n7084_), .B(\addr[13] ), .Y(_abc_41356_new_n7206_));
AND2X2 AND2X2_3481 ( .A(_abc_41356_new_n4117_), .B(raddrhold_13_), .Y(_abc_41356_new_n7207_));
AND2X2 AND2X2_3482 ( .A(_abc_41356_new_n3205_), .B(pc_13_), .Y(_abc_41356_new_n7208_));
AND2X2 AND2X2_3483 ( .A(_abc_41356_new_n3698_), .B(waddrhold_13_), .Y(_abc_41356_new_n7209_));
AND2X2 AND2X2_3484 ( .A(_abc_41356_new_n7211_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7212_));
AND2X2 AND2X2_3485 ( .A(_abc_41356_new_n7084_), .B(\addr[14] ), .Y(_abc_41356_new_n7214_));
AND2X2 AND2X2_3486 ( .A(_abc_41356_new_n5295_), .B(waddrhold_14_), .Y(_abc_41356_new_n7215_));
AND2X2 AND2X2_3487 ( .A(_abc_41356_new_n7175_), .B(pc_14_), .Y(_abc_41356_new_n7216_));
AND2X2 AND2X2_3488 ( .A(_abc_41356_new_n4811_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7217_));
AND2X2 AND2X2_3489 ( .A(_abc_41356_new_n7084_), .B(\addr[15] ), .Y(_abc_41356_new_n7221_));
AND2X2 AND2X2_349 ( .A(_abc_41356_new_n526_), .B(regfil_7__7_), .Y(_abc_41356_new_n1157_));
AND2X2 AND2X2_3490 ( .A(_abc_41356_new_n3205_), .B(pc_15_), .Y(_abc_41356_new_n7222_));
AND2X2 AND2X2_3491 ( .A(_abc_41356_new_n3698_), .B(waddrhold_15_), .Y(_abc_41356_new_n7223_));
AND2X2 AND2X2_3492 ( .A(_abc_41356_new_n7225_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7226_));
AND2X2 AND2X2_3493 ( .A(_abc_41356_new_n713_), .B(_abc_41356_new_n607_), .Y(_abc_41356_new_n7228_));
AND2X2 AND2X2_3494 ( .A(_abc_41356_new_n715_), .B(_abc_41356_new_n716_), .Y(_abc_41356_new_n7229_));
AND2X2 AND2X2_3495 ( .A(_abc_41356_new_n509_), .B(readio), .Y(_abc_41356_new_n7231_));
AND2X2 AND2X2_3496 ( .A(_abc_41356_new_n7230_), .B(_abc_41356_new_n7231_), .Y(_abc_41356_new_n7232_));
AND2X2 AND2X2_3497 ( .A(_abc_41356_new_n7066_), .B(_abc_41356_new_n7065_), .Y(_abc_41356_new_n7234_));
AND2X2 AND2X2_3498 ( .A(_abc_41356_new_n7234_), .B(inta), .Y(_abc_41356_new_n7235_));
AND2X2 AND2X2_3499 ( .A(_abc_41356_new_n4117_), .B(intcyc), .Y(_abc_41356_new_n7237_));
AND2X2 AND2X2_35 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n554_), .Y(_abc_41356_new_n555_));
AND2X2 AND2X2_350 ( .A(_abc_41356_new_n1152_), .B(_abc_41356_new_n1160_), .Y(_abc_41356_new_n1161_));
AND2X2 AND2X2_3500 ( .A(_abc_41356_new_n3205_), .B(_abc_41356_new_n3202_), .Y(_abc_41356_new_n7238_));
AND2X2 AND2X2_3501 ( .A(_abc_41356_new_n7240_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7241_));
AND2X2 AND2X2_3502 ( .A(_abc_41356_new_n7236_), .B(_abc_41356_new_n7241_), .Y(_0inta_0_0_));
AND2X2 AND2X2_3503 ( .A(_abc_41356_new_n1227_), .B(_abc_41356_new_n607_), .Y(_abc_41356_new_n7243_));
AND2X2 AND2X2_3504 ( .A(_abc_41356_new_n5842_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n7244_));
AND2X2 AND2X2_3505 ( .A(_abc_41356_new_n509_), .B(writeio), .Y(_abc_41356_new_n7247_));
AND2X2 AND2X2_3506 ( .A(_abc_41356_new_n7246_), .B(_abc_41356_new_n7247_), .Y(_abc_41356_new_n7248_));
AND2X2 AND2X2_3507 ( .A(_abc_41356_new_n7250_), .B(_abc_41356_new_n3553_), .Y(_abc_41356_new_n7251_));
AND2X2 AND2X2_3508 ( .A(_abc_41356_new_n7251_), .B(_abc_41356_new_n3489_), .Y(_abc_41356_new_n7252_));
AND2X2 AND2X2_3509 ( .A(_abc_41356_new_n3489_), .B(_abc_41356_new_n3554_), .Y(_abc_41356_new_n7253_));
AND2X2 AND2X2_351 ( .A(_abc_41356_new_n1161_), .B(_abc_41356_new_n614_), .Y(_abc_41356_new_n1162_));
AND2X2 AND2X2_3510 ( .A(_abc_41356_new_n7250_), .B(statesel_3_), .Y(_abc_41356_new_n7254_));
AND2X2 AND2X2_3511 ( .A(_abc_41356_new_n3487_), .B(_abc_41356_new_n7254_), .Y(_abc_41356_new_n7255_));
AND2X2 AND2X2_3512 ( .A(_abc_41356_new_n7258_), .B(_abc_41356_new_n3608_), .Y(_abc_41356_new_n7259_));
AND2X2 AND2X2_3513 ( .A(_abc_41356_new_n7260_), .B(statesel_5_), .Y(_abc_41356_new_n7261_));
AND2X2 AND2X2_3514 ( .A(_abc_41356_new_n7263_), .B(_abc_41356_new_n3487_), .Y(_abc_41356_new_n7264_));
AND2X2 AND2X2_3515 ( .A(_abc_41356_new_n7264_), .B(_abc_41356_new_n7262_), .Y(_abc_41356_new_n7265_));
AND2X2 AND2X2_3516 ( .A(_abc_41356_new_n3489_), .B(_abc_41356_new_n7250_), .Y(_abc_41356_new_n7266_));
AND2X2 AND2X2_3517 ( .A(_abc_41356_new_n7268_), .B(_abc_41356_new_n7261_), .Y(_abc_41356_new_n7269_));
AND2X2 AND2X2_3518 ( .A(_abc_41356_new_n3449_), .B(_abc_41356_new_n3488_), .Y(_abc_41356_new_n7270_));
AND2X2 AND2X2_3519 ( .A(statesel_4_), .B(statesel_5_), .Y(_abc_41356_new_n7271_));
AND2X2 AND2X2_352 ( .A(_abc_41356_new_n606_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n1163_));
AND2X2 AND2X2_3520 ( .A(_abc_41356_new_n7271_), .B(_abc_41356_new_n7250_), .Y(_abc_41356_new_n7272_));
AND2X2 AND2X2_3521 ( .A(_abc_41356_new_n7272_), .B(_abc_41356_new_n7270_), .Y(_abc_41356_new_n7273_));
AND2X2 AND2X2_3522 ( .A(_abc_41356_new_n7262_), .B(_abc_41356_new_n7263_), .Y(_abc_41356_new_n7274_));
AND2X2 AND2X2_3523 ( .A(_abc_41356_new_n7260_), .B(_abc_41356_new_n3594_), .Y(_abc_41356_new_n7276_));
AND2X2 AND2X2_3524 ( .A(_abc_41356_new_n7276_), .B(_abc_41356_new_n3449_), .Y(_abc_41356_new_n7277_));
AND2X2 AND2X2_3525 ( .A(_abc_41356_new_n7275_), .B(_abc_41356_new_n7277_), .Y(_abc_41356_new_n7278_));
AND2X2 AND2X2_3526 ( .A(_abc_41356_new_n3454_), .B(_abc_41356_new_n7282_), .Y(_abc_41356_new_n7283_));
AND2X2 AND2X2_3527 ( .A(_abc_41356_new_n516_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7285_));
AND2X2 AND2X2_3528 ( .A(_abc_41356_new_n4128_), .B(_abc_41356_new_n7285_), .Y(_abc_41356_new_n7286_));
AND2X2 AND2X2_3529 ( .A(_abc_41356_new_n7291_), .B(_abc_41356_new_n4156_), .Y(_abc_41356_new_n7292_));
AND2X2 AND2X2_353 ( .A(_abc_41356_new_n509_), .B(rdatahold_7_), .Y(_abc_41356_new_n1164_));
AND2X2 AND2X2_3530 ( .A(_abc_41356_new_n525_), .B(_abc_41356_new_n3279_), .Y(_abc_41356_new_n7295_));
AND2X2 AND2X2_3531 ( .A(_abc_41356_new_n4160_), .B(_abc_41356_new_n7295_), .Y(_abc_41356_new_n7296_));
AND2X2 AND2X2_3532 ( .A(_abc_41356_new_n7298_), .B(opcode_5_), .Y(_abc_41356_new_n7299_));
AND2X2 AND2X2_3533 ( .A(_abc_41356_new_n7300_), .B(_abc_41356_new_n7297_), .Y(_abc_41356_new_n7301_));
AND2X2 AND2X2_3534 ( .A(_abc_41356_new_n545_), .B(zero), .Y(_abc_41356_new_n7303_));
AND2X2 AND2X2_3535 ( .A(_abc_41356_new_n7305_), .B(_abc_41356_new_n576_), .Y(_abc_41356_new_n7306_));
AND2X2 AND2X2_3536 ( .A(_abc_41356_new_n7306_), .B(_abc_41356_new_n7304_), .Y(_abc_41356_new_n7307_));
AND2X2 AND2X2_3537 ( .A(_abc_41356_new_n682_), .B(_abc_41356_new_n7298_), .Y(_abc_41356_new_n7308_));
AND2X2 AND2X2_3538 ( .A(_abc_41356_new_n7310_), .B(_abc_41356_new_n7302_), .Y(_abc_41356_new_n7311_));
AND2X2 AND2X2_3539 ( .A(_abc_41356_new_n7292_), .B(_abc_41356_new_n7312_), .Y(_abc_41356_new_n7313_));
AND2X2 AND2X2_354 ( .A(_abc_41356_new_n1163_), .B(_abc_41356_new_n1164_), .Y(_abc_41356_new_n1165_));
AND2X2 AND2X2_3540 ( .A(_abc_41356_new_n3600_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7315_));
AND2X2 AND2X2_3541 ( .A(_abc_41356_new_n683_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7316_));
AND2X2 AND2X2_3542 ( .A(_abc_41356_new_n7316_), .B(_abc_41356_new_n4183_), .Y(_abc_41356_new_n7317_));
AND2X2 AND2X2_3543 ( .A(_abc_41356_new_n1233_), .B(opcode_5_), .Y(_abc_41356_new_n7318_));
AND2X2 AND2X2_3544 ( .A(_abc_41356_new_n7319_), .B(_abc_41356_new_n7321_), .Y(_abc_41356_new_n7322_));
AND2X2 AND2X2_3545 ( .A(_abc_41356_new_n7323_), .B(_abc_41356_new_n7318_), .Y(_abc_41356_new_n7324_));
AND2X2 AND2X2_3546 ( .A(_abc_41356_new_n7324_), .B(_abc_41356_new_n7293_), .Y(_abc_41356_new_n7325_));
AND2X2 AND2X2_3547 ( .A(_abc_41356_new_n7314_), .B(_abc_41356_new_n7328_), .Y(_abc_41356_new_n7329_));
AND2X2 AND2X2_3548 ( .A(_abc_41356_new_n7287_), .B(_abc_41356_new_n7329_), .Y(_abc_41356_new_n7330_));
AND2X2 AND2X2_3549 ( .A(_abc_41356_new_n7331_), .B(_abc_41356_new_n7284_), .Y(_abc_41356_new_n7332_));
AND2X2 AND2X2_355 ( .A(_abc_41356_new_n612_), .B(alu_res_7_), .Y(_abc_41356_new_n1166_));
AND2X2 AND2X2_3550 ( .A(_abc_41356_new_n7334_), .B(_abc_41356_new_n2928_), .Y(_abc_41356_new_n7335_));
AND2X2 AND2X2_3551 ( .A(_abc_41356_new_n3454_), .B(_abc_41356_new_n7271_), .Y(_abc_41356_new_n7337_));
AND2X2 AND2X2_3552 ( .A(_abc_41356_new_n7340_), .B(_abc_41356_new_n7336_), .Y(_abc_41356_new_n7341_));
AND2X2 AND2X2_3553 ( .A(_abc_41356_new_n7270_), .B(_abc_41356_new_n3580_), .Y(_abc_41356_new_n7343_));
AND2X2 AND2X2_3554 ( .A(_abc_41356_new_n7349_), .B(_abc_41356_new_n7345_), .Y(_abc_41356_new_n7350_));
AND2X2 AND2X2_3555 ( .A(_abc_41356_new_n7351_), .B(_abc_41356_new_n5414_), .Y(_abc_41356_new_n7352_));
AND2X2 AND2X2_3556 ( .A(_abc_41356_new_n7353_), .B(_abc_41356_new_n7354_), .Y(_abc_41356_new_n7355_));
AND2X2 AND2X2_3557 ( .A(_abc_41356_new_n7352_), .B(_abc_41356_new_n7355_), .Y(_abc_41356_new_n7356_));
AND2X2 AND2X2_3558 ( .A(_abc_41356_new_n7341_), .B(_abc_41356_new_n7356_), .Y(_abc_41356_new_n7357_));
AND2X2 AND2X2_3559 ( .A(_abc_41356_new_n7357_), .B(_abc_41356_new_n7332_), .Y(_abc_41356_new_n7358_));
AND2X2 AND2X2_356 ( .A(_abc_41356_new_n1168_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n1169_));
AND2X2 AND2X2_3560 ( .A(_abc_41356_new_n3454_), .B(_abc_41356_new_n7261_), .Y(_abc_41356_new_n7359_));
AND2X2 AND2X2_3561 ( .A(_abc_41356_new_n7251_), .B(_abc_41356_new_n3520_), .Y(_abc_41356_new_n7361_));
AND2X2 AND2X2_3562 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n4827_), .Y(_abc_41356_new_n7366_));
AND2X2 AND2X2_3563 ( .A(_abc_41356_new_n6535_), .B(_abc_41356_new_n7366_), .Y(_abc_41356_new_n7367_));
AND2X2 AND2X2_3564 ( .A(_abc_41356_new_n6521_), .B(_abc_41356_new_n7367_), .Y(_abc_41356_new_n7368_));
AND2X2 AND2X2_3565 ( .A(_abc_41356_new_n7365_), .B(_abc_41356_new_n7368_), .Y(_abc_41356_new_n7369_));
AND2X2 AND2X2_3566 ( .A(_abc_41356_new_n4130_), .B(_abc_41356_new_n7369_), .Y(_abc_41356_new_n7370_));
AND2X2 AND2X2_3567 ( .A(_abc_41356_new_n3317_), .B(_abc_41356_new_n607_), .Y(_abc_41356_new_n7372_));
AND2X2 AND2X2_3568 ( .A(_abc_41356_new_n7374_), .B(_abc_41356_new_n3321_), .Y(_abc_41356_new_n7375_));
AND2X2 AND2X2_3569 ( .A(_abc_41356_new_n7371_), .B(_abc_41356_new_n7375_), .Y(_abc_41356_new_n7376_));
AND2X2 AND2X2_357 ( .A(_abc_41356_new_n595_), .B(rdatahold_7_), .Y(_abc_41356_new_n1170_));
AND2X2 AND2X2_3570 ( .A(_abc_41356_new_n7364_), .B(_abc_41356_new_n7376_), .Y(_abc_41356_new_n7377_));
AND2X2 AND2X2_3571 ( .A(_abc_41356_new_n7377_), .B(_abc_41356_new_n7363_), .Y(_abc_41356_new_n7378_));
AND2X2 AND2X2_3572 ( .A(_abc_41356_new_n3489_), .B(_abc_41356_new_n3580_), .Y(_abc_41356_new_n7379_));
AND2X2 AND2X2_3573 ( .A(_abc_41356_new_n7380_), .B(_abc_41356_new_n7260_), .Y(_abc_41356_new_n7381_));
AND2X2 AND2X2_3574 ( .A(_abc_41356_new_n3580_), .B(_abc_41356_new_n3488_), .Y(_abc_41356_new_n7382_));
AND2X2 AND2X2_3575 ( .A(_abc_41356_new_n7362_), .B(_abc_41356_new_n7383_), .Y(_abc_41356_new_n7384_));
AND2X2 AND2X2_3576 ( .A(_abc_41356_new_n7389_), .B(_abc_41356_new_n7388_), .Y(_abc_41356_new_n7390_));
AND2X2 AND2X2_3577 ( .A(_abc_41356_new_n7339_), .B(_abc_41356_new_n7392_), .Y(_abc_41356_new_n7393_));
AND2X2 AND2X2_3578 ( .A(_abc_41356_new_n7391_), .B(_abc_41356_new_n7394_), .Y(_abc_41356_new_n7395_));
AND2X2 AND2X2_3579 ( .A(_abc_41356_new_n7395_), .B(_abc_41356_new_n7386_), .Y(_abc_41356_new_n7396_));
AND2X2 AND2X2_358 ( .A(_abc_41356_new_n1175_), .B(_abc_41356_new_n724_), .Y(_abc_41356_new_n1176_));
AND2X2 AND2X2_3580 ( .A(_abc_41356_new_n7400_), .B(_abc_41356_new_n7402_), .Y(_abc_41356_new_n7403_));
AND2X2 AND2X2_3581 ( .A(_abc_41356_new_n7398_), .B(_abc_41356_new_n7403_), .Y(_abc_41356_new_n7404_));
AND2X2 AND2X2_3582 ( .A(_abc_41356_new_n7397_), .B(_abc_41356_new_n7405_), .Y(_abc_41356_new_n7406_));
AND2X2 AND2X2_3583 ( .A(_abc_41356_new_n7276_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n7407_));
AND2X2 AND2X2_3584 ( .A(_abc_41356_new_n3451_), .B(_abc_41356_new_n7407_), .Y(_abc_41356_new_n7408_));
AND2X2 AND2X2_3585 ( .A(_abc_41356_new_n7408_), .B(_abc_41356_new_n7343_), .Y(_abc_41356_new_n7409_));
AND2X2 AND2X2_3586 ( .A(_abc_41356_new_n7270_), .B(_abc_41356_new_n3554_), .Y(_abc_41356_new_n7410_));
AND2X2 AND2X2_3587 ( .A(_abc_41356_new_n7337_), .B(_abc_41356_new_n7410_), .Y(_abc_41356_new_n7411_));
AND2X2 AND2X2_3588 ( .A(_abc_41356_new_n7413_), .B(_abc_41356_new_n7406_), .Y(_abc_41356_new_n7414_));
AND2X2 AND2X2_3589 ( .A(_abc_41356_new_n7378_), .B(_abc_41356_new_n7414_), .Y(_abc_41356_new_n7415_));
AND2X2 AND2X2_359 ( .A(_abc_41356_new_n1174_), .B(_abc_41356_new_n1176_), .Y(_abc_41356_new_n1177_));
AND2X2 AND2X2_3590 ( .A(_abc_41356_new_n715_), .B(_abc_41356_new_n3445_), .Y(_abc_41356_new_n7416_));
AND2X2 AND2X2_3591 ( .A(_abc_41356_new_n607_), .B(_abc_41356_new_n611_), .Y(_abc_41356_new_n7417_));
AND2X2 AND2X2_3592 ( .A(_abc_41356_new_n7421_), .B(_abc_41356_new_n7419_), .Y(_abc_41356_new_n7422_));
AND2X2 AND2X2_3593 ( .A(_abc_41356_new_n7251_), .B(_abc_41356_new_n7261_), .Y(_abc_41356_new_n7423_));
AND2X2 AND2X2_3594 ( .A(_abc_41356_new_n7423_), .B(_abc_41356_new_n7270_), .Y(_abc_41356_new_n7424_));
AND2X2 AND2X2_3595 ( .A(_abc_41356_new_n3487_), .B(_abc_41356_new_n3554_), .Y(_abc_41356_new_n7425_));
AND2X2 AND2X2_3596 ( .A(_abc_41356_new_n7425_), .B(_abc_41356_new_n3608_), .Y(_abc_41356_new_n7426_));
AND2X2 AND2X2_3597 ( .A(_abc_41356_new_n3454_), .B(_abc_41356_new_n7427_), .Y(_abc_41356_new_n7428_));
AND2X2 AND2X2_3598 ( .A(_abc_41356_new_n7058_), .B(_abc_41356_new_n3445_), .Y(_abc_41356_new_n7430_));
AND2X2 AND2X2_3599 ( .A(_abc_41356_new_n7244_), .B(_abc_41356_new_n717_), .Y(_abc_41356_new_n7433_));
AND2X2 AND2X2_36 ( .A(opcode_4_), .B(carry), .Y(_abc_41356_new_n556_));
AND2X2 AND2X2_360 ( .A(_abc_41356_new_n1178_), .B(_abc_41356_new_n1179_), .Y(_abc_41356_new_n1180_));
AND2X2 AND2X2_3600 ( .A(_abc_41356_new_n7432_), .B(_abc_41356_new_n7434_), .Y(_abc_41356_new_n7435_));
AND2X2 AND2X2_3601 ( .A(_abc_41356_new_n7429_), .B(_abc_41356_new_n7435_), .Y(_abc_41356_new_n7436_));
AND2X2 AND2X2_3602 ( .A(_abc_41356_new_n7436_), .B(_abc_41356_new_n7422_), .Y(_abc_41356_new_n7437_));
AND2X2 AND2X2_3603 ( .A(_abc_41356_new_n7415_), .B(_abc_41356_new_n7437_), .Y(_abc_41356_new_n7438_));
AND2X2 AND2X2_3604 ( .A(_abc_41356_new_n7438_), .B(_abc_41356_new_n7358_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_0_));
AND2X2 AND2X2_3605 ( .A(_abc_41356_new_n7440_), .B(_abc_41356_new_n7444_), .Y(_abc_41356_new_n7445_));
AND2X2 AND2X2_3606 ( .A(_abc_41356_new_n7251_), .B(_abc_41356_new_n3487_), .Y(_abc_41356_new_n7447_));
AND2X2 AND2X2_3607 ( .A(_abc_41356_new_n7254_), .B(_abc_41356_new_n3520_), .Y(_abc_41356_new_n7449_));
AND2X2 AND2X2_3608 ( .A(_abc_41356_new_n7448_), .B(_abc_41356_new_n7450_), .Y(_abc_41356_new_n7451_));
AND2X2 AND2X2_3609 ( .A(_abc_41356_new_n7453_), .B(_abc_41356_new_n5412_), .Y(_abc_41356_new_n7454_));
AND2X2 AND2X2_361 ( .A(_abc_41356_new_n712_), .B(_abc_41356_new_n1180_), .Y(_abc_41356_new_n1181_));
AND2X2 AND2X2_3610 ( .A(_abc_41356_new_n7244_), .B(_abc_41356_new_n3445_), .Y(_abc_41356_new_n7455_));
AND2X2 AND2X2_3611 ( .A(_abc_41356_new_n7454_), .B(_abc_41356_new_n7457_), .Y(_abc_41356_new_n7458_));
AND2X2 AND2X2_3612 ( .A(_abc_41356_new_n7337_), .B(_abc_41356_new_n7361_), .Y(_abc_41356_new_n7459_));
AND2X2 AND2X2_3613 ( .A(_abc_41356_new_n509_), .B(_abc_41356_new_n501_), .Y(_abc_41356_new_n7464_));
AND2X2 AND2X2_3614 ( .A(_abc_41356_new_n709_), .B(_abc_41356_new_n7464_), .Y(_abc_41356_new_n7465_));
AND2X2 AND2X2_3615 ( .A(_abc_41356_new_n7467_), .B(_abc_41356_new_n7466_), .Y(_abc_41356_new_n7468_));
AND2X2 AND2X2_3616 ( .A(_abc_41356_new_n7463_), .B(_abc_41356_new_n7468_), .Y(_abc_41356_new_n7469_));
AND2X2 AND2X2_3617 ( .A(_abc_41356_new_n7461_), .B(_abc_41356_new_n7469_), .Y(_abc_41356_new_n7470_));
AND2X2 AND2X2_3618 ( .A(_abc_41356_new_n7460_), .B(_abc_41356_new_n7470_), .Y(_abc_41356_new_n7471_));
AND2X2 AND2X2_3619 ( .A(_abc_41356_new_n7471_), .B(_abc_41356_new_n7458_), .Y(_abc_41356_new_n7472_));
AND2X2 AND2X2_362 ( .A(_abc_41356_new_n714_), .B(alu_res_7_), .Y(_abc_41356_new_n1182_));
AND2X2 AND2X2_3620 ( .A(_abc_41356_new_n7472_), .B(_abc_41356_new_n7445_), .Y(_abc_41356_new_n7473_));
AND2X2 AND2X2_3621 ( .A(_abc_41356_new_n7358_), .B(_abc_41356_new_n7414_), .Y(_abc_41356_new_n7474_));
AND2X2 AND2X2_3622 ( .A(_abc_41356_new_n7474_), .B(_abc_41356_new_n7473_), .Y(_abc_41356_new_n7475_));
AND2X2 AND2X2_3623 ( .A(_abc_41356_new_n7337_), .B(_abc_41356_new_n7343_), .Y(_abc_41356_new_n7477_));
AND2X2 AND2X2_3624 ( .A(_abc_41356_new_n7479_), .B(_abc_41356_new_n7276_), .Y(_abc_41356_new_n7480_));
AND2X2 AND2X2_3625 ( .A(_abc_41356_new_n7270_), .B(_abc_41356_new_n7254_), .Y(_abc_41356_new_n7481_));
AND2X2 AND2X2_3626 ( .A(_abc_41356_new_n7481_), .B(_abc_41356_new_n3608_), .Y(_abc_41356_new_n7482_));
AND2X2 AND2X2_3627 ( .A(_abc_41356_new_n3581_), .B(_abc_41356_new_n7261_), .Y(_abc_41356_new_n7487_));
AND2X2 AND2X2_3628 ( .A(_abc_41356_new_n7486_), .B(_abc_41356_new_n7488_), .Y(_abc_41356_new_n7489_));
AND2X2 AND2X2_3629 ( .A(_abc_41356_new_n7484_), .B(_abc_41356_new_n7489_), .Y(_abc_41356_new_n7490_));
AND2X2 AND2X2_363 ( .A(_abc_41356_new_n512_), .B(rdatahold_7_), .Y(_abc_41356_new_n1183_));
AND2X2 AND2X2_3630 ( .A(_abc_41356_new_n7359_), .B(_abc_41356_new_n7481_), .Y(_abc_41356_new_n7492_));
AND2X2 AND2X2_3631 ( .A(_abc_41356_new_n7493_), .B(_abc_41356_new_n7491_), .Y(_abc_41356_new_n7494_));
AND2X2 AND2X2_3632 ( .A(_abc_41356_new_n7494_), .B(_abc_41356_new_n7478_), .Y(_abc_41356_new_n7495_));
AND2X2 AND2X2_3633 ( .A(_abc_41356_new_n4184_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n7496_));
AND2X2 AND2X2_3634 ( .A(_abc_41356_new_n7497_), .B(_abc_41356_new_n7499_), .Y(_abc_41356_new_n7500_));
AND2X2 AND2X2_3635 ( .A(_abc_41356_new_n7434_), .B(_abc_41356_new_n7467_), .Y(_abc_41356_new_n7502_));
AND2X2 AND2X2_3636 ( .A(_abc_41356_new_n7501_), .B(_abc_41356_new_n7502_), .Y(_abc_41356_new_n7503_));
AND2X2 AND2X2_3637 ( .A(_abc_41356_new_n7454_), .B(_abc_41356_new_n7503_), .Y(_abc_41356_new_n7504_));
AND2X2 AND2X2_3638 ( .A(_abc_41356_new_n7341_), .B(_abc_41356_new_n7504_), .Y(_abc_41356_new_n7505_));
AND2X2 AND2X2_3639 ( .A(_abc_41356_new_n7505_), .B(_abc_41356_new_n7445_), .Y(_abc_41356_new_n7506_));
AND2X2 AND2X2_364 ( .A(_abc_41356_new_n718_), .B(\data[7] ), .Y(_abc_41356_new_n1184_));
AND2X2 AND2X2_3640 ( .A(_abc_41356_new_n7506_), .B(_abc_41356_new_n7495_), .Y(_abc_41356_new_n7507_));
AND2X2 AND2X2_3641 ( .A(_abc_41356_new_n7507_), .B(_abc_41356_new_n7415_), .Y(_abc_41356_new_n7508_));
AND2X2 AND2X2_3642 ( .A(_abc_41356_new_n7363_), .B(_abc_41356_new_n7352_), .Y(_abc_41356_new_n7510_));
AND2X2 AND2X2_3643 ( .A(_abc_41356_new_n7510_), .B(_abc_41356_new_n7422_), .Y(_abc_41356_new_n7511_));
AND2X2 AND2X2_3644 ( .A(_abc_41356_new_n7337_), .B(_abc_41356_new_n7253_), .Y(_abc_41356_new_n7515_));
AND2X2 AND2X2_3645 ( .A(_abc_41356_new_n7516_), .B(_abc_41356_new_n7514_), .Y(_abc_41356_new_n7517_));
AND2X2 AND2X2_3646 ( .A(_abc_41356_new_n7461_), .B(_abc_41356_new_n7518_), .Y(_abc_41356_new_n7519_));
AND2X2 AND2X2_3647 ( .A(_abc_41356_new_n7491_), .B(_abc_41356_new_n7434_), .Y(_abc_41356_new_n7520_));
AND2X2 AND2X2_3648 ( .A(_abc_41356_new_n7520_), .B(_abc_41356_new_n7519_), .Y(_abc_41356_new_n7521_));
AND2X2 AND2X2_3649 ( .A(_abc_41356_new_n7517_), .B(_abc_41356_new_n7521_), .Y(_abc_41356_new_n7522_));
AND2X2 AND2X2_365 ( .A(_abc_41356_new_n530_), .B(opcode_4_), .Y(_abc_41356_new_n1188_));
AND2X2 AND2X2_3650 ( .A(_abc_41356_new_n7458_), .B(_abc_41356_new_n7406_), .Y(_abc_41356_new_n7523_));
AND2X2 AND2X2_3651 ( .A(_abc_41356_new_n7522_), .B(_abc_41356_new_n7523_), .Y(_abc_41356_new_n7524_));
AND2X2 AND2X2_3652 ( .A(_abc_41356_new_n7524_), .B(_abc_41356_new_n7511_), .Y(_abc_41356_new_n7525_));
AND2X2 AND2X2_3653 ( .A(_abc_41356_new_n3454_), .B(_abc_41356_new_n7483_), .Y(_abc_41356_new_n7527_));
AND2X2 AND2X2_3654 ( .A(_abc_41356_new_n7058_), .B(_abc_41356_new_n717_), .Y(_abc_41356_new_n7533_));
AND2X2 AND2X2_3655 ( .A(_abc_41356_new_n7359_), .B(_abc_41356_new_n7379_), .Y(_abc_41356_new_n7545_));
AND2X2 AND2X2_3656 ( .A(_abc_41356_new_n7548_), .B(_abc_41356_new_n3490_), .Y(_abc_41356_new_n7549_));
AND2X2 AND2X2_3657 ( .A(_abc_41356_new_n7337_), .B(_abc_41356_new_n7549_), .Y(_abc_41356_new_n7550_));
AND2X2 AND2X2_3658 ( .A(_abc_41356_new_n3345_), .B(ei), .Y(_abc_41356_new_n7554_));
AND2X2 AND2X2_3659 ( .A(_abc_41356_new_n7556_), .B(_abc_41356_new_n7554_), .Y(_abc_41356_new_n7557_));
AND2X2 AND2X2_366 ( .A(_abc_41356_new_n1188_), .B(carry), .Y(_abc_41356_new_n1189_));
AND2X2 AND2X2_3660 ( .A(_abc_41356_new_n7558_), .B(ei), .Y(_abc_41356_new_n7559_));
AND2X2 AND2X2_3661 ( .A(_abc_41356_new_n3205_), .B(_abc_41356_new_n7560_), .Y(_abc_41356_new_n7561_));
AND2X2 AND2X2_3662 ( .A(alu_oprb_7_), .B(alu_opra_7_), .Y(alu__abc_40887_new_n34_));
AND2X2 AND2X2_3663 ( .A(alu__abc_40887_new_n35_), .B(alu__abc_40887_new_n33_), .Y(alu__abc_40887_new_n36_));
AND2X2 AND2X2_3664 ( .A(alu_oprb_6_), .B(alu_opra_6_), .Y(alu__abc_40887_new_n38_));
AND2X2 AND2X2_3665 ( .A(alu__abc_40887_new_n40_), .B(alu__abc_40887_new_n41_), .Y(alu__abc_40887_new_n42_));
AND2X2 AND2X2_3666 ( .A(alu__abc_40887_new_n43_), .B(alu__abc_40887_new_n39_), .Y(alu__abc_40887_new_n44_));
AND2X2 AND2X2_3667 ( .A(alu_oprb_1_), .B(alu_opra_1_), .Y(alu__abc_40887_new_n46_));
AND2X2 AND2X2_3668 ( .A(alu__abc_40887_new_n47_), .B(alu__abc_40887_new_n48_), .Y(alu__abc_40887_new_n49_));
AND2X2 AND2X2_3669 ( .A(alu_oprb_0_), .B(alu_opra_0_), .Y(alu__abc_40887_new_n50_));
AND2X2 AND2X2_367 ( .A(_abc_41356_new_n1109_), .B(_abc_41356_new_n1117_), .Y(_abc_41356_new_n1191_));
AND2X2 AND2X2_3670 ( .A(alu__abc_40887_new_n49_), .B(alu__abc_40887_new_n50_), .Y(alu__abc_40887_new_n51_));
AND2X2 AND2X2_3671 ( .A(alu_oprb_2_), .B(alu_opra_2_), .Y(alu__abc_40887_new_n53_));
AND2X2 AND2X2_3672 ( .A(alu__abc_40887_new_n55_), .B(alu__abc_40887_new_n56_), .Y(alu__abc_40887_new_n57_));
AND2X2 AND2X2_3673 ( .A(alu__abc_40887_new_n58_), .B(alu__abc_40887_new_n54_), .Y(alu__abc_40887_new_n59_));
AND2X2 AND2X2_3674 ( .A(alu_oprb_3_), .B(alu_opra_3_), .Y(alu__abc_40887_new_n60_));
AND2X2 AND2X2_3675 ( .A(alu__abc_40887_new_n61_), .B(alu__abc_40887_new_n62_), .Y(alu__abc_40887_new_n63_));
AND2X2 AND2X2_3676 ( .A(alu__abc_40887_new_n59_), .B(alu__abc_40887_new_n63_), .Y(alu__abc_40887_new_n64_));
AND2X2 AND2X2_3677 ( .A(alu__abc_40887_new_n52_), .B(alu__abc_40887_new_n64_), .Y(alu__abc_40887_new_n65_));
AND2X2 AND2X2_3678 ( .A(alu__abc_40887_new_n63_), .B(alu__abc_40887_new_n53_), .Y(alu__abc_40887_new_n66_));
AND2X2 AND2X2_3679 ( .A(alu_oprb_4_), .B(alu_opra_4_), .Y(alu__abc_40887_new_n69_));
AND2X2 AND2X2_368 ( .A(_abc_41356_new_n1193_), .B(_abc_41356_new_n698_), .Y(_abc_41356_new_n1194_));
AND2X2 AND2X2_3680 ( .A(alu__abc_40887_new_n71_), .B(alu__abc_40887_new_n72_), .Y(alu__abc_40887_new_n73_));
AND2X2 AND2X2_3681 ( .A(alu__abc_40887_new_n74_), .B(alu__abc_40887_new_n70_), .Y(alu__abc_40887_new_n75_));
AND2X2 AND2X2_3682 ( .A(alu__abc_40887_new_n76_), .B(alu__abc_40887_new_n77_), .Y(alu__abc_40887_new_n78_));
AND2X2 AND2X2_3683 ( .A(alu_oprb_5_), .B(alu_opra_5_), .Y(alu__abc_40887_new_n80_));
AND2X2 AND2X2_3684 ( .A(alu__abc_40887_new_n79_), .B(alu__abc_40887_new_n81_), .Y(alu__abc_40887_new_n82_));
AND2X2 AND2X2_3685 ( .A(alu__abc_40887_new_n75_), .B(alu__abc_40887_new_n82_), .Y(alu__abc_40887_new_n83_));
AND2X2 AND2X2_3686 ( .A(alu__abc_40887_new_n68_), .B(alu__abc_40887_new_n83_), .Y(alu__abc_40887_new_n84_));
AND2X2 AND2X2_3687 ( .A(alu__abc_40887_new_n82_), .B(alu__abc_40887_new_n69_), .Y(alu__abc_40887_new_n86_));
AND2X2 AND2X2_3688 ( .A(alu__abc_40887_new_n87_), .B(alu__abc_40887_new_n81_), .Y(alu__abc_40887_new_n88_));
AND2X2 AND2X2_3689 ( .A(alu__abc_40887_new_n85_), .B(alu__abc_40887_new_n88_), .Y(alu__abc_40887_new_n89_));
AND2X2 AND2X2_369 ( .A(_abc_41356_new_n1194_), .B(_abc_41356_new_n1192_), .Y(_abc_41356_new_n1195_));
AND2X2 AND2X2_3690 ( .A(alu__abc_40887_new_n90_), .B(alu__abc_40887_new_n39_), .Y(alu__abc_40887_new_n91_));
AND2X2 AND2X2_3691 ( .A(alu__abc_40887_new_n92_), .B(alu__abc_40887_new_n37_), .Y(alu__abc_40887_new_n93_));
AND2X2 AND2X2_3692 ( .A(alu__abc_40887_new_n91_), .B(alu__abc_40887_new_n36_), .Y(alu__abc_40887_new_n94_));
AND2X2 AND2X2_3693 ( .A(alu__abc_40887_new_n89_), .B(alu__abc_40887_new_n45_), .Y(alu__abc_40887_new_n98_));
AND2X2 AND2X2_3694 ( .A(alu__abc_40887_new_n68_), .B(alu__abc_40887_new_n75_), .Y(alu__abc_40887_new_n101_));
AND2X2 AND2X2_3695 ( .A(alu__abc_40887_new_n103_), .B(alu__abc_40887_new_n70_), .Y(alu__abc_40887_new_n104_));
AND2X2 AND2X2_3696 ( .A(alu__abc_40887_new_n102_), .B(alu__abc_40887_new_n104_), .Y(alu__abc_40887_new_n105_));
AND2X2 AND2X2_3697 ( .A(alu__abc_40887_new_n85_), .B(alu__abc_40887_new_n87_), .Y(alu__abc_40887_new_n107_));
AND2X2 AND2X2_3698 ( .A(alu__abc_40887_new_n106_), .B(alu__abc_40887_new_n107_), .Y(alu__abc_40887_new_n108_));
AND2X2 AND2X2_3699 ( .A(alu__abc_40887_new_n52_), .B(alu__abc_40887_new_n59_), .Y(alu__abc_40887_new_n109_));
AND2X2 AND2X2_37 ( .A(_abc_41356_new_n534_), .B(regfil_7__7_), .Y(_abc_41356_new_n557_));
AND2X2 AND2X2_370 ( .A(_abc_41356_new_n555_), .B(regfil_7__6_), .Y(_abc_41356_new_n1196_));
AND2X2 AND2X2_3700 ( .A(alu__abc_40887_new_n110_), .B(alu__abc_40887_new_n63_), .Y(alu__abc_40887_new_n111_));
AND2X2 AND2X2_3701 ( .A(alu__abc_40887_new_n112_), .B(alu__abc_40887_new_n113_), .Y(alu__abc_40887_new_n114_));
AND2X2 AND2X2_3702 ( .A(alu__abc_40887_new_n116_), .B(alu__abc_40887_new_n117_), .Y(alu__abc_40887_new_n118_));
AND2X2 AND2X2_3703 ( .A(alu__abc_40887_new_n119_), .B(alu__abc_40887_new_n115_), .Y(alu__abc_40887_new_n120_));
AND2X2 AND2X2_3704 ( .A(alu__abc_40887_new_n120_), .B(alu_cin), .Y(alu__abc_40887_new_n121_));
AND2X2 AND2X2_3705 ( .A(alu__abc_40887_new_n121_), .B(alu__abc_40887_new_n49_), .Y(alu__abc_40887_new_n122_));
AND2X2 AND2X2_3706 ( .A(alu__abc_40887_new_n123_), .B(alu__abc_40887_new_n124_), .Y(alu__abc_40887_new_n125_));
AND2X2 AND2X2_3707 ( .A(alu__abc_40887_new_n125_), .B(alu__abc_40887_new_n122_), .Y(alu__abc_40887_new_n126_));
AND2X2 AND2X2_3708 ( .A(alu__abc_40887_new_n114_), .B(alu__abc_40887_new_n126_), .Y(alu__abc_40887_new_n127_));
AND2X2 AND2X2_3709 ( .A(alu__abc_40887_new_n102_), .B(alu__abc_40887_new_n128_), .Y(alu__abc_40887_new_n129_));
AND2X2 AND2X2_371 ( .A(_abc_41356_new_n530_), .B(_abc_41356_new_n534_), .Y(_abc_41356_new_n1197_));
AND2X2 AND2X2_3710 ( .A(alu__abc_40887_new_n127_), .B(alu__abc_40887_new_n129_), .Y(alu__abc_40887_new_n130_));
AND2X2 AND2X2_3711 ( .A(alu__abc_40887_new_n130_), .B(alu__abc_40887_new_n108_), .Y(alu__abc_40887_new_n131_));
AND2X2 AND2X2_3712 ( .A(alu__abc_40887_new_n100_), .B(alu__abc_40887_new_n131_), .Y(alu__abc_40887_new_n132_));
AND2X2 AND2X2_3713 ( .A(alu__abc_40887_new_n96_), .B(alu__abc_40887_new_n133_), .Y(alu__abc_40887_new_n134_));
AND2X2 AND2X2_3714 ( .A(alu__abc_40887_new_n136_), .B(alu_sel_0_), .Y(alu__abc_40887_new_n137_));
AND2X2 AND2X2_3715 ( .A(alu__abc_40887_new_n137_), .B(alu__abc_40887_new_n135_), .Y(alu__abc_40887_new_n138_));
AND2X2 AND2X2_3716 ( .A(alu__abc_40887_new_n95_), .B(alu__abc_40887_new_n132_), .Y(alu__abc_40887_new_n140_));
AND2X2 AND2X2_3717 ( .A(alu_sel_1_), .B(alu_sel_0_), .Y(alu__abc_40887_new_n144_));
AND2X2 AND2X2_3718 ( .A(alu__abc_40887_new_n144_), .B(alu__abc_40887_new_n135_), .Y(alu__abc_40887_new_n145_));
AND2X2 AND2X2_3719 ( .A(alu__abc_40887_new_n146_), .B(alu_opra_3_), .Y(alu__abc_40887_new_n147_));
AND2X2 AND2X2_372 ( .A(_abc_41356_new_n1197_), .B(_abc_41356_new_n533_), .Y(_abc_41356_new_n1201_));
AND2X2 AND2X2_3720 ( .A(alu__abc_40887_new_n55_), .B(alu_opra_2_), .Y(alu__abc_40887_new_n149_));
AND2X2 AND2X2_3721 ( .A(alu__abc_40887_new_n148_), .B(alu__abc_40887_new_n149_), .Y(alu__abc_40887_new_n150_));
AND2X2 AND2X2_3722 ( .A(alu__abc_40887_new_n153_), .B(alu_opra_1_), .Y(alu__abc_40887_new_n154_));
AND2X2 AND2X2_3723 ( .A(alu__abc_40887_new_n117_), .B(alu_oprb_0_), .Y(alu__abc_40887_new_n156_));
AND2X2 AND2X2_3724 ( .A(alu__abc_40887_new_n157_), .B(alu__abc_40887_new_n155_), .Y(alu__abc_40887_new_n158_));
AND2X2 AND2X2_3725 ( .A(alu__abc_40887_new_n152_), .B(alu__abc_40887_new_n160_), .Y(alu__abc_40887_new_n161_));
AND2X2 AND2X2_3726 ( .A(alu__abc_40887_new_n71_), .B(alu_opra_4_), .Y(alu__abc_40887_new_n164_));
AND2X2 AND2X2_3727 ( .A(alu__abc_40887_new_n103_), .B(alu__abc_40887_new_n164_), .Y(alu__abc_40887_new_n165_));
AND2X2 AND2X2_3728 ( .A(alu__abc_40887_new_n76_), .B(alu_opra_5_), .Y(alu__abc_40887_new_n166_));
AND2X2 AND2X2_3729 ( .A(alu__abc_40887_new_n163_), .B(alu__abc_40887_new_n168_), .Y(alu__abc_40887_new_n169_));
AND2X2 AND2X2_373 ( .A(_abc_41356_new_n1202_), .B(_abc_41356_new_n1200_), .Y(_abc_41356_new_n1203_));
AND2X2 AND2X2_3730 ( .A(alu__abc_40887_new_n40_), .B(alu_opra_6_), .Y(alu__abc_40887_new_n171_));
AND2X2 AND2X2_3731 ( .A(alu__abc_40887_new_n170_), .B(alu__abc_40887_new_n172_), .Y(alu__abc_40887_new_n173_));
AND2X2 AND2X2_3732 ( .A(alu__abc_40887_new_n173_), .B(alu__abc_40887_new_n36_), .Y(alu__abc_40887_new_n175_));
AND2X2 AND2X2_3733 ( .A(alu__abc_40887_new_n176_), .B(alu__abc_40887_new_n174_), .Y(alu__abc_40887_new_n177_));
AND2X2 AND2X2_3734 ( .A(alu__abc_40887_new_n169_), .B(alu__abc_40887_new_n44_), .Y(alu__abc_40887_new_n179_));
AND2X2 AND2X2_3735 ( .A(alu__abc_40887_new_n180_), .B(alu__abc_40887_new_n170_), .Y(alu__abc_40887_new_n181_));
AND2X2 AND2X2_3736 ( .A(alu__abc_40887_new_n153_), .B(alu__abc_40887_new_n184_), .Y(alu__abc_40887_new_n185_));
AND2X2 AND2X2_3737 ( .A(alu__abc_40887_new_n186_), .B(alu__abc_40887_new_n187_), .Y(alu__abc_40887_new_n188_));
AND2X2 AND2X2_3738 ( .A(alu__abc_40887_new_n190_), .B(alu__abc_40887_new_n148_), .Y(alu__abc_40887_new_n191_));
AND2X2 AND2X2_3739 ( .A(alu__abc_40887_new_n189_), .B(alu__abc_40887_new_n191_), .Y(alu__abc_40887_new_n192_));
AND2X2 AND2X2_374 ( .A(_abc_41356_new_n1199_), .B(_abc_41356_new_n1203_), .Y(_abc_41356_new_n1204_));
AND2X2 AND2X2_3740 ( .A(alu__abc_40887_new_n193_), .B(alu__abc_40887_new_n183_), .Y(alu__abc_40887_new_n194_));
AND2X2 AND2X2_3741 ( .A(alu__abc_40887_new_n163_), .B(alu__abc_40887_new_n197_), .Y(alu__abc_40887_new_n198_));
AND2X2 AND2X2_3742 ( .A(alu__abc_40887_new_n196_), .B(alu__abc_40887_new_n198_), .Y(alu__abc_40887_new_n199_));
AND2X2 AND2X2_3743 ( .A(alu__abc_40887_new_n161_), .B(alu__abc_40887_new_n75_), .Y(alu__abc_40887_new_n201_));
AND2X2 AND2X2_3744 ( .A(alu__abc_40887_new_n189_), .B(alu__abc_40887_new_n190_), .Y(alu__abc_40887_new_n203_));
AND2X2 AND2X2_3745 ( .A(alu__abc_40887_new_n204_), .B(alu__abc_40887_new_n148_), .Y(alu__abc_40887_new_n205_));
AND2X2 AND2X2_3746 ( .A(alu__abc_40887_new_n206_), .B(alu__abc_40887_new_n207_), .Y(alu__abc_40887_new_n208_));
AND2X2 AND2X2_3747 ( .A(alu__abc_40887_new_n208_), .B(alu__abc_40887_new_n63_), .Y(alu__abc_40887_new_n209_));
AND2X2 AND2X2_3748 ( .A(alu__abc_40887_new_n158_), .B(alu__abc_40887_new_n59_), .Y(alu__abc_40887_new_n211_));
AND2X2 AND2X2_3749 ( .A(alu__abc_40887_new_n49_), .B(alu__abc_40887_new_n156_), .Y(alu__abc_40887_new_n215_));
AND2X2 AND2X2_375 ( .A(_abc_41356_new_n604_), .B(_abc_41356_new_n672_), .Y(_abc_41356_new_n1207_));
AND2X2 AND2X2_3750 ( .A(alu__abc_40887_new_n219_), .B(alu__abc_40887_new_n212_), .Y(alu__abc_40887_new_n220_));
AND2X2 AND2X2_3751 ( .A(alu__abc_40887_new_n210_), .B(alu__abc_40887_new_n220_), .Y(alu__abc_40887_new_n221_));
AND2X2 AND2X2_3752 ( .A(alu__abc_40887_new_n221_), .B(alu__abc_40887_new_n202_), .Y(alu__abc_40887_new_n222_));
AND2X2 AND2X2_3753 ( .A(alu__abc_40887_new_n222_), .B(alu__abc_40887_new_n200_), .Y(alu__abc_40887_new_n223_));
AND2X2 AND2X2_3754 ( .A(alu__abc_40887_new_n182_), .B(alu__abc_40887_new_n223_), .Y(alu__abc_40887_new_n224_));
AND2X2 AND2X2_3755 ( .A(alu__abc_40887_new_n178_), .B(alu__abc_40887_new_n224_), .Y(alu__abc_40887_new_n225_));
AND2X2 AND2X2_3756 ( .A(alu__abc_40887_new_n226_), .B(alu__abc_40887_new_n177_), .Y(alu__abc_40887_new_n227_));
AND2X2 AND2X2_3757 ( .A(alu__abc_40887_new_n228_), .B(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n229_));
AND2X2 AND2X2_3758 ( .A(alu__abc_40887_new_n136_), .B(alu__abc_40887_new_n230_), .Y(alu__abc_40887_new_n231_));
AND2X2 AND2X2_3759 ( .A(alu__abc_40887_new_n231_), .B(alu__abc_40887_new_n135_), .Y(alu__abc_40887_new_n232_));
AND2X2 AND2X2_376 ( .A(_abc_41356_new_n1208_), .B(_abc_41356_new_n668_), .Y(_abc_41356_new_n1209_));
AND2X2 AND2X2_3760 ( .A(alu__abc_40887_new_n95_), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n233_));
AND2X2 AND2X2_3761 ( .A(alu__abc_40887_new_n230_), .B(alu_sel_1_), .Y(alu__abc_40887_new_n234_));
AND2X2 AND2X2_3762 ( .A(alu__abc_40887_new_n234_), .B(alu__abc_40887_new_n135_), .Y(alu__abc_40887_new_n235_));
AND2X2 AND2X2_3763 ( .A(alu__abc_40887_new_n144_), .B(alu_sel_2_), .Y(alu__abc_40887_new_n236_));
AND2X2 AND2X2_3764 ( .A(alu__abc_40887_new_n177_), .B(alu__abc_40887_new_n237_), .Y(alu__abc_40887_new_n238_));
AND2X2 AND2X2_3765 ( .A(alu__abc_40887_new_n234_), .B(alu_sel_2_), .Y(alu__abc_40887_new_n239_));
AND2X2 AND2X2_3766 ( .A(alu__abc_40887_new_n239_), .B(alu__abc_40887_new_n33_), .Y(alu__abc_40887_new_n240_));
AND2X2 AND2X2_3767 ( .A(alu__abc_40887_new_n231_), .B(alu_sel_2_), .Y(alu__abc_40887_new_n241_));
AND2X2 AND2X2_3768 ( .A(alu__abc_40887_new_n241_), .B(alu__abc_40887_new_n34_), .Y(alu__abc_40887_new_n242_));
AND2X2 AND2X2_3769 ( .A(alu__abc_40887_new_n137_), .B(alu_sel_2_), .Y(alu__abc_40887_new_n243_));
AND2X2 AND2X2_377 ( .A(_abc_41356_new_n688_), .B(_abc_41356_new_n1210_), .Y(_abc_41356_new_n1211_));
AND2X2 AND2X2_3770 ( .A(alu__abc_40887_new_n36_), .B(alu__abc_40887_new_n243_), .Y(alu__abc_40887_new_n244_));
AND2X2 AND2X2_3771 ( .A(alu__abc_40887_new_n251_), .B(alu__abc_40887_new_n99_), .Y(alu__abc_40887_new_n252_));
AND2X2 AND2X2_3772 ( .A(alu__abc_40887_new_n133_), .B(alu__abc_40887_new_n138_), .Y(alu__abc_40887_new_n254_));
AND2X2 AND2X2_3773 ( .A(alu__abc_40887_new_n254_), .B(alu__abc_40887_new_n253_), .Y(alu__abc_40887_new_n255_));
AND2X2 AND2X2_3774 ( .A(alu__abc_40887_new_n257_), .B(alu__abc_40887_new_n256_), .Y(alu__abc_40887_new_n258_));
AND2X2 AND2X2_3775 ( .A(alu__abc_40887_new_n263_), .B(alu__abc_40887_new_n181_), .Y(alu__abc_40887_new_n264_));
AND2X2 AND2X2_3776 ( .A(alu__abc_40887_new_n265_), .B(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n266_));
AND2X2 AND2X2_3777 ( .A(alu__abc_40887_new_n100_), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n267_));
AND2X2 AND2X2_3778 ( .A(alu__abc_40887_new_n181_), .B(alu__abc_40887_new_n237_), .Y(alu__abc_40887_new_n268_));
AND2X2 AND2X2_3779 ( .A(alu__abc_40887_new_n44_), .B(alu__abc_40887_new_n243_), .Y(alu__abc_40887_new_n269_));
AND2X2 AND2X2_378 ( .A(_abc_41356_new_n1211_), .B(_abc_41356_new_n1209_), .Y(_abc_41356_new_n1212_));
AND2X2 AND2X2_3780 ( .A(alu__abc_40887_new_n239_), .B(alu__abc_40887_new_n43_), .Y(alu__abc_40887_new_n270_));
AND2X2 AND2X2_3781 ( .A(alu__abc_40887_new_n241_), .B(alu__abc_40887_new_n38_), .Y(alu__abc_40887_new_n271_));
AND2X2 AND2X2_3782 ( .A(alu__abc_40887_new_n281_), .B(alu__abc_40887_new_n280_), .Y(alu__abc_40887_new_n282_));
AND2X2 AND2X2_3783 ( .A(alu__abc_40887_new_n284_), .B(alu__abc_40887_new_n283_), .Y(alu__abc_40887_new_n285_));
AND2X2 AND2X2_3784 ( .A(alu__abc_40887_new_n285_), .B(alu__abc_40887_new_n142_), .Y(alu__abc_40887_new_n286_));
AND2X2 AND2X2_3785 ( .A(alu__abc_40887_new_n278_), .B(alu__abc_40887_new_n288_), .Y(alu__abc_40887_new_n289_));
AND2X2 AND2X2_3786 ( .A(alu__abc_40887_new_n186_), .B(alu__abc_40887_new_n115_), .Y(alu__abc_40887_new_n290_));
AND2X2 AND2X2_3787 ( .A(alu__abc_40887_new_n291_), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n292_));
AND2X2 AND2X2_3788 ( .A(alu__abc_40887_new_n217_), .B(alu__abc_40887_new_n214_), .Y(alu__abc_40887_new_n294_));
AND2X2 AND2X2_3789 ( .A(alu__abc_40887_new_n295_), .B(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n296_));
AND2X2 AND2X2_379 ( .A(_abc_41356_new_n599_), .B(_abc_41356_new_n535_), .Y(_abc_41356_new_n1215_));
AND2X2 AND2X2_3790 ( .A(alu__abc_40887_new_n291_), .B(alu__abc_40887_new_n297_), .Y(alu__abc_40887_new_n298_));
AND2X2 AND2X2_3791 ( .A(alu__abc_40887_new_n300_), .B(alu__abc_40887_new_n138_), .Y(alu__abc_40887_new_n301_));
AND2X2 AND2X2_3792 ( .A(alu__abc_40887_new_n301_), .B(alu__abc_40887_new_n299_), .Y(alu__abc_40887_new_n302_));
AND2X2 AND2X2_3793 ( .A(alu__abc_40887_new_n217_), .B(alu__abc_40887_new_n237_), .Y(alu__abc_40887_new_n303_));
AND2X2 AND2X2_3794 ( .A(alu__abc_40887_new_n49_), .B(alu__abc_40887_new_n243_), .Y(alu__abc_40887_new_n304_));
AND2X2 AND2X2_3795 ( .A(alu__abc_40887_new_n239_), .B(alu__abc_40887_new_n48_), .Y(alu__abc_40887_new_n305_));
AND2X2 AND2X2_3796 ( .A(alu__abc_40887_new_n231_), .B(alu__abc_40887_new_n46_), .Y(alu__abc_40887_new_n306_));
AND2X2 AND2X2_3797 ( .A(alu__abc_40887_new_n312_), .B(alu__abc_40887_new_n293_), .Y(alu__abc_40887_new_n313_));
AND2X2 AND2X2_3798 ( .A(alu__abc_40887_new_n317_), .B(alu__abc_40887_new_n316_), .Y(alu__abc_40887_new_n318_));
AND2X2 AND2X2_3799 ( .A(alu__abc_40887_new_n315_), .B(alu__abc_40887_new_n318_), .Y(alu__abc_40887_new_n319_));
AND2X2 AND2X2_38 ( .A(_abc_41356_new_n555_), .B(_abc_41356_new_n558_), .Y(_abc_41356_new_n559_));
AND2X2 AND2X2_380 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n1215_), .Y(_abc_41356_new_n1216_));
AND2X2 AND2X2_3800 ( .A(alu__abc_40887_new_n314_), .B(alu__abc_40887_new_n213_), .Y(alu__abc_40887_new_n321_));
AND2X2 AND2X2_3801 ( .A(alu__abc_40887_new_n139_), .B(alu__abc_40887_new_n279_), .Y(alu__abc_40887_new_n322_));
AND2X2 AND2X2_3802 ( .A(alu__abc_40887_new_n241_), .B(alu__abc_40887_new_n50_), .Y(alu__abc_40887_new_n325_));
AND2X2 AND2X2_3803 ( .A(alu__abc_40887_new_n239_), .B(alu__abc_40887_new_n119_), .Y(alu__abc_40887_new_n326_));
AND2X2 AND2X2_3804 ( .A(alu__abc_40887_new_n324_), .B(alu__abc_40887_new_n328_), .Y(alu__abc_40887_new_n329_));
AND2X2 AND2X2_3805 ( .A(alu__abc_40887_new_n329_), .B(alu__abc_40887_new_n320_), .Y(alu__abc_40887_new_n330_));
AND2X2 AND2X2_3806 ( .A(alu__abc_40887_new_n313_), .B(alu__abc_40887_new_n331_), .Y(alu__abc_40887_new_n332_));
AND2X2 AND2X2_3807 ( .A(alu__abc_40887_new_n338_), .B(alu__abc_40887_new_n339_), .Y(alu__abc_40887_new_n340_));
AND2X2 AND2X2_3808 ( .A(alu__abc_40887_new_n342_), .B(alu__abc_40887_new_n138_), .Y(alu__abc_40887_new_n343_));
AND2X2 AND2X2_3809 ( .A(alu__abc_40887_new_n343_), .B(alu__abc_40887_new_n341_), .Y(alu__abc_40887_new_n344_));
AND2X2 AND2X2_381 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n535_), .Y(_abc_41356_new_n1218_));
AND2X2 AND2X2_3810 ( .A(alu__abc_40887_new_n258_), .B(alu__abc_40887_new_n259_), .Y(alu__abc_40887_new_n345_));
AND2X2 AND2X2_3811 ( .A(alu__abc_40887_new_n346_), .B(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n347_));
AND2X2 AND2X2_3812 ( .A(alu__abc_40887_new_n114_), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n348_));
AND2X2 AND2X2_3813 ( .A(alu__abc_40887_new_n258_), .B(alu__abc_40887_new_n237_), .Y(alu__abc_40887_new_n349_));
AND2X2 AND2X2_3814 ( .A(alu__abc_40887_new_n63_), .B(alu__abc_40887_new_n243_), .Y(alu__abc_40887_new_n350_));
AND2X2 AND2X2_3815 ( .A(alu__abc_40887_new_n241_), .B(alu__abc_40887_new_n60_), .Y(alu__abc_40887_new_n351_));
AND2X2 AND2X2_3816 ( .A(alu__abc_40887_new_n239_), .B(alu__abc_40887_new_n62_), .Y(alu__abc_40887_new_n352_));
AND2X2 AND2X2_3817 ( .A(alu__abc_40887_new_n359_), .B(alu__abc_40887_new_n218_), .Y(alu__abc_40887_new_n360_));
AND2X2 AND2X2_3818 ( .A(alu__abc_40887_new_n361_), .B(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n362_));
AND2X2 AND2X2_3819 ( .A(alu__abc_40887_new_n363_), .B(alu__abc_40887_new_n300_), .Y(alu__abc_40887_new_n364_));
AND2X2 AND2X2_382 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n1218_), .Y(_abc_41356_new_n1219_));
AND2X2 AND2X2_3820 ( .A(alu__abc_40887_new_n339_), .B(alu__abc_40887_new_n138_), .Y(alu__abc_40887_new_n366_));
AND2X2 AND2X2_3821 ( .A(alu__abc_40887_new_n366_), .B(alu__abc_40887_new_n365_), .Y(alu__abc_40887_new_n367_));
AND2X2 AND2X2_3822 ( .A(alu__abc_40887_new_n359_), .B(alu__abc_40887_new_n237_), .Y(alu__abc_40887_new_n368_));
AND2X2 AND2X2_3823 ( .A(alu__abc_40887_new_n125_), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n369_));
AND2X2 AND2X2_3824 ( .A(alu__abc_40887_new_n239_), .B(alu__abc_40887_new_n58_), .Y(alu__abc_40887_new_n370_));
AND2X2 AND2X2_3825 ( .A(alu__abc_40887_new_n241_), .B(alu__abc_40887_new_n53_), .Y(alu__abc_40887_new_n371_));
AND2X2 AND2X2_3826 ( .A(alu__abc_40887_new_n59_), .B(alu__abc_40887_new_n243_), .Y(alu__abc_40887_new_n372_));
AND2X2 AND2X2_3827 ( .A(alu__abc_40887_new_n358_), .B(alu__abc_40887_new_n378_), .Y(alu__abc_40887_new_n381_));
AND2X2 AND2X2_3828 ( .A(alu__abc_40887_new_n384_), .B(alu__abc_40887_new_n379_), .Y(alu__abc_40887_new_n385_));
AND2X2 AND2X2_3829 ( .A(alu__abc_40887_new_n383_), .B(alu__abc_40887_new_n386_), .Y(alu__abc_40887_new_n387_));
AND2X2 AND2X2_383 ( .A(_abc_41356_new_n1217_), .B(_abc_41356_new_n1220_), .Y(_abc_41356_new_n1221_));
AND2X2 AND2X2_3830 ( .A(alu__abc_40887_new_n393_), .B(alu__abc_40887_new_n199_), .Y(alu__abc_40887_new_n394_));
AND2X2 AND2X2_3831 ( .A(alu__abc_40887_new_n395_), .B(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n396_));
AND2X2 AND2X2_3832 ( .A(alu__abc_40887_new_n199_), .B(alu__abc_40887_new_n237_), .Y(alu__abc_40887_new_n397_));
AND2X2 AND2X2_3833 ( .A(alu__abc_40887_new_n82_), .B(alu__abc_40887_new_n243_), .Y(alu__abc_40887_new_n398_));
AND2X2 AND2X2_3834 ( .A(alu__abc_40887_new_n239_), .B(alu__abc_40887_new_n79_), .Y(alu__abc_40887_new_n399_));
AND2X2 AND2X2_3835 ( .A(alu__abc_40887_new_n241_), .B(alu__abc_40887_new_n80_), .Y(alu__abc_40887_new_n401_));
AND2X2 AND2X2_3836 ( .A(alu__abc_40887_new_n407_), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n408_));
AND2X2 AND2X2_3837 ( .A(alu__abc_40887_new_n406_), .B(alu__abc_40887_new_n409_), .Y(alu__abc_40887_new_n410_));
AND2X2 AND2X2_3838 ( .A(alu__abc_40887_new_n342_), .B(alu__abc_40887_new_n411_), .Y(alu__abc_40887_new_n412_));
AND2X2 AND2X2_3839 ( .A(alu__abc_40887_new_n260_), .B(alu__abc_40887_new_n261_), .Y(alu__abc_40887_new_n415_));
AND2X2 AND2X2_384 ( .A(_abc_41356_new_n521_), .B(_abc_41356_new_n605_), .Y(_abc_41356_new_n1222_));
AND2X2 AND2X2_3840 ( .A(alu__abc_40887_new_n416_), .B(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n417_));
AND2X2 AND2X2_3841 ( .A(alu__abc_40887_new_n129_), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n418_));
AND2X2 AND2X2_3842 ( .A(alu__abc_40887_new_n261_), .B(alu__abc_40887_new_n237_), .Y(alu__abc_40887_new_n419_));
AND2X2 AND2X2_3843 ( .A(alu__abc_40887_new_n75_), .B(alu__abc_40887_new_n243_), .Y(alu__abc_40887_new_n420_));
AND2X2 AND2X2_3844 ( .A(alu__abc_40887_new_n239_), .B(alu__abc_40887_new_n74_), .Y(alu__abc_40887_new_n421_));
AND2X2 AND2X2_3845 ( .A(alu__abc_40887_new_n241_), .B(alu__abc_40887_new_n69_), .Y(alu__abc_40887_new_n423_));
AND2X2 AND2X2_3846 ( .A(alu__abc_40887_new_n428_), .B(alu__abc_40887_new_n414_), .Y(alu__abc_40887_new_n429_));
AND2X2 AND2X2_3847 ( .A(alu__abc_40887_new_n410_), .B(alu__abc_40887_new_n430_), .Y(alu__abc_40887_new_n431_));
AND2X2 AND2X2_3848 ( .A(alu__abc_40887_new_n263_), .B(alu__abc_40887_new_n432_), .Y(alu__abc_40887_new_n433_));
AND2X2 AND2X2_3849 ( .A(alu__abc_40887_new_n434_), .B(alu__abc_40887_new_n435_), .Y(alu__abc_40887_new_n436_));
AND2X2 AND2X2_385 ( .A(_abc_41356_new_n519_), .B(_abc_41356_new_n1222_), .Y(_abc_41356_new_n1223_));
AND2X2 AND2X2_3850 ( .A(alu__abc_40887_new_n436_), .B(alu__abc_40887_new_n391_), .Y(alu__abc_40887_new_n437_));
AND2X2 AND2X2_3851 ( .A(alu__abc_40887_new_n438_), .B(alu__abc_40887_new_n429_), .Y(alu__abc_40887_new_n439_));
AND2X2 AND2X2_3852 ( .A(alu__abc_40887_new_n442_), .B(alu__abc_40887_new_n443_), .Y(alu__abc_40887_new_n444_));
AND2X2 AND2X2_3853 ( .A(alu__abc_40887_new_n446_), .B(alu__abc_40887_new_n445_), .Y(alu__abc_40887_new_n447_));
AND2X2 AND2X2_3854 ( .A(alu__abc_40887_new_n441_), .B(alu__abc_40887_new_n448_), .Y(alu__abc_40887_new_n449_));
AND2X2 AND2X2_3855 ( .A(alu__abc_40887_new_n449_), .B(alu__abc_40887_new_n289_), .Y(alu__abc_40887_new_n450_));
AND2X2 AND2X2_3856 ( .A(alu__abc_40887_new_n286_), .B(alu__abc_40887_new_n287_), .Y(alu__abc_40887_new_n451_));
AND2X2 AND2X2_3857 ( .A(alu_sout), .B(alu__abc_40887_new_n277_), .Y(alu__abc_40887_new_n452_));
AND2X2 AND2X2_3858 ( .A(alu__abc_40887_new_n447_), .B(alu__abc_40887_new_n444_), .Y(alu__abc_40887_new_n454_));
AND2X2 AND2X2_3859 ( .A(alu__abc_40887_new_n440_), .B(alu__abc_40887_new_n387_), .Y(alu__abc_40887_new_n455_));
AND2X2 AND2X2_386 ( .A(_abc_41356_new_n509_), .B(_abc_41356_new_n590_), .Y(_abc_41356_new_n1224_));
AND2X2 AND2X2_3860 ( .A(alu__abc_40887_new_n456_), .B(alu__abc_40887_new_n453_), .Y(alu__abc_40887_new_n457_));
AND2X2 AND2X2_3861 ( .A(alu__abc_40887_new_n380_), .B(alu__abc_40887_new_n334_), .Y(alu__abc_40887_new_n459_));
AND2X2 AND2X2_3862 ( .A(alu__abc_40887_new_n439_), .B(alu__abc_40887_new_n459_), .Y(alu__abc_40887_new_n460_));
AND2X2 AND2X2_3863 ( .A(alu__abc_40887_new_n451_), .B(alu__abc_40887_new_n460_), .Y(alu_zout));
AND2X2 AND2X2_3864 ( .A(alu__abc_40887_new_n331_), .B(alu__abc_40887_new_n462_), .Y(alu__abc_40887_new_n463_));
AND2X2 AND2X2_3865 ( .A(alu__abc_40887_new_n236_), .B(alu_opra_0_), .Y(alu__abc_40887_new_n464_));
AND2X2 AND2X2_3866 ( .A(alu__abc_40887_new_n313_), .B(alu__abc_40887_new_n462_), .Y(alu__abc_40887_new_n466_));
AND2X2 AND2X2_3867 ( .A(alu__abc_40887_new_n236_), .B(alu_opra_1_), .Y(alu__abc_40887_new_n467_));
AND2X2 AND2X2_3868 ( .A(alu__abc_40887_new_n236_), .B(alu_opra_2_), .Y(alu__abc_40887_new_n469_));
AND2X2 AND2X2_3869 ( .A(alu__abc_40887_new_n378_), .B(alu__abc_40887_new_n462_), .Y(alu__abc_40887_new_n470_));
AND2X2 AND2X2_387 ( .A(_abc_41356_new_n1224_), .B(popdes_1_), .Y(_abc_41356_new_n1225_));
AND2X2 AND2X2_3870 ( .A(alu__abc_40887_new_n236_), .B(alu_opra_3_), .Y(alu__abc_40887_new_n472_));
AND2X2 AND2X2_3871 ( .A(alu__abc_40887_new_n358_), .B(alu__abc_40887_new_n462_), .Y(alu__abc_40887_new_n473_));
AND2X2 AND2X2_3872 ( .A(alu__abc_40887_new_n236_), .B(alu_opra_4_), .Y(alu__abc_40887_new_n475_));
AND2X2 AND2X2_3873 ( .A(alu__abc_40887_new_n430_), .B(alu__abc_40887_new_n462_), .Y(alu__abc_40887_new_n476_));
AND2X2 AND2X2_3874 ( .A(alu__abc_40887_new_n236_), .B(alu_opra_5_), .Y(alu__abc_40887_new_n478_));
AND2X2 AND2X2_3875 ( .A(alu__abc_40887_new_n410_), .B(alu__abc_40887_new_n462_), .Y(alu__abc_40887_new_n479_));
AND2X2 AND2X2_3876 ( .A(alu__abc_40887_new_n236_), .B(alu_opra_6_), .Y(alu__abc_40887_new_n481_));
AND2X2 AND2X2_3877 ( .A(alu__abc_40887_new_n277_), .B(alu__abc_40887_new_n462_), .Y(alu__abc_40887_new_n482_));
AND2X2 AND2X2_3878 ( .A(alu__abc_40887_new_n236_), .B(alu_opra_7_), .Y(alu__abc_40887_new_n484_));
AND2X2 AND2X2_3879 ( .A(alu_sout), .B(alu__abc_40887_new_n462_), .Y(alu__abc_40887_new_n485_));
AND2X2 AND2X2_388 ( .A(_abc_41356_new_n508_), .B(_abc_41356_new_n1225_), .Y(_abc_41356_new_n1226_));
AND2X2 AND2X2_3880 ( .A(alu__abc_40887_new_n174_), .B(alu__abc_40887_new_n488_), .Y(alu__abc_40887_new_n489_));
AND2X2 AND2X2_3881 ( .A(alu__abc_40887_new_n225_), .B(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n490_));
AND2X2 AND2X2_3882 ( .A(alu__abc_40887_new_n491_), .B(alu__abc_40887_new_n492_), .Y(alu__abc_40887_new_n493_));
AND2X2 AND2X2_3883 ( .A(alu__abc_40887_new_n140_), .B(alu__abc_40887_new_n138_), .Y(alu__abc_40887_new_n494_));
AND2X2 AND2X2_3884 ( .A(alu__abc_40887_new_n92_), .B(alu__abc_40887_new_n33_), .Y(alu__abc_40887_new_n495_));
AND2X2 AND2X2_3885 ( .A(alu__abc_40887_new_n135_), .B(alu__abc_40887_new_n136_), .Y(alu__abc_40887_new_n497_));
AND2X2 AND2X2_3886 ( .A(alu__abc_40887_new_n496_), .B(alu__abc_40887_new_n497_), .Y(alu__abc_40887_new_n498_));
AND2X2 AND2X2_389 ( .A(_abc_41356_new_n587_), .B(_abc_41356_new_n707_), .Y(_abc_41356_new_n1227_));
AND2X2 AND2X2_39 ( .A(_abc_41356_new_n561_), .B(_abc_41356_new_n532_), .Y(_abc_41356_new_n562_));
AND2X2 AND2X2_390 ( .A(_abc_41356_new_n519_), .B(_abc_41356_new_n1227_), .Y(_abc_41356_new_n1228_));
AND2X2 AND2X2_391 ( .A(opcode_6_), .B(opcode_7_), .Y(_abc_41356_new_n1232_));
AND2X2 AND2X2_392 ( .A(_abc_41356_new_n1232_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n1233_));
AND2X2 AND2X2_393 ( .A(_abc_41356_new_n676_), .B(_abc_41356_new_n1233_), .Y(_abc_41356_new_n1234_));
AND2X2 AND2X2_394 ( .A(_abc_41356_new_n1234_), .B(_abc_41356_new_n1215_), .Y(_abc_41356_new_n1235_));
AND2X2 AND2X2_395 ( .A(_abc_41356_new_n598_), .B(_abc_41356_new_n616_), .Y(_abc_41356_new_n1237_));
AND2X2 AND2X2_396 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n1237_), .Y(_abc_41356_new_n1238_));
AND2X2 AND2X2_397 ( .A(_abc_41356_new_n1239_), .B(_abc_41356_new_n1236_), .Y(_abc_41356_new_n1240_));
AND2X2 AND2X2_398 ( .A(_abc_41356_new_n1231_), .B(_abc_41356_new_n1240_), .Y(_abc_41356_new_n1241_));
AND2X2 AND2X2_399 ( .A(_abc_41356_new_n1241_), .B(_abc_41356_new_n1221_), .Y(_abc_41356_new_n1242_));
AND2X2 AND2X2_4 ( .A(_abc_41356_new_n504_), .B(_abc_41356_new_n506_), .Y(_abc_41356_new_n507_));
AND2X2 AND2X2_40 ( .A(_abc_41356_new_n512_), .B(_abc_41356_new_n564_), .Y(_abc_41356_new_n565_));
AND2X2 AND2X2_400 ( .A(_abc_41356_new_n1243_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n1244_));
AND2X2 AND2X2_401 ( .A(_abc_41356_new_n1214_), .B(_abc_41356_new_n1244_), .Y(_abc_41356_new_n1245_));
AND2X2 AND2X2_402 ( .A(_abc_41356_new_n1230_), .B(rdatahold_0_), .Y(_abc_41356_new_n1246_));
AND2X2 AND2X2_403 ( .A(_abc_41356_new_n1249_), .B(_abc_41356_new_n1248_), .Y(_abc_41356_new_n1250_));
AND2X2 AND2X2_404 ( .A(_abc_41356_new_n1258_), .B(_abc_41356_new_n1259_), .Y(_abc_41356_new_n1260_));
AND2X2 AND2X2_405 ( .A(_abc_41356_new_n1260_), .B(_abc_41356_new_n1257_), .Y(_abc_41356_new_n1261_));
AND2X2 AND2X2_406 ( .A(_abc_41356_new_n1261_), .B(_abc_41356_new_n1256_), .Y(_abc_41356_new_n1262_));
AND2X2 AND2X2_407 ( .A(_abc_41356_new_n1262_), .B(_abc_41356_new_n1255_), .Y(_abc_41356_new_n1263_));
AND2X2 AND2X2_408 ( .A(_abc_41356_new_n1263_), .B(_abc_41356_new_n1254_), .Y(_abc_41356_new_n1264_));
AND2X2 AND2X2_409 ( .A(_abc_41356_new_n1264_), .B(_abc_41356_new_n1253_), .Y(_abc_41356_new_n1265_));
AND2X2 AND2X2_41 ( .A(_abc_41356_new_n563_), .B(_abc_41356_new_n566_), .Y(_abc_41356_new_n567_));
AND2X2 AND2X2_410 ( .A(_abc_41356_new_n1265_), .B(_abc_41356_new_n1252_), .Y(_abc_41356_new_n1266_));
AND2X2 AND2X2_411 ( .A(_abc_41356_new_n1266_), .B(_abc_41356_new_n1251_), .Y(_abc_41356_new_n1267_));
AND2X2 AND2X2_412 ( .A(_abc_41356_new_n1269_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n1270_));
AND2X2 AND2X2_413 ( .A(_abc_41356_new_n1270_), .B(_abc_41356_new_n1268_), .Y(_abc_41356_new_n1271_));
AND2X2 AND2X2_414 ( .A(regfil_5__0_), .B(regfil_5__1_), .Y(_abc_41356_new_n1273_));
AND2X2 AND2X2_415 ( .A(_abc_41356_new_n1273_), .B(regfil_5__2_), .Y(_abc_41356_new_n1274_));
AND2X2 AND2X2_416 ( .A(_abc_41356_new_n1274_), .B(regfil_5__3_), .Y(_abc_41356_new_n1275_));
AND2X2 AND2X2_417 ( .A(regfil_5__7_), .B(regfil_5__6_), .Y(_abc_41356_new_n1276_));
AND2X2 AND2X2_418 ( .A(regfil_5__5_), .B(regfil_5__4_), .Y(_abc_41356_new_n1277_));
AND2X2 AND2X2_419 ( .A(_abc_41356_new_n1276_), .B(_abc_41356_new_n1277_), .Y(_abc_41356_new_n1278_));
AND2X2 AND2X2_42 ( .A(regfil_1__0_), .B(regfil_1__1_), .Y(_abc_41356_new_n568_));
AND2X2 AND2X2_420 ( .A(_abc_41356_new_n1275_), .B(_abc_41356_new_n1278_), .Y(_abc_41356_new_n1279_));
AND2X2 AND2X2_421 ( .A(_abc_41356_new_n1279_), .B(regfil_4__0_), .Y(_abc_41356_new_n1281_));
AND2X2 AND2X2_422 ( .A(_abc_41356_new_n1282_), .B(_abc_41356_new_n1280_), .Y(_abc_41356_new_n1283_));
AND2X2 AND2X2_423 ( .A(_abc_41356_new_n1237_), .B(_abc_41356_new_n681_), .Y(_abc_41356_new_n1286_));
AND2X2 AND2X2_424 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n1286_), .Y(_abc_41356_new_n1287_));
AND2X2 AND2X2_425 ( .A(regfil_5__1_), .B(sp_1_), .Y(_abc_41356_new_n1288_));
AND2X2 AND2X2_426 ( .A(_abc_41356_new_n1289_), .B(_abc_41356_new_n1290_), .Y(_abc_41356_new_n1291_));
AND2X2 AND2X2_427 ( .A(regfil_5__0_), .B(sp_0_), .Y(_abc_41356_new_n1292_));
AND2X2 AND2X2_428 ( .A(_abc_41356_new_n1291_), .B(_abc_41356_new_n1292_), .Y(_abc_41356_new_n1293_));
AND2X2 AND2X2_429 ( .A(_abc_41356_new_n1294_), .B(_abc_41356_new_n1289_), .Y(_abc_41356_new_n1295_));
AND2X2 AND2X2_43 ( .A(_abc_41356_new_n568_), .B(regfil_1__2_), .Y(_abc_41356_new_n569_));
AND2X2 AND2X2_430 ( .A(regfil_5__2_), .B(sp_2_), .Y(_abc_41356_new_n1297_));
AND2X2 AND2X2_431 ( .A(_abc_41356_new_n1257_), .B(_abc_41356_new_n1298_), .Y(_abc_41356_new_n1299_));
AND2X2 AND2X2_432 ( .A(regfil_5__3_), .B(sp_3_), .Y(_abc_41356_new_n1302_));
AND2X2 AND2X2_433 ( .A(_abc_41356_new_n1256_), .B(_abc_41356_new_n1303_), .Y(_abc_41356_new_n1304_));
AND2X2 AND2X2_434 ( .A(_abc_41356_new_n1301_), .B(_abc_41356_new_n1306_), .Y(_abc_41356_new_n1307_));
AND2X2 AND2X2_435 ( .A(_abc_41356_new_n1296_), .B(_abc_41356_new_n1307_), .Y(_abc_41356_new_n1308_));
AND2X2 AND2X2_436 ( .A(_abc_41356_new_n1306_), .B(_abc_41356_new_n1297_), .Y(_abc_41356_new_n1309_));
AND2X2 AND2X2_437 ( .A(regfil_5__7_), .B(sp_7_), .Y(_abc_41356_new_n1312_));
AND2X2 AND2X2_438 ( .A(_abc_41356_new_n1252_), .B(_abc_41356_new_n1314_), .Y(_abc_41356_new_n1315_));
AND2X2 AND2X2_439 ( .A(_abc_41356_new_n1316_), .B(_abc_41356_new_n1313_), .Y(_abc_41356_new_n1317_));
AND2X2 AND2X2_44 ( .A(_abc_41356_new_n569_), .B(regfil_1__3_), .Y(_abc_41356_new_n570_));
AND2X2 AND2X2_440 ( .A(regfil_5__6_), .B(sp_6_), .Y(_abc_41356_new_n1318_));
AND2X2 AND2X2_441 ( .A(_abc_41356_new_n1253_), .B(_abc_41356_new_n1319_), .Y(_abc_41356_new_n1320_));
AND2X2 AND2X2_442 ( .A(_abc_41356_new_n1322_), .B(_abc_41356_new_n1317_), .Y(_abc_41356_new_n1323_));
AND2X2 AND2X2_443 ( .A(regfil_5__4_), .B(sp_4_), .Y(_abc_41356_new_n1324_));
AND2X2 AND2X2_444 ( .A(_abc_41356_new_n1255_), .B(_abc_41356_new_n1325_), .Y(_abc_41356_new_n1326_));
AND2X2 AND2X2_445 ( .A(regfil_5__5_), .B(sp_5_), .Y(_abc_41356_new_n1329_));
AND2X2 AND2X2_446 ( .A(_abc_41356_new_n1254_), .B(_abc_41356_new_n1331_), .Y(_abc_41356_new_n1332_));
AND2X2 AND2X2_447 ( .A(_abc_41356_new_n1333_), .B(_abc_41356_new_n1330_), .Y(_abc_41356_new_n1334_));
AND2X2 AND2X2_448 ( .A(_abc_41356_new_n1328_), .B(_abc_41356_new_n1334_), .Y(_abc_41356_new_n1335_));
AND2X2 AND2X2_449 ( .A(_abc_41356_new_n1323_), .B(_abc_41356_new_n1335_), .Y(_abc_41356_new_n1336_));
AND2X2 AND2X2_45 ( .A(_abc_41356_new_n570_), .B(regfil_1__4_), .Y(_abc_41356_new_n571_));
AND2X2 AND2X2_450 ( .A(_abc_41356_new_n1311_), .B(_abc_41356_new_n1336_), .Y(_abc_41356_new_n1337_));
AND2X2 AND2X2_451 ( .A(_abc_41356_new_n1316_), .B(_abc_41356_new_n1318_), .Y(_abc_41356_new_n1338_));
AND2X2 AND2X2_452 ( .A(_abc_41356_new_n1334_), .B(_abc_41356_new_n1324_), .Y(_abc_41356_new_n1340_));
AND2X2 AND2X2_453 ( .A(_abc_41356_new_n1341_), .B(_abc_41356_new_n1323_), .Y(_abc_41356_new_n1342_));
AND2X2 AND2X2_454 ( .A(_abc_41356_new_n1251_), .B(_abc_41356_new_n1345_), .Y(_abc_41356_new_n1346_));
AND2X2 AND2X2_455 ( .A(regfil_4__0_), .B(sp_8_), .Y(_abc_41356_new_n1347_));
AND2X2 AND2X2_456 ( .A(_abc_41356_new_n1344_), .B(_abc_41356_new_n1349_), .Y(_abc_41356_new_n1350_));
AND2X2 AND2X2_457 ( .A(_abc_41356_new_n1351_), .B(_abc_41356_new_n1352_), .Y(_abc_41356_new_n1353_));
AND2X2 AND2X2_458 ( .A(_abc_41356_new_n1353_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n1354_));
AND2X2 AND2X2_459 ( .A(regfil_5__3_), .B(regfil_3__3_), .Y(_abc_41356_new_n1355_));
AND2X2 AND2X2_46 ( .A(_abc_41356_new_n571_), .B(regfil_1__5_), .Y(_abc_41356_new_n572_));
AND2X2 AND2X2_460 ( .A(_abc_41356_new_n1256_), .B(_abc_41356_new_n1356_), .Y(_abc_41356_new_n1357_));
AND2X2 AND2X2_461 ( .A(regfil_5__2_), .B(regfil_3__2_), .Y(_abc_41356_new_n1360_));
AND2X2 AND2X2_462 ( .A(_abc_41356_new_n1359_), .B(_abc_41356_new_n1360_), .Y(_abc_41356_new_n1361_));
AND2X2 AND2X2_463 ( .A(regfil_5__1_), .B(regfil_3__1_), .Y(_abc_41356_new_n1363_));
AND2X2 AND2X2_464 ( .A(regfil_3__0_), .B(regfil_5__0_), .Y(_abc_41356_new_n1364_));
AND2X2 AND2X2_465 ( .A(_abc_41356_new_n1365_), .B(_abc_41356_new_n1366_), .Y(_abc_41356_new_n1367_));
AND2X2 AND2X2_466 ( .A(_abc_41356_new_n1367_), .B(_abc_41356_new_n1364_), .Y(_abc_41356_new_n1368_));
AND2X2 AND2X2_467 ( .A(_abc_41356_new_n1257_), .B(_abc_41356_new_n1370_), .Y(_abc_41356_new_n1371_));
AND2X2 AND2X2_468 ( .A(_abc_41356_new_n1359_), .B(_abc_41356_new_n1373_), .Y(_abc_41356_new_n1374_));
AND2X2 AND2X2_469 ( .A(_abc_41356_new_n1369_), .B(_abc_41356_new_n1374_), .Y(_abc_41356_new_n1375_));
AND2X2 AND2X2_47 ( .A(_abc_41356_new_n572_), .B(regfil_1__6_), .Y(_abc_41356_new_n573_));
AND2X2 AND2X2_470 ( .A(regfil_5__7_), .B(regfil_3__7_), .Y(_abc_41356_new_n1377_));
AND2X2 AND2X2_471 ( .A(_abc_41356_new_n1378_), .B(_abc_41356_new_n1379_), .Y(_abc_41356_new_n1380_));
AND2X2 AND2X2_472 ( .A(regfil_5__6_), .B(regfil_3__6_), .Y(_abc_41356_new_n1381_));
AND2X2 AND2X2_473 ( .A(_abc_41356_new_n1382_), .B(_abc_41356_new_n1383_), .Y(_abc_41356_new_n1384_));
AND2X2 AND2X2_474 ( .A(_abc_41356_new_n1380_), .B(_abc_41356_new_n1384_), .Y(_abc_41356_new_n1385_));
AND2X2 AND2X2_475 ( .A(regfil_5__5_), .B(regfil_3__5_), .Y(_abc_41356_new_n1386_));
AND2X2 AND2X2_476 ( .A(_abc_41356_new_n1387_), .B(_abc_41356_new_n1388_), .Y(_abc_41356_new_n1389_));
AND2X2 AND2X2_477 ( .A(regfil_5__4_), .B(regfil_3__4_), .Y(_abc_41356_new_n1390_));
AND2X2 AND2X2_478 ( .A(_abc_41356_new_n1391_), .B(_abc_41356_new_n1392_), .Y(_abc_41356_new_n1393_));
AND2X2 AND2X2_479 ( .A(_abc_41356_new_n1389_), .B(_abc_41356_new_n1393_), .Y(_abc_41356_new_n1394_));
AND2X2 AND2X2_48 ( .A(_abc_41356_new_n573_), .B(regfil_1__7_), .Y(_abc_41356_new_n574_));
AND2X2 AND2X2_480 ( .A(_abc_41356_new_n1385_), .B(_abc_41356_new_n1394_), .Y(_abc_41356_new_n1395_));
AND2X2 AND2X2_481 ( .A(_abc_41356_new_n1376_), .B(_abc_41356_new_n1395_), .Y(_abc_41356_new_n1396_));
AND2X2 AND2X2_482 ( .A(_abc_41356_new_n1397_), .B(_abc_41356_new_n1388_), .Y(_abc_41356_new_n1398_));
AND2X2 AND2X2_483 ( .A(_abc_41356_new_n1385_), .B(_abc_41356_new_n1398_), .Y(_abc_41356_new_n1399_));
AND2X2 AND2X2_484 ( .A(_abc_41356_new_n1379_), .B(_abc_41356_new_n1381_), .Y(_abc_41356_new_n1400_));
AND2X2 AND2X2_485 ( .A(_abc_41356_new_n1405_), .B(_abc_41356_new_n1251_), .Y(_abc_41356_new_n1406_));
AND2X2 AND2X2_486 ( .A(regfil_2__0_), .B(regfil_4__0_), .Y(_abc_41356_new_n1407_));
AND2X2 AND2X2_487 ( .A(_abc_41356_new_n1409_), .B(_abc_41356_new_n1411_), .Y(_abc_41356_new_n1412_));
AND2X2 AND2X2_488 ( .A(_abc_41356_new_n525_), .B(opcode_4_), .Y(_abc_41356_new_n1413_));
AND2X2 AND2X2_489 ( .A(_abc_41356_new_n1237_), .B(_abc_41356_new_n1413_), .Y(_abc_41356_new_n1414_));
AND2X2 AND2X2_49 ( .A(_abc_41356_new_n534_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n576_));
AND2X2 AND2X2_490 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n1414_), .Y(_abc_41356_new_n1415_));
AND2X2 AND2X2_491 ( .A(_abc_41356_new_n1412_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n1416_));
AND2X2 AND2X2_492 ( .A(_abc_41356_new_n1237_), .B(_abc_41356_new_n535_), .Y(_abc_41356_new_n1417_));
AND2X2 AND2X2_493 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n1417_), .Y(_abc_41356_new_n1418_));
AND2X2 AND2X2_494 ( .A(regfil_1__1_), .B(regfil_5__1_), .Y(_abc_41356_new_n1419_));
AND2X2 AND2X2_495 ( .A(regfil_1__0_), .B(regfil_5__0_), .Y(_abc_41356_new_n1421_));
AND2X2 AND2X2_496 ( .A(_abc_41356_new_n648_), .B(_abc_41356_new_n1259_), .Y(_abc_41356_new_n1423_));
AND2X2 AND2X2_497 ( .A(_abc_41356_new_n1425_), .B(_abc_41356_new_n1420_), .Y(_abc_41356_new_n1426_));
AND2X2 AND2X2_498 ( .A(regfil_1__3_), .B(regfil_5__3_), .Y(_abc_41356_new_n1427_));
AND2X2 AND2X2_499 ( .A(_abc_41356_new_n645_), .B(_abc_41356_new_n1256_), .Y(_abc_41356_new_n1428_));
AND2X2 AND2X2_5 ( .A(_abc_41356_new_n507_), .B(_abc_41356_new_n502_), .Y(_abc_41356_new_n508_));
AND2X2 AND2X2_50 ( .A(_abc_41356_new_n545_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n578_));
AND2X2 AND2X2_500 ( .A(regfil_1__2_), .B(regfil_5__2_), .Y(_abc_41356_new_n1431_));
AND2X2 AND2X2_501 ( .A(_abc_41356_new_n646_), .B(_abc_41356_new_n1257_), .Y(_abc_41356_new_n1432_));
AND2X2 AND2X2_502 ( .A(_abc_41356_new_n1430_), .B(_abc_41356_new_n1434_), .Y(_abc_41356_new_n1435_));
AND2X2 AND2X2_503 ( .A(_abc_41356_new_n1438_), .B(_abc_41356_new_n1431_), .Y(_abc_41356_new_n1439_));
AND2X2 AND2X2_504 ( .A(_abc_41356_new_n1437_), .B(_abc_41356_new_n1441_), .Y(_abc_41356_new_n1442_));
AND2X2 AND2X2_505 ( .A(regfil_1__7_), .B(regfil_5__7_), .Y(_abc_41356_new_n1443_));
AND2X2 AND2X2_506 ( .A(_abc_41356_new_n1444_), .B(_abc_41356_new_n1445_), .Y(_abc_41356_new_n1446_));
AND2X2 AND2X2_507 ( .A(regfil_1__6_), .B(regfil_5__6_), .Y(_abc_41356_new_n1447_));
AND2X2 AND2X2_508 ( .A(_abc_41356_new_n1448_), .B(_abc_41356_new_n1449_), .Y(_abc_41356_new_n1450_));
AND2X2 AND2X2_509 ( .A(_abc_41356_new_n1446_), .B(_abc_41356_new_n1450_), .Y(_abc_41356_new_n1451_));
AND2X2 AND2X2_51 ( .A(_abc_41356_new_n578_), .B(_abc_41356_new_n526_), .Y(_abc_41356_new_n579_));
AND2X2 AND2X2_510 ( .A(regfil_1__4_), .B(regfil_5__4_), .Y(_abc_41356_new_n1452_));
AND2X2 AND2X2_511 ( .A(_abc_41356_new_n1453_), .B(_abc_41356_new_n1454_), .Y(_abc_41356_new_n1455_));
AND2X2 AND2X2_512 ( .A(regfil_1__5_), .B(regfil_5__5_), .Y(_abc_41356_new_n1456_));
AND2X2 AND2X2_513 ( .A(_abc_41356_new_n1457_), .B(_abc_41356_new_n1458_), .Y(_abc_41356_new_n1459_));
AND2X2 AND2X2_514 ( .A(_abc_41356_new_n1455_), .B(_abc_41356_new_n1459_), .Y(_abc_41356_new_n1460_));
AND2X2 AND2X2_515 ( .A(_abc_41356_new_n1451_), .B(_abc_41356_new_n1460_), .Y(_abc_41356_new_n1461_));
AND2X2 AND2X2_516 ( .A(_abc_41356_new_n1464_), .B(_abc_41356_new_n1458_), .Y(_abc_41356_new_n1465_));
AND2X2 AND2X2_517 ( .A(_abc_41356_new_n1451_), .B(_abc_41356_new_n1465_), .Y(_abc_41356_new_n1466_));
AND2X2 AND2X2_518 ( .A(_abc_41356_new_n1445_), .B(_abc_41356_new_n1447_), .Y(_abc_41356_new_n1467_));
AND2X2 AND2X2_519 ( .A(_abc_41356_new_n1463_), .B(_abc_41356_new_n1470_), .Y(_abc_41356_new_n1471_));
AND2X2 AND2X2_52 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n576_), .Y(_abc_41356_new_n580_));
AND2X2 AND2X2_520 ( .A(_abc_41356_new_n644_), .B(_abc_41356_new_n1251_), .Y(_abc_41356_new_n1473_));
AND2X2 AND2X2_521 ( .A(regfil_0__0_), .B(regfil_4__0_), .Y(_abc_41356_new_n1474_));
AND2X2 AND2X2_522 ( .A(_abc_41356_new_n1472_), .B(_abc_41356_new_n1476_), .Y(_abc_41356_new_n1477_));
AND2X2 AND2X2_523 ( .A(_abc_41356_new_n1478_), .B(_abc_41356_new_n1479_), .Y(_abc_41356_new_n1480_));
AND2X2 AND2X2_524 ( .A(_abc_41356_new_n1237_), .B(_abc_41356_new_n576_), .Y(_abc_41356_new_n1481_));
AND2X2 AND2X2_525 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n1481_), .Y(_abc_41356_new_n1482_));
AND2X2 AND2X2_526 ( .A(_abc_41356_new_n1480_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n1483_));
AND2X2 AND2X2_527 ( .A(_abc_41356_new_n1418_), .B(_abc_41356_new_n1252_), .Y(_abc_41356_new_n1486_));
AND2X2 AND2X2_528 ( .A(_abc_41356_new_n1485_), .B(_abc_41356_new_n1487_), .Y(_abc_41356_new_n1488_));
AND2X2 AND2X2_529 ( .A(_abc_41356_new_n1490_), .B(_abc_41356_new_n1284_), .Y(_abc_41356_new_n1491_));
AND2X2 AND2X2_53 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n580_), .Y(_abc_41356_new_n581_));
AND2X2 AND2X2_530 ( .A(_abc_41356_new_n1491_), .B(_abc_41356_new_n1272_), .Y(_abc_41356_new_n1492_));
AND2X2 AND2X2_531 ( .A(_abc_41356_new_n1493_), .B(_abc_41356_new_n1250_), .Y(_abc_41356_new_n1494_));
AND2X2 AND2X2_532 ( .A(_abc_41356_new_n1497_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n1498_));
AND2X2 AND2X2_533 ( .A(_abc_41356_new_n1496_), .B(_abc_41356_new_n1498_), .Y(_abc_41356_new_n1499_));
AND2X2 AND2X2_534 ( .A(_abc_41356_new_n1230_), .B(rdatahold_1_), .Y(_abc_41356_new_n1500_));
AND2X2 AND2X2_535 ( .A(_abc_41356_new_n1502_), .B(_abc_41356_new_n1248_), .Y(_abc_41356_new_n1503_));
AND2X2 AND2X2_536 ( .A(_abc_41356_new_n1267_), .B(_abc_41356_new_n1504_), .Y(_abc_41356_new_n1505_));
AND2X2 AND2X2_537 ( .A(_abc_41356_new_n1268_), .B(regfil_4__1_), .Y(_abc_41356_new_n1506_));
AND2X2 AND2X2_538 ( .A(_abc_41356_new_n1507_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n1508_));
AND2X2 AND2X2_539 ( .A(_abc_41356_new_n1281_), .B(regfil_4__1_), .Y(_abc_41356_new_n1511_));
AND2X2 AND2X2_54 ( .A(_abc_41356_new_n574_), .B(regfil_0__0_), .Y(_abc_41356_new_n582_));
AND2X2 AND2X2_540 ( .A(_abc_41356_new_n1512_), .B(_abc_41356_new_n1510_), .Y(_abc_41356_new_n1513_));
AND2X2 AND2X2_541 ( .A(_abc_41356_new_n1504_), .B(_abc_41356_new_n1515_), .Y(_abc_41356_new_n1516_));
AND2X2 AND2X2_542 ( .A(regfil_4__1_), .B(sp_9_), .Y(_abc_41356_new_n1517_));
AND2X2 AND2X2_543 ( .A(_abc_41356_new_n1349_), .B(_abc_41356_new_n1519_), .Y(_abc_41356_new_n1520_));
AND2X2 AND2X2_544 ( .A(_abc_41356_new_n1344_), .B(_abc_41356_new_n1520_), .Y(_abc_41356_new_n1521_));
AND2X2 AND2X2_545 ( .A(_abc_41356_new_n1524_), .B(_abc_41356_new_n1522_), .Y(_abc_41356_new_n1525_));
AND2X2 AND2X2_546 ( .A(_abc_41356_new_n1519_), .B(_abc_41356_new_n1347_), .Y(_abc_41356_new_n1526_));
AND2X2 AND2X2_547 ( .A(_abc_41356_new_n1287_), .B(_abc_41356_new_n1527_), .Y(_abc_41356_new_n1528_));
AND2X2 AND2X2_548 ( .A(_abc_41356_new_n1525_), .B(_abc_41356_new_n1528_), .Y(_abc_41356_new_n1529_));
AND2X2 AND2X2_549 ( .A(_abc_41356_new_n1403_), .B(_abc_41356_new_n1410_), .Y(_abc_41356_new_n1530_));
AND2X2 AND2X2_55 ( .A(_abc_41356_new_n583_), .B(_abc_41356_new_n581_), .Y(_abc_41356_new_n584_));
AND2X2 AND2X2_550 ( .A(regfil_2__1_), .B(regfil_4__1_), .Y(_abc_41356_new_n1531_));
AND2X2 AND2X2_551 ( .A(_abc_41356_new_n1532_), .B(_abc_41356_new_n1504_), .Y(_abc_41356_new_n1533_));
AND2X2 AND2X2_552 ( .A(_abc_41356_new_n1410_), .B(_abc_41356_new_n1535_), .Y(_abc_41356_new_n1538_));
AND2X2 AND2X2_553 ( .A(_abc_41356_new_n1403_), .B(_abc_41356_new_n1538_), .Y(_abc_41356_new_n1539_));
AND2X2 AND2X2_554 ( .A(_abc_41356_new_n1535_), .B(_abc_41356_new_n1407_), .Y(_abc_41356_new_n1541_));
AND2X2 AND2X2_555 ( .A(_abc_41356_new_n1540_), .B(_abc_41356_new_n1542_), .Y(_abc_41356_new_n1543_));
AND2X2 AND2X2_556 ( .A(_abc_41356_new_n1543_), .B(_abc_41356_new_n1537_), .Y(_abc_41356_new_n1544_));
AND2X2 AND2X2_557 ( .A(_abc_41356_new_n1544_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n1545_));
AND2X2 AND2X2_558 ( .A(_abc_41356_new_n1546_), .B(_abc_41356_new_n1504_), .Y(_abc_41356_new_n1547_));
AND2X2 AND2X2_559 ( .A(regfil_0__1_), .B(regfil_4__1_), .Y(_abc_41356_new_n1548_));
AND2X2 AND2X2_56 ( .A(_abc_41356_new_n584_), .B(_abc_41356_new_n575_), .Y(_abc_41356_new_n585_));
AND2X2 AND2X2_560 ( .A(_abc_41356_new_n1476_), .B(_abc_41356_new_n1550_), .Y(_abc_41356_new_n1551_));
AND2X2 AND2X2_561 ( .A(_abc_41356_new_n1550_), .B(_abc_41356_new_n1474_), .Y(_abc_41356_new_n1556_));
AND2X2 AND2X2_562 ( .A(_abc_41356_new_n1482_), .B(_abc_41356_new_n1557_), .Y(_abc_41356_new_n1558_));
AND2X2 AND2X2_563 ( .A(_abc_41356_new_n1555_), .B(_abc_41356_new_n1558_), .Y(_abc_41356_new_n1559_));
AND2X2 AND2X2_564 ( .A(_abc_41356_new_n1559_), .B(_abc_41356_new_n1553_), .Y(_abc_41356_new_n1560_));
AND2X2 AND2X2_565 ( .A(_abc_41356_new_n1418_), .B(_abc_41356_new_n1251_), .Y(_abc_41356_new_n1563_));
AND2X2 AND2X2_566 ( .A(_abc_41356_new_n1562_), .B(_abc_41356_new_n1564_), .Y(_abc_41356_new_n1565_));
AND2X2 AND2X2_567 ( .A(_abc_41356_new_n1567_), .B(_abc_41356_new_n1514_), .Y(_abc_41356_new_n1568_));
AND2X2 AND2X2_568 ( .A(_abc_41356_new_n1569_), .B(_abc_41356_new_n1503_), .Y(_abc_41356_new_n1570_));
AND2X2 AND2X2_569 ( .A(_abc_41356_new_n1573_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n1574_));
AND2X2 AND2X2_57 ( .A(_abc_41356_new_n586_), .B(state_3_), .Y(_abc_41356_new_n587_));
AND2X2 AND2X2_570 ( .A(_abc_41356_new_n1572_), .B(_abc_41356_new_n1574_), .Y(_abc_41356_new_n1575_));
AND2X2 AND2X2_571 ( .A(_abc_41356_new_n1230_), .B(rdatahold_2_), .Y(_abc_41356_new_n1576_));
AND2X2 AND2X2_572 ( .A(_abc_41356_new_n1578_), .B(_abc_41356_new_n1248_), .Y(_abc_41356_new_n1579_));
AND2X2 AND2X2_573 ( .A(_abc_41356_new_n1505_), .B(_abc_41356_new_n1580_), .Y(_abc_41356_new_n1581_));
AND2X2 AND2X2_574 ( .A(_abc_41356_new_n1583_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n1584_));
AND2X2 AND2X2_575 ( .A(_abc_41356_new_n1584_), .B(_abc_41356_new_n1582_), .Y(_abc_41356_new_n1585_));
AND2X2 AND2X2_576 ( .A(_abc_41356_new_n1511_), .B(regfil_4__2_), .Y(_abc_41356_new_n1588_));
AND2X2 AND2X2_577 ( .A(_abc_41356_new_n1589_), .B(_abc_41356_new_n1587_), .Y(_abc_41356_new_n1590_));
AND2X2 AND2X2_578 ( .A(_abc_41356_new_n1527_), .B(_abc_41356_new_n1592_), .Y(_abc_41356_new_n1593_));
AND2X2 AND2X2_579 ( .A(_abc_41356_new_n1522_), .B(_abc_41356_new_n1593_), .Y(_abc_41356_new_n1594_));
AND2X2 AND2X2_58 ( .A(_abc_41356_new_n521_), .B(_abc_41356_new_n587_), .Y(_abc_41356_new_n588_));
AND2X2 AND2X2_580 ( .A(_abc_41356_new_n1580_), .B(_abc_41356_new_n1596_), .Y(_abc_41356_new_n1597_));
AND2X2 AND2X2_581 ( .A(regfil_4__2_), .B(sp_10_), .Y(_abc_41356_new_n1598_));
AND2X2 AND2X2_582 ( .A(_abc_41356_new_n1595_), .B(_abc_41356_new_n1600_), .Y(_abc_41356_new_n1601_));
AND2X2 AND2X2_583 ( .A(_abc_41356_new_n1602_), .B(_abc_41356_new_n1603_), .Y(_abc_41356_new_n1604_));
AND2X2 AND2X2_584 ( .A(_abc_41356_new_n1604_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n1605_));
AND2X2 AND2X2_585 ( .A(_abc_41356_new_n1608_), .B(_abc_41356_new_n1580_), .Y(_abc_41356_new_n1609_));
AND2X2 AND2X2_586 ( .A(regfil_2__2_), .B(regfil_4__2_), .Y(_abc_41356_new_n1610_));
AND2X2 AND2X2_587 ( .A(_abc_41356_new_n1607_), .B(_abc_41356_new_n1612_), .Y(_abc_41356_new_n1613_));
AND2X2 AND2X2_588 ( .A(_abc_41356_new_n1614_), .B(_abc_41356_new_n1615_), .Y(_abc_41356_new_n1616_));
AND2X2 AND2X2_589 ( .A(_abc_41356_new_n1616_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n1617_));
AND2X2 AND2X2_59 ( .A(_abc_41356_new_n519_), .B(_abc_41356_new_n588_), .Y(_abc_41356_new_n589_));
AND2X2 AND2X2_590 ( .A(_abc_41356_new_n1553_), .B(_abc_41356_new_n1619_), .Y(_abc_41356_new_n1620_));
AND2X2 AND2X2_591 ( .A(_abc_41356_new_n1621_), .B(_abc_41356_new_n1580_), .Y(_abc_41356_new_n1622_));
AND2X2 AND2X2_592 ( .A(regfil_0__2_), .B(regfil_4__2_), .Y(_abc_41356_new_n1623_));
AND2X2 AND2X2_593 ( .A(_abc_41356_new_n1628_), .B(_abc_41356_new_n1625_), .Y(_abc_41356_new_n1629_));
AND2X2 AND2X2_594 ( .A(_abc_41356_new_n1629_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n1630_));
AND2X2 AND2X2_595 ( .A(_abc_41356_new_n1418_), .B(_abc_41356_new_n1504_), .Y(_abc_41356_new_n1633_));
AND2X2 AND2X2_596 ( .A(_abc_41356_new_n1632_), .B(_abc_41356_new_n1634_), .Y(_abc_41356_new_n1635_));
AND2X2 AND2X2_597 ( .A(_abc_41356_new_n1637_), .B(_abc_41356_new_n1591_), .Y(_abc_41356_new_n1638_));
AND2X2 AND2X2_598 ( .A(_abc_41356_new_n1638_), .B(_abc_41356_new_n1586_), .Y(_abc_41356_new_n1639_));
AND2X2 AND2X2_599 ( .A(_abc_41356_new_n1640_), .B(_abc_41356_new_n1579_), .Y(_abc_41356_new_n1641_));
AND2X2 AND2X2_6 ( .A(popdes_0_), .B(popdes_1_), .Y(_abc_41356_new_n510_));
AND2X2 AND2X2_60 ( .A(_abc_41356_new_n590_), .B(_abc_41356_new_n591_), .Y(_abc_41356_new_n592_));
AND2X2 AND2X2_600 ( .A(_abc_41356_new_n1644_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n1645_));
AND2X2 AND2X2_601 ( .A(_abc_41356_new_n1643_), .B(_abc_41356_new_n1645_), .Y(_abc_41356_new_n1646_));
AND2X2 AND2X2_602 ( .A(_abc_41356_new_n1230_), .B(rdatahold_3_), .Y(_abc_41356_new_n1647_));
AND2X2 AND2X2_603 ( .A(_abc_41356_new_n1649_), .B(_abc_41356_new_n1248_), .Y(_abc_41356_new_n1650_));
AND2X2 AND2X2_604 ( .A(_abc_41356_new_n1652_), .B(_abc_41356_new_n1653_), .Y(_abc_41356_new_n1654_));
AND2X2 AND2X2_605 ( .A(regfil_4__3_), .B(sp_11_), .Y(_abc_41356_new_n1656_));
AND2X2 AND2X2_606 ( .A(_abc_41356_new_n1655_), .B(_abc_41356_new_n1657_), .Y(_abc_41356_new_n1658_));
AND2X2 AND2X2_607 ( .A(_abc_41356_new_n1651_), .B(_abc_41356_new_n1659_), .Y(_abc_41356_new_n1660_));
AND2X2 AND2X2_608 ( .A(_abc_41356_new_n1661_), .B(_abc_41356_new_n1658_), .Y(_abc_41356_new_n1662_));
AND2X2 AND2X2_609 ( .A(_abc_41356_new_n1663_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n1664_));
AND2X2 AND2X2_61 ( .A(_abc_41356_new_n592_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n593_));
AND2X2 AND2X2_610 ( .A(regfil_2__3_), .B(regfil_4__3_), .Y(_abc_41356_new_n1667_));
AND2X2 AND2X2_611 ( .A(_abc_41356_new_n1669_), .B(_abc_41356_new_n1652_), .Y(_abc_41356_new_n1670_));
AND2X2 AND2X2_612 ( .A(_abc_41356_new_n1671_), .B(_abc_41356_new_n1668_), .Y(_abc_41356_new_n1672_));
AND2X2 AND2X2_613 ( .A(_abc_41356_new_n1676_), .B(_abc_41356_new_n1673_), .Y(_abc_41356_new_n1677_));
AND2X2 AND2X2_614 ( .A(_abc_41356_new_n1625_), .B(_abc_41356_new_n1679_), .Y(_abc_41356_new_n1680_));
AND2X2 AND2X2_615 ( .A(regfil_0__3_), .B(regfil_4__3_), .Y(_abc_41356_new_n1682_));
AND2X2 AND2X2_616 ( .A(_abc_41356_new_n1684_), .B(_abc_41356_new_n1652_), .Y(_abc_41356_new_n1685_));
AND2X2 AND2X2_617 ( .A(_abc_41356_new_n1686_), .B(_abc_41356_new_n1683_), .Y(_abc_41356_new_n1687_));
AND2X2 AND2X2_618 ( .A(_abc_41356_new_n1688_), .B(_abc_41356_new_n1690_), .Y(_abc_41356_new_n1691_));
AND2X2 AND2X2_619 ( .A(_abc_41356_new_n1691_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n1692_));
AND2X2 AND2X2_62 ( .A(_abc_41356_new_n508_), .B(_abc_41356_new_n593_), .Y(_abc_41356_new_n594_));
AND2X2 AND2X2_620 ( .A(_abc_41356_new_n1693_), .B(_abc_41356_new_n1678_), .Y(_abc_41356_new_n1694_));
AND2X2 AND2X2_621 ( .A(_abc_41356_new_n1418_), .B(regfil_4__2_), .Y(_abc_41356_new_n1695_));
AND2X2 AND2X2_622 ( .A(_abc_41356_new_n1588_), .B(regfil_4__3_), .Y(_abc_41356_new_n1699_));
AND2X2 AND2X2_623 ( .A(_abc_41356_new_n1700_), .B(_abc_41356_new_n1698_), .Y(_abc_41356_new_n1701_));
AND2X2 AND2X2_624 ( .A(_abc_41356_new_n1701_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n1702_));
AND2X2 AND2X2_625 ( .A(_abc_41356_new_n1582_), .B(regfil_4__3_), .Y(_abc_41356_new_n1705_));
AND2X2 AND2X2_626 ( .A(_abc_41356_new_n1581_), .B(_abc_41356_new_n1652_), .Y(_abc_41356_new_n1706_));
AND2X2 AND2X2_627 ( .A(_abc_41356_new_n1707_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n1708_));
AND2X2 AND2X2_628 ( .A(_abc_41356_new_n1704_), .B(_abc_41356_new_n1710_), .Y(_abc_41356_new_n1711_));
AND2X2 AND2X2_629 ( .A(_abc_41356_new_n1712_), .B(_abc_41356_new_n1650_), .Y(_abc_41356_new_n1713_));
AND2X2 AND2X2_63 ( .A(_abc_41356_new_n577_), .B(opcode_3_), .Y(_abc_41356_new_n598_));
AND2X2 AND2X2_630 ( .A(_abc_41356_new_n1716_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n1717_));
AND2X2 AND2X2_631 ( .A(_abc_41356_new_n1715_), .B(_abc_41356_new_n1717_), .Y(_abc_41356_new_n1718_));
AND2X2 AND2X2_632 ( .A(_abc_41356_new_n1230_), .B(rdatahold_4_), .Y(_abc_41356_new_n1719_));
AND2X2 AND2X2_633 ( .A(_abc_41356_new_n1721_), .B(_abc_41356_new_n1248_), .Y(_abc_41356_new_n1722_));
AND2X2 AND2X2_634 ( .A(_abc_41356_new_n1706_), .B(_abc_41356_new_n1723_), .Y(_abc_41356_new_n1724_));
AND2X2 AND2X2_635 ( .A(_abc_41356_new_n1707_), .B(regfil_4__4_), .Y(_abc_41356_new_n1725_));
AND2X2 AND2X2_636 ( .A(_abc_41356_new_n1726_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n1727_));
AND2X2 AND2X2_637 ( .A(_abc_41356_new_n1600_), .B(_abc_41356_new_n1658_), .Y(_abc_41356_new_n1729_));
AND2X2 AND2X2_638 ( .A(_abc_41356_new_n1520_), .B(_abc_41356_new_n1729_), .Y(_abc_41356_new_n1730_));
AND2X2 AND2X2_639 ( .A(_abc_41356_new_n1344_), .B(_abc_41356_new_n1730_), .Y(_abc_41356_new_n1731_));
AND2X2 AND2X2_64 ( .A(_abc_41356_new_n598_), .B(_abc_41356_new_n526_), .Y(_abc_41356_new_n599_));
AND2X2 AND2X2_640 ( .A(_abc_41356_new_n1732_), .B(_abc_41356_new_n1729_), .Y(_abc_41356_new_n1733_));
AND2X2 AND2X2_641 ( .A(_abc_41356_new_n1655_), .B(_abc_41356_new_n1598_), .Y(_abc_41356_new_n1734_));
AND2X2 AND2X2_642 ( .A(_abc_41356_new_n1723_), .B(_abc_41356_new_n1738_), .Y(_abc_41356_new_n1739_));
AND2X2 AND2X2_643 ( .A(regfil_4__4_), .B(sp_12_), .Y(_abc_41356_new_n1740_));
AND2X2 AND2X2_644 ( .A(_abc_41356_new_n1737_), .B(_abc_41356_new_n1742_), .Y(_abc_41356_new_n1743_));
AND2X2 AND2X2_645 ( .A(_abc_41356_new_n1744_), .B(_abc_41356_new_n1745_), .Y(_abc_41356_new_n1746_));
AND2X2 AND2X2_646 ( .A(_abc_41356_new_n1746_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n1747_));
AND2X2 AND2X2_647 ( .A(_abc_41356_new_n1748_), .B(_abc_41356_new_n1723_), .Y(_abc_41356_new_n1749_));
AND2X2 AND2X2_648 ( .A(regfil_0__4_), .B(regfil_4__4_), .Y(_abc_41356_new_n1750_));
AND2X2 AND2X2_649 ( .A(_abc_41356_new_n1686_), .B(_abc_41356_new_n1623_), .Y(_abc_41356_new_n1753_));
AND2X2 AND2X2_65 ( .A(_abc_41356_new_n599_), .B(_abc_41356_new_n576_), .Y(_abc_41356_new_n600_));
AND2X2 AND2X2_650 ( .A(_abc_41356_new_n1627_), .B(_abc_41356_new_n1687_), .Y(_abc_41356_new_n1755_));
AND2X2 AND2X2_651 ( .A(_abc_41356_new_n1618_), .B(_abc_41356_new_n1755_), .Y(_abc_41356_new_n1756_));
AND2X2 AND2X2_652 ( .A(_abc_41356_new_n1551_), .B(_abc_41356_new_n1755_), .Y(_abc_41356_new_n1759_));
AND2X2 AND2X2_653 ( .A(_abc_41356_new_n1761_), .B(_abc_41356_new_n1758_), .Y(_abc_41356_new_n1762_));
AND2X2 AND2X2_654 ( .A(_abc_41356_new_n1763_), .B(_abc_41356_new_n1752_), .Y(_abc_41356_new_n1764_));
AND2X2 AND2X2_655 ( .A(_abc_41356_new_n1765_), .B(_abc_41356_new_n1766_), .Y(_abc_41356_new_n1767_));
AND2X2 AND2X2_656 ( .A(_abc_41356_new_n1767_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n1768_));
AND2X2 AND2X2_657 ( .A(_abc_41356_new_n1612_), .B(_abc_41356_new_n1672_), .Y(_abc_41356_new_n1769_));
AND2X2 AND2X2_658 ( .A(_abc_41356_new_n1538_), .B(_abc_41356_new_n1769_), .Y(_abc_41356_new_n1770_));
AND2X2 AND2X2_659 ( .A(_abc_41356_new_n1403_), .B(_abc_41356_new_n1770_), .Y(_abc_41356_new_n1771_));
AND2X2 AND2X2_66 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n600_), .Y(_abc_41356_new_n601_));
AND2X2 AND2X2_660 ( .A(_abc_41356_new_n1606_), .B(_abc_41356_new_n1769_), .Y(_abc_41356_new_n1772_));
AND2X2 AND2X2_661 ( .A(_abc_41356_new_n1671_), .B(_abc_41356_new_n1610_), .Y(_abc_41356_new_n1773_));
AND2X2 AND2X2_662 ( .A(_abc_41356_new_n1777_), .B(_abc_41356_new_n1723_), .Y(_abc_41356_new_n1778_));
AND2X2 AND2X2_663 ( .A(regfil_2__4_), .B(regfil_4__4_), .Y(_abc_41356_new_n1779_));
AND2X2 AND2X2_664 ( .A(_abc_41356_new_n1776_), .B(_abc_41356_new_n1781_), .Y(_abc_41356_new_n1782_));
AND2X2 AND2X2_665 ( .A(_abc_41356_new_n1783_), .B(_abc_41356_new_n1784_), .Y(_abc_41356_new_n1785_));
AND2X2 AND2X2_666 ( .A(_abc_41356_new_n1785_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n1786_));
AND2X2 AND2X2_667 ( .A(_abc_41356_new_n1418_), .B(_abc_41356_new_n1652_), .Y(_abc_41356_new_n1789_));
AND2X2 AND2X2_668 ( .A(_abc_41356_new_n1788_), .B(_abc_41356_new_n1790_), .Y(_abc_41356_new_n1791_));
AND2X2 AND2X2_669 ( .A(_abc_41356_new_n1275_), .B(regfil_5__4_), .Y(_abc_41356_new_n1795_));
AND2X2 AND2X2_67 ( .A(_abc_41356_new_n597_), .B(_abc_41356_new_n602_), .Y(_abc_41356_new_n603_));
AND2X2 AND2X2_670 ( .A(_abc_41356_new_n1795_), .B(regfil_5__5_), .Y(_abc_41356_new_n1796_));
AND2X2 AND2X2_671 ( .A(_abc_41356_new_n1796_), .B(regfil_5__6_), .Y(_abc_41356_new_n1797_));
AND2X2 AND2X2_672 ( .A(_abc_41356_new_n1797_), .B(regfil_5__7_), .Y(_abc_41356_new_n1798_));
AND2X2 AND2X2_673 ( .A(_abc_41356_new_n1798_), .B(regfil_4__0_), .Y(_abc_41356_new_n1799_));
AND2X2 AND2X2_674 ( .A(_abc_41356_new_n1799_), .B(regfil_4__1_), .Y(_abc_41356_new_n1800_));
AND2X2 AND2X2_675 ( .A(_abc_41356_new_n1800_), .B(regfil_4__2_), .Y(_abc_41356_new_n1801_));
AND2X2 AND2X2_676 ( .A(_abc_41356_new_n1801_), .B(regfil_4__3_), .Y(_abc_41356_new_n1802_));
AND2X2 AND2X2_677 ( .A(_abc_41356_new_n1802_), .B(regfil_4__4_), .Y(_abc_41356_new_n1803_));
AND2X2 AND2X2_678 ( .A(_abc_41356_new_n1804_), .B(_abc_41356_new_n1794_), .Y(_abc_41356_new_n1805_));
AND2X2 AND2X2_679 ( .A(_abc_41356_new_n1793_), .B(_abc_41356_new_n1806_), .Y(_abc_41356_new_n1807_));
AND2X2 AND2X2_68 ( .A(_abc_41356_new_n603_), .B(_abc_41356_new_n596_), .Y(_abc_41356_new_n604_));
AND2X2 AND2X2_680 ( .A(_abc_41356_new_n1808_), .B(_abc_41356_new_n1722_), .Y(_abc_41356_new_n1809_));
AND2X2 AND2X2_681 ( .A(_abc_41356_new_n1812_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n1813_));
AND2X2 AND2X2_682 ( .A(_abc_41356_new_n1811_), .B(_abc_41356_new_n1813_), .Y(_abc_41356_new_n1814_));
AND2X2 AND2X2_683 ( .A(_abc_41356_new_n1230_), .B(rdatahold_5_), .Y(_abc_41356_new_n1815_));
AND2X2 AND2X2_684 ( .A(_abc_41356_new_n1817_), .B(_abc_41356_new_n1248_), .Y(_abc_41356_new_n1818_));
AND2X2 AND2X2_685 ( .A(_abc_41356_new_n1724_), .B(_abc_41356_new_n1819_), .Y(_abc_41356_new_n1820_));
AND2X2 AND2X2_686 ( .A(_abc_41356_new_n1821_), .B(regfil_4__5_), .Y(_abc_41356_new_n1822_));
AND2X2 AND2X2_687 ( .A(_abc_41356_new_n1823_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n1824_));
AND2X2 AND2X2_688 ( .A(_abc_41356_new_n1819_), .B(_abc_41356_new_n1826_), .Y(_abc_41356_new_n1827_));
AND2X2 AND2X2_689 ( .A(regfil_4__5_), .B(sp_13_), .Y(_abc_41356_new_n1828_));
AND2X2 AND2X2_69 ( .A(state_3_), .B(state_2_), .Y(_abc_41356_new_n605_));
AND2X2 AND2X2_690 ( .A(_abc_41356_new_n1830_), .B(_abc_41356_new_n1740_), .Y(_abc_41356_new_n1831_));
AND2X2 AND2X2_691 ( .A(_abc_41356_new_n1742_), .B(_abc_41356_new_n1830_), .Y(_abc_41356_new_n1835_));
AND2X2 AND2X2_692 ( .A(_abc_41356_new_n1737_), .B(_abc_41356_new_n1835_), .Y(_abc_41356_new_n1836_));
AND2X2 AND2X2_693 ( .A(_abc_41356_new_n1834_), .B(_abc_41356_new_n1837_), .Y(_abc_41356_new_n1838_));
AND2X2 AND2X2_694 ( .A(_abc_41356_new_n1838_), .B(_abc_41356_new_n1832_), .Y(_abc_41356_new_n1839_));
AND2X2 AND2X2_695 ( .A(_abc_41356_new_n1839_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n1840_));
AND2X2 AND2X2_696 ( .A(_abc_41356_new_n1418_), .B(regfil_4__4_), .Y(_abc_41356_new_n1841_));
AND2X2 AND2X2_697 ( .A(_abc_41356_new_n1842_), .B(_abc_41356_new_n1819_), .Y(_abc_41356_new_n1843_));
AND2X2 AND2X2_698 ( .A(regfil_2__5_), .B(regfil_4__5_), .Y(_abc_41356_new_n1844_));
AND2X2 AND2X2_699 ( .A(_abc_41356_new_n1781_), .B(_abc_41356_new_n1846_), .Y(_abc_41356_new_n1849_));
AND2X2 AND2X2_7 ( .A(_abc_41356_new_n510_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n511_));
AND2X2 AND2X2_70 ( .A(_abc_41356_new_n506_), .B(_abc_41356_new_n605_), .Y(_abc_41356_new_n606_));
AND2X2 AND2X2_700 ( .A(_abc_41356_new_n1776_), .B(_abc_41356_new_n1849_), .Y(_abc_41356_new_n1850_));
AND2X2 AND2X2_701 ( .A(_abc_41356_new_n1848_), .B(_abc_41356_new_n1851_), .Y(_abc_41356_new_n1852_));
AND2X2 AND2X2_702 ( .A(_abc_41356_new_n1846_), .B(_abc_41356_new_n1779_), .Y(_abc_41356_new_n1853_));
AND2X2 AND2X2_703 ( .A(_abc_41356_new_n1415_), .B(_abc_41356_new_n1854_), .Y(_abc_41356_new_n1855_));
AND2X2 AND2X2_704 ( .A(_abc_41356_new_n1852_), .B(_abc_41356_new_n1855_), .Y(_abc_41356_new_n1856_));
AND2X2 AND2X2_705 ( .A(_abc_41356_new_n1857_), .B(_abc_41356_new_n1819_), .Y(_abc_41356_new_n1858_));
AND2X2 AND2X2_706 ( .A(regfil_0__5_), .B(regfil_4__5_), .Y(_abc_41356_new_n1859_));
AND2X2 AND2X2_707 ( .A(_abc_41356_new_n1752_), .B(_abc_41356_new_n1861_), .Y(_abc_41356_new_n1862_));
AND2X2 AND2X2_708 ( .A(_abc_41356_new_n1861_), .B(_abc_41356_new_n1750_), .Y(_abc_41356_new_n1867_));
AND2X2 AND2X2_709 ( .A(_abc_41356_new_n1482_), .B(_abc_41356_new_n1868_), .Y(_abc_41356_new_n1869_));
AND2X2 AND2X2_71 ( .A(_abc_41356_new_n502_), .B(_abc_41356_new_n509_), .Y(_abc_41356_new_n607_));
AND2X2 AND2X2_710 ( .A(_abc_41356_new_n1866_), .B(_abc_41356_new_n1869_), .Y(_abc_41356_new_n1870_));
AND2X2 AND2X2_711 ( .A(_abc_41356_new_n1870_), .B(_abc_41356_new_n1864_), .Y(_abc_41356_new_n1871_));
AND2X2 AND2X2_712 ( .A(_abc_41356_new_n1803_), .B(regfil_4__5_), .Y(_abc_41356_new_n1877_));
AND2X2 AND2X2_713 ( .A(_abc_41356_new_n1878_), .B(_abc_41356_new_n1876_), .Y(_abc_41356_new_n1879_));
AND2X2 AND2X2_714 ( .A(_abc_41356_new_n1875_), .B(_abc_41356_new_n1880_), .Y(_abc_41356_new_n1881_));
AND2X2 AND2X2_715 ( .A(_abc_41356_new_n1882_), .B(_abc_41356_new_n1818_), .Y(_abc_41356_new_n1883_));
AND2X2 AND2X2_716 ( .A(_abc_41356_new_n1886_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n1887_));
AND2X2 AND2X2_717 ( .A(_abc_41356_new_n1885_), .B(_abc_41356_new_n1887_), .Y(_abc_41356_new_n1888_));
AND2X2 AND2X2_718 ( .A(_abc_41356_new_n1230_), .B(rdatahold_6_), .Y(_abc_41356_new_n1889_));
AND2X2 AND2X2_719 ( .A(_abc_41356_new_n1891_), .B(_abc_41356_new_n1248_), .Y(_abc_41356_new_n1892_));
AND2X2 AND2X2_72 ( .A(_abc_41356_new_n606_), .B(_abc_41356_new_n607_), .Y(_abc_41356_new_n608_));
AND2X2 AND2X2_720 ( .A(_abc_41356_new_n1820_), .B(_abc_41356_new_n1893_), .Y(_abc_41356_new_n1894_));
AND2X2 AND2X2_721 ( .A(_abc_41356_new_n1895_), .B(regfil_4__6_), .Y(_abc_41356_new_n1896_));
AND2X2 AND2X2_722 ( .A(_abc_41356_new_n1897_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n1898_));
AND2X2 AND2X2_723 ( .A(_abc_41356_new_n1893_), .B(_abc_41356_new_n1902_), .Y(_abc_41356_new_n1903_));
AND2X2 AND2X2_724 ( .A(regfil_4__6_), .B(sp_14_), .Y(_abc_41356_new_n1904_));
AND2X2 AND2X2_725 ( .A(_abc_41356_new_n1901_), .B(_abc_41356_new_n1906_), .Y(_abc_41356_new_n1908_));
AND2X2 AND2X2_726 ( .A(_abc_41356_new_n1909_), .B(_abc_41356_new_n1907_), .Y(_abc_41356_new_n1910_));
AND2X2 AND2X2_727 ( .A(_abc_41356_new_n1910_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n1911_));
AND2X2 AND2X2_728 ( .A(_abc_41356_new_n1864_), .B(_abc_41356_new_n1913_), .Y(_abc_41356_new_n1914_));
AND2X2 AND2X2_729 ( .A(_abc_41356_new_n1076_), .B(_abc_41356_new_n1893_), .Y(_abc_41356_new_n1916_));
AND2X2 AND2X2_73 ( .A(state_1_), .B(state_0_), .Y(_abc_41356_new_n610_));
AND2X2 AND2X2_730 ( .A(regfil_0__6_), .B(regfil_4__6_), .Y(_abc_41356_new_n1917_));
AND2X2 AND2X2_731 ( .A(_abc_41356_new_n1920_), .B(_abc_41356_new_n1921_), .Y(_abc_41356_new_n1922_));
AND2X2 AND2X2_732 ( .A(_abc_41356_new_n1922_), .B(_abc_41356_new_n1482_), .Y(_abc_41356_new_n1923_));
AND2X2 AND2X2_733 ( .A(_abc_41356_new_n1926_), .B(_abc_41356_new_n1893_), .Y(_abc_41356_new_n1927_));
AND2X2 AND2X2_734 ( .A(regfil_2__6_), .B(regfil_4__6_), .Y(_abc_41356_new_n1928_));
AND2X2 AND2X2_735 ( .A(_abc_41356_new_n1925_), .B(_abc_41356_new_n1930_), .Y(_abc_41356_new_n1931_));
AND2X2 AND2X2_736 ( .A(_abc_41356_new_n1932_), .B(_abc_41356_new_n1933_), .Y(_abc_41356_new_n1934_));
AND2X2 AND2X2_737 ( .A(_abc_41356_new_n1934_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n1935_));
AND2X2 AND2X2_738 ( .A(_abc_41356_new_n1418_), .B(_abc_41356_new_n1819_), .Y(_abc_41356_new_n1938_));
AND2X2 AND2X2_739 ( .A(_abc_41356_new_n1937_), .B(_abc_41356_new_n1939_), .Y(_abc_41356_new_n1940_));
AND2X2 AND2X2_74 ( .A(_abc_41356_new_n504_), .B(_abc_41356_new_n610_), .Y(_abc_41356_new_n611_));
AND2X2 AND2X2_740 ( .A(_abc_41356_new_n1877_), .B(regfil_4__6_), .Y(_abc_41356_new_n1944_));
AND2X2 AND2X2_741 ( .A(_abc_41356_new_n1945_), .B(_abc_41356_new_n1943_), .Y(_abc_41356_new_n1946_));
AND2X2 AND2X2_742 ( .A(_abc_41356_new_n1942_), .B(_abc_41356_new_n1947_), .Y(_abc_41356_new_n1948_));
AND2X2 AND2X2_743 ( .A(_abc_41356_new_n1949_), .B(_abc_41356_new_n1892_), .Y(_abc_41356_new_n1950_));
AND2X2 AND2X2_744 ( .A(_abc_41356_new_n1213_), .B(regfil_4__7_), .Y(_abc_41356_new_n1952_));
AND2X2 AND2X2_745 ( .A(_abc_41356_new_n1173_), .B(_abc_41356_new_n1212_), .Y(_abc_41356_new_n1953_));
AND2X2 AND2X2_746 ( .A(_abc_41356_new_n1954_), .B(_abc_41356_new_n1242_), .Y(_abc_41356_new_n1955_));
AND2X2 AND2X2_747 ( .A(_abc_41356_new_n1230_), .B(rdatahold_7_), .Y(_abc_41356_new_n1956_));
AND2X2 AND2X2_748 ( .A(_abc_41356_new_n1958_), .B(_abc_41356_new_n1248_), .Y(_abc_41356_new_n1959_));
AND2X2 AND2X2_749 ( .A(_abc_41356_new_n1963_), .B(_abc_41356_new_n1960_), .Y(_abc_41356_new_n1964_));
AND2X2 AND2X2_75 ( .A(_abc_41356_new_n519_), .B(_abc_41356_new_n611_), .Y(_abc_41356_new_n612_));
AND2X2 AND2X2_750 ( .A(_abc_41356_new_n1961_), .B(_abc_41356_new_n1967_), .Y(_abc_41356_new_n1968_));
AND2X2 AND2X2_751 ( .A(regfil_4__7_), .B(sp_15_), .Y(_abc_41356_new_n1969_));
AND2X2 AND2X2_752 ( .A(_abc_41356_new_n1966_), .B(_abc_41356_new_n1970_), .Y(_abc_41356_new_n1971_));
AND2X2 AND2X2_753 ( .A(_abc_41356_new_n1972_), .B(_abc_41356_new_n1973_), .Y(_abc_41356_new_n1974_));
AND2X2 AND2X2_754 ( .A(_abc_41356_new_n1975_), .B(_abc_41356_new_n1287_), .Y(_abc_41356_new_n1976_));
AND2X2 AND2X2_755 ( .A(_abc_41356_new_n535_), .B(regfil_4__6_), .Y(_abc_41356_new_n1977_));
AND2X2 AND2X2_756 ( .A(_abc_41356_new_n1237_), .B(_abc_41356_new_n1977_), .Y(_abc_41356_new_n1978_));
AND2X2 AND2X2_757 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n1978_), .Y(_abc_41356_new_n1979_));
AND2X2 AND2X2_758 ( .A(_abc_41356_new_n1134_), .B(_abc_41356_new_n1961_), .Y(_abc_41356_new_n1980_));
AND2X2 AND2X2_759 ( .A(regfil_0__7_), .B(regfil_4__7_), .Y(_abc_41356_new_n1981_));
AND2X2 AND2X2_76 ( .A(_abc_41356_new_n609_), .B(_abc_41356_new_n613_), .Y(_abc_41356_new_n614_));
AND2X2 AND2X2_760 ( .A(_abc_41356_new_n1915_), .B(_abc_41356_new_n1919_), .Y(_abc_41356_new_n1984_));
AND2X2 AND2X2_761 ( .A(_abc_41356_new_n1238_), .B(_abc_41356_new_n576_), .Y(_abc_41356_new_n1988_));
AND2X2 AND2X2_762 ( .A(_abc_41356_new_n1988_), .B(_abc_41356_new_n1990_), .Y(_abc_41356_new_n1991_));
AND2X2 AND2X2_763 ( .A(_abc_41356_new_n1987_), .B(_abc_41356_new_n1991_), .Y(_abc_41356_new_n1992_));
AND2X2 AND2X2_764 ( .A(_abc_41356_new_n1986_), .B(_abc_41356_new_n1992_), .Y(_abc_41356_new_n1993_));
AND2X2 AND2X2_765 ( .A(_abc_41356_new_n1996_), .B(_abc_41356_new_n1961_), .Y(_abc_41356_new_n1997_));
AND2X2 AND2X2_766 ( .A(regfil_2__7_), .B(regfil_4__7_), .Y(_abc_41356_new_n1998_));
AND2X2 AND2X2_767 ( .A(_abc_41356_new_n1238_), .B(_abc_41356_new_n1413_), .Y(_abc_41356_new_n2001_));
AND2X2 AND2X2_768 ( .A(_abc_41356_new_n2003_), .B(_abc_41356_new_n2001_), .Y(_abc_41356_new_n2004_));
AND2X2 AND2X2_769 ( .A(_abc_41356_new_n2004_), .B(_abc_41356_new_n2000_), .Y(_abc_41356_new_n2005_));
AND2X2 AND2X2_77 ( .A(_abc_41356_new_n615_), .B(opcode_0_), .Y(_abc_41356_new_n616_));
AND2X2 AND2X2_770 ( .A(_abc_41356_new_n1944_), .B(regfil_4__7_), .Y(_abc_41356_new_n2009_));
AND2X2 AND2X2_771 ( .A(_abc_41356_new_n2011_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n2012_));
AND2X2 AND2X2_772 ( .A(_abc_41356_new_n2012_), .B(_abc_41356_new_n2010_), .Y(_abc_41356_new_n2013_));
AND2X2 AND2X2_773 ( .A(_abc_41356_new_n2015_), .B(_abc_41356_new_n1965_), .Y(_abc_41356_new_n2016_));
AND2X2 AND2X2_774 ( .A(_abc_41356_new_n2017_), .B(_abc_41356_new_n1959_), .Y(_abc_41356_new_n2018_));
AND2X2 AND2X2_775 ( .A(_abc_41356_new_n2021_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n2023_));
AND2X2 AND2X2_776 ( .A(_abc_41356_new_n2024_), .B(wdatahold2_0_), .Y(_abc_41356_new_n2025_));
AND2X2 AND2X2_777 ( .A(_abc_41356_new_n578_), .B(_abc_41356_new_n623_), .Y(_abc_41356_new_n2026_));
AND2X2 AND2X2_778 ( .A(_abc_41356_new_n2026_), .B(_abc_41356_new_n535_), .Y(_abc_41356_new_n2027_));
AND2X2 AND2X2_779 ( .A(_abc_41356_new_n2030_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n2031_));
AND2X2 AND2X2_78 ( .A(_abc_41356_new_n616_), .B(regfil_1__0_), .Y(_abc_41356_new_n617_));
AND2X2 AND2X2_780 ( .A(_abc_41356_new_n2031_), .B(_abc_41356_new_n2029_), .Y(_abc_41356_new_n2032_));
AND2X2 AND2X2_781 ( .A(_abc_41356_new_n2033_), .B(pc_2_), .Y(_abc_41356_new_n2034_));
AND2X2 AND2X2_782 ( .A(_abc_41356_new_n2034_), .B(pc_3_), .Y(_abc_41356_new_n2035_));
AND2X2 AND2X2_783 ( .A(pc_5_), .B(pc_4_), .Y(_abc_41356_new_n2036_));
AND2X2 AND2X2_784 ( .A(pc_7_), .B(pc_6_), .Y(_abc_41356_new_n2037_));
AND2X2 AND2X2_785 ( .A(_abc_41356_new_n2036_), .B(_abc_41356_new_n2037_), .Y(_abc_41356_new_n2038_));
AND2X2 AND2X2_786 ( .A(_abc_41356_new_n2035_), .B(_abc_41356_new_n2038_), .Y(_abc_41356_new_n2039_));
AND2X2 AND2X2_787 ( .A(_abc_41356_new_n2039_), .B(pc_8_), .Y(_abc_41356_new_n2040_));
AND2X2 AND2X2_788 ( .A(_abc_41356_new_n2042_), .B(_abc_41356_new_n2041_), .Y(_abc_41356_new_n2043_));
AND2X2 AND2X2_789 ( .A(_abc_41356_new_n619_), .B(opcode_2_), .Y(_abc_41356_new_n2046_));
AND2X2 AND2X2_79 ( .A(_abc_41356_new_n615_), .B(_abc_41356_new_n618_), .Y(_abc_41356_new_n619_));
AND2X2 AND2X2_790 ( .A(_abc_41356_new_n616_), .B(_abc_41356_new_n527_), .Y(_abc_41356_new_n2047_));
AND2X2 AND2X2_791 ( .A(_abc_41356_new_n2047_), .B(_abc_41356_new_n576_), .Y(_abc_41356_new_n2048_));
AND2X2 AND2X2_792 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n2050_), .Y(_abc_41356_new_n2051_));
AND2X2 AND2X2_793 ( .A(_abc_41356_new_n2045_), .B(_abc_41356_new_n2052_), .Y(_abc_41356_new_n2053_));
AND2X2 AND2X2_794 ( .A(_abc_41356_new_n547_), .B(opcode_5_), .Y(_abc_41356_new_n2055_));
AND2X2 AND2X2_795 ( .A(_abc_41356_new_n2056_), .B(_abc_41356_new_n528_), .Y(_abc_41356_new_n2057_));
AND2X2 AND2X2_796 ( .A(_abc_41356_new_n2061_), .B(_abc_41356_new_n2054_), .Y(_abc_41356_new_n2062_));
AND2X2 AND2X2_797 ( .A(_abc_41356_new_n546_), .B(_abc_41356_new_n616_), .Y(_abc_41356_new_n2065_));
AND2X2 AND2X2_798 ( .A(_abc_41356_new_n2064_), .B(_abc_41356_new_n2066_), .Y(_abc_41356_new_n2067_));
AND2X2 AND2X2_799 ( .A(_abc_41356_new_n2067_), .B(_abc_41356_new_n2063_), .Y(_abc_41356_new_n2068_));
AND2X2 AND2X2_8 ( .A(_abc_41356_new_n508_), .B(_abc_41356_new_n511_), .Y(_abc_41356_new_n512_));
AND2X2 AND2X2_80 ( .A(_abc_41356_new_n619_), .B(regfil_0__0_), .Y(_abc_41356_new_n620_));
AND2X2 AND2X2_800 ( .A(_abc_41356_new_n2062_), .B(_abc_41356_new_n2068_), .Y(_abc_41356_new_n2069_));
AND2X2 AND2X2_801 ( .A(pc_2_), .B(pc_1_), .Y(_abc_41356_new_n2070_));
AND2X2 AND2X2_802 ( .A(_abc_41356_new_n2070_), .B(pc_3_), .Y(_abc_41356_new_n2071_));
AND2X2 AND2X2_803 ( .A(_abc_41356_new_n2071_), .B(pc_0_), .Y(_abc_41356_new_n2072_));
AND2X2 AND2X2_804 ( .A(_abc_41356_new_n2072_), .B(_abc_41356_new_n2038_), .Y(_abc_41356_new_n2073_));
AND2X2 AND2X2_805 ( .A(_abc_41356_new_n2074_), .B(_abc_41356_new_n2041_), .Y(_abc_41356_new_n2075_));
AND2X2 AND2X2_806 ( .A(_abc_41356_new_n2073_), .B(pc_8_), .Y(_abc_41356_new_n2076_));
AND2X2 AND2X2_807 ( .A(_abc_41356_new_n2078_), .B(_abc_41356_new_n2060_), .Y(_abc_41356_new_n2079_));
AND2X2 AND2X2_808 ( .A(_abc_41356_new_n2051_), .B(intcyc), .Y(_abc_41356_new_n2080_));
AND2X2 AND2X2_809 ( .A(_abc_41356_new_n681_), .B(regfil_7__0_), .Y(_abc_41356_new_n2081_));
AND2X2 AND2X2_81 ( .A(_abc_41356_new_n526_), .B(regfil_3__0_), .Y(_abc_41356_new_n622_));
AND2X2 AND2X2_810 ( .A(_abc_41356_new_n535_), .B(regfil_4__0_), .Y(_abc_41356_new_n2082_));
AND2X2 AND2X2_811 ( .A(opcode_4_), .B(regfil_2__0_), .Y(_abc_41356_new_n2084_));
AND2X2 AND2X2_812 ( .A(_abc_41356_new_n534_), .B(regfil_0__0_), .Y(_abc_41356_new_n2085_));
AND2X2 AND2X2_813 ( .A(_abc_41356_new_n2086_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n2087_));
AND2X2 AND2X2_814 ( .A(_abc_41356_new_n2088_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n2089_));
AND2X2 AND2X2_815 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n2082_), .Y(_abc_41356_new_n2090_));
AND2X2 AND2X2_816 ( .A(_abc_41356_new_n2097_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2098_));
AND2X2 AND2X2_817 ( .A(_abc_41356_new_n2098_), .B(_abc_41356_new_n2095_), .Y(_abc_41356_new_n2099_));
AND2X2 AND2X2_818 ( .A(_abc_41356_new_n2100_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2101_));
AND2X2 AND2X2_819 ( .A(_abc_41356_new_n2024_), .B(wdatahold2_1_), .Y(_abc_41356_new_n2103_));
AND2X2 AND2X2_82 ( .A(_abc_41356_new_n618_), .B(opcode_1_), .Y(_abc_41356_new_n623_));
AND2X2 AND2X2_820 ( .A(_abc_41356_new_n2105_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n2106_));
AND2X2 AND2X2_821 ( .A(_abc_41356_new_n2106_), .B(_abc_41356_new_n2104_), .Y(_abc_41356_new_n2107_));
AND2X2 AND2X2_822 ( .A(_abc_41356_new_n2040_), .B(pc_9_), .Y(_abc_41356_new_n2108_));
AND2X2 AND2X2_823 ( .A(_abc_41356_new_n2109_), .B(_abc_41356_new_n2110_), .Y(_abc_41356_new_n2111_));
AND2X2 AND2X2_824 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n2112_), .Y(_abc_41356_new_n2113_));
AND2X2 AND2X2_825 ( .A(_abc_41356_new_n2111_), .B(_abc_41356_new_n2114_), .Y(_abc_41356_new_n2115_));
AND2X2 AND2X2_826 ( .A(_abc_41356_new_n2076_), .B(pc_9_), .Y(_abc_41356_new_n2117_));
AND2X2 AND2X2_827 ( .A(_abc_41356_new_n2118_), .B(_abc_41356_new_n2116_), .Y(_abc_41356_new_n2119_));
AND2X2 AND2X2_828 ( .A(_abc_41356_new_n2119_), .B(_abc_41356_new_n2060_), .Y(_abc_41356_new_n2120_));
AND2X2 AND2X2_829 ( .A(_abc_41356_new_n2121_), .B(_abc_41356_new_n535_), .Y(_abc_41356_new_n2122_));
AND2X2 AND2X2_83 ( .A(_abc_41356_new_n623_), .B(regfil_2__0_), .Y(_abc_41356_new_n624_));
AND2X2 AND2X2_830 ( .A(_abc_41356_new_n2122_), .B(regfil_4__1_), .Y(_abc_41356_new_n2123_));
AND2X2 AND2X2_831 ( .A(_abc_41356_new_n681_), .B(regfil_7__1_), .Y(_abc_41356_new_n2124_));
AND2X2 AND2X2_832 ( .A(opcode_4_), .B(regfil_2__1_), .Y(_abc_41356_new_n2125_));
AND2X2 AND2X2_833 ( .A(_abc_41356_new_n534_), .B(regfil_0__1_), .Y(_abc_41356_new_n2126_));
AND2X2 AND2X2_834 ( .A(_abc_41356_new_n2127_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n2128_));
AND2X2 AND2X2_835 ( .A(_abc_41356_new_n2129_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n2130_));
AND2X2 AND2X2_836 ( .A(_abc_41356_new_n2113_), .B(intcyc), .Y(_abc_41356_new_n2131_));
AND2X2 AND2X2_837 ( .A(_abc_41356_new_n2137_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2138_));
AND2X2 AND2X2_838 ( .A(_abc_41356_new_n2136_), .B(_abc_41356_new_n2138_), .Y(_abc_41356_new_n2139_));
AND2X2 AND2X2_839 ( .A(_abc_41356_new_n2140_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2141_));
AND2X2 AND2X2_84 ( .A(_abc_41356_new_n616_), .B(regfil_5__0_), .Y(_abc_41356_new_n628_));
AND2X2 AND2X2_840 ( .A(_abc_41356_new_n2024_), .B(wdatahold2_2_), .Y(_abc_41356_new_n2143_));
AND2X2 AND2X2_841 ( .A(_abc_41356_new_n2145_), .B(_abc_41356_new_n2144_), .Y(_abc_41356_new_n2146_));
AND2X2 AND2X2_842 ( .A(_abc_41356_new_n2146_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n2147_));
AND2X2 AND2X2_843 ( .A(_abc_41356_new_n2108_), .B(pc_10_), .Y(_abc_41356_new_n2148_));
AND2X2 AND2X2_844 ( .A(_abc_41356_new_n2109_), .B(_abc_41356_new_n2149_), .Y(_abc_41356_new_n2150_));
AND2X2 AND2X2_845 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n2153_), .Y(_abc_41356_new_n2154_));
AND2X2 AND2X2_846 ( .A(_abc_41356_new_n2152_), .B(_abc_41356_new_n2155_), .Y(_abc_41356_new_n2156_));
AND2X2 AND2X2_847 ( .A(_abc_41356_new_n2118_), .B(_abc_41356_new_n2149_), .Y(_abc_41356_new_n2157_));
AND2X2 AND2X2_848 ( .A(_abc_41356_new_n2117_), .B(pc_10_), .Y(_abc_41356_new_n2158_));
AND2X2 AND2X2_849 ( .A(_abc_41356_new_n2160_), .B(_abc_41356_new_n2060_), .Y(_abc_41356_new_n2161_));
AND2X2 AND2X2_85 ( .A(_abc_41356_new_n623_), .B(regfil_6__0_), .Y(_abc_41356_new_n630_));
AND2X2 AND2X2_850 ( .A(_abc_41356_new_n681_), .B(regfil_7__2_), .Y(_abc_41356_new_n2162_));
AND2X2 AND2X2_851 ( .A(opcode_4_), .B(regfil_2__2_), .Y(_abc_41356_new_n2163_));
AND2X2 AND2X2_852 ( .A(_abc_41356_new_n534_), .B(regfil_0__2_), .Y(_abc_41356_new_n2164_));
AND2X2 AND2X2_853 ( .A(_abc_41356_new_n2165_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n2166_));
AND2X2 AND2X2_854 ( .A(_abc_41356_new_n2167_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n2168_));
AND2X2 AND2X2_855 ( .A(_abc_41356_new_n2154_), .B(intcyc), .Y(_abc_41356_new_n2169_));
AND2X2 AND2X2_856 ( .A(_abc_41356_new_n535_), .B(regfil_4__2_), .Y(_abc_41356_new_n2170_));
AND2X2 AND2X2_857 ( .A(_abc_41356_new_n2121_), .B(_abc_41356_new_n2170_), .Y(_abc_41356_new_n2171_));
AND2X2 AND2X2_858 ( .A(_abc_41356_new_n2177_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2178_));
AND2X2 AND2X2_859 ( .A(_abc_41356_new_n2176_), .B(_abc_41356_new_n2178_), .Y(_abc_41356_new_n2179_));
AND2X2 AND2X2_86 ( .A(_abc_41356_new_n619_), .B(regfil_4__0_), .Y(_abc_41356_new_n631_));
AND2X2 AND2X2_860 ( .A(_abc_41356_new_n2180_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2181_));
AND2X2 AND2X2_861 ( .A(_abc_41356_new_n2024_), .B(wdatahold2_3_), .Y(_abc_41356_new_n2183_));
AND2X2 AND2X2_862 ( .A(_abc_41356_new_n2185_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n2186_));
AND2X2 AND2X2_863 ( .A(_abc_41356_new_n2186_), .B(_abc_41356_new_n2184_), .Y(_abc_41356_new_n2187_));
AND2X2 AND2X2_864 ( .A(_abc_41356_new_n2148_), .B(pc_11_), .Y(_abc_41356_new_n2188_));
AND2X2 AND2X2_865 ( .A(_abc_41356_new_n2189_), .B(_abc_41356_new_n2190_), .Y(_abc_41356_new_n2191_));
AND2X2 AND2X2_866 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n2192_), .Y(_abc_41356_new_n2193_));
AND2X2 AND2X2_867 ( .A(_abc_41356_new_n2191_), .B(_abc_41356_new_n2194_), .Y(_abc_41356_new_n2195_));
AND2X2 AND2X2_868 ( .A(_abc_41356_new_n2158_), .B(pc_11_), .Y(_abc_41356_new_n2197_));
AND2X2 AND2X2_869 ( .A(_abc_41356_new_n2198_), .B(_abc_41356_new_n2196_), .Y(_abc_41356_new_n2199_));
AND2X2 AND2X2_87 ( .A(_abc_41356_new_n526_), .B(regfil_7__0_), .Y(_abc_41356_new_n632_));
AND2X2 AND2X2_870 ( .A(_abc_41356_new_n2199_), .B(_abc_41356_new_n2060_), .Y(_abc_41356_new_n2200_));
AND2X2 AND2X2_871 ( .A(_abc_41356_new_n2122_), .B(regfil_4__3_), .Y(_abc_41356_new_n2201_));
AND2X2 AND2X2_872 ( .A(_abc_41356_new_n681_), .B(regfil_7__3_), .Y(_abc_41356_new_n2202_));
AND2X2 AND2X2_873 ( .A(opcode_4_), .B(regfil_2__3_), .Y(_abc_41356_new_n2203_));
AND2X2 AND2X2_874 ( .A(_abc_41356_new_n534_), .B(regfil_0__3_), .Y(_abc_41356_new_n2204_));
AND2X2 AND2X2_875 ( .A(_abc_41356_new_n2205_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n2206_));
AND2X2 AND2X2_876 ( .A(_abc_41356_new_n2207_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n2208_));
AND2X2 AND2X2_877 ( .A(_abc_41356_new_n2193_), .B(intcyc), .Y(_abc_41356_new_n2209_));
AND2X2 AND2X2_878 ( .A(_abc_41356_new_n2215_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2216_));
AND2X2 AND2X2_879 ( .A(_abc_41356_new_n2214_), .B(_abc_41356_new_n2216_), .Y(_abc_41356_new_n2217_));
AND2X2 AND2X2_88 ( .A(_abc_41356_new_n627_), .B(_abc_41356_new_n635_), .Y(_abc_41356_new_n636_));
AND2X2 AND2X2_880 ( .A(_abc_41356_new_n2218_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2219_));
AND2X2 AND2X2_881 ( .A(_abc_41356_new_n2024_), .B(wdatahold2_4_), .Y(_abc_41356_new_n2221_));
AND2X2 AND2X2_882 ( .A(_abc_41356_new_n2223_), .B(_abc_41356_new_n2222_), .Y(_abc_41356_new_n2224_));
AND2X2 AND2X2_883 ( .A(_abc_41356_new_n2224_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n2225_));
AND2X2 AND2X2_884 ( .A(_abc_41356_new_n2188_), .B(pc_12_), .Y(_abc_41356_new_n2226_));
AND2X2 AND2X2_885 ( .A(_abc_41356_new_n2189_), .B(_abc_41356_new_n2227_), .Y(_abc_41356_new_n2228_));
AND2X2 AND2X2_886 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n2231_), .Y(_abc_41356_new_n2232_));
AND2X2 AND2X2_887 ( .A(_abc_41356_new_n2230_), .B(_abc_41356_new_n2233_), .Y(_abc_41356_new_n2234_));
AND2X2 AND2X2_888 ( .A(_abc_41356_new_n2198_), .B(_abc_41356_new_n2227_), .Y(_abc_41356_new_n2235_));
AND2X2 AND2X2_889 ( .A(_abc_41356_new_n2197_), .B(pc_12_), .Y(_abc_41356_new_n2236_));
AND2X2 AND2X2_89 ( .A(_abc_41356_new_n636_), .B(_abc_41356_new_n614_), .Y(_abc_41356_new_n637_));
AND2X2 AND2X2_890 ( .A(_abc_41356_new_n2238_), .B(_abc_41356_new_n2060_), .Y(_abc_41356_new_n2239_));
AND2X2 AND2X2_891 ( .A(_abc_41356_new_n681_), .B(regfil_7__4_), .Y(_abc_41356_new_n2240_));
AND2X2 AND2X2_892 ( .A(opcode_4_), .B(regfil_2__4_), .Y(_abc_41356_new_n2241_));
AND2X2 AND2X2_893 ( .A(_abc_41356_new_n534_), .B(regfil_0__4_), .Y(_abc_41356_new_n2242_));
AND2X2 AND2X2_894 ( .A(_abc_41356_new_n2243_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n2244_));
AND2X2 AND2X2_895 ( .A(_abc_41356_new_n2245_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n2246_));
AND2X2 AND2X2_896 ( .A(_abc_41356_new_n2232_), .B(intcyc), .Y(_abc_41356_new_n2247_));
AND2X2 AND2X2_897 ( .A(_abc_41356_new_n535_), .B(regfil_4__4_), .Y(_abc_41356_new_n2248_));
AND2X2 AND2X2_898 ( .A(_abc_41356_new_n2121_), .B(_abc_41356_new_n2248_), .Y(_abc_41356_new_n2249_));
AND2X2 AND2X2_899 ( .A(_abc_41356_new_n2255_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2256_));
AND2X2 AND2X2_9 ( .A(_abc_41356_new_n514_), .B(_abc_41356_new_n515_), .Y(_abc_41356_new_n516_));
AND2X2 AND2X2_90 ( .A(_abc_41356_new_n612_), .B(alu_res_0_), .Y(_abc_41356_new_n638_));
AND2X2 AND2X2_900 ( .A(_abc_41356_new_n2254_), .B(_abc_41356_new_n2256_), .Y(_abc_41356_new_n2257_));
AND2X2 AND2X2_901 ( .A(_abc_41356_new_n2258_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2259_));
AND2X2 AND2X2_902 ( .A(_abc_41356_new_n2024_), .B(wdatahold2_5_), .Y(_abc_41356_new_n2261_));
AND2X2 AND2X2_903 ( .A(_abc_41356_new_n2263_), .B(_abc_41356_new_n2262_), .Y(_abc_41356_new_n2264_));
AND2X2 AND2X2_904 ( .A(_abc_41356_new_n2264_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n2265_));
AND2X2 AND2X2_905 ( .A(_abc_41356_new_n2226_), .B(pc_13_), .Y(_abc_41356_new_n2266_));
AND2X2 AND2X2_906 ( .A(_abc_41356_new_n2267_), .B(_abc_41356_new_n2268_), .Y(_abc_41356_new_n2269_));
AND2X2 AND2X2_907 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n2270_), .Y(_abc_41356_new_n2271_));
AND2X2 AND2X2_908 ( .A(_abc_41356_new_n2269_), .B(_abc_41356_new_n2272_), .Y(_abc_41356_new_n2273_));
AND2X2 AND2X2_909 ( .A(_abc_41356_new_n2236_), .B(pc_13_), .Y(_abc_41356_new_n2275_));
AND2X2 AND2X2_91 ( .A(_abc_41356_new_n639_), .B(_abc_41356_new_n604_), .Y(_abc_41356_new_n640_));
AND2X2 AND2X2_910 ( .A(_abc_41356_new_n2276_), .B(_abc_41356_new_n2274_), .Y(_abc_41356_new_n2277_));
AND2X2 AND2X2_911 ( .A(_abc_41356_new_n2277_), .B(_abc_41356_new_n2060_), .Y(_abc_41356_new_n2278_));
AND2X2 AND2X2_912 ( .A(_abc_41356_new_n2122_), .B(regfil_4__5_), .Y(_abc_41356_new_n2279_));
AND2X2 AND2X2_913 ( .A(_abc_41356_new_n2271_), .B(intcyc), .Y(_abc_41356_new_n2280_));
AND2X2 AND2X2_914 ( .A(_abc_41356_new_n681_), .B(regfil_7__5_), .Y(_abc_41356_new_n2281_));
AND2X2 AND2X2_915 ( .A(opcode_4_), .B(regfil_2__5_), .Y(_abc_41356_new_n2282_));
AND2X2 AND2X2_916 ( .A(_abc_41356_new_n534_), .B(regfil_0__5_), .Y(_abc_41356_new_n2283_));
AND2X2 AND2X2_917 ( .A(_abc_41356_new_n2284_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n2285_));
AND2X2 AND2X2_918 ( .A(_abc_41356_new_n2286_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n2287_));
AND2X2 AND2X2_919 ( .A(_abc_41356_new_n2293_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2294_));
AND2X2 AND2X2_92 ( .A(_abc_41356_new_n642_), .B(rdatahold_0_), .Y(_abc_41356_new_n643_));
AND2X2 AND2X2_920 ( .A(_abc_41356_new_n2292_), .B(_abc_41356_new_n2294_), .Y(_abc_41356_new_n2295_));
AND2X2 AND2X2_921 ( .A(_abc_41356_new_n2296_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2297_));
AND2X2 AND2X2_922 ( .A(_abc_41356_new_n2024_), .B(wdatahold2_6_), .Y(_abc_41356_new_n2299_));
AND2X2 AND2X2_923 ( .A(_abc_41356_new_n2301_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n2302_));
AND2X2 AND2X2_924 ( .A(_abc_41356_new_n2302_), .B(_abc_41356_new_n2300_), .Y(_abc_41356_new_n2303_));
AND2X2 AND2X2_925 ( .A(_abc_41356_new_n2266_), .B(pc_14_), .Y(_abc_41356_new_n2304_));
AND2X2 AND2X2_926 ( .A(_abc_41356_new_n2305_), .B(_abc_41356_new_n2306_), .Y(_abc_41356_new_n2307_));
AND2X2 AND2X2_927 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n2308_), .Y(_abc_41356_new_n2309_));
AND2X2 AND2X2_928 ( .A(_abc_41356_new_n2307_), .B(_abc_41356_new_n2310_), .Y(_abc_41356_new_n2311_));
AND2X2 AND2X2_929 ( .A(_abc_41356_new_n2275_), .B(pc_14_), .Y(_abc_41356_new_n2313_));
AND2X2 AND2X2_93 ( .A(_abc_41356_new_n647_), .B(_abc_41356_new_n648_), .Y(_abc_41356_new_n649_));
AND2X2 AND2X2_930 ( .A(_abc_41356_new_n2314_), .B(_abc_41356_new_n2312_), .Y(_abc_41356_new_n2315_));
AND2X2 AND2X2_931 ( .A(_abc_41356_new_n2315_), .B(_abc_41356_new_n2060_), .Y(_abc_41356_new_n2316_));
AND2X2 AND2X2_932 ( .A(_abc_41356_new_n681_), .B(regfil_7__6_), .Y(_abc_41356_new_n2317_));
AND2X2 AND2X2_933 ( .A(opcode_4_), .B(regfil_2__6_), .Y(_abc_41356_new_n2318_));
AND2X2 AND2X2_934 ( .A(_abc_41356_new_n534_), .B(regfil_0__6_), .Y(_abc_41356_new_n2319_));
AND2X2 AND2X2_935 ( .A(_abc_41356_new_n2320_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n2321_));
AND2X2 AND2X2_936 ( .A(_abc_41356_new_n2322_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n2323_));
AND2X2 AND2X2_937 ( .A(_abc_41356_new_n2309_), .B(intcyc), .Y(_abc_41356_new_n2324_));
AND2X2 AND2X2_938 ( .A(_abc_41356_new_n2121_), .B(_abc_41356_new_n1977_), .Y(_abc_41356_new_n2325_));
AND2X2 AND2X2_939 ( .A(_abc_41356_new_n2331_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2332_));
AND2X2 AND2X2_94 ( .A(_abc_41356_new_n649_), .B(_abc_41356_new_n646_), .Y(_abc_41356_new_n650_));
AND2X2 AND2X2_940 ( .A(_abc_41356_new_n2330_), .B(_abc_41356_new_n2332_), .Y(_abc_41356_new_n2333_));
AND2X2 AND2X2_941 ( .A(_abc_41356_new_n2334_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2335_));
AND2X2 AND2X2_942 ( .A(_abc_41356_new_n2024_), .B(wdatahold2_7_), .Y(_abc_41356_new_n2337_));
AND2X2 AND2X2_943 ( .A(_abc_41356_new_n2339_), .B(_abc_41356_new_n2338_), .Y(_abc_41356_new_n2340_));
AND2X2 AND2X2_944 ( .A(_abc_41356_new_n2340_), .B(_abc_41356_new_n516_), .Y(_abc_41356_new_n2341_));
AND2X2 AND2X2_945 ( .A(_abc_41356_new_n2304_), .B(pc_15_), .Y(_abc_41356_new_n2343_));
AND2X2 AND2X2_946 ( .A(_abc_41356_new_n2344_), .B(_abc_41356_new_n2342_), .Y(_abc_41356_new_n2345_));
AND2X2 AND2X2_947 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n2346_), .Y(_abc_41356_new_n2347_));
AND2X2 AND2X2_948 ( .A(_abc_41356_new_n2345_), .B(_abc_41356_new_n2348_), .Y(_abc_41356_new_n2349_));
AND2X2 AND2X2_949 ( .A(_abc_41356_new_n2313_), .B(pc_15_), .Y(_abc_41356_new_n2351_));
AND2X2 AND2X2_95 ( .A(_abc_41356_new_n650_), .B(_abc_41356_new_n645_), .Y(_abc_41356_new_n651_));
AND2X2 AND2X2_950 ( .A(_abc_41356_new_n2352_), .B(_abc_41356_new_n2350_), .Y(_abc_41356_new_n2353_));
AND2X2 AND2X2_951 ( .A(_abc_41356_new_n2353_), .B(_abc_41356_new_n2060_), .Y(_abc_41356_new_n2354_));
AND2X2 AND2X2_952 ( .A(_abc_41356_new_n2122_), .B(regfil_4__7_), .Y(_abc_41356_new_n2355_));
AND2X2 AND2X2_953 ( .A(_abc_41356_new_n2347_), .B(intcyc), .Y(_abc_41356_new_n2356_));
AND2X2 AND2X2_954 ( .A(_abc_41356_new_n681_), .B(regfil_7__7_), .Y(_abc_41356_new_n2357_));
AND2X2 AND2X2_955 ( .A(opcode_4_), .B(regfil_2__7_), .Y(_abc_41356_new_n2358_));
AND2X2 AND2X2_956 ( .A(_abc_41356_new_n534_), .B(regfil_0__7_), .Y(_abc_41356_new_n2359_));
AND2X2 AND2X2_957 ( .A(_abc_41356_new_n2360_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n2361_));
AND2X2 AND2X2_958 ( .A(_abc_41356_new_n2362_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n2363_));
AND2X2 AND2X2_959 ( .A(_abc_41356_new_n2369_), .B(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2370_));
AND2X2 AND2X2_96 ( .A(_abc_41356_new_n657_), .B(_abc_41356_new_n644_), .Y(_abc_41356_new_n658_));
AND2X2 AND2X2_960 ( .A(_abc_41356_new_n2368_), .B(_abc_41356_new_n2370_), .Y(_abc_41356_new_n2371_));
AND2X2 AND2X2_961 ( .A(_abc_41356_new_n2372_), .B(_abc_41356_new_n523_), .Y(_abc_41356_new_n2373_));
AND2X2 AND2X2_962 ( .A(_abc_41356_new_n526_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n2376_));
AND2X2 AND2X2_963 ( .A(_abc_41356_new_n2376_), .B(_abc_41356_new_n1413_), .Y(_abc_41356_new_n2377_));
AND2X2 AND2X2_964 ( .A(_abc_41356_new_n524_), .B(_abc_41356_new_n2377_), .Y(_abc_41356_new_n2378_));
AND2X2 AND2X2_965 ( .A(_abc_41356_new_n2378_), .B(_abc_41356_new_n2375_), .Y(_abc_41356_new_n2379_));
AND2X2 AND2X2_966 ( .A(_abc_41356_new_n2380_), .B(_abc_41356_new_n2381_), .Y(_abc_41356_new_n2382_));
AND2X2 AND2X2_967 ( .A(_abc_41356_new_n2383_), .B(_abc_41356_new_n1207_), .Y(_abc_41356_new_n2384_));
AND2X2 AND2X2_968 ( .A(_abc_41356_new_n694_), .B(_abc_41356_new_n2384_), .Y(_abc_41356_new_n2385_));
AND2X2 AND2X2_969 ( .A(_abc_41356_new_n506_), .B(_abc_41356_new_n587_), .Y(_abc_41356_new_n2388_));
AND2X2 AND2X2_97 ( .A(_abc_41356_new_n656_), .B(regfil_0__0_), .Y(_abc_41356_new_n659_));
AND2X2 AND2X2_970 ( .A(_abc_41356_new_n519_), .B(_abc_41356_new_n2388_), .Y(_abc_41356_new_n2389_));
AND2X2 AND2X2_971 ( .A(_abc_41356_new_n509_), .B(_abc_41356_new_n591_), .Y(_abc_41356_new_n2390_));
AND2X2 AND2X2_972 ( .A(_abc_41356_new_n2390_), .B(popdes_0_), .Y(_abc_41356_new_n2391_));
AND2X2 AND2X2_973 ( .A(_abc_41356_new_n508_), .B(_abc_41356_new_n2391_), .Y(_abc_41356_new_n2392_));
AND2X2 AND2X2_974 ( .A(_abc_41356_new_n2397_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2398_));
AND2X2 AND2X2_975 ( .A(_abc_41356_new_n2387_), .B(_abc_41356_new_n2398_), .Y(_abc_41356_new_n2399_));
AND2X2 AND2X2_976 ( .A(_abc_41356_new_n2393_), .B(rdatahold2_0_), .Y(_abc_41356_new_n2400_));
AND2X2 AND2X2_977 ( .A(_abc_41356_new_n2404_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2405_));
AND2X2 AND2X2_978 ( .A(_abc_41356_new_n2403_), .B(_abc_41356_new_n2405_), .Y(_abc_41356_new_n2406_));
AND2X2 AND2X2_979 ( .A(_abc_41356_new_n2393_), .B(rdatahold2_1_), .Y(_abc_41356_new_n2407_));
AND2X2 AND2X2_98 ( .A(_abc_41356_new_n660_), .B(_abc_41356_new_n601_), .Y(_abc_41356_new_n661_));
AND2X2 AND2X2_980 ( .A(regfil_3__0_), .B(regfil_3__1_), .Y(_abc_41356_new_n2408_));
AND2X2 AND2X2_981 ( .A(_abc_41356_new_n2375_), .B(_abc_41356_new_n2409_), .Y(_abc_41356_new_n2410_));
AND2X2 AND2X2_982 ( .A(_abc_41356_new_n2378_), .B(opcode_3_), .Y(_abc_41356_new_n2412_));
AND2X2 AND2X2_983 ( .A(_abc_41356_new_n2412_), .B(_abc_41356_new_n2411_), .Y(_abc_41356_new_n2413_));
AND2X2 AND2X2_984 ( .A(_abc_41356_new_n2378_), .B(_abc_41356_new_n545_), .Y(_abc_41356_new_n2415_));
AND2X2 AND2X2_985 ( .A(_abc_41356_new_n2415_), .B(_abc_41356_new_n2414_), .Y(_abc_41356_new_n2416_));
AND2X2 AND2X2_986 ( .A(_abc_41356_new_n508_), .B(_abc_41356_new_n591_), .Y(_abc_41356_new_n2419_));
AND2X2 AND2X2_987 ( .A(_abc_41356_new_n509_), .B(popdes_0_), .Y(_abc_41356_new_n2420_));
AND2X2 AND2X2_988 ( .A(_abc_41356_new_n2419_), .B(_abc_41356_new_n2420_), .Y(_abc_41356_new_n2421_));
AND2X2 AND2X2_989 ( .A(_abc_41356_new_n2423_), .B(_abc_41356_new_n2422_), .Y(_abc_41356_new_n2424_));
AND2X2 AND2X2_99 ( .A(_abc_41356_new_n614_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n665_));
AND2X2 AND2X2_990 ( .A(_abc_41356_new_n2418_), .B(_abc_41356_new_n2424_), .Y(_abc_41356_new_n2425_));
AND2X2 AND2X2_991 ( .A(_abc_41356_new_n2429_), .B(_abc_41356_new_n2396_), .Y(_abc_41356_new_n2430_));
AND2X2 AND2X2_992 ( .A(_abc_41356_new_n2428_), .B(_abc_41356_new_n2430_), .Y(_abc_41356_new_n2431_));
AND2X2 AND2X2_993 ( .A(_abc_41356_new_n2393_), .B(rdatahold2_2_), .Y(_abc_41356_new_n2432_));
AND2X2 AND2X2_994 ( .A(_abc_41356_new_n2410_), .B(_abc_41356_new_n1370_), .Y(_abc_41356_new_n2433_));
AND2X2 AND2X2_995 ( .A(_abc_41356_new_n2434_), .B(regfil_3__2_), .Y(_abc_41356_new_n2435_));
AND2X2 AND2X2_996 ( .A(_abc_41356_new_n2412_), .B(_abc_41356_new_n2436_), .Y(_abc_41356_new_n2437_));
AND2X2 AND2X2_997 ( .A(_abc_41356_new_n2408_), .B(regfil_3__2_), .Y(_abc_41356_new_n2439_));
AND2X2 AND2X2_998 ( .A(_abc_41356_new_n2440_), .B(_abc_41356_new_n2438_), .Y(_abc_41356_new_n2441_));
AND2X2 AND2X2_999 ( .A(_abc_41356_new_n2415_), .B(_abc_41356_new_n2441_), .Y(_abc_41356_new_n2442_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_0_), .Q(state_0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_3_), .Q(regfil_4__3_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(clock), .D(_0sp_15_0__8_), .Q(sp_8_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(clock), .D(_0sp_15_0__9_), .Q(sp_9_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(clock), .D(_0sp_15_0__10_), .Q(sp_10_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(clock), .D(_0sp_15_0__11_), .Q(sp_11_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(clock), .D(_0sp_15_0__12_), .Q(sp_12_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(clock), .D(_0sp_15_0__13_), .Q(sp_13_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(clock), .D(_0sp_15_0__14_), .Q(sp_14_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(clock), .D(_0sp_15_0__15_), .Q(sp_15_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(clock), .D(_0regd_2_0__0_), .Q(regd_0_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(clock), .D(_0regd_2_0__1_), .Q(regd_1_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_4_), .Q(regfil_4__4_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(clock), .D(_0regd_2_0__2_), .Q(regd_2_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(clock), .D(_0datao_7_0__0_), .Q(\data[0] ));
DFFPOSX1 DFFPOSX1_112 ( .CLK(clock), .D(_0datao_7_0__1_), .Q(\data[1] ));
DFFPOSX1 DFFPOSX1_113 ( .CLK(clock), .D(_0datao_7_0__2_), .Q(\data[2] ));
DFFPOSX1 DFFPOSX1_114 ( .CLK(clock), .D(_0datao_7_0__3_), .Q(\data[3] ));
DFFPOSX1 DFFPOSX1_115 ( .CLK(clock), .D(_0datao_7_0__4_), .Q(\data[4] ));
DFFPOSX1 DFFPOSX1_116 ( .CLK(clock), .D(_0datao_7_0__5_), .Q(\data[5] ));
DFFPOSX1 DFFPOSX1_117 ( .CLK(clock), .D(_0datao_7_0__6_), .Q(\data[6] ));
DFFPOSX1 DFFPOSX1_118 ( .CLK(clock), .D(_0datao_7_0__7_), .Q(\data[7] ));
DFFPOSX1 DFFPOSX1_119 ( .CLK(clock), .D(_0waddrhold_15_0__0_), .Q(waddrhold_0_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_5_), .Q(regfil_4__5_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(clock), .D(_0waddrhold_15_0__1_), .Q(waddrhold_1_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(clock), .D(_0waddrhold_15_0__2_), .Q(waddrhold_2_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(clock), .D(_0waddrhold_15_0__3_), .Q(waddrhold_3_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(clock), .D(_0waddrhold_15_0__4_), .Q(waddrhold_4_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(clock), .D(_0waddrhold_15_0__5_), .Q(waddrhold_5_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(clock), .D(_0waddrhold_15_0__6_), .Q(waddrhold_6_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(clock), .D(_0waddrhold_15_0__7_), .Q(waddrhold_7_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(clock), .D(_0waddrhold_15_0__8_), .Q(waddrhold_8_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(clock), .D(_0waddrhold_15_0__9_), .Q(waddrhold_9_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(clock), .D(_0waddrhold_15_0__10_), .Q(waddrhold_10_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_6_), .Q(regfil_4__6_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(clock), .D(_0waddrhold_15_0__11_), .Q(waddrhold_11_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(clock), .D(_0waddrhold_15_0__12_), .Q(waddrhold_12_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(clock), .D(_0waddrhold_15_0__13_), .Q(waddrhold_13_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(clock), .D(_0waddrhold_15_0__14_), .Q(waddrhold_14_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(clock), .D(_0waddrhold_15_0__15_), .Q(waddrhold_15_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(clock), .D(_0raddrhold_15_0__0_), .Q(raddrhold_0_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(clock), .D(_0raddrhold_15_0__1_), .Q(raddrhold_1_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(clock), .D(_0raddrhold_15_0__2_), .Q(raddrhold_2_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(clock), .D(_0raddrhold_15_0__3_), .Q(raddrhold_3_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(clock), .D(_0raddrhold_15_0__4_), .Q(raddrhold_4_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_7_), .Q(regfil_4__7_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(clock), .D(_0raddrhold_15_0__5_), .Q(raddrhold_5_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(clock), .D(_0raddrhold_15_0__6_), .Q(raddrhold_6_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(clock), .D(_0raddrhold_15_0__7_), .Q(raddrhold_7_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(clock), .D(_0raddrhold_15_0__8_), .Q(raddrhold_8_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(clock), .D(_0raddrhold_15_0__9_), .Q(raddrhold_9_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(clock), .D(_0raddrhold_15_0__10_), .Q(raddrhold_10_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(clock), .D(_0raddrhold_15_0__11_), .Q(raddrhold_11_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(clock), .D(_0raddrhold_15_0__12_), .Q(raddrhold_12_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(clock), .D(_0raddrhold_15_0__13_), .Q(raddrhold_13_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(clock), .D(_0raddrhold_15_0__14_), .Q(raddrhold_14_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_0_), .Q(regfil_5__0_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(clock), .D(_0raddrhold_15_0__15_), .Q(raddrhold_15_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(clock), .D(_0wdatahold_7_0__0_), .Q(wdatahold_0_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(clock), .D(_0wdatahold_7_0__1_), .Q(wdatahold_1_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(clock), .D(_0wdatahold_7_0__2_), .Q(wdatahold_2_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(clock), .D(_0wdatahold_7_0__3_), .Q(wdatahold_3_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(clock), .D(_0wdatahold_7_0__4_), .Q(wdatahold_4_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(clock), .D(_0wdatahold_7_0__5_), .Q(wdatahold_5_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(clock), .D(_0wdatahold_7_0__6_), .Q(wdatahold_6_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(clock), .D(_0wdatahold_7_0__7_), .Q(wdatahold_7_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(clock), .D(_0wdatahold2_7_0__0_), .Q(wdatahold2_0_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_1_), .Q(regfil_5__1_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(clock), .D(_0wdatahold2_7_0__1_), .Q(wdatahold2_1_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(clock), .D(_0wdatahold2_7_0__2_), .Q(wdatahold2_2_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(clock), .D(_0wdatahold2_7_0__3_), .Q(wdatahold2_3_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(clock), .D(_0wdatahold2_7_0__4_), .Q(wdatahold2_4_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(clock), .D(_0wdatahold2_7_0__5_), .Q(wdatahold2_5_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(clock), .D(_0wdatahold2_7_0__6_), .Q(wdatahold2_6_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(clock), .D(_0wdatahold2_7_0__7_), .Q(wdatahold2_7_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(clock), .D(_0rdatahold_7_0__0_), .Q(rdatahold_0_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(clock), .D(_0rdatahold_7_0__1_), .Q(rdatahold_1_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(clock), .D(_0rdatahold_7_0__2_), .Q(rdatahold_2_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_2_), .Q(regfil_5__2_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(clock), .D(_0rdatahold_7_0__3_), .Q(rdatahold_3_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(clock), .D(_0rdatahold_7_0__4_), .Q(rdatahold_4_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(clock), .D(_0rdatahold_7_0__5_), .Q(rdatahold_5_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(clock), .D(_0rdatahold_7_0__6_), .Q(rdatahold_6_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(clock), .D(_0rdatahold_7_0__7_), .Q(rdatahold_7_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(clock), .D(_0rdatahold2_7_0__0_), .Q(rdatahold2_0_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(clock), .D(_0rdatahold2_7_0__1_), .Q(rdatahold2_1_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(clock), .D(_0rdatahold2_7_0__2_), .Q(rdatahold2_2_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(clock), .D(_0rdatahold2_7_0__3_), .Q(rdatahold2_3_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(clock), .D(_0rdatahold2_7_0__4_), .Q(rdatahold2_4_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_3_), .Q(regfil_5__3_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(clock), .D(_0rdatahold2_7_0__5_), .Q(rdatahold2_5_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(clock), .D(_0rdatahold2_7_0__6_), .Q(rdatahold2_6_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(clock), .D(_0rdatahold2_7_0__7_), .Q(rdatahold2_7_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(clock), .D(_0popdes_1_0__0_), .Q(popdes_0_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(clock), .D(_0popdes_1_0__1_), .Q(popdes_1_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(clock), .D(_0statesel_5_0__0_), .Q(statesel_0_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(clock), .D(_0statesel_5_0__1_), .Q(statesel_1_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(clock), .D(_0statesel_5_0__2_), .Q(statesel_2_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(clock), .D(_0statesel_5_0__3_), .Q(statesel_3_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(clock), .D(_0statesel_5_0__4_), .Q(statesel_4_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_4_), .Q(regfil_5__4_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(clock), .D(_0statesel_5_0__5_), .Q(statesel_5_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(clock), .D(_0eienb_0_0_), .Q(eienb));
DFFPOSX1 DFFPOSX1_192 ( .CLK(clock), .D(_0opcode_7_0__0_), .Q(opcode_0_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(clock), .D(_0opcode_7_0__1_), .Q(opcode_1_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(clock), .D(_0opcode_7_0__2_), .Q(opcode_2_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(clock), .D(_0opcode_7_0__3_), .Q(opcode_3_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(clock), .D(_0opcode_7_0__4_), .Q(opcode_4_));
DFFPOSX1 DFFPOSX1_197 ( .CLK(clock), .D(_0opcode_7_0__5_), .Q(opcode_5_));
DFFPOSX1 DFFPOSX1_198 ( .CLK(clock), .D(_0opcode_7_0__6_), .Q(opcode_6_));
DFFPOSX1 DFFPOSX1_199 ( .CLK(clock), .D(_0opcode_7_0__7_), .Q(opcode_7_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_1_), .Q(state_1_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_5_), .Q(regfil_5__5_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(clock), .D(_0carry_0_0_), .Q(carry));
DFFPOSX1 DFFPOSX1_201 ( .CLK(clock), .D(_0auxcar_0_0_), .Q(auxcar));
DFFPOSX1 DFFPOSX1_202 ( .CLK(clock), .D(_0sign_0_0_), .Q(sign));
DFFPOSX1 DFFPOSX1_203 ( .CLK(clock), .D(_0zero_0_0_), .Q(zero));
DFFPOSX1 DFFPOSX1_204 ( .CLK(clock), .D(_0parity_0_0_), .Q(parity));
DFFPOSX1 DFFPOSX1_205 ( .CLK(clock), .D(_0ei_0_0_), .Q(ei));
DFFPOSX1 DFFPOSX1_206 ( .CLK(clock), .D(_0intcyc_0_0_), .Q(intcyc));
DFFPOSX1 DFFPOSX1_207 ( .CLK(clock), .D(_0aluopra_7_0__0_), .Q(alu_opra_0_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(clock), .D(_0aluopra_7_0__1_), .Q(alu_opra_1_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(clock), .D(_0aluopra_7_0__2_), .Q(alu_opra_2_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_6_), .Q(regfil_5__6_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(clock), .D(_0aluopra_7_0__3_), .Q(alu_opra_3_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(clock), .D(_0aluopra_7_0__4_), .Q(alu_opra_4_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(clock), .D(_0aluopra_7_0__5_), .Q(alu_opra_5_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(clock), .D(_0aluopra_7_0__6_), .Q(alu_opra_6_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(clock), .D(_0aluopra_7_0__7_), .Q(alu_opra_7_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(clock), .D(_0aluoprb_7_0__0_), .Q(alu_oprb_0_));
DFFPOSX1 DFFPOSX1_216 ( .CLK(clock), .D(_0aluoprb_7_0__1_), .Q(alu_oprb_1_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(clock), .D(_0aluoprb_7_0__2_), .Q(alu_oprb_2_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(clock), .D(_0aluoprb_7_0__3_), .Q(alu_oprb_3_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(clock), .D(_0aluoprb_7_0__4_), .Q(alu_oprb_4_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_7_), .Q(regfil_5__7_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(clock), .D(_0aluoprb_7_0__5_), .Q(alu_oprb_5_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(clock), .D(_0aluoprb_7_0__6_), .Q(alu_oprb_6_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(clock), .D(_0aluoprb_7_0__7_), .Q(alu_oprb_7_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(clock), .D(_0alucin_0_0_), .Q(alu_cin));
DFFPOSX1 DFFPOSX1_224 ( .CLK(clock), .D(_0alusel_2_0__0_), .Q(alu_sel_0_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(clock), .D(_0alusel_2_0__1_), .Q(alu_sel_1_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(clock), .D(_0alusel_2_0__2_), .Q(alu_sel_2_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_0_), .Q(regfil_7__0_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_1_), .Q(regfil_7__1_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_2_), .Q(regfil_7__2_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_0_), .Q(regfil_1__0_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_3_), .Q(regfil_7__3_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_4_), .Q(regfil_7__4_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_5_), .Q(regfil_7__5_));
DFFPOSX1 DFFPOSX1_233 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_6_), .Q(regfil_7__6_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_7_), .Q(regfil_7__7_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_0_), .Q(regfil_3__0_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_1_), .Q(regfil_3__1_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_2_), .Q(regfil_3__2_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_3_), .Q(regfil_3__3_));
DFFPOSX1 DFFPOSX1_239 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_4_), .Q(regfil_3__4_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_1_), .Q(regfil_1__1_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_5_), .Q(regfil_3__5_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_6_), .Q(regfil_3__6_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_7_), .Q(regfil_3__7_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_2_), .Q(regfil_1__2_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_3_), .Q(regfil_1__3_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_4_), .Q(regfil_1__4_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_5_), .Q(regfil_1__5_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_6_), .Q(regfil_1__6_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_2_), .Q(state_2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_7_), .Q(regfil_1__7_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_0_), .Q(regfil_6__0_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_1_), .Q(regfil_6__1_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_2_), .Q(regfil_6__2_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_3_), .Q(regfil_6__3_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_4_), .Q(regfil_6__4_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_5_), .Q(regfil_6__5_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_6_), .Q(regfil_6__6_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_6__0__0__y_16185_7_), .Q(regfil_6__7_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_0_), .Q(regfil_2__0_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_3_), .Q(state_3_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_1_), .Q(regfil_2__1_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_2_), .Q(regfil_2__2_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_3_), .Q(regfil_2__3_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_4_), .Q(regfil_2__4_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_5_), .Q(regfil_2__5_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_6_), .Q(regfil_2__6_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_7_), .Q(regfil_2__7_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_0_), .Q(regfil_0__0_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_1_), .Q(regfil_0__1_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_2_), .Q(regfil_0__2_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_4_), .Q(state_4_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_3_), .Q(regfil_0__3_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_4_), .Q(regfil_0__4_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_5_), .Q(regfil_0__5_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_6_), .Q(regfil_0__6_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_0__0__0__y_15937_7_), .Q(regfil_0__7_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clock), .D(_0writeio_0_0_), .Q(writeio));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clock), .D(_0inta_0_0_), .Q(inta));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clock), .D(_0readio_0_0_), .Q(readio));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clock), .D(_0addr_15_0__0_), .Q(\addr[0] ));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clock), .D(_0addr_15_0__1_), .Q(\addr[1] ));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_5_), .Q(state_5_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clock), .D(_0addr_15_0__2_), .Q(\addr[2] ));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clock), .D(_0addr_15_0__3_), .Q(\addr[3] ));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clock), .D(_0addr_15_0__4_), .Q(\addr[4] ));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clock), .D(_0addr_15_0__5_), .Q(\addr[5] ));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clock), .D(_0addr_15_0__6_), .Q(\addr[6] ));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clock), .D(_0addr_15_0__7_), .Q(\addr[7] ));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clock), .D(_0addr_15_0__8_), .Q(\addr[8] ));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clock), .D(_0addr_15_0__9_), .Q(\addr[9] ));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clock), .D(_0addr_15_0__10_), .Q(\addr[10] ));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clock), .D(_0addr_15_0__11_), .Q(\addr[11] ));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_0_), .Q(regfil_4__0_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clock), .D(_0addr_15_0__12_), .Q(\addr[12] ));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clock), .D(_0addr_15_0__13_), .Q(\addr[13] ));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clock), .D(_0addr_15_0__14_), .Q(\addr[14] ));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clock), .D(_0addr_15_0__15_), .Q(\addr[15] ));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clock), .D(_0readmem_0_0_), .Q(readmem));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clock), .D(_0writemem_0_0_), .Q(writemem));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clock), .D(_0pc_15_0__0_), .Q(pc_0_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clock), .D(_0pc_15_0__1_), .Q(pc_1_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clock), .D(_0pc_15_0__2_), .Q(pc_2_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clock), .D(_0pc_15_0__3_), .Q(pc_3_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_1_), .Q(regfil_4__1_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clock), .D(_0pc_15_0__4_), .Q(pc_4_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(clock), .D(_0pc_15_0__5_), .Q(pc_5_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(clock), .D(_0pc_15_0__6_), .Q(pc_6_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(clock), .D(_0pc_15_0__7_), .Q(pc_7_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(clock), .D(_0pc_15_0__8_), .Q(pc_8_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(clock), .D(_0pc_15_0__9_), .Q(pc_9_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(clock), .D(_0pc_15_0__10_), .Q(pc_10_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(clock), .D(_0pc_15_0__11_), .Q(pc_11_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(clock), .D(_0pc_15_0__12_), .Q(pc_12_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(clock), .D(_0pc_15_0__13_), .Q(pc_13_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_2_), .Q(regfil_4__2_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(clock), .D(_0pc_15_0__14_), .Q(pc_14_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(clock), .D(_0pc_15_0__15_), .Q(pc_15_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(clock), .D(_0sp_15_0__0_), .Q(sp_0_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(clock), .D(_0sp_15_0__1_), .Q(sp_1_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(clock), .D(_0sp_15_0__2_), .Q(sp_2_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(clock), .D(_0sp_15_0__3_), .Q(sp_3_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(clock), .D(_0sp_15_0__4_), .Q(sp_4_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(clock), .D(_0sp_15_0__5_), .Q(sp_5_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(clock), .D(_0sp_15_0__6_), .Q(sp_6_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(clock), .D(_0sp_15_0__7_), .Q(sp_7_));
INVX1 INVX1_1 ( .A(state_5_), .Y(_abc_41356_new_n501_));
INVX1 INVX1_10 ( .A(opcode_5_), .Y(_abc_41356_new_n525_));
INVX1 INVX1_100 ( .A(_abc_41356_new_n1123_), .Y(_abc_41356_new_n1124_));
INVX1 INVX1_101 ( .A(alu_res_6_), .Y(_abc_41356_new_n1125_));
INVX1 INVX1_102 ( .A(_abc_41356_new_n1127_), .Y(_abc_41356_new_n1128_));
INVX1 INVX1_103 ( .A(_abc_41356_new_n1132_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_6_));
INVX1 INVX1_104 ( .A(regfil_0__7_), .Y(_abc_41356_new_n1134_));
INVX1 INVX1_105 ( .A(_abc_41356_new_n1136_), .Y(_abc_41356_new_n1137_));
INVX1 INVX1_106 ( .A(_abc_41356_new_n1139_), .Y(_abc_41356_new_n1140_));
INVX1 INVX1_107 ( .A(_abc_41356_new_n704_), .Y(_abc_41356_new_n1178_));
INVX1 INVX1_108 ( .A(_abc_41356_new_n1191_), .Y(_abc_41356_new_n1192_));
INVX1 INVX1_109 ( .A(_abc_41356_new_n1188_), .Y(_abc_41356_new_n1200_));
INVX1 INVX1_11 ( .A(_abc_41356_new_n531_), .Y(_abc_41356_new_n532_));
INVX1 INVX1_110 ( .A(_abc_41356_new_n1201_), .Y(_abc_41356_new_n1202_));
INVX1 INVX1_111 ( .A(_abc_41356_new_n1207_), .Y(_abc_41356_new_n1208_));
INVX1 INVX1_112 ( .A(_abc_41356_new_n693_), .Y(_abc_41356_new_n1210_));
INVX1 INVX1_113 ( .A(_abc_41356_new_n1212_), .Y(_abc_41356_new_n1213_));
INVX1 INVX1_114 ( .A(_abc_41356_new_n1216_), .Y(_abc_41356_new_n1217_));
INVX1 INVX1_115 ( .A(_abc_41356_new_n1219_), .Y(_abc_41356_new_n1220_));
INVX1 INVX1_116 ( .A(_abc_41356_new_n1230_), .Y(_abc_41356_new_n1231_));
INVX1 INVX1_117 ( .A(_abc_41356_new_n1235_), .Y(_abc_41356_new_n1236_));
INVX1 INVX1_118 ( .A(_abc_41356_new_n1238_), .Y(_abc_41356_new_n1239_));
INVX1 INVX1_119 ( .A(_abc_41356_new_n1229_), .Y(_abc_41356_new_n1248_));
INVX1 INVX1_12 ( .A(regfil_7__0_), .Y(_abc_41356_new_n533_));
INVX1 INVX1_120 ( .A(regfil_4__0_), .Y(_abc_41356_new_n1251_));
INVX1 INVX1_121 ( .A(regfil_5__7_), .Y(_abc_41356_new_n1252_));
INVX1 INVX1_122 ( .A(regfil_5__6_), .Y(_abc_41356_new_n1253_));
INVX1 INVX1_123 ( .A(regfil_5__5_), .Y(_abc_41356_new_n1254_));
INVX1 INVX1_124 ( .A(regfil_5__4_), .Y(_abc_41356_new_n1255_));
INVX1 INVX1_125 ( .A(regfil_5__3_), .Y(_abc_41356_new_n1256_));
INVX1 INVX1_126 ( .A(regfil_5__2_), .Y(_abc_41356_new_n1257_));
INVX1 INVX1_127 ( .A(regfil_5__0_), .Y(_abc_41356_new_n1258_));
INVX1 INVX1_128 ( .A(regfil_5__1_), .Y(_abc_41356_new_n1259_));
INVX1 INVX1_129 ( .A(_abc_41356_new_n1267_), .Y(_abc_41356_new_n1268_));
INVX1 INVX1_13 ( .A(opcode_4_), .Y(_abc_41356_new_n534_));
INVX1 INVX1_130 ( .A(_abc_41356_new_n1271_), .Y(_abc_41356_new_n1272_));
INVX1 INVX1_131 ( .A(_abc_41356_new_n1281_), .Y(_abc_41356_new_n1282_));
INVX1 INVX1_132 ( .A(_abc_41356_new_n1221_), .Y(_abc_41356_new_n1285_));
INVX1 INVX1_133 ( .A(_abc_41356_new_n1288_), .Y(_abc_41356_new_n1289_));
INVX1 INVX1_134 ( .A(_abc_41356_new_n1293_), .Y(_abc_41356_new_n1294_));
INVX1 INVX1_135 ( .A(_abc_41356_new_n1295_), .Y(_abc_41356_new_n1296_));
INVX1 INVX1_136 ( .A(sp_2_), .Y(_abc_41356_new_n1298_));
INVX1 INVX1_137 ( .A(_abc_41356_new_n1300_), .Y(_abc_41356_new_n1301_));
INVX1 INVX1_138 ( .A(sp_3_), .Y(_abc_41356_new_n1303_));
INVX1 INVX1_139 ( .A(_abc_41356_new_n1305_), .Y(_abc_41356_new_n1306_));
INVX1 INVX1_14 ( .A(regfil_7__3_), .Y(_abc_41356_new_n539_));
INVX1 INVX1_140 ( .A(_abc_41356_new_n1312_), .Y(_abc_41356_new_n1313_));
INVX1 INVX1_141 ( .A(sp_7_), .Y(_abc_41356_new_n1314_));
INVX1 INVX1_142 ( .A(_abc_41356_new_n1315_), .Y(_abc_41356_new_n1316_));
INVX1 INVX1_143 ( .A(sp_6_), .Y(_abc_41356_new_n1319_));
INVX1 INVX1_144 ( .A(_abc_41356_new_n1321_), .Y(_abc_41356_new_n1322_));
INVX1 INVX1_145 ( .A(sp_4_), .Y(_abc_41356_new_n1325_));
INVX1 INVX1_146 ( .A(_abc_41356_new_n1327_), .Y(_abc_41356_new_n1328_));
INVX1 INVX1_147 ( .A(_abc_41356_new_n1329_), .Y(_abc_41356_new_n1330_));
INVX1 INVX1_148 ( .A(sp_5_), .Y(_abc_41356_new_n1331_));
INVX1 INVX1_149 ( .A(_abc_41356_new_n1332_), .Y(_abc_41356_new_n1333_));
INVX1 INVX1_15 ( .A(regfil_7__2_), .Y(_abc_41356_new_n540_));
INVX1 INVX1_150 ( .A(sp_8_), .Y(_abc_41356_new_n1345_));
INVX1 INVX1_151 ( .A(_abc_41356_new_n1348_), .Y(_abc_41356_new_n1349_));
INVX1 INVX1_152 ( .A(_abc_41356_new_n1350_), .Y(_abc_41356_new_n1351_));
INVX1 INVX1_153 ( .A(regfil_3__3_), .Y(_abc_41356_new_n1356_));
INVX1 INVX1_154 ( .A(_abc_41356_new_n1358_), .Y(_abc_41356_new_n1359_));
INVX1 INVX1_155 ( .A(_abc_41356_new_n1363_), .Y(_abc_41356_new_n1365_));
INVX1 INVX1_156 ( .A(regfil_3__2_), .Y(_abc_41356_new_n1370_));
INVX1 INVX1_157 ( .A(_abc_41356_new_n1372_), .Y(_abc_41356_new_n1373_));
INVX1 INVX1_158 ( .A(_abc_41356_new_n1377_), .Y(_abc_41356_new_n1378_));
INVX1 INVX1_159 ( .A(_abc_41356_new_n1381_), .Y(_abc_41356_new_n1382_));
INVX1 INVX1_16 ( .A(_abc_41356_new_n542_), .Y(_abc_41356_new_n543_));
INVX1 INVX1_160 ( .A(_abc_41356_new_n1386_), .Y(_abc_41356_new_n1387_));
INVX1 INVX1_161 ( .A(_abc_41356_new_n1390_), .Y(_abc_41356_new_n1391_));
INVX1 INVX1_162 ( .A(_abc_41356_new_n1403_), .Y(_abc_41356_new_n1404_));
INVX1 INVX1_163 ( .A(regfil_2__0_), .Y(_abc_41356_new_n1405_));
INVX1 INVX1_164 ( .A(_abc_41356_new_n1408_), .Y(_abc_41356_new_n1410_));
INVX1 INVX1_165 ( .A(_abc_41356_new_n1419_), .Y(_abc_41356_new_n1420_));
INVX1 INVX1_166 ( .A(_abc_41356_new_n1421_), .Y(_abc_41356_new_n1422_));
INVX1 INVX1_167 ( .A(_abc_41356_new_n1429_), .Y(_abc_41356_new_n1430_));
INVX1 INVX1_168 ( .A(_abc_41356_new_n1433_), .Y(_abc_41356_new_n1434_));
INVX1 INVX1_169 ( .A(_abc_41356_new_n1435_), .Y(_abc_41356_new_n1436_));
INVX1 INVX1_17 ( .A(opcode_3_), .Y(_abc_41356_new_n545_));
INVX1 INVX1_170 ( .A(_abc_41356_new_n1428_), .Y(_abc_41356_new_n1438_));
INVX1 INVX1_171 ( .A(_abc_41356_new_n1440_), .Y(_abc_41356_new_n1441_));
INVX1 INVX1_172 ( .A(_abc_41356_new_n1443_), .Y(_abc_41356_new_n1444_));
INVX1 INVX1_173 ( .A(_abc_41356_new_n1447_), .Y(_abc_41356_new_n1448_));
INVX1 INVX1_174 ( .A(_abc_41356_new_n1452_), .Y(_abc_41356_new_n1453_));
INVX1 INVX1_175 ( .A(_abc_41356_new_n1456_), .Y(_abc_41356_new_n1457_));
INVX1 INVX1_176 ( .A(_abc_41356_new_n1461_), .Y(_abc_41356_new_n1462_));
INVX1 INVX1_177 ( .A(_abc_41356_new_n1469_), .Y(_abc_41356_new_n1470_));
INVX1 INVX1_178 ( .A(_abc_41356_new_n1471_), .Y(_abc_41356_new_n1472_));
INVX1 INVX1_179 ( .A(_abc_41356_new_n1475_), .Y(_abc_41356_new_n1476_));
INVX1 INVX1_18 ( .A(rdatahold_0_), .Y(_abc_41356_new_n564_));
INVX1 INVX1_180 ( .A(_abc_41356_new_n1477_), .Y(_abc_41356_new_n1478_));
INVX1 INVX1_181 ( .A(_abc_41356_new_n1486_), .Y(_abc_41356_new_n1487_));
INVX1 INVX1_182 ( .A(regfil_4__1_), .Y(_abc_41356_new_n1504_));
INVX1 INVX1_183 ( .A(_abc_41356_new_n1511_), .Y(_abc_41356_new_n1512_));
INVX1 INVX1_184 ( .A(sp_9_), .Y(_abc_41356_new_n1515_));
INVX1 INVX1_185 ( .A(_abc_41356_new_n1518_), .Y(_abc_41356_new_n1519_));
INVX1 INVX1_186 ( .A(_abc_41356_new_n1521_), .Y(_abc_41356_new_n1522_));
INVX1 INVX1_187 ( .A(_abc_41356_new_n1526_), .Y(_abc_41356_new_n1527_));
INVX1 INVX1_188 ( .A(regfil_2__1_), .Y(_abc_41356_new_n1532_));
INVX1 INVX1_189 ( .A(_abc_41356_new_n1534_), .Y(_abc_41356_new_n1535_));
INVX1 INVX1_19 ( .A(_abc_41356_new_n565_), .Y(_abc_41356_new_n566_));
INVX1 INVX1_190 ( .A(_abc_41356_new_n1539_), .Y(_abc_41356_new_n1540_));
INVX1 INVX1_191 ( .A(_abc_41356_new_n1541_), .Y(_abc_41356_new_n1542_));
INVX1 INVX1_192 ( .A(regfil_0__1_), .Y(_abc_41356_new_n1546_));
INVX1 INVX1_193 ( .A(_abc_41356_new_n1549_), .Y(_abc_41356_new_n1550_));
INVX1 INVX1_194 ( .A(_abc_41356_new_n1551_), .Y(_abc_41356_new_n1552_));
INVX1 INVX1_195 ( .A(_abc_41356_new_n1556_), .Y(_abc_41356_new_n1557_));
INVX1 INVX1_196 ( .A(_abc_41356_new_n1563_), .Y(_abc_41356_new_n1564_));
INVX1 INVX1_197 ( .A(regfil_4__2_), .Y(_abc_41356_new_n1580_));
INVX1 INVX1_198 ( .A(_abc_41356_new_n1581_), .Y(_abc_41356_new_n1582_));
INVX1 INVX1_199 ( .A(_abc_41356_new_n1585_), .Y(_abc_41356_new_n1586_));
INVX1 INVX1_2 ( .A(state_3_), .Y(_abc_41356_new_n503_));
INVX1 INVX1_20 ( .A(opcode_2_), .Y(_abc_41356_new_n577_));
INVX1 INVX1_200 ( .A(_abc_41356_new_n1588_), .Y(_abc_41356_new_n1589_));
INVX1 INVX1_201 ( .A(_abc_41356_new_n1517_), .Y(_abc_41356_new_n1592_));
INVX1 INVX1_202 ( .A(_abc_41356_new_n1594_), .Y(_abc_41356_new_n1595_));
INVX1 INVX1_203 ( .A(sp_10_), .Y(_abc_41356_new_n1596_));
INVX1 INVX1_204 ( .A(_abc_41356_new_n1599_), .Y(_abc_41356_new_n1600_));
INVX1 INVX1_205 ( .A(_abc_41356_new_n1601_), .Y(_abc_41356_new_n1602_));
INVX1 INVX1_206 ( .A(regfil_2__2_), .Y(_abc_41356_new_n1608_));
INVX1 INVX1_207 ( .A(_abc_41356_new_n1611_), .Y(_abc_41356_new_n1612_));
INVX1 INVX1_208 ( .A(_abc_41356_new_n1613_), .Y(_abc_41356_new_n1614_));
INVX1 INVX1_209 ( .A(_abc_41356_new_n1618_), .Y(_abc_41356_new_n1619_));
INVX1 INVX1_21 ( .A(_abc_41356_new_n582_), .Y(_abc_41356_new_n583_));
INVX1 INVX1_210 ( .A(regfil_0__2_), .Y(_abc_41356_new_n1621_));
INVX1 INVX1_211 ( .A(_abc_41356_new_n1620_), .Y(_abc_41356_new_n1626_));
INVX1 INVX1_212 ( .A(_abc_41356_new_n1624_), .Y(_abc_41356_new_n1627_));
INVX1 INVX1_213 ( .A(_abc_41356_new_n1633_), .Y(_abc_41356_new_n1634_));
INVX1 INVX1_214 ( .A(regfil_4__3_), .Y(_abc_41356_new_n1652_));
INVX1 INVX1_215 ( .A(sp_11_), .Y(_abc_41356_new_n1653_));
INVX1 INVX1_216 ( .A(_abc_41356_new_n1654_), .Y(_abc_41356_new_n1655_));
INVX1 INVX1_217 ( .A(_abc_41356_new_n1656_), .Y(_abc_41356_new_n1657_));
INVX1 INVX1_218 ( .A(_abc_41356_new_n1658_), .Y(_abc_41356_new_n1659_));
INVX1 INVX1_219 ( .A(_abc_41356_new_n1651_), .Y(_abc_41356_new_n1661_));
INVX1 INVX1_22 ( .A(state_2_), .Y(_abc_41356_new_n586_));
INVX1 INVX1_220 ( .A(_abc_41356_new_n1415_), .Y(_abc_41356_new_n1665_));
INVX1 INVX1_221 ( .A(_abc_41356_new_n1667_), .Y(_abc_41356_new_n1668_));
INVX1 INVX1_222 ( .A(regfil_2__3_), .Y(_abc_41356_new_n1669_));
INVX1 INVX1_223 ( .A(_abc_41356_new_n1670_), .Y(_abc_41356_new_n1671_));
INVX1 INVX1_224 ( .A(_abc_41356_new_n1666_), .Y(_abc_41356_new_n1674_));
INVX1 INVX1_225 ( .A(_abc_41356_new_n1672_), .Y(_abc_41356_new_n1675_));
INVX1 INVX1_226 ( .A(_abc_41356_new_n1623_), .Y(_abc_41356_new_n1679_));
INVX1 INVX1_227 ( .A(_abc_41356_new_n1680_), .Y(_abc_41356_new_n1681_));
INVX1 INVX1_228 ( .A(_abc_41356_new_n1682_), .Y(_abc_41356_new_n1683_));
INVX1 INVX1_229 ( .A(regfil_0__3_), .Y(_abc_41356_new_n1684_));
INVX1 INVX1_23 ( .A(popdes_0_), .Y(_abc_41356_new_n590_));
INVX1 INVX1_230 ( .A(_abc_41356_new_n1685_), .Y(_abc_41356_new_n1686_));
INVX1 INVX1_231 ( .A(_abc_41356_new_n1687_), .Y(_abc_41356_new_n1689_));
INVX1 INVX1_232 ( .A(_abc_41356_new_n1699_), .Y(_abc_41356_new_n1700_));
INVX1 INVX1_233 ( .A(_abc_41356_new_n1706_), .Y(_abc_41356_new_n1707_));
INVX1 INVX1_234 ( .A(_abc_41356_new_n1708_), .Y(_abc_41356_new_n1709_));
INVX1 INVX1_235 ( .A(regfil_4__4_), .Y(_abc_41356_new_n1723_));
INVX1 INVX1_236 ( .A(_abc_41356_new_n1593_), .Y(_abc_41356_new_n1732_));
INVX1 INVX1_237 ( .A(sp_12_), .Y(_abc_41356_new_n1738_));
INVX1 INVX1_238 ( .A(_abc_41356_new_n1741_), .Y(_abc_41356_new_n1742_));
INVX1 INVX1_239 ( .A(_abc_41356_new_n1743_), .Y(_abc_41356_new_n1744_));
INVX1 INVX1_24 ( .A(popdes_1_), .Y(_abc_41356_new_n591_));
INVX1 INVX1_240 ( .A(regfil_0__4_), .Y(_abc_41356_new_n1748_));
INVX1 INVX1_241 ( .A(_abc_41356_new_n1751_), .Y(_abc_41356_new_n1752_));
INVX1 INVX1_242 ( .A(_abc_41356_new_n1757_), .Y(_abc_41356_new_n1758_));
INVX1 INVX1_243 ( .A(_abc_41356_new_n1759_), .Y(_abc_41356_new_n1760_));
INVX1 INVX1_244 ( .A(_abc_41356_new_n1762_), .Y(_abc_41356_new_n1763_));
INVX1 INVX1_245 ( .A(_abc_41356_new_n1764_), .Y(_abc_41356_new_n1765_));
INVX1 INVX1_246 ( .A(regfil_2__4_), .Y(_abc_41356_new_n1777_));
INVX1 INVX1_247 ( .A(_abc_41356_new_n1780_), .Y(_abc_41356_new_n1781_));
INVX1 INVX1_248 ( .A(_abc_41356_new_n1782_), .Y(_abc_41356_new_n1783_));
INVX1 INVX1_249 ( .A(_abc_41356_new_n1789_), .Y(_abc_41356_new_n1790_));
INVX1 INVX1_25 ( .A(_abc_41356_new_n595_), .Y(_abc_41356_new_n596_));
INVX1 INVX1_250 ( .A(_abc_41356_new_n1803_), .Y(_abc_41356_new_n1804_));
INVX1 INVX1_251 ( .A(regfil_4__5_), .Y(_abc_41356_new_n1819_));
INVX1 INVX1_252 ( .A(_abc_41356_new_n1724_), .Y(_abc_41356_new_n1821_));
INVX1 INVX1_253 ( .A(sp_13_), .Y(_abc_41356_new_n1826_));
INVX1 INVX1_254 ( .A(_abc_41356_new_n1829_), .Y(_abc_41356_new_n1830_));
INVX1 INVX1_255 ( .A(_abc_41356_new_n1831_), .Y(_abc_41356_new_n1832_));
INVX1 INVX1_256 ( .A(_abc_41356_new_n1836_), .Y(_abc_41356_new_n1837_));
INVX1 INVX1_257 ( .A(regfil_2__5_), .Y(_abc_41356_new_n1842_));
INVX1 INVX1_258 ( .A(_abc_41356_new_n1845_), .Y(_abc_41356_new_n1846_));
INVX1 INVX1_259 ( .A(_abc_41356_new_n1850_), .Y(_abc_41356_new_n1851_));
INVX1 INVX1_26 ( .A(_abc_41356_new_n581_), .Y(_abc_41356_new_n597_));
INVX1 INVX1_260 ( .A(_abc_41356_new_n1853_), .Y(_abc_41356_new_n1854_));
INVX1 INVX1_261 ( .A(regfil_0__5_), .Y(_abc_41356_new_n1857_));
INVX1 INVX1_262 ( .A(_abc_41356_new_n1860_), .Y(_abc_41356_new_n1861_));
INVX1 INVX1_263 ( .A(_abc_41356_new_n1862_), .Y(_abc_41356_new_n1863_));
INVX1 INVX1_264 ( .A(_abc_41356_new_n1867_), .Y(_abc_41356_new_n1868_));
INVX1 INVX1_265 ( .A(_abc_41356_new_n1877_), .Y(_abc_41356_new_n1878_));
INVX1 INVX1_266 ( .A(regfil_4__6_), .Y(_abc_41356_new_n1893_));
INVX1 INVX1_267 ( .A(_abc_41356_new_n1820_), .Y(_abc_41356_new_n1895_));
INVX1 INVX1_268 ( .A(sp_14_), .Y(_abc_41356_new_n1902_));
INVX1 INVX1_269 ( .A(_abc_41356_new_n1905_), .Y(_abc_41356_new_n1906_));
INVX1 INVX1_27 ( .A(_abc_41356_new_n601_), .Y(_abc_41356_new_n602_));
INVX1 INVX1_270 ( .A(_abc_41356_new_n1908_), .Y(_abc_41356_new_n1909_));
INVX1 INVX1_271 ( .A(_abc_41356_new_n1912_), .Y(_abc_41356_new_n1913_));
INVX1 INVX1_272 ( .A(_abc_41356_new_n1914_), .Y(_abc_41356_new_n1915_));
INVX1 INVX1_273 ( .A(_abc_41356_new_n1918_), .Y(_abc_41356_new_n1919_));
INVX1 INVX1_274 ( .A(regfil_2__6_), .Y(_abc_41356_new_n1926_));
INVX1 INVX1_275 ( .A(_abc_41356_new_n1929_), .Y(_abc_41356_new_n1930_));
INVX1 INVX1_276 ( .A(_abc_41356_new_n1931_), .Y(_abc_41356_new_n1932_));
INVX1 INVX1_277 ( .A(_abc_41356_new_n1938_), .Y(_abc_41356_new_n1939_));
INVX1 INVX1_278 ( .A(_abc_41356_new_n1944_), .Y(_abc_41356_new_n1945_));
INVX1 INVX1_279 ( .A(regfil_4__7_), .Y(_abc_41356_new_n1961_));
INVX1 INVX1_28 ( .A(_abc_41356_new_n608_), .Y(_abc_41356_new_n609_));
INVX1 INVX1_280 ( .A(_abc_41356_new_n1894_), .Y(_abc_41356_new_n1962_));
INVX1 INVX1_281 ( .A(sp_15_), .Y(_abc_41356_new_n1967_));
INVX1 INVX1_282 ( .A(_abc_41356_new_n1966_), .Y(_abc_41356_new_n1972_));
INVX1 INVX1_283 ( .A(_abc_41356_new_n1970_), .Y(_abc_41356_new_n1973_));
INVX1 INVX1_284 ( .A(_abc_41356_new_n1982_), .Y(_abc_41356_new_n1983_));
INVX1 INVX1_285 ( .A(_abc_41356_new_n1917_), .Y(_abc_41356_new_n1989_));
INVX1 INVX1_286 ( .A(_abc_41356_new_n1994_), .Y(_abc_41356_new_n1995_));
INVX1 INVX1_287 ( .A(regfil_2__7_), .Y(_abc_41356_new_n1996_));
INVX1 INVX1_288 ( .A(_abc_41356_new_n1999_), .Y(_abc_41356_new_n2002_));
INVX1 INVX1_289 ( .A(_abc_41356_new_n2009_), .Y(_abc_41356_new_n2010_));
INVX1 INVX1_29 ( .A(_abc_41356_new_n612_), .Y(_abc_41356_new_n613_));
INVX1 INVX1_290 ( .A(_abc_41356_new_n523_), .Y(_abc_41356_new_n2020_));
INVX1 INVX1_291 ( .A(_abc_41356_new_n516_), .Y(_abc_41356_new_n2021_));
INVX1 INVX1_292 ( .A(_abc_41356_new_n1232_), .Y(_abc_41356_new_n2022_));
INVX1 INVX1_293 ( .A(_abc_41356_new_n2027_), .Y(_abc_41356_new_n2028_));
INVX1 INVX1_294 ( .A(pc_8_), .Y(_abc_41356_new_n2041_));
INVX1 INVX1_295 ( .A(_abc_41356_new_n2039_), .Y(_abc_41356_new_n2042_));
INVX1 INVX1_296 ( .A(_abc_41356_new_n2044_), .Y(_abc_41356_new_n2045_));
INVX1 INVX1_297 ( .A(intcyc), .Y(_abc_41356_new_n2049_));
INVX1 INVX1_298 ( .A(_abc_41356_new_n2046_), .Y(_abc_41356_new_n2054_));
INVX1 INVX1_299 ( .A(_abc_41356_new_n535_), .Y(_abc_41356_new_n2056_));
INVX1 INVX1_3 ( .A(state_1_), .Y(_abc_41356_new_n505_));
INVX1 INVX1_30 ( .A(opcode_1_), .Y(_abc_41356_new_n615_));
INVX1 INVX1_300 ( .A(_abc_41356_new_n2060_), .Y(_abc_41356_new_n2061_));
INVX1 INVX1_301 ( .A(_abc_41356_new_n1218_), .Y(_abc_41356_new_n2063_));
INVX1 INVX1_302 ( .A(_abc_41356_new_n2048_), .Y(_abc_41356_new_n2064_));
INVX1 INVX1_303 ( .A(_abc_41356_new_n2065_), .Y(_abc_41356_new_n2066_));
INVX1 INVX1_304 ( .A(_abc_41356_new_n2073_), .Y(_abc_41356_new_n2074_));
INVX1 INVX1_305 ( .A(_abc_41356_new_n2077_), .Y(_abc_41356_new_n2078_));
INVX1 INVX1_306 ( .A(_abc_41356_new_n2069_), .Y(_abc_41356_new_n2096_));
INVX1 INVX1_307 ( .A(_abc_41356_new_n2108_), .Y(_abc_41356_new_n2109_));
INVX1 INVX1_308 ( .A(_abc_41356_new_n2117_), .Y(_abc_41356_new_n2118_));
INVX1 INVX1_309 ( .A(pc_10_), .Y(_abc_41356_new_n2149_));
INVX1 INVX1_31 ( .A(opcode_0_), .Y(_abc_41356_new_n618_));
INVX1 INVX1_310 ( .A(_abc_41356_new_n2151_), .Y(_abc_41356_new_n2152_));
INVX1 INVX1_311 ( .A(_abc_41356_new_n2159_), .Y(_abc_41356_new_n2160_));
INVX1 INVX1_312 ( .A(_abc_41356_new_n2188_), .Y(_abc_41356_new_n2189_));
INVX1 INVX1_313 ( .A(_abc_41356_new_n2197_), .Y(_abc_41356_new_n2198_));
INVX1 INVX1_314 ( .A(pc_12_), .Y(_abc_41356_new_n2227_));
INVX1 INVX1_315 ( .A(_abc_41356_new_n2229_), .Y(_abc_41356_new_n2230_));
INVX1 INVX1_316 ( .A(_abc_41356_new_n2237_), .Y(_abc_41356_new_n2238_));
INVX1 INVX1_317 ( .A(_abc_41356_new_n2266_), .Y(_abc_41356_new_n2267_));
INVX1 INVX1_318 ( .A(_abc_41356_new_n2275_), .Y(_abc_41356_new_n2276_));
INVX1 INVX1_319 ( .A(_abc_41356_new_n2304_), .Y(_abc_41356_new_n2305_));
INVX1 INVX1_32 ( .A(regfil_0__0_), .Y(_abc_41356_new_n644_));
INVX1 INVX1_320 ( .A(_abc_41356_new_n2313_), .Y(_abc_41356_new_n2314_));
INVX1 INVX1_321 ( .A(_abc_41356_new_n2343_), .Y(_abc_41356_new_n2344_));
INVX1 INVX1_322 ( .A(_abc_41356_new_n2351_), .Y(_abc_41356_new_n2352_));
INVX1 INVX1_323 ( .A(regfil_3__0_), .Y(_abc_41356_new_n2375_));
INVX1 INVX1_324 ( .A(_abc_41356_new_n668_), .Y(_abc_41356_new_n2383_));
INVX1 INVX1_325 ( .A(_abc_41356_new_n2385_), .Y(_abc_41356_new_n2386_));
INVX1 INVX1_326 ( .A(_abc_41356_new_n2395_), .Y(_abc_41356_new_n2396_));
INVX1 INVX1_327 ( .A(regfil_3__1_), .Y(_abc_41356_new_n2409_));
INVX1 INVX1_328 ( .A(_abc_41356_new_n2411_), .Y(_abc_41356_new_n2414_));
INVX1 INVX1_329 ( .A(_abc_41356_new_n2421_), .Y(_abc_41356_new_n2422_));
INVX1 INVX1_33 ( .A(regfil_1__3_), .Y(_abc_41356_new_n645_));
INVX1 INVX1_330 ( .A(_abc_41356_new_n2410_), .Y(_abc_41356_new_n2434_));
INVX1 INVX1_331 ( .A(_abc_41356_new_n2439_), .Y(_abc_41356_new_n2440_));
INVX1 INVX1_332 ( .A(_abc_41356_new_n2433_), .Y(_abc_41356_new_n2454_));
INVX1 INVX1_333 ( .A(_abc_41356_new_n2459_), .Y(_abc_41356_new_n2460_));
INVX1 INVX1_334 ( .A(_abc_41356_new_n2453_), .Y(_abc_41356_new_n2473_));
INVX1 INVX1_335 ( .A(_abc_41356_new_n2474_), .Y(_abc_41356_new_n2475_));
INVX1 INVX1_336 ( .A(_abc_41356_new_n2480_), .Y(_abc_41356_new_n2481_));
INVX1 INVX1_337 ( .A(_abc_41356_new_n2494_), .Y(_abc_41356_new_n2495_));
INVX1 INVX1_338 ( .A(_abc_41356_new_n2499_), .Y(_abc_41356_new_n2500_));
INVX1 INVX1_339 ( .A(_abc_41356_new_n2514_), .Y(_abc_41356_new_n2515_));
INVX1 INVX1_34 ( .A(regfil_1__2_), .Y(_abc_41356_new_n646_));
INVX1 INVX1_340 ( .A(_abc_41356_new_n2519_), .Y(_abc_41356_new_n2520_));
INVX1 INVX1_341 ( .A(_abc_41356_new_n2534_), .Y(_abc_41356_new_n2535_));
INVX1 INVX1_342 ( .A(_abc_41356_new_n2540_), .Y(_abc_41356_new_n2541_));
INVX1 INVX1_343 ( .A(_abc_41356_new_n2550_), .Y(_abc_41356_new_n2551_));
INVX1 INVX1_344 ( .A(_abc_41356_new_n2556_), .Y(_abc_41356_new_n2557_));
INVX1 INVX1_345 ( .A(_abc_41356_new_n2567_), .Y(_abc_41356_new_n2569_));
INVX1 INVX1_346 ( .A(_abc_41356_new_n649_), .Y(_abc_41356_new_n2580_));
INVX1 INVX1_347 ( .A(_abc_41356_new_n569_), .Y(_abc_41356_new_n2584_));
INVX1 INVX1_348 ( .A(_abc_41356_new_n650_), .Y(_abc_41356_new_n2596_));
INVX1 INVX1_349 ( .A(_abc_41356_new_n570_), .Y(_abc_41356_new_n2600_));
INVX1 INVX1_35 ( .A(regfil_1__0_), .Y(_abc_41356_new_n647_));
INVX1 INVX1_350 ( .A(_abc_41356_new_n653_), .Y(_abc_41356_new_n2612_));
INVX1 INVX1_351 ( .A(_abc_41356_new_n571_), .Y(_abc_41356_new_n2616_));
INVX1 INVX1_352 ( .A(_abc_41356_new_n654_), .Y(_abc_41356_new_n2628_));
INVX1 INVX1_353 ( .A(_abc_41356_new_n572_), .Y(_abc_41356_new_n2632_));
INVX1 INVX1_354 ( .A(_abc_41356_new_n655_), .Y(_abc_41356_new_n2645_));
INVX1 INVX1_355 ( .A(_abc_41356_new_n573_), .Y(_abc_41356_new_n2650_));
INVX1 INVX1_356 ( .A(_abc_41356_new_n574_), .Y(_abc_41356_new_n2665_));
INVX1 INVX1_357 ( .A(_abc_41356_new_n2671_), .Y(_abc_41356_new_n2672_));
INVX1 INVX1_358 ( .A(_abc_41356_new_n2697_), .Y(_abc_41356_new_n2698_));
INVX1 INVX1_359 ( .A(_abc_41356_new_n2704_), .Y(_abc_41356_new_n2705_));
INVX1 INVX1_36 ( .A(regfil_1__1_), .Y(_abc_41356_new_n648_));
INVX1 INVX1_360 ( .A(_abc_41356_new_n2710_), .Y(_abc_41356_new_n2711_));
INVX1 INVX1_361 ( .A(_abc_41356_new_n2724_), .Y(_abc_41356_new_n2725_));
INVX1 INVX1_362 ( .A(_abc_41356_new_n2730_), .Y(_abc_41356_new_n2731_));
INVX1 INVX1_363 ( .A(_abc_41356_new_n2744_), .Y(_abc_41356_new_n2745_));
INVX1 INVX1_364 ( .A(_abc_41356_new_n2750_), .Y(_abc_41356_new_n2751_));
INVX1 INVX1_365 ( .A(_abc_41356_new_n2764_), .Y(_abc_41356_new_n2765_));
INVX1 INVX1_366 ( .A(_abc_41356_new_n2769_), .Y(_abc_41356_new_n2770_));
INVX1 INVX1_367 ( .A(_abc_41356_new_n2786_), .Y(_abc_41356_new_n2787_));
INVX1 INVX1_368 ( .A(_abc_41356_new_n2791_), .Y(_abc_41356_new_n2792_));
INVX1 INVX1_369 ( .A(_abc_41356_new_n2808_), .Y(_abc_41356_new_n2809_));
INVX1 INVX1_37 ( .A(_abc_41356_new_n651_), .Y(_abc_41356_new_n652_));
INVX1 INVX1_370 ( .A(_abc_41356_new_n2813_), .Y(_abc_41356_new_n2814_));
INVX1 INVX1_371 ( .A(_abc_41356_new_n2831_), .Y(_abc_41356_new_n2832_));
INVX1 INVX1_372 ( .A(_abc_41356_new_n2835_), .Y(_abc_41356_new_n2836_));
INVX1 INVX1_373 ( .A(_abc_41356_new_n1173_), .Y(_abc_41356_new_n2847_));
INVX1 INVX1_374 ( .A(rdatahold_7_), .Y(_abc_41356_new_n2852_));
INVX1 INVX1_375 ( .A(_abc_41356_new_n2393_), .Y(_abc_41356_new_n2853_));
INVX1 INVX1_376 ( .A(_abc_41356_new_n2855_), .Y(_abc_41356_new_n2856_));
INVX1 INVX1_377 ( .A(_abc_41356_new_n2857_), .Y(_abc_41356_new_n2858_));
INVX1 INVX1_378 ( .A(_abc_41356_new_n2412_), .Y(_abc_41356_new_n2861_));
INVX1 INVX1_379 ( .A(_abc_41356_new_n2833_), .Y(_abc_41356_new_n2863_));
INVX1 INVX1_38 ( .A(_abc_41356_new_n656_), .Y(_abc_41356_new_n657_));
INVX1 INVX1_380 ( .A(_abc_41356_new_n2872_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_7_));
INVX1 INVX1_381 ( .A(_abc_41356_new_n2874_), .Y(_abc_41356_new_n2875_));
INVX1 INVX1_382 ( .A(_abc_41356_new_n2876_), .Y(_abc_41356_new_n2877_));
INVX1 INVX1_383 ( .A(_abc_41356_new_n679_), .Y(_abc_41356_new_n2878_));
INVX1 INVX1_384 ( .A(_abc_41356_new_n2883_), .Y(_abc_41356_new_n2884_));
INVX1 INVX1_385 ( .A(_abc_41356_new_n2886_), .Y(_abc_41356_new_n2887_));
INVX1 INVX1_386 ( .A(_abc_41356_new_n2888_), .Y(_abc_41356_new_n2889_));
INVX1 INVX1_387 ( .A(_abc_41356_new_n2890_), .Y(_abc_41356_new_n2891_));
INVX1 INVX1_388 ( .A(_abc_41356_new_n2879_), .Y(_abc_41356_new_n2906_));
INVX1 INVX1_389 ( .A(_abc_41356_new_n2880_), .Y(_abc_41356_new_n2909_));
INVX1 INVX1_39 ( .A(_abc_41356_new_n665_), .Y(_abc_41356_new_n666_));
INVX1 INVX1_390 ( .A(_abc_41356_new_n2919_), .Y(_abc_41356_new_n2921_));
INVX1 INVX1_391 ( .A(_abc_41356_new_n2924_), .Y(_abc_41356_new_n2925_));
INVX1 INVX1_392 ( .A(_abc_41356_new_n2927_), .Y(_abc_41356_new_n2928_));
INVX1 INVX1_393 ( .A(_abc_41356_new_n2929_), .Y(_abc_41356_new_n2930_));
INVX1 INVX1_394 ( .A(_abc_41356_new_n2931_), .Y(_abc_41356_new_n2933_));
INVX1 INVX1_395 ( .A(_abc_41356_new_n2939_), .Y(_abc_41356_new_n2940_));
INVX1 INVX1_396 ( .A(_abc_41356_new_n3015_), .Y(_abc_41356_new_n3017_));
INVX1 INVX1_397 ( .A(_abc_41356_new_n2926_), .Y(_abc_41356_new_n3200_));
INVX1 INVX1_398 ( .A(_abc_41356_new_n518_), .Y(_abc_41356_new_n3201_));
INVX1 INVX1_399 ( .A(_abc_41356_new_n508_), .Y(_abc_41356_new_n3209_));
INVX1 INVX1_4 ( .A(reset), .Y(_abc_41356_new_n509_));
INVX1 INVX1_40 ( .A(_abc_41356_new_n670_), .Y(_abc_41356_new_n671_));
INVX1 INVX1_400 ( .A(_abc_41356_new_n3212_), .Y(_abc_41356_new_n3213_));
INVX1 INVX1_401 ( .A(_abc_41356_new_n510_), .Y(_abc_41356_new_n3219_));
INVX1 INVX1_402 ( .A(rdatahold2_7_), .Y(_abc_41356_new_n3236_));
INVX1 INVX1_403 ( .A(_abc_41356_new_n3237_), .Y(_abc_41356_new_n3238_));
INVX1 INVX1_404 ( .A(_abc_41356_new_n549_), .Y(_abc_41356_new_n3248_));
INVX1 INVX1_405 ( .A(_abc_41356_new_n676_), .Y(_abc_41356_new_n3265_));
INVX1 INVX1_406 ( .A(_abc_41356_new_n711_), .Y(_abc_41356_new_n3268_));
INVX1 INVX1_407 ( .A(_abc_41356_new_n1997_), .Y(_abc_41356_new_n3276_));
INVX1 INVX1_408 ( .A(carry), .Y(_abc_41356_new_n3279_));
INVX1 INVX1_409 ( .A(_abc_41356_new_n1968_), .Y(_abc_41356_new_n3291_));
INVX1 INVX1_41 ( .A(_abc_41356_new_n604_), .Y(_abc_41356_new_n674_));
INVX1 INVX1_410 ( .A(_abc_41356_new_n1237_), .Y(_abc_41356_new_n3295_));
INVX1 INVX1_411 ( .A(_abc_41356_new_n2058_), .Y(_abc_41356_new_n3296_));
INVX1 INVX1_412 ( .A(_abc_41356_new_n3319_), .Y(_abc_41356_new_n3321_));
INVX1 INVX1_413 ( .A(_abc_41356_new_n3205_), .Y(_abc_41356_new_n3345_));
INVX1 INVX1_414 ( .A(_abc_41356_new_n1481_), .Y(_abc_41356_new_n3353_));
INVX1 INVX1_415 ( .A(_abc_41356_new_n3354_), .Y(_abc_41356_new_n3355_));
INVX1 INVX1_416 ( .A(_abc_41356_new_n2377_), .Y(_abc_41356_new_n3357_));
INVX1 INVX1_417 ( .A(_abc_41356_new_n3361_), .Y(_abc_41356_new_n3362_));
INVX1 INVX1_418 ( .A(_abc_41356_new_n2994_), .Y(_abc_41356_new_n3366_));
INVX1 INVX1_419 ( .A(_abc_41356_new_n3378_), .Y(_abc_41356_new_n3379_));
INVX1 INVX1_42 ( .A(_abc_41356_new_n614_), .Y(_abc_41356_new_n675_));
INVX1 INVX1_420 ( .A(_abc_41356_new_n3364_), .Y(_abc_41356_new_n3384_));
INVX1 INVX1_421 ( .A(_abc_41356_new_n3365_), .Y(_abc_41356_new_n3386_));
INVX1 INVX1_422 ( .A(_abc_41356_new_n3400_), .Y(_abc_41356_new_n3401_));
INVX1 INVX1_423 ( .A(_abc_41356_new_n3408_), .Y(_abc_41356_new_n3409_));
INVX1 INVX1_424 ( .A(_abc_41356_new_n3438_), .Y(_abc_41356_new_n3439_));
INVX1 INVX1_425 ( .A(_abc_41356_new_n3440_), .Y(_abc_41356_new_n3441_));
INVX1 INVX1_426 ( .A(statesel_0_), .Y(_abc_41356_new_n3449_));
INVX1 INVX1_427 ( .A(_abc_41356_new_n3451_), .Y(_abc_41356_new_n3452_));
INVX1 INVX1_428 ( .A(_abc_41356_new_n3453_), .Y(_abc_41356_new_n3454_));
INVX1 INVX1_429 ( .A(_abc_41356_new_n3411_), .Y(_abc_41356_new_n3475_));
INVX1 INVX1_43 ( .A(_abc_41356_new_n677_), .Y(_abc_41356_new_n678_));
INVX1 INVX1_430 ( .A(statesel_1_), .Y(_abc_41356_new_n3488_));
INVX1 INVX1_431 ( .A(_abc_41356_new_n3494_), .Y(_abc_41356_new_n3495_));
INVX1 INVX1_432 ( .A(_abc_41356_new_n3521_), .Y(_abc_41356_new_n3522_));
INVX1 INVX1_433 ( .A(_abc_41356_new_n3356_), .Y(_abc_41356_new_n3533_));
INVX1 INVX1_434 ( .A(_abc_41356_new_n3380_), .Y(_abc_41356_new_n3534_));
INVX1 INVX1_435 ( .A(statesel_3_), .Y(_abc_41356_new_n3553_));
INVX1 INVX1_436 ( .A(_abc_41356_new_n3360_), .Y(_abc_41356_new_n3566_));
INVX1 INVX1_437 ( .A(_abc_41356_new_n3583_), .Y(_abc_41356_new_n3584_));
INVX1 INVX1_438 ( .A(statesel_5_), .Y(_abc_41356_new_n3594_));
INVX1 INVX1_439 ( .A(_abc_41356_new_n3595_), .Y(_abc_41356_new_n3596_));
INVX1 INVX1_44 ( .A(_abc_41356_new_n682_), .Y(_abc_41356_new_n683_));
INVX1 INVX1_440 ( .A(_abc_41356_new_n3615_), .Y(_abc_41356_new_n3616_));
INVX1 INVX1_441 ( .A(_abc_41356_new_n3625_), .Y(_abc_41356_new_n3626_));
INVX1 INVX1_442 ( .A(rdatahold_1_), .Y(_abc_41356_new_n3629_));
INVX1 INVX1_443 ( .A(_abc_41356_new_n3630_), .Y(_abc_41356_new_n3631_));
INVX1 INVX1_444 ( .A(_abc_41356_new_n3634_), .Y(_abc_41356_new_n3635_));
INVX1 INVX1_445 ( .A(_abc_41356_new_n3638_), .Y(_abc_41356_new_n3639_));
INVX1 INVX1_446 ( .A(rdatahold_4_), .Y(_abc_41356_new_n3642_));
INVX1 INVX1_447 ( .A(_abc_41356_new_n3643_), .Y(_abc_41356_new_n3644_));
INVX1 INVX1_448 ( .A(_abc_41356_new_n3647_), .Y(_abc_41356_new_n3648_));
INVX1 INVX1_449 ( .A(_abc_41356_new_n3651_), .Y(_abc_41356_new_n3652_));
INVX1 INVX1_45 ( .A(_abc_41356_new_n689_), .Y(_abc_41356_new_n690_));
INVX1 INVX1_450 ( .A(_abc_41356_new_n3655_), .Y(_abc_41356_new_n3656_));
INVX1 INVX1_451 ( .A(\data[0] ), .Y(_abc_41356_new_n3659_));
INVX1 INVX1_452 ( .A(_abc_41356_new_n3660_), .Y(_abc_41356_new_n3661_));
INVX1 INVX1_453 ( .A(\data[1] ), .Y(_abc_41356_new_n3664_));
INVX1 INVX1_454 ( .A(_abc_41356_new_n3665_), .Y(_abc_41356_new_n3666_));
INVX1 INVX1_455 ( .A(\data[2] ), .Y(_abc_41356_new_n3669_));
INVX1 INVX1_456 ( .A(_abc_41356_new_n3670_), .Y(_abc_41356_new_n3671_));
INVX1 INVX1_457 ( .A(\data[3] ), .Y(_abc_41356_new_n3674_));
INVX1 INVX1_458 ( .A(_abc_41356_new_n3675_), .Y(_abc_41356_new_n3676_));
INVX1 INVX1_459 ( .A(\data[4] ), .Y(_abc_41356_new_n3679_));
INVX1 INVX1_46 ( .A(_abc_41356_new_n695_), .Y(_abc_41356_new_n696_));
INVX1 INVX1_460 ( .A(_abc_41356_new_n3680_), .Y(_abc_41356_new_n3681_));
INVX1 INVX1_461 ( .A(\data[5] ), .Y(_abc_41356_new_n3684_));
INVX1 INVX1_462 ( .A(_abc_41356_new_n3685_), .Y(_abc_41356_new_n3686_));
INVX1 INVX1_463 ( .A(\data[6] ), .Y(_abc_41356_new_n3689_));
INVX1 INVX1_464 ( .A(_abc_41356_new_n3690_), .Y(_abc_41356_new_n3691_));
INVX1 INVX1_465 ( .A(\data[7] ), .Y(_abc_41356_new_n3694_));
INVX1 INVX1_466 ( .A(_abc_41356_new_n3695_), .Y(_abc_41356_new_n3696_));
INVX1 INVX1_467 ( .A(_abc_41356_new_n3698_), .Y(_abc_41356_new_n3699_));
INVX1 INVX1_468 ( .A(_abc_41356_new_n3430_), .Y(_abc_41356_new_n3701_));
INVX1 INVX1_469 ( .A(_abc_41356_new_n3427_), .Y(_abc_41356_new_n3702_));
INVX1 INVX1_47 ( .A(regfil_7__6_), .Y(_abc_41356_new_n700_));
INVX1 INVX1_470 ( .A(_abc_41356_new_n2026_), .Y(_abc_41356_new_n3710_));
INVX1 INVX1_471 ( .A(pc_0_), .Y(_abc_41356_new_n3723_));
INVX1 INVX1_472 ( .A(_abc_41356_new_n2062_), .Y(_abc_41356_new_n3724_));
INVX1 INVX1_473 ( .A(_abc_41356_new_n576_), .Y(_abc_41356_new_n3735_));
INVX1 INVX1_474 ( .A(_abc_41356_new_n3760_), .Y(_abc_41356_new_n3761_));
INVX1 INVX1_475 ( .A(_abc_41356_new_n3762_), .Y(_abc_41356_new_n3764_));
INVX1 INVX1_476 ( .A(pc_2_), .Y(_abc_41356_new_n3811_));
INVX1 INVX1_477 ( .A(_abc_41356_new_n3813_), .Y(_abc_41356_new_n3814_));
INVX1 INVX1_478 ( .A(pc_1_), .Y(_abc_41356_new_n3817_));
INVX1 INVX1_479 ( .A(_abc_41356_new_n3820_), .Y(_abc_41356_new_n3821_));
INVX1 INVX1_48 ( .A(regfil_7__5_), .Y(_abc_41356_new_n701_));
INVX1 INVX1_480 ( .A(_abc_41356_new_n2072_), .Y(_abc_41356_new_n3877_));
INVX1 INVX1_481 ( .A(_abc_41356_new_n2035_), .Y(_abc_41356_new_n3881_));
INVX1 INVX1_482 ( .A(_abc_41356_new_n3926_), .Y(_abc_41356_new_n3927_));
INVX1 INVX1_483 ( .A(_abc_41356_new_n3931_), .Y(_abc_41356_new_n3932_));
INVX1 INVX1_484 ( .A(pc_5_), .Y(_abc_41356_new_n3980_));
INVX1 INVX1_485 ( .A(_abc_41356_new_n3982_), .Y(_abc_41356_new_n3983_));
INVX1 INVX1_486 ( .A(_abc_41356_new_n3987_), .Y(_abc_41356_new_n3988_));
INVX1 INVX1_487 ( .A(_abc_41356_new_n4020_), .Y(_abc_41356_new_n4021_));
INVX1 INVX1_488 ( .A(_abc_41356_new_n4025_), .Y(_abc_41356_new_n4026_));
INVX1 INVX1_489 ( .A(pc_7_), .Y(_abc_41356_new_n4072_));
INVX1 INVX1_49 ( .A(_abc_41356_new_n702_), .Y(_abc_41356_new_n703_));
INVX1 INVX1_490 ( .A(_abc_41356_new_n4074_), .Y(_abc_41356_new_n4075_));
INVX1 INVX1_491 ( .A(_abc_41356_new_n4117_), .Y(_abc_41356_new_n4118_));
INVX1 INVX1_492 ( .A(_abc_41356_new_n3424_), .Y(_abc_41356_new_n4119_));
INVX1 INVX1_493 ( .A(_abc_41356_new_n4124_), .Y(_abc_41356_new_n4125_));
INVX1 INVX1_494 ( .A(_abc_41356_new_n4126_), .Y(_abc_41356_new_n4127_));
INVX1 INVX1_495 ( .A(_abc_41356_new_n4128_), .Y(_abc_41356_new_n4129_));
INVX1 INVX1_496 ( .A(_abc_41356_new_n4131_), .Y(_abc_41356_new_n4132_));
INVX1 INVX1_497 ( .A(_abc_41356_new_n4130_), .Y(_abc_41356_new_n4143_));
INVX1 INVX1_498 ( .A(_abc_41356_new_n4148_), .Y(_abc_41356_new_n4149_));
INVX1 INVX1_499 ( .A(_abc_41356_new_n2989_), .Y(_abc_41356_new_n4151_));
INVX1 INVX1_5 ( .A(regfil_7__1_), .Y(_abc_41356_new_n513_));
INVX1 INVX1_50 ( .A(waitr), .Y(_abc_41356_new_n716_));
INVX1 INVX1_500 ( .A(_abc_41356_new_n4158_), .Y(_abc_41356_new_n4159_));
INVX1 INVX1_501 ( .A(_abc_41356_new_n2997_), .Y(_abc_41356_new_n4160_));
INVX1 INVX1_502 ( .A(_abc_41356_new_n2992_), .Y(_abc_41356_new_n4161_));
INVX1 INVX1_503 ( .A(_abc_41356_new_n4162_), .Y(_abc_41356_new_n4163_));
INVX1 INVX1_504 ( .A(_abc_41356_new_n4164_), .Y(_abc_41356_new_n4165_));
INVX1 INVX1_505 ( .A(_abc_41356_new_n4168_), .Y(_abc_41356_new_n4173_));
INVX1 INVX1_506 ( .A(_abc_41356_new_n4170_), .Y(_abc_41356_new_n4175_));
INVX1 INVX1_507 ( .A(_abc_41356_new_n4184_), .Y(_abc_41356_new_n4185_));
INVX1 INVX1_508 ( .A(raddrhold_0_), .Y(_abc_41356_new_n4196_));
INVX1 INVX1_509 ( .A(_abc_41356_new_n4202_), .Y(_abc_41356_new_n4203_));
INVX1 INVX1_51 ( .A(_abc_41356_new_n723_), .Y(_abc_41356_new_n724_));
INVX1 INVX1_510 ( .A(_abc_41356_new_n4238_), .Y(_abc_41356_new_n4239_));
INVX1 INVX1_511 ( .A(_abc_41356_new_n4245_), .Y(_abc_41356_new_n4246_));
INVX1 INVX1_512 ( .A(_abc_41356_new_n4282_), .Y(_abc_41356_new_n4283_));
INVX1 INVX1_513 ( .A(_abc_41356_new_n4289_), .Y(_abc_41356_new_n4290_));
INVX1 INVX1_514 ( .A(_abc_41356_new_n4321_), .Y(_abc_41356_new_n4322_));
INVX1 INVX1_515 ( .A(_abc_41356_new_n4332_), .Y(_abc_41356_new_n4333_));
INVX1 INVX1_516 ( .A(_abc_41356_new_n4364_), .Y(_abc_41356_new_n4365_));
INVX1 INVX1_517 ( .A(_abc_41356_new_n4375_), .Y(_abc_41356_new_n4376_));
INVX1 INVX1_518 ( .A(_abc_41356_new_n4407_), .Y(_abc_41356_new_n4408_));
INVX1 INVX1_519 ( .A(_abc_41356_new_n4418_), .Y(_abc_41356_new_n4419_));
INVX1 INVX1_52 ( .A(_abc_41356_new_n736_), .Y(_abc_41356_new_n737_));
INVX1 INVX1_520 ( .A(_abc_41356_new_n4449_), .Y(_abc_41356_new_n4450_));
INVX1 INVX1_521 ( .A(_abc_41356_new_n4460_), .Y(_abc_41356_new_n4461_));
INVX1 INVX1_522 ( .A(_abc_41356_new_n4492_), .Y(_abc_41356_new_n4493_));
INVX1 INVX1_523 ( .A(_abc_41356_new_n4503_), .Y(_abc_41356_new_n4504_));
INVX1 INVX1_524 ( .A(_abc_41356_new_n4533_), .Y(_abc_41356_new_n4534_));
INVX1 INVX1_525 ( .A(_abc_41356_new_n4544_), .Y(_abc_41356_new_n4545_));
INVX1 INVX1_526 ( .A(_abc_41356_new_n4574_), .Y(_abc_41356_new_n4575_));
INVX1 INVX1_527 ( .A(_abc_41356_new_n4592_), .Y(_abc_41356_new_n4593_));
INVX1 INVX1_528 ( .A(_abc_41356_new_n4617_), .Y(_abc_41356_new_n4618_));
INVX1 INVX1_529 ( .A(_abc_41356_new_n4627_), .Y(_abc_41356_new_n4628_));
INVX1 INVX1_53 ( .A(_abc_41356_new_n658_), .Y(_abc_41356_new_n738_));
INVX1 INVX1_530 ( .A(_abc_41356_new_n4657_), .Y(_abc_41356_new_n4658_));
INVX1 INVX1_531 ( .A(_abc_41356_new_n4667_), .Y(_abc_41356_new_n4668_));
INVX1 INVX1_532 ( .A(_abc_41356_new_n4692_), .Y(_abc_41356_new_n4693_));
INVX1 INVX1_533 ( .A(_abc_41356_new_n4704_), .Y(_abc_41356_new_n4705_));
INVX1 INVX1_534 ( .A(_abc_41356_new_n4731_), .Y(_abc_41356_new_n4732_));
INVX1 INVX1_535 ( .A(_abc_41356_new_n4741_), .Y(_abc_41356_new_n4742_));
INVX1 INVX1_536 ( .A(_abc_41356_new_n4769_), .Y(_abc_41356_new_n4770_));
INVX1 INVX1_537 ( .A(_abc_41356_new_n4781_), .Y(_abc_41356_new_n4782_));
INVX1 INVX1_538 ( .A(raddrhold_15_), .Y(_abc_41356_new_n4810_));
INVX1 INVX1_539 ( .A(_abc_41356_new_n3433_), .Y(_abc_41356_new_n4819_));
INVX1 INVX1_54 ( .A(_abc_41356_new_n743_), .Y(_abc_41356_new_n744_));
INVX1 INVX1_540 ( .A(_abc_41356_new_n3414_), .Y(_abc_41356_new_n4827_));
INVX1 INVX1_541 ( .A(waddrhold_0_), .Y(_abc_41356_new_n4848_));
INVX1 INVX1_542 ( .A(sp_1_), .Y(_abc_41356_new_n4857_));
INVX1 INVX1_543 ( .A(_abc_41356_new_n3358_), .Y(_abc_41356_new_n4858_));
INVX1 INVX1_544 ( .A(_abc_41356_new_n3363_), .Y(_abc_41356_new_n4859_));
INVX1 INVX1_545 ( .A(_abc_41356_new_n4883_), .Y(_abc_41356_new_n4884_));
INVX1 INVX1_546 ( .A(_abc_41356_new_n4920_), .Y(_abc_41356_new_n4921_));
INVX1 INVX1_547 ( .A(_abc_41356_new_n4894_), .Y(_abc_41356_new_n4930_));
INVX1 INVX1_548 ( .A(_abc_41356_new_n4956_), .Y(_abc_41356_new_n4957_));
INVX1 INVX1_549 ( .A(_abc_41356_new_n4967_), .Y(_abc_41356_new_n4969_));
INVX1 INVX1_55 ( .A(_abc_41356_new_n790_), .Y(_abc_41356_new_n791_));
INVX1 INVX1_550 ( .A(_abc_41356_new_n4995_), .Y(_abc_41356_new_n4996_));
INVX1 INVX1_551 ( .A(_abc_41356_new_n4968_), .Y(_abc_41356_new_n5005_));
INVX1 INVX1_552 ( .A(_abc_41356_new_n5032_), .Y(_abc_41356_new_n5033_));
INVX1 INVX1_553 ( .A(_abc_41356_new_n5007_), .Y(_abc_41356_new_n5043_));
INVX1 INVX1_554 ( .A(_abc_41356_new_n5069_), .Y(_abc_41356_new_n5070_));
INVX1 INVX1_555 ( .A(_abc_41356_new_n5042_), .Y(_abc_41356_new_n5079_));
INVX1 INVX1_556 ( .A(_abc_41356_new_n5106_), .Y(_abc_41356_new_n5107_));
INVX1 INVX1_557 ( .A(_abc_41356_new_n5081_), .Y(_abc_41356_new_n5117_));
INVX1 INVX1_558 ( .A(_abc_41356_new_n5143_), .Y(_abc_41356_new_n5144_));
INVX1 INVX1_559 ( .A(_abc_41356_new_n5116_), .Y(_abc_41356_new_n5153_));
INVX1 INVX1_56 ( .A(_abc_41356_new_n796_), .Y(_abc_41356_new_n797_));
INVX1 INVX1_560 ( .A(_abc_41356_new_n5180_), .Y(_abc_41356_new_n5181_));
INVX1 INVX1_561 ( .A(_abc_41356_new_n5155_), .Y(_abc_41356_new_n5191_));
INVX1 INVX1_562 ( .A(_abc_41356_new_n5217_), .Y(_abc_41356_new_n5218_));
INVX1 INVX1_563 ( .A(_abc_41356_new_n5190_), .Y(_abc_41356_new_n5227_));
INVX1 INVX1_564 ( .A(_abc_41356_new_n5254_), .Y(_abc_41356_new_n5255_));
INVX1 INVX1_565 ( .A(_abc_41356_new_n5229_), .Y(_abc_41356_new_n5267_));
INVX1 INVX1_566 ( .A(_abc_41356_new_n5292_), .Y(_abc_41356_new_n5293_));
INVX1 INVX1_567 ( .A(_abc_41356_new_n5266_), .Y(_abc_41356_new_n5304_));
INVX1 INVX1_568 ( .A(_abc_41356_new_n5332_), .Y(_abc_41356_new_n5333_));
INVX1 INVX1_569 ( .A(_abc_41356_new_n5306_), .Y(_abc_41356_new_n5342_));
INVX1 INVX1_57 ( .A(rdatahold_2_), .Y(_abc_41356_new_n829_));
INVX1 INVX1_570 ( .A(_abc_41356_new_n5369_), .Y(_abc_41356_new_n5370_));
INVX1 INVX1_571 ( .A(_abc_41356_new_n5341_), .Y(_abc_41356_new_n5379_));
INVX1 INVX1_572 ( .A(_abc_41356_new_n5404_), .Y(_abc_41356_new_n5405_));
INVX1 INVX1_573 ( .A(_abc_41356_new_n5295_), .Y(_abc_41356_new_n5412_));
INVX1 INVX1_574 ( .A(_abc_41356_new_n5413_), .Y(_abc_41356_new_n5414_));
INVX1 INVX1_575 ( .A(_abc_41356_new_n3396_), .Y(_abc_41356_new_n5466_));
INVX1 INVX1_576 ( .A(_abc_41356_new_n5495_), .Y(_abc_41356_new_n5496_));
INVX1 INVX1_577 ( .A(_abc_41356_new_n1292_), .Y(_abc_41356_new_n5504_));
INVX1 INVX1_578 ( .A(_abc_41356_new_n1364_), .Y(_abc_41356_new_n5508_));
INVX1 INVX1_579 ( .A(_abc_41356_new_n1424_), .Y(_abc_41356_new_n5538_));
INVX1 INVX1_58 ( .A(_abc_41356_new_n830_), .Y(_abc_41356_new_n831_));
INVX1 INVX1_580 ( .A(_abc_41356_new_n1368_), .Y(_abc_41356_new_n5542_));
INVX1 INVX1_581 ( .A(_abc_41356_new_n5549_), .Y(_abc_41356_new_n5550_));
INVX1 INVX1_582 ( .A(_abc_41356_new_n1261_), .Y(_abc_41356_new_n5563_));
INVX1 INVX1_583 ( .A(_abc_41356_new_n5566_), .Y(_abc_41356_new_n5567_));
INVX1 INVX1_584 ( .A(_abc_41356_new_n1273_), .Y(_abc_41356_new_n5568_));
INVX1 INVX1_585 ( .A(_abc_41356_new_n5571_), .Y(_abc_41356_new_n5572_));
INVX1 INVX1_586 ( .A(_abc_41356_new_n5573_), .Y(_abc_41356_new_n5574_));
INVX1 INVX1_587 ( .A(_abc_41356_new_n1426_), .Y(_abc_41356_new_n5578_));
INVX1 INVX1_588 ( .A(_abc_41356_new_n5580_), .Y(_abc_41356_new_n5581_));
INVX1 INVX1_589 ( .A(_abc_41356_new_n5584_), .Y(_abc_41356_new_n5585_));
INVX1 INVX1_59 ( .A(_abc_41356_new_n833_), .Y(_abc_41356_new_n834_));
INVX1 INVX1_590 ( .A(_abc_41356_new_n5591_), .Y(_abc_41356_new_n5592_));
INVX1 INVX1_591 ( .A(_abc_41356_new_n1297_), .Y(_abc_41356_new_n5612_));
INVX1 INVX1_592 ( .A(_abc_41356_new_n5613_), .Y(_abc_41356_new_n5614_));
INVX1 INVX1_593 ( .A(_abc_41356_new_n1431_), .Y(_abc_41356_new_n5621_));
INVX1 INVX1_594 ( .A(_abc_41356_new_n5622_), .Y(_abc_41356_new_n5623_));
INVX1 INVX1_595 ( .A(_abc_41356_new_n1360_), .Y(_abc_41356_new_n5629_));
INVX1 INVX1_596 ( .A(_abc_41356_new_n5630_), .Y(_abc_41356_new_n5632_));
INVX1 INVX1_597 ( .A(_abc_41356_new_n1274_), .Y(_abc_41356_new_n5639_));
INVX1 INVX1_598 ( .A(_abc_41356_new_n5642_), .Y(_abc_41356_new_n5643_));
INVX1 INVX1_599 ( .A(_abc_41356_new_n1262_), .Y(_abc_41356_new_n5655_));
INVX1 INVX1_6 ( .A(opcode_6_), .Y(_abc_41356_new_n514_));
INVX1 INVX1_60 ( .A(_abc_41356_new_n851_), .Y(_abc_41356_new_n852_));
INVX1 INVX1_600 ( .A(_abc_41356_new_n5661_), .Y(_abc_41356_new_n5662_));
INVX1 INVX1_601 ( .A(_abc_41356_new_n1442_), .Y(_abc_41356_new_n5665_));
INVX1 INVX1_602 ( .A(_abc_41356_new_n5666_), .Y(_abc_41356_new_n5667_));
INVX1 INVX1_603 ( .A(_abc_41356_new_n5673_), .Y(_abc_41356_new_n5674_));
INVX1 INVX1_604 ( .A(_abc_41356_new_n5676_), .Y(_abc_41356_new_n5677_));
INVX1 INVX1_605 ( .A(_abc_41356_new_n1275_), .Y(_abc_41356_new_n5683_));
INVX1 INVX1_606 ( .A(_abc_41356_new_n5686_), .Y(_abc_41356_new_n5687_));
INVX1 INVX1_607 ( .A(_abc_41356_new_n1263_), .Y(_abc_41356_new_n5699_));
INVX1 INVX1_608 ( .A(_abc_41356_new_n1324_), .Y(_abc_41356_new_n5704_));
INVX1 INVX1_609 ( .A(_abc_41356_new_n1334_), .Y(_abc_41356_new_n5706_));
INVX1 INVX1_61 ( .A(_abc_41356_new_n857_), .Y(_abc_41356_new_n858_));
INVX1 INVX1_610 ( .A(_abc_41356_new_n5705_), .Y(_abc_41356_new_n5708_));
INVX1 INVX1_611 ( .A(_abc_41356_new_n5713_), .Y(_abc_41356_new_n5714_));
INVX1 INVX1_612 ( .A(_abc_41356_new_n1389_), .Y(_abc_41356_new_n5716_));
INVX1 INVX1_613 ( .A(_abc_41356_new_n5720_), .Y(_abc_41356_new_n5721_));
INVX1 INVX1_614 ( .A(_abc_41356_new_n1459_), .Y(_abc_41356_new_n5723_));
INVX1 INVX1_615 ( .A(_abc_41356_new_n1796_), .Y(_abc_41356_new_n5732_));
INVX1 INVX1_616 ( .A(_abc_41356_new_n1264_), .Y(_abc_41356_new_n5748_));
INVX1 INVX1_617 ( .A(_abc_41356_new_n5755_), .Y(_abc_41356_new_n5756_));
INVX1 INVX1_618 ( .A(_abc_41356_new_n5763_), .Y(_abc_41356_new_n5764_));
INVX1 INVX1_619 ( .A(_abc_41356_new_n5769_), .Y(_abc_41356_new_n5770_));
INVX1 INVX1_62 ( .A(rdatahold_3_), .Y(_abc_41356_new_n890_));
INVX1 INVX1_620 ( .A(_abc_41356_new_n5775_), .Y(_abc_41356_new_n5776_));
INVX1 INVX1_621 ( .A(_abc_41356_new_n1797_), .Y(_abc_41356_new_n5781_));
INVX1 INVX1_622 ( .A(_abc_41356_new_n1265_), .Y(_abc_41356_new_n5798_));
INVX1 INVX1_623 ( .A(_abc_41356_new_n1317_), .Y(_abc_41356_new_n5805_));
INVX1 INVX1_624 ( .A(_abc_41356_new_n5803_), .Y(_abc_41356_new_n5806_));
INVX1 INVX1_625 ( .A(_abc_41356_new_n5812_), .Y(_abc_41356_new_n5813_));
INVX1 INVX1_626 ( .A(_abc_41356_new_n1446_), .Y(_abc_41356_new_n5815_));
INVX1 INVX1_627 ( .A(_abc_41356_new_n1380_), .Y(_abc_41356_new_n5822_));
INVX1 INVX1_628 ( .A(_abc_41356_new_n5820_), .Y(_abc_41356_new_n5823_));
INVX1 INVX1_629 ( .A(_abc_41356_new_n1279_), .Y(_abc_41356_new_n5830_));
INVX1 INVX1_63 ( .A(_abc_41356_new_n891_), .Y(_abc_41356_new_n892_));
INVX1 INVX1_630 ( .A(_abc_41356_new_n5840_), .Y(_abc_41356_new_n5841_));
INVX1 INVX1_631 ( .A(_abc_41356_new_n5843_), .Y(_abc_41356_new_n5844_));
INVX1 INVX1_632 ( .A(_abc_41356_new_n1286_), .Y(_abc_41356_new_n5849_));
INVX1 INVX1_633 ( .A(_abc_41356_new_n2023_), .Y(_abc_41356_new_n5853_));
INVX1 INVX1_634 ( .A(_abc_41356_new_n5854_), .Y(_abc_41356_new_n5855_));
INVX1 INVX1_635 ( .A(_abc_41356_new_n5856_), .Y(_abc_41356_new_n5857_));
INVX1 INVX1_636 ( .A(_abc_41356_new_n5863_), .Y(_abc_41356_new_n5864_));
INVX1 INVX1_637 ( .A(_abc_41356_new_n3349_), .Y(_abc_41356_new_n5882_));
INVX1 INVX1_638 ( .A(sp_0_), .Y(_abc_41356_new_n5883_));
INVX1 INVX1_639 ( .A(_abc_41356_new_n5884_), .Y(_abc_41356_new_n5885_));
INVX1 INVX1_64 ( .A(regfil_7__4_), .Y(_abc_41356_new_n893_));
INVX1 INVX1_640 ( .A(_abc_41356_new_n5886_), .Y(_abc_41356_new_n5887_));
INVX1 INVX1_641 ( .A(_abc_41356_new_n5891_), .Y(_abc_41356_new_n5892_));
INVX1 INVX1_642 ( .A(_abc_41356_new_n5896_), .Y(_abc_41356_new_n5897_));
INVX1 INVX1_643 ( .A(_abc_41356_new_n4896_), .Y(_abc_41356_new_n5912_));
INVX1 INVX1_644 ( .A(_abc_41356_new_n5920_), .Y(_abc_41356_new_n5921_));
INVX1 INVX1_645 ( .A(_abc_41356_new_n5946_), .Y(_abc_41356_new_n5947_));
INVX1 INVX1_646 ( .A(_abc_41356_new_n5962_), .Y(_abc_41356_new_n5963_));
INVX1 INVX1_647 ( .A(_abc_41356_new_n5984_), .Y(_abc_41356_new_n5985_));
INVX1 INVX1_648 ( .A(_abc_41356_new_n5995_), .Y(_abc_41356_new_n5997_));
INVX1 INVX1_649 ( .A(_abc_41356_new_n6002_), .Y(_abc_41356_new_n6003_));
INVX1 INVX1_65 ( .A(_abc_41356_new_n894_), .Y(_abc_41356_new_n895_));
INVX1 INVX1_650 ( .A(_abc_41356_new_n6027_), .Y(_abc_41356_new_n6028_));
INVX1 INVX1_651 ( .A(_abc_41356_new_n6036_), .Y(_abc_41356_new_n6037_));
INVX1 INVX1_652 ( .A(_abc_41356_new_n5996_), .Y(_abc_41356_new_n6041_));
INVX1 INVX1_653 ( .A(_abc_41356_new_n6066_), .Y(_abc_41356_new_n6067_));
INVX1 INVX1_654 ( .A(_abc_41356_new_n6075_), .Y(_abc_41356_new_n6076_));
INVX1 INVX1_655 ( .A(_abc_41356_new_n6098_), .Y(_abc_41356_new_n6099_));
INVX1 INVX1_656 ( .A(_abc_41356_new_n6109_), .Y(_abc_41356_new_n6110_));
INVX1 INVX1_657 ( .A(_abc_41356_new_n6061_), .Y(_abc_41356_new_n6113_));
INVX1 INVX1_658 ( .A(_abc_41356_new_n6136_), .Y(_abc_41356_new_n6137_));
INVX1 INVX1_659 ( .A(_abc_41356_new_n6148_), .Y(_abc_41356_new_n6149_));
INVX1 INVX1_66 ( .A(_abc_41356_new_n896_), .Y(_abc_41356_new_n897_));
INVX1 INVX1_660 ( .A(_abc_41356_new_n6117_), .Y(_abc_41356_new_n6152_));
INVX1 INVX1_661 ( .A(_abc_41356_new_n6175_), .Y(_abc_41356_new_n6176_));
INVX1 INVX1_662 ( .A(_abc_41356_new_n6156_), .Y(_abc_41356_new_n6180_));
INVX1 INVX1_663 ( .A(_abc_41356_new_n6182_), .Y(_abc_41356_new_n6183_));
INVX1 INVX1_664 ( .A(_abc_41356_new_n6193_), .Y(_abc_41356_new_n6194_));
INVX1 INVX1_665 ( .A(_abc_41356_new_n6219_), .Y(_abc_41356_new_n6220_));
INVX1 INVX1_666 ( .A(_abc_41356_new_n6218_), .Y(_abc_41356_new_n6227_));
INVX1 INVX1_667 ( .A(_abc_41356_new_n6213_), .Y(_abc_41356_new_n6249_));
INVX1 INVX1_668 ( .A(_abc_41356_new_n6258_), .Y(_abc_41356_new_n6259_));
INVX1 INVX1_669 ( .A(_abc_41356_new_n6263_), .Y(_abc_41356_new_n6264_));
INVX1 INVX1_67 ( .A(_abc_41356_new_n902_), .Y(_abc_41356_new_n903_));
INVX1 INVX1_670 ( .A(_abc_41356_new_n6288_), .Y(_abc_41356_new_n6289_));
INVX1 INVX1_671 ( .A(_abc_41356_new_n6248_), .Y(_abc_41356_new_n6299_));
INVX1 INVX1_672 ( .A(_abc_41356_new_n6304_), .Y(_abc_41356_new_n6305_));
INVX1 INVX1_673 ( .A(_abc_41356_new_n6324_), .Y(_abc_41356_new_n6325_));
INVX1 INVX1_674 ( .A(_abc_41356_new_n6298_), .Y(_abc_41356_new_n6329_));
INVX1 INVX1_675 ( .A(_abc_41356_new_n6323_), .Y(_abc_41356_new_n6338_));
INVX1 INVX1_676 ( .A(_abc_41356_new_n6363_), .Y(_abc_41356_new_n6364_));
INVX1 INVX1_677 ( .A(_abc_41356_new_n6331_), .Y(_abc_41356_new_n6369_));
INVX1 INVX1_678 ( .A(_abc_41356_new_n6362_), .Y(_abc_41356_new_n6377_));
INVX1 INVX1_679 ( .A(_abc_41356_new_n6436_), .Y(_abc_41356_new_n6438_));
INVX1 INVX1_68 ( .A(_abc_41356_new_n918_), .Y(_abc_41356_new_n919_));
INVX1 INVX1_680 ( .A(_abc_41356_new_n6462_), .Y(_abc_41356_new_n6463_));
INVX1 INVX1_681 ( .A(_abc_41356_new_n6476_), .Y(_abc_41356_new_n6477_));
INVX1 INVX1_682 ( .A(_abc_41356_new_n6481_), .Y(_abc_41356_new_n6482_));
INVX1 INVX1_683 ( .A(_abc_41356_new_n6486_), .Y(_abc_41356_new_n6487_));
INVX1 INVX1_684 ( .A(_abc_41356_new_n3368_), .Y(_abc_41356_new_n6488_));
INVX1 INVX1_685 ( .A(_abc_41356_new_n6489_), .Y(_abc_41356_new_n6490_));
INVX1 INVX1_686 ( .A(_abc_41356_new_n1417_), .Y(_abc_41356_new_n6494_));
INVX1 INVX1_687 ( .A(_abc_41356_new_n6504_), .Y(_abc_41356_new_n6505_));
INVX1 INVX1_688 ( .A(_abc_41356_new_n681_), .Y(_abc_41356_new_n6513_));
INVX1 INVX1_689 ( .A(_abc_41356_new_n6517_), .Y(_abc_41356_new_n6518_));
INVX1 INVX1_69 ( .A(_abc_41356_new_n924_), .Y(_abc_41356_new_n925_));
INVX1 INVX1_690 ( .A(_abc_41356_new_n2057_), .Y(_abc_41356_new_n6519_));
INVX1 INVX1_691 ( .A(_abc_41356_new_n6529_), .Y(_abc_41356_new_n6530_));
INVX1 INVX1_692 ( .A(_abc_41356_new_n548_), .Y(_abc_41356_new_n6532_));
INVX1 INVX1_693 ( .A(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6533_));
INVX1 INVX1_694 ( .A(_abc_41356_new_n6537_), .Y(_abc_41356_new_n6538_));
INVX1 INVX1_695 ( .A(_abc_41356_new_n6577_), .Y(_abc_41356_new_n6578_));
INVX1 INVX1_696 ( .A(_abc_41356_new_n6590_), .Y(_abc_41356_new_n6591_));
INVX1 INVX1_697 ( .A(_abc_41356_new_n3879_), .Y(_abc_41356_new_n6598_));
INVX1 INVX1_698 ( .A(_abc_41356_new_n3883_), .Y(_abc_41356_new_n6600_));
INVX1 INVX1_699 ( .A(pc_3_), .Y(_abc_41356_new_n6602_));
INVX1 INVX1_7 ( .A(opcode_7_), .Y(_abc_41356_new_n515_));
INVX1 INVX1_70 ( .A(_abc_41356_new_n957_), .Y(_abc_41356_new_n958_));
INVX1 INVX1_700 ( .A(_abc_41356_new_n2070_), .Y(_abc_41356_new_n6603_));
INVX1 INVX1_701 ( .A(_abc_41356_new_n6613_), .Y(_abc_41356_new_n6614_));
INVX1 INVX1_702 ( .A(_abc_41356_new_n6616_), .Y(_abc_41356_new_n6617_));
INVX1 INVX1_703 ( .A(_abc_41356_new_n528_), .Y(_abc_41356_new_n6619_));
INVX1 INVX1_704 ( .A(_abc_41356_new_n6620_), .Y(_abc_41356_new_n6621_));
INVX1 INVX1_705 ( .A(_abc_41356_new_n6628_), .Y(_abc_41356_new_n6629_));
INVX1 INVX1_706 ( .A(_abc_41356_new_n6631_), .Y(_abc_41356_new_n6632_));
INVX1 INVX1_707 ( .A(_abc_41356_new_n6641_), .Y(_abc_41356_new_n6642_));
INVX1 INVX1_708 ( .A(_abc_41356_new_n6685_), .Y(_abc_41356_new_n6686_));
INVX1 INVX1_709 ( .A(_abc_41356_new_n6688_), .Y(_abc_41356_new_n6689_));
INVX1 INVX1_71 ( .A(_abc_41356_new_n698_), .Y(_abc_41356_new_n959_));
INVX1 INVX1_710 ( .A(_abc_41356_new_n6691_), .Y(_abc_41356_new_n6692_));
INVX1 INVX1_711 ( .A(_abc_41356_new_n6700_), .Y(_abc_41356_new_n6701_));
INVX1 INVX1_712 ( .A(_abc_41356_new_n6703_), .Y(_abc_41356_new_n6704_));
INVX1 INVX1_713 ( .A(_abc_41356_new_n4023_), .Y(_abc_41356_new_n6711_));
INVX1 INVX1_714 ( .A(_abc_41356_new_n4028_), .Y(_abc_41356_new_n6713_));
INVX1 INVX1_715 ( .A(pc_6_), .Y(_abc_41356_new_n6716_));
INVX1 INVX1_716 ( .A(_abc_41356_new_n6675_), .Y(_abc_41356_new_n6717_));
INVX1 INVX1_717 ( .A(_abc_41356_new_n6727_), .Y(_abc_41356_new_n6728_));
INVX1 INVX1_718 ( .A(_abc_41356_new_n6740_), .Y(_abc_41356_new_n6741_));
INVX1 INVX1_719 ( .A(_abc_41356_new_n6749_), .Y(_abc_41356_new_n6750_));
INVX1 INVX1_72 ( .A(_abc_41356_new_n963_), .Y(_abc_41356_new_n964_));
INVX1 INVX1_720 ( .A(_abc_41356_new_n6751_), .Y(_abc_41356_new_n6752_));
INVX1 INVX1_721 ( .A(_abc_41356_new_n6755_), .Y(_abc_41356_new_n6756_));
INVX1 INVX1_722 ( .A(_abc_41356_new_n6763_), .Y(_abc_41356_new_n6764_));
INVX1 INVX1_723 ( .A(_abc_41356_new_n6765_), .Y(_abc_41356_new_n6766_));
INVX1 INVX1_724 ( .A(_abc_41356_new_n6768_), .Y(_abc_41356_new_n6769_));
INVX1 INVX1_725 ( .A(_abc_41356_new_n6770_), .Y(_abc_41356_new_n6771_));
INVX1 INVX1_726 ( .A(_abc_41356_new_n6777_), .Y(_abc_41356_new_n6778_));
INVX1 INVX1_727 ( .A(_abc_41356_new_n6780_), .Y(_abc_41356_new_n6781_));
INVX1 INVX1_728 ( .A(_abc_41356_new_n6800_), .Y(_abc_41356_new_n6801_));
INVX1 INVX1_729 ( .A(_abc_41356_new_n6806_), .Y(_abc_41356_new_n6807_));
INVX1 INVX1_73 ( .A(_abc_41356_new_n899_), .Y(_abc_41356_new_n965_));
INVX1 INVX1_730 ( .A(_abc_41356_new_n6814_), .Y(_abc_41356_new_n6815_));
INVX1 INVX1_731 ( .A(pc_9_), .Y(_abc_41356_new_n6823_));
INVX1 INVX1_732 ( .A(_abc_41356_new_n6791_), .Y(_abc_41356_new_n6824_));
INVX1 INVX1_733 ( .A(_abc_41356_new_n2111_), .Y(_abc_41356_new_n6829_));
INVX1 INVX1_734 ( .A(_abc_41356_new_n2119_), .Y(_abc_41356_new_n6831_));
INVX1 INVX1_735 ( .A(_abc_41356_new_n6838_), .Y(_abc_41356_new_n6839_));
INVX1 INVX1_736 ( .A(_abc_41356_new_n6844_), .Y(_abc_41356_new_n6845_));
INVX1 INVX1_737 ( .A(_abc_41356_new_n6852_), .Y(_abc_41356_new_n6853_));
INVX1 INVX1_738 ( .A(_abc_41356_new_n6822_), .Y(_abc_41356_new_n6861_));
INVX1 INVX1_739 ( .A(_abc_41356_new_n6873_), .Y(_abc_41356_new_n6874_));
INVX1 INVX1_74 ( .A(_abc_41356_new_n970_), .Y(_abc_41356_new_n971_));
INVX1 INVX1_740 ( .A(_abc_41356_new_n6886_), .Y(_abc_41356_new_n6887_));
INVX1 INVX1_741 ( .A(_abc_41356_new_n6894_), .Y(_abc_41356_new_n6895_));
INVX1 INVX1_742 ( .A(_abc_41356_new_n6897_), .Y(_abc_41356_new_n6898_));
INVX1 INVX1_743 ( .A(_abc_41356_new_n2191_), .Y(_abc_41356_new_n6900_));
INVX1 INVX1_744 ( .A(_abc_41356_new_n2199_), .Y(_abc_41356_new_n6902_));
INVX1 INVX1_745 ( .A(pc_11_), .Y(_abc_41356_new_n6906_));
INVX1 INVX1_746 ( .A(_abc_41356_new_n6908_), .Y(_abc_41356_new_n6909_));
INVX1 INVX1_747 ( .A(_abc_41356_new_n6938_), .Y(_abc_41356_new_n6939_));
INVX1 INVX1_748 ( .A(_abc_41356_new_n6932_), .Y(_abc_41356_new_n6945_));
INVX1 INVX1_749 ( .A(_abc_41356_new_n6963_), .Y(_abc_41356_new_n6964_));
INVX1 INVX1_75 ( .A(_abc_41356_new_n972_), .Y(_abc_41356_new_n973_));
INVX1 INVX1_750 ( .A(_abc_41356_new_n6996_), .Y(_abc_41356_new_n6997_));
INVX1 INVX1_751 ( .A(_abc_41356_new_n7028_), .Y(_abc_41356_new_n7029_));
INVX1 INVX1_752 ( .A(_abc_41356_new_n7058_), .Y(_abc_41356_new_n7059_));
INVX1 INVX1_753 ( .A(_abc_41356_new_n3318_), .Y(_abc_41356_new_n7064_));
INVX1 INVX1_754 ( .A(_abc_41356_new_n7066_), .Y(_abc_41356_new_n7067_));
INVX1 INVX1_755 ( .A(_abc_41356_new_n7065_), .Y(_abc_41356_new_n7068_));
INVX1 INVX1_756 ( .A(_abc_41356_new_n3204_), .Y(_abc_41356_new_n7072_));
INVX1 INVX1_757 ( .A(_abc_41356_new_n7080_), .Y(_abc_41356_new_n7081_));
INVX1 INVX1_758 ( .A(_abc_41356_new_n7229_), .Y(_abc_41356_new_n7230_));
INVX1 INVX1_759 ( .A(_abc_41356_new_n7244_), .Y(_abc_41356_new_n7245_));
INVX1 INVX1_76 ( .A(alu_res_4_), .Y(_abc_41356_new_n974_));
INVX1 INVX1_760 ( .A(statesel_2_), .Y(_abc_41356_new_n7250_));
INVX1 INVX1_761 ( .A(statesel_4_), .Y(_abc_41356_new_n7260_));
INVX1 INVX1_762 ( .A(_abc_41356_new_n3554_), .Y(_abc_41356_new_n7262_));
INVX1 INVX1_763 ( .A(_abc_41356_new_n7254_), .Y(_abc_41356_new_n7263_));
INVX1 INVX1_764 ( .A(_abc_41356_new_n7274_), .Y(_abc_41356_new_n7275_));
INVX1 INVX1_765 ( .A(_abc_41356_new_n7283_), .Y(_abc_41356_new_n7284_));
INVX1 INVX1_766 ( .A(_abc_41356_new_n7286_), .Y(_abc_41356_new_n7287_));
INVX1 INVX1_767 ( .A(_abc_41356_new_n1233_), .Y(_abc_41356_new_n7288_));
INVX1 INVX1_768 ( .A(_abc_41356_new_n7290_), .Y(_abc_41356_new_n7291_));
INVX1 INVX1_769 ( .A(_abc_41356_new_n7293_), .Y(_abc_41356_new_n7294_));
INVX1 INVX1_77 ( .A(_abc_41356_new_n714_), .Y(_abc_41356_new_n975_));
INVX1 INVX1_770 ( .A(_abc_41356_new_n7295_), .Y(_abc_41356_new_n7297_));
INVX1 INVX1_771 ( .A(sign), .Y(_abc_41356_new_n7298_));
INVX1 INVX1_772 ( .A(_abc_41356_new_n7303_), .Y(_abc_41356_new_n7304_));
INVX1 INVX1_773 ( .A(_abc_41356_new_n7309_), .Y(_abc_41356_new_n7310_));
INVX1 INVX1_774 ( .A(parity), .Y(_abc_41356_new_n7320_));
INVX1 INVX1_775 ( .A(_abc_41356_new_n7322_), .Y(_abc_41356_new_n7323_));
INVX1 INVX1_776 ( .A(_abc_41356_new_n7327_), .Y(_abc_41356_new_n7328_));
INVX1 INVX1_777 ( .A(_abc_41356_new_n3391_), .Y(_abc_41356_new_n7333_));
INVX1 INVX1_778 ( .A(_abc_41356_new_n7337_), .Y(_abc_41356_new_n7338_));
INVX1 INVX1_779 ( .A(_abc_41356_new_n7261_), .Y(_abc_41356_new_n7342_));
INVX1 INVX1_78 ( .A(_abc_41356_new_n977_), .Y(_abc_41356_new_n978_));
INVX1 INVX1_780 ( .A(_abc_41356_new_n7343_), .Y(_abc_41356_new_n7344_));
INVX1 INVX1_781 ( .A(_abc_41356_new_n7276_), .Y(_abc_41356_new_n7346_));
INVX1 INVX1_782 ( .A(_abc_41356_new_n3489_), .Y(_abc_41356_new_n7347_));
INVX1 INVX1_783 ( .A(_abc_41356_new_n550_), .Y(_abc_41356_new_n7353_));
INVX1 INVX1_784 ( .A(_abc_41356_new_n7175_), .Y(_abc_41356_new_n7354_));
INVX1 INVX1_785 ( .A(_abc_41356_new_n7359_), .Y(_abc_41356_new_n7360_));
INVX1 INVX1_786 ( .A(_abc_41356_new_n7361_), .Y(_abc_41356_new_n7362_));
INVX1 INVX1_787 ( .A(_abc_41356_new_n6526_), .Y(_abc_41356_new_n7365_));
INVX1 INVX1_788 ( .A(_abc_41356_new_n7370_), .Y(_abc_41356_new_n7371_));
INVX1 INVX1_789 ( .A(_abc_41356_new_n7373_), .Y(_abc_41356_new_n7374_));
INVX1 INVX1_79 ( .A(_abc_41356_new_n982_), .Y(_abc_41356_new_n983_));
INVX1 INVX1_790 ( .A(_abc_41356_new_n7379_), .Y(_abc_41356_new_n7380_));
INVX1 INVX1_791 ( .A(_abc_41356_new_n7382_), .Y(_abc_41356_new_n7383_));
INVX1 INVX1_792 ( .A(_abc_41356_new_n7271_), .Y(_abc_41356_new_n7387_));
INVX1 INVX1_793 ( .A(_abc_41356_new_n7252_), .Y(_abc_41356_new_n7388_));
INVX1 INVX1_794 ( .A(_abc_41356_new_n7264_), .Y(_abc_41356_new_n7389_));
INVX1 INVX1_795 ( .A(_abc_41356_new_n7253_), .Y(_abc_41356_new_n7392_));
INVX1 INVX1_796 ( .A(_abc_41356_new_n680_), .Y(_abc_41356_new_n7399_));
INVX1 INVX1_797 ( .A(_abc_41356_new_n7285_), .Y(_abc_41356_new_n7401_));
INVX1 INVX1_798 ( .A(_abc_41356_new_n7412_), .Y(_abc_41356_new_n7413_));
INVX1 INVX1_799 ( .A(_abc_41356_new_n7418_), .Y(_abc_41356_new_n7419_));
INVX1 INVX1_8 ( .A(state_4_), .Y(_abc_41356_new_n517_));
INVX1 INVX1_80 ( .A(_abc_41356_new_n985_), .Y(_abc_41356_new_n986_));
INVX1 INVX1_800 ( .A(_abc_41356_new_n7408_), .Y(_abc_41356_new_n7420_));
INVX1 INVX1_801 ( .A(_abc_41356_new_n7428_), .Y(_abc_41356_new_n7429_));
INVX1 INVX1_802 ( .A(_abc_41356_new_n7431_), .Y(_abc_41356_new_n7432_));
INVX1 INVX1_803 ( .A(_abc_41356_new_n7433_), .Y(_abc_41356_new_n7434_));
INVX1 INVX1_804 ( .A(_abc_41356_new_n7316_), .Y(_abc_41356_new_n7441_));
INVX1 INVX1_805 ( .A(_abc_41356_new_n3001_), .Y(_abc_41356_new_n7442_));
INVX1 INVX1_806 ( .A(_abc_41356_new_n3608_), .Y(_abc_41356_new_n7446_));
INVX1 INVX1_807 ( .A(_abc_41356_new_n7447_), .Y(_abc_41356_new_n7448_));
INVX1 INVX1_808 ( .A(_abc_41356_new_n7449_), .Y(_abc_41356_new_n7450_));
INVX1 INVX1_809 ( .A(_abc_41356_new_n7456_), .Y(_abc_41356_new_n7457_));
INVX1 INVX1_81 ( .A(_abc_41356_new_n991_), .Y(_abc_41356_new_n992_));
INVX1 INVX1_810 ( .A(_abc_41356_new_n7459_), .Y(_abc_41356_new_n7460_));
INVX1 INVX1_811 ( .A(_abc_41356_new_n3445_), .Y(_abc_41356_new_n7462_));
INVX1 INVX1_812 ( .A(_abc_41356_new_n7465_), .Y(_abc_41356_new_n7466_));
INVX1 INVX1_813 ( .A(_abc_41356_new_n7228_), .Y(_abc_41356_new_n7467_));
INVX1 INVX1_814 ( .A(_abc_41356_new_n7475_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_1_));
INVX1 INVX1_815 ( .A(_abc_41356_new_n7477_), .Y(_abc_41356_new_n7478_));
INVX1 INVX1_816 ( .A(_abc_41356_new_n7483_), .Y(_abc_41356_new_n7484_));
INVX1 INVX1_817 ( .A(_abc_41356_new_n3555_), .Y(_abc_41356_new_n7485_));
INVX1 INVX1_818 ( .A(_abc_41356_new_n7487_), .Y(_abc_41356_new_n7488_));
INVX1 INVX1_819 ( .A(_abc_41356_new_n7492_), .Y(_abc_41356_new_n7493_));
INVX1 INVX1_82 ( .A(rdatahold_5_), .Y(_abc_41356_new_n1024_));
INVX1 INVX1_820 ( .A(_abc_41356_new_n7496_), .Y(_abc_41356_new_n7497_));
INVX1 INVX1_821 ( .A(_abc_41356_new_n507_), .Y(_abc_41356_new_n7498_));
INVX1 INVX1_822 ( .A(_abc_41356_new_n7508_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_2_));
INVX1 INVX1_823 ( .A(_abc_41356_new_n3556_), .Y(_abc_41356_new_n7512_));
INVX1 INVX1_824 ( .A(_abc_41356_new_n7407_), .Y(_abc_41356_new_n7513_));
INVX1 INVX1_825 ( .A(_abc_41356_new_n7515_), .Y(_abc_41356_new_n7516_));
INVX1 INVX1_826 ( .A(_abc_41356_new_n7409_), .Y(_abc_41356_new_n7518_));
INVX1 INVX1_827 ( .A(_abc_41356_new_n7525_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_3_));
INVX1 INVX1_828 ( .A(_abc_41356_new_n7453_), .Y(_abc_41356_new_n7528_));
INVX1 INVX1_829 ( .A(_abc_41356_new_n7502_), .Y(_abc_41356_new_n7531_));
INVX1 INVX1_83 ( .A(_abc_41356_new_n1025_), .Y(_abc_41356_new_n1026_));
INVX1 INVX1_830 ( .A(_abc_41356_new_n7332_), .Y(_abc_41356_new_n7542_));
INVX1 INVX1_831 ( .A(_abc_41356_new_n6089_), .Y(_abc_41356_new_n7555_));
INVX1 INVX1_832 ( .A(intr), .Y(_abc_41356_new_n7558_));
INVX1 INVX1_833 ( .A(alu__abc_40887_new_n34_), .Y(alu__abc_40887_new_n35_));
INVX1 INVX1_834 ( .A(alu__abc_40887_new_n36_), .Y(alu__abc_40887_new_n37_));
INVX1 INVX1_835 ( .A(alu__abc_40887_new_n38_), .Y(alu__abc_40887_new_n39_));
INVX1 INVX1_836 ( .A(alu_oprb_6_), .Y(alu__abc_40887_new_n40_));
INVX1 INVX1_837 ( .A(alu_opra_6_), .Y(alu__abc_40887_new_n41_));
INVX1 INVX1_838 ( .A(alu__abc_40887_new_n42_), .Y(alu__abc_40887_new_n43_));
INVX1 INVX1_839 ( .A(alu__abc_40887_new_n44_), .Y(alu__abc_40887_new_n45_));
INVX1 INVX1_84 ( .A(_abc_41356_new_n530_), .Y(_abc_41356_new_n1029_));
INVX1 INVX1_840 ( .A(alu__abc_40887_new_n46_), .Y(alu__abc_40887_new_n47_));
INVX1 INVX1_841 ( .A(alu__abc_40887_new_n53_), .Y(alu__abc_40887_new_n54_));
INVX1 INVX1_842 ( .A(alu_oprb_2_), .Y(alu__abc_40887_new_n55_));
INVX1 INVX1_843 ( .A(alu_opra_2_), .Y(alu__abc_40887_new_n56_));
INVX1 INVX1_844 ( .A(alu__abc_40887_new_n57_), .Y(alu__abc_40887_new_n58_));
INVX1 INVX1_845 ( .A(alu__abc_40887_new_n60_), .Y(alu__abc_40887_new_n61_));
INVX1 INVX1_846 ( .A(alu__abc_40887_new_n69_), .Y(alu__abc_40887_new_n70_));
INVX1 INVX1_847 ( .A(alu_oprb_4_), .Y(alu__abc_40887_new_n71_));
INVX1 INVX1_848 ( .A(alu_opra_4_), .Y(alu__abc_40887_new_n72_));
INVX1 INVX1_849 ( .A(alu__abc_40887_new_n73_), .Y(alu__abc_40887_new_n74_));
INVX1 INVX1_85 ( .A(_abc_41356_new_n1030_), .Y(_abc_41356_new_n1031_));
INVX1 INVX1_850 ( .A(alu_oprb_5_), .Y(alu__abc_40887_new_n76_));
INVX1 INVX1_851 ( .A(alu_opra_5_), .Y(alu__abc_40887_new_n77_));
INVX1 INVX1_852 ( .A(alu__abc_40887_new_n78_), .Y(alu__abc_40887_new_n79_));
INVX1 INVX1_853 ( .A(alu__abc_40887_new_n80_), .Y(alu__abc_40887_new_n81_));
INVX1 INVX1_854 ( .A(alu__abc_40887_new_n84_), .Y(alu__abc_40887_new_n85_));
INVX1 INVX1_855 ( .A(alu__abc_40887_new_n86_), .Y(alu__abc_40887_new_n87_));
INVX1 INVX1_856 ( .A(alu__abc_40887_new_n91_), .Y(alu__abc_40887_new_n92_));
INVX1 INVX1_857 ( .A(alu__abc_40887_new_n95_), .Y(alu__abc_40887_new_n96_));
INVX1 INVX1_858 ( .A(alu__abc_40887_new_n90_), .Y(alu__abc_40887_new_n97_));
INVX1 INVX1_859 ( .A(alu__abc_40887_new_n99_), .Y(alu__abc_40887_new_n100_));
INVX1 INVX1_86 ( .A(_abc_41356_new_n1033_), .Y(_abc_41356_new_n1034_));
INVX1 INVX1_860 ( .A(alu__abc_40887_new_n101_), .Y(alu__abc_40887_new_n102_));
INVX1 INVX1_861 ( .A(alu__abc_40887_new_n82_), .Y(alu__abc_40887_new_n103_));
INVX1 INVX1_862 ( .A(alu__abc_40887_new_n105_), .Y(alu__abc_40887_new_n106_));
INVX1 INVX1_863 ( .A(alu__abc_40887_new_n111_), .Y(alu__abc_40887_new_n112_));
INVX1 INVX1_864 ( .A(alu__abc_40887_new_n50_), .Y(alu__abc_40887_new_n115_));
INVX1 INVX1_865 ( .A(alu_oprb_0_), .Y(alu__abc_40887_new_n116_));
INVX1 INVX1_866 ( .A(alu_opra_0_), .Y(alu__abc_40887_new_n117_));
INVX1 INVX1_867 ( .A(alu__abc_40887_new_n118_), .Y(alu__abc_40887_new_n119_));
INVX1 INVX1_868 ( .A(alu__abc_40887_new_n109_), .Y(alu__abc_40887_new_n123_));
INVX1 INVX1_869 ( .A(alu__abc_40887_new_n132_), .Y(alu__abc_40887_new_n133_));
INVX1 INVX1_87 ( .A(_abc_41356_new_n1035_), .Y(_abc_41356_new_n1036_));
INVX1 INVX1_870 ( .A(alu_sel_2_), .Y(alu__abc_40887_new_n135_));
INVX1 INVX1_871 ( .A(alu_sel_1_), .Y(alu__abc_40887_new_n136_));
INVX1 INVX1_872 ( .A(alu__abc_40887_new_n138_), .Y(alu__abc_40887_new_n139_));
INVX1 INVX1_873 ( .A(alu__abc_40887_new_n142_), .Y(alu__abc_40887_new_n143_));
INVX1 INVX1_874 ( .A(alu_oprb_3_), .Y(alu__abc_40887_new_n146_));
INVX1 INVX1_875 ( .A(alu__abc_40887_new_n63_), .Y(alu__abc_40887_new_n148_));
INVX1 INVX1_876 ( .A(alu__abc_40887_new_n151_), .Y(alu__abc_40887_new_n152_));
INVX1 INVX1_877 ( .A(alu_oprb_1_), .Y(alu__abc_40887_new_n153_));
INVX1 INVX1_878 ( .A(alu__abc_40887_new_n154_), .Y(alu__abc_40887_new_n155_));
INVX1 INVX1_879 ( .A(alu__abc_40887_new_n167_), .Y(alu__abc_40887_new_n168_));
INVX1 INVX1_88 ( .A(regfil_0__6_), .Y(_abc_41356_new_n1076_));
INVX1 INVX1_880 ( .A(alu__abc_40887_new_n171_), .Y(alu__abc_40887_new_n172_));
INVX1 INVX1_881 ( .A(alu__abc_40887_new_n175_), .Y(alu__abc_40887_new_n176_));
INVX1 INVX1_882 ( .A(alu__abc_40887_new_n177_), .Y(alu__abc_40887_new_n178_));
INVX1 INVX1_883 ( .A(alu__abc_40887_new_n179_), .Y(alu__abc_40887_new_n180_));
INVX1 INVX1_884 ( .A(alu__abc_40887_new_n181_), .Y(alu__abc_40887_new_n182_));
INVX1 INVX1_885 ( .A(alu__abc_40887_new_n75_), .Y(alu__abc_40887_new_n183_));
INVX1 INVX1_886 ( .A(alu_opra_1_), .Y(alu__abc_40887_new_n184_));
INVX1 INVX1_887 ( .A(alu__abc_40887_new_n156_), .Y(alu__abc_40887_new_n187_));
INVX1 INVX1_888 ( .A(alu__abc_40887_new_n59_), .Y(alu__abc_40887_new_n190_));
INVX1 INVX1_889 ( .A(alu__abc_40887_new_n165_), .Y(alu__abc_40887_new_n197_));
INVX1 INVX1_89 ( .A(_abc_41356_new_n1080_), .Y(_abc_41356_new_n1081_));
INVX1 INVX1_890 ( .A(alu__abc_40887_new_n199_), .Y(alu__abc_40887_new_n200_));
INVX1 INVX1_891 ( .A(alu__abc_40887_new_n149_), .Y(alu__abc_40887_new_n207_));
INVX1 INVX1_892 ( .A(alu_cin), .Y(alu__abc_40887_new_n213_));
INVX1 INVX1_893 ( .A(alu__abc_40887_new_n216_), .Y(alu__abc_40887_new_n217_));
INVX1 INVX1_894 ( .A(alu__abc_40887_new_n218_), .Y(alu__abc_40887_new_n219_));
INVX1 INVX1_895 ( .A(alu__abc_40887_new_n224_), .Y(alu__abc_40887_new_n226_));
INVX1 INVX1_896 ( .A(alu_sel_0_), .Y(alu__abc_40887_new_n230_));
INVX1 INVX1_897 ( .A(alu__abc_40887_new_n131_), .Y(alu__abc_40887_new_n251_));
INVX1 INVX1_898 ( .A(alu__abc_40887_new_n252_), .Y(alu__abc_40887_new_n253_));
INVX1 INVX1_899 ( .A(alu__abc_40887_new_n220_), .Y(alu__abc_40887_new_n259_));
INVX1 INVX1_9 ( .A(state_0_), .Y(_abc_41356_new_n520_));
INVX1 INVX1_90 ( .A(_abc_41356_new_n603_), .Y(_abc_41356_new_n1082_));
INVX1 INVX1_900 ( .A(alu__abc_40887_new_n202_), .Y(alu__abc_40887_new_n261_));
INVX1 INVX1_901 ( .A(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n279_));
INVX1 INVX1_902 ( .A(alu__abc_40887_new_n227_), .Y(alu__abc_40887_new_n281_));
INVX1 INVX1_903 ( .A(alu__abc_40887_new_n248_), .Y(alu__abc_40887_new_n284_));
INVX1 INVX1_904 ( .A(alu__abc_40887_new_n277_), .Y(alu__abc_40887_new_n287_));
INVX1 INVX1_905 ( .A(alu__abc_40887_new_n292_), .Y(alu__abc_40887_new_n293_));
INVX1 INVX1_906 ( .A(alu__abc_40887_new_n121_), .Y(alu__abc_40887_new_n297_));
INVX1 INVX1_907 ( .A(alu__abc_40887_new_n298_), .Y(alu__abc_40887_new_n299_));
INVX1 INVX1_908 ( .A(alu__abc_40887_new_n122_), .Y(alu__abc_40887_new_n300_));
INVX1 INVX1_909 ( .A(alu__abc_40887_new_n120_), .Y(alu__abc_40887_new_n314_));
INVX1 INVX1_91 ( .A(_abc_41356_new_n1083_), .Y(_abc_41356_new_n1084_));
INVX1 INVX1_910 ( .A(alu__abc_40887_new_n237_), .Y(alu__abc_40887_new_n315_));
INVX1 INVX1_911 ( .A(alu__abc_40887_new_n243_), .Y(alu__abc_40887_new_n316_));
INVX1 INVX1_912 ( .A(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n317_));
INVX1 INVX1_913 ( .A(alu__abc_40887_new_n327_), .Y(alu__abc_40887_new_n328_));
INVX1 INVX1_914 ( .A(alu__abc_40887_new_n330_), .Y(alu__abc_40887_new_n331_));
INVX1 INVX1_915 ( .A(alu__abc_40887_new_n333_), .Y(alu__abc_40887_new_n334_));
INVX1 INVX1_916 ( .A(alu__abc_40887_new_n335_), .Y(alu__abc_40887_new_n336_));
INVX1 INVX1_917 ( .A(alu__abc_40887_new_n113_), .Y(alu__abc_40887_new_n337_));
INVX1 INVX1_918 ( .A(alu__abc_40887_new_n126_), .Y(alu__abc_40887_new_n339_));
INVX1 INVX1_919 ( .A(alu__abc_40887_new_n340_), .Y(alu__abc_40887_new_n341_));
INVX1 INVX1_92 ( .A(_abc_41356_new_n1091_), .Y(_abc_41356_new_n1092_));
INVX1 INVX1_920 ( .A(alu__abc_40887_new_n127_), .Y(alu__abc_40887_new_n342_));
INVX1 INVX1_921 ( .A(alu__abc_40887_new_n212_), .Y(alu__abc_40887_new_n359_));
INVX1 INVX1_922 ( .A(alu__abc_40887_new_n125_), .Y(alu__abc_40887_new_n363_));
INVX1 INVX1_923 ( .A(alu__abc_40887_new_n364_), .Y(alu__abc_40887_new_n365_));
INVX1 INVX1_924 ( .A(alu__abc_40887_new_n379_), .Y(alu__abc_40887_new_n380_));
INVX1 INVX1_925 ( .A(alu__abc_40887_new_n381_), .Y(alu__abc_40887_new_n384_));
INVX1 INVX1_926 ( .A(alu__abc_40887_new_n388_), .Y(alu__abc_40887_new_n389_));
INVX1 INVX1_927 ( .A(alu__abc_40887_new_n391_), .Y(alu__abc_40887_new_n392_));
INVX1 INVX1_928 ( .A(alu__abc_40887_new_n108_), .Y(alu__abc_40887_new_n407_));
INVX1 INVX1_929 ( .A(alu__abc_40887_new_n408_), .Y(alu__abc_40887_new_n409_));
INVX1 INVX1_93 ( .A(rdatahold_6_), .Y(_abc_41356_new_n1097_));
INVX1 INVX1_930 ( .A(alu__abc_40887_new_n129_), .Y(alu__abc_40887_new_n411_));
INVX1 INVX1_931 ( .A(alu__abc_40887_new_n427_), .Y(alu__abc_40887_new_n428_));
INVX1 INVX1_932 ( .A(alu__abc_40887_new_n429_), .Y(alu__abc_40887_new_n430_));
INVX1 INVX1_933 ( .A(alu__abc_40887_new_n404_), .Y(alu__abc_40887_new_n435_));
INVX1 INVX1_934 ( .A(alu__abc_40887_new_n236_), .Y(alu__abc_40887_new_n462_));
INVX1 INVX1_935 ( .A(alu_opra_7_), .Y(alu__abc_40887_new_n487_));
INVX1 INVX1_94 ( .A(_abc_41356_new_n512_), .Y(_abc_41356_new_n1099_));
INVX1 INVX1_95 ( .A(_abc_41356_new_n555_), .Y(_abc_41356_new_n1103_));
INVX1 INVX1_96 ( .A(_abc_41356_new_n1104_), .Y(_abc_41356_new_n1105_));
INVX1 INVX1_97 ( .A(_abc_41356_new_n1107_), .Y(_abc_41356_new_n1108_));
INVX1 INVX1_98 ( .A(_abc_41356_new_n1109_), .Y(_abc_41356_new_n1110_));
INVX1 INVX1_99 ( .A(regfil_7__7_), .Y(_abc_41356_new_n1117_));
OR2X2 OR2X2_1 ( .A(_abc_41356_new_n541_), .B(_abc_41356_new_n539_), .Y(_abc_41356_new_n542_));
OR2X2 OR2X2_10 ( .A(_abc_41356_new_n620_), .B(_abc_41356_new_n617_), .Y(_abc_41356_new_n621_));
OR2X2 OR2X2_100 ( .A(_abc_41356_new_n862_), .B(_abc_41356_new_n863_), .Y(_abc_41356_new_n864_));
OR2X2 OR2X2_1000 ( .A(_abc_41356_new_n3411_), .B(statesel_0_), .Y(_abc_41356_new_n3412_));
OR2X2 OR2X2_1001 ( .A(_abc_41356_new_n3369_), .B(_abc_41356_new_n3408_), .Y(_abc_41356_new_n3415_));
OR2X2 OR2X2_1002 ( .A(_abc_41356_new_n3415_), .B(_abc_41356_new_n3414_), .Y(_abc_41356_new_n3416_));
OR2X2 OR2X2_1003 ( .A(_abc_41356_new_n3417_), .B(_abc_41356_new_n3413_), .Y(_abc_41356_new_n3418_));
OR2X2 OR2X2_1004 ( .A(_abc_41356_new_n3407_), .B(_abc_41356_new_n3418_), .Y(_abc_41356_new_n3419_));
OR2X2 OR2X2_1005 ( .A(_abc_41356_new_n3419_), .B(_abc_41356_new_n3390_), .Y(_abc_41356_new_n3420_));
OR2X2 OR2X2_1006 ( .A(_abc_41356_new_n3014_), .B(_abc_41356_new_n1163_), .Y(_abc_41356_new_n3422_));
OR2X2 OR2X2_1007 ( .A(_abc_41356_new_n3425_), .B(_abc_41356_new_n3427_), .Y(_abc_41356_new_n3428_));
OR2X2 OR2X2_1008 ( .A(_abc_41356_new_n3428_), .B(_abc_41356_new_n3424_), .Y(_abc_41356_new_n3429_));
OR2X2 OR2X2_1009 ( .A(_abc_41356_new_n3430_), .B(_abc_41356_new_n3432_), .Y(_abc_41356_new_n3433_));
OR2X2 OR2X2_101 ( .A(_abc_41356_new_n866_), .B(_abc_41356_new_n865_), .Y(_abc_41356_new_n867_));
OR2X2 OR2X2_1010 ( .A(_abc_41356_new_n3434_), .B(_abc_41356_new_n2924_), .Y(_abc_41356_new_n3435_));
OR2X2 OR2X2_1011 ( .A(_abc_41356_new_n3435_), .B(_abc_41356_new_n3433_), .Y(_abc_41356_new_n3436_));
OR2X2 OR2X2_1012 ( .A(_abc_41356_new_n3436_), .B(_abc_41356_new_n3429_), .Y(_abc_41356_new_n3437_));
OR2X2 OR2X2_1013 ( .A(_abc_41356_new_n3437_), .B(_abc_41356_new_n3422_), .Y(_abc_41356_new_n3438_));
OR2X2 OR2X2_1014 ( .A(_abc_41356_new_n3443_), .B(reset), .Y(_abc_41356_new_n3444_));
OR2X2 OR2X2_1015 ( .A(_abc_41356_new_n3444_), .B(_abc_41356_new_n3446_), .Y(_abc_41356_new_n3447_));
OR2X2 OR2X2_1016 ( .A(_abc_41356_new_n3438_), .B(_abc_41356_new_n3450_), .Y(_abc_41356_new_n3451_));
OR2X2 OR2X2_1017 ( .A(_abc_41356_new_n3452_), .B(reset), .Y(_abc_41356_new_n3453_));
OR2X2 OR2X2_1018 ( .A(_abc_41356_new_n3448_), .B(_abc_41356_new_n3455_), .Y(_abc_41356_new_n3456_));
OR2X2 OR2X2_1019 ( .A(_abc_41356_new_n3421_), .B(_abc_41356_new_n3456_), .Y(_0statesel_5_0__0_));
OR2X2 OR2X2_102 ( .A(_abc_41356_new_n864_), .B(_abc_41356_new_n867_), .Y(_abc_41356_new_n868_));
OR2X2 OR2X2_1020 ( .A(_abc_41356_new_n3378_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n3459_));
OR2X2 OR2X2_1021 ( .A(_abc_41356_new_n3458_), .B(_abc_41356_new_n3459_), .Y(_abc_41356_new_n3460_));
OR2X2 OR2X2_1022 ( .A(_abc_41356_new_n3401_), .B(_abc_41356_new_n3462_), .Y(_abc_41356_new_n3463_));
OR2X2 OR2X2_1023 ( .A(_abc_41356_new_n3408_), .B(_abc_41356_new_n3466_), .Y(_abc_41356_new_n3467_));
OR2X2 OR2X2_1024 ( .A(_abc_41356_new_n3467_), .B(_abc_41356_new_n3465_), .Y(_abc_41356_new_n3468_));
OR2X2 OR2X2_1025 ( .A(_abc_41356_new_n3468_), .B(_abc_41356_new_n3373_), .Y(_abc_41356_new_n3469_));
OR2X2 OR2X2_1026 ( .A(_abc_41356_new_n3464_), .B(_abc_41356_new_n3469_), .Y(_abc_41356_new_n3470_));
OR2X2 OR2X2_1027 ( .A(_abc_41356_new_n677_), .B(statesel_1_), .Y(_abc_41356_new_n3472_));
OR2X2 OR2X2_1028 ( .A(_abc_41356_new_n3408_), .B(statesel_1_), .Y(_abc_41356_new_n3474_));
OR2X2 OR2X2_1029 ( .A(_abc_41356_new_n3477_), .B(_abc_41356_new_n3473_), .Y(_abc_41356_new_n3478_));
OR2X2 OR2X2_103 ( .A(_abc_41356_new_n868_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n869_));
OR2X2 OR2X2_1030 ( .A(_abc_41356_new_n3471_), .B(_abc_41356_new_n3478_), .Y(_abc_41356_new_n3479_));
OR2X2 OR2X2_1031 ( .A(_abc_41356_new_n3461_), .B(_abc_41356_new_n3479_), .Y(_abc_41356_new_n3480_));
OR2X2 OR2X2_1032 ( .A(_abc_41356_new_n3481_), .B(_abc_41356_new_n3483_), .Y(_abc_41356_new_n3484_));
OR2X2 OR2X2_1033 ( .A(_abc_41356_new_n3487_), .B(_abc_41356_new_n3489_), .Y(_abc_41356_new_n3490_));
OR2X2 OR2X2_1034 ( .A(_abc_41356_new_n3491_), .B(_abc_41356_new_n3486_), .Y(_abc_41356_new_n3492_));
OR2X2 OR2X2_1035 ( .A(_abc_41356_new_n3485_), .B(_abc_41356_new_n3492_), .Y(_0statesel_5_0__1_));
OR2X2 OR2X2_1036 ( .A(_abc_41356_new_n3378_), .B(_abc_41356_new_n3495_), .Y(_abc_41356_new_n3496_));
OR2X2 OR2X2_1037 ( .A(_abc_41356_new_n3384_), .B(_abc_41356_new_n3496_), .Y(_abc_41356_new_n3497_));
OR2X2 OR2X2_1038 ( .A(_abc_41356_new_n3498_), .B(_abc_41356_new_n3497_), .Y(_abc_41356_new_n3499_));
OR2X2 OR2X2_1039 ( .A(_abc_41356_new_n682_), .B(statesel_2_), .Y(_abc_41356_new_n3501_));
OR2X2 OR2X2_104 ( .A(_abc_41356_new_n870_), .B(_abc_41356_new_n871_), .Y(_abc_41356_new_n872_));
OR2X2 OR2X2_1040 ( .A(_abc_41356_new_n3394_), .B(_abc_41356_new_n677_), .Y(_abc_41356_new_n3504_));
OR2X2 OR2X2_1041 ( .A(_abc_41356_new_n3504_), .B(_abc_41356_new_n3503_), .Y(_abc_41356_new_n3505_));
OR2X2 OR2X2_1042 ( .A(_abc_41356_new_n3502_), .B(_abc_41356_new_n3505_), .Y(_abc_41356_new_n3506_));
OR2X2 OR2X2_1043 ( .A(_abc_41356_new_n3400_), .B(statesel_2_), .Y(_abc_41356_new_n3507_));
OR2X2 OR2X2_1044 ( .A(_abc_41356_new_n3510_), .B(_abc_41356_new_n3391_), .Y(_abc_41356_new_n3511_));
OR2X2 OR2X2_1045 ( .A(_abc_41356_new_n3509_), .B(_abc_41356_new_n3512_), .Y(_abc_41356_new_n3513_));
OR2X2 OR2X2_1046 ( .A(_abc_41356_new_n3500_), .B(_abc_41356_new_n3513_), .Y(_abc_41356_new_n3514_));
OR2X2 OR2X2_1047 ( .A(_abc_41356_new_n3515_), .B(_abc_41356_new_n3516_), .Y(_abc_41356_new_n3517_));
OR2X2 OR2X2_1048 ( .A(_abc_41356_new_n3523_), .B(_abc_41356_new_n3524_), .Y(_abc_41356_new_n3525_));
OR2X2 OR2X2_1049 ( .A(_abc_41356_new_n3520_), .B(statesel_2_), .Y(_abc_41356_new_n3526_));
OR2X2 OR2X2_105 ( .A(_abc_41356_new_n874_), .B(_abc_41356_new_n873_), .Y(_abc_41356_new_n875_));
OR2X2 OR2X2_1050 ( .A(_abc_41356_new_n3519_), .B(_abc_41356_new_n3528_), .Y(_abc_41356_new_n3529_));
OR2X2 OR2X2_1051 ( .A(_abc_41356_new_n3518_), .B(_abc_41356_new_n3529_), .Y(_0statesel_5_0__2_));
OR2X2 OR2X2_1052 ( .A(_abc_41356_new_n3534_), .B(_abc_41356_new_n3533_), .Y(_abc_41356_new_n3535_));
OR2X2 OR2X2_1053 ( .A(_abc_41356_new_n3532_), .B(_abc_41356_new_n3535_), .Y(_abc_41356_new_n3536_));
OR2X2 OR2X2_1054 ( .A(_abc_41356_new_n3395_), .B(_abc_41356_new_n677_), .Y(_abc_41356_new_n3538_));
OR2X2 OR2X2_1055 ( .A(_abc_41356_new_n3538_), .B(_abc_41356_new_n3465_), .Y(_abc_41356_new_n3539_));
OR2X2 OR2X2_1056 ( .A(_abc_41356_new_n682_), .B(statesel_3_), .Y(_abc_41356_new_n3540_));
OR2X2 OR2X2_1057 ( .A(_abc_41356_new_n3541_), .B(_abc_41356_new_n3539_), .Y(_abc_41356_new_n3542_));
OR2X2 OR2X2_1058 ( .A(_abc_41356_new_n3400_), .B(statesel_3_), .Y(_abc_41356_new_n3543_));
OR2X2 OR2X2_1059 ( .A(_abc_41356_new_n3546_), .B(statesel_3_), .Y(_abc_41356_new_n3547_));
OR2X2 OR2X2_106 ( .A(_abc_41356_new_n872_), .B(_abc_41356_new_n875_), .Y(_abc_41356_new_n876_));
OR2X2 OR2X2_1060 ( .A(_abc_41356_new_n3510_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n3548_));
OR2X2 OR2X2_1061 ( .A(_abc_41356_new_n3545_), .B(_abc_41356_new_n3549_), .Y(_abc_41356_new_n3550_));
OR2X2 OR2X2_1062 ( .A(_abc_41356_new_n3537_), .B(_abc_41356_new_n3550_), .Y(_abc_41356_new_n3551_));
OR2X2 OR2X2_1063 ( .A(_abc_41356_new_n3482_), .B(_abc_41356_new_n3557_), .Y(_abc_41356_new_n3558_));
OR2X2 OR2X2_1064 ( .A(_abc_41356_new_n3523_), .B(_abc_41356_new_n3558_), .Y(_abc_41356_new_n3559_));
OR2X2 OR2X2_1065 ( .A(_abc_41356_new_n3560_), .B(_abc_41356_new_n3556_), .Y(_abc_41356_new_n3561_));
OR2X2 OR2X2_1066 ( .A(_abc_41356_new_n3552_), .B(_abc_41356_new_n3561_), .Y(_abc_41356_new_n3562_));
OR2X2 OR2X2_1067 ( .A(_abc_41356_new_n3563_), .B(_abc_41356_new_n3531_), .Y(_0statesel_5_0__3_));
OR2X2 OR2X2_1068 ( .A(_abc_41356_new_n3567_), .B(_abc_41356_new_n3566_), .Y(_abc_41356_new_n3568_));
OR2X2 OR2X2_1069 ( .A(_abc_41356_new_n3403_), .B(_abc_41356_new_n3548_), .Y(_abc_41356_new_n3570_));
OR2X2 OR2X2_107 ( .A(_abc_41356_new_n876_), .B(opcode_2_), .Y(_abc_41356_new_n877_));
OR2X2 OR2X2_1070 ( .A(_abc_41356_new_n3392_), .B(_abc_41356_new_n3572_), .Y(_abc_41356_new_n3573_));
OR2X2 OR2X2_1071 ( .A(_abc_41356_new_n3574_), .B(_abc_41356_new_n3546_), .Y(_abc_41356_new_n3575_));
OR2X2 OR2X2_1072 ( .A(_abc_41356_new_n3571_), .B(_abc_41356_new_n3575_), .Y(_abc_41356_new_n3576_));
OR2X2 OR2X2_1073 ( .A(_abc_41356_new_n3576_), .B(_abc_41356_new_n3569_), .Y(_abc_41356_new_n3577_));
OR2X2 OR2X2_1074 ( .A(_abc_41356_new_n3581_), .B(statesel_4_), .Y(_abc_41356_new_n3582_));
OR2X2 OR2X2_1075 ( .A(_abc_41356_new_n3585_), .B(_abc_41356_new_n3586_), .Y(_abc_41356_new_n3587_));
OR2X2 OR2X2_1076 ( .A(_abc_41356_new_n3588_), .B(_abc_41356_new_n3579_), .Y(_abc_41356_new_n3589_));
OR2X2 OR2X2_1077 ( .A(_abc_41356_new_n3578_), .B(_abc_41356_new_n3589_), .Y(_abc_41356_new_n3590_));
OR2X2 OR2X2_1078 ( .A(_abc_41356_new_n3591_), .B(_abc_41356_new_n3565_), .Y(_0statesel_5_0__4_));
OR2X2 OR2X2_1079 ( .A(_abc_41356_new_n3599_), .B(_abc_41356_new_n3546_), .Y(_abc_41356_new_n3600_));
OR2X2 OR2X2_108 ( .A(_abc_41356_new_n879_), .B(_abc_41356_new_n880_), .Y(_abc_41356_new_n881_));
OR2X2 OR2X2_1080 ( .A(_abc_41356_new_n3598_), .B(_abc_41356_new_n3600_), .Y(_abc_41356_new_n3601_));
OR2X2 OR2X2_1081 ( .A(_abc_41356_new_n3597_), .B(_abc_41356_new_n3601_), .Y(_abc_41356_new_n3602_));
OR2X2 OR2X2_1082 ( .A(_abc_41356_new_n3604_), .B(_abc_41356_new_n3482_), .Y(_abc_41356_new_n3605_));
OR2X2 OR2X2_1083 ( .A(_abc_41356_new_n3585_), .B(_abc_41356_new_n3605_), .Y(_abc_41356_new_n3606_));
OR2X2 OR2X2_1084 ( .A(_abc_41356_new_n3607_), .B(_abc_41356_new_n3610_), .Y(_abc_41356_new_n3611_));
OR2X2 OR2X2_1085 ( .A(_abc_41356_new_n3603_), .B(_abc_41356_new_n3611_), .Y(_abc_41356_new_n3612_));
OR2X2 OR2X2_1086 ( .A(_abc_41356_new_n3613_), .B(_abc_41356_new_n3593_), .Y(_0statesel_5_0__5_));
OR2X2 OR2X2_1087 ( .A(_abc_41356_new_n3616_), .B(opcode_4_), .Y(_abc_41356_new_n3617_));
OR2X2 OR2X2_1088 ( .A(_abc_41356_new_n3615_), .B(popdes_0_), .Y(_abc_41356_new_n3618_));
OR2X2 OR2X2_1089 ( .A(_abc_41356_new_n3616_), .B(opcode_5_), .Y(_abc_41356_new_n3620_));
OR2X2 OR2X2_109 ( .A(_abc_41356_new_n882_), .B(_abc_41356_new_n861_), .Y(_abc_41356_new_n883_));
OR2X2 OR2X2_1090 ( .A(_abc_41356_new_n3615_), .B(popdes_1_), .Y(_abc_41356_new_n3621_));
OR2X2 OR2X2_1091 ( .A(_abc_41356_new_n3623_), .B(rdatahold2_0_), .Y(_abc_41356_new_n3624_));
OR2X2 OR2X2_1092 ( .A(_abc_41356_new_n3623_), .B(rdatahold2_1_), .Y(_abc_41356_new_n3628_));
OR2X2 OR2X2_1093 ( .A(_abc_41356_new_n3623_), .B(rdatahold2_2_), .Y(_abc_41356_new_n3633_));
OR2X2 OR2X2_1094 ( .A(_abc_41356_new_n3623_), .B(rdatahold2_3_), .Y(_abc_41356_new_n3637_));
OR2X2 OR2X2_1095 ( .A(_abc_41356_new_n3623_), .B(rdatahold2_4_), .Y(_abc_41356_new_n3641_));
OR2X2 OR2X2_1096 ( .A(_abc_41356_new_n3623_), .B(rdatahold2_5_), .Y(_abc_41356_new_n3646_));
OR2X2 OR2X2_1097 ( .A(_abc_41356_new_n3623_), .B(rdatahold2_6_), .Y(_abc_41356_new_n3650_));
OR2X2 OR2X2_1098 ( .A(_abc_41356_new_n3623_), .B(rdatahold2_7_), .Y(_abc_41356_new_n3654_));
OR2X2 OR2X2_1099 ( .A(_abc_41356_new_n3623_), .B(rdatahold_0_), .Y(_abc_41356_new_n3658_));
OR2X2 OR2X2_11 ( .A(_abc_41356_new_n624_), .B(_abc_41356_new_n622_), .Y(_abc_41356_new_n625_));
OR2X2 OR2X2_110 ( .A(_abc_41356_new_n860_), .B(_abc_41356_new_n883_), .Y(_abc_41356_new_n884_));
OR2X2 OR2X2_1100 ( .A(_abc_41356_new_n3623_), .B(rdatahold_1_), .Y(_abc_41356_new_n3663_));
OR2X2 OR2X2_1101 ( .A(_abc_41356_new_n3623_), .B(rdatahold_2_), .Y(_abc_41356_new_n3668_));
OR2X2 OR2X2_1102 ( .A(_abc_41356_new_n3623_), .B(rdatahold_3_), .Y(_abc_41356_new_n3673_));
OR2X2 OR2X2_1103 ( .A(_abc_41356_new_n3623_), .B(rdatahold_4_), .Y(_abc_41356_new_n3678_));
OR2X2 OR2X2_1104 ( .A(_abc_41356_new_n3623_), .B(rdatahold_5_), .Y(_abc_41356_new_n3683_));
OR2X2 OR2X2_1105 ( .A(_abc_41356_new_n3623_), .B(rdatahold_6_), .Y(_abc_41356_new_n3688_));
OR2X2 OR2X2_1106 ( .A(_abc_41356_new_n3623_), .B(rdatahold_7_), .Y(_abc_41356_new_n3693_));
OR2X2 OR2X2_1107 ( .A(_abc_41356_new_n3704_), .B(reset), .Y(_abc_41356_new_n3705_));
OR2X2 OR2X2_1108 ( .A(_abc_41356_new_n3707_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n3708_));
OR2X2 OR2X2_1109 ( .A(_abc_41356_new_n3712_), .B(_abc_41356_new_n3711_), .Y(_abc_41356_new_n3713_));
OR2X2 OR2X2_111 ( .A(_abc_41356_new_n855_), .B(_abc_41356_new_n884_), .Y(_abc_41356_new_n885_));
OR2X2 OR2X2_1110 ( .A(_abc_41356_new_n3713_), .B(_abc_41356_new_n3710_), .Y(_abc_41356_new_n3714_));
OR2X2 OR2X2_1111 ( .A(_abc_41356_new_n2026_), .B(wdatahold_0_), .Y(_abc_41356_new_n3715_));
OR2X2 OR2X2_1112 ( .A(_abc_41356_new_n636_), .B(_abc_41356_new_n3475_), .Y(_abc_41356_new_n3718_));
OR2X2 OR2X2_1113 ( .A(_abc_41356_new_n3411_), .B(wdatahold_0_), .Y(_abc_41356_new_n3719_));
OR2X2 OR2X2_1114 ( .A(_abc_41356_new_n3721_), .B(_abc_41356_new_n3717_), .Y(_abc_41356_new_n3722_));
OR2X2 OR2X2_1115 ( .A(_abc_41356_new_n3727_), .B(_abc_41356_new_n3726_), .Y(_abc_41356_new_n3728_));
OR2X2 OR2X2_1116 ( .A(_abc_41356_new_n3711_), .B(_abc_41356_new_n3730_), .Y(_abc_41356_new_n3731_));
OR2X2 OR2X2_1117 ( .A(_abc_41356_new_n534_), .B(regfil_3__0_), .Y(_abc_41356_new_n3732_));
OR2X2 OR2X2_1118 ( .A(_abc_41356_new_n3731_), .B(_abc_41356_new_n3733_), .Y(_abc_41356_new_n3734_));
OR2X2 OR2X2_1119 ( .A(_abc_41356_new_n3735_), .B(regfil_1__0_), .Y(_abc_41356_new_n3736_));
OR2X2 OR2X2_112 ( .A(_abc_41356_new_n885_), .B(_abc_41356_new_n696_), .Y(_abc_41356_new_n886_));
OR2X2 OR2X2_1120 ( .A(_abc_41356_new_n3737_), .B(_abc_41356_new_n3738_), .Y(_abc_41356_new_n3739_));
OR2X2 OR2X2_1121 ( .A(_abc_41356_new_n3740_), .B(_abc_41356_new_n3729_), .Y(_abc_41356_new_n3741_));
OR2X2 OR2X2_1122 ( .A(_abc_41356_new_n3725_), .B(_abc_41356_new_n3741_), .Y(_abc_41356_new_n3742_));
OR2X2 OR2X2_1123 ( .A(_abc_41356_new_n3743_), .B(_abc_41356_new_n3722_), .Y(_abc_41356_new_n3744_));
OR2X2 OR2X2_1124 ( .A(_abc_41356_new_n3744_), .B(_abc_41356_new_n3709_), .Y(_abc_41356_new_n3745_));
OR2X2 OR2X2_1125 ( .A(_abc_41356_new_n3748_), .B(_abc_41356_new_n3749_), .Y(_abc_41356_new_n3750_));
OR2X2 OR2X2_1126 ( .A(_abc_41356_new_n3750_), .B(_abc_41356_new_n3747_), .Y(_abc_41356_new_n3751_));
OR2X2 OR2X2_1127 ( .A(_abc_41356_new_n3746_), .B(_abc_41356_new_n3751_), .Y(_abc_41356_new_n3752_));
OR2X2 OR2X2_1128 ( .A(_abc_41356_new_n3753_), .B(_abc_41356_new_n3706_), .Y(_0wdatahold_7_0__0_));
OR2X2 OR2X2_1129 ( .A(_abc_41356_new_n3476_), .B(_abc_41356_new_n3756_), .Y(_abc_41356_new_n3757_));
OR2X2 OR2X2_113 ( .A(_abc_41356_new_n695_), .B(regfil_7__3_), .Y(_abc_41356_new_n887_));
OR2X2 OR2X2_1130 ( .A(_abc_41356_new_n3707_), .B(_abc_41356_new_n3757_), .Y(_abc_41356_new_n3758_));
OR2X2 OR2X2_1131 ( .A(_abc_41356_new_n3764_), .B(intcyc), .Y(_abc_41356_new_n3765_));
OR2X2 OR2X2_1132 ( .A(_abc_41356_new_n2049_), .B(pc_1_), .Y(_abc_41356_new_n3766_));
OR2X2 OR2X2_1133 ( .A(_abc_41356_new_n3768_), .B(_abc_41356_new_n3769_), .Y(_abc_41356_new_n3770_));
OR2X2 OR2X2_1134 ( .A(_abc_41356_new_n681_), .B(_abc_41356_new_n3774_), .Y(_abc_41356_new_n3775_));
OR2X2 OR2X2_1135 ( .A(_abc_41356_new_n3773_), .B(_abc_41356_new_n3775_), .Y(_abc_41356_new_n3776_));
OR2X2 OR2X2_1136 ( .A(_abc_41356_new_n3777_), .B(_abc_41356_new_n3771_), .Y(_abc_41356_new_n3778_));
OR2X2 OR2X2_1137 ( .A(_abc_41356_new_n3779_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n3780_));
OR2X2 OR2X2_1138 ( .A(_abc_41356_new_n3770_), .B(_abc_41356_new_n3781_), .Y(_abc_41356_new_n3782_));
OR2X2 OR2X2_1139 ( .A(_abc_41356_new_n3782_), .B(_abc_41356_new_n3763_), .Y(_abc_41356_new_n3783_));
OR2X2 OR2X2_114 ( .A(_abc_41356_new_n899_), .B(_abc_41356_new_n898_), .Y(_abc_41356_new_n900_));
OR2X2 OR2X2_1140 ( .A(_abc_41356_new_n3786_), .B(_abc_41356_new_n3788_), .Y(_abc_41356_new_n3789_));
OR2X2 OR2X2_1141 ( .A(_abc_41356_new_n3792_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n3793_));
OR2X2 OR2X2_1142 ( .A(_abc_41356_new_n3793_), .B(_abc_41356_new_n3790_), .Y(_abc_41356_new_n3794_));
OR2X2 OR2X2_1143 ( .A(_abc_41356_new_n3785_), .B(_abc_41356_new_n3794_), .Y(_abc_41356_new_n3795_));
OR2X2 OR2X2_1144 ( .A(_abc_41356_new_n3795_), .B(_abc_41356_new_n3759_), .Y(_abc_41356_new_n3796_));
OR2X2 OR2X2_1145 ( .A(_abc_41356_new_n2887_), .B(wdatahold_1_), .Y(_abc_41356_new_n3797_));
OR2X2 OR2X2_1146 ( .A(_abc_41356_new_n3801_), .B(_abc_41356_new_n3802_), .Y(_abc_41356_new_n3803_));
OR2X2 OR2X2_1147 ( .A(_abc_41356_new_n3803_), .B(_abc_41356_new_n3800_), .Y(_abc_41356_new_n3804_));
OR2X2 OR2X2_1148 ( .A(_abc_41356_new_n3799_), .B(_abc_41356_new_n3804_), .Y(_abc_41356_new_n3805_));
OR2X2 OR2X2_1149 ( .A(_abc_41356_new_n3806_), .B(_abc_41356_new_n3755_), .Y(_0wdatahold_7_0__1_));
OR2X2 OR2X2_115 ( .A(_abc_41356_new_n904_), .B(_abc_41356_new_n555_), .Y(_abc_41356_new_n905_));
OR2X2 OR2X2_1150 ( .A(_abc_41356_new_n3812_), .B(_abc_41356_new_n3810_), .Y(_abc_41356_new_n3813_));
OR2X2 OR2X2_1151 ( .A(_abc_41356_new_n2049_), .B(pc_2_), .Y(_abc_41356_new_n3816_));
OR2X2 OR2X2_1152 ( .A(_abc_41356_new_n3819_), .B(_abc_41356_new_n2034_), .Y(_abc_41356_new_n3820_));
OR2X2 OR2X2_1153 ( .A(_abc_41356_new_n3821_), .B(intcyc), .Y(_abc_41356_new_n3822_));
OR2X2 OR2X2_1154 ( .A(_abc_41356_new_n534_), .B(regfil_3__2_), .Y(_abc_41356_new_n3827_));
OR2X2 OR2X2_1155 ( .A(_abc_41356_new_n3828_), .B(_abc_41356_new_n3826_), .Y(_abc_41356_new_n3829_));
OR2X2 OR2X2_1156 ( .A(_abc_41356_new_n3829_), .B(_abc_41356_new_n3825_), .Y(_abc_41356_new_n3830_));
OR2X2 OR2X2_1157 ( .A(_abc_41356_new_n3735_), .B(regfil_1__2_), .Y(_abc_41356_new_n3831_));
OR2X2 OR2X2_1158 ( .A(_abc_41356_new_n3834_), .B(_abc_41356_new_n3835_), .Y(_abc_41356_new_n3836_));
OR2X2 OR2X2_1159 ( .A(_abc_41356_new_n3836_), .B(_abc_41356_new_n3833_), .Y(_abc_41356_new_n3837_));
OR2X2 OR2X2_116 ( .A(_abc_41356_new_n906_), .B(_abc_41356_new_n530_), .Y(_abc_41356_new_n907_));
OR2X2 OR2X2_1160 ( .A(_abc_41356_new_n3837_), .B(_abc_41356_new_n3824_), .Y(_abc_41356_new_n3838_));
OR2X2 OR2X2_1161 ( .A(_abc_41356_new_n3838_), .B(_abc_41356_new_n3815_), .Y(_abc_41356_new_n3839_));
OR2X2 OR2X2_1162 ( .A(_abc_41356_new_n3809_), .B(_abc_41356_new_n3839_), .Y(_abc_41356_new_n3840_));
OR2X2 OR2X2_1163 ( .A(_abc_41356_new_n3843_), .B(_abc_41356_new_n3826_), .Y(_abc_41356_new_n3844_));
OR2X2 OR2X2_1164 ( .A(_abc_41356_new_n3844_), .B(_abc_41356_new_n3710_), .Y(_abc_41356_new_n3845_));
OR2X2 OR2X2_1165 ( .A(_abc_41356_new_n2026_), .B(wdatahold_2_), .Y(_abc_41356_new_n3846_));
OR2X2 OR2X2_1166 ( .A(_abc_41356_new_n3476_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n3849_));
OR2X2 OR2X2_1167 ( .A(_abc_41356_new_n3850_), .B(_abc_41356_new_n3848_), .Y(_abc_41356_new_n3851_));
OR2X2 OR2X2_1168 ( .A(_abc_41356_new_n3851_), .B(_abc_41356_new_n3842_), .Y(_abc_41356_new_n3852_));
OR2X2 OR2X2_1169 ( .A(_abc_41356_new_n3841_), .B(_abc_41356_new_n3852_), .Y(_abc_41356_new_n3853_));
OR2X2 OR2X2_117 ( .A(_abc_41356_new_n908_), .B(_abc_41356_new_n512_), .Y(_abc_41356_new_n909_));
OR2X2 OR2X2_1170 ( .A(_abc_41356_new_n3856_), .B(_abc_41356_new_n3857_), .Y(_abc_41356_new_n3858_));
OR2X2 OR2X2_1171 ( .A(_abc_41356_new_n3858_), .B(_abc_41356_new_n3855_), .Y(_abc_41356_new_n3859_));
OR2X2 OR2X2_1172 ( .A(_abc_41356_new_n3854_), .B(_abc_41356_new_n3859_), .Y(_abc_41356_new_n3860_));
OR2X2 OR2X2_1173 ( .A(_abc_41356_new_n3861_), .B(_abc_41356_new_n3808_), .Y(_0wdatahold_7_0__2_));
OR2X2 OR2X2_1174 ( .A(_abc_41356_new_n3866_), .B(_abc_41356_new_n3865_), .Y(_abc_41356_new_n3867_));
OR2X2 OR2X2_1175 ( .A(_abc_41356_new_n3867_), .B(_abc_41356_new_n3710_), .Y(_abc_41356_new_n3868_));
OR2X2 OR2X2_1176 ( .A(_abc_41356_new_n2026_), .B(wdatahold_3_), .Y(_abc_41356_new_n3869_));
OR2X2 OR2X2_1177 ( .A(_abc_41356_new_n878_), .B(_abc_41356_new_n3475_), .Y(_abc_41356_new_n3872_));
OR2X2 OR2X2_1178 ( .A(_abc_41356_new_n3411_), .B(wdatahold_3_), .Y(_abc_41356_new_n3873_));
OR2X2 OR2X2_1179 ( .A(_abc_41356_new_n3875_), .B(_abc_41356_new_n3871_), .Y(_abc_41356_new_n3876_));
OR2X2 OR2X2_118 ( .A(_abc_41356_new_n913_), .B(_abc_41356_new_n912_), .Y(_abc_41356_new_n914_));
OR2X2 OR2X2_1180 ( .A(_abc_41356_new_n3810_), .B(pc_3_), .Y(_abc_41356_new_n3878_));
OR2X2 OR2X2_1181 ( .A(_abc_41356_new_n2034_), .B(pc_3_), .Y(_abc_41356_new_n3882_));
OR2X2 OR2X2_1182 ( .A(_abc_41356_new_n3883_), .B(intcyc), .Y(_abc_41356_new_n3884_));
OR2X2 OR2X2_1183 ( .A(_abc_41356_new_n2049_), .B(pc_3_), .Y(_abc_41356_new_n3885_));
OR2X2 OR2X2_1184 ( .A(_abc_41356_new_n534_), .B(regfil_3__3_), .Y(_abc_41356_new_n3889_));
OR2X2 OR2X2_1185 ( .A(_abc_41356_new_n3890_), .B(_abc_41356_new_n3865_), .Y(_abc_41356_new_n3891_));
OR2X2 OR2X2_1186 ( .A(_abc_41356_new_n3735_), .B(regfil_1__3_), .Y(_abc_41356_new_n3892_));
OR2X2 OR2X2_1187 ( .A(_abc_41356_new_n3894_), .B(_abc_41356_new_n3895_), .Y(_abc_41356_new_n3896_));
OR2X2 OR2X2_1188 ( .A(_abc_41356_new_n3896_), .B(_abc_41356_new_n3888_), .Y(_abc_41356_new_n3897_));
OR2X2 OR2X2_1189 ( .A(_abc_41356_new_n3897_), .B(_abc_41356_new_n3887_), .Y(_abc_41356_new_n3898_));
OR2X2 OR2X2_119 ( .A(_abc_41356_new_n914_), .B(_abc_41356_new_n911_), .Y(_abc_41356_new_n915_));
OR2X2 OR2X2_1190 ( .A(_abc_41356_new_n3898_), .B(_abc_41356_new_n3880_), .Y(_abc_41356_new_n3899_));
OR2X2 OR2X2_1191 ( .A(_abc_41356_new_n3900_), .B(_abc_41356_new_n3876_), .Y(_abc_41356_new_n3901_));
OR2X2 OR2X2_1192 ( .A(_abc_41356_new_n3864_), .B(_abc_41356_new_n3901_), .Y(_abc_41356_new_n3902_));
OR2X2 OR2X2_1193 ( .A(_abc_41356_new_n3905_), .B(_abc_41356_new_n3906_), .Y(_abc_41356_new_n3907_));
OR2X2 OR2X2_1194 ( .A(_abc_41356_new_n3907_), .B(_abc_41356_new_n3904_), .Y(_abc_41356_new_n3908_));
OR2X2 OR2X2_1195 ( .A(_abc_41356_new_n3903_), .B(_abc_41356_new_n3908_), .Y(_abc_41356_new_n3909_));
OR2X2 OR2X2_1196 ( .A(_abc_41356_new_n3910_), .B(_abc_41356_new_n3863_), .Y(_0wdatahold_7_0__3_));
OR2X2 OR2X2_1197 ( .A(_abc_41356_new_n3915_), .B(_abc_41356_new_n3914_), .Y(_abc_41356_new_n3916_));
OR2X2 OR2X2_1198 ( .A(_abc_41356_new_n3916_), .B(_abc_41356_new_n3710_), .Y(_abc_41356_new_n3917_));
OR2X2 OR2X2_1199 ( .A(_abc_41356_new_n2026_), .B(wdatahold_4_), .Y(_abc_41356_new_n3918_));
OR2X2 OR2X2_12 ( .A(_abc_41356_new_n621_), .B(_abc_41356_new_n625_), .Y(_abc_41356_new_n626_));
OR2X2 OR2X2_120 ( .A(_abc_41356_new_n910_), .B(_abc_41356_new_n915_), .Y(_abc_41356_new_n916_));
OR2X2 OR2X2_1200 ( .A(_abc_41356_new_n945_), .B(_abc_41356_new_n3475_), .Y(_abc_41356_new_n3921_));
OR2X2 OR2X2_1201 ( .A(_abc_41356_new_n3411_), .B(wdatahold_4_), .Y(_abc_41356_new_n3922_));
OR2X2 OR2X2_1202 ( .A(_abc_41356_new_n3924_), .B(_abc_41356_new_n3920_), .Y(_abc_41356_new_n3925_));
OR2X2 OR2X2_1203 ( .A(_abc_41356_new_n2072_), .B(pc_4_), .Y(_abc_41356_new_n3928_));
OR2X2 OR2X2_1204 ( .A(_abc_41356_new_n2035_), .B(pc_4_), .Y(_abc_41356_new_n3933_));
OR2X2 OR2X2_1205 ( .A(_abc_41356_new_n3934_), .B(intcyc), .Y(_abc_41356_new_n3935_));
OR2X2 OR2X2_1206 ( .A(_abc_41356_new_n2049_), .B(pc_4_), .Y(_abc_41356_new_n3936_));
OR2X2 OR2X2_1207 ( .A(_abc_41356_new_n3914_), .B(_abc_41356_new_n3940_), .Y(_abc_41356_new_n3941_));
OR2X2 OR2X2_1208 ( .A(_abc_41356_new_n534_), .B(regfil_3__4_), .Y(_abc_41356_new_n3942_));
OR2X2 OR2X2_1209 ( .A(_abc_41356_new_n3941_), .B(_abc_41356_new_n3943_), .Y(_abc_41356_new_n3944_));
OR2X2 OR2X2_121 ( .A(_abc_41356_new_n889_), .B(_abc_41356_new_n916_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_3_));
OR2X2 OR2X2_1210 ( .A(_abc_41356_new_n3735_), .B(regfil_1__4_), .Y(_abc_41356_new_n3945_));
OR2X2 OR2X2_1211 ( .A(_abc_41356_new_n3947_), .B(_abc_41356_new_n3948_), .Y(_abc_41356_new_n3949_));
OR2X2 OR2X2_1212 ( .A(_abc_41356_new_n3949_), .B(_abc_41356_new_n3939_), .Y(_abc_41356_new_n3950_));
OR2X2 OR2X2_1213 ( .A(_abc_41356_new_n3950_), .B(_abc_41356_new_n3938_), .Y(_abc_41356_new_n3951_));
OR2X2 OR2X2_1214 ( .A(_abc_41356_new_n3951_), .B(_abc_41356_new_n3930_), .Y(_abc_41356_new_n3952_));
OR2X2 OR2X2_1215 ( .A(_abc_41356_new_n3953_), .B(_abc_41356_new_n3925_), .Y(_abc_41356_new_n3954_));
OR2X2 OR2X2_1216 ( .A(_abc_41356_new_n3913_), .B(_abc_41356_new_n3954_), .Y(_abc_41356_new_n3955_));
OR2X2 OR2X2_1217 ( .A(_abc_41356_new_n3958_), .B(_abc_41356_new_n3959_), .Y(_abc_41356_new_n3960_));
OR2X2 OR2X2_1218 ( .A(_abc_41356_new_n3960_), .B(_abc_41356_new_n3957_), .Y(_abc_41356_new_n3961_));
OR2X2 OR2X2_1219 ( .A(_abc_41356_new_n3956_), .B(_abc_41356_new_n3961_), .Y(_abc_41356_new_n3962_));
OR2X2 OR2X2_122 ( .A(_abc_41356_new_n851_), .B(regfil_0__4_), .Y(_abc_41356_new_n918_));
OR2X2 OR2X2_1220 ( .A(_abc_41356_new_n3963_), .B(_abc_41356_new_n3912_), .Y(_0wdatahold_7_0__4_));
OR2X2 OR2X2_1221 ( .A(_abc_41356_new_n3968_), .B(_abc_41356_new_n3967_), .Y(_abc_41356_new_n3969_));
OR2X2 OR2X2_1222 ( .A(_abc_41356_new_n3969_), .B(_abc_41356_new_n3710_), .Y(_abc_41356_new_n3970_));
OR2X2 OR2X2_1223 ( .A(_abc_41356_new_n2026_), .B(wdatahold_5_), .Y(_abc_41356_new_n3971_));
OR2X2 OR2X2_1224 ( .A(_abc_41356_new_n1012_), .B(_abc_41356_new_n3475_), .Y(_abc_41356_new_n3974_));
OR2X2 OR2X2_1225 ( .A(_abc_41356_new_n3411_), .B(wdatahold_5_), .Y(_abc_41356_new_n3975_));
OR2X2 OR2X2_1226 ( .A(_abc_41356_new_n3977_), .B(_abc_41356_new_n3973_), .Y(_abc_41356_new_n3978_));
OR2X2 OR2X2_1227 ( .A(_abc_41356_new_n3981_), .B(_abc_41356_new_n3979_), .Y(_abc_41356_new_n3982_));
OR2X2 OR2X2_1228 ( .A(_abc_41356_new_n3986_), .B(_abc_41356_new_n3985_), .Y(_abc_41356_new_n3987_));
OR2X2 OR2X2_1229 ( .A(_abc_41356_new_n2049_), .B(pc_5_), .Y(_abc_41356_new_n3989_));
OR2X2 OR2X2_123 ( .A(_abc_41356_new_n919_), .B(_abc_41356_new_n920_), .Y(_abc_41356_new_n921_));
OR2X2 OR2X2_1230 ( .A(_abc_41356_new_n3988_), .B(_abc_41356_new_n3991_), .Y(_abc_41356_new_n3992_));
OR2X2 OR2X2_1231 ( .A(_abc_41356_new_n3990_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n3993_));
OR2X2 OR2X2_1232 ( .A(_abc_41356_new_n534_), .B(regfil_3__5_), .Y(_abc_41356_new_n3995_));
OR2X2 OR2X2_1233 ( .A(_abc_41356_new_n3996_), .B(_abc_41356_new_n3967_), .Y(_abc_41356_new_n3997_));
OR2X2 OR2X2_1234 ( .A(_abc_41356_new_n3735_), .B(regfil_1__5_), .Y(_abc_41356_new_n3998_));
OR2X2 OR2X2_1235 ( .A(_abc_41356_new_n4000_), .B(_abc_41356_new_n4001_), .Y(_abc_41356_new_n4002_));
OR2X2 OR2X2_1236 ( .A(_abc_41356_new_n3994_), .B(_abc_41356_new_n4002_), .Y(_abc_41356_new_n4003_));
OR2X2 OR2X2_1237 ( .A(_abc_41356_new_n4003_), .B(_abc_41356_new_n3984_), .Y(_abc_41356_new_n4004_));
OR2X2 OR2X2_1238 ( .A(_abc_41356_new_n4005_), .B(_abc_41356_new_n3978_), .Y(_abc_41356_new_n4006_));
OR2X2 OR2X2_1239 ( .A(_abc_41356_new_n4006_), .B(_abc_41356_new_n3966_), .Y(_abc_41356_new_n4007_));
OR2X2 OR2X2_124 ( .A(_abc_41356_new_n857_), .B(regfil_0__4_), .Y(_abc_41356_new_n923_));
OR2X2 OR2X2_1240 ( .A(_abc_41356_new_n4010_), .B(_abc_41356_new_n4011_), .Y(_abc_41356_new_n4012_));
OR2X2 OR2X2_1241 ( .A(_abc_41356_new_n4012_), .B(_abc_41356_new_n4009_), .Y(_abc_41356_new_n4013_));
OR2X2 OR2X2_1242 ( .A(_abc_41356_new_n4008_), .B(_abc_41356_new_n4013_), .Y(_abc_41356_new_n4014_));
OR2X2 OR2X2_1243 ( .A(_abc_41356_new_n4015_), .B(_abc_41356_new_n3965_), .Y(_0wdatahold_7_0__5_));
OR2X2 OR2X2_1244 ( .A(_abc_41356_new_n3707_), .B(_abc_41356_new_n3849_), .Y(_abc_41356_new_n4018_));
OR2X2 OR2X2_1245 ( .A(_abc_41356_new_n3979_), .B(pc_6_), .Y(_abc_41356_new_n4022_));
OR2X2 OR2X2_1246 ( .A(_abc_41356_new_n3985_), .B(pc_6_), .Y(_abc_41356_new_n4027_));
OR2X2 OR2X2_1247 ( .A(_abc_41356_new_n4029_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n4030_));
OR2X2 OR2X2_1248 ( .A(_abc_41356_new_n534_), .B(regfil_3__6_), .Y(_abc_41356_new_n4034_));
OR2X2 OR2X2_1249 ( .A(_abc_41356_new_n4035_), .B(_abc_41356_new_n4033_), .Y(_abc_41356_new_n4036_));
OR2X2 OR2X2_125 ( .A(_abc_41356_new_n930_), .B(_abc_41356_new_n929_), .Y(_abc_41356_new_n931_));
OR2X2 OR2X2_1250 ( .A(_abc_41356_new_n4036_), .B(_abc_41356_new_n4032_), .Y(_abc_41356_new_n4037_));
OR2X2 OR2X2_1251 ( .A(_abc_41356_new_n3735_), .B(regfil_1__6_), .Y(_abc_41356_new_n4038_));
OR2X2 OR2X2_1252 ( .A(_abc_41356_new_n4043_), .B(_abc_41356_new_n4041_), .Y(_abc_41356_new_n4044_));
OR2X2 OR2X2_1253 ( .A(_abc_41356_new_n4040_), .B(_abc_41356_new_n4044_), .Y(_abc_41356_new_n4045_));
OR2X2 OR2X2_1254 ( .A(_abc_41356_new_n4031_), .B(_abc_41356_new_n4045_), .Y(_abc_41356_new_n4046_));
OR2X2 OR2X2_1255 ( .A(_abc_41356_new_n4046_), .B(_abc_41356_new_n4024_), .Y(_abc_41356_new_n4047_));
OR2X2 OR2X2_1256 ( .A(_abc_41356_new_n4049_), .B(_abc_41356_new_n4033_), .Y(_abc_41356_new_n4050_));
OR2X2 OR2X2_1257 ( .A(_abc_41356_new_n4050_), .B(_abc_41356_new_n3710_), .Y(_abc_41356_new_n4051_));
OR2X2 OR2X2_1258 ( .A(_abc_41356_new_n2026_), .B(wdatahold_6_), .Y(_abc_41356_new_n4052_));
OR2X2 OR2X2_1259 ( .A(_abc_41356_new_n4055_), .B(_abc_41356_new_n4054_), .Y(_abc_41356_new_n4056_));
OR2X2 OR2X2_126 ( .A(_abc_41356_new_n933_), .B(_abc_41356_new_n932_), .Y(_abc_41356_new_n934_));
OR2X2 OR2X2_1260 ( .A(_abc_41356_new_n4048_), .B(_abc_41356_new_n4056_), .Y(_abc_41356_new_n4057_));
OR2X2 OR2X2_1261 ( .A(_abc_41356_new_n4019_), .B(_abc_41356_new_n4057_), .Y(_abc_41356_new_n4058_));
OR2X2 OR2X2_1262 ( .A(_abc_41356_new_n4061_), .B(_abc_41356_new_n4062_), .Y(_abc_41356_new_n4063_));
OR2X2 OR2X2_1263 ( .A(_abc_41356_new_n4063_), .B(_abc_41356_new_n4060_), .Y(_abc_41356_new_n4064_));
OR2X2 OR2X2_1264 ( .A(_abc_41356_new_n4059_), .B(_abc_41356_new_n4064_), .Y(_abc_41356_new_n4065_));
OR2X2 OR2X2_1265 ( .A(_abc_41356_new_n4066_), .B(_abc_41356_new_n4017_), .Y(_0wdatahold_7_0__6_));
OR2X2 OR2X2_1266 ( .A(_abc_41356_new_n4025_), .B(pc_7_), .Y(_abc_41356_new_n4069_));
OR2X2 OR2X2_1267 ( .A(_abc_41356_new_n4073_), .B(_abc_41356_new_n2073_), .Y(_abc_41356_new_n4074_));
OR2X2 OR2X2_1268 ( .A(_abc_41356_new_n4077_), .B(_abc_41356_new_n4079_), .Y(_abc_41356_new_n4080_));
OR2X2 OR2X2_1269 ( .A(_abc_41356_new_n534_), .B(regfil_3__7_), .Y(_abc_41356_new_n4081_));
OR2X2 OR2X2_127 ( .A(_abc_41356_new_n931_), .B(_abc_41356_new_n934_), .Y(_abc_41356_new_n935_));
OR2X2 OR2X2_1270 ( .A(_abc_41356_new_n4080_), .B(_abc_41356_new_n4082_), .Y(_abc_41356_new_n4083_));
OR2X2 OR2X2_1271 ( .A(_abc_41356_new_n3735_), .B(regfil_1__7_), .Y(_abc_41356_new_n4084_));
OR2X2 OR2X2_1272 ( .A(_abc_41356_new_n4086_), .B(_abc_41356_new_n4088_), .Y(_abc_41356_new_n4089_));
OR2X2 OR2X2_1273 ( .A(_abc_41356_new_n4089_), .B(_abc_41356_new_n4078_), .Y(_abc_41356_new_n4090_));
OR2X2 OR2X2_1274 ( .A(_abc_41356_new_n4076_), .B(_abc_41356_new_n4090_), .Y(_abc_41356_new_n4091_));
OR2X2 OR2X2_1275 ( .A(_abc_41356_new_n4091_), .B(_abc_41356_new_n4071_), .Y(_abc_41356_new_n4092_));
OR2X2 OR2X2_1276 ( .A(_abc_41356_new_n4094_), .B(_abc_41356_new_n4077_), .Y(_abc_41356_new_n4095_));
OR2X2 OR2X2_1277 ( .A(_abc_41356_new_n4095_), .B(_abc_41356_new_n3710_), .Y(_abc_41356_new_n4096_));
OR2X2 OR2X2_1278 ( .A(_abc_41356_new_n2026_), .B(wdatahold_7_), .Y(_abc_41356_new_n4097_));
OR2X2 OR2X2_1279 ( .A(_abc_41356_new_n1161_), .B(_abc_41356_new_n3475_), .Y(_abc_41356_new_n4100_));
OR2X2 OR2X2_128 ( .A(_abc_41356_new_n935_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n936_));
OR2X2 OR2X2_1280 ( .A(_abc_41356_new_n3411_), .B(wdatahold_7_), .Y(_abc_41356_new_n4101_));
OR2X2 OR2X2_1281 ( .A(_abc_41356_new_n4103_), .B(_abc_41356_new_n4099_), .Y(_abc_41356_new_n4104_));
OR2X2 OR2X2_1282 ( .A(_abc_41356_new_n4105_), .B(_abc_41356_new_n4104_), .Y(_abc_41356_new_n4106_));
OR2X2 OR2X2_1283 ( .A(_abc_41356_new_n4106_), .B(_abc_41356_new_n4093_), .Y(_abc_41356_new_n4107_));
OR2X2 OR2X2_1284 ( .A(_abc_41356_new_n4110_), .B(_abc_41356_new_n4111_), .Y(_abc_41356_new_n4112_));
OR2X2 OR2X2_1285 ( .A(_abc_41356_new_n4112_), .B(_abc_41356_new_n4109_), .Y(_abc_41356_new_n4113_));
OR2X2 OR2X2_1286 ( .A(_abc_41356_new_n4108_), .B(_abc_41356_new_n4113_), .Y(_abc_41356_new_n4114_));
OR2X2 OR2X2_1287 ( .A(_abc_41356_new_n4115_), .B(_abc_41356_new_n4068_), .Y(_0wdatahold_7_0__7_));
OR2X2 OR2X2_1288 ( .A(_abc_41356_new_n4121_), .B(reset), .Y(_abc_41356_new_n4122_));
OR2X2 OR2X2_1289 ( .A(_abc_41356_new_n3392_), .B(_abc_41356_new_n3361_), .Y(_abc_41356_new_n4124_));
OR2X2 OR2X2_129 ( .A(_abc_41356_new_n937_), .B(opcode_2_), .Y(_abc_41356_new_n938_));
OR2X2 OR2X2_1290 ( .A(_abc_41356_new_n4127_), .B(_abc_41356_new_n3373_), .Y(_abc_41356_new_n4128_));
OR2X2 OR2X2_1291 ( .A(_abc_41356_new_n682_), .B(raddrhold_0_), .Y(_abc_41356_new_n4134_));
OR2X2 OR2X2_1292 ( .A(opcode_4_), .B(regfil_1__0_), .Y(_abc_41356_new_n4137_));
OR2X2 OR2X2_1293 ( .A(_abc_41356_new_n4136_), .B(_abc_41356_new_n4139_), .Y(_abc_41356_new_n4140_));
OR2X2 OR2X2_1294 ( .A(_abc_41356_new_n4140_), .B(_abc_41356_new_n4135_), .Y(_abc_41356_new_n4141_));
OR2X2 OR2X2_1295 ( .A(_abc_41356_new_n4141_), .B(_abc_41356_new_n4130_), .Y(_abc_41356_new_n4142_));
OR2X2 OR2X2_1296 ( .A(_abc_41356_new_n4143_), .B(raddrhold_0_), .Y(_abc_41356_new_n4144_));
OR2X2 OR2X2_1297 ( .A(_abc_41356_new_n3355_), .B(_abc_41356_new_n4152_), .Y(_abc_41356_new_n4153_));
OR2X2 OR2X2_1298 ( .A(_abc_41356_new_n4153_), .B(_abc_41356_new_n4147_), .Y(_abc_41356_new_n4154_));
OR2X2 OR2X2_1299 ( .A(_abc_41356_new_n4176_), .B(_abc_41356_new_n4174_), .Y(_abc_41356_new_n4177_));
OR2X2 OR2X2_13 ( .A(_abc_41356_new_n626_), .B(opcode_2_), .Y(_abc_41356_new_n627_));
OR2X2 OR2X2_130 ( .A(_abc_41356_new_n940_), .B(_abc_41356_new_n941_), .Y(_abc_41356_new_n942_));
OR2X2 OR2X2_1300 ( .A(_abc_41356_new_n4177_), .B(_abc_41356_new_n4172_), .Y(_abc_41356_new_n4178_));
OR2X2 OR2X2_1301 ( .A(_abc_41356_new_n4181_), .B(_abc_41356_new_n4180_), .Y(_abc_41356_new_n4182_));
OR2X2 OR2X2_1302 ( .A(_abc_41356_new_n4188_), .B(_abc_41356_new_n4189_), .Y(_abc_41356_new_n4190_));
OR2X2 OR2X2_1303 ( .A(_abc_41356_new_n4190_), .B(_abc_41356_new_n4187_), .Y(_abc_41356_new_n4191_));
OR2X2 OR2X2_1304 ( .A(_abc_41356_new_n4179_), .B(_abc_41356_new_n4191_), .Y(_abc_41356_new_n4192_));
OR2X2 OR2X2_1305 ( .A(_abc_41356_new_n4192_), .B(_abc_41356_new_n4146_), .Y(_abc_41356_new_n4193_));
OR2X2 OR2X2_1306 ( .A(_abc_41356_new_n4195_), .B(_abc_41356_new_n4197_), .Y(_abc_41356_new_n4198_));
OR2X2 OR2X2_1307 ( .A(_abc_41356_new_n4194_), .B(_abc_41356_new_n4198_), .Y(_abc_41356_new_n4199_));
OR2X2 OR2X2_1308 ( .A(_abc_41356_new_n4200_), .B(_abc_41356_new_n4123_), .Y(_0raddrhold_15_0__0_));
OR2X2 OR2X2_1309 ( .A(_abc_41356_new_n682_), .B(raddrhold_1_), .Y(_abc_41356_new_n4204_));
OR2X2 OR2X2_131 ( .A(_abc_41356_new_n942_), .B(_abc_41356_new_n939_), .Y(_abc_41356_new_n943_));
OR2X2 OR2X2_1310 ( .A(_abc_41356_new_n3772_), .B(_abc_41356_new_n3774_), .Y(_abc_41356_new_n4208_));
OR2X2 OR2X2_1311 ( .A(_abc_41356_new_n4207_), .B(_abc_41356_new_n4209_), .Y(_abc_41356_new_n4210_));
OR2X2 OR2X2_1312 ( .A(_abc_41356_new_n4210_), .B(_abc_41356_new_n4206_), .Y(_abc_41356_new_n4211_));
OR2X2 OR2X2_1313 ( .A(_abc_41356_new_n4211_), .B(_abc_41356_new_n4130_), .Y(_abc_41356_new_n4212_));
OR2X2 OR2X2_1314 ( .A(_abc_41356_new_n4143_), .B(raddrhold_1_), .Y(_abc_41356_new_n4213_));
OR2X2 OR2X2_1315 ( .A(_abc_41356_new_n4217_), .B(_abc_41356_new_n4218_), .Y(_abc_41356_new_n4219_));
OR2X2 OR2X2_1316 ( .A(_abc_41356_new_n4219_), .B(_abc_41356_new_n4216_), .Y(_abc_41356_new_n4220_));
OR2X2 OR2X2_1317 ( .A(_abc_41356_new_n4223_), .B(_abc_41356_new_n4222_), .Y(_abc_41356_new_n4224_));
OR2X2 OR2X2_1318 ( .A(_abc_41356_new_n4226_), .B(_abc_41356_new_n4227_), .Y(_abc_41356_new_n4228_));
OR2X2 OR2X2_1319 ( .A(_abc_41356_new_n4228_), .B(_abc_41356_new_n4225_), .Y(_abc_41356_new_n4229_));
OR2X2 OR2X2_132 ( .A(_abc_41356_new_n943_), .B(_abc_41356_new_n938_), .Y(_abc_41356_new_n944_));
OR2X2 OR2X2_1320 ( .A(_abc_41356_new_n4221_), .B(_abc_41356_new_n4229_), .Y(_abc_41356_new_n4230_));
OR2X2 OR2X2_1321 ( .A(_abc_41356_new_n4230_), .B(_abc_41356_new_n4215_), .Y(_abc_41356_new_n4231_));
OR2X2 OR2X2_1322 ( .A(_abc_41356_new_n4232_), .B(_abc_41356_new_n4233_), .Y(_abc_41356_new_n4234_));
OR2X2 OR2X2_1323 ( .A(raddrhold_0_), .B(raddrhold_1_), .Y(_abc_41356_new_n4237_));
OR2X2 OR2X2_1324 ( .A(_abc_41356_new_n4236_), .B(_abc_41356_new_n4242_), .Y(_abc_41356_new_n4243_));
OR2X2 OR2X2_1325 ( .A(_abc_41356_new_n4235_), .B(_abc_41356_new_n4243_), .Y(_0raddrhold_15_0__1_));
OR2X2 OR2X2_1326 ( .A(_abc_41356_new_n682_), .B(raddrhold_2_), .Y(_abc_41356_new_n4248_));
OR2X2 OR2X2_1327 ( .A(opcode_4_), .B(regfil_1__2_), .Y(_abc_41356_new_n4251_));
OR2X2 OR2X2_1328 ( .A(_abc_41356_new_n4250_), .B(_abc_41356_new_n4253_), .Y(_abc_41356_new_n4254_));
OR2X2 OR2X2_1329 ( .A(_abc_41356_new_n4254_), .B(_abc_41356_new_n4249_), .Y(_abc_41356_new_n4255_));
OR2X2 OR2X2_133 ( .A(_abc_41356_new_n946_), .B(_abc_41356_new_n947_), .Y(_abc_41356_new_n948_));
OR2X2 OR2X2_1330 ( .A(_abc_41356_new_n4255_), .B(_abc_41356_new_n4130_), .Y(_abc_41356_new_n4256_));
OR2X2 OR2X2_1331 ( .A(_abc_41356_new_n4143_), .B(raddrhold_2_), .Y(_abc_41356_new_n4257_));
OR2X2 OR2X2_1332 ( .A(_abc_41356_new_n4261_), .B(_abc_41356_new_n4262_), .Y(_abc_41356_new_n4263_));
OR2X2 OR2X2_1333 ( .A(_abc_41356_new_n4263_), .B(_abc_41356_new_n4260_), .Y(_abc_41356_new_n4264_));
OR2X2 OR2X2_1334 ( .A(_abc_41356_new_n4267_), .B(_abc_41356_new_n4266_), .Y(_abc_41356_new_n4268_));
OR2X2 OR2X2_1335 ( .A(_abc_41356_new_n4270_), .B(_abc_41356_new_n4271_), .Y(_abc_41356_new_n4272_));
OR2X2 OR2X2_1336 ( .A(_abc_41356_new_n4272_), .B(_abc_41356_new_n4269_), .Y(_abc_41356_new_n4273_));
OR2X2 OR2X2_1337 ( .A(_abc_41356_new_n4265_), .B(_abc_41356_new_n4273_), .Y(_abc_41356_new_n4274_));
OR2X2 OR2X2_1338 ( .A(_abc_41356_new_n4274_), .B(_abc_41356_new_n4259_), .Y(_abc_41356_new_n4275_));
OR2X2 OR2X2_1339 ( .A(_abc_41356_new_n4276_), .B(_abc_41356_new_n4277_), .Y(_abc_41356_new_n4278_));
OR2X2 OR2X2_134 ( .A(_abc_41356_new_n949_), .B(_abc_41356_new_n928_), .Y(_abc_41356_new_n950_));
OR2X2 OR2X2_1340 ( .A(_abc_41356_new_n4238_), .B(raddrhold_2_), .Y(_abc_41356_new_n4281_));
OR2X2 OR2X2_1341 ( .A(_abc_41356_new_n4280_), .B(_abc_41356_new_n4285_), .Y(_abc_41356_new_n4286_));
OR2X2 OR2X2_1342 ( .A(_abc_41356_new_n4279_), .B(_abc_41356_new_n4286_), .Y(_0raddrhold_15_0__2_));
OR2X2 OR2X2_1343 ( .A(_abc_41356_new_n682_), .B(raddrhold_3_), .Y(_abc_41356_new_n4292_));
OR2X2 OR2X2_1344 ( .A(opcode_4_), .B(regfil_1__3_), .Y(_abc_41356_new_n4295_));
OR2X2 OR2X2_1345 ( .A(_abc_41356_new_n4294_), .B(_abc_41356_new_n4297_), .Y(_abc_41356_new_n4298_));
OR2X2 OR2X2_1346 ( .A(_abc_41356_new_n4298_), .B(_abc_41356_new_n4293_), .Y(_abc_41356_new_n4299_));
OR2X2 OR2X2_1347 ( .A(_abc_41356_new_n4299_), .B(_abc_41356_new_n4130_), .Y(_abc_41356_new_n4300_));
OR2X2 OR2X2_1348 ( .A(_abc_41356_new_n4143_), .B(raddrhold_3_), .Y(_abc_41356_new_n4301_));
OR2X2 OR2X2_1349 ( .A(_abc_41356_new_n4305_), .B(_abc_41356_new_n4306_), .Y(_abc_41356_new_n4307_));
OR2X2 OR2X2_135 ( .A(_abc_41356_new_n927_), .B(_abc_41356_new_n950_), .Y(_abc_41356_new_n951_));
OR2X2 OR2X2_1350 ( .A(_abc_41356_new_n4307_), .B(_abc_41356_new_n4304_), .Y(_abc_41356_new_n4308_));
OR2X2 OR2X2_1351 ( .A(_abc_41356_new_n4311_), .B(_abc_41356_new_n4310_), .Y(_abc_41356_new_n4312_));
OR2X2 OR2X2_1352 ( .A(_abc_41356_new_n4314_), .B(_abc_41356_new_n4315_), .Y(_abc_41356_new_n4316_));
OR2X2 OR2X2_1353 ( .A(_abc_41356_new_n4316_), .B(_abc_41356_new_n4313_), .Y(_abc_41356_new_n4317_));
OR2X2 OR2X2_1354 ( .A(_abc_41356_new_n4309_), .B(_abc_41356_new_n4317_), .Y(_abc_41356_new_n4318_));
OR2X2 OR2X2_1355 ( .A(_abc_41356_new_n4318_), .B(_abc_41356_new_n4303_), .Y(_abc_41356_new_n4319_));
OR2X2 OR2X2_1356 ( .A(_abc_41356_new_n4282_), .B(raddrhold_3_), .Y(_abc_41356_new_n4323_));
OR2X2 OR2X2_1357 ( .A(_abc_41356_new_n4325_), .B(_abc_41356_new_n4326_), .Y(_abc_41356_new_n4327_));
OR2X2 OR2X2_1358 ( .A(_abc_41356_new_n4320_), .B(_abc_41356_new_n4327_), .Y(_abc_41356_new_n4328_));
OR2X2 OR2X2_1359 ( .A(_abc_41356_new_n4329_), .B(_abc_41356_new_n4288_), .Y(_0raddrhold_15_0__3_));
OR2X2 OR2X2_136 ( .A(_abc_41356_new_n922_), .B(_abc_41356_new_n951_), .Y(_abc_41356_new_n952_));
OR2X2 OR2X2_1360 ( .A(_abc_41356_new_n682_), .B(raddrhold_4_), .Y(_abc_41356_new_n4335_));
OR2X2 OR2X2_1361 ( .A(opcode_4_), .B(regfil_1__4_), .Y(_abc_41356_new_n4338_));
OR2X2 OR2X2_1362 ( .A(_abc_41356_new_n4337_), .B(_abc_41356_new_n4340_), .Y(_abc_41356_new_n4341_));
OR2X2 OR2X2_1363 ( .A(_abc_41356_new_n4341_), .B(_abc_41356_new_n4336_), .Y(_abc_41356_new_n4342_));
OR2X2 OR2X2_1364 ( .A(_abc_41356_new_n4342_), .B(_abc_41356_new_n4130_), .Y(_abc_41356_new_n4343_));
OR2X2 OR2X2_1365 ( .A(_abc_41356_new_n4143_), .B(raddrhold_4_), .Y(_abc_41356_new_n4344_));
OR2X2 OR2X2_1366 ( .A(_abc_41356_new_n4348_), .B(_abc_41356_new_n4349_), .Y(_abc_41356_new_n4350_));
OR2X2 OR2X2_1367 ( .A(_abc_41356_new_n4350_), .B(_abc_41356_new_n4347_), .Y(_abc_41356_new_n4351_));
OR2X2 OR2X2_1368 ( .A(_abc_41356_new_n4354_), .B(_abc_41356_new_n4353_), .Y(_abc_41356_new_n4355_));
OR2X2 OR2X2_1369 ( .A(_abc_41356_new_n4357_), .B(_abc_41356_new_n4358_), .Y(_abc_41356_new_n4359_));
OR2X2 OR2X2_137 ( .A(_abc_41356_new_n952_), .B(_abc_41356_new_n696_), .Y(_abc_41356_new_n953_));
OR2X2 OR2X2_1370 ( .A(_abc_41356_new_n4359_), .B(_abc_41356_new_n4356_), .Y(_abc_41356_new_n4360_));
OR2X2 OR2X2_1371 ( .A(_abc_41356_new_n4352_), .B(_abc_41356_new_n4360_), .Y(_abc_41356_new_n4361_));
OR2X2 OR2X2_1372 ( .A(_abc_41356_new_n4361_), .B(_abc_41356_new_n4346_), .Y(_abc_41356_new_n4362_));
OR2X2 OR2X2_1373 ( .A(_abc_41356_new_n4321_), .B(raddrhold_4_), .Y(_abc_41356_new_n4366_));
OR2X2 OR2X2_1374 ( .A(_abc_41356_new_n4368_), .B(_abc_41356_new_n4369_), .Y(_abc_41356_new_n4370_));
OR2X2 OR2X2_1375 ( .A(_abc_41356_new_n4363_), .B(_abc_41356_new_n4370_), .Y(_abc_41356_new_n4371_));
OR2X2 OR2X2_1376 ( .A(_abc_41356_new_n4372_), .B(_abc_41356_new_n4331_), .Y(_0raddrhold_15_0__4_));
OR2X2 OR2X2_1377 ( .A(_abc_41356_new_n682_), .B(raddrhold_5_), .Y(_abc_41356_new_n4378_));
OR2X2 OR2X2_1378 ( .A(opcode_4_), .B(regfil_1__5_), .Y(_abc_41356_new_n4381_));
OR2X2 OR2X2_1379 ( .A(_abc_41356_new_n4380_), .B(_abc_41356_new_n4383_), .Y(_abc_41356_new_n4384_));
OR2X2 OR2X2_138 ( .A(_abc_41356_new_n695_), .B(regfil_7__4_), .Y(_abc_41356_new_n954_));
OR2X2 OR2X2_1380 ( .A(_abc_41356_new_n4384_), .B(_abc_41356_new_n4379_), .Y(_abc_41356_new_n4385_));
OR2X2 OR2X2_1381 ( .A(_abc_41356_new_n4385_), .B(_abc_41356_new_n4130_), .Y(_abc_41356_new_n4386_));
OR2X2 OR2X2_1382 ( .A(_abc_41356_new_n4143_), .B(raddrhold_5_), .Y(_abc_41356_new_n4387_));
OR2X2 OR2X2_1383 ( .A(_abc_41356_new_n4391_), .B(_abc_41356_new_n4392_), .Y(_abc_41356_new_n4393_));
OR2X2 OR2X2_1384 ( .A(_abc_41356_new_n4393_), .B(_abc_41356_new_n4390_), .Y(_abc_41356_new_n4394_));
OR2X2 OR2X2_1385 ( .A(_abc_41356_new_n4397_), .B(_abc_41356_new_n4396_), .Y(_abc_41356_new_n4398_));
OR2X2 OR2X2_1386 ( .A(_abc_41356_new_n4400_), .B(_abc_41356_new_n4401_), .Y(_abc_41356_new_n4402_));
OR2X2 OR2X2_1387 ( .A(_abc_41356_new_n4402_), .B(_abc_41356_new_n4399_), .Y(_abc_41356_new_n4403_));
OR2X2 OR2X2_1388 ( .A(_abc_41356_new_n4395_), .B(_abc_41356_new_n4403_), .Y(_abc_41356_new_n4404_));
OR2X2 OR2X2_1389 ( .A(_abc_41356_new_n4404_), .B(_abc_41356_new_n4389_), .Y(_abc_41356_new_n4405_));
OR2X2 OR2X2_139 ( .A(_abc_41356_new_n899_), .B(regfil_7__4_), .Y(_abc_41356_new_n960_));
OR2X2 OR2X2_1390 ( .A(_abc_41356_new_n4364_), .B(raddrhold_5_), .Y(_abc_41356_new_n4409_));
OR2X2 OR2X2_1391 ( .A(_abc_41356_new_n4411_), .B(_abc_41356_new_n4412_), .Y(_abc_41356_new_n4413_));
OR2X2 OR2X2_1392 ( .A(_abc_41356_new_n4406_), .B(_abc_41356_new_n4413_), .Y(_abc_41356_new_n4414_));
OR2X2 OR2X2_1393 ( .A(_abc_41356_new_n4415_), .B(_abc_41356_new_n4374_), .Y(_0raddrhold_15_0__5_));
OR2X2 OR2X2_1394 ( .A(_abc_41356_new_n4130_), .B(_abc_41356_new_n4420_), .Y(_abc_41356_new_n4421_));
OR2X2 OR2X2_1395 ( .A(opcode_4_), .B(regfil_1__6_), .Y(_abc_41356_new_n4424_));
OR2X2 OR2X2_1396 ( .A(_abc_41356_new_n4427_), .B(_abc_41356_new_n4426_), .Y(_abc_41356_new_n4428_));
OR2X2 OR2X2_1397 ( .A(_abc_41356_new_n4423_), .B(_abc_41356_new_n4428_), .Y(_abc_41356_new_n4429_));
OR2X2 OR2X2_1398 ( .A(_abc_41356_new_n4422_), .B(_abc_41356_new_n4429_), .Y(_abc_41356_new_n4430_));
OR2X2 OR2X2_1399 ( .A(_abc_41356_new_n4433_), .B(_abc_41356_new_n4434_), .Y(_abc_41356_new_n4435_));
OR2X2 OR2X2_14 ( .A(_abc_41356_new_n628_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n629_));
OR2X2 OR2X2_140 ( .A(_abc_41356_new_n960_), .B(_abc_41356_new_n959_), .Y(_abc_41356_new_n961_));
OR2X2 OR2X2_1400 ( .A(_abc_41356_new_n4435_), .B(_abc_41356_new_n4432_), .Y(_abc_41356_new_n4436_));
OR2X2 OR2X2_1401 ( .A(_abc_41356_new_n4439_), .B(_abc_41356_new_n4438_), .Y(_abc_41356_new_n4440_));
OR2X2 OR2X2_1402 ( .A(_abc_41356_new_n4442_), .B(_abc_41356_new_n4443_), .Y(_abc_41356_new_n4444_));
OR2X2 OR2X2_1403 ( .A(_abc_41356_new_n4444_), .B(_abc_41356_new_n4441_), .Y(_abc_41356_new_n4445_));
OR2X2 OR2X2_1404 ( .A(_abc_41356_new_n4437_), .B(_abc_41356_new_n4445_), .Y(_abc_41356_new_n4446_));
OR2X2 OR2X2_1405 ( .A(_abc_41356_new_n4446_), .B(_abc_41356_new_n4431_), .Y(_abc_41356_new_n4447_));
OR2X2 OR2X2_1406 ( .A(_abc_41356_new_n4407_), .B(raddrhold_6_), .Y(_abc_41356_new_n4451_));
OR2X2 OR2X2_1407 ( .A(_abc_41356_new_n4453_), .B(_abc_41356_new_n4454_), .Y(_abc_41356_new_n4455_));
OR2X2 OR2X2_1408 ( .A(_abc_41356_new_n4448_), .B(_abc_41356_new_n4455_), .Y(_abc_41356_new_n4456_));
OR2X2 OR2X2_1409 ( .A(_abc_41356_new_n4457_), .B(_abc_41356_new_n4417_), .Y(_0raddrhold_15_0__6_));
OR2X2 OR2X2_141 ( .A(_abc_41356_new_n699_), .B(_abc_41356_new_n893_), .Y(_abc_41356_new_n966_));
OR2X2 OR2X2_1410 ( .A(_abc_41356_new_n682_), .B(raddrhold_7_), .Y(_abc_41356_new_n4463_));
OR2X2 OR2X2_1411 ( .A(opcode_4_), .B(regfil_1__7_), .Y(_abc_41356_new_n4466_));
OR2X2 OR2X2_1412 ( .A(_abc_41356_new_n4465_), .B(_abc_41356_new_n4468_), .Y(_abc_41356_new_n4469_));
OR2X2 OR2X2_1413 ( .A(_abc_41356_new_n4469_), .B(_abc_41356_new_n4464_), .Y(_abc_41356_new_n4470_));
OR2X2 OR2X2_1414 ( .A(_abc_41356_new_n4470_), .B(_abc_41356_new_n4130_), .Y(_abc_41356_new_n4471_));
OR2X2 OR2X2_1415 ( .A(_abc_41356_new_n4143_), .B(raddrhold_7_), .Y(_abc_41356_new_n4472_));
OR2X2 OR2X2_1416 ( .A(_abc_41356_new_n4476_), .B(_abc_41356_new_n4477_), .Y(_abc_41356_new_n4478_));
OR2X2 OR2X2_1417 ( .A(_abc_41356_new_n4478_), .B(_abc_41356_new_n4475_), .Y(_abc_41356_new_n4479_));
OR2X2 OR2X2_1418 ( .A(_abc_41356_new_n4482_), .B(_abc_41356_new_n4481_), .Y(_abc_41356_new_n4483_));
OR2X2 OR2X2_1419 ( .A(_abc_41356_new_n4485_), .B(_abc_41356_new_n4486_), .Y(_abc_41356_new_n4487_));
OR2X2 OR2X2_142 ( .A(_abc_41356_new_n965_), .B(_abc_41356_new_n966_), .Y(_abc_41356_new_n967_));
OR2X2 OR2X2_1420 ( .A(_abc_41356_new_n4487_), .B(_abc_41356_new_n4484_), .Y(_abc_41356_new_n4488_));
OR2X2 OR2X2_1421 ( .A(_abc_41356_new_n4480_), .B(_abc_41356_new_n4488_), .Y(_abc_41356_new_n4489_));
OR2X2 OR2X2_1422 ( .A(_abc_41356_new_n4489_), .B(_abc_41356_new_n4474_), .Y(_abc_41356_new_n4490_));
OR2X2 OR2X2_1423 ( .A(_abc_41356_new_n4449_), .B(raddrhold_7_), .Y(_abc_41356_new_n4494_));
OR2X2 OR2X2_1424 ( .A(_abc_41356_new_n4496_), .B(_abc_41356_new_n4497_), .Y(_abc_41356_new_n4498_));
OR2X2 OR2X2_1425 ( .A(_abc_41356_new_n4491_), .B(_abc_41356_new_n4498_), .Y(_abc_41356_new_n4499_));
OR2X2 OR2X2_1426 ( .A(_abc_41356_new_n4500_), .B(_abc_41356_new_n4459_), .Y(_0raddrhold_15_0__7_));
OR2X2 OR2X2_1427 ( .A(_abc_41356_new_n682_), .B(raddrhold_8_), .Y(_abc_41356_new_n4506_));
OR2X2 OR2X2_1428 ( .A(_abc_41356_new_n4508_), .B(_abc_41356_new_n4509_), .Y(_abc_41356_new_n4510_));
OR2X2 OR2X2_1429 ( .A(_abc_41356_new_n4510_), .B(_abc_41356_new_n4507_), .Y(_abc_41356_new_n4511_));
OR2X2 OR2X2_143 ( .A(_abc_41356_new_n975_), .B(_abc_41356_new_n974_), .Y(_abc_41356_new_n976_));
OR2X2 OR2X2_1430 ( .A(_abc_41356_new_n4511_), .B(_abc_41356_new_n4130_), .Y(_abc_41356_new_n4512_));
OR2X2 OR2X2_1431 ( .A(_abc_41356_new_n4143_), .B(raddrhold_8_), .Y(_abc_41356_new_n4513_));
OR2X2 OR2X2_1432 ( .A(_abc_41356_new_n4517_), .B(_abc_41356_new_n4518_), .Y(_abc_41356_new_n4519_));
OR2X2 OR2X2_1433 ( .A(_abc_41356_new_n4519_), .B(_abc_41356_new_n4516_), .Y(_abc_41356_new_n4520_));
OR2X2 OR2X2_1434 ( .A(_abc_41356_new_n4523_), .B(_abc_41356_new_n4522_), .Y(_abc_41356_new_n4524_));
OR2X2 OR2X2_1435 ( .A(_abc_41356_new_n4526_), .B(_abc_41356_new_n4527_), .Y(_abc_41356_new_n4528_));
OR2X2 OR2X2_1436 ( .A(_abc_41356_new_n4528_), .B(_abc_41356_new_n4525_), .Y(_abc_41356_new_n4529_));
OR2X2 OR2X2_1437 ( .A(_abc_41356_new_n4521_), .B(_abc_41356_new_n4529_), .Y(_abc_41356_new_n4530_));
OR2X2 OR2X2_1438 ( .A(_abc_41356_new_n4530_), .B(_abc_41356_new_n4515_), .Y(_abc_41356_new_n4531_));
OR2X2 OR2X2_1439 ( .A(_abc_41356_new_n4492_), .B(raddrhold_8_), .Y(_abc_41356_new_n4535_));
OR2X2 OR2X2_144 ( .A(_abc_41356_new_n956_), .B(_abc_41356_new_n983_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_4_));
OR2X2 OR2X2_1440 ( .A(_abc_41356_new_n4537_), .B(_abc_41356_new_n4538_), .Y(_abc_41356_new_n4539_));
OR2X2 OR2X2_1441 ( .A(_abc_41356_new_n4532_), .B(_abc_41356_new_n4539_), .Y(_abc_41356_new_n4540_));
OR2X2 OR2X2_1442 ( .A(_abc_41356_new_n4541_), .B(_abc_41356_new_n4502_), .Y(_0raddrhold_15_0__8_));
OR2X2 OR2X2_1443 ( .A(_abc_41356_new_n682_), .B(raddrhold_9_), .Y(_abc_41356_new_n4547_));
OR2X2 OR2X2_1444 ( .A(_abc_41356_new_n4549_), .B(_abc_41356_new_n4550_), .Y(_abc_41356_new_n4551_));
OR2X2 OR2X2_1445 ( .A(_abc_41356_new_n4551_), .B(_abc_41356_new_n4548_), .Y(_abc_41356_new_n4552_));
OR2X2 OR2X2_1446 ( .A(_abc_41356_new_n4552_), .B(_abc_41356_new_n4130_), .Y(_abc_41356_new_n4553_));
OR2X2 OR2X2_1447 ( .A(_abc_41356_new_n4143_), .B(raddrhold_9_), .Y(_abc_41356_new_n4554_));
OR2X2 OR2X2_1448 ( .A(_abc_41356_new_n4558_), .B(_abc_41356_new_n4559_), .Y(_abc_41356_new_n4560_));
OR2X2 OR2X2_1449 ( .A(_abc_41356_new_n4560_), .B(_abc_41356_new_n4557_), .Y(_abc_41356_new_n4561_));
OR2X2 OR2X2_145 ( .A(_abc_41356_new_n918_), .B(regfil_0__5_), .Y(_abc_41356_new_n985_));
OR2X2 OR2X2_1450 ( .A(_abc_41356_new_n4564_), .B(_abc_41356_new_n4563_), .Y(_abc_41356_new_n4565_));
OR2X2 OR2X2_1451 ( .A(_abc_41356_new_n4567_), .B(_abc_41356_new_n4568_), .Y(_abc_41356_new_n4569_));
OR2X2 OR2X2_1452 ( .A(_abc_41356_new_n4569_), .B(_abc_41356_new_n4566_), .Y(_abc_41356_new_n4570_));
OR2X2 OR2X2_1453 ( .A(_abc_41356_new_n4562_), .B(_abc_41356_new_n4570_), .Y(_abc_41356_new_n4571_));
OR2X2 OR2X2_1454 ( .A(_abc_41356_new_n4571_), .B(_abc_41356_new_n4556_), .Y(_abc_41356_new_n4572_));
OR2X2 OR2X2_1455 ( .A(_abc_41356_new_n4533_), .B(raddrhold_9_), .Y(_abc_41356_new_n4576_));
OR2X2 OR2X2_1456 ( .A(_abc_41356_new_n4578_), .B(_abc_41356_new_n4579_), .Y(_abc_41356_new_n4580_));
OR2X2 OR2X2_1457 ( .A(_abc_41356_new_n4573_), .B(_abc_41356_new_n4580_), .Y(_abc_41356_new_n4581_));
OR2X2 OR2X2_1458 ( .A(_abc_41356_new_n4582_), .B(_abc_41356_new_n4543_), .Y(_0raddrhold_15_0__9_));
OR2X2 OR2X2_1459 ( .A(_abc_41356_new_n4586_), .B(_abc_41356_new_n4587_), .Y(_abc_41356_new_n4588_));
OR2X2 OR2X2_146 ( .A(_abc_41356_new_n986_), .B(_abc_41356_new_n987_), .Y(_abc_41356_new_n988_));
OR2X2 OR2X2_1460 ( .A(_abc_41356_new_n4588_), .B(_abc_41356_new_n4585_), .Y(_abc_41356_new_n4589_));
OR2X2 OR2X2_1461 ( .A(_abc_41356_new_n682_), .B(raddrhold_10_), .Y(_abc_41356_new_n4594_));
OR2X2 OR2X2_1462 ( .A(_abc_41356_new_n4596_), .B(_abc_41356_new_n4597_), .Y(_abc_41356_new_n4598_));
OR2X2 OR2X2_1463 ( .A(_abc_41356_new_n4130_), .B(_abc_41356_new_n4598_), .Y(_abc_41356_new_n4599_));
OR2X2 OR2X2_1464 ( .A(_abc_41356_new_n4599_), .B(_abc_41356_new_n4591_), .Y(_abc_41356_new_n4600_));
OR2X2 OR2X2_1465 ( .A(_abc_41356_new_n4143_), .B(raddrhold_10_), .Y(_abc_41356_new_n4601_));
OR2X2 OR2X2_1466 ( .A(_abc_41356_new_n4605_), .B(_abc_41356_new_n4604_), .Y(_abc_41356_new_n4606_));
OR2X2 OR2X2_1467 ( .A(_abc_41356_new_n4608_), .B(_abc_41356_new_n4609_), .Y(_abc_41356_new_n4610_));
OR2X2 OR2X2_1468 ( .A(_abc_41356_new_n4610_), .B(_abc_41356_new_n4607_), .Y(_abc_41356_new_n4611_));
OR2X2 OR2X2_1469 ( .A(_abc_41356_new_n4603_), .B(_abc_41356_new_n4611_), .Y(_abc_41356_new_n4612_));
OR2X2 OR2X2_147 ( .A(_abc_41356_new_n924_), .B(regfil_0__5_), .Y(_abc_41356_new_n990_));
OR2X2 OR2X2_1470 ( .A(_abc_41356_new_n4612_), .B(_abc_41356_new_n4590_), .Y(_abc_41356_new_n4613_));
OR2X2 OR2X2_1471 ( .A(_abc_41356_new_n4574_), .B(raddrhold_10_), .Y(_abc_41356_new_n4616_));
OR2X2 OR2X2_1472 ( .A(_abc_41356_new_n4620_), .B(_abc_41356_new_n4615_), .Y(_abc_41356_new_n4621_));
OR2X2 OR2X2_1473 ( .A(_abc_41356_new_n4614_), .B(_abc_41356_new_n4621_), .Y(_abc_41356_new_n4622_));
OR2X2 OR2X2_1474 ( .A(_abc_41356_new_n4623_), .B(_abc_41356_new_n4584_), .Y(_0raddrhold_15_0__10_));
OR2X2 OR2X2_1475 ( .A(_abc_41356_new_n682_), .B(raddrhold_11_), .Y(_abc_41356_new_n4629_));
OR2X2 OR2X2_1476 ( .A(_abc_41356_new_n4631_), .B(_abc_41356_new_n4632_), .Y(_abc_41356_new_n4633_));
OR2X2 OR2X2_1477 ( .A(_abc_41356_new_n4626_), .B(_abc_41356_new_n4633_), .Y(_abc_41356_new_n4634_));
OR2X2 OR2X2_1478 ( .A(_abc_41356_new_n4638_), .B(_abc_41356_new_n4637_), .Y(_abc_41356_new_n4639_));
OR2X2 OR2X2_1479 ( .A(_abc_41356_new_n4186_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4640_));
OR2X2 OR2X2_148 ( .A(_abc_41356_new_n996_), .B(_abc_41356_new_n997_), .Y(_abc_41356_new_n998_));
OR2X2 OR2X2_1480 ( .A(_abc_41356_new_n4636_), .B(_abc_41356_new_n4641_), .Y(_abc_41356_new_n4642_));
OR2X2 OR2X2_1481 ( .A(_abc_41356_new_n4643_), .B(_abc_41356_new_n4644_), .Y(_abc_41356_new_n4645_));
OR2X2 OR2X2_1482 ( .A(_abc_41356_new_n4648_), .B(_abc_41356_new_n4184_), .Y(_abc_41356_new_n4649_));
OR2X2 OR2X2_1483 ( .A(_abc_41356_new_n4649_), .B(_abc_41356_new_n4647_), .Y(_abc_41356_new_n4650_));
OR2X2 OR2X2_1484 ( .A(_abc_41356_new_n4651_), .B(_abc_41356_new_n4646_), .Y(_abc_41356_new_n4652_));
OR2X2 OR2X2_1485 ( .A(_abc_41356_new_n4652_), .B(_abc_41356_new_n4642_), .Y(_abc_41356_new_n4653_));
OR2X2 OR2X2_1486 ( .A(_abc_41356_new_n4617_), .B(raddrhold_11_), .Y(_abc_41356_new_n4656_));
OR2X2 OR2X2_1487 ( .A(_abc_41356_new_n4660_), .B(_abc_41356_new_n4655_), .Y(_abc_41356_new_n4661_));
OR2X2 OR2X2_1488 ( .A(_abc_41356_new_n4654_), .B(_abc_41356_new_n4661_), .Y(_abc_41356_new_n4662_));
OR2X2 OR2X2_1489 ( .A(_abc_41356_new_n4663_), .B(_abc_41356_new_n4625_), .Y(_0raddrhold_15_0__11_));
OR2X2 OR2X2_149 ( .A(_abc_41356_new_n1000_), .B(_abc_41356_new_n999_), .Y(_abc_41356_new_n1001_));
OR2X2 OR2X2_1490 ( .A(_abc_41356_new_n682_), .B(raddrhold_12_), .Y(_abc_41356_new_n4669_));
OR2X2 OR2X2_1491 ( .A(_abc_41356_new_n4671_), .B(_abc_41356_new_n4672_), .Y(_abc_41356_new_n4673_));
OR2X2 OR2X2_1492 ( .A(_abc_41356_new_n4666_), .B(_abc_41356_new_n4673_), .Y(_abc_41356_new_n4674_));
OR2X2 OR2X2_1493 ( .A(_abc_41356_new_n4674_), .B(_abc_41356_new_n4675_), .Y(_abc_41356_new_n4676_));
OR2X2 OR2X2_1494 ( .A(_abc_41356_new_n4679_), .B(_abc_41356_new_n4678_), .Y(_abc_41356_new_n4680_));
OR2X2 OR2X2_1495 ( .A(_abc_41356_new_n4683_), .B(_abc_41356_new_n4682_), .Y(_abc_41356_new_n4684_));
OR2X2 OR2X2_1496 ( .A(_abc_41356_new_n4647_), .B(_abc_41356_new_n4184_), .Y(_abc_41356_new_n4686_));
OR2X2 OR2X2_1497 ( .A(_abc_41356_new_n4687_), .B(_abc_41356_new_n4685_), .Y(_abc_41356_new_n4688_));
OR2X2 OR2X2_1498 ( .A(_abc_41356_new_n4688_), .B(_abc_41356_new_n4681_), .Y(_abc_41356_new_n4689_));
OR2X2 OR2X2_1499 ( .A(_abc_41356_new_n4689_), .B(_abc_41356_new_n4677_), .Y(_abc_41356_new_n4690_));
OR2X2 OR2X2_15 ( .A(_abc_41356_new_n631_), .B(_abc_41356_new_n632_), .Y(_abc_41356_new_n633_));
OR2X2 OR2X2_150 ( .A(_abc_41356_new_n998_), .B(_abc_41356_new_n1001_), .Y(_abc_41356_new_n1002_));
OR2X2 OR2X2_1500 ( .A(_abc_41356_new_n4657_), .B(raddrhold_12_), .Y(_abc_41356_new_n4694_));
OR2X2 OR2X2_1501 ( .A(_abc_41356_new_n4696_), .B(_abc_41356_new_n4697_), .Y(_abc_41356_new_n4698_));
OR2X2 OR2X2_1502 ( .A(_abc_41356_new_n4691_), .B(_abc_41356_new_n4698_), .Y(_abc_41356_new_n4699_));
OR2X2 OR2X2_1503 ( .A(_abc_41356_new_n4700_), .B(_abc_41356_new_n4665_), .Y(_0raddrhold_15_0__12_));
OR2X2 OR2X2_1504 ( .A(_abc_41356_new_n682_), .B(raddrhold_13_), .Y(_abc_41356_new_n4706_));
OR2X2 OR2X2_1505 ( .A(_abc_41356_new_n4708_), .B(_abc_41356_new_n4709_), .Y(_abc_41356_new_n4710_));
OR2X2 OR2X2_1506 ( .A(_abc_41356_new_n4703_), .B(_abc_41356_new_n4710_), .Y(_abc_41356_new_n4711_));
OR2X2 OR2X2_1507 ( .A(_abc_41356_new_n4713_), .B(_abc_41356_new_n4714_), .Y(_abc_41356_new_n4715_));
OR2X2 OR2X2_1508 ( .A(_abc_41356_new_n4647_), .B(_abc_41356_new_n4648_), .Y(_abc_41356_new_n4717_));
OR2X2 OR2X2_1509 ( .A(_abc_41356_new_n4721_), .B(_abc_41356_new_n4720_), .Y(_abc_41356_new_n4722_));
OR2X2 OR2X2_151 ( .A(_abc_41356_new_n1002_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n1003_));
OR2X2 OR2X2_1510 ( .A(_abc_41356_new_n4723_), .B(_abc_41356_new_n4719_), .Y(_abc_41356_new_n4724_));
OR2X2 OR2X2_1511 ( .A(_abc_41356_new_n4718_), .B(_abc_41356_new_n4724_), .Y(_abc_41356_new_n4725_));
OR2X2 OR2X2_1512 ( .A(_abc_41356_new_n4725_), .B(_abc_41356_new_n4716_), .Y(_abc_41356_new_n4726_));
OR2X2 OR2X2_1513 ( .A(_abc_41356_new_n4726_), .B(_abc_41356_new_n4712_), .Y(_abc_41356_new_n4727_));
OR2X2 OR2X2_1514 ( .A(_abc_41356_new_n4692_), .B(raddrhold_13_), .Y(_abc_41356_new_n4730_));
OR2X2 OR2X2_1515 ( .A(_abc_41356_new_n4734_), .B(_abc_41356_new_n4729_), .Y(_abc_41356_new_n4735_));
OR2X2 OR2X2_1516 ( .A(_abc_41356_new_n4728_), .B(_abc_41356_new_n4735_), .Y(_abc_41356_new_n4736_));
OR2X2 OR2X2_1517 ( .A(_abc_41356_new_n4737_), .B(_abc_41356_new_n4702_), .Y(_0raddrhold_15_0__13_));
OR2X2 OR2X2_1518 ( .A(_abc_41356_new_n682_), .B(raddrhold_14_), .Y(_abc_41356_new_n4743_));
OR2X2 OR2X2_1519 ( .A(_abc_41356_new_n4745_), .B(_abc_41356_new_n4746_), .Y(_abc_41356_new_n4747_));
OR2X2 OR2X2_152 ( .A(_abc_41356_new_n1004_), .B(_abc_41356_new_n1005_), .Y(_abc_41356_new_n1006_));
OR2X2 OR2X2_1520 ( .A(_abc_41356_new_n4130_), .B(_abc_41356_new_n4747_), .Y(_abc_41356_new_n4748_));
OR2X2 OR2X2_1521 ( .A(_abc_41356_new_n4740_), .B(_abc_41356_new_n4748_), .Y(_abc_41356_new_n4749_));
OR2X2 OR2X2_1522 ( .A(_abc_41356_new_n4143_), .B(raddrhold_14_), .Y(_abc_41356_new_n4750_));
OR2X2 OR2X2_1523 ( .A(_abc_41356_new_n4754_), .B(_abc_41356_new_n4755_), .Y(_abc_41356_new_n4756_));
OR2X2 OR2X2_1524 ( .A(_abc_41356_new_n4756_), .B(_abc_41356_new_n4753_), .Y(_abc_41356_new_n4757_));
OR2X2 OR2X2_1525 ( .A(_abc_41356_new_n4761_), .B(_abc_41356_new_n4760_), .Y(_abc_41356_new_n4762_));
OR2X2 OR2X2_1526 ( .A(_abc_41356_new_n4763_), .B(_abc_41356_new_n4759_), .Y(_abc_41356_new_n4764_));
OR2X2 OR2X2_1527 ( .A(_abc_41356_new_n4758_), .B(_abc_41356_new_n4764_), .Y(_abc_41356_new_n4765_));
OR2X2 OR2X2_1528 ( .A(_abc_41356_new_n4765_), .B(_abc_41356_new_n4752_), .Y(_abc_41356_new_n4766_));
OR2X2 OR2X2_1529 ( .A(_abc_41356_new_n4731_), .B(raddrhold_14_), .Y(_abc_41356_new_n4771_));
OR2X2 OR2X2_153 ( .A(_abc_41356_new_n1008_), .B(_abc_41356_new_n1007_), .Y(_abc_41356_new_n1009_));
OR2X2 OR2X2_1530 ( .A(_abc_41356_new_n4773_), .B(_abc_41356_new_n4768_), .Y(_abc_41356_new_n4774_));
OR2X2 OR2X2_1531 ( .A(_abc_41356_new_n4767_), .B(_abc_41356_new_n4774_), .Y(_abc_41356_new_n4775_));
OR2X2 OR2X2_1532 ( .A(_abc_41356_new_n4776_), .B(_abc_41356_new_n4739_), .Y(_0raddrhold_15_0__14_));
OR2X2 OR2X2_1533 ( .A(_abc_41356_new_n682_), .B(raddrhold_15_), .Y(_abc_41356_new_n4780_));
OR2X2 OR2X2_1534 ( .A(_abc_41356_new_n4784_), .B(_abc_41356_new_n4785_), .Y(_abc_41356_new_n4786_));
OR2X2 OR2X2_1535 ( .A(_abc_41356_new_n4130_), .B(_abc_41356_new_n4786_), .Y(_abc_41356_new_n4787_));
OR2X2 OR2X2_1536 ( .A(_abc_41356_new_n4779_), .B(_abc_41356_new_n4787_), .Y(_abc_41356_new_n4788_));
OR2X2 OR2X2_1537 ( .A(_abc_41356_new_n4143_), .B(raddrhold_15_), .Y(_abc_41356_new_n4789_));
OR2X2 OR2X2_1538 ( .A(_abc_41356_new_n4793_), .B(_abc_41356_new_n4794_), .Y(_abc_41356_new_n4795_));
OR2X2 OR2X2_1539 ( .A(_abc_41356_new_n4792_), .B(_abc_41356_new_n4795_), .Y(_abc_41356_new_n4796_));
OR2X2 OR2X2_154 ( .A(_abc_41356_new_n1006_), .B(_abc_41356_new_n1009_), .Y(_abc_41356_new_n1010_));
OR2X2 OR2X2_1540 ( .A(_abc_41356_new_n4800_), .B(_abc_41356_new_n4799_), .Y(_abc_41356_new_n4801_));
OR2X2 OR2X2_1541 ( .A(_abc_41356_new_n4802_), .B(_abc_41356_new_n4798_), .Y(_abc_41356_new_n4803_));
OR2X2 OR2X2_1542 ( .A(_abc_41356_new_n4797_), .B(_abc_41356_new_n4803_), .Y(_abc_41356_new_n4804_));
OR2X2 OR2X2_1543 ( .A(_abc_41356_new_n4804_), .B(_abc_41356_new_n4791_), .Y(_abc_41356_new_n4805_));
OR2X2 OR2X2_1544 ( .A(_abc_41356_new_n4813_), .B(_abc_41356_new_n4809_), .Y(_abc_41356_new_n4814_));
OR2X2 OR2X2_1545 ( .A(_abc_41356_new_n4808_), .B(_abc_41356_new_n4814_), .Y(_abc_41356_new_n4815_));
OR2X2 OR2X2_1546 ( .A(_abc_41356_new_n4806_), .B(_abc_41356_new_n4815_), .Y(_abc_41356_new_n4816_));
OR2X2 OR2X2_1547 ( .A(_abc_41356_new_n4817_), .B(_abc_41356_new_n4778_), .Y(_0raddrhold_15_0__15_));
OR2X2 OR2X2_1548 ( .A(_abc_41356_new_n4820_), .B(reset), .Y(_abc_41356_new_n4821_));
OR2X2 OR2X2_1549 ( .A(_abc_41356_new_n2096_), .B(waddrhold_0_), .Y(_abc_41356_new_n4823_));
OR2X2 OR2X2_155 ( .A(_abc_41356_new_n1010_), .B(opcode_2_), .Y(_abc_41356_new_n1011_));
OR2X2 OR2X2_1550 ( .A(_abc_41356_new_n2069_), .B(sp_0_), .Y(_abc_41356_new_n4824_));
OR2X2 OR2X2_1551 ( .A(_abc_41356_new_n4829_), .B(_abc_41356_new_n4183_), .Y(_abc_41356_new_n4830_));
OR2X2 OR2X2_1552 ( .A(_abc_41356_new_n682_), .B(waddrhold_0_), .Y(_abc_41356_new_n4834_));
OR2X2 OR2X2_1553 ( .A(_abc_41356_new_n4836_), .B(_abc_41356_new_n4837_), .Y(_abc_41356_new_n4838_));
OR2X2 OR2X2_1554 ( .A(_abc_41356_new_n4839_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4840_));
OR2X2 OR2X2_1555 ( .A(_abc_41356_new_n4840_), .B(_abc_41356_new_n4833_), .Y(_abc_41356_new_n4841_));
OR2X2 OR2X2_1556 ( .A(_abc_41356_new_n4841_), .B(_abc_41356_new_n4831_), .Y(_abc_41356_new_n4842_));
OR2X2 OR2X2_1557 ( .A(_abc_41356_new_n4826_), .B(_abc_41356_new_n4842_), .Y(_abc_41356_new_n4843_));
OR2X2 OR2X2_1558 ( .A(_abc_41356_new_n2887_), .B(waddrhold_0_), .Y(_abc_41356_new_n4844_));
OR2X2 OR2X2_1559 ( .A(_abc_41356_new_n4849_), .B(_abc_41356_new_n4850_), .Y(_abc_41356_new_n4851_));
OR2X2 OR2X2_156 ( .A(_abc_41356_new_n1013_), .B(_abc_41356_new_n1014_), .Y(_abc_41356_new_n1015_));
OR2X2 OR2X2_1560 ( .A(_abc_41356_new_n4851_), .B(_abc_41356_new_n4847_), .Y(_abc_41356_new_n4852_));
OR2X2 OR2X2_1561 ( .A(_abc_41356_new_n4846_), .B(_abc_41356_new_n4852_), .Y(_abc_41356_new_n4853_));
OR2X2 OR2X2_1562 ( .A(_abc_41356_new_n4854_), .B(_abc_41356_new_n4822_), .Y(_0waddrhold_15_0__0_));
OR2X2 OR2X2_1563 ( .A(_abc_41356_new_n4859_), .B(_abc_41356_new_n4858_), .Y(_abc_41356_new_n4860_));
OR2X2 OR2X2_1564 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n4862_), .Y(_abc_41356_new_n4863_));
OR2X2 OR2X2_1565 ( .A(_abc_41356_new_n4861_), .B(_abc_41356_new_n4863_), .Y(_abc_41356_new_n4864_));
OR2X2 OR2X2_1566 ( .A(_abc_41356_new_n2096_), .B(waddrhold_1_), .Y(_abc_41356_new_n4865_));
OR2X2 OR2X2_1567 ( .A(_abc_41356_new_n682_), .B(waddrhold_1_), .Y(_abc_41356_new_n4871_));
OR2X2 OR2X2_1568 ( .A(_abc_41356_new_n4873_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4874_));
OR2X2 OR2X2_1569 ( .A(_abc_41356_new_n4874_), .B(_abc_41356_new_n4870_), .Y(_abc_41356_new_n4875_));
OR2X2 OR2X2_157 ( .A(_abc_41356_new_n1016_), .B(_abc_41356_new_n995_), .Y(_abc_41356_new_n1017_));
OR2X2 OR2X2_1570 ( .A(_abc_41356_new_n4875_), .B(_abc_41356_new_n4868_), .Y(_abc_41356_new_n4876_));
OR2X2 OR2X2_1571 ( .A(_abc_41356_new_n4867_), .B(_abc_41356_new_n4876_), .Y(_abc_41356_new_n4877_));
OR2X2 OR2X2_1572 ( .A(_abc_41356_new_n2887_), .B(waddrhold_1_), .Y(_abc_41356_new_n4878_));
OR2X2 OR2X2_1573 ( .A(waddrhold_0_), .B(waddrhold_1_), .Y(_abc_41356_new_n4885_));
OR2X2 OR2X2_1574 ( .A(_abc_41356_new_n4887_), .B(_abc_41356_new_n4882_), .Y(_abc_41356_new_n4888_));
OR2X2 OR2X2_1575 ( .A(_abc_41356_new_n4888_), .B(_abc_41356_new_n4881_), .Y(_abc_41356_new_n4889_));
OR2X2 OR2X2_1576 ( .A(_abc_41356_new_n4880_), .B(_abc_41356_new_n4889_), .Y(_abc_41356_new_n4890_));
OR2X2 OR2X2_1577 ( .A(_abc_41356_new_n4891_), .B(_abc_41356_new_n4856_), .Y(_0waddrhold_15_0__1_));
OR2X2 OR2X2_1578 ( .A(_abc_41356_new_n4894_), .B(_abc_41356_new_n4895_), .Y(_abc_41356_new_n4896_));
OR2X2 OR2X2_1579 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n4898_), .Y(_abc_41356_new_n4899_));
OR2X2 OR2X2_158 ( .A(_abc_41356_new_n994_), .B(_abc_41356_new_n1017_), .Y(_abc_41356_new_n1018_));
OR2X2 OR2X2_1580 ( .A(_abc_41356_new_n4897_), .B(_abc_41356_new_n4899_), .Y(_abc_41356_new_n4900_));
OR2X2 OR2X2_1581 ( .A(_abc_41356_new_n2096_), .B(waddrhold_2_), .Y(_abc_41356_new_n4901_));
OR2X2 OR2X2_1582 ( .A(_abc_41356_new_n682_), .B(waddrhold_2_), .Y(_abc_41356_new_n4907_));
OR2X2 OR2X2_1583 ( .A(_abc_41356_new_n4909_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4910_));
OR2X2 OR2X2_1584 ( .A(_abc_41356_new_n4910_), .B(_abc_41356_new_n4906_), .Y(_abc_41356_new_n4911_));
OR2X2 OR2X2_1585 ( .A(_abc_41356_new_n4911_), .B(_abc_41356_new_n4904_), .Y(_abc_41356_new_n4912_));
OR2X2 OR2X2_1586 ( .A(_abc_41356_new_n4903_), .B(_abc_41356_new_n4912_), .Y(_abc_41356_new_n4913_));
OR2X2 OR2X2_1587 ( .A(_abc_41356_new_n2887_), .B(waddrhold_2_), .Y(_abc_41356_new_n4914_));
OR2X2 OR2X2_1588 ( .A(_abc_41356_new_n4883_), .B(waddrhold_2_), .Y(_abc_41356_new_n4919_));
OR2X2 OR2X2_1589 ( .A(_abc_41356_new_n4923_), .B(_abc_41356_new_n4918_), .Y(_abc_41356_new_n4924_));
OR2X2 OR2X2_159 ( .A(_abc_41356_new_n989_), .B(_abc_41356_new_n1018_), .Y(_abc_41356_new_n1019_));
OR2X2 OR2X2_1590 ( .A(_abc_41356_new_n4924_), .B(_abc_41356_new_n4917_), .Y(_abc_41356_new_n4925_));
OR2X2 OR2X2_1591 ( .A(_abc_41356_new_n4916_), .B(_abc_41356_new_n4925_), .Y(_abc_41356_new_n4926_));
OR2X2 OR2X2_1592 ( .A(_abc_41356_new_n4927_), .B(_abc_41356_new_n4893_), .Y(_0waddrhold_15_0__2_));
OR2X2 OR2X2_1593 ( .A(_abc_41356_new_n4930_), .B(_abc_41356_new_n1303_), .Y(_abc_41356_new_n4931_));
OR2X2 OR2X2_1594 ( .A(_abc_41356_new_n4894_), .B(sp_3_), .Y(_abc_41356_new_n4932_));
OR2X2 OR2X2_1595 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n4935_), .Y(_abc_41356_new_n4936_));
OR2X2 OR2X2_1596 ( .A(_abc_41356_new_n4934_), .B(_abc_41356_new_n4936_), .Y(_abc_41356_new_n4937_));
OR2X2 OR2X2_1597 ( .A(_abc_41356_new_n2096_), .B(waddrhold_3_), .Y(_abc_41356_new_n4938_));
OR2X2 OR2X2_1598 ( .A(_abc_41356_new_n682_), .B(waddrhold_3_), .Y(_abc_41356_new_n4944_));
OR2X2 OR2X2_1599 ( .A(_abc_41356_new_n4946_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4947_));
OR2X2 OR2X2_16 ( .A(_abc_41356_new_n633_), .B(_abc_41356_new_n630_), .Y(_abc_41356_new_n634_));
OR2X2 OR2X2_160 ( .A(_abc_41356_new_n1019_), .B(_abc_41356_new_n696_), .Y(_abc_41356_new_n1020_));
OR2X2 OR2X2_1600 ( .A(_abc_41356_new_n4947_), .B(_abc_41356_new_n4943_), .Y(_abc_41356_new_n4948_));
OR2X2 OR2X2_1601 ( .A(_abc_41356_new_n4948_), .B(_abc_41356_new_n4941_), .Y(_abc_41356_new_n4949_));
OR2X2 OR2X2_1602 ( .A(_abc_41356_new_n4940_), .B(_abc_41356_new_n4949_), .Y(_abc_41356_new_n4950_));
OR2X2 OR2X2_1603 ( .A(_abc_41356_new_n2887_), .B(waddrhold_3_), .Y(_abc_41356_new_n4951_));
OR2X2 OR2X2_1604 ( .A(_abc_41356_new_n4920_), .B(waddrhold_3_), .Y(_abc_41356_new_n4958_));
OR2X2 OR2X2_1605 ( .A(_abc_41356_new_n4960_), .B(_abc_41356_new_n4955_), .Y(_abc_41356_new_n4961_));
OR2X2 OR2X2_1606 ( .A(_abc_41356_new_n4961_), .B(_abc_41356_new_n4954_), .Y(_abc_41356_new_n4962_));
OR2X2 OR2X2_1607 ( .A(_abc_41356_new_n4953_), .B(_abc_41356_new_n4962_), .Y(_abc_41356_new_n4963_));
OR2X2 OR2X2_1608 ( .A(_abc_41356_new_n4964_), .B(_abc_41356_new_n4929_), .Y(_0waddrhold_15_0__3_));
OR2X2 OR2X2_1609 ( .A(_abc_41356_new_n4970_), .B(_abc_41356_new_n4968_), .Y(_abc_41356_new_n4971_));
OR2X2 OR2X2_161 ( .A(_abc_41356_new_n695_), .B(regfil_7__5_), .Y(_abc_41356_new_n1021_));
OR2X2 OR2X2_1610 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n4973_), .Y(_abc_41356_new_n4974_));
OR2X2 OR2X2_1611 ( .A(_abc_41356_new_n4972_), .B(_abc_41356_new_n4974_), .Y(_abc_41356_new_n4975_));
OR2X2 OR2X2_1612 ( .A(_abc_41356_new_n2096_), .B(waddrhold_4_), .Y(_abc_41356_new_n4976_));
OR2X2 OR2X2_1613 ( .A(_abc_41356_new_n682_), .B(waddrhold_4_), .Y(_abc_41356_new_n4982_));
OR2X2 OR2X2_1614 ( .A(_abc_41356_new_n4984_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n4985_));
OR2X2 OR2X2_1615 ( .A(_abc_41356_new_n4985_), .B(_abc_41356_new_n4981_), .Y(_abc_41356_new_n4986_));
OR2X2 OR2X2_1616 ( .A(_abc_41356_new_n4986_), .B(_abc_41356_new_n4979_), .Y(_abc_41356_new_n4987_));
OR2X2 OR2X2_1617 ( .A(_abc_41356_new_n4978_), .B(_abc_41356_new_n4987_), .Y(_abc_41356_new_n4988_));
OR2X2 OR2X2_1618 ( .A(_abc_41356_new_n2887_), .B(waddrhold_4_), .Y(_abc_41356_new_n4989_));
OR2X2 OR2X2_1619 ( .A(_abc_41356_new_n4993_), .B(_abc_41356_new_n4992_), .Y(_abc_41356_new_n4994_));
OR2X2 OR2X2_162 ( .A(_abc_41356_new_n1027_), .B(_abc_41356_new_n512_), .Y(_abc_41356_new_n1028_));
OR2X2 OR2X2_1620 ( .A(_abc_41356_new_n4956_), .B(waddrhold_4_), .Y(_abc_41356_new_n4997_));
OR2X2 OR2X2_1621 ( .A(_abc_41356_new_n4999_), .B(_abc_41356_new_n4994_), .Y(_abc_41356_new_n5000_));
OR2X2 OR2X2_1622 ( .A(_abc_41356_new_n4991_), .B(_abc_41356_new_n5000_), .Y(_abc_41356_new_n5001_));
OR2X2 OR2X2_1623 ( .A(_abc_41356_new_n5002_), .B(_abc_41356_new_n4966_), .Y(_0waddrhold_15_0__4_));
OR2X2 OR2X2_1624 ( .A(_abc_41356_new_n5006_), .B(_abc_41356_new_n5007_), .Y(_abc_41356_new_n5008_));
OR2X2 OR2X2_1625 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5010_), .Y(_abc_41356_new_n5011_));
OR2X2 OR2X2_1626 ( .A(_abc_41356_new_n5009_), .B(_abc_41356_new_n5011_), .Y(_abc_41356_new_n5012_));
OR2X2 OR2X2_1627 ( .A(_abc_41356_new_n2096_), .B(waddrhold_5_), .Y(_abc_41356_new_n5013_));
OR2X2 OR2X2_1628 ( .A(_abc_41356_new_n682_), .B(waddrhold_5_), .Y(_abc_41356_new_n5019_));
OR2X2 OR2X2_1629 ( .A(_abc_41356_new_n5021_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5022_));
OR2X2 OR2X2_163 ( .A(_abc_41356_new_n1039_), .B(_abc_41356_new_n555_), .Y(_abc_41356_new_n1040_));
OR2X2 OR2X2_1630 ( .A(_abc_41356_new_n5022_), .B(_abc_41356_new_n5018_), .Y(_abc_41356_new_n5023_));
OR2X2 OR2X2_1631 ( .A(_abc_41356_new_n5023_), .B(_abc_41356_new_n5016_), .Y(_abc_41356_new_n5024_));
OR2X2 OR2X2_1632 ( .A(_abc_41356_new_n5015_), .B(_abc_41356_new_n5024_), .Y(_abc_41356_new_n5025_));
OR2X2 OR2X2_1633 ( .A(_abc_41356_new_n2887_), .B(waddrhold_5_), .Y(_abc_41356_new_n5026_));
OR2X2 OR2X2_1634 ( .A(_abc_41356_new_n5030_), .B(_abc_41356_new_n5029_), .Y(_abc_41356_new_n5031_));
OR2X2 OR2X2_1635 ( .A(_abc_41356_new_n4995_), .B(waddrhold_5_), .Y(_abc_41356_new_n5034_));
OR2X2 OR2X2_1636 ( .A(_abc_41356_new_n5036_), .B(_abc_41356_new_n5031_), .Y(_abc_41356_new_n5037_));
OR2X2 OR2X2_1637 ( .A(_abc_41356_new_n5028_), .B(_abc_41356_new_n5037_), .Y(_abc_41356_new_n5038_));
OR2X2 OR2X2_1638 ( .A(_abc_41356_new_n5039_), .B(_abc_41356_new_n5004_), .Y(_0waddrhold_15_0__5_));
OR2X2 OR2X2_1639 ( .A(_abc_41356_new_n5044_), .B(_abc_41356_new_n5042_), .Y(_abc_41356_new_n5045_));
OR2X2 OR2X2_164 ( .A(_abc_41356_new_n1038_), .B(_abc_41356_new_n1040_), .Y(_abc_41356_new_n1041_));
OR2X2 OR2X2_1640 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5047_), .Y(_abc_41356_new_n5048_));
OR2X2 OR2X2_1641 ( .A(_abc_41356_new_n5046_), .B(_abc_41356_new_n5048_), .Y(_abc_41356_new_n5049_));
OR2X2 OR2X2_1642 ( .A(_abc_41356_new_n2096_), .B(waddrhold_6_), .Y(_abc_41356_new_n5050_));
OR2X2 OR2X2_1643 ( .A(_abc_41356_new_n682_), .B(waddrhold_6_), .Y(_abc_41356_new_n5056_));
OR2X2 OR2X2_1644 ( .A(_abc_41356_new_n5058_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5059_));
OR2X2 OR2X2_1645 ( .A(_abc_41356_new_n5059_), .B(_abc_41356_new_n5055_), .Y(_abc_41356_new_n5060_));
OR2X2 OR2X2_1646 ( .A(_abc_41356_new_n5060_), .B(_abc_41356_new_n5053_), .Y(_abc_41356_new_n5061_));
OR2X2 OR2X2_1647 ( .A(_abc_41356_new_n5052_), .B(_abc_41356_new_n5061_), .Y(_abc_41356_new_n5062_));
OR2X2 OR2X2_1648 ( .A(_abc_41356_new_n2887_), .B(waddrhold_6_), .Y(_abc_41356_new_n5063_));
OR2X2 OR2X2_1649 ( .A(_abc_41356_new_n5067_), .B(_abc_41356_new_n5066_), .Y(_abc_41356_new_n5068_));
OR2X2 OR2X2_165 ( .A(_abc_41356_new_n1042_), .B(_abc_41356_new_n1028_), .Y(_abc_41356_new_n1043_));
OR2X2 OR2X2_1650 ( .A(_abc_41356_new_n5032_), .B(waddrhold_6_), .Y(_abc_41356_new_n5071_));
OR2X2 OR2X2_1651 ( .A(_abc_41356_new_n5073_), .B(_abc_41356_new_n5068_), .Y(_abc_41356_new_n5074_));
OR2X2 OR2X2_1652 ( .A(_abc_41356_new_n5065_), .B(_abc_41356_new_n5074_), .Y(_abc_41356_new_n5075_));
OR2X2 OR2X2_1653 ( .A(_abc_41356_new_n5076_), .B(_abc_41356_new_n5041_), .Y(_0waddrhold_15_0__6_));
OR2X2 OR2X2_1654 ( .A(_abc_41356_new_n5080_), .B(_abc_41356_new_n5081_), .Y(_abc_41356_new_n5082_));
OR2X2 OR2X2_1655 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5084_), .Y(_abc_41356_new_n5085_));
OR2X2 OR2X2_1656 ( .A(_abc_41356_new_n5083_), .B(_abc_41356_new_n5085_), .Y(_abc_41356_new_n5086_));
OR2X2 OR2X2_1657 ( .A(_abc_41356_new_n2096_), .B(waddrhold_7_), .Y(_abc_41356_new_n5087_));
OR2X2 OR2X2_1658 ( .A(_abc_41356_new_n682_), .B(waddrhold_7_), .Y(_abc_41356_new_n5093_));
OR2X2 OR2X2_1659 ( .A(_abc_41356_new_n5095_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5096_));
OR2X2 OR2X2_166 ( .A(_abc_41356_new_n1047_), .B(_abc_41356_new_n1046_), .Y(_abc_41356_new_n1048_));
OR2X2 OR2X2_1660 ( .A(_abc_41356_new_n5096_), .B(_abc_41356_new_n5092_), .Y(_abc_41356_new_n5097_));
OR2X2 OR2X2_1661 ( .A(_abc_41356_new_n5097_), .B(_abc_41356_new_n5090_), .Y(_abc_41356_new_n5098_));
OR2X2 OR2X2_1662 ( .A(_abc_41356_new_n5089_), .B(_abc_41356_new_n5098_), .Y(_abc_41356_new_n5099_));
OR2X2 OR2X2_1663 ( .A(_abc_41356_new_n2887_), .B(waddrhold_7_), .Y(_abc_41356_new_n5100_));
OR2X2 OR2X2_1664 ( .A(_abc_41356_new_n5104_), .B(_abc_41356_new_n5103_), .Y(_abc_41356_new_n5105_));
OR2X2 OR2X2_1665 ( .A(_abc_41356_new_n5069_), .B(waddrhold_7_), .Y(_abc_41356_new_n5108_));
OR2X2 OR2X2_1666 ( .A(_abc_41356_new_n5110_), .B(_abc_41356_new_n5105_), .Y(_abc_41356_new_n5111_));
OR2X2 OR2X2_1667 ( .A(_abc_41356_new_n5102_), .B(_abc_41356_new_n5111_), .Y(_abc_41356_new_n5112_));
OR2X2 OR2X2_1668 ( .A(_abc_41356_new_n5113_), .B(_abc_41356_new_n5078_), .Y(_0waddrhold_15_0__7_));
OR2X2 OR2X2_1669 ( .A(_abc_41356_new_n5118_), .B(_abc_41356_new_n5116_), .Y(_abc_41356_new_n5119_));
OR2X2 OR2X2_167 ( .A(_abc_41356_new_n1048_), .B(_abc_41356_new_n1045_), .Y(_abc_41356_new_n1049_));
OR2X2 OR2X2_1670 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5121_), .Y(_abc_41356_new_n5122_));
OR2X2 OR2X2_1671 ( .A(_abc_41356_new_n5120_), .B(_abc_41356_new_n5122_), .Y(_abc_41356_new_n5123_));
OR2X2 OR2X2_1672 ( .A(_abc_41356_new_n2096_), .B(waddrhold_8_), .Y(_abc_41356_new_n5124_));
OR2X2 OR2X2_1673 ( .A(_abc_41356_new_n682_), .B(waddrhold_8_), .Y(_abc_41356_new_n5130_));
OR2X2 OR2X2_1674 ( .A(_abc_41356_new_n5132_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5133_));
OR2X2 OR2X2_1675 ( .A(_abc_41356_new_n5133_), .B(_abc_41356_new_n5129_), .Y(_abc_41356_new_n5134_));
OR2X2 OR2X2_1676 ( .A(_abc_41356_new_n5134_), .B(_abc_41356_new_n5127_), .Y(_abc_41356_new_n5135_));
OR2X2 OR2X2_1677 ( .A(_abc_41356_new_n5126_), .B(_abc_41356_new_n5135_), .Y(_abc_41356_new_n5136_));
OR2X2 OR2X2_1678 ( .A(_abc_41356_new_n2887_), .B(waddrhold_8_), .Y(_abc_41356_new_n5137_));
OR2X2 OR2X2_1679 ( .A(_abc_41356_new_n5141_), .B(_abc_41356_new_n5140_), .Y(_abc_41356_new_n5142_));
OR2X2 OR2X2_168 ( .A(_abc_41356_new_n1044_), .B(_abc_41356_new_n1049_), .Y(_abc_41356_new_n1050_));
OR2X2 OR2X2_1680 ( .A(_abc_41356_new_n5106_), .B(waddrhold_8_), .Y(_abc_41356_new_n5145_));
OR2X2 OR2X2_1681 ( .A(_abc_41356_new_n5147_), .B(_abc_41356_new_n5142_), .Y(_abc_41356_new_n5148_));
OR2X2 OR2X2_1682 ( .A(_abc_41356_new_n5139_), .B(_abc_41356_new_n5148_), .Y(_abc_41356_new_n5149_));
OR2X2 OR2X2_1683 ( .A(_abc_41356_new_n5150_), .B(_abc_41356_new_n5115_), .Y(_0waddrhold_15_0__8_));
OR2X2 OR2X2_1684 ( .A(_abc_41356_new_n5154_), .B(_abc_41356_new_n5155_), .Y(_abc_41356_new_n5156_));
OR2X2 OR2X2_1685 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5158_), .Y(_abc_41356_new_n5159_));
OR2X2 OR2X2_1686 ( .A(_abc_41356_new_n5157_), .B(_abc_41356_new_n5159_), .Y(_abc_41356_new_n5160_));
OR2X2 OR2X2_1687 ( .A(_abc_41356_new_n2096_), .B(waddrhold_9_), .Y(_abc_41356_new_n5161_));
OR2X2 OR2X2_1688 ( .A(_abc_41356_new_n682_), .B(waddrhold_9_), .Y(_abc_41356_new_n5167_));
OR2X2 OR2X2_1689 ( .A(_abc_41356_new_n5169_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5170_));
OR2X2 OR2X2_169 ( .A(_abc_41356_new_n1023_), .B(_abc_41356_new_n1050_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_5_));
OR2X2 OR2X2_1690 ( .A(_abc_41356_new_n5170_), .B(_abc_41356_new_n5166_), .Y(_abc_41356_new_n5171_));
OR2X2 OR2X2_1691 ( .A(_abc_41356_new_n5171_), .B(_abc_41356_new_n5164_), .Y(_abc_41356_new_n5172_));
OR2X2 OR2X2_1692 ( .A(_abc_41356_new_n5163_), .B(_abc_41356_new_n5172_), .Y(_abc_41356_new_n5173_));
OR2X2 OR2X2_1693 ( .A(_abc_41356_new_n2887_), .B(waddrhold_9_), .Y(_abc_41356_new_n5174_));
OR2X2 OR2X2_1694 ( .A(_abc_41356_new_n5178_), .B(_abc_41356_new_n5177_), .Y(_abc_41356_new_n5179_));
OR2X2 OR2X2_1695 ( .A(_abc_41356_new_n5143_), .B(waddrhold_9_), .Y(_abc_41356_new_n5182_));
OR2X2 OR2X2_1696 ( .A(_abc_41356_new_n5184_), .B(_abc_41356_new_n5179_), .Y(_abc_41356_new_n5185_));
OR2X2 OR2X2_1697 ( .A(_abc_41356_new_n5176_), .B(_abc_41356_new_n5185_), .Y(_abc_41356_new_n5186_));
OR2X2 OR2X2_1698 ( .A(_abc_41356_new_n5187_), .B(_abc_41356_new_n5152_), .Y(_0waddrhold_15_0__9_));
OR2X2 OR2X2_1699 ( .A(_abc_41356_new_n5192_), .B(_abc_41356_new_n5190_), .Y(_abc_41356_new_n5193_));
OR2X2 OR2X2_17 ( .A(_abc_41356_new_n634_), .B(_abc_41356_new_n629_), .Y(_abc_41356_new_n635_));
OR2X2 OR2X2_170 ( .A(_abc_41356_new_n1053_), .B(_abc_41356_new_n1054_), .Y(_abc_41356_new_n1055_));
OR2X2 OR2X2_1700 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5195_), .Y(_abc_41356_new_n5196_));
OR2X2 OR2X2_1701 ( .A(_abc_41356_new_n5194_), .B(_abc_41356_new_n5196_), .Y(_abc_41356_new_n5197_));
OR2X2 OR2X2_1702 ( .A(_abc_41356_new_n2096_), .B(waddrhold_10_), .Y(_abc_41356_new_n5198_));
OR2X2 OR2X2_1703 ( .A(_abc_41356_new_n682_), .B(waddrhold_10_), .Y(_abc_41356_new_n5204_));
OR2X2 OR2X2_1704 ( .A(_abc_41356_new_n5206_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5207_));
OR2X2 OR2X2_1705 ( .A(_abc_41356_new_n5207_), .B(_abc_41356_new_n5203_), .Y(_abc_41356_new_n5208_));
OR2X2 OR2X2_1706 ( .A(_abc_41356_new_n5208_), .B(_abc_41356_new_n5201_), .Y(_abc_41356_new_n5209_));
OR2X2 OR2X2_1707 ( .A(_abc_41356_new_n5200_), .B(_abc_41356_new_n5209_), .Y(_abc_41356_new_n5210_));
OR2X2 OR2X2_1708 ( .A(_abc_41356_new_n2887_), .B(waddrhold_10_), .Y(_abc_41356_new_n5211_));
OR2X2 OR2X2_1709 ( .A(_abc_41356_new_n5215_), .B(_abc_41356_new_n5214_), .Y(_abc_41356_new_n5216_));
OR2X2 OR2X2_171 ( .A(_abc_41356_new_n1057_), .B(_abc_41356_new_n1056_), .Y(_abc_41356_new_n1058_));
OR2X2 OR2X2_1710 ( .A(_abc_41356_new_n5180_), .B(waddrhold_10_), .Y(_abc_41356_new_n5219_));
OR2X2 OR2X2_1711 ( .A(_abc_41356_new_n5221_), .B(_abc_41356_new_n5216_), .Y(_abc_41356_new_n5222_));
OR2X2 OR2X2_1712 ( .A(_abc_41356_new_n5213_), .B(_abc_41356_new_n5222_), .Y(_abc_41356_new_n5223_));
OR2X2 OR2X2_1713 ( .A(_abc_41356_new_n5224_), .B(_abc_41356_new_n5189_), .Y(_0waddrhold_15_0__10_));
OR2X2 OR2X2_1714 ( .A(_abc_41356_new_n5228_), .B(_abc_41356_new_n5229_), .Y(_abc_41356_new_n5230_));
OR2X2 OR2X2_1715 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5232_), .Y(_abc_41356_new_n5233_));
OR2X2 OR2X2_1716 ( .A(_abc_41356_new_n5231_), .B(_abc_41356_new_n5233_), .Y(_abc_41356_new_n5234_));
OR2X2 OR2X2_1717 ( .A(_abc_41356_new_n2096_), .B(waddrhold_11_), .Y(_abc_41356_new_n5235_));
OR2X2 OR2X2_1718 ( .A(_abc_41356_new_n682_), .B(waddrhold_11_), .Y(_abc_41356_new_n5241_));
OR2X2 OR2X2_1719 ( .A(_abc_41356_new_n5243_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5244_));
OR2X2 OR2X2_172 ( .A(_abc_41356_new_n1055_), .B(_abc_41356_new_n1058_), .Y(_abc_41356_new_n1059_));
OR2X2 OR2X2_1720 ( .A(_abc_41356_new_n5244_), .B(_abc_41356_new_n5240_), .Y(_abc_41356_new_n5245_));
OR2X2 OR2X2_1721 ( .A(_abc_41356_new_n5245_), .B(_abc_41356_new_n5238_), .Y(_abc_41356_new_n5246_));
OR2X2 OR2X2_1722 ( .A(_abc_41356_new_n5237_), .B(_abc_41356_new_n5246_), .Y(_abc_41356_new_n5247_));
OR2X2 OR2X2_1723 ( .A(_abc_41356_new_n2887_), .B(waddrhold_11_), .Y(_abc_41356_new_n5248_));
OR2X2 OR2X2_1724 ( .A(_abc_41356_new_n5252_), .B(_abc_41356_new_n5251_), .Y(_abc_41356_new_n5253_));
OR2X2 OR2X2_1725 ( .A(_abc_41356_new_n5217_), .B(waddrhold_11_), .Y(_abc_41356_new_n5256_));
OR2X2 OR2X2_1726 ( .A(_abc_41356_new_n5258_), .B(_abc_41356_new_n5253_), .Y(_abc_41356_new_n5259_));
OR2X2 OR2X2_1727 ( .A(_abc_41356_new_n5250_), .B(_abc_41356_new_n5259_), .Y(_abc_41356_new_n5260_));
OR2X2 OR2X2_1728 ( .A(_abc_41356_new_n5261_), .B(_abc_41356_new_n5226_), .Y(_0waddrhold_15_0__11_));
OR2X2 OR2X2_1729 ( .A(_abc_41356_new_n5264_), .B(_abc_41356_new_n5263_), .Y(_abc_41356_new_n5265_));
OR2X2 OR2X2_173 ( .A(_abc_41356_new_n1059_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n1060_));
OR2X2 OR2X2_1730 ( .A(_abc_41356_new_n5268_), .B(_abc_41356_new_n5266_), .Y(_abc_41356_new_n5269_));
OR2X2 OR2X2_1731 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5271_), .Y(_abc_41356_new_n5272_));
OR2X2 OR2X2_1732 ( .A(_abc_41356_new_n5270_), .B(_abc_41356_new_n5272_), .Y(_abc_41356_new_n5273_));
OR2X2 OR2X2_1733 ( .A(_abc_41356_new_n2096_), .B(waddrhold_12_), .Y(_abc_41356_new_n5274_));
OR2X2 OR2X2_1734 ( .A(_abc_41356_new_n682_), .B(waddrhold_12_), .Y(_abc_41356_new_n5278_));
OR2X2 OR2X2_1735 ( .A(_abc_41356_new_n5282_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5283_));
OR2X2 OR2X2_1736 ( .A(_abc_41356_new_n5280_), .B(_abc_41356_new_n5283_), .Y(_abc_41356_new_n5284_));
OR2X2 OR2X2_1737 ( .A(_abc_41356_new_n5284_), .B(_abc_41356_new_n5277_), .Y(_abc_41356_new_n5285_));
OR2X2 OR2X2_1738 ( .A(_abc_41356_new_n5276_), .B(_abc_41356_new_n5285_), .Y(_abc_41356_new_n5286_));
OR2X2 OR2X2_1739 ( .A(_abc_41356_new_n2887_), .B(waddrhold_12_), .Y(_abc_41356_new_n5287_));
OR2X2 OR2X2_174 ( .A(_abc_41356_new_n1061_), .B(_abc_41356_new_n1062_), .Y(_abc_41356_new_n1063_));
OR2X2 OR2X2_1740 ( .A(_abc_41356_new_n5289_), .B(_abc_41356_new_n5265_), .Y(_abc_41356_new_n5290_));
OR2X2 OR2X2_1741 ( .A(_abc_41356_new_n5254_), .B(waddrhold_12_), .Y(_abc_41356_new_n5294_));
OR2X2 OR2X2_1742 ( .A(_abc_41356_new_n5297_), .B(_abc_41356_new_n5298_), .Y(_abc_41356_new_n5299_));
OR2X2 OR2X2_1743 ( .A(_abc_41356_new_n5291_), .B(_abc_41356_new_n5299_), .Y(_0waddrhold_15_0__12_));
OR2X2 OR2X2_1744 ( .A(_abc_41356_new_n5302_), .B(_abc_41356_new_n5301_), .Y(_abc_41356_new_n5303_));
OR2X2 OR2X2_1745 ( .A(_abc_41356_new_n5305_), .B(_abc_41356_new_n5306_), .Y(_abc_41356_new_n5307_));
OR2X2 OR2X2_1746 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5309_), .Y(_abc_41356_new_n5310_));
OR2X2 OR2X2_1747 ( .A(_abc_41356_new_n5308_), .B(_abc_41356_new_n5310_), .Y(_abc_41356_new_n5311_));
OR2X2 OR2X2_1748 ( .A(_abc_41356_new_n2096_), .B(waddrhold_13_), .Y(_abc_41356_new_n5312_));
OR2X2 OR2X2_1749 ( .A(_abc_41356_new_n682_), .B(waddrhold_13_), .Y(_abc_41356_new_n5318_));
OR2X2 OR2X2_175 ( .A(_abc_41356_new_n1065_), .B(_abc_41356_new_n1064_), .Y(_abc_41356_new_n1066_));
OR2X2 OR2X2_1750 ( .A(_abc_41356_new_n5320_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5321_));
OR2X2 OR2X2_1751 ( .A(_abc_41356_new_n5321_), .B(_abc_41356_new_n5317_), .Y(_abc_41356_new_n5322_));
OR2X2 OR2X2_1752 ( .A(_abc_41356_new_n5322_), .B(_abc_41356_new_n5315_), .Y(_abc_41356_new_n5323_));
OR2X2 OR2X2_1753 ( .A(_abc_41356_new_n5314_), .B(_abc_41356_new_n5323_), .Y(_abc_41356_new_n5324_));
OR2X2 OR2X2_1754 ( .A(_abc_41356_new_n2887_), .B(waddrhold_13_), .Y(_abc_41356_new_n5325_));
OR2X2 OR2X2_1755 ( .A(_abc_41356_new_n5327_), .B(_abc_41356_new_n5303_), .Y(_abc_41356_new_n5328_));
OR2X2 OR2X2_1756 ( .A(_abc_41356_new_n5292_), .B(waddrhold_13_), .Y(_abc_41356_new_n5331_));
OR2X2 OR2X2_1757 ( .A(_abc_41356_new_n5335_), .B(_abc_41356_new_n5330_), .Y(_abc_41356_new_n5336_));
OR2X2 OR2X2_1758 ( .A(_abc_41356_new_n5329_), .B(_abc_41356_new_n5336_), .Y(_0waddrhold_15_0__13_));
OR2X2 OR2X2_1759 ( .A(_abc_41356_new_n5339_), .B(_abc_41356_new_n5338_), .Y(_abc_41356_new_n5340_));
OR2X2 OR2X2_176 ( .A(_abc_41356_new_n1063_), .B(_abc_41356_new_n1066_), .Y(_abc_41356_new_n1067_));
OR2X2 OR2X2_1760 ( .A(_abc_41356_new_n5343_), .B(_abc_41356_new_n5341_), .Y(_abc_41356_new_n5344_));
OR2X2 OR2X2_1761 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5346_), .Y(_abc_41356_new_n5347_));
OR2X2 OR2X2_1762 ( .A(_abc_41356_new_n5345_), .B(_abc_41356_new_n5347_), .Y(_abc_41356_new_n5348_));
OR2X2 OR2X2_1763 ( .A(_abc_41356_new_n2096_), .B(waddrhold_14_), .Y(_abc_41356_new_n5349_));
OR2X2 OR2X2_1764 ( .A(_abc_41356_new_n682_), .B(waddrhold_14_), .Y(_abc_41356_new_n5355_));
OR2X2 OR2X2_1765 ( .A(_abc_41356_new_n5357_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5358_));
OR2X2 OR2X2_1766 ( .A(_abc_41356_new_n5358_), .B(_abc_41356_new_n5354_), .Y(_abc_41356_new_n5359_));
OR2X2 OR2X2_1767 ( .A(_abc_41356_new_n5359_), .B(_abc_41356_new_n5352_), .Y(_abc_41356_new_n5360_));
OR2X2 OR2X2_1768 ( .A(_abc_41356_new_n5351_), .B(_abc_41356_new_n5360_), .Y(_abc_41356_new_n5361_));
OR2X2 OR2X2_1769 ( .A(_abc_41356_new_n2887_), .B(waddrhold_14_), .Y(_abc_41356_new_n5362_));
OR2X2 OR2X2_177 ( .A(_abc_41356_new_n1067_), .B(opcode_2_), .Y(_abc_41356_new_n1068_));
OR2X2 OR2X2_1770 ( .A(_abc_41356_new_n5364_), .B(_abc_41356_new_n5340_), .Y(_abc_41356_new_n5365_));
OR2X2 OR2X2_1771 ( .A(_abc_41356_new_n5332_), .B(waddrhold_14_), .Y(_abc_41356_new_n5367_));
OR2X2 OR2X2_1772 ( .A(_abc_41356_new_n5371_), .B(_abc_41356_new_n5368_), .Y(_abc_41356_new_n5372_));
OR2X2 OR2X2_1773 ( .A(_abc_41356_new_n5366_), .B(_abc_41356_new_n5373_), .Y(_0waddrhold_15_0__14_));
OR2X2 OR2X2_1774 ( .A(_abc_41356_new_n5376_), .B(_abc_41356_new_n5375_), .Y(_abc_41356_new_n5377_));
OR2X2 OR2X2_1775 ( .A(_abc_41356_new_n5341_), .B(sp_15_), .Y(_abc_41356_new_n5378_));
OR2X2 OR2X2_1776 ( .A(_abc_41356_new_n5379_), .B(_abc_41356_new_n1967_), .Y(_abc_41356_new_n5380_));
OR2X2 OR2X2_1777 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n5383_), .Y(_abc_41356_new_n5384_));
OR2X2 OR2X2_1778 ( .A(_abc_41356_new_n5382_), .B(_abc_41356_new_n5384_), .Y(_abc_41356_new_n5385_));
OR2X2 OR2X2_1779 ( .A(_abc_41356_new_n2096_), .B(waddrhold_15_), .Y(_abc_41356_new_n5386_));
OR2X2 OR2X2_178 ( .A(_abc_41356_new_n1071_), .B(_abc_41356_new_n1072_), .Y(_abc_41356_new_n1073_));
OR2X2 OR2X2_1780 ( .A(_abc_41356_new_n682_), .B(waddrhold_15_), .Y(_abc_41356_new_n5392_));
OR2X2 OR2X2_1781 ( .A(_abc_41356_new_n5394_), .B(_abc_41356_new_n2886_), .Y(_abc_41356_new_n5395_));
OR2X2 OR2X2_1782 ( .A(_abc_41356_new_n5395_), .B(_abc_41356_new_n5391_), .Y(_abc_41356_new_n5396_));
OR2X2 OR2X2_1783 ( .A(_abc_41356_new_n5396_), .B(_abc_41356_new_n5389_), .Y(_abc_41356_new_n5397_));
OR2X2 OR2X2_1784 ( .A(_abc_41356_new_n5388_), .B(_abc_41356_new_n5397_), .Y(_abc_41356_new_n5398_));
OR2X2 OR2X2_1785 ( .A(_abc_41356_new_n2887_), .B(waddrhold_15_), .Y(_abc_41356_new_n5399_));
OR2X2 OR2X2_1786 ( .A(_abc_41356_new_n5401_), .B(_abc_41356_new_n5377_), .Y(_abc_41356_new_n5402_));
OR2X2 OR2X2_1787 ( .A(_abc_41356_new_n5369_), .B(waddrhold_15_), .Y(_abc_41356_new_n5406_));
OR2X2 OR2X2_1788 ( .A(_abc_41356_new_n5408_), .B(_abc_41356_new_n5409_), .Y(_abc_41356_new_n5410_));
OR2X2 OR2X2_1789 ( .A(_abc_41356_new_n5403_), .B(_abc_41356_new_n5410_), .Y(_0waddrhold_15_0__15_));
OR2X2 OR2X2_179 ( .A(_abc_41356_new_n1070_), .B(_abc_41356_new_n1073_), .Y(_abc_41356_new_n1074_));
OR2X2 OR2X2_1790 ( .A(_abc_41356_new_n5417_), .B(_abc_41356_new_n5418_), .Y(_abc_41356_new_n5419_));
OR2X2 OR2X2_1791 ( .A(_abc_41356_new_n5416_), .B(_abc_41356_new_n5419_), .Y(_0datao_7_0__0_));
OR2X2 OR2X2_1792 ( .A(_abc_41356_new_n5422_), .B(_abc_41356_new_n5423_), .Y(_abc_41356_new_n5424_));
OR2X2 OR2X2_1793 ( .A(_abc_41356_new_n5421_), .B(_abc_41356_new_n5424_), .Y(_0datao_7_0__1_));
OR2X2 OR2X2_1794 ( .A(_abc_41356_new_n5427_), .B(_abc_41356_new_n5428_), .Y(_abc_41356_new_n5429_));
OR2X2 OR2X2_1795 ( .A(_abc_41356_new_n5426_), .B(_abc_41356_new_n5429_), .Y(_0datao_7_0__2_));
OR2X2 OR2X2_1796 ( .A(_abc_41356_new_n5432_), .B(_abc_41356_new_n5433_), .Y(_abc_41356_new_n5434_));
OR2X2 OR2X2_1797 ( .A(_abc_41356_new_n5431_), .B(_abc_41356_new_n5434_), .Y(_0datao_7_0__3_));
OR2X2 OR2X2_1798 ( .A(_abc_41356_new_n5437_), .B(_abc_41356_new_n5438_), .Y(_abc_41356_new_n5439_));
OR2X2 OR2X2_1799 ( .A(_abc_41356_new_n5436_), .B(_abc_41356_new_n5439_), .Y(_0datao_7_0__4_));
OR2X2 OR2X2_18 ( .A(_abc_41356_new_n637_), .B(_abc_41356_new_n638_), .Y(_abc_41356_new_n639_));
OR2X2 OR2X2_180 ( .A(_abc_41356_new_n1077_), .B(_abc_41356_new_n1078_), .Y(_abc_41356_new_n1079_));
OR2X2 OR2X2_1800 ( .A(_abc_41356_new_n5442_), .B(_abc_41356_new_n5443_), .Y(_abc_41356_new_n5444_));
OR2X2 OR2X2_1801 ( .A(_abc_41356_new_n5441_), .B(_abc_41356_new_n5444_), .Y(_0datao_7_0__5_));
OR2X2 OR2X2_1802 ( .A(_abc_41356_new_n5447_), .B(_abc_41356_new_n5448_), .Y(_abc_41356_new_n5449_));
OR2X2 OR2X2_1803 ( .A(_abc_41356_new_n5446_), .B(_abc_41356_new_n5449_), .Y(_0datao_7_0__6_));
OR2X2 OR2X2_1804 ( .A(_abc_41356_new_n5452_), .B(_abc_41356_new_n5453_), .Y(_abc_41356_new_n5454_));
OR2X2 OR2X2_1805 ( .A(_abc_41356_new_n5451_), .B(_abc_41356_new_n5454_), .Y(_0datao_7_0__7_));
OR2X2 OR2X2_1806 ( .A(_abc_41356_new_n2020_), .B(opcode_7_), .Y(_abc_41356_new_n5456_));
OR2X2 OR2X2_1807 ( .A(_abc_41356_new_n5458_), .B(regd_0_), .Y(_abc_41356_new_n5459_));
OR2X2 OR2X2_1808 ( .A(_abc_41356_new_n3410_), .B(_abc_41356_new_n5460_), .Y(_abc_41356_new_n5461_));
OR2X2 OR2X2_1809 ( .A(_abc_41356_new_n3396_), .B(_abc_41356_new_n5463_), .Y(_abc_41356_new_n5464_));
OR2X2 OR2X2_181 ( .A(_abc_41356_new_n985_), .B(regfil_0__6_), .Y(_abc_41356_new_n1083_));
OR2X2 OR2X2_1810 ( .A(_abc_41356_new_n5464_), .B(regd_0_), .Y(_abc_41356_new_n5465_));
OR2X2 OR2X2_1811 ( .A(_abc_41356_new_n5466_), .B(opcode_3_), .Y(_abc_41356_new_n5467_));
OR2X2 OR2X2_1812 ( .A(_abc_41356_new_n5462_), .B(_abc_41356_new_n5469_), .Y(_abc_41356_new_n5470_));
OR2X2 OR2X2_1813 ( .A(_abc_41356_new_n5471_), .B(_abc_41356_new_n5457_), .Y(_0regd_2_0__0_));
OR2X2 OR2X2_1814 ( .A(_abc_41356_new_n5458_), .B(regd_1_), .Y(_abc_41356_new_n5474_));
OR2X2 OR2X2_1815 ( .A(_abc_41356_new_n5464_), .B(regd_1_), .Y(_abc_41356_new_n5477_));
OR2X2 OR2X2_1816 ( .A(_abc_41356_new_n5466_), .B(opcode_4_), .Y(_abc_41356_new_n5478_));
OR2X2 OR2X2_1817 ( .A(_abc_41356_new_n5476_), .B(_abc_41356_new_n5480_), .Y(_abc_41356_new_n5481_));
OR2X2 OR2X2_1818 ( .A(_abc_41356_new_n5482_), .B(_abc_41356_new_n5473_), .Y(_0regd_2_0__1_));
OR2X2 OR2X2_1819 ( .A(_abc_41356_new_n5458_), .B(regd_2_), .Y(_abc_41356_new_n5485_));
OR2X2 OR2X2_182 ( .A(_abc_41356_new_n1085_), .B(_abc_41356_new_n602_), .Y(_abc_41356_new_n1086_));
OR2X2 OR2X2_1820 ( .A(_abc_41356_new_n5464_), .B(regd_2_), .Y(_abc_41356_new_n5488_));
OR2X2 OR2X2_1821 ( .A(_abc_41356_new_n5466_), .B(opcode_5_), .Y(_abc_41356_new_n5489_));
OR2X2 OR2X2_1822 ( .A(_abc_41356_new_n5487_), .B(_abc_41356_new_n5491_), .Y(_abc_41356_new_n5492_));
OR2X2 OR2X2_1823 ( .A(_abc_41356_new_n5493_), .B(_abc_41356_new_n5484_), .Y(_0regd_2_0__2_));
OR2X2 OR2X2_1824 ( .A(_abc_41356_new_n663_), .B(_abc_41356_new_n5496_), .Y(_abc_41356_new_n5497_));
OR2X2 OR2X2_1825 ( .A(_abc_41356_new_n5495_), .B(regfil_5__0_), .Y(_abc_41356_new_n5498_));
OR2X2 OR2X2_1826 ( .A(_abc_41356_new_n1236_), .B(regfil_3__0_), .Y(_abc_41356_new_n5502_));
OR2X2 OR2X2_1827 ( .A(regfil_5__0_), .B(sp_0_), .Y(_abc_41356_new_n5505_));
OR2X2 OR2X2_1828 ( .A(regfil_3__0_), .B(regfil_5__0_), .Y(_abc_41356_new_n5509_));
OR2X2 OR2X2_1829 ( .A(regfil_1__0_), .B(regfil_5__0_), .Y(_abc_41356_new_n5512_));
OR2X2 OR2X2_183 ( .A(_abc_41356_new_n1086_), .B(_abc_41356_new_n1084_), .Y(_abc_41356_new_n1087_));
OR2X2 OR2X2_1830 ( .A(_abc_41356_new_n5511_), .B(_abc_41356_new_n5514_), .Y(_abc_41356_new_n5515_));
OR2X2 OR2X2_1831 ( .A(_abc_41356_new_n5515_), .B(_abc_41356_new_n5507_), .Y(_abc_41356_new_n5516_));
OR2X2 OR2X2_1832 ( .A(_abc_41356_new_n5517_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n5518_));
OR2X2 OR2X2_1833 ( .A(_abc_41356_new_n5518_), .B(_abc_41356_new_n5516_), .Y(_abc_41356_new_n5519_));
OR2X2 OR2X2_1834 ( .A(_abc_41356_new_n5520_), .B(_abc_41356_new_n5501_), .Y(_abc_41356_new_n5521_));
OR2X2 OR2X2_1835 ( .A(_abc_41356_new_n5500_), .B(_abc_41356_new_n5521_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_0_));
OR2X2 OR2X2_1836 ( .A(_abc_41356_new_n771_), .B(_abc_41356_new_n5496_), .Y(_abc_41356_new_n5524_));
OR2X2 OR2X2_1837 ( .A(_abc_41356_new_n5495_), .B(regfil_5__1_), .Y(_abc_41356_new_n5525_));
OR2X2 OR2X2_1838 ( .A(_abc_41356_new_n1236_), .B(regfil_3__1_), .Y(_abc_41356_new_n5528_));
OR2X2 OR2X2_1839 ( .A(_abc_41356_new_n1260_), .B(_abc_41356_new_n1273_), .Y(_abc_41356_new_n5529_));
OR2X2 OR2X2_184 ( .A(_abc_41356_new_n1089_), .B(_abc_41356_new_n1075_), .Y(_abc_41356_new_n1090_));
OR2X2 OR2X2_1840 ( .A(_abc_41356_new_n5530_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n5531_));
OR2X2 OR2X2_1841 ( .A(_abc_41356_new_n1291_), .B(_abc_41356_new_n1292_), .Y(_abc_41356_new_n5532_));
OR2X2 OR2X2_1842 ( .A(_abc_41356_new_n5534_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n5535_));
OR2X2 OR2X2_1843 ( .A(_abc_41356_new_n5538_), .B(_abc_41356_new_n1421_), .Y(_abc_41356_new_n5539_));
OR2X2 OR2X2_1844 ( .A(_abc_41356_new_n1367_), .B(_abc_41356_new_n1364_), .Y(_abc_41356_new_n5543_));
OR2X2 OR2X2_1845 ( .A(_abc_41356_new_n5541_), .B(_abc_41356_new_n5545_), .Y(_abc_41356_new_n5546_));
OR2X2 OR2X2_1846 ( .A(_abc_41356_new_n5546_), .B(_abc_41356_new_n5536_), .Y(_abc_41356_new_n5547_));
OR2X2 OR2X2_1847 ( .A(_abc_41356_new_n5547_), .B(_abc_41356_new_n5535_), .Y(_abc_41356_new_n5548_));
OR2X2 OR2X2_1848 ( .A(_abc_41356_new_n5552_), .B(_abc_41356_new_n5531_), .Y(_abc_41356_new_n5553_));
OR2X2 OR2X2_1849 ( .A(_abc_41356_new_n5527_), .B(_abc_41356_new_n5554_), .Y(_abc_41356_new_n5555_));
OR2X2 OR2X2_185 ( .A(_abc_41356_new_n1090_), .B(_abc_41356_new_n1052_), .Y(_abc_41356_new_n1091_));
OR2X2 OR2X2_1850 ( .A(_abc_41356_new_n5555_), .B(_abc_41356_new_n5523_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_1_));
OR2X2 OR2X2_1851 ( .A(_abc_41356_new_n5558_), .B(_abc_41356_new_n5557_), .Y(_abc_41356_new_n5559_));
OR2X2 OR2X2_1852 ( .A(_abc_41356_new_n1236_), .B(regfil_3__2_), .Y(_abc_41356_new_n5562_));
OR2X2 OR2X2_1853 ( .A(_abc_41356_new_n1260_), .B(_abc_41356_new_n1257_), .Y(_abc_41356_new_n5564_));
OR2X2 OR2X2_1854 ( .A(_abc_41356_new_n5569_), .B(_abc_41356_new_n1274_), .Y(_abc_41356_new_n5570_));
OR2X2 OR2X2_1855 ( .A(_abc_41356_new_n1296_), .B(_abc_41356_new_n1301_), .Y(_abc_41356_new_n5575_));
OR2X2 OR2X2_1856 ( .A(_abc_41356_new_n5578_), .B(_abc_41356_new_n1434_), .Y(_abc_41356_new_n5579_));
OR2X2 OR2X2_1857 ( .A(_abc_41356_new_n1369_), .B(_abc_41356_new_n1373_), .Y(_abc_41356_new_n5586_));
OR2X2 OR2X2_1858 ( .A(_abc_41356_new_n5588_), .B(_abc_41356_new_n1418_), .Y(_abc_41356_new_n5589_));
OR2X2 OR2X2_1859 ( .A(_abc_41356_new_n5589_), .B(_abc_41356_new_n5583_), .Y(_abc_41356_new_n5590_));
OR2X2 OR2X2_186 ( .A(_abc_41356_new_n1094_), .B(_abc_41356_new_n723_), .Y(_abc_41356_new_n1095_));
OR2X2 OR2X2_1860 ( .A(_abc_41356_new_n5593_), .B(_abc_41356_new_n5577_), .Y(_abc_41356_new_n5594_));
OR2X2 OR2X2_1861 ( .A(_abc_41356_new_n5594_), .B(_abc_41356_new_n1285_), .Y(_abc_41356_new_n5595_));
OR2X2 OR2X2_1862 ( .A(_abc_41356_new_n5597_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n5598_));
OR2X2 OR2X2_1863 ( .A(_abc_41356_new_n5599_), .B(_abc_41356_new_n5561_), .Y(_abc_41356_new_n5600_));
OR2X2 OR2X2_1864 ( .A(_abc_41356_new_n5600_), .B(_abc_41356_new_n5560_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_2_));
OR2X2 OR2X2_1865 ( .A(_abc_41356_new_n885_), .B(_abc_41356_new_n5496_), .Y(_abc_41356_new_n5602_));
OR2X2 OR2X2_1866 ( .A(_abc_41356_new_n5495_), .B(regfil_5__3_), .Y(_abc_41356_new_n5603_));
OR2X2 OR2X2_1867 ( .A(_abc_41356_new_n1236_), .B(regfil_3__3_), .Y(_abc_41356_new_n5607_));
OR2X2 OR2X2_1868 ( .A(_abc_41356_new_n5608_), .B(_abc_41356_new_n1262_), .Y(_abc_41356_new_n5609_));
OR2X2 OR2X2_1869 ( .A(_abc_41356_new_n5610_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n5611_));
OR2X2 OR2X2_187 ( .A(_abc_41356_new_n1093_), .B(_abc_41356_new_n1095_), .Y(_abc_41356_new_n1096_));
OR2X2 OR2X2_1870 ( .A(_abc_41356_new_n5614_), .B(_abc_41356_new_n1306_), .Y(_abc_41356_new_n5615_));
OR2X2 OR2X2_1871 ( .A(_abc_41356_new_n5613_), .B(_abc_41356_new_n1305_), .Y(_abc_41356_new_n5616_));
OR2X2 OR2X2_1872 ( .A(_abc_41356_new_n5618_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n5619_));
OR2X2 OR2X2_1873 ( .A(_abc_41356_new_n5623_), .B(_abc_41356_new_n1430_), .Y(_abc_41356_new_n5624_));
OR2X2 OR2X2_1874 ( .A(_abc_41356_new_n5622_), .B(_abc_41356_new_n1429_), .Y(_abc_41356_new_n5626_));
OR2X2 OR2X2_1875 ( .A(_abc_41356_new_n5630_), .B(_abc_41356_new_n1358_), .Y(_abc_41356_new_n5631_));
OR2X2 OR2X2_1876 ( .A(_abc_41356_new_n5632_), .B(_abc_41356_new_n1359_), .Y(_abc_41356_new_n5633_));
OR2X2 OR2X2_1877 ( .A(_abc_41356_new_n5628_), .B(_abc_41356_new_n5635_), .Y(_abc_41356_new_n5636_));
OR2X2 OR2X2_1878 ( .A(_abc_41356_new_n5636_), .B(_abc_41356_new_n5620_), .Y(_abc_41356_new_n5637_));
OR2X2 OR2X2_1879 ( .A(_abc_41356_new_n5637_), .B(_abc_41356_new_n5619_), .Y(_abc_41356_new_n5638_));
OR2X2 OR2X2_188 ( .A(_abc_41356_new_n1100_), .B(_abc_41356_new_n555_), .Y(_abc_41356_new_n1101_));
OR2X2 OR2X2_1880 ( .A(_abc_41356_new_n5640_), .B(_abc_41356_new_n1275_), .Y(_abc_41356_new_n5641_));
OR2X2 OR2X2_1881 ( .A(_abc_41356_new_n5644_), .B(_abc_41356_new_n5611_), .Y(_abc_41356_new_n5645_));
OR2X2 OR2X2_1882 ( .A(_abc_41356_new_n5646_), .B(_abc_41356_new_n5606_), .Y(_abc_41356_new_n5647_));
OR2X2 OR2X2_1883 ( .A(_abc_41356_new_n5647_), .B(_abc_41356_new_n5605_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_3_));
OR2X2 OR2X2_1884 ( .A(_abc_41356_new_n952_), .B(_abc_41356_new_n5496_), .Y(_abc_41356_new_n5649_));
OR2X2 OR2X2_1885 ( .A(_abc_41356_new_n5495_), .B(regfil_5__4_), .Y(_abc_41356_new_n5650_));
OR2X2 OR2X2_1886 ( .A(_abc_41356_new_n1236_), .B(regfil_3__4_), .Y(_abc_41356_new_n5654_));
OR2X2 OR2X2_1887 ( .A(_abc_41356_new_n5656_), .B(_abc_41356_new_n1263_), .Y(_abc_41356_new_n5657_));
OR2X2 OR2X2_1888 ( .A(_abc_41356_new_n5658_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n5659_));
OR2X2 OR2X2_1889 ( .A(_abc_41356_new_n1376_), .B(_abc_41356_new_n1393_), .Y(_abc_41356_new_n5660_));
OR2X2 OR2X2_189 ( .A(_abc_41356_new_n1111_), .B(_abc_41356_new_n1112_), .Y(_abc_41356_new_n1113_));
OR2X2 OR2X2_1890 ( .A(_abc_41356_new_n5665_), .B(_abc_41356_new_n1455_), .Y(_abc_41356_new_n5668_));
OR2X2 OR2X2_1891 ( .A(_abc_41356_new_n5670_), .B(_abc_41356_new_n1418_), .Y(_abc_41356_new_n5671_));
OR2X2 OR2X2_1892 ( .A(_abc_41356_new_n5671_), .B(_abc_41356_new_n5664_), .Y(_abc_41356_new_n5672_));
OR2X2 OR2X2_1893 ( .A(_abc_41356_new_n1311_), .B(_abc_41356_new_n1328_), .Y(_abc_41356_new_n5678_));
OR2X2 OR2X2_1894 ( .A(_abc_41356_new_n5680_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n5681_));
OR2X2 OR2X2_1895 ( .A(_abc_41356_new_n5675_), .B(_abc_41356_new_n5681_), .Y(_abc_41356_new_n5682_));
OR2X2 OR2X2_1896 ( .A(_abc_41356_new_n5684_), .B(_abc_41356_new_n1795_), .Y(_abc_41356_new_n5685_));
OR2X2 OR2X2_1897 ( .A(_abc_41356_new_n5688_), .B(_abc_41356_new_n5659_), .Y(_abc_41356_new_n5689_));
OR2X2 OR2X2_1898 ( .A(_abc_41356_new_n5690_), .B(_abc_41356_new_n5653_), .Y(_abc_41356_new_n5691_));
OR2X2 OR2X2_1899 ( .A(_abc_41356_new_n5691_), .B(_abc_41356_new_n5652_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_4_));
OR2X2 OR2X2_19 ( .A(_abc_41356_new_n585_), .B(_abc_41356_new_n640_), .Y(_abc_41356_new_n641_));
OR2X2 OR2X2_190 ( .A(_abc_41356_new_n1114_), .B(_abc_41356_new_n1102_), .Y(_abc_41356_new_n1115_));
OR2X2 OR2X2_1900 ( .A(_abc_41356_new_n1019_), .B(_abc_41356_new_n5496_), .Y(_abc_41356_new_n5693_));
OR2X2 OR2X2_1901 ( .A(_abc_41356_new_n5495_), .B(regfil_5__5_), .Y(_abc_41356_new_n5694_));
OR2X2 OR2X2_1902 ( .A(_abc_41356_new_n1236_), .B(regfil_3__5_), .Y(_abc_41356_new_n5698_));
OR2X2 OR2X2_1903 ( .A(_abc_41356_new_n5700_), .B(_abc_41356_new_n1264_), .Y(_abc_41356_new_n5701_));
OR2X2 OR2X2_1904 ( .A(_abc_41356_new_n5702_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n5703_));
OR2X2 OR2X2_1905 ( .A(_abc_41356_new_n5705_), .B(_abc_41356_new_n5706_), .Y(_abc_41356_new_n5707_));
OR2X2 OR2X2_1906 ( .A(_abc_41356_new_n5708_), .B(_abc_41356_new_n1334_), .Y(_abc_41356_new_n5709_));
OR2X2 OR2X2_1907 ( .A(_abc_41356_new_n5711_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n5712_));
OR2X2 OR2X2_1908 ( .A(_abc_41356_new_n5714_), .B(_abc_41356_new_n1389_), .Y(_abc_41356_new_n5715_));
OR2X2 OR2X2_1909 ( .A(_abc_41356_new_n5713_), .B(_abc_41356_new_n5716_), .Y(_abc_41356_new_n5717_));
OR2X2 OR2X2_191 ( .A(_abc_41356_new_n1116_), .B(_abc_41356_new_n1118_), .Y(_abc_41356_new_n1119_));
OR2X2 OR2X2_1910 ( .A(_abc_41356_new_n5718_), .B(_abc_41356_new_n1665_), .Y(_abc_41356_new_n5719_));
OR2X2 OR2X2_1911 ( .A(_abc_41356_new_n5721_), .B(_abc_41356_new_n1459_), .Y(_abc_41356_new_n5722_));
OR2X2 OR2X2_1912 ( .A(_abc_41356_new_n5720_), .B(_abc_41356_new_n5723_), .Y(_abc_41356_new_n5724_));
OR2X2 OR2X2_1913 ( .A(_abc_41356_new_n5726_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n5727_));
OR2X2 OR2X2_1914 ( .A(_abc_41356_new_n5728_), .B(_abc_41356_new_n5729_), .Y(_abc_41356_new_n5730_));
OR2X2 OR2X2_1915 ( .A(_abc_41356_new_n5730_), .B(_abc_41356_new_n5712_), .Y(_abc_41356_new_n5731_));
OR2X2 OR2X2_1916 ( .A(_abc_41356_new_n1795_), .B(regfil_5__5_), .Y(_abc_41356_new_n5733_));
OR2X2 OR2X2_1917 ( .A(_abc_41356_new_n5734_), .B(_abc_41356_new_n1220_), .Y(_abc_41356_new_n5735_));
OR2X2 OR2X2_1918 ( .A(_abc_41356_new_n5737_), .B(_abc_41356_new_n5703_), .Y(_abc_41356_new_n5738_));
OR2X2 OR2X2_1919 ( .A(_abc_41356_new_n5739_), .B(_abc_41356_new_n5697_), .Y(_abc_41356_new_n5740_));
OR2X2 OR2X2_192 ( .A(_abc_41356_new_n1120_), .B(_abc_41356_new_n1098_), .Y(_abc_41356_new_n1121_));
OR2X2 OR2X2_1920 ( .A(_abc_41356_new_n5740_), .B(_abc_41356_new_n5696_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_5_));
OR2X2 OR2X2_1921 ( .A(_abc_41356_new_n1091_), .B(_abc_41356_new_n5496_), .Y(_abc_41356_new_n5743_));
OR2X2 OR2X2_1922 ( .A(_abc_41356_new_n5495_), .B(regfil_5__6_), .Y(_abc_41356_new_n5744_));
OR2X2 OR2X2_1923 ( .A(_abc_41356_new_n1236_), .B(regfil_3__6_), .Y(_abc_41356_new_n5747_));
OR2X2 OR2X2_1924 ( .A(_abc_41356_new_n5749_), .B(_abc_41356_new_n1265_), .Y(_abc_41356_new_n5750_));
OR2X2 OR2X2_1925 ( .A(_abc_41356_new_n5751_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n5752_));
OR2X2 OR2X2_1926 ( .A(_abc_41356_new_n5753_), .B(_abc_41356_new_n1398_), .Y(_abc_41356_new_n5754_));
OR2X2 OR2X2_1927 ( .A(_abc_41356_new_n5754_), .B(_abc_41356_new_n1384_), .Y(_abc_41356_new_n5757_));
OR2X2 OR2X2_1928 ( .A(_abc_41356_new_n5760_), .B(_abc_41356_new_n1465_), .Y(_abc_41356_new_n5761_));
OR2X2 OR2X2_1929 ( .A(_abc_41356_new_n5761_), .B(_abc_41356_new_n1450_), .Y(_abc_41356_new_n5762_));
OR2X2 OR2X2_193 ( .A(_abc_41356_new_n702_), .B(_abc_41356_new_n1106_), .Y(_abc_41356_new_n1122_));
OR2X2 OR2X2_1930 ( .A(_abc_41356_new_n5766_), .B(_abc_41356_new_n1418_), .Y(_abc_41356_new_n5767_));
OR2X2 OR2X2_1931 ( .A(_abc_41356_new_n5767_), .B(_abc_41356_new_n5759_), .Y(_abc_41356_new_n5768_));
OR2X2 OR2X2_1932 ( .A(_abc_41356_new_n5772_), .B(_abc_41356_new_n1341_), .Y(_abc_41356_new_n5773_));
OR2X2 OR2X2_1933 ( .A(_abc_41356_new_n5773_), .B(_abc_41356_new_n1322_), .Y(_abc_41356_new_n5774_));
OR2X2 OR2X2_1934 ( .A(_abc_41356_new_n5778_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n5779_));
OR2X2 OR2X2_1935 ( .A(_abc_41356_new_n5771_), .B(_abc_41356_new_n5779_), .Y(_abc_41356_new_n5780_));
OR2X2 OR2X2_1936 ( .A(_abc_41356_new_n1796_), .B(regfil_5__6_), .Y(_abc_41356_new_n5782_));
OR2X2 OR2X2_1937 ( .A(_abc_41356_new_n5783_), .B(_abc_41356_new_n1220_), .Y(_abc_41356_new_n5784_));
OR2X2 OR2X2_1938 ( .A(_abc_41356_new_n5785_), .B(_abc_41356_new_n5752_), .Y(_abc_41356_new_n5786_));
OR2X2 OR2X2_1939 ( .A(_abc_41356_new_n5746_), .B(_abc_41356_new_n5787_), .Y(_abc_41356_new_n5788_));
OR2X2 OR2X2_194 ( .A(_abc_41356_new_n975_), .B(_abc_41356_new_n1125_), .Y(_abc_41356_new_n1126_));
OR2X2 OR2X2_1940 ( .A(_abc_41356_new_n5788_), .B(_abc_41356_new_n5742_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_6_));
OR2X2 OR2X2_1941 ( .A(_abc_41356_new_n5791_), .B(_abc_41356_new_n5790_), .Y(_abc_41356_new_n5792_));
OR2X2 OR2X2_1942 ( .A(_abc_41356_new_n5793_), .B(_abc_41356_new_n5794_), .Y(_abc_41356_new_n5795_));
OR2X2 OR2X2_1943 ( .A(_abc_41356_new_n1236_), .B(regfil_3__7_), .Y(_abc_41356_new_n5796_));
OR2X2 OR2X2_1944 ( .A(_abc_41356_new_n5799_), .B(_abc_41356_new_n1266_), .Y(_abc_41356_new_n5800_));
OR2X2 OR2X2_1945 ( .A(_abc_41356_new_n5801_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n5802_));
OR2X2 OR2X2_1946 ( .A(_abc_41356_new_n5775_), .B(_abc_41356_new_n1318_), .Y(_abc_41356_new_n5803_));
OR2X2 OR2X2_1947 ( .A(_abc_41356_new_n5803_), .B(_abc_41356_new_n1317_), .Y(_abc_41356_new_n5804_));
OR2X2 OR2X2_1948 ( .A(_abc_41356_new_n5806_), .B(_abc_41356_new_n5805_), .Y(_abc_41356_new_n5807_));
OR2X2 OR2X2_1949 ( .A(_abc_41356_new_n5809_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n5810_));
OR2X2 OR2X2_195 ( .A(_abc_41356_new_n1078_), .B(_abc_41356_new_n1134_), .Y(_abc_41356_new_n1135_));
OR2X2 OR2X2_1950 ( .A(_abc_41356_new_n5813_), .B(_abc_41356_new_n1446_), .Y(_abc_41356_new_n5814_));
OR2X2 OR2X2_1951 ( .A(_abc_41356_new_n5812_), .B(_abc_41356_new_n5815_), .Y(_abc_41356_new_n5816_));
OR2X2 OR2X2_1952 ( .A(_abc_41356_new_n5818_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n5819_));
OR2X2 OR2X2_1953 ( .A(_abc_41356_new_n5824_), .B(_abc_41356_new_n5821_), .Y(_abc_41356_new_n5825_));
OR2X2 OR2X2_1954 ( .A(_abc_41356_new_n5825_), .B(_abc_41356_new_n1665_), .Y(_abc_41356_new_n5826_));
OR2X2 OR2X2_1955 ( .A(_abc_41356_new_n5827_), .B(_abc_41356_new_n5811_), .Y(_abc_41356_new_n5828_));
OR2X2 OR2X2_1956 ( .A(_abc_41356_new_n5828_), .B(_abc_41356_new_n5810_), .Y(_abc_41356_new_n5829_));
OR2X2 OR2X2_1957 ( .A(_abc_41356_new_n1797_), .B(regfil_5__7_), .Y(_abc_41356_new_n5831_));
OR2X2 OR2X2_1958 ( .A(_abc_41356_new_n5832_), .B(_abc_41356_new_n1220_), .Y(_abc_41356_new_n5833_));
OR2X2 OR2X2_1959 ( .A(_abc_41356_new_n5834_), .B(_abc_41356_new_n5802_), .Y(_abc_41356_new_n5835_));
OR2X2 OR2X2_196 ( .A(_abc_41356_new_n1138_), .B(_abc_41356_new_n597_), .Y(_abc_41356_new_n1139_));
OR2X2 OR2X2_1960 ( .A(_abc_41356_new_n5795_), .B(_abc_41356_new_n5836_), .Y(_abc_36060_memoryregfil_wrmux_5__3__0__y_16171_7_));
OR2X2 OR2X2_1961 ( .A(_abc_41356_new_n5838_), .B(_abc_41356_new_n5839_), .Y(_abc_41356_new_n5840_));
OR2X2 OR2X2_1962 ( .A(_abc_41356_new_n5846_), .B(reset), .Y(_abc_41356_new_n5847_));
OR2X2 OR2X2_1963 ( .A(_abc_41356_new_n5851_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n5852_));
OR2X2 OR2X2_1964 ( .A(_abc_41356_new_n5858_), .B(sp_0_), .Y(_abc_41356_new_n5859_));
OR2X2 OR2X2_1965 ( .A(_abc_41356_new_n5860_), .B(_abc_41356_new_n5850_), .Y(_abc_41356_new_n5861_));
OR2X2 OR2X2_1966 ( .A(_abc_41356_new_n5868_), .B(_abc_41356_new_n5867_), .Y(_abc_41356_new_n5869_));
OR2X2 OR2X2_1967 ( .A(_abc_41356_new_n5866_), .B(_abc_41356_new_n5869_), .Y(_abc_41356_new_n5870_));
OR2X2 OR2X2_1968 ( .A(_abc_41356_new_n5871_), .B(_abc_41356_new_n5848_), .Y(_0sp_15_0__0_));
OR2X2 OR2X2_1969 ( .A(_abc_41356_new_n5877_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n5878_));
OR2X2 OR2X2_197 ( .A(_abc_41356_new_n1142_), .B(_abc_41356_new_n1141_), .Y(_abc_41356_new_n1143_));
OR2X2 OR2X2_1970 ( .A(_abc_41356_new_n5879_), .B(_abc_41356_new_n5878_), .Y(_abc_41356_new_n5880_));
OR2X2 OR2X2_1971 ( .A(_abc_41356_new_n5880_), .B(_abc_41356_new_n5876_), .Y(_abc_41356_new_n5881_));
OR2X2 OR2X2_1972 ( .A(_abc_41356_new_n5882_), .B(_abc_41356_new_n5888_), .Y(_abc_41356_new_n5889_));
OR2X2 OR2X2_1973 ( .A(_abc_41356_new_n5854_), .B(_abc_41356_new_n4857_), .Y(_abc_41356_new_n5893_));
OR2X2 OR2X2_1974 ( .A(_abc_41356_new_n5853_), .B(sp_1_), .Y(_abc_41356_new_n5898_));
OR2X2 OR2X2_1975 ( .A(_abc_41356_new_n5903_), .B(_abc_41356_new_n5902_), .Y(_abc_41356_new_n5904_));
OR2X2 OR2X2_1976 ( .A(_abc_41356_new_n5901_), .B(_abc_41356_new_n5904_), .Y(_abc_41356_new_n5905_));
OR2X2 OR2X2_1977 ( .A(_abc_41356_new_n5906_), .B(_abc_41356_new_n5873_), .Y(_0sp_15_0__1_));
OR2X2 OR2X2_1978 ( .A(_abc_41356_new_n5913_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n5914_));
OR2X2 OR2X2_1979 ( .A(_abc_41356_new_n5914_), .B(_abc_41356_new_n5911_), .Y(_abc_41356_new_n5915_));
OR2X2 OR2X2_198 ( .A(_abc_41356_new_n1146_), .B(_abc_41356_new_n1145_), .Y(_abc_41356_new_n1147_));
OR2X2 OR2X2_1980 ( .A(_abc_41356_new_n5910_), .B(_abc_41356_new_n5915_), .Y(_abc_41356_new_n5916_));
OR2X2 OR2X2_1981 ( .A(_abc_41356_new_n5916_), .B(_abc_41356_new_n5909_), .Y(_abc_41356_new_n5917_));
OR2X2 OR2X2_1982 ( .A(_abc_41356_new_n5886_), .B(sp_2_), .Y(_abc_41356_new_n5918_));
OR2X2 OR2X2_1983 ( .A(_abc_41356_new_n5919_), .B(_abc_41356_new_n5922_), .Y(_abc_41356_new_n5923_));
OR2X2 OR2X2_1984 ( .A(_abc_41356_new_n5926_), .B(_abc_41356_new_n5925_), .Y(_abc_41356_new_n5927_));
OR2X2 OR2X2_1985 ( .A(_abc_41356_new_n5928_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n5929_));
OR2X2 OR2X2_1986 ( .A(_abc_41356_new_n5924_), .B(_abc_41356_new_n5929_), .Y(_abc_41356_new_n5930_));
OR2X2 OR2X2_1987 ( .A(_abc_41356_new_n5853_), .B(sp_2_), .Y(_abc_41356_new_n5931_));
OR2X2 OR2X2_1988 ( .A(_abc_41356_new_n5937_), .B(_abc_41356_new_n5936_), .Y(_abc_41356_new_n5938_));
OR2X2 OR2X2_1989 ( .A(_abc_41356_new_n5938_), .B(_abc_41356_new_n5935_), .Y(_abc_41356_new_n5939_));
OR2X2 OR2X2_199 ( .A(_abc_41356_new_n1149_), .B(_abc_41356_new_n1148_), .Y(_abc_41356_new_n1150_));
OR2X2 OR2X2_1990 ( .A(_abc_41356_new_n5934_), .B(_abc_41356_new_n5939_), .Y(_abc_41356_new_n5940_));
OR2X2 OR2X2_1991 ( .A(_abc_41356_new_n5941_), .B(_abc_41356_new_n5908_), .Y(_0sp_15_0__2_));
OR2X2 OR2X2_1992 ( .A(_abc_41356_new_n4895_), .B(sp_3_), .Y(_abc_41356_new_n5948_));
OR2X2 OR2X2_1993 ( .A(_abc_41356_new_n5951_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n5952_));
OR2X2 OR2X2_1994 ( .A(_abc_41356_new_n5952_), .B(_abc_41356_new_n5950_), .Y(_abc_41356_new_n5953_));
OR2X2 OR2X2_1995 ( .A(_abc_41356_new_n5945_), .B(_abc_41356_new_n5953_), .Y(_abc_41356_new_n5954_));
OR2X2 OR2X2_1996 ( .A(_abc_41356_new_n5954_), .B(_abc_41356_new_n5944_), .Y(_abc_41356_new_n5955_));
OR2X2 OR2X2_1997 ( .A(_abc_41356_new_n4931_), .B(sp_0_), .Y(_abc_41356_new_n5956_));
OR2X2 OR2X2_1998 ( .A(_abc_41356_new_n5925_), .B(sp_3_), .Y(_abc_41356_new_n5957_));
OR2X2 OR2X2_1999 ( .A(_abc_41356_new_n5960_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n5961_));
OR2X2 OR2X2_2 ( .A(_abc_41356_new_n543_), .B(auxcar), .Y(_abc_41356_new_n544_));
OR2X2 OR2X2_20 ( .A(_abc_41356_new_n595_), .B(_abc_41356_new_n608_), .Y(_abc_41356_new_n642_));
OR2X2 OR2X2_200 ( .A(_abc_41356_new_n1147_), .B(_abc_41356_new_n1150_), .Y(_abc_41356_new_n1151_));
OR2X2 OR2X2_2000 ( .A(_abc_41356_new_n5920_), .B(sp_3_), .Y(_abc_41356_new_n5964_));
OR2X2 OR2X2_2001 ( .A(_abc_41356_new_n5961_), .B(_abc_41356_new_n5966_), .Y(_abc_41356_new_n5967_));
OR2X2 OR2X2_2002 ( .A(_abc_41356_new_n5967_), .B(_abc_41356_new_n5959_), .Y(_abc_41356_new_n5968_));
OR2X2 OR2X2_2003 ( .A(_abc_41356_new_n5853_), .B(sp_3_), .Y(_abc_41356_new_n5969_));
OR2X2 OR2X2_2004 ( .A(_abc_41356_new_n5974_), .B(_abc_41356_new_n5975_), .Y(_abc_41356_new_n5976_));
OR2X2 OR2X2_2005 ( .A(_abc_41356_new_n5976_), .B(_abc_41356_new_n5973_), .Y(_abc_41356_new_n5977_));
OR2X2 OR2X2_2006 ( .A(_abc_41356_new_n5972_), .B(_abc_41356_new_n5977_), .Y(_abc_41356_new_n5978_));
OR2X2 OR2X2_2007 ( .A(_abc_41356_new_n5979_), .B(_abc_41356_new_n5943_), .Y(_0sp_15_0__3_));
OR2X2 OR2X2_2008 ( .A(_abc_41356_new_n5946_), .B(sp_4_), .Y(_abc_41356_new_n5986_));
OR2X2 OR2X2_2009 ( .A(_abc_41356_new_n5989_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n5990_));
OR2X2 OR2X2_201 ( .A(_abc_41356_new_n1151_), .B(opcode_2_), .Y(_abc_41356_new_n1152_));
OR2X2 OR2X2_2010 ( .A(_abc_41356_new_n5990_), .B(_abc_41356_new_n5988_), .Y(_abc_41356_new_n5991_));
OR2X2 OR2X2_2011 ( .A(_abc_41356_new_n5983_), .B(_abc_41356_new_n5991_), .Y(_abc_41356_new_n5992_));
OR2X2 OR2X2_2012 ( .A(_abc_41356_new_n5992_), .B(_abc_41356_new_n5982_), .Y(_abc_41356_new_n5993_));
OR2X2 OR2X2_2013 ( .A(_abc_41356_new_n5998_), .B(_abc_41356_new_n5996_), .Y(_abc_41356_new_n5999_));
OR2X2 OR2X2_2014 ( .A(_abc_41356_new_n6000_), .B(_abc_41356_new_n5994_), .Y(_abc_41356_new_n6001_));
OR2X2 OR2X2_2015 ( .A(_abc_41356_new_n5962_), .B(sp_4_), .Y(_abc_41356_new_n6004_));
OR2X2 OR2X2_2016 ( .A(_abc_41356_new_n6006_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6007_));
OR2X2 OR2X2_2017 ( .A(_abc_41356_new_n6001_), .B(_abc_41356_new_n6007_), .Y(_abc_41356_new_n6008_));
OR2X2 OR2X2_2018 ( .A(_abc_41356_new_n5853_), .B(sp_4_), .Y(_abc_41356_new_n6009_));
OR2X2 OR2X2_2019 ( .A(_abc_41356_new_n6013_), .B(_abc_41356_new_n6014_), .Y(_abc_41356_new_n6015_));
OR2X2 OR2X2_202 ( .A(_abc_41356_new_n1153_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n1154_));
OR2X2 OR2X2_2020 ( .A(_abc_41356_new_n6015_), .B(_abc_41356_new_n6016_), .Y(_abc_41356_new_n6017_));
OR2X2 OR2X2_2021 ( .A(_abc_41356_new_n6012_), .B(_abc_41356_new_n6017_), .Y(_abc_41356_new_n6018_));
OR2X2 OR2X2_2022 ( .A(_abc_41356_new_n6019_), .B(_abc_41356_new_n5981_), .Y(_0sp_15_0__4_));
OR2X2 OR2X2_2023 ( .A(_abc_41356_new_n5875_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6022_));
OR2X2 OR2X2_2024 ( .A(_abc_41356_new_n6023_), .B(_abc_41356_new_n5856_), .Y(_abc_41356_new_n6024_));
OR2X2 OR2X2_2025 ( .A(_abc_41356_new_n5984_), .B(sp_5_), .Y(_abc_41356_new_n6029_));
OR2X2 OR2X2_2026 ( .A(_abc_41356_new_n6031_), .B(_abc_41356_new_n6032_), .Y(_abc_41356_new_n6033_));
OR2X2 OR2X2_2027 ( .A(_abc_41356_new_n6026_), .B(_abc_41356_new_n6033_), .Y(_abc_41356_new_n6034_));
OR2X2 OR2X2_2028 ( .A(_abc_41356_new_n6002_), .B(sp_5_), .Y(_abc_41356_new_n6038_));
OR2X2 OR2X2_2029 ( .A(_abc_41356_new_n6041_), .B(_abc_41356_new_n1331_), .Y(_abc_41356_new_n6042_));
OR2X2 OR2X2_203 ( .A(_abc_41356_new_n1156_), .B(_abc_41356_new_n1157_), .Y(_abc_41356_new_n1158_));
OR2X2 OR2X2_2030 ( .A(_abc_41356_new_n5996_), .B(sp_5_), .Y(_abc_41356_new_n6043_));
OR2X2 OR2X2_2031 ( .A(_abc_41356_new_n6045_), .B(_abc_41356_new_n6040_), .Y(_abc_41356_new_n6046_));
OR2X2 OR2X2_2032 ( .A(_abc_41356_new_n6035_), .B(_abc_41356_new_n6047_), .Y(_abc_41356_new_n6048_));
OR2X2 OR2X2_2033 ( .A(_abc_41356_new_n6025_), .B(_abc_41356_new_n6048_), .Y(_abc_41356_new_n6049_));
OR2X2 OR2X2_2034 ( .A(_abc_41356_new_n6052_), .B(_abc_41356_new_n6053_), .Y(_abc_41356_new_n6054_));
OR2X2 OR2X2_2035 ( .A(_abc_41356_new_n6054_), .B(_abc_41356_new_n6051_), .Y(_abc_41356_new_n6055_));
OR2X2 OR2X2_2036 ( .A(_abc_41356_new_n6050_), .B(_abc_41356_new_n6055_), .Y(_abc_41356_new_n6056_));
OR2X2 OR2X2_2037 ( .A(_abc_41356_new_n6057_), .B(_abc_41356_new_n6021_), .Y(_0sp_15_0__5_));
OR2X2 OR2X2_2038 ( .A(_abc_41356_new_n5043_), .B(sp_0_), .Y(_abc_41356_new_n6062_));
OR2X2 OR2X2_2039 ( .A(_abc_41356_new_n6063_), .B(_abc_41356_new_n6061_), .Y(_abc_41356_new_n6064_));
OR2X2 OR2X2_204 ( .A(_abc_41356_new_n1158_), .B(_abc_41356_new_n1155_), .Y(_abc_41356_new_n1159_));
OR2X2 OR2X2_2040 ( .A(_abc_41356_new_n6036_), .B(sp_6_), .Y(_abc_41356_new_n6068_));
OR2X2 OR2X2_2041 ( .A(_abc_41356_new_n6065_), .B(_abc_41356_new_n6070_), .Y(_abc_41356_new_n6071_));
OR2X2 OR2X2_2042 ( .A(_abc_41356_new_n6060_), .B(_abc_41356_new_n6072_), .Y(_abc_41356_new_n6073_));
OR2X2 OR2X2_2043 ( .A(_abc_41356_new_n6027_), .B(sp_6_), .Y(_abc_41356_new_n6077_));
OR2X2 OR2X2_2044 ( .A(_abc_41356_new_n6080_), .B(_abc_41356_new_n6081_), .Y(_abc_41356_new_n6082_));
OR2X2 OR2X2_2045 ( .A(_abc_41356_new_n6082_), .B(_abc_41356_new_n6079_), .Y(_abc_41356_new_n6083_));
OR2X2 OR2X2_2046 ( .A(_abc_41356_new_n6085_), .B(_abc_41356_new_n6086_), .Y(_abc_41356_new_n6087_));
OR2X2 OR2X2_2047 ( .A(_abc_41356_new_n6084_), .B(_abc_41356_new_n6087_), .Y(_abc_41356_new_n6088_));
OR2X2 OR2X2_2048 ( .A(_abc_41356_new_n6090_), .B(_abc_41356_new_n6083_), .Y(_abc_41356_new_n6091_));
OR2X2 OR2X2_2049 ( .A(_abc_41356_new_n6074_), .B(_abc_41356_new_n6091_), .Y(_abc_41356_new_n6092_));
OR2X2 OR2X2_205 ( .A(_abc_41356_new_n1159_), .B(_abc_41356_new_n1154_), .Y(_abc_41356_new_n1160_));
OR2X2 OR2X2_2050 ( .A(_abc_41356_new_n6093_), .B(_abc_41356_new_n6059_), .Y(_0sp_15_0__6_));
OR2X2 OR2X2_2051 ( .A(_abc_41356_new_n6075_), .B(sp_7_), .Y(_abc_41356_new_n6100_));
OR2X2 OR2X2_2052 ( .A(_abc_41356_new_n6103_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6104_));
OR2X2 OR2X2_2053 ( .A(_abc_41356_new_n6102_), .B(_abc_41356_new_n6104_), .Y(_abc_41356_new_n6105_));
OR2X2 OR2X2_2054 ( .A(_abc_41356_new_n6097_), .B(_abc_41356_new_n6105_), .Y(_abc_41356_new_n6106_));
OR2X2 OR2X2_2055 ( .A(_abc_41356_new_n6106_), .B(_abc_41356_new_n6096_), .Y(_abc_41356_new_n6107_));
OR2X2 OR2X2_2056 ( .A(_abc_41356_new_n6066_), .B(sp_7_), .Y(_abc_41356_new_n6108_));
OR2X2 OR2X2_2057 ( .A(_abc_41356_new_n6114_), .B(_abc_41356_new_n5855_), .Y(_abc_41356_new_n6115_));
OR2X2 OR2X2_2058 ( .A(_abc_41356_new_n6118_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6119_));
OR2X2 OR2X2_2059 ( .A(_abc_41356_new_n6116_), .B(_abc_41356_new_n6119_), .Y(_abc_41356_new_n6120_));
OR2X2 OR2X2_206 ( .A(_abc_41356_new_n1166_), .B(_abc_41356_new_n1165_), .Y(_abc_41356_new_n1167_));
OR2X2 OR2X2_2060 ( .A(_abc_41356_new_n6120_), .B(_abc_41356_new_n6112_), .Y(_abc_41356_new_n6121_));
OR2X2 OR2X2_2061 ( .A(_abc_41356_new_n5853_), .B(sp_7_), .Y(_abc_41356_new_n6122_));
OR2X2 OR2X2_2062 ( .A(_abc_41356_new_n6127_), .B(_abc_41356_new_n6128_), .Y(_abc_41356_new_n6129_));
OR2X2 OR2X2_2063 ( .A(_abc_41356_new_n6129_), .B(_abc_41356_new_n6126_), .Y(_abc_41356_new_n6130_));
OR2X2 OR2X2_2064 ( .A(_abc_41356_new_n6125_), .B(_abc_41356_new_n6130_), .Y(_abc_41356_new_n6131_));
OR2X2 OR2X2_2065 ( .A(_abc_41356_new_n6132_), .B(_abc_41356_new_n6095_), .Y(_0sp_15_0__7_));
OR2X2 OR2X2_2066 ( .A(_abc_41356_new_n6098_), .B(sp_8_), .Y(_abc_41356_new_n6138_));
OR2X2 OR2X2_2067 ( .A(_abc_41356_new_n6142_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6143_));
OR2X2 OR2X2_2068 ( .A(_abc_41356_new_n6141_), .B(_abc_41356_new_n6143_), .Y(_abc_41356_new_n6144_));
OR2X2 OR2X2_2069 ( .A(_abc_41356_new_n6144_), .B(_abc_41356_new_n6140_), .Y(_abc_41356_new_n6145_));
OR2X2 OR2X2_207 ( .A(_abc_41356_new_n1162_), .B(_abc_41356_new_n1167_), .Y(_abc_41356_new_n1168_));
OR2X2 OR2X2_2070 ( .A(_abc_41356_new_n6145_), .B(_abc_41356_new_n6135_), .Y(_abc_41356_new_n6146_));
OR2X2 OR2X2_2071 ( .A(_abc_41356_new_n6109_), .B(sp_8_), .Y(_abc_41356_new_n6147_));
OR2X2 OR2X2_2072 ( .A(_abc_41356_new_n6153_), .B(_abc_41356_new_n5855_), .Y(_abc_41356_new_n6154_));
OR2X2 OR2X2_2073 ( .A(_abc_41356_new_n6157_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6158_));
OR2X2 OR2X2_2074 ( .A(_abc_41356_new_n6155_), .B(_abc_41356_new_n6158_), .Y(_abc_41356_new_n6159_));
OR2X2 OR2X2_2075 ( .A(_abc_41356_new_n6159_), .B(_abc_41356_new_n6151_), .Y(_abc_41356_new_n6160_));
OR2X2 OR2X2_2076 ( .A(_abc_41356_new_n5853_), .B(sp_8_), .Y(_abc_41356_new_n6161_));
OR2X2 OR2X2_2077 ( .A(_abc_41356_new_n6166_), .B(_abc_41356_new_n6167_), .Y(_abc_41356_new_n6168_));
OR2X2 OR2X2_2078 ( .A(_abc_41356_new_n6168_), .B(_abc_41356_new_n6165_), .Y(_abc_41356_new_n6169_));
OR2X2 OR2X2_2079 ( .A(_abc_41356_new_n6164_), .B(_abc_41356_new_n6169_), .Y(_abc_41356_new_n6170_));
OR2X2 OR2X2_208 ( .A(_abc_41356_new_n1169_), .B(_abc_41356_new_n1170_), .Y(_abc_41356_new_n1171_));
OR2X2 OR2X2_2080 ( .A(_abc_41356_new_n6171_), .B(_abc_41356_new_n6134_), .Y(_0sp_15_0__8_));
OR2X2 OR2X2_2081 ( .A(_abc_41356_new_n6148_), .B(sp_9_), .Y(_abc_41356_new_n6174_));
OR2X2 OR2X2_2082 ( .A(_abc_41356_new_n6157_), .B(sp_9_), .Y(_abc_41356_new_n6179_));
OR2X2 OR2X2_2083 ( .A(_abc_41356_new_n6181_), .B(_abc_41356_new_n6183_), .Y(_abc_41356_new_n6184_));
OR2X2 OR2X2_2084 ( .A(_abc_41356_new_n6185_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6186_));
OR2X2 OR2X2_2085 ( .A(_abc_41356_new_n6186_), .B(_abc_41356_new_n6178_), .Y(_abc_41356_new_n6187_));
OR2X2 OR2X2_2086 ( .A(_abc_41356_new_n6189_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6190_));
OR2X2 OR2X2_2087 ( .A(_abc_41356_new_n6188_), .B(_abc_41356_new_n6190_), .Y(_abc_41356_new_n6191_));
OR2X2 OR2X2_2088 ( .A(_abc_41356_new_n6136_), .B(sp_9_), .Y(_abc_41356_new_n6195_));
OR2X2 OR2X2_2089 ( .A(_abc_41356_new_n6197_), .B(_abc_41356_new_n6192_), .Y(_abc_41356_new_n6198_));
OR2X2 OR2X2_209 ( .A(_abc_41356_new_n1144_), .B(_abc_41356_new_n1171_), .Y(_abc_41356_new_n1172_));
OR2X2 OR2X2_2090 ( .A(_abc_41356_new_n6191_), .B(_abc_41356_new_n6198_), .Y(_abc_41356_new_n6199_));
OR2X2 OR2X2_2091 ( .A(_abc_41356_new_n5853_), .B(sp_9_), .Y(_abc_41356_new_n6200_));
OR2X2 OR2X2_2092 ( .A(_abc_41356_new_n6205_), .B(_abc_41356_new_n6206_), .Y(_abc_41356_new_n6207_));
OR2X2 OR2X2_2093 ( .A(_abc_41356_new_n6207_), .B(_abc_41356_new_n6204_), .Y(_abc_41356_new_n6208_));
OR2X2 OR2X2_2094 ( .A(_abc_41356_new_n6203_), .B(_abc_41356_new_n6208_), .Y(_abc_41356_new_n6209_));
OR2X2 OR2X2_2095 ( .A(_abc_41356_new_n6210_), .B(_abc_41356_new_n6173_), .Y(_0sp_15_0__9_));
OR2X2 OR2X2_2096 ( .A(_abc_41356_new_n5191_), .B(sp_0_), .Y(_abc_41356_new_n6214_));
OR2X2 OR2X2_2097 ( .A(_abc_41356_new_n6215_), .B(_abc_41356_new_n6213_), .Y(_abc_41356_new_n6216_));
OR2X2 OR2X2_2098 ( .A(_abc_41356_new_n6175_), .B(sp_10_), .Y(_abc_41356_new_n6221_));
OR2X2 OR2X2_2099 ( .A(_abc_41356_new_n6217_), .B(_abc_41356_new_n6223_), .Y(_abc_41356_new_n6224_));
OR2X2 OR2X2_21 ( .A(_abc_41356_new_n652_), .B(regfil_1__4_), .Y(_abc_41356_new_n653_));
OR2X2 OR2X2_210 ( .A(_abc_41356_new_n1172_), .B(_abc_41356_new_n1140_), .Y(_abc_41356_new_n1173_));
OR2X2 OR2X2_2100 ( .A(_abc_41356_new_n6193_), .B(sp_10_), .Y(_abc_41356_new_n6228_));
OR2X2 OR2X2_2101 ( .A(_abc_41356_new_n6232_), .B(_abc_41356_new_n6231_), .Y(_abc_41356_new_n6233_));
OR2X2 OR2X2_2102 ( .A(_abc_41356_new_n6233_), .B(_abc_41356_new_n6230_), .Y(_abc_41356_new_n6234_));
OR2X2 OR2X2_2103 ( .A(_abc_41356_new_n6235_), .B(_abc_41356_new_n6226_), .Y(_abc_41356_new_n6236_));
OR2X2 OR2X2_2104 ( .A(_abc_41356_new_n6236_), .B(_abc_41356_new_n6225_), .Y(_abc_41356_new_n6237_));
OR2X2 OR2X2_2105 ( .A(_abc_41356_new_n6241_), .B(_abc_41356_new_n6240_), .Y(_abc_41356_new_n6242_));
OR2X2 OR2X2_2106 ( .A(_abc_41356_new_n6242_), .B(_abc_41356_new_n6239_), .Y(_abc_41356_new_n6243_));
OR2X2 OR2X2_2107 ( .A(_abc_41356_new_n6238_), .B(_abc_41356_new_n6243_), .Y(_abc_41356_new_n6244_));
OR2X2 OR2X2_2108 ( .A(_abc_41356_new_n6245_), .B(_abc_41356_new_n6212_), .Y(_0sp_15_0__10_));
OR2X2 OR2X2_2109 ( .A(_abc_41356_new_n6250_), .B(_abc_41356_new_n6248_), .Y(_abc_41356_new_n6251_));
OR2X2 OR2X2_211 ( .A(_abc_41356_new_n1173_), .B(_abc_41356_new_n696_), .Y(_abc_41356_new_n1174_));
OR2X2 OR2X2_2110 ( .A(_abc_41356_new_n6253_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6254_));
OR2X2 OR2X2_2111 ( .A(_abc_41356_new_n6252_), .B(_abc_41356_new_n6254_), .Y(_abc_41356_new_n6255_));
OR2X2 OR2X2_2112 ( .A(_abc_41356_new_n6219_), .B(sp_11_), .Y(_abc_41356_new_n6256_));
OR2X2 OR2X2_2113 ( .A(_abc_41356_new_n6255_), .B(_abc_41356_new_n6261_), .Y(_abc_41356_new_n6262_));
OR2X2 OR2X2_2114 ( .A(_abc_41356_new_n6218_), .B(sp_11_), .Y(_abc_41356_new_n6265_));
OR2X2 OR2X2_2115 ( .A(_abc_41356_new_n6270_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6271_));
OR2X2 OR2X2_2116 ( .A(_abc_41356_new_n6269_), .B(_abc_41356_new_n6271_), .Y(_abc_41356_new_n6272_));
OR2X2 OR2X2_2117 ( .A(_abc_41356_new_n6268_), .B(_abc_41356_new_n6272_), .Y(_abc_41356_new_n6273_));
OR2X2 OR2X2_2118 ( .A(_abc_41356_new_n6273_), .B(_abc_41356_new_n6267_), .Y(_abc_41356_new_n6274_));
OR2X2 OR2X2_2119 ( .A(_abc_41356_new_n5853_), .B(sp_11_), .Y(_abc_41356_new_n6275_));
OR2X2 OR2X2_212 ( .A(_abc_41356_new_n695_), .B(regfil_7__7_), .Y(_abc_41356_new_n1175_));
OR2X2 OR2X2_2120 ( .A(_abc_41356_new_n6280_), .B(_abc_41356_new_n6281_), .Y(_abc_41356_new_n6282_));
OR2X2 OR2X2_2121 ( .A(_abc_41356_new_n6282_), .B(_abc_41356_new_n6279_), .Y(_abc_41356_new_n6283_));
OR2X2 OR2X2_2122 ( .A(_abc_41356_new_n6278_), .B(_abc_41356_new_n6283_), .Y(_abc_41356_new_n6284_));
OR2X2 OR2X2_2123 ( .A(_abc_41356_new_n6285_), .B(_abc_41356_new_n6247_), .Y(_0sp_15_0__11_));
OR2X2 OR2X2_2124 ( .A(_abc_41356_new_n6263_), .B(sp_12_), .Y(_abc_41356_new_n6290_));
OR2X2 OR2X2_2125 ( .A(_abc_41356_new_n6294_), .B(_abc_41356_new_n6293_), .Y(_abc_41356_new_n6295_));
OR2X2 OR2X2_2126 ( .A(_abc_41356_new_n6295_), .B(_abc_41356_new_n6292_), .Y(_abc_41356_new_n6296_));
OR2X2 OR2X2_2127 ( .A(_abc_41356_new_n6300_), .B(_abc_41356_new_n6298_), .Y(_abc_41356_new_n6301_));
OR2X2 OR2X2_2128 ( .A(_abc_41356_new_n6258_), .B(sp_12_), .Y(_abc_41356_new_n6303_));
OR2X2 OR2X2_2129 ( .A(_abc_41356_new_n6302_), .B(_abc_41356_new_n6307_), .Y(_abc_41356_new_n6308_));
OR2X2 OR2X2_213 ( .A(_abc_41356_new_n703_), .B(regfil_7__7_), .Y(_abc_41356_new_n1179_));
OR2X2 OR2X2_2130 ( .A(_abc_41356_new_n6309_), .B(_abc_41356_new_n6310_), .Y(_abc_41356_new_n6311_));
OR2X2 OR2X2_2131 ( .A(_abc_41356_new_n6311_), .B(_abc_41356_new_n6297_), .Y(_abc_41356_new_n6312_));
OR2X2 OR2X2_2132 ( .A(_abc_41356_new_n6315_), .B(_abc_41356_new_n6316_), .Y(_abc_41356_new_n6317_));
OR2X2 OR2X2_2133 ( .A(_abc_41356_new_n6317_), .B(_abc_41356_new_n6314_), .Y(_abc_41356_new_n6318_));
OR2X2 OR2X2_2134 ( .A(_abc_41356_new_n6313_), .B(_abc_41356_new_n6318_), .Y(_abc_41356_new_n6319_));
OR2X2 OR2X2_2135 ( .A(_abc_41356_new_n6320_), .B(_abc_41356_new_n6287_), .Y(_0sp_15_0__12_));
OR2X2 OR2X2_2136 ( .A(_abc_41356_new_n6304_), .B(sp_13_), .Y(_abc_41356_new_n6326_));
OR2X2 OR2X2_2137 ( .A(_abc_41356_new_n6330_), .B(_abc_41356_new_n6331_), .Y(_abc_41356_new_n6332_));
OR2X2 OR2X2_2138 ( .A(_abc_41356_new_n6334_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6335_));
OR2X2 OR2X2_2139 ( .A(_abc_41356_new_n6333_), .B(_abc_41356_new_n6335_), .Y(_abc_41356_new_n6336_));
OR2X2 OR2X2_214 ( .A(_abc_41356_new_n1183_), .B(_abc_41356_new_n1184_), .Y(_abc_41356_new_n1185_));
OR2X2 OR2X2_2140 ( .A(_abc_41356_new_n6336_), .B(_abc_41356_new_n6328_), .Y(_abc_41356_new_n6337_));
OR2X2 OR2X2_2141 ( .A(_abc_41356_new_n6288_), .B(sp_13_), .Y(_abc_41356_new_n6339_));
OR2X2 OR2X2_2142 ( .A(_abc_41356_new_n6344_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6345_));
OR2X2 OR2X2_2143 ( .A(_abc_41356_new_n6343_), .B(_abc_41356_new_n6345_), .Y(_abc_41356_new_n6346_));
OR2X2 OR2X2_2144 ( .A(_abc_41356_new_n6342_), .B(_abc_41356_new_n6346_), .Y(_abc_41356_new_n6347_));
OR2X2 OR2X2_2145 ( .A(_abc_41356_new_n6347_), .B(_abc_41356_new_n6341_), .Y(_abc_41356_new_n6348_));
OR2X2 OR2X2_2146 ( .A(_abc_41356_new_n5853_), .B(sp_13_), .Y(_abc_41356_new_n6349_));
OR2X2 OR2X2_2147 ( .A(_abc_41356_new_n6354_), .B(_abc_41356_new_n6355_), .Y(_abc_41356_new_n6356_));
OR2X2 OR2X2_2148 ( .A(_abc_41356_new_n6356_), .B(_abc_41356_new_n6353_), .Y(_abc_41356_new_n6357_));
OR2X2 OR2X2_2149 ( .A(_abc_41356_new_n6352_), .B(_abc_41356_new_n6357_), .Y(_abc_41356_new_n6358_));
OR2X2 OR2X2_215 ( .A(_abc_41356_new_n1185_), .B(_abc_41356_new_n1182_), .Y(_abc_41356_new_n1186_));
OR2X2 OR2X2_2150 ( .A(_abc_41356_new_n6359_), .B(_abc_41356_new_n6322_), .Y(_0sp_15_0__13_));
OR2X2 OR2X2_2151 ( .A(_abc_41356_new_n6324_), .B(sp_14_), .Y(_abc_41356_new_n6365_));
OR2X2 OR2X2_2152 ( .A(_abc_41356_new_n6370_), .B(_abc_41356_new_n6368_), .Y(_abc_41356_new_n6371_));
OR2X2 OR2X2_2153 ( .A(_abc_41356_new_n6373_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6374_));
OR2X2 OR2X2_2154 ( .A(_abc_41356_new_n6372_), .B(_abc_41356_new_n6374_), .Y(_abc_41356_new_n6375_));
OR2X2 OR2X2_2155 ( .A(_abc_41356_new_n6375_), .B(_abc_41356_new_n6367_), .Y(_abc_41356_new_n6376_));
OR2X2 OR2X2_2156 ( .A(_abc_41356_new_n6323_), .B(sp_14_), .Y(_abc_41356_new_n6378_));
OR2X2 OR2X2_2157 ( .A(_abc_41356_new_n6383_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6384_));
OR2X2 OR2X2_2158 ( .A(_abc_41356_new_n6382_), .B(_abc_41356_new_n6384_), .Y(_abc_41356_new_n6385_));
OR2X2 OR2X2_2159 ( .A(_abc_41356_new_n6381_), .B(_abc_41356_new_n6385_), .Y(_abc_41356_new_n6386_));
OR2X2 OR2X2_216 ( .A(_abc_41356_new_n1186_), .B(_abc_41356_new_n1181_), .Y(_abc_41356_new_n1187_));
OR2X2 OR2X2_2160 ( .A(_abc_41356_new_n6386_), .B(_abc_41356_new_n6380_), .Y(_abc_41356_new_n6387_));
OR2X2 OR2X2_2161 ( .A(_abc_41356_new_n5853_), .B(sp_14_), .Y(_abc_41356_new_n6388_));
OR2X2 OR2X2_2162 ( .A(_abc_41356_new_n6393_), .B(_abc_41356_new_n6394_), .Y(_abc_41356_new_n6395_));
OR2X2 OR2X2_2163 ( .A(_abc_41356_new_n6395_), .B(_abc_41356_new_n6392_), .Y(_abc_41356_new_n6396_));
OR2X2 OR2X2_2164 ( .A(_abc_41356_new_n6391_), .B(_abc_41356_new_n6396_), .Y(_abc_41356_new_n6397_));
OR2X2 OR2X2_2165 ( .A(_abc_41356_new_n6398_), .B(_abc_41356_new_n6361_), .Y(_0sp_15_0__14_));
OR2X2 OR2X2_2166 ( .A(_abc_41356_new_n6401_), .B(_abc_41356_new_n6402_), .Y(_abc_41356_new_n6403_));
OR2X2 OR2X2_2167 ( .A(_abc_41356_new_n6368_), .B(sp_15_), .Y(_abc_41356_new_n6405_));
OR2X2 OR2X2_2168 ( .A(_abc_41356_new_n5380_), .B(sp_0_), .Y(_abc_41356_new_n6406_));
OR2X2 OR2X2_2169 ( .A(_abc_41356_new_n6409_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6410_));
OR2X2 OR2X2_217 ( .A(_abc_41356_new_n1187_), .B(_abc_41356_new_n1189_), .Y(_abc_41356_new_n1190_));
OR2X2 OR2X2_2170 ( .A(_abc_41356_new_n6408_), .B(_abc_41356_new_n6410_), .Y(_abc_41356_new_n6411_));
OR2X2 OR2X2_2171 ( .A(_abc_41356_new_n6411_), .B(_abc_41356_new_n6404_), .Y(_abc_41356_new_n6412_));
OR2X2 OR2X2_2172 ( .A(_abc_41356_new_n6413_), .B(_abc_41356_new_n6414_), .Y(_abc_41356_new_n6415_));
OR2X2 OR2X2_2173 ( .A(_abc_41356_new_n6419_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6420_));
OR2X2 OR2X2_2174 ( .A(_abc_41356_new_n6418_), .B(_abc_41356_new_n6420_), .Y(_abc_41356_new_n6421_));
OR2X2 OR2X2_2175 ( .A(_abc_41356_new_n6417_), .B(_abc_41356_new_n6421_), .Y(_abc_41356_new_n6422_));
OR2X2 OR2X2_2176 ( .A(_abc_41356_new_n6422_), .B(_abc_41356_new_n6416_), .Y(_abc_41356_new_n6423_));
OR2X2 OR2X2_2177 ( .A(_abc_41356_new_n5853_), .B(sp_15_), .Y(_abc_41356_new_n6424_));
OR2X2 OR2X2_2178 ( .A(_abc_41356_new_n6429_), .B(_abc_41356_new_n6430_), .Y(_abc_41356_new_n6431_));
OR2X2 OR2X2_2179 ( .A(_abc_41356_new_n6431_), .B(_abc_41356_new_n6428_), .Y(_abc_41356_new_n6432_));
OR2X2 OR2X2_218 ( .A(_abc_41356_new_n1109_), .B(_abc_41356_new_n1117_), .Y(_abc_41356_new_n1193_));
OR2X2 OR2X2_2180 ( .A(_abc_41356_new_n6427_), .B(_abc_41356_new_n6432_), .Y(_abc_41356_new_n6433_));
OR2X2 OR2X2_2181 ( .A(_abc_41356_new_n6434_), .B(_abc_41356_new_n6400_), .Y(_0sp_15_0__15_));
OR2X2 OR2X2_2182 ( .A(_abc_41356_new_n6436_), .B(regfil_0__0_), .Y(_abc_41356_new_n6437_));
OR2X2 OR2X2_2183 ( .A(_abc_41356_new_n663_), .B(_abc_41356_new_n6438_), .Y(_abc_41356_new_n6439_));
OR2X2 OR2X2_2184 ( .A(_abc_41356_new_n6436_), .B(regfil_0__1_), .Y(_abc_41356_new_n6441_));
OR2X2 OR2X2_2185 ( .A(_abc_41356_new_n771_), .B(_abc_41356_new_n6438_), .Y(_abc_41356_new_n6442_));
OR2X2 OR2X2_2186 ( .A(_abc_41356_new_n6436_), .B(regfil_0__2_), .Y(_abc_41356_new_n6444_));
OR2X2 OR2X2_2187 ( .A(_abc_41356_new_n824_), .B(_abc_41356_new_n6438_), .Y(_abc_41356_new_n6445_));
OR2X2 OR2X2_2188 ( .A(_abc_41356_new_n6436_), .B(regfil_0__3_), .Y(_abc_41356_new_n6447_));
OR2X2 OR2X2_2189 ( .A(_abc_41356_new_n885_), .B(_abc_41356_new_n6438_), .Y(_abc_41356_new_n6448_));
OR2X2 OR2X2_219 ( .A(_abc_41356_new_n1196_), .B(_abc_41356_new_n1197_), .Y(_abc_41356_new_n1198_));
OR2X2 OR2X2_2190 ( .A(_abc_41356_new_n6436_), .B(regfil_0__4_), .Y(_abc_41356_new_n6450_));
OR2X2 OR2X2_2191 ( .A(_abc_41356_new_n952_), .B(_abc_41356_new_n6438_), .Y(_abc_41356_new_n6451_));
OR2X2 OR2X2_2192 ( .A(_abc_41356_new_n6436_), .B(regfil_0__5_), .Y(_abc_41356_new_n6453_));
OR2X2 OR2X2_2193 ( .A(_abc_41356_new_n1019_), .B(_abc_41356_new_n6438_), .Y(_abc_41356_new_n6454_));
OR2X2 OR2X2_2194 ( .A(_abc_41356_new_n6436_), .B(regfil_0__6_), .Y(_abc_41356_new_n6456_));
OR2X2 OR2X2_2195 ( .A(_abc_41356_new_n1091_), .B(_abc_41356_new_n6438_), .Y(_abc_41356_new_n6457_));
OR2X2 OR2X2_2196 ( .A(_abc_41356_new_n6436_), .B(regfil_0__7_), .Y(_abc_41356_new_n6459_));
OR2X2 OR2X2_2197 ( .A(_abc_41356_new_n1173_), .B(_abc_41356_new_n6438_), .Y(_abc_41356_new_n6460_));
OR2X2 OR2X2_2198 ( .A(_abc_41356_new_n4148_), .B(_abc_41356_new_n677_), .Y(_abc_41356_new_n6462_));
OR2X2 OR2X2_2199 ( .A(_abc_41356_new_n6464_), .B(_abc_41356_new_n6465_), .Y(_abc_41356_new_n6466_));
OR2X2 OR2X2_22 ( .A(_abc_41356_new_n653_), .B(regfil_1__5_), .Y(_abc_41356_new_n654_));
OR2X2 OR2X2_220 ( .A(_abc_41356_new_n1195_), .B(_abc_41356_new_n1198_), .Y(_abc_41356_new_n1199_));
OR2X2 OR2X2_2200 ( .A(_abc_41356_new_n6467_), .B(_abc_41356_new_n6468_), .Y(_abc_41356_new_n6469_));
OR2X2 OR2X2_2201 ( .A(_abc_41356_new_n1413_), .B(_abc_41356_new_n535_), .Y(_abc_41356_new_n6473_));
OR2X2 OR2X2_2202 ( .A(_abc_41356_new_n6474_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n6475_));
OR2X2 OR2X2_2203 ( .A(_abc_41356_new_n6475_), .B(_abc_41356_new_n6472_), .Y(_abc_41356_new_n6476_));
OR2X2 OR2X2_2204 ( .A(_abc_41356_new_n1414_), .B(_abc_41356_new_n5890_), .Y(_abc_41356_new_n6480_));
OR2X2 OR2X2_2205 ( .A(_abc_41356_new_n6480_), .B(_abc_41356_new_n6479_), .Y(_abc_41356_new_n6481_));
OR2X2 OR2X2_2206 ( .A(_abc_41356_new_n6490_), .B(pc_0_), .Y(_abc_41356_new_n6491_));
OR2X2 OR2X2_2207 ( .A(_abc_41356_new_n6487_), .B(_abc_41356_new_n6491_), .Y(_abc_41356_new_n6492_));
OR2X2 OR2X2_2208 ( .A(_abc_41356_new_n3495_), .B(_abc_41356_new_n3723_), .Y(_abc_41356_new_n6493_));
OR2X2 OR2X2_2209 ( .A(_abc_41356_new_n6498_), .B(_abc_41356_new_n6493_), .Y(_abc_41356_new_n6499_));
OR2X2 OR2X2_221 ( .A(_abc_41356_new_n1204_), .B(_abc_41356_new_n1190_), .Y(_abc_41356_new_n1205_));
OR2X2 OR2X2_2210 ( .A(_abc_41356_new_n6500_), .B(_abc_41356_new_n6471_), .Y(_abc_41356_new_n6501_));
OR2X2 OR2X2_2211 ( .A(_abc_41356_new_n5840_), .B(_abc_41356_new_n6503_), .Y(_abc_41356_new_n6504_));
OR2X2 OR2X2_2212 ( .A(_abc_41356_new_n6507_), .B(_abc_41356_new_n6508_), .Y(_abc_41356_new_n6509_));
OR2X2 OR2X2_2213 ( .A(_abc_41356_new_n6502_), .B(_abc_41356_new_n6509_), .Y(_abc_41356_new_n6510_));
OR2X2 OR2X2_2214 ( .A(_abc_41356_new_n6510_), .B(_abc_41356_new_n6470_), .Y(_abc_41356_new_n6511_));
OR2X2 OR2X2_2215 ( .A(_abc_41356_new_n554_), .B(_abc_41356_new_n6515_), .Y(_abc_41356_new_n6516_));
OR2X2 OR2X2_2216 ( .A(_abc_41356_new_n6516_), .B(_abc_41356_new_n6514_), .Y(_abc_41356_new_n6517_));
OR2X2 OR2X2_2217 ( .A(_abc_41356_new_n4158_), .B(_abc_41356_new_n536_), .Y(_abc_41356_new_n6522_));
OR2X2 OR2X2_2218 ( .A(_abc_41356_new_n6522_), .B(_abc_41356_new_n4164_), .Y(_abc_41356_new_n6523_));
OR2X2 OR2X2_2219 ( .A(_abc_41356_new_n3299_), .B(_abc_41356_new_n3349_), .Y(_abc_41356_new_n6524_));
OR2X2 OR2X2_222 ( .A(_abc_41356_new_n1177_), .B(_abc_41356_new_n1205_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_7_));
OR2X2 OR2X2_2220 ( .A(_abc_41356_new_n6524_), .B(_abc_41356_new_n2377_), .Y(_abc_41356_new_n6525_));
OR2X2 OR2X2_2221 ( .A(_abc_41356_new_n6523_), .B(_abc_41356_new_n6525_), .Y(_abc_41356_new_n6526_));
OR2X2 OR2X2_2222 ( .A(_abc_41356_new_n3393_), .B(_abc_41356_new_n6479_), .Y(_abc_41356_new_n6527_));
OR2X2 OR2X2_2223 ( .A(_abc_41356_new_n6475_), .B(_abc_41356_new_n6527_), .Y(_abc_41356_new_n6528_));
OR2X2 OR2X2_2224 ( .A(_abc_41356_new_n6526_), .B(_abc_41356_new_n6528_), .Y(_abc_41356_new_n6529_));
OR2X2 OR2X2_2225 ( .A(_abc_41356_new_n6540_), .B(_abc_41356_new_n6541_), .Y(_abc_41356_new_n6542_));
OR2X2 OR2X2_2226 ( .A(_abc_41356_new_n6542_), .B(_abc_41356_new_n4148_), .Y(_abc_41356_new_n6543_));
OR2X2 OR2X2_2227 ( .A(_abc_41356_new_n6539_), .B(_abc_41356_new_n6543_), .Y(_abc_41356_new_n6544_));
OR2X2 OR2X2_2228 ( .A(_abc_41356_new_n4149_), .B(pc_1_), .Y(_abc_41356_new_n6545_));
OR2X2 OR2X2_2229 ( .A(_abc_41356_new_n6553_), .B(_abc_41356_new_n6552_), .Y(_abc_41356_new_n6554_));
OR2X2 OR2X2_223 ( .A(_abc_41356_new_n663_), .B(_abc_41356_new_n1213_), .Y(_abc_41356_new_n1214_));
OR2X2 OR2X2_2230 ( .A(_abc_41356_new_n6554_), .B(_abc_41356_new_n6551_), .Y(_abc_41356_new_n6555_));
OR2X2 OR2X2_2231 ( .A(_abc_41356_new_n6550_), .B(_abc_41356_new_n6555_), .Y(_abc_41356_new_n6556_));
OR2X2 OR2X2_2232 ( .A(_abc_41356_new_n6556_), .B(_abc_41356_new_n6549_), .Y(_abc_41356_new_n6557_));
OR2X2 OR2X2_2233 ( .A(_abc_41356_new_n6558_), .B(_abc_41356_new_n6548_), .Y(_abc_41356_new_n6559_));
OR2X2 OR2X2_2234 ( .A(_abc_41356_new_n6559_), .B(_abc_41356_new_n6547_), .Y(_abc_41356_new_n6560_));
OR2X2 OR2X2_2235 ( .A(_abc_41356_new_n6562_), .B(_abc_41356_new_n6563_), .Y(_abc_41356_new_n6564_));
OR2X2 OR2X2_2236 ( .A(_abc_41356_new_n6561_), .B(_abc_41356_new_n6564_), .Y(_abc_41356_new_n6565_));
OR2X2 OR2X2_2237 ( .A(_abc_41356_new_n6537_), .B(_abc_41356_new_n3813_), .Y(_abc_41356_new_n6567_));
OR2X2 OR2X2_2238 ( .A(_abc_41356_new_n4125_), .B(_abc_41356_new_n3820_), .Y(_abc_41356_new_n6568_));
OR2X2 OR2X2_2239 ( .A(_abc_41356_new_n3818_), .B(_abc_41356_new_n2070_), .Y(_abc_41356_new_n6569_));
OR2X2 OR2X2_224 ( .A(_abc_41356_new_n1226_), .B(_abc_41356_new_n1228_), .Y(_abc_41356_new_n1229_));
OR2X2 OR2X2_2240 ( .A(_abc_41356_new_n678_), .B(_abc_41356_new_n6569_), .Y(_abc_41356_new_n6570_));
OR2X2 OR2X2_2241 ( .A(_abc_41356_new_n6574_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6575_));
OR2X2 OR2X2_2242 ( .A(_abc_41356_new_n6573_), .B(_abc_41356_new_n6575_), .Y(_abc_41356_new_n6576_));
OR2X2 OR2X2_2243 ( .A(_abc_41356_new_n6486_), .B(_abc_41356_new_n3813_), .Y(_abc_41356_new_n6579_));
OR2X2 OR2X2_2244 ( .A(_abc_41356_new_n3494_), .B(_abc_41356_new_n6569_), .Y(_abc_41356_new_n6580_));
OR2X2 OR2X2_2245 ( .A(_abc_41356_new_n6494_), .B(_abc_41356_new_n1257_), .Y(_abc_41356_new_n6581_));
OR2X2 OR2X2_2246 ( .A(_abc_41356_new_n6489_), .B(_abc_41356_new_n3820_), .Y(_abc_41356_new_n6582_));
OR2X2 OR2X2_2247 ( .A(_abc_41356_new_n6586_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6587_));
OR2X2 OR2X2_2248 ( .A(_abc_41356_new_n5853_), .B(_abc_41356_new_n3813_), .Y(_abc_41356_new_n6588_));
OR2X2 OR2X2_2249 ( .A(_abc_41356_new_n6593_), .B(_abc_41356_new_n6594_), .Y(_abc_41356_new_n6595_));
OR2X2 OR2X2_225 ( .A(_abc_41356_new_n1229_), .B(_abc_41356_new_n1223_), .Y(_abc_41356_new_n1230_));
OR2X2 OR2X2_2250 ( .A(_abc_41356_new_n6592_), .B(_abc_41356_new_n6595_), .Y(_abc_41356_new_n6596_));
OR2X2 OR2X2_2251 ( .A(_abc_41356_new_n6537_), .B(_abc_41356_new_n6598_), .Y(_abc_41356_new_n6599_));
OR2X2 OR2X2_2252 ( .A(_abc_41356_new_n4125_), .B(_abc_41356_new_n6600_), .Y(_abc_41356_new_n6601_));
OR2X2 OR2X2_2253 ( .A(_abc_41356_new_n6604_), .B(_abc_41356_new_n2071_), .Y(_abc_41356_new_n6605_));
OR2X2 OR2X2_2254 ( .A(_abc_41356_new_n6605_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n6606_));
OR2X2 OR2X2_2255 ( .A(_abc_41356_new_n6610_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6611_));
OR2X2 OR2X2_2256 ( .A(_abc_41356_new_n6609_), .B(_abc_41356_new_n6611_), .Y(_abc_41356_new_n6612_));
OR2X2 OR2X2_2257 ( .A(_abc_41356_new_n6486_), .B(_abc_41356_new_n6598_), .Y(_abc_41356_new_n6615_));
OR2X2 OR2X2_2258 ( .A(_abc_41356_new_n3494_), .B(_abc_41356_new_n6605_), .Y(_abc_41356_new_n6618_));
OR2X2 OR2X2_2259 ( .A(_abc_41356_new_n6626_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6627_));
OR2X2 OR2X2_226 ( .A(_abc_41356_new_n1212_), .B(regfil_4__0_), .Y(_abc_41356_new_n1243_));
OR2X2 OR2X2_2260 ( .A(_abc_41356_new_n6634_), .B(_abc_41356_new_n6635_), .Y(_abc_41356_new_n6636_));
OR2X2 OR2X2_2261 ( .A(_abc_41356_new_n6633_), .B(_abc_41356_new_n6636_), .Y(_abc_41356_new_n6637_));
OR2X2 OR2X2_2262 ( .A(_abc_41356_new_n2071_), .B(pc_4_), .Y(_abc_41356_new_n6643_));
OR2X2 OR2X2_2263 ( .A(_abc_41356_new_n6645_), .B(_abc_41356_new_n4148_), .Y(_abc_41356_new_n6646_));
OR2X2 OR2X2_2264 ( .A(_abc_41356_new_n6640_), .B(_abc_41356_new_n6646_), .Y(_abc_41356_new_n6647_));
OR2X2 OR2X2_2265 ( .A(_abc_41356_new_n6639_), .B(_abc_41356_new_n6647_), .Y(_abc_41356_new_n6648_));
OR2X2 OR2X2_2266 ( .A(_abc_41356_new_n4149_), .B(pc_4_), .Y(_abc_41356_new_n6649_));
OR2X2 OR2X2_2267 ( .A(_abc_41356_new_n6651_), .B(_abc_41356_new_n6652_), .Y(_abc_41356_new_n6653_));
OR2X2 OR2X2_2268 ( .A(_abc_41356_new_n6659_), .B(_abc_41356_new_n6660_), .Y(_abc_41356_new_n6661_));
OR2X2 OR2X2_2269 ( .A(_abc_41356_new_n6661_), .B(_abc_41356_new_n6658_), .Y(_abc_41356_new_n6662_));
OR2X2 OR2X2_227 ( .A(_abc_41356_new_n1245_), .B(_abc_41356_new_n1246_), .Y(_abc_41356_new_n1247_));
OR2X2 OR2X2_2270 ( .A(_abc_41356_new_n6662_), .B(_abc_41356_new_n6657_), .Y(_abc_41356_new_n6663_));
OR2X2 OR2X2_2271 ( .A(_abc_41356_new_n6656_), .B(_abc_41356_new_n6663_), .Y(_abc_41356_new_n6664_));
OR2X2 OR2X2_2272 ( .A(_abc_41356_new_n6664_), .B(_abc_41356_new_n6655_), .Y(_abc_41356_new_n6665_));
OR2X2 OR2X2_2273 ( .A(_abc_41356_new_n6667_), .B(_abc_41356_new_n6668_), .Y(_abc_41356_new_n6669_));
OR2X2 OR2X2_2274 ( .A(_abc_41356_new_n6666_), .B(_abc_41356_new_n6669_), .Y(_abc_41356_new_n6670_));
OR2X2 OR2X2_2275 ( .A(_abc_41356_new_n6654_), .B(_abc_41356_new_n6670_), .Y(_abc_41356_new_n6671_));
OR2X2 OR2X2_2276 ( .A(_abc_41356_new_n6537_), .B(_abc_41356_new_n3982_), .Y(_abc_41356_new_n6673_));
OR2X2 OR2X2_2277 ( .A(_abc_41356_new_n4125_), .B(_abc_41356_new_n3987_), .Y(_abc_41356_new_n6674_));
OR2X2 OR2X2_2278 ( .A(_abc_41356_new_n6676_), .B(_abc_41356_new_n6675_), .Y(_abc_41356_new_n6677_));
OR2X2 OR2X2_2279 ( .A(_abc_41356_new_n6677_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n6678_));
OR2X2 OR2X2_228 ( .A(_abc_41356_new_n1236_), .B(regfil_2__0_), .Y(_abc_41356_new_n1249_));
OR2X2 OR2X2_2280 ( .A(_abc_41356_new_n6682_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6683_));
OR2X2 OR2X2_2281 ( .A(_abc_41356_new_n6681_), .B(_abc_41356_new_n6683_), .Y(_abc_41356_new_n6684_));
OR2X2 OR2X2_2282 ( .A(_abc_41356_new_n6486_), .B(_abc_41356_new_n3982_), .Y(_abc_41356_new_n6687_));
OR2X2 OR2X2_2283 ( .A(_abc_41356_new_n2061_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n6690_));
OR2X2 OR2X2_2284 ( .A(_abc_41356_new_n6677_), .B(_abc_41356_new_n3494_), .Y(_abc_41356_new_n6693_));
OR2X2 OR2X2_2285 ( .A(_abc_41356_new_n6698_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6699_));
OR2X2 OR2X2_2286 ( .A(_abc_41356_new_n6706_), .B(_abc_41356_new_n6707_), .Y(_abc_41356_new_n6708_));
OR2X2 OR2X2_2287 ( .A(_abc_41356_new_n6705_), .B(_abc_41356_new_n6708_), .Y(_abc_41356_new_n6709_));
OR2X2 OR2X2_2288 ( .A(_abc_41356_new_n6537_), .B(_abc_41356_new_n6711_), .Y(_abc_41356_new_n6712_));
OR2X2 OR2X2_2289 ( .A(_abc_41356_new_n6713_), .B(_abc_41356_new_n4125_), .Y(_abc_41356_new_n6714_));
OR2X2 OR2X2_229 ( .A(_abc_41356_new_n1266_), .B(_abc_41356_new_n1251_), .Y(_abc_41356_new_n1269_));
OR2X2 OR2X2_2290 ( .A(_abc_41356_new_n6718_), .B(_abc_41356_new_n6715_), .Y(_abc_41356_new_n6719_));
OR2X2 OR2X2_2291 ( .A(_abc_41356_new_n6719_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n6720_));
OR2X2 OR2X2_2292 ( .A(_abc_41356_new_n6724_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6725_));
OR2X2 OR2X2_2293 ( .A(_abc_41356_new_n6723_), .B(_abc_41356_new_n6725_), .Y(_abc_41356_new_n6726_));
OR2X2 OR2X2_2294 ( .A(_abc_41356_new_n6486_), .B(_abc_41356_new_n6711_), .Y(_abc_41356_new_n6729_));
OR2X2 OR2X2_2295 ( .A(_abc_41356_new_n6713_), .B(_abc_41356_new_n6489_), .Y(_abc_41356_new_n6730_));
OR2X2 OR2X2_2296 ( .A(_abc_41356_new_n6494_), .B(_abc_41356_new_n1253_), .Y(_abc_41356_new_n6731_));
OR2X2 OR2X2_2297 ( .A(_abc_41356_new_n6719_), .B(_abc_41356_new_n3494_), .Y(_abc_41356_new_n6732_));
OR2X2 OR2X2_2298 ( .A(_abc_41356_new_n6736_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6737_));
OR2X2 OR2X2_2299 ( .A(_abc_41356_new_n6711_), .B(_abc_41356_new_n5853_), .Y(_abc_41356_new_n6738_));
OR2X2 OR2X2_23 ( .A(_abc_41356_new_n654_), .B(regfil_1__6_), .Y(_abc_41356_new_n655_));
OR2X2 OR2X2_230 ( .A(_abc_41356_new_n1279_), .B(regfil_4__0_), .Y(_abc_41356_new_n1280_));
OR2X2 OR2X2_2300 ( .A(_abc_41356_new_n6743_), .B(_abc_41356_new_n6744_), .Y(_abc_41356_new_n6745_));
OR2X2 OR2X2_2301 ( .A(_abc_41356_new_n6742_), .B(_abc_41356_new_n6745_), .Y(_abc_41356_new_n6746_));
OR2X2 OR2X2_2302 ( .A(_abc_41356_new_n6537_), .B(_abc_41356_new_n4074_), .Y(_abc_41356_new_n6748_));
OR2X2 OR2X2_2303 ( .A(_abc_41356_new_n6715_), .B(pc_7_), .Y(_abc_41356_new_n6753_));
OR2X2 OR2X2_2304 ( .A(_abc_41356_new_n6760_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6761_));
OR2X2 OR2X2_2305 ( .A(_abc_41356_new_n6759_), .B(_abc_41356_new_n6761_), .Y(_abc_41356_new_n6762_));
OR2X2 OR2X2_2306 ( .A(_abc_41356_new_n6486_), .B(_abc_41356_new_n4074_), .Y(_abc_41356_new_n6767_));
OR2X2 OR2X2_2307 ( .A(_abc_41356_new_n6775_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6776_));
OR2X2 OR2X2_2308 ( .A(_abc_41356_new_n6783_), .B(_abc_41356_new_n6784_), .Y(_abc_41356_new_n6785_));
OR2X2 OR2X2_2309 ( .A(_abc_41356_new_n6782_), .B(_abc_41356_new_n6785_), .Y(_abc_41356_new_n6786_));
OR2X2 OR2X2_231 ( .A(_abc_41356_new_n1283_), .B(_abc_41356_new_n1220_), .Y(_abc_41356_new_n1284_));
OR2X2 OR2X2_2310 ( .A(_abc_41356_new_n6537_), .B(_abc_41356_new_n2077_), .Y(_abc_41356_new_n6788_));
OR2X2 OR2X2_2311 ( .A(_abc_41356_new_n4125_), .B(_abc_41356_new_n2044_), .Y(_abc_41356_new_n6789_));
OR2X2 OR2X2_2312 ( .A(_abc_41356_new_n6790_), .B(_abc_41356_new_n6791_), .Y(_abc_41356_new_n6792_));
OR2X2 OR2X2_2313 ( .A(_abc_41356_new_n6792_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n6793_));
OR2X2 OR2X2_2314 ( .A(_abc_41356_new_n6797_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6798_));
OR2X2 OR2X2_2315 ( .A(_abc_41356_new_n6796_), .B(_abc_41356_new_n6798_), .Y(_abc_41356_new_n6799_));
OR2X2 OR2X2_2316 ( .A(_abc_41356_new_n2044_), .B(_abc_41356_new_n6489_), .Y(_abc_41356_new_n6802_));
OR2X2 OR2X2_2317 ( .A(_abc_41356_new_n6792_), .B(_abc_41356_new_n3494_), .Y(_abc_41356_new_n6803_));
OR2X2 OR2X2_2318 ( .A(_abc_41356_new_n6486_), .B(_abc_41356_new_n2077_), .Y(_abc_41356_new_n6805_));
OR2X2 OR2X2_2319 ( .A(_abc_41356_new_n6810_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6811_));
OR2X2 OR2X2_232 ( .A(regfil_5__1_), .B(sp_1_), .Y(_abc_41356_new_n1290_));
OR2X2 OR2X2_2320 ( .A(_abc_41356_new_n2077_), .B(_abc_41356_new_n5853_), .Y(_abc_41356_new_n6812_));
OR2X2 OR2X2_2321 ( .A(_abc_41356_new_n6817_), .B(_abc_41356_new_n6818_), .Y(_abc_41356_new_n6819_));
OR2X2 OR2X2_2322 ( .A(_abc_41356_new_n6816_), .B(_abc_41356_new_n6819_), .Y(_abc_41356_new_n6820_));
OR2X2 OR2X2_2323 ( .A(_abc_41356_new_n6825_), .B(_abc_41356_new_n6822_), .Y(_abc_41356_new_n6826_));
OR2X2 OR2X2_2324 ( .A(_abc_41356_new_n6826_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n6827_));
OR2X2 OR2X2_2325 ( .A(_abc_41356_new_n6829_), .B(_abc_41356_new_n4125_), .Y(_abc_41356_new_n6830_));
OR2X2 OR2X2_2326 ( .A(_abc_41356_new_n6537_), .B(_abc_41356_new_n6831_), .Y(_abc_41356_new_n6832_));
OR2X2 OR2X2_2327 ( .A(_abc_41356_new_n6835_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6836_));
OR2X2 OR2X2_2328 ( .A(_abc_41356_new_n6834_), .B(_abc_41356_new_n6836_), .Y(_abc_41356_new_n6837_));
OR2X2 OR2X2_2329 ( .A(_abc_41356_new_n6829_), .B(_abc_41356_new_n6489_), .Y(_abc_41356_new_n6840_));
OR2X2 OR2X2_233 ( .A(_abc_41356_new_n1299_), .B(_abc_41356_new_n1297_), .Y(_abc_41356_new_n1300_));
OR2X2 OR2X2_2330 ( .A(_abc_41356_new_n6826_), .B(_abc_41356_new_n3494_), .Y(_abc_41356_new_n6841_));
OR2X2 OR2X2_2331 ( .A(_abc_41356_new_n6486_), .B(_abc_41356_new_n6831_), .Y(_abc_41356_new_n6843_));
OR2X2 OR2X2_2332 ( .A(_abc_41356_new_n6848_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6849_));
OR2X2 OR2X2_2333 ( .A(_abc_41356_new_n6831_), .B(_abc_41356_new_n5853_), .Y(_abc_41356_new_n6850_));
OR2X2 OR2X2_2334 ( .A(_abc_41356_new_n6855_), .B(_abc_41356_new_n6856_), .Y(_abc_41356_new_n6857_));
OR2X2 OR2X2_2335 ( .A(_abc_41356_new_n6854_), .B(_abc_41356_new_n6857_), .Y(_abc_41356_new_n6858_));
OR2X2 OR2X2_2336 ( .A(_abc_41356_new_n6862_), .B(_abc_41356_new_n6860_), .Y(_abc_41356_new_n6863_));
OR2X2 OR2X2_2337 ( .A(_abc_41356_new_n6863_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n6864_));
OR2X2 OR2X2_2338 ( .A(_abc_41356_new_n6537_), .B(_abc_41356_new_n2159_), .Y(_abc_41356_new_n6865_));
OR2X2 OR2X2_2339 ( .A(_abc_41356_new_n2151_), .B(_abc_41356_new_n4125_), .Y(_abc_41356_new_n6866_));
OR2X2 OR2X2_234 ( .A(_abc_41356_new_n1304_), .B(_abc_41356_new_n1302_), .Y(_abc_41356_new_n1305_));
OR2X2 OR2X2_2340 ( .A(_abc_41356_new_n6870_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n6871_));
OR2X2 OR2X2_2341 ( .A(_abc_41356_new_n6869_), .B(_abc_41356_new_n6871_), .Y(_abc_41356_new_n6872_));
OR2X2 OR2X2_2342 ( .A(_abc_41356_new_n6494_), .B(_abc_41356_new_n1580_), .Y(_abc_41356_new_n6875_));
OR2X2 OR2X2_2343 ( .A(_abc_41356_new_n2151_), .B(_abc_41356_new_n6489_), .Y(_abc_41356_new_n6876_));
OR2X2 OR2X2_2344 ( .A(_abc_41356_new_n6863_), .B(_abc_41356_new_n3494_), .Y(_abc_41356_new_n6877_));
OR2X2 OR2X2_2345 ( .A(_abc_41356_new_n6486_), .B(_abc_41356_new_n2159_), .Y(_abc_41356_new_n6878_));
OR2X2 OR2X2_2346 ( .A(_abc_41356_new_n6882_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n6883_));
OR2X2 OR2X2_2347 ( .A(_abc_41356_new_n2159_), .B(_abc_41356_new_n5853_), .Y(_abc_41356_new_n6884_));
OR2X2 OR2X2_2348 ( .A(_abc_41356_new_n6889_), .B(_abc_41356_new_n6890_), .Y(_abc_41356_new_n6891_));
OR2X2 OR2X2_2349 ( .A(_abc_41356_new_n6888_), .B(_abc_41356_new_n6891_), .Y(_abc_41356_new_n6892_));
OR2X2 OR2X2_235 ( .A(_abc_41356_new_n1309_), .B(_abc_41356_new_n1302_), .Y(_abc_41356_new_n1310_));
OR2X2 OR2X2_2350 ( .A(_abc_41356_new_n6860_), .B(pc_11_), .Y(_abc_41356_new_n6896_));
OR2X2 OR2X2_2351 ( .A(_abc_41356_new_n6898_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n6899_));
OR2X2 OR2X2_2352 ( .A(_abc_41356_new_n6900_), .B(_abc_41356_new_n4125_), .Y(_abc_41356_new_n6901_));
OR2X2 OR2X2_2353 ( .A(_abc_41356_new_n6537_), .B(_abc_41356_new_n6902_), .Y(_abc_41356_new_n6903_));
OR2X2 OR2X2_2354 ( .A(_abc_41356_new_n4149_), .B(_abc_41356_new_n6906_), .Y(_abc_41356_new_n6907_));
OR2X2 OR2X2_2355 ( .A(_abc_41356_new_n6913_), .B(_abc_41356_new_n6914_), .Y(_abc_41356_new_n6915_));
OR2X2 OR2X2_2356 ( .A(_abc_41356_new_n6917_), .B(_abc_41356_new_n6916_), .Y(_abc_41356_new_n6918_));
OR2X2 OR2X2_2357 ( .A(_abc_41356_new_n6915_), .B(_abc_41356_new_n6918_), .Y(_abc_41356_new_n6919_));
OR2X2 OR2X2_2358 ( .A(_abc_41356_new_n6919_), .B(_abc_41356_new_n6912_), .Y(_abc_41356_new_n6920_));
OR2X2 OR2X2_2359 ( .A(_abc_41356_new_n6921_), .B(_abc_41356_new_n6911_), .Y(_abc_41356_new_n6922_));
OR2X2 OR2X2_236 ( .A(_abc_41356_new_n1308_), .B(_abc_41356_new_n1310_), .Y(_abc_41356_new_n1311_));
OR2X2 OR2X2_2360 ( .A(_abc_41356_new_n6910_), .B(_abc_41356_new_n6922_), .Y(_abc_41356_new_n6923_));
OR2X2 OR2X2_2361 ( .A(_abc_41356_new_n6925_), .B(_abc_41356_new_n6926_), .Y(_abc_41356_new_n6927_));
OR2X2 OR2X2_2362 ( .A(_abc_41356_new_n6924_), .B(_abc_41356_new_n6927_), .Y(_abc_41356_new_n6928_));
OR2X2 OR2X2_2363 ( .A(_abc_41356_new_n6930_), .B(_abc_41356_new_n6931_), .Y(_abc_41356_new_n6932_));
OR2X2 OR2X2_2364 ( .A(_abc_41356_new_n6932_), .B(_abc_41356_new_n678_), .Y(_abc_41356_new_n6933_));
OR2X2 OR2X2_2365 ( .A(_abc_41356_new_n2229_), .B(_abc_41356_new_n4125_), .Y(_abc_41356_new_n6934_));
OR2X2 OR2X2_2366 ( .A(_abc_41356_new_n6537_), .B(_abc_41356_new_n2237_), .Y(_abc_41356_new_n6935_));
OR2X2 OR2X2_2367 ( .A(_abc_41356_new_n4149_), .B(pc_12_), .Y(_abc_41356_new_n6940_));
OR2X2 OR2X2_2368 ( .A(_abc_41356_new_n6949_), .B(_abc_41356_new_n6948_), .Y(_abc_41356_new_n6950_));
OR2X2 OR2X2_2369 ( .A(_abc_41356_new_n6950_), .B(_abc_41356_new_n6947_), .Y(_abc_41356_new_n6951_));
OR2X2 OR2X2_237 ( .A(_abc_41356_new_n1320_), .B(_abc_41356_new_n1318_), .Y(_abc_41356_new_n1321_));
OR2X2 OR2X2_2370 ( .A(_abc_41356_new_n6951_), .B(_abc_41356_new_n6946_), .Y(_abc_41356_new_n6952_));
OR2X2 OR2X2_2371 ( .A(_abc_41356_new_n6952_), .B(_abc_41356_new_n6944_), .Y(_abc_41356_new_n6953_));
OR2X2 OR2X2_2372 ( .A(_abc_41356_new_n6954_), .B(_abc_41356_new_n6943_), .Y(_abc_41356_new_n6955_));
OR2X2 OR2X2_2373 ( .A(_abc_41356_new_n6955_), .B(_abc_41356_new_n6942_), .Y(_abc_41356_new_n6956_));
OR2X2 OR2X2_2374 ( .A(_abc_41356_new_n6958_), .B(_abc_41356_new_n6959_), .Y(_abc_41356_new_n6960_));
OR2X2 OR2X2_2375 ( .A(_abc_41356_new_n6957_), .B(_abc_41356_new_n6960_), .Y(_abc_41356_new_n6961_));
OR2X2 OR2X2_2376 ( .A(_abc_41356_new_n6931_), .B(pc_13_), .Y(_abc_41356_new_n6965_));
OR2X2 OR2X2_2377 ( .A(_abc_41356_new_n6969_), .B(_abc_41356_new_n6968_), .Y(_abc_41356_new_n6970_));
OR2X2 OR2X2_2378 ( .A(_abc_41356_new_n6970_), .B(_abc_41356_new_n4148_), .Y(_abc_41356_new_n6971_));
OR2X2 OR2X2_2379 ( .A(_abc_41356_new_n6971_), .B(_abc_41356_new_n6967_), .Y(_abc_41356_new_n6972_));
OR2X2 OR2X2_238 ( .A(_abc_41356_new_n1326_), .B(_abc_41356_new_n1324_), .Y(_abc_41356_new_n1327_));
OR2X2 OR2X2_2380 ( .A(_abc_41356_new_n4149_), .B(pc_13_), .Y(_abc_41356_new_n6973_));
OR2X2 OR2X2_2381 ( .A(_abc_41356_new_n6978_), .B(_abc_41356_new_n6979_), .Y(_abc_41356_new_n6980_));
OR2X2 OR2X2_2382 ( .A(_abc_41356_new_n6981_), .B(_abc_41356_new_n6982_), .Y(_abc_41356_new_n6983_));
OR2X2 OR2X2_2383 ( .A(_abc_41356_new_n6980_), .B(_abc_41356_new_n6983_), .Y(_abc_41356_new_n6984_));
OR2X2 OR2X2_2384 ( .A(_abc_41356_new_n6984_), .B(_abc_41356_new_n6977_), .Y(_abc_41356_new_n6985_));
OR2X2 OR2X2_2385 ( .A(_abc_41356_new_n6986_), .B(_abc_41356_new_n6976_), .Y(_abc_41356_new_n6987_));
OR2X2 OR2X2_2386 ( .A(_abc_41356_new_n6987_), .B(_abc_41356_new_n6975_), .Y(_abc_41356_new_n6988_));
OR2X2 OR2X2_2387 ( .A(_abc_41356_new_n6990_), .B(_abc_41356_new_n6991_), .Y(_abc_41356_new_n6992_));
OR2X2 OR2X2_2388 ( .A(_abc_41356_new_n6989_), .B(_abc_41356_new_n6992_), .Y(_abc_41356_new_n6993_));
OR2X2 OR2X2_2389 ( .A(_abc_41356_new_n6963_), .B(pc_14_), .Y(_abc_41356_new_n6998_));
OR2X2 OR2X2_239 ( .A(_abc_41356_new_n1338_), .B(_abc_41356_new_n1312_), .Y(_abc_41356_new_n1339_));
OR2X2 OR2X2_2390 ( .A(_abc_41356_new_n7001_), .B(_abc_41356_new_n4148_), .Y(_abc_41356_new_n7002_));
OR2X2 OR2X2_2391 ( .A(_abc_41356_new_n7002_), .B(_abc_41356_new_n7000_), .Y(_abc_41356_new_n7003_));
OR2X2 OR2X2_2392 ( .A(_abc_41356_new_n7003_), .B(_abc_41356_new_n6995_), .Y(_abc_41356_new_n7004_));
OR2X2 OR2X2_2393 ( .A(_abc_41356_new_n4149_), .B(pc_14_), .Y(_abc_41356_new_n7005_));
OR2X2 OR2X2_2394 ( .A(_abc_41356_new_n7012_), .B(_abc_41356_new_n1978_), .Y(_abc_41356_new_n7013_));
OR2X2 OR2X2_2395 ( .A(_abc_41356_new_n7011_), .B(_abc_41356_new_n7013_), .Y(_abc_41356_new_n7014_));
OR2X2 OR2X2_2396 ( .A(_abc_41356_new_n7014_), .B(_abc_41356_new_n7010_), .Y(_abc_41356_new_n7015_));
OR2X2 OR2X2_2397 ( .A(_abc_41356_new_n7015_), .B(_abc_41356_new_n7009_), .Y(_abc_41356_new_n7016_));
OR2X2 OR2X2_2398 ( .A(_abc_41356_new_n7017_), .B(_abc_41356_new_n7008_), .Y(_abc_41356_new_n7018_));
OR2X2 OR2X2_2399 ( .A(_abc_41356_new_n7018_), .B(_abc_41356_new_n7007_), .Y(_abc_41356_new_n7019_));
OR2X2 OR2X2_24 ( .A(_abc_41356_new_n655_), .B(regfil_1__7_), .Y(_abc_41356_new_n656_));
OR2X2 OR2X2_240 ( .A(_abc_41356_new_n1340_), .B(_abc_41356_new_n1329_), .Y(_abc_41356_new_n1341_));
OR2X2 OR2X2_2400 ( .A(_abc_41356_new_n7021_), .B(_abc_41356_new_n7022_), .Y(_abc_41356_new_n7023_));
OR2X2 OR2X2_2401 ( .A(_abc_41356_new_n7020_), .B(_abc_41356_new_n7023_), .Y(_abc_41356_new_n7024_));
OR2X2 OR2X2_2402 ( .A(_abc_41356_new_n6996_), .B(pc_15_), .Y(_abc_41356_new_n7027_));
OR2X2 OR2X2_2403 ( .A(_abc_41356_new_n7031_), .B(_abc_41356_new_n7032_), .Y(_abc_41356_new_n7033_));
OR2X2 OR2X2_2404 ( .A(_abc_41356_new_n7033_), .B(_abc_41356_new_n7026_), .Y(_abc_41356_new_n7034_));
OR2X2 OR2X2_2405 ( .A(_abc_41356_new_n7034_), .B(_abc_41356_new_n4148_), .Y(_abc_41356_new_n7035_));
OR2X2 OR2X2_2406 ( .A(_abc_41356_new_n4149_), .B(pc_15_), .Y(_abc_41356_new_n7036_));
OR2X2 OR2X2_2407 ( .A(_abc_41356_new_n7042_), .B(_abc_41356_new_n3282_), .Y(_abc_41356_new_n7043_));
OR2X2 OR2X2_2408 ( .A(_abc_41356_new_n7041_), .B(_abc_41356_new_n7043_), .Y(_abc_41356_new_n7044_));
OR2X2 OR2X2_2409 ( .A(_abc_41356_new_n7044_), .B(_abc_41356_new_n7040_), .Y(_abc_41356_new_n7045_));
OR2X2 OR2X2_241 ( .A(_abc_41356_new_n1342_), .B(_abc_41356_new_n1339_), .Y(_abc_41356_new_n1343_));
OR2X2 OR2X2_2410 ( .A(_abc_41356_new_n7045_), .B(_abc_41356_new_n7039_), .Y(_abc_41356_new_n7046_));
OR2X2 OR2X2_2411 ( .A(_abc_41356_new_n7047_), .B(_abc_41356_new_n7048_), .Y(_abc_41356_new_n7049_));
OR2X2 OR2X2_2412 ( .A(_abc_41356_new_n7049_), .B(_abc_41356_new_n7038_), .Y(_abc_41356_new_n7050_));
OR2X2 OR2X2_2413 ( .A(_abc_41356_new_n7052_), .B(_abc_41356_new_n7053_), .Y(_abc_41356_new_n7054_));
OR2X2 OR2X2_2414 ( .A(_abc_41356_new_n7051_), .B(_abc_41356_new_n7054_), .Y(_abc_41356_new_n7055_));
OR2X2 OR2X2_2415 ( .A(_abc_41356_new_n7059_), .B(waitr), .Y(_abc_41356_new_n7060_));
OR2X2 OR2X2_2416 ( .A(_abc_41356_new_n7062_), .B(_abc_41356_new_n7057_), .Y(_0writemem_0_0_));
OR2X2 OR2X2_2417 ( .A(_abc_41356_new_n7069_), .B(_abc_41356_new_n7067_), .Y(_abc_41356_new_n7070_));
OR2X2 OR2X2_2418 ( .A(_abc_41356_new_n7070_), .B(_abc_41356_new_n7065_), .Y(_abc_41356_new_n7071_));
OR2X2 OR2X2_2419 ( .A(_abc_41356_new_n7072_), .B(_abc_41356_new_n7073_), .Y(_abc_41356_new_n7074_));
OR2X2 OR2X2_242 ( .A(_abc_41356_new_n1337_), .B(_abc_41356_new_n1343_), .Y(_abc_41356_new_n1344_));
OR2X2 OR2X2_2420 ( .A(_abc_41356_new_n7074_), .B(readmem), .Y(_abc_41356_new_n7075_));
OR2X2 OR2X2_2421 ( .A(_abc_41356_new_n7078_), .B(_abc_41356_new_n7079_), .Y(_abc_41356_new_n7080_));
OR2X2 OR2X2_2422 ( .A(_abc_41356_new_n7083_), .B(reset), .Y(_abc_41356_new_n7084_));
OR2X2 OR2X2_2423 ( .A(_abc_41356_new_n7088_), .B(_abc_41356_new_n7087_), .Y(_abc_41356_new_n7089_));
OR2X2 OR2X2_2424 ( .A(_abc_41356_new_n7089_), .B(_abc_41356_new_n7090_), .Y(_abc_41356_new_n7091_));
OR2X2 OR2X2_2425 ( .A(_abc_41356_new_n7091_), .B(_abc_41356_new_n7086_), .Y(_abc_41356_new_n7092_));
OR2X2 OR2X2_2426 ( .A(_abc_41356_new_n7085_), .B(_abc_41356_new_n7093_), .Y(_0addr_15_0__0_));
OR2X2 OR2X2_2427 ( .A(_abc_41356_new_n7098_), .B(_abc_41356_new_n7097_), .Y(_abc_41356_new_n7099_));
OR2X2 OR2X2_2428 ( .A(_abc_41356_new_n7099_), .B(_abc_41356_new_n7100_), .Y(_abc_41356_new_n7101_));
OR2X2 OR2X2_2429 ( .A(_abc_41356_new_n7101_), .B(_abc_41356_new_n7096_), .Y(_abc_41356_new_n7102_));
OR2X2 OR2X2_243 ( .A(_abc_41356_new_n1346_), .B(_abc_41356_new_n1347_), .Y(_abc_41356_new_n1348_));
OR2X2 OR2X2_2430 ( .A(_abc_41356_new_n7095_), .B(_abc_41356_new_n7103_), .Y(_0addr_15_0__1_));
OR2X2 OR2X2_2431 ( .A(_abc_41356_new_n7108_), .B(_abc_41356_new_n7107_), .Y(_abc_41356_new_n7109_));
OR2X2 OR2X2_2432 ( .A(_abc_41356_new_n7109_), .B(_abc_41356_new_n7110_), .Y(_abc_41356_new_n7111_));
OR2X2 OR2X2_2433 ( .A(_abc_41356_new_n7111_), .B(_abc_41356_new_n7106_), .Y(_abc_41356_new_n7112_));
OR2X2 OR2X2_2434 ( .A(_abc_41356_new_n7105_), .B(_abc_41356_new_n7113_), .Y(_0addr_15_0__2_));
OR2X2 OR2X2_2435 ( .A(_abc_41356_new_n7118_), .B(_abc_41356_new_n7117_), .Y(_abc_41356_new_n7119_));
OR2X2 OR2X2_2436 ( .A(_abc_41356_new_n7119_), .B(_abc_41356_new_n7120_), .Y(_abc_41356_new_n7121_));
OR2X2 OR2X2_2437 ( .A(_abc_41356_new_n7121_), .B(_abc_41356_new_n7116_), .Y(_abc_41356_new_n7122_));
OR2X2 OR2X2_2438 ( .A(_abc_41356_new_n7115_), .B(_abc_41356_new_n7123_), .Y(_0addr_15_0__3_));
OR2X2 OR2X2_2439 ( .A(_abc_41356_new_n7128_), .B(_abc_41356_new_n7127_), .Y(_abc_41356_new_n7129_));
OR2X2 OR2X2_244 ( .A(_abc_41356_new_n1344_), .B(_abc_41356_new_n1349_), .Y(_abc_41356_new_n1352_));
OR2X2 OR2X2_2440 ( .A(_abc_41356_new_n7129_), .B(_abc_41356_new_n7130_), .Y(_abc_41356_new_n7131_));
OR2X2 OR2X2_2441 ( .A(_abc_41356_new_n7131_), .B(_abc_41356_new_n7126_), .Y(_abc_41356_new_n7132_));
OR2X2 OR2X2_2442 ( .A(_abc_41356_new_n7125_), .B(_abc_41356_new_n7133_), .Y(_0addr_15_0__4_));
OR2X2 OR2X2_2443 ( .A(_abc_41356_new_n7138_), .B(_abc_41356_new_n7137_), .Y(_abc_41356_new_n7139_));
OR2X2 OR2X2_2444 ( .A(_abc_41356_new_n7139_), .B(_abc_41356_new_n7140_), .Y(_abc_41356_new_n7141_));
OR2X2 OR2X2_2445 ( .A(_abc_41356_new_n7141_), .B(_abc_41356_new_n7136_), .Y(_abc_41356_new_n7142_));
OR2X2 OR2X2_2446 ( .A(_abc_41356_new_n7135_), .B(_abc_41356_new_n7143_), .Y(_0addr_15_0__5_));
OR2X2 OR2X2_2447 ( .A(_abc_41356_new_n7148_), .B(_abc_41356_new_n7147_), .Y(_abc_41356_new_n7149_));
OR2X2 OR2X2_2448 ( .A(_abc_41356_new_n7149_), .B(_abc_41356_new_n7150_), .Y(_abc_41356_new_n7151_));
OR2X2 OR2X2_2449 ( .A(_abc_41356_new_n7151_), .B(_abc_41356_new_n7146_), .Y(_abc_41356_new_n7152_));
OR2X2 OR2X2_245 ( .A(_abc_41356_new_n1357_), .B(_abc_41356_new_n1355_), .Y(_abc_41356_new_n1358_));
OR2X2 OR2X2_2450 ( .A(_abc_41356_new_n7145_), .B(_abc_41356_new_n7153_), .Y(_0addr_15_0__6_));
OR2X2 OR2X2_2451 ( .A(_abc_41356_new_n7158_), .B(_abc_41356_new_n7157_), .Y(_abc_41356_new_n7159_));
OR2X2 OR2X2_2452 ( .A(_abc_41356_new_n7159_), .B(_abc_41356_new_n7160_), .Y(_abc_41356_new_n7161_));
OR2X2 OR2X2_2453 ( .A(_abc_41356_new_n7161_), .B(_abc_41356_new_n7156_), .Y(_abc_41356_new_n7162_));
OR2X2 OR2X2_2454 ( .A(_abc_41356_new_n7155_), .B(_abc_41356_new_n7163_), .Y(_0addr_15_0__7_));
OR2X2 OR2X2_2455 ( .A(_abc_41356_new_n7168_), .B(_abc_41356_new_n7167_), .Y(_abc_41356_new_n7169_));
OR2X2 OR2X2_2456 ( .A(_abc_41356_new_n7169_), .B(_abc_41356_new_n7166_), .Y(_abc_41356_new_n7170_));
OR2X2 OR2X2_2457 ( .A(_abc_41356_new_n7165_), .B(_abc_41356_new_n7171_), .Y(_0addr_15_0__8_));
OR2X2 OR2X2_2458 ( .A(_abc_41356_new_n7176_), .B(_abc_41356_new_n7178_), .Y(_abc_41356_new_n7179_));
OR2X2 OR2X2_2459 ( .A(_abc_41356_new_n7179_), .B(_abc_41356_new_n7174_), .Y(_abc_41356_new_n7180_));
OR2X2 OR2X2_246 ( .A(_abc_41356_new_n1361_), .B(_abc_41356_new_n1355_), .Y(_abc_41356_new_n1362_));
OR2X2 OR2X2_2460 ( .A(_abc_41356_new_n7173_), .B(_abc_41356_new_n7180_), .Y(_0addr_15_0__9_));
OR2X2 OR2X2_2461 ( .A(_abc_41356_new_n7184_), .B(_abc_41356_new_n7186_), .Y(_abc_41356_new_n7187_));
OR2X2 OR2X2_2462 ( .A(_abc_41356_new_n7187_), .B(_abc_41356_new_n7183_), .Y(_abc_41356_new_n7188_));
OR2X2 OR2X2_2463 ( .A(_abc_41356_new_n7182_), .B(_abc_41356_new_n7188_), .Y(_0addr_15_0__10_));
OR2X2 OR2X2_2464 ( .A(_abc_41356_new_n7192_), .B(_abc_41356_new_n7194_), .Y(_abc_41356_new_n7195_));
OR2X2 OR2X2_2465 ( .A(_abc_41356_new_n7195_), .B(_abc_41356_new_n7191_), .Y(_abc_41356_new_n7196_));
OR2X2 OR2X2_2466 ( .A(_abc_41356_new_n7190_), .B(_abc_41356_new_n7196_), .Y(_0addr_15_0__11_));
OR2X2 OR2X2_2467 ( .A(_abc_41356_new_n7200_), .B(_abc_41356_new_n7201_), .Y(_abc_41356_new_n7202_));
OR2X2 OR2X2_2468 ( .A(_abc_41356_new_n7202_), .B(_abc_41356_new_n7199_), .Y(_abc_41356_new_n7203_));
OR2X2 OR2X2_2469 ( .A(_abc_41356_new_n7198_), .B(_abc_41356_new_n7204_), .Y(_0addr_15_0__12_));
OR2X2 OR2X2_247 ( .A(regfil_5__1_), .B(regfil_3__1_), .Y(_abc_41356_new_n1366_));
OR2X2 OR2X2_2470 ( .A(_abc_41356_new_n7208_), .B(_abc_41356_new_n7209_), .Y(_abc_41356_new_n7210_));
OR2X2 OR2X2_2471 ( .A(_abc_41356_new_n7210_), .B(_abc_41356_new_n7207_), .Y(_abc_41356_new_n7211_));
OR2X2 OR2X2_2472 ( .A(_abc_41356_new_n7206_), .B(_abc_41356_new_n7212_), .Y(_0addr_15_0__13_));
OR2X2 OR2X2_2473 ( .A(_abc_41356_new_n7217_), .B(_abc_41356_new_n7216_), .Y(_abc_41356_new_n7218_));
OR2X2 OR2X2_2474 ( .A(_abc_41356_new_n7218_), .B(_abc_41356_new_n7215_), .Y(_abc_41356_new_n7219_));
OR2X2 OR2X2_2475 ( .A(_abc_41356_new_n7214_), .B(_abc_41356_new_n7219_), .Y(_0addr_15_0__14_));
OR2X2 OR2X2_2476 ( .A(_abc_41356_new_n7222_), .B(_abc_41356_new_n7223_), .Y(_abc_41356_new_n7224_));
OR2X2 OR2X2_2477 ( .A(_abc_41356_new_n7224_), .B(_abc_41356_new_n4807_), .Y(_abc_41356_new_n7225_));
OR2X2 OR2X2_2478 ( .A(_abc_41356_new_n7221_), .B(_abc_41356_new_n7226_), .Y(_0addr_15_0__15_));
OR2X2 OR2X2_2479 ( .A(_abc_41356_new_n7232_), .B(_abc_41356_new_n7228_), .Y(_0readio_0_0_));
OR2X2 OR2X2_248 ( .A(_abc_41356_new_n1368_), .B(_abc_41356_new_n1363_), .Y(_abc_41356_new_n1369_));
OR2X2 OR2X2_2480 ( .A(_abc_41356_new_n7070_), .B(_abc_41356_new_n7235_), .Y(_abc_41356_new_n7236_));
OR2X2 OR2X2_2481 ( .A(_abc_41356_new_n7238_), .B(inta), .Y(_abc_41356_new_n7239_));
OR2X2 OR2X2_2482 ( .A(_abc_41356_new_n7239_), .B(_abc_41356_new_n7237_), .Y(_abc_41356_new_n7240_));
OR2X2 OR2X2_2483 ( .A(_abc_41356_new_n7245_), .B(waitr), .Y(_abc_41356_new_n7246_));
OR2X2 OR2X2_2484 ( .A(_abc_41356_new_n7248_), .B(_abc_41356_new_n7243_), .Y(_0writeio_0_0_));
OR2X2 OR2X2_2485 ( .A(_abc_41356_new_n7253_), .B(_abc_41356_new_n7255_), .Y(_abc_41356_new_n7256_));
OR2X2 OR2X2_2486 ( .A(_abc_41356_new_n7256_), .B(_abc_41356_new_n3555_), .Y(_abc_41356_new_n7257_));
OR2X2 OR2X2_2487 ( .A(_abc_41356_new_n7257_), .B(_abc_41356_new_n7252_), .Y(_abc_41356_new_n7258_));
OR2X2 OR2X2_2488 ( .A(_abc_41356_new_n3555_), .B(_abc_41356_new_n7266_), .Y(_abc_41356_new_n7267_));
OR2X2 OR2X2_2489 ( .A(_abc_41356_new_n7265_), .B(_abc_41356_new_n7267_), .Y(_abc_41356_new_n7268_));
OR2X2 OR2X2_249 ( .A(_abc_41356_new_n1371_), .B(_abc_41356_new_n1360_), .Y(_abc_41356_new_n1372_));
OR2X2 OR2X2_2490 ( .A(_abc_41356_new_n7278_), .B(_abc_41356_new_n7273_), .Y(_abc_41356_new_n7279_));
OR2X2 OR2X2_2491 ( .A(_abc_41356_new_n7279_), .B(_abc_41356_new_n3609_), .Y(_abc_41356_new_n7280_));
OR2X2 OR2X2_2492 ( .A(_abc_41356_new_n7280_), .B(_abc_41356_new_n7269_), .Y(_abc_41356_new_n7281_));
OR2X2 OR2X2_2493 ( .A(_abc_41356_new_n7281_), .B(_abc_41356_new_n7259_), .Y(_abc_41356_new_n7282_));
OR2X2 OR2X2_2494 ( .A(_abc_41356_new_n2048_), .B(_abc_41356_new_n3779_), .Y(_abc_41356_new_n7289_));
OR2X2 OR2X2_2495 ( .A(_abc_41356_new_n3495_), .B(_abc_41356_new_n7289_), .Y(_abc_41356_new_n7290_));
OR2X2 OR2X2_2496 ( .A(_abc_41356_new_n3368_), .B(_abc_41356_new_n619_), .Y(_abc_41356_new_n7293_));
OR2X2 OR2X2_2497 ( .A(_abc_41356_new_n4151_), .B(_abc_41356_new_n7299_), .Y(_abc_41356_new_n7300_));
OR2X2 OR2X2_2498 ( .A(_abc_41356_new_n7301_), .B(_abc_41356_new_n7296_), .Y(_abc_41356_new_n7302_));
OR2X2 OR2X2_2499 ( .A(_abc_41356_new_n545_), .B(zero), .Y(_abc_41356_new_n7305_));
OR2X2 OR2X2_25 ( .A(_abc_41356_new_n658_), .B(_abc_41356_new_n659_), .Y(_abc_41356_new_n660_));
OR2X2 OR2X2_250 ( .A(_abc_41356_new_n1375_), .B(_abc_41356_new_n1362_), .Y(_abc_41356_new_n1376_));
OR2X2 OR2X2_2500 ( .A(_abc_41356_new_n7307_), .B(_abc_41356_new_n7308_), .Y(_abc_41356_new_n7309_));
OR2X2 OR2X2_2501 ( .A(_abc_41356_new_n7311_), .B(_abc_41356_new_n7294_), .Y(_abc_41356_new_n7312_));
OR2X2 OR2X2_2502 ( .A(_abc_41356_new_n7313_), .B(_abc_41356_new_n7288_), .Y(_abc_41356_new_n7314_));
OR2X2 OR2X2_2503 ( .A(_abc_41356_new_n3366_), .B(parity), .Y(_abc_41356_new_n7319_));
OR2X2 OR2X2_2504 ( .A(_abc_41356_new_n4161_), .B(_abc_41356_new_n7320_), .Y(_abc_41356_new_n7321_));
OR2X2 OR2X2_2505 ( .A(_abc_41356_new_n7325_), .B(_abc_41356_new_n7317_), .Y(_abc_41356_new_n7326_));
OR2X2 OR2X2_2506 ( .A(_abc_41356_new_n7326_), .B(_abc_41356_new_n7315_), .Y(_abc_41356_new_n7327_));
OR2X2 OR2X2_2507 ( .A(_abc_41356_new_n7330_), .B(_abc_41356_new_n3265_), .Y(_abc_41356_new_n7331_));
OR2X2 OR2X2_2508 ( .A(_abc_41356_new_n7333_), .B(_abc_41356_new_n3265_), .Y(_abc_41356_new_n7334_));
OR2X2 OR2X2_2509 ( .A(_abc_41356_new_n7335_), .B(reset), .Y(_abc_41356_new_n7336_));
OR2X2 OR2X2_251 ( .A(regfil_5__7_), .B(regfil_3__7_), .Y(_abc_41356_new_n1379_));
OR2X2 OR2X2_2510 ( .A(_abc_41356_new_n7263_), .B(_abc_41356_new_n3488_), .Y(_abc_41356_new_n7339_));
OR2X2 OR2X2_2511 ( .A(_abc_41356_new_n7338_), .B(_abc_41356_new_n7339_), .Y(_abc_41356_new_n7340_));
OR2X2 OR2X2_2512 ( .A(_abc_41356_new_n7344_), .B(_abc_41356_new_n7342_), .Y(_abc_41356_new_n7345_));
OR2X2 OR2X2_2513 ( .A(_abc_41356_new_n7347_), .B(_abc_41356_new_n7263_), .Y(_abc_41356_new_n7348_));
OR2X2 OR2X2_2514 ( .A(_abc_41356_new_n7348_), .B(_abc_41356_new_n7346_), .Y(_abc_41356_new_n7349_));
OR2X2 OR2X2_2515 ( .A(_abc_41356_new_n3453_), .B(_abc_41356_new_n7350_), .Y(_abc_41356_new_n7351_));
OR2X2 OR2X2_2516 ( .A(_abc_41356_new_n7360_), .B(_abc_41356_new_n7362_), .Y(_abc_41356_new_n7363_));
OR2X2 OR2X2_2517 ( .A(_abc_41356_new_n7338_), .B(_abc_41356_new_n7348_), .Y(_abc_41356_new_n7364_));
OR2X2 OR2X2_2518 ( .A(_abc_41356_new_n3446_), .B(_abc_41356_new_n7372_), .Y(_abc_41356_new_n7373_));
OR2X2 OR2X2_2519 ( .A(_abc_41356_new_n7384_), .B(statesel_5_), .Y(_abc_41356_new_n7385_));
OR2X2 OR2X2_252 ( .A(regfil_5__6_), .B(regfil_3__6_), .Y(_abc_41356_new_n1383_));
OR2X2 OR2X2_2520 ( .A(_abc_41356_new_n7385_), .B(_abc_41356_new_n7381_), .Y(_abc_41356_new_n7386_));
OR2X2 OR2X2_2521 ( .A(_abc_41356_new_n7390_), .B(_abc_41356_new_n7387_), .Y(_abc_41356_new_n7391_));
OR2X2 OR2X2_2522 ( .A(_abc_41356_new_n7393_), .B(_abc_41356_new_n7342_), .Y(_abc_41356_new_n7394_));
OR2X2 OR2X2_2523 ( .A(_abc_41356_new_n3453_), .B(_abc_41356_new_n7396_), .Y(_abc_41356_new_n7397_));
OR2X2 OR2X2_2524 ( .A(_abc_41356_new_n3363_), .B(_abc_41356_new_n7288_), .Y(_abc_41356_new_n7398_));
OR2X2 OR2X2_2525 ( .A(_abc_41356_new_n3475_), .B(_abc_41356_new_n7399_), .Y(_abc_41356_new_n7400_));
OR2X2 OR2X2_2526 ( .A(_abc_41356_new_n4827_), .B(_abc_41356_new_n7401_), .Y(_abc_41356_new_n7402_));
OR2X2 OR2X2_2527 ( .A(_abc_41356_new_n7404_), .B(_abc_41356_new_n3265_), .Y(_abc_41356_new_n7405_));
OR2X2 OR2X2_2528 ( .A(_abc_41356_new_n7411_), .B(_abc_41356_new_n7409_), .Y(_abc_41356_new_n7412_));
OR2X2 OR2X2_2529 ( .A(_abc_41356_new_n7416_), .B(_abc_41356_new_n7417_), .Y(_abc_41356_new_n7418_));
OR2X2 OR2X2_253 ( .A(regfil_5__5_), .B(regfil_3__5_), .Y(_abc_41356_new_n1388_));
OR2X2 OR2X2_2530 ( .A(_abc_41356_new_n7420_), .B(_abc_41356_new_n7392_), .Y(_abc_41356_new_n7421_));
OR2X2 OR2X2_2531 ( .A(_abc_41356_new_n7424_), .B(_abc_41356_new_n7426_), .Y(_abc_41356_new_n7427_));
OR2X2 OR2X2_2532 ( .A(_abc_41356_new_n7430_), .B(_abc_41356_new_n7057_), .Y(_abc_41356_new_n7431_));
OR2X2 OR2X2_2533 ( .A(_abc_41356_new_n7338_), .B(_abc_41356_new_n7380_), .Y(_abc_41356_new_n7440_));
OR2X2 OR2X2_2534 ( .A(_abc_41356_new_n3265_), .B(_abc_41356_new_n7442_), .Y(_abc_41356_new_n7443_));
OR2X2 OR2X2_2535 ( .A(_abc_41356_new_n7443_), .B(_abc_41356_new_n7441_), .Y(_abc_41356_new_n7444_));
OR2X2 OR2X2_2536 ( .A(_abc_41356_new_n7451_), .B(_abc_41356_new_n7446_), .Y(_abc_41356_new_n7452_));
OR2X2 OR2X2_2537 ( .A(_abc_41356_new_n3453_), .B(_abc_41356_new_n7452_), .Y(_abc_41356_new_n7453_));
OR2X2 OR2X2_2538 ( .A(_abc_41356_new_n7455_), .B(_abc_41356_new_n7243_), .Y(_abc_41356_new_n7456_));
OR2X2 OR2X2_2539 ( .A(_abc_41356_new_n7420_), .B(_abc_41356_new_n7450_), .Y(_abc_41356_new_n7461_));
OR2X2 OR2X2_254 ( .A(regfil_5__4_), .B(regfil_3__4_), .Y(_abc_41356_new_n1392_));
OR2X2 OR2X2_2540 ( .A(_abc_41356_new_n7064_), .B(_abc_41356_new_n7462_), .Y(_abc_41356_new_n7463_));
OR2X2 OR2X2_2541 ( .A(_abc_41356_new_n7447_), .B(_abc_41356_new_n3581_), .Y(_abc_41356_new_n7479_));
OR2X2 OR2X2_2542 ( .A(_abc_41356_new_n7480_), .B(_abc_41356_new_n7482_), .Y(_abc_41356_new_n7483_));
OR2X2 OR2X2_2543 ( .A(_abc_41356_new_n7485_), .B(_abc_41356_new_n7387_), .Y(_abc_41356_new_n7486_));
OR2X2 OR2X2_2544 ( .A(_abc_41356_new_n3453_), .B(_abc_41356_new_n7490_), .Y(_abc_41356_new_n7491_));
OR2X2 OR2X2_2545 ( .A(_abc_41356_new_n3203_), .B(_abc_41356_new_n7498_), .Y(_abc_41356_new_n7499_));
OR2X2 OR2X2_2546 ( .A(_abc_41356_new_n7500_), .B(reset), .Y(_abc_41356_new_n7501_));
OR2X2 OR2X2_2547 ( .A(_abc_41356_new_n7512_), .B(_abc_41356_new_n7513_), .Y(_abc_41356_new_n7514_));
OR2X2 OR2X2_2548 ( .A(_abc_41356_new_n7431_), .B(_abc_41356_new_n7418_), .Y(_abc_41356_new_n7529_));
OR2X2 OR2X2_2549 ( .A(_abc_41356_new_n7529_), .B(_abc_41356_new_n7373_), .Y(_abc_41356_new_n7530_));
OR2X2 OR2X2_255 ( .A(_abc_41356_new_n1386_), .B(_abc_41356_new_n1390_), .Y(_abc_41356_new_n1397_));
OR2X2 OR2X2_2550 ( .A(_abc_41356_new_n7456_), .B(_abc_41356_new_n4241_), .Y(_abc_41356_new_n7532_));
OR2X2 OR2X2_2551 ( .A(_abc_41356_new_n7533_), .B(_abc_41356_new_n5413_), .Y(_abc_41356_new_n7534_));
OR2X2 OR2X2_2552 ( .A(_abc_41356_new_n7532_), .B(_abc_41356_new_n7534_), .Y(_abc_41356_new_n7535_));
OR2X2 OR2X2_2553 ( .A(_abc_41356_new_n7535_), .B(_abc_41356_new_n7531_), .Y(_abc_41356_new_n7536_));
OR2X2 OR2X2_2554 ( .A(_abc_41356_new_n7536_), .B(_abc_41356_new_n7530_), .Y(_abc_41356_new_n7537_));
OR2X2 OR2X2_2555 ( .A(_abc_41356_new_n7528_), .B(_abc_41356_new_n7537_), .Y(_abc_41356_new_n7538_));
OR2X2 OR2X2_2556 ( .A(_abc_41356_new_n7538_), .B(_abc_41356_new_n7527_), .Y(_abc_41356_new_n7539_));
OR2X2 OR2X2_2557 ( .A(_abc_41356_new_n7515_), .B(_abc_41356_new_n7492_), .Y(_abc_41356_new_n7540_));
OR2X2 OR2X2_2558 ( .A(_abc_41356_new_n7539_), .B(_abc_41356_new_n7540_), .Y(_abc_41356_new_n7541_));
OR2X2 OR2X2_2559 ( .A(_abc_41356_new_n7542_), .B(_abc_41356_new_n7412_), .Y(_abc_41356_new_n7543_));
OR2X2 OR2X2_256 ( .A(_abc_41356_new_n1400_), .B(_abc_41356_new_n1377_), .Y(_abc_41356_new_n1401_));
OR2X2 OR2X2_2560 ( .A(_abc_41356_new_n7541_), .B(_abc_41356_new_n7543_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_4_));
OR2X2 OR2X2_2561 ( .A(_abc_41356_new_n7428_), .B(_abc_41356_new_n550_), .Y(_abc_41356_new_n7546_));
OR2X2 OR2X2_2562 ( .A(_abc_41356_new_n7546_), .B(_abc_41356_new_n7545_), .Y(_abc_41356_new_n7547_));
OR2X2 OR2X2_2563 ( .A(_abc_41356_new_n7382_), .B(_abc_41356_new_n7254_), .Y(_abc_41356_new_n7548_));
OR2X2 OR2X2_2564 ( .A(_abc_41356_new_n7459_), .B(_abc_41356_new_n7477_), .Y(_abc_41356_new_n7551_));
OR2X2 OR2X2_2565 ( .A(_abc_41356_new_n7551_), .B(_abc_41356_new_n7550_), .Y(_abc_41356_new_n7552_));
OR2X2 OR2X2_2566 ( .A(_abc_41356_new_n7552_), .B(_abc_41356_new_n7547_), .Y(_abc_36060_auto_fsm_map_cc_170_map_fsm_12881_5_));
OR2X2 OR2X2_2567 ( .A(_abc_41356_new_n7555_), .B(_abc_41356_new_n6533_), .Y(_abc_41356_new_n7556_));
OR2X2 OR2X2_2568 ( .A(_abc_41356_new_n7559_), .B(eienb), .Y(_abc_41356_new_n7560_));
OR2X2 OR2X2_2569 ( .A(_abc_41356_new_n7561_), .B(reset), .Y(_abc_41356_new_n7562_));
OR2X2 OR2X2_257 ( .A(_abc_41356_new_n1399_), .B(_abc_41356_new_n1401_), .Y(_abc_41356_new_n1402_));
OR2X2 OR2X2_2570 ( .A(_abc_41356_new_n7557_), .B(_abc_41356_new_n7562_), .Y(_0ei_0_0_));
OR2X2 OR2X2_2571 ( .A(alu_oprb_7_), .B(alu_opra_7_), .Y(alu__abc_40887_new_n33_));
OR2X2 OR2X2_2572 ( .A(alu_oprb_1_), .B(alu_opra_1_), .Y(alu__abc_40887_new_n48_));
OR2X2 OR2X2_2573 ( .A(alu__abc_40887_new_n51_), .B(alu__abc_40887_new_n46_), .Y(alu__abc_40887_new_n52_));
OR2X2 OR2X2_2574 ( .A(alu_oprb_3_), .B(alu_opra_3_), .Y(alu__abc_40887_new_n62_));
OR2X2 OR2X2_2575 ( .A(alu__abc_40887_new_n66_), .B(alu__abc_40887_new_n60_), .Y(alu__abc_40887_new_n67_));
OR2X2 OR2X2_2576 ( .A(alu__abc_40887_new_n65_), .B(alu__abc_40887_new_n67_), .Y(alu__abc_40887_new_n68_));
OR2X2 OR2X2_2577 ( .A(alu__abc_40887_new_n89_), .B(alu__abc_40887_new_n45_), .Y(alu__abc_40887_new_n90_));
OR2X2 OR2X2_2578 ( .A(alu__abc_40887_new_n93_), .B(alu__abc_40887_new_n94_), .Y(alu__abc_40887_new_n95_));
OR2X2 OR2X2_2579 ( .A(alu__abc_40887_new_n97_), .B(alu__abc_40887_new_n98_), .Y(alu__abc_40887_new_n99_));
OR2X2 OR2X2_258 ( .A(_abc_41356_new_n1396_), .B(_abc_41356_new_n1402_), .Y(_abc_41356_new_n1403_));
OR2X2 OR2X2_2580 ( .A(alu__abc_40887_new_n109_), .B(alu__abc_40887_new_n53_), .Y(alu__abc_40887_new_n110_));
OR2X2 OR2X2_2581 ( .A(alu__abc_40887_new_n110_), .B(alu__abc_40887_new_n63_), .Y(alu__abc_40887_new_n113_));
OR2X2 OR2X2_2582 ( .A(alu__abc_40887_new_n52_), .B(alu__abc_40887_new_n59_), .Y(alu__abc_40887_new_n124_));
OR2X2 OR2X2_2583 ( .A(alu__abc_40887_new_n68_), .B(alu__abc_40887_new_n75_), .Y(alu__abc_40887_new_n128_));
OR2X2 OR2X2_2584 ( .A(alu__abc_40887_new_n140_), .B(alu__abc_40887_new_n139_), .Y(alu__abc_40887_new_n141_));
OR2X2 OR2X2_2585 ( .A(alu__abc_40887_new_n141_), .B(alu__abc_40887_new_n134_), .Y(alu__abc_40887_new_n142_));
OR2X2 OR2X2_2586 ( .A(alu__abc_40887_new_n150_), .B(alu__abc_40887_new_n147_), .Y(alu__abc_40887_new_n151_));
OR2X2 OR2X2_2587 ( .A(alu__abc_40887_new_n49_), .B(alu__abc_40887_new_n156_), .Y(alu__abc_40887_new_n157_));
OR2X2 OR2X2_2588 ( .A(alu__abc_40887_new_n59_), .B(alu__abc_40887_new_n63_), .Y(alu__abc_40887_new_n159_));
OR2X2 OR2X2_2589 ( .A(alu__abc_40887_new_n158_), .B(alu__abc_40887_new_n159_), .Y(alu__abc_40887_new_n160_));
OR2X2 OR2X2_259 ( .A(_abc_41356_new_n1406_), .B(_abc_41356_new_n1407_), .Y(_abc_41356_new_n1408_));
OR2X2 OR2X2_2590 ( .A(alu__abc_40887_new_n75_), .B(alu__abc_40887_new_n82_), .Y(alu__abc_40887_new_n162_));
OR2X2 OR2X2_2591 ( .A(alu__abc_40887_new_n161_), .B(alu__abc_40887_new_n162_), .Y(alu__abc_40887_new_n163_));
OR2X2 OR2X2_2592 ( .A(alu__abc_40887_new_n165_), .B(alu__abc_40887_new_n166_), .Y(alu__abc_40887_new_n167_));
OR2X2 OR2X2_2593 ( .A(alu__abc_40887_new_n169_), .B(alu__abc_40887_new_n44_), .Y(alu__abc_40887_new_n170_));
OR2X2 OR2X2_2594 ( .A(alu__abc_40887_new_n173_), .B(alu__abc_40887_new_n36_), .Y(alu__abc_40887_new_n174_));
OR2X2 OR2X2_2595 ( .A(alu__abc_40887_new_n185_), .B(alu__abc_40887_new_n46_), .Y(alu__abc_40887_new_n186_));
OR2X2 OR2X2_2596 ( .A(alu__abc_40887_new_n188_), .B(alu__abc_40887_new_n154_), .Y(alu__abc_40887_new_n189_));
OR2X2 OR2X2_2597 ( .A(alu__abc_40887_new_n192_), .B(alu__abc_40887_new_n151_), .Y(alu__abc_40887_new_n193_));
OR2X2 OR2X2_2598 ( .A(alu__abc_40887_new_n103_), .B(alu__abc_40887_new_n164_), .Y(alu__abc_40887_new_n195_));
OR2X2 OR2X2_2599 ( .A(alu__abc_40887_new_n194_), .B(alu__abc_40887_new_n195_), .Y(alu__abc_40887_new_n196_));
OR2X2 OR2X2_26 ( .A(_abc_41356_new_n661_), .B(_abc_41356_new_n643_), .Y(_abc_41356_new_n662_));
OR2X2 OR2X2_260 ( .A(_abc_41356_new_n1404_), .B(_abc_41356_new_n1408_), .Y(_abc_41356_new_n1409_));
OR2X2 OR2X2_2600 ( .A(alu__abc_40887_new_n194_), .B(alu__abc_40887_new_n201_), .Y(alu__abc_40887_new_n202_));
OR2X2 OR2X2_2601 ( .A(alu__abc_40887_new_n203_), .B(alu__abc_40887_new_n149_), .Y(alu__abc_40887_new_n204_));
OR2X2 OR2X2_2602 ( .A(alu__abc_40887_new_n158_), .B(alu__abc_40887_new_n59_), .Y(alu__abc_40887_new_n206_));
OR2X2 OR2X2_2603 ( .A(alu__abc_40887_new_n205_), .B(alu__abc_40887_new_n209_), .Y(alu__abc_40887_new_n210_));
OR2X2 OR2X2_2604 ( .A(alu__abc_40887_new_n203_), .B(alu__abc_40887_new_n211_), .Y(alu__abc_40887_new_n212_));
OR2X2 OR2X2_2605 ( .A(alu__abc_40887_new_n120_), .B(alu__abc_40887_new_n213_), .Y(alu__abc_40887_new_n214_));
OR2X2 OR2X2_2606 ( .A(alu__abc_40887_new_n188_), .B(alu__abc_40887_new_n215_), .Y(alu__abc_40887_new_n216_));
OR2X2 OR2X2_2607 ( .A(alu__abc_40887_new_n217_), .B(alu__abc_40887_new_n214_), .Y(alu__abc_40887_new_n218_));
OR2X2 OR2X2_2608 ( .A(alu__abc_40887_new_n225_), .B(alu__abc_40887_new_n227_), .Y(alu__abc_40887_new_n228_));
OR2X2 OR2X2_2609 ( .A(alu__abc_40887_new_n235_), .B(alu__abc_40887_new_n236_), .Y(alu__abc_40887_new_n237_));
OR2X2 OR2X2_261 ( .A(_abc_41356_new_n1403_), .B(_abc_41356_new_n1410_), .Y(_abc_41356_new_n1411_));
OR2X2 OR2X2_2610 ( .A(alu__abc_40887_new_n242_), .B(alu__abc_40887_new_n244_), .Y(alu__abc_40887_new_n245_));
OR2X2 OR2X2_2611 ( .A(alu__abc_40887_new_n245_), .B(alu__abc_40887_new_n240_), .Y(alu__abc_40887_new_n246_));
OR2X2 OR2X2_2612 ( .A(alu__abc_40887_new_n238_), .B(alu__abc_40887_new_n246_), .Y(alu__abc_40887_new_n247_));
OR2X2 OR2X2_2613 ( .A(alu__abc_40887_new_n247_), .B(alu__abc_40887_new_n233_), .Y(alu__abc_40887_new_n248_));
OR2X2 OR2X2_2614 ( .A(alu__abc_40887_new_n229_), .B(alu__abc_40887_new_n248_), .Y(alu__abc_40887_new_n249_));
OR2X2 OR2X2_2615 ( .A(alu__abc_40887_new_n249_), .B(alu__abc_40887_new_n143_), .Y(alu_sout));
OR2X2 OR2X2_2616 ( .A(alu__abc_40887_new_n208_), .B(alu__abc_40887_new_n63_), .Y(alu__abc_40887_new_n256_));
OR2X2 OR2X2_2617 ( .A(alu__abc_40887_new_n204_), .B(alu__abc_40887_new_n148_), .Y(alu__abc_40887_new_n257_));
OR2X2 OR2X2_2618 ( .A(alu__abc_40887_new_n258_), .B(alu__abc_40887_new_n259_), .Y(alu__abc_40887_new_n260_));
OR2X2 OR2X2_2619 ( .A(alu__abc_40887_new_n199_), .B(alu__abc_40887_new_n261_), .Y(alu__abc_40887_new_n262_));
OR2X2 OR2X2_262 ( .A(_abc_41356_new_n1423_), .B(_abc_41356_new_n1419_), .Y(_abc_41356_new_n1424_));
OR2X2 OR2X2_2620 ( .A(alu__abc_40887_new_n262_), .B(alu__abc_40887_new_n260_), .Y(alu__abc_40887_new_n263_));
OR2X2 OR2X2_2621 ( .A(alu__abc_40887_new_n264_), .B(alu__abc_40887_new_n224_), .Y(alu__abc_40887_new_n265_));
OR2X2 OR2X2_2622 ( .A(alu__abc_40887_new_n271_), .B(alu__abc_40887_new_n270_), .Y(alu__abc_40887_new_n272_));
OR2X2 OR2X2_2623 ( .A(alu__abc_40887_new_n272_), .B(alu__abc_40887_new_n269_), .Y(alu__abc_40887_new_n273_));
OR2X2 OR2X2_2624 ( .A(alu__abc_40887_new_n268_), .B(alu__abc_40887_new_n273_), .Y(alu__abc_40887_new_n274_));
OR2X2 OR2X2_2625 ( .A(alu__abc_40887_new_n267_), .B(alu__abc_40887_new_n274_), .Y(alu__abc_40887_new_n275_));
OR2X2 OR2X2_2626 ( .A(alu__abc_40887_new_n266_), .B(alu__abc_40887_new_n275_), .Y(alu__abc_40887_new_n276_));
OR2X2 OR2X2_2627 ( .A(alu__abc_40887_new_n276_), .B(alu__abc_40887_new_n255_), .Y(alu__abc_40887_new_n277_));
OR2X2 OR2X2_2628 ( .A(alu_sout), .B(alu__abc_40887_new_n277_), .Y(alu__abc_40887_new_n278_));
OR2X2 OR2X2_2629 ( .A(alu__abc_40887_new_n226_), .B(alu__abc_40887_new_n177_), .Y(alu__abc_40887_new_n280_));
OR2X2 OR2X2_263 ( .A(_abc_41356_new_n1424_), .B(_abc_41356_new_n1422_), .Y(_abc_41356_new_n1425_));
OR2X2 OR2X2_2630 ( .A(alu__abc_40887_new_n282_), .B(alu__abc_40887_new_n279_), .Y(alu__abc_40887_new_n283_));
OR2X2 OR2X2_2631 ( .A(alu__abc_40887_new_n286_), .B(alu__abc_40887_new_n287_), .Y(alu__abc_40887_new_n288_));
OR2X2 OR2X2_2632 ( .A(alu__abc_40887_new_n290_), .B(alu__abc_40887_new_n51_), .Y(alu__abc_40887_new_n291_));
OR2X2 OR2X2_2633 ( .A(alu__abc_40887_new_n219_), .B(alu__abc_40887_new_n294_), .Y(alu__abc_40887_new_n295_));
OR2X2 OR2X2_2634 ( .A(alu__abc_40887_new_n232_), .B(alu__abc_40887_new_n306_), .Y(alu__abc_40887_new_n307_));
OR2X2 OR2X2_2635 ( .A(alu__abc_40887_new_n307_), .B(alu__abc_40887_new_n305_), .Y(alu__abc_40887_new_n308_));
OR2X2 OR2X2_2636 ( .A(alu__abc_40887_new_n308_), .B(alu__abc_40887_new_n304_), .Y(alu__abc_40887_new_n309_));
OR2X2 OR2X2_2637 ( .A(alu__abc_40887_new_n303_), .B(alu__abc_40887_new_n309_), .Y(alu__abc_40887_new_n310_));
OR2X2 OR2X2_2638 ( .A(alu__abc_40887_new_n302_), .B(alu__abc_40887_new_n310_), .Y(alu__abc_40887_new_n311_));
OR2X2 OR2X2_2639 ( .A(alu__abc_40887_new_n296_), .B(alu__abc_40887_new_n311_), .Y(alu__abc_40887_new_n312_));
OR2X2 OR2X2_264 ( .A(_abc_41356_new_n1428_), .B(_abc_41356_new_n1427_), .Y(_abc_41356_new_n1429_));
OR2X2 OR2X2_2640 ( .A(alu__abc_40887_new_n319_), .B(alu__abc_40887_new_n314_), .Y(alu__abc_40887_new_n320_));
OR2X2 OR2X2_2641 ( .A(alu__abc_40887_new_n121_), .B(alu__abc_40887_new_n322_), .Y(alu__abc_40887_new_n323_));
OR2X2 OR2X2_2642 ( .A(alu__abc_40887_new_n323_), .B(alu__abc_40887_new_n321_), .Y(alu__abc_40887_new_n324_));
OR2X2 OR2X2_2643 ( .A(alu__abc_40887_new_n325_), .B(alu__abc_40887_new_n326_), .Y(alu__abc_40887_new_n327_));
OR2X2 OR2X2_2644 ( .A(alu__abc_40887_new_n313_), .B(alu__abc_40887_new_n331_), .Y(alu__abc_40887_new_n333_));
OR2X2 OR2X2_2645 ( .A(alu__abc_40887_new_n334_), .B(alu__abc_40887_new_n332_), .Y(alu__abc_40887_new_n335_));
OR2X2 OR2X2_2646 ( .A(alu__abc_40887_new_n337_), .B(alu__abc_40887_new_n111_), .Y(alu__abc_40887_new_n338_));
OR2X2 OR2X2_2647 ( .A(alu__abc_40887_new_n221_), .B(alu__abc_40887_new_n345_), .Y(alu__abc_40887_new_n346_));
OR2X2 OR2X2_2648 ( .A(alu__abc_40887_new_n351_), .B(alu__abc_40887_new_n352_), .Y(alu__abc_40887_new_n353_));
OR2X2 OR2X2_2649 ( .A(alu__abc_40887_new_n353_), .B(alu__abc_40887_new_n350_), .Y(alu__abc_40887_new_n354_));
OR2X2 OR2X2_265 ( .A(_abc_41356_new_n1432_), .B(_abc_41356_new_n1431_), .Y(_abc_41356_new_n1433_));
OR2X2 OR2X2_2650 ( .A(alu__abc_40887_new_n349_), .B(alu__abc_40887_new_n354_), .Y(alu__abc_40887_new_n355_));
OR2X2 OR2X2_2651 ( .A(alu__abc_40887_new_n355_), .B(alu__abc_40887_new_n348_), .Y(alu__abc_40887_new_n356_));
OR2X2 OR2X2_2652 ( .A(alu__abc_40887_new_n356_), .B(alu__abc_40887_new_n347_), .Y(alu__abc_40887_new_n357_));
OR2X2 OR2X2_2653 ( .A(alu__abc_40887_new_n357_), .B(alu__abc_40887_new_n344_), .Y(alu__abc_40887_new_n358_));
OR2X2 OR2X2_2654 ( .A(alu__abc_40887_new_n360_), .B(alu__abc_40887_new_n220_), .Y(alu__abc_40887_new_n361_));
OR2X2 OR2X2_2655 ( .A(alu__abc_40887_new_n372_), .B(alu__abc_40887_new_n371_), .Y(alu__abc_40887_new_n373_));
OR2X2 OR2X2_2656 ( .A(alu__abc_40887_new_n373_), .B(alu__abc_40887_new_n370_), .Y(alu__abc_40887_new_n374_));
OR2X2 OR2X2_2657 ( .A(alu__abc_40887_new_n369_), .B(alu__abc_40887_new_n374_), .Y(alu__abc_40887_new_n375_));
OR2X2 OR2X2_2658 ( .A(alu__abc_40887_new_n375_), .B(alu__abc_40887_new_n368_), .Y(alu__abc_40887_new_n376_));
OR2X2 OR2X2_2659 ( .A(alu__abc_40887_new_n367_), .B(alu__abc_40887_new_n376_), .Y(alu__abc_40887_new_n377_));
OR2X2 OR2X2_266 ( .A(_abc_41356_new_n1436_), .B(_abc_41356_new_n1426_), .Y(_abc_41356_new_n1437_));
OR2X2 OR2X2_2660 ( .A(alu__abc_40887_new_n377_), .B(alu__abc_40887_new_n362_), .Y(alu__abc_40887_new_n378_));
OR2X2 OR2X2_2661 ( .A(alu__abc_40887_new_n358_), .B(alu__abc_40887_new_n378_), .Y(alu__abc_40887_new_n379_));
OR2X2 OR2X2_2662 ( .A(alu__abc_40887_new_n380_), .B(alu__abc_40887_new_n381_), .Y(alu__abc_40887_new_n382_));
OR2X2 OR2X2_2663 ( .A(alu__abc_40887_new_n382_), .B(alu__abc_40887_new_n336_), .Y(alu__abc_40887_new_n383_));
OR2X2 OR2X2_2664 ( .A(alu__abc_40887_new_n385_), .B(alu__abc_40887_new_n335_), .Y(alu__abc_40887_new_n386_));
OR2X2 OR2X2_2665 ( .A(alu__abc_40887_new_n130_), .B(alu__abc_40887_new_n108_), .Y(alu__abc_40887_new_n388_));
OR2X2 OR2X2_2666 ( .A(alu__abc_40887_new_n131_), .B(alu__abc_40887_new_n139_), .Y(alu__abc_40887_new_n390_));
OR2X2 OR2X2_2667 ( .A(alu__abc_40887_new_n390_), .B(alu__abc_40887_new_n389_), .Y(alu__abc_40887_new_n391_));
OR2X2 OR2X2_2668 ( .A(alu__abc_40887_new_n260_), .B(alu__abc_40887_new_n261_), .Y(alu__abc_40887_new_n393_));
OR2X2 OR2X2_2669 ( .A(alu__abc_40887_new_n394_), .B(alu__abc_40887_new_n223_), .Y(alu__abc_40887_new_n395_));
OR2X2 OR2X2_267 ( .A(_abc_41356_new_n1439_), .B(_abc_41356_new_n1427_), .Y(_abc_41356_new_n1440_));
OR2X2 OR2X2_2670 ( .A(alu__abc_40887_new_n398_), .B(alu__abc_40887_new_n399_), .Y(alu__abc_40887_new_n400_));
OR2X2 OR2X2_2671 ( .A(alu__abc_40887_new_n401_), .B(alu__abc_40887_new_n232_), .Y(alu__abc_40887_new_n402_));
OR2X2 OR2X2_2672 ( .A(alu__abc_40887_new_n400_), .B(alu__abc_40887_new_n402_), .Y(alu__abc_40887_new_n403_));
OR2X2 OR2X2_2673 ( .A(alu__abc_40887_new_n397_), .B(alu__abc_40887_new_n403_), .Y(alu__abc_40887_new_n404_));
OR2X2 OR2X2_2674 ( .A(alu__abc_40887_new_n396_), .B(alu__abc_40887_new_n404_), .Y(alu__abc_40887_new_n405_));
OR2X2 OR2X2_2675 ( .A(alu__abc_40887_new_n405_), .B(alu__abc_40887_new_n392_), .Y(alu__abc_40887_new_n406_));
OR2X2 OR2X2_2676 ( .A(alu__abc_40887_new_n130_), .B(alu__abc_40887_new_n139_), .Y(alu__abc_40887_new_n413_));
OR2X2 OR2X2_2677 ( .A(alu__abc_40887_new_n413_), .B(alu__abc_40887_new_n412_), .Y(alu__abc_40887_new_n414_));
OR2X2 OR2X2_2678 ( .A(alu__abc_40887_new_n415_), .B(alu__abc_40887_new_n222_), .Y(alu__abc_40887_new_n416_));
OR2X2 OR2X2_2679 ( .A(alu__abc_40887_new_n420_), .B(alu__abc_40887_new_n421_), .Y(alu__abc_40887_new_n422_));
OR2X2 OR2X2_268 ( .A(regfil_1__7_), .B(regfil_5__7_), .Y(_abc_41356_new_n1445_));
OR2X2 OR2X2_2680 ( .A(alu__abc_40887_new_n422_), .B(alu__abc_40887_new_n423_), .Y(alu__abc_40887_new_n424_));
OR2X2 OR2X2_2681 ( .A(alu__abc_40887_new_n419_), .B(alu__abc_40887_new_n424_), .Y(alu__abc_40887_new_n425_));
OR2X2 OR2X2_2682 ( .A(alu__abc_40887_new_n425_), .B(alu__abc_40887_new_n418_), .Y(alu__abc_40887_new_n426_));
OR2X2 OR2X2_2683 ( .A(alu__abc_40887_new_n417_), .B(alu__abc_40887_new_n426_), .Y(alu__abc_40887_new_n427_));
OR2X2 OR2X2_2684 ( .A(alu__abc_40887_new_n222_), .B(alu__abc_40887_new_n200_), .Y(alu__abc_40887_new_n432_));
OR2X2 OR2X2_2685 ( .A(alu__abc_40887_new_n433_), .B(alu__abc_40887_new_n279_), .Y(alu__abc_40887_new_n434_));
OR2X2 OR2X2_2686 ( .A(alu__abc_40887_new_n437_), .B(alu__abc_40887_new_n408_), .Y(alu__abc_40887_new_n438_));
OR2X2 OR2X2_2687 ( .A(alu__abc_40887_new_n431_), .B(alu__abc_40887_new_n439_), .Y(alu__abc_40887_new_n440_));
OR2X2 OR2X2_2688 ( .A(alu__abc_40887_new_n440_), .B(alu__abc_40887_new_n387_), .Y(alu__abc_40887_new_n441_));
OR2X2 OR2X2_2689 ( .A(alu__abc_40887_new_n382_), .B(alu__abc_40887_new_n335_), .Y(alu__abc_40887_new_n442_));
OR2X2 OR2X2_269 ( .A(regfil_1__6_), .B(regfil_5__6_), .Y(_abc_41356_new_n1449_));
OR2X2 OR2X2_2690 ( .A(alu__abc_40887_new_n385_), .B(alu__abc_40887_new_n336_), .Y(alu__abc_40887_new_n443_));
OR2X2 OR2X2_2691 ( .A(alu__abc_40887_new_n438_), .B(alu__abc_40887_new_n429_), .Y(alu__abc_40887_new_n445_));
OR2X2 OR2X2_2692 ( .A(alu__abc_40887_new_n410_), .B(alu__abc_40887_new_n430_), .Y(alu__abc_40887_new_n446_));
OR2X2 OR2X2_2693 ( .A(alu__abc_40887_new_n447_), .B(alu__abc_40887_new_n444_), .Y(alu__abc_40887_new_n448_));
OR2X2 OR2X2_2694 ( .A(alu__abc_40887_new_n452_), .B(alu__abc_40887_new_n451_), .Y(alu__abc_40887_new_n453_));
OR2X2 OR2X2_2695 ( .A(alu__abc_40887_new_n454_), .B(alu__abc_40887_new_n455_), .Y(alu__abc_40887_new_n456_));
OR2X2 OR2X2_2696 ( .A(alu__abc_40887_new_n457_), .B(alu__abc_40887_new_n450_), .Y(alu_parity));
OR2X2 OR2X2_2697 ( .A(alu__abc_40887_new_n463_), .B(alu__abc_40887_new_n464_), .Y(alu_res_0_));
OR2X2 OR2X2_2698 ( .A(alu__abc_40887_new_n466_), .B(alu__abc_40887_new_n467_), .Y(alu_res_1_));
OR2X2 OR2X2_2699 ( .A(alu__abc_40887_new_n470_), .B(alu__abc_40887_new_n469_), .Y(alu_res_2_));
OR2X2 OR2X2_27 ( .A(_abc_41356_new_n662_), .B(_abc_41356_new_n641_), .Y(_abc_41356_new_n663_));
OR2X2 OR2X2_270 ( .A(regfil_1__4_), .B(regfil_5__4_), .Y(_abc_41356_new_n1454_));
OR2X2 OR2X2_2700 ( .A(alu__abc_40887_new_n473_), .B(alu__abc_40887_new_n472_), .Y(alu_res_3_));
OR2X2 OR2X2_2701 ( .A(alu__abc_40887_new_n476_), .B(alu__abc_40887_new_n475_), .Y(alu_res_4_));
OR2X2 OR2X2_2702 ( .A(alu__abc_40887_new_n479_), .B(alu__abc_40887_new_n478_), .Y(alu_res_5_));
OR2X2 OR2X2_2703 ( .A(alu__abc_40887_new_n482_), .B(alu__abc_40887_new_n481_), .Y(alu_res_6_));
OR2X2 OR2X2_2704 ( .A(alu__abc_40887_new_n485_), .B(alu__abc_40887_new_n484_), .Y(alu_res_7_));
OR2X2 OR2X2_2705 ( .A(alu__abc_40887_new_n487_), .B(alu_oprb_7_), .Y(alu__abc_40887_new_n488_));
OR2X2 OR2X2_2706 ( .A(alu__abc_40887_new_n490_), .B(alu__abc_40887_new_n489_), .Y(alu__abc_40887_new_n491_));
OR2X2 OR2X2_2707 ( .A(alu__abc_40887_new_n237_), .B(alu__abc_40887_new_n145_), .Y(alu__abc_40887_new_n492_));
OR2X2 OR2X2_2708 ( .A(alu__abc_40887_new_n495_), .B(alu__abc_40887_new_n34_), .Y(alu__abc_40887_new_n496_));
OR2X2 OR2X2_2709 ( .A(alu__abc_40887_new_n494_), .B(alu__abc_40887_new_n498_), .Y(alu__abc_40887_new_n499_));
OR2X2 OR2X2_271 ( .A(regfil_1__5_), .B(regfil_5__5_), .Y(_abc_41356_new_n1458_));
OR2X2 OR2X2_2710 ( .A(alu__abc_40887_new_n493_), .B(alu__abc_40887_new_n499_), .Y(alu_cout));
OR2X2 OR2X2_272 ( .A(_abc_41356_new_n1442_), .B(_abc_41356_new_n1462_), .Y(_abc_41356_new_n1463_));
OR2X2 OR2X2_273 ( .A(_abc_41356_new_n1452_), .B(_abc_41356_new_n1456_), .Y(_abc_41356_new_n1464_));
OR2X2 OR2X2_274 ( .A(_abc_41356_new_n1467_), .B(_abc_41356_new_n1443_), .Y(_abc_41356_new_n1468_));
OR2X2 OR2X2_275 ( .A(_abc_41356_new_n1466_), .B(_abc_41356_new_n1468_), .Y(_abc_41356_new_n1469_));
OR2X2 OR2X2_276 ( .A(_abc_41356_new_n1473_), .B(_abc_41356_new_n1474_), .Y(_abc_41356_new_n1475_));
OR2X2 OR2X2_277 ( .A(_abc_41356_new_n1472_), .B(_abc_41356_new_n1476_), .Y(_abc_41356_new_n1479_));
OR2X2 OR2X2_278 ( .A(_abc_41356_new_n1483_), .B(_abc_41356_new_n1418_), .Y(_abc_41356_new_n1484_));
OR2X2 OR2X2_279 ( .A(_abc_41356_new_n1484_), .B(_abc_41356_new_n1416_), .Y(_abc_41356_new_n1485_));
OR2X2 OR2X2_28 ( .A(_abc_41356_new_n614_), .B(regd_2_), .Y(_abc_41356_new_n664_));
OR2X2 OR2X2_280 ( .A(_abc_41356_new_n1488_), .B(_abc_41356_new_n1354_), .Y(_abc_41356_new_n1489_));
OR2X2 OR2X2_281 ( .A(_abc_41356_new_n1489_), .B(_abc_41356_new_n1285_), .Y(_abc_41356_new_n1490_));
OR2X2 OR2X2_282 ( .A(_abc_41356_new_n1492_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n1493_));
OR2X2 OR2X2_283 ( .A(_abc_41356_new_n1494_), .B(_abc_41356_new_n1247_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_0_));
OR2X2 OR2X2_284 ( .A(_abc_41356_new_n771_), .B(_abc_41356_new_n1213_), .Y(_abc_41356_new_n1496_));
OR2X2 OR2X2_285 ( .A(_abc_41356_new_n1212_), .B(regfil_4__1_), .Y(_abc_41356_new_n1497_));
OR2X2 OR2X2_286 ( .A(_abc_41356_new_n1499_), .B(_abc_41356_new_n1500_), .Y(_abc_41356_new_n1501_));
OR2X2 OR2X2_287 ( .A(_abc_41356_new_n1236_), .B(regfil_2__1_), .Y(_abc_41356_new_n1502_));
OR2X2 OR2X2_288 ( .A(_abc_41356_new_n1506_), .B(_abc_41356_new_n1505_), .Y(_abc_41356_new_n1507_));
OR2X2 OR2X2_289 ( .A(_abc_41356_new_n1508_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n1509_));
OR2X2 OR2X2_29 ( .A(_abc_41356_new_n614_), .B(regd_1_), .Y(_abc_41356_new_n669_));
OR2X2 OR2X2_290 ( .A(_abc_41356_new_n1281_), .B(regfil_4__1_), .Y(_abc_41356_new_n1510_));
OR2X2 OR2X2_291 ( .A(_abc_41356_new_n1513_), .B(_abc_41356_new_n1220_), .Y(_abc_41356_new_n1514_));
OR2X2 OR2X2_292 ( .A(_abc_41356_new_n1516_), .B(_abc_41356_new_n1517_), .Y(_abc_41356_new_n1518_));
OR2X2 OR2X2_293 ( .A(_abc_41356_new_n1519_), .B(_abc_41356_new_n1347_), .Y(_abc_41356_new_n1523_));
OR2X2 OR2X2_294 ( .A(_abc_41356_new_n1350_), .B(_abc_41356_new_n1523_), .Y(_abc_41356_new_n1524_));
OR2X2 OR2X2_295 ( .A(_abc_41356_new_n1533_), .B(_abc_41356_new_n1531_), .Y(_abc_41356_new_n1534_));
OR2X2 OR2X2_296 ( .A(_abc_41356_new_n1535_), .B(_abc_41356_new_n1407_), .Y(_abc_41356_new_n1536_));
OR2X2 OR2X2_297 ( .A(_abc_41356_new_n1530_), .B(_abc_41356_new_n1536_), .Y(_abc_41356_new_n1537_));
OR2X2 OR2X2_298 ( .A(_abc_41356_new_n1547_), .B(_abc_41356_new_n1548_), .Y(_abc_41356_new_n1549_));
OR2X2 OR2X2_299 ( .A(_abc_41356_new_n1471_), .B(_abc_41356_new_n1552_), .Y(_abc_41356_new_n1553_));
OR2X2 OR2X2_3 ( .A(_abc_41356_new_n552_), .B(_abc_41356_new_n538_), .Y(_abc_41356_new_n553_));
OR2X2 OR2X2_30 ( .A(_abc_41356_new_n675_), .B(_abc_41356_new_n686_), .Y(_abc_41356_new_n687_));
OR2X2 OR2X2_300 ( .A(_abc_41356_new_n1550_), .B(_abc_41356_new_n1474_), .Y(_abc_41356_new_n1554_));
OR2X2 OR2X2_301 ( .A(_abc_41356_new_n1477_), .B(_abc_41356_new_n1554_), .Y(_abc_41356_new_n1555_));
OR2X2 OR2X2_302 ( .A(_abc_41356_new_n1560_), .B(_abc_41356_new_n1418_), .Y(_abc_41356_new_n1561_));
OR2X2 OR2X2_303 ( .A(_abc_41356_new_n1561_), .B(_abc_41356_new_n1545_), .Y(_abc_41356_new_n1562_));
OR2X2 OR2X2_304 ( .A(_abc_41356_new_n1565_), .B(_abc_41356_new_n1529_), .Y(_abc_41356_new_n1566_));
OR2X2 OR2X2_305 ( .A(_abc_41356_new_n1566_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n1567_));
OR2X2 OR2X2_306 ( .A(_abc_41356_new_n1568_), .B(_abc_41356_new_n1509_), .Y(_abc_41356_new_n1569_));
OR2X2 OR2X2_307 ( .A(_abc_41356_new_n1570_), .B(_abc_41356_new_n1501_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_1_));
OR2X2 OR2X2_308 ( .A(_abc_41356_new_n824_), .B(_abc_41356_new_n1213_), .Y(_abc_41356_new_n1572_));
OR2X2 OR2X2_309 ( .A(_abc_41356_new_n1212_), .B(regfil_4__2_), .Y(_abc_41356_new_n1573_));
OR2X2 OR2X2_31 ( .A(_abc_41356_new_n674_), .B(_abc_41356_new_n687_), .Y(_abc_41356_new_n688_));
OR2X2 OR2X2_310 ( .A(_abc_41356_new_n1575_), .B(_abc_41356_new_n1576_), .Y(_abc_41356_new_n1577_));
OR2X2 OR2X2_311 ( .A(_abc_41356_new_n1236_), .B(regfil_2__2_), .Y(_abc_41356_new_n1578_));
OR2X2 OR2X2_312 ( .A(_abc_41356_new_n1505_), .B(_abc_41356_new_n1580_), .Y(_abc_41356_new_n1583_));
OR2X2 OR2X2_313 ( .A(_abc_41356_new_n1511_), .B(regfil_4__2_), .Y(_abc_41356_new_n1587_));
OR2X2 OR2X2_314 ( .A(_abc_41356_new_n1590_), .B(_abc_41356_new_n1220_), .Y(_abc_41356_new_n1591_));
OR2X2 OR2X2_315 ( .A(_abc_41356_new_n1597_), .B(_abc_41356_new_n1598_), .Y(_abc_41356_new_n1599_));
OR2X2 OR2X2_316 ( .A(_abc_41356_new_n1595_), .B(_abc_41356_new_n1600_), .Y(_abc_41356_new_n1603_));
OR2X2 OR2X2_317 ( .A(_abc_41356_new_n1541_), .B(_abc_41356_new_n1531_), .Y(_abc_41356_new_n1606_));
OR2X2 OR2X2_318 ( .A(_abc_41356_new_n1539_), .B(_abc_41356_new_n1606_), .Y(_abc_41356_new_n1607_));
OR2X2 OR2X2_319 ( .A(_abc_41356_new_n1609_), .B(_abc_41356_new_n1610_), .Y(_abc_41356_new_n1611_));
OR2X2 OR2X2_32 ( .A(_abc_41356_new_n614_), .B(regd_0_), .Y(_abc_41356_new_n691_));
OR2X2 OR2X2_320 ( .A(_abc_41356_new_n1607_), .B(_abc_41356_new_n1612_), .Y(_abc_41356_new_n1615_));
OR2X2 OR2X2_321 ( .A(_abc_41356_new_n1556_), .B(_abc_41356_new_n1548_), .Y(_abc_41356_new_n1618_));
OR2X2 OR2X2_322 ( .A(_abc_41356_new_n1622_), .B(_abc_41356_new_n1623_), .Y(_abc_41356_new_n1624_));
OR2X2 OR2X2_323 ( .A(_abc_41356_new_n1620_), .B(_abc_41356_new_n1624_), .Y(_abc_41356_new_n1625_));
OR2X2 OR2X2_324 ( .A(_abc_41356_new_n1626_), .B(_abc_41356_new_n1627_), .Y(_abc_41356_new_n1628_));
OR2X2 OR2X2_325 ( .A(_abc_41356_new_n1630_), .B(_abc_41356_new_n1418_), .Y(_abc_41356_new_n1631_));
OR2X2 OR2X2_326 ( .A(_abc_41356_new_n1631_), .B(_abc_41356_new_n1617_), .Y(_abc_41356_new_n1632_));
OR2X2 OR2X2_327 ( .A(_abc_41356_new_n1635_), .B(_abc_41356_new_n1605_), .Y(_abc_41356_new_n1636_));
OR2X2 OR2X2_328 ( .A(_abc_41356_new_n1636_), .B(_abc_41356_new_n1285_), .Y(_abc_41356_new_n1637_));
OR2X2 OR2X2_329 ( .A(_abc_41356_new_n1639_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n1640_));
OR2X2 OR2X2_33 ( .A(_abc_41356_new_n663_), .B(_abc_41356_new_n696_), .Y(_abc_41356_new_n697_));
OR2X2 OR2X2_330 ( .A(_abc_41356_new_n1641_), .B(_abc_41356_new_n1577_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_2_));
OR2X2 OR2X2_331 ( .A(_abc_41356_new_n885_), .B(_abc_41356_new_n1213_), .Y(_abc_41356_new_n1643_));
OR2X2 OR2X2_332 ( .A(_abc_41356_new_n1212_), .B(regfil_4__3_), .Y(_abc_41356_new_n1644_));
OR2X2 OR2X2_333 ( .A(_abc_41356_new_n1646_), .B(_abc_41356_new_n1647_), .Y(_abc_41356_new_n1648_));
OR2X2 OR2X2_334 ( .A(_abc_41356_new_n1236_), .B(regfil_2__3_), .Y(_abc_41356_new_n1649_));
OR2X2 OR2X2_335 ( .A(_abc_41356_new_n1601_), .B(_abc_41356_new_n1598_), .Y(_abc_41356_new_n1651_));
OR2X2 OR2X2_336 ( .A(_abc_41356_new_n1662_), .B(_abc_41356_new_n1660_), .Y(_abc_41356_new_n1663_));
OR2X2 OR2X2_337 ( .A(_abc_41356_new_n1613_), .B(_abc_41356_new_n1610_), .Y(_abc_41356_new_n1666_));
OR2X2 OR2X2_338 ( .A(_abc_41356_new_n1666_), .B(_abc_41356_new_n1672_), .Y(_abc_41356_new_n1673_));
OR2X2 OR2X2_339 ( .A(_abc_41356_new_n1674_), .B(_abc_41356_new_n1675_), .Y(_abc_41356_new_n1676_));
OR2X2 OR2X2_34 ( .A(_abc_41356_new_n551_), .B(_abc_41356_new_n537_), .Y(_abc_41356_new_n698_));
OR2X2 OR2X2_340 ( .A(_abc_41356_new_n1677_), .B(_abc_41356_new_n1665_), .Y(_abc_41356_new_n1678_));
OR2X2 OR2X2_341 ( .A(_abc_41356_new_n1681_), .B(_abc_41356_new_n1687_), .Y(_abc_41356_new_n1688_));
OR2X2 OR2X2_342 ( .A(_abc_41356_new_n1680_), .B(_abc_41356_new_n1689_), .Y(_abc_41356_new_n1690_));
OR2X2 OR2X2_343 ( .A(_abc_41356_new_n1692_), .B(_abc_41356_new_n1415_), .Y(_abc_41356_new_n1693_));
OR2X2 OR2X2_344 ( .A(_abc_41356_new_n1694_), .B(_abc_41356_new_n1695_), .Y(_abc_41356_new_n1696_));
OR2X2 OR2X2_345 ( .A(_abc_41356_new_n1696_), .B(_abc_41356_new_n1664_), .Y(_abc_41356_new_n1697_));
OR2X2 OR2X2_346 ( .A(_abc_41356_new_n1588_), .B(regfil_4__3_), .Y(_abc_41356_new_n1698_));
OR2X2 OR2X2_347 ( .A(_abc_41356_new_n1702_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n1703_));
OR2X2 OR2X2_348 ( .A(_abc_41356_new_n1697_), .B(_abc_41356_new_n1703_), .Y(_abc_41356_new_n1704_));
OR2X2 OR2X2_349 ( .A(_abc_41356_new_n1709_), .B(_abc_41356_new_n1705_), .Y(_abc_41356_new_n1710_));
OR2X2 OR2X2_35 ( .A(_abc_41356_new_n530_), .B(_abc_41356_new_n555_), .Y(_abc_41356_new_n699_));
OR2X2 OR2X2_350 ( .A(_abc_41356_new_n1711_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n1712_));
OR2X2 OR2X2_351 ( .A(_abc_41356_new_n1713_), .B(_abc_41356_new_n1648_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_3_));
OR2X2 OR2X2_352 ( .A(_abc_41356_new_n952_), .B(_abc_41356_new_n1213_), .Y(_abc_41356_new_n1715_));
OR2X2 OR2X2_353 ( .A(_abc_41356_new_n1212_), .B(regfil_4__4_), .Y(_abc_41356_new_n1716_));
OR2X2 OR2X2_354 ( .A(_abc_41356_new_n1718_), .B(_abc_41356_new_n1719_), .Y(_abc_41356_new_n1720_));
OR2X2 OR2X2_355 ( .A(_abc_41356_new_n1236_), .B(regfil_2__4_), .Y(_abc_41356_new_n1721_));
OR2X2 OR2X2_356 ( .A(_abc_41356_new_n1725_), .B(_abc_41356_new_n1724_), .Y(_abc_41356_new_n1726_));
OR2X2 OR2X2_357 ( .A(_abc_41356_new_n1727_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n1728_));
OR2X2 OR2X2_358 ( .A(_abc_41356_new_n1734_), .B(_abc_41356_new_n1656_), .Y(_abc_41356_new_n1735_));
OR2X2 OR2X2_359 ( .A(_abc_41356_new_n1733_), .B(_abc_41356_new_n1735_), .Y(_abc_41356_new_n1736_));
OR2X2 OR2X2_36 ( .A(_abc_41356_new_n704_), .B(carry), .Y(_abc_41356_new_n705_));
OR2X2 OR2X2_360 ( .A(_abc_41356_new_n1731_), .B(_abc_41356_new_n1736_), .Y(_abc_41356_new_n1737_));
OR2X2 OR2X2_361 ( .A(_abc_41356_new_n1739_), .B(_abc_41356_new_n1740_), .Y(_abc_41356_new_n1741_));
OR2X2 OR2X2_362 ( .A(_abc_41356_new_n1737_), .B(_abc_41356_new_n1742_), .Y(_abc_41356_new_n1745_));
OR2X2 OR2X2_363 ( .A(_abc_41356_new_n1749_), .B(_abc_41356_new_n1750_), .Y(_abc_41356_new_n1751_));
OR2X2 OR2X2_364 ( .A(_abc_41356_new_n1753_), .B(_abc_41356_new_n1682_), .Y(_abc_41356_new_n1754_));
OR2X2 OR2X2_365 ( .A(_abc_41356_new_n1756_), .B(_abc_41356_new_n1754_), .Y(_abc_41356_new_n1757_));
OR2X2 OR2X2_366 ( .A(_abc_41356_new_n1471_), .B(_abc_41356_new_n1760_), .Y(_abc_41356_new_n1761_));
OR2X2 OR2X2_367 ( .A(_abc_41356_new_n1763_), .B(_abc_41356_new_n1752_), .Y(_abc_41356_new_n1766_));
OR2X2 OR2X2_368 ( .A(_abc_41356_new_n1773_), .B(_abc_41356_new_n1667_), .Y(_abc_41356_new_n1774_));
OR2X2 OR2X2_369 ( .A(_abc_41356_new_n1772_), .B(_abc_41356_new_n1774_), .Y(_abc_41356_new_n1775_));
OR2X2 OR2X2_37 ( .A(_abc_41356_new_n718_), .B(_abc_41356_new_n714_), .Y(_abc_41356_new_n719_));
OR2X2 OR2X2_370 ( .A(_abc_41356_new_n1771_), .B(_abc_41356_new_n1775_), .Y(_abc_41356_new_n1776_));
OR2X2 OR2X2_371 ( .A(_abc_41356_new_n1778_), .B(_abc_41356_new_n1779_), .Y(_abc_41356_new_n1780_));
OR2X2 OR2X2_372 ( .A(_abc_41356_new_n1776_), .B(_abc_41356_new_n1781_), .Y(_abc_41356_new_n1784_));
OR2X2 OR2X2_373 ( .A(_abc_41356_new_n1786_), .B(_abc_41356_new_n1418_), .Y(_abc_41356_new_n1787_));
OR2X2 OR2X2_374 ( .A(_abc_41356_new_n1787_), .B(_abc_41356_new_n1768_), .Y(_abc_41356_new_n1788_));
OR2X2 OR2X2_375 ( .A(_abc_41356_new_n1791_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n1792_));
OR2X2 OR2X2_376 ( .A(_abc_41356_new_n1792_), .B(_abc_41356_new_n1747_), .Y(_abc_41356_new_n1793_));
OR2X2 OR2X2_377 ( .A(_abc_41356_new_n1699_), .B(regfil_4__4_), .Y(_abc_41356_new_n1794_));
OR2X2 OR2X2_378 ( .A(_abc_41356_new_n1805_), .B(_abc_41356_new_n1220_), .Y(_abc_41356_new_n1806_));
OR2X2 OR2X2_379 ( .A(_abc_41356_new_n1807_), .B(_abc_41356_new_n1728_), .Y(_abc_41356_new_n1808_));
OR2X2 OR2X2_38 ( .A(_abc_41356_new_n719_), .B(_abc_41356_new_n512_), .Y(_abc_41356_new_n720_));
OR2X2 OR2X2_380 ( .A(_abc_41356_new_n1809_), .B(_abc_41356_new_n1720_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_4_));
OR2X2 OR2X2_381 ( .A(_abc_41356_new_n1019_), .B(_abc_41356_new_n1213_), .Y(_abc_41356_new_n1811_));
OR2X2 OR2X2_382 ( .A(_abc_41356_new_n1212_), .B(regfil_4__5_), .Y(_abc_41356_new_n1812_));
OR2X2 OR2X2_383 ( .A(_abc_41356_new_n1814_), .B(_abc_41356_new_n1815_), .Y(_abc_41356_new_n1816_));
OR2X2 OR2X2_384 ( .A(_abc_41356_new_n1236_), .B(regfil_2__5_), .Y(_abc_41356_new_n1817_));
OR2X2 OR2X2_385 ( .A(_abc_41356_new_n1822_), .B(_abc_41356_new_n1820_), .Y(_abc_41356_new_n1823_));
OR2X2 OR2X2_386 ( .A(_abc_41356_new_n1824_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n1825_));
OR2X2 OR2X2_387 ( .A(_abc_41356_new_n1827_), .B(_abc_41356_new_n1828_), .Y(_abc_41356_new_n1829_));
OR2X2 OR2X2_388 ( .A(_abc_41356_new_n1830_), .B(_abc_41356_new_n1740_), .Y(_abc_41356_new_n1833_));
OR2X2 OR2X2_389 ( .A(_abc_41356_new_n1743_), .B(_abc_41356_new_n1833_), .Y(_abc_41356_new_n1834_));
OR2X2 OR2X2_39 ( .A(_abc_41356_new_n720_), .B(_abc_41356_new_n712_), .Y(_abc_41356_new_n721_));
OR2X2 OR2X2_390 ( .A(_abc_41356_new_n1843_), .B(_abc_41356_new_n1844_), .Y(_abc_41356_new_n1845_));
OR2X2 OR2X2_391 ( .A(_abc_41356_new_n1846_), .B(_abc_41356_new_n1779_), .Y(_abc_41356_new_n1847_));
OR2X2 OR2X2_392 ( .A(_abc_41356_new_n1782_), .B(_abc_41356_new_n1847_), .Y(_abc_41356_new_n1848_));
OR2X2 OR2X2_393 ( .A(_abc_41356_new_n1858_), .B(_abc_41356_new_n1859_), .Y(_abc_41356_new_n1860_));
OR2X2 OR2X2_394 ( .A(_abc_41356_new_n1762_), .B(_abc_41356_new_n1863_), .Y(_abc_41356_new_n1864_));
OR2X2 OR2X2_395 ( .A(_abc_41356_new_n1861_), .B(_abc_41356_new_n1750_), .Y(_abc_41356_new_n1865_));
OR2X2 OR2X2_396 ( .A(_abc_41356_new_n1764_), .B(_abc_41356_new_n1865_), .Y(_abc_41356_new_n1866_));
OR2X2 OR2X2_397 ( .A(_abc_41356_new_n1871_), .B(_abc_41356_new_n1856_), .Y(_abc_41356_new_n1872_));
OR2X2 OR2X2_398 ( .A(_abc_41356_new_n1872_), .B(_abc_41356_new_n1841_), .Y(_abc_41356_new_n1873_));
OR2X2 OR2X2_399 ( .A(_abc_41356_new_n1873_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n1874_));
OR2X2 OR2X2_4 ( .A(_abc_41356_new_n557_), .B(_abc_41356_new_n556_), .Y(_abc_41356_new_n558_));
OR2X2 OR2X2_40 ( .A(_abc_41356_new_n721_), .B(_abc_41356_new_n699_), .Y(_abc_41356_new_n722_));
OR2X2 OR2X2_400 ( .A(_abc_41356_new_n1874_), .B(_abc_41356_new_n1840_), .Y(_abc_41356_new_n1875_));
OR2X2 OR2X2_401 ( .A(_abc_41356_new_n1803_), .B(regfil_4__5_), .Y(_abc_41356_new_n1876_));
OR2X2 OR2X2_402 ( .A(_abc_41356_new_n1879_), .B(_abc_41356_new_n1220_), .Y(_abc_41356_new_n1880_));
OR2X2 OR2X2_403 ( .A(_abc_41356_new_n1881_), .B(_abc_41356_new_n1825_), .Y(_abc_41356_new_n1882_));
OR2X2 OR2X2_404 ( .A(_abc_41356_new_n1883_), .B(_abc_41356_new_n1816_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_5_));
OR2X2 OR2X2_405 ( .A(_abc_41356_new_n1091_), .B(_abc_41356_new_n1213_), .Y(_abc_41356_new_n1885_));
OR2X2 OR2X2_406 ( .A(_abc_41356_new_n1212_), .B(regfil_4__6_), .Y(_abc_41356_new_n1886_));
OR2X2 OR2X2_407 ( .A(_abc_41356_new_n1888_), .B(_abc_41356_new_n1889_), .Y(_abc_41356_new_n1890_));
OR2X2 OR2X2_408 ( .A(_abc_41356_new_n1236_), .B(regfil_2__6_), .Y(_abc_41356_new_n1891_));
OR2X2 OR2X2_409 ( .A(_abc_41356_new_n1896_), .B(_abc_41356_new_n1894_), .Y(_abc_41356_new_n1897_));
OR2X2 OR2X2_41 ( .A(_abc_41356_new_n722_), .B(_abc_41356_new_n698_), .Y(_abc_41356_new_n723_));
OR2X2 OR2X2_410 ( .A(_abc_41356_new_n1898_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n1899_));
OR2X2 OR2X2_411 ( .A(_abc_41356_new_n1831_), .B(_abc_41356_new_n1828_), .Y(_abc_41356_new_n1900_));
OR2X2 OR2X2_412 ( .A(_abc_41356_new_n1836_), .B(_abc_41356_new_n1900_), .Y(_abc_41356_new_n1901_));
OR2X2 OR2X2_413 ( .A(_abc_41356_new_n1903_), .B(_abc_41356_new_n1904_), .Y(_abc_41356_new_n1905_));
OR2X2 OR2X2_414 ( .A(_abc_41356_new_n1901_), .B(_abc_41356_new_n1906_), .Y(_abc_41356_new_n1907_));
OR2X2 OR2X2_415 ( .A(_abc_41356_new_n1867_), .B(_abc_41356_new_n1859_), .Y(_abc_41356_new_n1912_));
OR2X2 OR2X2_416 ( .A(_abc_41356_new_n1916_), .B(_abc_41356_new_n1917_), .Y(_abc_41356_new_n1918_));
OR2X2 OR2X2_417 ( .A(_abc_41356_new_n1915_), .B(_abc_41356_new_n1919_), .Y(_abc_41356_new_n1920_));
OR2X2 OR2X2_418 ( .A(_abc_41356_new_n1914_), .B(_abc_41356_new_n1918_), .Y(_abc_41356_new_n1921_));
OR2X2 OR2X2_419 ( .A(_abc_41356_new_n1853_), .B(_abc_41356_new_n1844_), .Y(_abc_41356_new_n1924_));
OR2X2 OR2X2_42 ( .A(_abc_41356_new_n695_), .B(regfil_7__0_), .Y(_abc_41356_new_n725_));
OR2X2 OR2X2_420 ( .A(_abc_41356_new_n1850_), .B(_abc_41356_new_n1924_), .Y(_abc_41356_new_n1925_));
OR2X2 OR2X2_421 ( .A(_abc_41356_new_n1927_), .B(_abc_41356_new_n1928_), .Y(_abc_41356_new_n1929_));
OR2X2 OR2X2_422 ( .A(_abc_41356_new_n1925_), .B(_abc_41356_new_n1930_), .Y(_abc_41356_new_n1933_));
OR2X2 OR2X2_423 ( .A(_abc_41356_new_n1935_), .B(_abc_41356_new_n1418_), .Y(_abc_41356_new_n1936_));
OR2X2 OR2X2_424 ( .A(_abc_41356_new_n1936_), .B(_abc_41356_new_n1923_), .Y(_abc_41356_new_n1937_));
OR2X2 OR2X2_425 ( .A(_abc_41356_new_n1940_), .B(_abc_41356_new_n1219_), .Y(_abc_41356_new_n1941_));
OR2X2 OR2X2_426 ( .A(_abc_41356_new_n1941_), .B(_abc_41356_new_n1911_), .Y(_abc_41356_new_n1942_));
OR2X2 OR2X2_427 ( .A(_abc_41356_new_n1877_), .B(regfil_4__6_), .Y(_abc_41356_new_n1943_));
OR2X2 OR2X2_428 ( .A(_abc_41356_new_n1946_), .B(_abc_41356_new_n1220_), .Y(_abc_41356_new_n1947_));
OR2X2 OR2X2_429 ( .A(_abc_41356_new_n1948_), .B(_abc_41356_new_n1899_), .Y(_abc_41356_new_n1949_));
OR2X2 OR2X2_43 ( .A(_abc_41356_new_n730_), .B(_abc_41356_new_n729_), .Y(_abc_41356_new_n731_));
OR2X2 OR2X2_430 ( .A(_abc_41356_new_n1950_), .B(_abc_41356_new_n1890_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_6_));
OR2X2 OR2X2_431 ( .A(_abc_41356_new_n1953_), .B(_abc_41356_new_n1952_), .Y(_abc_41356_new_n1954_));
OR2X2 OR2X2_432 ( .A(_abc_41356_new_n1955_), .B(_abc_41356_new_n1956_), .Y(_abc_41356_new_n1957_));
OR2X2 OR2X2_433 ( .A(_abc_41356_new_n1236_), .B(regfil_2__7_), .Y(_abc_41356_new_n1958_));
OR2X2 OR2X2_434 ( .A(_abc_41356_new_n1894_), .B(regfil_4__7_), .Y(_abc_41356_new_n1960_));
OR2X2 OR2X2_435 ( .A(_abc_41356_new_n1962_), .B(_abc_41356_new_n1961_), .Y(_abc_41356_new_n1963_));
OR2X2 OR2X2_436 ( .A(_abc_41356_new_n1964_), .B(_abc_41356_new_n1217_), .Y(_abc_41356_new_n1965_));
OR2X2 OR2X2_437 ( .A(_abc_41356_new_n1908_), .B(_abc_41356_new_n1904_), .Y(_abc_41356_new_n1966_));
OR2X2 OR2X2_438 ( .A(_abc_41356_new_n1968_), .B(_abc_41356_new_n1969_), .Y(_abc_41356_new_n1970_));
OR2X2 OR2X2_439 ( .A(_abc_41356_new_n1974_), .B(_abc_41356_new_n1971_), .Y(_abc_41356_new_n1975_));
OR2X2 OR2X2_44 ( .A(_abc_41356_new_n731_), .B(_abc_41356_new_n728_), .Y(_abc_41356_new_n732_));
OR2X2 OR2X2_440 ( .A(_abc_41356_new_n1980_), .B(_abc_41356_new_n1981_), .Y(_abc_41356_new_n1982_));
OR2X2 OR2X2_441 ( .A(_abc_41356_new_n1984_), .B(_abc_41356_new_n1917_), .Y(_abc_41356_new_n1985_));
OR2X2 OR2X2_442 ( .A(_abc_41356_new_n1985_), .B(_abc_41356_new_n1983_), .Y(_abc_41356_new_n1986_));
OR2X2 OR2X2_443 ( .A(_abc_41356_new_n1921_), .B(_abc_41356_new_n1982_), .Y(_abc_41356_new_n1987_));
OR2X2 OR2X2_444 ( .A(_abc_41356_new_n1982_), .B(_abc_41356_new_n1989_), .Y(_abc_41356_new_n1990_));
OR2X2 OR2X2_445 ( .A(_abc_41356_new_n1931_), .B(_abc_41356_new_n1928_), .Y(_abc_41356_new_n1994_));
OR2X2 OR2X2_446 ( .A(_abc_41356_new_n1997_), .B(_abc_41356_new_n1998_), .Y(_abc_41356_new_n1999_));
OR2X2 OR2X2_447 ( .A(_abc_41356_new_n1995_), .B(_abc_41356_new_n1999_), .Y(_abc_41356_new_n2000_));
OR2X2 OR2X2_448 ( .A(_abc_41356_new_n1994_), .B(_abc_41356_new_n2002_), .Y(_abc_41356_new_n2003_));
OR2X2 OR2X2_449 ( .A(_abc_41356_new_n2005_), .B(_abc_41356_new_n1993_), .Y(_abc_41356_new_n2006_));
OR2X2 OR2X2_45 ( .A(_abc_41356_new_n727_), .B(_abc_41356_new_n732_), .Y(_abc_41356_new_n733_));
OR2X2 OR2X2_450 ( .A(_abc_41356_new_n2006_), .B(_abc_41356_new_n1979_), .Y(_abc_41356_new_n2007_));
OR2X2 OR2X2_451 ( .A(_abc_41356_new_n2007_), .B(_abc_41356_new_n1976_), .Y(_abc_41356_new_n2008_));
OR2X2 OR2X2_452 ( .A(_abc_41356_new_n1944_), .B(regfil_4__7_), .Y(_abc_41356_new_n2011_));
OR2X2 OR2X2_453 ( .A(_abc_41356_new_n2013_), .B(_abc_41356_new_n1216_), .Y(_abc_41356_new_n2014_));
OR2X2 OR2X2_454 ( .A(_abc_41356_new_n2008_), .B(_abc_41356_new_n2014_), .Y(_abc_41356_new_n2015_));
OR2X2 OR2X2_455 ( .A(_abc_41356_new_n2016_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n2017_));
OR2X2 OR2X2_456 ( .A(_abc_41356_new_n2018_), .B(_abc_41356_new_n1957_), .Y(_abc_36060_memoryregfil_wrmux_4__4__0__y_16147_7_));
OR2X2 OR2X2_457 ( .A(_abc_41356_new_n2020_), .B(_abc_41356_new_n2023_), .Y(_abc_41356_new_n2024_));
OR2X2 OR2X2_458 ( .A(_abc_41356_new_n2028_), .B(regfil_4__0_), .Y(_abc_41356_new_n2029_));
OR2X2 OR2X2_459 ( .A(_abc_41356_new_n2027_), .B(wdatahold2_0_), .Y(_abc_41356_new_n2030_));
OR2X2 OR2X2_46 ( .A(_abc_41356_new_n733_), .B(_abc_41356_new_n567_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_0_));
OR2X2 OR2X2_460 ( .A(pc_1_), .B(pc_0_), .Y(_abc_41356_new_n2033_));
OR2X2 OR2X2_461 ( .A(_abc_41356_new_n2043_), .B(_abc_41356_new_n2040_), .Y(_abc_41356_new_n2044_));
OR2X2 OR2X2_462 ( .A(_abc_41356_new_n2049_), .B(pc_8_), .Y(_abc_41356_new_n2050_));
OR2X2 OR2X2_463 ( .A(_abc_41356_new_n2051_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n2052_));
OR2X2 OR2X2_464 ( .A(_abc_41356_new_n554_), .B(_abc_41356_new_n2057_), .Y(_abc_41356_new_n2058_));
OR2X2 OR2X2_465 ( .A(_abc_41356_new_n2058_), .B(_abc_41356_new_n2055_), .Y(_abc_41356_new_n2059_));
OR2X2 OR2X2_466 ( .A(_abc_41356_new_n2059_), .B(_abc_41356_new_n536_), .Y(_abc_41356_new_n2060_));
OR2X2 OR2X2_467 ( .A(_abc_41356_new_n2075_), .B(_abc_41356_new_n2076_), .Y(_abc_41356_new_n2077_));
OR2X2 OR2X2_468 ( .A(_abc_41356_new_n2082_), .B(_abc_41356_new_n2081_), .Y(_abc_41356_new_n2083_));
OR2X2 OR2X2_469 ( .A(_abc_41356_new_n2085_), .B(_abc_41356_new_n2084_), .Y(_abc_41356_new_n2086_));
OR2X2 OR2X2_47 ( .A(regfil_0__0_), .B(regfil_0__1_), .Y(_abc_41356_new_n735_));
OR2X2 OR2X2_470 ( .A(_abc_41356_new_n2083_), .B(_abc_41356_new_n2087_), .Y(_abc_41356_new_n2088_));
OR2X2 OR2X2_471 ( .A(_abc_41356_new_n2089_), .B(_abc_41356_new_n2090_), .Y(_abc_41356_new_n2091_));
OR2X2 OR2X2_472 ( .A(_abc_41356_new_n2091_), .B(_abc_41356_new_n2080_), .Y(_abc_41356_new_n2092_));
OR2X2 OR2X2_473 ( .A(_abc_41356_new_n2079_), .B(_abc_41356_new_n2092_), .Y(_abc_41356_new_n2093_));
OR2X2 OR2X2_474 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n2093_), .Y(_abc_41356_new_n2094_));
OR2X2 OR2X2_475 ( .A(_abc_41356_new_n2094_), .B(_abc_41356_new_n2053_), .Y(_abc_41356_new_n2095_));
OR2X2 OR2X2_476 ( .A(_abc_41356_new_n2096_), .B(wdatahold2_0_), .Y(_abc_41356_new_n2097_));
OR2X2 OR2X2_477 ( .A(_abc_41356_new_n2099_), .B(_abc_41356_new_n2032_), .Y(_abc_41356_new_n2100_));
OR2X2 OR2X2_478 ( .A(_abc_41356_new_n2101_), .B(_abc_41356_new_n2025_), .Y(_0wdatahold2_7_0__0_));
OR2X2 OR2X2_479 ( .A(_abc_41356_new_n2028_), .B(regfil_4__1_), .Y(_abc_41356_new_n2104_));
OR2X2 OR2X2_48 ( .A(_abc_41356_new_n656_), .B(_abc_41356_new_n735_), .Y(_abc_41356_new_n736_));
OR2X2 OR2X2_480 ( .A(_abc_41356_new_n2027_), .B(wdatahold2_1_), .Y(_abc_41356_new_n2105_));
OR2X2 OR2X2_481 ( .A(_abc_41356_new_n2040_), .B(pc_9_), .Y(_abc_41356_new_n2110_));
OR2X2 OR2X2_482 ( .A(_abc_41356_new_n2049_), .B(pc_9_), .Y(_abc_41356_new_n2112_));
OR2X2 OR2X2_483 ( .A(_abc_41356_new_n2113_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n2114_));
OR2X2 OR2X2_484 ( .A(_abc_41356_new_n2076_), .B(pc_9_), .Y(_abc_41356_new_n2116_));
OR2X2 OR2X2_485 ( .A(_abc_41356_new_n579_), .B(_abc_41356_new_n2065_), .Y(_abc_41356_new_n2121_));
OR2X2 OR2X2_486 ( .A(_abc_41356_new_n2126_), .B(_abc_41356_new_n2125_), .Y(_abc_41356_new_n2127_));
OR2X2 OR2X2_487 ( .A(_abc_41356_new_n2128_), .B(_abc_41356_new_n2124_), .Y(_abc_41356_new_n2129_));
OR2X2 OR2X2_488 ( .A(_abc_41356_new_n2130_), .B(_abc_41356_new_n2131_), .Y(_abc_41356_new_n2132_));
OR2X2 OR2X2_489 ( .A(_abc_41356_new_n2132_), .B(_abc_41356_new_n2123_), .Y(_abc_41356_new_n2133_));
OR2X2 OR2X2_49 ( .A(_abc_41356_new_n739_), .B(_abc_41356_new_n737_), .Y(_abc_41356_new_n740_));
OR2X2 OR2X2_490 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n2133_), .Y(_abc_41356_new_n2134_));
OR2X2 OR2X2_491 ( .A(_abc_41356_new_n2134_), .B(_abc_41356_new_n2120_), .Y(_abc_41356_new_n2135_));
OR2X2 OR2X2_492 ( .A(_abc_41356_new_n2135_), .B(_abc_41356_new_n2115_), .Y(_abc_41356_new_n2136_));
OR2X2 OR2X2_493 ( .A(_abc_41356_new_n2096_), .B(wdatahold2_1_), .Y(_abc_41356_new_n2137_));
OR2X2 OR2X2_494 ( .A(_abc_41356_new_n2139_), .B(_abc_41356_new_n2107_), .Y(_abc_41356_new_n2140_));
OR2X2 OR2X2_495 ( .A(_abc_41356_new_n2141_), .B(_abc_41356_new_n2103_), .Y(_0wdatahold2_7_0__1_));
OR2X2 OR2X2_496 ( .A(_abc_41356_new_n2027_), .B(wdatahold2_2_), .Y(_abc_41356_new_n2144_));
OR2X2 OR2X2_497 ( .A(_abc_41356_new_n2028_), .B(regfil_4__2_), .Y(_abc_41356_new_n2145_));
OR2X2 OR2X2_498 ( .A(_abc_41356_new_n2150_), .B(_abc_41356_new_n2148_), .Y(_abc_41356_new_n2151_));
OR2X2 OR2X2_499 ( .A(_abc_41356_new_n2049_), .B(pc_10_), .Y(_abc_41356_new_n2153_));
OR2X2 OR2X2_5 ( .A(_abc_41356_new_n559_), .B(_abc_41356_new_n530_), .Y(_abc_41356_new_n560_));
OR2X2 OR2X2_50 ( .A(_abc_41356_new_n582_), .B(regfil_0__1_), .Y(_abc_41356_new_n742_));
OR2X2 OR2X2_500 ( .A(_abc_41356_new_n2154_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n2155_));
OR2X2 OR2X2_501 ( .A(_abc_41356_new_n2157_), .B(_abc_41356_new_n2158_), .Y(_abc_41356_new_n2159_));
OR2X2 OR2X2_502 ( .A(_abc_41356_new_n2164_), .B(_abc_41356_new_n2163_), .Y(_abc_41356_new_n2165_));
OR2X2 OR2X2_503 ( .A(_abc_41356_new_n2166_), .B(_abc_41356_new_n2162_), .Y(_abc_41356_new_n2167_));
OR2X2 OR2X2_504 ( .A(_abc_41356_new_n2169_), .B(_abc_41356_new_n2171_), .Y(_abc_41356_new_n2172_));
OR2X2 OR2X2_505 ( .A(_abc_41356_new_n2172_), .B(_abc_41356_new_n2168_), .Y(_abc_41356_new_n2173_));
OR2X2 OR2X2_506 ( .A(_abc_41356_new_n2069_), .B(_abc_41356_new_n2173_), .Y(_abc_41356_new_n2174_));
OR2X2 OR2X2_507 ( .A(_abc_41356_new_n2174_), .B(_abc_41356_new_n2161_), .Y(_abc_41356_new_n2175_));
OR2X2 OR2X2_508 ( .A(_abc_41356_new_n2175_), .B(_abc_41356_new_n2156_), .Y(_abc_41356_new_n2176_));
OR2X2 OR2X2_509 ( .A(_abc_41356_new_n2096_), .B(wdatahold2_2_), .Y(_abc_41356_new_n2177_));
OR2X2 OR2X2_51 ( .A(_abc_41356_new_n748_), .B(_abc_41356_new_n749_), .Y(_abc_41356_new_n750_));
OR2X2 OR2X2_510 ( .A(_abc_41356_new_n2179_), .B(_abc_41356_new_n2147_), .Y(_abc_41356_new_n2180_));
OR2X2 OR2X2_511 ( .A(_abc_41356_new_n2181_), .B(_abc_41356_new_n2143_), .Y(_0wdatahold2_7_0__2_));
OR2X2 OR2X2_512 ( .A(_abc_41356_new_n2028_), .B(regfil_4__3_), .Y(_abc_41356_new_n2184_));
OR2X2 OR2X2_513 ( .A(_abc_41356_new_n2027_), .B(wdatahold2_3_), .Y(_abc_41356_new_n2185_));
OR2X2 OR2X2_514 ( .A(_abc_41356_new_n2148_), .B(pc_11_), .Y(_abc_41356_new_n2190_));
OR2X2 OR2X2_515 ( .A(_abc_41356_new_n2049_), .B(pc_11_), .Y(_abc_41356_new_n2192_));
OR2X2 OR2X2_516 ( .A(_abc_41356_new_n2193_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n2194_));
OR2X2 OR2X2_517 ( .A(_abc_41356_new_n2158_), .B(pc_11_), .Y(_abc_41356_new_n2196_));
OR2X2 OR2X2_518 ( .A(_abc_41356_new_n2204_), .B(_abc_41356_new_n2203_), .Y(_abc_41356_new_n2205_));
OR2X2 OR2X2_519 ( .A(_abc_41356_new_n2206_), .B(_abc_41356_new_n2202_), .Y(_abc_41356_new_n2207_));
OR2X2 OR2X2_52 ( .A(_abc_41356_new_n752_), .B(_abc_41356_new_n751_), .Y(_abc_41356_new_n753_));
OR2X2 OR2X2_520 ( .A(_abc_41356_new_n2208_), .B(_abc_41356_new_n2209_), .Y(_abc_41356_new_n2210_));
OR2X2 OR2X2_521 ( .A(_abc_41356_new_n2210_), .B(_abc_41356_new_n2201_), .Y(_abc_41356_new_n2211_));
OR2X2 OR2X2_522 ( .A(_abc_41356_new_n2200_), .B(_abc_41356_new_n2211_), .Y(_abc_41356_new_n2212_));
OR2X2 OR2X2_523 ( .A(_abc_41356_new_n2212_), .B(_abc_41356_new_n2195_), .Y(_abc_41356_new_n2213_));
OR2X2 OR2X2_524 ( .A(_abc_41356_new_n2213_), .B(_abc_41356_new_n2069_), .Y(_abc_41356_new_n2214_));
OR2X2 OR2X2_525 ( .A(_abc_41356_new_n2096_), .B(wdatahold2_3_), .Y(_abc_41356_new_n2215_));
OR2X2 OR2X2_526 ( .A(_abc_41356_new_n2217_), .B(_abc_41356_new_n2187_), .Y(_abc_41356_new_n2218_));
OR2X2 OR2X2_527 ( .A(_abc_41356_new_n2219_), .B(_abc_41356_new_n2183_), .Y(_0wdatahold2_7_0__3_));
OR2X2 OR2X2_528 ( .A(_abc_41356_new_n2027_), .B(wdatahold2_4_), .Y(_abc_41356_new_n2222_));
OR2X2 OR2X2_529 ( .A(_abc_41356_new_n2028_), .B(regfil_4__4_), .Y(_abc_41356_new_n2223_));
OR2X2 OR2X2_53 ( .A(_abc_41356_new_n750_), .B(_abc_41356_new_n753_), .Y(_abc_41356_new_n754_));
OR2X2 OR2X2_530 ( .A(_abc_41356_new_n2228_), .B(_abc_41356_new_n2226_), .Y(_abc_41356_new_n2229_));
OR2X2 OR2X2_531 ( .A(_abc_41356_new_n2049_), .B(pc_12_), .Y(_abc_41356_new_n2231_));
OR2X2 OR2X2_532 ( .A(_abc_41356_new_n2232_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n2233_));
OR2X2 OR2X2_533 ( .A(_abc_41356_new_n2235_), .B(_abc_41356_new_n2236_), .Y(_abc_41356_new_n2237_));
OR2X2 OR2X2_534 ( .A(_abc_41356_new_n2242_), .B(_abc_41356_new_n2241_), .Y(_abc_41356_new_n2243_));
OR2X2 OR2X2_535 ( .A(_abc_41356_new_n2244_), .B(_abc_41356_new_n2240_), .Y(_abc_41356_new_n2245_));
OR2X2 OR2X2_536 ( .A(_abc_41356_new_n2247_), .B(_abc_41356_new_n2249_), .Y(_abc_41356_new_n2250_));
OR2X2 OR2X2_537 ( .A(_abc_41356_new_n2250_), .B(_abc_41356_new_n2246_), .Y(_abc_41356_new_n2251_));
OR2X2 OR2X2_538 ( .A(_abc_41356_new_n2239_), .B(_abc_41356_new_n2251_), .Y(_abc_41356_new_n2252_));
OR2X2 OR2X2_539 ( .A(_abc_41356_new_n2252_), .B(_abc_41356_new_n2234_), .Y(_abc_41356_new_n2253_));
OR2X2 OR2X2_54 ( .A(_abc_41356_new_n754_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n755_));
OR2X2 OR2X2_540 ( .A(_abc_41356_new_n2253_), .B(_abc_41356_new_n2069_), .Y(_abc_41356_new_n2254_));
OR2X2 OR2X2_541 ( .A(_abc_41356_new_n2096_), .B(wdatahold2_4_), .Y(_abc_41356_new_n2255_));
OR2X2 OR2X2_542 ( .A(_abc_41356_new_n2257_), .B(_abc_41356_new_n2225_), .Y(_abc_41356_new_n2258_));
OR2X2 OR2X2_543 ( .A(_abc_41356_new_n2259_), .B(_abc_41356_new_n2221_), .Y(_0wdatahold2_7_0__4_));
OR2X2 OR2X2_544 ( .A(_abc_41356_new_n2027_), .B(wdatahold2_5_), .Y(_abc_41356_new_n2262_));
OR2X2 OR2X2_545 ( .A(_abc_41356_new_n2028_), .B(regfil_4__5_), .Y(_abc_41356_new_n2263_));
OR2X2 OR2X2_546 ( .A(_abc_41356_new_n2226_), .B(pc_13_), .Y(_abc_41356_new_n2268_));
OR2X2 OR2X2_547 ( .A(_abc_41356_new_n2049_), .B(pc_13_), .Y(_abc_41356_new_n2270_));
OR2X2 OR2X2_548 ( .A(_abc_41356_new_n2271_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n2272_));
OR2X2 OR2X2_549 ( .A(_abc_41356_new_n2236_), .B(pc_13_), .Y(_abc_41356_new_n2274_));
OR2X2 OR2X2_55 ( .A(_abc_41356_new_n756_), .B(_abc_41356_new_n757_), .Y(_abc_41356_new_n758_));
OR2X2 OR2X2_550 ( .A(_abc_41356_new_n2283_), .B(_abc_41356_new_n2282_), .Y(_abc_41356_new_n2284_));
OR2X2 OR2X2_551 ( .A(_abc_41356_new_n2285_), .B(_abc_41356_new_n2281_), .Y(_abc_41356_new_n2286_));
OR2X2 OR2X2_552 ( .A(_abc_41356_new_n2287_), .B(_abc_41356_new_n2280_), .Y(_abc_41356_new_n2288_));
OR2X2 OR2X2_553 ( .A(_abc_41356_new_n2288_), .B(_abc_41356_new_n2279_), .Y(_abc_41356_new_n2289_));
OR2X2 OR2X2_554 ( .A(_abc_41356_new_n2278_), .B(_abc_41356_new_n2289_), .Y(_abc_41356_new_n2290_));
OR2X2 OR2X2_555 ( .A(_abc_41356_new_n2290_), .B(_abc_41356_new_n2273_), .Y(_abc_41356_new_n2291_));
OR2X2 OR2X2_556 ( .A(_abc_41356_new_n2291_), .B(_abc_41356_new_n2069_), .Y(_abc_41356_new_n2292_));
OR2X2 OR2X2_557 ( .A(_abc_41356_new_n2096_), .B(wdatahold2_5_), .Y(_abc_41356_new_n2293_));
OR2X2 OR2X2_558 ( .A(_abc_41356_new_n2295_), .B(_abc_41356_new_n2265_), .Y(_abc_41356_new_n2296_));
OR2X2 OR2X2_559 ( .A(_abc_41356_new_n2297_), .B(_abc_41356_new_n2261_), .Y(_0wdatahold2_7_0__5_));
OR2X2 OR2X2_56 ( .A(_abc_41356_new_n760_), .B(_abc_41356_new_n759_), .Y(_abc_41356_new_n761_));
OR2X2 OR2X2_560 ( .A(_abc_41356_new_n2028_), .B(regfil_4__6_), .Y(_abc_41356_new_n2300_));
OR2X2 OR2X2_561 ( .A(_abc_41356_new_n2027_), .B(wdatahold2_6_), .Y(_abc_41356_new_n2301_));
OR2X2 OR2X2_562 ( .A(_abc_41356_new_n2266_), .B(pc_14_), .Y(_abc_41356_new_n2306_));
OR2X2 OR2X2_563 ( .A(_abc_41356_new_n2049_), .B(pc_14_), .Y(_abc_41356_new_n2308_));
OR2X2 OR2X2_564 ( .A(_abc_41356_new_n2309_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n2310_));
OR2X2 OR2X2_565 ( .A(_abc_41356_new_n2275_), .B(pc_14_), .Y(_abc_41356_new_n2312_));
OR2X2 OR2X2_566 ( .A(_abc_41356_new_n2319_), .B(_abc_41356_new_n2318_), .Y(_abc_41356_new_n2320_));
OR2X2 OR2X2_567 ( .A(_abc_41356_new_n2321_), .B(_abc_41356_new_n2317_), .Y(_abc_41356_new_n2322_));
OR2X2 OR2X2_568 ( .A(_abc_41356_new_n2324_), .B(_abc_41356_new_n2325_), .Y(_abc_41356_new_n2326_));
OR2X2 OR2X2_569 ( .A(_abc_41356_new_n2326_), .B(_abc_41356_new_n2323_), .Y(_abc_41356_new_n2327_));
OR2X2 OR2X2_57 ( .A(_abc_41356_new_n758_), .B(_abc_41356_new_n761_), .Y(_abc_41356_new_n762_));
OR2X2 OR2X2_570 ( .A(_abc_41356_new_n2316_), .B(_abc_41356_new_n2327_), .Y(_abc_41356_new_n2328_));
OR2X2 OR2X2_571 ( .A(_abc_41356_new_n2328_), .B(_abc_41356_new_n2311_), .Y(_abc_41356_new_n2329_));
OR2X2 OR2X2_572 ( .A(_abc_41356_new_n2329_), .B(_abc_41356_new_n2069_), .Y(_abc_41356_new_n2330_));
OR2X2 OR2X2_573 ( .A(_abc_41356_new_n2096_), .B(wdatahold2_6_), .Y(_abc_41356_new_n2331_));
OR2X2 OR2X2_574 ( .A(_abc_41356_new_n2333_), .B(_abc_41356_new_n2303_), .Y(_abc_41356_new_n2334_));
OR2X2 OR2X2_575 ( .A(_abc_41356_new_n2335_), .B(_abc_41356_new_n2299_), .Y(_0wdatahold2_7_0__6_));
OR2X2 OR2X2_576 ( .A(_abc_41356_new_n2027_), .B(wdatahold2_7_), .Y(_abc_41356_new_n2338_));
OR2X2 OR2X2_577 ( .A(_abc_41356_new_n2028_), .B(regfil_4__7_), .Y(_abc_41356_new_n2339_));
OR2X2 OR2X2_578 ( .A(_abc_41356_new_n2304_), .B(pc_15_), .Y(_abc_41356_new_n2342_));
OR2X2 OR2X2_579 ( .A(_abc_41356_new_n2049_), .B(pc_15_), .Y(_abc_41356_new_n2346_));
OR2X2 OR2X2_58 ( .A(_abc_41356_new_n762_), .B(opcode_2_), .Y(_abc_41356_new_n763_));
OR2X2 OR2X2_580 ( .A(_abc_41356_new_n2347_), .B(_abc_41356_new_n2046_), .Y(_abc_41356_new_n2348_));
OR2X2 OR2X2_581 ( .A(_abc_41356_new_n2313_), .B(pc_15_), .Y(_abc_41356_new_n2350_));
OR2X2 OR2X2_582 ( .A(_abc_41356_new_n2359_), .B(_abc_41356_new_n2358_), .Y(_abc_41356_new_n2360_));
OR2X2 OR2X2_583 ( .A(_abc_41356_new_n2361_), .B(_abc_41356_new_n2357_), .Y(_abc_41356_new_n2362_));
OR2X2 OR2X2_584 ( .A(_abc_41356_new_n2363_), .B(_abc_41356_new_n2356_), .Y(_abc_41356_new_n2364_));
OR2X2 OR2X2_585 ( .A(_abc_41356_new_n2364_), .B(_abc_41356_new_n2355_), .Y(_abc_41356_new_n2365_));
OR2X2 OR2X2_586 ( .A(_abc_41356_new_n2354_), .B(_abc_41356_new_n2365_), .Y(_abc_41356_new_n2366_));
OR2X2 OR2X2_587 ( .A(_abc_41356_new_n2366_), .B(_abc_41356_new_n2349_), .Y(_abc_41356_new_n2367_));
OR2X2 OR2X2_588 ( .A(_abc_41356_new_n2367_), .B(_abc_41356_new_n2069_), .Y(_abc_41356_new_n2368_));
OR2X2 OR2X2_589 ( .A(_abc_41356_new_n2096_), .B(wdatahold2_7_), .Y(_abc_41356_new_n2369_));
OR2X2 OR2X2_59 ( .A(_abc_41356_new_n765_), .B(_abc_41356_new_n766_), .Y(_abc_41356_new_n767_));
OR2X2 OR2X2_590 ( .A(_abc_41356_new_n2371_), .B(_abc_41356_new_n2341_), .Y(_abc_41356_new_n2372_));
OR2X2 OR2X2_591 ( .A(_abc_41356_new_n2373_), .B(_abc_41356_new_n2337_), .Y(_0wdatahold2_7_0__7_));
OR2X2 OR2X2_592 ( .A(_abc_41356_new_n2379_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n2380_));
OR2X2 OR2X2_593 ( .A(_abc_41356_new_n1236_), .B(regfil_5__0_), .Y(_abc_41356_new_n2381_));
OR2X2 OR2X2_594 ( .A(_abc_41356_new_n663_), .B(_abc_41356_new_n2386_), .Y(_abc_41356_new_n2387_));
OR2X2 OR2X2_595 ( .A(_abc_41356_new_n2392_), .B(_abc_41356_new_n2389_), .Y(_abc_41356_new_n2393_));
OR2X2 OR2X2_596 ( .A(_abc_41356_new_n2378_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n2394_));
OR2X2 OR2X2_597 ( .A(_abc_41356_new_n2394_), .B(_abc_41356_new_n2393_), .Y(_abc_41356_new_n2395_));
OR2X2 OR2X2_598 ( .A(_abc_41356_new_n2385_), .B(regfil_3__0_), .Y(_abc_41356_new_n2397_));
OR2X2 OR2X2_599 ( .A(_abc_41356_new_n2399_), .B(_abc_41356_new_n2400_), .Y(_abc_41356_new_n2401_));
OR2X2 OR2X2_6 ( .A(_abc_41356_new_n553_), .B(_abc_41356_new_n560_), .Y(_abc_41356_new_n561_));
OR2X2 OR2X2_60 ( .A(_abc_41356_new_n768_), .B(_abc_41356_new_n747_), .Y(_abc_41356_new_n769_));
OR2X2 OR2X2_600 ( .A(_abc_41356_new_n2401_), .B(_abc_41356_new_n2382_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_0_));
OR2X2 OR2X2_601 ( .A(_abc_41356_new_n771_), .B(_abc_41356_new_n2386_), .Y(_abc_41356_new_n2403_));
OR2X2 OR2X2_602 ( .A(_abc_41356_new_n2385_), .B(regfil_3__1_), .Y(_abc_41356_new_n2404_));
OR2X2 OR2X2_603 ( .A(_abc_41356_new_n2410_), .B(_abc_41356_new_n2408_), .Y(_abc_41356_new_n2411_));
OR2X2 OR2X2_604 ( .A(_abc_41356_new_n2416_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n2417_));
OR2X2 OR2X2_605 ( .A(_abc_41356_new_n2417_), .B(_abc_41356_new_n2413_), .Y(_abc_41356_new_n2418_));
OR2X2 OR2X2_606 ( .A(_abc_41356_new_n1236_), .B(regfil_5__1_), .Y(_abc_41356_new_n2423_));
OR2X2 OR2X2_607 ( .A(_abc_41356_new_n2425_), .B(_abc_41356_new_n2407_), .Y(_abc_41356_new_n2426_));
OR2X2 OR2X2_608 ( .A(_abc_41356_new_n2406_), .B(_abc_41356_new_n2426_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_1_));
OR2X2 OR2X2_609 ( .A(_abc_41356_new_n824_), .B(_abc_41356_new_n2386_), .Y(_abc_41356_new_n2428_));
OR2X2 OR2X2_61 ( .A(_abc_41356_new_n746_), .B(_abc_41356_new_n769_), .Y(_abc_41356_new_n770_));
OR2X2 OR2X2_610 ( .A(_abc_41356_new_n2385_), .B(regfil_3__2_), .Y(_abc_41356_new_n2429_));
OR2X2 OR2X2_611 ( .A(_abc_41356_new_n2435_), .B(_abc_41356_new_n2433_), .Y(_abc_41356_new_n2436_));
OR2X2 OR2X2_612 ( .A(_abc_41356_new_n2408_), .B(regfil_3__2_), .Y(_abc_41356_new_n2438_));
OR2X2 OR2X2_613 ( .A(_abc_41356_new_n2437_), .B(_abc_41356_new_n2442_), .Y(_abc_41356_new_n2443_));
OR2X2 OR2X2_614 ( .A(_abc_41356_new_n2443_), .B(_abc_41356_new_n2444_), .Y(_abc_41356_new_n2445_));
OR2X2 OR2X2_615 ( .A(_abc_41356_new_n2445_), .B(_abc_41356_new_n2432_), .Y(_abc_41356_new_n2446_));
OR2X2 OR2X2_616 ( .A(_abc_41356_new_n2431_), .B(_abc_41356_new_n2446_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_2_));
OR2X2 OR2X2_617 ( .A(_abc_41356_new_n885_), .B(_abc_41356_new_n2386_), .Y(_abc_41356_new_n2448_));
OR2X2 OR2X2_618 ( .A(_abc_41356_new_n2385_), .B(regfil_3__3_), .Y(_abc_41356_new_n2449_));
OR2X2 OR2X2_619 ( .A(_abc_41356_new_n2455_), .B(_abc_41356_new_n2453_), .Y(_abc_41356_new_n2456_));
OR2X2 OR2X2_62 ( .A(_abc_41356_new_n741_), .B(_abc_41356_new_n770_), .Y(_abc_41356_new_n771_));
OR2X2 OR2X2_620 ( .A(_abc_41356_new_n2439_), .B(regfil_3__3_), .Y(_abc_41356_new_n2458_));
OR2X2 OR2X2_621 ( .A(_abc_41356_new_n2457_), .B(_abc_41356_new_n2462_), .Y(_abc_41356_new_n2463_));
OR2X2 OR2X2_622 ( .A(_abc_41356_new_n2463_), .B(_abc_41356_new_n2464_), .Y(_abc_41356_new_n2465_));
OR2X2 OR2X2_623 ( .A(_abc_41356_new_n2465_), .B(_abc_41356_new_n2452_), .Y(_abc_41356_new_n2466_));
OR2X2 OR2X2_624 ( .A(_abc_41356_new_n2451_), .B(_abc_41356_new_n2466_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_3_));
OR2X2 OR2X2_625 ( .A(_abc_41356_new_n952_), .B(_abc_41356_new_n2386_), .Y(_abc_41356_new_n2468_));
OR2X2 OR2X2_626 ( .A(_abc_41356_new_n2385_), .B(regfil_3__4_), .Y(_abc_41356_new_n2469_));
OR2X2 OR2X2_627 ( .A(_abc_41356_new_n2473_), .B(regfil_3__4_), .Y(_abc_41356_new_n2474_));
OR2X2 OR2X2_628 ( .A(_abc_41356_new_n2475_), .B(_abc_41356_new_n2476_), .Y(_abc_41356_new_n2477_));
OR2X2 OR2X2_629 ( .A(_abc_41356_new_n2459_), .B(regfil_3__4_), .Y(_abc_41356_new_n2479_));
OR2X2 OR2X2_63 ( .A(_abc_41356_new_n771_), .B(_abc_41356_new_n696_), .Y(_abc_41356_new_n772_));
OR2X2 OR2X2_630 ( .A(_abc_41356_new_n2478_), .B(_abc_41356_new_n2483_), .Y(_abc_41356_new_n2484_));
OR2X2 OR2X2_631 ( .A(_abc_41356_new_n2484_), .B(_abc_41356_new_n2485_), .Y(_abc_41356_new_n2486_));
OR2X2 OR2X2_632 ( .A(_abc_41356_new_n2486_), .B(_abc_41356_new_n2472_), .Y(_abc_41356_new_n2487_));
OR2X2 OR2X2_633 ( .A(_abc_41356_new_n2471_), .B(_abc_41356_new_n2487_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_4_));
OR2X2 OR2X2_634 ( .A(_abc_41356_new_n1019_), .B(_abc_41356_new_n2386_), .Y(_abc_41356_new_n2489_));
OR2X2 OR2X2_635 ( .A(_abc_41356_new_n2385_), .B(regfil_3__5_), .Y(_abc_41356_new_n2490_));
OR2X2 OR2X2_636 ( .A(_abc_41356_new_n2474_), .B(regfil_3__5_), .Y(_abc_41356_new_n2494_));
OR2X2 OR2X2_637 ( .A(_abc_41356_new_n2495_), .B(_abc_41356_new_n2496_), .Y(_abc_41356_new_n2497_));
OR2X2 OR2X2_638 ( .A(_abc_41356_new_n2480_), .B(regfil_3__5_), .Y(_abc_41356_new_n2501_));
OR2X2 OR2X2_639 ( .A(_abc_41356_new_n2498_), .B(_abc_41356_new_n2503_), .Y(_abc_41356_new_n2504_));
OR2X2 OR2X2_64 ( .A(_abc_41356_new_n695_), .B(regfil_7__1_), .Y(_abc_41356_new_n773_));
OR2X2 OR2X2_640 ( .A(_abc_41356_new_n2504_), .B(_abc_41356_new_n2505_), .Y(_abc_41356_new_n2506_));
OR2X2 OR2X2_641 ( .A(_abc_41356_new_n2506_), .B(_abc_41356_new_n2493_), .Y(_abc_41356_new_n2507_));
OR2X2 OR2X2_642 ( .A(_abc_41356_new_n2492_), .B(_abc_41356_new_n2507_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_5_));
OR2X2 OR2X2_643 ( .A(_abc_41356_new_n1091_), .B(_abc_41356_new_n2386_), .Y(_abc_41356_new_n2509_));
OR2X2 OR2X2_644 ( .A(_abc_41356_new_n2385_), .B(regfil_3__6_), .Y(_abc_41356_new_n2510_));
OR2X2 OR2X2_645 ( .A(_abc_41356_new_n2494_), .B(regfil_3__6_), .Y(_abc_41356_new_n2514_));
OR2X2 OR2X2_646 ( .A(_abc_41356_new_n2515_), .B(_abc_41356_new_n2516_), .Y(_abc_41356_new_n2517_));
OR2X2 OR2X2_647 ( .A(_abc_41356_new_n2499_), .B(regfil_3__6_), .Y(_abc_41356_new_n2521_));
OR2X2 OR2X2_648 ( .A(_abc_41356_new_n2518_), .B(_abc_41356_new_n2523_), .Y(_abc_41356_new_n2524_));
OR2X2 OR2X2_649 ( .A(_abc_41356_new_n2524_), .B(_abc_41356_new_n2525_), .Y(_abc_41356_new_n2526_));
OR2X2 OR2X2_65 ( .A(_abc_41356_new_n778_), .B(_abc_41356_new_n777_), .Y(_abc_41356_new_n779_));
OR2X2 OR2X2_650 ( .A(_abc_41356_new_n2526_), .B(_abc_41356_new_n2513_), .Y(_abc_41356_new_n2527_));
OR2X2 OR2X2_651 ( .A(_abc_41356_new_n2512_), .B(_abc_41356_new_n2527_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_6_));
OR2X2 OR2X2_652 ( .A(_abc_41356_new_n1173_), .B(_abc_41356_new_n2386_), .Y(_abc_41356_new_n2529_));
OR2X2 OR2X2_653 ( .A(_abc_41356_new_n2385_), .B(regfil_3__7_), .Y(_abc_41356_new_n2530_));
OR2X2 OR2X2_654 ( .A(_abc_41356_new_n2514_), .B(regfil_3__7_), .Y(_abc_41356_new_n2534_));
OR2X2 OR2X2_655 ( .A(_abc_41356_new_n2535_), .B(_abc_41356_new_n2536_), .Y(_abc_41356_new_n2537_));
OR2X2 OR2X2_656 ( .A(_abc_41356_new_n2519_), .B(regfil_3__7_), .Y(_abc_41356_new_n2539_));
OR2X2 OR2X2_657 ( .A(_abc_41356_new_n2538_), .B(_abc_41356_new_n2543_), .Y(_abc_41356_new_n2544_));
OR2X2 OR2X2_658 ( .A(_abc_41356_new_n2544_), .B(_abc_41356_new_n2545_), .Y(_abc_41356_new_n2546_));
OR2X2 OR2X2_659 ( .A(_abc_41356_new_n2546_), .B(_abc_41356_new_n2533_), .Y(_abc_41356_new_n2547_));
OR2X2 OR2X2_66 ( .A(_abc_41356_new_n779_), .B(_abc_41356_new_n776_), .Y(_abc_41356_new_n780_));
OR2X2 OR2X2_660 ( .A(_abc_41356_new_n2532_), .B(_abc_41356_new_n2547_), .Y(_abc_36060_memoryregfil_wrmux_3__2__0__y_16089_7_));
OR2X2 OR2X2_661 ( .A(_abc_41356_new_n663_), .B(_abc_41356_new_n2551_), .Y(_abc_41356_new_n2552_));
OR2X2 OR2X2_662 ( .A(_abc_41356_new_n2550_), .B(regfil_1__0_), .Y(_abc_41356_new_n2553_));
OR2X2 OR2X2_663 ( .A(_abc_41356_new_n2559_), .B(_abc_41356_new_n2560_), .Y(_abc_41356_new_n2561_));
OR2X2 OR2X2_664 ( .A(_abc_41356_new_n2555_), .B(_abc_41356_new_n2561_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_0_));
OR2X2 OR2X2_665 ( .A(_abc_41356_new_n771_), .B(_abc_41356_new_n2551_), .Y(_abc_41356_new_n2563_));
OR2X2 OR2X2_666 ( .A(_abc_41356_new_n2550_), .B(regfil_1__1_), .Y(_abc_41356_new_n2564_));
OR2X2 OR2X2_667 ( .A(_abc_41356_new_n649_), .B(_abc_41356_new_n568_), .Y(_abc_41356_new_n2567_));
OR2X2 OR2X2_668 ( .A(_abc_41356_new_n581_), .B(_abc_41356_new_n2567_), .Y(_abc_41356_new_n2568_));
OR2X2 OR2X2_669 ( .A(_abc_41356_new_n601_), .B(_abc_41356_new_n2569_), .Y(_abc_41356_new_n2570_));
OR2X2 OR2X2_67 ( .A(_abc_41356_new_n783_), .B(_abc_41356_new_n784_), .Y(_abc_41356_new_n785_));
OR2X2 OR2X2_670 ( .A(_abc_41356_new_n2572_), .B(_abc_41356_new_n2573_), .Y(_abc_41356_new_n2574_));
OR2X2 OR2X2_671 ( .A(_abc_41356_new_n2566_), .B(_abc_41356_new_n2574_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_1_));
OR2X2 OR2X2_672 ( .A(_abc_41356_new_n824_), .B(_abc_41356_new_n2551_), .Y(_abc_41356_new_n2576_));
OR2X2 OR2X2_673 ( .A(_abc_41356_new_n2550_), .B(regfil_1__2_), .Y(_abc_41356_new_n2577_));
OR2X2 OR2X2_674 ( .A(_abc_41356_new_n2581_), .B(_abc_41356_new_n650_), .Y(_abc_41356_new_n2582_));
OR2X2 OR2X2_675 ( .A(_abc_41356_new_n568_), .B(regfil_1__2_), .Y(_abc_41356_new_n2585_));
OR2X2 OR2X2_676 ( .A(_abc_41356_new_n2583_), .B(_abc_41356_new_n2587_), .Y(_abc_41356_new_n2588_));
OR2X2 OR2X2_677 ( .A(_abc_41356_new_n2588_), .B(_abc_41356_new_n2589_), .Y(_abc_41356_new_n2590_));
OR2X2 OR2X2_678 ( .A(_abc_41356_new_n2579_), .B(_abc_41356_new_n2590_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_2_));
OR2X2 OR2X2_679 ( .A(_abc_41356_new_n885_), .B(_abc_41356_new_n2551_), .Y(_abc_41356_new_n2592_));
OR2X2 OR2X2_68 ( .A(_abc_41356_new_n785_), .B(_abc_41356_new_n782_), .Y(_abc_41356_new_n786_));
OR2X2 OR2X2_680 ( .A(_abc_41356_new_n2550_), .B(regfil_1__3_), .Y(_abc_41356_new_n2593_));
OR2X2 OR2X2_681 ( .A(_abc_41356_new_n2597_), .B(_abc_41356_new_n651_), .Y(_abc_41356_new_n2598_));
OR2X2 OR2X2_682 ( .A(_abc_41356_new_n569_), .B(regfil_1__3_), .Y(_abc_41356_new_n2601_));
OR2X2 OR2X2_683 ( .A(_abc_41356_new_n2599_), .B(_abc_41356_new_n2603_), .Y(_abc_41356_new_n2604_));
OR2X2 OR2X2_684 ( .A(_abc_41356_new_n2604_), .B(_abc_41356_new_n2605_), .Y(_abc_41356_new_n2606_));
OR2X2 OR2X2_685 ( .A(_abc_41356_new_n2595_), .B(_abc_41356_new_n2606_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_3_));
OR2X2 OR2X2_686 ( .A(_abc_41356_new_n952_), .B(_abc_41356_new_n2551_), .Y(_abc_41356_new_n2608_));
OR2X2 OR2X2_687 ( .A(_abc_41356_new_n2550_), .B(regfil_1__4_), .Y(_abc_41356_new_n2609_));
OR2X2 OR2X2_688 ( .A(_abc_41356_new_n2612_), .B(_abc_41356_new_n2613_), .Y(_abc_41356_new_n2614_));
OR2X2 OR2X2_689 ( .A(_abc_41356_new_n570_), .B(regfil_1__4_), .Y(_abc_41356_new_n2617_));
OR2X2 OR2X2_69 ( .A(_abc_41356_new_n786_), .B(_abc_41356_new_n781_), .Y(_abc_41356_new_n787_));
OR2X2 OR2X2_690 ( .A(_abc_41356_new_n2615_), .B(_abc_41356_new_n2619_), .Y(_abc_41356_new_n2620_));
OR2X2 OR2X2_691 ( .A(_abc_41356_new_n2620_), .B(_abc_41356_new_n2621_), .Y(_abc_41356_new_n2622_));
OR2X2 OR2X2_692 ( .A(_abc_41356_new_n2611_), .B(_abc_41356_new_n2622_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_4_));
OR2X2 OR2X2_693 ( .A(_abc_41356_new_n1019_), .B(_abc_41356_new_n2551_), .Y(_abc_41356_new_n2624_));
OR2X2 OR2X2_694 ( .A(_abc_41356_new_n2550_), .B(regfil_1__5_), .Y(_abc_41356_new_n2625_));
OR2X2 OR2X2_695 ( .A(_abc_41356_new_n2628_), .B(_abc_41356_new_n2629_), .Y(_abc_41356_new_n2630_));
OR2X2 OR2X2_696 ( .A(_abc_41356_new_n571_), .B(regfil_1__5_), .Y(_abc_41356_new_n2633_));
OR2X2 OR2X2_697 ( .A(_abc_41356_new_n2631_), .B(_abc_41356_new_n2635_), .Y(_abc_41356_new_n2636_));
OR2X2 OR2X2_698 ( .A(_abc_41356_new_n2636_), .B(_abc_41356_new_n2637_), .Y(_abc_41356_new_n2638_));
OR2X2 OR2X2_699 ( .A(_abc_41356_new_n2627_), .B(_abc_41356_new_n2638_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_5_));
OR2X2 OR2X2_7 ( .A(_abc_41356_new_n562_), .B(_abc_41356_new_n512_), .Y(_abc_41356_new_n563_));
OR2X2 OR2X2_70 ( .A(_abc_41356_new_n780_), .B(_abc_41356_new_n787_), .Y(_abc_41356_new_n788_));
OR2X2 OR2X2_700 ( .A(_abc_41356_new_n1091_), .B(_abc_41356_new_n2551_), .Y(_abc_41356_new_n2640_));
OR2X2 OR2X2_701 ( .A(_abc_41356_new_n2550_), .B(regfil_1__6_), .Y(_abc_41356_new_n2641_));
OR2X2 OR2X2_702 ( .A(_abc_41356_new_n2645_), .B(_abc_41356_new_n2646_), .Y(_abc_41356_new_n2647_));
OR2X2 OR2X2_703 ( .A(_abc_41356_new_n572_), .B(regfil_1__6_), .Y(_abc_41356_new_n2649_));
OR2X2 OR2X2_704 ( .A(_abc_41356_new_n2648_), .B(_abc_41356_new_n2652_), .Y(_abc_41356_new_n2653_));
OR2X2 OR2X2_705 ( .A(_abc_41356_new_n2653_), .B(_abc_41356_new_n2644_), .Y(_abc_41356_new_n2654_));
OR2X2 OR2X2_706 ( .A(_abc_41356_new_n2643_), .B(_abc_41356_new_n2654_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_6_));
OR2X2 OR2X2_707 ( .A(_abc_41356_new_n1173_), .B(_abc_41356_new_n2551_), .Y(_abc_41356_new_n2656_));
OR2X2 OR2X2_708 ( .A(_abc_41356_new_n2550_), .B(regfil_1__7_), .Y(_abc_41356_new_n2657_));
OR2X2 OR2X2_709 ( .A(_abc_41356_new_n657_), .B(_abc_41356_new_n2661_), .Y(_abc_41356_new_n2662_));
OR2X2 OR2X2_71 ( .A(_abc_41356_new_n775_), .B(_abc_41356_new_n788_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_1_));
OR2X2 OR2X2_710 ( .A(_abc_41356_new_n573_), .B(regfil_1__7_), .Y(_abc_41356_new_n2664_));
OR2X2 OR2X2_711 ( .A(_abc_41356_new_n2663_), .B(_abc_41356_new_n2667_), .Y(_abc_41356_new_n2668_));
OR2X2 OR2X2_712 ( .A(_abc_41356_new_n2668_), .B(_abc_41356_new_n2660_), .Y(_abc_41356_new_n2669_));
OR2X2 OR2X2_713 ( .A(_abc_41356_new_n2659_), .B(_abc_41356_new_n2669_), .Y(_abc_36060_memoryregfil_wrmux_1__1__0__y_16001_7_));
OR2X2 OR2X2_714 ( .A(_abc_41356_new_n663_), .B(_abc_41356_new_n2672_), .Y(_abc_41356_new_n2673_));
OR2X2 OR2X2_715 ( .A(_abc_41356_new_n2671_), .B(regfil_6__0_), .Y(_abc_41356_new_n2674_));
OR2X2 OR2X2_716 ( .A(_abc_41356_new_n771_), .B(_abc_41356_new_n2672_), .Y(_abc_41356_new_n2676_));
OR2X2 OR2X2_717 ( .A(_abc_41356_new_n2671_), .B(regfil_6__1_), .Y(_abc_41356_new_n2677_));
OR2X2 OR2X2_718 ( .A(_abc_41356_new_n824_), .B(_abc_41356_new_n2672_), .Y(_abc_41356_new_n2679_));
OR2X2 OR2X2_719 ( .A(_abc_41356_new_n2671_), .B(regfil_6__2_), .Y(_abc_41356_new_n2680_));
OR2X2 OR2X2_72 ( .A(_abc_41356_new_n736_), .B(regfil_0__2_), .Y(_abc_41356_new_n790_));
OR2X2 OR2X2_720 ( .A(_abc_41356_new_n885_), .B(_abc_41356_new_n2672_), .Y(_abc_41356_new_n2682_));
OR2X2 OR2X2_721 ( .A(_abc_41356_new_n2671_), .B(regfil_6__3_), .Y(_abc_41356_new_n2683_));
OR2X2 OR2X2_722 ( .A(_abc_41356_new_n952_), .B(_abc_41356_new_n2672_), .Y(_abc_41356_new_n2685_));
OR2X2 OR2X2_723 ( .A(_abc_41356_new_n2671_), .B(regfil_6__4_), .Y(_abc_41356_new_n2686_));
OR2X2 OR2X2_724 ( .A(_abc_41356_new_n1019_), .B(_abc_41356_new_n2672_), .Y(_abc_41356_new_n2688_));
OR2X2 OR2X2_725 ( .A(_abc_41356_new_n2671_), .B(regfil_6__5_), .Y(_abc_41356_new_n2689_));
OR2X2 OR2X2_726 ( .A(_abc_41356_new_n1091_), .B(_abc_41356_new_n2672_), .Y(_abc_41356_new_n2691_));
OR2X2 OR2X2_727 ( .A(_abc_41356_new_n2671_), .B(regfil_6__6_), .Y(_abc_41356_new_n2692_));
OR2X2 OR2X2_728 ( .A(_abc_41356_new_n1173_), .B(_abc_41356_new_n2672_), .Y(_abc_41356_new_n2694_));
OR2X2 OR2X2_729 ( .A(_abc_41356_new_n2671_), .B(regfil_6__7_), .Y(_abc_41356_new_n2695_));
OR2X2 OR2X2_73 ( .A(_abc_41356_new_n791_), .B(_abc_41356_new_n792_), .Y(_abc_41356_new_n793_));
OR2X2 OR2X2_730 ( .A(_abc_41356_new_n663_), .B(_abc_41356_new_n2698_), .Y(_abc_41356_new_n2699_));
OR2X2 OR2X2_731 ( .A(_abc_41356_new_n2697_), .B(regfil_2__0_), .Y(_abc_41356_new_n2700_));
OR2X2 OR2X2_732 ( .A(_abc_41356_new_n2534_), .B(regfil_2__0_), .Y(_abc_41356_new_n2704_));
OR2X2 OR2X2_733 ( .A(_abc_41356_new_n2705_), .B(_abc_41356_new_n2706_), .Y(_abc_41356_new_n2707_));
OR2X2 OR2X2_734 ( .A(_abc_41356_new_n2540_), .B(regfil_2__0_), .Y(_abc_41356_new_n2709_));
OR2X2 OR2X2_735 ( .A(_abc_41356_new_n2708_), .B(_abc_41356_new_n2713_), .Y(_abc_41356_new_n2714_));
OR2X2 OR2X2_736 ( .A(_abc_41356_new_n2714_), .B(_abc_41356_new_n2715_), .Y(_abc_41356_new_n2716_));
OR2X2 OR2X2_737 ( .A(_abc_41356_new_n2716_), .B(_abc_41356_new_n2703_), .Y(_abc_41356_new_n2717_));
OR2X2 OR2X2_738 ( .A(_abc_41356_new_n2702_), .B(_abc_41356_new_n2717_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_0_));
OR2X2 OR2X2_739 ( .A(_abc_41356_new_n771_), .B(_abc_41356_new_n2698_), .Y(_abc_41356_new_n2719_));
OR2X2 OR2X2_74 ( .A(_abc_41356_new_n743_), .B(regfil_0__2_), .Y(_abc_41356_new_n795_));
OR2X2 OR2X2_740 ( .A(_abc_41356_new_n2697_), .B(regfil_2__1_), .Y(_abc_41356_new_n2720_));
OR2X2 OR2X2_741 ( .A(_abc_41356_new_n2704_), .B(regfil_2__1_), .Y(_abc_41356_new_n2724_));
OR2X2 OR2X2_742 ( .A(_abc_41356_new_n2725_), .B(_abc_41356_new_n2726_), .Y(_abc_41356_new_n2727_));
OR2X2 OR2X2_743 ( .A(_abc_41356_new_n2710_), .B(regfil_2__1_), .Y(_abc_41356_new_n2729_));
OR2X2 OR2X2_744 ( .A(_abc_41356_new_n2728_), .B(_abc_41356_new_n2733_), .Y(_abc_41356_new_n2734_));
OR2X2 OR2X2_745 ( .A(_abc_41356_new_n2734_), .B(_abc_41356_new_n2735_), .Y(_abc_41356_new_n2736_));
OR2X2 OR2X2_746 ( .A(_abc_41356_new_n2736_), .B(_abc_41356_new_n2723_), .Y(_abc_41356_new_n2737_));
OR2X2 OR2X2_747 ( .A(_abc_41356_new_n2722_), .B(_abc_41356_new_n2737_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_1_));
OR2X2 OR2X2_748 ( .A(_abc_41356_new_n824_), .B(_abc_41356_new_n2698_), .Y(_abc_41356_new_n2739_));
OR2X2 OR2X2_749 ( .A(_abc_41356_new_n2697_), .B(regfil_2__2_), .Y(_abc_41356_new_n2740_));
OR2X2 OR2X2_75 ( .A(_abc_41356_new_n802_), .B(_abc_41356_new_n801_), .Y(_abc_41356_new_n803_));
OR2X2 OR2X2_750 ( .A(_abc_41356_new_n2724_), .B(regfil_2__2_), .Y(_abc_41356_new_n2744_));
OR2X2 OR2X2_751 ( .A(_abc_41356_new_n2745_), .B(_abc_41356_new_n2746_), .Y(_abc_41356_new_n2747_));
OR2X2 OR2X2_752 ( .A(_abc_41356_new_n2730_), .B(regfil_2__2_), .Y(_abc_41356_new_n2749_));
OR2X2 OR2X2_753 ( .A(_abc_41356_new_n2748_), .B(_abc_41356_new_n2753_), .Y(_abc_41356_new_n2754_));
OR2X2 OR2X2_754 ( .A(_abc_41356_new_n2754_), .B(_abc_41356_new_n2755_), .Y(_abc_41356_new_n2756_));
OR2X2 OR2X2_755 ( .A(_abc_41356_new_n2756_), .B(_abc_41356_new_n2743_), .Y(_abc_41356_new_n2757_));
OR2X2 OR2X2_756 ( .A(_abc_41356_new_n2757_), .B(_abc_41356_new_n2742_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_2_));
OR2X2 OR2X2_757 ( .A(_abc_41356_new_n885_), .B(_abc_41356_new_n2698_), .Y(_abc_41356_new_n2759_));
OR2X2 OR2X2_758 ( .A(_abc_41356_new_n2697_), .B(regfil_2__3_), .Y(_abc_41356_new_n2760_));
OR2X2 OR2X2_759 ( .A(_abc_41356_new_n2750_), .B(regfil_2__3_), .Y(_abc_41356_new_n2766_));
OR2X2 OR2X2_76 ( .A(_abc_41356_new_n805_), .B(_abc_41356_new_n804_), .Y(_abc_41356_new_n806_));
OR2X2 OR2X2_760 ( .A(_abc_41356_new_n2744_), .B(regfil_2__3_), .Y(_abc_41356_new_n2769_));
OR2X2 OR2X2_761 ( .A(_abc_41356_new_n2770_), .B(_abc_41356_new_n2771_), .Y(_abc_41356_new_n2772_));
OR2X2 OR2X2_762 ( .A(_abc_41356_new_n2773_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n2774_));
OR2X2 OR2X2_763 ( .A(_abc_41356_new_n2774_), .B(_abc_41356_new_n2768_), .Y(_abc_41356_new_n2775_));
OR2X2 OR2X2_764 ( .A(_abc_41356_new_n1236_), .B(regfil_4__3_), .Y(_abc_41356_new_n2776_));
OR2X2 OR2X2_765 ( .A(_abc_41356_new_n2778_), .B(_abc_41356_new_n2763_), .Y(_abc_41356_new_n2779_));
OR2X2 OR2X2_766 ( .A(_abc_41356_new_n2779_), .B(_abc_41356_new_n2762_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_3_));
OR2X2 OR2X2_767 ( .A(_abc_41356_new_n952_), .B(_abc_41356_new_n2698_), .Y(_abc_41356_new_n2781_));
OR2X2 OR2X2_768 ( .A(_abc_41356_new_n2697_), .B(regfil_2__4_), .Y(_abc_41356_new_n2782_));
OR2X2 OR2X2_769 ( .A(_abc_41356_new_n2764_), .B(regfil_2__4_), .Y(_abc_41356_new_n2788_));
OR2X2 OR2X2_77 ( .A(_abc_41356_new_n803_), .B(_abc_41356_new_n806_), .Y(_abc_41356_new_n807_));
OR2X2 OR2X2_770 ( .A(_abc_41356_new_n2769_), .B(regfil_2__4_), .Y(_abc_41356_new_n2791_));
OR2X2 OR2X2_771 ( .A(_abc_41356_new_n2792_), .B(_abc_41356_new_n2793_), .Y(_abc_41356_new_n2794_));
OR2X2 OR2X2_772 ( .A(_abc_41356_new_n2795_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n2796_));
OR2X2 OR2X2_773 ( .A(_abc_41356_new_n2796_), .B(_abc_41356_new_n2790_), .Y(_abc_41356_new_n2797_));
OR2X2 OR2X2_774 ( .A(_abc_41356_new_n1236_), .B(regfil_4__4_), .Y(_abc_41356_new_n2798_));
OR2X2 OR2X2_775 ( .A(_abc_41356_new_n2800_), .B(_abc_41356_new_n2785_), .Y(_abc_41356_new_n2801_));
OR2X2 OR2X2_776 ( .A(_abc_41356_new_n2801_), .B(_abc_41356_new_n2784_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_4_));
OR2X2 OR2X2_777 ( .A(_abc_41356_new_n1019_), .B(_abc_41356_new_n2698_), .Y(_abc_41356_new_n2803_));
OR2X2 OR2X2_778 ( .A(_abc_41356_new_n2697_), .B(regfil_2__5_), .Y(_abc_41356_new_n2804_));
OR2X2 OR2X2_779 ( .A(_abc_41356_new_n2786_), .B(regfil_2__5_), .Y(_abc_41356_new_n2810_));
OR2X2 OR2X2_78 ( .A(_abc_41356_new_n807_), .B(opcode_2_), .Y(_abc_41356_new_n808_));
OR2X2 OR2X2_780 ( .A(_abc_41356_new_n2791_), .B(regfil_2__5_), .Y(_abc_41356_new_n2813_));
OR2X2 OR2X2_781 ( .A(_abc_41356_new_n2814_), .B(_abc_41356_new_n2815_), .Y(_abc_41356_new_n2816_));
OR2X2 OR2X2_782 ( .A(_abc_41356_new_n2817_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n2818_));
OR2X2 OR2X2_783 ( .A(_abc_41356_new_n2818_), .B(_abc_41356_new_n2812_), .Y(_abc_41356_new_n2819_));
OR2X2 OR2X2_784 ( .A(_abc_41356_new_n1236_), .B(regfil_4__5_), .Y(_abc_41356_new_n2820_));
OR2X2 OR2X2_785 ( .A(_abc_41356_new_n2822_), .B(_abc_41356_new_n2807_), .Y(_abc_41356_new_n2823_));
OR2X2 OR2X2_786 ( .A(_abc_41356_new_n2823_), .B(_abc_41356_new_n2806_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_5_));
OR2X2 OR2X2_787 ( .A(_abc_41356_new_n1091_), .B(_abc_41356_new_n2698_), .Y(_abc_41356_new_n2825_));
OR2X2 OR2X2_788 ( .A(_abc_41356_new_n2697_), .B(regfil_2__6_), .Y(_abc_41356_new_n2826_));
OR2X2 OR2X2_789 ( .A(_abc_41356_new_n2808_), .B(regfil_2__6_), .Y(_abc_41356_new_n2830_));
OR2X2 OR2X2_79 ( .A(_abc_41356_new_n809_), .B(_abc_41356_new_n577_), .Y(_abc_41356_new_n810_));
OR2X2 OR2X2_790 ( .A(_abc_41356_new_n2813_), .B(regfil_2__6_), .Y(_abc_41356_new_n2835_));
OR2X2 OR2X2_791 ( .A(_abc_41356_new_n2836_), .B(_abc_41356_new_n2837_), .Y(_abc_41356_new_n2838_));
OR2X2 OR2X2_792 ( .A(_abc_41356_new_n2839_), .B(_abc_41356_new_n1235_), .Y(_abc_41356_new_n2840_));
OR2X2 OR2X2_793 ( .A(_abc_41356_new_n2840_), .B(_abc_41356_new_n2834_), .Y(_abc_41356_new_n2841_));
OR2X2 OR2X2_794 ( .A(_abc_41356_new_n1236_), .B(regfil_4__6_), .Y(_abc_41356_new_n2842_));
OR2X2 OR2X2_795 ( .A(_abc_41356_new_n2844_), .B(_abc_41356_new_n2829_), .Y(_abc_41356_new_n2845_));
OR2X2 OR2X2_796 ( .A(_abc_41356_new_n2828_), .B(_abc_41356_new_n2845_), .Y(_abc_36060_memoryregfil_wrmux_2__1__0__y_16043_6_));
OR2X2 OR2X2_797 ( .A(_abc_41356_new_n2849_), .B(_abc_41356_new_n2395_), .Y(_abc_41356_new_n2850_));
OR2X2 OR2X2_798 ( .A(_abc_41356_new_n2848_), .B(_abc_41356_new_n2850_), .Y(_abc_41356_new_n2851_));
OR2X2 OR2X2_799 ( .A(_abc_41356_new_n2853_), .B(_abc_41356_new_n2852_), .Y(_abc_41356_new_n2854_));
OR2X2 OR2X2_8 ( .A(_abc_41356_new_n574_), .B(regfil_0__0_), .Y(_abc_41356_new_n575_));
OR2X2 OR2X2_80 ( .A(_abc_41356_new_n812_), .B(_abc_41356_new_n813_), .Y(_abc_41356_new_n814_));
OR2X2 OR2X2_800 ( .A(_abc_41356_new_n2836_), .B(_abc_41356_new_n2861_), .Y(_abc_41356_new_n2862_));
OR2X2 OR2X2_801 ( .A(_abc_41356_new_n2860_), .B(_abc_41356_new_n2865_), .Y(_abc_41356_new_n2866_));
OR2X2 OR2X2_802 ( .A(_abc_41356_new_n2868_), .B(_abc_41356_new_n2421_), .Y(_abc_41356_new_n2869_));
OR2X2 OR2X2_803 ( .A(_abc_41356_new_n2867_), .B(_abc_41356_new_n2869_), .Y(_abc_41356_new_n2870_));
OR2X2 OR2X2_804 ( .A(_abc_41356_new_n677_), .B(_abc_41356_new_n2022_), .Y(_abc_41356_new_n2881_));
OR2X2 OR2X2_805 ( .A(_abc_41356_new_n2020_), .B(_abc_41356_new_n2881_), .Y(_abc_41356_new_n2882_));
OR2X2 OR2X2_806 ( .A(_abc_41356_new_n2885_), .B(_abc_41356_new_n2893_), .Y(_0alusel_2_0__0_));
OR2X2 OR2X2_807 ( .A(_abc_41356_new_n678_), .B(opcode_4_), .Y(_abc_41356_new_n2895_));
OR2X2 OR2X2_808 ( .A(_abc_41356_new_n677_), .B(alu_sel_1_), .Y(_abc_41356_new_n2896_));
OR2X2 OR2X2_809 ( .A(_abc_41356_new_n2874_), .B(alu_sel_1_), .Y(_abc_41356_new_n2899_));
OR2X2 OR2X2_81 ( .A(_abc_41356_new_n814_), .B(_abc_41356_new_n811_), .Y(_abc_41356_new_n815_));
OR2X2 OR2X2_810 ( .A(_abc_41356_new_n2901_), .B(_abc_41356_new_n2902_), .Y(_abc_41356_new_n2903_));
OR2X2 OR2X2_811 ( .A(_abc_41356_new_n2903_), .B(_abc_41356_new_n2898_), .Y(_abc_41356_new_n2904_));
OR2X2 OR2X2_812 ( .A(_abc_41356_new_n2905_), .B(_abc_41356_new_n2907_), .Y(_0alusel_2_0__1_));
OR2X2 OR2X2_813 ( .A(_abc_41356_new_n677_), .B(alu_sel_2_), .Y(_abc_41356_new_n2912_));
OR2X2 OR2X2_814 ( .A(_abc_41356_new_n2913_), .B(_abc_41356_new_n2911_), .Y(_abc_41356_new_n2914_));
OR2X2 OR2X2_815 ( .A(_abc_41356_new_n678_), .B(opcode_5_), .Y(_abc_41356_new_n2915_));
OR2X2 OR2X2_816 ( .A(_abc_41356_new_n2910_), .B(_abc_41356_new_n2917_), .Y(_0alusel_2_0__2_));
OR2X2 OR2X2_817 ( .A(_abc_41356_new_n2919_), .B(alu_cin), .Y(_abc_41356_new_n2920_));
OR2X2 OR2X2_818 ( .A(_abc_41356_new_n2921_), .B(carry), .Y(_abc_41356_new_n2922_));
OR2X2 OR2X2_819 ( .A(_abc_41356_new_n636_), .B(_abc_41356_new_n2887_), .Y(_abc_41356_new_n2936_));
OR2X2 OR2X2_82 ( .A(_abc_41356_new_n815_), .B(_abc_41356_new_n810_), .Y(_abc_41356_new_n816_));
OR2X2 OR2X2_820 ( .A(_abc_41356_new_n2935_), .B(_abc_41356_new_n2937_), .Y(_abc_41356_new_n2938_));
OR2X2 OR2X2_821 ( .A(_abc_41356_new_n2876_), .B(opcode_6_), .Y(_abc_41356_new_n2939_));
OR2X2 OR2X2_822 ( .A(_abc_41356_new_n2940_), .B(alu_oprb_0_), .Y(_abc_41356_new_n2941_));
OR2X2 OR2X2_823 ( .A(_abc_41356_new_n2942_), .B(_abc_41356_new_n2932_), .Y(_0aluoprb_7_0__0_));
OR2X2 OR2X2_824 ( .A(_abc_41356_new_n2934_), .B(_abc_41356_new_n2944_), .Y(_abc_41356_new_n2945_));
OR2X2 OR2X2_825 ( .A(_abc_41356_new_n2949_), .B(_abc_41356_new_n2947_), .Y(_abc_41356_new_n2950_));
OR2X2 OR2X2_826 ( .A(_abc_41356_new_n2946_), .B(_abc_41356_new_n2950_), .Y(_0aluoprb_7_0__1_));
OR2X2 OR2X2_827 ( .A(_abc_41356_new_n2954_), .B(_abc_41356_new_n2953_), .Y(_abc_41356_new_n2955_));
OR2X2 OR2X2_828 ( .A(_abc_41356_new_n2952_), .B(_abc_41356_new_n2955_), .Y(_0aluoprb_7_0__2_));
OR2X2 OR2X2_829 ( .A(_abc_41356_new_n2957_), .B(_abc_41356_new_n2958_), .Y(_abc_41356_new_n2959_));
OR2X2 OR2X2_83 ( .A(_abc_41356_new_n818_), .B(_abc_41356_new_n819_), .Y(_abc_41356_new_n820_));
OR2X2 OR2X2_830 ( .A(_abc_41356_new_n2961_), .B(_abc_41356_new_n2962_), .Y(_abc_41356_new_n2963_));
OR2X2 OR2X2_831 ( .A(_abc_41356_new_n2963_), .B(_abc_41356_new_n2960_), .Y(_0aluoprb_7_0__3_));
OR2X2 OR2X2_832 ( .A(_abc_41356_new_n2967_), .B(_abc_41356_new_n2966_), .Y(_abc_41356_new_n2968_));
OR2X2 OR2X2_833 ( .A(_abc_41356_new_n2965_), .B(_abc_41356_new_n2968_), .Y(_0aluoprb_7_0__4_));
OR2X2 OR2X2_834 ( .A(_abc_41356_new_n2972_), .B(_abc_41356_new_n2971_), .Y(_abc_41356_new_n2973_));
OR2X2 OR2X2_835 ( .A(_abc_41356_new_n2970_), .B(_abc_41356_new_n2973_), .Y(_0aluoprb_7_0__5_));
OR2X2 OR2X2_836 ( .A(_abc_41356_new_n2975_), .B(_abc_41356_new_n2976_), .Y(_abc_41356_new_n2977_));
OR2X2 OR2X2_837 ( .A(_abc_41356_new_n2980_), .B(_abc_41356_new_n2979_), .Y(_abc_41356_new_n2981_));
OR2X2 OR2X2_838 ( .A(_abc_41356_new_n2981_), .B(_abc_41356_new_n2978_), .Y(_0aluoprb_7_0__6_));
OR2X2 OR2X2_839 ( .A(_abc_41356_new_n2985_), .B(_abc_41356_new_n2984_), .Y(_abc_41356_new_n2986_));
OR2X2 OR2X2_84 ( .A(_abc_41356_new_n821_), .B(_abc_41356_new_n800_), .Y(_abc_41356_new_n822_));
OR2X2 OR2X2_840 ( .A(_abc_41356_new_n2983_), .B(_abc_41356_new_n2986_), .Y(_0aluoprb_7_0__7_));
OR2X2 OR2X2_841 ( .A(_abc_41356_new_n2990_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n2991_));
OR2X2 OR2X2_842 ( .A(_abc_41356_new_n2995_), .B(_abc_41356_new_n2993_), .Y(_abc_41356_new_n2996_));
OR2X2 OR2X2_843 ( .A(_abc_41356_new_n2996_), .B(_abc_41356_new_n2998_), .Y(_abc_41356_new_n2999_));
OR2X2 OR2X2_844 ( .A(_abc_41356_new_n2999_), .B(_abc_41356_new_n2991_), .Y(_abc_41356_new_n3000_));
OR2X2 OR2X2_845 ( .A(_abc_41356_new_n3002_), .B(opcode_5_), .Y(_abc_41356_new_n3003_));
OR2X2 OR2X2_846 ( .A(_abc_41356_new_n3005_), .B(_abc_41356_new_n3006_), .Y(_abc_41356_new_n3007_));
OR2X2 OR2X2_847 ( .A(_abc_41356_new_n3007_), .B(_abc_41356_new_n3004_), .Y(_abc_41356_new_n3008_));
OR2X2 OR2X2_848 ( .A(_abc_41356_new_n3008_), .B(_abc_41356_new_n3003_), .Y(_abc_41356_new_n3009_));
OR2X2 OR2X2_849 ( .A(_abc_41356_new_n3011_), .B(_abc_41356_new_n2988_), .Y(_abc_41356_new_n3012_));
OR2X2 OR2X2_85 ( .A(_abc_41356_new_n799_), .B(_abc_41356_new_n822_), .Y(_abc_41356_new_n823_));
OR2X2 OR2X2_850 ( .A(_abc_41356_new_n3020_), .B(_abc_41356_new_n3018_), .Y(_abc_41356_new_n3021_));
OR2X2 OR2X2_851 ( .A(_abc_41356_new_n3022_), .B(_abc_41356_new_n3016_), .Y(_abc_41356_new_n3023_));
OR2X2 OR2X2_852 ( .A(_abc_41356_new_n3013_), .B(_abc_41356_new_n3023_), .Y(_0aluopra_7_0__0_));
OR2X2 OR2X2_853 ( .A(_abc_41356_new_n3026_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3027_));
OR2X2 OR2X2_854 ( .A(_abc_41356_new_n3029_), .B(_abc_41356_new_n3028_), .Y(_abc_41356_new_n3030_));
OR2X2 OR2X2_855 ( .A(_abc_41356_new_n3030_), .B(_abc_41356_new_n3031_), .Y(_abc_41356_new_n3032_));
OR2X2 OR2X2_856 ( .A(_abc_41356_new_n3032_), .B(_abc_41356_new_n3027_), .Y(_abc_41356_new_n3033_));
OR2X2 OR2X2_857 ( .A(_abc_41356_new_n3034_), .B(opcode_5_), .Y(_abc_41356_new_n3035_));
OR2X2 OR2X2_858 ( .A(_abc_41356_new_n3037_), .B(_abc_41356_new_n3038_), .Y(_abc_41356_new_n3039_));
OR2X2 OR2X2_859 ( .A(_abc_41356_new_n3039_), .B(_abc_41356_new_n3036_), .Y(_abc_41356_new_n3040_));
OR2X2 OR2X2_86 ( .A(_abc_41356_new_n794_), .B(_abc_41356_new_n823_), .Y(_abc_41356_new_n824_));
OR2X2 OR2X2_860 ( .A(_abc_41356_new_n3040_), .B(_abc_41356_new_n3035_), .Y(_abc_41356_new_n3041_));
OR2X2 OR2X2_861 ( .A(_abc_41356_new_n3043_), .B(_abc_41356_new_n3025_), .Y(_abc_41356_new_n3044_));
OR2X2 OR2X2_862 ( .A(_abc_41356_new_n3047_), .B(_abc_41356_new_n3046_), .Y(_abc_41356_new_n3048_));
OR2X2 OR2X2_863 ( .A(_abc_41356_new_n3045_), .B(_abc_41356_new_n3048_), .Y(_0aluopra_7_0__1_));
OR2X2 OR2X2_864 ( .A(_abc_41356_new_n3051_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3052_));
OR2X2 OR2X2_865 ( .A(_abc_41356_new_n3054_), .B(_abc_41356_new_n3053_), .Y(_abc_41356_new_n3055_));
OR2X2 OR2X2_866 ( .A(_abc_41356_new_n3055_), .B(_abc_41356_new_n3056_), .Y(_abc_41356_new_n3057_));
OR2X2 OR2X2_867 ( .A(_abc_41356_new_n3057_), .B(_abc_41356_new_n3052_), .Y(_abc_41356_new_n3058_));
OR2X2 OR2X2_868 ( .A(_abc_41356_new_n3059_), .B(opcode_5_), .Y(_abc_41356_new_n3060_));
OR2X2 OR2X2_869 ( .A(_abc_41356_new_n3062_), .B(_abc_41356_new_n3063_), .Y(_abc_41356_new_n3064_));
OR2X2 OR2X2_87 ( .A(_abc_41356_new_n824_), .B(_abc_41356_new_n696_), .Y(_abc_41356_new_n825_));
OR2X2 OR2X2_870 ( .A(_abc_41356_new_n3064_), .B(_abc_41356_new_n3061_), .Y(_abc_41356_new_n3065_));
OR2X2 OR2X2_871 ( .A(_abc_41356_new_n3065_), .B(_abc_41356_new_n3060_), .Y(_abc_41356_new_n3066_));
OR2X2 OR2X2_872 ( .A(_abc_41356_new_n3068_), .B(_abc_41356_new_n3050_), .Y(_abc_41356_new_n3069_));
OR2X2 OR2X2_873 ( .A(_abc_41356_new_n3072_), .B(_abc_41356_new_n3071_), .Y(_abc_41356_new_n3073_));
OR2X2 OR2X2_874 ( .A(_abc_41356_new_n3070_), .B(_abc_41356_new_n3073_), .Y(_0aluopra_7_0__2_));
OR2X2 OR2X2_875 ( .A(_abc_41356_new_n3076_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3077_));
OR2X2 OR2X2_876 ( .A(_abc_41356_new_n3079_), .B(_abc_41356_new_n3078_), .Y(_abc_41356_new_n3080_));
OR2X2 OR2X2_877 ( .A(_abc_41356_new_n3080_), .B(_abc_41356_new_n3081_), .Y(_abc_41356_new_n3082_));
OR2X2 OR2X2_878 ( .A(_abc_41356_new_n3082_), .B(_abc_41356_new_n3077_), .Y(_abc_41356_new_n3083_));
OR2X2 OR2X2_879 ( .A(_abc_41356_new_n3084_), .B(opcode_5_), .Y(_abc_41356_new_n3085_));
OR2X2 OR2X2_88 ( .A(_abc_41356_new_n695_), .B(regfil_7__2_), .Y(_abc_41356_new_n826_));
OR2X2 OR2X2_880 ( .A(_abc_41356_new_n3087_), .B(_abc_41356_new_n3088_), .Y(_abc_41356_new_n3089_));
OR2X2 OR2X2_881 ( .A(_abc_41356_new_n3089_), .B(_abc_41356_new_n3086_), .Y(_abc_41356_new_n3090_));
OR2X2 OR2X2_882 ( .A(_abc_41356_new_n3090_), .B(_abc_41356_new_n3085_), .Y(_abc_41356_new_n3091_));
OR2X2 OR2X2_883 ( .A(_abc_41356_new_n3093_), .B(_abc_41356_new_n3075_), .Y(_abc_41356_new_n3094_));
OR2X2 OR2X2_884 ( .A(_abc_41356_new_n3097_), .B(_abc_41356_new_n3096_), .Y(_abc_41356_new_n3098_));
OR2X2 OR2X2_885 ( .A(_abc_41356_new_n3095_), .B(_abc_41356_new_n3098_), .Y(_0aluopra_7_0__3_));
OR2X2 OR2X2_886 ( .A(_abc_41356_new_n3101_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3102_));
OR2X2 OR2X2_887 ( .A(_abc_41356_new_n3104_), .B(_abc_41356_new_n3103_), .Y(_abc_41356_new_n3105_));
OR2X2 OR2X2_888 ( .A(_abc_41356_new_n3105_), .B(_abc_41356_new_n3106_), .Y(_abc_41356_new_n3107_));
OR2X2 OR2X2_889 ( .A(_abc_41356_new_n3107_), .B(_abc_41356_new_n3102_), .Y(_abc_41356_new_n3108_));
OR2X2 OR2X2_89 ( .A(_abc_41356_new_n835_), .B(_abc_41356_new_n836_), .Y(_abc_41356_new_n837_));
OR2X2 OR2X2_890 ( .A(_abc_41356_new_n3109_), .B(opcode_5_), .Y(_abc_41356_new_n3110_));
OR2X2 OR2X2_891 ( .A(_abc_41356_new_n3112_), .B(_abc_41356_new_n3113_), .Y(_abc_41356_new_n3114_));
OR2X2 OR2X2_892 ( .A(_abc_41356_new_n3114_), .B(_abc_41356_new_n3111_), .Y(_abc_41356_new_n3115_));
OR2X2 OR2X2_893 ( .A(_abc_41356_new_n3115_), .B(_abc_41356_new_n3110_), .Y(_abc_41356_new_n3116_));
OR2X2 OR2X2_894 ( .A(_abc_41356_new_n3118_), .B(_abc_41356_new_n3100_), .Y(_abc_41356_new_n3119_));
OR2X2 OR2X2_895 ( .A(_abc_41356_new_n3122_), .B(_abc_41356_new_n3121_), .Y(_abc_41356_new_n3123_));
OR2X2 OR2X2_896 ( .A(_abc_41356_new_n3120_), .B(_abc_41356_new_n3123_), .Y(_0aluopra_7_0__4_));
OR2X2 OR2X2_897 ( .A(_abc_41356_new_n3126_), .B(opcode_5_), .Y(_abc_41356_new_n3127_));
OR2X2 OR2X2_898 ( .A(_abc_41356_new_n3129_), .B(_abc_41356_new_n3130_), .Y(_abc_41356_new_n3131_));
OR2X2 OR2X2_899 ( .A(_abc_41356_new_n3131_), .B(_abc_41356_new_n3128_), .Y(_abc_41356_new_n3132_));
OR2X2 OR2X2_9 ( .A(_abc_41356_new_n594_), .B(_abc_41356_new_n589_), .Y(_abc_41356_new_n595_));
OR2X2 OR2X2_90 ( .A(_abc_41356_new_n838_), .B(_abc_41356_new_n832_), .Y(_abc_41356_new_n839_));
OR2X2 OR2X2_900 ( .A(_abc_41356_new_n3132_), .B(_abc_41356_new_n3127_), .Y(_abc_41356_new_n3133_));
OR2X2 OR2X2_901 ( .A(_abc_41356_new_n3134_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3135_));
OR2X2 OR2X2_902 ( .A(_abc_41356_new_n3137_), .B(_abc_41356_new_n3136_), .Y(_abc_41356_new_n3138_));
OR2X2 OR2X2_903 ( .A(_abc_41356_new_n3138_), .B(_abc_41356_new_n3139_), .Y(_abc_41356_new_n3140_));
OR2X2 OR2X2_904 ( .A(_abc_41356_new_n3140_), .B(_abc_41356_new_n3135_), .Y(_abc_41356_new_n3141_));
OR2X2 OR2X2_905 ( .A(_abc_41356_new_n3143_), .B(_abc_41356_new_n3125_), .Y(_abc_41356_new_n3144_));
OR2X2 OR2X2_906 ( .A(_abc_41356_new_n3147_), .B(_abc_41356_new_n3146_), .Y(_abc_41356_new_n3148_));
OR2X2 OR2X2_907 ( .A(_abc_41356_new_n3145_), .B(_abc_41356_new_n3148_), .Y(_0aluopra_7_0__5_));
OR2X2 OR2X2_908 ( .A(_abc_41356_new_n3151_), .B(opcode_5_), .Y(_abc_41356_new_n3152_));
OR2X2 OR2X2_909 ( .A(_abc_41356_new_n3154_), .B(_abc_41356_new_n3155_), .Y(_abc_41356_new_n3156_));
OR2X2 OR2X2_91 ( .A(_abc_41356_new_n840_), .B(_abc_41356_new_n512_), .Y(_abc_41356_new_n841_));
OR2X2 OR2X2_910 ( .A(_abc_41356_new_n3156_), .B(_abc_41356_new_n3153_), .Y(_abc_41356_new_n3157_));
OR2X2 OR2X2_911 ( .A(_abc_41356_new_n3157_), .B(_abc_41356_new_n3152_), .Y(_abc_41356_new_n3158_));
OR2X2 OR2X2_912 ( .A(_abc_41356_new_n3159_), .B(_abc_41356_new_n525_), .Y(_abc_41356_new_n3160_));
OR2X2 OR2X2_913 ( .A(_abc_41356_new_n3162_), .B(_abc_41356_new_n3161_), .Y(_abc_41356_new_n3163_));
OR2X2 OR2X2_914 ( .A(_abc_41356_new_n3163_), .B(_abc_41356_new_n3164_), .Y(_abc_41356_new_n3165_));
OR2X2 OR2X2_915 ( .A(_abc_41356_new_n3165_), .B(_abc_41356_new_n3160_), .Y(_abc_41356_new_n3166_));
OR2X2 OR2X2_916 ( .A(_abc_41356_new_n3168_), .B(_abc_41356_new_n3150_), .Y(_abc_41356_new_n3169_));
OR2X2 OR2X2_917 ( .A(_abc_41356_new_n3172_), .B(_abc_41356_new_n3171_), .Y(_abc_41356_new_n3173_));
OR2X2 OR2X2_918 ( .A(_abc_41356_new_n3170_), .B(_abc_41356_new_n3173_), .Y(_0aluopra_7_0__6_));
OR2X2 OR2X2_919 ( .A(_abc_41356_new_n3176_), .B(_abc_41356_new_n3177_), .Y(_abc_41356_new_n3178_));
OR2X2 OR2X2_92 ( .A(_abc_41356_new_n839_), .B(_abc_41356_new_n841_), .Y(_abc_41356_new_n842_));
OR2X2 OR2X2_920 ( .A(_abc_41356_new_n3180_), .B(_abc_41356_new_n3179_), .Y(_abc_41356_new_n3181_));
OR2X2 OR2X2_921 ( .A(_abc_41356_new_n3178_), .B(_abc_41356_new_n3181_), .Y(_abc_41356_new_n3182_));
OR2X2 OR2X2_922 ( .A(_abc_41356_new_n3184_), .B(_abc_41356_new_n3185_), .Y(_abc_41356_new_n3186_));
OR2X2 OR2X2_923 ( .A(_abc_41356_new_n3187_), .B(_abc_41356_new_n3188_), .Y(_abc_41356_new_n3189_));
OR2X2 OR2X2_924 ( .A(_abc_41356_new_n3189_), .B(_abc_41356_new_n3186_), .Y(_abc_41356_new_n3190_));
OR2X2 OR2X2_925 ( .A(_abc_41356_new_n3183_), .B(_abc_41356_new_n3191_), .Y(_abc_41356_new_n3192_));
OR2X2 OR2X2_926 ( .A(_abc_41356_new_n3193_), .B(_abc_41356_new_n3175_), .Y(_abc_41356_new_n3194_));
OR2X2 OR2X2_927 ( .A(_abc_41356_new_n3197_), .B(_abc_41356_new_n3196_), .Y(_abc_41356_new_n3198_));
OR2X2 OR2X2_928 ( .A(_abc_41356_new_n3195_), .B(_abc_41356_new_n3198_), .Y(_0aluopra_7_0__7_));
OR2X2 OR2X2_929 ( .A(_abc_41356_new_n3201_), .B(_abc_41356_new_n3202_), .Y(_abc_41356_new_n3203_));
OR2X2 OR2X2_93 ( .A(_abc_41356_new_n846_), .B(_abc_41356_new_n845_), .Y(_abc_41356_new_n847_));
OR2X2 OR2X2_930 ( .A(_abc_41356_new_n3203_), .B(_abc_41356_new_n3200_), .Y(_abc_41356_new_n3204_));
OR2X2 OR2X2_931 ( .A(_abc_41356_new_n3205_), .B(intcyc), .Y(_abc_41356_new_n3206_));
OR2X2 OR2X2_932 ( .A(_abc_41356_new_n3211_), .B(_abc_41356_new_n3210_), .Y(_abc_41356_new_n3212_));
OR2X2 OR2X2_933 ( .A(_abc_41356_new_n3214_), .B(reset), .Y(_abc_41356_new_n3215_));
OR2X2 OR2X2_934 ( .A(_abc_41356_new_n3220_), .B(_abc_41356_new_n3218_), .Y(_abc_41356_new_n3221_));
OR2X2 OR2X2_935 ( .A(_abc_41356_new_n3217_), .B(_abc_41356_new_n3222_), .Y(_abc_41356_new_n3223_));
OR2X2 OR2X2_936 ( .A(_abc_41356_new_n3216_), .B(_abc_41356_new_n3224_), .Y(_0parity_0_0_));
OR2X2 OR2X2_937 ( .A(_abc_41356_new_n3229_), .B(_abc_41356_new_n3228_), .Y(_abc_41356_new_n3230_));
OR2X2 OR2X2_938 ( .A(_abc_41356_new_n3227_), .B(_abc_41356_new_n3231_), .Y(_abc_41356_new_n3232_));
OR2X2 OR2X2_939 ( .A(_abc_41356_new_n3226_), .B(_abc_41356_new_n3233_), .Y(_0zero_0_0_));
OR2X2 OR2X2_94 ( .A(_abc_41356_new_n847_), .B(_abc_41356_new_n844_), .Y(_abc_41356_new_n848_));
OR2X2 OR2X2_940 ( .A(_abc_41356_new_n510_), .B(sign), .Y(_abc_41356_new_n3239_));
OR2X2 OR2X2_941 ( .A(_abc_41356_new_n3243_), .B(_abc_41356_new_n3242_), .Y(_abc_41356_new_n3244_));
OR2X2 OR2X2_942 ( .A(_abc_41356_new_n3244_), .B(_abc_41356_new_n3241_), .Y(_abc_41356_new_n3245_));
OR2X2 OR2X2_943 ( .A(_abc_41356_new_n3235_), .B(_abc_41356_new_n3246_), .Y(_0sign_0_0_));
OR2X2 OR2X2_944 ( .A(_abc_41356_new_n3249_), .B(_abc_41356_new_n3248_), .Y(_abc_41356_new_n3250_));
OR2X2 OR2X2_945 ( .A(_abc_41356_new_n549_), .B(auxcar), .Y(_abc_41356_new_n3251_));
OR2X2 OR2X2_946 ( .A(_abc_41356_new_n3254_), .B(_abc_41356_new_n3255_), .Y(_abc_41356_new_n3256_));
OR2X2 OR2X2_947 ( .A(_abc_41356_new_n3258_), .B(_abc_41356_new_n3257_), .Y(_abc_41356_new_n3259_));
OR2X2 OR2X2_948 ( .A(_abc_41356_new_n3253_), .B(_abc_41356_new_n3259_), .Y(_abc_41356_new_n3260_));
OR2X2 OR2X2_949 ( .A(_abc_41356_new_n3261_), .B(_abc_41356_new_n3263_), .Y(_0auxcar_0_0_));
OR2X2 OR2X2_95 ( .A(_abc_41356_new_n843_), .B(_abc_41356_new_n848_), .Y(_abc_41356_new_n849_));
OR2X2 OR2X2_950 ( .A(_abc_41356_new_n3266_), .B(reset), .Y(_abc_41356_new_n3267_));
OR2X2 OR2X2_951 ( .A(_abc_41356_new_n3272_), .B(_abc_41356_new_n1981_), .Y(_abc_41356_new_n3273_));
OR2X2 OR2X2_952 ( .A(_abc_41356_new_n1994_), .B(_abc_41356_new_n1998_), .Y(_abc_41356_new_n3275_));
OR2X2 OR2X2_953 ( .A(_abc_41356_new_n3282_), .B(_abc_41356_new_n3281_), .Y(_abc_41356_new_n3283_));
OR2X2 OR2X2_954 ( .A(_abc_41356_new_n3285_), .B(_abc_41356_new_n3284_), .Y(_abc_41356_new_n3286_));
OR2X2 OR2X2_955 ( .A(_abc_41356_new_n3283_), .B(_abc_41356_new_n3286_), .Y(_abc_41356_new_n3287_));
OR2X2 OR2X2_956 ( .A(_abc_41356_new_n3278_), .B(_abc_41356_new_n3287_), .Y(_abc_41356_new_n3288_));
OR2X2 OR2X2_957 ( .A(_abc_41356_new_n3274_), .B(_abc_41356_new_n3288_), .Y(_abc_41356_new_n3289_));
OR2X2 OR2X2_958 ( .A(_abc_41356_new_n1966_), .B(_abc_41356_new_n1969_), .Y(_abc_41356_new_n3290_));
OR2X2 OR2X2_959 ( .A(_abc_41356_new_n3289_), .B(_abc_41356_new_n3293_), .Y(_abc_41356_new_n3294_));
OR2X2 OR2X2_96 ( .A(_abc_41356_new_n828_), .B(_abc_41356_new_n849_), .Y(_abc_36060_memoryregfil_wrmux_7__4__0__y_16247_2_));
OR2X2 OR2X2_960 ( .A(_abc_41356_new_n3299_), .B(_abc_41356_new_n2021_), .Y(_abc_41356_new_n3300_));
OR2X2 OR2X2_961 ( .A(_abc_41356_new_n3298_), .B(_abc_41356_new_n3300_), .Y(_abc_41356_new_n3301_));
OR2X2 OR2X2_962 ( .A(_abc_41356_new_n3294_), .B(_abc_41356_new_n3301_), .Y(_abc_41356_new_n3302_));
OR2X2 OR2X2_963 ( .A(_abc_41356_new_n516_), .B(carry), .Y(_abc_41356_new_n3303_));
OR2X2 OR2X2_964 ( .A(_abc_41356_new_n3306_), .B(_abc_41356_new_n3307_), .Y(_abc_41356_new_n3308_));
OR2X2 OR2X2_965 ( .A(_abc_41356_new_n3309_), .B(_abc_41356_new_n3310_), .Y(_abc_41356_new_n3311_));
OR2X2 OR2X2_966 ( .A(_abc_41356_new_n3308_), .B(_abc_41356_new_n3312_), .Y(_abc_41356_new_n3313_));
OR2X2 OR2X2_967 ( .A(_abc_41356_new_n3305_), .B(_abc_41356_new_n3313_), .Y(_abc_41356_new_n3314_));
OR2X2 OR2X2_968 ( .A(_abc_41356_new_n3315_), .B(_abc_41356_new_n3271_), .Y(_0carry_0_0_));
OR2X2 OR2X2_969 ( .A(_abc_41356_new_n3319_), .B(opcode_0_), .Y(_abc_41356_new_n3320_));
OR2X2 OR2X2_97 ( .A(_abc_41356_new_n790_), .B(regfil_0__3_), .Y(_abc_41356_new_n851_));
OR2X2 OR2X2_970 ( .A(_abc_41356_new_n3321_), .B(\data[0] ), .Y(_abc_41356_new_n3322_));
OR2X2 OR2X2_971 ( .A(_abc_41356_new_n3325_), .B(_abc_41356_new_n3324_), .Y(_0opcode_7_0__1_));
OR2X2 OR2X2_972 ( .A(_abc_41356_new_n3319_), .B(opcode_2_), .Y(_abc_41356_new_n3327_));
OR2X2 OR2X2_973 ( .A(_abc_41356_new_n3321_), .B(\data[2] ), .Y(_abc_41356_new_n3328_));
OR2X2 OR2X2_974 ( .A(_abc_41356_new_n3331_), .B(_abc_41356_new_n3330_), .Y(_0opcode_7_0__3_));
OR2X2 OR2X2_975 ( .A(_abc_41356_new_n3319_), .B(opcode_4_), .Y(_abc_41356_new_n3333_));
OR2X2 OR2X2_976 ( .A(_abc_41356_new_n3321_), .B(\data[4] ), .Y(_abc_41356_new_n3334_));
OR2X2 OR2X2_977 ( .A(_abc_41356_new_n3319_), .B(opcode_5_), .Y(_abc_41356_new_n3336_));
OR2X2 OR2X2_978 ( .A(_abc_41356_new_n3321_), .B(\data[5] ), .Y(_abc_41356_new_n3337_));
OR2X2 OR2X2_979 ( .A(_abc_41356_new_n3340_), .B(_abc_41356_new_n3339_), .Y(_0opcode_7_0__6_));
OR2X2 OR2X2_98 ( .A(_abc_41356_new_n852_), .B(_abc_41356_new_n853_), .Y(_abc_41356_new_n854_));
OR2X2 OR2X2_980 ( .A(_abc_41356_new_n3343_), .B(_abc_41356_new_n3342_), .Y(_0opcode_7_0__7_));
OR2X2 OR2X2_981 ( .A(_abc_41356_new_n3346_), .B(_abc_41356_new_n676_), .Y(_abc_41356_new_n3347_));
OR2X2 OR2X2_982 ( .A(_abc_41356_new_n3350_), .B(_abc_41356_new_n3348_), .Y(_abc_41356_new_n3351_));
OR2X2 OR2X2_983 ( .A(_abc_41356_new_n3369_), .B(_abc_41356_new_n580_), .Y(_abc_41356_new_n3370_));
OR2X2 OR2X2_984 ( .A(_abc_41356_new_n2027_), .B(_abc_41356_new_n3373_), .Y(_abc_41356_new_n3374_));
OR2X2 OR2X2_985 ( .A(_abc_41356_new_n3374_), .B(_abc_41356_new_n3371_), .Y(_abc_41356_new_n3375_));
OR2X2 OR2X2_986 ( .A(_abc_41356_new_n3375_), .B(_abc_41356_new_n3370_), .Y(_abc_41356_new_n3376_));
OR2X2 OR2X2_987 ( .A(_abc_41356_new_n3376_), .B(_abc_41356_new_n3377_), .Y(_abc_41356_new_n3378_));
OR2X2 OR2X2_988 ( .A(_abc_41356_new_n3386_), .B(_abc_41356_new_n3385_), .Y(_abc_41356_new_n3387_));
OR2X2 OR2X2_989 ( .A(_abc_41356_new_n3384_), .B(_abc_41356_new_n3387_), .Y(_abc_41356_new_n3388_));
OR2X2 OR2X2_99 ( .A(_abc_41356_new_n796_), .B(regfil_0__3_), .Y(_abc_41356_new_n856_));
OR2X2 OR2X2_990 ( .A(_abc_41356_new_n3383_), .B(_abc_41356_new_n3388_), .Y(_abc_41356_new_n3389_));
OR2X2 OR2X2_991 ( .A(_abc_41356_new_n3369_), .B(_abc_41356_new_n2027_), .Y(_abc_41356_new_n3392_));
OR2X2 OR2X2_992 ( .A(_abc_41356_new_n677_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n3396_));
OR2X2 OR2X2_993 ( .A(_abc_41356_new_n3396_), .B(_abc_41356_new_n3395_), .Y(_abc_41356_new_n3397_));
OR2X2 OR2X2_994 ( .A(_abc_41356_new_n3397_), .B(_abc_41356_new_n3394_), .Y(_abc_41356_new_n3398_));
OR2X2 OR2X2_995 ( .A(_abc_41356_new_n3398_), .B(_abc_41356_new_n3393_), .Y(_abc_41356_new_n3399_));
OR2X2 OR2X2_996 ( .A(_abc_41356_new_n3399_), .B(_abc_41356_new_n3392_), .Y(_abc_41356_new_n3400_));
OR2X2 OR2X2_997 ( .A(_abc_41356_new_n3401_), .B(_abc_41356_new_n2874_), .Y(_abc_41356_new_n3402_));
OR2X2 OR2X2_998 ( .A(_abc_41356_new_n3401_), .B(_abc_41356_new_n683_), .Y(_abc_41356_new_n3404_));
OR2X2 OR2X2_999 ( .A(_abc_41356_new_n3405_), .B(_abc_41356_new_n3391_), .Y(_abc_41356_new_n3406_));


endmodule