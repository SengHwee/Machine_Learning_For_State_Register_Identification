module b06_reset(clock, RESET_G, nRESET_G, EQL, CONT_EQL, CC_MUX_REG_2_, CC_MUX_REG_1_, USCITE_REG_2_, USCITE_REG_1_, ENABLE_COUNT_REG, ACKOUT_REG);
  output ACKOUT_REG;
  output CC_MUX_REG_1_;
  output CC_MUX_REG_2_;
  input CONT_EQL;
  output ENABLE_COUNT_REG;
  input EQL;
  input RESET_G;
  wire STATE_REG_0_;
  wire STATE_REG_1_;
  wire STATE_REG_2_;
  output USCITE_REG_1_;
  output USCITE_REG_2_;
  wire _abc_317_n15;
  wire _abc_317_n16;
  wire _abc_317_n17;
  wire _abc_317_n18;
  wire _abc_317_n19;
  wire _abc_317_n20;
  wire _abc_317_n21;
  wire _abc_317_n22;
  wire _abc_317_n23_1;
  wire _abc_317_n24;
  wire _abc_317_n25;
  wire _abc_317_n27;
  wire _abc_317_n28;
  wire _abc_317_n29_1;
  wire _abc_317_n30;
  wire _abc_317_n31;
  wire _abc_317_n32;
  wire _abc_317_n33;
  wire _abc_317_n34;
  wire _abc_317_n35_1;
  wire _abc_317_n36;
  wire _abc_317_n38;
  wire _abc_317_n39_1;
  wire _abc_317_n40;
  wire _abc_317_n41;
  wire _abc_317_n42_1;
  wire _abc_317_n43;
  wire _abc_317_n44_1;
  wire _abc_317_n46;
  wire _abc_317_n47;
  wire _abc_317_n48_1;
  wire _abc_317_n49;
  wire _abc_317_n50;
  wire _abc_317_n51;
  wire _abc_317_n52;
  wire _abc_317_n53;
  wire _abc_317_n55;
  wire _abc_317_n56;
  wire _abc_317_n57;
  wire _abc_317_n58;
  wire _abc_317_n59;
  wire _abc_317_n61;
  wire _abc_317_n62;
  wire _abc_317_n64;
  wire _abc_317_n66;
  wire _abc_317_n67;
  wire _abc_317_n68;
  wire _abc_317_n69;
  wire _abc_317_n70;
  input clock;
  wire n22;
  wire n26;
  wire n31;
  wire n36;
  wire n41;
  wire n45;
  wire n49;
  wire n53;
  input nRESET_G;
  AND2X2 AND2X2_1 ( .A(_abc_317_n19), .B(_abc_317_n16), .Y(_abc_317_n20) );
  AND2X2 AND2X2_10 ( .A(_abc_317_n41), .B(_abc_317_n43), .Y(_abc_317_n44_1) );
  AND2X2 AND2X2_11 ( .A(STATE_REG_1_), .B(EQL), .Y(_abc_317_n46) );
  AND2X2 AND2X2_12 ( .A(_abc_317_n46), .B(_abc_317_n27), .Y(_abc_317_n47) );
  AND2X2 AND2X2_13 ( .A(_abc_317_n17), .B(nRESET_G), .Y(_abc_317_n49) );
  AND2X2 AND2X2_14 ( .A(STATE_REG_2_), .B(STATE_REG_0_), .Y(_abc_317_n50) );
  AND2X2 AND2X2_15 ( .A(_abc_317_n49), .B(_abc_317_n51), .Y(_abc_317_n52) );
  AND2X2 AND2X2_16 ( .A(_abc_317_n52), .B(_abc_317_n48_1), .Y(_abc_317_n53) );
  AND2X2 AND2X2_17 ( .A(_abc_317_n55), .B(nRESET_G), .Y(_abc_317_n56) );
  AND2X2 AND2X2_18 ( .A(_abc_317_n38), .B(_abc_317_n57), .Y(_abc_317_n58) );
  AND2X2 AND2X2_19 ( .A(_abc_317_n58), .B(_abc_317_n56), .Y(_abc_317_n59) );
  AND2X2 AND2X2_2 ( .A(_abc_317_n23_1), .B(_abc_317_n22), .Y(_abc_317_n24) );
  AND2X2 AND2X2_20 ( .A(_abc_317_n19), .B(_abc_317_n61), .Y(_abc_317_n62) );
  AND2X2 AND2X2_21 ( .A(_abc_317_n46), .B(STATE_REG_2_), .Y(_abc_317_n64) );
  AND2X2 AND2X2_22 ( .A(_abc_317_n50), .B(STATE_REG_1_), .Y(_abc_317_n67) );
  AND2X2 AND2X2_23 ( .A(_abc_317_n68), .B(nRESET_G), .Y(_abc_317_n69) );
  AND2X2 AND2X2_24 ( .A(_abc_317_n69), .B(_abc_317_n66), .Y(_abc_317_n70) );
  AND2X2 AND2X2_3 ( .A(_abc_317_n27), .B(STATE_REG_2_), .Y(_abc_317_n28) );
  AND2X2 AND2X2_4 ( .A(_abc_317_n15), .B(_abc_317_n22), .Y(_abc_317_n29_1) );
  AND2X2 AND2X2_5 ( .A(_abc_317_n29_1), .B(_abc_317_n28), .Y(_abc_317_n30) );
  AND2X2 AND2X2_6 ( .A(_abc_317_n33), .B(STATE_REG_0_), .Y(_abc_317_n34) );
  AND2X2 AND2X2_7 ( .A(_abc_317_n32), .B(_abc_317_n35_1), .Y(_abc_317_n36) );
  AND2X2 AND2X2_8 ( .A(_abc_317_n34), .B(_abc_317_n15), .Y(_abc_317_n40) );
  AND2X2 AND2X2_9 ( .A(EQL), .B(nRESET_G), .Y(_abc_317_n42_1) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n41), .Q(CC_MUX_REG_2_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n45), .Q(CC_MUX_REG_1_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n49), .Q(USCITE_REG_2_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n53), .Q(USCITE_REG_1_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n22), .Q(ACKOUT_REG) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n26), .Q(STATE_REG_2_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n31), .Q(STATE_REG_1_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n36), .Q(STATE_REG_0_) );
  INVX1 INVX1_1 ( .A(STATE_REG_1_), .Y(_abc_317_n15) );
  INVX1 INVX1_10 ( .A(_abc_317_n53), .Y(n45) );
  INVX1 INVX1_11 ( .A(_abc_317_n40), .Y(_abc_317_n55) );
  INVX1 INVX1_12 ( .A(_abc_317_n47), .Y(_abc_317_n57) );
  INVX1 INVX1_13 ( .A(_abc_317_n59), .Y(n41) );
  INVX1 INVX1_14 ( .A(_abc_317_n70), .Y(n22) );
  INVX1 INVX1_2 ( .A(_abc_317_n17), .Y(_abc_317_n18) );
  INVX1 INVX1_3 ( .A(nRESET_G), .Y(_abc_317_n21) );
  INVX1 INVX1_4 ( .A(EQL), .Y(_abc_317_n22) );
  INVX1 INVX1_5 ( .A(STATE_REG_0_), .Y(_abc_317_n27) );
  INVX1 INVX1_6 ( .A(STATE_REG_2_), .Y(_abc_317_n33) );
  INVX1 INVX1_7 ( .A(_abc_317_n38), .Y(_abc_317_n39_1) );
  INVX1 INVX1_8 ( .A(_abc_317_n42_1), .Y(_abc_317_n43) );
  INVX1 INVX1_9 ( .A(_abc_317_n50), .Y(_abc_317_n51) );
  OR2X2 OR2X2_1 ( .A(_abc_317_n15), .B(STATE_REG_0_), .Y(_abc_317_n16) );
  OR2X2 OR2X2_10 ( .A(_abc_317_n36), .B(_abc_317_n31), .Y(n31) );
  OR2X2 OR2X2_11 ( .A(_abc_317_n24), .B(_abc_317_n33), .Y(_abc_317_n38) );
  OR2X2 OR2X2_12 ( .A(_abc_317_n40), .B(_abc_317_n21), .Y(_abc_317_n41) );
  OR2X2 OR2X2_13 ( .A(_abc_317_n44_1), .B(_abc_317_n39_1), .Y(n26) );
  OR2X2 OR2X2_14 ( .A(_abc_317_n47), .B(_abc_317_n29_1), .Y(_abc_317_n48_1) );
  OR2X2 OR2X2_15 ( .A(_abc_317_n17), .B(_abc_317_n15), .Y(_abc_317_n61) );
  OR2X2 OR2X2_16 ( .A(_abc_317_n62), .B(_abc_317_n43), .Y(n53) );
  OR2X2 OR2X2_17 ( .A(_abc_317_n31), .B(_abc_317_n64), .Y(n49) );
  OR2X2 OR2X2_18 ( .A(_abc_317_n61), .B(EQL), .Y(_abc_317_n66) );
  OR2X2 OR2X2_19 ( .A(_abc_317_n67), .B(CONT_EQL), .Y(_abc_317_n68) );
  OR2X2 OR2X2_2 ( .A(STATE_REG_2_), .B(STATE_REG_0_), .Y(_abc_317_n17) );
  OR2X2 OR2X2_3 ( .A(_abc_317_n18), .B(STATE_REG_1_), .Y(_abc_317_n19) );
  OR2X2 OR2X2_4 ( .A(STATE_REG_0_), .B(STATE_REG_1_), .Y(_abc_317_n23_1) );
  OR2X2 OR2X2_5 ( .A(_abc_317_n24), .B(_abc_317_n21), .Y(_abc_317_n25) );
  OR2X2 OR2X2_6 ( .A(_abc_317_n20), .B(_abc_317_n25), .Y(n36) );
  OR2X2 OR2X2_7 ( .A(_abc_317_n30), .B(_abc_317_n21), .Y(_abc_317_n31) );
  OR2X2 OR2X2_8 ( .A(_abc_317_n18), .B(EQL), .Y(_abc_317_n32) );
  OR2X2 OR2X2_9 ( .A(_abc_317_n34), .B(STATE_REG_1_), .Y(_abc_317_n35_1) );
endmodule